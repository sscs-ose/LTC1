** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/MUX_TB.sch
**.subckt MUX_TB
V1 VSS GND 0
.save i(v1)
V2 VDD VSS 3.3
.save i(v2)
V3 SEL VSS pulse(0 3.3 0 100p 100p 100n 200n)
.save i(v3)
C1 OUT VSS 50f m=1
V4 A VSS 0
.save i(v4)
V5 B VSS 3.3
.save i(v5)
x1 VDD VSS A B SEL OUT pex_Mux2x1
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.include pex_Mux2x1.spice
.control
save all
*dc v3 0 3.3 0.1

tran 10p 1u
plot v(A) v(B)+3.5 v(SEL)+7 v(OUT)+10.5
*write test_nfet_03v3.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
