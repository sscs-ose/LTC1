magic
tech gf180mcuD
magscale 1 10
timestamp 1714565245
<< nwell >>
rect 8578 11491 8995 11493
rect 8561 11488 8995 11491
rect 35448 -7135 35605 -7054
rect 34288 -8979 34546 -8905
rect 37498 -8979 37754 -8906
<< pwell >>
rect -1655 14936 1868 15545
rect 2266 14920 4018 15522
rect -1972 11532 2228 12319
rect -1972 10320 2228 11104
rect 25669 10957 25993 11253
rect 25669 9223 25993 9500
<< nsubdiff >>
rect 35448 -7135 35605 -7054
rect 34288 -8979 34546 -8905
rect 37498 -8979 37754 -8906
<< metal1 >>
rect -734 55462 -180 55520
rect 4523 55463 5059 55511
rect 2762 54729 2988 54776
rect 8386 54369 8903 54424
rect -2698 52726 -2423 52744
rect -2698 52674 -2669 52726
rect -2617 52724 -2423 52726
rect -2617 52674 -2505 52724
rect -2698 52672 -2505 52674
rect -2453 52672 -2423 52724
rect -2698 52639 -2423 52672
rect -3477 52612 -2423 52639
rect -3477 52599 -2503 52612
rect -3477 52547 -2669 52599
rect -2617 52560 -2503 52599
rect -2451 52560 -2423 52612
rect -2617 52547 -2423 52560
rect -3477 52491 -2423 52547
rect -2698 52472 -2423 52491
rect -2698 52461 -2498 52472
rect -2698 52409 -2669 52461
rect -2617 52420 -2498 52461
rect -2446 52420 -2423 52472
rect -2617 52409 -2423 52420
rect -2698 52394 -2423 52409
rect 9089 48634 9166 48762
rect -1113 48238 -1066 48601
rect -2388 44200 -2113 44218
rect -2388 44148 -2359 44200
rect -2307 44198 -2113 44200
rect -2307 44148 -2195 44198
rect -2388 44146 -2195 44148
rect -2143 44146 -2113 44198
rect -2388 44086 -2113 44146
rect -2388 44073 -2193 44086
rect -3246 44021 -2359 44073
rect -2307 44034 -2193 44073
rect -2141 44034 -2113 44086
rect -2307 44021 -2113 44034
rect -3246 43946 -2113 44021
rect -3246 43935 -2188 43946
rect -3246 43925 -2359 43935
rect -2388 43883 -2359 43925
rect -2307 43894 -2188 43935
rect -2136 43894 -2113 43946
rect -2307 43883 -2113 43894
rect -2388 43868 -2113 43883
rect -2381 43659 -2106 43677
rect -2381 43607 -2352 43659
rect -2300 43657 -2106 43659
rect -2300 43607 -2188 43657
rect -2381 43605 -2188 43607
rect -2136 43605 -2106 43657
rect -2381 43547 -2106 43605
rect -3246 43545 -2106 43547
rect -3246 43532 -2186 43545
rect -3246 43480 -2352 43532
rect -2300 43493 -2186 43532
rect -2134 43493 -2106 43545
rect -2300 43480 -2106 43493
rect -3246 43405 -2106 43480
rect -3246 43399 -2181 43405
rect -2381 43394 -2181 43399
rect -2381 43342 -2352 43394
rect -2300 43353 -2181 43394
rect -2129 43353 -2106 43405
rect -2300 43342 -2106 43353
rect -2381 43327 -2106 43342
rect 7285 41464 7336 42465
rect 7526 40566 7997 40618
rect 61 39776 236 39866
rect 4351 39720 4955 39766
rect -2489 36766 -2214 36784
rect -2489 36714 -2460 36766
rect -2408 36764 -2214 36766
rect -2408 36714 -2296 36764
rect -2489 36712 -2296 36714
rect -2244 36712 -2214 36764
rect -2489 36680 -2214 36712
rect -3157 36652 -2214 36680
rect -3157 36639 -2294 36652
rect -3157 36587 -2460 36639
rect -2408 36600 -2294 36639
rect -2242 36600 -2214 36652
rect -2408 36587 -2214 36600
rect -3157 36532 -2214 36587
rect -2489 36512 -2214 36532
rect -2489 36501 -2289 36512
rect -2489 36449 -2460 36501
rect -2408 36460 -2289 36501
rect -2237 36460 -2214 36512
rect -2408 36449 -2214 36460
rect -2489 36434 -2214 36449
rect 2010 28025 2740 28118
rect 2010 28017 2609 28025
rect 2010 27965 2043 28017
rect 2095 28014 2419 28017
rect 2095 27965 2222 28014
rect 2010 27962 2222 27965
rect 2274 27965 2419 28014
rect 2471 27973 2609 28017
rect 2661 27973 2740 28025
rect 2471 27965 2740 27973
rect 2274 27962 2740 27965
rect 2010 27890 2740 27962
rect 2010 27838 2046 27890
rect 2098 27882 2609 27890
rect 2098 27879 2411 27882
rect 2098 27838 2222 27879
rect 2010 27827 2222 27838
rect 2274 27830 2411 27879
rect 2463 27838 2609 27882
rect 2661 27838 2740 27890
rect 2463 27830 2740 27838
rect 2274 27827 2740 27830
rect 2010 27720 2740 27827
rect 5020 26011 5999 26363
rect -3588 25040 -3261 25051
rect -3588 24988 -3571 25040
rect -3519 24988 -3451 25040
rect -3399 24988 -3331 25040
rect -3279 24988 -3261 25040
rect -3588 24965 -3261 24988
rect -3896 24920 -3261 24965
rect -3896 24868 -3571 24920
rect -3519 24868 -3451 24920
rect -3399 24868 -3331 24920
rect -3279 24868 -3261 24920
rect -3896 24824 -3261 24868
rect -3588 24800 -3261 24824
rect -3588 24748 -3571 24800
rect -3519 24748 -3451 24800
rect -3399 24748 -3331 24800
rect -3279 24748 -3261 24800
rect -3588 24732 -3261 24748
rect -1788 23765 -968 23954
rect -15701 22681 -2908 23203
rect 5647 23168 5999 26011
rect 2715 22816 11131 23168
rect -16303 20819 -5921 21327
rect -6429 19580 -5921 20819
rect -3430 21220 -2908 22681
rect -3430 20698 20375 21220
rect -6429 19524 16649 19580
rect -6429 19472 14140 19524
rect 14192 19472 14311 19524
rect 14363 19472 14482 19524
rect 14534 19472 14653 19524
rect 14705 19472 14824 19524
rect 14876 19472 14995 19524
rect 15047 19472 15166 19524
rect 15218 19472 15337 19524
rect 15389 19472 15508 19524
rect 15560 19472 15679 19524
rect 15731 19472 15850 19524
rect 15902 19472 16021 19524
rect 16073 19472 16192 19524
rect 16244 19472 16363 19524
rect 16415 19472 16534 19524
rect 16586 19472 16649 19524
rect -6429 19359 16649 19472
rect -6429 19307 14140 19359
rect 14192 19307 14311 19359
rect 14363 19307 14482 19359
rect 14534 19307 14653 19359
rect 14705 19307 14824 19359
rect 14876 19307 14995 19359
rect 15047 19307 15166 19359
rect 15218 19307 15337 19359
rect 15389 19307 15508 19359
rect 15560 19307 15679 19359
rect 15731 19307 15850 19359
rect 15902 19307 16021 19359
rect 16073 19307 16192 19359
rect 16244 19307 16363 19359
rect 16415 19307 16534 19359
rect 16586 19307 16649 19359
rect -6429 19194 16649 19307
rect -15247 18808 -10439 19168
rect -6429 19142 14140 19194
rect 14192 19142 14311 19194
rect 14363 19142 14482 19194
rect 14534 19142 14653 19194
rect 14705 19142 14824 19194
rect 14876 19142 14995 19194
rect 15047 19142 15166 19194
rect 15218 19142 15337 19194
rect 15389 19142 15508 19194
rect 15560 19142 15679 19194
rect 15731 19142 15850 19194
rect 15902 19142 16021 19194
rect 16073 19142 16192 19194
rect 16244 19142 16363 19194
rect 16415 19142 16534 19194
rect 16586 19142 16649 19194
rect -6429 19073 16649 19142
rect -6429 19072 13608 19073
rect 14077 19031 16649 19073
rect 19853 19560 20375 20698
rect 19853 19038 24914 19560
rect -15247 18756 -13882 18808
rect -13830 18756 -13758 18808
rect -13706 18756 -13634 18808
rect -13582 18756 -13510 18808
rect -13458 18756 -10439 18808
rect -15247 18684 -10439 18756
rect -15247 18632 -13882 18684
rect -13830 18632 -13758 18684
rect -13706 18632 -13634 18684
rect -13582 18632 -13510 18684
rect -13458 18632 -10439 18684
rect -15247 18560 -10439 18632
rect -15247 18508 -13882 18560
rect -13830 18508 -13758 18560
rect -13706 18508 -13634 18560
rect -13582 18508 -13510 18560
rect -13458 18508 -10439 18560
rect -15247 18441 -10439 18508
rect -17257 18436 -10439 18441
rect -17257 18384 -13882 18436
rect -13830 18384 -13758 18436
rect -13706 18384 -13634 18436
rect -13582 18384 -13510 18436
rect -13458 18384 -10439 18436
rect -17257 17722 -10439 18384
rect -17257 17670 -13966 17722
rect -13914 17670 -13842 17722
rect -13790 17670 -13718 17722
rect -13666 17670 -13594 17722
rect -13542 17714 -10439 17722
rect -13542 17670 -12463 17714
rect -17257 17662 -12463 17670
rect -12411 17662 -12339 17714
rect -12287 17662 -12215 17714
rect -12163 17662 -12091 17714
rect -12039 17662 -10439 17714
rect -17257 17598 -10439 17662
rect -17257 17546 -13966 17598
rect -13914 17546 -13842 17598
rect -13790 17546 -13718 17598
rect -13666 17546 -13594 17598
rect -13542 17590 -10439 17598
rect -13542 17546 -12463 17590
rect -17257 17538 -12463 17546
rect -12411 17538 -12339 17590
rect -12287 17538 -12215 17590
rect -12163 17538 -12091 17590
rect -12039 17538 -10439 17590
rect -17257 17474 -10439 17538
rect -17257 17449 -13966 17474
rect -15247 17422 -13966 17449
rect -13914 17422 -13842 17474
rect -13790 17422 -13718 17474
rect -13666 17422 -13594 17474
rect -13542 17466 -10439 17474
rect -13542 17422 -12463 17466
rect -15247 17414 -12463 17422
rect -12411 17414 -12339 17466
rect -12287 17414 -12215 17466
rect -12163 17414 -12091 17466
rect -12039 17414 -10439 17466
rect -15247 17350 -10439 17414
rect -15247 17298 -13966 17350
rect -13914 17298 -13842 17350
rect -13790 17298 -13718 17350
rect -13666 17298 -13594 17350
rect -13542 17342 -10439 17350
rect -13542 17298 -12463 17342
rect -15247 17290 -12463 17298
rect -12411 17290 -12339 17342
rect -12287 17290 -12215 17342
rect -12163 17290 -12091 17342
rect -12039 17290 -10439 17342
rect -15247 16941 -10439 17290
rect -5404 18033 23162 18506
rect -5404 15562 -4931 18033
rect 9800 17596 10310 17660
rect 9800 17544 9836 17596
rect 9888 17544 9964 17596
rect 10016 17593 10310 17596
rect 10016 17544 10115 17593
rect 9800 17541 10115 17544
rect 10167 17541 10310 17593
rect 9800 17482 10310 17541
rect 7638 17437 10310 17482
rect 7638 17385 9834 17437
rect 9886 17435 10181 17437
rect 9886 17385 10005 17435
rect 7638 17383 10005 17385
rect 10057 17385 10181 17435
rect 10233 17385 10310 17437
rect 10057 17383 10310 17385
rect 7638 17338 10310 17383
rect 7638 16685 7782 17338
rect 9800 17274 10310 17338
rect 9800 17258 10197 17274
rect 9800 17253 10048 17258
rect 9800 17201 9846 17253
rect 9898 17206 10048 17253
rect 10100 17222 10197 17258
rect 10249 17222 10310 17274
rect 10100 17206 10310 17222
rect 9898 17201 10310 17206
rect 9800 17160 10310 17201
rect 4098 16541 7782 16685
rect 9750 16933 10260 16990
rect 9750 16926 10054 16933
rect 9750 16923 9923 16926
rect 9750 16871 9795 16923
rect 9847 16874 9923 16923
rect 9975 16881 10054 16926
rect 10106 16881 10260 16933
rect 9975 16874 10260 16881
rect 9847 16871 10260 16874
rect 9750 16749 10260 16871
rect 9750 16744 10107 16749
rect 9750 16726 9959 16744
rect 9750 16674 9790 16726
rect 9842 16692 9959 16726
rect 10011 16697 10107 16744
rect 10159 16697 10260 16749
rect 10011 16692 10260 16697
rect 9842 16674 10260 16692
rect 9750 16616 10260 16674
rect 9750 16606 10141 16616
rect 9750 16575 9964 16606
rect 9750 16523 9767 16575
rect 9819 16554 9964 16575
rect 10016 16564 10141 16606
rect 10193 16564 10260 16616
rect 10016 16554 10260 16564
rect 9819 16523 10260 16554
rect 9750 16490 10260 16523
rect 1520 15970 1593 16058
rect 1320 15880 1398 15964
rect -17080 15089 -4931 15562
rect 1740 15510 1998 15563
rect 1863 15507 1996 15510
rect 9778 15355 9980 16490
rect 1530 15295 2126 15296
rect 1530 15240 2128 15295
rect 1532 15239 2128 15240
rect 3928 15153 9980 15355
rect 13774 16462 14012 16506
rect 22689 16495 23162 18033
rect 13774 16312 21382 16462
rect 3968 14741 4219 14775
rect 3968 14689 4007 14741
rect 4059 14689 4134 14741
rect 4186 14689 4219 14741
rect 3968 14651 4219 14689
rect 11733 14403 11992 14405
rect 2167 13969 7519 14172
rect -16003 13352 -12360 13755
rect -17855 13273 -12360 13352
rect -17855 13252 -14237 13273
rect -17855 13200 -15546 13252
rect -15494 13200 -15422 13252
rect -15370 13200 -15298 13252
rect -15246 13200 -15174 13252
rect -15122 13221 -14237 13252
rect -14185 13221 -14113 13273
rect -14061 13221 -13989 13273
rect -13937 13221 -13865 13273
rect -13813 13221 -12360 13273
rect -15122 13200 -12360 13221
rect -17855 13149 -12360 13200
rect -17855 13128 -14237 13149
rect -17855 13076 -15546 13128
rect -15494 13076 -15422 13128
rect -15370 13076 -15298 13128
rect -15246 13076 -15174 13128
rect -15122 13097 -14237 13128
rect -14185 13097 -14113 13149
rect -14061 13097 -13989 13149
rect -13937 13097 -13865 13149
rect -13813 13097 -12360 13149
rect -15122 13076 -12360 13097
rect -17855 13025 -12360 13076
rect -17855 13004 -14237 13025
rect -17855 12952 -15546 13004
rect -15494 12952 -15422 13004
rect -15370 12952 -15298 13004
rect -15246 12952 -15174 13004
rect -15122 12973 -14237 13004
rect -14185 12973 -14113 13025
rect -14061 12973 -13989 13025
rect -13937 12973 -13865 13025
rect -13813 12973 -12360 13025
rect -15122 12952 -12360 12973
rect -17855 12901 -12360 12952
rect -17855 12880 -14237 12901
rect -17855 12828 -15546 12880
rect -15494 12828 -15422 12880
rect -15370 12828 -15298 12880
rect -15246 12828 -15174 12880
rect -15122 12849 -14237 12880
rect -14185 12849 -14113 12901
rect -14061 12849 -13989 12901
rect -13937 12849 -13865 12901
rect -13813 12849 -12360 12901
rect -15122 12828 -12360 12849
rect -17855 12710 -12360 12828
rect -16003 12531 -12360 12710
rect 5930 11533 6133 13969
rect 6482 11515 6685 13969
rect 7316 11533 7519 13969
rect 9781 13966 11992 14403
rect 9781 11862 10218 13966
rect 11532 13843 11992 13966
rect 10844 13450 11116 13516
rect 10844 13398 10858 13450
rect 10910 13398 10996 13450
rect 11048 13398 11116 13450
rect 10844 13323 11116 13398
rect 10844 13271 10861 13323
rect 10913 13321 11116 13323
rect 10913 13271 11000 13321
rect 10844 13269 11000 13271
rect 11052 13269 11116 13321
rect 10844 13252 11116 13269
rect 10844 13212 11222 13252
rect 12351 13241 12512 13253
rect 10844 13179 11335 13212
rect 12222 13195 12512 13241
rect 12351 13184 12512 13195
rect 10844 13170 11000 13179
rect 10844 13118 10860 13170
rect 10912 13127 11000 13170
rect 11052 13140 11335 13179
rect 11052 13127 11222 13140
rect 10912 13118 11222 13127
rect 10844 13100 11222 13118
rect 10999 12899 11286 12914
rect 10999 12862 12306 12899
rect 10999 12810 11046 12862
rect 11098 12810 11184 12862
rect 11236 12810 12306 12862
rect 10999 12754 12306 12810
rect 10999 12730 11286 12754
rect 10999 12678 11173 12730
rect 11225 12678 11286 12730
rect 10999 12626 11286 12678
rect 12387 12469 12512 13184
rect 12257 12415 12529 12469
rect 12257 12363 12271 12415
rect 12323 12363 12409 12415
rect 12461 12363 12529 12415
rect 12257 12288 12529 12363
rect 12257 12236 12274 12288
rect 12326 12286 12529 12288
rect 12326 12236 12413 12286
rect 12257 12234 12413 12236
rect 12465 12234 12529 12286
rect 12257 12217 12529 12234
rect 12257 12144 12533 12217
rect 12257 12135 12413 12144
rect 12257 12083 12273 12135
rect 12325 12092 12413 12135
rect 12465 12092 12533 12144
rect 12325 12083 12533 12092
rect 12257 12065 12533 12083
rect 8578 11665 8995 11731
rect 8578 11662 8876 11665
rect 8578 11661 8731 11662
rect 8578 11609 8609 11661
rect 8661 11610 8731 11661
rect 8783 11613 8876 11662
rect 8928 11613 8995 11665
rect 8783 11610 8995 11613
rect 8661 11609 8995 11610
rect 8578 11550 8995 11609
rect 9781 11564 12433 11862
rect 8578 11549 8746 11550
rect 8578 11497 8615 11549
rect 8667 11498 8746 11549
rect 8798 11498 8885 11550
rect 8937 11498 8995 11550
rect 8667 11497 8995 11498
rect 8578 11491 8995 11497
rect 9959 11492 12433 11564
rect 8561 11488 8995 11491
rect 1646 10690 2266 10779
rect 2407 10345 2529 10437
rect -9592 9631 -8737 9680
rect -9592 9579 -9354 9631
rect -9302 9579 -8805 9631
rect -8753 9579 -8737 9631
rect -9592 9519 -8737 9579
rect -9574 8915 -8717 8964
rect -9574 8863 -9334 8915
rect -9282 8863 -8785 8915
rect -8733 8863 -8717 8915
rect -9574 8803 -8717 8863
rect -488 7484 -184 10115
rect 11236 9990 11632 10070
rect 11236 9979 11521 9990
rect 11236 9927 11344 9979
rect 11396 9938 11521 9979
rect 11573 9938 11632 9990
rect 11396 9927 11632 9938
rect 11236 9858 11632 9927
rect 11236 9848 11414 9858
rect 11236 9796 11278 9848
rect 11330 9806 11414 9848
rect 11466 9853 11632 9858
rect 11466 9806 11561 9853
rect 11330 9801 11561 9806
rect 11613 9801 11632 9853
rect 11330 9796 11632 9801
rect 11236 9772 11632 9796
rect 3173 9217 5247 9311
rect 3173 9045 3267 9217
rect 2329 8964 3267 9045
rect 2329 8912 2389 8964
rect 2441 8912 2711 8964
rect 2763 8912 3267 8964
rect 2329 8790 3267 8912
rect 12063 8509 12433 11492
rect 11423 7982 11671 8029
rect 11423 7930 11440 7982
rect 11492 7930 11574 7982
rect 11626 7930 11671 7982
rect 11423 7894 11671 7930
rect 12747 7909 13129 7920
rect 11423 7874 11740 7894
rect 11423 7868 11837 7874
rect 11423 7816 11435 7868
rect 11487 7856 11837 7868
rect 11487 7816 11564 7856
rect 11423 7804 11564 7816
rect 11616 7804 11837 7856
rect 12692 7851 13129 7909
rect 11423 7802 11837 7804
rect 11423 7782 11740 7802
rect 12747 7798 13129 7851
rect 11423 7781 11671 7782
rect 5341 7484 5645 7666
rect -488 7366 5645 7484
rect -1513 7255 5645 7366
rect 10977 7473 11090 7643
rect 10977 7360 11833 7473
rect 13007 7311 13129 7798
rect -1513 7252 1047 7255
rect -1513 7231 644 7252
rect -1513 7179 137 7231
rect 189 7200 644 7231
rect 696 7203 1047 7252
rect 1099 7203 5645 7255
rect 696 7200 5645 7203
rect 189 7180 5645 7200
rect 12940 7305 13192 7311
rect 12940 7253 12966 7305
rect 13018 7253 13102 7305
rect 13154 7253 13192 7305
rect 12940 7192 13192 7253
rect 189 7179 1309 7180
rect -1513 6968 1309 7179
rect 12940 7140 12961 7192
rect 13013 7185 13192 7192
rect 13013 7140 13097 7185
rect -1513 6961 910 6968
rect -1513 6923 511 6961
rect -1513 6871 95 6923
rect 147 6909 511 6923
rect 563 6916 910 6961
rect 962 6916 1309 6968
rect 563 6909 1309 6916
rect 147 6871 1309 6909
rect 8560 7073 9108 7137
rect 12940 7133 13097 7140
rect 13149 7133 13192 7185
rect 12940 7111 13192 7133
rect 8560 7068 8953 7073
rect 8560 7016 8598 7068
rect 8650 7016 8741 7068
rect 8793 7021 8953 7068
rect 9005 7021 9108 7073
rect 8793 7016 9108 7021
rect 8560 6956 9108 7016
rect 8560 6904 8598 6956
rect 8650 6904 8746 6956
rect 8798 6904 8984 6956
rect 9036 6904 9108 6956
rect 8560 6879 9108 6904
rect -1513 6646 1309 6871
rect -1513 6632 998 6646
rect -1513 6608 644 6632
rect -1513 6604 266 6608
rect -1513 6552 -7 6604
rect 45 6556 266 6604
rect 318 6580 644 6608
rect 696 6594 998 6632
rect 1050 6594 1309 6646
rect 696 6580 1309 6594
rect 318 6556 1309 6580
rect 45 6552 1309 6556
rect -1513 6250 1309 6552
rect -1513 6187 1298 6250
rect -1513 6135 620 6187
rect 672 6135 1298 6187
rect -1513 5811 1298 6135
rect 12397 5486 12483 5488
rect 12397 5403 12791 5486
rect 12397 5392 12679 5403
rect 12397 5340 12502 5392
rect 12554 5351 12679 5392
rect 12731 5351 12791 5403
rect 12554 5340 12791 5351
rect 12397 5271 12791 5340
rect 12397 5261 12572 5271
rect 12397 5209 12436 5261
rect 12488 5219 12572 5261
rect 12624 5266 12791 5271
rect 12624 5219 12719 5266
rect 12488 5214 12719 5219
rect 12771 5214 12791 5266
rect 12488 5209 12791 5214
rect 12397 5185 12791 5209
rect -9554 4579 6428 4675
rect 4463 3808 5878 3909
rect 4463 3805 5616 3808
rect 4463 3784 5213 3805
rect 4463 3732 4706 3784
rect 4758 3753 5213 3784
rect 5265 3756 5616 3805
rect 5668 3756 5878 3808
rect 5265 3753 5878 3756
rect 4758 3732 5878 3753
rect 4463 3521 5878 3732
rect 4463 3514 5479 3521
rect 4463 3476 5080 3514
rect 4463 3424 4664 3476
rect 4716 3462 5080 3476
rect 5132 3469 5479 3514
rect 5531 3469 5878 3521
rect 5132 3462 5878 3469
rect 4716 3424 5878 3462
rect 4463 3199 5878 3424
rect 4463 3185 5567 3199
rect 4463 3161 5213 3185
rect 4463 3157 4835 3161
rect 4463 3105 4562 3157
rect 4614 3109 4835 3157
rect 4887 3133 5213 3161
rect 5265 3147 5567 3185
rect 5619 3147 5878 3199
rect 5265 3133 5878 3147
rect 4887 3109 5878 3133
rect 4614 3105 5878 3109
rect 4463 3077 5878 3105
rect 4463 2954 6454 3077
rect 4463 2905 5878 2954
rect 13774 2751 14012 16312
rect -9407 2513 14012 2751
rect 16352 15363 19534 15786
rect 16352 2170 16775 15363
rect 17927 14293 18154 14470
rect 17890 14268 18200 14293
rect 17890 14008 17931 14268
rect 18191 14008 18200 14268
rect 17890 13943 18200 14008
rect 17890 13787 17919 13943
rect 18179 13787 18200 13943
rect 17890 13738 18200 13787
rect 19111 14167 19534 15363
rect 19111 14115 19181 14167
rect 19233 14115 19412 14167
rect 19464 14115 19534 14167
rect 20406 14143 20600 14210
rect 20393 14129 20705 14143
rect 19111 13953 19534 14115
rect 19111 13901 19179 13953
rect 19231 13901 19401 13953
rect 19453 13901 19534 13953
rect 19111 13731 19534 13901
rect 20370 14091 20705 14129
rect 20370 13831 20393 14091
rect 20653 13831 20705 14091
rect 20370 13811 20705 13831
rect 19111 13723 19389 13731
rect 19111 13671 19178 13723
rect 19230 13679 19389 13723
rect 19441 13679 19534 13731
rect 19230 13671 19534 13679
rect 19111 13591 19534 13671
rect 21232 13292 21382 16312
rect 22689 16431 23393 16495
rect 22689 16379 22822 16431
rect 22874 16379 22942 16431
rect 22994 16379 23062 16431
rect 23114 16379 23182 16431
rect 23234 16379 23302 16431
rect 23354 16379 23393 16431
rect 22689 16311 23393 16379
rect 22689 16259 22822 16311
rect 22874 16259 22942 16311
rect 22994 16259 23062 16311
rect 23114 16259 23182 16311
rect 23234 16259 23302 16311
rect 23354 16259 23393 16311
rect 22689 16210 23393 16259
rect 22079 15270 22652 15272
rect 21918 15250 22652 15270
rect 21918 15198 22094 15250
rect 22146 15198 22214 15250
rect 22266 15198 22334 15250
rect 22386 15198 22454 15250
rect 22506 15198 22574 15250
rect 22626 15198 22652 15250
rect 21918 15130 22652 15198
rect 21918 15078 22094 15130
rect 22146 15078 22214 15130
rect 22266 15078 22334 15130
rect 22386 15078 22454 15130
rect 22506 15078 22574 15130
rect 22626 15078 22652 15130
rect 21918 15051 22652 15078
rect 21918 15049 22491 15051
rect 22045 14662 22661 14694
rect 21999 14632 22694 14662
rect 21999 14580 22063 14632
rect 22115 14580 22183 14632
rect 22235 14580 22303 14632
rect 22355 14580 22423 14632
rect 22475 14580 22543 14632
rect 22595 14580 22694 14632
rect 21999 14512 22694 14580
rect 21999 14470 22063 14512
rect 22045 14460 22063 14470
rect 22115 14460 22183 14512
rect 22235 14460 22303 14512
rect 22355 14460 22423 14512
rect 22475 14460 22543 14512
rect 22595 14470 22694 14512
rect 22595 14460 22661 14470
rect 22045 14427 22661 14460
rect 24392 14135 24914 19038
rect 95781 18452 96117 18466
rect 95781 18400 95813 18452
rect 95865 18400 95933 18452
rect 95985 18400 96053 18452
rect 96105 18400 96117 18452
rect 95781 18396 96117 18400
rect 95781 18332 96232 18396
rect 95781 18280 95813 18332
rect 95865 18280 95933 18332
rect 95985 18280 96053 18332
rect 96105 18280 96232 18332
rect 95781 18236 96232 18280
rect 95781 18212 96117 18236
rect 95781 18160 95813 18212
rect 95865 18160 95933 18212
rect 95985 18160 96053 18212
rect 96105 18160 96117 18212
rect 95781 18126 96117 18160
rect 26344 16826 26987 16880
rect 26344 16802 26428 16826
rect 26285 16774 26428 16802
rect 26480 16774 26548 16826
rect 26600 16774 26668 16826
rect 26720 16774 26788 16826
rect 26840 16774 26908 16826
rect 26960 16774 26987 16826
rect 26285 16706 26987 16774
rect 26285 16654 26428 16706
rect 26480 16654 26548 16706
rect 26600 16654 26668 16706
rect 26720 16654 26788 16706
rect 26840 16654 26908 16706
rect 26960 16654 26987 16706
rect 26285 16626 26987 16654
rect 26344 16591 26987 16626
rect 95893 16826 96229 16840
rect 95893 16774 95925 16826
rect 95977 16774 96045 16826
rect 96097 16774 96165 16826
rect 96217 16774 96229 16826
rect 95893 16770 96229 16774
rect 95893 16706 96344 16770
rect 95893 16654 95925 16706
rect 95977 16654 96045 16706
rect 96097 16654 96165 16706
rect 96217 16654 96344 16706
rect 95893 16610 96344 16654
rect 95893 16586 96229 16610
rect 95893 16534 95925 16586
rect 95977 16534 96045 16586
rect 96097 16534 96165 16586
rect 96217 16534 96229 16586
rect 95893 16489 96229 16534
rect 66781 15482 88697 15857
rect 22087 14087 24914 14135
rect 21918 14084 24914 14087
rect 21918 13928 22116 14084
rect 22272 13928 22498 14084
rect 22654 13928 22917 14084
rect 23073 13928 24914 14084
rect 21918 13926 24914 13928
rect 22087 13910 24914 13926
rect 28009 14158 45862 14382
rect 28009 14106 37935 14158
rect 37987 14106 38055 14158
rect 38107 14106 38175 14158
rect 38227 14106 38295 14158
rect 38347 14106 38415 14158
rect 38467 14106 45862 14158
rect 28009 14038 45862 14106
rect 28009 13986 37935 14038
rect 37987 13986 38055 14038
rect 38107 13986 38175 14038
rect 38227 13986 38295 14038
rect 38347 13986 38415 14038
rect 38467 13986 45862 14038
rect 28009 13917 45862 13986
rect 22087 13904 24841 13910
rect 21938 13658 22849 13700
rect 21833 13616 22849 13658
rect 21833 13564 22006 13616
rect 22058 13564 22429 13616
rect 22481 13564 22720 13616
rect 22772 13564 22849 13616
rect 21833 13522 22849 13564
rect 21938 13497 22849 13522
rect 21232 13239 22530 13292
rect 21232 13187 21838 13239
rect 21890 13187 22077 13239
rect 22129 13187 22410 13239
rect 22462 13187 22530 13239
rect 21232 13142 22530 13187
rect 28009 13000 28474 13917
rect 29826 13325 30426 13389
rect 29826 13323 29830 13325
rect 29802 13273 29830 13323
rect 29882 13273 29950 13325
rect 30002 13273 30070 13325
rect 30122 13273 30190 13325
rect 30242 13273 30310 13325
rect 30362 13323 30426 13325
rect 30362 13273 31638 13323
rect 29802 13205 31638 13273
rect 29802 13153 29830 13205
rect 29882 13153 29950 13205
rect 30002 13153 30070 13205
rect 30122 13153 30190 13205
rect 30242 13153 30310 13205
rect 30362 13153 31638 13205
rect 29802 13134 31638 13153
rect 28009 12882 28470 13000
rect 22767 12489 24077 12615
rect 25831 12525 28470 12882
rect 22767 12487 23800 12489
rect 22767 12486 23246 12487
rect 22823 12412 22947 12486
rect 23122 12412 23246 12486
rect 23406 12412 23530 12487
rect 23676 12412 23800 12487
rect 23953 12412 24077 12489
rect 25830 12503 28470 12525
rect 25830 12433 26744 12503
rect 24624 12412 24967 12413
rect 25540 12412 25770 12413
rect 25830 12412 26545 12433
rect 22793 11960 26545 12412
rect 23396 11515 23551 11668
rect 26224 11549 26277 11586
rect 22449 11211 22560 11220
rect 19654 11188 19738 11204
rect 19654 11136 19670 11188
rect 19722 11136 19738 11188
rect 19654 11121 19738 11136
rect 19895 11193 19979 11209
rect 19895 11141 19911 11193
rect 19963 11141 19979 11193
rect 19895 11126 19979 11141
rect 20134 11195 20218 11211
rect 20134 11143 20150 11195
rect 20202 11143 20218 11195
rect 20134 11139 20218 11143
rect 20206 11128 20218 11139
rect 20361 11195 20445 11211
rect 20361 11143 20377 11195
rect 20429 11143 20445 11195
rect 20361 11128 20445 11143
rect 22449 11167 22956 11211
rect 22449 11115 22481 11167
rect 22533 11115 22956 11167
rect 22449 11110 22956 11115
rect 22449 11023 22560 11110
rect 22449 10971 22476 11023
rect 22528 10971 22560 11023
rect 22449 10942 22560 10971
rect 23689 10953 23771 11033
rect 18271 9770 18472 10580
rect 21819 10516 22140 10575
rect 21819 10334 22833 10516
rect 31449 10181 31638 13134
rect 31886 11708 32351 13917
rect 44097 13320 44562 13917
rect 45397 13320 45862 13917
rect 64769 13772 65603 13916
rect 64769 13720 64929 13772
rect 64981 13768 65603 13772
rect 64981 13720 65188 13768
rect 64769 13718 65188 13720
rect 47691 13716 65188 13718
rect 65240 13716 65603 13768
rect 47691 13703 65603 13716
rect 47691 13651 65429 13703
rect 65481 13651 65603 13703
rect 47691 13621 65603 13651
rect 47691 13569 64933 13621
rect 64985 13591 65603 13621
rect 64985 13569 65200 13591
rect 47691 13539 65200 13569
rect 65252 13550 65603 13591
rect 65252 13539 65424 13550
rect 47691 13498 65424 13539
rect 65476 13498 65603 13550
rect 47691 13454 65603 13498
rect 47691 13452 65190 13454
rect 47691 13400 64932 13452
rect 64984 13402 65190 13452
rect 65242 13407 65603 13454
rect 65242 13402 65422 13407
rect 64984 13400 65422 13402
rect 47691 13355 65422 13400
rect 65474 13355 65603 13407
rect 47691 13277 65603 13355
rect 47691 13225 64982 13277
rect 65034 13272 65603 13277
rect 65034 13225 65184 13272
rect 47691 13220 65184 13225
rect 65236 13260 65603 13272
rect 65236 13220 65347 13260
rect 47691 13208 65347 13220
rect 65399 13208 65603 13260
rect 47691 13149 65603 13208
rect 41677 12634 41885 12734
rect 41677 12582 41755 12634
rect 41807 12582 41885 12634
rect 41677 12384 41885 12582
rect 41677 12332 41755 12384
rect 41807 12378 41885 12384
rect 41807 12332 42113 12378
rect 41677 12160 42113 12332
rect 41677 12108 41755 12160
rect 41807 12108 42113 12160
rect 41677 12061 42113 12108
rect 33300 11005 33380 11085
rect 33768 11014 33853 11090
rect 37793 10784 38571 10840
rect 37793 10732 37877 10784
rect 37929 10732 37997 10784
rect 38049 10732 38117 10784
rect 38169 10732 38237 10784
rect 38289 10732 38357 10784
rect 38409 10732 38571 10784
rect 37793 10664 38571 10732
rect 37793 10612 37877 10664
rect 37929 10612 37997 10664
rect 38049 10612 38117 10664
rect 38169 10612 38237 10664
rect 38289 10612 38357 10664
rect 38409 10612 38571 10664
rect 37793 10547 38571 10612
rect 19888 9897 22600 10122
rect 31449 10073 32313 10181
rect 31449 9975 31638 10073
rect 28770 9909 28848 9964
rect 29009 9914 29087 9964
rect 29248 9916 29326 9964
rect 29474 9916 29552 9964
rect 22373 9505 22600 9897
rect 28768 9893 28852 9909
rect 28768 9841 28784 9893
rect 28836 9841 28852 9893
rect 28768 9826 28852 9841
rect 29009 9898 29093 9914
rect 29009 9846 29025 9898
rect 29077 9846 29093 9898
rect 29009 9831 29093 9846
rect 29248 9900 29332 9916
rect 29248 9848 29264 9900
rect 29316 9848 29332 9900
rect 29248 9833 29332 9848
rect 29474 9900 29559 9916
rect 29474 9848 29491 9900
rect 29543 9848 29559 9900
rect 29474 9833 29559 9848
rect 28770 9794 28848 9826
rect 29009 9794 29087 9831
rect 29248 9794 29326 9833
rect 29474 9794 29552 9833
rect 22373 9472 22743 9505
rect 22373 9390 22985 9472
rect 22373 9358 22743 9390
rect 19614 9158 19692 9209
rect 19853 9163 19931 9209
rect 20318 9165 20396 9209
rect 19612 9142 19696 9158
rect 19612 9090 19628 9142
rect 19680 9090 19696 9142
rect 19612 9075 19696 9090
rect 19853 9147 19937 9163
rect 19853 9095 19869 9147
rect 19921 9095 19937 9147
rect 19853 9080 19937 9095
rect 20092 9149 20176 9153
rect 20092 9097 20108 9149
rect 20160 9097 20176 9149
rect 20092 9082 20176 9097
rect 20318 9149 20403 9165
rect 20318 9097 20335 9149
rect 20387 9097 20403 9149
rect 20318 9082 20403 9097
rect 19614 9039 19692 9075
rect 19853 9039 19931 9080
rect 20092 9039 20170 9082
rect 20318 9039 20396 9082
rect 26167 8889 26249 8932
rect 28228 8584 28434 9476
rect 30473 8717 30883 9048
rect 26351 8450 26523 8578
rect 22178 8009 22619 8152
rect 18490 7270 18630 7690
rect 22476 7354 22619 8009
rect 22865 7922 22989 8384
rect 23323 7922 23447 8384
rect 24418 7922 24542 8396
rect 25281 7922 25405 8393
rect 25975 7922 26099 8413
rect 26224 8326 26523 8450
rect 26343 8324 26523 8326
rect 26351 7922 26523 8324
rect 22840 7881 26523 7922
rect 22840 7879 23419 7881
rect 22840 7874 23180 7879
rect 22840 7822 22939 7874
rect 22991 7827 23180 7874
rect 23232 7829 23419 7879
rect 23471 7829 23646 7881
rect 23698 7829 26523 7881
rect 23232 7827 26523 7829
rect 22991 7822 26523 7827
rect 22840 7798 26523 7822
rect 26351 7706 26523 7798
rect 22476 7211 26978 7354
rect 28714 6915 28792 6970
rect 28953 6920 29031 6970
rect 29192 6922 29270 6970
rect 29418 6922 29496 6970
rect 28712 6899 28796 6915
rect 17937 6751 18038 6809
rect 20377 6789 22546 6850
rect 28712 6847 28728 6899
rect 28780 6847 28796 6899
rect 28712 6832 28796 6847
rect 28953 6904 29037 6920
rect 28953 6852 28969 6904
rect 29021 6852 29037 6904
rect 28953 6837 29037 6852
rect 29192 6906 29276 6922
rect 29192 6854 29208 6906
rect 29260 6854 29276 6906
rect 29192 6839 29276 6854
rect 29418 6906 29503 6922
rect 29418 6854 29435 6906
rect 29487 6854 29503 6906
rect 29418 6839 29503 6854
rect 28714 6800 28792 6832
rect 28953 6800 29031 6837
rect 29192 6800 29270 6839
rect 29418 6800 29496 6839
rect 17937 6711 19507 6751
rect 20377 6737 22134 6789
rect 22186 6737 22430 6789
rect 22482 6737 22546 6789
rect 17937 6670 19508 6711
rect 17937 6646 18072 6670
rect 17938 6618 18072 6646
rect 18124 6618 18192 6670
rect 18244 6618 18312 6670
rect 18364 6618 18432 6670
rect 18484 6618 18552 6670
rect 18604 6618 18672 6670
rect 18724 6618 18792 6670
rect 18844 6618 18912 6670
rect 18964 6618 19032 6670
rect 19084 6618 19152 6670
rect 19204 6618 19272 6670
rect 19324 6618 19392 6670
rect 19444 6618 19508 6670
rect 17938 6585 19508 6618
rect 20377 6705 22546 6737
rect 20377 6083 20564 6705
rect 22083 6683 22546 6705
rect 18154 6014 20564 6083
rect 18154 6011 18892 6014
rect 18154 5959 18232 6011
rect 18284 6009 18892 6011
rect 18284 5959 18410 6009
rect 18154 5957 18410 5959
rect 18462 6008 18892 6009
rect 18462 5957 18651 6008
rect 18154 5956 18651 5957
rect 18703 5962 18892 6008
rect 18944 5962 20564 6014
rect 18703 5956 20564 5962
rect 18154 5896 20564 5956
rect 27871 5059 28268 6488
rect 28962 6257 29078 6331
rect 31485 6257 31602 9975
rect 32011 9879 32303 9911
rect 32011 9827 32075 9879
rect 32127 9827 32303 9879
rect 32011 9792 32303 9827
rect 33754 9608 33830 9683
rect 33953 8907 34341 9396
rect 36812 8907 37200 10205
rect 33953 8519 37200 8907
rect 28962 6141 31602 6257
rect 32225 5373 32329 5795
rect 35051 5043 35609 8519
rect 47691 8399 48260 13149
rect 64769 13020 65603 13149
rect 47690 8228 48260 8399
rect 47690 8176 47793 8228
rect 47845 8176 47949 8228
rect 48001 8176 48260 8228
rect 47690 7940 48260 8176
rect 50084 9609 57840 9830
rect 50084 7719 50305 9609
rect 53921 9316 54794 9377
rect 53921 9315 54374 9316
rect 53921 9314 54252 9315
rect 53921 9262 54014 9314
rect 54066 9262 54133 9314
rect 54185 9263 54252 9314
rect 54304 9264 54374 9315
rect 54426 9315 54794 9316
rect 54426 9264 54492 9315
rect 54304 9263 54492 9264
rect 54544 9263 54794 9315
rect 54185 9262 54794 9263
rect 53921 9199 54794 9262
rect 53921 9197 54374 9199
rect 53921 9196 54254 9197
rect 53921 9144 54014 9196
rect 54066 9144 54133 9196
rect 54185 9145 54254 9196
rect 54306 9147 54374 9197
rect 54426 9195 54794 9199
rect 54426 9147 54493 9195
rect 54306 9145 54493 9147
rect 54185 9144 54493 9145
rect 53921 9143 54493 9144
rect 54545 9143 54794 9195
rect 53921 9088 54794 9143
rect 43227 7112 43321 7123
rect 46153 7119 46241 7356
rect 46418 7119 46522 7356
rect 46706 7119 46809 7356
rect 46908 7188 47005 7356
rect 50084 7338 50292 7719
rect 46908 7119 47009 7188
rect 48084 7130 50292 7338
rect 57619 7531 57840 9609
rect 61491 9323 62361 9385
rect 61491 9322 61944 9323
rect 61491 9321 61822 9322
rect 61491 9269 61584 9321
rect 61636 9269 61703 9321
rect 61755 9270 61822 9321
rect 61874 9271 61944 9322
rect 61996 9322 62361 9323
rect 61996 9271 62062 9322
rect 61874 9270 62062 9271
rect 62114 9270 62361 9322
rect 61755 9269 62361 9270
rect 61491 9206 62361 9269
rect 61491 9204 61944 9206
rect 61491 9203 61824 9204
rect 61491 9151 61584 9203
rect 61636 9151 61703 9203
rect 61755 9152 61824 9203
rect 61876 9154 61944 9204
rect 61996 9202 62361 9206
rect 61996 9154 62063 9202
rect 61876 9152 62063 9154
rect 61755 9151 62063 9152
rect 61491 9150 62063 9151
rect 62115 9150 62361 9202
rect 61491 9099 62361 9150
rect 58049 7531 58270 8320
rect 66783 7933 67158 15482
rect 57619 7310 58270 7531
rect 43227 7111 43449 7112
rect 43820 7111 43992 7112
rect 43227 7104 44714 7111
rect 43227 6948 43285 7104
rect 43441 6948 43828 7104
rect 43984 6948 44538 7104
rect 44694 6948 44714 7104
rect 46136 7078 47059 7119
rect 46136 7073 46937 7078
rect 46136 7021 46195 7073
rect 46247 7070 46937 7073
rect 46247 7068 46721 7070
rect 46247 7021 46441 7068
rect 46136 7016 46441 7021
rect 46493 7018 46721 7068
rect 46773 7026 46937 7070
rect 46989 7026 47059 7078
rect 46773 7018 47059 7026
rect 46493 7016 47059 7018
rect 46136 6961 47059 7016
rect 43227 6941 44714 6948
rect 43227 6940 43449 6941
rect 43820 6940 43992 6941
rect 43227 6919 43321 6940
rect 38263 6633 39669 6671
rect 38263 6608 39913 6633
rect 38263 6452 39342 6608
rect 39498 6452 39913 6608
rect 38263 6430 39913 6452
rect 38287 6427 39913 6430
rect 38287 6418 39669 6427
rect 38287 6414 38493 6418
rect 43759 6074 44718 6127
rect 43759 6022 43825 6074
rect 43877 6061 44718 6074
rect 43877 6022 44074 6061
rect 43759 6009 44074 6022
rect 44126 6060 44718 6061
rect 44126 6056 44530 6060
rect 44126 6009 44308 6056
rect 43759 6004 44308 6009
rect 44360 6008 44530 6056
rect 44582 6008 44718 6060
rect 44360 6004 44718 6008
rect 43759 5971 44718 6004
rect 40396 4708 42297 5056
rect 30400 4487 30604 4659
rect 27094 4405 27485 4463
rect 27094 4353 27149 4405
rect 27201 4353 27381 4405
rect 27433 4353 27485 4405
rect 27094 4209 27485 4353
rect 30400 4435 30470 4487
rect 30522 4435 30604 4487
rect 30400 4263 30604 4435
rect 27094 4157 27146 4209
rect 27198 4157 27381 4209
rect 27433 4157 27485 4209
rect 27094 4108 27485 4157
rect 30300 4226 30604 4263
rect 42800 4230 42910 4490
rect 30300 4174 30470 4226
rect 30522 4174 30604 4226
rect 43290 4210 43400 4470
rect 30300 4138 30604 4174
rect 30400 4129 30604 4138
rect 27110 3940 27240 4108
rect 48084 2343 48292 7130
rect 50084 6664 50292 7130
rect 56775 6803 57334 6920
rect 56775 6797 57017 6803
rect 56775 6792 56834 6797
rect 56251 6745 56834 6792
rect 56886 6751 57017 6797
rect 57069 6751 57204 6803
rect 57256 6751 57334 6803
rect 56886 6745 57334 6751
rect 56251 6721 57334 6745
rect 56775 6641 57334 6721
rect 58049 6680 58270 7310
rect 66784 6887 67156 7933
rect 64336 6799 67156 6887
rect 64234 6728 67156 6799
rect 64336 6639 67156 6728
rect 56294 5050 58424 5232
rect 53695 4662 54568 4724
rect 53695 4661 54148 4662
rect 53695 4660 54026 4661
rect 53695 4608 53788 4660
rect 53840 4608 53907 4660
rect 53959 4609 54026 4660
rect 54078 4610 54148 4661
rect 54200 4661 54568 4662
rect 54200 4610 54266 4661
rect 54078 4609 54266 4610
rect 54318 4609 54568 4661
rect 53959 4608 54568 4609
rect 53695 4545 54568 4608
rect 53695 4543 54148 4545
rect 53695 4542 54028 4543
rect 53695 4490 53788 4542
rect 53840 4490 53907 4542
rect 53959 4491 54028 4542
rect 54080 4493 54148 4543
rect 54200 4541 54568 4545
rect 54200 4493 54267 4541
rect 54080 4491 54267 4493
rect 53959 4490 54267 4491
rect 53695 4489 54267 4490
rect 54319 4489 54568 4541
rect 53695 4412 54568 4489
rect 53695 4319 54344 4412
rect 53701 4315 54344 4319
rect 53701 4314 54194 4315
rect 50335 2374 50478 3627
rect 48076 2220 48292 2343
rect 50081 2231 50478 2374
rect -9320 1747 16775 2170
rect -3741 1437 -447 1445
rect -9031 1372 -447 1437
rect -9031 1358 -3106 1372
rect -9031 1098 -3695 1358
rect -3435 1112 -3106 1358
rect -2846 1112 -447 1372
rect -3435 1098 -447 1112
rect -9031 1076 -447 1098
rect -3741 1068 -447 1076
rect 47945 1007 48083 1256
rect 50081 1007 50224 2231
rect 50335 1992 50478 2231
rect 56852 2118 57411 2224
rect 56403 2107 57411 2118
rect 56403 2101 57094 2107
rect 56403 2049 56911 2101
rect 56963 2055 57094 2101
rect 57146 2055 57281 2107
rect 57333 2055 57411 2107
rect 56963 2049 57411 2055
rect 56403 2041 57411 2049
rect 56852 1945 57411 2041
rect 47943 864 50224 1007
rect -2319 300 931 372
rect -2789 299 931 300
rect -2789 287 -1728 299
rect -9055 285 -1728 287
rect -9055 25 -2317 285
rect -2057 39 -1728 285
rect -1468 39 931 299
rect -2057 25 931 39
rect -9055 24 931 25
rect -2789 14 931 24
rect -2319 -5 931 14
rect -9000 -259 3075 -188
rect 51096 -229 51474 450
rect 60742 -72 61120 5177
rect 60575 -221 61286 -72
rect 60575 -229 60991 -221
rect -9000 -311 2727 -259
rect 2779 -261 3075 -259
rect 2779 -311 2891 -261
rect -9000 -313 2891 -311
rect 2943 -313 3075 -261
rect -9000 -373 3075 -313
rect -9000 -386 2893 -373
rect -9000 -438 2727 -386
rect 2779 -425 2893 -386
rect 2945 -425 3075 -373
rect 2779 -438 3075 -425
rect -9000 -513 3075 -438
rect -9000 -524 2898 -513
rect -9000 -576 2727 -524
rect 2779 -565 2898 -524
rect 2950 -565 3075 -513
rect 2779 -576 3075 -565
rect -9000 -634 3075 -576
rect 47417 -245 60991 -229
rect 47417 -297 60715 -245
rect 60767 -273 60991 -245
rect 61043 -273 61286 -221
rect 60767 -297 61286 -273
rect 47417 -480 61286 -297
rect 47417 -483 61143 -480
rect 47417 -535 60677 -483
rect 60729 -484 61143 -483
rect 60729 -535 60900 -484
rect 47417 -536 60900 -535
rect 60952 -532 61143 -484
rect 61195 -532 61286 -480
rect 60952 -536 61286 -532
rect 47417 -607 61286 -536
rect 60575 -608 61286 -607
rect 4778 -990 5148 -932
rect 4778 -1042 4828 -990
rect 4880 -992 5148 -990
rect 4880 -1042 4992 -992
rect 4778 -1044 4992 -1042
rect 5044 -1044 5148 -992
rect 4778 -1072 5148 -1044
rect -9081 -1104 5148 -1072
rect -9081 -1117 4994 -1104
rect -9081 -1169 4828 -1117
rect 4880 -1156 4994 -1117
rect 5046 -1156 5148 -1104
rect 4880 -1169 5148 -1156
rect -9081 -1237 5148 -1169
rect 4778 -1244 5148 -1237
rect 4778 -1255 4999 -1244
rect 4778 -1307 4828 -1255
rect 4880 -1296 4999 -1255
rect 5051 -1296 5148 -1244
rect 4880 -1307 5148 -1296
rect 4778 -1338 5148 -1307
rect 4844 -1524 5214 -1512
rect -9098 -1556 5214 -1524
rect -9098 -1569 5060 -1556
rect -9098 -1621 4894 -1569
rect 4946 -1608 5060 -1569
rect 5112 -1608 5214 -1556
rect 4946 -1621 5214 -1608
rect -9098 -1689 5214 -1621
rect 18080 -1534 18860 -1470
rect 18080 -1541 18702 -1534
rect 18080 -1546 18452 -1541
rect 18080 -1598 18145 -1546
rect 18197 -1593 18452 -1546
rect 18504 -1586 18702 -1541
rect 18754 -1586 18860 -1534
rect 18504 -1593 18860 -1586
rect 18197 -1598 18860 -1593
rect 18080 -1660 18860 -1598
rect 4844 -1696 5214 -1689
rect 4844 -1707 5065 -1696
rect 4844 -1759 4894 -1707
rect 4946 -1748 5065 -1707
rect 5117 -1748 5214 -1696
rect 4946 -1759 5214 -1748
rect 4844 -1790 5214 -1759
rect 66784 -2176 67156 6639
rect 88322 -822 88697 15482
rect 95755 15638 96091 15652
rect 95755 15586 95787 15638
rect 95839 15586 95907 15638
rect 95959 15586 96027 15638
rect 96079 15586 96091 15638
rect 95755 15582 96091 15586
rect 95755 15518 96206 15582
rect 95755 15466 95787 15518
rect 95839 15466 95907 15518
rect 95959 15466 96027 15518
rect 96079 15466 96206 15518
rect 95755 15422 96206 15466
rect 95755 15398 96091 15422
rect 95755 15346 95787 15398
rect 95839 15346 95907 15398
rect 95959 15346 96027 15398
rect 96079 15346 96091 15398
rect 95755 15301 96091 15346
rect 95584 14604 96107 14621
rect 95584 14552 95801 14604
rect 95853 14552 95921 14604
rect 95973 14552 96041 14604
rect 96093 14552 96107 14604
rect 95584 14548 96107 14552
rect 95584 14484 96220 14548
rect 95584 14432 95801 14484
rect 95853 14432 95921 14484
rect 95973 14432 96041 14484
rect 96093 14432 96220 14484
rect 95584 14388 96220 14432
rect 95584 14364 96107 14388
rect 95584 14312 95801 14364
rect 95853 14312 95921 14364
rect 95973 14312 96041 14364
rect 96093 14312 96107 14364
rect 95584 14267 96107 14312
rect 98848 4719 99160 4739
rect 98848 4667 98889 4719
rect 98941 4713 99160 4719
rect 98941 4667 99064 4713
rect 98848 4661 99064 4667
rect 99116 4661 99160 4713
rect 98848 4660 99160 4661
rect 98848 4564 99482 4660
rect 98848 4560 99065 4564
rect 98848 4508 98887 4560
rect 98939 4512 99065 4560
rect 99117 4512 99482 4564
rect 98939 4508 99482 4512
rect 98848 4440 99482 4508
rect 98848 4395 99160 4440
rect 98848 4343 98890 4395
rect 98942 4390 99160 4395
rect 98942 4343 99078 4390
rect 98848 4338 99078 4343
rect 99130 4338 99160 4390
rect 91327 4255 92059 4316
rect 98848 4305 99160 4338
rect 91327 4254 91780 4255
rect 91327 4253 91658 4254
rect 91327 4201 91420 4253
rect 91472 4201 91539 4253
rect 91591 4202 91658 4253
rect 91710 4203 91780 4254
rect 91832 4254 92059 4255
rect 91832 4203 91898 4254
rect 91710 4202 91898 4203
rect 91950 4202 92059 4254
rect 91591 4201 92059 4202
rect 91327 4138 92059 4201
rect 91327 4136 91780 4138
rect 91327 4135 91660 4136
rect 91327 4083 91420 4135
rect 91472 4083 91539 4135
rect 91591 4084 91660 4135
rect 91712 4086 91780 4136
rect 91832 4134 92059 4138
rect 91832 4086 91899 4134
rect 91712 4084 91899 4086
rect 91591 4083 91899 4084
rect 91327 4082 91899 4083
rect 91951 4082 92059 4134
rect 91327 4051 92059 4082
rect 95089 2666 95620 2970
rect 95089 2614 95236 2666
rect 95288 2614 95356 2666
rect 95408 2614 95476 2666
rect 95528 2614 95620 2666
rect 95089 2546 95620 2614
rect 95089 2494 95236 2546
rect 95288 2494 95356 2546
rect 95408 2494 95476 2546
rect 95528 2494 95620 2546
rect 95089 2426 95620 2494
rect 95089 2374 95236 2426
rect 95288 2374 95356 2426
rect 95408 2374 95476 2426
rect 95528 2374 95620 2426
rect 95089 2270 95620 2374
rect 89920 -212 90106 119
rect 89820 -271 90211 -212
rect 89820 -278 90095 -271
rect 89820 -330 89881 -278
rect 89933 -323 90095 -278
rect 90147 -323 90211 -271
rect 89933 -330 90211 -323
rect 89820 -472 90211 -330
rect 89820 -524 89878 -472
rect 89930 -524 90086 -472
rect 90138 -524 90211 -472
rect 89820 -564 90211 -524
rect 4506 -2253 4874 -2240
rect 4506 -2305 4796 -2253
rect 4848 -2305 4874 -2253
rect 4506 -2330 4874 -2305
rect -8967 -2356 4874 -2330
rect -8967 -2408 4547 -2356
rect 4599 -2408 4687 -2356
rect 4739 -2408 4874 -2356
rect -8967 -2441 4874 -2408
rect 4506 -2477 4874 -2441
rect 4506 -2529 4549 -2477
rect 4601 -2480 4874 -2477
rect 4601 -2529 4695 -2480
rect 4506 -2532 4695 -2529
rect 4747 -2485 4874 -2480
rect 4747 -2532 4815 -2485
rect 4506 -2537 4815 -2532
rect 4867 -2537 4874 -2485
rect 4506 -2563 4874 -2537
rect 21848 -2548 67156 -2176
rect 87273 -1197 88697 -822
rect 5001 -2620 5371 -2608
rect -8872 -2652 5371 -2620
rect -8872 -2665 5217 -2652
rect -8872 -2717 5051 -2665
rect 5103 -2704 5217 -2665
rect 5269 -2704 5371 -2652
rect 5103 -2717 5371 -2704
rect -8872 -2785 5371 -2717
rect 5001 -2792 5371 -2785
rect 5001 -2803 5222 -2792
rect 5001 -2855 5051 -2803
rect 5103 -2844 5222 -2803
rect 5274 -2844 5371 -2792
rect 5103 -2855 5371 -2844
rect 5001 -2886 5371 -2855
rect 4905 -3038 5275 -3026
rect -8855 -3070 5275 -3038
rect -8855 -3083 5121 -3070
rect -8855 -3135 4955 -3083
rect 5007 -3122 5121 -3083
rect 5173 -3122 5275 -3070
rect 5007 -3135 5275 -3122
rect -8855 -3203 5275 -3135
rect 4905 -3210 5275 -3203
rect 4905 -3221 5126 -3210
rect 4905 -3273 4955 -3221
rect 5007 -3262 5126 -3221
rect 5178 -3262 5275 -3210
rect 5007 -3273 5275 -3262
rect 4905 -3304 5275 -3273
rect 4882 -3452 5252 -3440
rect -8942 -3484 5252 -3452
rect -8942 -3497 5098 -3484
rect -8942 -3549 4932 -3497
rect 4984 -3536 5098 -3497
rect 5150 -3536 5252 -3484
rect 4984 -3549 5252 -3536
rect -8942 -3617 5252 -3549
rect 4882 -3624 5252 -3617
rect 4882 -3635 5103 -3624
rect 4882 -3687 4932 -3635
rect 4984 -3676 5103 -3635
rect 5155 -3676 5252 -3624
rect 4984 -3687 5252 -3676
rect 4882 -3718 5252 -3687
rect 4928 -3931 5298 -3919
rect -8977 -3963 5298 -3931
rect -8977 -3976 5144 -3963
rect -8977 -4028 4978 -3976
rect 5030 -4015 5144 -3976
rect 5196 -4015 5298 -3963
rect 5030 -4028 5298 -4015
rect -8977 -4096 5298 -4028
rect 4928 -4103 5298 -4096
rect 4928 -4114 5149 -4103
rect 4928 -4166 4978 -4114
rect 5030 -4155 5149 -4114
rect 5201 -4155 5298 -4103
rect 5030 -4166 5298 -4155
rect 4928 -4197 5298 -4166
rect 5033 -4474 5403 -4462
rect -8942 -4506 5403 -4474
rect -8942 -4519 5249 -4506
rect -8942 -4571 5083 -4519
rect 5135 -4558 5249 -4519
rect 5301 -4558 5403 -4506
rect 5135 -4571 5403 -4558
rect -8942 -4639 5403 -4571
rect 5033 -4646 5403 -4639
rect 5033 -4657 5254 -4646
rect 5033 -4709 5083 -4657
rect 5135 -4698 5254 -4657
rect 5306 -4698 5403 -4646
rect 5135 -4709 5403 -4698
rect 5033 -4740 5403 -4709
rect 18482 -5517 18859 -3258
rect 20039 -3510 20131 -3484
rect 21848 -3510 22220 -2548
rect 20039 -3680 22220 -3510
rect 87273 -4550 87648 -1197
rect 98576 -1966 98937 -1953
rect 98576 -2018 98635 -1966
rect 98687 -1967 98937 -1966
rect 98687 -2018 98809 -1967
rect 98576 -2019 98809 -2018
rect 98861 -2019 98937 -1967
rect 98576 -2020 98937 -2019
rect 98576 -2132 99239 -2020
rect 98576 -2184 98636 -2132
rect 98688 -2135 99239 -2132
rect 98688 -2137 98937 -2135
rect 98688 -2184 98834 -2137
rect 98576 -2189 98834 -2184
rect 98886 -2189 98937 -2137
rect 98576 -2221 98937 -2189
rect 98546 -2863 98907 -2850
rect 98546 -2915 98605 -2863
rect 98657 -2864 98907 -2863
rect 98657 -2915 98779 -2864
rect 98546 -2916 98779 -2915
rect 98831 -2916 98907 -2864
rect 98546 -2917 98907 -2916
rect 98546 -3029 99209 -2917
rect 98546 -3081 98606 -3029
rect 98658 -3032 99209 -3029
rect 98658 -3034 98907 -3032
rect 98658 -3081 98804 -3034
rect 98546 -3086 98804 -3081
rect 98856 -3086 98907 -3034
rect 98546 -3118 98907 -3086
rect 98538 -3346 98899 -3333
rect 98538 -3398 98597 -3346
rect 98649 -3347 98899 -3346
rect 98649 -3398 98771 -3347
rect 98538 -3399 98771 -3398
rect 98823 -3399 98899 -3347
rect 98538 -3400 98899 -3399
rect 98538 -3512 99201 -3400
rect 98538 -3564 98598 -3512
rect 98650 -3515 99201 -3512
rect 98650 -3517 98899 -3515
rect 98650 -3564 98796 -3517
rect 98538 -3569 98796 -3564
rect 98848 -3569 98899 -3517
rect 98538 -3601 98899 -3569
rect 98576 -3898 98937 -3885
rect 98576 -3950 98635 -3898
rect 98687 -3899 98937 -3898
rect 98687 -3950 98809 -3899
rect 98576 -3951 98809 -3950
rect 98861 -3951 98937 -3899
rect 98576 -3952 98937 -3951
rect 98576 -4064 99239 -3952
rect 98576 -4116 98636 -4064
rect 98688 -4067 99239 -4064
rect 98688 -4069 98937 -4067
rect 98688 -4116 98834 -4069
rect 98576 -4121 98834 -4116
rect 98886 -4121 98937 -4069
rect 98576 -4153 98937 -4121
rect 87090 -4724 87760 -4550
rect 87090 -4776 87136 -4724
rect 87188 -4776 87256 -4724
rect 87308 -4776 87376 -4724
rect 87428 -4776 87760 -4724
rect 87090 -4844 87760 -4776
rect 87090 -4896 87136 -4844
rect 87188 -4896 87256 -4844
rect 87308 -4896 87376 -4844
rect 87428 -4896 87760 -4844
rect 87090 -4964 87760 -4896
rect 87090 -5016 87136 -4964
rect 87188 -5016 87256 -4964
rect 87308 -5016 87376 -4964
rect 87428 -5016 87760 -4964
rect 87090 -5090 87760 -5016
rect 35448 -7135 35605 -7054
rect 46331 -7299 48908 -7093
rect 6386 -8123 6433 -7467
rect 13089 -7874 13136 -7507
rect 28743 -7995 28833 -7665
rect 57536 -8443 57583 -7347
rect 64239 -8183 64286 -7477
rect 79893 -8205 79983 -7375
rect 98574 -7474 98910 -7460
rect 98574 -7526 98606 -7474
rect 98658 -7526 98726 -7474
rect 98778 -7526 98846 -7474
rect 98898 -7526 98910 -7474
rect 98574 -7530 98910 -7526
rect 98574 -7594 99250 -7530
rect 98574 -7646 98606 -7594
rect 98658 -7646 98726 -7594
rect 98778 -7646 98846 -7594
rect 98898 -7646 99250 -7594
rect 98574 -7690 99250 -7646
rect 98574 -7714 98910 -7690
rect 98574 -7766 98606 -7714
rect 98658 -7766 98726 -7714
rect 98778 -7766 98846 -7714
rect 98898 -7766 98910 -7714
rect 98574 -7800 98910 -7766
rect 54726 -8904 56321 -8804
rect 34288 -8979 34546 -8905
rect 37498 -8979 37754 -8906
rect 48724 -9293 48793 -9131
rect 48405 -9341 48793 -9293
rect 48405 -9393 48446 -9341
rect 48498 -9353 48793 -9341
rect 48498 -9393 48585 -9353
rect 48405 -9405 48585 -9393
rect 48637 -9405 48793 -9353
rect 48405 -9457 48793 -9405
rect 48405 -9509 48440 -9457
rect 48492 -9478 48793 -9457
rect 48492 -9509 48588 -9478
rect 48405 -9530 48588 -9509
rect 48640 -9530 48793 -9478
rect 48405 -9571 48793 -9530
rect 48405 -9623 48443 -9571
rect 48495 -9594 48793 -9571
rect 48495 -9623 48588 -9594
rect 48405 -9646 48588 -9623
rect 48640 -9646 48793 -9594
rect 48405 -9663 48793 -9646
rect 13833 -10333 13879 -9997
rect 48724 -10104 48793 -9663
rect 52279 -11322 53565 -11166
rect 52279 -11368 53571 -11322
rect 52279 -11371 53319 -11368
rect 52279 -11379 53077 -11371
rect 52279 -11381 52808 -11379
rect 52279 -11394 52553 -11381
rect 52279 -11446 52348 -11394
rect 52400 -11433 52553 -11394
rect 52605 -11431 52808 -11381
rect 52860 -11423 53077 -11379
rect 53129 -11420 53319 -11371
rect 53371 -11420 53571 -11368
rect 53129 -11423 53571 -11420
rect 52860 -11431 53571 -11423
rect 52605 -11433 53571 -11431
rect 52400 -11446 53571 -11433
rect 52279 -11550 53571 -11446
rect 52279 -11551 53406 -11550
rect 52279 -11563 53247 -11551
rect 52279 -11566 53034 -11563
rect 52279 -11576 52789 -11566
rect 52279 -11584 52556 -11576
rect 52279 -11636 52350 -11584
rect 52402 -11628 52556 -11584
rect 52608 -11618 52789 -11576
rect 52841 -11615 53034 -11566
rect 53086 -11603 53247 -11563
rect 53299 -11602 53406 -11551
rect 53458 -11602 53571 -11550
rect 53299 -11603 53571 -11602
rect 53086 -11615 53571 -11603
rect 52841 -11618 53571 -11615
rect 52608 -11628 53571 -11618
rect 52402 -11636 53571 -11628
rect 13098 -12624 13146 -12186
rect 28843 -12493 28889 -11707
rect 52279 -11736 53571 -11636
rect 52279 -11744 53355 -11736
rect 52279 -11754 53157 -11744
rect 52279 -11757 52918 -11754
rect 52279 -11759 52707 -11757
rect 52279 -11760 52509 -11759
rect 52279 -11812 52341 -11760
rect 52393 -11811 52509 -11760
rect 52561 -11809 52707 -11759
rect 52759 -11806 52918 -11757
rect 52970 -11796 53157 -11754
rect 53209 -11788 53355 -11744
rect 53407 -11788 53571 -11736
rect 53209 -11796 53571 -11788
rect 52970 -11806 53571 -11796
rect 52759 -11809 53571 -11806
rect 52561 -11811 53571 -11809
rect 52393 -11812 53571 -11811
rect 52279 -11848 53571 -11812
rect 56118 -13869 56321 -8904
rect 64983 -10117 65030 -10037
rect 64983 -10164 65333 -10117
rect 64983 -10343 65030 -10164
rect 64248 -12534 64296 -11606
rect 79993 -12443 80039 -11737
rect 48789 -14156 56323 -13869
rect 48789 -14208 49199 -14156
rect 49251 -14208 49319 -14156
rect 49371 -14208 49439 -14156
rect 49491 -14208 56323 -14156
rect 48789 -14276 56323 -14208
rect 48789 -14328 49199 -14276
rect 49251 -14328 49319 -14276
rect 49371 -14328 49439 -14276
rect 49491 -14328 56323 -14276
rect 48789 -14514 56323 -14328
rect 25725 -14613 27275 -14562
rect 14185 -16057 14240 -15620
rect 27991 -15636 28043 -14884
rect 19853 -16443 19978 -16366
rect 28905 -18073 28951 -17807
rect 42594 -18574 45406 -18222
rect 52080 -31258 52856 -14514
rect 77165 -14593 77995 -14542
rect 65335 -15997 65390 -15493
rect 65336 -16516 65388 -15997
rect 79141 -16316 79193 -14894
rect 79617 -17833 80103 -17787
rect 80055 -18003 80101 -17833
rect 93784 -18554 96726 -18202
rect -25406 -32034 52856 -31258
<< via1 >>
rect -2669 52674 -2617 52726
rect -2505 52672 -2453 52724
rect -2669 52547 -2617 52599
rect -2503 52560 -2451 52612
rect -2669 52409 -2617 52461
rect -2498 52420 -2446 52472
rect -2359 44148 -2307 44200
rect -2195 44146 -2143 44198
rect -2359 44021 -2307 44073
rect -2193 44034 -2141 44086
rect -2359 43883 -2307 43935
rect -2188 43894 -2136 43946
rect -2352 43607 -2300 43659
rect -2188 43605 -2136 43657
rect -2352 43480 -2300 43532
rect -2186 43493 -2134 43545
rect -2352 43342 -2300 43394
rect -2181 43353 -2129 43405
rect -2460 36714 -2408 36766
rect -2296 36712 -2244 36764
rect -2460 36587 -2408 36639
rect -2294 36600 -2242 36652
rect -2460 36449 -2408 36501
rect -2289 36460 -2237 36512
rect 2043 27965 2095 28017
rect 2222 27962 2274 28014
rect 2419 27965 2471 28017
rect 2609 27973 2661 28025
rect 2046 27838 2098 27890
rect 2222 27827 2274 27879
rect 2411 27830 2463 27882
rect 2609 27838 2661 27890
rect -3571 24988 -3519 25040
rect -3451 24988 -3399 25040
rect -3331 24988 -3279 25040
rect -3571 24868 -3519 24920
rect -3451 24868 -3399 24920
rect -3331 24868 -3279 24920
rect -3571 24748 -3519 24800
rect -3451 24748 -3399 24800
rect -3331 24748 -3279 24800
rect 14140 19472 14192 19524
rect 14311 19472 14363 19524
rect 14482 19472 14534 19524
rect 14653 19472 14705 19524
rect 14824 19472 14876 19524
rect 14995 19472 15047 19524
rect 15166 19472 15218 19524
rect 15337 19472 15389 19524
rect 15508 19472 15560 19524
rect 15679 19472 15731 19524
rect 15850 19472 15902 19524
rect 16021 19472 16073 19524
rect 16192 19472 16244 19524
rect 16363 19472 16415 19524
rect 16534 19472 16586 19524
rect 14140 19307 14192 19359
rect 14311 19307 14363 19359
rect 14482 19307 14534 19359
rect 14653 19307 14705 19359
rect 14824 19307 14876 19359
rect 14995 19307 15047 19359
rect 15166 19307 15218 19359
rect 15337 19307 15389 19359
rect 15508 19307 15560 19359
rect 15679 19307 15731 19359
rect 15850 19307 15902 19359
rect 16021 19307 16073 19359
rect 16192 19307 16244 19359
rect 16363 19307 16415 19359
rect 16534 19307 16586 19359
rect 14140 19142 14192 19194
rect 14311 19142 14363 19194
rect 14482 19142 14534 19194
rect 14653 19142 14705 19194
rect 14824 19142 14876 19194
rect 14995 19142 15047 19194
rect 15166 19142 15218 19194
rect 15337 19142 15389 19194
rect 15508 19142 15560 19194
rect 15679 19142 15731 19194
rect 15850 19142 15902 19194
rect 16021 19142 16073 19194
rect 16192 19142 16244 19194
rect 16363 19142 16415 19194
rect 16534 19142 16586 19194
rect -13882 18756 -13830 18808
rect -13758 18756 -13706 18808
rect -13634 18756 -13582 18808
rect -13510 18756 -13458 18808
rect -13882 18632 -13830 18684
rect -13758 18632 -13706 18684
rect -13634 18632 -13582 18684
rect -13510 18632 -13458 18684
rect -13882 18508 -13830 18560
rect -13758 18508 -13706 18560
rect -13634 18508 -13582 18560
rect -13510 18508 -13458 18560
rect -13882 18384 -13830 18436
rect -13758 18384 -13706 18436
rect -13634 18384 -13582 18436
rect -13510 18384 -13458 18436
rect -13966 17670 -13914 17722
rect -13842 17670 -13790 17722
rect -13718 17670 -13666 17722
rect -13594 17670 -13542 17722
rect -12463 17662 -12411 17714
rect -12339 17662 -12287 17714
rect -12215 17662 -12163 17714
rect -12091 17662 -12039 17714
rect -13966 17546 -13914 17598
rect -13842 17546 -13790 17598
rect -13718 17546 -13666 17598
rect -13594 17546 -13542 17598
rect -12463 17538 -12411 17590
rect -12339 17538 -12287 17590
rect -12215 17538 -12163 17590
rect -12091 17538 -12039 17590
rect -13966 17422 -13914 17474
rect -13842 17422 -13790 17474
rect -13718 17422 -13666 17474
rect -13594 17422 -13542 17474
rect -12463 17414 -12411 17466
rect -12339 17414 -12287 17466
rect -12215 17414 -12163 17466
rect -12091 17414 -12039 17466
rect -13966 17298 -13914 17350
rect -13842 17298 -13790 17350
rect -13718 17298 -13666 17350
rect -13594 17298 -13542 17350
rect -12463 17290 -12411 17342
rect -12339 17290 -12287 17342
rect -12215 17290 -12163 17342
rect -12091 17290 -12039 17342
rect 9836 17544 9888 17596
rect 9964 17544 10016 17596
rect 10115 17541 10167 17593
rect 9834 17385 9886 17437
rect 10005 17383 10057 17435
rect 10181 17385 10233 17437
rect 9846 17201 9898 17253
rect 10048 17206 10100 17258
rect 10197 17222 10249 17274
rect 9795 16871 9847 16923
rect 9923 16874 9975 16926
rect 10054 16881 10106 16933
rect 9790 16674 9842 16726
rect 9959 16692 10011 16744
rect 10107 16697 10159 16749
rect 9767 16523 9819 16575
rect 9964 16554 10016 16606
rect 10141 16564 10193 16616
rect 4007 14689 4059 14741
rect 4134 14689 4186 14741
rect -15546 13200 -15494 13252
rect -15422 13200 -15370 13252
rect -15298 13200 -15246 13252
rect -15174 13200 -15122 13252
rect -14237 13221 -14185 13273
rect -14113 13221 -14061 13273
rect -13989 13221 -13937 13273
rect -13865 13221 -13813 13273
rect -15546 13076 -15494 13128
rect -15422 13076 -15370 13128
rect -15298 13076 -15246 13128
rect -15174 13076 -15122 13128
rect -14237 13097 -14185 13149
rect -14113 13097 -14061 13149
rect -13989 13097 -13937 13149
rect -13865 13097 -13813 13149
rect -15546 12952 -15494 13004
rect -15422 12952 -15370 13004
rect -15298 12952 -15246 13004
rect -15174 12952 -15122 13004
rect -14237 12973 -14185 13025
rect -14113 12973 -14061 13025
rect -13989 12973 -13937 13025
rect -13865 12973 -13813 13025
rect -15546 12828 -15494 12880
rect -15422 12828 -15370 12880
rect -15298 12828 -15246 12880
rect -15174 12828 -15122 12880
rect -14237 12849 -14185 12901
rect -14113 12849 -14061 12901
rect -13989 12849 -13937 12901
rect -13865 12849 -13813 12901
rect 10858 13398 10910 13450
rect 10996 13398 11048 13450
rect 10861 13271 10913 13323
rect 11000 13269 11052 13321
rect 10860 13118 10912 13170
rect 11000 13127 11052 13179
rect 11046 12810 11098 12862
rect 11184 12810 11236 12862
rect 11173 12678 11225 12730
rect 12271 12363 12323 12415
rect 12409 12363 12461 12415
rect 12274 12236 12326 12288
rect 12413 12234 12465 12286
rect 12273 12083 12325 12135
rect 12413 12092 12465 12144
rect 8609 11609 8661 11661
rect 8731 11610 8783 11662
rect 8876 11613 8928 11665
rect 8615 11497 8667 11549
rect 8746 11498 8798 11550
rect 8885 11498 8937 11550
rect -9354 9579 -9302 9631
rect -8805 9579 -8753 9631
rect -9334 8863 -9282 8915
rect -8785 8863 -8733 8915
rect 11344 9927 11396 9979
rect 11521 9938 11573 9990
rect 11278 9796 11330 9848
rect 11414 9806 11466 9858
rect 11561 9801 11613 9853
rect 2389 8912 2441 8964
rect 2711 8912 2763 8964
rect 11440 7930 11492 7982
rect 11574 7930 11626 7982
rect 11435 7816 11487 7868
rect 11564 7804 11616 7856
rect 137 7179 189 7231
rect 644 7200 696 7252
rect 1047 7203 1099 7255
rect 12966 7253 13018 7305
rect 13102 7253 13154 7305
rect 12961 7140 13013 7192
rect 95 6871 147 6923
rect 511 6909 563 6961
rect 910 6916 962 6968
rect 13097 7133 13149 7185
rect 8598 7016 8650 7068
rect 8741 7016 8793 7068
rect 8953 7021 9005 7073
rect 8598 6904 8650 6956
rect 8746 6904 8798 6956
rect 8984 6904 9036 6956
rect -7 6552 45 6604
rect 266 6556 318 6608
rect 644 6580 696 6632
rect 998 6594 1050 6646
rect 620 6135 672 6187
rect 12502 5340 12554 5392
rect 12679 5351 12731 5403
rect 12436 5209 12488 5261
rect 12572 5219 12624 5271
rect 12719 5214 12771 5266
rect 4706 3732 4758 3784
rect 5213 3753 5265 3805
rect 5616 3756 5668 3808
rect 4664 3424 4716 3476
rect 5080 3462 5132 3514
rect 5479 3469 5531 3521
rect 4562 3105 4614 3157
rect 4835 3109 4887 3161
rect 5213 3133 5265 3185
rect 5567 3147 5619 3199
rect 17931 14008 18191 14268
rect 17919 13787 18179 13943
rect 19181 14115 19233 14167
rect 19412 14115 19464 14167
rect 19179 13901 19231 13953
rect 19401 13901 19453 13953
rect 20393 13831 20653 14091
rect 19178 13671 19230 13723
rect 19389 13679 19441 13731
rect 22822 16379 22874 16431
rect 22942 16379 22994 16431
rect 23062 16379 23114 16431
rect 23182 16379 23234 16431
rect 23302 16379 23354 16431
rect 22822 16259 22874 16311
rect 22942 16259 22994 16311
rect 23062 16259 23114 16311
rect 23182 16259 23234 16311
rect 23302 16259 23354 16311
rect 22094 15198 22146 15250
rect 22214 15198 22266 15250
rect 22334 15198 22386 15250
rect 22454 15198 22506 15250
rect 22574 15198 22626 15250
rect 22094 15078 22146 15130
rect 22214 15078 22266 15130
rect 22334 15078 22386 15130
rect 22454 15078 22506 15130
rect 22574 15078 22626 15130
rect 22063 14580 22115 14632
rect 22183 14580 22235 14632
rect 22303 14580 22355 14632
rect 22423 14580 22475 14632
rect 22543 14580 22595 14632
rect 22063 14460 22115 14512
rect 22183 14460 22235 14512
rect 22303 14460 22355 14512
rect 22423 14460 22475 14512
rect 22543 14460 22595 14512
rect 95813 18400 95865 18452
rect 95933 18400 95985 18452
rect 96053 18400 96105 18452
rect 95813 18280 95865 18332
rect 95933 18280 95985 18332
rect 96053 18280 96105 18332
rect 95813 18160 95865 18212
rect 95933 18160 95985 18212
rect 96053 18160 96105 18212
rect 26428 16774 26480 16826
rect 26548 16774 26600 16826
rect 26668 16774 26720 16826
rect 26788 16774 26840 16826
rect 26908 16774 26960 16826
rect 26428 16654 26480 16706
rect 26548 16654 26600 16706
rect 26668 16654 26720 16706
rect 26788 16654 26840 16706
rect 26908 16654 26960 16706
rect 95925 16774 95977 16826
rect 96045 16774 96097 16826
rect 96165 16774 96217 16826
rect 95925 16654 95977 16706
rect 96045 16654 96097 16706
rect 96165 16654 96217 16706
rect 95925 16534 95977 16586
rect 96045 16534 96097 16586
rect 96165 16534 96217 16586
rect 22116 13928 22272 14084
rect 22498 13928 22654 14084
rect 22917 13928 23073 14084
rect 37935 14106 37987 14158
rect 38055 14106 38107 14158
rect 38175 14106 38227 14158
rect 38295 14106 38347 14158
rect 38415 14106 38467 14158
rect 37935 13986 37987 14038
rect 38055 13986 38107 14038
rect 38175 13986 38227 14038
rect 38295 13986 38347 14038
rect 38415 13986 38467 14038
rect 22006 13564 22058 13616
rect 22429 13564 22481 13616
rect 22720 13564 22772 13616
rect 21838 13187 21890 13239
rect 22077 13187 22129 13239
rect 22410 13187 22462 13239
rect 29830 13273 29882 13325
rect 29950 13273 30002 13325
rect 30070 13273 30122 13325
rect 30190 13273 30242 13325
rect 30310 13273 30362 13325
rect 29830 13153 29882 13205
rect 29950 13153 30002 13205
rect 30070 13153 30122 13205
rect 30190 13153 30242 13205
rect 30310 13153 30362 13205
rect 19670 11136 19722 11188
rect 19911 11141 19963 11193
rect 20150 11143 20202 11195
rect 20377 11143 20429 11195
rect 22481 11115 22533 11167
rect 22476 10971 22528 11023
rect 64929 13720 64981 13772
rect 65188 13716 65240 13768
rect 65429 13651 65481 13703
rect 64933 13569 64985 13621
rect 65200 13539 65252 13591
rect 65424 13498 65476 13550
rect 64932 13400 64984 13452
rect 65190 13402 65242 13454
rect 65422 13355 65474 13407
rect 64982 13225 65034 13277
rect 65184 13220 65236 13272
rect 65347 13208 65399 13260
rect 41755 12582 41807 12634
rect 41755 12332 41807 12384
rect 41755 12108 41807 12160
rect 37877 10732 37929 10784
rect 37997 10732 38049 10784
rect 38117 10732 38169 10784
rect 38237 10732 38289 10784
rect 38357 10732 38409 10784
rect 37877 10612 37929 10664
rect 37997 10612 38049 10664
rect 38117 10612 38169 10664
rect 38237 10612 38289 10664
rect 38357 10612 38409 10664
rect 28784 9841 28836 9893
rect 29025 9846 29077 9898
rect 29264 9848 29316 9900
rect 29491 9848 29543 9900
rect 19628 9090 19680 9142
rect 19869 9095 19921 9147
rect 20108 9097 20160 9149
rect 20335 9097 20387 9149
rect 22939 7822 22991 7874
rect 23180 7827 23232 7879
rect 23419 7829 23471 7881
rect 23646 7829 23698 7881
rect 28728 6847 28780 6899
rect 28969 6852 29021 6904
rect 29208 6854 29260 6906
rect 29435 6854 29487 6906
rect 22134 6737 22186 6789
rect 22430 6737 22482 6789
rect 18072 6618 18124 6670
rect 18192 6618 18244 6670
rect 18312 6618 18364 6670
rect 18432 6618 18484 6670
rect 18552 6618 18604 6670
rect 18672 6618 18724 6670
rect 18792 6618 18844 6670
rect 18912 6618 18964 6670
rect 19032 6618 19084 6670
rect 19152 6618 19204 6670
rect 19272 6618 19324 6670
rect 19392 6618 19444 6670
rect 18232 5959 18284 6011
rect 18410 5957 18462 6009
rect 18651 5956 18703 6008
rect 18892 5962 18944 6014
rect 32075 9827 32127 9879
rect 47793 8176 47845 8228
rect 47949 8176 48001 8228
rect 54014 9262 54066 9314
rect 54133 9262 54185 9314
rect 54252 9263 54304 9315
rect 54374 9264 54426 9316
rect 54492 9263 54544 9315
rect 54014 9144 54066 9196
rect 54133 9144 54185 9196
rect 54254 9145 54306 9197
rect 54374 9147 54426 9199
rect 54493 9143 54545 9195
rect 61584 9269 61636 9321
rect 61703 9269 61755 9321
rect 61822 9270 61874 9322
rect 61944 9271 61996 9323
rect 62062 9270 62114 9322
rect 61584 9151 61636 9203
rect 61703 9151 61755 9203
rect 61824 9152 61876 9204
rect 61944 9154 61996 9206
rect 62063 9150 62115 9202
rect 43285 6948 43441 7104
rect 43828 6948 43984 7104
rect 44538 6948 44694 7104
rect 46195 7021 46247 7073
rect 46441 7016 46493 7068
rect 46721 7018 46773 7070
rect 46937 7026 46989 7078
rect 39342 6452 39498 6608
rect 43825 6022 43877 6074
rect 44074 6009 44126 6061
rect 44308 6004 44360 6056
rect 44530 6008 44582 6060
rect 27149 4353 27201 4405
rect 27381 4353 27433 4405
rect 30470 4435 30522 4487
rect 27146 4157 27198 4209
rect 27381 4157 27433 4209
rect 30470 4174 30522 4226
rect 56834 6745 56886 6797
rect 57017 6751 57069 6803
rect 57204 6751 57256 6803
rect 53788 4608 53840 4660
rect 53907 4608 53959 4660
rect 54026 4609 54078 4661
rect 54148 4610 54200 4662
rect 54266 4609 54318 4661
rect 53788 4490 53840 4542
rect 53907 4490 53959 4542
rect 54028 4491 54080 4543
rect 54148 4493 54200 4545
rect 54267 4489 54319 4541
rect -3695 1098 -3435 1358
rect -3106 1112 -2846 1372
rect 56911 2049 56963 2101
rect 57094 2055 57146 2107
rect 57281 2055 57333 2107
rect -2317 25 -2057 285
rect -1728 39 -1468 299
rect 2727 -311 2779 -259
rect 2891 -313 2943 -261
rect 2727 -438 2779 -386
rect 2893 -425 2945 -373
rect 2727 -576 2779 -524
rect 2898 -565 2950 -513
rect 60715 -297 60767 -245
rect 60991 -273 61043 -221
rect 60677 -535 60729 -483
rect 60900 -536 60952 -484
rect 61143 -532 61195 -480
rect 4828 -1042 4880 -990
rect 4992 -1044 5044 -992
rect 4828 -1169 4880 -1117
rect 4994 -1156 5046 -1104
rect 4828 -1307 4880 -1255
rect 4999 -1296 5051 -1244
rect 4894 -1621 4946 -1569
rect 5060 -1608 5112 -1556
rect 18145 -1598 18197 -1546
rect 18452 -1593 18504 -1541
rect 18702 -1586 18754 -1534
rect 4894 -1759 4946 -1707
rect 5065 -1748 5117 -1696
rect 95787 15586 95839 15638
rect 95907 15586 95959 15638
rect 96027 15586 96079 15638
rect 95787 15466 95839 15518
rect 95907 15466 95959 15518
rect 96027 15466 96079 15518
rect 95787 15346 95839 15398
rect 95907 15346 95959 15398
rect 96027 15346 96079 15398
rect 95801 14552 95853 14604
rect 95921 14552 95973 14604
rect 96041 14552 96093 14604
rect 95801 14432 95853 14484
rect 95921 14432 95973 14484
rect 96041 14432 96093 14484
rect 95801 14312 95853 14364
rect 95921 14312 95973 14364
rect 96041 14312 96093 14364
rect 98889 4667 98941 4719
rect 99064 4661 99116 4713
rect 98887 4508 98939 4560
rect 99065 4512 99117 4564
rect 98890 4343 98942 4395
rect 99078 4338 99130 4390
rect 91420 4201 91472 4253
rect 91539 4201 91591 4253
rect 91658 4202 91710 4254
rect 91780 4203 91832 4255
rect 91898 4202 91950 4254
rect 91420 4083 91472 4135
rect 91539 4083 91591 4135
rect 91660 4084 91712 4136
rect 91780 4086 91832 4138
rect 91899 4082 91951 4134
rect 95236 2614 95288 2666
rect 95356 2614 95408 2666
rect 95476 2614 95528 2666
rect 95236 2494 95288 2546
rect 95356 2494 95408 2546
rect 95476 2494 95528 2546
rect 95236 2374 95288 2426
rect 95356 2374 95408 2426
rect 95476 2374 95528 2426
rect 89881 -330 89933 -278
rect 90095 -323 90147 -271
rect 89878 -524 89930 -472
rect 90086 -524 90138 -472
rect 4796 -2305 4848 -2253
rect 4547 -2408 4599 -2356
rect 4687 -2408 4739 -2356
rect 4549 -2529 4601 -2477
rect 4695 -2532 4747 -2480
rect 4815 -2537 4867 -2485
rect 5051 -2717 5103 -2665
rect 5217 -2704 5269 -2652
rect 5051 -2855 5103 -2803
rect 5222 -2844 5274 -2792
rect 4955 -3135 5007 -3083
rect 5121 -3122 5173 -3070
rect 4955 -3273 5007 -3221
rect 5126 -3262 5178 -3210
rect 4932 -3549 4984 -3497
rect 5098 -3536 5150 -3484
rect 4932 -3687 4984 -3635
rect 5103 -3676 5155 -3624
rect 4978 -4028 5030 -3976
rect 5144 -4015 5196 -3963
rect 4978 -4166 5030 -4114
rect 5149 -4155 5201 -4103
rect 5083 -4571 5135 -4519
rect 5249 -4558 5301 -4506
rect 5083 -4709 5135 -4657
rect 5254 -4698 5306 -4646
rect 98635 -2018 98687 -1966
rect 98809 -2019 98861 -1967
rect 98636 -2184 98688 -2132
rect 98834 -2189 98886 -2137
rect 98605 -2915 98657 -2863
rect 98779 -2916 98831 -2864
rect 98606 -3081 98658 -3029
rect 98804 -3086 98856 -3034
rect 98597 -3398 98649 -3346
rect 98771 -3399 98823 -3347
rect 98598 -3564 98650 -3512
rect 98796 -3569 98848 -3517
rect 98635 -3950 98687 -3898
rect 98809 -3951 98861 -3899
rect 98636 -4116 98688 -4064
rect 98834 -4121 98886 -4069
rect 87136 -4776 87188 -4724
rect 87256 -4776 87308 -4724
rect 87376 -4776 87428 -4724
rect 87136 -4896 87188 -4844
rect 87256 -4896 87308 -4844
rect 87376 -4896 87428 -4844
rect 87136 -5016 87188 -4964
rect 87256 -5016 87308 -4964
rect 87376 -5016 87428 -4964
rect 98606 -7526 98658 -7474
rect 98726 -7526 98778 -7474
rect 98846 -7526 98898 -7474
rect 98606 -7646 98658 -7594
rect 98726 -7646 98778 -7594
rect 98846 -7646 98898 -7594
rect 98606 -7766 98658 -7714
rect 98726 -7766 98778 -7714
rect 98846 -7766 98898 -7714
rect 48446 -9393 48498 -9341
rect 48585 -9405 48637 -9353
rect 48440 -9509 48492 -9457
rect 48588 -9530 48640 -9478
rect 48443 -9623 48495 -9571
rect 48588 -9646 48640 -9594
rect 52348 -11446 52400 -11394
rect 52553 -11433 52605 -11381
rect 52808 -11431 52860 -11379
rect 53077 -11423 53129 -11371
rect 53319 -11420 53371 -11368
rect 52350 -11636 52402 -11584
rect 52556 -11628 52608 -11576
rect 52789 -11618 52841 -11566
rect 53034 -11615 53086 -11563
rect 53247 -11603 53299 -11551
rect 53406 -11602 53458 -11550
rect 52341 -11812 52393 -11760
rect 52509 -11811 52561 -11759
rect 52707 -11809 52759 -11757
rect 52918 -11806 52970 -11754
rect 53157 -11796 53209 -11744
rect 53355 -11788 53407 -11736
rect 49199 -14208 49251 -14156
rect 49319 -14208 49371 -14156
rect 49439 -14208 49491 -14156
rect 49199 -14328 49251 -14276
rect 49319 -14328 49371 -14276
rect 49439 -14328 49491 -14276
<< metal2 >>
rect -2698 52728 -2423 52744
rect -2698 52672 -2671 52728
rect -2615 52726 -2423 52728
rect -2615 52672 -2507 52726
rect -2698 52670 -2507 52672
rect -2451 52670 -2423 52726
rect -2698 52614 -2423 52670
rect -2698 52601 -2505 52614
rect -2698 52545 -2671 52601
rect -2615 52558 -2505 52601
rect -2449 52558 -2423 52614
rect -2615 52545 -2423 52558
rect -2698 52474 -2423 52545
rect -2698 52463 -2500 52474
rect -2698 52407 -2671 52463
rect -2615 52418 -2500 52463
rect -2444 52418 -2423 52474
rect -2615 52407 -2423 52418
rect -2698 52394 -2423 52407
rect -2388 44202 -2113 44218
rect -2388 44146 -2361 44202
rect -2305 44200 -2113 44202
rect -2305 44146 -2197 44200
rect -2388 44144 -2197 44146
rect -2141 44144 -2113 44200
rect -2388 44088 -2113 44144
rect -2388 44075 -2195 44088
rect -2388 44019 -2361 44075
rect -2305 44032 -2195 44075
rect -2139 44032 -2113 44088
rect -2305 44019 -2113 44032
rect -2388 43948 -2113 44019
rect -2388 43937 -2190 43948
rect -2388 43881 -2361 43937
rect -2305 43892 -2190 43937
rect -2134 43892 -2113 43948
rect -2305 43881 -2113 43892
rect -2388 43868 -2113 43881
rect -2381 43661 -2106 43677
rect -2381 43605 -2354 43661
rect -2298 43659 -2106 43661
rect -2298 43605 -2190 43659
rect -2381 43603 -2190 43605
rect -2134 43603 -2106 43659
rect -2381 43547 -2106 43603
rect -2381 43534 -2188 43547
rect -2381 43478 -2354 43534
rect -2298 43491 -2188 43534
rect -2132 43491 -2106 43547
rect -2298 43478 -2106 43491
rect -2381 43407 -2106 43478
rect -2381 43396 -2183 43407
rect -2381 43340 -2354 43396
rect -2298 43351 -2183 43396
rect -2127 43351 -2106 43407
rect -2298 43340 -2106 43351
rect -2381 43327 -2106 43340
rect -2489 36768 -2214 36784
rect -2489 36712 -2462 36768
rect -2406 36766 -2214 36768
rect -2406 36712 -2298 36766
rect -2489 36710 -2298 36712
rect -2242 36710 -2214 36766
rect -2489 36654 -2214 36710
rect -2489 36641 -2296 36654
rect -2489 36585 -2462 36641
rect -2406 36598 -2296 36641
rect -2240 36598 -2214 36654
rect -2406 36585 -2214 36598
rect -2489 36514 -2214 36585
rect -2489 36503 -2291 36514
rect -2489 36447 -2462 36503
rect -2406 36458 -2291 36503
rect -2235 36458 -2214 36514
rect -2406 36447 -2214 36458
rect -2489 36434 -2214 36447
rect 2010 28027 2740 28118
rect 2010 28019 2607 28027
rect 2010 27963 2041 28019
rect 2097 28016 2417 28019
rect 2097 27963 2220 28016
rect 2010 27960 2220 27963
rect 2276 27963 2417 28016
rect 2473 27971 2607 28019
rect 2663 27971 2740 28027
rect 2473 27963 2740 27971
rect 2276 27960 2740 27963
rect 2010 27892 2740 27960
rect 2010 27836 2044 27892
rect 2100 27884 2607 27892
rect 2100 27881 2409 27884
rect 2100 27836 2220 27881
rect 2010 27825 2220 27836
rect 2276 27828 2409 27881
rect 2465 27836 2607 27884
rect 2663 27836 2740 27892
rect 2465 27828 2740 27836
rect 2276 27825 2740 27828
rect 2010 27720 2740 27825
rect -3588 25044 -3261 25051
rect -3592 25043 -3165 25044
rect -3592 25040 -1026 25043
rect -3592 24988 -3571 25040
rect -3519 24988 -3451 25040
rect -3399 24988 -3331 25040
rect -3279 24988 -1026 25040
rect -3592 24951 -1026 24988
rect -3592 24920 -464 24951
rect -3592 24868 -3571 24920
rect -3519 24868 -3451 24920
rect -3399 24868 -3331 24920
rect -3279 24868 -464 24920
rect -3592 24840 -464 24868
rect -3592 24800 -1026 24840
rect -3592 24748 -3571 24800
rect -3519 24748 -3451 24800
rect -3399 24748 -3331 24800
rect -3279 24748 -1026 24800
rect -3592 24732 -3165 24748
rect -1775 20749 -1405 23311
rect 8582 21777 9071 21859
rect 8582 21757 8980 21777
rect 8582 21701 8765 21757
rect 8821 21721 8980 21757
rect 9036 21721 9071 21777
rect 8821 21701 9071 21721
rect 8582 21604 9071 21701
rect 8582 21594 8916 21604
rect 8582 21538 8654 21594
rect 8710 21548 8916 21594
rect 8972 21548 9071 21604
rect 8710 21538 9071 21548
rect 8582 21353 9071 21538
rect 8582 21343 8892 21353
rect 8582 21287 8672 21343
rect 8728 21297 8892 21343
rect 8948 21297 9071 21353
rect 8728 21287 9071 21297
rect 8582 21236 9071 21287
rect -265 20749 1066 20974
rect -1794 20711 1066 20749
rect -1794 20691 377 20711
rect -1794 20635 162 20691
rect 218 20655 377 20691
rect 433 20655 1066 20711
rect 218 20635 1066 20655
rect -1794 20538 1066 20635
rect -1794 20528 313 20538
rect -1794 20472 51 20528
rect 107 20482 313 20528
rect 369 20482 1066 20538
rect 107 20472 1066 20482
rect -1794 20340 1066 20472
rect -265 20287 1066 20340
rect -265 20277 289 20287
rect -265 20221 69 20277
rect 125 20231 289 20277
rect 345 20231 1066 20287
rect 125 20221 1066 20231
rect -265 19888 1066 20221
rect -15247 18862 -10439 19168
rect -15247 18808 -12465 18862
rect -15247 18756 -13882 18808
rect -13830 18756 -13758 18808
rect -13706 18756 -13634 18808
rect -13582 18756 -13510 18808
rect -13458 18806 -12465 18808
rect -12409 18806 -12341 18862
rect -12285 18806 -12217 18862
rect -12161 18806 -12093 18862
rect -12037 18810 -10439 18862
rect -12037 18806 -10918 18810
rect -13458 18756 -10918 18806
rect -15247 18754 -10918 18756
rect -10862 18754 -10794 18810
rect -10738 18754 -10670 18810
rect -10614 18754 -10546 18810
rect -10490 18754 -10439 18810
rect -15247 18738 -10439 18754
rect -15247 18684 -12465 18738
rect -15247 18632 -13882 18684
rect -13830 18632 -13758 18684
rect -13706 18632 -13634 18684
rect -13582 18632 -13510 18684
rect -13458 18682 -12465 18684
rect -12409 18682 -12341 18738
rect -12285 18682 -12217 18738
rect -12161 18682 -12093 18738
rect -12037 18686 -10439 18738
rect -12037 18682 -10918 18686
rect -13458 18632 -10918 18682
rect -15247 18630 -10918 18632
rect -10862 18630 -10794 18686
rect -10738 18630 -10670 18686
rect -10614 18630 -10546 18686
rect -10490 18630 -10439 18686
rect -15247 18614 -10439 18630
rect -15247 18560 -12465 18614
rect -15247 18508 -13882 18560
rect -13830 18508 -13758 18560
rect -13706 18508 -13634 18560
rect -13582 18508 -13510 18560
rect -13458 18558 -12465 18560
rect -12409 18558 -12341 18614
rect -12285 18558 -12217 18614
rect -12161 18558 -12093 18614
rect -12037 18562 -10439 18614
rect -12037 18558 -10918 18562
rect -13458 18508 -10918 18558
rect -15247 18506 -10918 18508
rect -10862 18506 -10794 18562
rect -10738 18506 -10670 18562
rect -10614 18506 -10546 18562
rect -10490 18506 -10439 18562
rect -15247 18490 -10439 18506
rect -15247 18436 -12465 18490
rect -15247 18384 -13882 18436
rect -13830 18384 -13758 18436
rect -13706 18384 -13634 18436
rect -13582 18384 -13510 18436
rect -13458 18434 -12465 18436
rect -12409 18434 -12341 18490
rect -12285 18434 -12217 18490
rect -12161 18434 -12093 18490
rect -12037 18438 -10439 18490
rect -12037 18434 -10918 18438
rect -13458 18384 -10918 18434
rect -15247 18382 -10918 18384
rect -10862 18382 -10794 18438
rect -10738 18382 -10670 18438
rect -10614 18382 -10546 18438
rect -10490 18382 -10439 18438
rect -15247 17722 -10439 18382
rect -15247 17670 -13966 17722
rect -13914 17670 -13842 17722
rect -13790 17670 -13718 17722
rect -13666 17670 -13594 17722
rect -13542 17714 -10439 17722
rect -13542 17670 -12463 17714
rect -15247 17662 -12463 17670
rect -12411 17662 -12339 17714
rect -12287 17662 -12215 17714
rect -12163 17662 -12091 17714
rect -12039 17662 -10439 17714
rect -15247 17598 -10439 17662
rect -15247 17546 -13966 17598
rect -13914 17546 -13842 17598
rect -13790 17546 -13718 17598
rect -13666 17546 -13594 17598
rect -13542 17590 -10439 17598
rect -13542 17546 -12463 17590
rect -15247 17538 -12463 17546
rect -12411 17538 -12339 17590
rect -12287 17538 -12215 17590
rect -12163 17538 -12091 17590
rect -12039 17538 -10439 17590
rect -15247 17474 -10439 17538
rect -15247 17422 -13966 17474
rect -13914 17422 -13842 17474
rect -13790 17422 -13718 17474
rect -13666 17422 -13594 17474
rect -13542 17466 -10439 17474
rect -13542 17422 -12463 17466
rect -15247 17414 -12463 17422
rect -12411 17414 -12339 17466
rect -12287 17414 -12215 17466
rect -12163 17414 -12091 17466
rect -12039 17414 -10439 17466
rect -15247 17350 -10439 17414
rect -15247 17298 -13966 17350
rect -13914 17298 -13842 17350
rect -13790 17298 -13718 17350
rect -13666 17298 -13594 17350
rect -13542 17342 -10439 17350
rect -13542 17298 -12463 17342
rect -15247 17290 -12463 17298
rect -12411 17290 -12339 17342
rect -12287 17290 -12215 17342
rect -12163 17290 -12091 17342
rect -12039 17290 -10439 17342
rect -15247 16941 -10439 17290
rect 2458 16522 2515 16888
rect -198 15447 -142 15448
rect -298 15391 -132 15447
rect -198 15252 -142 15391
rect 2503 15111 2561 15299
rect 3968 14743 4219 14775
rect 3968 14687 4005 14743
rect 4061 14687 4132 14743
rect 4188 14687 4219 14743
rect 3968 14651 4219 14687
rect 1122 14386 1678 14442
rect 2080 14352 2136 14528
rect 919 13812 975 14048
rect -16003 13290 -12360 13755
rect -16003 13275 -13209 13290
rect -16003 13252 -14239 13275
rect -16003 13200 -15546 13252
rect -15494 13200 -15422 13252
rect -15370 13200 -15298 13252
rect -15246 13200 -15174 13252
rect -15122 13219 -14239 13252
rect -14183 13219 -14115 13275
rect -14059 13219 -13991 13275
rect -13935 13219 -13867 13275
rect -13811 13234 -13209 13275
rect -13153 13234 -13085 13290
rect -13029 13234 -12961 13290
rect -12905 13234 -12837 13290
rect -12781 13234 -12360 13290
rect -13811 13219 -12360 13234
rect -15122 13200 -12360 13219
rect -16003 13166 -12360 13200
rect -16003 13151 -13209 13166
rect -16003 13128 -14239 13151
rect -16003 13076 -15546 13128
rect -15494 13076 -15422 13128
rect -15370 13076 -15298 13128
rect -15246 13076 -15174 13128
rect -15122 13095 -14239 13128
rect -14183 13095 -14115 13151
rect -14059 13095 -13991 13151
rect -13935 13095 -13867 13151
rect -13811 13110 -13209 13151
rect -13153 13110 -13085 13166
rect -13029 13110 -12961 13166
rect -12905 13110 -12837 13166
rect -12781 13110 -12360 13166
rect -13811 13095 -12360 13110
rect -15122 13076 -12360 13095
rect -16003 13042 -12360 13076
rect -16003 13027 -13209 13042
rect -16003 13004 -14239 13027
rect -16003 12952 -15546 13004
rect -15494 12952 -15422 13004
rect -15370 12952 -15298 13004
rect -15246 12952 -15174 13004
rect -15122 12971 -14239 13004
rect -14183 12971 -14115 13027
rect -14059 12971 -13991 13027
rect -13935 12971 -13867 13027
rect -13811 12986 -13209 13027
rect -13153 12986 -13085 13042
rect -13029 12986 -12961 13042
rect -12905 12986 -12837 13042
rect -12781 12986 -12360 13042
rect -13811 12971 -12360 12986
rect -15122 12952 -12360 12971
rect -16003 12918 -12360 12952
rect -16003 12903 -13209 12918
rect -16003 12880 -14239 12903
rect -16003 12828 -15546 12880
rect -15494 12828 -15422 12880
rect -15370 12828 -15298 12880
rect -15246 12828 -15174 12880
rect -15122 12847 -14239 12880
rect -14183 12847 -14115 12903
rect -14059 12847 -13991 12903
rect -13935 12847 -13867 12903
rect -13811 12862 -13209 12903
rect -13153 12862 -13085 12918
rect -13029 12862 -12961 12918
rect -12905 12862 -12837 12918
rect -12781 12862 -12360 12918
rect -13811 12847 -12360 12862
rect -15122 12828 -12360 12847
rect -16003 12531 -12360 12828
rect 1943 11782 1999 12188
rect 8582 11731 8987 21236
rect 41677 20265 44259 20474
rect 14077 19524 16649 19580
rect 14077 19472 14140 19524
rect 14192 19472 14311 19524
rect 14363 19472 14482 19524
rect 14534 19472 14653 19524
rect 14705 19472 14824 19524
rect 14876 19472 14995 19524
rect 15047 19472 15166 19524
rect 15218 19472 15337 19524
rect 15389 19472 15508 19524
rect 15560 19472 15679 19524
rect 15731 19472 15850 19524
rect 15902 19472 16021 19524
rect 16073 19472 16192 19524
rect 16244 19472 16363 19524
rect 16415 19472 16534 19524
rect 16586 19472 16649 19524
rect 14077 19370 16649 19472
rect 14077 19359 23289 19370
rect 14077 19307 14140 19359
rect 14192 19307 14311 19359
rect 14363 19307 14482 19359
rect 14534 19307 14653 19359
rect 14705 19307 14824 19359
rect 14876 19307 14995 19359
rect 15047 19307 15166 19359
rect 15218 19307 15337 19359
rect 15389 19307 15508 19359
rect 15560 19307 15679 19359
rect 15731 19307 15850 19359
rect 15902 19307 16021 19359
rect 16073 19307 16192 19359
rect 16244 19307 16363 19359
rect 16415 19307 16534 19359
rect 16586 19307 23289 19359
rect 14077 19194 23289 19307
rect 14077 19142 14140 19194
rect 14192 19142 14311 19194
rect 14363 19142 14482 19194
rect 14534 19142 14653 19194
rect 14705 19142 14824 19194
rect 14876 19142 14995 19194
rect 15047 19142 15166 19194
rect 15218 19142 15337 19194
rect 15389 19142 15508 19194
rect 15560 19142 15679 19194
rect 15731 19142 15850 19194
rect 15902 19142 16021 19194
rect 16073 19142 16192 19194
rect 16244 19142 16363 19194
rect 16415 19142 16534 19194
rect 16586 19142 23289 19194
rect 14077 19031 23289 19142
rect 22950 18662 23289 19031
rect 22949 18577 23289 18662
rect 22949 18238 29869 18577
rect 9800 17596 10310 17660
rect 9800 17544 9836 17596
rect 9888 17544 9964 17596
rect 10016 17593 10310 17596
rect 10016 17544 10115 17593
rect 9800 17541 10115 17544
rect 10167 17541 10310 17593
rect 9800 17470 10310 17541
rect 9800 17437 21600 17470
rect 9800 17385 9834 17437
rect 9886 17435 10181 17437
rect 9886 17385 10005 17435
rect 9800 17383 10005 17385
rect 10057 17385 10181 17435
rect 10233 17385 21600 17437
rect 10057 17383 21600 17385
rect 9800 17274 21600 17383
rect 9800 17258 10197 17274
rect 9800 17253 10048 17258
rect 9800 17201 9846 17253
rect 9898 17206 10048 17253
rect 10100 17222 10197 17258
rect 10249 17250 21600 17274
rect 10249 17222 10310 17250
rect 10100 17206 10310 17222
rect 9898 17201 10310 17206
rect 9800 17160 10310 17201
rect 9750 16933 10260 16990
rect 9750 16926 10054 16933
rect 9750 16923 9923 16926
rect 9750 16871 9795 16923
rect 9847 16874 9923 16923
rect 9975 16881 10054 16926
rect 10106 16914 10260 16933
rect 10106 16881 20684 16914
rect 9975 16874 20684 16881
rect 9847 16871 20684 16874
rect 9750 16749 20684 16871
rect 9750 16744 10107 16749
rect 9750 16726 9959 16744
rect 9750 16674 9790 16726
rect 9842 16692 9959 16726
rect 10011 16697 10107 16744
rect 10159 16697 20684 16749
rect 10011 16692 20684 16697
rect 9842 16674 20684 16692
rect 9750 16646 20684 16674
rect 9750 16616 10260 16646
rect 9750 16606 10141 16616
rect 9750 16575 9964 16606
rect 9750 16523 9767 16575
rect 9819 16554 9964 16575
rect 10016 16564 10141 16606
rect 10193 16564 10260 16616
rect 10016 16554 10260 16564
rect 9819 16523 10260 16554
rect 9750 16490 10260 16523
rect 12240 16138 19962 16431
rect 12240 14461 12533 16138
rect 19669 15309 19962 16138
rect 20416 15743 20684 16646
rect 21380 16087 21600 17250
rect 26344 16826 26987 16880
rect 26344 16774 26428 16826
rect 26480 16774 26548 16826
rect 26600 16774 26668 16826
rect 26720 16774 26788 16826
rect 26840 16774 26908 16826
rect 26960 16799 26987 16826
rect 29530 16799 29869 18238
rect 26960 16774 37528 16799
rect 26344 16706 37528 16774
rect 26344 16654 26428 16706
rect 26480 16654 26548 16706
rect 26600 16654 26668 16706
rect 26720 16654 26788 16706
rect 26840 16654 26908 16706
rect 26960 16654 37528 16706
rect 26344 16594 37528 16654
rect 26344 16591 26987 16594
rect 22735 16494 23393 16495
rect 22735 16431 36567 16494
rect 22735 16379 22822 16431
rect 22874 16379 22942 16431
rect 22994 16379 23062 16431
rect 23114 16379 23182 16431
rect 23234 16379 23302 16431
rect 23354 16379 36567 16431
rect 22735 16311 36567 16379
rect 22735 16259 22822 16311
rect 22874 16259 22942 16311
rect 22994 16259 23062 16311
rect 23114 16259 23182 16311
rect 23234 16259 23302 16311
rect 23354 16289 36567 16311
rect 23354 16259 23393 16289
rect 22735 16210 23393 16259
rect 21380 15884 35629 16087
rect 20416 15712 24234 15743
rect 20416 15506 33629 15712
rect 20416 15475 24234 15506
rect 19669 15286 23314 15309
rect 19669 15250 31910 15286
rect 19669 15198 22094 15250
rect 22146 15198 22214 15250
rect 22266 15198 22334 15250
rect 22386 15198 22454 15250
rect 22506 15198 22574 15250
rect 22626 15198 31910 15250
rect 19669 15130 31910 15198
rect 10823 14168 12533 14461
rect 12941 14846 19271 15094
rect 19669 15078 22094 15130
rect 22146 15078 22214 15130
rect 22266 15078 22334 15130
rect 22386 15078 22454 15130
rect 22506 15078 22574 15130
rect 22626 15078 31910 15130
rect 19669 15039 31910 15078
rect 19669 15016 23314 15039
rect 10823 13450 11116 14168
rect 10823 13398 10858 13450
rect 10910 13398 10996 13450
rect 11048 13398 11116 13450
rect 10823 13323 11116 13398
rect 10823 13271 10861 13323
rect 10913 13321 11116 13323
rect 10913 13271 11000 13321
rect 10823 13269 11000 13271
rect 11052 13269 11116 13321
rect 10823 13179 11116 13269
rect 10823 13170 11000 13179
rect 10823 13118 10860 13170
rect 10912 13127 11000 13170
rect 11052 13127 11116 13179
rect 10912 13118 11116 13127
rect 10823 13099 11116 13118
rect 10999 12864 11286 12914
rect 10999 12808 11044 12864
rect 11100 12808 11182 12864
rect 11238 12808 11286 12864
rect 10999 12732 11286 12808
rect 10999 12728 11171 12732
rect 10999 12672 11044 12728
rect 11100 12676 11171 12728
rect 11227 12676 11286 12732
rect 11100 12672 11286 12676
rect 10999 12626 11286 12672
rect 12236 12459 12529 12469
rect 12236 12415 12533 12459
rect 12236 12363 12271 12415
rect 12323 12363 12409 12415
rect 12461 12363 12533 12415
rect 12236 12288 12533 12363
rect 12236 12236 12274 12288
rect 12326 12286 12533 12288
rect 12326 12236 12413 12286
rect 12236 12234 12413 12236
rect 12465 12234 12533 12286
rect 12236 12144 12533 12234
rect 12236 12135 12413 12144
rect 12236 12083 12273 12135
rect 12325 12092 12413 12135
rect 12465 12092 12533 12144
rect 12325 12083 12533 12092
rect 12236 12064 12533 12083
rect 8578 11667 8995 11731
rect 8578 11664 8873 11667
rect 8578 11663 8727 11664
rect 8578 11607 8607 11663
rect 8663 11608 8727 11663
rect 8783 11611 8873 11664
rect 8929 11611 8995 11667
rect 8783 11608 8995 11611
rect 8663 11607 8995 11608
rect 8578 11552 8995 11607
rect 8578 11496 8612 11552
rect 8668 11496 8743 11552
rect 8799 11496 8883 11552
rect 8939 11496 8995 11552
rect 8578 11488 8995 11496
rect 2211 10352 2759 10425
rect -9408 9642 -8737 9680
rect 2686 9642 2759 10352
rect 11239 10062 11632 10070
rect 12240 10062 12533 12064
rect 11238 10056 12533 10062
rect 11236 9990 12533 10056
rect 11236 9979 11521 9990
rect 11236 9927 11344 9979
rect 11396 9938 11521 9979
rect 11573 9938 12533 9990
rect 11396 9927 12533 9938
rect 11236 9858 12533 9927
rect 11236 9848 11414 9858
rect 11236 9796 11278 9848
rect 11330 9806 11414 9848
rect 11466 9853 12533 9858
rect 11466 9806 11561 9853
rect 11330 9801 11561 9806
rect 11613 9801 12533 9853
rect 11330 9796 12533 9801
rect 11236 9772 12533 9796
rect 11238 9769 12533 9772
rect -9408 9631 2759 9642
rect -9408 9579 -9354 9631
rect -9302 9579 -8805 9631
rect -8753 9579 2759 9631
rect -9408 9569 2759 9579
rect -9408 9519 -8737 9569
rect 2329 9019 3267 9045
rect -9415 8964 3267 9019
rect -9415 8915 2389 8964
rect -9415 8863 -9334 8915
rect -9282 8863 -8785 8915
rect -8733 8912 2389 8915
rect 2441 8912 2711 8964
rect 2763 8912 3267 8964
rect -8733 8863 3267 8912
rect -9415 8790 3267 8863
rect 12941 8826 13189 14846
rect 19023 14678 19271 14846
rect 22059 14694 22659 14696
rect 22045 14678 22661 14694
rect 19023 14632 30057 14678
rect 19023 14580 22063 14632
rect 22115 14580 22183 14632
rect 22235 14580 22303 14632
rect 22355 14580 22423 14632
rect 22475 14580 22543 14632
rect 22595 14580 30057 14632
rect 19023 14512 30057 14580
rect 19023 14460 22063 14512
rect 22115 14460 22183 14512
rect 22235 14460 22303 14512
rect 22355 14460 22423 14512
rect 22475 14460 22543 14512
rect 22595 14460 30057 14512
rect 19023 14430 30057 14460
rect 22045 14427 22661 14430
rect 17357 14268 18262 14318
rect 17357 14180 17931 14268
rect 17357 14160 17795 14180
rect 17357 14104 17580 14160
rect 17636 14124 17795 14160
rect 17851 14124 17931 14180
rect 17636 14104 17931 14124
rect 17357 14008 17931 14104
rect 18191 14008 18262 14268
rect 17357 14007 18262 14008
rect 17357 13997 17731 14007
rect 17357 13941 17469 13997
rect 17525 13951 17731 13997
rect 17787 13951 18262 14007
rect 17525 13945 18262 13951
rect 17525 13943 17920 13945
rect 17976 13943 18262 13945
rect 17525 13941 17919 13943
rect 17357 13787 17919 13941
rect 18179 13787 18262 13943
rect 17357 13756 18262 13787
rect 17357 13746 17707 13756
rect 17357 13690 17487 13746
rect 17543 13700 17707 13746
rect 17763 13700 18262 13756
rect 17543 13695 18262 13700
rect 17543 13690 17924 13695
rect 17357 13639 17924 13690
rect 17980 13639 18262 13695
rect 17357 13551 18262 13639
rect 19111 14167 19532 14279
rect 19111 14115 19181 14167
rect 19233 14115 19412 14167
rect 19464 14115 19532 14167
rect 19111 13953 19532 14115
rect 19111 13901 19179 13953
rect 19231 13901 19401 13953
rect 19453 13901 19532 13953
rect 19111 13731 19532 13901
rect 20130 14145 20656 14238
rect 20130 14104 20725 14145
rect 20130 14094 20480 14104
rect 20130 14038 20260 14094
rect 20316 14091 20480 14094
rect 20536 14091 20725 14104
rect 20316 14038 20393 14091
rect 20130 13905 20393 14038
rect 20130 13849 20251 13905
rect 20307 13849 20393 13905
rect 20130 13831 20393 13849
rect 20653 13831 20725 14091
rect 22087 14087 23144 14135
rect 22087 14084 28904 14087
rect 22087 13928 22116 14084
rect 22272 13928 22498 14084
rect 22654 13928 22917 14084
rect 23073 13928 28904 14084
rect 22087 13926 28904 13928
rect 22087 13904 23144 13926
rect 20130 13787 20725 13831
rect 19111 13723 19389 13731
rect 19111 13671 19178 13723
rect 19230 13679 19389 13723
rect 19441 13679 19532 13731
rect 19230 13671 19532 13679
rect 19111 13591 19532 13671
rect 11423 8578 13189 8826
rect 13467 13461 13922 13516
rect 17357 13495 17705 13551
rect 17761 13495 18262 13551
rect 17357 13461 18262 13495
rect 13467 13285 18262 13461
rect 13467 13116 18226 13285
rect 11423 7982 11671 8578
rect 11423 7930 11440 7982
rect 11492 7930 11574 7982
rect 11626 7930 11671 7982
rect 11423 7868 11671 7930
rect 11423 7816 11435 7868
rect 11487 7856 11671 7868
rect 11487 7816 11564 7856
rect 11423 7804 11564 7816
rect 11616 7804 11671 7856
rect 11423 7781 11671 7804
rect -1513 7356 1298 7366
rect -1513 7255 1309 7356
rect -1513 7252 1047 7255
rect -1513 7231 644 7252
rect -1513 7214 137 7231
rect -1513 7186 -260 7214
rect -1513 7130 -1242 7186
rect -1186 7158 -260 7186
rect -204 7179 137 7214
rect 189 7200 644 7231
rect 696 7203 1047 7252
rect 1099 7203 1309 7255
rect 696 7200 1309 7203
rect 189 7179 1309 7200
rect -204 7158 1309 7179
rect -1186 7130 1309 7158
rect 12940 7305 13192 7311
rect 12940 7253 12966 7305
rect 13018 7253 13102 7305
rect 13154 7253 13192 7305
rect 12940 7192 13192 7253
rect 12940 7140 12961 7192
rect 13013 7185 13192 7192
rect 13013 7140 13097 7185
rect -1513 6968 1309 7130
rect -1513 6961 910 6968
rect -1513 6923 511 6961
rect -1513 6871 95 6923
rect 147 6909 511 6923
rect 563 6916 910 6961
rect 962 6916 1309 6968
rect 563 6909 1309 6916
rect 147 6871 1309 6909
rect 8560 7075 9108 7137
rect 12940 7133 13097 7140
rect 13149 7133 13192 7185
rect 12940 7111 13192 7133
rect 8560 7068 8951 7075
rect 8560 7012 8590 7068
rect 8650 7016 8731 7068
rect 8793 7019 8951 7068
rect 9007 7019 9108 7075
rect 8793 7016 9108 7019
rect 8646 7012 8731 7016
rect 8787 7012 9108 7016
rect 8560 6958 9108 7012
rect 8560 6902 8596 6958
rect 8652 6956 9108 6958
rect 8652 6953 8746 6956
rect 8798 6953 8984 6956
rect 8652 6902 8737 6953
rect 8798 6904 8977 6953
rect 9036 6904 9108 6956
rect 8560 6897 8737 6902
rect 8793 6897 8977 6904
rect 9033 6897 9108 6904
rect 8560 6879 9108 6897
rect -1513 6861 1309 6871
rect -1513 6805 -404 6861
rect -348 6805 1309 6861
rect -1513 6724 1309 6805
rect -1513 6668 -989 6724
rect -933 6668 1309 6724
rect -1513 6646 1309 6668
rect -1513 6632 998 6646
rect -1513 6608 644 6632
rect -1513 6604 266 6608
rect -1513 6552 -7 6604
rect 45 6556 266 6604
rect 318 6580 644 6608
rect 696 6594 998 6632
rect 1050 6594 1309 6646
rect 696 6580 1309 6594
rect 318 6556 1309 6580
rect 45 6552 1309 6556
rect -1513 6370 1309 6552
rect -1513 6314 -440 6370
rect -384 6314 1309 6370
rect -1513 6240 1309 6314
rect -1513 6184 -996 6240
rect -940 6187 1309 6240
rect -940 6184 620 6187
rect -1513 6135 620 6184
rect 672 6135 1309 6187
rect -1513 5879 1309 6135
rect -1513 5811 1298 5879
rect -1500 3460 -1072 5811
rect 12397 5486 12483 5488
rect 12397 5469 12848 5486
rect 12382 5466 12848 5469
rect 12941 5466 13189 7111
rect 12382 5403 13189 5466
rect 12382 5392 12679 5403
rect 12382 5340 12502 5392
rect 12554 5351 12679 5392
rect 12731 5351 13189 5403
rect 12554 5340 13189 5351
rect 12382 5271 13189 5340
rect 12382 5261 12572 5271
rect 12382 5209 12436 5261
rect 12488 5219 12572 5261
rect 12624 5266 13189 5271
rect 12624 5219 12719 5266
rect 12488 5214 12719 5219
rect 12771 5218 13189 5266
rect 12771 5214 12848 5218
rect 12488 5209 12848 5214
rect 12382 5176 12848 5209
rect -1531 3336 -1072 3460
rect 4463 3808 5878 3909
rect 4463 3805 5616 3808
rect 4463 3784 5213 3805
rect 4463 3732 4706 3784
rect 4758 3753 5213 3784
rect 5265 3756 5616 3805
rect 5668 3756 5878 3808
rect 5265 3753 5878 3756
rect 4758 3732 5878 3753
rect 4463 3521 5878 3732
rect 4463 3514 5479 3521
rect 4463 3476 5080 3514
rect 4463 3424 4664 3476
rect 4716 3462 5080 3476
rect 5132 3469 5479 3514
rect 5531 3469 5878 3521
rect 5132 3462 5878 3469
rect 4716 3424 5878 3462
rect 4463 3336 5878 3424
rect -1531 3199 6122 3336
rect -1531 3185 5567 3199
rect -1531 3161 5213 3185
rect -1531 3157 4835 3161
rect -1531 3105 4562 3157
rect 4614 3109 4835 3157
rect 4887 3133 5213 3161
rect 5265 3147 5567 3185
rect 5619 3147 6122 3199
rect 5265 3133 6122 3147
rect 4887 3109 6122 3133
rect 4614 3105 6122 3109
rect -1531 2908 6122 3105
rect -1531 1445 -1103 2908
rect 4463 2905 5878 2908
rect -3741 1372 -447 1445
rect -3741 1358 -3106 1372
rect -3741 1098 -3695 1358
rect -3435 1112 -3106 1358
rect -2846 1334 -447 1372
rect -2846 1174 -1958 1334
rect -1798 1322 -447 1334
rect -1798 1174 -1368 1322
rect -2846 1162 -1368 1174
rect -1208 1308 -447 1322
rect -1208 1162 -693 1308
rect -2846 1148 -693 1162
rect -533 1148 -447 1308
rect -2846 1112 -447 1148
rect -3435 1098 -447 1112
rect -3741 1068 -447 1098
rect -2319 300 931 372
rect -2789 299 931 300
rect -2789 285 -1728 299
rect -2789 25 -2317 285
rect -2057 39 -1728 285
rect -1468 261 931 299
rect -1468 101 -580 261
rect -420 249 931 261
rect -420 101 10 249
rect -1468 89 10 101
rect 170 235 931 249
rect 170 89 685 235
rect -1468 75 685 89
rect 845 75 931 235
rect -1468 39 931 75
rect -2057 25 931 39
rect -2789 14 931 25
rect -2319 -5 931 14
rect 2197 -257 3075 -188
rect 2197 -313 2725 -257
rect 2781 -259 3075 -257
rect 2781 -313 2889 -259
rect 2197 -315 2889 -313
rect 2945 -315 3075 -259
rect 2197 -371 3075 -315
rect 2197 -384 2891 -371
rect 2197 -440 2725 -384
rect 2781 -427 2891 -384
rect 2947 -427 3075 -371
rect 2781 -440 3075 -427
rect 2197 -511 3075 -440
rect 2197 -522 2896 -511
rect 2197 -578 2725 -522
rect 2781 -567 2896 -522
rect 2952 -567 3075 -511
rect 2781 -578 3075 -567
rect 2197 -634 3075 -578
rect 4778 -988 5148 -932
rect 4778 -1044 4826 -988
rect 4882 -990 5148 -988
rect 4882 -1044 4990 -990
rect 4778 -1046 4990 -1044
rect 5046 -1046 5148 -990
rect 4778 -1102 5148 -1046
rect 4778 -1115 4992 -1102
rect 4778 -1171 4826 -1115
rect 4882 -1158 4992 -1115
rect 5048 -1158 5148 -1102
rect 4882 -1171 5148 -1158
rect 4778 -1242 5148 -1171
rect 4778 -1253 4997 -1242
rect 4778 -1309 4826 -1253
rect 4882 -1298 4997 -1253
rect 5053 -1298 5148 -1242
rect 4882 -1309 5148 -1298
rect 4778 -1338 5148 -1309
rect 4844 -1554 5214 -1512
rect 4844 -1567 5058 -1554
rect 4844 -1623 4892 -1567
rect 4948 -1610 5058 -1567
rect 5114 -1610 5214 -1554
rect 4948 -1623 5214 -1610
rect 4844 -1694 5214 -1623
rect 4844 -1705 5063 -1694
rect 4844 -1761 4892 -1705
rect 4948 -1750 5063 -1705
rect 5119 -1750 5214 -1694
rect 4948 -1761 5214 -1750
rect 4844 -1790 5214 -1761
rect 4506 -2253 4874 -2240
rect 4506 -2305 4796 -2253
rect 4848 -2255 4874 -2253
rect 4848 -2305 11467 -2255
rect 4506 -2356 11467 -2305
rect 4506 -2408 4547 -2356
rect 4599 -2408 4687 -2356
rect 4739 -2408 11467 -2356
rect 4506 -2455 11467 -2408
rect 4506 -2477 4874 -2455
rect 4506 -2529 4549 -2477
rect 4601 -2480 4874 -2477
rect 4601 -2529 4695 -2480
rect 4506 -2532 4695 -2529
rect 4747 -2485 4874 -2480
rect 4747 -2532 4815 -2485
rect 4506 -2537 4815 -2532
rect 4867 -2537 4874 -2485
rect 4506 -2563 4874 -2537
rect 5001 -2650 5371 -2608
rect 5001 -2663 5215 -2650
rect 5001 -2719 5049 -2663
rect 5105 -2706 5215 -2663
rect 5271 -2706 5371 -2650
rect 5105 -2719 5371 -2706
rect 5001 -2790 5371 -2719
rect 5001 -2801 5220 -2790
rect 5001 -2857 5049 -2801
rect 5105 -2846 5220 -2801
rect 5276 -2846 5371 -2790
rect 5105 -2857 5371 -2846
rect 5001 -2886 5371 -2857
rect 4905 -3068 5275 -3026
rect 4905 -3081 5119 -3068
rect 4905 -3137 4953 -3081
rect 5009 -3124 5119 -3081
rect 5175 -3124 5275 -3068
rect 5009 -3137 5275 -3124
rect 4905 -3208 5275 -3137
rect 4905 -3219 5124 -3208
rect 4905 -3275 4953 -3219
rect 5009 -3264 5124 -3219
rect 5180 -3264 5275 -3208
rect 5009 -3275 5275 -3264
rect 4905 -3304 5275 -3275
rect 4882 -3482 5252 -3440
rect 4882 -3495 5096 -3482
rect 4882 -3551 4930 -3495
rect 4986 -3538 5096 -3495
rect 5152 -3538 5252 -3482
rect 4986 -3551 5252 -3538
rect 4882 -3622 5252 -3551
rect 4882 -3633 5101 -3622
rect 4882 -3689 4930 -3633
rect 4986 -3678 5101 -3633
rect 5157 -3678 5252 -3622
rect 4986 -3689 5252 -3678
rect 4882 -3718 5252 -3689
rect 11285 -3874 11467 -2455
rect 13467 -3380 13922 13116
rect 17908 12969 18198 13116
rect 19228 12977 19380 13591
rect 20406 12980 20725 13787
rect 21938 13658 22849 13700
rect 25430 13658 26138 13671
rect 21938 13618 26138 13658
rect 21938 13616 25520 13618
rect 21938 13564 22006 13616
rect 22058 13564 22429 13616
rect 22481 13564 22720 13616
rect 22772 13564 25520 13616
rect 21938 13562 25520 13564
rect 25576 13562 25708 13618
rect 25764 13562 25903 13618
rect 25959 13562 26138 13618
rect 21938 13522 26138 13562
rect 21938 13497 22849 13522
rect 25430 13504 26138 13522
rect 25430 13503 26015 13504
rect 21799 13290 22548 13292
rect 21799 13239 25263 13290
rect 21799 13187 21838 13239
rect 21890 13187 22077 13239
rect 22129 13187 22410 13239
rect 22462 13187 25263 13239
rect 21799 13142 25263 13187
rect 22003 13130 25263 13142
rect 17908 12820 18711 12969
rect 19228 12825 19543 12977
rect 19391 12008 19543 12825
rect 20406 12807 22149 12980
rect 21976 12098 22149 12807
rect 25103 12633 25263 13130
rect 25103 12473 28368 12633
rect 21863 11925 22149 12098
rect 27026 11727 27558 11886
rect 28208 11854 28368 12473
rect 28743 12234 28904 13926
rect 29809 13377 30057 14430
rect 29808 13325 30422 13377
rect 29808 13273 29830 13325
rect 29882 13273 29950 13325
rect 30002 13273 30070 13325
rect 30122 13273 30190 13325
rect 30242 13273 30310 13325
rect 30362 13273 30422 13325
rect 29808 13205 30422 13273
rect 29808 13153 29830 13205
rect 29882 13153 29950 13205
rect 30002 13153 30070 13205
rect 30122 13153 30190 13205
rect 30242 13153 30310 13205
rect 30362 13153 30422 13205
rect 29808 13140 30422 13153
rect 28743 12073 30776 12234
rect 30615 11894 30776 12073
rect 23388 11515 23551 11668
rect 27026 11650 27185 11727
rect 28208 11694 30139 11854
rect 30615 11733 30983 11894
rect 26304 11491 27236 11650
rect 19654 11190 19738 11204
rect 19654 11134 19668 11190
rect 19724 11134 19738 11190
rect 19654 11121 19738 11134
rect 19895 11195 19979 11209
rect 19895 11139 19909 11195
rect 19965 11139 19979 11195
rect 19895 11126 19979 11139
rect 20120 11197 20230 11220
rect 20120 11141 20148 11197
rect 20204 11141 20230 11197
rect 20120 11110 20230 11141
rect 20361 11197 20445 11211
rect 20361 11141 20375 11197
rect 20431 11141 20445 11197
rect 20361 11128 20445 11141
rect 22449 11208 22560 11220
rect 22449 11167 22574 11208
rect 21983 11113 22080 11125
rect 22449 11115 22481 11167
rect 22533 11115 22574 11167
rect 22449 11113 22574 11115
rect 21983 11072 22574 11113
rect 21983 11023 22575 11072
rect 21983 10971 22476 11023
rect 22528 10971 22575 11023
rect 21983 10919 22575 10971
rect 21984 10918 22575 10919
rect 27077 11032 27236 11491
rect 27077 10873 27324 11032
rect 29660 10913 29767 11694
rect 30822 10849 30983 11733
rect 31663 9951 31910 15039
rect 33423 12307 33629 15506
rect 33149 12101 33629 12307
rect 33423 11895 33629 12101
rect 28768 9895 28852 9909
rect 28768 9839 28782 9895
rect 28838 9839 28852 9895
rect 28768 9826 28852 9839
rect 29009 9900 29093 9914
rect 29009 9844 29023 9900
rect 29079 9844 29093 9900
rect 29009 9831 29093 9844
rect 29248 9902 29332 9916
rect 29248 9846 29262 9902
rect 29318 9846 29332 9902
rect 29248 9833 29332 9846
rect 29475 9902 29559 9916
rect 29475 9846 29489 9902
rect 29545 9846 29559 9902
rect 29475 9833 29559 9846
rect 30909 9879 32327 9951
rect 35426 9902 35629 15884
rect 36362 11499 36567 16289
rect 37323 12528 37528 16594
rect 41677 15783 41886 20265
rect 48755 18466 96067 18473
rect 48755 18452 96117 18466
rect 48755 18400 95813 18452
rect 95865 18400 95933 18452
rect 95985 18400 96053 18452
rect 96105 18400 96117 18452
rect 48755 18332 96117 18400
rect 48755 18280 95813 18332
rect 95865 18280 95933 18332
rect 95985 18280 96053 18332
rect 96105 18280 96117 18332
rect 48755 18212 96117 18280
rect 48755 18160 95813 18212
rect 95865 18160 95933 18212
rect 95985 18160 96053 18212
rect 96105 18160 96117 18212
rect 48755 18126 96117 18160
rect 48755 18118 96067 18126
rect 37851 14158 38494 14212
rect 37851 14106 37935 14158
rect 37987 14106 38055 14158
rect 38107 14106 38175 14158
rect 38227 14106 38295 14158
rect 38347 14106 38415 14158
rect 38467 14106 38494 14158
rect 37851 14038 38494 14106
rect 37851 13986 37935 14038
rect 37987 13986 38055 14038
rect 38107 13986 38175 14038
rect 38227 13986 38295 14038
rect 38347 13986 38415 14038
rect 38467 13986 38494 14038
rect 37851 13923 38494 13986
rect 37852 10840 37971 13923
rect 38108 10840 38227 13923
rect 38374 10840 38493 13923
rect 41677 12634 41885 15783
rect 39735 12603 41562 12604
rect 39735 12349 41564 12603
rect 37793 10784 38571 10840
rect 37793 10732 37877 10784
rect 37929 10732 37997 10784
rect 38049 10732 38117 10784
rect 38169 10732 38237 10784
rect 38289 10732 38357 10784
rect 38409 10732 38571 10784
rect 37793 10664 38571 10732
rect 37793 10612 37877 10664
rect 37929 10612 37997 10664
rect 38049 10612 38117 10664
rect 38169 10612 38237 10664
rect 38289 10612 38357 10664
rect 38409 10612 38571 10664
rect 37793 10547 38571 10612
rect 38124 10314 38319 10344
rect 30909 9827 32075 9879
rect 32127 9827 32327 9879
rect 30909 9794 32327 9827
rect 34743 9821 35629 9902
rect 31663 9749 31910 9794
rect 32011 9792 32327 9794
rect 32170 9693 32327 9792
rect 35426 9791 35629 9821
rect 38116 9812 38319 10314
rect 35450 9784 35605 9791
rect 35021 9697 35271 9715
rect 34756 9668 35271 9697
rect 34756 9620 35439 9668
rect 34858 9581 35439 9620
rect 38116 9581 38311 9812
rect 34858 9492 38311 9581
rect 29769 9190 31596 9392
rect 35150 9389 38311 9492
rect 35367 9386 38311 9389
rect 41307 9609 41564 12349
rect 41677 12582 41755 12634
rect 41807 12582 41885 12634
rect 41677 12384 41885 12582
rect 41677 12332 41755 12384
rect 41807 12378 41885 12384
rect 41807 12332 42111 12378
rect 41677 12160 42111 12332
rect 41677 12108 41755 12160
rect 41807 12108 42111 12160
rect 41677 12061 42111 12108
rect 19612 9144 19696 9158
rect 19612 9088 19626 9144
rect 19682 9088 19696 9144
rect 19612 9075 19696 9088
rect 19853 9149 19937 9163
rect 19853 9093 19867 9149
rect 19923 9093 19937 9149
rect 19853 9080 19937 9093
rect 20060 9151 20200 9180
rect 20060 9095 20106 9151
rect 20162 9095 20200 9151
rect 20060 9070 20200 9095
rect 20319 9151 20403 9165
rect 20319 9095 20333 9151
rect 20389 9095 20403 9151
rect 20319 9082 20403 9095
rect 26250 8881 27154 9033
rect 29769 8898 29971 9190
rect 30473 9032 30883 9048
rect 30473 9019 30667 9032
rect 30473 8963 30535 9019
rect 30591 8976 30667 9019
rect 30723 9031 30883 9032
rect 30723 8976 30792 9031
rect 30591 8975 30792 8976
rect 30848 8975 30883 9031
rect 30591 8963 30883 8975
rect 30473 8922 30883 8963
rect 30473 8906 30665 8922
rect 21824 8205 22125 8362
rect 14535 7961 18323 8019
rect 14535 7905 14587 7961
rect 14643 7905 14803 7961
rect 14859 7947 18323 7961
rect 14859 7905 15062 7947
rect 14535 7838 15062 7905
rect 14535 7782 14589 7838
rect 14645 7833 15062 7838
rect 14645 7782 14803 7833
rect 14535 7777 14803 7782
rect 14859 7777 15062 7833
rect 14535 7720 15062 7777
rect 19342 7505 19505 8018
rect 21968 7600 22125 8205
rect 27002 8017 27154 8881
rect 29614 8696 30098 8898
rect 30473 8850 30532 8906
rect 30588 8866 30665 8906
rect 30721 8866 30792 8922
rect 30848 8866 30883 8922
rect 30588 8850 30883 8866
rect 30473 8795 30883 8850
rect 30473 8793 30654 8795
rect 30473 8737 30529 8793
rect 30585 8739 30654 8793
rect 30710 8739 30792 8795
rect 30848 8739 30883 8795
rect 30585 8737 30883 8739
rect 30473 8717 30883 8737
rect 22923 7876 23007 7890
rect 22923 7820 22937 7876
rect 22993 7820 23007 7876
rect 22923 7807 23007 7820
rect 23164 7881 23248 7895
rect 23164 7825 23178 7881
rect 23234 7825 23248 7881
rect 23164 7812 23248 7825
rect 23403 7883 23487 7897
rect 23403 7827 23417 7883
rect 23473 7827 23487 7883
rect 23403 7814 23487 7827
rect 23630 7883 23714 7897
rect 23630 7827 23644 7883
rect 23700 7827 23714 7883
rect 27002 7865 27262 8017
rect 23630 7814 23714 7827
rect 19076 7342 19505 7505
rect 21969 7489 22125 7600
rect 21177 7488 22125 7489
rect 19076 6798 19239 7342
rect 20972 7320 22125 7488
rect 15116 6670 19536 6798
rect 15116 6618 18072 6670
rect 18124 6618 18192 6670
rect 18244 6618 18312 6670
rect 18364 6618 18432 6670
rect 18484 6618 18552 6670
rect 18604 6618 18672 6670
rect 18724 6618 18792 6670
rect 18844 6618 18912 6670
rect 18964 6618 19032 6670
rect 19084 6618 19152 6670
rect 19204 6618 19272 6670
rect 19324 6618 19392 6670
rect 19444 6618 19536 6670
rect 15116 6535 19536 6618
rect 15116 6265 15379 6535
rect 15019 6153 15419 6265
rect 15019 5993 15167 6153
rect 15327 5993 15419 6153
rect 20972 6253 21508 7320
rect 22083 6789 26596 6907
rect 28712 6901 28796 6915
rect 28712 6845 28726 6901
rect 28782 6845 28796 6901
rect 28712 6832 28796 6845
rect 28953 6906 29037 6920
rect 28953 6850 28967 6906
rect 29023 6850 29037 6906
rect 28953 6837 29037 6850
rect 29192 6908 29276 6922
rect 29192 6852 29206 6908
rect 29262 6852 29276 6908
rect 29192 6839 29276 6852
rect 29419 6908 29503 6922
rect 29419 6852 29433 6908
rect 29489 6852 29503 6908
rect 29419 6839 29503 6852
rect 22083 6737 22134 6789
rect 22186 6737 22430 6789
rect 22482 6737 26596 6789
rect 22083 6705 26596 6737
rect 22083 6683 22546 6705
rect 15019 5444 15419 5993
rect 18154 6016 19195 6083
rect 18154 6013 18890 6016
rect 18154 5957 18230 6013
rect 18286 6011 18890 6013
rect 18286 5957 18408 6011
rect 18464 6010 18890 6011
rect 18154 5955 18408 5957
rect 18464 5955 18649 6010
rect 18705 5960 18890 6010
rect 18946 5960 19195 6016
rect 18154 5954 18649 5955
rect 18705 5954 19195 5960
rect 18154 5896 19195 5954
rect 20972 5718 22844 6253
rect 15019 5284 15167 5444
rect 15327 5284 15419 5444
rect 15019 4632 15419 5284
rect 15019 4472 15167 4632
rect 15327 4472 15419 4632
rect 15019 4270 15419 4472
rect 18271 -774 18995 -726
rect 18271 -830 18331 -774
rect 18387 -830 18995 -774
rect 18271 -916 18995 -830
rect 18271 -935 18795 -916
rect 18271 -991 18536 -935
rect 18592 -972 18795 -935
rect 18851 -972 18995 -916
rect 18592 -991 18995 -972
rect 18271 -1063 18995 -991
rect 18080 -1531 18860 -1470
rect 18080 -1534 18706 -1531
rect 18080 -1541 18702 -1534
rect 18080 -1544 18452 -1541
rect 18504 -1544 18702 -1541
rect 18080 -1600 18143 -1544
rect 18199 -1600 18452 -1544
rect 18508 -1586 18702 -1544
rect 18508 -1587 18706 -1586
rect 18762 -1587 18860 -1531
rect 18508 -1600 18860 -1587
rect 18080 -1660 18860 -1600
rect 22309 -2588 22844 5718
rect 26394 5828 26596 6705
rect 31394 5828 31596 9190
rect 38043 7647 38298 9386
rect 41307 9354 48122 9609
rect 47867 8400 48122 9354
rect 47690 8252 48122 8400
rect 47690 8228 48258 8252
rect 47690 8176 47793 8228
rect 47845 8176 47949 8228
rect 48001 8176 48258 8228
rect 47690 8137 48258 8176
rect 47690 7940 48260 8137
rect 47852 7647 48122 7648
rect 38043 7392 48122 7647
rect 44110 7124 44460 7130
rect 43227 7106 44715 7124
rect 43227 6946 43283 7106
rect 43443 6946 43826 7106
rect 43986 6946 44536 7106
rect 44696 6946 44715 7106
rect 46136 7080 47059 7119
rect 46136 7075 46935 7080
rect 46136 7019 46193 7075
rect 46249 7072 46935 7075
rect 46249 7070 46719 7072
rect 46249 7019 46439 7070
rect 46136 7014 46439 7019
rect 46495 7016 46719 7070
rect 46775 7024 46935 7072
rect 46991 7024 47059 7080
rect 47852 7063 48122 7392
rect 46775 7016 47059 7024
rect 46495 7014 47059 7016
rect 46136 6961 47059 7014
rect 43227 6919 44715 6946
rect 44110 6850 44480 6919
rect 44110 6810 44460 6850
rect 38263 6610 39669 6671
rect 38263 6450 38310 6610
rect 38470 6608 39669 6610
rect 38470 6452 39342 6608
rect 39498 6452 39669 6608
rect 38470 6450 39669 6452
rect 38263 6430 39669 6450
rect 38287 6418 39669 6430
rect 38287 6414 38493 6418
rect 43759 6076 44718 6127
rect 43759 6020 43823 6076
rect 43879 6063 44718 6076
rect 43879 6020 44072 6063
rect 44128 6062 44718 6063
rect 43759 6007 44072 6020
rect 44128 6058 44528 6062
rect 44128 6007 44306 6058
rect 43759 6002 44306 6007
rect 44362 6006 44528 6058
rect 44584 6006 44718 6062
rect 44362 6002 44718 6006
rect 43759 5971 44718 6002
rect 26394 5626 31596 5828
rect 27261 4463 27365 4884
rect 30400 4489 30604 4659
rect 27094 4407 27485 4463
rect 27094 4351 27147 4407
rect 27203 4351 27379 4407
rect 27435 4351 27485 4407
rect 27094 4211 27485 4351
rect 27094 4155 27144 4211
rect 27200 4155 27379 4211
rect 27435 4155 27485 4211
rect 27094 4108 27485 4155
rect 30400 4433 30468 4489
rect 30524 4433 30604 4489
rect 30400 4228 30604 4433
rect 30400 4172 30468 4228
rect 30524 4172 30604 4228
rect 30400 4129 30604 4172
rect 42506 3896 42578 4557
rect 43641 4181 43717 4559
rect 47853 4548 48122 7063
rect 45792 4279 48122 4548
rect 48835 4181 49030 18118
rect 43641 4105 49030 4181
rect 49748 16826 96229 16841
rect 49748 16774 95925 16826
rect 95977 16774 96045 16826
rect 96097 16774 96165 16826
rect 96217 16774 96229 16826
rect 49748 16706 96229 16774
rect 49748 16654 95925 16706
rect 95977 16654 96045 16706
rect 96097 16654 96165 16706
rect 96217 16654 96229 16706
rect 49748 16586 96229 16654
rect 49748 16534 95925 16586
rect 95977 16534 96045 16586
rect 96097 16534 96165 16586
rect 96217 16534 96229 16586
rect 49748 16489 96229 16534
rect 49748 4178 50100 16489
rect 56872 15638 96169 15678
rect 56872 15586 95787 15638
rect 95839 15586 95907 15638
rect 95959 15586 96027 15638
rect 96079 15586 96169 15638
rect 56872 15518 96169 15586
rect 56872 15466 95787 15518
rect 95839 15466 95907 15518
rect 95959 15466 96027 15518
rect 96079 15466 96169 15518
rect 56872 15398 96169 15466
rect 56872 15346 95787 15398
rect 95839 15346 95907 15398
rect 95959 15346 96027 15398
rect 96079 15346 96169 15398
rect 56872 15281 96169 15346
rect 53921 9318 54794 9377
rect 53921 9317 54372 9318
rect 53921 9314 54248 9317
rect 53921 9258 54012 9314
rect 54068 9258 54131 9314
rect 54187 9261 54248 9314
rect 54304 9262 54372 9317
rect 54428 9317 54794 9318
rect 54428 9262 54489 9317
rect 54304 9261 54489 9262
rect 54545 9261 54794 9317
rect 54187 9258 54794 9261
rect 53921 9204 54794 9258
rect 53921 9200 54373 9204
rect 53921 9198 54253 9200
rect 53921 9142 54012 9198
rect 54068 9142 54130 9198
rect 54186 9144 54253 9198
rect 54309 9148 54373 9200
rect 54429 9197 54794 9204
rect 54429 9148 54491 9197
rect 54309 9147 54374 9148
rect 54426 9147 54491 9148
rect 54309 9144 54491 9147
rect 54186 9142 54491 9144
rect 53921 9141 54491 9142
rect 54547 9141 54794 9197
rect 53921 9088 54794 9141
rect 56872 6920 57269 15281
rect 95584 14604 96107 14621
rect 95584 14595 95801 14604
rect 62288 14552 95801 14595
rect 95853 14552 95921 14604
rect 95973 14552 96041 14604
rect 96093 14552 96107 14604
rect 62288 14484 96107 14552
rect 62288 14432 95801 14484
rect 95853 14432 95921 14484
rect 95973 14432 96041 14484
rect 96093 14432 96107 14484
rect 62288 14364 96107 14432
rect 62288 14312 95801 14364
rect 95853 14312 95921 14364
rect 95973 14312 96041 14364
rect 96093 14312 96107 14364
rect 62288 14299 96107 14312
rect 62297 11311 62576 14299
rect 95584 14267 96107 14299
rect 64769 13772 65603 13916
rect 64769 13720 64929 13772
rect 64981 13768 65603 13772
rect 64981 13720 65188 13768
rect 64769 13716 65188 13720
rect 65240 13759 65603 13768
rect 65240 13716 71106 13759
rect 64769 13703 71106 13716
rect 64769 13651 65429 13703
rect 65481 13651 71106 13703
rect 64769 13621 71106 13651
rect 64769 13569 64933 13621
rect 64985 13591 71106 13621
rect 64985 13569 65200 13591
rect 64769 13539 65200 13569
rect 65252 13550 71106 13591
rect 65252 13539 65424 13550
rect 64769 13498 65424 13539
rect 65476 13498 71106 13550
rect 64769 13454 71106 13498
rect 64769 13452 65190 13454
rect 64769 13400 64932 13452
rect 64984 13402 65190 13452
rect 65242 13407 71106 13454
rect 65242 13402 65422 13407
rect 64984 13400 65422 13402
rect 64769 13355 65422 13400
rect 65474 13355 71106 13407
rect 64769 13318 71106 13355
rect 64769 13277 65603 13318
rect 64769 13225 64982 13277
rect 65034 13272 65603 13277
rect 65034 13225 65184 13272
rect 64769 13220 65184 13225
rect 65236 13260 65603 13272
rect 65236 13220 65347 13260
rect 64769 13208 65347 13220
rect 65399 13208 65603 13260
rect 64769 13020 65603 13208
rect 62297 11032 65851 11311
rect 61491 9325 62361 9385
rect 61491 9324 61942 9325
rect 61491 9321 61818 9324
rect 61491 9265 61582 9321
rect 61638 9265 61701 9321
rect 61757 9268 61818 9321
rect 61874 9269 61942 9324
rect 61998 9324 62361 9325
rect 61998 9269 62059 9324
rect 61874 9268 62059 9269
rect 62115 9268 62361 9324
rect 61757 9265 62361 9268
rect 61491 9211 62361 9265
rect 61491 9207 61943 9211
rect 61491 9205 61823 9207
rect 61491 9149 61582 9205
rect 61638 9149 61700 9205
rect 61756 9151 61823 9205
rect 61879 9155 61943 9207
rect 61999 9204 62361 9211
rect 61999 9155 62061 9204
rect 61879 9154 61944 9155
rect 61996 9154 62061 9155
rect 61879 9151 62061 9154
rect 61756 9149 62061 9151
rect 61491 9148 62061 9149
rect 62117 9148 62361 9204
rect 61491 9099 62361 9148
rect 56775 6803 57334 6920
rect 56775 6797 57017 6803
rect 56775 6745 56834 6797
rect 56886 6751 57017 6797
rect 57069 6751 57204 6803
rect 57256 6751 57334 6803
rect 56886 6745 57334 6751
rect 56775 6641 57334 6745
rect 53695 4664 54568 4724
rect 53695 4663 54146 4664
rect 53695 4660 54022 4663
rect 53695 4604 53786 4660
rect 53842 4604 53905 4660
rect 53961 4607 54022 4660
rect 54078 4608 54146 4663
rect 54202 4663 54568 4664
rect 54202 4608 54263 4663
rect 54078 4607 54263 4608
rect 54319 4607 54568 4663
rect 53961 4604 54568 4607
rect 53695 4550 54568 4604
rect 53695 4546 54147 4550
rect 53695 4544 54027 4546
rect 53695 4488 53786 4544
rect 53842 4488 53904 4544
rect 53960 4490 54027 4544
rect 54083 4494 54147 4546
rect 54203 4543 54568 4550
rect 54203 4494 54265 4543
rect 54083 4493 54148 4494
rect 54200 4493 54265 4494
rect 54083 4490 54265 4493
rect 53960 4488 54265 4490
rect 53695 4487 54265 4488
rect 54321 4487 54568 4543
rect 53695 4412 54568 4487
rect 53695 4319 54344 4412
rect 53701 4315 54344 4319
rect 53701 4314 54194 4315
rect 49747 3896 50102 4178
rect 42506 3824 50102 3896
rect 49747 3823 50102 3824
rect 65572 2224 65851 11032
rect 98848 4723 99160 4739
rect 98848 4667 98889 4723
rect 98945 4717 99160 4723
rect 98945 4667 99064 4717
rect 98848 4661 99064 4667
rect 99120 4661 99160 4717
rect 98848 4568 99160 4661
rect 98848 4564 99065 4568
rect 98848 4508 98887 4564
rect 98943 4512 99065 4564
rect 99121 4512 99160 4568
rect 98943 4508 99160 4512
rect 98848 4399 99160 4508
rect 98848 4343 98890 4399
rect 98946 4394 99160 4399
rect 98946 4343 99078 4394
rect 98848 4338 99078 4343
rect 99134 4338 99160 4394
rect 91327 4257 92059 4316
rect 98848 4305 99160 4338
rect 91327 4256 91778 4257
rect 91327 4253 91654 4256
rect 91327 4197 91418 4253
rect 91474 4197 91537 4253
rect 91593 4200 91654 4253
rect 91710 4201 91778 4256
rect 91834 4256 92059 4257
rect 91834 4201 91895 4256
rect 91710 4200 91895 4201
rect 91951 4200 92059 4256
rect 91593 4197 92059 4200
rect 91327 4143 92059 4197
rect 91327 4139 91779 4143
rect 91327 4137 91659 4139
rect 91327 4081 91418 4137
rect 91474 4081 91536 4137
rect 91592 4083 91659 4137
rect 91715 4087 91779 4139
rect 91835 4136 92059 4143
rect 91835 4087 91897 4136
rect 91715 4086 91780 4087
rect 91832 4086 91897 4087
rect 91715 4083 91897 4086
rect 91592 4081 91897 4083
rect 91327 4080 91897 4081
rect 91953 4080 92059 4136
rect 91327 4051 92059 4080
rect 95089 2785 95620 2970
rect 95089 2666 96818 2785
rect 95089 2614 95236 2666
rect 95288 2614 95356 2666
rect 95408 2614 95476 2666
rect 95528 2614 96818 2666
rect 95089 2546 96818 2614
rect 95089 2494 95236 2546
rect 95288 2494 95356 2546
rect 95408 2494 95476 2546
rect 95528 2494 96818 2546
rect 95089 2426 96818 2494
rect 95089 2374 95236 2426
rect 95288 2374 95356 2426
rect 95408 2374 95476 2426
rect 95528 2390 96818 2426
rect 95528 2374 95620 2390
rect 95089 2270 95620 2374
rect 56852 2107 65851 2224
rect 56852 2101 57094 2107
rect 56852 2049 56911 2101
rect 56963 2055 57094 2101
rect 57146 2055 57281 2107
rect 57333 2055 65851 2107
rect 56963 2049 65851 2055
rect 56852 1945 65851 2049
rect 94369 368 94922 651
rect 60575 -221 61286 -72
rect 60575 -245 60991 -221
rect 60575 -297 60715 -245
rect 60767 -273 60991 -245
rect 61043 -273 61286 -221
rect 60767 -279 61286 -273
rect 89820 -271 90211 -212
rect 89820 -274 90095 -271
rect 86535 -278 90095 -274
rect 60767 -297 74020 -279
rect 60575 -480 74020 -297
rect 60575 -483 61143 -480
rect 60575 -535 60677 -483
rect 60729 -484 61143 -483
rect 60729 -535 60900 -484
rect 60575 -536 60900 -535
rect 60952 -532 61143 -484
rect 61195 -532 74020 -480
rect 86535 -330 89881 -278
rect 89933 -323 90095 -278
rect 90147 -323 90211 -271
rect 89933 -330 90211 -323
rect 86535 -472 90211 -330
rect 86535 -505 89878 -472
rect 60952 -536 74020 -532
rect 60575 -541 74020 -536
rect 89820 -524 89878 -505
rect 89930 -524 90086 -472
rect 90138 -524 90211 -472
rect 60575 -608 61286 -541
rect 89820 -564 90211 -524
rect 22309 -3123 47333 -2588
rect 13467 -3705 17126 -3380
rect 17805 -3874 17987 -3316
rect 4928 -3961 5298 -3919
rect 4928 -3974 5142 -3961
rect 4928 -4030 4976 -3974
rect 5032 -4017 5142 -3974
rect 5198 -4017 5298 -3961
rect 5032 -4030 5298 -4017
rect 4928 -4101 5298 -4030
rect 11285 -4056 17987 -3874
rect 11296 -4081 17960 -4056
rect 4928 -4112 5147 -4101
rect 4928 -4168 4976 -4112
rect 5032 -4157 5147 -4112
rect 5203 -4157 5298 -4101
rect 5032 -4168 5298 -4157
rect 4928 -4197 5298 -4168
rect 5033 -4504 5403 -4462
rect 5033 -4517 5247 -4504
rect 5033 -4573 5081 -4517
rect 5137 -4560 5247 -4517
rect 5303 -4560 5403 -4504
rect 5137 -4573 5403 -4560
rect 5033 -4644 5403 -4573
rect 5033 -4655 5252 -4644
rect 5033 -4711 5081 -4655
rect 5137 -4700 5252 -4655
rect 5308 -4700 5403 -4644
rect 5137 -4711 5403 -4700
rect 5033 -4740 5403 -4711
rect 46962 -5017 47332 -3123
rect 87090 -4722 87760 -4550
rect 87090 -4778 87132 -4722
rect 87188 -4778 87252 -4722
rect 87308 -4778 87372 -4722
rect 87428 -4778 87760 -4722
rect 87090 -4842 87760 -4778
rect 87090 -4898 87132 -4842
rect 87188 -4898 87252 -4842
rect 87308 -4898 87372 -4842
rect 87428 -4898 87760 -4842
rect 87090 -4962 87760 -4898
rect 45298 -5387 48300 -5017
rect 87090 -5018 87134 -4962
rect 87190 -5018 87252 -4962
rect 87308 -5018 87372 -4962
rect 87428 -5018 87760 -4962
rect 87090 -5090 87760 -5018
rect 47930 -9293 48300 -5387
rect 94639 -7468 94922 368
rect 96448 -5325 96818 2390
rect 98576 -1962 98937 -1953
rect 98576 -2018 98635 -1962
rect 98691 -1963 98937 -1962
rect 98691 -2018 98809 -1963
rect 98576 -2019 98809 -2018
rect 98865 -2019 98937 -1963
rect 98576 -2128 98937 -2019
rect 98576 -2184 98636 -2128
rect 98692 -2133 98937 -2128
rect 98692 -2184 98834 -2133
rect 98576 -2189 98834 -2184
rect 98890 -2189 98937 -2133
rect 98576 -2221 98937 -2189
rect 98546 -2859 98907 -2850
rect 98546 -2915 98605 -2859
rect 98661 -2860 98907 -2859
rect 98661 -2915 98779 -2860
rect 98546 -2916 98779 -2915
rect 98835 -2916 98907 -2860
rect 98546 -3025 98907 -2916
rect 98546 -3081 98606 -3025
rect 98662 -3030 98907 -3025
rect 98662 -3081 98804 -3030
rect 98546 -3086 98804 -3081
rect 98860 -3086 98907 -3030
rect 98546 -3118 98907 -3086
rect 98538 -3342 98899 -3333
rect 98538 -3398 98597 -3342
rect 98653 -3343 98899 -3342
rect 98653 -3398 98771 -3343
rect 98538 -3399 98771 -3398
rect 98827 -3399 98899 -3343
rect 98538 -3508 98899 -3399
rect 98538 -3564 98598 -3508
rect 98654 -3513 98899 -3508
rect 98654 -3564 98796 -3513
rect 98538 -3569 98796 -3564
rect 98852 -3569 98899 -3513
rect 98538 -3601 98899 -3569
rect 98576 -3894 98937 -3885
rect 98576 -3950 98635 -3894
rect 98691 -3895 98937 -3894
rect 98691 -3950 98809 -3895
rect 98576 -3951 98809 -3950
rect 98865 -3951 98937 -3895
rect 98576 -4060 98937 -3951
rect 98576 -4116 98636 -4060
rect 98692 -4065 98937 -4060
rect 98692 -4116 98834 -4065
rect 98576 -4121 98834 -4116
rect 98890 -4121 98937 -4065
rect 98576 -4153 98937 -4121
rect 98574 -7468 98910 -7460
rect 94639 -7474 98910 -7468
rect 94639 -7526 98606 -7474
rect 98658 -7526 98726 -7474
rect 98778 -7526 98846 -7474
rect 98898 -7526 98910 -7474
rect 94639 -7594 98910 -7526
rect 94639 -7646 98606 -7594
rect 98658 -7646 98726 -7594
rect 98778 -7646 98846 -7594
rect 98898 -7646 98910 -7594
rect 94639 -7714 98910 -7646
rect 94639 -7751 98606 -7714
rect 98574 -7766 98606 -7751
rect 98658 -7766 98726 -7714
rect 98778 -7766 98846 -7714
rect 98898 -7766 98910 -7714
rect 98574 -7800 98910 -7766
rect 47930 -9341 48775 -9293
rect 47930 -9393 48446 -9341
rect 48498 -9353 48775 -9341
rect 48498 -9393 48585 -9353
rect 47930 -9405 48585 -9393
rect 48637 -9405 48775 -9353
rect 47930 -9457 48775 -9405
rect 47930 -9509 48440 -9457
rect 48492 -9478 48775 -9457
rect 48492 -9509 48588 -9478
rect 47930 -9530 48588 -9509
rect 48640 -9530 48775 -9478
rect 47930 -9571 48775 -9530
rect 47930 -9623 48443 -9571
rect 48495 -9594 48775 -9571
rect 48495 -9623 48588 -9594
rect 47930 -9646 48588 -9623
rect 48640 -9646 48775 -9594
rect 47930 -9663 48775 -9646
rect 52279 -11322 53565 -11166
rect 52279 -11366 53571 -11322
rect 52279 -11369 53317 -11366
rect 52279 -11377 53075 -11369
rect 52279 -11379 52806 -11377
rect 52279 -11392 52551 -11379
rect 52279 -11448 52346 -11392
rect 52402 -11435 52551 -11392
rect 52607 -11433 52806 -11379
rect 52862 -11425 53075 -11377
rect 53131 -11422 53317 -11369
rect 53373 -11422 53571 -11366
rect 53131 -11425 53571 -11422
rect 52862 -11433 53571 -11425
rect 52607 -11435 53571 -11433
rect 52402 -11448 53571 -11435
rect 52279 -11548 53571 -11448
rect 52279 -11549 53404 -11548
rect 52279 -11561 53245 -11549
rect 52279 -11564 53032 -11561
rect 52279 -11574 52787 -11564
rect 52279 -11582 52554 -11574
rect 52279 -11638 52348 -11582
rect 52404 -11630 52554 -11582
rect 52610 -11620 52787 -11574
rect 52843 -11617 53032 -11564
rect 53088 -11605 53245 -11561
rect 53301 -11604 53404 -11549
rect 53460 -11604 53571 -11548
rect 53301 -11605 53571 -11604
rect 53088 -11617 53571 -11605
rect 52843 -11620 53571 -11617
rect 52610 -11630 53571 -11620
rect 52404 -11638 53571 -11630
rect 52279 -11734 53571 -11638
rect 52279 -11742 53353 -11734
rect 52279 -11752 53155 -11742
rect 52279 -11755 52916 -11752
rect 52279 -11757 52705 -11755
rect 52279 -11758 52507 -11757
rect 52279 -11814 52339 -11758
rect 52395 -11813 52507 -11758
rect 52563 -11811 52705 -11757
rect 52761 -11808 52916 -11755
rect 52972 -11798 53155 -11752
rect 53211 -11790 53353 -11742
rect 53409 -11790 53571 -11734
rect 53211 -11798 53571 -11790
rect 52972 -11808 53571 -11798
rect 52761 -11811 53571 -11808
rect 52563 -11813 53571 -11811
rect 52395 -11814 53571 -11813
rect 52279 -11848 53571 -11814
rect 48991 -14156 49554 -14074
rect 48991 -14208 49199 -14156
rect 49251 -14208 49319 -14156
rect 49371 -14208 49439 -14156
rect 49491 -14208 49554 -14156
rect 48991 -14276 49554 -14208
rect 48991 -14328 49199 -14276
rect 49251 -14328 49319 -14276
rect 49371 -14328 49439 -14276
rect 49491 -14328 49554 -14276
rect 48991 -14450 49554 -14328
<< via2 >>
rect -2671 52726 -2615 52728
rect -2671 52674 -2669 52726
rect -2669 52674 -2617 52726
rect -2617 52674 -2615 52726
rect -2671 52672 -2615 52674
rect -2507 52724 -2451 52726
rect -2507 52672 -2505 52724
rect -2505 52672 -2453 52724
rect -2453 52672 -2451 52724
rect -2507 52670 -2451 52672
rect -2505 52612 -2449 52614
rect -2671 52599 -2615 52601
rect -2671 52547 -2669 52599
rect -2669 52547 -2617 52599
rect -2617 52547 -2615 52599
rect -2505 52560 -2503 52612
rect -2503 52560 -2451 52612
rect -2451 52560 -2449 52612
rect -2505 52558 -2449 52560
rect -2671 52545 -2615 52547
rect -2500 52472 -2444 52474
rect -2671 52461 -2615 52463
rect -2671 52409 -2669 52461
rect -2669 52409 -2617 52461
rect -2617 52409 -2615 52461
rect -2500 52420 -2498 52472
rect -2498 52420 -2446 52472
rect -2446 52420 -2444 52472
rect -2500 52418 -2444 52420
rect -2671 52407 -2615 52409
rect -2361 44200 -2305 44202
rect -2361 44148 -2359 44200
rect -2359 44148 -2307 44200
rect -2307 44148 -2305 44200
rect -2361 44146 -2305 44148
rect -2197 44198 -2141 44200
rect -2197 44146 -2195 44198
rect -2195 44146 -2143 44198
rect -2143 44146 -2141 44198
rect -2197 44144 -2141 44146
rect -2195 44086 -2139 44088
rect -2361 44073 -2305 44075
rect -2361 44021 -2359 44073
rect -2359 44021 -2307 44073
rect -2307 44021 -2305 44073
rect -2195 44034 -2193 44086
rect -2193 44034 -2141 44086
rect -2141 44034 -2139 44086
rect -2195 44032 -2139 44034
rect -2361 44019 -2305 44021
rect -2190 43946 -2134 43948
rect -2361 43935 -2305 43937
rect -2361 43883 -2359 43935
rect -2359 43883 -2307 43935
rect -2307 43883 -2305 43935
rect -2190 43894 -2188 43946
rect -2188 43894 -2136 43946
rect -2136 43894 -2134 43946
rect -2190 43892 -2134 43894
rect -2361 43881 -2305 43883
rect -2354 43659 -2298 43661
rect -2354 43607 -2352 43659
rect -2352 43607 -2300 43659
rect -2300 43607 -2298 43659
rect -2354 43605 -2298 43607
rect -2190 43657 -2134 43659
rect -2190 43605 -2188 43657
rect -2188 43605 -2136 43657
rect -2136 43605 -2134 43657
rect -2190 43603 -2134 43605
rect -2188 43545 -2132 43547
rect -2354 43532 -2298 43534
rect -2354 43480 -2352 43532
rect -2352 43480 -2300 43532
rect -2300 43480 -2298 43532
rect -2188 43493 -2186 43545
rect -2186 43493 -2134 43545
rect -2134 43493 -2132 43545
rect -2188 43491 -2132 43493
rect -2354 43478 -2298 43480
rect -2183 43405 -2127 43407
rect -2354 43394 -2298 43396
rect -2354 43342 -2352 43394
rect -2352 43342 -2300 43394
rect -2300 43342 -2298 43394
rect -2183 43353 -2181 43405
rect -2181 43353 -2129 43405
rect -2129 43353 -2127 43405
rect -2183 43351 -2127 43353
rect -2354 43340 -2298 43342
rect -2462 36766 -2406 36768
rect -2462 36714 -2460 36766
rect -2460 36714 -2408 36766
rect -2408 36714 -2406 36766
rect -2462 36712 -2406 36714
rect -2298 36764 -2242 36766
rect -2298 36712 -2296 36764
rect -2296 36712 -2244 36764
rect -2244 36712 -2242 36764
rect -2298 36710 -2242 36712
rect -2296 36652 -2240 36654
rect -2462 36639 -2406 36641
rect -2462 36587 -2460 36639
rect -2460 36587 -2408 36639
rect -2408 36587 -2406 36639
rect -2296 36600 -2294 36652
rect -2294 36600 -2242 36652
rect -2242 36600 -2240 36652
rect -2296 36598 -2240 36600
rect -2462 36585 -2406 36587
rect -2291 36512 -2235 36514
rect -2462 36501 -2406 36503
rect -2462 36449 -2460 36501
rect -2460 36449 -2408 36501
rect -2408 36449 -2406 36501
rect -2291 36460 -2289 36512
rect -2289 36460 -2237 36512
rect -2237 36460 -2235 36512
rect -2291 36458 -2235 36460
rect -2462 36447 -2406 36449
rect 2607 28025 2663 28027
rect 2041 28017 2097 28019
rect 2041 27965 2043 28017
rect 2043 27965 2095 28017
rect 2095 27965 2097 28017
rect 2417 28017 2473 28019
rect 2041 27963 2097 27965
rect 2220 28014 2276 28016
rect 2220 27962 2222 28014
rect 2222 27962 2274 28014
rect 2274 27962 2276 28014
rect 2417 27965 2419 28017
rect 2419 27965 2471 28017
rect 2471 27965 2473 28017
rect 2607 27973 2609 28025
rect 2609 27973 2661 28025
rect 2661 27973 2663 28025
rect 2607 27971 2663 27973
rect 2417 27963 2473 27965
rect 2220 27960 2276 27962
rect 2044 27890 2100 27892
rect 2044 27838 2046 27890
rect 2046 27838 2098 27890
rect 2098 27838 2100 27890
rect 2607 27890 2663 27892
rect 2409 27882 2465 27884
rect 2044 27836 2100 27838
rect 2220 27879 2276 27881
rect 2220 27827 2222 27879
rect 2222 27827 2274 27879
rect 2274 27827 2276 27879
rect 2409 27830 2411 27882
rect 2411 27830 2463 27882
rect 2463 27830 2465 27882
rect 2607 27838 2609 27890
rect 2609 27838 2661 27890
rect 2661 27838 2663 27890
rect 2607 27836 2663 27838
rect 2409 27828 2465 27830
rect 2220 27825 2276 27827
rect 8765 21701 8821 21757
rect 8980 21721 9036 21777
rect 8654 21538 8710 21594
rect 8916 21548 8972 21604
rect 8672 21287 8728 21343
rect 8892 21297 8948 21353
rect 162 20635 218 20691
rect 377 20655 433 20711
rect 51 20472 107 20528
rect 313 20482 369 20538
rect 69 20221 125 20277
rect 289 20231 345 20287
rect -12465 18806 -12409 18862
rect -12341 18806 -12285 18862
rect -12217 18806 -12161 18862
rect -12093 18806 -12037 18862
rect -10918 18754 -10862 18810
rect -10794 18754 -10738 18810
rect -10670 18754 -10614 18810
rect -10546 18754 -10490 18810
rect -12465 18682 -12409 18738
rect -12341 18682 -12285 18738
rect -12217 18682 -12161 18738
rect -12093 18682 -12037 18738
rect -10918 18630 -10862 18686
rect -10794 18630 -10738 18686
rect -10670 18630 -10614 18686
rect -10546 18630 -10490 18686
rect -12465 18558 -12409 18614
rect -12341 18558 -12285 18614
rect -12217 18558 -12161 18614
rect -12093 18558 -12037 18614
rect -10918 18506 -10862 18562
rect -10794 18506 -10738 18562
rect -10670 18506 -10614 18562
rect -10546 18506 -10490 18562
rect -12465 18434 -12409 18490
rect -12341 18434 -12285 18490
rect -12217 18434 -12161 18490
rect -12093 18434 -12037 18490
rect -10918 18382 -10862 18438
rect -10794 18382 -10738 18438
rect -10670 18382 -10614 18438
rect -10546 18382 -10490 18438
rect 4005 14741 4061 14743
rect 4005 14689 4007 14741
rect 4007 14689 4059 14741
rect 4059 14689 4061 14741
rect 4005 14687 4061 14689
rect 4132 14741 4188 14743
rect 4132 14689 4134 14741
rect 4134 14689 4186 14741
rect 4186 14689 4188 14741
rect 4132 14687 4188 14689
rect -14239 13273 -14183 13275
rect -14239 13221 -14237 13273
rect -14237 13221 -14185 13273
rect -14185 13221 -14183 13273
rect -14239 13219 -14183 13221
rect -14115 13273 -14059 13275
rect -14115 13221 -14113 13273
rect -14113 13221 -14061 13273
rect -14061 13221 -14059 13273
rect -14115 13219 -14059 13221
rect -13991 13273 -13935 13275
rect -13991 13221 -13989 13273
rect -13989 13221 -13937 13273
rect -13937 13221 -13935 13273
rect -13991 13219 -13935 13221
rect -13867 13273 -13811 13275
rect -13867 13221 -13865 13273
rect -13865 13221 -13813 13273
rect -13813 13221 -13811 13273
rect -13209 13234 -13153 13290
rect -13085 13234 -13029 13290
rect -12961 13234 -12905 13290
rect -12837 13234 -12781 13290
rect -13867 13219 -13811 13221
rect -14239 13149 -14183 13151
rect -14239 13097 -14237 13149
rect -14237 13097 -14185 13149
rect -14185 13097 -14183 13149
rect -14239 13095 -14183 13097
rect -14115 13149 -14059 13151
rect -14115 13097 -14113 13149
rect -14113 13097 -14061 13149
rect -14061 13097 -14059 13149
rect -14115 13095 -14059 13097
rect -13991 13149 -13935 13151
rect -13991 13097 -13989 13149
rect -13989 13097 -13937 13149
rect -13937 13097 -13935 13149
rect -13991 13095 -13935 13097
rect -13867 13149 -13811 13151
rect -13867 13097 -13865 13149
rect -13865 13097 -13813 13149
rect -13813 13097 -13811 13149
rect -13209 13110 -13153 13166
rect -13085 13110 -13029 13166
rect -12961 13110 -12905 13166
rect -12837 13110 -12781 13166
rect -13867 13095 -13811 13097
rect -14239 13025 -14183 13027
rect -14239 12973 -14237 13025
rect -14237 12973 -14185 13025
rect -14185 12973 -14183 13025
rect -14239 12971 -14183 12973
rect -14115 13025 -14059 13027
rect -14115 12973 -14113 13025
rect -14113 12973 -14061 13025
rect -14061 12973 -14059 13025
rect -14115 12971 -14059 12973
rect -13991 13025 -13935 13027
rect -13991 12973 -13989 13025
rect -13989 12973 -13937 13025
rect -13937 12973 -13935 13025
rect -13991 12971 -13935 12973
rect -13867 13025 -13811 13027
rect -13867 12973 -13865 13025
rect -13865 12973 -13813 13025
rect -13813 12973 -13811 13025
rect -13209 12986 -13153 13042
rect -13085 12986 -13029 13042
rect -12961 12986 -12905 13042
rect -12837 12986 -12781 13042
rect -13867 12971 -13811 12973
rect -14239 12901 -14183 12903
rect -14239 12849 -14237 12901
rect -14237 12849 -14185 12901
rect -14185 12849 -14183 12901
rect -14239 12847 -14183 12849
rect -14115 12901 -14059 12903
rect -14115 12849 -14113 12901
rect -14113 12849 -14061 12901
rect -14061 12849 -14059 12901
rect -14115 12847 -14059 12849
rect -13991 12901 -13935 12903
rect -13991 12849 -13989 12901
rect -13989 12849 -13937 12901
rect -13937 12849 -13935 12901
rect -13991 12847 -13935 12849
rect -13867 12901 -13811 12903
rect -13867 12849 -13865 12901
rect -13865 12849 -13813 12901
rect -13813 12849 -13811 12901
rect -13209 12862 -13153 12918
rect -13085 12862 -13029 12918
rect -12961 12862 -12905 12918
rect -12837 12862 -12781 12918
rect -13867 12847 -13811 12849
rect 11044 12862 11100 12864
rect 11044 12810 11046 12862
rect 11046 12810 11098 12862
rect 11098 12810 11100 12862
rect 11044 12808 11100 12810
rect 11182 12862 11238 12864
rect 11182 12810 11184 12862
rect 11184 12810 11236 12862
rect 11236 12810 11238 12862
rect 11182 12808 11238 12810
rect 11171 12730 11227 12732
rect 11044 12672 11100 12728
rect 11171 12678 11173 12730
rect 11173 12678 11225 12730
rect 11225 12678 11227 12730
rect 11171 12676 11227 12678
rect 8873 11665 8929 11667
rect 8607 11661 8663 11663
rect 8607 11609 8609 11661
rect 8609 11609 8661 11661
rect 8661 11609 8663 11661
rect 8607 11607 8663 11609
rect 8727 11662 8783 11664
rect 8727 11610 8731 11662
rect 8731 11610 8783 11662
rect 8873 11613 8876 11665
rect 8876 11613 8928 11665
rect 8928 11613 8929 11665
rect 8873 11611 8929 11613
rect 8727 11608 8783 11610
rect 8612 11549 8668 11552
rect 8612 11497 8615 11549
rect 8615 11497 8667 11549
rect 8667 11497 8668 11549
rect 8612 11496 8668 11497
rect 8743 11550 8799 11552
rect 8743 11498 8746 11550
rect 8746 11498 8798 11550
rect 8798 11498 8799 11550
rect 8743 11496 8799 11498
rect 8883 11550 8939 11552
rect 8883 11498 8885 11550
rect 8885 11498 8937 11550
rect 8937 11498 8939 11550
rect 8883 11496 8939 11498
rect 17580 14104 17636 14160
rect 17795 14124 17851 14180
rect 18056 14056 18112 14112
rect 17469 13941 17525 13997
rect 17731 13951 17787 14007
rect 17920 13943 17976 13945
rect 17920 13889 17976 13943
rect 17487 13690 17543 13746
rect 17707 13700 17763 13756
rect 17924 13639 17980 13695
rect 20260 14038 20316 14094
rect 20480 14091 20536 14104
rect 20480 14048 20536 14091
rect 20251 13849 20307 13905
rect 20478 13843 20534 13899
rect 17705 13495 17761 13551
rect -1242 7130 -1186 7186
rect -260 7158 -204 7214
rect 8951 7073 9007 7075
rect 8590 7016 8598 7068
rect 8598 7016 8646 7068
rect 8731 7016 8741 7068
rect 8741 7016 8787 7068
rect 8951 7021 8953 7073
rect 8953 7021 9005 7073
rect 9005 7021 9007 7073
rect 8951 7019 9007 7021
rect 8590 7012 8646 7016
rect 8731 7012 8787 7016
rect 8596 6956 8652 6958
rect 8596 6904 8598 6956
rect 8598 6904 8650 6956
rect 8650 6904 8652 6956
rect 8596 6902 8652 6904
rect 8737 6904 8746 6953
rect 8746 6904 8793 6953
rect 8977 6904 8984 6953
rect 8984 6904 9033 6953
rect 8737 6897 8793 6904
rect 8977 6897 9033 6904
rect -404 6805 -348 6861
rect -989 6668 -933 6724
rect -440 6314 -384 6370
rect -996 6184 -940 6240
rect -1958 1174 -1798 1334
rect -1368 1162 -1208 1322
rect -693 1148 -533 1308
rect -580 101 -420 261
rect 10 89 170 249
rect 685 75 845 235
rect 2725 -259 2781 -257
rect 2725 -311 2727 -259
rect 2727 -311 2779 -259
rect 2779 -311 2781 -259
rect 2725 -313 2781 -311
rect 2889 -261 2945 -259
rect 2889 -313 2891 -261
rect 2891 -313 2943 -261
rect 2943 -313 2945 -261
rect 2889 -315 2945 -313
rect 2891 -373 2947 -371
rect 2725 -386 2781 -384
rect 2725 -438 2727 -386
rect 2727 -438 2779 -386
rect 2779 -438 2781 -386
rect 2891 -425 2893 -373
rect 2893 -425 2945 -373
rect 2945 -425 2947 -373
rect 2891 -427 2947 -425
rect 2725 -440 2781 -438
rect 2896 -513 2952 -511
rect 2725 -524 2781 -522
rect 2725 -576 2727 -524
rect 2727 -576 2779 -524
rect 2779 -576 2781 -524
rect 2896 -565 2898 -513
rect 2898 -565 2950 -513
rect 2950 -565 2952 -513
rect 2896 -567 2952 -565
rect 2725 -578 2781 -576
rect 4826 -990 4882 -988
rect 4826 -1042 4828 -990
rect 4828 -1042 4880 -990
rect 4880 -1042 4882 -990
rect 4826 -1044 4882 -1042
rect 4990 -992 5046 -990
rect 4990 -1044 4992 -992
rect 4992 -1044 5044 -992
rect 5044 -1044 5046 -992
rect 4990 -1046 5046 -1044
rect 4992 -1104 5048 -1102
rect 4826 -1117 4882 -1115
rect 4826 -1169 4828 -1117
rect 4828 -1169 4880 -1117
rect 4880 -1169 4882 -1117
rect 4992 -1156 4994 -1104
rect 4994 -1156 5046 -1104
rect 5046 -1156 5048 -1104
rect 4992 -1158 5048 -1156
rect 4826 -1171 4882 -1169
rect 4997 -1244 5053 -1242
rect 4826 -1255 4882 -1253
rect 4826 -1307 4828 -1255
rect 4828 -1307 4880 -1255
rect 4880 -1307 4882 -1255
rect 4997 -1296 4999 -1244
rect 4999 -1296 5051 -1244
rect 5051 -1296 5053 -1244
rect 4997 -1298 5053 -1296
rect 4826 -1309 4882 -1307
rect 5058 -1556 5114 -1554
rect 4892 -1569 4948 -1567
rect 4892 -1621 4894 -1569
rect 4894 -1621 4946 -1569
rect 4946 -1621 4948 -1569
rect 5058 -1608 5060 -1556
rect 5060 -1608 5112 -1556
rect 5112 -1608 5114 -1556
rect 5058 -1610 5114 -1608
rect 4892 -1623 4948 -1621
rect 5063 -1696 5119 -1694
rect 4892 -1707 4948 -1705
rect 4892 -1759 4894 -1707
rect 4894 -1759 4946 -1707
rect 4946 -1759 4948 -1707
rect 5063 -1748 5065 -1696
rect 5065 -1748 5117 -1696
rect 5117 -1748 5119 -1696
rect 5063 -1750 5119 -1748
rect 4892 -1761 4948 -1759
rect 5215 -2652 5271 -2650
rect 5049 -2665 5105 -2663
rect 5049 -2717 5051 -2665
rect 5051 -2717 5103 -2665
rect 5103 -2717 5105 -2665
rect 5215 -2704 5217 -2652
rect 5217 -2704 5269 -2652
rect 5269 -2704 5271 -2652
rect 5215 -2706 5271 -2704
rect 5049 -2719 5105 -2717
rect 5220 -2792 5276 -2790
rect 5049 -2803 5105 -2801
rect 5049 -2855 5051 -2803
rect 5051 -2855 5103 -2803
rect 5103 -2855 5105 -2803
rect 5220 -2844 5222 -2792
rect 5222 -2844 5274 -2792
rect 5274 -2844 5276 -2792
rect 5220 -2846 5276 -2844
rect 5049 -2857 5105 -2855
rect 5119 -3070 5175 -3068
rect 4953 -3083 5009 -3081
rect 4953 -3135 4955 -3083
rect 4955 -3135 5007 -3083
rect 5007 -3135 5009 -3083
rect 5119 -3122 5121 -3070
rect 5121 -3122 5173 -3070
rect 5173 -3122 5175 -3070
rect 5119 -3124 5175 -3122
rect 4953 -3137 5009 -3135
rect 5124 -3210 5180 -3208
rect 4953 -3221 5009 -3219
rect 4953 -3273 4955 -3221
rect 4955 -3273 5007 -3221
rect 5007 -3273 5009 -3221
rect 5124 -3262 5126 -3210
rect 5126 -3262 5178 -3210
rect 5178 -3262 5180 -3210
rect 5124 -3264 5180 -3262
rect 4953 -3275 5009 -3273
rect 5096 -3484 5152 -3482
rect 4930 -3497 4986 -3495
rect 4930 -3549 4932 -3497
rect 4932 -3549 4984 -3497
rect 4984 -3549 4986 -3497
rect 5096 -3536 5098 -3484
rect 5098 -3536 5150 -3484
rect 5150 -3536 5152 -3484
rect 5096 -3538 5152 -3536
rect 4930 -3551 4986 -3549
rect 5101 -3624 5157 -3622
rect 4930 -3635 4986 -3633
rect 4930 -3687 4932 -3635
rect 4932 -3687 4984 -3635
rect 4984 -3687 4986 -3635
rect 5101 -3676 5103 -3624
rect 5103 -3676 5155 -3624
rect 5155 -3676 5157 -3624
rect 5101 -3678 5157 -3676
rect 4930 -3689 4986 -3687
rect 25520 13562 25576 13618
rect 25708 13562 25764 13618
rect 25903 13562 25959 13618
rect 19668 11188 19724 11190
rect 19668 11136 19670 11188
rect 19670 11136 19722 11188
rect 19722 11136 19724 11188
rect 19668 11134 19724 11136
rect 19909 11193 19965 11195
rect 19909 11141 19911 11193
rect 19911 11141 19963 11193
rect 19963 11141 19965 11193
rect 19909 11139 19965 11141
rect 20148 11195 20204 11197
rect 20148 11143 20150 11195
rect 20150 11143 20202 11195
rect 20202 11143 20204 11195
rect 20148 11141 20204 11143
rect 20375 11195 20431 11197
rect 20375 11143 20377 11195
rect 20377 11143 20429 11195
rect 20429 11143 20431 11195
rect 20375 11141 20431 11143
rect 28782 9893 28838 9895
rect 28782 9841 28784 9893
rect 28784 9841 28836 9893
rect 28836 9841 28838 9893
rect 28782 9839 28838 9841
rect 29023 9898 29079 9900
rect 29023 9846 29025 9898
rect 29025 9846 29077 9898
rect 29077 9846 29079 9898
rect 29023 9844 29079 9846
rect 29262 9900 29318 9902
rect 29262 9848 29264 9900
rect 29264 9848 29316 9900
rect 29316 9848 29318 9900
rect 29262 9846 29318 9848
rect 29489 9900 29545 9902
rect 29489 9848 29491 9900
rect 29491 9848 29543 9900
rect 29543 9848 29545 9900
rect 29489 9846 29545 9848
rect 19626 9142 19682 9144
rect 19626 9090 19628 9142
rect 19628 9090 19680 9142
rect 19680 9090 19682 9142
rect 19626 9088 19682 9090
rect 19867 9147 19923 9149
rect 19867 9095 19869 9147
rect 19869 9095 19921 9147
rect 19921 9095 19923 9147
rect 19867 9093 19923 9095
rect 20106 9149 20162 9151
rect 20106 9097 20108 9149
rect 20108 9097 20160 9149
rect 20160 9097 20162 9149
rect 20106 9095 20162 9097
rect 20333 9149 20389 9151
rect 20333 9097 20335 9149
rect 20335 9097 20387 9149
rect 20387 9097 20389 9149
rect 20333 9095 20389 9097
rect 30535 8963 30591 9019
rect 30667 8976 30723 9032
rect 30792 8975 30848 9031
rect 14587 7905 14643 7961
rect 14803 7905 14859 7961
rect 14589 7782 14645 7838
rect 14803 7777 14859 7833
rect 30532 8850 30588 8906
rect 30665 8866 30721 8922
rect 30792 8866 30848 8922
rect 30529 8737 30585 8793
rect 30654 8739 30710 8795
rect 30792 8739 30848 8795
rect 22937 7874 22993 7876
rect 22937 7822 22939 7874
rect 22939 7822 22991 7874
rect 22991 7822 22993 7874
rect 22937 7820 22993 7822
rect 23178 7879 23234 7881
rect 23178 7827 23180 7879
rect 23180 7827 23232 7879
rect 23232 7827 23234 7879
rect 23178 7825 23234 7827
rect 23417 7881 23473 7883
rect 23417 7829 23419 7881
rect 23419 7829 23471 7881
rect 23471 7829 23473 7881
rect 23417 7827 23473 7829
rect 23644 7881 23700 7883
rect 23644 7829 23646 7881
rect 23646 7829 23698 7881
rect 23698 7829 23700 7881
rect 23644 7827 23700 7829
rect 15167 5993 15327 6153
rect 28726 6899 28782 6901
rect 28726 6847 28728 6899
rect 28728 6847 28780 6899
rect 28780 6847 28782 6899
rect 28726 6845 28782 6847
rect 28967 6904 29023 6906
rect 28967 6852 28969 6904
rect 28969 6852 29021 6904
rect 29021 6852 29023 6904
rect 28967 6850 29023 6852
rect 29206 6906 29262 6908
rect 29206 6854 29208 6906
rect 29208 6854 29260 6906
rect 29260 6854 29262 6906
rect 29206 6852 29262 6854
rect 29433 6906 29489 6908
rect 29433 6854 29435 6906
rect 29435 6854 29487 6906
rect 29487 6854 29489 6906
rect 29433 6852 29489 6854
rect 18890 6014 18946 6016
rect 18230 6011 18286 6013
rect 18230 5959 18232 6011
rect 18232 5959 18284 6011
rect 18284 5959 18286 6011
rect 18230 5957 18286 5959
rect 18408 6009 18464 6011
rect 18408 5957 18410 6009
rect 18410 5957 18462 6009
rect 18462 5957 18464 6009
rect 18408 5955 18464 5957
rect 18649 6008 18705 6010
rect 18649 5956 18651 6008
rect 18651 5956 18703 6008
rect 18703 5956 18705 6008
rect 18890 5962 18892 6014
rect 18892 5962 18944 6014
rect 18944 5962 18946 6014
rect 18890 5960 18946 5962
rect 18649 5954 18705 5956
rect 15167 5284 15327 5444
rect 15167 4472 15327 4632
rect 18331 -830 18387 -774
rect 18536 -991 18592 -935
rect 18795 -972 18851 -916
rect 18706 -1534 18762 -1531
rect 18143 -1546 18199 -1544
rect 18143 -1598 18145 -1546
rect 18145 -1598 18197 -1546
rect 18197 -1598 18199 -1546
rect 18143 -1600 18199 -1598
rect 18452 -1593 18504 -1544
rect 18504 -1593 18508 -1544
rect 18706 -1586 18754 -1534
rect 18754 -1586 18762 -1534
rect 18706 -1587 18762 -1586
rect 18452 -1600 18508 -1593
rect 43283 7104 43443 7106
rect 43283 6948 43285 7104
rect 43285 6948 43441 7104
rect 43441 6948 43443 7104
rect 43283 6946 43443 6948
rect 43826 7104 43986 7106
rect 43826 6948 43828 7104
rect 43828 6948 43984 7104
rect 43984 6948 43986 7104
rect 43826 6946 43986 6948
rect 44536 7104 44696 7106
rect 44536 6948 44538 7104
rect 44538 6948 44694 7104
rect 44694 6948 44696 7104
rect 44536 6946 44696 6948
rect 46935 7078 46991 7080
rect 46193 7073 46249 7075
rect 46193 7021 46195 7073
rect 46195 7021 46247 7073
rect 46247 7021 46249 7073
rect 46719 7070 46775 7072
rect 46193 7019 46249 7021
rect 46439 7068 46495 7070
rect 46439 7016 46441 7068
rect 46441 7016 46493 7068
rect 46493 7016 46495 7068
rect 46719 7018 46721 7070
rect 46721 7018 46773 7070
rect 46773 7018 46775 7070
rect 46935 7026 46937 7078
rect 46937 7026 46989 7078
rect 46989 7026 46991 7078
rect 46935 7024 46991 7026
rect 46719 7016 46775 7018
rect 46439 7014 46495 7016
rect 38310 6450 38470 6610
rect 43823 6074 43879 6076
rect 43823 6022 43825 6074
rect 43825 6022 43877 6074
rect 43877 6022 43879 6074
rect 43823 6020 43879 6022
rect 44072 6061 44128 6063
rect 44072 6009 44074 6061
rect 44074 6009 44126 6061
rect 44126 6009 44128 6061
rect 44528 6060 44584 6062
rect 44072 6007 44128 6009
rect 44306 6056 44362 6058
rect 44306 6004 44308 6056
rect 44308 6004 44360 6056
rect 44360 6004 44362 6056
rect 44528 6008 44530 6060
rect 44530 6008 44582 6060
rect 44582 6008 44584 6060
rect 44528 6006 44584 6008
rect 44306 6002 44362 6004
rect 27147 4405 27203 4407
rect 27147 4353 27149 4405
rect 27149 4353 27201 4405
rect 27201 4353 27203 4405
rect 27147 4351 27203 4353
rect 27379 4405 27435 4407
rect 27379 4353 27381 4405
rect 27381 4353 27433 4405
rect 27433 4353 27435 4405
rect 27379 4351 27435 4353
rect 27144 4209 27200 4211
rect 27144 4157 27146 4209
rect 27146 4157 27198 4209
rect 27198 4157 27200 4209
rect 27144 4155 27200 4157
rect 27379 4209 27435 4211
rect 27379 4157 27381 4209
rect 27381 4157 27433 4209
rect 27433 4157 27435 4209
rect 27379 4155 27435 4157
rect 30468 4487 30524 4489
rect 30468 4435 30470 4487
rect 30470 4435 30522 4487
rect 30522 4435 30524 4487
rect 30468 4433 30524 4435
rect 30468 4226 30524 4228
rect 30468 4174 30470 4226
rect 30470 4174 30522 4226
rect 30522 4174 30524 4226
rect 30468 4172 30524 4174
rect 54248 9315 54304 9317
rect 54012 9262 54014 9314
rect 54014 9262 54066 9314
rect 54066 9262 54068 9314
rect 54012 9258 54068 9262
rect 54131 9262 54133 9314
rect 54133 9262 54185 9314
rect 54185 9262 54187 9314
rect 54131 9258 54187 9262
rect 54248 9263 54252 9315
rect 54252 9263 54304 9315
rect 54248 9261 54304 9263
rect 54372 9316 54428 9318
rect 54372 9264 54374 9316
rect 54374 9264 54426 9316
rect 54426 9264 54428 9316
rect 54372 9262 54428 9264
rect 54489 9315 54545 9317
rect 54489 9263 54492 9315
rect 54492 9263 54544 9315
rect 54544 9263 54545 9315
rect 54489 9261 54545 9263
rect 54012 9196 54068 9198
rect 54012 9144 54014 9196
rect 54014 9144 54066 9196
rect 54066 9144 54068 9196
rect 54012 9142 54068 9144
rect 54130 9196 54186 9198
rect 54130 9144 54133 9196
rect 54133 9144 54185 9196
rect 54185 9144 54186 9196
rect 54253 9197 54309 9200
rect 54253 9145 54254 9197
rect 54254 9145 54306 9197
rect 54306 9145 54309 9197
rect 54373 9199 54429 9204
rect 54373 9148 54374 9199
rect 54374 9148 54426 9199
rect 54426 9148 54429 9199
rect 54491 9195 54547 9197
rect 54253 9144 54309 9145
rect 54130 9142 54186 9144
rect 54491 9143 54493 9195
rect 54493 9143 54545 9195
rect 54545 9143 54547 9195
rect 54491 9141 54547 9143
rect 61818 9322 61874 9324
rect 61582 9269 61584 9321
rect 61584 9269 61636 9321
rect 61636 9269 61638 9321
rect 61582 9265 61638 9269
rect 61701 9269 61703 9321
rect 61703 9269 61755 9321
rect 61755 9269 61757 9321
rect 61701 9265 61757 9269
rect 61818 9270 61822 9322
rect 61822 9270 61874 9322
rect 61818 9268 61874 9270
rect 61942 9323 61998 9325
rect 61942 9271 61944 9323
rect 61944 9271 61996 9323
rect 61996 9271 61998 9323
rect 61942 9269 61998 9271
rect 62059 9322 62115 9324
rect 62059 9270 62062 9322
rect 62062 9270 62114 9322
rect 62114 9270 62115 9322
rect 62059 9268 62115 9270
rect 61582 9203 61638 9205
rect 61582 9151 61584 9203
rect 61584 9151 61636 9203
rect 61636 9151 61638 9203
rect 61582 9149 61638 9151
rect 61700 9203 61756 9205
rect 61700 9151 61703 9203
rect 61703 9151 61755 9203
rect 61755 9151 61756 9203
rect 61823 9204 61879 9207
rect 61823 9152 61824 9204
rect 61824 9152 61876 9204
rect 61876 9152 61879 9204
rect 61943 9206 61999 9211
rect 61943 9155 61944 9206
rect 61944 9155 61996 9206
rect 61996 9155 61999 9206
rect 62061 9202 62117 9204
rect 61823 9151 61879 9152
rect 61700 9149 61756 9151
rect 62061 9150 62063 9202
rect 62063 9150 62115 9202
rect 62115 9150 62117 9202
rect 62061 9148 62117 9150
rect 54022 4661 54078 4663
rect 53786 4608 53788 4660
rect 53788 4608 53840 4660
rect 53840 4608 53842 4660
rect 53786 4604 53842 4608
rect 53905 4608 53907 4660
rect 53907 4608 53959 4660
rect 53959 4608 53961 4660
rect 53905 4604 53961 4608
rect 54022 4609 54026 4661
rect 54026 4609 54078 4661
rect 54022 4607 54078 4609
rect 54146 4662 54202 4664
rect 54146 4610 54148 4662
rect 54148 4610 54200 4662
rect 54200 4610 54202 4662
rect 54146 4608 54202 4610
rect 54263 4661 54319 4663
rect 54263 4609 54266 4661
rect 54266 4609 54318 4661
rect 54318 4609 54319 4661
rect 54263 4607 54319 4609
rect 53786 4542 53842 4544
rect 53786 4490 53788 4542
rect 53788 4490 53840 4542
rect 53840 4490 53842 4542
rect 53786 4488 53842 4490
rect 53904 4542 53960 4544
rect 53904 4490 53907 4542
rect 53907 4490 53959 4542
rect 53959 4490 53960 4542
rect 54027 4543 54083 4546
rect 54027 4491 54028 4543
rect 54028 4491 54080 4543
rect 54080 4491 54083 4543
rect 54147 4545 54203 4550
rect 54147 4494 54148 4545
rect 54148 4494 54200 4545
rect 54200 4494 54203 4545
rect 54265 4541 54321 4543
rect 54027 4490 54083 4491
rect 53904 4488 53960 4490
rect 54265 4489 54267 4541
rect 54267 4489 54319 4541
rect 54319 4489 54321 4541
rect 54265 4487 54321 4489
rect 98889 4719 98945 4723
rect 98889 4667 98941 4719
rect 98941 4667 98945 4719
rect 99064 4713 99120 4717
rect 99064 4661 99116 4713
rect 99116 4661 99120 4713
rect 99065 4564 99121 4568
rect 98887 4560 98943 4564
rect 98887 4508 98939 4560
rect 98939 4508 98943 4560
rect 99065 4512 99117 4564
rect 99117 4512 99121 4564
rect 98890 4395 98946 4399
rect 98890 4343 98942 4395
rect 98942 4343 98946 4395
rect 99078 4390 99134 4394
rect 99078 4338 99130 4390
rect 99130 4338 99134 4390
rect 91654 4254 91710 4256
rect 91418 4201 91420 4253
rect 91420 4201 91472 4253
rect 91472 4201 91474 4253
rect 91418 4197 91474 4201
rect 91537 4201 91539 4253
rect 91539 4201 91591 4253
rect 91591 4201 91593 4253
rect 91537 4197 91593 4201
rect 91654 4202 91658 4254
rect 91658 4202 91710 4254
rect 91654 4200 91710 4202
rect 91778 4255 91834 4257
rect 91778 4203 91780 4255
rect 91780 4203 91832 4255
rect 91832 4203 91834 4255
rect 91778 4201 91834 4203
rect 91895 4254 91951 4256
rect 91895 4202 91898 4254
rect 91898 4202 91950 4254
rect 91950 4202 91951 4254
rect 91895 4200 91951 4202
rect 91418 4135 91474 4137
rect 91418 4083 91420 4135
rect 91420 4083 91472 4135
rect 91472 4083 91474 4135
rect 91418 4081 91474 4083
rect 91536 4135 91592 4137
rect 91536 4083 91539 4135
rect 91539 4083 91591 4135
rect 91591 4083 91592 4135
rect 91659 4136 91715 4139
rect 91659 4084 91660 4136
rect 91660 4084 91712 4136
rect 91712 4084 91715 4136
rect 91779 4138 91835 4143
rect 91779 4087 91780 4138
rect 91780 4087 91832 4138
rect 91832 4087 91835 4138
rect 91897 4134 91953 4136
rect 91659 4083 91715 4084
rect 91536 4081 91592 4083
rect 91897 4082 91899 4134
rect 91899 4082 91951 4134
rect 91951 4082 91953 4134
rect 91897 4080 91953 4082
rect 5142 -3963 5198 -3961
rect 4976 -3976 5032 -3974
rect 4976 -4028 4978 -3976
rect 4978 -4028 5030 -3976
rect 5030 -4028 5032 -3976
rect 5142 -4015 5144 -3963
rect 5144 -4015 5196 -3963
rect 5196 -4015 5198 -3963
rect 5142 -4017 5198 -4015
rect 4976 -4030 5032 -4028
rect 5147 -4103 5203 -4101
rect 4976 -4114 5032 -4112
rect 4976 -4166 4978 -4114
rect 4978 -4166 5030 -4114
rect 5030 -4166 5032 -4114
rect 5147 -4155 5149 -4103
rect 5149 -4155 5201 -4103
rect 5201 -4155 5203 -4103
rect 5147 -4157 5203 -4155
rect 4976 -4168 5032 -4166
rect 5247 -4506 5303 -4504
rect 5081 -4519 5137 -4517
rect 5081 -4571 5083 -4519
rect 5083 -4571 5135 -4519
rect 5135 -4571 5137 -4519
rect 5247 -4558 5249 -4506
rect 5249 -4558 5301 -4506
rect 5301 -4558 5303 -4506
rect 5247 -4560 5303 -4558
rect 5081 -4573 5137 -4571
rect 5252 -4646 5308 -4644
rect 5081 -4657 5137 -4655
rect 5081 -4709 5083 -4657
rect 5083 -4709 5135 -4657
rect 5135 -4709 5137 -4657
rect 5252 -4698 5254 -4646
rect 5254 -4698 5306 -4646
rect 5306 -4698 5308 -4646
rect 5252 -4700 5308 -4698
rect 5081 -4711 5137 -4709
rect 87132 -4724 87188 -4722
rect 87132 -4776 87136 -4724
rect 87136 -4776 87188 -4724
rect 87132 -4778 87188 -4776
rect 87252 -4724 87308 -4722
rect 87252 -4776 87256 -4724
rect 87256 -4776 87308 -4724
rect 87252 -4778 87308 -4776
rect 87372 -4724 87428 -4722
rect 87372 -4776 87376 -4724
rect 87376 -4776 87428 -4724
rect 87372 -4778 87428 -4776
rect 87132 -4844 87188 -4842
rect 87132 -4896 87136 -4844
rect 87136 -4896 87188 -4844
rect 87132 -4898 87188 -4896
rect 87252 -4844 87308 -4842
rect 87252 -4896 87256 -4844
rect 87256 -4896 87308 -4844
rect 87252 -4898 87308 -4896
rect 87372 -4844 87428 -4842
rect 87372 -4896 87376 -4844
rect 87376 -4896 87428 -4844
rect 87372 -4898 87428 -4896
rect 87134 -4964 87190 -4962
rect 87134 -5016 87136 -4964
rect 87136 -5016 87188 -4964
rect 87188 -5016 87190 -4964
rect 87134 -5018 87190 -5016
rect 87252 -4964 87308 -4962
rect 87252 -5016 87256 -4964
rect 87256 -5016 87308 -4964
rect 87252 -5018 87308 -5016
rect 87372 -4964 87428 -4962
rect 87372 -5016 87376 -4964
rect 87376 -5016 87428 -4964
rect 87372 -5018 87428 -5016
rect 98635 -1966 98691 -1962
rect 98635 -2018 98687 -1966
rect 98687 -2018 98691 -1966
rect 98809 -1967 98865 -1963
rect 98809 -2019 98861 -1967
rect 98861 -2019 98865 -1967
rect 98636 -2132 98692 -2128
rect 98636 -2184 98688 -2132
rect 98688 -2184 98692 -2132
rect 98834 -2137 98890 -2133
rect 98834 -2189 98886 -2137
rect 98886 -2189 98890 -2137
rect 98605 -2863 98661 -2859
rect 98605 -2915 98657 -2863
rect 98657 -2915 98661 -2863
rect 98779 -2864 98835 -2860
rect 98779 -2916 98831 -2864
rect 98831 -2916 98835 -2864
rect 98606 -3029 98662 -3025
rect 98606 -3081 98658 -3029
rect 98658 -3081 98662 -3029
rect 98804 -3034 98860 -3030
rect 98804 -3086 98856 -3034
rect 98856 -3086 98860 -3034
rect 98597 -3346 98653 -3342
rect 98597 -3398 98649 -3346
rect 98649 -3398 98653 -3346
rect 98771 -3347 98827 -3343
rect 98771 -3399 98823 -3347
rect 98823 -3399 98827 -3347
rect 98598 -3512 98654 -3508
rect 98598 -3564 98650 -3512
rect 98650 -3564 98654 -3512
rect 98796 -3517 98852 -3513
rect 98796 -3569 98848 -3517
rect 98848 -3569 98852 -3517
rect 98635 -3898 98691 -3894
rect 98635 -3950 98687 -3898
rect 98687 -3950 98691 -3898
rect 98809 -3899 98865 -3895
rect 98809 -3951 98861 -3899
rect 98861 -3951 98865 -3899
rect 98636 -4064 98692 -4060
rect 98636 -4116 98688 -4064
rect 98688 -4116 98692 -4064
rect 98834 -4069 98890 -4065
rect 98834 -4121 98886 -4069
rect 98886 -4121 98890 -4069
rect 53317 -11368 53373 -11366
rect 53075 -11371 53131 -11369
rect 52806 -11379 52862 -11377
rect 52551 -11381 52607 -11379
rect 52346 -11394 52402 -11392
rect 52346 -11446 52348 -11394
rect 52348 -11446 52400 -11394
rect 52400 -11446 52402 -11394
rect 52551 -11433 52553 -11381
rect 52553 -11433 52605 -11381
rect 52605 -11433 52607 -11381
rect 52806 -11431 52808 -11379
rect 52808 -11431 52860 -11379
rect 52860 -11431 52862 -11379
rect 53075 -11423 53077 -11371
rect 53077 -11423 53129 -11371
rect 53129 -11423 53131 -11371
rect 53317 -11420 53319 -11368
rect 53319 -11420 53371 -11368
rect 53371 -11420 53373 -11368
rect 53317 -11422 53373 -11420
rect 53075 -11425 53131 -11423
rect 52806 -11433 52862 -11431
rect 52551 -11435 52607 -11433
rect 52346 -11448 52402 -11446
rect 53245 -11551 53301 -11549
rect 53032 -11563 53088 -11561
rect 52787 -11566 52843 -11564
rect 52554 -11576 52610 -11574
rect 52348 -11584 52404 -11582
rect 52348 -11636 52350 -11584
rect 52350 -11636 52402 -11584
rect 52402 -11636 52404 -11584
rect 52554 -11628 52556 -11576
rect 52556 -11628 52608 -11576
rect 52608 -11628 52610 -11576
rect 52787 -11618 52789 -11566
rect 52789 -11618 52841 -11566
rect 52841 -11618 52843 -11566
rect 53032 -11615 53034 -11563
rect 53034 -11615 53086 -11563
rect 53086 -11615 53088 -11563
rect 53245 -11603 53247 -11551
rect 53247 -11603 53299 -11551
rect 53299 -11603 53301 -11551
rect 53245 -11605 53301 -11603
rect 53404 -11550 53460 -11548
rect 53404 -11602 53406 -11550
rect 53406 -11602 53458 -11550
rect 53458 -11602 53460 -11550
rect 53404 -11604 53460 -11602
rect 53032 -11617 53088 -11615
rect 52787 -11620 52843 -11618
rect 52554 -11630 52610 -11628
rect 52348 -11638 52404 -11636
rect 53353 -11736 53409 -11734
rect 53155 -11744 53211 -11742
rect 52916 -11754 52972 -11752
rect 52705 -11757 52761 -11755
rect 52339 -11760 52395 -11758
rect 52339 -11812 52341 -11760
rect 52341 -11812 52393 -11760
rect 52393 -11812 52395 -11760
rect 52339 -11814 52395 -11812
rect 52507 -11759 52563 -11757
rect 52507 -11811 52509 -11759
rect 52509 -11811 52561 -11759
rect 52561 -11811 52563 -11759
rect 52705 -11809 52707 -11757
rect 52707 -11809 52759 -11757
rect 52759 -11809 52761 -11757
rect 52916 -11806 52918 -11754
rect 52918 -11806 52970 -11754
rect 52970 -11806 52972 -11754
rect 53155 -11796 53157 -11744
rect 53157 -11796 53209 -11744
rect 53209 -11796 53211 -11744
rect 53353 -11788 53355 -11736
rect 53355 -11788 53407 -11736
rect 53407 -11788 53409 -11736
rect 53353 -11790 53409 -11788
rect 53155 -11798 53211 -11796
rect 52916 -11808 52972 -11806
rect 52705 -11811 52761 -11809
rect 52507 -11813 52563 -11811
<< metal3 >>
rect -2499 60654 -2287 62719
rect -2499 60442 -1911 60654
rect -2698 52728 -2423 52744
rect -2698 52672 -2671 52728
rect -2615 52726 -2423 52728
rect -2615 52672 -2507 52726
rect -2698 52670 -2507 52672
rect -2451 52670 -2423 52726
rect -2698 52614 -2423 52670
rect -2698 52601 -2505 52614
rect -2698 52545 -2671 52601
rect -2615 52558 -2505 52601
rect -2449 52575 -2423 52614
rect -2449 52558 861 52575
rect -2615 52545 861 52558
rect -2698 52474 861 52545
rect -2698 52463 -2500 52474
rect -2698 52407 -2671 52463
rect -2615 52418 -2500 52463
rect -2444 52418 861 52474
rect -2615 52407 861 52418
rect -2698 52399 861 52407
rect -2698 52394 -2423 52399
rect -2135 50814 -1964 52180
rect -2388 44202 -2113 44218
rect -2388 44146 -2361 44202
rect -2305 44200 -2113 44202
rect -2305 44146 -2197 44200
rect -2388 44144 -2197 44146
rect -2141 44144 -2113 44200
rect -2388 44088 -2113 44144
rect -2388 44075 -2195 44088
rect -2388 44019 -2361 44075
rect -2305 44032 -2195 44075
rect -2139 44032 -2113 44088
rect -2305 44019 -2113 44032
rect -2388 43948 -2113 44019
rect -2388 43937 -2190 43948
rect -2388 43881 -2361 43937
rect -2305 43892 -2190 43937
rect -2134 43933 -2113 43948
rect 1490 43933 1578 44198
rect -2134 43892 1578 43933
rect -2305 43881 1578 43892
rect -2388 43868 1578 43881
rect -2336 43845 1578 43868
rect -2336 43798 -2269 43845
rect 1490 43798 1578 43845
rect -2381 43661 -2106 43677
rect -2381 43605 -2354 43661
rect -2298 43659 -2106 43661
rect -2298 43605 -2190 43659
rect -2381 43603 -2190 43605
rect -2134 43603 -2106 43659
rect -2381 43547 -2106 43603
rect -2381 43534 -2188 43547
rect -2381 43478 -2354 43534
rect -2298 43491 -2188 43534
rect -2132 43491 -2106 43547
rect -2298 43478 -2106 43491
rect -2381 43407 -2106 43478
rect -2381 43396 -2183 43407
rect -2381 43340 -2354 43396
rect -2298 43351 -2183 43396
rect -2127 43351 -2106 43407
rect -2298 43340 -2106 43351
rect -2381 43327 -2106 43340
rect -2489 36768 -2214 36784
rect -2489 36712 -2462 36768
rect -2406 36766 -2214 36768
rect -2406 36712 -2298 36766
rect -2489 36710 -2298 36712
rect -2242 36710 -2214 36766
rect -2489 36654 -2214 36710
rect -2489 36641 -2296 36654
rect -2489 36585 -2462 36641
rect -2406 36598 -2296 36641
rect -2240 36598 -2214 36654
rect -2406 36585 -2214 36598
rect -2489 36514 -2214 36585
rect -2489 36503 -2291 36514
rect -2489 36447 -2462 36503
rect -2406 36458 -2291 36503
rect -2235 36458 -2214 36514
rect -2406 36447 -2214 36458
rect -2489 36434 -2214 36447
rect 6888 32662 7411 33451
rect -4689 32139 7411 32662
rect -15247 18862 -10439 19168
rect -15247 18806 -12465 18862
rect -12409 18806 -12341 18862
rect -12285 18806 -12217 18862
rect -12161 18806 -12093 18862
rect -12037 18858 -10439 18862
rect -4689 18858 -4166 32139
rect 2010 28027 2740 28118
rect 2010 28019 2607 28027
rect 2010 27963 2041 28019
rect 2097 28016 2417 28019
rect 2097 27963 2220 28016
rect 2010 27960 2220 27963
rect 2276 27963 2417 28016
rect 2473 27971 2607 28019
rect 2663 27971 2740 28027
rect 2473 27963 2740 27971
rect 2276 27960 2740 27963
rect 2010 27892 2740 27960
rect 2010 27836 2044 27892
rect 2100 27884 2607 27892
rect 2100 27881 2409 27884
rect 2100 27836 2220 27881
rect 2010 27825 2220 27836
rect 2276 27828 2409 27881
rect 2465 27836 2607 27884
rect 2663 27836 2740 27892
rect 2465 27828 2740 27836
rect 2276 27825 2740 27828
rect 2010 27720 2740 27825
rect 2011 21918 2709 27720
rect 2011 21777 22718 21918
rect 2011 21757 8980 21777
rect 2011 21701 8765 21757
rect 8821 21721 8980 21757
rect 9036 21721 22718 21777
rect 8821 21701 22718 21721
rect 2011 21604 22718 21701
rect 2011 21594 8916 21604
rect 2011 21538 8654 21594
rect 8710 21548 8916 21594
rect 8972 21548 22718 21604
rect 8710 21538 22718 21548
rect 2011 21353 22718 21538
rect 2011 21343 8892 21353
rect 2011 21287 8672 21343
rect 8728 21297 8892 21343
rect 8948 21297 22718 21353
rect 8728 21287 22718 21297
rect 2011 21220 22718 21287
rect -265 20781 1066 20974
rect -265 20711 20745 20781
rect -265 20691 377 20711
rect -265 20635 162 20691
rect 218 20655 377 20691
rect 433 20655 20745 20711
rect 218 20635 20745 20655
rect -265 20538 20745 20635
rect -265 20528 313 20538
rect -265 20472 51 20528
rect 107 20482 313 20528
rect 369 20482 20745 20538
rect 107 20472 20745 20482
rect -265 20287 20745 20472
rect -265 20277 289 20287
rect -265 20221 69 20277
rect 125 20231 289 20277
rect 345 20231 20745 20287
rect 125 20221 20745 20231
rect -265 20107 20745 20221
rect -265 19888 1066 20107
rect -12037 18810 17883 18858
rect -12037 18806 -10918 18810
rect -15247 18754 -10918 18806
rect -10862 18754 -10794 18810
rect -10738 18754 -10670 18810
rect -10614 18754 -10546 18810
rect -10490 18754 17883 18810
rect -15247 18738 17883 18754
rect -15247 18682 -12465 18738
rect -12409 18682 -12341 18738
rect -12285 18682 -12217 18738
rect -12161 18682 -12093 18738
rect -12037 18686 17883 18738
rect -12037 18682 -10918 18686
rect -15247 18630 -10918 18682
rect -10862 18630 -10794 18686
rect -10738 18630 -10670 18686
rect -10614 18630 -10546 18686
rect -10490 18630 17883 18686
rect -15247 18614 17883 18630
rect -15247 18558 -12465 18614
rect -12409 18558 -12341 18614
rect -12285 18558 -12217 18614
rect -12161 18558 -12093 18614
rect -12037 18562 17883 18614
rect -12037 18558 -10918 18562
rect -15247 18506 -10918 18558
rect -10862 18506 -10794 18562
rect -10738 18506 -10670 18562
rect -10614 18506 -10546 18562
rect -10490 18506 17883 18562
rect -15247 18490 17883 18506
rect -15247 18434 -12465 18490
rect -12409 18434 -12341 18490
rect -12285 18434 -12217 18490
rect -12161 18434 -12093 18490
rect -12037 18438 17883 18490
rect -12037 18434 -10918 18438
rect -15247 18382 -10918 18434
rect -10862 18382 -10794 18438
rect -10738 18382 -10670 18438
rect -10614 18382 -10546 18438
rect -10490 18382 17883 18438
rect -15247 18335 17883 18382
rect -15247 16941 -10439 18335
rect 3978 14775 4746 14777
rect 3968 14743 4746 14775
rect 3968 14687 4005 14743
rect 4061 14687 4132 14743
rect 4188 14687 4746 14743
rect 3968 14653 4746 14687
rect 3968 14651 4219 14653
rect -16003 13566 -12360 13755
rect -16003 13290 3454 13566
rect -16003 13275 -13209 13290
rect -16003 13219 -14239 13275
rect -14183 13219 -14115 13275
rect -14059 13219 -13991 13275
rect -13935 13219 -13867 13275
rect -13811 13234 -13209 13275
rect -13153 13234 -13085 13290
rect -13029 13234 -12961 13290
rect -12905 13234 -12837 13290
rect -12781 13266 3454 13290
rect -12781 13234 -12360 13266
rect -13811 13219 -12360 13234
rect -16003 13166 -12360 13219
rect -16003 13151 -13209 13166
rect -16003 13095 -14239 13151
rect -14183 13095 -14115 13151
rect -14059 13095 -13991 13151
rect -13935 13095 -13867 13151
rect -13811 13110 -13209 13151
rect -13153 13110 -13085 13166
rect -13029 13110 -12961 13166
rect -12905 13110 -12837 13166
rect -12781 13110 -12360 13166
rect -13811 13095 -12360 13110
rect -16003 13042 -12360 13095
rect -16003 13027 -13209 13042
rect -16003 12971 -14239 13027
rect -14183 12971 -14115 13027
rect -14059 12971 -13991 13027
rect -13935 12971 -13867 13027
rect -13811 12986 -13209 13027
rect -13153 12986 -13085 13042
rect -13029 12986 -12961 13042
rect -12905 12986 -12837 13042
rect -12781 12986 -12360 13042
rect -13811 12971 -12360 12986
rect -16003 12918 -12360 12971
rect -16003 12903 -13209 12918
rect -16003 12847 -14239 12903
rect -14183 12847 -14115 12903
rect -14059 12847 -13991 12903
rect -13935 12847 -13867 12903
rect -13811 12862 -13209 12903
rect -13153 12862 -13085 12918
rect -13029 12862 -12961 12918
rect -12905 12862 -12837 12918
rect -12781 12862 -12360 12918
rect -13811 12847 -12360 12862
rect -16003 12531 -12360 12847
rect 3190 12470 3419 13266
rect 4622 12876 4746 14653
rect 17360 14316 17883 18335
rect 17360 14180 18261 14316
rect 17360 14160 17795 14180
rect 17360 14104 17580 14160
rect 17636 14124 17795 14160
rect 17851 14124 18261 14180
rect 17636 14112 18261 14124
rect 17636 14104 18056 14112
rect 17360 14056 18056 14104
rect 18112 14056 18261 14112
rect 17360 14007 18261 14056
rect 17360 13997 17731 14007
rect 17360 13941 17469 13997
rect 17525 13951 17731 13997
rect 17787 13951 18261 14007
rect 17525 13945 18261 13951
rect 17525 13941 17920 13945
rect 17360 13889 17920 13941
rect 17976 13889 18261 13945
rect 17360 13756 18261 13889
rect 17360 13746 17707 13756
rect 17360 13690 17487 13746
rect 17543 13700 17707 13746
rect 17763 13700 18261 13756
rect 20071 14104 20745 20107
rect 22020 17766 22718 21220
rect 22020 17741 49711 17766
rect 22020 17109 91956 17741
rect 22020 17094 55075 17109
rect 22020 17068 49711 17094
rect 20071 14094 20480 14104
rect 20071 14038 20260 14094
rect 20316 14048 20480 14094
rect 20536 14048 20745 14104
rect 20316 14038 20745 14048
rect 20071 13905 20745 14038
rect 20071 13849 20251 13905
rect 20307 13899 20745 13905
rect 20307 13849 20478 13899
rect 20071 13843 20478 13849
rect 20534 13843 20745 13899
rect 20071 13708 20745 13843
rect 17543 13695 18261 13700
rect 17543 13690 17924 13695
rect 17360 13639 17924 13690
rect 17980 13639 18261 13695
rect 26035 13671 26139 13672
rect 25430 13657 26202 13671
rect 17360 13551 18261 13639
rect 17360 13495 17705 13551
rect 17761 13495 18261 13551
rect 17360 13289 18261 13495
rect 25426 13618 26202 13657
rect 25426 13562 25520 13618
rect 25576 13562 25708 13618
rect 25764 13562 25903 13618
rect 25959 13562 26202 13618
rect 25426 13428 26202 13562
rect 10999 12876 11286 12914
rect 4622 12864 11286 12876
rect 4622 12808 11044 12864
rect 11100 12808 11182 12864
rect 11238 12808 11286 12864
rect 4622 12752 11286 12808
rect 10999 12732 11286 12752
rect 10999 12728 11171 12732
rect 10999 12672 11044 12728
rect 11100 12676 11171 12728
rect 11227 12676 11286 12732
rect 11100 12672 11286 12676
rect 10999 12626 11286 12672
rect 25973 12470 26202 13428
rect 3190 12241 26202 12470
rect 8578 11667 8996 11732
rect 8578 11664 8873 11667
rect 8578 11663 8727 11664
rect 8578 11607 8607 11663
rect 8663 11608 8727 11663
rect 8783 11611 8873 11664
rect 8929 11611 8996 11667
rect 8783 11608 8996 11611
rect 8663 11607 8996 11608
rect 8578 11552 8996 11607
rect 8578 11496 8612 11552
rect 8668 11496 8743 11552
rect 8799 11496 8883 11552
rect 8939 11496 8996 11552
rect 8578 11488 8996 11496
rect -1513 7214 1298 7366
rect -1513 7186 -260 7214
rect -1513 7130 -1242 7186
rect -1186 7158 -260 7186
rect -204 7158 1298 7214
rect -1186 7130 1298 7158
rect 8648 7137 8897 11488
rect 19634 11244 19861 11247
rect 19622 11197 20513 11244
rect 19622 11195 20148 11197
rect 19622 11190 19909 11195
rect 19622 11134 19668 11190
rect 19724 11139 19909 11190
rect 19965 11141 20148 11195
rect 20204 11141 20375 11197
rect 20431 11141 20513 11197
rect 19965 11139 20513 11141
rect 19724 11134 20513 11139
rect 19622 11090 20513 11134
rect 19634 9198 19861 11090
rect 20286 9198 20513 11090
rect 19580 9187 19979 9198
rect 20206 9187 20513 9198
rect 19580 9151 20513 9187
rect 19580 9149 20106 9151
rect 19580 9144 19867 9149
rect 19580 9088 19626 9144
rect 19682 9093 19867 9144
rect 19923 9095 20106 9149
rect 20162 9095 20333 9151
rect 20389 9095 20513 9151
rect 19923 9093 20513 9095
rect 19682 9088 20513 9093
rect 19580 9044 20513 9088
rect 14286 7961 15062 8019
rect 14286 7905 14587 7961
rect 14643 7905 14803 7961
rect 14859 7905 15062 7961
rect 14286 7838 15062 7905
rect 14286 7782 14589 7838
rect 14645 7833 15062 7838
rect 14645 7782 14803 7833
rect 14286 7777 14803 7782
rect 14859 7777 15062 7833
rect 14286 7720 15062 7777
rect 20286 8003 20513 9044
rect 25973 9080 26202 12241
rect 28727 10002 32041 10065
rect 28718 9902 32041 10002
rect 28718 9900 29262 9902
rect 28718 9895 29023 9900
rect 28718 9839 28782 9895
rect 28838 9844 29023 9895
rect 29079 9846 29262 9900
rect 29318 9846 29489 9902
rect 29545 9846 32041 9902
rect 29079 9844 32041 9846
rect 28838 9839 32041 9844
rect 28718 9814 32041 9839
rect 28718 9777 29681 9814
rect 30509 9080 30918 9085
rect 25973 9032 30918 9080
rect 25973 9019 30667 9032
rect 25973 8963 30535 9019
rect 30591 8976 30667 9019
rect 30723 9031 30918 9032
rect 30723 8976 30792 9031
rect 30591 8975 30792 8976
rect 30848 8975 30918 9031
rect 30591 8963 30918 8975
rect 25973 8922 30918 8963
rect 25973 8906 30665 8922
rect 25973 8851 30532 8906
rect 30355 8850 30532 8851
rect 30588 8866 30665 8906
rect 30721 8866 30792 8922
rect 30848 8866 30918 8922
rect 30588 8850 30918 8866
rect 30355 8795 30918 8850
rect 30355 8793 30654 8795
rect 30355 8737 30529 8793
rect 30585 8739 30654 8793
rect 30710 8739 30792 8795
rect 30848 8739 30918 8795
rect 30585 8737 30918 8739
rect 30355 8672 30918 8737
rect 20286 7955 20641 8003
rect 20286 7883 26699 7955
rect 20286 7881 23417 7883
rect 20286 7876 23178 7881
rect 20286 7820 22937 7876
rect 22993 7825 23178 7876
rect 23234 7827 23417 7881
rect 23473 7827 23644 7883
rect 23700 7827 26699 7883
rect 23234 7825 26699 7827
rect 22993 7820 26699 7825
rect 20286 7728 26699 7820
rect -1513 7062 1298 7130
rect -1513 7006 -700 7062
rect -644 7006 1298 7062
rect -1513 6983 1298 7006
rect -1513 6927 -1287 6983
rect -1231 6927 1298 6983
rect -1513 6861 1298 6927
rect 8560 7075 9108 7137
rect 8560 7068 8951 7075
rect 8560 7012 8590 7068
rect 8646 7012 8731 7068
rect 8787 7019 8951 7068
rect 9007 7019 9108 7075
rect 8787 7012 9108 7019
rect 8560 6958 9108 7012
rect 8560 6902 8596 6958
rect 8652 6953 9108 6958
rect 8652 6902 8737 6953
rect 8560 6897 8737 6902
rect 8793 6897 8977 6953
rect 9033 6897 9108 6953
rect 8560 6879 9108 6897
rect -1513 6805 -404 6861
rect -348 6825 1298 6861
rect -348 6805 -13 6825
rect -1513 6769 -13 6805
rect 43 6769 1298 6825
rect -1513 6724 1298 6769
rect -1513 6668 -989 6724
rect -933 6668 1298 6724
rect -1513 6525 1298 6668
rect -1513 6482 -750 6525
rect -1513 6426 -1301 6482
rect -1245 6469 -750 6482
rect -694 6469 1298 6525
rect -1245 6426 1298 6469
rect -1513 6370 1298 6426
rect -1513 6314 -440 6370
rect -384 6314 1298 6370
rect -1513 6240 1298 6314
rect -1513 6184 -996 6240
rect -940 6203 1298 6240
rect -940 6184 610 6203
rect -1513 6147 610 6184
rect 666 6147 1298 6203
rect -1513 6145 1298 6147
rect -1513 6117 -714 6145
rect -1513 6061 -1319 6117
rect -1263 6089 -714 6117
rect -658 6109 1298 6145
rect -658 6089 -70 6109
rect -1263 6061 -70 6089
rect -1513 6053 -70 6061
rect -14 6053 1298 6109
rect -1513 5811 1298 6053
rect -3741 1435 -447 1445
rect 14286 1435 14585 7720
rect 15019 6153 15419 6265
rect 15019 5993 15167 6153
rect 15327 5993 15419 6153
rect 15019 5444 15419 5993
rect 15019 5284 15167 5444
rect 15327 5284 15419 5444
rect 15019 4632 15419 5284
rect 15019 4472 15167 4632
rect 15327 4472 15419 4632
rect 15019 4270 15419 4472
rect 16013 6016 19210 6142
rect 16013 6013 18890 6016
rect 16013 5957 18230 6013
rect 18286 6011 18890 6013
rect 18286 5957 18408 6011
rect 16013 5955 18408 5957
rect 18464 6010 18890 6011
rect 18464 5955 18649 6010
rect 16013 5954 18649 5955
rect 18705 5960 18890 6010
rect 18946 5960 19210 6016
rect 18705 5954 19210 5960
rect 16013 5893 19210 5954
rect -3741 1334 14585 1435
rect -3741 1174 -1958 1334
rect -1798 1322 14585 1334
rect -1798 1174 -1368 1322
rect -3741 1162 -1368 1174
rect -1208 1308 14585 1322
rect -1208 1162 -693 1308
rect -3741 1148 -693 1162
rect -533 1148 14585 1308
rect -3741 1136 14585 1148
rect -3741 1068 -447 1136
rect -2319 300 931 372
rect -2789 287 931 300
rect 15116 287 15379 4270
rect -2789 261 15379 287
rect -2789 101 -580 261
rect -420 249 15379 261
rect -420 101 10 249
rect -2789 89 10 101
rect 170 235 15379 249
rect 170 89 685 235
rect -2789 75 685 89
rect 845 75 15379 235
rect -2789 24 15379 75
rect -2789 14 931 24
rect -2319 -5 931 14
rect 2197 -257 3075 -188
rect 2197 -313 2725 -257
rect 2781 -259 3075 -257
rect 2781 -313 2889 -259
rect 2197 -315 2889 -313
rect 2945 -298 3075 -259
rect 16013 -298 16262 5893
rect 20318 352 20641 7728
rect 26472 6980 26699 7728
rect 31790 6980 32041 9814
rect 49039 9313 49671 17068
rect 53921 9318 54794 9377
rect 53921 9317 54372 9318
rect 53921 9314 54248 9317
rect 53921 9313 54012 9314
rect 49039 9258 54012 9313
rect 54068 9258 54131 9314
rect 54187 9261 54248 9314
rect 54304 9262 54372 9317
rect 54428 9317 54794 9318
rect 54428 9262 54489 9317
rect 54304 9261 54489 9262
rect 54545 9313 54794 9317
rect 61491 9325 62361 9385
rect 61491 9324 61942 9325
rect 61491 9321 61818 9324
rect 61491 9313 61582 9321
rect 54545 9265 61582 9313
rect 61638 9265 61701 9321
rect 61757 9268 61818 9321
rect 61874 9269 61942 9324
rect 61998 9324 62361 9325
rect 61998 9269 62059 9324
rect 61874 9268 62059 9269
rect 62115 9313 62361 9324
rect 62115 9268 62375 9313
rect 61757 9265 62375 9268
rect 54545 9261 62375 9265
rect 54187 9258 62375 9261
rect 49039 9211 62375 9258
rect 49039 9207 61943 9211
rect 49039 9205 61823 9207
rect 49039 9204 61582 9205
rect 49039 9200 54373 9204
rect 49039 9198 54253 9200
rect 49039 9142 54012 9198
rect 54068 9142 54130 9198
rect 54186 9144 54253 9198
rect 54309 9148 54373 9200
rect 54429 9197 61582 9204
rect 54429 9148 54491 9197
rect 54309 9144 54491 9148
rect 54186 9142 54491 9144
rect 49039 9141 54491 9142
rect 54547 9149 61582 9197
rect 61638 9149 61700 9205
rect 61756 9151 61823 9205
rect 61879 9155 61943 9207
rect 61999 9204 62375 9211
rect 61999 9155 62061 9204
rect 61879 9151 62061 9155
rect 61756 9149 62061 9151
rect 54547 9148 62061 9149
rect 62117 9148 62375 9204
rect 54547 9141 62375 9148
rect 49039 9087 62375 9141
rect 26472 6908 32041 6980
rect 26472 6906 29206 6908
rect 26472 6901 28967 6906
rect 26472 6845 28726 6901
rect 28782 6850 28967 6901
rect 29023 6852 29206 6906
rect 29262 6852 29433 6908
rect 29489 6852 32041 6908
rect 29023 6850 32041 6852
rect 28782 6845 32041 6850
rect 26472 6753 32041 6845
rect 27167 4463 27415 6753
rect 31790 6741 32041 6753
rect 32327 7125 32533 7128
rect 32327 7124 43272 7125
rect 44110 7124 44460 7130
rect 32327 7106 44715 7124
rect 32327 6946 43283 7106
rect 43443 6946 43826 7106
rect 43986 6946 44536 7106
rect 44696 6946 44715 7106
rect 46136 7080 47059 7119
rect 46136 7075 46935 7080
rect 46136 7019 46193 7075
rect 46249 7072 46935 7075
rect 46249 7070 46719 7072
rect 46249 7019 46439 7070
rect 46136 7014 46439 7019
rect 46495 7016 46719 7070
rect 46775 7024 46935 7072
rect 46991 7024 47059 7080
rect 46775 7016 47059 7024
rect 46495 7014 47059 7016
rect 46136 6961 47059 7014
rect 32327 6919 44715 6946
rect 30400 5978 30606 5983
rect 32327 5978 32533 6919
rect 38287 6610 38493 6919
rect 44110 6850 44480 6919
rect 44110 6810 44460 6850
rect 38287 6450 38310 6610
rect 38470 6450 38493 6610
rect 38287 6414 38493 6450
rect 46593 6195 46752 6961
rect 46519 6163 47743 6195
rect 46512 6130 47745 6163
rect 30400 5772 32533 5978
rect 43759 6076 47745 6130
rect 43759 6020 43823 6076
rect 43879 6063 47745 6076
rect 43879 6020 44072 6063
rect 43759 6007 44072 6020
rect 44128 6062 47745 6063
rect 44128 6058 44528 6062
rect 44128 6007 44306 6058
rect 43759 6002 44306 6007
rect 44362 6006 44528 6058
rect 44584 6006 47745 6062
rect 44362 6002 47745 6006
rect 43759 5971 47745 6002
rect 46512 5937 47745 5971
rect 46519 5906 47743 5937
rect 30400 4489 30606 5772
rect 27094 4407 27485 4463
rect 27094 4351 27147 4407
rect 27203 4351 27379 4407
rect 27435 4351 27485 4407
rect 27094 4211 27485 4351
rect 27094 4155 27144 4211
rect 27200 4155 27379 4211
rect 27435 4155 27485 4211
rect 27094 4108 27485 4155
rect 30400 4433 30468 4489
rect 30524 4433 30606 4489
rect 30400 4228 30606 4433
rect 30400 4172 30468 4228
rect 30524 4172 30606 4228
rect 30400 4129 30606 4172
rect 47454 3849 47743 5906
rect 49039 4545 49671 9087
rect 91324 4952 91956 17109
rect 53695 4664 54568 4724
rect 53695 4663 54146 4664
rect 53695 4660 54022 4663
rect 53695 4604 53786 4660
rect 53842 4604 53905 4660
rect 53961 4607 54022 4660
rect 54078 4608 54146 4663
rect 54202 4663 54568 4664
rect 54202 4608 54263 4663
rect 54078 4607 54263 4608
rect 54319 4607 54568 4663
rect 53961 4604 54568 4607
rect 53695 4550 54568 4604
rect 53695 4546 54147 4550
rect 53695 4545 54027 4546
rect 49039 4544 54027 4545
rect 49039 4488 53786 4544
rect 53842 4488 53904 4544
rect 53960 4490 54027 4544
rect 54083 4494 54147 4546
rect 54203 4545 54568 4550
rect 91324 4723 99215 4952
rect 91324 4667 98889 4723
rect 98945 4717 99215 4723
rect 98945 4667 99064 4717
rect 91324 4661 99064 4667
rect 99120 4661 99215 4717
rect 91324 4568 99215 4661
rect 91324 4564 99065 4568
rect 54203 4543 57420 4545
rect 54203 4494 54265 4543
rect 54083 4490 54265 4494
rect 53960 4488 54265 4490
rect 49039 4487 54265 4488
rect 54321 4487 57420 4543
rect 49039 4319 57420 4487
rect 49039 4304 49671 4319
rect 49161 4303 49588 4304
rect 49161 3849 49588 3854
rect 47454 3560 49588 3849
rect 17589 29 20641 352
rect 2945 -315 16262 -298
rect 2197 -371 16262 -315
rect 2197 -384 2891 -371
rect 2197 -440 2725 -384
rect 2781 -427 2891 -384
rect 2947 -427 16262 -371
rect 2781 -440 16262 -427
rect 2197 -511 16262 -440
rect 2197 -522 2896 -511
rect 2197 -578 2725 -522
rect 2781 -567 2896 -522
rect 2952 -547 16262 -511
rect 2952 -567 3075 -547
rect 2781 -578 3075 -567
rect 2197 -634 3075 -578
rect 4778 -988 5148 -932
rect 4778 -1044 4826 -988
rect 4882 -990 5148 -988
rect 4882 -1044 4990 -990
rect 4778 -1046 4990 -1044
rect 5046 -1004 5148 -990
rect 5046 -1046 15958 -1004
rect 4778 -1102 15958 -1046
rect 4778 -1115 4992 -1102
rect 4778 -1171 4826 -1115
rect 4882 -1158 4992 -1115
rect 5048 -1158 15958 -1102
rect 4882 -1171 15958 -1158
rect 4778 -1242 15958 -1171
rect 4778 -1253 4997 -1242
rect 4778 -1309 4826 -1253
rect 4882 -1298 4997 -1253
rect 5053 -1298 15958 -1242
rect 4882 -1309 15958 -1298
rect 4778 -1321 15958 -1309
rect 4778 -1338 5148 -1321
rect 4844 -1554 14921 -1512
rect 4844 -1567 5058 -1554
rect 4844 -1623 4892 -1567
rect 4948 -1610 5058 -1567
rect 5114 -1610 14921 -1554
rect 4948 -1623 14921 -1610
rect 4844 -1694 14921 -1623
rect 4844 -1705 5063 -1694
rect 4844 -1761 4892 -1705
rect 4948 -1750 5063 -1705
rect 5119 -1750 14921 -1694
rect 4948 -1756 14921 -1750
rect 4948 -1761 5222 -1756
rect 4844 -1773 5222 -1761
rect 4844 -1790 5214 -1773
rect 14677 -2260 14921 -1756
rect 15641 -1813 15958 -1321
rect 17649 -1459 17851 29
rect 18284 -774 21310 -725
rect 18284 -830 18331 -774
rect 18387 -830 21310 -774
rect 18284 -916 21310 -830
rect 18284 -935 18795 -916
rect 18284 -991 18536 -935
rect 18592 -972 18795 -935
rect 18851 -972 21310 -916
rect 18592 -991 21310 -972
rect 18284 -1061 21310 -991
rect 20974 -1269 21310 -1061
rect 17649 -1531 18861 -1459
rect 17649 -1544 18706 -1531
rect 17649 -1600 18143 -1544
rect 18199 -1600 18452 -1544
rect 18508 -1587 18706 -1544
rect 18762 -1587 18861 -1531
rect 18508 -1600 18861 -1587
rect 17649 -1661 18861 -1600
rect 20974 -1605 26713 -1269
rect 15641 -2130 25855 -1813
rect 24985 -2260 25196 -2248
rect 14677 -2504 25212 -2260
rect 5001 -2623 5379 -2608
rect 4971 -2650 24848 -2623
rect 4971 -2663 5215 -2650
rect 4971 -2719 5049 -2663
rect 5105 -2706 5215 -2663
rect 5271 -2706 24848 -2650
rect 5105 -2719 24848 -2706
rect 4971 -2774 24848 -2719
rect 5001 -2790 5379 -2774
rect 5001 -2801 5220 -2790
rect 5001 -2857 5049 -2801
rect 5105 -2846 5220 -2801
rect 5276 -2846 5379 -2790
rect 5105 -2857 5379 -2846
rect 5001 -2869 5379 -2857
rect 5001 -2886 5371 -2869
rect 4975 -3026 16639 -2983
rect 4905 -3068 16639 -3026
rect 4905 -3081 5119 -3068
rect 4905 -3137 4953 -3081
rect 5009 -3124 5119 -3081
rect 5175 -3124 16639 -3068
rect 5009 -3137 16639 -3124
rect 4905 -3208 16639 -3137
rect 4905 -3219 5124 -3208
rect 4905 -3275 4953 -3219
rect 5009 -3264 5124 -3219
rect 5180 -3232 16639 -3208
rect 5180 -3264 5283 -3232
rect 5009 -3275 5283 -3264
rect 4905 -3287 5283 -3275
rect 4905 -3304 5275 -3287
rect 4882 -3462 5260 -3440
rect 4882 -3482 16212 -3462
rect 4882 -3495 5096 -3482
rect 4882 -3551 4930 -3495
rect 4986 -3538 5096 -3495
rect 5152 -3538 16212 -3482
rect 4986 -3551 16212 -3538
rect 4882 -3622 16212 -3551
rect 4882 -3633 5101 -3622
rect 4882 -3689 4930 -3633
rect 4986 -3678 5101 -3633
rect 5157 -3643 16212 -3622
rect 5157 -3678 5260 -3643
rect 4986 -3689 5260 -3678
rect 4882 -3701 5260 -3689
rect 4882 -3718 5252 -3701
rect 5001 -3919 7452 -3878
rect 4928 -3961 7452 -3919
rect 4928 -3974 5142 -3961
rect 4928 -4030 4976 -3974
rect 5032 -4017 5142 -3974
rect 5198 -4017 7452 -3961
rect 5032 -4030 7452 -4017
rect 4928 -4101 7452 -4030
rect 4928 -4112 5147 -4101
rect 4928 -4168 4976 -4112
rect 5032 -4157 5147 -4112
rect 5203 -4103 7452 -4101
rect 5203 -4157 5306 -4103
rect 5032 -4168 5306 -4157
rect 4928 -4180 5306 -4168
rect 4928 -4197 5298 -4180
rect 7227 -4372 7452 -4103
rect 5070 -4462 6102 -4418
rect 5033 -4504 6102 -4462
rect 5033 -4517 5247 -4504
rect 5033 -4573 5081 -4517
rect 5137 -4560 5247 -4517
rect 5303 -4560 6102 -4504
rect 5137 -4573 6102 -4560
rect 5033 -4630 6102 -4573
rect 5033 -4644 5411 -4630
rect 5033 -4655 5252 -4644
rect 5033 -4711 5081 -4655
rect 5137 -4700 5252 -4655
rect 5308 -4700 5411 -4644
rect 5137 -4711 5411 -4700
rect 5033 -4723 5411 -4711
rect 5033 -4740 5403 -4723
rect 16031 -5048 16212 -3643
rect 16390 -5174 16639 -3232
rect 24697 -5269 24848 -2774
rect 24985 -5303 25196 -2504
rect 25538 -3786 25855 -2130
rect 26377 -2241 26713 -1605
rect 49161 -1981 49588 3560
rect 57127 213 57420 4319
rect 91324 4508 98887 4564
rect 98943 4512 99065 4564
rect 99121 4512 99215 4568
rect 98943 4508 99215 4512
rect 91324 4399 99215 4508
rect 91324 4343 98890 4399
rect 98946 4394 99215 4399
rect 98946 4343 99078 4394
rect 91324 4338 99078 4343
rect 99134 4338 99215 4394
rect 91324 4320 99215 4338
rect 91324 4257 92059 4320
rect 98838 4305 99160 4320
rect 91324 4256 91778 4257
rect 91324 4253 91654 4256
rect 91324 4197 91418 4253
rect 91474 4197 91537 4253
rect 91593 4200 91654 4253
rect 91710 4201 91778 4256
rect 91834 4256 92059 4257
rect 91834 4201 91895 4256
rect 91710 4200 91895 4201
rect 91951 4200 92059 4256
rect 91593 4197 92059 4200
rect 91324 4143 92059 4197
rect 91324 4139 91779 4143
rect 91324 4137 91659 4139
rect 91324 4081 91418 4137
rect 91474 4081 91536 4137
rect 91592 4083 91659 4137
rect 91715 4087 91779 4139
rect 91835 4136 92059 4143
rect 91835 4087 91897 4136
rect 91715 4083 91897 4087
rect 91592 4081 91897 4083
rect 91324 4080 91897 4081
rect 91953 4080 92059 4136
rect 91324 4051 92059 4080
rect 91324 4026 91956 4051
rect 55465 -151 57420 213
rect 26377 -2577 36376 -2241
rect 49161 -2408 51945 -1981
rect 25538 -4103 32240 -3786
rect 31923 -5255 32240 -4103
rect 36040 -6541 36376 -2577
rect 51518 -4201 51945 -2408
rect 51284 -4246 52067 -4201
rect 51284 -4273 51585 -4246
rect 51284 -4329 51344 -4273
rect 51400 -4302 51585 -4273
rect 51641 -4277 52067 -4246
rect 51641 -4302 51860 -4277
rect 51400 -4329 51860 -4302
rect 51284 -4333 51860 -4329
rect 51916 -4333 52067 -4277
rect 51284 -4396 52067 -4333
rect 51284 -4415 51571 -4396
rect 51284 -4471 51328 -4415
rect 51384 -4452 51571 -4415
rect 51627 -4427 52067 -4396
rect 51627 -4452 51833 -4427
rect 51384 -4471 51833 -4452
rect 51284 -4483 51833 -4471
rect 51889 -4483 52067 -4427
rect 51284 -4573 52067 -4483
rect 51284 -4577 51559 -4573
rect 51284 -4633 51313 -4577
rect 51369 -4629 51559 -4577
rect 51615 -4577 52067 -4573
rect 51615 -4629 51867 -4577
rect 51369 -4633 51867 -4629
rect 51923 -4633 52067 -4577
rect 51284 -4719 52067 -4633
rect 36093 -14454 36324 -6662
rect 52279 -11322 53565 -11166
rect 52279 -11366 53571 -11322
rect 52279 -11369 53317 -11366
rect 52279 -11377 53075 -11369
rect 52279 -11379 52806 -11377
rect 52279 -11392 52551 -11379
rect 52279 -11448 52346 -11392
rect 52402 -11435 52551 -11392
rect 52607 -11433 52806 -11379
rect 52862 -11425 53075 -11377
rect 53131 -11422 53317 -11369
rect 53373 -11422 53571 -11366
rect 53131 -11425 53571 -11422
rect 52862 -11433 53571 -11425
rect 52607 -11435 53571 -11433
rect 52402 -11448 53571 -11435
rect 52279 -11479 53571 -11448
rect 55465 -11479 55829 -151
rect 67147 -1962 98964 -1936
rect 67147 -2018 98635 -1962
rect 98691 -1963 98964 -1962
rect 98691 -2018 98809 -1963
rect 67147 -2019 98809 -2018
rect 98865 -2019 98964 -1963
rect 67147 -2128 98964 -2019
rect 67147 -2184 98636 -2128
rect 98692 -2133 98964 -2128
rect 98692 -2184 98834 -2133
rect 67147 -2189 98834 -2184
rect 98890 -2189 98964 -2133
rect 67147 -2230 98964 -2189
rect 67147 -4968 67396 -2230
rect 98546 -2859 98907 -2850
rect 98546 -2905 98605 -2859
rect 75818 -2915 98605 -2905
rect 98661 -2860 98907 -2859
rect 98661 -2915 98779 -2860
rect 75818 -2916 98779 -2915
rect 98835 -2916 98907 -2860
rect 75818 -3025 98907 -2916
rect 75818 -3081 98606 -3025
rect 98662 -3030 98907 -3025
rect 98662 -3081 98804 -3030
rect 75818 -3086 98804 -3081
rect 98860 -3086 98907 -3030
rect 75818 -3114 98907 -3086
rect 57040 -5286 59498 -5074
rect 75848 -5104 75996 -3114
rect 98546 -3118 98907 -3114
rect 76086 -3342 98994 -3305
rect 76086 -3398 98597 -3342
rect 98653 -3343 98994 -3342
rect 98653 -3398 98771 -3343
rect 76086 -3399 98771 -3398
rect 98827 -3399 98994 -3343
rect 76086 -3508 98994 -3399
rect 76086 -3564 98598 -3508
rect 98654 -3513 98994 -3508
rect 98654 -3564 98796 -3513
rect 76086 -3569 98796 -3564
rect 98852 -3569 98994 -3513
rect 76086 -3614 98994 -3569
rect 67579 -5310 68894 -5139
rect 75883 -5179 75961 -5104
rect 76158 -5181 76323 -3614
rect 98576 -3892 98937 -3885
rect 83093 -3894 99108 -3892
rect 83093 -3950 98635 -3894
rect 98691 -3895 99108 -3894
rect 98691 -3950 98809 -3895
rect 83093 -3951 98809 -3950
rect 98865 -3951 99108 -3895
rect 83093 -4060 99108 -3951
rect 83093 -4116 98636 -4060
rect 98692 -4065 99108 -4060
rect 98692 -4116 98834 -4065
rect 83093 -4121 98834 -4116
rect 98890 -4121 99108 -4065
rect 83093 -4168 99108 -4121
rect 83093 -5156 83369 -4168
rect 87090 -4722 87760 -4550
rect 87090 -4778 87132 -4722
rect 87188 -4778 87252 -4722
rect 87308 -4778 87372 -4722
rect 87428 -4778 87760 -4722
rect 87090 -4842 87760 -4778
rect 87090 -4898 87132 -4842
rect 87188 -4898 87252 -4842
rect 87308 -4898 87372 -4842
rect 87428 -4898 87760 -4842
rect 87090 -4962 87760 -4898
rect 87090 -5018 87134 -4962
rect 87190 -5018 87252 -4962
rect 87308 -5018 87372 -4962
rect 87428 -5018 87760 -4962
rect 87090 -5090 87760 -5018
rect 52279 -11548 55829 -11479
rect 52279 -11549 53404 -11548
rect 52279 -11561 53245 -11549
rect 52279 -11564 53032 -11561
rect 52279 -11574 52787 -11564
rect 52279 -11582 52554 -11574
rect 52279 -11638 52348 -11582
rect 52404 -11630 52554 -11582
rect 52610 -11620 52787 -11574
rect 52843 -11617 53032 -11564
rect 53088 -11605 53245 -11561
rect 53301 -11604 53404 -11549
rect 53460 -11604 55829 -11548
rect 53301 -11605 55829 -11604
rect 53088 -11617 55829 -11605
rect 52843 -11620 55829 -11617
rect 52610 -11630 55829 -11620
rect 52404 -11638 55829 -11630
rect 52279 -11734 55829 -11638
rect 52279 -11742 53353 -11734
rect 52279 -11752 53155 -11742
rect 52279 -11755 52916 -11752
rect 52279 -11757 52705 -11755
rect 52279 -11758 52507 -11757
rect 52279 -11814 52339 -11758
rect 52395 -11813 52507 -11758
rect 52563 -11811 52705 -11757
rect 52761 -11808 52916 -11755
rect 52972 -11798 53155 -11752
rect 53211 -11790 53353 -11742
rect 53409 -11790 55829 -11734
rect 53211 -11798 55829 -11790
rect 52972 -11808 55829 -11798
rect 52761 -11811 55829 -11808
rect 52563 -11813 55829 -11811
rect 52395 -11814 55829 -11813
rect 52279 -11843 55829 -11814
rect 52279 -11848 53571 -11843
rect 87243 -14434 87474 -5992
rect 34855 -14685 36324 -14454
rect 78405 -14665 87474 -14434
<< via3 >>
rect -700 7006 -644 7062
rect -1287 6927 -1231 6983
rect -13 6769 43 6825
rect -1301 6426 -1245 6482
rect -750 6469 -694 6525
rect 610 6147 666 6203
rect -1319 6061 -1263 6117
rect -714 6089 -658 6145
rect -70 6053 -14 6109
rect 51344 -4329 51400 -4273
rect 51585 -4302 51641 -4246
rect 51860 -4333 51916 -4277
rect 51328 -4471 51384 -4415
rect 51571 -4452 51627 -4396
rect 51833 -4483 51889 -4427
rect 51313 -4633 51369 -4577
rect 51559 -4629 51615 -4573
rect 51867 -4633 51923 -4577
<< metal4 >>
rect -7940 41508 -7091 41515
rect -7940 41159 -2689 41508
rect -7940 40575 -2522 41159
rect -7940 -27439 -7091 40575
rect -1377 7366 -914 29105
rect -1513 7062 1298 7366
rect -1513 7006 -700 7062
rect -644 7006 1298 7062
rect -1513 6983 1298 7006
rect -1513 6927 -1287 6983
rect -1231 6927 1298 6983
rect -1513 6825 1298 6927
rect -1513 6769 -13 6825
rect 43 6769 1298 6825
rect -1513 6525 1298 6769
rect -1513 6482 -750 6525
rect -1513 6426 -1301 6482
rect -1245 6469 -750 6482
rect -694 6469 1298 6525
rect -1245 6426 1298 6469
rect -1513 6203 1298 6426
rect -1513 6147 610 6203
rect 666 6147 1298 6203
rect -1513 6145 1298 6147
rect -1513 6117 -714 6145
rect -1513 6061 -1319 6117
rect -1263 6089 -714 6117
rect -658 6109 1298 6145
rect -658 6089 -70 6109
rect -1263 6061 -70 6089
rect -1513 6053 -70 6061
rect -14 6053 1298 6109
rect -1513 5811 1298 6053
rect -1377 -5477 -914 5811
rect 51271 -4204 52095 -4173
rect 27683 -4246 64047 -4204
rect 27683 -4273 51585 -4246
rect 27683 -4329 51344 -4273
rect 51400 -4302 51585 -4273
rect 51641 -4277 64047 -4246
rect 51641 -4302 51860 -4277
rect 51400 -4329 51860 -4302
rect 27683 -4333 51860 -4329
rect 51916 -4333 64047 -4277
rect 27683 -4396 64047 -4333
rect 27683 -4415 51571 -4396
rect 27683 -4471 51328 -4415
rect 51384 -4452 51571 -4415
rect 51627 -4427 64047 -4396
rect 51627 -4452 51833 -4427
rect 51384 -4471 51833 -4452
rect 27683 -4483 51833 -4471
rect 51889 -4483 64047 -4427
rect 27683 -4573 64047 -4483
rect 27683 -4577 51559 -4573
rect 27683 -4633 51313 -4577
rect 51369 -4629 51559 -4577
rect 51615 -4577 64047 -4573
rect 51615 -4629 51867 -4577
rect 51369 -4633 51867 -4629
rect 51923 -4633 64047 -4577
rect 27683 -4710 64047 -4633
rect 27683 -4719 28790 -4710
rect 28900 -4719 29370 -4710
rect 29480 -4719 64047 -4710
rect -1377 -5956 8303 -5477
rect -1377 -8482 -914 -5956
rect 39504 -25347 59472 -24884
rect 11279 -27389 12128 -26499
rect 21483 -27389 22332 -26499
rect 11279 -27439 22332 -27389
rect -7940 -27686 22332 -27439
rect 28864 -27686 29713 -26251
rect 62449 -27498 66334 -26649
rect 62449 -27686 63298 -27498
rect -7940 -28288 63298 -27686
rect 21483 -28535 63298 -28288
rect 65485 -27544 66334 -27498
rect 72203 -27544 73052 -26649
rect 65485 -27594 73052 -27544
rect 80015 -27594 80864 -26550
rect 65485 -28393 80864 -27594
rect 72203 -28443 80864 -28393
<< metal5 >>
rect 95553 96750 98008 97088
rect 97670 -190 98008 96750
rect 85331 -528 98008 -190
use 7b_divider_magic  7b_divider_magic_0
timestamp 1713971633
transform 1 0 57381 0 1 -16876
box -441 -10214 40218 12749
use 7b_divider_magic  7b_divider_magic_1
timestamp 1713971633
transform 0 -1 9619 -1 0 62378
box -441 -10214 40218 12749
use 7b_divider_magic  7b_divider_magic_2
timestamp 1713971633
transform 1 0 6231 0 1 -16896
box -441 -10214 40218 12749
use A_MUX  A_MUX_0
timestamp 1713185578
transform 1 0 42495 0 1 4782
box -285 -452 3979 2227
use A_MUX  A_MUX_1
timestamp 1713185578
transform 1 0 18282 0 -1 12510
box -285 -452 3979 2227
use A_MUX  A_MUX_2
timestamp 1713185578
transform 1 0 18240 0 1 7818
box -285 -452 3979 2227
use A_MUX  A_MUX_3
timestamp 1713185578
transform -1 0 30924 0 -1 11425
box -285 -452 3979 2227
use A_MUX  A_MUX_4
timestamp 1713185578
transform -1 0 30867 0 -1 8419
box -285 -452 3979 2227
use A_MUX  A_MUX_5
timestamp 1713185578
transform 1 0 16712 0 1 -3124
box -285 -452 3979 2227
use A_MUX  A_MUX_6
timestamp 1713185578
transform 1 0 36417 0 -1 12138
box -285 -452 3979 2227
use cap_11p  cap_11p_0
timestamp 1713185578
transform 1 0 94240 0 1 13088
box -26450 -13708 -6739 632
use cap_240p  cap_240p_0
timestamp 1713185578
transform 1 0 89483 0 -1 28277
box -68140 -68970 6839 8429
use CP_1  CP_1_0
timestamp 1713185578
transform 1 0 33105 0 1 10459
box -1133 -1188 2101 1774
use Current_Mirror_Top  Current_Mirror_Top_0
timestamp 1713185578
transform -1 0 2228 0 1 10249
box -1992 -209 4486 7070
use INV_2  INV_2_0
timestamp 1713185578
transform 1 0 11673 0 1 7901
box 21 -485 1081 648
use INV_2  INV_2_1
timestamp 1713185578
transform 1 0 11228 0 1 13239
box 21 -485 1081 648
use PFD_T2  PFD_T2_0
timestamp 1713275964
transform 1 0 22661 0 1 8437
box -28 -113 4062 3793
use RES_74k  RES_74k_0
timestamp 1713358893
transform 1 0 38279 0 1 8429
box 3672 -1154 9606 4970
use Tappered_Buffer  Tappered_Buffer_0
timestamp 1713185578
transform 1 0 50570 0 1 3553
box -161 -3147 5956 944
use Tappered_Buffer  Tappered_Buffer_1
timestamp 1713185578
transform 1 0 50390 0 1 8230
box -161 -3147 5956 944
use Tappered_Buffer  Tappered_Buffer_2
timestamp 1713185578
transform 1 0 58351 0 1 8237
box -161 -3147 5956 944
use Tappered_Buffer  Tappered_Buffer_3
timestamp 1713185578
transform -1 0 94996 0 1 3197
box -161 -3147 5956 944
use Tappered_Buffer  Tappered_Buffer_5
timestamp 1713185578
transform 1 0 48878 0 -1 -10328
box -161 -3147 5956 944
use Tappered_Buffer  Tappered_Buffer_6
timestamp 1713185578
transform -1 0 4941 0 1 26954
box -161 -3147 5956 944
use Tappered_Buffer  Tappered_Buffer_7
timestamp 1713185578
transform -1 0 11108 0 1 10738
box -161 -3147 5956 944
use Tappered_Buffer  Tappered_Buffer_8
timestamp 1713185578
transform -1 0 12287 0 1 6101
box -161 -3147 5956 944
use VCO_DFF_C  VCO_DFF_C_0
timestamp 1713971361
transform 1 0 24282 0 1 -1600
box -90 -27 23932 7176
<< labels >>
flabel metal1 s 1578 15993 1578 15993 0 FreeSans 750 180 0 0 G_source_up
port 1 nsew
flabel metal1 s 1382 15902 1382 15902 0 FreeSans 750 180 0 0 G_source_dn
port 2 nsew
flabel metal1 s 1916 15531 1916 15531 0 FreeSans 750 180 0 0 G_sink_up
port 3 nsew
flabel metal1 s 1919 15268 1919 15268 0 FreeSans 750 180 0 0 G_sink_dn
port 4 nsew
flabel metal1 s 22036 6756 22036 6756 0 FreeSans 2500 0 0 0 S3
port 5 nsew
flabel metal1 s 21788 13207 21788 13207 0 FreeSans 2500 0 0 0 S2
port 6 nsew
flabel metal1 s 19290 14218 19290 14218 0 FreeSans 2500 0 0 0 S1
port 7 nsew
flabel metal1 s 17988 6714 17988 6714 0 FreeSans 2500 0 0 0 S6
port 8 nsew
flabel metal1 s 21995 13993 21995 13993 0 FreeSans 2500 0 0 0 UP_INPUT
port 9 nsew
flabel metal1 s 21858 13590 21858 13590 0 FreeSans 2500 0 0 0 DN_INPUT
port 10 nsew
flabel metal1 s 18022 14399 18022 14399 0 FreeSans 2500 0 0 0 F_IN
port 11 nsew
flabel metal1 s 30024 14122 30024 14122 0 FreeSans 2500 0 0 0 VDD
port 12 nsew
flabel metal1 s 42870 4240 42870 4240 0 FreeSans 2500 0 0 0 VCTRL_IN
port 13 nsew
flabel metal1 s 43370 4280 43370 4280 0 FreeSans 2500 0 0 0 S4
port 14 nsew
flabel metal1 s 26249 11574 26249 11574 0 FreeSans 2500 0 0 0 UP1
port 15 nsew
flabel metal1 s 26214 8908 26214 8908 0 FreeSans 2500 0 0 0 DN1
port 16 nsew
flabel metal1 s 22703 16344 22703 16344 0 FreeSans 2500 0 0 0 LF_OFFCHIP
port 17 nsew
flabel metal1 s 26307 16690 26307 16690 0 FreeSans 2500 0 0 0 S5
port 18 nsew
flabel metal1 s 56568 6749 56568 6749 0 FreeSans 2500 0 0 0 OUTB
port 19 nsew
flabel metal1 s 56817 2078 56817 2078 0 FreeSans 2500 0 0 0 OUT
port 20 nsew
flabel metal1 s 99070 -7610 99070 -7610 0 FreeSans 2500 0 0 0 OUT1
port 21 nsew
flabel metal1 s 99137 -2090 99137 -2090 0 FreeSans 2500 0 0 0 D13
port 22 nsew
flabel metal1 s 99090 -2966 99090 -2966 0 FreeSans 2500 0 0 0 D12
port 23 nsew
flabel metal1 s 99146 -3471 99146 -3471 0 FreeSans 2500 0 0 0 D14
port 24 nsew
flabel metal1 s 99171 -4022 99171 -4022 0 FreeSans 2500 0 0 0 D15
port 25 nsew
flabel metal1 s 4423 -2365 4423 -2365 0 FreeSans 2500 0 0 0 S7
port 26 nsew
flabel metal1 s 4793 -4573 4793 -4573 0 FreeSans 2500 0 0 0 D4
port 27 nsew
flabel metal1 s 4742 -4063 4742 -4063 0 FreeSans 2500 0 0 0 D6
port 28 nsew
flabel metal1 s 4675 -3537 4675 -3537 0 FreeSans 2500 0 0 0 D1
port 29 nsew
flabel metal1 s 4723 -3078 4723 -3078 0 FreeSans 2500 0 0 0 D5
port 30 nsew
flabel metal1 s 4752 -2715 4752 -2715 0 FreeSans 2500 0 0 0 D0
port 31 nsew
flabel metal1 s 4646 -1595 4646 -1595 0 FreeSans 2500 0 0 0 D2
port 32 nsew
flabel metal1 s 4579 -1155 4579 -1155 0 FreeSans 2500 0 0 0 D3
port 33 nsew
flabel metal1 s -3395 52547 -3395 52547 0 FreeSans 2500 0 0 0 D8
port 34 nsew
flabel metal1 s -3154 44010 -3154 44010 0 FreeSans 2500 0 0 0 D7
port 35 nsew
flabel metal1 s -3184 43467 -3184 43467 0 FreeSans 2500 0 0 0 D9
port 36 nsew
flabel metal1 s -3049 36634 -3049 36634 0 FreeSans 2500 0 0 0 D10
port 37 nsew
flabel metal1 s -3814 24857 -3814 24857 0 FreeSans 2500 0 0 0 PRE_SCALAR
port 38 nsew
flabel metal1 s 4188 9245 4188 9245 0 FreeSans 2500 0 0 0 UP_OUT
port 39 nsew
flabel metal1 s 5730 4634 5730 4634 0 FreeSans 2500 0 0 0 DN_OUT
port 40 nsew
flabel metal2 s 21999 15127 21999 15127 0 FreeSans 2500 0 0 0 UP
port 41 nsew
flabel metal2 s 22016 14545 22016 14545 0 FreeSans 2500 0 0 0 DN
port 42 nsew
flabel metal1 s 99365 4556 99365 4556 0 FreeSans 2500 0 0 0 VDD_TEST
port 43 nsew
flabel metal1 s 39830 6510 39830 6510 0 FreeSans 2500 0 0 0 VCTRL_OBV
port 44 nsew
flabel metal1 s 13110 -7700 13110 -7700 0 FreeSans 2500 0 0 0 Q02
port 45 nsew
flabel metal1 s 13860 -10180 13860 -10180 0 FreeSans 2500 0 0 0 Q07
port 46 nsew
flabel metal1 s 28770 -7800 28770 -7800 0 FreeSans 2500 0 0 0 Q01
port 47 nsew
flabel metal1 s 14210 -15910 14210 -15910 0 FreeSans 2500 0 0 0 Q05
port 48 nsew
flabel metal1 s 13110 -12310 13110 -12310 0 FreeSans 2500 0 0 0 Q06
port 49 nsew
flabel metal1 s 28860 -12250 28860 -12250 0 FreeSans 2500 0 0 0 Q03
port 50 nsew
flabel metal1 s 28010 -15010 28010 -15010 0 FreeSans 2500 0 0 0 Q04
port 51 nsew
flabel metal1 s 28920 -18000 28920 -18000 0 FreeSans 2500 0 0 0 P02
port 52 nsew
flabel metal1 s 6410 -8020 6410 -8020 0 FreeSans 2500 0 0 0 LD0
port 53 nsew
flabel metal1 s 43780 -18390 43780 -18390 0 FreeSans 2500 0 0 0 OUT01
port 54 nsew
flabel metal1 s 95190 -18410 95190 -18410 0 FreeSans 5000 0 0 0 OUT11
port 55 nsew
flabel metal1 s 57550 -8180 57550 -8180 0 FreeSans 5000 0 0 0 LD1
port 56 nsew
flabel metal1 s 64250 -7650 64250 -7650 0 FreeSans 5000 0 0 0 Q12
port 57 nsew
flabel metal1 s 79910 -7950 79910 -7950 0 FreeSans 5000 0 0 0 Q11
port 58 nsew
flabel metal1 s 64260 -11900 64260 -11900 0 FreeSans 5000 0 0 0 Q16
port 59 nsew
flabel metal1 s 80010 -12090 80010 -12090 0 FreeSans 5000 0 0 0 Q13
port 60 nsew
flabel metal1 s 65360 -15960 65360 -15960 0 FreeSans 5000 0 0 0 Q15
port 61 nsew
flabel metal1 s 79160 -15880 79160 -15880 0 FreeSans 5000 0 0 0 Q14
port 62 nsew
flabel metal1 s 65000 -10230 65000 -10230 0 FreeSans 5000 0 0 0 Q17
port 63 nsew
flabel metal1 s 80070 -17980 80070 -17980 0 FreeSans 5000 0 0 0 P12
port 64 nsew
flabel metal1 s 8667 22935 8667 22935 0 FreeSans 5000 0 0 0 OUT21
port 65 nsew
flabel metal1 s 4687 55482 4687 55482 0 FreeSans 5000 0 0 0 Q26
port 66 nsew
flabel metal1 s 2862 54749 2862 54749 0 FreeSans 5000 0 0 0 Q27
port 67 nsew
flabel metal1 s 8628 54398 8628 54398 0 FreeSans 5000 0 0 0 Q25
port 68 nsew
flabel metal1 s -561 55487 -561 55487 0 FreeSans 5000 0 0 0 Q22
port 69 nsew
flabel metal1 s -1095 48432 -1095 48432 0 FreeSans 5000 0 0 0 LD2
port 70 nsew
flabel metal1 s 137 39812 137 39812 0 FreeSans 5000 0 0 0 Q21
port 71 nsew
flabel metal1 s 4469 39744 4469 39744 0 FreeSans 5000 0 0 0 Q23
port 72 nsew
flabel metal1 s 7673 40583 7673 40583 0 FreeSans 5000 0 0 0 Q24
port 73 nsew
flabel metal1 s 48873 -14249 48873 -14249 0 FreeSans 2500 0 0 0 DIV_OUT
port 74 nsew
flabel metal1 s 2488 10382 2488 10382 0 FreeSans 2500 0 0 0 ITAIL
port 75 nsew
flabel metal1 s 5149 16633 5149 16633 0 FreeSans 2500 0 0 0 ITAIL_SRC
port 76 nsew
flabel metal1 s 5143 15231 5143 15231 0 FreeSans 2500 0 0 0 ITAIL_SINK
port 77 nsew
flabel metal2 s 2480 16670 2480 16670 0 FreeSans 2500 0 0 0 A0
port 78 nsew
flabel metal2 s 2530 15190 2530 15190 0 FreeSans 2500 0 0 0 A3
port 79 nsew
flabel metal2 s 2100 14450 2100 14450 0 FreeSans 2500 0 0 0 G1_2
port 80 nsew
flabel metal2 s 1230 14410 1230 14410 0 FreeSans 2500 0 0 0 SD0_1
port 81 nsew
flabel metal2 s 1970 11950 1970 11950 0 FreeSans 2500 0 0 0 SD2_1
port 82 nsew
flabel metal1 s 1720 10740 1720 10740 0 FreeSans 2500 0 0 0 G2_1
port 83 nsew
flabel metal2 s 940 13900 940 13900 0 FreeSans 2500 0 0 0 G1_1
port 84 nsew
flabel metal2 s -170 15280 -170 15280 0 FreeSans 2500 0 0 0 SD01
port 85 nsew
flabel metal1 s 50943 -423 50943 -423 0 FreeSans 2000 0 0 0 VSS
port 86 nsew
<< end >>
