* NGSPICE file created from pll_1_mag.ext - technology: gf180mcuC

.subckt pmos_3p3_M8SWPS a_n28_n124# a_n116_n80# a_28_n80# w_n202_n210#
X0 a_28_n80# a_n28_n124# a_n116_n80# w_n202_n210# pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
.ends

.subckt nmos_3p3_5QNVWA a_n116_n44# a_28_n44# a_n28_n88# VSUBS
X0 a_28_n44# a_n28_n88# a_n116_n44# VSUBS nfet_03v3 ad=0.194p pd=1.76u as=0.194p ps=1.76u w=0.44u l=0.28u
.ends

.subckt nand2_mag IN2 IN1 VSS OUT m1_186_70# VDD
Xpmos_3p3_M8SWPS_0 IN1 OUT VDD VDD pmos_3p3_M8SWPS
Xpmos_3p3_M8SWPS_1 IN2 VDD OUT VDD pmos_3p3_M8SWPS
Xnmos_3p3_5QNVWA_0 VSS m1_186_70# IN2 VSS nmos_3p3_5QNVWA
Xnmos_3p3_5QNVWA_1 m1_186_70# OUT IN1 VSS nmos_3p3_5QNVWA
.ends

.subckt nmos_3p3_VGTVWA a_n116_n66# a_28_n66# a_n28_n110# VSUBS
X0 a_28_n66# a_n28_n110# a_n116_n66# VSUBS nfet_03v3 ad=0.29p pd=2.2u as=0.29p ps=2.2u w=0.66u l=0.28u
.ends

.subckt nand3_mag IN3 IN2 IN1 nmos_3p3_VGTVWA_1/a_28_n66# VSS nmos_3p3_VGTVWA_0/a_28_n66#
+ OUT VDD
Xnmos_3p3_VGTVWA_0 nmos_3p3_VGTVWA_1/a_28_n66# nmos_3p3_VGTVWA_0/a_28_n66# IN2 VSS
+ nmos_3p3_VGTVWA
Xnmos_3p3_VGTVWA_1 VSS nmos_3p3_VGTVWA_1/a_28_n66# IN3 VSS nmos_3p3_VGTVWA
Xnmos_3p3_VGTVWA_2 nmos_3p3_VGTVWA_0/a_28_n66# OUT IN1 VSS nmos_3p3_VGTVWA
Xpmos_3p3_M8SWPS_0 IN1 VDD OUT VDD pmos_3p3_M8SWPS
Xpmos_3p3_M8SWPS_1 IN3 VDD OUT VDD pmos_3p3_M8SWPS
Xpmos_3p3_M8SWPS_2 IN2 OUT VDD VDD pmos_3p3_M8SWPS
.ends

.subckt pmos_3p3_MQGBLR a_n28_n124# a_n116_n80# a_28_n80# w_n202_n210#
X0 a_28_n80# a_n28_n124# a_n116_n80# w_n202_n210# pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
.ends

.subckt nmos_3p3_DDNVWA a_n120_n36# a_28_n22# a_n28_n66# VSUBS
X0 a_28_n22# a_n28_n66# a_n120_n36# VSUBS nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
.ends

.subckt GF_INV_MAG VDD VSS IN OUT
Xpmos_3p3_MQGBLR_0 IN VDD OUT VDD pmos_3p3_MQGBLR
Xnmos_3p3_DDNVWA_0 VSS OUT IN VSS nmos_3p3_DDNVWA
.ends

.subckt JK_FF_mag RST J K nand2_mag_1/m1_186_70# nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ nand2_mag_3/m1_186_70# nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66# nand2_mag_2/m1_186_70#
+ nand2_mag_4/m1_186_70# nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66# nand2_mag_4/IN2 nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# nand2_mag_1/IN2 nand3_mag_2/OUT nand3_mag_0/OUT
+ CLK QB nand3_mag_1/IN1 nand2_mag_3/IN1 nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66# nand2_mag_0/m1_186_70#
+ Q nand3_mag_1/OUT VDD VSS
Xnand2_mag_1 nand2_mag_1/IN2 QB VSS Q nand2_mag_1/m1_186_70# VDD nand2_mag
Xnand3_mag_2 J CLK Q nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66# VSS nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66#
+ nand3_mag_2/OUT VDD nand3_mag
Xnand2_mag_2 nand3_mag_0/OUT nand3_mag_1/OUT VSS nand3_mag_1/IN1 nand2_mag_2/m1_186_70#
+ VDD nand2_mag
Xnand2_mag_3 nand3_mag_1/OUT nand2_mag_3/IN1 VSS nand2_mag_4/IN2 nand2_mag_3/m1_186_70#
+ VDD nand2_mag
Xnand2_mag_4 nand2_mag_4/IN2 Q VSS QB nand2_mag_4/m1_186_70# VDD nand2_mag
XGF_INV_MAG_0 VDD VSS CLK nand2_mag_3/IN1 GF_INV_MAG
Xnand3_mag_0 K CLK QB nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66# VSS nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ nand3_mag_0/OUT VDD nand3_mag
Xnand2_mag_0 nand3_mag_1/IN1 nand2_mag_3/IN1 VSS nand2_mag_1/IN2 nand2_mag_0/m1_186_70#
+ VDD nand2_mag
Xnand3_mag_1 nand3_mag_2/OUT RST nand3_mag_1/IN1 nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ VSS nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66# nand3_mag_1/OUT VDD nand3_mag
.ends

.subckt pmos_3p3_M8QNDR w_n202_n290# a_28_n160# a_n116_n160# a_n28_n204#
X0 a_28_n160# a_n28_n204# a_n116_n160# w_n202_n290# pfet_03v3 ad=0.704p pd=4.08u as=0.704p ps=4.08u w=1.6u l=0.28u
.ends

.subckt pmos_3p3_M4YALR w_n202_n290# a_28_n160# a_n116_n160# a_n28_n204#
X0 a_28_n160# a_n28_n204# a_n116_n160# w_n202_n290# pfet_03v3 ad=0.704p pd=4.08u as=0.704p ps=4.08u w=1.6u l=0.28u
.ends

.subckt or_2_mag VSS VDD IN2 IN1 OUT
Xpmos_3p3_M8QNDR_0 VDD pmos_3p3_M8QNDR_0/a_28_n160# VDD IN2 pmos_3p3_M8QNDR
XGF_INV_MAG_1 VDD VSS GF_INV_MAG_1/IN OUT GF_INV_MAG
Xpmos_3p3_M4YALR_0 VDD GF_INV_MAG_1/IN pmos_3p3_M8QNDR_0/a_28_n160# IN1 pmos_3p3_M4YALR
Xnmos_3p3_DDNVWA_0 GF_INV_MAG_1/IN VSS IN1 VSS nmos_3p3_DDNVWA
Xnmos_3p3_DDNVWA_1 VSS GF_INV_MAG_1/IN IN2 VSS nmos_3p3_DDNVWA
.ends

.subckt and2_mag IN2 IN1 OUT VSS VDD
Xpmos_3p3_M8SWPS_0 IN1 GF_INV_MAG_0/IN VDD VDD pmos_3p3_M8SWPS
Xpmos_3p3_M8SWPS_1 IN2 VDD GF_INV_MAG_0/IN VDD pmos_3p3_M8SWPS
XGF_INV_MAG_0 VDD VSS GF_INV_MAG_0/IN OUT GF_INV_MAG
Xnmos_3p3_5QNVWA_0 VSS m1_186_70# IN2 VSS nmos_3p3_5QNVWA
Xnmos_3p3_5QNVWA_1 m1_186_70# GF_INV_MAG_0/IN IN1 VSS nmos_3p3_5QNVWA
.ends

.subckt pmos_3p3_MW53B7 a_n188_n80# a_n100_n124# a_100_n80# w_n274_n210#
X0 a_100_n80# a_n100_n124# a_n188_n80# w_n274_n210# pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
.ends

.subckt nmos_3p3_MGBSF7 a_100_n22# a_n100_n66# a_n192_n36# VSUBS
X0 a_100_n22# a_n100_n66# a_n192_n36# VSUBS nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
.ends

.subckt Inverter_delayed_mag VDD VSS IN OUT
Xpmos_3p3_MW53B7_0 VDD IN OUT VDD pmos_3p3_MW53B7
Xnmos_3p3_MGBSF7_0 OUT IN VSS VSS nmos_3p3_MGBSF7
.ends

.subckt Buffer_delayed_mag IN OUT VSS VDD
Xpmos_3p3_MW53B7_0 VDD IN Inverter_delayed_mag_0/IN VDD pmos_3p3_MW53B7
XInverter_delayed_mag_0 VDD VSS Inverter_delayed_mag_0/IN OUT Inverter_delayed_mag
Xnmos_3p3_MGBSF7_0 Inverter_delayed_mag_0/IN IN VSS VSS nmos_3p3_MGBSF7
.ends

.subckt pmos_3p3_MYFUKR a_28_n240# a_n28_n284# a_n116_n240# w_n202_n370#
X0 a_28_n240# a_n28_n284# a_n116_n240# w_n202_n370# pfet_03v3 ad=1.06p pd=5.68u as=1.06p ps=5.68u w=2.4u l=0.28u
.ends

.subckt nor_3_mag IN3 IN2 IN1 OUT VSS VDD
Xnmos_3p3_DDNVWA_2 OUT VSS IN2 VSS nmos_3p3_DDNVWA
Xpmos_3p3_MYFUKR_0 OUT IN1 pmos_3p3_MYFUKR_2/a_28_n240# VDD pmos_3p3_MYFUKR
Xpmos_3p3_MYFUKR_1 pmos_3p3_MYFUKR_1/a_28_n240# IN3 VDD VDD pmos_3p3_MYFUKR
Xpmos_3p3_MYFUKR_2 pmos_3p3_MYFUKR_2/a_28_n240# IN2 pmos_3p3_MYFUKR_1/a_28_n240# VDD
+ pmos_3p3_MYFUKR
Xnmos_3p3_DDNVWA_0 VSS OUT IN1 VSS nmos_3p3_DDNVWA
Xnmos_3p3_DDNVWA_1 VSS OUT IN3 VSS nmos_3p3_DDNVWA
.ends

.subckt CLK_DIV_11_mag_new CLK Vdiv11 Q3 Q2 Q1 Q0 RST VDD VSS
XJK_FF_mag_1 RST JK_FF_mag_1/K JK_FF_mag_1/K m1_7762_3820# m1_5915_5036# m1_7352_4917#
+ m1_6081_3939# m1_6634_3820# m1_7916_4917# m1_6799_5036# JK_FF_mag_1/nand2_mag_4/IN2
+ m1_5921_3939# m1_6075_5036# JK_FF_mag_1/nand2_mag_1/IN2 JK_FF_mag_1/nand3_mag_2/OUT
+ JK_FF_mag_1/nand3_mag_0/OUT CLK JK_FF_mag_1/QB JK_FF_mag_1/nand3_mag_1/IN1 JK_FF_mag_1/nand2_mag_3/IN1
+ m1_6639_5036# m1_7198_3820# Q2 JK_FF_mag_1/nand3_mag_1/OUT VDD VSS JK_FF_mag
XJK_FF_mag_0 RST JK_FF_mag_0/K JK_FF_mag_0/K m1_4627_3818# m1_2780_5034# m1_4217_4915#
+ m1_2946_3937# m1_3499_3818# m1_4781_4915# m1_3664_5034# JK_FF_mag_0/nand2_mag_4/IN2
+ m1_2786_3937# m1_2940_5034# JK_FF_mag_0/nand2_mag_1/IN2 JK_FF_mag_0/nand3_mag_2/OUT
+ JK_FF_mag_0/nand3_mag_0/OUT CLK or_2_mag_3/IN2 JK_FF_mag_0/nand3_mag_1/IN1 JK_FF_mag_0/nand2_mag_3/IN1
+ m1_3504_5034# m1_4063_3818# Q3 JK_FF_mag_0/nand3_mag_1/OUT VDD VSS JK_FF_mag
XJK_FF_mag_2 RST JK_FF_mag_2/K JK_FF_mag_2/K m1_10876_3818# m1_9029_5034# m1_10466_4915#
+ m1_9195_3937# m1_9748_3818# m1_11030_4915# m1_9913_5034# JK_FF_mag_2/nand2_mag_4/IN2
+ m1_9035_3937# m1_9189_5034# JK_FF_mag_2/nand2_mag_1/IN2 JK_FF_mag_2/nand3_mag_2/OUT
+ JK_FF_mag_2/nand3_mag_0/OUT CLK or_2_mag_3/IN1 JK_FF_mag_2/nand3_mag_1/IN1 JK_FF_mag_2/nand2_mag_3/IN1
+ m1_9753_5034# m1_10312_3818# Q1 JK_FF_mag_2/nand3_mag_1/OUT VDD VSS JK_FF_mag
XJK_FF_mag_3 RST JK_FF_mag_3/K JK_FF_mag_3/K m1_14035_3822# m1_12188_5038# m1_13625_4919#
+ m1_12354_3941# m1_12907_3822# m1_14189_4919# m1_13072_5038# JK_FF_mag_3/nand2_mag_4/IN2
+ m1_12194_3941# m1_12348_5038# JK_FF_mag_3/nand2_mag_1/IN2 JK_FF_mag_3/nand3_mag_2/OUT
+ JK_FF_mag_3/nand3_mag_0/OUT CLK JK_FF_mag_3/QB JK_FF_mag_3/nand3_mag_1/IN1 JK_FF_mag_3/nand2_mag_3/IN1
+ m1_12912_5038# m1_13471_3822# Q0 JK_FF_mag_3/nand3_mag_1/OUT VDD VSS JK_FF_mag
XGF_INV_MAG_0 VDD VSS nand3_mag_0/OUT or_2_mag_0/IN2 GF_INV_MAG
XGF_INV_MAG_1 VDD VSS nand3_mag_1/OUT GF_INV_MAG_1/OUT GF_INV_MAG
XGF_INV_MAG_2 VDD VSS nor_3_mag_0/OUT Vdiv11 GF_INV_MAG
Xor_2_mag_0 VSS VDD or_2_mag_0/IN2 or_2_mag_0/IN1 JK_FF_mag_0/K or_2_mag
Xor_2_mag_1 VSS VDD Q0 or_2_mag_1/IN1 JK_FF_mag_2/K or_2_mag
Xor_2_mag_3 VSS VDD or_2_mag_3/IN2 or_2_mag_3/IN1 JK_FF_mag_3/K or_2_mag
Xand2_mag_0 Q1 Q3 or_2_mag_0/IN1 VSS VDD and2_mag
Xand2_mag_1 Q0 Q1 JK_FF_mag_1/K VSS VDD and2_mag
Xand2_mag_2 Q1 Q3 or_2_mag_1/IN1 VSS VDD and2_mag
Xand2_mag_3 Q1 and2_mag_3/IN1 and2_mag_3/OUT VSS VDD and2_mag
XBuffer_delayed_mag_1 GF_INV_MAG_1/OUT nor_3_mag_0/IN3 VSS VDD Buffer_delayed_mag
XBuffer_delayed_mag_0 Q2 and2_mag_3/IN1 VSS VDD Buffer_delayed_mag
Xnor_3_mag_0 nor_3_mag_0/IN3 and2_mag_3/OUT Q3 nor_3_mag_0/OUT VSS VDD nor_3_mag
Xnand3_mag_0 Q1 Q0 Q2 nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66# VSS nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ nand3_mag_0/OUT VDD nand3_mag
Xnand3_mag_1 and2_mag_3/IN1 Q0 CLK nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66# VSS nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ nand3_mag_1/OUT VDD nand3_mag
.ends

.subckt CLK_div_10_mag RST CLK VDD Q0 Q1 Q2 Q3 Vdiv10 VSS
XJK_FF_mag_0 RST VDD JK_FF_mag_0/K JK_FF_mag_0/nand2_mag_1/m1_186_70# JK_FF_mag_0/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_0/nand2_mag_3/m1_186_70# JK_FF_mag_0/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_0/nand2_mag_2/m1_186_70# JK_FF_mag_0/nand2_mag_4/m1_186_70# JK_FF_mag_0/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_0/nand2_mag_4/IN2 JK_FF_mag_0/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_0/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_0/nand2_mag_1/IN2
+ JK_FF_mag_0/nand3_mag_2/OUT JK_FF_mag_0/nand3_mag_0/OUT Q0 JK_FF_mag_2/K JK_FF_mag_0/nand3_mag_1/IN1
+ JK_FF_mag_0/nand2_mag_3/IN1 JK_FF_mag_0/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_0/nand2_mag_0/m1_186_70# Q3 JK_FF_mag_0/nand3_mag_1/OUT VDD VSS JK_FF_mag
XJK_FF_mag_1 RST VDD VDD JK_FF_mag_1/nand2_mag_1/m1_186_70# JK_FF_mag_1/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_1/nand2_mag_3/m1_186_70# JK_FF_mag_1/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_1/nand2_mag_2/m1_186_70# JK_FF_mag_1/nand2_mag_4/m1_186_70# JK_FF_mag_1/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_1/nand2_mag_4/IN2 JK_FF_mag_1/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_1/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_1/nand2_mag_1/IN2
+ JK_FF_mag_1/nand3_mag_2/OUT JK_FF_mag_1/nand3_mag_0/OUT CLK JK_FF_mag_1/QB JK_FF_mag_1/nand3_mag_1/IN1
+ JK_FF_mag_1/nand2_mag_3/IN1 JK_FF_mag_1/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_1/nand2_mag_0/m1_186_70# Q0 JK_FF_mag_1/nand3_mag_1/OUT VDD VSS JK_FF_mag
XJK_FF_mag_2 RST VDD JK_FF_mag_2/K JK_FF_mag_2/nand2_mag_1/m1_186_70# JK_FF_mag_2/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_2/nand2_mag_3/m1_186_70# JK_FF_mag_2/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_2/nand2_mag_2/m1_186_70# JK_FF_mag_2/nand2_mag_4/m1_186_70# JK_FF_mag_2/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_2/nand2_mag_4/IN2 JK_FF_mag_2/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_2/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_2/nand2_mag_1/IN2
+ JK_FF_mag_2/nand3_mag_2/OUT JK_FF_mag_2/nand3_mag_0/OUT Q0 JK_FF_mag_2/QB JK_FF_mag_2/nand3_mag_1/IN1
+ JK_FF_mag_2/nand2_mag_3/IN1 JK_FF_mag_2/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_2/nand2_mag_0/m1_186_70# Q1 JK_FF_mag_2/nand3_mag_1/OUT VDD VSS JK_FF_mag
XJK_FF_mag_3 RST VDD VDD JK_FF_mag_3/nand2_mag_1/m1_186_70# JK_FF_mag_3/nand3_mag_2/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_3/nand2_mag_3/m1_186_70# JK_FF_mag_3/nand3_mag_0/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_3/nand2_mag_2/m1_186_70# JK_FF_mag_3/nand2_mag_4/m1_186_70# JK_FF_mag_3/nand3_mag_1/nmos_3p3_VGTVWA_0/a_28_n66#
+ JK_FF_mag_3/nand2_mag_4/IN2 JK_FF_mag_3/nand3_mag_0/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_3/nand3_mag_2/nmos_3p3_VGTVWA_0/a_28_n66# JK_FF_mag_3/nand2_mag_1/IN2
+ JK_FF_mag_3/nand3_mag_2/OUT JK_FF_mag_3/nand3_mag_0/OUT Q1 JK_FF_mag_3/QB JK_FF_mag_3/nand3_mag_1/IN1
+ JK_FF_mag_3/nand2_mag_3/IN1 JK_FF_mag_3/nand3_mag_1/nmos_3p3_VGTVWA_1/a_28_n66#
+ JK_FF_mag_3/nand2_mag_0/m1_186_70# Q2 JK_FF_mag_3/nand3_mag_1/OUT VDD VSS JK_FF_mag
Xand2_mag_0 Q1 Q2 and2_mag_0/OUT VSS VDD and2_mag
Xand2_mag_1 Q0 Q2 and2_mag_1/OUT VSS VDD and2_mag
Xand2_mag_2 Q2 Q1 JK_FF_mag_0/K VSS VDD and2_mag
XBuffer_delayed_mag_0 and2_mag_1/OUT nor_3_mag_0/IN3 VSS VDD Buffer_delayed_mag
Xnor_3_mag_0 nor_3_mag_0/IN3 and2_mag_0/OUT Q3 Vdiv10 VSS VDD nor_3_mag
.ends

.subckt CLK_div_110_mag VDD CLK Vdiv110 RST VSS
XCLK_DIV_11_mag_new_0 CLK CLK_div_10_mag_0/CLK CLK_DIV_11_mag_new_0/Q3 CLK_DIV_11_mag_new_0/Q2
+ CLK_DIV_11_mag_new_0/Q1 CLK_DIV_11_mag_new_0/Q0 RST VDD VSS CLK_DIV_11_mag_new
XCLK_div_10_mag_0 RST CLK_div_10_mag_0/CLK VDD CLK_div_10_mag_0/Q0 CLK_div_10_mag_0/Q1
+ CLK_div_10_mag_0/Q2 CLK_div_10_mag_0/Q3 Vdiv110 VSS CLK_div_10_mag
.ends

.subckt inv_my_mag VDD VSS IN OUT
Xpmos_3p3_MQGBLR_0 IN VDD OUT VDD pmos_3p3_MQGBLR
Xnmos_3p3_DDNVWA_0 VSS OUT IN VSS nmos_3p3_DDNVWA
.ends

.subckt nand2 VDD IN2 IN1 OUT VSS
Xpmos_3p3_M8SWPS_0 IN1 OUT VDD VDD pmos_3p3_M8SWPS
Xpmos_3p3_M8SWPS_1 IN2 VDD OUT VDD pmos_3p3_M8SWPS
Xnmos_3p3_5QNVWA_0 VSS m1_186_70# IN2 VSS nmos_3p3_5QNVWA
Xnmos_3p3_5QNVWA_1 m1_186_70# OUT IN1 VSS nmos_3p3_5QNVWA
.ends

.subckt inv VDD VSS IN OUT
Xpmos_3p3_MQGBLR_0 IN VDD OUT VDD pmos_3p3_MQGBLR
Xnmos_3p3_DDNVWA_0 VSS OUT IN VSS nmos_3p3_DDNVWA
.ends

.subckt DFF_ D RST CLK Q QB nand2_4/IN2 VDD VSS
Xnand2_6 VDD Q nand2_7/IN1 QB VSS nand2
Xnand2_7 VDD D nand2_7/IN1 nand2_7/OUT VSS nand2
Xinv_my_mag_0 VDD VSS inv_0/IN inv_0/OUT inv_my_mag
Xinv_0 VDD VSS inv_0/IN inv_0/OUT inv
Xnand2_0 VDD CLK RST nand2_5/IN2 VSS nand2
Xnand2_1 VDD inv_0/OUT nand2_5/IN2 nand2_4/IN2 VSS nand2
Xnand2_2 VDD nand2_4/IN2 nand2_7/OUT nand2_3/IN2 VSS nand2
Xnand2_3 VDD nand2_3/IN2 RST inv_0/IN VSS nand2
Xnand2_4 VDD nand2_4/IN2 QB Q VSS nand2
Xnand2_5 VDD nand2_5/IN2 inv_0/IN nand2_7/IN1 VSS nand2
.ends

.subckt nmos_3p3_5GGST2 a_n52_n50# a_n212_n50# a_52_n94# a_108_n50# a_n356_n50# a_268_n50#
+ a_n108_n94# a_n268_n94# a_212_n94# VSUBS
X0 a_108_n50# a_52_n94# a_n52_n50# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X1 a_268_n50# a_212_n94# a_108_n50# VSUBS nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X2 a_n52_n50# a_n108_n94# a_n212_n50# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X3 a_n212_n50# a_n268_n94# a_n356_n50# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
.ends

.subckt pmos_3p3_MWXUAR a_212_n144# a_268_n100# a_n268_n144# a_n356_n100# a_n52_n100#
+ a_n212_n100# w_n442_n230# a_108_n100# a_52_n144# a_n108_n144#
X0 a_n52_n100# a_n108_n144# a_n212_n100# w_n442_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_n212_n100# a_n268_n144# a_n356_n100# w_n442_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X2 a_108_n100# a_52_n144# a_n52_n100# w_n442_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_268_n100# a_212_n144# a_108_n100# w_n442_n230# pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt buffer_loading_mag VDD VSS OUT IN
Xnmos_3p3_5GGST2_0 VSS a_876_227# IN a_876_227# VSS VSS IN IN IN VSS nmos_3p3_5GGST2
Xpmos_3p3_MWXUAR_0 IN VDD IN VDD VDD a_876_227# VDD a_876_227# IN IN pmos_3p3_MWXUAR
X0 OUT a_876_227# VDD VDD pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 OUT a_876_227# VSS VSS nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X2 OUT a_876_227# VDD VDD pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X3 VSS a_876_227# OUT VSS nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X4 VDD a_876_227# OUT VDD pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X5 OUT a_876_227# VSS VSS nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X6 VSS a_876_227# OUT VSS nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X7 VDD a_876_227# OUT VDD pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt nmos_3p3_EA23U2 a_122_n100# a_n52_n100# a_n122_n144# a_296_n100# a_n226_n100#
+ a_n296_n144# a_n384_n100# a_52_n144# a_226_n144# VSUBS
X0 a_296_n100# a_226_n144# a_122_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.35u
X1 a_n226_n100# a_n296_n144# a_n384_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.35u
X2 a_n52_n100# a_n122_n144# a_n226_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X3 a_122_n100# a_52_n144# a_n52_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
.ends

.subckt pmos_3p3_M6H3WS a_n52_n50# a_n384_n50# a_296_n50# a_226_n94# a_n296_n94# w_n470_n180#
+ a_52_n94# a_n226_n50# a_122_n50# a_n122_n94#
X0 a_n52_n50# a_n122_n94# a_n226_n50# w_n470_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X1 a_122_n50# a_52_n94# a_n52_n50# w_n470_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X2 a_296_n50# a_226_n94# a_122_n50# w_n470_n180# pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.35u
X3 a_n226_n50# a_n296_n94# a_n384_n50# w_n470_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.35u
.ends

.subckt gf_inv_mag VDD VSS OUT IN
Xnmos_3p3_EA23U2_0 OUT VSS IN VSS OUT IN VSS IN IN VSS nmos_3p3_EA23U2
Xpmos_3p3_M6H3WS_0 VDD VDD VDD IN IN VDD IN OUT OUT IN pmos_3p3_M6H3WS
.ends

.subckt buffer_mag VDD OUT IN VSS
Xgf_inv_mag_0 VDD VSS gf_inv_mag_1/IN IN gf_inv_mag
Xgf_inv_mag_1 VDD VSS OUT gf_inv_mag_1/IN gf_inv_mag
.ends

.subckt PFD_layout PD PU VREF VDIV VDD VSS
Xinv_my_mag_0 VDD VSS VREF inv_0/OUT inv_my_mag
Xinv_my_mag_1 VDD VSS VDIV inv_1/OUT inv_my_mag
XDFF__0 VDD DFF__1/RST inv_1/OUT DFF__0/Q DFF__0/QB DFF__0/nand2_4/IN2 VDD VSS DFF_
XDFF__1 VDD DFF__1/RST inv_0/OUT DFF__1/Q DFF__1/QB DFF__1/nand2_4/IN2 VDD VSS DFF_
Xbuffer_loading_mag_0 VDD VSS PU DFF__1/Q buffer_loading_mag
Xbuffer_loading_mag_1 VDD VSS PD DFF__0/Q buffer_loading_mag
Xinv_0 VDD VSS VREF inv_0/OUT inv
Xinv_1 VDD VSS VDIV inv_1/OUT inv
Xbuffer_mag_0 VDD DFF__1/RST nand2_0/OUT VSS buffer_mag
Xnand2_0 VDD DFF__0/Q DFF__1/Q nand2_0/OUT VSS nand2
.ends

.subckt mim_2p0fF_WS3THJ m4_n4490_n4370# m4_n4370_n4250#
X0 m4_n4370_n4250# m4_n4490_n4370# cap_mim_2f0_m4m5_noshield c_width=42.5u c_length=42.5u
.ends

.subckt cap3p_layout Pp Nn
Xmim_2p0fF_WS3THJ_0 Nn Pp mim_2p0fF_WS3THJ
.ends

.subckt ppolyf_u_TPG873 a_1000_n1102# a_280_1000# a_n440_1000# a_n920_n1102# a_n440_n1102#
+ a_520_n1102# a_40_1000# a_n200_1000# a_n1160_1000# a_n200_n1102# a_n1160_n1102#
+ w_n1344_n1286# a_1000_1000# a_760_1000# a_n680_n1102# a_n920_1000# a_760_n1102#
+ a_520_1000# a_280_n1102# a_n680_1000# a_40_n1102#
X0 a_n680_1000# a_n680_n1102# w_n1344_n1286# ppolyf_u r_width=0.8u r_length=10u
X1 a_n920_1000# a_n920_n1102# w_n1344_n1286# ppolyf_u r_width=0.8u r_length=10u
X2 a_280_1000# a_280_n1102# w_n1344_n1286# ppolyf_u r_width=0.8u r_length=10u
X3 a_520_1000# a_520_n1102# w_n1344_n1286# ppolyf_u r_width=0.8u r_length=10u
X4 a_40_1000# a_40_n1102# w_n1344_n1286# ppolyf_u r_width=0.8u r_length=10u
X5 a_n1160_1000# a_n1160_n1102# w_n1344_n1286# ppolyf_u r_width=0.8u r_length=10u
X6 a_760_1000# a_760_n1102# w_n1344_n1286# ppolyf_u r_width=0.8u r_length=10u
X7 a_1000_1000# a_1000_n1102# w_n1344_n1286# ppolyf_u r_width=0.8u r_length=10u
X8 a_n200_1000# a_n200_n1102# w_n1344_n1286# ppolyf_u r_width=0.8u r_length=10u
X9 a_n440_1000# a_n440_n1102# w_n1344_n1286# ppolyf_u r_width=0.8u r_length=10u
.ends

.subckt res_48k_mag A B VDD
Xppolyf_u_TPG873_0 m1_n2577_205# m1_n3297_2306# m1_n3777_2306# m1_n4497_204# m1_n4017_204#
+ m1_n3057_204# m1_n3297_2306# m1_n3777_2306# A m1_n3537_204# m1_n4497_204# VDD B
+ m1_n2817_2306# m1_n4017_204# m1_n4257_2306# m1_n2577_205# m1_n2817_2306# m1_n3057_204#
+ m1_n4257_2306# m1_n3537_204# ppolyf_u_TPG873
.ends

.subckt mim_2p0fF_Q67PCK m4_5681_n21380# m4_11295_n21380# m4_n16775_n21380# m4_n22389_n21380#
+ m4_n11041_n21260# m4_17029_n21260# m4_5801_n21260# m4_11415_n21260# m4_67_n21380#
+ m4_n16655_n21260# m4_187_n21260# m4_n5547_n21380# m4_n22269_n21260# m4_16909_n21380#
+ m4_n11161_n21380# m4_n5427_n21260#
X0 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X1 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X2 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X3 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X4 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X5 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X6 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X7 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X8 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X9 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X10 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X11 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X12 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X13 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X14 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X15 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X16 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X17 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X18 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X19 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X20 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X21 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X22 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X23 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X24 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X25 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X26 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X27 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X28 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X29 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X30 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X31 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X32 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X33 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X34 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X35 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X36 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X37 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X38 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X39 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X40 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X41 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X42 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X43 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X44 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X45 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X46 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X47 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X48 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X49 m4_17029_n21260# m4_16909_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X50 m4_n11041_n21260# m4_n11161_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X51 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X52 m4_5801_n21260# m4_5681_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X53 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X54 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X55 m4_n16655_n21260# m4_n16775_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X56 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X57 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X58 m4_n5427_n21260# m4_n5547_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X59 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X60 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X61 m4_187_n21260# m4_67_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X62 m4_n22269_n21260# m4_n22389_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X63 m4_11415_n21260# m4_11295_n21380# cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
.ends

.subckt cap80p_mag P N
Xmim_2p0fF_Q67PCK_0 N N N N P P P P N P P N P N N P mim_2p0fF_Q67PCK
.ends

.subckt LF_mag VSS VDD VCNTL
Xcap3p_layout_0 VCNTL VSS cap3p_layout
Xres_48k_mag_0 VCNTL cap80p_mag_0/P VDD res_48k_mag
Xcap80p_mag_0 cap80p_mag_0/P VSS cap80p_mag
.ends

.subckt nmos_3p3_GYTGVN a_n260_n36# a_168_n28# a_56_n72# a_n168_n72# a_n56_n28# VSUBS
X0 a_n56_n28# a_n168_n72# a_n260_n36# VSUBS nfet_03v3 ad=92.8f pd=0.92u as=0.158p ps=1.64u w=0.28u l=0.56u
X1 a_168_n28# a_56_n72# a_n56_n28# VSUBS nfet_03v3 ad=0.158p pd=1.64u as=92.8f ps=0.92u w=0.28u l=0.56u
.ends

.subckt pmos_3p3_HVHFD7 a_n52_n50# w_n338_n180# a_52_n94# a_164_n50# a_n252_n50# a_n164_n94#
X0 a_164_n50# a_52_n94# a_n52_n50# w_n338_n180# pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.56u
X1 a_n52_n50# a_n164_n94# a_n252_n50# w_n338_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.56u
.ends

.subckt CP_mag VDD VSS VCNTL PU PD IPD_ IPD+
Xnmos_3p3_GYTGVN_0 m1_1391_990# m1_1391_990# PD PD VCNTL VSS nmos_3p3_GYTGVN
Xnmos_3p3_GYTGVN_1 VSS VSS IPD+ IPD+ IPD+ VSS nmos_3p3_GYTGVN
Xnmos_3p3_GYTGVN_2 VSS VSS IPD+ IPD+ m1_1391_990# VSS nmos_3p3_GYTGVN
Xpmos_3p3_HVHFD7_0 m1_1376_1265# VDD IPD_ VDD VDD IPD_ pmos_3p3_HVHFD7
Xpmos_3p3_HVHFD7_1 VCNTL VDD inv_0/OUT m1_1376_1265# m1_1376_1265# inv_0/OUT pmos_3p3_HVHFD7
Xpmos_3p3_HVHFD7_2 IPD_ VDD IPD_ VDD VDD IPD_ pmos_3p3_HVHFD7
Xinv_0 VDD VSS PU inv_0/OUT inv
.ends

.subckt nmos_3p3_9MTZEK a_n52_n70# a_52_n114# a_n122_n114# a_n210_n70# a_122_n70#
+ VSUBS
X0 a_n52_n70# a_n122_n114# a_n210_n70# VSUBS nfet_03v3 ad=0.182p pd=1.22u as=0.308p ps=2.28u w=0.7u l=0.35u
X1 a_122_n70# a_52_n114# a_n52_n70# VSUBS nfet_03v3 ad=0.308p pd=2.28u as=0.182p ps=1.22u w=0.7u l=0.35u
.ends

.subckt pmos_3p3_585UPK a_52_n184# a_122_n140# a_n52_n140# a_n122_n184# a_n210_n140#
+ w_n296_n270#
X0 a_122_n140# a_52_n184# a_n52_n140# w_n296_n270# pfet_03v3 ad=0.616p pd=3.68u as=0.364p ps=1.92u w=1.4u l=0.35u
X1 a_n52_n140# a_n122_n184# a_n210_n140# w_n296_n270# pfet_03v3 ad=0.364p pd=1.92u as=0.616p ps=3.68u w=1.4u l=0.35u
.ends

.subckt GF_INV4 VDD IN OUT VSS
Xnmos_3p3_9MTZEK_0 OUT IN IN VSS VSS VSS nmos_3p3_9MTZEK
Xpmos_3p3_585UPK_0 IN VDD OUT IN VDD VDD pmos_3p3_585UPK
.ends

.subckt pmos_3p3_ZB3RD7 a_268_n144# a_n52_n100# a_n468_n100# a_164_n100# a_380_n100#
+ a_n164_n144# a_n380_n144# a_52_n144# a_n268_n100# w_n554_n230#
X0 a_n268_n100# a_n380_n144# a_n468_n100# w_n554_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X1 a_380_n100# a_268_n144# a_164_n100# w_n554_n230# pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X2 a_164_n100# a_52_n144# a_n52_n100# w_n554_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X3 a_n52_n100# a_n164_n144# a_n268_n100# w_n554_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
.ends

.subckt nmos_3p3_FSHHD6 a_n52_n100# a_164_n100# a_n164_n144# a_n252_n100# a_52_n144#
+ VSUBS
X0 a_164_n100# a_52_n144# a_n52_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X1 a_n52_n100# a_n164_n144# a_n252_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
.ends

.subckt nmos_3p3_VMHHD6 a_268_n144# a_n52_n100# a_n468_n100# a_164_n100# a_380_n100#
+ a_n164_n144# a_n380_n144# a_52_n144# a_n268_n100# VSUBS
X0 a_n268_n100# a_n380_n144# a_n468_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X1 a_380_n100# a_268_n144# a_164_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X2 a_164_n100# a_52_n144# a_n52_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X3 a_n52_n100# a_n164_n144# a_n268_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
.ends

.subckt nmos_3p3_QNHHD6 a_56_n100# a_n56_n144# a_n144_n100# VSUBS
X0 a_56_n100# a_n56_n144# a_n144_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.56u
.ends

.subckt Delay_Cell_mag OUT OUTB EN VCONT INB IN VSS VDD
Xpmos_3p3_ZB3RD7_5 OUT VDD VDD OUTB VDD OUT OUT OUT OUTB VDD pmos_3p3_ZB3RD7
Xpmos_3p3_ZB3RD7_4 OUTB VDD VDD OUT VDD OUTB OUTB OUTB OUT VDD pmos_3p3_ZB3RD7
Xnmos_3p3_FSHHD6_0 a_562_n2079# VSS EN VSS EN VSS nmos_3p3_FSHHD6
Xnmos_3p3_VMHHD6_0 VCONT VSS VSS a_2095_n808# VSS VCONT VCONT VCONT a_2095_n808# VSS
+ nmos_3p3_VMHHD6
Xnmos_3p3_VMHHD6_2 INB a_562_n2079# a_562_n2079# OUTB a_562_n2079# INB INB INB OUTB
+ VSS nmos_3p3_VMHHD6
Xnmos_3p3_VMHHD6_1 IN a_562_n2079# a_562_n2079# OUT a_562_n2079# IN IN IN OUT VSS
+ nmos_3p3_VMHHD6
Xnmos_3p3_QNHHD6_0 a_562_n2079# a_562_n2079# a_562_n2079# VSS nmos_3p3_QNHHD6
Xnmos_3p3_QNHHD6_1 a_562_n2079# a_562_n2079# a_562_n2079# VSS nmos_3p3_QNHHD6
Xpmos_3p3_ZB3RD7_0 a_2095_n808# VDD VDD a_2095_n808# VDD a_2095_n808# a_2095_n808#
+ a_2095_n808# a_2095_n808# VDD pmos_3p3_ZB3RD7
Xpmos_3p3_ZB3RD7_1 OUT m1_277_n67# m1_277_n67# OUT m1_277_n67# OUT OUT OUT OUT VDD
+ pmos_3p3_ZB3RD7
Xpmos_3p3_ZB3RD7_2 OUTB m1_277_n67# m1_277_n67# OUTB m1_277_n67# OUTB OUTB OUTB OUTB
+ VDD pmos_3p3_ZB3RD7
Xpmos_3p3_ZB3RD7_3 a_2095_n808# m1_277_n67# m1_277_n67# VDD m1_277_n67# a_2095_n808#
+ a_2095_n808# a_2095_n808# VDD VDD pmos_3p3_ZB3RD7
.ends

.subckt nmos_3p3_AQSZEK a_n123_n70# a_35_n70# a_n35_n114# VSUBS
X0 a_35_n70# a_n35_n114# a_n123_n70# VSUBS nfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.35u
.ends

.subckt pmos_3p3_HBGRPK w_n213_n166# a_35_n35# a_n35_n79# a_n127_n36#
X0 a_35_n35# a_n35_n79# a_n127_n36# w_n213_n166# pfet_03v3 ad=0.165p pd=1.64u as=0.165p ps=1.64u w=0.35u l=0.35u
.ends

.subckt GF_INV1 VDD IN OUT VSS
Xnmos_3p3_AQSZEK_0 VSS OUT IN VSS nmos_3p3_AQSZEK
Xpmos_3p3_HBGRPK_0 VDD OUT IN VDD pmos_3p3_HBGRPK
.ends

.subckt pmos_3p3_MD4UPK a_52_n324# a_226_n324# a_122_n280# a_n52_n280# a_296_n280#
+ w_n470_n410# a_n226_n280# a_n384_n280# a_n122_n324# a_n296_n324#
X0 a_296_n280# a_226_n324# a_122_n280# w_n470_n410# pfet_03v3 ad=1.23p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.35u
X1 a_n226_n280# a_n296_n324# a_n384_n280# w_n470_n410# pfet_03v3 ad=0.728p pd=3.32u as=1.23p ps=6.48u w=2.8u l=0.35u
X2 a_122_n280# a_52_n324# a_n52_n280# w_n470_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.35u
X3 a_n52_n280# a_n122_n324# a_n226_n280# w_n470_n410# pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.35u
.ends

.subckt nmos_3p3_S7UZWU a_52_n184# a_226_n184# a_122_n140# a_n52_n140# a_n122_n184#
+ a_296_n140# a_n226_n140# a_n296_n184# a_n384_n140# VSUBS
X0 a_n226_n140# a_n296_n184# a_n384_n140# VSUBS nfet_03v3 ad=0.364p pd=1.92u as=0.616p ps=3.68u w=1.4u l=0.35u
X1 a_122_n140# a_52_n184# a_n52_n140# VSUBS nfet_03v3 ad=0.364p pd=1.92u as=0.364p ps=1.92u w=1.4u l=0.35u
X2 a_n52_n140# a_n122_n184# a_n226_n140# VSUBS nfet_03v3 ad=0.364p pd=1.92u as=0.364p ps=1.92u w=1.4u l=0.35u
X3 a_296_n140# a_226_n184# a_122_n140# VSUBS nfet_03v3 ad=0.616p pd=3.68u as=0.364p ps=1.92u w=1.4u l=0.35u
.ends

.subckt GF_INV16 VDD IN OUT VSS
Xpmos_3p3_MD4UPK_0 IN IN OUT VDD VDD VDD OUT VDD IN IN pmos_3p3_MD4UPK
Xnmos_3p3_S7UZWU_0 IN IN OUT VSS IN VSS OUT IN VSS VSS nmos_3p3_S7UZWU
.ends

.subckt pmos_3p3_HDJZPK a_n52_n50# a_n384_n50# a_296_n50# a_226_n94# a_n296_n94# w_n470_n180#
+ a_52_n94# a_n226_n50# a_122_n50# a_n122_n94#
X0 a_n52_n50# a_n122_n94# a_n226_n50# w_n470_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X1 a_122_n50# a_52_n94# a_n52_n50# w_n470_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X2 a_296_n50# a_226_n94# a_122_n50# w_n470_n180# pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.35u
X3 a_n226_n50# a_n296_n94# a_n384_n50# w_n470_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.35u
.ends

.subckt nmos_3p3_VDSZE6 a_122_n100# a_n52_n100# a_n122_n144# a_296_n100# a_n226_n100#
+ a_n296_n144# a_n384_n100# a_52_n144# a_226_n144# VSUBS
X0 a_296_n100# a_226_n144# a_122_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.35u
X1 a_n226_n100# a_n296_n144# a_n384_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.35u
X2 a_n52_n100# a_n122_n144# a_n226_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X3 a_122_n100# a_52_n144# a_n52_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
.ends

.subckt Stage_INV IN OUT VDD VSS
Xpmos_3p3_HDJZPK_0 VDD VDD VDD IN IN VDD IN OUT OUT IN pmos_3p3_HDJZPK
Xnmos_3p3_VDSZE6_0 OUT VSS IN VSS OUT IN VSS IN IN VSS nmos_3p3_VDSZE6
.ends

.subckt VCO_mag EN VCONT OUT OUTB VDD VSS
XGF_INV4_0 VDD GF_INV4_0/IN GF_INV4_0/OUT VSS GF_INV4
XGF_INV4_1 VDD GF_INV4_1/IN GF_INV4_1/OUT VSS GF_INV4
XDelay_Cell_mag_0 Delay_Cell_mag_3/INB Delay_Cell_mag_3/IN EN VCONT Stage_INV_0/OUT
+ Stage_INV_1/OUT VSS VDD Delay_Cell_mag
XGF_INV1_1 VDD GF_INV1_1/IN GF_INV4_1/IN VSS GF_INV1
XGF_INV1_0 VDD GF_INV1_0/IN GF_INV4_0/IN VSS GF_INV1
XDelay_Cell_mag_1 Delay_Cell_mag_2/INB Delay_Cell_mag_2/IN EN VCONT GF_INV1_0/IN GF_INV1_1/IN
+ VSS VDD Delay_Cell_mag
XGF_INV16_2 VDD GF_INV4_0/OUT OUT VSS GF_INV16
XGF_INV16_1 VDD GF_INV4_1/OUT OUTB VSS GF_INV16
XStage_INV_0 Stage_INV_0/IN Stage_INV_0/OUT VDD VSS Stage_INV
XDelay_Cell_mag_2 Stage_INV_0/IN Stage_INV_1/IN EN VCONT Delay_Cell_mag_2/INB Delay_Cell_mag_2/IN
+ VSS VDD Delay_Cell_mag
XDelay_Cell_mag_3 GF_INV1_0/IN GF_INV1_1/IN EN VCONT Delay_Cell_mag_3/INB Delay_Cell_mag_3/IN
+ VSS VDD Delay_Cell_mag
XStage_INV_1 Stage_INV_1/IN Stage_INV_1/OUT VDD VSS Stage_INV
.ends

.subckt pmos_3p3_Q354KU a_212_n144# a_268_n100# a_n692_n100# a_n268_n144# a_372_n144#
+ a_428_n100# a_n52_n100# a_n428_n144# a_532_n144# a_588_n100# w_n922_n230# a_n212_n100#
+ a_n588_n144# a_692_n144# a_748_n100# a_n372_n100# a_n748_n144# a_108_n100# a_52_n144#
+ a_n836_n100# a_n532_n100# a_n108_n144#
X0 a_n52_n100# a_n108_n144# a_n212_n100# w_n922_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_588_n100# a_532_n144# a_428_n100# w_n922_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 a_n212_n100# a_n268_n144# a_n372_n100# w_n922_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_n692_n100# a_n748_n144# a_n836_n100# w_n922_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X4 a_748_n100# a_692_n144# a_588_n100# w_n922_n230# pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X5 a_108_n100# a_52_n144# a_n52_n100# w_n922_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X6 a_268_n100# a_212_n144# a_108_n100# w_n922_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X7 a_n372_n100# a_n428_n144# a_n532_n100# w_n922_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X8 a_428_n100# a_372_n144# a_268_n100# w_n922_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X9 a_n532_n100# a_n588_n144# a_n692_n100# w_n922_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt nmos_3p3_W9BEG7 a_212_n144# a_268_n100# a_n692_n100# a_n268_n144# a_372_n144#
+ a_428_n100# a_n52_n100# a_n428_n144# a_532_n144# a_588_n100# a_n212_n100# a_n588_n144#
+ a_692_n144# a_748_n100# a_n372_n100# a_n748_n144# a_108_n100# a_52_n144# a_n836_n100#
+ a_n532_n100# a_n108_n144# VSUBS
X0 a_n52_n100# a_n108_n144# a_n212_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_588_n100# a_532_n144# a_428_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 a_n212_n100# a_n268_n144# a_n372_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_n692_n100# a_n748_n144# a_n836_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X4 a_748_n100# a_692_n144# a_588_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X5 a_108_n100# a_52_n144# a_n52_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X6 a_268_n100# a_212_n144# a_108_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X7 a_n372_n100# a_n428_n144# a_n532_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X8 a_428_n100# a_372_n144# a_268_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X9 a_n532_n100# a_n588_n144# a_n692_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt Transmission_gate_mag CLK VDD VIN VOUT VSS
Xinv_my_mag_0 VDD VSS CLK inv_my_mag_0/OUT inv_my_mag
Xpmos_3p3_Q354KU_0 inv_my_mag_0/OUT VOUT VOUT inv_my_mag_0/OUT inv_my_mag_0/OUT VIN
+ VOUT inv_my_mag_0/OUT inv_my_mag_0/OUT VOUT VDD VIN inv_my_mag_0/OUT inv_my_mag_0/OUT
+ VIN VOUT inv_my_mag_0/OUT VIN inv_my_mag_0/OUT VIN VIN inv_my_mag_0/OUT pmos_3p3_Q354KU
Xnmos_3p3_W9BEG7_0 CLK VOUT VOUT CLK CLK VIN VOUT CLK CLK VOUT VIN CLK CLK VIN VOUT
+ CLK VIN CLK VIN VIN CLK VSS nmos_3p3_W9BEG7
.ends

.subckt a2x1mux_mag IN1 IN2 SEL VOUT VDD VSS
Xinv_my_mag_0 VDD VSS SEL inv_my_mag_0/OUT inv_my_mag
XTransmission_gate_mag_0 inv_my_mag_0/OUT VDD IN1 VOUT VSS Transmission_gate_mag
XTransmission_gate_mag_1 SEL VDD IN2 VOUT VSS Transmission_gate_mag
.ends

.subckt pll_1_mag EN VDD_VCO Vref IPD_ IPD+ LP_ext RST_DIV pu pd VSS VDD VCO_op VCO_op_bar
XCLK_div_110_mag_0 VDD VCO_op PFD_layout_0/VDIV RST_DIV VSS CLK_div_110_mag
XPFD_layout_0 pd pu Vref PFD_layout_0/VDIV VDD VSS PFD_layout
XLF_mag_0 VSS VDD LF_mag_0/VCNTL LF_mag
XCP_mag_0 VDD VSS CP_mag_0/VCNTL pu pd IPD_ IPD+ CP_mag
XVCO_mag_0 EN CP_mag_0/VCNTL VCO_op VCO_op_bar VDD_VCO VSS VCO_mag
Xa2x1mux_mag_0 LP_ext LF_mag_0/VCNTL a2x1mux_mag_0/SEL CP_mag_0/VCNTL VDD VSS a2x1mux_mag
.ends

