magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1262 -1046 1262 1046
<< metal1 >>
rect -262 40 262 46
rect -262 14 -256 40
rect -230 14 -202 40
rect -176 14 -148 40
rect -122 14 -94 40
rect -68 14 -40 40
rect -14 14 14 40
rect 40 14 68 40
rect 94 14 122 40
rect 148 14 176 40
rect 202 14 230 40
rect 256 14 262 40
rect -262 -14 262 14
rect -262 -40 -256 -14
rect -230 -40 -202 -14
rect -176 -40 -148 -14
rect -122 -40 -94 -14
rect -68 -40 -40 -14
rect -14 -40 14 -14
rect 40 -40 68 -14
rect 94 -40 122 -14
rect 148 -40 176 -14
rect 202 -40 230 -14
rect 256 -40 262 -14
rect -262 -46 262 -40
<< via1 >>
rect -256 14 -230 40
rect -202 14 -176 40
rect -148 14 -122 40
rect -94 14 -68 40
rect -40 14 -14 40
rect 14 14 40 40
rect 68 14 94 40
rect 122 14 148 40
rect 176 14 202 40
rect 230 14 256 40
rect -256 -40 -230 -14
rect -202 -40 -176 -14
rect -148 -40 -122 -14
rect -94 -40 -68 -14
rect -40 -40 -14 -14
rect 14 -40 40 -14
rect 68 -40 94 -14
rect 122 -40 148 -14
rect 176 -40 202 -14
rect 230 -40 256 -14
<< metal2 >>
rect -262 40 262 46
rect -262 14 -256 40
rect -230 14 -202 40
rect -176 14 -148 40
rect -122 14 -94 40
rect -68 14 -40 40
rect -14 14 14 40
rect 40 14 68 40
rect 94 14 122 40
rect 148 14 176 40
rect 202 14 230 40
rect 256 14 262 40
rect -262 -14 262 14
rect -262 -40 -256 -14
rect -230 -40 -202 -14
rect -176 -40 -148 -14
rect -122 -40 -94 -14
rect -68 -40 -40 -14
rect -14 -40 14 -14
rect 40 -40 68 -14
rect 94 -40 122 -14
rect 148 -40 176 -14
rect 202 -40 230 -14
rect 256 -40 262 -14
rect -262 -46 262 -40
<< end >>
