magic
tech gf180mcuC
magscale 1 10
timestamp 1693911244
<< nwell >>
rect -282 -1902 282 1902
<< pmos >>
rect -108 1172 -52 1772
rect 52 1172 108 1772
rect -108 436 -52 1036
rect 52 436 108 1036
rect -108 -300 -52 300
rect 52 -300 108 300
rect -108 -1036 -52 -436
rect 52 -1036 108 -436
rect -108 -1772 -52 -1172
rect 52 -1772 108 -1172
<< pdiff >>
rect -196 1759 -108 1772
rect -196 1185 -183 1759
rect -137 1185 -108 1759
rect -196 1172 -108 1185
rect -52 1759 52 1772
rect -52 1185 -23 1759
rect 23 1185 52 1759
rect -52 1172 52 1185
rect 108 1759 196 1772
rect 108 1185 137 1759
rect 183 1185 196 1759
rect 108 1172 196 1185
rect -196 1023 -108 1036
rect -196 449 -183 1023
rect -137 449 -108 1023
rect -196 436 -108 449
rect -52 1023 52 1036
rect -52 449 -23 1023
rect 23 449 52 1023
rect -52 436 52 449
rect 108 1023 196 1036
rect 108 449 137 1023
rect 183 449 196 1023
rect 108 436 196 449
rect -196 287 -108 300
rect -196 -287 -183 287
rect -137 -287 -108 287
rect -196 -300 -108 -287
rect -52 287 52 300
rect -52 -287 -23 287
rect 23 -287 52 287
rect -52 -300 52 -287
rect 108 287 196 300
rect 108 -287 137 287
rect 183 -287 196 287
rect 108 -300 196 -287
rect -196 -449 -108 -436
rect -196 -1023 -183 -449
rect -137 -1023 -108 -449
rect -196 -1036 -108 -1023
rect -52 -449 52 -436
rect -52 -1023 -23 -449
rect 23 -1023 52 -449
rect -52 -1036 52 -1023
rect 108 -449 196 -436
rect 108 -1023 137 -449
rect 183 -1023 196 -449
rect 108 -1036 196 -1023
rect -196 -1185 -108 -1172
rect -196 -1759 -183 -1185
rect -137 -1759 -108 -1185
rect -196 -1772 -108 -1759
rect -52 -1185 52 -1172
rect -52 -1759 -23 -1185
rect 23 -1759 52 -1185
rect -52 -1772 52 -1759
rect 108 -1185 196 -1172
rect 108 -1759 137 -1185
rect 183 -1759 196 -1185
rect 108 -1772 196 -1759
<< pdiffc >>
rect -183 1185 -137 1759
rect -23 1185 23 1759
rect 137 1185 183 1759
rect -183 449 -137 1023
rect -23 449 23 1023
rect 137 449 183 1023
rect -183 -287 -137 287
rect -23 -287 23 287
rect 137 -287 183 287
rect -183 -1023 -137 -449
rect -23 -1023 23 -449
rect 137 -1023 183 -449
rect -183 -1759 -137 -1185
rect -23 -1759 23 -1185
rect 137 -1759 183 -1185
<< polysilicon >>
rect -108 1772 -52 1816
rect 52 1772 108 1816
rect -108 1128 -52 1172
rect 52 1128 108 1172
rect -108 1036 -52 1080
rect 52 1036 108 1080
rect -108 392 -52 436
rect 52 392 108 436
rect -108 300 -52 344
rect 52 300 108 344
rect -108 -344 -52 -300
rect 52 -344 108 -300
rect -108 -436 -52 -392
rect 52 -436 108 -392
rect -108 -1080 -52 -1036
rect 52 -1080 108 -1036
rect -108 -1172 -52 -1128
rect 52 -1172 108 -1128
rect -108 -1816 -52 -1772
rect 52 -1816 108 -1772
<< metal1 >>
rect -183 1759 -137 1770
rect -183 1174 -137 1185
rect -23 1759 23 1770
rect -23 1174 23 1185
rect 137 1759 183 1770
rect 137 1174 183 1185
rect -183 1023 -137 1034
rect -183 438 -137 449
rect -23 1023 23 1034
rect -23 438 23 449
rect 137 1023 183 1034
rect 137 438 183 449
rect -183 287 -137 298
rect -183 -298 -137 -287
rect -23 287 23 298
rect -23 -298 23 -287
rect 137 287 183 298
rect 137 -298 183 -287
rect -183 -449 -137 -438
rect -183 -1034 -137 -1023
rect -23 -449 23 -438
rect -23 -1034 23 -1023
rect 137 -449 183 -438
rect 137 -1034 183 -1023
rect -183 -1185 -137 -1174
rect -183 -1770 -137 -1759
rect -23 -1185 23 -1174
rect -23 -1770 23 -1759
rect 137 -1185 183 -1174
rect 137 -1770 183 -1759
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 3 l 0.280 m 5 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
