magic
tech gf180mcuC
magscale 1 10
timestamp 1690287175
<< nwell >>
rect 75 2351 639 2861
rect 838 2351 1402 2861
rect 1649 2351 2213 2861
rect 75 1380 639 1890
rect 838 1380 1402 1890
rect 1649 1380 2213 1890
rect 75 405 639 915
rect 838 404 1402 914
rect 1649 404 2213 914
<< pwell >>
rect 366 2323 426 2324
rect 1129 2323 1189 2324
rect 1940 2323 2000 2324
rect 366 2279 429 2323
rect 1129 2279 1192 2323
rect 1940 2279 2003 2323
rect 137 2043 577 2279
rect 900 2043 1340 2279
rect 1711 2043 2151 2279
rect 366 1352 426 1353
rect 1129 1352 1189 1353
rect 1940 1352 2000 1353
rect 366 1308 429 1352
rect 1129 1308 1192 1352
rect 1940 1308 2003 1352
rect 137 1072 577 1308
rect 900 1072 1340 1308
rect 1711 1072 2151 1308
rect 366 377 426 378
rect 366 333 429 377
rect 1129 376 1189 377
rect 1940 376 2000 377
rect 137 97 577 333
rect 1129 332 1192 376
rect 1940 332 2003 376
rect 900 96 1340 332
rect 1711 96 2151 332
<< nmos >>
rect 249 2111 305 2211
rect 409 2111 465 2211
rect 1012 2111 1068 2211
rect 1172 2111 1228 2211
rect 1823 2111 1879 2211
rect 1983 2111 2039 2211
rect 249 1140 305 1240
rect 409 1140 465 1240
rect 1012 1140 1068 1240
rect 1172 1140 1228 1240
rect 1823 1140 1879 1240
rect 1983 1140 2039 1240
rect 249 165 305 265
rect 409 165 465 265
rect 1012 164 1068 264
rect 1172 164 1228 264
rect 1823 164 1879 264
rect 1983 164 2039 264
<< pmos >>
rect 249 2481 305 2581
rect 409 2481 465 2581
rect 1012 2481 1068 2581
rect 1172 2481 1228 2581
rect 1823 2481 1879 2581
rect 1983 2481 2039 2581
rect 249 1510 305 1610
rect 409 1510 465 1610
rect 1012 1510 1068 1610
rect 1172 1510 1228 1610
rect 1823 1510 1879 1610
rect 1983 1510 2039 1610
rect 249 535 305 635
rect 409 535 465 635
rect 1012 534 1068 634
rect 1172 534 1228 634
rect 1823 534 1879 634
rect 1983 534 2039 634
<< ndiff >>
rect 161 2198 249 2211
rect 161 2124 174 2198
rect 220 2124 249 2198
rect 161 2111 249 2124
rect 305 2198 409 2211
rect 305 2124 334 2198
rect 380 2124 409 2198
rect 305 2111 409 2124
rect 465 2198 553 2211
rect 465 2124 494 2198
rect 540 2124 553 2198
rect 465 2111 553 2124
rect 924 2198 1012 2211
rect 924 2124 937 2198
rect 983 2124 1012 2198
rect 924 2111 1012 2124
rect 1068 2198 1172 2211
rect 1068 2124 1097 2198
rect 1143 2124 1172 2198
rect 1068 2111 1172 2124
rect 1228 2198 1316 2211
rect 1228 2124 1257 2198
rect 1303 2124 1316 2198
rect 1228 2111 1316 2124
rect 1735 2198 1823 2211
rect 1735 2124 1748 2198
rect 1794 2124 1823 2198
rect 1735 2111 1823 2124
rect 1879 2198 1983 2211
rect 1879 2124 1908 2198
rect 1954 2124 1983 2198
rect 1879 2111 1983 2124
rect 2039 2198 2127 2211
rect 2039 2124 2068 2198
rect 2114 2124 2127 2198
rect 2039 2111 2127 2124
rect 161 1227 249 1240
rect 161 1153 174 1227
rect 220 1153 249 1227
rect 161 1140 249 1153
rect 305 1227 409 1240
rect 305 1153 334 1227
rect 380 1153 409 1227
rect 305 1140 409 1153
rect 465 1227 553 1240
rect 465 1153 494 1227
rect 540 1153 553 1227
rect 465 1140 553 1153
rect 924 1227 1012 1240
rect 924 1153 937 1227
rect 983 1153 1012 1227
rect 924 1140 1012 1153
rect 1068 1227 1172 1240
rect 1068 1153 1097 1227
rect 1143 1153 1172 1227
rect 1068 1140 1172 1153
rect 1228 1227 1316 1240
rect 1228 1153 1257 1227
rect 1303 1153 1316 1227
rect 1228 1140 1316 1153
rect 1735 1227 1823 1240
rect 1735 1153 1748 1227
rect 1794 1153 1823 1227
rect 1735 1140 1823 1153
rect 1879 1227 1983 1240
rect 1879 1153 1908 1227
rect 1954 1153 1983 1227
rect 1879 1140 1983 1153
rect 2039 1227 2127 1240
rect 2039 1153 2068 1227
rect 2114 1153 2127 1227
rect 2039 1140 2127 1153
rect 161 252 249 265
rect 161 178 174 252
rect 220 178 249 252
rect 161 165 249 178
rect 305 252 409 265
rect 305 178 334 252
rect 380 178 409 252
rect 305 165 409 178
rect 465 252 553 265
rect 465 178 494 252
rect 540 178 553 252
rect 465 165 553 178
rect 924 251 1012 264
rect 924 177 937 251
rect 983 177 1012 251
rect 924 164 1012 177
rect 1068 251 1172 264
rect 1068 177 1097 251
rect 1143 177 1172 251
rect 1068 164 1172 177
rect 1228 251 1316 264
rect 1228 177 1257 251
rect 1303 177 1316 251
rect 1228 164 1316 177
rect 1735 251 1823 264
rect 1735 177 1748 251
rect 1794 177 1823 251
rect 1735 164 1823 177
rect 1879 251 1983 264
rect 1879 177 1908 251
rect 1954 177 1983 251
rect 1879 164 1983 177
rect 2039 251 2127 264
rect 2039 177 2068 251
rect 2114 177 2127 251
rect 2039 164 2127 177
<< pdiff >>
rect 161 2568 249 2581
rect 161 2494 174 2568
rect 220 2494 249 2568
rect 161 2481 249 2494
rect 305 2568 409 2581
rect 305 2494 334 2568
rect 380 2494 409 2568
rect 305 2481 409 2494
rect 465 2568 553 2581
rect 465 2494 494 2568
rect 540 2494 553 2568
rect 465 2481 553 2494
rect 924 2568 1012 2581
rect 924 2494 937 2568
rect 983 2494 1012 2568
rect 924 2481 1012 2494
rect 1068 2568 1172 2581
rect 1068 2494 1097 2568
rect 1143 2494 1172 2568
rect 1068 2481 1172 2494
rect 1228 2568 1316 2581
rect 1228 2494 1257 2568
rect 1303 2494 1316 2568
rect 1228 2481 1316 2494
rect 1735 2568 1823 2581
rect 1735 2494 1748 2568
rect 1794 2494 1823 2568
rect 1735 2481 1823 2494
rect 1879 2568 1983 2581
rect 1879 2494 1908 2568
rect 1954 2494 1983 2568
rect 1879 2481 1983 2494
rect 2039 2568 2127 2581
rect 2039 2494 2068 2568
rect 2114 2494 2127 2568
rect 2039 2481 2127 2494
rect 161 1597 249 1610
rect 161 1523 174 1597
rect 220 1523 249 1597
rect 161 1510 249 1523
rect 305 1597 409 1610
rect 305 1523 334 1597
rect 380 1523 409 1597
rect 305 1510 409 1523
rect 465 1597 553 1610
rect 465 1523 494 1597
rect 540 1523 553 1597
rect 465 1510 553 1523
rect 924 1597 1012 1610
rect 924 1523 937 1597
rect 983 1523 1012 1597
rect 924 1510 1012 1523
rect 1068 1597 1172 1610
rect 1068 1523 1097 1597
rect 1143 1523 1172 1597
rect 1068 1510 1172 1523
rect 1228 1597 1316 1610
rect 1228 1523 1257 1597
rect 1303 1523 1316 1597
rect 1228 1510 1316 1523
rect 1735 1597 1823 1610
rect 1735 1523 1748 1597
rect 1794 1523 1823 1597
rect 1735 1510 1823 1523
rect 1879 1597 1983 1610
rect 1879 1523 1908 1597
rect 1954 1523 1983 1597
rect 1879 1510 1983 1523
rect 2039 1597 2127 1610
rect 2039 1523 2068 1597
rect 2114 1523 2127 1597
rect 2039 1510 2127 1523
rect 161 622 249 635
rect 161 548 174 622
rect 220 548 249 622
rect 161 535 249 548
rect 305 622 409 635
rect 305 548 334 622
rect 380 548 409 622
rect 305 535 409 548
rect 465 622 553 635
rect 465 548 494 622
rect 540 548 553 622
rect 465 535 553 548
rect 924 621 1012 634
rect 924 547 937 621
rect 983 547 1012 621
rect 924 534 1012 547
rect 1068 621 1172 634
rect 1068 547 1097 621
rect 1143 547 1172 621
rect 1068 534 1172 547
rect 1228 621 1316 634
rect 1228 547 1257 621
rect 1303 547 1316 621
rect 1228 534 1316 547
rect 1735 621 1823 634
rect 1735 547 1748 621
rect 1794 547 1823 621
rect 1735 534 1823 547
rect 1879 621 1983 634
rect 1879 547 1908 621
rect 1954 547 1983 621
rect 1879 534 1983 547
rect 2039 621 2127 634
rect 2039 547 2068 621
rect 2114 547 2127 621
rect 2039 534 2127 547
<< ndiffc >>
rect 174 2124 220 2198
rect 334 2124 380 2198
rect 494 2124 540 2198
rect 937 2124 983 2198
rect 1097 2124 1143 2198
rect 1257 2124 1303 2198
rect 1748 2124 1794 2198
rect 1908 2124 1954 2198
rect 2068 2124 2114 2198
rect 174 1153 220 1227
rect 334 1153 380 1227
rect 494 1153 540 1227
rect 937 1153 983 1227
rect 1097 1153 1143 1227
rect 1257 1153 1303 1227
rect 1748 1153 1794 1227
rect 1908 1153 1954 1227
rect 2068 1153 2114 1227
rect 174 178 220 252
rect 334 178 380 252
rect 494 178 540 252
rect 937 177 983 251
rect 1097 177 1143 251
rect 1257 177 1303 251
rect 1748 177 1794 251
rect 1908 177 1954 251
rect 2068 177 2114 251
<< pdiffc >>
rect 174 2494 220 2568
rect 334 2494 380 2568
rect 494 2494 540 2568
rect 937 2494 983 2568
rect 1097 2494 1143 2568
rect 1257 2494 1303 2568
rect 1748 2494 1794 2568
rect 1908 2494 1954 2568
rect 2068 2494 2114 2568
rect 174 1523 220 1597
rect 334 1523 380 1597
rect 494 1523 540 1597
rect 937 1523 983 1597
rect 1097 1523 1143 1597
rect 1257 1523 1303 1597
rect 1748 1523 1794 1597
rect 1908 1523 1954 1597
rect 2068 1523 2114 1597
rect 174 548 220 622
rect 334 548 380 622
rect 494 548 540 622
rect 937 547 983 621
rect 1097 547 1143 621
rect 1257 547 1303 621
rect 1748 547 1794 621
rect 1908 547 1954 621
rect 2068 547 2114 621
<< psubdiff >>
rect 87 2017 641 2033
rect 87 1969 118 2017
rect 587 1969 641 2017
rect 87 1951 641 1969
rect 850 2017 1404 2033
rect 850 1969 881 2017
rect 1350 1969 1404 2017
rect 850 1951 1404 1969
rect 1661 2017 2215 2033
rect 1661 1969 1692 2017
rect 2161 1969 2215 2017
rect 1661 1951 2215 1969
rect 87 1046 641 1062
rect 87 998 118 1046
rect 587 998 641 1046
rect 87 980 641 998
rect 850 1046 1404 1062
rect 850 998 881 1046
rect 1350 998 1404 1046
rect 850 980 1404 998
rect 1661 1046 2215 1062
rect 1661 998 1692 1046
rect 2161 998 2215 1046
rect 1661 980 2215 998
rect 87 71 641 87
rect 87 23 118 71
rect 587 23 641 71
rect 87 5 641 23
rect 850 70 1404 86
rect 850 22 881 70
rect 1350 22 1404 70
rect 850 4 1404 22
rect 1661 70 2215 86
rect 1661 22 1692 70
rect 2161 22 2215 70
rect 1661 4 2215 22
<< nsubdiff >>
rect 153 2815 559 2835
rect 153 2759 190 2815
rect 502 2759 559 2815
rect 153 2738 559 2759
rect 916 2815 1322 2835
rect 916 2759 953 2815
rect 1265 2759 1322 2815
rect 916 2738 1322 2759
rect 1727 2815 2133 2835
rect 1727 2759 1764 2815
rect 2076 2759 2133 2815
rect 1727 2738 2133 2759
rect 153 1844 559 1864
rect 153 1788 190 1844
rect 502 1788 559 1844
rect 153 1767 559 1788
rect 916 1844 1322 1864
rect 916 1788 953 1844
rect 1265 1788 1322 1844
rect 916 1767 1322 1788
rect 1727 1844 2133 1864
rect 1727 1788 1764 1844
rect 2076 1788 2133 1844
rect 1727 1767 2133 1788
rect 153 869 559 889
rect 153 813 190 869
rect 502 813 559 869
rect 153 792 559 813
rect 916 868 1322 888
rect 916 812 953 868
rect 1265 812 1322 868
rect 916 791 1322 812
rect 1727 868 2133 888
rect 1727 812 1764 868
rect 2076 812 2133 868
rect 1727 791 2133 812
<< psubdiffcont >>
rect 118 1969 587 2017
rect 881 1969 1350 2017
rect 1692 1969 2161 2017
rect 118 998 587 1046
rect 881 998 1350 1046
rect 1692 998 2161 1046
rect 118 23 587 71
rect 881 22 1350 70
rect 1692 22 2161 70
<< nsubdiffcont >>
rect 190 2759 502 2815
rect 953 2759 1265 2815
rect 1764 2759 2076 2815
rect 190 1788 502 1844
rect 953 1788 1265 1844
rect 1764 1788 2076 1844
rect 190 813 502 869
rect 953 812 1265 868
rect 1764 812 2076 868
<< polysilicon >>
rect 249 2581 305 2625
rect 409 2581 465 2625
rect 1012 2581 1068 2625
rect 1172 2581 1228 2625
rect 1823 2581 1879 2625
rect 1983 2581 2039 2625
rect 249 2437 305 2481
rect 175 2423 305 2437
rect 175 2364 189 2423
rect 252 2364 305 2423
rect 175 2349 305 2364
rect 249 2211 305 2349
rect 409 2336 465 2481
rect 1012 2437 1068 2481
rect 938 2423 1068 2437
rect 938 2364 952 2423
rect 1015 2364 1068 2423
rect 938 2349 1068 2364
rect 353 2323 465 2336
rect 353 2264 366 2323
rect 429 2264 465 2323
rect 353 2251 465 2264
rect 409 2211 465 2251
rect 1012 2211 1068 2349
rect 1172 2336 1228 2481
rect 1823 2437 1879 2481
rect 1749 2423 1879 2437
rect 1749 2364 1763 2423
rect 1826 2364 1879 2423
rect 1749 2349 1879 2364
rect 1116 2323 1228 2336
rect 1116 2264 1129 2323
rect 1192 2264 1228 2323
rect 1116 2251 1228 2264
rect 1172 2211 1228 2251
rect 1823 2211 1879 2349
rect 1983 2336 2039 2481
rect 1927 2323 2039 2336
rect 1927 2264 1940 2323
rect 2003 2264 2039 2323
rect 1927 2251 2039 2264
rect 1983 2211 2039 2251
rect 249 2067 305 2111
rect 409 2067 465 2111
rect 1012 2067 1068 2111
rect 1172 2067 1228 2111
rect 1823 2067 1879 2111
rect 1983 2067 2039 2111
rect 249 1610 305 1654
rect 409 1610 465 1654
rect 1012 1610 1068 1654
rect 1172 1610 1228 1654
rect 1823 1610 1879 1654
rect 1983 1610 2039 1654
rect 249 1466 305 1510
rect 175 1452 305 1466
rect 175 1393 189 1452
rect 252 1393 305 1452
rect 175 1378 305 1393
rect 249 1240 305 1378
rect 409 1365 465 1510
rect 1012 1466 1068 1510
rect 938 1452 1068 1466
rect 938 1393 952 1452
rect 1015 1393 1068 1452
rect 938 1378 1068 1393
rect 353 1352 465 1365
rect 353 1293 366 1352
rect 429 1293 465 1352
rect 353 1280 465 1293
rect 409 1240 465 1280
rect 1012 1240 1068 1378
rect 1172 1365 1228 1510
rect 1823 1466 1879 1510
rect 1749 1452 1879 1466
rect 1749 1393 1763 1452
rect 1826 1393 1879 1452
rect 1749 1378 1879 1393
rect 1116 1352 1228 1365
rect 1116 1293 1129 1352
rect 1192 1293 1228 1352
rect 1116 1280 1228 1293
rect 1172 1240 1228 1280
rect 1823 1240 1879 1378
rect 1983 1365 2039 1510
rect 1927 1352 2039 1365
rect 1927 1293 1940 1352
rect 2003 1293 2039 1352
rect 1927 1280 2039 1293
rect 1983 1240 2039 1280
rect 249 1096 305 1140
rect 409 1096 465 1140
rect 1012 1096 1068 1140
rect 1172 1096 1228 1140
rect 1823 1096 1879 1140
rect 1983 1096 2039 1140
rect 249 635 305 679
rect 409 635 465 679
rect 1012 634 1068 678
rect 1172 634 1228 678
rect 1823 634 1879 678
rect 1983 634 2039 678
rect 249 491 305 535
rect 175 477 305 491
rect 175 418 189 477
rect 252 418 305 477
rect 175 403 305 418
rect 249 265 305 403
rect 409 390 465 535
rect 1012 490 1068 534
rect 938 476 1068 490
rect 938 417 952 476
rect 1015 417 1068 476
rect 938 402 1068 417
rect 353 377 465 390
rect 353 318 366 377
rect 429 318 465 377
rect 353 305 465 318
rect 409 265 465 305
rect 1012 264 1068 402
rect 1172 389 1228 534
rect 1823 490 1879 534
rect 1749 476 1879 490
rect 1749 417 1763 476
rect 1826 417 1879 476
rect 1749 402 1879 417
rect 1116 376 1228 389
rect 1116 317 1129 376
rect 1192 317 1228 376
rect 1116 304 1228 317
rect 1172 264 1228 304
rect 1823 264 1879 402
rect 1983 389 2039 534
rect 1927 376 2039 389
rect 1927 317 1940 376
rect 2003 317 2039 376
rect 1927 304 2039 317
rect 1983 264 2039 304
rect 249 121 305 165
rect 409 121 465 165
rect 1012 120 1068 164
rect 1172 120 1228 164
rect 1823 120 1879 164
rect 1983 120 2039 164
<< polycontact >>
rect 189 2364 252 2423
rect 952 2364 1015 2423
rect 366 2264 429 2323
rect 1763 2364 1826 2423
rect 1129 2264 1192 2323
rect 1940 2264 2003 2323
rect 189 1393 252 1452
rect 952 1393 1015 1452
rect 366 1293 429 1352
rect 1763 1393 1826 1452
rect 1129 1293 1192 1352
rect 1940 1293 2003 1352
rect 189 418 252 477
rect 952 417 1015 476
rect 366 318 429 377
rect 1763 417 1826 476
rect 1129 317 1192 376
rect 1940 317 2003 376
<< metal1 >>
rect 75 2845 639 2861
rect 838 2845 1402 2861
rect 1649 2845 2213 2861
rect -304 2802 -208 2817
rect 75 2815 2213 2845
rect 75 2802 190 2815
rect -304 2735 -289 2802
rect -222 2759 190 2802
rect 502 2759 953 2815
rect 1265 2759 1764 2815
rect 2076 2759 2213 2815
rect -222 2735 2213 2759
rect -304 2729 -208 2735
rect 75 2730 2213 2735
rect 75 2711 639 2730
rect 838 2711 1402 2730
rect 1649 2711 2213 2730
rect 171 2568 222 2711
rect 171 2494 174 2568
rect 220 2494 222 2568
rect 171 2492 222 2494
rect 334 2568 380 2579
rect 174 2483 220 2492
rect 334 2441 380 2494
rect 494 2568 540 2711
rect 494 2483 540 2494
rect 934 2568 985 2711
rect 934 2494 937 2568
rect 983 2494 985 2568
rect 934 2492 985 2494
rect 1097 2568 1143 2579
rect 937 2483 983 2492
rect 1097 2441 1143 2494
rect 1257 2568 1303 2711
rect 1257 2483 1303 2494
rect 1745 2568 1796 2711
rect 1745 2494 1748 2568
rect 1794 2494 1796 2568
rect 1745 2492 1796 2494
rect 1908 2568 1954 2579
rect 1748 2483 1794 2492
rect 1908 2441 1954 2494
rect 2068 2568 2114 2711
rect 2068 2483 2114 2494
rect 334 2437 443 2441
rect 1097 2437 1206 2441
rect 1908 2437 2017 2441
rect 2280 2437 2361 2451
rect 175 2423 264 2437
rect 175 2395 189 2423
rect 74 2364 189 2395
rect 252 2364 264 2423
rect 334 2395 883 2437
rect 938 2423 1027 2437
rect 938 2395 952 2423
rect 410 2391 952 2395
rect 74 2349 264 2364
rect 74 2301 120 2349
rect 355 2323 440 2334
rect 355 2301 366 2323
rect 74 2264 366 2301
rect 429 2264 440 2323
rect 74 2255 440 2264
rect 174 2198 220 2209
rect 334 2208 380 2209
rect 174 2044 220 2124
rect 321 2198 388 2208
rect 321 2124 334 2198
rect 380 2124 388 2198
rect 321 2110 388 2124
rect 494 2198 540 2391
rect 837 2364 952 2391
rect 1015 2364 1027 2423
rect 1097 2401 1402 2437
rect 1749 2427 1838 2437
rect 1097 2395 1314 2401
rect 1173 2391 1314 2395
rect 837 2349 1027 2364
rect 837 2301 883 2349
rect 1257 2345 1314 2391
rect 1370 2391 1402 2401
rect 1738 2423 1838 2427
rect 1738 2421 1763 2423
rect 1738 2395 1749 2421
rect 1370 2345 1380 2391
rect 1648 2365 1749 2395
rect 1648 2364 1763 2365
rect 1826 2364 1838 2423
rect 1908 2435 2426 2437
rect 1908 2395 2293 2435
rect 1984 2391 2293 2395
rect 1648 2349 1838 2364
rect 1118 2323 1203 2334
rect 1118 2301 1129 2323
rect 837 2264 1129 2301
rect 1192 2264 1203 2323
rect 837 2255 1203 2264
rect 1257 2333 1380 2345
rect 494 2113 540 2124
rect 937 2198 983 2209
rect 1097 2208 1143 2209
rect 937 2044 983 2124
rect 1084 2198 1151 2208
rect 1084 2124 1097 2198
rect 1143 2124 1151 2198
rect 1084 2110 1151 2124
rect 1257 2198 1303 2333
rect 1929 2323 2014 2334
rect 1599 2301 1681 2302
rect 1929 2301 1940 2323
rect 1599 2264 1940 2301
rect 2003 2264 2014 2323
rect 1599 2208 1615 2264
rect 1671 2255 2014 2264
rect 1671 2208 1681 2255
rect 1599 2197 1681 2208
rect 1748 2198 1794 2209
rect 1908 2208 1954 2209
rect 1257 2113 1303 2124
rect 1748 2044 1794 2124
rect 1895 2198 1962 2208
rect 1895 2124 1908 2198
rect 1954 2124 1962 2198
rect 1895 2110 1962 2124
rect 2068 2198 2114 2391
rect 2280 2379 2293 2391
rect 2349 2391 2426 2435
rect 2349 2379 2361 2391
rect 2280 2369 2361 2379
rect 2068 2113 2114 2124
rect -111 2028 -25 2042
rect 51 2037 667 2044
rect 814 2037 1430 2044
rect 1625 2037 2241 2044
rect 51 2028 2241 2037
rect -111 2027 2241 2028
rect -111 1962 -99 2027
rect -34 2017 2241 2027
rect -34 1969 118 2017
rect 587 1970 881 2017
rect 587 1969 667 1970
rect -34 1962 667 1969
rect -111 1961 667 1962
rect -111 1955 -25 1961
rect 51 1946 667 1961
rect 814 1969 881 1970
rect 1350 1970 1692 2017
rect 1350 1969 1430 1970
rect 814 1946 1430 1969
rect 1625 1969 1692 1970
rect 2161 1969 2241 2017
rect 1625 1946 2241 1969
rect -304 1871 -194 1872
rect 75 1871 639 1890
rect 838 1871 1402 1890
rect 1649 1871 2213 1890
rect -304 1851 2213 1871
rect -304 1784 -289 1851
rect -222 1844 2213 1851
rect -222 1788 190 1844
rect 502 1788 953 1844
rect 1265 1788 1764 1844
rect 2076 1788 2213 1844
rect -222 1784 2213 1788
rect -304 1756 2213 1784
rect 75 1740 639 1756
rect 838 1740 1402 1756
rect 1649 1740 2213 1756
rect 171 1597 222 1740
rect 171 1523 174 1597
rect 220 1523 222 1597
rect 171 1521 222 1523
rect 334 1597 380 1608
rect 174 1512 220 1521
rect 334 1470 380 1523
rect 494 1597 540 1740
rect 687 1625 765 1635
rect 687 1571 699 1625
rect 753 1621 765 1625
rect 753 1575 883 1621
rect 753 1571 765 1575
rect 687 1559 765 1571
rect 494 1512 540 1523
rect 334 1466 443 1470
rect 175 1452 264 1466
rect 175 1424 189 1452
rect 74 1393 189 1424
rect 252 1393 264 1452
rect 334 1424 639 1466
rect 410 1420 639 1424
rect 74 1378 264 1393
rect 74 1330 120 1378
rect 355 1352 440 1363
rect 355 1330 366 1352
rect 74 1293 366 1330
rect 429 1293 440 1352
rect 74 1284 440 1293
rect 174 1227 220 1238
rect 334 1237 380 1238
rect 174 1073 220 1153
rect 321 1227 388 1237
rect 321 1153 334 1227
rect 380 1153 388 1227
rect 321 1139 388 1153
rect 494 1227 540 1420
rect 593 1213 639 1420
rect 837 1424 883 1575
rect 934 1597 985 1740
rect 934 1523 937 1597
rect 983 1523 985 1597
rect 934 1521 985 1523
rect 1097 1597 1143 1608
rect 937 1512 983 1521
rect 1097 1470 1143 1523
rect 1257 1597 1303 1740
rect 1745 1597 1796 1740
rect 1893 1669 1971 1681
rect 1893 1615 1905 1669
rect 1959 1615 1971 1669
rect 1893 1603 1971 1615
rect 1257 1512 1303 1523
rect 1560 1573 1643 1588
rect 1560 1519 1574 1573
rect 1628 1519 1643 1573
rect 1745 1523 1748 1597
rect 1794 1523 1796 1597
rect 1745 1521 1796 1523
rect 1908 1597 1955 1603
rect 1954 1592 1955 1597
rect 2068 1597 2114 1740
rect 1560 1504 1643 1519
rect 1748 1512 1794 1521
rect 1097 1466 1206 1470
rect 938 1452 1027 1466
rect 938 1424 952 1452
rect 837 1393 952 1424
rect 1015 1393 1027 1452
rect 1097 1437 1402 1466
rect 1097 1424 1321 1437
rect 1173 1420 1321 1424
rect 837 1378 1027 1393
rect 1257 1383 1321 1420
rect 1375 1420 1402 1437
rect 1578 1424 1624 1504
rect 1908 1470 1954 1523
rect 2068 1512 2114 1523
rect 1908 1466 2017 1470
rect 1749 1452 1838 1466
rect 1749 1424 1763 1452
rect 1375 1383 1387 1420
rect 1257 1377 1387 1383
rect 1578 1393 1763 1424
rect 1826 1393 1838 1452
rect 1908 1424 2244 1466
rect 1984 1420 2244 1424
rect 1578 1378 1838 1393
rect 1118 1352 1203 1363
rect 816 1330 886 1332
rect 1118 1330 1129 1352
rect 816 1319 1129 1330
rect 816 1263 826 1319
rect 882 1293 1129 1319
rect 1192 1293 1203 1352
rect 882 1284 1203 1293
rect 1257 1330 1303 1377
rect 1929 1352 2014 1363
rect 1929 1330 1940 1352
rect 1257 1293 1940 1330
rect 2003 1293 2014 1352
rect 1257 1284 2014 1293
rect 882 1263 886 1284
rect 816 1251 886 1263
rect 937 1227 983 1238
rect 1097 1237 1143 1238
rect 593 1204 696 1213
rect 593 1154 630 1204
rect 494 1142 540 1153
rect 618 1150 630 1154
rect 684 1150 696 1204
rect 618 1141 696 1150
rect 937 1073 983 1153
rect 1084 1227 1151 1237
rect 1084 1153 1097 1227
rect 1143 1153 1151 1227
rect 1084 1139 1151 1153
rect 1257 1227 1303 1284
rect 1257 1142 1303 1153
rect 1748 1227 1794 1238
rect 1908 1237 1954 1238
rect 1748 1073 1794 1153
rect 1895 1227 1962 1237
rect 1895 1153 1908 1227
rect 1954 1153 1962 1227
rect 1895 1139 1962 1153
rect 2068 1227 2114 1420
rect 2198 1410 2244 1420
rect 2198 1364 2343 1410
rect 2068 1142 2114 1153
rect 51 1064 667 1073
rect 814 1064 1430 1073
rect 1625 1064 2241 1073
rect -110 1057 -29 1064
rect 51 1057 2241 1064
rect -110 1056 2241 1057
rect -110 991 -98 1056
rect -33 1046 2241 1056
rect -33 998 118 1046
rect 587 998 881 1046
rect 1350 998 1692 1046
rect 2161 998 2241 1046
rect -33 997 2241 998
rect -33 991 667 997
rect -110 990 667 991
rect -110 986 -29 990
rect 51 975 667 990
rect 814 975 1430 997
rect 1625 975 2241 997
rect 75 883 639 915
rect 838 883 1402 914
rect 1649 883 2213 914
rect -299 869 2213 883
rect -299 843 190 869
rect -299 775 -289 843
rect -222 813 190 843
rect 502 868 2213 869
rect 502 813 953 868
rect -222 812 953 813
rect 1265 812 1764 868
rect 2076 812 2213 868
rect -222 775 2213 812
rect -299 768 2213 775
rect -299 767 -208 768
rect -299 763 -210 767
rect 75 765 639 768
rect 171 622 222 765
rect 171 548 174 622
rect 220 548 222 622
rect 171 546 222 548
rect 334 622 380 633
rect 174 537 220 546
rect 334 495 380 548
rect 494 622 540 765
rect 838 764 1402 768
rect 1649 764 2213 768
rect 494 537 540 548
rect 934 621 985 764
rect 934 547 937 621
rect 983 547 985 621
rect 934 545 985 547
rect 1097 621 1143 632
rect 937 536 983 545
rect 749 514 824 526
rect 334 491 443 495
rect 175 477 264 491
rect 175 449 189 477
rect 74 418 189 449
rect 252 418 264 477
rect 334 449 639 491
rect 410 445 639 449
rect 749 460 758 514
rect 812 460 824 514
rect 1097 494 1143 547
rect 1257 621 1303 764
rect 1257 536 1303 547
rect 1745 621 1796 764
rect 1745 547 1748 621
rect 1794 547 1796 621
rect 1745 545 1796 547
rect 1908 621 1954 632
rect 1748 536 1794 545
rect 1908 494 1954 547
rect 2068 621 2114 764
rect 2068 536 2114 547
rect 1097 490 1206 494
rect 1908 490 2017 494
rect 749 448 824 460
rect 938 476 1027 490
rect 938 448 952 476
rect 74 403 264 418
rect 74 355 120 403
rect 355 377 440 388
rect 355 355 366 377
rect 74 318 366 355
rect 429 318 440 377
rect 74 309 440 318
rect 174 252 220 263
rect 334 262 380 263
rect 174 98 220 178
rect 321 252 388 262
rect 321 178 334 252
rect 380 178 388 252
rect 321 164 388 178
rect 494 252 540 445
rect 593 354 639 445
rect 762 417 952 448
rect 1015 417 1027 476
rect 1097 463 1402 490
rect 1097 448 1320 463
rect 1173 444 1320 448
rect 762 402 1027 417
rect 1257 409 1320 444
rect 1374 444 1402 463
rect 1749 476 1838 490
rect 1749 448 1763 476
rect 1374 409 1386 444
rect 1257 396 1386 409
rect 1648 417 1763 448
rect 1826 417 1838 476
rect 1908 455 2213 490
rect 1908 448 2125 455
rect 1984 444 2125 448
rect 1648 402 1838 417
rect 1118 376 1203 387
rect 1118 354 1129 376
rect 593 317 1129 354
rect 1192 317 1203 376
rect 593 308 1203 317
rect 494 167 540 178
rect 937 251 983 262
rect 1097 261 1143 262
rect -111 86 -18 96
rect 51 86 667 98
rect 937 97 983 177
rect 1084 251 1151 261
rect 1084 177 1097 251
rect 1143 177 1151 251
rect 1084 163 1151 177
rect 1257 251 1303 396
rect 1648 380 1694 402
rect 2068 401 2125 444
rect 2179 444 2213 455
rect 2179 401 2189 444
rect 2068 389 2189 401
rect 1586 373 1694 380
rect 1586 319 1599 373
rect 1653 354 1694 373
rect 1929 376 2014 387
rect 1929 354 1940 376
rect 1653 319 1940 354
rect 1586 317 1940 319
rect 2003 317 2014 376
rect 1586 308 2014 317
rect 1586 305 1655 308
rect 1257 166 1303 177
rect 1748 251 1794 262
rect 1908 261 1954 262
rect 1748 97 1794 177
rect 1895 251 1962 261
rect 1895 177 1908 251
rect 1954 177 1962 251
rect 1895 163 1962 177
rect 2068 251 2114 389
rect 2068 166 2114 177
rect 814 86 1430 97
rect 1625 86 2241 97
rect -111 19 -99 86
rect -32 71 2241 86
rect -32 23 118 71
rect 587 70 2241 71
rect 587 23 881 70
rect -32 22 881 23
rect 1350 22 1692 70
rect 2161 22 2241 70
rect -32 19 2241 22
rect -111 7 -18 19
rect 51 0 667 19
rect 814 -1 1430 19
rect 1625 -1 2241 19
<< via1 >>
rect -289 2735 -222 2802
rect 1314 2345 1370 2401
rect 1749 2365 1763 2421
rect 1763 2365 1805 2421
rect 1615 2208 1671 2264
rect 2293 2379 2349 2435
rect -99 1962 -34 2027
rect -289 1784 -222 1851
rect 699 1571 753 1625
rect 1905 1615 1959 1669
rect 1574 1519 1628 1573
rect 1321 1383 1375 1437
rect 826 1263 882 1319
rect 630 1150 684 1204
rect -98 991 -33 1056
rect -289 775 -222 843
rect 758 460 812 514
rect 1320 409 1374 463
rect 2125 401 2179 455
rect 1599 319 1653 373
rect -99 19 -32 86
<< metal2 >>
rect -304 2802 -208 2817
rect -304 2735 -289 2802
rect -222 2735 -208 2802
rect -304 2729 -208 2735
rect -289 1872 -222 2729
rect 1749 2430 2180 2456
rect 1738 2421 2180 2430
rect 1304 2401 1380 2410
rect 697 2345 1314 2401
rect 1370 2345 1380 2401
rect 1738 2365 1749 2421
rect 1805 2400 2180 2421
rect 1805 2365 1819 2400
rect 1738 2349 1819 2365
rect -111 2027 -25 2042
rect -111 1962 -99 2027
rect -34 1962 -25 2027
rect -111 1955 -25 1962
rect -304 1851 -194 1872
rect -304 1784 -289 1851
rect -222 1784 -194 1851
rect -304 1756 -194 1784
rect -289 883 -222 1756
rect -99 1064 -32 1955
rect 697 1659 753 2345
rect 1304 2333 1380 2345
rect 1599 2293 1681 2302
rect 1599 2264 1960 2293
rect 1599 2208 1615 2264
rect 1671 2237 1960 2264
rect 1671 2208 1681 2237
rect 1599 2197 1681 2208
rect 1904 1681 1960 2237
rect 1893 1669 1971 1681
rect 697 1635 754 1659
rect 687 1625 765 1635
rect 687 1571 699 1625
rect 753 1571 765 1625
rect 1893 1615 1905 1669
rect 1959 1615 1971 1669
rect 1893 1603 1971 1615
rect 687 1559 765 1571
rect 1560 1574 1643 1588
rect 1560 1518 1573 1574
rect 1629 1518 1643 1574
rect 1560 1504 1643 1518
rect 1303 1437 1387 1449
rect 1303 1383 1321 1437
rect 1375 1383 1387 1437
rect 1303 1377 1387 1383
rect 1320 1346 1377 1377
rect 816 1319 886 1332
rect 816 1263 826 1319
rect 882 1263 1002 1319
rect 816 1251 886 1263
rect 616 1204 699 1214
rect 616 1191 630 1204
rect 548 1150 630 1191
rect 684 1150 699 1204
rect 548 1140 699 1150
rect 548 1135 660 1140
rect -110 1056 -29 1064
rect -110 991 -98 1056
rect -33 991 -29 1056
rect -110 986 -29 991
rect -299 843 -210 883
rect -299 775 -289 843
rect -222 775 -210 843
rect -299 763 -210 775
rect -99 96 -32 986
rect 548 640 604 1135
rect 548 584 813 640
rect 757 526 813 584
rect 749 514 824 526
rect 749 460 758 514
rect 812 460 824 514
rect 749 448 824 460
rect 946 464 1002 1263
rect 1321 1127 1377 1346
rect 1321 1071 1654 1127
rect 1303 464 1386 466
rect 946 463 1386 464
rect 946 409 1320 463
rect 1374 409 1386 463
rect 946 408 1386 409
rect 1303 396 1386 408
rect 1598 380 1654 1071
rect 2124 460 2180 2400
rect 2280 2435 2361 2451
rect 2280 2379 2293 2435
rect 2349 2379 2361 2435
rect 2280 2369 2361 2379
rect 2293 1583 2349 2369
rect 2284 1574 2360 1583
rect 2284 1518 2293 1574
rect 2349 1518 2360 1574
rect 2284 1506 2360 1518
rect 2112 455 2189 460
rect 2112 401 2125 455
rect 2179 401 2189 455
rect 2112 389 2189 401
rect 1586 373 1655 380
rect 1586 319 1599 373
rect 1653 319 1655 373
rect 1586 305 1655 319
rect -111 86 -18 96
rect -111 19 -99 86
rect -32 19 -18 86
rect -111 7 -18 19
<< via2 >>
rect 1573 1573 1629 1574
rect 1573 1519 1574 1573
rect 1574 1519 1628 1573
rect 1628 1519 1629 1573
rect 1573 1518 1629 1519
rect 2293 1518 2349 1574
<< metal3 >>
rect 1560 1574 1643 1588
rect 2284 1574 2360 1583
rect 1560 1518 1573 1574
rect 1629 1518 2293 1574
rect 2349 1518 2360 1574
rect 1560 1504 1643 1518
rect 2284 1506 2360 1518
<< labels >>
flabel metal1 93 2328 93 2328 0 FreeSans 480 0 0 0 Ri-1
port 0 nsew
flabel metal1 1098 2792 1098 2792 0 FreeSans 480 0 0 0 VDD
port 1 nsew
flabel metal1 1102 2005 1102 2005 0 FreeSans 480 0 0 0 VSS
port 2 nsew
flabel metal1 2322 1385 2322 1385 0 FreeSans 480 0 0 0 Q
port 3 nsew
flabel metal1 2396 2412 2396 2412 0 FreeSans 480 0 0 0 QB
port 4 nsew
flabel metal1 93 1350 93 1350 0 FreeSans 480 0 0 0 Ci
port 5 nsew
flabel metal1 92 377 92 377 0 FreeSans 480 0 0 0 Ri
port 6 nsew
flabel nsubdiffcont 344 841 344 841 0 FreeSans 320 0 0 0 NAND_3.VDD
flabel psubdiffcont 353 49 353 49 0 FreeSans 320 0 0 0 NAND_3.VSS
flabel metal1 104 427 104 427 0 FreeSans 480 0 0 0 NAND_3.B
flabel metal1 107 329 107 329 0 FreeSans 480 0 0 0 NAND_3.A
flabel metal1 606 473 606 473 0 FreeSans 480 0 0 0 NAND_3.OUT
flabel nsubdiffcont 344 1816 344 1816 0 FreeSans 320 0 0 0 NAND_2.VDD
flabel psubdiffcont 353 1024 353 1024 0 FreeSans 320 0 0 0 NAND_2.VSS
flabel metal1 104 1402 104 1402 0 FreeSans 480 0 0 0 NAND_2.B
flabel metal1 107 1304 107 1304 0 FreeSans 480 0 0 0 NAND_2.A
flabel metal1 606 1448 606 1448 0 FreeSans 480 0 0 0 NAND_2.OUT
flabel nsubdiffcont 344 2787 344 2787 0 FreeSans 320 0 0 0 NAND_0.VDD
flabel psubdiffcont 353 1995 353 1995 0 FreeSans 320 0 0 0 NAND_0.VSS
flabel metal1 104 2373 104 2373 0 FreeSans 480 0 0 0 NAND_0.B
flabel metal1 107 2275 107 2275 0 FreeSans 480 0 0 0 NAND_0.A
flabel metal1 606 2419 606 2419 0 FreeSans 480 0 0 0 NAND_0.OUT
flabel nsubdiffcont 1107 840 1107 840 0 FreeSans 320 0 0 0 NAND_6.VDD
flabel psubdiffcont 1116 48 1116 48 0 FreeSans 320 0 0 0 NAND_6.VSS
flabel metal1 867 426 867 426 0 FreeSans 480 0 0 0 NAND_6.B
flabel metal1 870 328 870 328 0 FreeSans 480 0 0 0 NAND_6.A
flabel metal1 1369 472 1369 472 0 FreeSans 480 0 0 0 NAND_6.OUT
flabel nsubdiffcont 1107 1816 1107 1816 0 FreeSans 320 0 0 0 NAND_5.VDD
flabel psubdiffcont 1116 1024 1116 1024 0 FreeSans 320 0 0 0 NAND_5.VSS
flabel metal1 867 1402 867 1402 0 FreeSans 480 0 0 0 NAND_5.B
flabel metal1 870 1304 870 1304 0 FreeSans 480 0 0 0 NAND_5.A
flabel metal1 1369 1448 1369 1448 0 FreeSans 480 0 0 0 NAND_5.OUT
flabel nsubdiffcont 1107 2787 1107 2787 0 FreeSans 320 0 0 0 NAND_1.VDD
flabel psubdiffcont 1116 1995 1116 1995 0 FreeSans 320 0 0 0 NAND_1.VSS
flabel metal1 867 2373 867 2373 0 FreeSans 480 0 0 0 NAND_1.B
flabel metal1 870 2275 870 2275 0 FreeSans 480 0 0 0 NAND_1.A
flabel metal1 1369 2419 1369 2419 0 FreeSans 480 0 0 0 NAND_1.OUT
flabel nsubdiffcont 1918 840 1918 840 0 FreeSans 320 0 0 0 NAND_7.VDD
flabel psubdiffcont 1927 48 1927 48 0 FreeSans 320 0 0 0 NAND_7.VSS
flabel metal1 1678 426 1678 426 0 FreeSans 480 0 0 0 NAND_7.B
flabel metal1 1681 328 1681 328 0 FreeSans 480 0 0 0 NAND_7.A
flabel metal1 2180 472 2180 472 0 FreeSans 480 0 0 0 NAND_7.OUT
flabel nsubdiffcont 1918 1816 1918 1816 0 FreeSans 320 0 0 0 NAND_8.VDD
flabel psubdiffcont 1927 1024 1927 1024 0 FreeSans 320 0 0 0 NAND_8.VSS
flabel metal1 1678 1402 1678 1402 0 FreeSans 480 0 0 0 NAND_8.B
flabel metal1 1681 1304 1681 1304 0 FreeSans 480 0 0 0 NAND_8.A
flabel metal1 2180 1448 2180 1448 0 FreeSans 480 0 0 0 NAND_8.OUT
flabel nsubdiffcont 1918 2787 1918 2787 0 FreeSans 320 0 0 0 NAND_4.VDD
flabel psubdiffcont 1927 1995 1927 1995 0 FreeSans 320 0 0 0 NAND_4.VSS
flabel metal1 1678 2373 1678 2373 0 FreeSans 480 0 0 0 NAND_4.B
flabel metal1 1681 2275 1681 2275 0 FreeSans 480 0 0 0 NAND_4.A
flabel metal1 2180 2419 2180 2419 0 FreeSans 480 0 0 0 NAND_4.OUT
<< end >>
