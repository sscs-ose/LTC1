* NGSPICE file created from 7b_divider_magic_flat.ext - technology: gf180mcuC

.subckt pex_7b_divider_magic VDD LD D2_7 Q1 D2_6 Q2 D2_5 D2_4 Q3 Q4 D2_3 D2_2 Q5 D2_1 Q6 Q7 CLK VSS OUT1 P2
X0 a_2749_684# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A VDD.t150 VDD.t144 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1 VSS CLK.t0 a_16065_9774# VSS.t667 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B a_1209_7469# VDD.t143 VDD.t142 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X3 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B a_15865_3363# VSS.t729 VSS.t172 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X4 DFF_magic_0.tg_magic_0.IN CLK.t1 DFF_magic_0.tg_magic_3.OUT VSS.t666 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X5 7b_counter_0.3_inp_AND_magic_0.C Q3.t3 a_23207_5815# VDD.t2284 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X6 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t11 VSS.t728 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X7 a_1559_n1526# D2_4.t0 p2_gen_magic_0.xnor_magic_3.OUT VDD.t2045 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X8 a_30365_3514# P2.t6 a_30365_4922# VDD.t2219 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X9 VDD a_14556_n8142# p3_gen_magic_0.3_inp_AND_magic_0.B VDD.t1792 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X10 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT VDD.t1800 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X11 VDD Q3.t4 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT VDD.t2287 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X12 a_6725_2092# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B a_6725_684# VDD.t422 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X13 VDD p3_gen_magic_0.xnor_magic_1.B.t3 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT VDD.t2455 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X14 a_2749_2092# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B a_2749_684# VDD.t147 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X15 a_16065_2253# D2_3.t0 VSS.t1448 VSS.t625 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X16 VDD 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A a_17405_10149# VDD.t1033 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X17 p2_gen_magic_0.xnor_magic_1.OUT p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT a_1541_n4081# VDD.t1150 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X18 VDD a_23258_1746# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B VDD.t471 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X19 a_21381_3524# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B VSS.t53 VSS.t52 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X20 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A a_19841_9774# VDD.t170 VDD.t169 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X21 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT VDD.t1093 VDD.t1092 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X22 p3_gen_magic_0.xnor_magic_4.OUT Q2.t3 a_5054_n6471# VSS.t1406 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X23 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_6.t0 VDD.t1363 VDD.t1362 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X24 a_1541_n3597# D2_1.t0 p2_gen_magic_0.xnor_magic_1.OUT VDD.t1149 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X25 7b_counter_0.MDFF_5.LD a_29512_8496.t9 VDD.t1195 VDD.t1189 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X26 a_12174_n8579# p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p3_gen_magic_0.AND2_magic_1.A VDD.t1415 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X27 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A a_15865_4557# VSS.t93 VSS.t92 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X28 a_11279_8697# 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B a_11191_10149# VDD.t165 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X29 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B a_5185_2253# VDD.t1646 VDD.t1645 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X30 VDD a_19841_9774# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A VDD.t166 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X31 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t9 VDD.t1199 VDD.t1198 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X32 a_12931_7470# D2_2.t0 VSS.t1099 VSS.t619 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X33 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B a_1209_2253# VDD.t1748 VDD.t1747 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X34 a_18891_6886# 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_19152_5956# VDD.t1750 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X35 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A LD.t9 VSS.t1056 VSS.t1055 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X36 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_17405_8741# VDD.t577 VDD.t575 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X37 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5054_n1042# VDD.t770 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X38 a_26038_4932# 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_26126_3480# VDD.t776 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X39 a_1209_8579# D2_7.t0 VDD.t1958 VDD.t1957 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X40 VSS mux_magic_0.IN2.t5 divide_by_2_0.tg_magic_2.IN VSS.t1243 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X41 a_24059_4877# 7b_counter_0.MDFF_7.tspc2_magic_0.D VSS.t1353 VSS.t1352 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X42 7b_counter_0.MDFF_1.tspc2_magic_0.D a_17405_2092# VDD.t2328 VDD.t2327 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X43 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT CLK.t2 VSS.t665 VSS.t664 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X44 VDD 7b_counter_0.DFF_magic_0.Q.t6 DFF_magic_0.D VDD.t2047 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X45 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q1.t3 VDD.t2059 VDD.t2058 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X46 mux_magic_0.AND2_magic_0.A D2_1.t1 VDD.t1301 VDD.t1300 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X47 VDD 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t3 a_23560_3728# VDD.t1467 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X48 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK.t3 VDD.t2530 VDD.t2529 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X49 VSS p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.P3.t1 VSS.t30 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X50 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT CLK.t4 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t2 VSS.t663 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X51 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK.t5 VDD.t2528 VDD.t2527 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X52 VDD 7b_counter_0.MDFF_4.LD.t9 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A VDD.t1476 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X53 VDD 7b_counter_0.DFF_magic_0.Q.t7 7b_counter_0.DFF_magic_0.D VDD.t2050 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X54 a_19307_6886# 7b_counter_0.MDFF_6.tspc2_magic_0.CLK VSS.t1019 VSS.t1018 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X55 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t10 VSS.t900 VSS.t899 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X56 a_7215_10149# 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B a_7303_8697# VDD.t1442 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X57 a_4496_10093# 7b_counter_0.MDFF_3.tspc2_magic_0.D VDD.t1455 VDD.t1453 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X58 a_4651_9163# 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t3 VSS.t1164 VSS.t1163 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X59 a_23985_7877# 7b_counter_0.3_inp_AND_magic_0.B VDD.t1757 VDD.t1755 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X60 VSS 7b_counter_0.MDFF_4.LD.t11 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A VSS.t901 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X61 VSS CLK.t6 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VSS.t660 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X62 VSS 7b_counter_0.MDFF_4.LD.t12 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A VSS.t904 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X63 p3_gen_magic_0.3_inp_AND_magic_0.C a_16186_n8142# VSS.t1008 VSS.t1007 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X64 VSS D2_5.t0 a_1409_3363# VSS.t584 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X65 VSS divide_by_2_1.tg_magic_3.CLK.t3 divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT VSS.t1147 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X66 VSS a_11279_1124# 7b_counter_0.MDFF_4.tspc2_magic_0.D VSS.t708 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X67 VDD D2_5.t1 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT VDD.t2719 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X68 p2_gen_magic_0.AND2_magic_1.A D2_5.t2 a_12174_n3597# VDD.t441 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X69 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q3.t5 VSS.t1337 VSS.t1336 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X70 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t13 VSS.t908 VSS.t907 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X71 VDD 7b_counter_0.MDFF_4.LD.t14 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A VDD.t1479 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X72 a_15865_1059# 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A VDD.t592 VDD.t591 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X73 VDD 7b_counter_0.MDFF_4.LD.t15 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A VDD.t1482 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X74 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT Q6.t3 VDD.t2162 VDD.t2161 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X75 a_9059_n1973# p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_0.OUT VSS.t1010 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X76 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t16 VDD.t1486 VDD.t1485 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X77 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT VDD.t1743 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X78 a_1209_3363# D2_5.t3 VDD.t2723 VDD.t2722 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X79 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q2.t4 VDD.t2410 VDD.t2409 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X80 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t17 VDD.t1488 VDD.t1487 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X81 VDD 7b_counter_0.MDFF_4.LD.t18 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A VDD.t1489 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X82 a_22991_5815# Q1.t4 VDD.t2061 VDD.t2060 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X83 VDD divide_by_2_0.tg_magic_3.CLK.t5 divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT VDD.t1811 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X84 DFF_magic_0.tg_magic_2.IN DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT DFF_magic_0.tg_magic_2.OUT VDD.t1002 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X85 VDD a_12387_9730# 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A VDD.t1015 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X86 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK CLK.t7 VDD.t2526 VDD.t2525 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X87 a_2749_2092# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B a_2749_684# VDD.t372 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X88 a_4235_3947# 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t4 a_4496_4877# VDD.t2449 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X89 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t6 VSS.t1386 VSS.t1385 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X90 a_6725_684# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B a_6725_2092# VDD.t421 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X91 VDD a_5185_1059# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A VDD.t1688 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X92 VSS 7b_counter_0.MDFF_0.QB.t4 a_1409_4557# VSS.t1426 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X93 a_5185_7469# D2_7.t1 VDD.t1960 VDD.t1959 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X94 VDD 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A a_1209_6275# VDD.t1705 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X95 VSS p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT P2.t1 VSS.t1380 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X96 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A LD.t10 VSS.t1058 VSS.t1057 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X97 7b_counter_0.3_inp_AND_magic_0.VOUT 7b_counter_0.3_inp_AND_magic_0.VOUT 7b_counter_0.3_inp_AND_magic_0.VOUT VDD.t792 pfet_03v3 ad=0.493p pd=3.12u as=1.97p ps=12.5u w=1.12u l=0.56u
X98 a_15865_3363# 7b_counter_0.MDFF_4.LD.t19 a_16065_3363# VSS.t909 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X99 7b_counter_0.DFF_magic_0.tg_magic_0.IN 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.OUT VDD.t795 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X100 VSS 7b_counter_0.MDFF_5.LD.t10 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A VSS.t744 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X101 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.CLK.t6 VDD.t1815 VDD.t1814 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X102 a_8643_n1526# D2_2.t1 p2_gen_magic_0.xnor_magic_0.OUT VDD.t458 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X103 a_12387_8536# 7b_counter_0.MDFF_5.LD.t11 a_12931_8580# VSS.t747 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X104 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1559_n1042# VDD.t2046 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X105 p2_gen_magic_0.xnor_magic_1.OUT Q7.t3 a_1541_n3150# VSS.t845 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X106 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK CLK.t8 VSS.t655 VSS.t654 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X107 a_8825_1669# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t3 7b_counter_0.MDFF_4.QB.t3 VSS.t1514 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X108 VSS CLK.t9 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t1 VSS.t657 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X109 a_2749_8740# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B VSS.t48 VSS.t47 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X110 VDD p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5054_n5540# VDD.t75 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X111 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t12 VSS.t749 VSS.t748 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X112 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t6 VDD.t2021 VDD.t2020 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X113 a_16065_2253# 7b_counter_0.MDFF_4.LD.t20 a_15865_2253# VSS.t910 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X114 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B a_15865_3363# VDD.t1175 VDD.t1174 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X115 a_8411_3319# 7b_counter_0.MDFF_4.LD.t21 VDD.t1493 VDD.t1492 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X116 VDD 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A a_11191_684# VDD.t350 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X117 a_1409_1059# Q4.t3 VSS.t976 VSS.t975 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X118 VDD 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A a_12387_4513# VDD.t1437 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X119 a_11279_3480# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B a_11191_4932# VDD.t1144 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X120 VDD 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A a_11191_5901# VDD.t360 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X121 VDD OR_magic_2.A.t6 a_30365_4922# VDD.t2329 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X122 a_11292_n2115# p2_gen_magic_0.xnor_magic_4.OUT VDD.t773 VDD.t771 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X123 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.D VDD.t368 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X124 a_21381_3524# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B a_21381_4932# VDD.t78 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X125 VSS D2_7.t2 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT VSS.t1123 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X126 VSS CLK.t10 DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VSS.t652 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X127 p2_gen_magic_0.3_inp_AND_magic_0.A a_11292_n2115# VSS.t181 VSS.t180 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X128 VDD Q6.t4 a_21504_5904# VDD.t2163 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X129 a_15865_4557# 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A a_16065_4557# VSS.t160 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X130 VDD 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A a_26038_684# VDD.t1096 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X131 a_12387_9730# 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A a_12931_9774# VSS.t686 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X132 VDD p2_gen_magic_0.3_inp_AND_magic_0.C.t3 a_13353_n2115# VDD.t2714 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X133 a_5185_2253# D2_5.t4 VDD.t2725 VDD.t2724 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X134 a_13769_n2115# p2_gen_magic_0.3_inp_AND_magic_0.B a_13553_n2115# VSS.t689 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X135 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q1.t5 VSS.t1194 VSS.t1193 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X136 VSS a_26126_1124# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t0 VSS.t409 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X137 VDD 7b_counter_0.MDFF_4.LD.t22 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A VDD.t1494 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X138 VSS a_22150_1124# Q4.t0 VSS.t692 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X139 a_9212_739# 7b_counter_0.MDFF_4.tspc2_magic_0.D VSS.t1029 VSS.t1028 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X140 p3_gen_magic_0.3_inp_AND_magic_0.VOUT a_13353_n6613# VDD.t1134 VDD.t1132 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X141 VSS p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VSS.t725 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X142 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t7 7b_counter_0.DFF_magic_0.D VSS.t1173 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X143 VDD OR_magic_1.VOUT.t3 divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT VDD.t2495 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X144 a_24536_3947# a_24059_4877# a_23560_3728# VSS.t1355 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X145 VSS divide_by_2_0.tg_magic_1.IN.t12 divide_by_2_0.tg_magic_0.IN VSS.t860 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X146 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT VDD.t1799 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X147 VDD p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t12 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN VDD.t2241 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X148 VDD p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT a_1541_n4081# VDD.t808 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X149 VSS p2_gen_magic_0.xnor_magic_3.OUT.t4 a_11708_n2115# VSS.t1290 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X150 VSS 7b_counter_0.MDFF_0.tspc2_magic_0.D a_4235_3947# VSS.t457 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X151 mux_magic_0.IN2 divide_by_2_0.tg_magic_3.IN.t18 VDD.t11 VDD.t10 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X152 mux_magic_0.AND2_magic_0.A D2_1.t2 VDD.t1303 VDD.t1302 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X153 VSS a_11279_6341# 7b_counter_0.MDFF_5.tspc2_magic_0.D VSS.t460 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X154 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT VDD.t287 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X155 p3_gen_magic_0.3_inp_AND_magic_0.C a_16186_n8142# VDD.t1725 VDD.t1724 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X156 a_14756_n8142# p3_gen_magic_0.AND2_magic_1.A a_14556_n8142# VSS.t868 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X157 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.OUT VDD.t564 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X158 LD a_27567_8496.t9 VSS.t731 VSS.t730 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X159 LD a_27567_8496.t10 VDD.t1177 VDD.t1176 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X160 a_11492_n6613# p3_gen_magic_0.xnor_magic_4.OUT a_11708_n6613# VSS.t230 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X161 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B a_19841_8580# VDD.t1125 VDD.t1124 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X162 VSS D2_3.t1 a_16065_2253# VSS.t615 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X163 a_15865_7470# D2_1.t3 VDD.t1305 VDD.t1304 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X164 VDD Q1.t6 a_8643_n1526# VDD.t1731 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X165 7b_counter_0.MDFF_4.LD a_31440_8496.t9 VDD.t21 VDD.t20 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X166 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B a_23258_1746# VDD.t470 VDD.t469 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X167 VSS 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A a_21381_3524# VSS.t52 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X168 7b_counter_0.3_inp_AND_magic_0.C Q3.t6 a_23207_5815# VDD.t2290 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X169 VSS D2_6.t1 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT VSS.t836 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X170 a_17405_10149# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B a_17405_8741# VDD.t575 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X171 a_5452_n7648# p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_5.OUT.t4 VSS.t1009 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X172 a_5185_1059# 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A VDD.t574 VDD.t573 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X173 VDD 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A a_22062_684# VDD.t847 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X174 a_20041_8580# D2_1.t4 VSS.t792 VSS.t791 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X175 VDD 7b_counter_0.MDFF_4.LD.t23 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A VDD.t1497 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X176 VDD a_29512_8496.t10 7b_counter_0.MDFF_5.LD.t7 VDD.t1191 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X177 VDD Q4.t4 a_1209_1059# VDD.t1647 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X178 VDD divide_by_2_1.tg_magic_3.IN.t18 mux_magic_0.IN1.t5 VDD.t109 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X179 VSS p3_gen_magic_0.xnor_magic_3.OUT.t5 a_11708_n6613# VSS.t230 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X180 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_3.OUT VDD.t133 VDD.t132 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X181 VDD LD.t11 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A VDD.t1831 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X182 VDD D2_1.t5 p3_gen_magic_0.xnor_magic_1.B VDD.t1306 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X183 VDD 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A a_22062_684# VDD.t476 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X184 VDD CLK.t11 DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD.t2539 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X185 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A a_15865_6276# VDD.t2207 VDD.t2206 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X186 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_3.CLK.t7 divide_by_2_0.tg_magic_2.IN VSS.t1039 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X187 a_17405_2092# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B a_17405_684# VDD.t2218 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X188 VSS D2_2.t2 a_12931_7470# VSS.t612 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X189 p3_gen_magic_0.xnor_magic_6.OUT p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT a_8523_n8579# VDD.t65 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X190 VSS D2_3.t2 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT VSS.t1451 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X191 VSS D2_1.t6 mux_magic_0.AND2_magic_0.A VSS.t793 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X192 DFF_magic_0.D DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT DFF_magic_0.tg_magic_3.OUT VDD.t941 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X193 a_17405_7309# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_17405_5901# VDD.t629 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X194 VDD Q4.t5 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT VDD.t1650 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X195 VDD LD.t12 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A VDD.t1834 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X196 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A LD.t13 VDD.t1838 VDD.t1837 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X197 VDD 7b_counter_0.MDFF_4.QB.t4 a_12387_552# VDD.t1432 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X198 a_19841_4557# 7b_counter_0.MDFF_1.tspc2_magic_0.Q VDD.t652 VDD.t651 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X199 VDD 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A a_27234_4513# VDD.t1763 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X200 VSS p3_gen_magic_0.xnor_magic_1.B.t4 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT VSS.t1440 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X201 a_26126_3480# 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_26038_4932# VDD.t775 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X202 VDD 7b_counter_0.MDFF_0.tspc2_magic_0.D a_4496_4877# VDD.t876 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X203 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT CLK.t12 VDD.t2538 VDD.t2537 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X204 VSS p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VSS.t722 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X205 VSS CLK.t13 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VSS.t649 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X206 DFF_magic_0.tg_magic_2.IN OR_magic_2.A.t7 VDD.t2333 VDD.t2332 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X207 VDD D2_1.t7 mux_magic_0.AND2_magic_0.A VDD.t1309 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X208 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT Q6.t5 VSS.t1260 VSS.t1259 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X209 VSS Q5.t3 7b_counter_0.3_inp_AND_magic_0.A VSS.t122 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X210 a_20041_9774# 7b_counter_0.MDFF_6.tspc2_magic_0.Q VSS.t151 VSS.t150 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X211 DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_3.CLK.t6 DFF_magic_0.D.t6 VSS.t1498 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X212 VSS 7b_counter_0.MDFF_5.LD.t13 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A VSS.t750 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X213 VDD p3_gen_magic_0.3_inp_AND_magic_0.A a_13353_n6613# VDD.t902 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X214 a_23793_5904# Q5.t4 7b_counter_0.3_inp_AND_magic_0.A VDD.t220 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X215 OR_magic_2.A DFF_magic_0.tg_magic_2.OUT VDD.t1012 VDD.t1011 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X216 VSS divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_1.IN.t1 VSS.t82 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X217 VSS D2_2.t3 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT VSS.t1102 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X218 a_8825_1669# a_8713_1625# VSS.t244 VSS.t243 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X219 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t24 VSS.t912 VSS.t911 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X220 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t25 VSS.t913 VSS.t899 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X221 DFF_magic_0.tg_magic_0.IN DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT DFF_magic_0.tg_magic_3.OUT VDD.t762 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X222 divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.CLK.t4 VSS.t1151 VSS.t1150 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X223 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t26 VSS.t915 VSS.t914 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X224 VDD a_15865_2253# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B VDD.t334 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X225 a_8411_3319# D2_6.t2 VDD.t1365 VDD.t1364 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X226 VSS 7b_counter_0.MDFF_4.LD.t27 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A VSS.t901 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X227 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT VDD.t1742 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X228 a_7215_10149# 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B a_7303_8697# VDD.t1441 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X229 a_2749_8740# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B a_2749_10148# VDD.t69 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X230 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t28 VDD.t1501 VDD.t1500 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X231 VDD divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_1.IN.t4 VDD.t129 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X232 a_11191_10149# 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B a_11279_8697# VDD.t164 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X233 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT VDD.t1029 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X234 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B a_8411_8536# VDD.t447 VDD.t446 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X235 VDD D2_4.t1 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT VDD.t2254 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X236 mux_magic_0.AND2_magic_0.A D2_1.t8 VDD.t1312 VDD.t1300 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X237 VDD 7b_counter_0.MDFF_4.LD.t29 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A VDD.t1502 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X238 a_11191_684# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_11279_1124# VDD.t451 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X239 divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT OR_magic_1.VOUT.t4 VDD.t2499 VDD.t2498 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X240 a_11292_n2115# p2_gen_magic_0.xnor_magic_0.OUT a_11492_n2115# VSS.t180 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X241 VDD Q2.t5 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT VDD.t2411 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X242 a_5036_n8579# p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_5.OUT VDD.t759 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X243 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT D2_5.t5 VSS.t1535 VSS.t1534 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X244 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t12 VSS.t1556 VSS.t1555 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X245 a_13769_n2115# p2_gen_magic_0.3_inp_AND_magic_0.B a_13553_n2115# VSS.t689 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X246 a_24401_7877# 7b_counter_0.3_inp_AND_magic_0.B a_24185_7877# VSS.t1022 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X247 VDD a_1209_9773# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A VDD.t685 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X248 a_32616_n2458# mux_magic_0.IN2.t6 VDD.t2145 VDD.t2144 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X249 7b_counter_0.MDFF_6.tspc2_magic_0.Q 7b_counter_0.MDFF_6.QB.t4 VDD.t2247 VDD.t2246 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X250 VSS D2_4.t2 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT VSS.t1309 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X251 a_2749_4932# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A VDD.t677 VDD.t676 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X252 a_22991_5815# Q1.t7 VDD.t2065 VDD.t2064 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X253 a_5470_n1973# p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_4.OUT VSS.t158 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X254 VDD LD.t14 a_1209_7469# VDD.t1839 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X255 a_14556_n3644# p2_gen_magic_0.AND2_magic_1.A a_14756_n3644# VSS.t1031 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X256 VDD divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_1.IN.t8 VDD.t834 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X257 VSS p2_gen_magic_0.xnor_magic_3.OUT.t5 a_11708_n2115# VSS.t1290 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X258 a_9412_739# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t4 a_9212_739# VDD.t2708 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X259 a_23207_5815# Q2.t6 a_22991_5815# VDD.t2414 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X260 7b_counter_0.DFF_magic_0.tg_magic_2.IN 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_2.OUT VDD.t331 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X261 VDD CLK.t14 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD.t2534 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X262 VDD 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t8 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD.t2022 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X263 VSS 7b_counter_0.MDFF_5.LD.t14 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A VSS.t753 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X264 VDD D2_6.t3 a_8411_3319# VDD.t1366 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X265 a_15865_7470# 7b_counter_0.MDFF_5.LD.t15 VDD.t1201 VDD.t1200 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X266 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT Q6.t6 VDD.t2167 VDD.t2166 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X267 a_19152_5956# 7b_counter_0.MDFF_6.tspc2_magic_0.D VDD.t209 VDD.t207 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X268 7b_counter_0.DFF_magic_0.D 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.OUT VDD.t367 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X269 VDD p2_gen_magic_0.xnor_magic_5.OUT a_16186_n3644# VDD.t212 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X270 a_21381_4932# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A VDD.t860 VDD.t855 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X271 a_20171_6886# 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 7b_counter_0.MDFF_6.QB.t3 VSS.t1017 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X272 divide_by_2_0.tg_magic_2.IN mux_magic_0.IN2.t7 VDD.t2147 VDD.t2146 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X273 p3_gen_magic_0.AND2_magic_1.A Q4.t6 a_12174_n7648# VSS.t977 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X274 a_26038_684# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A VDD.t1099 VDD.t1096 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X275 a_26038_684# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B a_26126_1124# VDD.t1065 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X276 a_23672_3947# a_23560_3728# VSS.t1497 VSS.t1496 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X277 a_12387_3319# 7b_counter_0.MDFF_4.LD.t30 VDD.t1506 VDD.t1505 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X278 a_22062_684# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B a_22150_1124# VDD.t476 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X279 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT VSS.t683 VSS.t682 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X280 VDD LD.t15 a_1209_2253# VDD.t1842 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X281 VDD p3_gen_magic_0.xnor_magic_0.OUT a_11292_n6613# VDD.t1071 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X282 P2 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT VDD.t2375 VDD.t2374 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X283 VDD D2_4.t3 a_27234_3319# VDD.t2257 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X284 a_2749_10148# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A VDD.t694 VDD.t69 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X285 VDD LD.t16 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A VDD.t1834 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X286 VSS a_12387_5769# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A VSS.t200 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X287 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_4.t4 VSS.t1313 VSS.t1312 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X288 mux_magic_0.IN2 divide_by_2_0.tg_magic_3.IN.t19 VDD.t13 VDD.t12 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X289 VSS 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t5 a_9689_1669# VSS.t1515 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X290 a_12387_1746# 7b_counter_0.MDFF_4.LD.t31 a_12931_2253# VSS.t918 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X291 VDD Q3.t7 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT VDD.t2299 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X292 DFF_magic_0.tg_magic_0.IN DFF_magic_0.tg_magic_1.IN.t12 VDD.t55 VDD.t54 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X293 a_17405_10149# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A VDD.t1036 VDD.t863 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X294 VDD a_8713_1625# 7b_counter_0.MDFF_4.QB.t1 VDD.t461 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X295 a_24059_4877# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t4 a_24259_4877# VDD.t1470 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X296 7b_counter_0.3_inp_AND_magic_0.A Q5.t5 a_23793_5904# VDD.t221 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X297 a_1541_n8579# p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.OUT VDD.t370 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X298 7b_counter_0.MDFF_1.tspc2_magic_0.Q 7b_counter_0.MDFF_1.QB.t4 VDD.t84 VDD.t83 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X299 VDD D2_1.t9 a_19841_8580# VDD.t1313 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X300 VSS DFF_magic_0.tg_magic_2.OUT OR_magic_2.A.t1 VSS.t526 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X301 VDD 7b_counter_0.MDFF_5.LD.t16 a_15865_7470# VDD.t1202 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X302 a_32616_n1264# mux_magic_0.AND2_magic_0.A a_32816_n1264# VSS.t523 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X303 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q2.t7 VSS.t1408 VSS.t1407 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X304 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_2749_7308# VDD.t950 VDD.t949 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X305 7b_counter_0.3_inp_AND_magic_0.VOUT a_23985_7877# VDD.t1760 VDD.t1758 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X306 a_12931_1059# 7b_counter_0.MDFF_4.QB.t5 VSS.t873 VSS.t872 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X307 VDD D2_3.t3 a_15865_2253# VDD.t2465 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X308 VSS D2_1.t10 a_20041_8580# VSS.t796 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X309 p3_gen_magic_0.xnor_magic_4.OUT D2_3.t4 a_5054_n6024# VDD.t401 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X310 DFF_magic_0.tg_magic_3.OUT CLK.t15 DFF_magic_0.tg_magic_0.IN VSS.t648 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X311 a_9412_739# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t6 a_9212_739# VDD.t2709 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X312 mux_magic_0.IN1 divide_by_2_1.tg_magic_3.IN.t19 VDD.t113 VDD.t112 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X313 VSS D2_2.t4 a_9059_n6471# VSS.t1105 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X314 VSS Q3.t8 a_27778_1059# VSS.t1341 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X315 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t32 VDD.t1508 VDD.t1507 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X316 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A LD.t17 VDD.t1848 VDD.t1847 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X317 a_8523_n7648# p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT VSS.t46 VSS.t45 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X318 VSS divide_by_2_1.tg_magic_3.CLK.t5 divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT VSS.t1152 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X319 Q7 a_6725_7308# VSS.t70 VSS.t69 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X320 VDD Q2.t8 a_5054_n1526# VDD.t293 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X321 a_27234_3319# 7b_counter_0.MDFF_4.LD.t33 VDD.t1510 VDD.t1509 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X322 a_19152_1223# a_18891_1669# a_19307_1669# VSS.t63 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X323 VDD 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A a_19841_4557# VDD.t1718 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X324 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN VSS.t721 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X325 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_7.t3 VDD.t1962 VDD.t1961 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X326 p3_gen_magic_0.xnor_magic_5.OUT D2_7.t4 a_5036_n8095# VDD.t758 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X327 a_32616_n2458# D2_1.t11 a_32816_n2458# VSS.t799 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X328 VDD a_23560_3728# 7b_counter_0.MDFF_7.QB.t2 VDD.t2685 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X329 a_24401_7877# 7b_counter_0.3_inp_AND_magic_0.B a_24185_7877# VSS.t1022 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X330 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_6.t4 VSS.t840 VSS.t839 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X331 VDD CLK.t16 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD.t2531 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X332 VSS 7b_counter_0.3_inp_AND_magic_0.VOUT a_24003_10051# VSS.t416 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X333 a_12387_5769# 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A VDD.t561 VDD.t560 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X334 p3_gen_magic_0.AND2_magic_1.A p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_12174_n8579# VDD.t1414 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X335 VSS 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_20041_9774# VSS.t147 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X336 a_17405_5901# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_17405_7309# VDD.t628 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X337 a_16186_n3644# p2_gen_magic_0.xnor_magic_5.OUT a_16386_n3644# VSS.t119 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X338 VSS a_8411_3319# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B VSS.t174 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X339 VDD Q5.t6 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT VDD.t222 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X340 VDD Q6.t7 a_5036_n3597# VDD.t262 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X341 a_12931_8580# 7b_counter_0.MDFF_5.LD.t17 a_12387_8536# VSS.t756 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X342 VDD DFF_magic_0.tg_magic_2.OUT OR_magic_2.A.t4 VDD.t1008 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X343 p3_gen_magic_0.xnor_magic_3.OUT Q3.t9 a_1559_n6471# VSS.t1344 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X344 VDD 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A a_15865_9774# VDD.t499 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X345 a_7215_10149# 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A VDD.t516 VDD.t513 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X346 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_6.t5 VDD.t1370 VDD.t1369 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X347 VDD 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A a_11191_4932# VDD.t520 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X348 divide_by_2_0.tg_magic_2.IN mux_magic_0.IN2.t8 VSS.t1247 VSS.t1246 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X349 DFF_magic_0.tg_magic_1.IN CLK.t17 DFF_magic_0.tg_magic_2.OUT VSS.t647 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X350 a_27234_1746# 7b_counter_0.MDFF_4.LD.t34 a_27778_2253# VSS.t919 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X351 VDD divide_by_2_1.tg_magic_3.CLK.t6 divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT VDD.t1990 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X352 VDD a_8411_3319# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B VDD.t339 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X353 a_12387_552# 7b_counter_0.MDFF_4.QB.t6 VDD.t2019 VDD.t2018 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X354 a_12387_4513# Q5.t7 VDD.t226 VDD.t225 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X355 a_27778_1059# Q3.t10 VSS.t1346 VSS.t1345 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X356 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t35 VSS.t920 VSS.t914 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X357 Q5 a_6725_2092# VDD.t1032 VDD.t421 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X358 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B a_12387_8536# VDD.t569 VDD.t568 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X359 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT VDD.t665 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X360 divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT OR_magic_2.VOUT.t3 VSS.t378 VSS.t377 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X361 a_11279_8697# 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A VSS.t153 VSS.t152 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X362 a_18891_1669# 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_19152_739# VDD.t963 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X363 VSS a_8411_4513# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A VSS.t509 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X364 p3_gen_magic_0.xnor_magic_3.OUT D2_4.t5 a_1559_n6024# VDD.t408 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X365 a_12931_9774# 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A a_12387_9730# VSS.t685 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X366 p3_gen_magic_0.xnor_magic_6.OUT Q5.t8 a_8523_n7648# VSS.t125 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X367 VDD p3_gen_magic_0.AND2_magic_1.A a_14556_n8142# VDD.t1418 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X368 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT CLK.t18 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN VSS.t646 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X369 VDD 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 7b_counter_0.DFF_magic_0.Q.t5 VDD.t615 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X370 VDD OR_magic_1.VOUT.t5 divide_by_2_1.tg_magic_3.CLK VDD.t2500 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X371 a_5054_n1973# p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT VSS.t403 VSS.t402 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X372 7b_counter_0.3_inp_AND_magic_0.B Q6.t8 VSS.t1262 VSS.t1261 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X373 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN P2.t7 VDD.t2221 VDD.t2220 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X374 VDD 7b_counter_0.MDFF_4.LD.t36 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A VDD.t1511 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X375 VDD D2_2.t5 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT VDD.t1927 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X376 VDD p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.P3.t5 VDD.t43 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X377 VDD Q6.t9 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT VDD.t2170 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X378 VSS Q7.t4 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT VSS.t846 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X379 a_23258_552# 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A VDD.t307 VDD.t306 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X380 VSS Q5.t9 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT VSS.t126 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X381 VDD 7b_counter_0.MDFF_4.QB.t7 7b_counter_0.MDFF_4.tspc2_magic_0.Q VDD.t1429 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X382 divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.CLK.t8 VDD.t1817 VDD.t1816 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X383 VDD DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_1.IN.t5 VDD.t1048 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X384 p3_gen_magic_0.3_inp_AND_magic_0.VOUT CLK.t19 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT VSS.t645 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X385 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_2.IN VDD.t330 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X386 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q3.t11 VDD.t2292 VDD.t2291 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X387 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A a_12387_9730# VDD.t1014 VDD.t1013 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X388 VDD 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A a_19841_9774# VDD.t259 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X389 p3_gen_magic_0.3_inp_AND_magic_0.A p3_gen_magic_0.3_inp_AND_magic_0.A p3_gen_magic_0.3_inp_AND_magic_0.A VDD.t905 pfet_03v3 ad=0.493p pd=3.12u as=1.97p ps=12.5u w=1.12u l=0.56u
X390 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t18 VDD.t1206 VDD.t1205 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X391 VDD 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t5 VDD.t803 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X392 a_5385_6275# 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A a_5185_6275# VSS.t329 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X393 a_23352_n6798# p3_gen_magic_0.P3.t6 VSS.t886 VSS.t885 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X394 VDD 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A a_17405_684# VDD.t199 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X395 a_15865_1059# 7b_counter_0.MDFF_1.QB.t5 VDD.t86 VDD.t85 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X396 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_8643_n5540# VDD.t981 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X397 VDD D2_1.t12 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT VDD.t1316 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X398 VSS 7b_counter_0.MDFF_1.tspc2_magic_0.D a_18891_1669# VSS.t532 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X399 VDD 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_19152_6440# VDD.t204 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X400 VDD mux_magic_0.IN1.t6 a_32616_n1264# VDD.t2351 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X401 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t9 VDD.t2026 VDD.t2025 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X402 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT CLK.t20 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t1 VSS.t644 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X403 VDD Q6.t10 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT VDD.t2173 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X404 a_8713_6842# a_9212_5956# a_9689_6886# VSS.t364 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X405 divide_by_2_0.tg_magic_3.CLK OR_magic_2.VOUT.t4 VDD.t729 VDD.t728 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X406 a_17405_3524# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B a_17405_4932# VDD.t160 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X407 VSS 7b_counter_0.MDFF_7.QB.t4 7b_counter_0.MDFF_7.tspc2_magic_0.Q VSS.t0 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X408 7b_counter_0.MDFF_5.LD a_29512_8496.t11 VSS.t738 VSS.t737 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X409 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A a_1209_6275# VSS.t1004 VSS.t1003 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X410 VDD CLK.t21 a_12387_3319# VDD.t2542 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X411 7b_counter_0.MDFF_5.LD a_29512_8496.t12 VDD.t1188 VDD.t1187 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X412 a_19841_3363# 7b_counter_0.MDFF_4.LD.t37 a_20041_3363# VSS.t921 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X413 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT divide_by_2_1.tg_magic_1.IN.t8 VDD.t438 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X414 a_27234_3319# D2_4.t6 VDD.t2261 VDD.t2260 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X415 OUT1 a_34156_n2297# VDD.t440 VDD.t48 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X416 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t13 VDD.t2245 VDD.t2244 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X417 a_23352_n6798# p3_gen_magic_0.P3.t7 a_23352_n5390# VDD.t1456 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X418 a_9689_1669# a_9212_739# a_8713_1625# VSS.t701 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X419 VDD a_1209_4557# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A VDD.t707 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X420 VSS 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A a_17405_3524# VSS.t94 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X421 VDD 7b_counter_0.MDFF_5.LD.t19 a_12387_6963# VDD.t1207 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X422 VSS p3_gen_magic_0.xnor_magic_1.OUT.t4 a_16386_n8142# VSS.t35 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X423 VSS CLK.t22 DFF_magic_0.tg_magic_3.CLK.t1 VSS.t641 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X424 a_17405_8741# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B VSS.t451 VSS.t324 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X425 a_5385_7469# LD.t18 a_5185_7469# VSS.t1059 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X426 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_2749_2092# VSS.t259 VSS.t107 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X427 VDD LD.t19 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A VDD.t1849 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X428 a_24259_4877# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t5 a_24059_4877# VDD.t1471 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X429 7b_counter_0.MDFF_3.tspc2_magic_0.Q 7b_counter_0.MDFF_3.QB VSS.t323 VSS.t322 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X430 a_12174_n8095# Q4.t7 VDD.t1653 VDD.t636 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X431 VDD p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1559_n5540# VDD.t580 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X432 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT divide_by_2_0.tg_magic_0.IN VDD.t954 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X433 a_1559_n1973# p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT VSS.t1190 VSS.t1189 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X434 divide_by_2_1.tg_magic_3.IN OR_magic_1.VOUT.t6 divide_by_2_1.tg_magic_1.IN.t11 VSS.t1472 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X435 p2_gen_magic_0.3_inp_AND_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t7 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT VSS.t1387 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X436 a_11191_10149# 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A VDD.t284 VDD.t277 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X437 VSS CLK.t23 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK VSS.t638 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X438 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B a_1209_7469# VSS.t88 VSS.t87 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X439 a_14556_n3644# p2_gen_magic_0.xnor_magic_6.OUT VDD.t870 VDD.t869 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X440 a_19841_4557# 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A a_20041_4557# VSS.t1006 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X441 VDD 7b_counter_0.3_inp_AND_magic_0.C a_23985_7877# VDD.t31 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X442 VSS 7b_counter_0.MDFF_4.QB.t8 a_12931_1059# VSS.t1167 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X443 VDD LD.t20 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A VDD.t1852 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X444 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t8 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.t1 VSS.t1388 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X445 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_3.OUT VDD.t1047 VDD.t1046 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X446 a_27778_1059# 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A a_27234_552# VSS.t304 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X447 VDD p3_gen_magic_0.xnor_magic_3.OUT.t6 a_11292_n6613# VDD.t452 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X448 a_21381_8741# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B a_21381_10149# VDD.t171 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X449 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_3.CLK.t7 divide_by_2_1.tg_magic_2.IN VSS.t1155 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X450 a_23802_1059# 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A a_23258_552# VSS.t162 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X451 VDD DFF_magic_0.tg_magic_3.CLK.t7 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD.t2693 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X452 a_11708_n6613# p3_gen_magic_0.xnor_magic_4.OUT a_11492_n6613# VSS.t260 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X453 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_4.t7 VDD.t2263 VDD.t2262 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X454 VDD 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A a_11191_10149# VDD.t277 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X455 a_21504_5904# Q6.t11 VDD.t2177 VDD.t2176 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X456 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A a_5185_1059# VSS.t995 VSS.t994 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X457 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q2.t9 VDD.t2418 VDD.t2417 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X458 a_11708_n6613# p3_gen_magic_0.xnor_magic_4.OUT a_11492_n6613# VSS.t260 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X459 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t9 VDD.t2385 VDD.t2384 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X460 a_2749_4932# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B a_2749_3524# VDD.t181 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X461 VDD 7b_counter_0.MDFF_5.QB.t4 a_12387_5769# VDD.t924 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X462 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t13 VDD.t2750 VDD.t2749 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X463 VDD D2_3.t5 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT VDD.t2468 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X464 VSS a_12387_3319# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B VSS.t205 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X465 VDD 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A a_27234_552# VDD.t585 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X466 VDD OR_magic_2.VOUT.t5 divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT VDD.t730 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X467 7b_counter_0.MDFF_0.tspc2_magic_0.Q 7b_counter_0.MDFF_0.QB.t5 VDD.t2442 VDD.t2441 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X468 a_1957_n7648# p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_1.OUT.t1 VSS.t444 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X469 7b_counter_0.DFF_magic_0.tg_magic_2.IN 7b_counter_0.DFF_magic_0.Q.t8 VDD.t2054 VDD.t2053 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X470 divide_by_2_0.tg_magic_1.IN OR_magic_2.VOUT.t6 divide_by_2_0.tg_magic_3.IN.t3 VSS.t379 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X471 VDD p2_gen_magic_0.xnor_magic_0.OUT a_11292_n2115# VDD.t1736 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X472 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.CLK.t9 VSS.t1041 VSS.t1040 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X473 VDD a_19841_3363# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B VDD.t433 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X474 VDD OR_magic_2.A.t8 DFF_magic_0.tg_magic_2.IN VDD.t2334 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X475 a_2749_684# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B a_2749_2092# VDD.t371 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X476 a_23802_2253# D2_4.t8 VSS.t1315 VSS.t1314 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X477 VDD a_1209_1059# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A VDD.t121 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X478 VSS D2_7.t5 a_5452_n3150# VSS.t1126 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X479 VDD p3_gen_magic_0.P3.t8 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN VDD.t1457 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X480 VDD mux_magic_0.AND2_magic_0.A a_32616_n1264# VDD.t994 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X481 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t10 VDD.t2028 VDD.t2027 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X482 VSS a_7303_3480# Q6.t0 VSS.t273 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X483 VSS p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t14 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN VSS.t869 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X484 VDD D2_2.t6 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT VDD.t1930 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X485 VSS a_12387_4513# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A VSS.t703 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X486 a_17405_5901# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A VDD.t2214 VDD.t2211 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X487 a_18891_1669# 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_19152_739# VDD.t962 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X488 VDD a_12387_3319# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B VDD.t1068 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X489 7b_counter_0.MDFF_4.LD a_31440_8496.t10 VSS.t14 VSS.t13 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X490 a_1209_6275# 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A a_1409_6275# VSS.t1002 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X491 a_16186_n8142# p3_gen_magic_0.xnor_magic_5.OUT.t5 VDD.t105 VDD.t104 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X492 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT Q4.t8 VDD.t1655 VDD.t1654 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X493 7b_counter_0.MDFF_4.LD a_31440_8496.t11 VDD.t23 VDD.t22 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X494 divide_by_2_1.tg_magic_3.CLK OR_magic_1.VOUT.t7 VDD.t2504 VDD.t2503 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X495 VDD 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A a_11191_5901# VDD.t357 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X496 VDD p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD.t1168 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X497 VDD OR_magic_2.VOUT.t7 divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT VDD.t733 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X498 VSS a_4496_4393# a_5515_3947# VSS.t467 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X499 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_15865_7470# VSS.t699 VSS.t194 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X500 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q3.t12 VDD.t2294 VDD.t2293 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X501 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_3.OUT VSS.t545 VSS.t544 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X502 VDD 7b_counter_0.MDFF_0.QB.t6 a_1209_4557# VDD.t2443 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X503 a_12931_2253# 7b_counter_0.MDFF_4.LD.t38 a_12387_1746# VSS.t922 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X504 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_3.CLK.t8 divide_by_2_1.tg_magic_3.IN.t11 VSS.t1156 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X505 a_17405_4932# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A VDD.t162 VDD.t156 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X506 a_5515_9163# 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t4 7b_counter_0.MDFF_3.QB VSS.t1165 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X507 a_8643_n1973# p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT VSS.t239 VSS.t238 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X508 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_3.OUT VDD.t1045 VDD.t1044 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X509 a_17405_8741# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B a_17405_10149# VDD.t863 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X510 VDD D2_7.t6 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT VDD.t1963 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X511 7b_counter_0.DFF_magic_0.tg_magic_2.IN 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_2.OUT VDD.t329 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X512 mux_magic_0.IN2 divide_by_2_0.tg_magic_3.IN.t20 VSS.t9 VSS.t8 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X513 p2_gen_magic_0.xnor_magic_1.OUT D2_1.t13 a_1541_n3597# VDD.t1150 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X514 DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK.t24 VSS.t637 VSS.t636 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X515 a_8523_n8095# Q5.t10 VDD.t228 VDD.t227 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X516 p2_gen_magic_0.xnor_magic_5.OUT p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT a_5036_n4081# VDD.t399 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X517 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_3.OUT VDD.t802 VDD.t801 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X518 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_3.t6 VSS.t1455 VSS.t1454 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X519 a_1209_7469# LD.t21 a_1409_7469# VSS.t1060 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X520 a_2749_5900# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A VDD.t430 VDD.t427 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X521 a_16186_n3644# p2_gen_magic_0.xnor_magic_1.OUT.t5 VDD.t2405 VDD.t2404 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X522 VDD Q1.t8 a_12387_9730# VDD.t2066 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X523 a_8411_8536# 7b_counter_0.MDFF_5.LD.t20 a_8955_8580# VSS.t757 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X524 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT CLK.t25 VDD.t2546 VDD.t2545 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X525 a_32616_n1264# mux_magic_0.IN1.t7 VDD.t2355 VDD.t2354 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X526 VDD 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t11 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD.t2029 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X527 divide_by_2_0.tg_magic_0.IN OR_magic_2.VOUT.t8 divide_by_2_0.tg_magic_3.OUT VSS.t380 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X528 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B a_1209_8579# VDD.t323 VDD.t322 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X529 VSS a_27234_3319# 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B VSS.t245 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X530 a_20171_6886# a_19152_6440# VSS.t265 VSS.t264 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X531 a_9689_6886# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t3 VSS.t473 VSS.t472 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X532 VDD LD.t22 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A VDD.t1852 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X533 divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT OR_magic_1.VOUT.t8 VDD.t2506 VDD.t2505 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X534 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A a_27234_552# VDD.t545 VDD.t544 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X535 VDD OR_magic_1.VOUT.t9 divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT VDD.t2507 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X536 VDD 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A a_8411_4513# VDD.t600 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X537 VSS 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A a_6725_7308# VSS.t278 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X538 VDD 7b_counter_0.MDFF_7.tspc2_magic_0.Q a_23258_552# VDD.t725 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X539 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.IN.t3 VDD.t437 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X540 VSS mux_magic_0.IN1.t8 divide_by_2_1.tg_magic_2.IN VSS.t1368 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X541 VDD mux_magic_0.IN1.t9 divide_by_2_1.tg_magic_2.IN VDD.t2356 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X542 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_2.t7 VDD.t1934 VDD.t1933 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X543 a_1209_1059# 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A VDD.t815 VDD.t814 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X544 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_2.t8 VSS.t1109 VSS.t1108 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X545 a_5185_1059# 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A a_5385_1059# VSS.t299 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X546 VDD DFF_magic_0.D.t14 a_29512_8496.t3 VDD.t2117 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X547 VDD CLK.t26 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD.t2552 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X548 a_4235_9163# 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t5 a_4496_10093# VDD.t2010 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X549 a_8411_9730# 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A a_8955_9774# VSS.t188 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X550 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q7.t5 VDD.t1377 VDD.t1376 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X551 VDD a_12387_5769# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A VDD.t404 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X552 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT CLK.t27 VSS.t635 VSS.t634 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X553 VDD a_8411_9730# 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A VDD.t380 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X554 VSS a_27234_4513# 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A VSS.t340 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X555 a_5385_2253# LD.t23 a_5185_2253# VSS.t1061 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X556 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B a_1209_3363# VDD.t292 VDD.t291 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X557 divide_by_2_1.tg_magic_0.IN OR_magic_1.VOUT.t10 divide_by_2_1.tg_magic_3.OUT VSS.t1473 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X558 p2_gen_magic_0.3_inp_AND_magic_0.VOUT a_13353_n2115# VSS.t687 VSS.t401 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X559 p2_gen_magic_0.xnor_magic_0.OUT Q1.t9 a_8643_n1973# VSS.t1195 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X560 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT Q5.t11 VDD.t230 VDD.t229 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X561 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A LD.t24 VDD.t1858 VDD.t1857 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X562 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A LD.t25 VDD.t1860 VDD.t1859 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X563 a_12387_552# 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A VDD.t2383 VDD.t2382 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X564 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B a_1209_2253# VSS.t1012 VSS.t156 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X565 a_21381_10149# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A VDD.t177 VDD.t173 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X566 VDD 7b_counter_0.MDFF_4.LD.t39 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A VDD.t1514 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X567 a_6725_684# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A VDD.t1697 VDD.t1693 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X568 a_6725_7308# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B VSS.t277 VSS.t276 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X569 VDD p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD.t1165 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X570 a_12590_n3150# p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p2_gen_magic_0.AND2_magic_1.A VSS.t343 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X571 a_2749_7308# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B VSS.t540 VSS.t47 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X572 a_14756_n8142# p3_gen_magic_0.xnor_magic_6.OUT VSS.t496 VSS.t495 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X573 VDD p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT a_5036_n8579# VDD.t1728 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X574 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t40 VDD.t1518 VDD.t1517 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X575 VDD 7b_counter_0.MDFF_4.LD.t41 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A VDD.t1519 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X576 VDD a_7303_3480# Q6.t2 VDD.t526 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X577 VDD 7b_counter_0.MDFF_4.LD.t42 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A VDD.t1479 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X578 p2_gen_magic_0.xnor_magic_0.OUT D2_2.t9 a_8643_n1526# VDD.t457 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X579 a_13553_n6613# p3_gen_magic_0.3_inp_AND_magic_0.B a_13769_n6613# VSS.t471 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X580 VDD.t1062 VDD.t1061 VDD.t1062 VDD.t865 pfet_03v3 ad=0.493p pd=3.12u as=0 ps=0 w=1.12u l=0.56u
X581 divide_by_2_1.tg_magic_3.CLK OR_magic_1.VOUT.t11 VDD.t2511 VDD.t2510 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X582 VDD 7b_counter_0.MDFF_4.LD.t43 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A VDD.t1482 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X583 VDD D2_4.t9 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT VDD.t2264 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X584 VDD a_27234_1746# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B VDD.t466 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X585 a_15865_7470# 7b_counter_0.MDFF_5.LD.t21 a_16065_7470# VSS.t758 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X586 a_2749_3524# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B a_2749_4932# VDD.t180 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X587 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t44 VDD.t1526 VDD.t1485 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X588 p3_gen_magic_0.P3 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT VSS.t29 VSS.t28 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X589 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK.t28 VSS.t633 VSS.t632 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X590 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t45 VDD.t1527 VDD.t1487 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X591 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t11 VDD.t2692 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X592 a_16065_6276# 7b_counter_0.MDFF_6.QB.t5 VSS.t1303 VSS.t1302 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X593 VDD p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t15 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN VDD.t1421 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X594 divide_by_2_1.tg_magic_3.OUT OR_magic_1.VOUT.t12 divide_by_2_1.tg_magic_0.IN VSS.t1474 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X595 VDD a_4496_4393# 7b_counter_0.MDFF_0.QB.t3 VDD.t899 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X596 VDD p3_gen_magic_0.P3.t9 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN VDD.t1460 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X597 VDD 7b_counter_0.DFF_magic_0.Q.t9 7b_counter_0.DFF_magic_0.tg_magic_2.IN VDD.t2055 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X598 VSS p3_gen_magic_0.3_inp_AND_magic_0.C.t3 a_13769_n6613# VSS.t470 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X599 VSS 7b_counter_0.MDFF_3.QB a_1409_9773# VSS.t319 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X600 DFF_magic_0.tg_magic_2.OUT DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT DFF_magic_0.tg_magic_1.IN.t11 VDD.t2202 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X601 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_3.OUT VDD.t800 VDD.t799 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X602 7b_counter_0.3_inp_AND_magic_0.C Q3.t13 a_23207_5815# VDD.t2284 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X603 a_1409_8579# LD.t26 a_1209_8579# VSS.t1062 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X604 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK.t29 VDD.t2551 VDD.t2550 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X605 VDD p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD.t1162 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X606 a_13553_n2115# p2_gen_magic_0.3_inp_AND_magic_0.A a_13353_n2115# VSS.t400 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X607 VSS 7b_counter_0.MDFF_5.LD.t22 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A VSS.t744 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X608 VDD divide_by_2_0.tg_magic_1.IN.t13 divide_by_2_0.tg_magic_0.IN VDD.t1404 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X609 a_32616_n1264# mux_magic_0.AND2_magic_0.A VDD.t993 VDD.t992 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X610 a_6725_2092# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B a_6725_684# VDD.t420 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X611 DFF_magic_0.D 7b_counter_0.DFF_magic_0.Q.t10 VSS.t1192 VSS.t1191 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X612 VDD Q3.t14 a_1559_n1526# VDD.t603 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X613 VSS 7b_counter_0.MDFF_5.LD.t23 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A VSS.t761 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X614 a_12174_n4081# p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT VDD.t670 VDD.t669 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X615 VSS a_11279_3480# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t0 VSS.t708 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X616 VDD 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A a_21381_10149# VDD.t173 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X617 VSS p3_gen_magic_0.3_inp_AND_magic_0.C.t4 a_13769_n6613# VSS.t471 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X618 a_2749_2092# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B a_2749_684# VDD.t147 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X619 VSS OR_magic_2.A.t9 a_30365_3514# VSS.t1357 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X620 VDD DFF_magic_0.tg_magic_3.CLK.t8 DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD.t2696 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X621 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t24 VSS.t765 VSS.t764 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X622 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.B.t5 VDD.t2459 VDD.t2458 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X623 DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_3.CLK.t9 DFF_magic_0.D.t7 VSS.t1499 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X624 Q3 a_21381_3524# VDD.t82 VDD.t79 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X625 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t25 VSS.t766 VSS.t748 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X626 VSS D2_5.t6 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT VSS.t1536 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X627 a_1409_6275# Q6.t12 VSS.t1264 VSS.t1263 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X628 7b_counter_0.MDFF_3.tspc2_magic_0.D a_2749_8740# VDD.t72 VDD.t71 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X629 VSS a_31440_8496.t12 7b_counter_0.MDFF_4.LD.t3 VSS.t15 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X630 VDD a_31440_8496.t13 7b_counter_0.MDFF_4.LD.t4 VDD.t24 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X631 a_9412_5956# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t4 a_9212_5956# VDD.t908 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X632 VDD D2_7.t7 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT VDD.t1966 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X633 VSS p3_gen_magic_0.3_inp_AND_magic_0.C.t5 a_13769_n6613# VSS.t470 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X634 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.IN.t1 VDD.t563 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X635 VDD Q7.t6 a_1541_n3597# VDD.t808 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X636 divide_by_2_0.tg_magic_3.CLK OR_magic_2.VOUT.t9 VSS.t382 VSS.t381 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X637 a_1209_4557# 7b_counter_0.MDFF_0.QB.t7 VDD.t2447 VDD.t2446 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X638 Q1 a_21381_8741# VSS.t285 VSS.t284 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X639 P2 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT VSS.t1379 VSS.t1378 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X640 VDD 7b_counter_0.MDFF_4.LD.t46 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A VDD.t1528 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X641 VDD 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A a_5185_1059# VDD.t570 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X642 a_12387_6963# D2_2.t10 VDD.t1936 VDD.t1935 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X643 VSS 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A a_2749_2092# VSS.t89 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X644 VDD 7b_counter_0.MDFF_4.LD.t47 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A VDD.t1489 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X645 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_3.CLK.t9 divide_by_2_1.tg_magic_3.OUT VSS.t1157 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X646 7b_counter_0.MDFF_3.QB 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t6 a_5515_9163# VSS.t1166 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X647 a_22062_684# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A VDD.t850 VDD.t847 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X648 VDD 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A a_5185_6275# VDD.t640 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X649 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t48 VDD.t1534 VDD.t1533 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X650 7b_counter_0.MDFF_1.tspc2_magic_0.D a_17405_2092# VDD.t2326 VDD.t2325 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X651 VDD 7b_counter_0.MDFF_4.LD.t49 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A VDD.t1494 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X652 a_12174_n7648# p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT VSS.t866 VSS.t865 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X653 a_1409_7469# CLK.t30 VSS.t631 VSS.t630 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X654 7b_counter_0.MDFF_6.tspc2_magic_0.D a_17405_7309# VDD.t632 VDD.t631 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X655 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN CLK.t31 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT VSS.t629 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X656 a_8955_8580# D2_2.t11 VSS.t1111 VSS.t1110 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X657 divide_by_2_0.tg_magic_2.IN divide_by_2_0.tg_magic_3.CLK.t10 divide_by_2_0.tg_magic_3.IN.t13 VSS.t1042 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X658 VDD D2_6.t6 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT VDD.t1371 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X659 a_13353_n2115# p2_gen_magic_0.3_inp_AND_magic_0.A a_13553_n2115# VSS.t401 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X660 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q7.t7 VSS.t850 VSS.t849 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X661 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_12387_1746# VDD.t413 VDD.t412 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X662 a_1209_2253# LD.t27 a_1409_2253# VSS.t1063 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X663 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A LD.t28 VDD.t1861 VDD.t1859 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X664 VDD 7b_counter_0.MDFF_4.LD.t50 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A VDD.t1537 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X665 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A a_15865_4557# VDD.t155 VDD.t154 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X666 divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT OR_magic_1.VOUT.t13 VDD.t2513 VDD.t2512 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X667 a_8411_4513# 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A VDD.t599 VDD.t598 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X668 VDD LD.t29 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A VDD.t1862 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X669 VDD CLK.t32 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD.t2547 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X670 a_16386_n8142# p3_gen_magic_0.xnor_magic_1.OUT.t5 VSS.t39 VSS.t38 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X671 a_15865_8580# CLK.t33 VDD.t2556 VDD.t2555 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X672 a_4235_9163# 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t7 a_4496_10093# VDD.t2011 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X673 a_8939_n3150# p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_6.OUT VSS.t430 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X674 VDD 7b_counter_0.MDFF_4.LD.t51 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A VDD.t1497 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X675 7b_counter_0.MDFF_1.tspc2_magic_0.Q 7b_counter_0.MDFF_1.QB.t6 VDD.t88 VDD.t87 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X676 divide_by_2_1.tg_magic_2.IN divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.IN.t2 VDD.t99 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X677 a_5385_1059# 7b_counter_0.MDFF_0.tspc2_magic_0.Q VSS.t443 VSS.t442 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X678 VDD LD.t30 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A VDD.t1865 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X679 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN P2.t8 VSS.t1284 VSS.t1283 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X680 VSS a_26126_3480# 7b_counter_0.MDFF_7.tspc2_magic_0.D VSS.t409 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X681 a_8955_9774# 7b_counter_0.MDFF_5.tspc2_magic_0.Q VSS.t358 VSS.t357 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X682 VDD LD.t31 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A VDD.t1831 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X683 VDD 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A a_2749_4932# VDD.t672 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X684 a_22991_5815# Q1.t10 VDD.t2069 VDD.t2060 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X685 a_16065_6276# 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A a_15865_6276# VSS.t171 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X686 DFF_magic_0.tg_magic_2.IN DFF_magic_0.tg_magic_3.CLK.t10 DFF_magic_0.tg_magic_2.OUT VSS.t1500 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X687 a_7303_8697# 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B a_7215_10149# VDD.t1440 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X688 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_3.t7 VDD.t2472 VDD.t2471 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X689 a_23207_5815# Q2.t10 a_22991_5815# VDD.t2414 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X690 VDD a_11279_6341# 7b_counter_0.MDFF_5.tspc2_magic_0.D VDD.t549 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X691 VDD 7b_counter_0.MDFF_7.tspc2_magic_0.D a_24259_4877# VDD.t2318 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X692 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t10 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT VSS.t1389 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X693 VDD CLK.t34 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t4 VDD.t2566 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X694 VDD Q5.t12 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT VDD.t231 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X695 VSS D2_3.t8 a_5470_n6471# VSS.t1456 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X696 VSS 7b_counter_0.MDFF_5.LD.t26 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A VSS.t750 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X697 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t14 VSS.t1301 VSS.t1300 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X698 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A LD.t32 VSS.t1065 VSS.t1064 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X699 VSS a_23258_552# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A VSS.t518 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X700 a_13553_n2115# p2_gen_magic_0.3_inp_AND_magic_0.A a_13353_n2115# VSS.t400 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X701 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A a_1209_9773# VDD.t684 VDD.t683 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X702 a_8523_n4081# p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT VDD.t820 VDD.t240 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X703 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t10 VDD.t1715 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X704 VDD 7b_counter_0.MDFF_4.LD.t52 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A VDD.t1542 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X705 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK CLK.t35 VSS.t628 VSS.t627 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X706 a_17405_3524# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B a_17405_4932# VDD.t951 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X707 VDD 7b_counter_0.MDFF_4.LD.t53 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A VDD.t1545 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X708 VDD a_11279_3480# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t2 VDD.t1144 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X709 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t27 VDD.t1211 VDD.t1210 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X710 p2_gen_magic_0.xnor_magic_4.OUT Q2.t11 a_5054_n1973# VSS.t1409 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X711 a_30365_4922# OR_magic_2.A.t10 VDD.t2337 VDD.t2329 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X712 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t54 VDD.t1548 VDD.t1500 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X713 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A a_15865_9774# VDD.t506 VDD.t505 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X714 VDD a_15865_3363# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B VDD.t1171 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X715 a_19841_9774# 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A VDD.t258 VDD.t257 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X716 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B a_27234_1746# VDD.t465 VDD.t464 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X717 a_5515_3947# a_4496_4393# VSS.t466 VSS.t465 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X718 a_11292_n6613# p3_gen_magic_0.xnor_magic_4.OUT VDD.t491 VDD.t489 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X719 VDD CLK.t36 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD.t2563 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X720 VDD 7b_counter_0.MDFF_4.LD.t55 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A VDD.t1502 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X721 VSS 7b_counter_0.MDFF_6.QB.t6 a_16065_6276# VSS.t1304 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X722 VDD 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A a_26038_684# VDD.t1096 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X723 VSS 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_19307_6886# VSS.t1013 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X724 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT D2_5.t7 VDD.t2727 VDD.t2726 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X725 a_4496_4877# 7b_counter_0.MDFF_0.tspc2_magic_0.D VDD.t875 VDD.t871 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X726 7b_counter_0.DFF_magic_0.tg_magic_2.IN 7b_counter_0.DFF_magic_0.Q.t11 VDD.t2105 VDD.t2104 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X727 VDD CLK.t37 DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD.t2560 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X728 Q1 a_21381_8741# VDD.t548 VDD.t546 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X729 VDD 7b_counter_0.3_inp_AND_magic_0.VOUT 7b_counter_0.DFF_magic_0.D VDD.t789 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X730 VDD 7b_counter_0.MDFF_4.LD.t56 a_23258_1746# VDD.t1551 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X731 VDD divide_by_2_0.tg_magic_1.IN.t14 divide_by_2_0.tg_magic_0.IN VDD.t1407 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X732 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT DFF_magic_0.tg_magic_2.OUT VDD.t2201 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X733 a_19152_5956# 7b_counter_0.MDFF_6.tspc2_magic_0.D VDD.t208 VDD.t207 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X734 a_11279_1124# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A VSS.t178 VSS.t177 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X735 a_8955_8580# 7b_counter_0.MDFF_5.LD.t28 a_8411_8536# VSS.t769 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X736 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t29 VSS.t771 VSS.t770 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X737 VDD LD.t33 a_1209_8579# VDD.t1870 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X738 VSS 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t6 a_24536_3947# VSS.t889 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X739 a_1409_3363# LD.t34 a_1209_3363# VSS.t1066 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X740 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A a_15865_1059# VSS.t308 VSS.t307 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X741 VDD 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A a_7215_4932# VDD.t969 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X742 a_21381_10149# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B a_21381_8741# VDD.t546 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X743 p2_gen_magic_0.3_inp_AND_magic_0.C a_16186_n3644# VSS.t121 VSS.t120 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X744 a_23560_3728# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t7 VDD.t1473 VDD.t1472 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X745 VSS 7b_counter_0.MDFF_5.LD.t30 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A VSS.t753 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X746 VSS DFF_magic_0.D.t17 a_31440_8496.t1 VSS.t1228 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X747 VDD DFF_magic_0.D.t18 a_31440_8496.t7 VDD.t2122 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X748 a_8411_4513# 7b_counter_0.MDFF_4.tspc2_magic_0.Q VDD.t315 VDD.t314 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X749 a_34156_n889# mux_magic_0.OR_magic_0.A VDD.t826 VDD.t821 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X750 a_19841_8580# 7b_counter_0.MDFF_5.LD.t31 VDD.t1213 VDD.t1212 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X751 VSS D2_4.t10 a_1975_n6471# VSS.t1316 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X752 VDD DFF_magic_0.tg_magic_1.IN.t13 DFF_magic_0.tg_magic_0.IN VDD.t56 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X753 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q3.t15 VSS.t1335 VSS.t1334 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X754 p3_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT a_1541_n8579# VDD.t369 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X755 VDD 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t8 a_4496_9609# VDD.t1450 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X756 VSS 7b_counter_0.MDFF_3.tspc2_magic_0.D a_4235_9163# VSS.t882 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X757 a_15865_8580# 7b_counter_0.MDFF_5.LD.t32 VDD.t1215 VDD.t1214 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X758 VDD 7b_counter_0.3_inp_AND_magic_0.A a_23985_7877# VDD.t267 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X759 a_7303_8697# 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A VSS.t271 VSS.t270 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X760 a_8955_9774# 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A a_8411_9730# VSS.t187 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X761 VDD CLK.t38 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t3 VDD.t2557 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X762 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t57 VDD.t1555 VDD.t1554 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X763 a_9212_739# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t7 a_9412_739# VDD.t2710 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X764 7b_counter_0.3_inp_AND_magic_0.C Q3.t16 a_23207_5815# VDD.t2290 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X765 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_3.CLK.t10 divide_by_2_1.tg_magic_3.IN.t9 VSS.t1158 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X766 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t58 VDD.t1557 VDD.t1556 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X767 VDD 7b_counter_0.MDFF_4.LD.t59 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A VDD.t1558 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X768 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.CLK.t11 VDD.t1819 VDD.t1818 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X769 VDD 7b_counter_0.MDFF_4.LD.t60 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A VDD.t1561 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X770 VDD a_26126_3480# 7b_counter_0.MDFF_7.tspc2_magic_0.D VDD.t775 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X771 a_1409_4557# 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A a_1209_4557# VSS.t86 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X772 VDD LD.t35 a_5185_7469# VDD.t1873 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X773 a_1209_6275# 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A VDD.t1704 VDD.t1703 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X774 VDD a_15865_6276# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A VDD.t2203 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X775 VDD 7b_counter_0.MDFF_4.LD.t61 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A VDD.t1564 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X776 VDD Q1.t11 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT VDD.t2070 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X777 VDD LD.t36 a_1209_3363# VDD.t1876 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X778 a_16065_3363# CLK.t39 VSS.t626 VSS.t625 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X779 VDD p3_gen_magic_0.xnor_magic_6.OUT a_14556_n8142# VDD.t936 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X780 VSS D2_2.t12 a_8955_8580# VSS.t1112 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X781 VSS D2_6.t7 a_8939_n7648# VSS.t841 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X782 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5054_n5540# VDD.t401 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X783 a_11191_4932# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A VDD.t523 VDD.t520 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X784 7b_counter_0.DFF_magic_0.tg_magic_3.CLK CLK.t40 VSS.t624 VSS.t623 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X785 VDD CLK.t41 DFF_magic_0.tg_magic_3.CLK.t5 VDD.t2569 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X786 a_22150_1124# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A VSS.t446 VSS.t445 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X787 a_1409_2253# CLK.t42 VSS.t622 VSS.t621 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X788 VDD 7b_counter_0.MDFF_5.tspc2_magic_0.D a_9412_5956# VDD.t889 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X789 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN P2.t9 VDD.t2223 VDD.t2222 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X790 VSS DFF_magic_0.tg_magic_3.CLK.t11 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VSS.t1501 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X791 7b_counter_0.DFF_magic_0.tg_magic_0.IN 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t12 VDD.t915 VDD.t914 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X792 a_5036_n8095# Q6.t13 VDD.t2178 VDD.t1726 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X793 VDD 7b_counter_0.MDFF_4.tspc2_magic_0.Q a_8411_4513# VDD.t311 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X794 VDD CLK.t43 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t5 VDD.t2579 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X795 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT D2_5.t8 VDD.t2729 VDD.t2728 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X796 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A LD.t37 VDD.t1880 VDD.t1879 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X797 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_0.IN VDD.t794 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X798 a_17405_2092# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B VSS.t1282 VSS.t500 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X799 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t33 VSS.t775 VSS.t774 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X800 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT divide_by_2_0.tg_magic_1.IN.t11 VDD.t896 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X801 VDD 7b_counter_0.MDFF_5.LD.t34 a_15865_8580# VDD.t1216 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X802 a_12931_8580# CLK.t44 VSS.t620 VSS.t619 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X803 divide_by_2_0.tg_magic_2.IN divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.IN.t17 VDD.t999 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X804 VDD a_19152_1223# 7b_counter_0.MDFF_1.QB.t1 VDD.t94 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X805 a_16065_4557# Q2.t12 VSS.t1411 VSS.t1410 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X806 VSS D2_7.t8 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT VSS.t1129 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X807 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A LD.t38 VDD.t1882 VDD.t1881 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X808 VDD a_14556_n3644# p2_gen_magic_0.3_inp_AND_magic_0.B VDD.t680 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X809 VDD LD.t39 a_5185_2253# VDD.t1883 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X810 VSS 7b_counter_0.MDFF_5.tspc2_magic_0.Q a_8955_9774# VSS.t354 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X811 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A LD.t40 VDD.t1886 VDD.t1847 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X812 OR_magic_2.VOUT a_23352_n6798# VSS.t112 VSS.t111 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X813 VDD D2_1.t14 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT VDD.t1319 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X814 VDD CLK.t45 a_15865_3363# VDD.t2576 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X815 a_11191_684# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_11279_1124# VDD.t450 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X816 VSS Q4.t9 a_1409_1059# VSS.t978 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X817 VSS p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t4 VSS.t1036 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X818 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.t7 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.t6 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.t7 VDD.t865 pfet_03v3 ad=0.493p pd=3.12u as=0 ps=0 w=1.12u l=0.56u
X819 a_12387_4513# 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A VDD.t1436 VDD.t1435 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X820 a_11191_5901# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_11279_6341# VDD.t551 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X821 a_11279_6341# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A VSS.t179 VSS.t152 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X822 a_17405_10149# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A VDD.t1035 VDD.t1033 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X823 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_3.t9 VDD.t2474 VDD.t2473 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X824 VDD 7b_counter_0.MDFF_7.QB.t5 a_27234_4513# VDD.t0 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X825 VDD p2_gen_magic_0.xnor_magic_0.OUT a_11292_n2115# VDD.t1736 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X826 a_17405_684# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A VDD.t198 VDD.t197 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X827 DFF_magic_0.tg_magic_0.IN DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT DFF_magic_0.tg_magic_3.OUT VDD.t761 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X828 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_6.t8 VDD.t1375 VDD.t1374 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X829 VDD D2_4.t11 a_23258_1746# VDD.t2267 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X830 a_24259_4877# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t8 a_24059_4877# VDD.t1474 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X831 a_12931_9774# Q1.t12 VSS.t1197 VSS.t1196 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X832 a_1209_9773# 7b_counter_0.MDFF_3.QB VDD.t625 VDD.t624 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X833 a_1559_n1042# p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT VDD.t607 VDD.t606 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X834 OR_magic_2.VOUT a_23352_n6798# VDD.t192 VDD.t190 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X835 VDD Q7.t8 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT VDD.t1380 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X836 a_5036_n7648# p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT VSS.t399 VSS.t398 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X837 a_14756_n3644# p2_gen_magic_0.AND2_magic_1.A a_14556_n3644# VSS.t1030 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X838 a_2749_3524# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B a_2749_4932# VDD.t179 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X839 VDD divide_by_2_1.tg_magic_1.IN.t12 divide_by_2_1.tg_magic_0.IN VDD.t477 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X840 a_23207_5815# Q2.t13 a_22991_5815# VDD.t2414 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X841 VDD 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A a_23258_552# VDD.t303 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X842 a_23560_3728# a_24059_4877# a_24536_3947# VSS.t1354 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X843 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1559_n5540# VDD.t408 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X844 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_3.CLK.t12 divide_by_2_0.tg_magic_3.OUT VSS.t1043 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X845 VDD D2_1.t15 p3_gen_magic_0.xnor_magic_1.B VDD.t1322 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X846 a_22991_5815# Q1.t13 VDD.t2073 VDD.t2064 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X847 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_2.t13 VDD.t1938 VDD.t1937 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X848 p3_gen_magic_0.P3 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT VDD.t42 VDD.t41 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X849 a_15865_1059# 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A a_16065_1059# VSS.t306 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X850 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A LD.t41 VSS.t1068 VSS.t1067 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X851 a_17405_4932# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A VDD.t161 VDD.t160 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X852 a_12387_5769# 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A a_12931_6276# VSS.t294 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X853 a_2749_10148# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A VDD.t693 VDD.t692 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X854 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q1.t14 VDD.t2075 VDD.t2074 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X855 VSS a_27567_8496.t11 LD.t2 VSS.t732 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X856 VDD Q4.t10 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT VDD.t1656 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X857 VDD a_27567_8496.t12 LD.t3 VDD.t1178 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X858 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT Q5.t13 VSS.t130 VSS.t129 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X859 VDD 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t6 a_8713_6842# VDD.t886 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X860 VSS p2_gen_magic_0.xnor_magic_3.OUT.t6 a_11708_n2115# VSS.t405 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X861 Q7 a_6725_7308# VDD.t103 VDD.t102 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X862 VSS OR_magic_2.A.t11 DFF_magic_0.tg_magic_2.IN VSS.t1360 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X863 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT CLK.t46 VDD.t2575 VDD.t2574 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X864 VSS OR_magic_2.VOUT.t10 divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT VSS.t383 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X865 a_26038_684# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B a_26126_1124# VDD.t1065 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X866 a_27234_4513# 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A VDD.t1762 VDD.t1761 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X867 a_19307_6886# a_18891_6886# a_19152_6440# VSS.t1021 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X868 a_22062_684# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B a_22150_1124# VDD.t476 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X869 a_4496_4877# 7b_counter_0.MDFF_0.tspc2_magic_0.D VDD.t874 VDD.t873 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X870 VSS OR_magic_2.A.t12 a_23352_n6798# VSS.t1363 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X871 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT divide_by_2_1.tg_magic_0.IN VDD.t1137 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X872 VDD 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A a_7215_10149# VDD.t513 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X873 VDD p3_gen_magic_0.3_inp_AND_magic_0.C.t6 a_13353_n6613# VDD.t1987 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X874 VDD D2_5.t9 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT VDD.t2730 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X875 VSS D2_1.t16 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT VSS.t800 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X876 DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK.t47 VDD.t2573 VDD.t2572 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X877 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_17405_3524# VDD.t722 VDD.t720 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X878 VDD 7b_counter_0.MDFF_6.QB.t7 a_15865_6276# VDD.t2248 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X879 DFF_magic_0.tg_magic_2.OUT DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT DFF_magic_0.tg_magic_1.IN.t9 VDD.t2200 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X880 a_20041_3363# 7b_counter_0.MDFF_4.LD.t62 a_19841_3363# VSS.t923 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X881 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT Q6.t14 VDD.t2180 VDD.t2179 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X882 7b_counter_0.3_inp_AND_magic_0.A Q4.t11 VSS.t982 VSS.t981 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X883 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t35 VDD.t1220 VDD.t1219 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X884 VDD 7b_counter_0.MDFF_6.tspc2_magic_0.D a_19152_5956# VDD.t204 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X885 a_16065_3363# 7b_counter_0.MDFF_4.LD.t63 a_15865_3363# VSS.t910 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X886 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_4.t12 VDD.t2271 VDD.t2270 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X887 a_17405_7309# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B VSS.t325 VSS.t324 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X888 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A LD.t42 VDD.t1888 VDD.t1887 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X889 VDD p3_gen_magic_0.xnor_magic_1.OUT.t6 a_16186_n8142# VDD.t49 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X890 DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT DFF_magic_0.tg_magic_3.CLK.t12 VDD.t2700 VDD.t2699 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X891 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_3.OUT VSS.t81 VSS.t80 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X892 VDD p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT a_1541_n8579# VDD.t844 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X893 VSS 7b_counter_0.MDFF_4.QB.t9 7b_counter_0.MDFF_4.tspc2_magic_0.Q VSS.t1170 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X894 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t1 VDD.t664 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X895 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t11 VDD.t2387 VDD.t2386 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X896 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_17405_8741# VSS.t301 VSS.t300 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X897 7b_counter_0.DFF_magic_0.tg_magic_0.IN 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t13 VDD.t917 VDD.t916 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X898 VDD divide_by_2_1.tg_magic_3.CLK.t11 divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT VDD.t1993 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X899 a_7215_4932# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B a_7303_3480# VDD.t816 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X900 a_23352_n5390# OR_magic_2.A.t13 VDD.t2339 VDD.t2338 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X901 a_32816_n1264# mux_magic_0.AND2_magic_0.A a_32616_n1264# VSS.t522 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X902 VDD a_8411_4513# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A VDD.t966 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X903 a_1541_n7648# p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT VSS.t183 VSS.t182 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X904 VDD a_7303_8697# Q2.t2 VDD.t1445 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X905 7b_counter_0.3_inp_AND_magic_0.A Q5.t14 a_23793_5904# VDD.t221 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X906 VDD Q4.t12 a_12174_n8095# VDD.t633 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X907 a_20041_4557# 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A a_19841_4557# VSS.t1005 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X908 VSS 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B a_7303_8697# VSS.t876 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X909 a_16065_4557# 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A a_15865_4557# VSS.t159 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X910 mux_magic_0.AND2_magic_0.A D2_1.t17 VSS.t804 VSS.t803 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X911 VDD 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A a_11191_10149# VDD.t164 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X912 7b_counter_0.DFF_magic_0.tg_magic_0.IN CLK.t48 7b_counter_0.DFF_magic_0.tg_magic_3.OUT VSS.t618 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X913 mux_magic_0.OR_magic_0.B a_32616_n2458# VDD.t699 VDD.t698 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X914 a_2749_5900# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B a_2749_7308# VDD.t949 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X915 VSS Q1.t15 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT VSS.t1198 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X916 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.B.t6 VSS.t1444 VSS.t1443 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X917 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A a_23258_552# VDD.t986 VDD.t985 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X918 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT D2_5.t10 VSS.t1540 VSS.t1539 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X919 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t64 VDD.t1568 VDD.t1567 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X920 VDD a_27234_552# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A VDD.t541 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X921 VSS CLK.t49 a_16065_3363# VSS.t615 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X922 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t65 VDD.t1570 VDD.t1569 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X923 a_1209_7469# LD.t43 VDD.t1890 VDD.t1889 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X924 a_32816_n2458# D2_1.t18 a_32616_n2458# VSS.t805 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X925 VDD Q4.t13 a_23793_5904# VDD.t1661 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X926 a_11492_n6613# p3_gen_magic_0.xnor_magic_0.OUT a_11292_n6613# VSS.t675 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X927 a_8643_n1042# p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT VDD.t1735 VDD.t1734 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X928 VDD 7b_counter_0.MDFF_5.LD.t36 a_12387_8536# VDD.t1221 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X929 a_21504_5904# Q7.t9 7b_counter_0.3_inp_AND_magic_0.B VDD.t1383 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X930 a_24185_7877# 7b_counter_0.3_inp_AND_magic_0.A a_23985_7877# VSS.t146 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X931 VDD.t1060 VDD.t1059 VDD.t1060 VDD.t905 pfet_03v3 ad=0.493p pd=3.12u as=0 ps=0 w=1.12u l=0.56u
X932 VDD 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t14 7b_counter_0.DFF_magic_0.tg_magic_0.IN VDD.t918 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X933 VDD 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A a_11191_684# VDD.t347 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X934 7b_counter_0.DFF_magic_0.tg_magic_0.IN 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.OUT VDD.t793 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X935 VSS divide_by_2_0.tg_magic_3.CLK.t13 divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT VSS.t1044 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X936 VSS D2_5.t11 a_12590_n7648# VSS.t1541 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X937 VDD Q2.t14 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT VDD.t2419 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X938 VSS CLK.t50 a_12931_8580# VSS.t612 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X939 a_11492_n6613# p3_gen_magic_0.xnor_magic_0.OUT a_11292_n6613# VSS.t675 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X940 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A LD.t44 VDD.t1892 VDD.t1891 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X941 a_8523_n8095# D2_6.t9 p3_gen_magic_0.xnor_magic_6.OUT VDD.t64 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X942 divide_by_2_1.tg_magic_0.IN divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.OUT VDD.t1136 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X943 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A LD.t45 VSS.t1070 VSS.t1069 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X944 VSS Q2.t15 a_16065_4557# VSS.t1412 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X945 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A LD.t46 VSS.t1072 VSS.t1071 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X946 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK.t51 VDD.t2591 VDD.t2590 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X947 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t12 VDD.t2033 VDD.t2032 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X948 a_2749_10148# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B a_2749_8740# VDD.t68 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X949 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t37 VSS.t777 VSS.t776 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X950 divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT OR_magic_2.VOUT.t11 VDD.t737 VDD.t736 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X951 p2_gen_magic_0.3_inp_AND_magic_0.C a_16186_n3644# VDD.t219 VDD.t218 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X952 VSS a_12387_6963# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B VSS.t295 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X953 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT CLK.t52 VDD.t2589 VDD.t2588 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X954 a_11492_n2115# p2_gen_magic_0.xnor_magic_4.OUT a_11708_n2115# VSS.t405 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X955 a_1209_2253# LD.t47 VDD.t1894 VDD.t1893 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X956 VSS DFF_magic_0.tg_magic_1.IN.t14 DFF_magic_0.tg_magic_0.IN VSS.t40 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X957 VDD 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A a_26038_4932# VDD.t390 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X958 VDD Q5.t15 a_12387_4513# VDD.t234 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X959 a_34156_n2297# mux_magic_0.OR_magic_0.B VSS.t34 VSS.t33 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X960 7b_counter_0.MDFF_0.tspc2_magic_0.D a_2749_3524# VSS.t108 VSS.t107 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X961 a_27234_4513# 7b_counter_0.MDFF_7.QB.t6 VDD.t4 VDD.t3 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X962 p3_gen_magic_0.3_inp_AND_magic_0.A a_11292_n6613# VDD.t1078 VDD.t1076 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X963 DFF_magic_0.tg_magic_2.IN OR_magic_2.A.t14 VDD.t2341 VDD.t2340 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X964 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.D VDD.t366 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X965 VDD D2_1.t19 a_32616_n2458# VDD.t1325 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X966 a_5452_n3150# p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_5.OUT VSS.t144 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X967 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_4.t13 VSS.t1320 VSS.t1319 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X968 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_15865_7470# VDD.t1131 VDD.t1130 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X969 a_13353_n6613# p3_gen_magic_0.3_inp_AND_magic_0.B VDD.t1797 VDD.t1795 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X970 VDD 7b_counter_0.MDFF_7.QB.t7 7b_counter_0.MDFF_7.tspc2_magic_0.Q VDD.t5 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X971 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A a_5185_6275# VSS.t110 VSS.t109 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X972 a_23793_5904# Q4.t14 VDD.t1665 VDD.t1664 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X973 VSS Q1.t16 a_12931_9774# VSS.t1201 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X974 p3_gen_magic_0.3_inp_AND_magic_0.B a_14556_n8142# VSS.t1033 VSS.t1032 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X975 mux_magic_0.OR_magic_0.A a_32616_n1264# VSS.t498 VSS.t497 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X976 VSS p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t15 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN VSS.t1297 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X977 VSS divide_by_2_1.tg_magic_3.IN.t20 mux_magic_0.IN1.t1 VSS.t73 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X978 VSS Q7.t10 7b_counter_0.3_inp_AND_magic_0.B VSS.t851 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X979 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A LD.t48 VDD.t1895 VDD.t1887 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X980 VDD Q4.t15 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT VDD.t1666 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X981 VDD CLK.t53 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD.t2585 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X982 a_12931_2253# D2_6.t10 VSS.t844 VSS.t568 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X983 Q5 a_6725_2092# VSS.t536 VSS.t535 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X984 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK VDD.t1161 VDD.t1160 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X985 a_24536_3947# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t9 VSS.t893 VSS.t892 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X986 a_34156_n2297# mux_magic_0.OR_magic_0.B a_34156_n889# VDD.t46 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X987 DFF_magic_0.tg_magic_2.OUT DFF_magic_0.tg_magic_3.CLK.t13 DFF_magic_0.tg_magic_2.IN VSS.t1504 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X988 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B a_19841_3363# VDD.t432 VDD.t431 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X989 VDD 7b_counter_0.MDFF_5.tspc2_magic_0.Q a_8411_9730# VDD.t702 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X990 VSS CLK.t54 a_27778_2253# VSS.t609 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X991 a_15865_2253# D2_3.t10 VDD.t2476 VDD.t2475 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X992 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_17405_8741# VDD.t576 VDD.t575 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X993 VSS DFF_magic_0.D.t21 a_27567_8496.t1 VSS.t1233 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X994 VDD DFF_magic_0.D.t22 a_27567_8496.t7 VDD.t2127 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X995 LD a_27567_8496.t13 VSS.t736 VSS.t735 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X996 p2_gen_magic_0.xnor_magic_4.OUT D2_3.t11 a_5054_n1526# VDD.t770 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X997 LD a_27567_8496.t14 VDD.t1182 VDD.t1181 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X998 a_19841_8580# D2_1.t20 VDD.t1329 VDD.t1328 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X999 a_8713_6842# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t7 VDD.t911 VDD.t884 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1000 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B a_5185_7469# VSS.t1000 VSS.t999 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1001 VSS D2_2.t14 a_9059_n1973# VSS.t1115 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1002 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_7.t9 VDD.t1970 VDD.t1969 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1003 mux_magic_0.OR_magic_0.B a_32616_n2458# VSS.t353 VSS.t352 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1004 VDD 7b_counter_0.MDFF_7.tspc2_magic_0.D a_24259_4877# VDD.t1467 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1005 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT CLK.t55 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN VSS.t608 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1006 VDD Q5.t16 a_8523_n8095# VDD.t237 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1007 a_19307_1669# 7b_counter_0.MDFF_1.tspc2_magic_0.CLK VSS.t508 VSS.t507 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1008 a_5036_n4081# p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT VDD.t266 VDD.t265 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1009 a_7215_10149# 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B a_7303_8697# VDD.t510 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1010 VDD divide_by_2_1.tg_magic_3.IN.t21 mux_magic_0.IN1.t3 VDD.t114 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1011 p2_gen_magic_0.xnor_magic_5.OUT D2_7.t10 a_5036_n3597# VDD.t399 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1012 divide_by_2_1.tg_magic_0.IN divide_by_2_1.tg_magic_1.IN.t13 VDD.t481 VDD.t480 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1013 a_23352_n5390# OR_magic_2.A.t15 VDD.t2342 VDD.t1456 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1014 VDD CLK.t56 DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD.t2582 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1015 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_6.t11 VSS.t830 VSS.t829 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1016 VSS D2_1.t21 p3_gen_magic_0.xnor_magic_1.B VSS.t806 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1017 divide_by_2_1.tg_magic_2.IN mux_magic_0.IN1.t10 VDD.t2360 VDD.t2359 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1018 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B a_19841_8580# VSS.t696 VSS.t695 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1019 VDD divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_1.IN.t3 VDD.t126 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1020 VSS Q4.t16 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT VSS.t983 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1021 p2_gen_magic_0.xnor_magic_3.OUT Q3.t17 a_1559_n1973# VSS.t1333 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1022 a_24185_7877# 7b_counter_0.3_inp_AND_magic_0.A a_23985_7877# VSS.t146 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1023 a_27778_2253# CLK.t57 VSS.t607 VSS.t606 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1024 VDD a_19841_4557# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A VDD.t655 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1025 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK.t58 VDD.t2600 VDD.t2599 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1026 VDD a_11279_8697# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t2 VDD.t165 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1027 7b_counter_0.DFF_magic_0.tg_magic_1.IN CLK.t59 7b_counter_0.DFF_magic_0.tg_magic_2.OUT VSS.t605 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1028 OR_magic_2.A DFF_magic_0.tg_magic_2.OUT VDD.t1007 VDD.t1006 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1029 a_21381_3524# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B a_21381_4932# VDD.t80 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1030 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A a_8411_9730# VDD.t379 VDD.t378 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1031 VDD a_11279_1124# 7b_counter_0.MDFF_4.tspc2_magic_0.D VDD.t1772 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1032 VSS OR_magic_1.VOUT.t14 divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT VSS.t1475 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1033 VDD 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A a_12387_552# VDD.t2379 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1034 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A a_19841_9774# VSS.t101 VSS.t100 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1035 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t12 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN VSS.t1390 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1036 a_12387_3319# 7b_counter_0.MDFF_4.LD.t66 a_12931_3363# VSS.t918 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1037 a_11191_4932# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B a_11279_3480# VDD.t517 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1038 a_2749_7308# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B a_2749_5900# VDD.t1040 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1039 VDD p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD.t1157 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1040 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B a_8411_3319# VDD.t338 VDD.t337 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1041 7b_counter_0.DFF_magic_0.Q 7b_counter_0.DFF_magic_0.tg_magic_2.OUT VDD.t614 VDD.t613 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1042 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT VSS.t720 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1043 VDD a_12387_4513# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A VDD.t1140 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1044 p2_gen_magic_0.xnor_magic_3.OUT D2_4.t14 a_1559_n1526# VDD.t2046 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1045 VDD LD.t49 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A VDD.t1865 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1046 p3_gen_magic_0.3_inp_AND_magic_0.B a_14556_n8142# VDD.t1791 VDD.t1790 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1047 7b_counter_0.DFF_magic_0.tg_magic_2.IN 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t13 7b_counter_0.DFF_magic_0.tg_magic_2.OUT VSS.t1174 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1048 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.B.t7 VDD.t2461 VDD.t2460 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1049 VSS 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B a_11279_8697# VSS.t97 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1050 7b_counter_0.MDFF_0.tspc2_magic_0.D a_2749_3524# VDD.t184 VDD.t181 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1051 VDD 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_19841_9774# VDD.t274 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1052 a_5185_6275# 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A a_5385_6275# VSS.t328 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1053 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t38 VDD.t1225 VDD.t1224 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1054 VDD p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t7 VDD.t1089 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1055 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK VDD.t1156 VDD.t1155 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1056 VSS Q5.t17 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT VSS.t131 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1057 p2_gen_magic_0.AND2_magic_1.A Q4.t17 a_12174_n3150# VSS.t986 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1058 7b_counter_0.3_inp_AND_magic_0.C Q3.t18 a_23207_5815# VDD.t2284 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1059 7b_counter_0.3_inp_AND_magic_0.B Q7.t11 a_21504_5904# VDD.t1384 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1060 a_15865_9774# 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A VDD.t498 VDD.t497 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1061 7b_counter_0.MDFF_6.tspc2_magic_0.Q 7b_counter_0.MDFF_6.QB.t8 VSS.t1308 VSS.t1307 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1062 a_12387_4513# 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A a_12931_4557# VSS.t875 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1063 a_21504_5904# Q6.t15 VDD.t2181 VDD.t2176 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1064 divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT OR_magic_2.VOUT.t12 VDD.t739 VDD.t738 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1065 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q1.t17 VDD.t2077 VDD.t2076 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1066 a_21381_4932# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B a_21381_3524# VDD.t79 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1067 a_15865_2253# 7b_counter_0.MDFF_4.LD.t67 VDD.t1572 VDD.t1571 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1068 a_12931_6276# 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A a_12387_5769# VSS.t293 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1069 a_5054_n1042# p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT VDD.t297 VDD.t296 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1070 VDD 7b_counter_0.MDFF_5.LD.t39 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A VDD.t1226 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1071 VDD D2_3.t12 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT VDD.t2477 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1072 OR_magic_1.VOUT a_30365_3514# VDD.t979 VDD.t977 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1073 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN p3_gen_magic_0.P3.t10 VDD.t1464 VDD.t1463 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1074 a_5185_7469# LD.t50 a_5385_7469# VSS.t1073 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1075 a_6725_5900# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A VDD.t540 VDD.t537 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1076 a_1559_n6024# Q3.t19 VDD.t2302 VDD.t578 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1077 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A LD.t51 VSS.t1074 VSS.t1071 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1078 a_26038_4932# 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_26126_3480# VDD.t774 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1079 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN CLK.t60 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT VSS.t604 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1080 a_19152_6440# 7b_counter_0.MDFF_6.tspc2_magic_0.CLK VDD.t1752 VDD.t202 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1081 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t40 VDD.t1230 VDD.t1229 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1082 VDD D2_5.t12 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT VDD.t2733 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1083 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK VDD.t1154 VDD.t1153 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1084 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p2_gen_magic_0.3_inp_AND_magic_0.VOUT.t5 VDD.t318 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1085 VDD 7b_counter_0.MDFF_4.LD.t68 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A VDD.t1519 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1086 7b_counter_0.DFF_magic_0.D 7b_counter_0.DFF_magic_0.Q.t12 a_24003_10051# VSS.t1215 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1087 divide_by_2_0.tg_magic_0.IN divide_by_2_0.tg_magic_1.IN.t15 VDD.t1411 VDD.t1410 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1088 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT divide_by_2_0.tg_magic_2.IN VDD.t998 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1089 VDD p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT a_12174_n4081# VDD.t666 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1090 VSS p2_gen_magic_0.xnor_magic_1.OUT.t6 a_16386_n3644# VSS.t1401 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1091 VDD a_26126_1124# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t2 VDD.t1064 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1092 VDD a_22150_1124# Q4.t2 VDD.t475 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1093 a_1541_n8095# Q7.t12 VDD.t1385 VDD.t842 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1094 VDD 7b_counter_0.MDFF_4.LD.t69 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A VDD.t1575 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1095 a_20041_3363# D2_3.t13 VSS.t1460 VSS.t1459 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1096 VDD 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A a_17405_5901# VDD.t2211 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1097 a_8523_n3150# p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT VSS.t450 VSS.t449 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1098 a_27234_3319# 7b_counter_0.MDFF_4.LD.t70 a_27778_3363# VSS.t919 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1099 a_12174_n3597# Q4.t18 VDD.t1669 VDD.t669 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1100 DFF_magic_0.D DFF_magic_0.tg_magic_3.CLK.t14 DFF_magic_0.tg_magic_3.OUT VSS.t1505 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1101 VDD a_27234_3319# 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B VDD.t1081 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1102 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A a_12387_552# VDD.t647 VDD.t646 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1103 VDD 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A a_8411_9730# VDD.t375 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1104 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A a_1209_4557# VDD.t706 VDD.t705 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1105 VSS D2_6.t12 a_12931_2253# VSS.t548 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1106 VSS a_23560_3728# a_23672_3947# VSS.t1493 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1107 a_23985_7877# 7b_counter_0.3_inp_AND_magic_0.B VDD.t1756 VDD.t1755 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1108 a_12387_6963# 7b_counter_0.MDFF_5.LD.t41 VDD.t1232 VDD.t1231 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1109 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_7.t11 VDD.t1972 VDD.t1971 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1110 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A LD.t52 VDD.t1898 VDD.t1891 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1111 VDD D2_3.t14 a_19841_3363# VDD.t2480 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1112 DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT DFF_magic_0.tg_magic_0.IN VDD.t760 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1113 VDD p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT P2.t4 VDD.t2371 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1114 a_27778_2253# 7b_counter_0.MDFF_4.LD.t71 a_27234_1746# VSS.t924 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1115 VDD 7b_counter_0.MDFF_4.LD.t72 a_15865_2253# VDD.t1578 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1116 VSS a_4496_9609# a_5515_9163# VSS.t210 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1117 VDD p2_gen_magic_0.3_inp_AND_magic_0.C.t4 a_13353_n2115# VDD.t2714 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1118 a_23802_2253# 7b_counter_0.MDFF_4.LD.t73 a_23258_1746# VSS.t925 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1119 VSS 7b_counter_0.MDFF_5.LD.t42 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A VSS.t778 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1120 VDD 7b_counter_0.MDFF_5.LD.t43 a_19841_8580# VDD.t1233 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1121 divide_by_2_1.tg_magic_2.IN divide_by_2_1.tg_magic_3.CLK.t12 divide_by_2_1.tg_magic_3.IN.t13 VSS.t1159 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1122 a_6725_7308# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B a_6725_5900# VDD.t533 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1123 a_2749_7308# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B a_2749_5900# VDD.t423 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1124 a_20041_4557# 7b_counter_0.MDFF_1.tspc2_magic_0.Q VSS.t337 VSS.t336 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1125 a_27234_4513# 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A a_27778_4557# VSS.t1025 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1126 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B a_5185_2253# VSS.t974 VSS.t973 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1127 VDD 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A a_2749_5900# VDD.t427 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1128 a_22991_5815# Q1.t18 VDD.t2078 VDD.t2060 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1129 mux_magic_0.IN1 divide_by_2_1.tg_magic_3.IN.t22 VDD.t118 VDD.t117 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1130 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_6.t13 VDD.t1358 VDD.t1357 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1131 a_8523_n4081# p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_6.OUT VDD.t862 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1132 a_11708_n2115# p2_gen_magic_0.xnor_magic_4.OUT a_11492_n2115# VSS.t404 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1133 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t74 VDD.t1582 VDD.t1581 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1134 DFF_magic_0.tg_magic_2.IN OR_magic_2.A.t16 VSS.t1367 VSS.t1366 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1135 a_4496_10093# 7b_counter_0.MDFF_3.tspc2_magic_0.D VDD.t1454 VDD.t1453 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1136 VSS divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_1.IN.t4 VSS.t436 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1137 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A LD.t53 VDD.t1899 VDD.t1879 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1138 a_11191_10149# 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B a_11279_8697# VDD.t164 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1139 a_12387_8536# CLK.t61 VDD.t2598 VDD.t2597 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1140 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_7.t12 VSS.t1133 VSS.t1132 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1141 VDD p2_gen_magic_0.AND2_magic_1.A a_14556_n3644# VDD.t1787 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1142 p2_gen_magic_0.xnor_magic_6.OUT Q5.t18 a_8523_n3150# VSS.t134 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1143 a_30365_3514# P2.t10 a_30365_4922# VDD.t2219 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1144 p2_gen_magic_0.3_inp_AND_magic_0.A a_11292_n2115# VDD.t365 VDD.t363 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1145 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t75 VDD.t1583 VDD.t1533 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1146 a_9412_739# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t8 a_9212_739# VDD.t2708 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1147 p2_gen_magic_0.3_inp_AND_magic_0.VOUT a_13353_n2115# VDD.t1109 VDD.t1107 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1148 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN p3_gen_magic_0.P3.t11 VSS.t888 VSS.t887 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1149 a_13353_n2115# p2_gen_magic_0.3_inp_AND_magic_0.B VDD.t1112 VDD.t1110 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1150 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t76 VDD.t1585 VDD.t1584 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1151 7b_counter_0.DFF_magic_0.tg_magic_2.OUT CLK.t62 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t7 VSS.t603 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1152 a_34156_n889# mux_magic_0.OR_magic_0.B a_34156_n2297# VDD.t48 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1153 VDD D2_2.t15 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT VDD.t1939 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1154 VDD Q6.t16 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT VDD.t2182 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1155 VSS OR_magic_1.VOUT.t15 divide_by_2_1.tg_magic_3.CLK VSS.t1478 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1156 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t13 VDD.t2389 VDD.t2388 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1157 divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT OR_magic_1.VOUT.t16 VSS.t1482 VSS.t1481 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1158 LD a_27567_8496.t15 VDD.t1183 VDD.t1176 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1159 VDD 7b_counter_0.MDFF_5.LD.t44 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A VDD.t1236 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1160 VDD OR_magic_2.VOUT.t13 divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT VDD.t740 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1161 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK VSS.t719 VSS.t718 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1162 VDD 7b_counter_0.MDFF_5.LD.t45 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A VDD.t1226 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1163 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN VDD.t1798 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1164 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B a_12387_3319# VDD.t1067 VDD.t1066 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1165 a_8643_n6024# Q1.t19 VDD.t2079 VDD.t990 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1166 divide_by_2_0.tg_magic_0.IN divide_by_2_0.tg_magic_1.IN.t16 VSS.t864 VSS.t863 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1167 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q3.t20 VDD.t2296 VDD.t2295 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1168 VDD 7b_counter_0.MDFF_5.LD.t46 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A VDD.t1241 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1169 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t16 VDD.t2237 VDD.t2236 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1170 a_11191_5901# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_11279_6341# VDD.t550 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1171 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t14 7b_counter_0.DFF_magic_0.tg_magic_2.IN VSS.t1175 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1172 VSS 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A a_2749_3524# VSS.t89 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1173 7b_counter_0.MDFF_3.QB a_4496_9609# VDD.t418 VDD.t417 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1174 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t47 VDD.t1244 VDD.t1229 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1175 VSS 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t15 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VSS.t1176 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1176 VSS divide_by_2_1.tg_magic_1.IN.t14 divide_by_2_1.tg_magic_0.IN VSS.t254 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1177 VSS 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 7b_counter_0.DFF_magic_0.Q.t1 VSS.t314 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1178 VDD D2_6.t14 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT VDD.t1346 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1179 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B a_1209_8579# VSS.t169 VSS.t87 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1180 a_5385_6275# 7b_counter_0.MDFF_3.tspc2_magic_0.Q VSS.t292 VSS.t291 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1181 a_19152_739# 7b_counter_0.MDFF_1.tspc2_magic_0.D VDD.t1026 VDD.t1025 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1182 p3_gen_magic_0.xnor_magic_5.OUT Q6.t17 a_5036_n7648# VSS.t1265 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1183 VDD p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT a_8523_n4081# VDD.t249 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1184 a_20171_1669# 7b_counter_0.MDFF_1.tspc2_magic_0.CLK 7b_counter_0.MDFF_1.QB.t3 VSS.t506 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1185 a_11191_10149# 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B a_11279_8697# VDD.t163 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1186 VDD 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A a_12387_9730# VDD.t1104 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1187 VDD mux_magic_0.IN2.t9 divide_by_2_0.tg_magic_2.IN VDD.t2148 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1188 VDD OR_magic_1.VOUT.t17 divide_by_2_1.tg_magic_3.CLK VDD.t2514 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1189 VSS a_19152_6440# a_20171_6886# VSS.t261 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1190 VDD 7b_counter_0.MDFF_5.LD.t48 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A VDD.t1245 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1191 divide_by_2_0.tg_magic_0.IN OR_magic_2.VOUT.t14 divide_by_2_0.tg_magic_3.OUT VSS.t386 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1192 a_8523_n3597# Q5.t19 VDD.t241 VDD.t240 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1193 VSS 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A a_6725_2092# VSS.t996 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1194 VDD CLK.t63 a_15865_9774# VDD.t2594 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1195 7b_counter_0.MDFF_5.LD a_29512_8496.t13 VSS.t740 VSS.t739 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1196 7b_counter_0.MDFF_5.LD a_29512_8496.t14 VDD.t1190 VDD.t1189 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1197 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_3.t15 VSS.t1462 VSS.t1461 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1198 a_5054_n1042# p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_4.OUT VDD.t769 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1199 a_7215_4932# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A VDD.t974 VDD.t969 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1200 a_26126_1124# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B a_26038_684# VDD.t1064 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1201 VSS a_12387_552# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A VSS.t330 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1202 VDD p3_gen_magic_0.xnor_magic_0.OUT a_11292_n6613# VDD.t1071 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1203 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT Q4.t19 VDD.t1671 VDD.t1670 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1204 VDD Q1.t20 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT VDD.t2080 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1205 a_19152_739# 7b_counter_0.MDFF_1.tspc2_magic_0.D VDD.t1024 VDD.t1023 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1206 a_5385_7469# D2_7.t13 VSS.t1135 VSS.t1134 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1207 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK CLK.t64 VDD.t2593 VDD.t2592 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1208 DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK.t65 VDD.t2602 VDD.t2601 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1209 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK.t66 VSS.t602 VSS.t601 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1210 7b_counter_0.DFF_magic_0.D 7b_counter_0.3_inp_AND_magic_0.VOUT VDD.t788 VDD.t787 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1211 VDD 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t2 VDD.t796 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1212 VDD 7b_counter_0.MDFF_5.LD.t49 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A VDD.t1248 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1213 a_5185_2253# LD.t54 a_5385_2253# VSS.t1075 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1214 VDD p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t14 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD.t2390 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1215 divide_by_2_1.tg_magic_0.IN divide_by_2_1.tg_magic_1.IN.t15 VDD.t483 VDD.t482 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1216 VSS a_8713_6842# a_8825_6886# VSS.t367 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1217 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_2749_7308# VDD.t948 VDD.t947 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1218 VSS Q3.t21 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT VSS.t1338 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1219 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A a_12387_5769# VDD.t403 VDD.t402 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1220 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_2.t16 VSS.t1119 VSS.t1118 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1221 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT divide_by_2_1.tg_magic_1.IN.t6 VDD.t436 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1222 VSS D2_3.t16 a_20041_3363# VSS.t1463 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1223 VDD 7b_counter_0.MDFF_4.LD.t77 a_12387_1746# VDD.t1586 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1224 divide_by_2_1.tg_magic_2.IN mux_magic_0.IN1.t11 VSS.t1372 VSS.t1371 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1225 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_27234_3319# VDD.t1080 VDD.t1079 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1226 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN VDD.t1741 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1227 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT Q5.t20 VDD.t243 VDD.t242 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1228 a_11708_n2115# p2_gen_magic_0.xnor_magic_4.OUT a_11492_n2115# VSS.t404 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1229 a_6725_2092# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B VSS.t214 VSS.t213 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1230 VDD D2_2.t17 a_12387_6963# VDD.t1942 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1231 a_2749_2092# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B VSS.t184 VSS.t105 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1232 VDD D2_1.t22 mux_magic_0.AND2_magic_0.A VDD.t1309 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1233 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_4.t15 VDD.t2273 VDD.t2272 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1234 a_13353_n2115# p2_gen_magic_0.3_inp_AND_magic_0.B VDD.t1111 VDD.t1110 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1235 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q2.t16 VDD.t2423 VDD.t2422 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1236 p3_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT a_5036_n8579# VDD.t758 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1237 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B a_15865_8580# VSS.t195 VSS.t194 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1238 VDD divide_by_2_0.tg_magic_3.CLK.t14 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT VDD.t1820 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1239 a_1559_n1042# p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_3.OUT VDD.t2045 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1240 VSS 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_20041_4557# VSS.t333 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1241 VDD 7b_counter_0.MDFF_5.LD.t50 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A VDD.t1251 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1242 a_1957_n3150# p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_1.OUT.t0 VSS.t424 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1243 a_21381_3524# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B a_21381_4932# VDD.t78 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1244 a_12931_3363# 7b_counter_0.MDFF_4.LD.t78 a_12387_3319# VSS.t922 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1245 VDD 7b_counter_0.MDFF_5.LD.t51 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A VDD.t1236 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1246 a_14756_n3644# p2_gen_magic_0.xnor_magic_6.OUT VSS.t456 VSS.t455 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1247 VDD CLK.t67 DFF_magic_0.tg_magic_3.CLK.t4 VDD.t2606 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1248 VSS a_27234_552# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A VSS.t281 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1249 a_16065_7470# D2_1.t23 VSS.t809 VSS.t558 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1250 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t79 VDD.t1590 VDD.t1589 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1251 VDD a_15865_4557# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A VDD.t151 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1252 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT DFF_magic_0.tg_magic_3.CLK.t15 VSS.t1507 VSS.t1506 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1253 7b_counter_0.MDFF_1.tspc2_magic_0.D a_17405_2092# VSS.t1356 VSS.t370 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1254 a_21381_8741# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B VSS.t698 VSS.t697 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1255 VDD 7b_counter_0.MDFF_4.LD.t80 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A VDD.t1575 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1256 a_2749_4932# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A VDD.t673 VDD.t672 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1257 a_1209_8579# LD.t55 a_1409_8579# VSS.t1060 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1258 VDD 7b_counter_0.MDFF_5.tspc2_magic_0.D a_9412_5956# VDD.t889 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1259 a_12174_n8095# D2_5.t13 p3_gen_magic_0.AND2_magic_1.A VDD.t1415 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1260 a_23258_552# 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A a_23802_1059# VSS.t161 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1261 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t81 VDD.t1593 VDD.t1556 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1262 a_11279_3480# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A VSS.t272 VSS.t177 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1263 a_1409_9773# 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A a_1209_9773# VSS.t413 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1264 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A a_15865_9774# VSS.t269 VSS.t268 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1265 a_16186_n3644# p2_gen_magic_0.xnor_magic_5.OUT VDD.t211 VDD.t210 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1266 DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT DFF_magic_0.tg_magic_3.CLK.t16 VSS.t1509 VSS.t1508 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1267 VSS p2_gen_magic_0.3_inp_AND_magic_0.C.t5 a_13769_n2115# VSS.t688 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1268 VDD 7b_counter_0.MDFF_4.LD.t82 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A VDD.t1561 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1269 a_2749_4932# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A VDD.t671 VDD.t178 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1270 VDD 7b_counter_0.MDFF_4.LD.t83 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A VDD.t1564 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1271 a_23207_5815# Q2.t17 a_22991_5815# VDD.t2414 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1272 VDD Q7.t13 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT VDD.t1386 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1273 a_12931_4557# 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A a_12387_4513# VSS.t874 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1274 a_34156_n2297# mux_magic_0.OR_magic_0.B a_34156_n889# VDD.t47 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1275 VDD a_23258_552# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A VDD.t982 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1276 VDD 7b_counter_0.MDFF_4.LD.t84 a_27234_1746# VDD.t1598 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1277 a_1541_n4081# p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT VDD.t807 VDD.t806 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1278 VDD divide_by_2_0.tg_magic_3.IN.t21 mux_magic_0.IN2.t3 VDD.t14 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1279 VDD a_16186_n8142# p3_gen_magic_0.3_inp_AND_magic_0.C.t1 VDD.t1721 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1280 VSS p3_gen_magic_0.xnor_magic_6.OUT a_14756_n8142# VSS.t492 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1281 VDD D2_7.t14 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT VDD.t1973 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1282 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.IN.t0 VDD.t562 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1283 a_19152_739# 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_18891_1669# VDD.t961 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1284 a_11279_6341# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_11191_5901# VDD.t549 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1285 VSS Q2.t18 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT VSS.t1415 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1286 VDD 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A a_1209_9773# VDD.t784 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1287 VSS 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t1 VSS.t421 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1288 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t52 VSS.t781 VSS.t774 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1289 7b_counter_0.DFF_magic_0.tg_magic_2.IN 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t16 7b_counter_0.DFF_magic_0.tg_magic_2.OUT VSS.t1179 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1290 VDD p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t17 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN VDD.t2238 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1291 VDD 7b_counter_0.MDFF_5.LD.t53 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A VDD.t1248 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1292 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q7.t14 VDD.t1390 VDD.t1389 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1293 OR_magic_2.A DFF_magic_0.tg_magic_2.OUT VSS.t525 VSS.t524 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1294 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t17 VSS.t1181 VSS.t1180 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1295 VSS p2_gen_magic_0.3_inp_AND_magic_0.C.t6 a_13769_n2115# VSS.t1523 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1296 a_32816_n1264# mux_magic_0.IN1.t12 VSS.t1374 VSS.t1373 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1297 divide_by_2_1.tg_magic_0.IN divide_by_2_1.tg_magic_1.IN.t16 VSS.t258 VSS.t257 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1298 VSS 7b_counter_0.MDFF_5.LD.t54 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A VSS.t782 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1299 VSS 7b_counter_0.DFF_magic_0.Q.t13 7b_counter_0.DFF_magic_0.tg_magic_2.IN VSS.t1216 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1300 a_17405_4932# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B a_17405_3524# VDD.t720 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1301 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.IN.t17 VDD.t1768 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1302 VDD 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_19152_1223# VDD.t958 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1303 VSS Q6.t18 a_1409_6275# VSS.t1266 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1304 VDD 7b_counter_0.MDFF_5.LD.t55 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A VDD.t1258 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1305 7b_counter_0.MDFF_4.LD a_31440_8496.t14 VSS.t19 VSS.t18 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1306 7b_counter_0.MDFF_4.LD a_31440_8496.t15 VDD.t27 VDD.t20 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1307 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_3.CLK.t15 divide_by_2_0.tg_magic_3.IN.t10 VSS.t1047 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1308 a_8713_1625# a_9212_739# a_9689_1669# VSS.t700 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1309 VDD 7b_counter_0.MDFF_5.LD.t56 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A VDD.t1261 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1310 a_5054_n6024# Q2.t19 VDD.t2424 VDD.t73 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1311 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B a_1209_3363# VSS.t157 VSS.t156 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1312 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t57 VDD.t1264 VDD.t1210 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1313 mux_magic_0.AND2_magic_0.A D2_1.t24 VSS.t811 VSS.t810 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1314 VDD 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A a_1209_4557# VDD.t136 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1315 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t58 VDD.t1265 VDD.t1224 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1316 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_2.t18 VDD.t1946 VDD.t1945 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1317 VSS a_29512_8496.t15 7b_counter_0.MDFF_5.LD.t0 VSS.t741 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1318 VDD a_29512_8496.t16 7b_counter_0.MDFF_5.LD.t4 VDD.t1191 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1319 VDD a_12387_6963# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B VDD.t712 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1320 VDD 7b_counter_0.MDFF_1.QB.t7 a_15865_1059# VDD.t89 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1321 VSS OR_magic_1.VOUT.t18 divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT VSS.t1483 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1322 VDD 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A a_7215_4932# VDD.t816 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1323 a_4235_3947# 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t5 a_4496_4877# VDD.t2449 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1324 VDD CLK.t68 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD.t2603 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1325 a_5515_9163# a_4496_9609# VSS.t209 VSS.t208 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1326 VDD 7b_counter_0.MDFF_5.LD.t59 a_8411_8536# VDD.t1266 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1327 VDD 7b_counter_0.MDFF_5.tspc2_magic_0.D a_9412_5956# VDD.t886 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1328 VDD OR_magic_2.A.t17 DFF_magic_0.tg_magic_2.IN VDD.t2343 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1329 a_5185_6275# 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A VDD.t639 VDD.t638 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1330 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT VSS.t717 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1331 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q7.t15 VDD.t1392 VDD.t1391 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1332 a_17405_3524# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B VSS.t501 VSS.t500 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1333 a_32816_n2458# mux_magic_0.IN2.t10 VSS.t1249 VSS.t1248 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1334 VSS CLK.t69 a_1409_7469# VSS.t598 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1335 7b_counter_0.MDFF_6.tspc2_magic_0.D a_17405_7309# VSS.t326 VSS.t300 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1336 a_8643_n1042# p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_0.OUT VDD.t458 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1337 a_15865_8580# 7b_counter_0.MDFF_5.LD.t60 a_16065_8580# VSS.t758 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1338 a_24003_10051# 7b_counter_0.DFF_magic_0.Q.t14 7b_counter_0.DFF_magic_0.D VSS.t1219 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1339 a_12174_n8579# p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT VDD.t637 VDD.t636 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1340 a_26126_1124# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A VSS.t684 VSS.t192 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1341 a_5385_2253# D2_5.t14 VSS.t1545 VSS.t1544 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1342 a_16386_n3644# p2_gen_magic_0.xnor_magic_1.OUT.t7 VSS.t1405 VSS.t1404 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1343 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A a_1209_4557# VSS.t360 VSS.t359 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1344 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT Q5.t21 VDD.t245 VDD.t244 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1345 VDD a_1209_6275# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A VDD.t1710 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1346 a_8825_6886# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t8 7b_counter_0.MDFF_5.QB.t3 VSS.t475 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1347 VSS 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_5385_1059# VSS.t439 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1348 a_4651_3947# a_4235_3947# a_4496_4393# VSS.t155 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1349 a_16065_7470# 7b_counter_0.MDFF_5.LD.t61 a_15865_7470# VSS.t785 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1350 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK.t70 VSS.t597 VSS.t596 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1351 VDD 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A a_7215_10149# VDD.t510 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1352 VDD Q2.t20 a_15865_4557# VDD.t2425 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1353 VDD 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A a_11191_5901# VDD.t353 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1354 VDD OR_magic_1.VOUT.t19 divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT VDD.t2517 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1355 DFF_magic_0.tg_magic_2.OUT CLK.t71 DFF_magic_0.tg_magic_1.IN.t7 VSS.t595 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1356 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_2749_2092# VDD.t488 VDD.t371 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1357 a_21381_8741# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B a_21381_10149# VDD.t171 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1358 VSS p3_gen_magic_0.xnor_magic_1.B.t8 a_1957_n7648# VSS.t1445 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1359 VSS 7b_counter_0.MDFF_7.tspc2_magic_0.Q a_23802_1059# VSS.t374 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1360 a_15865_9774# 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A a_16065_9774# VSS.t267 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1361 divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.CLK.t13 VDD.t1997 VDD.t1996 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1362 VDD p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.P3.t3 VDD.t38 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1363 a_13553_n2115# p2_gen_magic_0.3_inp_AND_magic_0.B a_13769_n2115# VSS.t688 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1364 VDD D2_4.t16 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT VDD.t2274 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1365 VSS a_23258_1746# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B VSS.t248 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1366 VDD 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A a_11191_4932# VDD.t520 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1367 VDD mux_magic_0.IN2.t11 a_32616_n2458# VDD.t2151 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1368 a_27234_552# Q3.t22 VDD.t2298 VDD.t2297 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1369 VSS LD.t56 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A VSS.t1076 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1370 a_14556_n8142# p3_gen_magic_0.AND2_magic_1.A VDD.t1417 VDD.t1416 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1371 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN CLK.t72 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT VSS.t594 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1372 p3_gen_magic_0.3_inp_AND_magic_0.VOUT a_13353_n6613# VDD.t1133 VDD.t1132 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1373 a_9212_5956# 7b_counter_0.MDFF_5.tspc2_magic_0.D VSS.t464 VSS.t463 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1374 VSS D2_3.t17 a_5470_n1973# VSS.t1466 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1375 VDD mux_magic_0.IN1.t13 divide_by_2_1.tg_magic_2.IN VDD.t2361 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1376 a_21381_4932# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A VDD.t859 VDD.t855 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1377 VSS Q6.t19 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT VSS.t1269 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1378 DFF_magic_0.tg_magic_3.CLK CLK.t73 VDD.t2610 VDD.t2609 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1379 a_26038_4932# 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A VDD.t389 VDD.t383 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1380 DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK.t74 VSS.t593 VSS.t592 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1381 7b_counter_0.MDFF_0.tspc2_magic_0.Q 7b_counter_0.MDFF_0.QB.t8 VDD.t2448 VDD.t2441 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1382 VDD divide_by_2_0.tg_magic_3.CLK.t16 divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT VDD.t1823 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1383 VDD p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8643_n1042# VDD.t1731 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1384 a_11191_684# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A VDD.t346 VDD.t345 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1385 VSS D2_1.t25 a_16065_7470# VSS.t550 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1386 VSS 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t6 a_4651_3947# VSS.t1434 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1387 VDD 7b_counter_0.DFF_magic_0.Q.t15 DFF_magic_0.D VDD.t2106 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1388 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT CLK.t75 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t0 VSS.t591 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1389 VDD Q3.t23 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT VDD.t2303 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1390 a_9412_739# 7b_counter_0.MDFF_4.tspc2_magic_0.D VDD.t1784 VDD.t1783 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1391 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK.t76 VDD.t2616 VDD.t2615 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1392 VSS 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A a_21381_8741# VSS.t102 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1393 VDD LD.t57 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A VDD.t1849 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1394 VSS p2_gen_magic_0.3_inp_AND_magic_0.C.t7 a_13769_n2115# VSS.t1526 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1395 a_1409_8579# D2_7.t15 VSS.t1136 VSS.t630 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1396 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t85 VDD.t1602 VDD.t1601 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1397 7b_counter_0.MDFF_5.LD a_29512_8496.t17 VDD.t1194 VDD.t1187 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1398 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT D2_1.t26 VDD.t1333 VDD.t1332 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1399 VDD 7b_counter_0.MDFF_5.LD.t62 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A VDD.t1251 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1400 p3_gen_magic_0.xnor_magic_6.OUT D2_6.t15 a_8523_n8095# VDD.t65 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1401 a_17405_684# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A VDD.t196 VDD.t195 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1402 a_1209_3363# LD.t58 a_1409_3363# VSS.t1063 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1403 VSS p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t3 VSS.t679 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1404 a_17405_684# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A VDD.t194 VDD.t193 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1405 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t86 VDD.t1603 VDD.t1567 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1406 VDD OR_magic_2.VOUT.t15 divide_by_2_0.tg_magic_3.CLK.t2 VDD.t743 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1407 a_17405_5901# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A VDD.t2210 VDD.t2209 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1408 a_17405_7309# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_17405_5901# VDD.t627 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1409 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t87 VDD.t1604 VDD.t1569 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1410 VDD 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t7 a_4496_4393# VDD.t876 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1411 a_1209_8579# LD.t59 VDD.t1903 VDD.t1902 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1412 DFF_magic_0.tg_magic_0.IN DFF_magic_0.tg_magic_1.IN.t15 VSS.t44 VSS.t43 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1413 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B a_15865_2253# VSS.t173 VSS.t172 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1414 a_23352_n5390# p3_gen_magic_0.P3.t12 a_23352_n6798# VDD.t190 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1415 7b_counter_0.3_inp_AND_magic_0.VOUT a_23985_7877# VDD.t1759 VDD.t1758 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1416 a_23258_1746# 7b_counter_0.MDFF_4.LD.t88 VDD.t1606 VDD.t1605 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1417 VDD DFF_magic_0.tg_magic_1.IN.t16 DFF_magic_0.tg_magic_0.IN VDD.t59 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1418 a_17405_8741# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B a_17405_10149# VDD.t864 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1419 a_16386_n8142# p3_gen_magic_0.xnor_magic_5.OUT.t6 a_16186_n8142# VSS.t71 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1420 VDD p3_gen_magic_0.3_inp_AND_magic_0.A a_13353_n6613# VDD.t902 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1421 a_4235_3947# 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t8 a_4496_4877# VDD.t2452 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1422 VSS 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_11279_1124# VSS.t227 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1423 a_17405_3524# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B a_17405_4932# VDD.t160 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1424 a_12174_n3150# p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT VSS.t223 VSS.t222 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1425 a_4496_9609# 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t9 VDD.t2014 VDD.t1448 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1426 divide_by_2_0.tg_magic_0.IN divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.OUT VDD.t953 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1427 p3_gen_magic_0.xnor_magic_1.B D2_1.t27 VDD.t1335 VDD.t1334 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1428 VSS D2_4.t17 a_1975_n1973# VSS.t1321 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1429 a_1209_4557# 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A a_1409_4557# VSS.t85 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1430 a_8523_n8579# p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT VDD.t310 VDD.t227 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1431 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t15 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.t0 VSS.t1391 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1432 VDD Q6.t20 a_1209_6275# VDD.t2185 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1433 a_8825_6886# a_8713_6842# VSS.t366 VSS.t365 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1434 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A LD.t60 VSS.t1079 VSS.t1069 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1435 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t63 VSS.t787 VSS.t786 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1436 7b_counter_0.DFF_magic_0.tg_magic_2.IN 7b_counter_0.DFF_magic_0.Q.t16 VSS.t1221 VSS.t1220 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1437 a_23352_n6798# p3_gen_magic_0.P3.t13 a_23352_n5390# VDD.t1456 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1438 a_8411_3319# 7b_counter_0.MDFF_4.LD.t89 a_8955_3363# VSS.t926 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1439 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t64 VSS.t788 VSS.t776 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1440 a_23207_5815# Q2.t21 a_22991_5815# VDD.t2414 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1441 a_5054_n6024# D2_3.t18 p3_gen_magic_0.xnor_magic_4.OUT VDD.t400 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1442 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.OUT VDD.t1767 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1443 a_2749_5900# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A VDD.t426 VDD.t425 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1444 a_2749_8740# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B a_2749_10148# VDD.t67 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1445 a_20171_1669# a_19152_1223# VSS.t68 VSS.t67 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1446 DFF_magic_0.tg_magic_2.IN DFF_magic_0.tg_magic_3.CLK.t17 DFF_magic_0.tg_magic_2.OUT VSS.t1510 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1447 a_9689_1669# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t9 VSS.t1519 VSS.t1518 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1448 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t65 VDD.t1271 VDD.t1219 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1449 a_12387_1746# D2_6.t16 VDD.t1356 VDD.t1355 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1450 7b_counter_0.MDFF_3.tspc2_magic_0.D a_2749_8740# VSS.t50 VSS.t49 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1451 a_1209_3363# LD.t61 VDD.t1905 VDD.t1904 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1452 VDD 7b_counter_0.MDFF_5.LD.t66 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A VDD.t1272 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1453 a_6725_5900# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B a_6725_7308# VDD.t102 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1454 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT VSS.t716 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1455 a_7215_4932# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B a_7303_3480# VDD.t817 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1456 a_30365_3514# P2.t11 a_30365_4922# VDD.t2224 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1457 a_5036_n8095# D2_7.t16 p3_gen_magic_0.xnor_magic_5.OUT.t0 VDD.t759 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1458 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q2.t22 VDD.t2429 VDD.t2428 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1459 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK CLK.t77 VDD.t2614 VDD.t2613 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1460 7b_counter_0.3_inp_AND_magic_0.C Q3.t24 VSS.t1348 VSS.t1347 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1461 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B a_15865_8580# VDD.t397 VDD.t396 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1462 VSS CLK.t78 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VSS.t588 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1463 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN CLK.t79 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT VSS.t587 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1464 a_8411_8536# 7b_counter_0.MDFF_5.LD.t67 VDD.t1276 VDD.t1275 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1465 a_9412_5956# 7b_counter_0.MDFF_5.tspc2_magic_0.D VDD.t885 VDD.t884 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1466 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT divide_by_2_0.tg_magic_1.IN.t10 VDD.t895 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1467 VDD OR_magic_1.VOUT.t20 divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT VDD.t2520 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1468 a_5185_7469# LD.t62 VDD.t1907 VDD.t1906 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1469 VDD 7b_counter_0.MDFF_4.LD.t90 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A VDD.t1542 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1470 a_8411_4513# 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A a_8955_4557# VSS.t310 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1471 a_12174_n4081# p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.AND2_magic_1.A VDD.t442 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1472 a_21381_8741# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B a_21381_10149# VDD.t1126 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1473 a_5036_n3597# Q6.t21 VDD.t2188 VDD.t265 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1474 VDD p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t6 VDD.t1086 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1475 VDD OR_magic_2.A.t18 a_23352_n5390# VDD.t2338 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1476 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t91 VDD.t1609 VDD.t1581 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1477 a_1975_n6471# p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_3.OUT.t3 VSS.t302 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1478 VDD 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A a_11191_4932# VDD.t517 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1479 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_3.t19 VDD.t2484 VDD.t2483 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1480 VSS 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B a_26126_1124# VSS.t406 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1481 p3_gen_magic_0.xnor_magic_1.B D2_1.t28 VSS.t815 VSS.t814 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1482 a_15865_9774# CLK.t80 VDD.t2612 VDD.t2611 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1483 DFF_magic_0.tg_magic_3.CLK CLK.t81 VDD.t2618 VDD.t2617 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1484 VSS 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B a_22150_1124# VSS.t251 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1485 a_9412_5956# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t9 a_9212_5956# VDD.t912 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1486 VSS CLK.t82 a_1409_2253# VSS.t584 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1487 VDD a_1209_7469# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B VDD.t139 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1488 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t18 7b_counter_0.DFF_magic_0.D VSS.t1182 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1489 DFF_magic_0.tg_magic_2.OUT CLK.t83 DFF_magic_0.tg_magic_1.IN.t6 VSS.t583 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1490 VDD 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A a_1209_1059# VDD.t811 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1491 p3_gen_magic_0.xnor_magic_1.OUT Q7.t16 a_1541_n7648# VSS.t854 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1492 a_15865_3363# CLK.t84 VDD.t2625 VDD.t2624 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1493 divide_by_2_0.tg_magic_3.IN OR_magic_2.VOUT.t16 divide_by_2_0.tg_magic_1.IN.t1 VSS.t387 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1494 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT Q4.t20 VSS.t988 VSS.t987 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1495 a_1409_1059# 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A a_1209_1059# VSS.t426 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1496 a_4496_4393# a_4235_3947# a_4651_3947# VSS.t154 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1497 VDD Q5.t22 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT VDD.t246 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1498 a_22150_1124# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B a_22062_684# VDD.t475 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1499 7b_counter_0.DFF_magic_0.tg_magic_3.CLK CLK.t85 VDD.t2623 VDD.t2622 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1500 divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT OR_magic_1.VOUT.t21 VDD.t2524 VDD.t2523 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1501 VDD CLK.t86 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK VDD.t2619 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1502 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t0 VDD.t663 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1503 DFF_magic_0.tg_magic_2.IN DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT DFF_magic_0.tg_magic_2.OUT VDD.t1001 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1504 VSS OR_magic_2.VOUT.t17 divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT VSS.t388 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1505 a_21381_10149# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A VDD.t174 VDD.t173 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1506 7b_counter_0.MDFF_4.LD a_31440_8496.t16 VDD.t28 VDD.t22 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1507 VSS CLK.t87 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VSS.t580 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1508 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN p3_gen_magic_0.P3.t14 VDD.t1466 VDD.t1465 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1509 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT VDD.t286 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1510 a_6725_684# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A VDD.t1696 VDD.t420 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1511 a_1559_n6024# D2_4.t18 p3_gen_magic_0.xnor_magic_3.OUT VDD.t407 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1512 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_3.OUT VDD.t833 VDD.t832 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1513 a_5185_2253# LD.t63 VDD.t1909 VDD.t1908 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1514 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN CLK.t88 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT VSS.t579 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1515 VSS 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_11279_6341# VSS.t97 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1516 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t16 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT VSS.t1392 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1517 VSS 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t10 a_9689_6886# VSS.t476 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1518 a_15865_2253# 7b_counter_0.MDFF_4.LD.t92 a_16065_2253# VSS.t909 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1519 divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT OR_magic_2.VOUT.t18 VDD.t747 VDD.t746 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1520 a_12387_6963# 7b_counter_0.MDFF_5.LD.t68 a_12931_7470# VSS.t747 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1521 VDD a_1209_2253# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B VDD.t1744 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1522 a_16065_1059# 7b_counter_0.MDFF_1.QB.t8 VSS.t56 VSS.t55 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1523 VSS LD.t64 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A VSS.t1080 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1524 a_1541_n8095# p3_gen_magic_0.xnor_magic_1.B.t9 p3_gen_magic_0.xnor_magic_1.OUT VDD.t370 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1525 a_30365_4922# P2.t12 a_30365_3514# VDD.t977 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1526 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A a_19841_4557# VDD.t654 VDD.t653 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1527 VDD a_8713_6842# 7b_counter_0.MDFF_5.QB.t1 VDD.t717 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1528 VDD 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A a_26038_4932# VDD.t386 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1529 VDD LD.t65 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A VDD.t1862 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1530 a_19841_9774# 7b_counter_0.MDFF_6.tspc2_magic_0.Q VDD.t273 VDD.t272 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1531 VDD Q4.t21 a_23793_5904# VDD.t1661 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1532 DFF_magic_0.D 7b_counter_0.DFF_magic_0.Q.t17 VDD.t2110 VDD.t2109 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1533 a_21504_5904# Q7.t17 7b_counter_0.3_inp_AND_magic_0.B VDD.t1383 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1534 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT Q5.t23 VSS.t136 VSS.t135 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1535 VDD CLK.t89 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD.t2626 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1536 a_19152_5956# 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_18891_6886# VDD.t1751 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1537 VSS 7b_counter_0.MDFF_4.LD.t93 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A VSS.t927 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1538 VDD 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A a_2749_10148# VDD.t688 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1539 7b_counter_0.3_inp_AND_magic_0.C Q1.t21 VSS.t1205 VSS.t1204 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1540 VSS DFF_magic_0.tg_magic_3.CLK.t18 DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VSS.t1511 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1541 a_12931_6276# 7b_counter_0.MDFF_5.QB.t5 VSS.t485 VSS.t484 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1542 VSS 7b_counter_0.MDFF_4.LD.t94 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A VSS.t930 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1543 VSS p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t17 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VSS.t1393 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1544 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t95 VSS.t934 VSS.t933 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1545 a_15865_6276# 7b_counter_0.MDFF_6.QB.t9 VDD.t2252 VDD.t2251 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1546 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t7 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t6 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t7 VDD.t1052 pfet_03v3 ad=0.493p pd=3.12u as=0 ps=0 w=1.12u l=0.56u
X1547 a_1409_3363# D2_5.t15 VSS.t1546 VSS.t621 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1548 divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.CLK.t14 VSS.t1161 VSS.t1160 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1549 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t96 VSS.t936 VSS.t935 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1550 VDD p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5054_n1042# VDD.t293 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1551 7b_counter_0.MDFF_3.tspc2_magic_0.D a_2749_8740# VDD.t70 VDD.t68 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1552 a_19152_6440# a_18891_6886# a_19307_6886# VSS.t1020 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1553 a_8411_8536# D2_2.t19 VDD.t1948 VDD.t1947 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1554 VDD 7b_counter_0.3_inp_AND_magic_0.C a_23985_7877# VDD.t31 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1555 VDD a_15865_7470# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B VDD.t1127 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1556 Q3 a_21381_3524# VSS.t54 VSS.t52 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1557 a_1559_n5540# p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT VDD.t579 VDD.t578 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1558 p3_gen_magic_0.AND2_magic_1.A D2_5.t16 a_12174_n8095# VDD.t1414 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1559 7b_counter_0.DFF_magic_0.tg_magic_3.CLK CLK.t90 VDD.t2638 VDD.t2637 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1560 a_4496_10093# 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t10 a_4235_9163# VDD.t2015 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1561 a_19152_5956# 7b_counter_0.MDFF_6.tspc2_magic_0.D VDD.t203 VDD.t202 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1562 DFF_magic_0.tg_magic_0.IN CLK.t91 DFF_magic_0.tg_magic_3.OUT VSS.t578 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1563 a_4496_4877# 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t9 a_4235_3947# VDD.t2453 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1564 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t9 VSS.t715 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1565 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT VDD.t1028 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1566 a_23793_5904# Q4.t22 VDD.t1674 VDD.t1664 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1567 divide_by_2_0.tg_magic_2.IN divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.IN.t15 VDD.t997 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1568 VDD Q1.t22 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT VDD.t2083 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1569 VSS a_8411_8536# 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B VSS.t224 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1570 a_9059_n6471# p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_0.OUT VSS.t521 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1571 VDD p2_gen_magic_0.xnor_magic_6.OUT a_14556_n3644# VDD.t866 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1572 a_1409_4557# 7b_counter_0.MDFF_0.QB.t9 VSS.t1430 VSS.t1429 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1573 VSS D2_6.t17 a_8939_n3150# VSS.t826 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1574 a_1209_6275# Q6.t22 VDD.t2190 VDD.t2189 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1575 VDD Q4.t23 a_12174_n3597# VDD.t666 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1576 a_19841_3363# 7b_counter_0.MDFF_4.LD.t97 VDD.t1611 VDD.t1610 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1577 VDD 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A a_6725_684# VDD.t1693 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1578 VDD CLK.t92 a_1209_7469# VDD.t2634 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1579 a_5185_1059# 7b_counter_0.MDFF_0.tspc2_magic_0.Q VDD.t841 VDD.t840 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1580 divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.CLK.t15 VDD.t1999 VDD.t1998 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1581 a_8955_3363# D2_6.t18 VSS.t825 VSS.t824 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1582 VSS P2.t13 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN VSS.t1285 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1583 p2_gen_magic_0.3_inp_AND_magic_0.VOUT a_13353_n2115# VDD.t1108 VDD.t1107 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1584 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.IN.t15 VDD.t1766 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1585 a_15865_3363# 7b_counter_0.MDFF_4.LD.t98 VDD.t1613 VDD.t1612 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1586 a_26038_684# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B a_26126_1124# VDD.t1063 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1587 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A a_8411_4513# VDD.t965 VDD.t964 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1588 VSS Q1.t23 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT VSS.t1206 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1589 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT D2_1.t29 VSS.t817 VSS.t816 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1590 a_23985_7877# 7b_counter_0.3_inp_AND_magic_0.A a_24185_7877# VSS.t145 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1591 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT D2_5.t17 VDD.t2737 VDD.t2736 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1592 a_2749_684# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A VDD.t149 VDD.t144 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1593 VDD 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t19 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD.t2039 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1594 p2_gen_magic_0.3_inp_AND_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT VDD.t317 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1595 a_1209_9773# 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A VDD.t783 VDD.t782 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1596 a_6725_7308# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B a_6725_5900# VDD.t532 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1597 a_8643_n6024# D2_2.t20 p3_gen_magic_0.xnor_magic_0.OUT VDD.t980 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1598 7b_counter_0.DFF_magic_0.tg_magic_3.OUT CLK.t93 7b_counter_0.DFF_magic_0.tg_magic_0.IN VSS.t577 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1599 VDD D2_4.t19 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT VDD.t2277 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1600 a_30365_4922# OR_magic_2.A.t19 VDD.t2348 VDD.t2219 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1601 VSS a_8411_9730# 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A VSS.t189 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1602 VDD D2_2.t21 a_8411_8536# VDD.t1949 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1603 a_11292_n6613# p3_gen_magic_0.xnor_magic_0.OUT a_11492_n6613# VSS.t674 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1604 VDD Q2.t23 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT VDD.t2430 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1605 VSS 7b_counter_0.MDFF_4.LD.t99 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A VSS.t937 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1606 VDD p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t18 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD.t2393 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1607 VDD p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t16 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN VDD.t1424 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1608 a_8955_4557# 7b_counter_0.MDFF_4.tspc2_magic_0.Q VSS.t168 VSS.t167 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1609 a_13769_n6613# p3_gen_magic_0.3_inp_AND_magic_0.B a_13553_n6613# VSS.t471 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1610 VSS 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t20 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VSS.t1183 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1611 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_3.t20 VDD.t2486 VDD.t2485 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1612 a_23672_3947# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t10 7b_counter_0.MDFF_7.QB.t1 VSS.t894 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1613 VDD CLK.t94 a_1209_2253# VDD.t2631 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1614 p2_gen_magic_0.xnor_magic_6.OUT p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT a_8523_n4081# VDD.t861 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1615 a_16065_1059# 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A a_15865_1059# VSS.t305 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1616 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT CLK.t95 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t0 VSS.t576 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1617 VDD 7b_counter_0.MDFF_5.QB.t6 7b_counter_0.MDFF_5.tspc2_magic_0.Q VDD.t927 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1618 a_11492_n2115# p2_gen_magic_0.xnor_magic_0.OUT a_11292_n2115# VSS.t1011 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1619 a_12387_8536# 7b_counter_0.MDFF_5.LD.t69 VDD.t1278 VDD.t1277 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1620 p3_gen_magic_0.3_inp_AND_magic_0.A a_11292_n6613# VSS.t676 VSS.t674 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1621 VDD p2_gen_magic_0.xnor_magic_3.OUT.t7 a_11292_n2115# VDD.t2231 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1622 7b_counter_0.DFF_magic_0.D 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t21 7b_counter_0.DFF_magic_0.tg_magic_3.OUT VSS.t1186 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1623 VSS p3_gen_magic_0.xnor_magic_3.OUT.t7 a_11708_n6613# VSS.t233 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1624 a_8523_n3597# D2_6.t19 p2_gen_magic_0.xnor_magic_6.OUT VDD.t862 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1625 VDD 7b_counter_0.MDFF_3.tspc2_magic_0.D a_4496_10093# VDD.t1450 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1626 VDD 7b_counter_0.MDFF_4.tspc2_magic_0.D a_9412_739# VDD.t1778 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1627 VDD 7b_counter_0.MDFF_4.LD.t100 a_15865_3363# VDD.t1614 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1628 VDD a_15865_9774# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A VDD.t502 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1629 a_13769_n6613# p3_gen_magic_0.3_inp_AND_magic_0.B a_13553_n6613# VSS.t470 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1630 OUT1 a_34156_n2297# VSS.t221 VSS.t220 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1631 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT divide_by_2_1.tg_magic_2.IN VDD.t98 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1632 VDD a_11279_1124# 7b_counter_0.MDFF_4.tspc2_magic_0.D VDD.t1769 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1633 a_4651_3947# 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t10 VSS.t1438 VSS.t1437 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1634 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_3.OUT VSS.t435 VSS.t434 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1635 DFF_magic_0.D 7b_counter_0.DFF_magic_0.Q.t18 VDD.t2098 VDD.t2097 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1636 VDD Q7.t18 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT VDD.t1393 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1637 VDD a_11279_6341# 7b_counter_0.MDFF_5.tspc2_magic_0.D VDD.t879 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1638 a_5036_n3150# p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT VSS.t197 VSS.t196 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1639 VDD 7b_counter_0.MDFF_7.tspc2_magic_0.D a_24259_4877# VDD.t2318 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1640 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q1.t24 VSS.t1210 VSS.t1209 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1641 VSS 7b_counter_0.MDFF_6.tspc2_magic_0.D a_18891_6886# VSS.t115 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1642 VSS 7b_counter_0.MDFF_4.LD.t101 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A VSS.t940 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1643 VDD p2_gen_magic_0.3_inp_AND_magic_0.A a_13353_n2115# VDD.t763 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1644 VDD a_31440_8496.t17 7b_counter_0.MDFF_4.LD.t8 VDD.t24 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1645 VSS LD.t66 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A VSS.t1083 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1646 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT Q6.t23 VDD.t2192 VDD.t2191 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1647 DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK.t96 VDD.t2630 VDD.t2629 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1648 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_2.t22 VDD.t1953 VDD.t1952 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1649 VSS LD.t67 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A VSS.t1086 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1650 VSS p3_gen_magic_0.xnor_magic_3.OUT.t8 a_11708_n6613# VSS.t233 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1651 VDD.t1058 VDD.t1057 VDD.t1058 VDD.t766 pfet_03v3 ad=0.493p pd=3.12u as=0 ps=0 w=1.12u l=0.56u
X1652 a_17405_684# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B a_17405_2092# VDD.t2217 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1653 a_17405_4932# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A VDD.t159 VDD.t156 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1654 VDD a_15865_1059# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A VDD.t595 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1655 a_15865_6276# 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A VDD.t328 VDD.t327 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1656 VDD p3_gen_magic_0.xnor_magic_5.OUT.t7 a_16186_n8142# VDD.t106 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1657 VSS p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t19 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VSS.t1396 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1658 VSS 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t15 7b_counter_0.DFF_magic_0.tg_magic_0.IN VSS.t479 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1659 VDD Q4.t24 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT VDD.t1677 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1660 a_19841_8580# 7b_counter_0.MDFF_5.LD.t70 a_20041_8580# VSS.t789 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1661 divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT OR_magic_2.VOUT.t19 VDD.t749 VDD.t748 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1662 p2_gen_magic_0.3_inp_AND_magic_0.B a_14556_n3644# VSS.t347 VSS.t346 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1663 VDD divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_1.IN.t6 VDD.t829 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1664 OUT1 a_34156_n2297# VDD.t439 VDD.t48 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1665 VDD Q1.t25 a_8643_n6024# VDD.t987 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1666 VDD a_27234_4513# 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A VDD.t660 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1667 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A LD.t68 VDD.t1913 VDD.t1912 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1668 a_9689_6886# a_9212_5956# a_8713_6842# VSS.t363 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1669 VSS 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A a_17405_8741# VSS.t537 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1670 VDD D2_1.t30 a_15865_7470# VDD.t1336 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1671 VSS D2_6.t20 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT VSS.t831 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1672 DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT DFF_magic_0.D.t1 VDD.t940 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1673 a_8643_n5540# p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT VDD.t991 VDD.t990 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1674 VSS 7b_counter_0.MDFF_1.QB.t9 a_16065_1059# VSS.t57 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1675 VDD 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_19841_4557# VDD.t648 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1676 VSS 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_19307_1669# VSS.t502 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1677 VSS divide_by_2_0.tg_magic_3.IN.t22 mux_magic_0.IN2.t4 VSS.t10 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1678 VSS CLK.t97 DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VSS.t573 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1679 p2_gen_magic_0.3_inp_AND_magic_0.A a_11292_n2115# VDD.t364 VDD.t363 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1680 a_4496_4877# 7b_counter_0.MDFF_0.tspc2_magic_0.D VDD.t872 VDD.t871 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1681 VDD Q3.t25 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT VDD.t2306 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1682 Q3 a_21381_3524# VDD.t81 VDD.t79 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1683 mux_magic_0.IN1 divide_by_2_1.tg_magic_3.IN.t23 VSS.t77 VSS.t76 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1684 a_5036_n4081# p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_5.OUT VDD.t398 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1685 7b_counter_0.3_inp_AND_magic_0.B Q7.t19 a_21504_5904# VDD.t1384 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1686 VSS D2_3.t21 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT VSS.t1469 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1687 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_4.t20 VDD.t2281 VDD.t2280 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1688 VDD p2_gen_magic_0.xnor_magic_1.OUT.t8 a_16186_n3644# VDD.t2406 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1689 a_12387_9730# 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A VDD.t1103 VDD.t1102 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1690 divide_by_2_0.tg_magic_2.IN mux_magic_0.IN2.t12 VDD.t2155 VDD.t2154 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1691 7b_counter_0.MDFF_3.tspc2_magic_0.Q 7b_counter_0.MDFF_3.QB VDD.t623 VDD.t621 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1692 VDD CLK.t98 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD.t2645 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1693 divide_by_2_0.tg_magic_3.OUT OR_magic_2.VOUT.t20 divide_by_2_0.tg_magic_0.IN VSS.t391 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1694 a_19841_9774# 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A a_20041_9774# VSS.t143 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1695 divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.CLK.t16 VDD.t2001 VDD.t2000 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1696 VDD Q5.t24 a_8523_n3597# VDD.t249 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1697 a_23258_552# 7b_counter_0.MDFF_7.tspc2_magic_0.Q VDD.t724 VDD.t723 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1698 a_8955_3363# 7b_counter_0.MDFF_4.LD.t102 a_8411_3319# VSS.t943 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1699 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A LD.t69 VDD.t1915 VDD.t1914 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1700 VSS 7b_counter_0.MDFF_5.QB.t7 a_12931_6276# VSS.t486 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1701 VDD DFF_magic_0.tg_magic_2.OUT OR_magic_2.A.t2 VDD.t1003 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1702 VDD 7b_counter_0.MDFF_1.tspc2_magic_0.D a_19152_739# VDD.t1020 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1703 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t103 VSS.t945 VSS.t944 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1704 VDD p3_gen_magic_0.xnor_magic_3.OUT.t9 a_11292_n6613# VDD.t452 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1705 DFF_magic_0.tg_magic_3.CLK CLK.t99 VSS.t572 VSS.t571 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1706 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT Q6.t24 VSS.t1273 VSS.t1272 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1707 VDD 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A a_15865_6276# VDD.t324 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1708 VSS 7b_counter_0.MDFF_4.LD.t104 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A VSS.t927 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1709 VSS 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A a_2749_8740# VSS.t215 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1710 a_1541_n3150# p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT VSS.t712 VSS.t711 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1711 VSS 7b_counter_0.MDFF_4.LD.t105 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A VSS.t948 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1712 VDD 7b_counter_0.MDFF_5.LD.t71 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A VDD.t1258 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1713 7b_counter_0.3_inp_AND_magic_0.VOUT a_23985_7877# VSS.t1023 VSS.t145 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1714 a_24259_4877# 7b_counter_0.MDFF_7.tspc2_magic_0.D VDD.t2317 VDD.t1472 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1715 VDD a_26126_1124# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t1 VDD.t1064 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1716 VDD 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A a_6725_5900# VDD.t537 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1717 a_27234_552# 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A VDD.t584 VDD.t583 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1718 VDD a_22150_1124# Q4.t1 VDD.t475 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1719 VDD divide_by_2_1.tg_magic_1.IN.t17 divide_by_2_1.tg_magic_0.IN VDD.t484 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1720 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t106 VSS.t951 VSS.t935 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1721 VDD 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A a_11191_10149# VDD.t277 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1722 VSS D2_2.t23 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT VSS.t1120 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1723 VDD a_8411_8536# 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B VDD.t443 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1724 VDD Q6.t25 a_21504_5904# VDD.t2163 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1725 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK.t100 VDD.t2644 VDD.t2643 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1726 VSS Q4.t25 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT VSS.t989 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1727 VDD 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A a_11191_684# VDD.t342 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1728 a_7303_3480# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A VSS.t513 VSS.t512 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1729 DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK.t101 VDD.t2642 VDD.t2641 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1730 a_8955_4557# 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A a_8411_4513# VSS.t309 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1731 a_8411_9730# 7b_counter_0.MDFF_5.tspc2_magic_0.Q VDD.t701 VDD.t700 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1732 VSS a_12387_8536# 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B VSS.t295 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1733 a_21381_4932# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A VDD.t858 VDD.t78 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1734 VSS DFF_magic_0.D.t30 a_29512_8496.t7 VSS.t1240 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1735 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_3.OUT VDD.t125 VDD.t124 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1736 VDD DFF_magic_0.D.t31 a_29512_8496.t8 VDD.t2117 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1737 VDD Q5.t25 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT VDD.t252 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1738 a_11492_n2115# p2_gen_magic_0.xnor_magic_0.OUT a_11292_n2115# VSS.t1011 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1739 VDD divide_by_2_1.tg_magic_3.CLK.t17 divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT VDD.t2002 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1740 a_1209_7469# CLK.t102 VDD.t2640 VDD.t2639 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1741 VSS D2_6.t21 a_8955_3363# VSS.t821 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1742 VDD a_7303_3480# Q6.t1 VDD.t526 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1743 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A a_12387_4513# VDD.t1139 VDD.t1138 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1744 VDD 7b_counter_0.MDFF_4.tspc2_magic_0.D a_9412_739# VDD.t1778 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1745 a_1541_n4081# p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_1.OUT.t1 VDD.t1149 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1746 a_24185_7877# 7b_counter_0.3_inp_AND_magic_0.B a_24401_7877# VSS.t25 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1747 VSS D2_4.t21 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT VSS.t1324 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1748 VDD 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t16 7b_counter_0.DFF_magic_0.tg_magic_0.IN VDD.t921 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1749 VSS D2_5.t18 a_12590_n3150# VSS.t1547 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1750 VDD Q2.t24 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT VDD.t2433 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1751 a_5470_n6471# p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_4.OUT VSS.t51 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1752 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p2_gen_magic_0.3_inp_AND_magic_0.VOUT.t3 VDD.t316 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1753 VSS a_7303_8697# Q2.t0 VSS.t879 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1754 a_14556_n8142# p3_gen_magic_0.AND2_magic_1.A a_14756_n8142# VSS.t867 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1755 a_6725_5900# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A VDD.t536 VDD.t533 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1756 a_5036_n8579# p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT VDD.t1727 VDD.t1726 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1757 VSS a_12387_9730# 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A VSS.t529 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1758 7b_counter_0.DFF_magic_0.tg_magic_0.IN CLK.t103 7b_counter_0.DFF_magic_0.tg_magic_3.OUT VSS.t570 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1759 a_12931_3363# CLK.t104 VSS.t569 VSS.t568 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1760 a_2749_5900# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A VDD.t424 VDD.t423 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1761 a_18891_6886# 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_19152_5956# VDD.t1750 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1762 VDD a_32616_n1264# mux_magic_0.OR_magic_0.A VDD.t944 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1763 a_23207_5815# Q2.t25 a_22991_5815# VDD.t2414 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1764 VDD 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 7b_counter_0.DFF_magic_0.Q.t3 VDD.t610 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1765 VSS D2_4.t22 a_27778_3363# VSS.t609 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1766 7b_counter_0.3_inp_AND_magic_0.C Q3.t26 a_23207_5815# VDD.t2284 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1767 VSS 7b_counter_0.MDFF_4.tspc2_magic_0.Q a_8955_4557# VSS.t164 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1768 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t22 VSS.t1188 VSS.t1187 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1769 VDD 7b_counter_0.MDFF_4.LD.t107 a_12387_3319# VDD.t1617 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1770 VSS 7b_counter_0.MDFF_4.LD.t108 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A VSS.t937 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1771 VDD 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A a_22062_684# VDD.t847 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1772 a_12931_7470# 7b_counter_0.MDFF_5.LD.t72 a_12387_6963# VSS.t756 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1773 DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT DFF_magic_0.D.t0 VDD.t939 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1774 a_1209_2253# CLK.t105 VDD.t2649 VDD.t2648 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1775 VDD p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT P2.t3 VDD.t2368 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1776 VSS 7b_counter_0.MDFF_4.LD.t109 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A VSS.t954 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1777 a_17405_8741# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B a_17405_10149# VDD.t863 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1778 a_17405_10149# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A VDD.t1034 VDD.t1033 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1779 VDD CLK.t106 a_12387_8536# VDD.t2658 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1780 a_17405_2092# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B a_17405_684# VDD.t2216 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1781 VSS CLK.t107 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VSS.t565 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1782 VDD divide_by_2_1.tg_magic_3.CLK.t18 divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT VDD.t2005 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1783 a_12931_4557# Q5.t26 VSS.t138 VSS.t137 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1784 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK VDD.t1152 VDD.t1151 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1785 a_24259_4877# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t12 a_24059_4877# VDD.t1474 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1786 a_23793_5904# Q5.t27 7b_counter_0.3_inp_AND_magic_0.A VDD.t220 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1787 divide_by_2_0.tg_magic_0.IN divide_by_2_0.tg_magic_1.IN.t17 VDD.t1413 VDD.t1412 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1788 VSS 7b_counter_0.MDFF_7.QB.t8 a_27778_4557# VSS.t3 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1789 p2_gen_magic_0.AND2_magic_1.A p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_12174_n4081# VDD.t441 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1790 a_1559_n1526# Q3.t27 VDD.t2309 VDD.t606 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1791 divide_by_2_1.tg_magic_2.IN mux_magic_0.IN1.t14 VDD.t2365 VDD.t2364 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1792 a_21381_10149# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A VDD.t172 VDD.t171 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1793 divide_by_2_1.tg_magic_3.IN OR_magic_1.VOUT.t22 divide_by_2_1.tg_magic_1.IN.t10 VSS.t1486 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1794 VDD Q3.t28 a_27234_552# VDD.t2310 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1795 VDD DFF_magic_0.D.t32 a_31440_8496.t4 VDD.t2122 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1796 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A LD.t70 VDD.t1916 VDD.t1914 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1797 VDD p3_gen_magic_0.xnor_magic_1.B.t10 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT VDD.t2462 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1798 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A LD.t71 VSS.t1089 VSS.t1057 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1799 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A LD.t72 VSS.t1091 VSS.t1090 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1800 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t73 VDD.t1282 VDD.t1281 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1801 a_11279_1124# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_11191_684# VDD.t449 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1802 VSS 7b_counter_0.MDFF_4.LD.t110 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A VSS.t940 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1803 7b_counter_0.DFF_magic_0.tg_magic_0.IN 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t17 VSS.t483 VSS.t482 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1804 VDD Q6.t26 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT VDD.t2195 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1805 a_12387_552# 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A a_12931_1059# VSS.t1384 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1806 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B a_15865_2253# VDD.t333 VDD.t332 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1807 VSS LD.t73 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A VSS.t1086 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1808 a_27778_3363# D2_4.t23 VSS.t1329 VSS.t606 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1809 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_7.t17 VDD.t1977 VDD.t1976 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1810 a_2749_10148# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A VDD.t689 VDD.t688 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1811 a_1541_n3597# Q7.t20 VDD.t1396 VDD.t806 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1812 VDD 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t11 a_8713_1625# VDD.t1775 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1813 a_2749_3524# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B VSS.t106 VSS.t105 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1814 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A a_27234_4513# VDD.t659 VDD.t658 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1815 VSS OR_magic_2.VOUT.t21 divide_by_2_0.tg_magic_3.CLK.t2 VSS.t392 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1816 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q2.t26 VSS.t1419 VSS.t1418 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1817 VDD 7b_counter_0.MDFF_4.tspc2_magic_0.D a_9412_739# VDD.t1775 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1818 Q7 a_6725_7308# VDD.t101 VDD.t100 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1819 DFF_magic_0.tg_magic_2.OUT DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT DFF_magic_0.tg_magic_2.IN VDD.t1000 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1820 VDD DFF_magic_0.tg_magic_3.CLK.t19 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD.t2701 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1821 a_12387_9730# Q1.t26 VDD.t2089 VDD.t2088 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1822 a_19307_1669# a_18891_1669# a_19152_1223# VSS.t62 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1823 VDD 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A a_7215_4932# VDD.t969 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1824 a_2749_684# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A VDD.t148 VDD.t147 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1825 a_17405_2092# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B a_17405_684# VDD.t2215 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1826 VDD 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A a_12387_5769# VDD.t557 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1827 VDD Q2.t27 a_5054_n6024# VDD.t75 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1828 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A a_15865_1059# VDD.t594 VDD.t593 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1829 VDD 7b_counter_0.3_inp_AND_magic_0.A a_23985_7877# VDD.t267 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1830 a_27778_4557# 7b_counter_0.MDFF_7.QB.t9 VSS.t7 VSS.t6 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1831 a_19841_3363# D2_3.t22 VDD.t2488 VDD.t2487 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1832 P2 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT VDD.t2367 VDD.t2366 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1833 VDD 7b_counter_0.MDFF_4.LD.t111 a_27234_3319# VDD.t1620 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1834 a_14556_n8142# p3_gen_magic_0.xnor_magic_6.OUT VDD.t935 VDD.t934 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1835 a_5054_n5540# p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT VDD.t74 VDD.t73 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1836 divide_by_2_1.tg_magic_0.IN divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.OUT VDD.t1135 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1837 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_17405_3524# VSS.t371 VSS.t370 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1838 a_22991_5815# Q1.t27 VDD.t2090 VDD.t2060 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1839 VSS 7b_counter_0.3_inp_AND_magic_0.C a_24401_7877# VSS.t25 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1840 a_16186_n8142# p3_gen_magic_0.xnor_magic_5.OUT.t8 a_16386_n8142# VSS.t72 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1841 VDD Q6.t27 a_5036_n8095# VDD.t1728 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1842 p2_gen_magic_0.3_inp_AND_magic_0.A p2_gen_magic_0.3_inp_AND_magic_0.A p2_gen_magic_0.3_inp_AND_magic_0.A VDD.t766 pfet_03v3 ad=0.493p pd=3.12u as=1.97p ps=12.5u w=1.12u l=0.56u
X1843 VSS 7b_counter_0.MDFF_4.LD.t112 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A VSS.t959 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1844 VSS 7b_counter_0.MDFF_4.LD.t113 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A VSS.t948 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1845 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_8643_n1042# VDD.t457 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1846 VDD a_19841_8580# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B VDD.t1121 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1847 VDD a_7303_8697# Q2.t1 VDD.t1440 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1848 VDD 7b_counter_0.MDFF_5.LD.t74 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A VDD.t1241 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1849 VDD p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT a_12174_n8579# VDD.t633 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1850 VSS 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B a_7303_3480# VSS.t427 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1851 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_7.t18 VSS.t1138 VSS.t1137 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1852 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_2.OUT VDD.t2691 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1853 p2_gen_magic_0.3_inp_AND_magic_0.B a_14556_n3644# VDD.t679 VDD.t678 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1854 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT D2_1.t31 VDD.t1340 VDD.t1339 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1855 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT VSS.t1035 VSS.t1034 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1856 VDD 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A a_21381_4932# VDD.t855 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1857 a_27234_552# 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A a_27778_1059# VSS.t303 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1858 VDD.t1056 VDD.t1054 VDD.t1056 VDD.t1055 pfet_03v3 ad=0.493p pd=3.12u as=0 ps=0 w=1.12u l=0.56u
X1859 VDD D2_3.t23 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT VDD.t2489 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1860 VDD a_12387_8536# 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B VDD.t565 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1861 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN VDD.t285 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1862 VDD a_11279_3480# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t1 VDD.t1144 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1863 a_30365_4922# OR_magic_2.A.t20 VDD.t2349 VDD.t2329 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1864 a_5054_n6471# p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT VSS.t199 VSS.t198 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1865 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT VDD.t1810 VDD.t1809 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1866 a_8643_n1526# Q1.t28 VDD.t2091 VDD.t1734 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1867 p3_gen_magic_0.P3 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT VDD.t37 VDD.t36 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1868 VDD p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1559_n1042# VDD.t603 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1869 divide_by_2_1.tg_magic_3.CLK OR_magic_1.VOUT.t23 VSS.t1488 VSS.t1487 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1870 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A a_1209_9773# VSS.t349 VSS.t348 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1871 VDD p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t20 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD.t2396 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1872 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q1.t29 VDD.t2093 VDD.t2092 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1873 VSS a_11279_8697# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t0 VSS.t460 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1874 VSS D2_7.t19 a_5452_n7648# VSS.t1139 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1875 VSS Q7.t21 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT VSS.t855 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1876 VDD a_27567_8496.t16 LD.t7 VDD.t1178 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1877 p3_gen_magic_0.3_inp_AND_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT VDD.t1714 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1878 VSS 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_5385_6275# VSS.t288 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1879 VSS CLK.t108 a_12931_3363# VSS.t548 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1880 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t75 VDD.t1285 VDD.t1281 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1881 mux_magic_0.OR_magic_0.A a_32616_n1264# VDD.t943 VDD.t942 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1882 7b_counter_0.DFF_magic_0.Q 7b_counter_0.DFF_magic_0.tg_magic_2.OUT VDD.t609 VDD.t608 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1883 p3_gen_magic_0.xnor_magic_1.B D2_1.t32 VDD.t1342 VDD.t1341 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1884 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t17 VDD.t1428 VDD.t1427 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1885 VDD D2_2.t24 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT VDD.t1954 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1886 VDD D2_3.t24 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT VDD.t2492 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1887 a_27778_3363# 7b_counter_0.MDFF_4.LD.t114 a_27234_3319# VSS.t924 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1888 a_8523_n8579# p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_6.OUT VDD.t64 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1889 VDD 7b_counter_0.MDFF_4.QB.t10 7b_counter_0.MDFF_4.tspc2_magic_0.Q VDD.t1429 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1890 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t8 VDD.t1713 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1891 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT Q4.t26 VDD.t1681 VDD.t1680 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1892 OR_magic_2.VOUT a_23352_n6798# VDD.t191 VDD.t190 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1893 VDD p2_gen_magic_0.xnor_magic_3.OUT.t8 a_11292_n2115# VDD.t2231 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1894 VSS a_12387_1746# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B VSS.t205 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1895 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t115 VDD.t1623 VDD.t1554 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1896 divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.CLK.t17 VDD.t1827 VDD.t1826 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1897 a_18891_1669# 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_19152_739# VDD.t957 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1898 7b_counter_0.DFF_magic_0.Q 7b_counter_0.DFF_magic_0.tg_magic_2.OUT VSS.t313 VSS.t312 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1899 VDD D2_5.t19 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT VDD.t2738 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1900 a_2749_3524# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B a_2749_4932# VDD.t178 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1901 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q3.t29 VDD.t2314 VDD.t2313 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1902 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t116 VSS.t965 VSS.t964 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1903 VSS 7b_counter_0.3_inp_AND_magic_0.C a_24401_7877# VSS.t20 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1904 divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT OR_magic_2.VOUT.t22 VSS.t396 VSS.t395 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1905 VDD 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t23 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD.t2042 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1906 p3_gen_magic_0.3_inp_AND_magic_0.A a_11292_n6613# VDD.t1077 VDD.t1076 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1907 DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT DFF_magic_0.tg_magic_3.CLK.t20 VDD.t2705 VDD.t2704 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1908 a_6725_2092# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B a_6725_684# VDD.t419 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1909 VSS D2_7.t20 a_5385_7469# VSS.t1142 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1910 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A a_5185_1059# VDD.t1687 VDD.t1686 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1911 VSS Q5.t28 a_12931_4557# VSS.t139 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1912 7b_counter_0.MDFF_6.tspc2_magic_0.D a_17405_7309# VDD.t630 VDD.t628 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1913 a_13353_n6613# p3_gen_magic_0.3_inp_AND_magic_0.B VDD.t1796 VDD.t1795 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1914 a_26126_3480# 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A VSS.t193 VSS.t192 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1915 VDD 7b_counter_0.MDFF_7.QB.t10 7b_counter_0.MDFF_7.tspc2_magic_0.Q VDD.t5 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1916 VDD p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t7 VDD.t1806 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1917 VDD CLK.t109 DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD.t2655 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1918 a_27778_4557# 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A a_27234_4513# VSS.t1024 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1919 a_17405_7309# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_17405_5901# VDD.t626 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1920 divide_by_2_1.tg_magic_1.IN OR_magic_1.VOUT.t24 divide_by_2_1.tg_magic_3.IN.t6 VSS.t1489 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1921 a_18891_6886# 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_19152_5956# VDD.t1749 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1922 a_16186_n8142# p3_gen_magic_0.xnor_magic_1.OUT.t7 VDD.t53 VDD.t52 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1923 a_34156_n2297# mux_magic_0.OR_magic_0.B a_34156_n889# VDD.t46 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1924 a_4496_10093# 7b_counter_0.MDFF_3.tspc2_magic_0.D VDD.t1449 VDD.t1448 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1925 a_1559_n6471# p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT VSS.t204 VSS.t203 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1926 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN VDD.t1027 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1927 VSS Q3.t30 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT VSS.t1349 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1928 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A LD.t74 VDD.t1917 VDD.t1837 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1929 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A LD.t75 VSS.t1094 VSS.t1090 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1930 VDD a_26126_3480# 7b_counter_0.MDFF_7.tspc2_magic_0.D VDD.t777 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1931 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A LD.t76 VDD.t1919 VDD.t1918 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1932 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_17405_3524# VDD.t721 VDD.t720 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1933 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t76 VDD.t1287 VDD.t1286 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1934 VDD DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_1.IN.t2 VDD.t1041 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1935 a_8713_1625# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t12 VDD.t2713 VDD.t1783 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1936 VDD a_5185_6275# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A VDD.t187 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1937 divide_by_2_1.tg_magic_2.IN divide_by_2_1.tg_magic_3.CLK.t19 divide_by_2_1.tg_magic_3.IN.t12 VSS.t1162 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1938 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT DFF_magic_0.tg_magic_3.CLK.t21 VDD.t2707 VDD.t2706 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1939 7b_counter_0.MDFF_6.tspc2_magic_0.Q 7b_counter_0.MDFF_6.QB.t10 VDD.t2253 VDD.t2246 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1940 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_2749_7308# VSS.t499 VSS.t49 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1941 VDD p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT a_8523_n8579# VDD.t237 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1942 VDD divide_by_2_0.tg_magic_3.CLK.t18 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT VDD.t1828 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1943 a_7215_4932# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B a_7303_3480# VDD.t816 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1944 a_23352_n5390# OR_magic_2.A.t21 VDD.t2350 VDD.t2338 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1945 a_12387_1746# 7b_counter_0.MDFF_4.LD.t117 VDD.t1625 VDD.t1624 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1946 Q5 a_6725_2092# VDD.t1031 VDD.t1030 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1947 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_3.OUT VDD.t828 VDD.t827 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1948 VDD CLK.t110 a_27234_1746# VDD.t2652 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1949 a_5054_n5540# p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_4.OUT VDD.t400 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1950 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B a_19841_3363# VSS.t219 VSS.t218 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1951 VDD 7b_counter_0.MDFF_4.LD.t118 a_19841_3363# VDD.t1626 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1952 VSS a_27234_1746# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B VSS.t245 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1953 VDD P2.t14 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN VDD.t2225 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1954 VDD p2_gen_magic_0.3_inp_AND_magic_0.A a_13353_n2115# VDD.t763 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1955 VDD 7b_counter_0.DFF_magic_0.Q.t19 7b_counter_0.DFF_magic_0.tg_magic_2.IN VDD.t2099 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1956 a_1209_9773# 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A a_1409_9773# VSS.t412 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1957 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.IN.t6 VDD.t894 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1958 a_23258_1746# 7b_counter_0.MDFF_4.LD.t119 a_23802_2253# VSS.t966 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1959 divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.CLK.t19 VSS.t1049 VSS.t1048 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1960 VDD mux_magic_0.IN2.t13 divide_by_2_0.tg_magic_2.IN VDD.t2156 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1961 7b_counter_0.DFF_magic_0.tg_magic_2.OUT CLK.t111 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t6 VSS.t563 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1962 VDD a_11279_8697# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t1 VDD.t165 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1963 a_12590_n7648# p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p3_gen_magic_0.AND2_magic_1.A VSS.t327 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1964 VDD 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A a_2749_684# VDD.t144 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1965 a_1209_1059# Q4.t27 VDD.t1683 VDD.t1682 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1966 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_2749_2092# VDD.t487 VDD.t371 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1967 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK VSS.t714 VSS.t713 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1968 a_12174_n3597# D2_5.t20 p2_gen_magic_0.AND2_magic_1.A VDD.t442 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1969 a_22062_684# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B a_22150_1124# VDD.t474 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1970 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A a_19841_4557# VSS.t339 VSS.t338 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1971 a_11292_n6613# p3_gen_magic_0.xnor_magic_4.OUT VDD.t490 VDD.t489 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1972 mux_magic_0.AND2_magic_0.A D2_1.t33 VDD.t1343 VDD.t1302 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1973 VDD 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_5185_1059# VDD.t837 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1974 VDD OR_magic_2.VOUT.t23 divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT VDD.t750 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1975 a_2749_8740# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B a_2749_10148# VDD.t66 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1976 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t9 VDD.t2690 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1977 VDD 7b_counter_0.MDFF_4.LD.t120 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A VDD.t1528 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1978 a_12387_3319# CLK.t112 VDD.t2651 VDD.t2650 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1979 VDD divide_by_2_0.tg_magic_3.IN.t23 mux_magic_0.IN2 VDD.t17 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1980 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t11 VDD.t2378 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1981 a_11191_5901# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A VDD.t354 VDD.t353 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1982 a_9412_5956# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t11 a_9212_5956# VDD.t912 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1983 a_27234_1746# 7b_counter_0.MDFF_4.LD.t121 VDD.t1632 VDD.t1631 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1984 a_4651_9163# a_4235_9163# a_4496_9609# VSS.t186 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1985 Q1 a_21381_8741# VDD.t547 VDD.t546 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1986 VDD D2_6.t22 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT VDD.t1359 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1987 7b_counter_0.MDFF_0.tspc2_magic_0.Q 7b_counter_0.MDFF_0.QB.t10 VSS.t1432 VSS.t1431 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1988 VSS 7b_counter_0.3_inp_AND_magic_0.C a_24401_7877# VSS.t20 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1989 a_23802_1059# 7b_counter_0.MDFF_7.tspc2_magic_0.Q VSS.t373 VSS.t372 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1990 7b_counter_0.MDFF_3.tspc2_magic_0.Q 7b_counter_0.MDFF_3.QB VDD.t622 VDD.t621 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1991 VSS mux_magic_0.OR_magic_0.A a_34156_n2297# VSS.t431 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1992 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK CLK.t113 VDD.t2662 VDD.t2661 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1993 7b_counter_0.DFF_magic_0.D 7b_counter_0.DFF_magic_0.Q.t20 VDD.t2103 VDD.t2102 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1994 a_32616_n2458# D2_1.t34 VDD.t1345 VDD.t1344 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1995 VSS 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B a_11279_3480# VSS.t227 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1996 VDD 7b_counter_0.MDFF_3.QB a_1209_9773# VDD.t618 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1997 p2_gen_magic_0.xnor_magic_5.OUT Q6.t28 a_5036_n3150# VSS.t1274 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1998 VSS p2_gen_magic_0.xnor_magic_6.OUT a_14756_n3644# VSS.t452 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1999 VDD p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t6 VDD.t1803 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2000 a_34156_n889# mux_magic_0.OR_magic_0.A VDD.t825 VDD.t46 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2001 VSS Q2.t28 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT VSS.t1420 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2002 7b_counter_0.MDFF_1.tspc2_magic_0.Q 7b_counter_0.MDFF_1.QB.t10 VSS.t61 VSS.t60 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2003 VDD 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A a_26038_4932# VDD.t383 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2004 a_1559_n5540# p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_3.OUT.t1 VDD.t407 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2005 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t21 VDD.t2400 VDD.t2399 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2006 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_3.CLK.t20 divide_by_2_0.tg_magic_3.IN.t9 VSS.t1050 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2007 VDD DFF_magic_0.D.t34 a_27567_8496.t4 VDD.t2127 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2008 LD a_27567_8496.t17 VDD.t1186 VDD.t1181 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2009 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT Q4.t28 VDD.t1685 VDD.t1684 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2010 VSS CLK.t114 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t0 VSS.t560 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2011 a_1409_6275# 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A a_1209_6275# VSS.t1001 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2012 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A a_15865_6276# VSS.t1279 VSS.t1278 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X2013 VDD Q1.t30 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT VDD.t2094 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2014 a_8643_n6471# p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT VSS.t517 VSS.t516 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2015 a_34156_n889# mux_magic_0.OR_magic_0.A VDD.t824 VDD.t821 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2016 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A LD.t77 VDD.t1921 VDD.t1920 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2017 a_12931_1059# 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A a_12387_552# VSS.t1383 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2018 VDD a_1209_8579# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B VDD.t319 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2019 p3_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_1.B.t11 a_1541_n8095# VDD.t369 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2020 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A LD.t78 VDD.t1922 VDD.t1918 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2021 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_3.OUT VSS.t420 VSS.t419 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2022 VDD 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_5185_6275# VDD.t554 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2023 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t77 VDD.t1288 VDD.t1286 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2024 a_1209_4557# 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A VDD.t135 VDD.t134 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2025 a_5054_n1526# Q2.t29 VDD.t2438 VDD.t296 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2026 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_12387_6963# VDD.t711 VDD.t710 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2027 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT DFF_magic_0.tg_magic_3.CLK.t22 VDD.t2035 VDD.t2034 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2028 a_6725_5900# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A VDD.t535 VDD.t534 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2029 VDD D2_7.t21 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT VDD.t1978 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2030 VDD CLK.t115 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD.t2668 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2031 a_19152_1223# 7b_counter_0.MDFF_1.tspc2_magic_0.CLK VDD.t956 VDD.t955 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2032 VSS 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t11 a_4651_9163# VSS.t1529 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2033 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t78 VDD.t1290 VDD.t1289 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2034 VDD p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT a_5036_n4081# VDD.t262 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2035 OR_magic_1.VOUT a_30365_3514# VSS.t515 VSS.t514 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X2036 a_24003_10051# 7b_counter_0.3_inp_AND_magic_0.VOUT VSS.t415 VSS.t414 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2037 VDD 7b_counter_0.MDFF_5.LD.t79 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A VDD.t1261 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2038 VDD 7b_counter_0.MDFF_5.LD.t80 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A VDD.t1245 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2039 VSS 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_26126_3480# VSS.t406 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2040 a_1409_7469# LD.t79 a_1209_7469# VSS.t1062 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2041 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT Q5.t29 VDD.t256 VDD.t255 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2042 VDD DFF_magic_0.tg_magic_3.CLK.t23 DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD.t2036 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2043 a_16065_8580# CLK.t116 VSS.t559 VSS.t558 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2044 a_12387_5769# 7b_counter_0.MDFF_5.QB.t8 VDD.t931 VDD.t930 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2045 divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT OR_magic_1.VOUT.t25 VSS.t1491 VSS.t1490 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2046 DFF_magic_0.tg_magic_0.IN DFF_magic_0.tg_magic_1.IN.t17 VDD.t63 VDD.t62 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2047 VSS D2_5.t21 a_5385_2253# VSS.t1550 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2048 a_17405_5901# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A VDD.t2208 VDD.t627 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2049 a_1541_n8579# p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT VDD.t843 VDD.t842 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2050 VDD p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t22 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD.t2401 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2051 VDD a_1209_3363# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B VDD.t288 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2052 a_13353_n6613# p3_gen_magic_0.3_inp_AND_magic_0.A a_13553_n6613# VSS.t471 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2053 VDD D2_6.t23 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT VDD.t1349 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2054 VSS mux_magic_0.IN1.t15 a_32816_n1264# VSS.t1375 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2055 a_15865_4557# Q2.t30 VDD.t2440 VDD.t2439 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2056 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t10 VDD.t2377 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2057 VSS 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A a_17405_2092# VSS.t94 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2058 VSS D2_4.t24 a_23802_2253# VSS.t1330 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2059 VSS 7b_counter_0.MDFF_4.LD.t122 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A VSS.t967 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2060 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A a_5185_6275# VDD.t186 VDD.t185 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2061 VDD a_12387_552# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A VDD.t643 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2062 a_4235_9163# 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t12 a_4496_10093# VDD.t2011 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2063 p3_gen_magic_0.3_inp_AND_magic_0.VOUT a_13353_n6613# VSS.t702 VSS.t470 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2064 VDD a_5185_7469# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B VDD.t1700 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2065 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A a_1209_6275# VDD.t1709 VDD.t1708 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2066 a_6725_7308# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B a_6725_5900# VDD.t531 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2067 p3_gen_magic_0.xnor_magic_0.OUT Q1.t31 a_8643_n6471# VSS.t1211 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2068 VDD a_32616_n2458# mux_magic_0.OR_magic_0.B VDD.t695 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2069 a_5385_1059# 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A a_5185_1059# VSS.t298 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2070 a_16065_9774# CLK.t117 VSS.t557 VSS.t556 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2071 VDD a_19152_6440# 7b_counter_0.MDFF_6.QB.t0 VDD.t492 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2072 a_2749_7308# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B a_2749_5900# VDD.t1039 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2073 a_8939_n7648# p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_6.OUT VSS.t163 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2074 VDD 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A a_26038_684# VDD.t1065 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2075 a_11191_5901# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_11279_6341# VDD.t357 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2076 a_19152_739# 7b_counter_0.MDFF_1.tspc2_magic_0.D VDD.t1019 VDD.t1018 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2077 VDD D2_6.t24 a_12387_1746# VDD.t1352 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2078 VSS p3_gen_magic_0.P3.t15 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN VSS.t896 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2079 divide_by_2_0.tg_magic_2.IN divide_by_2_0.tg_magic_3.CLK.t21 divide_by_2_0.tg_magic_3.IN.t12 VSS.t1051 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2080 VDD P2.t15 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN VDD.t2228 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2081 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A LD.t80 VDD.t1923 VDD.t1881 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2082 VSS mux_magic_0.IN2.t14 a_32816_n2458# VSS.t1250 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2083 a_27234_1746# CLK.t118 VDD.t2667 VDD.t2666 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2084 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A a_1209_1059# VSS.t79 VSS.t78 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X2085 a_5515_3947# 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t11 7b_counter_0.MDFF_0.QB.t0 VSS.t1439 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2086 a_23258_1746# D2_4.t25 VDD.t2283 VDD.t2282 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2087 VSS CLK.t119 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VSS.t553 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2088 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t123 VDD.t1634 VDD.t1633 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2089 VDD a_15865_8580# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B VDD.t393 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2090 p3_gen_magic_0.xnor_magic_0.OUT D2_2.t25 a_8643_n6024# VDD.t981 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2091 VSS Q6.t29 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT VSS.t1275 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2092 a_11191_4932# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B a_11279_3480# VDD.t517 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2093 VDD 7b_counter_0.MDFF_5.LD.t81 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A VDD.t1272 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2094 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT VDD.t1085 VDD.t1084 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2095 VDD Q7.t22 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT VDD.t1397 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2096 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A LD.t81 VSS.t1096 VSS.t1095 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2097 a_8643_n5540# p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_0.OUT VDD.t980 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2098 a_1409_9773# 7b_counter_0.MDFF_3.QB VSS.t318 VSS.t317 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2099 VDD a_5185_2253# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B VDD.t1642 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2100 VDD 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A a_17405_4932# VDD.t156 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2101 a_13553_n6613# p3_gen_magic_0.3_inp_AND_magic_0.A a_13353_n6613# VSS.t471 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2102 a_15865_6276# 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A a_16065_6276# VSS.t170 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2103 VDD OR_magic_2.VOUT.t24 divide_by_2_0.tg_magic_3.CLK.t3 VDD.t753 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2104 VSS 7b_counter_0.DFF_magic_0.Q.t21 DFF_magic_0.D VSS.t1212 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2105 VDD.t1053 VDD.t1051 VDD.t1053 VDD.t1052 pfet_03v3 ad=0.493p pd=3.12u as=0 ps=0 w=1.12u l=0.56u
X2106 VDD D2_7.t22 a_1209_8579# VDD.t1981 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2107 VDD a_16186_n3644# p2_gen_magic_0.3_inp_AND_magic_0.C.t1 VDD.t215 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2108 divide_by_2_1.tg_magic_2.IN divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.IN.t0 VDD.t97 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2109 divide_by_2_1.tg_magic_0.IN OR_magic_1.VOUT.t26 divide_by_2_1.tg_magic_3.OUT VSS.t1492 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2110 a_30365_3514# P2.t16 VSS.t1289 VSS.t1288 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2111 VDD CLK.t120 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD.t2663 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2112 VDD CLK.t121 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD.t2671 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2113 p2_gen_magic_0.xnor_magic_6.OUT D2_6.t25 a_8523_n3597# VDD.t861 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2114 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT VDD.t2376 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2115 a_13553_n6613# p3_gen_magic_0.3_inp_AND_magic_0.A a_13353_n6613# VSS.t470 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2116 VDD 7b_counter_0.MDFF_5.QB.t9 7b_counter_0.MDFF_5.tspc2_magic_0.Q VDD.t927 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X2117 a_4496_4393# 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t12 VDD.t2454 VDD.t873 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2118 VSS D2_7.t23 a_1409_8579# VSS.t598 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2119 VDD Q3.t31 a_1559_n6024# VDD.t580 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2120 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q7.t23 VDD.t1401 VDD.t1400 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2121 VDD 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A a_7215_10149# VDD.t507 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2122 a_9212_5956# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t12 a_9412_5956# VDD.t913 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2123 a_4496_9609# a_4235_9163# a_4651_9163# VSS.t185 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2124 VDD p3_gen_magic_0.3_inp_AND_magic_0.C.t7 a_13353_n6613# VDD.t1987 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2125 VDD a_4496_9609# 7b_counter_0.MDFF_3.QB VDD.t414 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2126 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t124 VSS.t970 VSS.t907 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2127 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT D2_5.t22 VDD.t2742 VDD.t2741 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2128 divide_by_2_0.tg_magic_0.IN divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.OUT VDD.t952 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2129 VSS D2_5.t23 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT VSS.t1534 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2130 a_20041_8580# 7b_counter_0.MDFF_5.LD.t82 a_19841_8580# VSS.t790 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2131 VDD CLK.t122 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK VDD.t2682 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2132 VSS 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A a_17405_7309# VSS.t537 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2133 a_16386_n3644# p2_gen_magic_0.xnor_magic_5.OUT a_16186_n3644# VSS.t118 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2134 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT VDD.t1802 VDD.t1801 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2135 OR_magic_1.VOUT a_30365_3514# VDD.t978 VDD.t977 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X2136 a_16065_8580# 7b_counter_0.MDFF_5.LD.t83 a_15865_8580# VSS.t785 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2137 VDD mux_magic_0.OR_magic_0.A a_34156_n889# VDD.t821 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2138 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t23 VSS.t1400 VSS.t1399 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2139 VSS a_19152_1223# a_20171_1669# VSS.t64 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2140 VDD Q7.t24 a_1541_n8095# VDD.t844 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2141 a_26038_4932# 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_26126_3480# VDD.t386 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2142 VSS 7b_counter_0.MDFF_5.QB.t10 7b_counter_0.MDFF_5.tspc2_magic_0.Q VSS.t489 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2143 VDD D2_5.t24 a_1209_3363# VDD.t2743 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2144 a_8411_9730# 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A VDD.t374 VDD.t373 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2145 a_19841_4557# 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A VDD.t1717 VDD.t1716 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2146 divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.CLK.t20 VDD.t2009 VDD.t2008 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2147 a_15865_4557# 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A VDD.t302 VDD.t301 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2148 a_5054_n1526# D2_3.t25 p2_gen_magic_0.xnor_magic_4.OUT VDD.t769 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2149 VDD p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8643_n5540# VDD.t987 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2150 a_5185_6275# 7b_counter_0.MDFF_3.tspc2_magic_0.Q VDD.t553 VDD.t552 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2151 VSS DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_1.IN.t0 VSS.t541 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2152 a_20041_9774# 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A a_19841_9774# VSS.t142 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2153 VDD D2_7.t24 a_5185_7469# VDD.t1984 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2154 divide_by_2_0.tg_magic_3.CLK OR_magic_2.VOUT.t25 VDD.t757 VDD.t756 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2155 VSS LD.t82 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A VSS.t1083 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2156 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A LD.t83 VDD.t1924 VDD.t1920 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2157 a_16065_9774# 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A a_15865_9774# VSS.t266 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2158 VSS Q2.t31 7b_counter_0.3_inp_AND_magic_0.C VSS.t1423 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2159 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK.t123 VDD.t2681 VDD.t2680 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2160 VSS 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A a_2749_7308# VSS.t215 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2161 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q7.t25 VSS.t859 VSS.t858 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2162 a_5036_n3597# D2_7.t25 p2_gen_magic_0.xnor_magic_5.OUT VDD.t398 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2163 a_23352_n6798# p3_gen_magic_0.P3.t16 a_23352_n5390# VDD.t1475 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2164 VSS a_8713_1625# a_8825_1669# VSS.t240 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2165 a_6725_684# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A VDD.t1692 VDD.t1691 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2166 VDD a_12387_1746# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B VDD.t409 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2167 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A LD.t84 VDD.t1925 VDD.t1857 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2168 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t84 VDD.t1297 VDD.t1198 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2169 a_11191_684# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_11279_1124# VDD.t448 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2170 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A LD.t85 VDD.t1926 VDD.t1912 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2171 a_1209_1059# 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A a_1409_1059# VSS.t425 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2172 VDD 7b_counter_0.MDFF_4.LD.t125 a_8411_3319# VDD.t1635 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2173 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t85 VDD.t1298 VDD.t1205 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2174 VSS CLK.t124 a_16065_8580# VSS.t550 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2175 a_11191_4932# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B a_11279_3480# VDD.t1143 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2176 a_7303_3480# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B a_7215_4932# VDD.t526 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2177 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t86 VDD.t1299 VDD.t1289 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2178 VSS D2_1.t35 a_1957_n3150# VSS.t818 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2179 divide_by_2_0.tg_magic_3.IN OR_magic_2.VOUT.t26 divide_by_2_0.tg_magic_1.IN.t2 VSS.t397 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2180 a_11292_n2115# p2_gen_magic_0.xnor_magic_4.OUT VDD.t772 VDD.t771 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2181 VSS divide_by_2_0.tg_magic_3.CLK.t22 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT VSS.t1052 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X2182 VDD CLK.t125 a_15865_8580# VDD.t2677 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2183 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK.t126 VSS.t547 VSS.t546 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2184 a_1409_2253# LD.t86 a_1209_2253# VSS.t1066 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2185 a_1975_n1973# p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_3.OUT.t1 VSS.t311 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2186 VDD 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A a_15865_4557# VDD.t298 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2187 VDD CLK.t127 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t2 VDD.t2674 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2188 VDD D2_5.t25 a_5185_2253# VDD.t2746 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2189 a_14556_n3644# p2_gen_magic_0.AND2_magic_1.A VDD.t1786 VDD.t1785 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2190 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT Q4.t29 VSS.t993 VSS.t992 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X2191 VDD 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A a_15865_1059# VDD.t588 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2192 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A a_1209_1059# VDD.t120 VDD.t119 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2193 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B a_5185_7469# VDD.t1699 VDD.t1698 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X2194 7b_counter_0.MDFF_0.tspc2_magic_0.D a_2749_3524# VDD.t183 VDD.t182 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
R0 VDD.t2371 VDD.t2617 2420.69
R1 VDD.t2325 VDD.t955 1683.52
R2 VDD.t1023 VDD.t2217 1646.52
R3 VDD.t1371 VDD.t1684 1275.86
R4 VDD.t1349 VDD.t1670 1275.86
R5 VDD.t421 VDD.t1429 1199.13
R6 VDD.t927 VDD.t102 1198.41
R7 VDD.t1440 VDD.t621 1198.41
R8 VDD.t139 VDD.t425 1194.81
R9 VDD.t2092 VDD.t2492 1168.97
R10 VDD.t2477 VDD.t2076 1168.97
R11 VDD.t2730 VDD.t1785 1105.34
R12 VDD.t1416 VDD.t2719 1105.34
R13 VDD.t1055 VDD.t2097 1070.89
R14 VDD.t1334 VDD.t1721 1061.39
R15 VDD.t766 VDD.t763 1049.07
R16 VDD.t905 VDD.t902 1049.07
R17 VDD.t803 VDD.t2529 1046.14
R18 VDD.t829 VDD.t746 1046.14
R19 VDD.t1155 VDD.t1086 1046.14
R20 VDD.t1806 VDD.t2590 1046.14
R21 VDD.t2641 VDD.t1041 1046.14
R22 VDD.t126 VDD.t2523 1046.14
R23 VDD.t449 VDD.n1353 1034.06
R24 VDD.t680 VDD.t210 1007.33
R25 VDD.t1792 VDD.t104 1007.33
R26 VDD.n1353 VDD.t1769 1007.16
R27 VDD.t2274 VDD.t2409 1006.9
R28 VDD.t2166 VDD.t1319 1006.9
R29 VDD.t2264 VDD.t2428 1006.9
R30 VDD.t2455 VDD.t2191 1006.9
R31 VDD.t1973 VDD.t244 993.104
R32 VDD.t229 VDD.t1963 993.104
R33 VDD.t446 VDD.t507 958.63
R34 VDD.t1700 VDD.t534 958.63
R35 VDD.t334 VDD.t197 957.376
R36 VDD.t710 VDD.t360 957.376
R37 VDD.t1079 VDD.t390 957.376
R38 VDD.t1127 VDD.t2209 957.376
R39 VDD.t319 VDD.t692 957.376
R40 VDD.t288 VDD.t676 957.376
R41 VDD.t1691 VDD.t1642 957.376
R42 VDD.t342 VDD.t412 957.376
R43 VDD.n1364 VDD.t1601 921.26
R44 VDD.n1364 VDD.t1514 921.26
R45 VDD.t949 VDD.t1887 911.077
R46 VDD.t2246 VDD.t2163 900.633
R47 VDD.t1261 VDD.t165 864.109
R48 VDD.t1144 VDD.t1482 864.109
R49 VDD.t1064 VDD.t1489 864.109
R50 VDD.t1198 VDD.t575 864.109
R51 VDD.t371 VDD.t1891 864.109
R52 VDD.t720 VDD.t1567 864.109
R53 VDD.t962 VDD.t92 861.423
R54 VDD.t957 VDD.t83 842.491
R55 VDD.t1584 VDD.t591 842.491
R56 VDD.t1476 VDD.t2379 842.491
R57 VDD.n1277 VDD.t947 841.558
R58 VDD.t886 VDD.t549 806.37
R59 VDD.t775 VDD.t1467 806.37
R60 VDD.t202 VDD.t628 806.37
R61 VDD.t1448 VDD.t68 806.37
R62 VDD.t873 VDD.t181 806.37
R63 VDD.t2005 VDD.t2364 787.708
R64 VDD.t2340 VDD.t2036 787.708
R65 VDD.t2692 VDD.t608 787.708
R66 VDD.t2039 VDD.t2104 787.708
R67 VDD.t895 VDD.t10 787.708
R68 VDD.t1811 VDD.t2146 787.708
R69 VDD.t1463 VDD.t2663 787.708
R70 VDD.t36 VDD.t663 787.708
R71 VDD.t2401 VDD.t2220 787.708
R72 VDD.t2378 VDD.t2374 787.708
R73 VDD.t2202 VDD.t1006 787.708
R74 VDD.t438 VDD.t117 787.708
R75 VDD.t2498 VDD.t1135 782.313
R76 VDD.t97 VDD.t2008 782.313
R77 VDD.t761 VDD.t2601 782.313
R78 VDD.t1001 VDD.t2704 782.313
R79 VDD.t366 VDD.t2042 782.313
R80 VDD.t2690 VDD.t2563 782.313
R81 VDD.t2550 VDD.t795 782.313
R82 VDD.t331 VDD.t2032 782.313
R83 VDD.t563 VDD.t1828 782.313
R84 VDD.t896 VDD.t740 782.313
R85 VDD.t738 VDD.t952 782.313
R86 VDD.t999 VDD.t1826 782.313
R87 VDD.t1028 VDD.t2545 782.313
R88 VDD.t1742 VDD.t1153 782.313
R89 VDD.t2531 VDD.t1715 782.313
R90 VDD.t664 VDD.t1168 782.313
R91 VDD.t2599 VDD.t1799 782.313
R92 VDD.t286 VDD.t2384 782.313
R93 VDD.t316 VDD.t2390 782.313
R94 VDD.t2377 VDD.t2626 782.313
R95 VDD.t939 VDD.t2701 782.313
R96 VDD.t2539 VDD.t2200 782.313
R97 VDD.t1766 VDD.t1993 782.313
R98 VDD.t436 VDD.t2507 782.313
R99 VDD.n862 VDD.t792 776.163
R100 VDD.t1205 VDD.t1258 757.283
R101 VDD.n2425 VDD.t1445 757.01
R102 VDD.n1312 VDD.t100 757.01
R103 VDD.n546 VDD.t2327 755.245
R104 VDD.n1070 VDD.t879 755.245
R105 VDD.n782 VDD.t777 755.245
R106 VDD.n1023 VDD.t631 755.245
R107 VDD.n2416 VDD.t71 755.245
R108 VDD.n1256 VDD.t182 755.245
R109 VDD.n1166 VDD.t1030 755.245
R110 VDD.n245 VDD.t1772 755.245
R111 VDD.t2579 VDD.t2027 746.33
R112 VDD.t2682 VDD.t2537 746.33
R113 VDD.t2566 VDD.t2399 746.33
R114 VDD.t2034 VDD.t2606 746.33
R115 VDD.t753 VDD.t1814 741.497
R116 VDD.t2500 VDD.t2000 741.497
R117 VDD.n1045 VDD.n1040 720.605
R118 VDD.t2520 VDD.t480 713.571
R119 VDD.t62 VDD.t2655 713.571
R120 VDD.t2668 VDD.t916 713.571
R121 VDD.t730 VDD.t1410 713.571
R122 VDD.t2236 VDD.t1157 713.571
R123 VDD.t2585 VDD.t2749 713.571
R124 VDD.t368 VDD.t799 699.505
R125 VDD.t562 VDD.t832 699.505
R126 VDD.t1713 VDD.t1084 699.505
R127 VDD.t318 VDD.t1801 699.505
R128 VDD.t1044 VDD.t940 699.505
R129 VDD.t1768 VDD.t132 699.505
R130 VDD.t2094 VDD.t1731 684.721
R131 VDD.t293 VDD.t2411 684.721
R132 VDD.t2299 VDD.t603 684.721
R133 VDD.t808 VDD.t1397 684.721
R134 VDD.t262 VDD.t2173 684.721
R135 VDD.t246 VDD.t249 684.721
R136 VDD.t1677 VDD.t666 684.721
R137 VDD.t2306 VDD.t580 684.721
R138 VDD.t2080 VDD.t987 684.721
R139 VDD.t2430 VDD.t75 684.721
R140 VDD.t1386 VDD.t844 684.721
R141 VDD.t1728 VDD.t2195 684.721
R142 VDD.t231 VDD.t237 684.721
R143 VDD.t633 VDD.t1656 684.721
R144 VDD.t1918 VDD.t1703 669.359
R145 VDD.t1914 VDD.t638 669.359
R146 VDD.t375 VDD.t1241 669.359
R147 VDD.t1104 VDD.t1251 669.359
R148 VDD.t1437 VDD.t1497 669.359
R149 VDD.t600 VDD.t1519 669.359
R150 VDD.t557 VDD.t1236 669.359
R151 VDD.t303 VDD.t1542 669.359
R152 VDD.t1575 VDD.t585 669.359
R153 VDD.t1763 VDD.t1561 669.359
R154 VDD.t1229 VDD.t327 669.359
R155 VDD.t257 VDD.t1210 669.359
R156 VDD.t497 VDD.t1224 669.359
R157 VDD.t782 VDD.t1857 669.359
R158 VDD.t134 VDD.t1912 669.359
R159 VDD.t1837 VDD.t573 669.359
R160 VDD.t1920 VDD.t814 669.359
R161 VDD.t1485 VDD.t1716 669.359
R162 VDD.t1487 VDD.t301 669.359
R163 VDD.t1300 VDD.t992 669.359
R164 VDD.t1945 VDD.t458 634.721
R165 VDD.t769 VDD.t2483 634.721
R166 VDD.t2272 VDD.t2045 634.721
R167 VDD.t1332 VDD.t1149 634.721
R168 VDD.t1971 VDD.t398 634.721
R169 VDD.t862 VDD.t1374 634.721
R170 VDD.t442 VDD.t2726 634.721
R171 VDD.t980 VDD.t1933 634.721
R172 VDD.t400 VDD.t2471 634.721
R173 VDD.t407 VDD.t2262 634.721
R174 VDD.t2458 VDD.t370 634.721
R175 VDD.t759 VDD.t1961 634.721
R176 VDD.t1362 VDD.t64 634.721
R177 VDD.t1415 VDD.t2741 634.721
R178 VDD.n862 VDD.t1055 625
R179 VDD.t1693 VDD.t1688 621.245
R180 VDD.t187 VDD.t537 621.072
R181 VDD.t378 VDD.t513 621.072
R182 VDD.t1710 VDD.t427 613.875
R183 VDD.n1365 VDD.n1364 611.722
R184 VDD.n1364 VDD.n1363 611.722
R185 VDD.n545 VDD.t2325 606.742
R186 VDD.t2064 VDD.t1383 581.967
R187 VDD.t1189 VDD.t2125 572.513
R188 VDD.t1545 VDD.t1517 566.929
R189 VDD.t1601 VDD.t1545 566.929
R190 VDD.t1514 VDD.t1589 566.929
R191 VDD.t1589 VDD.t1537 566.929
R192 VDD.t425 VDD.t1039 561.039
R193 VDD.n1599 VDD.t99 549.321
R194 VDD.n1707 VDD.t1002 549.321
R195 VDD.n611 VDD.t329 549.321
R196 VDD.n1828 VDD.t997 549.321
R197 VDD.n1910 VDD.t1029 549.321
R198 VDD.n1737 VDD.t287 549.321
R199 VDD.n1354 VDD.t1769 534.769
R200 VDD.t2290 VDD.t1661 519.126
R201 VDD.t507 VDD.t1442 504.673
R202 VDD.t534 VDD.t531 504.673
R203 VDD.t197 VDD.t2216 503.497
R204 VDD.t360 VDD.t551 503.497
R205 VDD.t390 VDD.t774 503.497
R206 VDD.t2209 VDD.t629 503.497
R207 VDD.t692 VDD.t67 503.497
R208 VDD.t676 VDD.t179 503.497
R209 VDD.t422 VDD.t1691 503.497
R210 VDD.t451 VDD.t342 503.497
R211 VDD.t484 VDD.n1599 491.791
R212 VDD.t59 VDD.n1707 491.791
R213 VDD.t921 VDD.n611 491.791
R214 VDD.t1407 VDD.n1828 491.791
R215 VDD.t2238 VDD.n1910 491.791
R216 VDD.t1421 VDD.n1737 491.791
R217 VDD.t1176 VDD.n22 423.697
R218 VDD.t1171 VDD.n481 421.245
R219 VDD.t568 VDD.n2443 421.245
R220 VDD.n2443 VDD.t1013 421.245
R221 VDD.n2459 VDD.t1121 421.245
R222 VDD.n322 VDD.t1138 421.245
R223 VDD.n322 VDD.t1066 421.245
R224 VDD.n1337 VDD.t964 421.245
R225 VDD.n1337 VDD.t337 421.245
R226 VDD.n736 VDD.t464 421.245
R227 VDD.n769 VDD.t469 421.245
R228 VDD.n769 VDD.t985 421.245
R229 VDD.n736 VDD.t544 421.245
R230 VDD.n2455 VDD.t393 421.245
R231 VDD.n2459 VDD.t166 421.245
R232 VDD.n2455 VDD.t502 421.245
R233 VDD.t1744 VDD.n1203 421.245
R234 VDD.n1203 VDD.t121 421.245
R235 VDD.t433 VDD.n572 421.245
R236 VDD.n572 VDD.t655 421.245
R237 VDD.n481 VDD.t151 421.245
R238 VDD.n1679 VDD.t944 421.245
R239 VDD.t695 VDD.n1679 421.245
R240 VDD.n519 VDD.t199 413.92
R241 VDD.n1356 VDD.t345 413.92
R242 VDD.n521 VDD.n519 406.594
R243 VDD.n1357 VDD.n1356 406.594
R244 VDD.t94 VDD.t87 404.495
R245 VDD.t92 VDD.t94 404.495
R246 VDD.t1025 VDD.t962 404.495
R247 VDD.t958 VDD.t1025 404.495
R248 VDD.t2218 VDD.t195 404.495
R249 VDD.t787 VDD.t2050 402.986
R250 VDD.t2050 VDD.t2102 402.986
R251 VDD.n1061 VDD.n1060 402.747
R252 VDD.n668 VDD.n667 402.747
R253 VDD.n1021 VDD.n1020 402.747
R254 VDD.n2414 VDD.n2413 402.747
R255 VDD.n1254 VDD.n1253 402.747
R256 VDD.t1174 VDD.t1171 395.604
R257 VDD.t2576 VDD.t1174 395.604
R258 VDD.t2624 VDD.t1614 395.604
R259 VDD.t1614 VDD.t1612 395.604
R260 VDD.t332 VDD.t334 395.604
R261 VDD.t2465 VDD.t332 395.604
R262 VDD.t2475 VDD.t1578 395.604
R263 VDD.t1578 VDD.t1571 395.604
R264 VDD.t1708 VDD.t1710 395.604
R265 VDD.t2185 VDD.t1708 395.604
R266 VDD.t1705 VDD.t2189 395.604
R267 VDD.t1703 VDD.t1705 395.604
R268 VDD.t142 VDD.t139 395.604
R269 VDD.t2634 VDD.t142 395.604
R270 VDD.t2639 VDD.t1839 395.604
R271 VDD.t1839 VDD.t1889 395.604
R272 VDD.t185 VDD.t187 395.604
R273 VDD.t554 VDD.t185 395.604
R274 VDD.t640 VDD.t552 395.604
R275 VDD.t638 VDD.t640 395.604
R276 VDD.t1277 VDD.t1221 395.604
R277 VDD.t2658 VDD.t1277 395.604
R278 VDD.t2597 VDD.t565 395.604
R279 VDD.t565 VDD.t568 395.604
R280 VDD.t373 VDD.t375 395.604
R281 VDD.t702 VDD.t373 395.604
R282 VDD.t700 VDD.t380 395.604
R283 VDD.t380 VDD.t378 395.604
R284 VDD.t1102 VDD.t1104 395.604
R285 VDD.t2066 VDD.t1102 395.604
R286 VDD.t1015 VDD.t2088 395.604
R287 VDD.t1013 VDD.t1015 395.604
R288 VDD.t1124 VDD.t1121 395.604
R289 VDD.t1313 VDD.t1124 395.604
R290 VDD.t1328 VDD.t1233 395.604
R291 VDD.t1233 VDD.t1212 395.604
R292 VDD.t1435 VDD.t1437 395.604
R293 VDD.t234 VDD.t1435 395.604
R294 VDD.t225 VDD.t1140 395.604
R295 VDD.t1140 VDD.t1138 395.604
R296 VDD.t1505 VDD.t1617 395.604
R297 VDD.t2542 VDD.t1505 395.604
R298 VDD.t1068 VDD.t2650 395.604
R299 VDD.t1066 VDD.t1068 395.604
R300 VDD.t598 VDD.t600 395.604
R301 VDD.t311 VDD.t598 395.604
R302 VDD.t966 VDD.t314 395.604
R303 VDD.t964 VDD.t966 395.604
R304 VDD.t1492 VDD.t1635 395.604
R305 VDD.t1366 VDD.t1492 395.604
R306 VDD.t339 VDD.t1364 395.604
R307 VDD.t337 VDD.t339 395.604
R308 VDD.t1231 VDD.t1207 395.604
R309 VDD.t1942 VDD.t1231 395.604
R310 VDD.t1935 VDD.t712 395.604
R311 VDD.t712 VDD.t710 395.604
R312 VDD.t560 VDD.t924 395.604
R313 VDD.t404 VDD.t930 395.604
R314 VDD.t1631 VDD.t1598 395.604
R315 VDD.t2652 VDD.t1631 395.604
R316 VDD.t2666 VDD.t466 395.604
R317 VDD.t466 VDD.t464 395.604
R318 VDD.t1605 VDD.t1551 395.604
R319 VDD.t2267 VDD.t1605 395.604
R320 VDD.t471 VDD.t2282 395.604
R321 VDD.t469 VDD.t471 395.604
R322 VDD.t306 VDD.t303 395.604
R323 VDD.t725 VDD.t306 395.604
R324 VDD.t982 VDD.t723 395.604
R325 VDD.t985 VDD.t982 395.604
R326 VDD.t585 VDD.t583 395.604
R327 VDD.t583 VDD.t2310 395.604
R328 VDD.t541 VDD.t2297 395.604
R329 VDD.t544 VDD.t541 395.604
R330 VDD.t0 VDD.t1761 395.604
R331 VDD.t660 VDD.t3 395.604
R332 VDD.t1509 VDD.t1620 395.604
R333 VDD.t2257 VDD.t1509 395.604
R334 VDD.t2260 VDD.t1081 395.604
R335 VDD.t1081 VDD.t1079 395.604
R336 VDD.t1130 VDD.t1127 395.604
R337 VDD.t1336 VDD.t1130 395.604
R338 VDD.t1304 VDD.t1202 395.604
R339 VDD.t1202 VDD.t1200 395.604
R340 VDD.t2206 VDD.t2248 395.604
R341 VDD.t2251 VDD.t324 395.604
R342 VDD.t396 VDD.t393 395.604
R343 VDD.t2677 VDD.t396 395.604
R344 VDD.t2555 VDD.t1216 395.604
R345 VDD.t1216 VDD.t1214 395.604
R346 VDD.t166 VDD.t169 395.604
R347 VDD.t169 VDD.t274 395.604
R348 VDD.t272 VDD.t259 395.604
R349 VDD.t259 VDD.t257 395.604
R350 VDD.t502 VDD.t505 395.604
R351 VDD.t505 VDD.t2594 395.604
R352 VDD.t2611 VDD.t499 395.604
R353 VDD.t499 VDD.t497 395.604
R354 VDD.t1275 VDD.t1266 395.604
R355 VDD.t1949 VDD.t1275 395.604
R356 VDD.t1947 VDD.t443 395.604
R357 VDD.t443 VDD.t446 395.604
R358 VDD.t322 VDD.t319 395.604
R359 VDD.t1981 VDD.t322 395.604
R360 VDD.t1957 VDD.t1870 395.604
R361 VDD.t1870 VDD.t1902 395.604
R362 VDD.t683 VDD.t618 395.604
R363 VDD.t624 VDD.t784 395.604
R364 VDD.t1698 VDD.t1700 395.604
R365 VDD.t1984 VDD.t1698 395.604
R366 VDD.t1959 VDD.t1873 395.604
R367 VDD.t1873 VDD.t1906 395.604
R368 VDD.t291 VDD.t288 395.604
R369 VDD.t2743 VDD.t291 395.604
R370 VDD.t2722 VDD.t1876 395.604
R371 VDD.t1876 VDD.t1904 395.604
R372 VDD.t705 VDD.t2443 395.604
R373 VDD.t2446 VDD.t136 395.604
R374 VDD.t1747 VDD.t1744 395.604
R375 VDD.t2631 VDD.t1747 395.604
R376 VDD.t2648 VDD.t1842 395.604
R377 VDD.t1842 VDD.t1893 395.604
R378 VDD.t1688 VDD.t1686 395.604
R379 VDD.t1686 VDD.t837 395.604
R380 VDD.t570 VDD.t840 395.604
R381 VDD.t573 VDD.t570 395.604
R382 VDD.t121 VDD.t119 395.604
R383 VDD.t119 VDD.t1647 395.604
R384 VDD.t811 VDD.t1682 395.604
R385 VDD.t814 VDD.t811 395.604
R386 VDD.t1642 VDD.t1645 395.604
R387 VDD.t1645 VDD.t2746 395.604
R388 VDD.t2724 VDD.t1883 395.604
R389 VDD.t1883 VDD.t1908 395.604
R390 VDD.t1624 VDD.t1586 395.604
R391 VDD.t1352 VDD.t1624 395.604
R392 VDD.t409 VDD.t1355 395.604
R393 VDD.t412 VDD.t409 395.604
R394 VDD.t961 VDD.t957 395.604
R395 VDD.t1018 VDD.t963 395.604
R396 VDD.t1020 VDD.t1018 395.604
R397 VDD.t2217 VDD.t2215 395.604
R398 VDD.t199 VDD.t193 395.604
R399 VDD.t89 VDD.t593 395.604
R400 VDD.t588 VDD.t85 395.604
R401 VDD.t2382 VDD.t1432 395.604
R402 VDD.t2018 VDD.t643 395.604
R403 VDD.t345 VDD.t347 395.604
R404 VDD.t448 VDD.t449 395.604
R405 VDD.t431 VDD.t433 395.604
R406 VDD.t2480 VDD.t431 395.604
R407 VDD.t2487 VDD.t1626 395.604
R408 VDD.t1626 VDD.t1610 395.604
R409 VDD.t655 VDD.t653 395.604
R410 VDD.t653 VDD.t648 395.604
R411 VDD.t1718 VDD.t651 395.604
R412 VDD.t1716 VDD.t1718 395.604
R413 VDD.t151 VDD.t154 395.604
R414 VDD.t154 VDD.t2425 395.604
R415 VDD.t298 VDD.t2439 395.604
R416 VDD.t301 VDD.t298 395.604
R417 VDD.t218 VDD.t215 395.604
R418 VDD.t2406 VDD.t218 395.604
R419 VDD.t212 VDD.t2404 395.604
R420 VDD.t210 VDD.t212 395.604
R421 VDD.t678 VDD.t680 395.604
R422 VDD.t866 VDD.t678 395.604
R423 VDD.t1787 VDD.t869 395.604
R424 VDD.t1785 VDD.t1787 395.604
R425 VDD.t1721 VDD.t1724 395.604
R426 VDD.t1724 VDD.t49 395.604
R427 VDD.t106 VDD.t52 395.604
R428 VDD.t104 VDD.t106 395.604
R429 VDD.t1790 VDD.t1792 395.604
R430 VDD.t936 VDD.t1790 395.604
R431 VDD.t934 VDD.t1418 395.604
R432 VDD.t1418 VDD.t1416 395.604
R433 VDD.t944 VDD.t942 395.604
R434 VDD.t942 VDD.t2351 395.604
R435 VDD.t994 VDD.t2354 395.604
R436 VDD.t992 VDD.t994 395.604
R437 VDD.t698 VDD.t695 395.604
R438 VDD.t2151 VDD.t698 395.604
R439 VDD.t2144 VDD.t1325 395.604
R440 VDD.t1325 VDD.t1344 395.604
R441 VDD.t963 VDD.n505 390.111
R442 VDD.t1511 VDD.n1362 386.447
R443 VDD.n529 VDD.t1507 384.615
R444 VDD.n530 VDD.t1558 380.952
R445 VDD.t1633 VDD.n1361 380.952
R446 VDD.t482 VDD.t484 372.414
R447 VDD.t480 VDD.t477 372.414
R448 VDD.t2359 VDD.t2361 372.414
R449 VDD.t2364 VDD.t2356 372.414
R450 VDD.t54 VDD.t59 372.414
R451 VDD.t56 VDD.t62 372.414
R452 VDD.t2332 VDD.t2343 372.414
R453 VDD.t2334 VDD.t2340 372.414
R454 VDD.t1952 VDD.t1939 372.414
R455 VDD.t1930 VDD.t1945 372.414
R456 VDD.t2074 VDD.t2094 372.414
R457 VDD.t2083 VDD.t2092 372.414
R458 VDD.t2492 VDD.t2485 372.414
R459 VDD.t2483 VDD.t2468 372.414
R460 VDD.t2411 VDD.t2422 372.414
R461 VDD.t2409 VDD.t2433 372.414
R462 VDD.t2280 VDD.t2274 372.414
R463 VDD.t2254 VDD.t2272 372.414
R464 VDD.t2295 VDD.t2299 372.414
R465 VDD.t2287 VDD.t2293 372.414
R466 VDD.t2109 VDD.t2106 372.414
R467 VDD.t2097 VDD.t2047 372.414
R468 VDD.t2622 VDD.t2579 372.414
R469 VDD.t2674 VDD.t2637 372.414
R470 VDD.t613 VDD.t615 372.414
R471 VDD.t608 VDD.t610 372.414
R472 VDD.t914 VDD.t921 372.414
R473 VDD.t916 VDD.t918 372.414
R474 VDD.t2053 VDD.t2099 372.414
R475 VDD.t2104 VDD.t2055 372.414
R476 VDD.t1397 VDD.t1391 372.414
R477 VDD.t1393 VDD.t1400 372.414
R478 VDD.t2173 VDD.t2179 372.414
R479 VDD.t2182 VDD.t2166 372.414
R480 VDD.t1319 VDD.t1339 372.414
R481 VDD.t1316 VDD.t1332 372.414
R482 VDD.t255 VDD.t246 372.414
R483 VDD.t244 VDD.t222 372.414
R484 VDD.t1976 VDD.t1973 372.414
R485 VDD.t1966 VDD.t1971 372.414
R486 VDD.t1654 VDD.t1677 372.414
R487 VDD.t1684 VDD.t1666 372.414
R488 VDD.t1357 VDD.t1371 372.414
R489 VDD.t1374 VDD.t1359 372.414
R490 VDD.t2736 VDD.t2730 372.414
R491 VDD.t2726 VDD.t2738 372.414
R492 VDD.t12 VDD.t17 372.414
R493 VDD.t10 VDD.t14 372.414
R494 VDD.t1412 VDD.t1407 372.414
R495 VDD.t1410 VDD.t1404 372.414
R496 VDD.t2154 VDD.t2148 372.414
R497 VDD.t2146 VDD.t2156 372.414
R498 VDD.t1465 VDD.t1457 372.414
R499 VDD.t1460 VDD.t1463 372.414
R500 VDD.t2244 VDD.t2238 372.414
R501 VDD.t2241 VDD.t2236 372.414
R502 VDD.t2291 VDD.t2306 372.414
R503 VDD.t2303 VDD.t2313 372.414
R504 VDD.t1937 VDD.t1927 372.414
R505 VDD.t1933 VDD.t1954 372.414
R506 VDD.t2058 VDD.t2080 372.414
R507 VDD.t2076 VDD.t2070 372.414
R508 VDD.t2473 VDD.t2477 372.414
R509 VDD.t2471 VDD.t2489 372.414
R510 VDD.t2417 VDD.t2430 372.414
R511 VDD.t2428 VDD.t2419 372.414
R512 VDD.t2270 VDD.t2264 372.414
R513 VDD.t2262 VDD.t2277 372.414
R514 VDD.t1376 VDD.t1386 372.414
R515 VDD.t1380 VDD.t1389 372.414
R516 VDD.t2195 VDD.t2161 372.414
R517 VDD.t2191 VDD.t2170 372.414
R518 VDD.t2460 VDD.t2455 372.414
R519 VDD.t2462 VDD.t2458 372.414
R520 VDD.t242 VDD.t231 372.414
R521 VDD.t252 VDD.t229 372.414
R522 VDD.t1963 VDD.t1969 372.414
R523 VDD.t1961 VDD.t1978 372.414
R524 VDD.t1656 VDD.t1680 372.414
R525 VDD.t1670 VDD.t1650 372.414
R526 VDD.t1369 VDD.t1349 372.414
R527 VDD.t1346 VDD.t1362 372.414
R528 VDD.t2719 VDD.t2728 372.414
R529 VDD.t2741 VDD.t2733 372.414
R530 VDD.t1341 VDD.t1322 372.414
R531 VDD.t1306 VDD.t1334 372.414
R532 VDD.t2592 VDD.t2682 372.414
R533 VDD.t2619 VDD.t2661 372.414
R534 VDD.t41 VDD.t43 372.414
R535 VDD.t38 VDD.t36 372.414
R536 VDD.t1427 VDD.t1421 372.414
R537 VDD.t2749 VDD.t1424 372.414
R538 VDD.t2222 VDD.t2225 372.414
R539 VDD.t2220 VDD.t2228 372.414
R540 VDD.t2525 VDD.t2566 372.414
R541 VDD.t2557 VDD.t2613 372.414
R542 VDD.t2606 VDD.t2609 372.414
R543 VDD.t2617 VDD.t2569 372.414
R544 VDD.t2366 VDD.t2371 372.414
R545 VDD.t2374 VDD.t2368 372.414
R546 VDD.t1011 VDD.t1003 372.414
R547 VDD.t1006 VDD.t1008 372.414
R548 VDD.t112 VDD.t109 372.414
R549 VDD.t117 VDD.t114 372.414
R550 VDD.t801 VDD.t803 367.974
R551 VDD.t799 VDD.t796 367.974
R552 VDD.t827 VDD.t829 367.974
R553 VDD.t832 VDD.t834 367.974
R554 VDD.t1086 VDD.t1092 367.974
R555 VDD.t1084 VDD.t1089 367.974
R556 VDD.t1809 VDD.t1806 367.974
R557 VDD.t1801 VDD.t1803 367.974
R558 VDD.t1041 VDD.t1046 367.974
R559 VDD.t1048 VDD.t1044 367.974
R560 VDD.t124 VDD.t126 367.974
R561 VDD.t132 VDD.t129 367.974
R562 VDD.t2505 VDD.t2520 367.348
R563 VDD.t2495 VDD.t2498 367.348
R564 VDD.t1137 VDD.t1136 367.348
R565 VDD.t1996 VDD.t2005 367.348
R566 VDD.t2008 VDD.t1990 367.348
R567 VDD.t99 VDD.t98 367.348
R568 VDD.t2655 VDD.t2629 367.348
R569 VDD.t2601 VDD.t2560 367.348
R570 VDD.t760 VDD.t762 367.348
R571 VDD.t2036 VDD.t2699 367.348
R572 VDD.t2704 VDD.t2696 367.348
R573 VDD.t1000 VDD.t1002 367.348
R574 VDD.t367 VDD.t368 367.348
R575 VDD.t2042 VDD.t2025 367.348
R576 VDD.t2027 VDD.t2029 367.348
R577 VDD.t2691 VDD.t2692 367.348
R578 VDD.t2563 VDD.t2615 367.348
R579 VDD.t2529 VDD.t2671 367.348
R580 VDD.t2680 VDD.t2668 367.348
R581 VDD.t2547 VDD.t2550 367.348
R582 VDD.t794 VDD.t793 367.348
R583 VDD.t2020 VDD.t2039 367.348
R584 VDD.t2032 VDD.t2022 367.348
R585 VDD.t329 VDD.t330 367.348
R586 VDD.t564 VDD.t562 367.348
R587 VDD.t1828 VDD.t1818 367.348
R588 VDD.t1814 VDD.t1820 367.348
R589 VDD.t728 VDD.t753 367.348
R590 VDD.t743 VDD.t756 367.348
R591 VDD.t894 VDD.t895 367.348
R592 VDD.t740 VDD.t748 367.348
R593 VDD.t746 VDD.t733 367.348
R594 VDD.t736 VDD.t730 367.348
R595 VDD.t750 VDD.t738 367.348
R596 VDD.t954 VDD.t953 367.348
R597 VDD.t1816 VDD.t1811 367.348
R598 VDD.t1826 VDD.t1823 367.348
R599 VDD.t997 VDD.t998 367.348
R600 VDD.t2663 VDD.t2588 367.348
R601 VDD.t2545 VDD.t2645 367.348
R602 VDD.t1027 VDD.t1029 367.348
R603 VDD.t1157 VDD.t1151 367.348
R604 VDD.t1153 VDD.t1162 367.348
R605 VDD.t1741 VDD.t1743 367.348
R606 VDD.t1714 VDD.t1713 367.348
R607 VDD.t2574 VDD.t2531 367.348
R608 VDD.t2537 VDD.t2603 367.348
R609 VDD.t663 VDD.t665 367.348
R610 VDD.t1168 VDD.t1160 367.348
R611 VDD.t1165 VDD.t1155 367.348
R612 VDD.t2643 VDD.t2585 367.348
R613 VDD.t2552 VDD.t2599 367.348
R614 VDD.t1798 VDD.t1800 367.348
R615 VDD.t2386 VDD.t2401 367.348
R616 VDD.t2384 VDD.t2393 367.348
R617 VDD.t287 VDD.t285 367.348
R618 VDD.t317 VDD.t318 367.348
R619 VDD.t2390 VDD.t2388 367.348
R620 VDD.t2399 VDD.t2396 367.348
R621 VDD.t2376 VDD.t2378 367.348
R622 VDD.t2626 VDD.t2527 367.348
R623 VDD.t2590 VDD.t2534 367.348
R624 VDD.t940 VDD.t941 367.348
R625 VDD.t2701 VDD.t2706 367.348
R626 VDD.t2693 VDD.t2034 367.348
R627 VDD.t2201 VDD.t2202 367.348
R628 VDD.t2572 VDD.t2539 367.348
R629 VDD.t2582 VDD.t2641 367.348
R630 VDD.t1767 VDD.t1768 367.348
R631 VDD.t1993 VDD.t1998 367.348
R632 VDD.t2000 VDD.t2002 367.348
R633 VDD.t2503 VDD.t2500 367.348
R634 VDD.t2514 VDD.t2510 367.348
R635 VDD.t437 VDD.t438 367.348
R636 VDD.t2507 VDD.t2512 367.348
R637 VDD.t2523 VDD.t2517 367.348
R638 VDD.n2 VDD.t20 364.93
R639 VDD.n15 VDD.t1187 364.93
R640 VDD.n29 VDD.t1181 364.93
R641 VDD.n830 VDD.t367 360.545
R642 VDD.n819 VDD.t2691 360.545
R643 VDD.n1870 VDD.t564 360.545
R644 VDD.n1859 VDD.t894 360.545
R645 VDD.n1782 VDD.t1714 360.545
R646 VDD.t665 VDD.n2169 360.545
R647 VDD.n2208 VDD.t317 360.545
R648 VDD.n2197 VDD.t2376 360.545
R649 VDD.t941 VDD.n1547 360.545
R650 VDD.n1527 VDD.t2201 360.545
R651 VDD.n1648 VDD.t1767 360.545
R652 VDD.n1637 VDD.t437 360.545
R653 VDD.n1605 VDD.t1137 358.844
R654 VDD.t98 VDD.n1598 358.844
R655 VDD.n1719 VDD.t760 358.844
R656 VDD.n1703 VDD.t1000 358.844
R657 VDD.n793 VDD.t794 358.844
R658 VDD.t330 VDD.n610 358.844
R659 VDD.n1834 VDD.t954 358.844
R660 VDD.t998 VDD.n1827 358.844
R661 VDD.n1905 VDD.t1027 358.844
R662 VDD.n1922 VDD.t1741 358.844
R663 VDD.n1743 VDD.t1798 358.844
R664 VDD.t285 VDD.n1736 358.844
R665 VDD.t450 VDD.t350 357.616
R666 VDD.t2215 VDD.n514 353.481
R667 VDD.n1057 VDD.t402 342.491
R668 VDD.n664 VDD.t658 342.491
R669 VDD.t2203 VDD.n1019 342.491
R670 VDD.t685 VDD.n2412 342.491
R671 VDD.t707 VDD.n1252 342.491
R672 VDD.n522 VDD.t595 342.491
R673 VDD.n1358 VDD.t646 342.491
R674 VDD.t1107 VDD.t865 337.587
R675 VDD.t363 VDD.t766 337.587
R676 VDD.t1132 VDD.t1052 337.587
R677 VDD.t1076 VDD.t905 337.587
R678 VDD.n37 VDD.t789 296.642
R679 VDD.t1039 VDD.n1277 280.519
R680 VDD.t955 VDD.n544 256.555
R681 VDD.t1442 VDD.n2425 252.337
R682 VDD.n1312 VDD.t531 252.337
R683 VDD.t2216 VDD.n546 251.749
R684 VDD.n1070 VDD.t551 251.749
R685 VDD.t774 VDD.n782 251.749
R686 VDD.t629 VDD.n1023 251.749
R687 VDD.n2416 VDD.t67 251.749
R688 VDD.t179 VDD.n1256 251.749
R689 VDD.n1166 VDD.t422 251.749
R690 VDD.n245 VDD.t451 251.749
R691 VDD.n1052 VDD.t557 250.917
R692 VDD.n658 VDD.t1763 250.917
R693 VDD.t327 VDD.n1030 250.917
R694 VDD.n2410 VDD.t782 250.917
R695 VDD.n1250 VDD.t134 250.917
R696 VDD.n544 VDD.t1023 250.917
R697 VDD.t591 VDD.n528 250.917
R698 VDD.t2379 VDD.n1360 250.917
R699 VDD.t1852 VDD.t1918 233.011
R700 VDD.t1834 VDD.t1914 233.011
R701 VDD.t1241 VDD.t1219 233.011
R702 VDD.t1497 VDD.t1556 233.011
R703 VDD.t1519 VDD.t1500 233.011
R704 VDD.t1542 VDD.t1554 233.011
R705 VDD.t1581 VDD.t1575 233.011
R706 VDD.t1210 VDD.t1245 233.011
R707 VDD.t1224 VDD.t1272 233.011
R708 VDD.t1251 VDD.t1289 233.011
R709 VDD.t1849 VDD.t1837 233.011
R710 VDD.t1862 VDD.t1920 233.011
R711 VDD.t1564 VDD.t1485 233.011
R712 VDD.t1502 VDD.t1487 233.011
R713 VDD.t1309 VDD.t1300 233.011
R714 VDD.n123 VDD.t1261 227.617
R715 VDD.n306 VDD.t1479 227.617
R716 VDD.n1319 VDD.t1482 227.617
R717 VDD.n748 VDD.t1489 227.617
R718 VDD.n714 VDD.t1528 227.617
R719 VDD.n620 VDD.t1494 227.617
R720 VDD.n1046 VDD.t1226 227.617
R721 VDD.t1258 VDD.n2452 227.617
R722 VDD.n1106 VDD.t1859 226.537
R723 VDD.t1887 VDD.n1087 226.537
R724 VDD.n1037 VDD.t1286 226.537
R725 VDD.n2457 VDD.t1198 226.537
R726 VDD.n2453 VDD.t1205 226.537
R727 VDD.t1881 VDD.n2405 226.537
R728 VDD.t1847 VDD.n1264 226.537
R729 VDD.t1891 VDD.n1174 226.537
R730 VDD.n1193 VDD.t1879 226.537
R731 VDD.t1567 VDD.n452 226.537
R732 VDD.n471 VDD.t1569 226.537
R733 VDD.n1688 VDD.t1302 226.537
R734 VDD.t1758 VDD.n862 225.712
R735 VDD.n626 VDD.t1533 224.381
R736 VDD.n1051 VDD.t1281 224.381
R737 VDD.n2409 VDD.t1865 224.381
R738 VDD.t1831 VDD.n1263 224.381
R739 VDD.t477 VDD.n1601 215.518
R740 VDD.t2356 VDD.n1591 215.518
R741 VDD.n1708 VDD.t56 215.518
R742 VDD.n1692 VDD.t2334 215.518
R743 VDD.n1473 VDD.t1952 215.518
R744 VDD.n2233 VDD.t2074 215.518
R745 VDD.n2265 VDD.t2485 215.518
R746 VDD.n2269 VDD.t2422 215.518
R747 VDD.n2270 VDD.t2280 215.518
R748 VDD.n2274 VDD.t2295 215.518
R749 VDD.n861 VDD.t2109 215.518
R750 VDD.n838 VDD.t2622 215.518
R751 VDD.n818 VDD.t613 215.518
R752 VDD.t918 VDD.n613 215.518
R753 VDD.t2055 VDD.n603 215.518
R754 VDD.t1391 VDD.n2279 215.518
R755 VDD.t2179 VDD.n2282 215.518
R756 VDD.t1339 VDD.n2281 215.518
R757 VDD.n1414 VDD.t255 215.518
R758 VDD.n2284 VDD.t1976 215.518
R759 VDD.n1400 VDD.t1654 215.518
R760 VDD.n1404 VDD.t1357 215.518
R761 VDD.n1390 VDD.t2736 215.518
R762 VDD.n1858 VDD.t12 215.518
R763 VDD.t1404 VDD.n1830 215.518
R764 VDD.t2156 VDD.n1820 215.518
R765 VDD.n1894 VDD.t1460 215.518
R766 VDD.n1911 VDD.t2241 215.518
R767 VDD.n2002 VDD.t2291 215.518
R768 VDD.n1956 VDD.t1937 215.518
R769 VDD.n1963 VDD.t2058 215.518
R770 VDD.n1964 VDD.t2473 215.518
R771 VDD.n1994 VDD.t2417 215.518
R772 VDD.n1995 VDD.t2270 215.518
R773 VDD.n2130 VDD.t1376 215.518
R774 VDD.n2116 VDD.t2161 215.518
R775 VDD.n2117 VDD.t2460 215.518
R776 VDD.n2099 VDD.t242 215.518
R777 VDD.n2106 VDD.t1969 215.518
R778 VDD.n2085 VDD.t1680 215.518
R779 VDD.n2086 VDD.t1369 215.518
R780 VDD.n2075 VDD.t2728 215.518
R781 VDD.n2054 VDD.t1341 215.518
R782 VDD.n1790 VDD.t2592 215.518
R783 VDD.t1424 VDD.n1739 215.518
R784 VDD.t2228 VDD.n1729 215.518
R785 VDD.n2216 VDD.t2525 215.518
R786 VDD.n1723 VDD.t2609 215.518
R787 VDD.n2196 VDD.t2366 215.518
R788 VDD.n1526 VDD.t1011 215.518
R789 VDD.n1636 VDD.t112 215.518
R790 VDD.n829 VDD.t801 212.947
R791 VDD.n1869 VDD.t827 212.947
R792 VDD.t1092 VDD.n2167 212.947
R793 VDD.n2207 VDD.t1809 212.947
R794 VDD.t1046 VDD.n1548 212.947
R795 VDD.n1647 VDD.t124 212.947
R796 VDD.n1606 VDD.t2495 212.585
R797 VDD.t1990 VDD.n1595 212.585
R798 VDD.t2560 VDD.n1718 212.585
R799 VDD.t2696 VDD.n1702 212.585
R800 VDD.n837 VDD.t2025 212.585
R801 VDD.n823 VDD.t2615 212.585
R802 VDD.n794 VDD.t2547 212.585
R803 VDD.t2022 VDD.n607 212.585
R804 VDD.n1877 VDD.t1818 212.585
R805 VDD.n1878 VDD.t728 212.585
R806 VDD.n1863 VDD.t748 212.585
R807 VDD.n1835 VDD.t750 212.585
R808 VDD.t1823 VDD.n1824 212.585
R809 VDD.t2645 VDD.n1904 212.585
R810 VDD.t1162 VDD.n1921 212.585
R811 VDD.n1786 VDD.t2574 212.585
R812 VDD.t1160 VDD.n2168 212.585
R813 VDD.n1744 VDD.t2552 212.585
R814 VDD.t2393 VDD.n1733 212.585
R815 VDD.n2215 VDD.t2388 212.585
R816 VDD.n2201 VDD.t2527 212.585
R817 VDD.t2706 VDD.n1546 212.585
R818 VDD.n1549 VDD.t2572 212.585
R819 VDD.n1655 VDD.t1998 212.585
R820 VDD.n1656 VDD.t2503 212.585
R821 VDD.n1641 VDD.t2512 212.585
R822 VDD.t31 VDD.t1758 211.974
R823 VDD.t1755 VDD.t267 211.974
R824 VDD.t2714 VDD.t1107 211.974
R825 VDD.t763 VDD.t1110 211.974
R826 VDD.t2231 VDD.t363 211.974
R827 VDD.t771 VDD.t1736 211.974
R828 VDD.t1987 VDD.t1132 211.974
R829 VDD.t902 VDD.t1795 211.974
R830 VDD.t452 VDD.t1076 211.974
R831 VDD.t489 VDD.t1071 211.974
R832 VDD.t458 VDD.t457 209.101
R833 VDD.t1731 VDD.t1734 209.101
R834 VDD.t770 VDD.t769 209.101
R835 VDD.t296 VDD.t293 209.101
R836 VDD.t2045 VDD.t2046 209.101
R837 VDD.t603 VDD.t606 209.101
R838 VDD.t1149 VDD.t1150 209.101
R839 VDD.t806 VDD.t808 209.101
R840 VDD.t398 VDD.t399 209.101
R841 VDD.t265 VDD.t262 209.101
R842 VDD.t861 VDD.t862 209.101
R843 VDD.t249 VDD.t240 209.101
R844 VDD.t441 VDD.t442 209.101
R845 VDD.t666 VDD.t669 209.101
R846 VDD.t981 VDD.t980 209.101
R847 VDD.t987 VDD.t990 209.101
R848 VDD.t401 VDD.t400 209.101
R849 VDD.t75 VDD.t73 209.101
R850 VDD.t408 VDD.t407 209.101
R851 VDD.t580 VDD.t578 209.101
R852 VDD.t370 VDD.t369 209.101
R853 VDD.t844 VDD.t842 209.101
R854 VDD.t758 VDD.t759 209.101
R855 VDD.t1726 VDD.t1728 209.101
R856 VDD.t64 VDD.t65 209.101
R857 VDD.t237 VDD.t227 209.101
R858 VDD.t1414 VDD.t1415 209.101
R859 VDD.t636 VDD.t633 209.101
R860 VDD.t24 VDD.t22 204.739
R861 VDD.t20 VDD.t24 204.739
R862 VDD.t2122 VDD.t2120 204.739
R863 VDD.t2125 VDD.t2122 204.739
R864 VDD.t1191 VDD.t1189 204.739
R865 VDD.t1187 VDD.t1191 204.739
R866 VDD.t2117 VDD.t2115 204.739
R867 VDD.t2111 VDD.t2117 204.739
R868 VDD.t1178 VDD.t1176 204.739
R869 VDD.t1181 VDD.t1178 204.739
R870 VDD.t2113 VDD.t2127 204.739
R871 VDD.t2127 VDD.t2130 204.739
R872 VDD.n545 VDD.t2218 202.248
R873 VDD.n1353 VDD.t1775 200.87
R874 VDD.n482 VDD.t2576 197.803
R875 VDD.n482 VDD.t2624 197.803
R876 VDD.n547 VDD.t2465 197.803
R877 VDD.n547 VDD.t2475 197.803
R878 VDD.n1098 VDD.t2185 197.803
R879 VDD.t2189 VDD.n1098 197.803
R880 VDD.n1278 VDD.t2634 197.803
R881 VDD.n1278 VDD.t2639 197.803
R882 VDD.n1079 VDD.t554 197.803
R883 VDD.t552 VDD.n1079 197.803
R884 VDD.n2444 VDD.t2658 197.803
R885 VDD.n2444 VDD.t2597 197.803
R886 VDD.n158 VDD.t702 197.803
R887 VDD.n158 VDD.t700 197.803
R888 VDD.n2442 VDD.t2066 197.803
R889 VDD.t2088 VDD.n2442 197.803
R890 VDD.n425 VDD.t1313 197.803
R891 VDD.n425 VDD.t1328 197.803
R892 VDD.n307 VDD.t234 197.803
R893 VDD.n307 VDD.t225 197.803
R894 VDD.n321 VDD.t2542 197.803
R895 VDD.t2650 VDD.n321 197.803
R896 VDD.n1320 VDD.t311 197.803
R897 VDD.t314 VDD.n1320 197.803
R898 VDD.n1336 VDD.t1366 197.803
R899 VDD.t1364 VDD.n1336 197.803
R900 VDD.n360 VDD.t1942 197.803
R901 VDD.n360 VDD.t1935 197.803
R902 VDD.n1056 VDD.t924 197.803
R903 VDD.t930 VDD.n1056 197.803
R904 VDD.n724 VDD.t2652 197.803
R905 VDD.n724 VDD.t2666 197.803
R906 VDD.n768 VDD.t2267 197.803
R907 VDD.t2282 VDD.n768 197.803
R908 VDD.n749 VDD.t725 197.803
R909 VDD.t723 VDD.n749 197.803
R910 VDD.n735 VDD.t2310 197.803
R911 VDD.t2297 VDD.n735 197.803
R912 VDD.n663 VDD.t0 197.803
R913 VDD.t3 VDD.n663 197.803
R914 VDD.n783 VDD.t2257 197.803
R915 VDD.n783 VDD.t2260 197.803
R916 VDD.n1024 VDD.t1336 197.803
R917 VDD.n1024 VDD.t1304 197.803
R918 VDD.t2248 VDD.n1018 197.803
R919 VDD.n1018 VDD.t2251 197.803
R920 VDD.n82 VDD.t2677 197.803
R921 VDD.n82 VDD.t2555 197.803
R922 VDD.t274 VDD.n2458 197.803
R923 VDD.n2458 VDD.t272 197.803
R924 VDD.t2594 VDD.n2454 197.803
R925 VDD.n2454 VDD.t2611 197.803
R926 VDD.n2426 VDD.t1949 197.803
R927 VDD.n2426 VDD.t1947 197.803
R928 VDD.n2394 VDD.t1981 197.803
R929 VDD.n2394 VDD.t1957 197.803
R930 VDD.t618 VDD.n2411 197.803
R931 VDD.n2411 VDD.t624 197.803
R932 VDD.n1299 VDD.t1984 197.803
R933 VDD.n1299 VDD.t1959 197.803
R934 VDD.n1257 VDD.t2743 197.803
R935 VDD.n1257 VDD.t2722 197.803
R936 VDD.t2443 VDD.n1251 197.803
R937 VDD.n1251 VDD.t2446 197.803
R938 VDD.n1204 VDD.t2631 197.803
R939 VDD.n1204 VDD.t2648 197.803
R940 VDD.n1173 VDD.t837 197.803
R941 VDD.t840 VDD.n1173 197.803
R942 VDD.t1647 VDD.n1185 197.803
R943 VDD.t1682 VDD.n1185 197.803
R944 VDD.t2746 VDD.n1165 197.803
R945 VDD.n1165 VDD.t2724 197.803
R946 VDD.n244 VDD.t1352 197.803
R947 VDD.t1355 VDD.n244 197.803
R948 VDD.n525 VDD.t89 197.803
R949 VDD.t85 VDD.n525 197.803
R950 VDD.t1432 VDD.n1359 197.803
R951 VDD.n1359 VDD.t2018 197.803
R952 VDD.n573 VDD.t2480 197.803
R953 VDD.n573 VDD.t2487 197.803
R954 VDD.t648 VDD.n444 197.803
R955 VDD.t651 VDD.n444 197.803
R956 VDD.t2425 VDD.n463 197.803
R957 VDD.t2439 VDD.n463 197.803
R958 VDD.n1383 VDD.t2406 197.803
R959 VDD.t2404 VDD.n1383 197.803
R960 VDD.n1384 VDD.t866 197.803
R961 VDD.t869 VDD.n1384 197.803
R962 VDD.n2066 VDD.t49 197.803
R963 VDD.t52 VDD.n2066 197.803
R964 VDD.n2067 VDD.t936 197.803
R965 VDD.n2067 VDD.t934 197.803
R966 VDD.n1687 VDD.t2351 197.803
R967 VDD.t2354 VDD.n1687 197.803
R968 VDD.n1680 VDD.t2151 197.803
R969 VDD.n1680 VDD.t2144 197.803
R970 VDD.t221 VDD.t220 196.721
R971 VDD.t1661 VDD.t1664 196.721
R972 VDD.t2414 VDD.t2290 196.721
R973 VDD.t1383 VDD.t1384 196.721
R974 VDD.t2163 VDD.t2176 196.721
R975 VDD.n1061 VDD.t353 196.523
R976 VDD.n668 VDD.t383 196.523
R977 VDD.t2211 VDD.n1021 196.523
R978 VDD.t688 VDD.n2414 196.523
R979 VDD.t672 VDD.n1254 196.523
R980 VDD.n1354 VDD.t448 195.971
R981 VDD.t1248 VDD.n1036 193.096
R982 VDD.t884 VDD.t886 187.827
R983 VDD.t889 VDD.t884 187.827
R984 VDD.t912 VDD.t889 187.827
R985 VDD.t913 VDD.t908 187.827
R986 VDD.t717 VDD.t715 187.827
R987 VDD.t715 VDD.t927 187.827
R988 VDD.t353 VDD.t357 187.827
R989 VDD.t549 VDD.t550 187.827
R990 VDD.t383 VDD.t386 187.827
R991 VDD.t776 VDD.t775 187.827
R992 VDD.t1467 VDD.t1472 187.827
R993 VDD.t1472 VDD.t2318 187.827
R994 VDD.t2318 VDD.t1474 187.827
R995 VDD.t1470 VDD.t1471 187.827
R996 VDD.t2685 VDD.t2688 187.827
R997 VDD.t2688 VDD.t5 187.827
R998 VDD.t492 VDD.t2246 187.827
R999 VDD.t495 VDD.t492 187.827
R1000 VDD.t1751 VDD.t1749 187.827
R1001 VDD.t1750 VDD.t207 187.827
R1002 VDD.t207 VDD.t204 187.827
R1003 VDD.t204 VDD.t202 187.827
R1004 VDD.t628 VDD.t626 187.827
R1005 VDD.t627 VDD.t2211 187.827
R1006 VDD.t621 VDD.t414 187.827
R1007 VDD.t414 VDD.t417 187.827
R1008 VDD.t1453 VDD.t1450 187.827
R1009 VDD.t1450 VDD.t1448 187.827
R1010 VDD.t68 VDD.t66 187.827
R1011 VDD.t69 VDD.t688 187.827
R1012 VDD.t899 VDD.t2441 187.827
R1013 VDD.t897 VDD.t899 187.827
R1014 VDD.t871 VDD.t876 187.827
R1015 VDD.t876 VDD.t873 187.827
R1016 VDD.t181 VDD.t180 187.827
R1017 VDD.t178 VDD.t672 187.827
R1018 VDD.t1775 VDD.t1783 187.827
R1019 VDD.t1783 VDD.t1778 187.827
R1020 VDD.t1778 VDD.t2708 187.827
R1021 VDD.t2709 VDD.t2710 187.827
R1022 VDD.t459 VDD.t461 187.827
R1023 VDD.t1429 VDD.t459 187.827
R1024 VDD.t419 VDD.t421 187.827
R1025 VDD.t420 VDD.t1693 187.827
R1026 VDD.t513 VDD.t510 187.663
R1027 VDD.t1441 VDD.t1440 187.663
R1028 VDD.t102 VDD.t532 187.663
R1029 VDD.t537 VDD.t533 187.663
R1030 VDD.n1313 VDD.t912 186.088
R1031 VDD.t1474 VDD.n781 186.088
R1032 VDD.t2708 VDD.n1352 186.088
R1033 VDD.n999 VDD.t1750 185.218
R1034 VDD.t1040 VDD.t949 180.905
R1035 VDD.t427 VDD.t423 180.905
R1036 VDD.n245 VDD.t450 178.809
R1037 VDD.n22 VDD.t2111 164.929
R1038 VDD.n1355 VDD.n1354 157.51
R1039 VDD.n2417 VDD.t1453 157.392
R1040 VDD.n1601 VDD.t482 156.898
R1041 VDD.n1591 VDD.t2359 156.898
R1042 VDD.n1708 VDD.t54 156.898
R1043 VDD.n1692 VDD.t2332 156.898
R1044 VDD.n1473 VDD.t1930 156.898
R1045 VDD.n2233 VDD.t2083 156.898
R1046 VDD.t2468 VDD.n2265 156.898
R1047 VDD.t2433 VDD.n2269 156.898
R1048 VDD.n2270 VDD.t2254 156.898
R1049 VDD.n2274 VDD.t2287 156.898
R1050 VDD.t2047 VDD.n861 156.898
R1051 VDD.n838 VDD.t2674 156.898
R1052 VDD.t610 VDD.n818 156.898
R1053 VDD.n613 VDD.t914 156.898
R1054 VDD.n603 VDD.t2053 156.898
R1055 VDD.n2279 VDD.t1393 156.898
R1056 VDD.n2282 VDD.t2182 156.898
R1057 VDD.n2281 VDD.t1316 156.898
R1058 VDD.t222 VDD.n1414 156.898
R1059 VDD.n2284 VDD.t1966 156.898
R1060 VDD.t1666 VDD.n1400 156.898
R1061 VDD.t1359 VDD.n1404 156.898
R1062 VDD.t2738 VDD.n1390 156.898
R1063 VDD.t14 VDD.n1858 156.898
R1064 VDD.n1830 VDD.t1412 156.898
R1065 VDD.n1820 VDD.t2154 156.898
R1066 VDD.n1894 VDD.t1465 156.898
R1067 VDD.n1911 VDD.t2244 156.898
R1068 VDD.n2002 VDD.t2303 156.898
R1069 VDD.t1954 VDD.n1956 156.898
R1070 VDD.t2070 VDD.n1963 156.898
R1071 VDD.t2489 VDD.n1964 156.898
R1072 VDD.t2419 VDD.n1994 156.898
R1073 VDD.t2277 VDD.n1995 156.898
R1074 VDD.n2130 VDD.t1380 156.898
R1075 VDD.t2170 VDD.n2116 156.898
R1076 VDD.n2117 VDD.t2462 156.898
R1077 VDD.n2099 VDD.t252 156.898
R1078 VDD.t1978 VDD.n2106 156.898
R1079 VDD.t1650 VDD.n2085 156.898
R1080 VDD.n2086 VDD.t1346 156.898
R1081 VDD.t2733 VDD.n2075 156.898
R1082 VDD.n2054 VDD.t1306 156.898
R1083 VDD.n1790 VDD.t2619 156.898
R1084 VDD.n1739 VDD.t1427 156.898
R1085 VDD.n1729 VDD.t2222 156.898
R1086 VDD.n2216 VDD.t2557 156.898
R1087 VDD.t2569 VDD.n1723 156.898
R1088 VDD.t2368 VDD.n2196 156.898
R1089 VDD.t1008 VDD.n1526 156.898
R1090 VDD.t114 VDD.n1636 156.898
R1091 VDD.n1227 VDD.t871 155.653
R1092 VDD.t796 VDD.n829 155.026
R1093 VDD.t834 VDD.n1869 155.026
R1094 VDD.n2167 VDD.t1089 155.026
R1095 VDD.t1803 VDD.n2207 155.026
R1096 VDD.n1548 VDD.t1048 155.026
R1097 VDD.t129 VDD.n1647 155.026
R1098 VDD.n1606 VDD.t2505 154.762
R1099 VDD.n1595 VDD.t1996 154.762
R1100 VDD.n1718 VDD.t2629 154.762
R1101 VDD.n1702 VDD.t2699 154.762
R1102 VDD.t2029 VDD.n837 154.762
R1103 VDD.t2671 VDD.n823 154.762
R1104 VDD.n794 VDD.t2680 154.762
R1105 VDD.n607 VDD.t2020 154.762
R1106 VDD.t1820 VDD.n1877 154.762
R1107 VDD.n1878 VDD.t743 154.762
R1108 VDD.t733 VDD.n1863 154.762
R1109 VDD.n1835 VDD.t736 154.762
R1110 VDD.n1824 VDD.t1816 154.762
R1111 VDD.n1904 VDD.t2588 154.762
R1112 VDD.n1921 VDD.t1151 154.762
R1113 VDD.t2603 VDD.n1786 154.762
R1114 VDD.n2168 VDD.t1165 154.762
R1115 VDD.n1744 VDD.t2643 154.762
R1116 VDD.n1733 VDD.t2386 154.762
R1117 VDD.t2396 VDD.n2215 154.762
R1118 VDD.t2534 VDD.n2201 154.762
R1119 VDD.n1546 VDD.t2693 154.762
R1120 VDD.n1549 VDD.t2582 154.762
R1121 VDD.t2002 VDD.n1655 154.762
R1122 VDD.n1656 VDD.t2514 154.762
R1123 VDD.t2517 VDD.n1641 154.762
R1124 VDD.n544 VDD.t958 147.94
R1125 VDD.n2443 VDD.t277 145.662
R1126 VDD.t520 VDD.n322 145.662
R1127 VDD.t969 VDD.n1337 145.662
R1128 VDD.t847 VDD.n769 145.662
R1129 VDD.t1096 VDD.n736 145.662
R1130 VDD.t173 VDD.n2459 145.662
R1131 VDD.t1033 VDD.n2455 145.662
R1132 VDD.n1203 VDD.t144 145.662
R1133 VDD.n572 VDD.t855 145.662
R1134 VDD.n481 VDD.t156 145.662
R1135 VDD.n1679 VDD.t821 145.662
R1136 VDD.n2175 VDD.t41 144.828
R1137 VDD.n1052 VDD.t560 144.69
R1138 VDD.t1761 VDD.n658 144.69
R1139 VDD.n1030 VDD.t324 144.69
R1140 VDD.t784 VDD.n2410 144.69
R1141 VDD.t136 VDD.n1250 144.69
R1142 VDD.n544 VDD.t1020 144.69
R1143 VDD.n528 VDD.t588 144.69
R1144 VDD.n1360 VDD.t2382 144.69
R1145 VDD.n863 VDD.t31 143.279
R1146 VDD.n2227 VDD.t2714 143.279
R1147 VDD.n2228 VDD.t2231 143.279
R1148 VDD.n1937 VDD.t1987 143.279
R1149 VDD.n2146 VDD.t452 143.279
R1150 VDD.n2173 VDD.t38 137.931
R1151 VDD.n877 VDD.t2064 137.524
R1152 VDD.t2224 VDD.t977 136.796
R1153 VDD.t2219 VDD.t2329 136.796
R1154 VDD.t164 VDD.t277 136.796
R1155 VDD.t165 VDD.t163 136.796
R1156 VDD.t517 VDD.t520 136.796
R1157 VDD.t1143 VDD.t1144 136.796
R1158 VDD.t816 VDD.t969 136.796
R1159 VDD.t817 VDD.t526 136.796
R1160 VDD.t476 VDD.t847 136.796
R1161 VDD.t474 VDD.t475 136.796
R1162 VDD.t1065 VDD.t1096 136.796
R1163 VDD.t1063 VDD.t1064 136.796
R1164 VDD.t1126 VDD.t546 136.796
R1165 VDD.t171 VDD.t173 136.796
R1166 VDD.t575 VDD.t864 136.796
R1167 VDD.t863 VDD.t1033 136.796
R1168 VDD.t372 VDD.t371 136.796
R1169 VDD.t144 VDD.t147 136.796
R1170 VDD.t80 VDD.t79 136.796
R1171 VDD.t855 VDD.t78 136.796
R1172 VDD.t951 VDD.t720 136.796
R1173 VDD.t156 VDD.t160 136.796
R1174 VDD.t1475 VDD.t190 136.796
R1175 VDD.t1456 VDD.t2338 136.796
R1176 VDD.t47 VDD.t48 136.796
R1177 VDD.t821 VDD.t46 136.796
R1178 VDD.n876 VDD.t221 133.881
R1179 VDD.n998 VDD.t1384 133.881
R1180 VDD.n1569 VDD.t2224 122.23
R1181 VDD.t163 VDD.n116 122.23
R1182 VDD.n323 VDD.t1143 122.23
R1183 VDD.n1338 VDD.t817 122.23
R1184 VDD.n770 VDD.t474 122.23
R1185 VDD.n737 VDD.t1063 122.23
R1186 VDD.n2460 VDD.t1126 122.23
R1187 VDD.t864 VDD.n2456 122.23
R1188 VDD.n1177 VDD.t372 122.23
R1189 VDD.n436 VDD.t80 122.23
R1190 VDD.n455 VDD.t951 122.23
R1191 VDD.n1883 VDD.t1475 122.23
R1192 VDD.n1678 VDD.t47 122.23
R1193 VDD.t2414 VDD.t2284 116.947
R1194 VDD.t2414 VDD.t2060 116.947
R1195 VDD.n2232 VDD.t457 114.231
R1196 VDD.n2266 VDD.t770 114.231
R1197 VDD.n2273 VDD.t2046 114.231
R1198 VDD.t1150 VDD.n2280 114.231
R1199 VDD.t399 VDD.n2283 114.231
R1200 VDD.n1405 VDD.t861 114.231
R1201 VDD.n1391 VDD.t441 114.231
R1202 VDD.n1957 VDD.t981 114.231
R1203 VDD.n1993 VDD.t401 114.231
R1204 VDD.n1996 VDD.t408 114.231
R1205 VDD.n2129 VDD.t369 114.231
R1206 VDD.n2107 VDD.t758 114.231
R1207 VDD.n2098 VDD.t65 114.231
R1208 VDD.n2076 VDD.t1414 114.231
R1209 VDD.n2424 VDD.t2015 111.305
R1210 VDD.n1130 VDD.t2453 108.697
R1211 VDD.n37 VDD.t787 106.344
R1212 VDD.n1226 VDD.n1225 106.088
R1213 VDD.n2366 VDD.n2365 101.74
R1214 VDD.t1734 VDD.n2232 94.8698
R1215 VDD.n2266 VDD.t296 94.8698
R1216 VDD.t606 VDD.n2273 94.8698
R1217 VDD.n2280 VDD.t806 94.8698
R1218 VDD.n2283 VDD.t265 94.8698
R1219 VDD.t240 VDD.n1405 94.8698
R1220 VDD.t669 VDD.n1391 94.8698
R1221 VDD.t990 VDD.n1957 94.8698
R1222 VDD.t73 VDD.n1993 94.8698
R1223 VDD.t578 VDD.n1996 94.8698
R1224 VDD.t842 VDD.n2129 94.8698
R1225 VDD.n2107 VDD.t1726 94.8698
R1226 VDD.t227 VDD.n2098 94.8698
R1227 VDD.n2076 VDD.t636 94.8698
R1228 VDD.t550 VDD.n1070 93.9135
R1229 VDD.n782 VDD.t776 93.9135
R1230 VDD.n1023 VDD.t626 93.9135
R1231 VDD.t66 VDD.n2416 93.9135
R1232 VDD.n1256 VDD.t180 93.9135
R1233 VDD.n1166 VDD.t419 93.9135
R1234 VDD.n2425 VDD.t1441 93.832
R1235 VDD.t532 VDD.n1312 93.832
R1236 VDD.n1277 VDD.t1040 90.4528
R1237 VDD.t2011 VDD.n2366 83.4788
R1238 VDD.n1130 VDD.t2452 79.1309
R1239 VDD.t2449 VDD.n1226 79.1309
R1240 VDD.t2010 VDD.n2424 76.5222
R1241 VDD.n1070 VDD.n1069 73.9135
R1242 VDD.n782 VDD.n635 73.9135
R1243 VDD.n1023 VDD.n1022 73.9135
R1244 VDD.n2416 VDD.n2415 73.9135
R1245 VDD.n1256 VDD.n1255 73.9135
R1246 VDD.n1167 VDD.n1166 73.9135
R1247 VDD.n2425 VDD.n167 73.8493
R1248 VDD.n1312 VDD.n1311 73.8493
R1249 VDD.n1277 VDD.n1090 71.1898
R1250 VDD.t2120 VDD.n2 71.0905
R1251 VDD.t2115 VDD.n15 71.0905
R1252 VDD.n29 VDD.t2113 71.0905
R1253 VDD.n2175 VDD.n2174 70.6902
R1254 VDD.n863 VDD.t1755 68.6953
R1255 VDD.t1110 VDD.n2227 68.6953
R1256 VDD.n2228 VDD.t771 68.6953
R1257 VDD.t1795 VDD.n1937 68.6953
R1258 VDD.n2146 VDD.t489 68.6953
R1259 VDD.n546 VDD.n545 63.1204
R1260 VDD.t1664 VDD.n876 62.842
R1261 VDD.t2176 VDD.n998 62.842
R1262 VDD.n877 VDD.t2414 59.199
R1263 VDD.n1057 VDD.t404 53.1141
R1264 VDD.n664 VDD.t660 53.1141
R1265 VDD.n1019 VDD.t2206 53.1141
R1266 VDD.n2412 VDD.t683 53.1141
R1267 VDD.n1252 VDD.t705 53.1141
R1268 VDD.t593 VDD.n522 53.1141
R1269 VDD.t643 VDD.n1358 53.1141
R1270 VDD.n2230 VDD 44.41
R1271 VDD VDD.n2145 44.41
R1272 VDD.t193 VDD.n514 42.125
R1273 VDD.t347 VDD.n1355 42.125
R1274 VDD.n1227 VDD.t2449 32.1744
R1275 VDD.n1036 VDD.n376 31.2842
R1276 VDD.n1365 VDD.t1507 31.136
R1277 VDD.n1363 VDD.t1511 31.136
R1278 VDD.n2417 VDD.t2011 30.4353
R1279 VDD.t1494 VDD.n619 24.6392
R1280 VDD.n2407 VDD.t1881 24.6392
R1281 VDD.n1266 VDD.t1847 24.6392
R1282 VDD.t908 VDD.t717 24.3483
R1283 VDD.t1471 VDD.t2685 24.3483
R1284 VDD.t1749 VDD.t495 24.3483
R1285 VDD.t417 VDD.t2010 24.3483
R1286 VDD.t2452 VDD.t897 24.3483
R1287 VDD.t461 VDD.t2709 24.3483
R1288 VDD.n1060 VDD.t402 21.9785
R1289 VDD.n667 VDD.t658 21.9785
R1290 VDD.n1020 VDD.t2203 21.9785
R1291 VDD.n2413 VDD.t685 21.9785
R1292 VDD.n1253 VDD.t707 21.9785
R1293 VDD.t595 VDD.n521 21.9785
R1294 VDD.t646 VDD.n1357 21.9785
R1295 VDD.n1069 VDD.t357 20.0005
R1296 VDD.t386 VDD.n635 20.0005
R1297 VDD.n1022 VDD.t627 20.0005
R1298 VDD.n2415 VDD.t69 20.0005
R1299 VDD.n1255 VDD.t178 20.0005
R1300 VDD.n1167 VDD.t420 20.0005
R1301 VDD.n167 VDD.t510 19.9831
R1302 VDD.n1311 VDD.t533 19.9831
R1303 VDD.t423 VDD.n1090 19.2635
R1304 VDD.n2174 VDD.n2173 18.966
R1305 VDD.n1040 VDD.t1286 18.3392
R1306 VDD.t1226 VDD.n1045 18.3392
R1307 VDD.n2224 VDD.t1057 16.2823
R1308 VDD.n1500 VDD.t1061 16.2823
R1309 VDD.n2150 VDD.t1059 16.2823
R1310 VDD.n1924 VDD.t1051 16.2823
R1311 VDD.n843 VDD.t1054 16.2775
R1312 VDD.n530 VDD.t1584 14.6525
R1313 VDD.n1361 VDD.t1476 14.6525
R1314 VDD.n1569 VDD.t2219 14.5667
R1315 VDD.n116 VDD.t164 14.5667
R1316 VDD.n323 VDD.t517 14.5667
R1317 VDD.n1338 VDD.t816 14.5667
R1318 VDD.n770 VDD.t476 14.5667
R1319 VDD.n737 VDD.t1065 14.5667
R1320 VDD.n2460 VDD.t171 14.5667
R1321 VDD.n2456 VDD.t863 14.5667
R1322 VDD.t147 VDD.n1177 14.5667
R1323 VDD.t78 VDD.n436 14.5667
R1324 VDD.t160 VDD.n455 14.5667
R1325 VDD.n1883 VDD.t1456 14.5667
R1326 VDD.t46 VDD.n1678 14.5667
R1327 VDD.n1634 VDD 12.4951
R1328 VDD.n1454 VDD.t2294 12.4261
R1329 VDD.n2006 VDD.t2314 12.4261
R1330 VDD.n1455 VDD.n1451 12.3181
R1331 VDD.n2007 VDD.n2003 12.3181
R1332 VDD.n2467 VDD.n2466 11.1843
R1333 VDD.t1558 VDD.n529 10.9895
R1334 VDD.n1721 VDD.n1720 10.0532
R1335 VDD.n841 VDD.n840 9.49846
R1336 VDD.n869 VDD.n868 9.31626
R1337 VDD.n1362 VDD.t1633 9.15801
R1338 VDD.t1561 VDD.n626 8.63049
R1339 VDD.t1236 VDD.n1051 8.63049
R1340 VDD.t1857 VDD.n2409 8.63049
R1341 VDD.n1263 VDD.t1912 8.63049
R1342 VDD.t1135 VDD.n1605 8.5039
R1343 VDD.n1598 VDD.t97 8.5039
R1344 VDD.n1719 VDD.t761 8.5039
R1345 VDD.n1703 VDD.t1001 8.5039
R1346 VDD.t795 VDD.n793 8.5039
R1347 VDD.n610 VDD.t331 8.5039
R1348 VDD.t952 VDD.n1834 8.5039
R1349 VDD.n1827 VDD.t999 8.5039
R1350 VDD.n1905 VDD.t1028 8.5039
R1351 VDD.n1922 VDD.t1742 8.5039
R1352 VDD.t1799 VDD.n1743 8.5039
R1353 VDD.n1736 VDD.t286 8.5039
R1354 VDD.n779 VDD.n778 8.10277
R1355 VDD.n2430 VDD.n143 8.10232
R1356 VDD.n1350 VDD.n1349 8.10232
R1357 VDD.n1303 VDD.n177 8.10201
R1358 VDD.n1221 VDD.n1220 8.10201
R1359 VDD.n430 VDD.n429 8.10155
R1360 VDD.n577 VDD.n565 8.10155
R1361 VDD.n2194 VDD.n2193 7.99248
R1362 VDD.n1691 VDD.n1690 7.78414
R1363 VDD.n1881 VDD.n1804 7.7598
R1364 VDD.n2219 VDD.n1501 7.7598
R1365 VDD.n1727 VDD.t2375 7.64083
R1366 VDD.n1525 VDD.t1007 7.64083
R1367 VDD.n2194 VDD.n1724 7.5993
R1368 VDD.n1554 VDD.n1522 7.5993
R1369 VDD.n1660 VDD.n1659 7.58495
R1370 VDD.n815 VDD.n814 7.53174
R1371 VDD.n1855 VDD.n1854 7.53174
R1372 VDD.n1626 VDD.n1625 7.53174
R1373 VDD.n2277 VDD.n2276 7.44996
R1374 VDD.n2133 VDD.n2132 7.44996
R1375 VDD.n2463 VDD.n2462 7.31403
R1376 VDD.n2423 VDD.n168 6.99457
R1377 VDD.n2418 VDD.n178 6.99457
R1378 VDD.n2257 VDD.t2273 6.93712
R1379 VDD.n2241 VDD.n2240 6.93712
R1380 VDD.n1471 VDD.t1946 6.93712
R1381 VDD.n1987 VDD.t2263 6.93712
R1382 VDD.n1971 VDD.n1970 6.93712
R1383 VDD.n1953 VDD.t1934 6.93712
R1384 VDD.n1472 VDD.n1468 6.90536
R1385 VDD.n1954 VDD.n1950 6.90536
R1386 VDD.n2354 VDD.n181 6.87374
R1387 VDD.n1224 VDD.n1131 6.8344
R1388 VDD.n1228 VDD.n1129 6.8344
R1389 VDD.n830 VDD.t366 6.80322
R1390 VDD.n819 VDD.t2690 6.80322
R1391 VDD.n1870 VDD.t563 6.80322
R1392 VDD.n1859 VDD.t896 6.80322
R1393 VDD.t1715 VDD.n1782 6.80322
R1394 VDD.n2169 VDD.t664 6.80322
R1395 VDD.n2208 VDD.t316 6.80322
R1396 VDD.n2197 VDD.t2377 6.80322
R1397 VDD.n1547 VDD.t939 6.80322
R1398 VDD.t2200 VDD.n1527 6.80322
R1399 VDD.n1648 VDD.t1766 6.80322
R1400 VDD.n1637 VDD.t436 6.80322
R1401 VDD.n136 VDD.n134 6.76079
R1402 VDD.n678 VDD.n676 6.76079
R1403 VDD.n263 VDD.n261 6.76079
R1404 VDD.n404 VDD.t496 6.76023
R1405 VDD.n173 VDD.t418 6.76023
R1406 VDD.n1136 VDD.t898 6.76023
R1407 VDD.n501 VDD.t93 6.76023
R1408 VDD.n2420 VDD.n2356 6.7505
R1409 VDD.n2355 VDD.n180 6.7505
R1410 VDD.n1369 VDD.n1368 6.7505
R1411 VDD.n2314 VDD.n2313 6.7505
R1412 VDD.n1224 VDD.n1129 6.51406
R1413 VDD.n1106 VDD.t1852 6.47299
R1414 VDD.n1087 VDD.t1834 6.47299
R1415 VDD.n1037 VDD.t1248 6.47299
R1416 VDD.t1245 VDD.n2457 6.47299
R1417 VDD.t1272 VDD.n2453 6.47299
R1418 VDD.n2405 VDD.t1865 6.47299
R1419 VDD.n1264 VDD.t1831 6.47299
R1420 VDD.n1174 VDD.t1849 6.47299
R1421 VDD.n1193 VDD.t1862 6.47299
R1422 VDD.n452 VDD.t1564 6.47299
R1423 VDD.n471 VDD.t1502 6.47299
R1424 VDD.n1688 VDD.t1309 6.47299
R1425 VDD.n2190 VDD.n2189 6.46984
R1426 VDD.n1574 VDD.n1569 6.3005
R1427 VDD.n1624 VDD.n1591 6.3005
R1428 VDD.n1620 VDD.n1595 6.3005
R1429 VDD.n1617 VDD.n1598 6.3005
R1430 VDD VDD.n1599 6.3005
R1431 VDD.n1615 VDD.n1601 6.3005
R1432 VDD.n1611 VDD.n1606 6.3005
R1433 VDD.n1693 VDD.n1692 6.3005
R1434 VDD.n1702 VDD.n1701 6.3005
R1435 VDD.n1704 VDD.n1703 6.3005
R1436 VDD.n1707 VDD 6.3005
R1437 VDD.n1709 VDD.n1708 6.3005
R1438 VDD.n1718 VDD.n1717 6.3005
R1439 VDD.n1720 VDD.n1719 6.3005
R1440 VDD.n483 VDD.n482 6.3005
R1441 VDD.n548 VDD.n547 6.3005
R1442 VDD.n1279 VDD.n1278 6.3005
R1443 VDD.n2445 VDD.n2444 6.3005
R1444 VDD.n426 VDD.n425 6.3005
R1445 VDD.n306 VDD.n305 6.3005
R1446 VDD.n312 VDD.n307 6.3005
R1447 VDD.n321 VDD.n320 6.3005
R1448 VDD.n324 VDD.n323 6.3005
R1449 VDD.n1336 VDD.n1335 6.3005
R1450 VDD.n1342 VDD.n1338 6.3005
R1451 VDD.n1346 VDD.n1320 6.3005
R1452 VDD.n1319 VDD.n1318 6.3005
R1453 VDD.n1314 VDD.n1313 6.3005
R1454 VDD.n361 VDD.n360 6.3005
R1455 VDD.n1069 VDD.n1068 6.3005
R1456 VDD.n1062 VDD.n1061 6.3005
R1457 VDD.n1056 VDD.n1055 6.3005
R1458 VDD.n1053 VDD.n1052 6.3005
R1459 VDD.n1058 VDD.n1057 6.3005
R1460 VDD.n1060 VDD.n1059 6.3005
R1461 VDD.n864 VDD.n863 6.3005
R1462 VDD.n861 VDD.n860 6.3005
R1463 VDD.n839 VDD.n838 6.3005
R1464 VDD VDD.n830 6.3005
R1465 VDD.n837 VDD.n836 6.3005
R1466 VDD.n829 VDD.n828 6.3005
R1467 VDD.n823 VDD.n822 6.3005
R1468 VDD VDD.n819 6.3005
R1469 VDD.n818 VDD.n817 6.3005
R1470 VDD.n813 VDD.n603 6.3005
R1471 VDD.n809 VDD.n607 6.3005
R1472 VDD.n806 VDD.n610 6.3005
R1473 VDD VDD.n611 6.3005
R1474 VDD.n725 VDD.n724 6.3005
R1475 VDD.n768 VDD.n767 6.3005
R1476 VDD.n771 VDD.n770 6.3005
R1477 VDD.n715 VDD.n714 6.3005
R1478 VDD.n735 VDD.n734 6.3005
R1479 VDD.n738 VDD.n737 6.3005
R1480 VDD.n748 VDD.n747 6.3005
R1481 VDD.n775 VDD.n749 6.3005
R1482 VDD.n784 VDD.n783 6.3005
R1483 VDD.n781 VDD.n780 6.3005
R1484 VDD.n671 VDD.n635 6.3005
R1485 VDD.n669 VDD.n668 6.3005
R1486 VDD.n667 VDD.n666 6.3005
R1487 VDD.n665 VDD.n664 6.3005
R1488 VDD.n663 VDD.n662 6.3005
R1489 VDD.n658 VDD.n628 6.3005
R1490 VDD VDD.n626 6.3005
R1491 VDD.n790 VDD.n620 6.3005
R1492 VDD.n804 VDD.n613 6.3005
R1493 VDD.n799 VDD.n794 6.3005
R1494 VDD.n793 VDD.n587 6.3005
R1495 VDD.n876 VDD.n875 6.3005
R1496 VDD.n878 VDD.n877 6.3005
R1497 VDD.n1025 VDD.n1024 6.3005
R1498 VDD.n1047 VDD.n1046 6.3005
R1499 VDD.n1045 VDD.n1044 6.3005
R1500 VDD.n1051 VDD 6.3005
R1501 VDD.n1040 VDD.n1039 6.3005
R1502 VDD VDD.n1037 6.3005
R1503 VDD.n1035 VDD.n1034 6.3005
R1504 VDD.n1036 VDD.n1035 6.3005
R1505 VDD VDD.n377 6.3005
R1506 VDD.n377 VDD.n376 6.3005
R1507 VDD.n1030 VDD.n1029 6.3005
R1508 VDD.n1018 VDD.n1017 6.3005
R1509 VDD.n1019 VDD.n1013 6.3005
R1510 VDD.n1020 VDD.n1012 6.3005
R1511 VDD.n1021 VDD.n1009 6.3005
R1512 VDD.n1022 VDD.n1003 6.3005
R1513 VDD.n1000 VDD.n999 6.3005
R1514 VDD.n83 VDD.n82 6.3005
R1515 VDD VDD.n22 6.3005
R1516 VDD.n2469 VDD.n29 6.3005
R1517 VDD.n2465 VDD.n37 6.3005
R1518 VDD.n2461 VDD.n2460 6.3005
R1519 VDD.n2458 VDD.n51 6.3005
R1520 VDD.n2457 VDD 6.3005
R1521 VDD.n2456 VDD.n56 6.3005
R1522 VDD.n2454 VDD.n67 6.3005
R1523 VDD.n2453 VDD 6.3005
R1524 VDD.n2452 VDD.n2451 6.3005
R1525 VDD.n2442 VDD.n2441 6.3005
R1526 VDD.n2437 VDD.n116 6.3005
R1527 VDD.n2434 VDD.n123 6.3005
R1528 VDD.n159 VDD.n158 6.3005
R1529 VDD.n2427 VDD.n2426 6.3005
R1530 VDD.n167 VDD.n166 6.3005
R1531 VDD.n2395 VDD.n2394 6.3005
R1532 VDD.n2409 VDD 6.3005
R1533 VDD VDD.n2405 6.3005
R1534 VDD.n2410 VDD.n2387 6.3005
R1535 VDD.n2411 VDD.n2383 6.3005
R1536 VDD.n2412 VDD.n2379 6.3005
R1537 VDD.n2413 VDD.n2378 6.3005
R1538 VDD.n2414 VDD.n2375 6.3005
R1539 VDD.n2415 VDD.n2369 6.3005
R1540 VDD.n2419 VDD.n2418 6.3005
R1541 VDD.n2418 VDD.n2417 6.3005
R1542 VDD.n2423 VDD.n2422 6.3005
R1543 VDD.n2424 VDD.n2423 6.3005
R1544 VDD.n1300 VDD.n1299 6.3005
R1545 VDD.n1311 VDD.n1310 6.3005
R1546 VDD.n1306 VDD.n1079 6.3005
R1547 VDD VDD.n1087 6.3005
R1548 VDD.n1288 VDD.n1090 6.3005
R1549 VDD.n1284 VDD.n1098 6.3005
R1550 VDD VDD.n1106 6.3005
R1551 VDD.n1258 VDD.n1257 6.3005
R1552 VDD VDD.n1264 6.3005
R1553 VDD.n1263 VDD 6.3005
R1554 VDD.n1250 VDD.n1114 6.3005
R1555 VDD.n1251 VDD.n1249 6.3005
R1556 VDD.n1252 VDD.n1242 6.3005
R1557 VDD.n1253 VDD.n1241 6.3005
R1558 VDD.n1254 VDD.n1238 6.3005
R1559 VDD.n1255 VDD.n1232 6.3005
R1560 VDD.n1222 VDD.n1131 6.3005
R1561 VDD.n1131 VDD.n1130 6.3005
R1562 VDD.n1229 VDD.n1228 6.3005
R1563 VDD.n1228 VDD.n1227 6.3005
R1564 VDD.n1205 VDD.n1204 6.3005
R1565 VDD VDD.n1193 6.3005
R1566 VDD.n1210 VDD.n1185 6.3005
R1567 VDD.n1214 VDD.n1177 6.3005
R1568 VDD VDD.n1174 6.3005
R1569 VDD.n1173 VDD.n1172 6.3005
R1570 VDD.n1165 VDD.n1164 6.3005
R1571 VDD.n1168 VDD.n1167 6.3005
R1572 VDD.n1352 VDD.n1351 6.3005
R1573 VDD.n244 VDD.n243 6.3005
R1574 VDD.n1355 VDD.n231 6.3005
R1575 VDD.n1359 VDD.n216 6.3005
R1576 VDD.n1362 VDD.n205 6.3005
R1577 VDD.n1363 VDD.n204 6.3005
R1578 VDD.n1361 VDD 6.3005
R1579 VDD.n1360 VDD.n212 6.3005
R1580 VDD.n1358 VDD.n220 6.3005
R1581 VDD.n1357 VDD.n221 6.3005
R1582 VDD.n1356 VDD.n223 6.3005
R1583 VDD.n1367 VDD.n1365 6.3005
R1584 VDD VDD.n530 6.3005
R1585 VDD.n529 VDD 6.3005
R1586 VDD.n552 VDD.n528 6.3005
R1587 VDD.n554 VDD.n525 6.3005
R1588 VDD.n556 VDD.n522 6.3005
R1589 VDD.n557 VDD.n521 6.3005
R1590 VDD.n559 VDD.n519 6.3005
R1591 VDD.n561 VDD.n514 6.3005
R1592 VDD.n564 VDD.n505 6.3005
R1593 VDD.n574 VDD.n573 6.3005
R1594 VDD VDD.n471 6.3005
R1595 VDD.n488 VDD.n463 6.3005
R1596 VDD.n492 VDD.n455 6.3005
R1597 VDD VDD.n452 6.3005
R1598 VDD.n580 VDD.n444 6.3005
R1599 VDD.n584 VDD.n436 6.3005
R1600 VDD.n998 VDD 6.3005
R1601 VDD.n1383 VDD.n1382 6.3005
R1602 VDD.n2311 VDD.n1384 6.3005
R1603 VDD.n2306 VDD.n1390 6.3005
R1604 VDD.n2304 VDD.n1391 6.3005
R1605 VDD.n2300 VDD.n1400 6.3005
R1606 VDD.n2296 VDD.n1404 6.3005
R1607 VDD.n2294 VDD.n1405 6.3005
R1608 VDD.n2290 VDD.n1414 6.3005
R1609 VDD.n2286 VDD.n2284 6.3005
R1610 VDD.n2283 VDD.n1418 6.3005
R1611 VDD.n2282 VDD.n1430 6.3005
R1612 VDD.n2281 VDD.n1437 6.3005
R1613 VDD.n2280 VDD.n1439 6.3005
R1614 VDD.n2279 VDD.n2278 6.3005
R1615 VDD.n2275 VDD.n2274 6.3005
R1616 VDD.n2267 VDD.n2266 6.3005
R1617 VDD.n2232 VDD.n2231 6.3005
R1618 VDD.n1474 VDD.n1473 6.3005
R1619 VDD.n2234 VDD.n2233 6.3005
R1620 VDD.n2265 VDD.n2264 6.3005
R1621 VDD.n2269 VDD.n2268 6.3005
R1622 VDD.n2271 VDD.n2270 6.3005
R1623 VDD.n2273 VDD.n2272 6.3005
R1624 VDD.n2229 VDD.n2228 6.3005
R1625 VDD.n2227 VDD.n2226 6.3005
R1626 VDD VDD.n1870 6.3005
R1627 VDD.n1877 VDD.n1876 6.3005
R1628 VDD.n1879 VDD.n1878 6.3005
R1629 VDD.n1869 VDD.n1868 6.3005
R1630 VDD.n1863 VDD.n1862 6.3005
R1631 VDD VDD.n1859 6.3005
R1632 VDD.n1858 VDD.n1857 6.3005
R1633 VDD.n1853 VDD.n1820 6.3005
R1634 VDD.n1849 VDD.n1824 6.3005
R1635 VDD.n1846 VDD.n1827 6.3005
R1636 VDD VDD.n1828 6.3005
R1637 VDD.n1844 VDD.n1830 6.3005
R1638 VDD.n1840 VDD.n1835 6.3005
R1639 VDD.n1834 VDD.n1804 6.3005
R1640 VDD.n1884 VDD.n1883 6.3005
R1641 VDD.n2055 VDD.n2054 6.3005
R1642 VDD.n2066 VDD.n2065 6.3005
R1643 VDD.n2068 VDD.n2067 6.3005
R1644 VDD.n2075 VDD.n2074 6.3005
R1645 VDD.n2077 VDD.n2076 6.3005
R1646 VDD.n2085 VDD.n2084 6.3005
R1647 VDD.n2087 VDD.n2086 6.3005
R1648 VDD.n2098 VDD.n2097 6.3005
R1649 VDD.n2100 VDD.n2099 6.3005
R1650 VDD.n2106 VDD.n2105 6.3005
R1651 VDD.n2108 VDD.n2107 6.3005
R1652 VDD.n2116 VDD.n2115 6.3005
R1653 VDD.n2118 VDD.n2117 6.3005
R1654 VDD.n2129 VDD.n2128 6.3005
R1655 VDD.n2131 VDD.n2130 6.3005
R1656 VDD.n2136 VDD.n1996 6.3005
R1657 VDD.n2139 VDD.n1993 6.3005
R1658 VDD.n2144 VDD.n1957 6.3005
R1659 VDD.n1956 VDD.n1955 6.3005
R1660 VDD.n2142 VDD.n1963 6.3005
R1661 VDD.n2141 VDD.n1964 6.3005
R1662 VDD.n2138 VDD.n1994 6.3005
R1663 VDD.n2137 VDD.n1995 6.3005
R1664 VDD.n2134 VDD.n2002 6.3005
R1665 VDD.n2147 VDD.n2146 6.3005
R1666 VDD.n2152 VDD.n1937 6.3005
R1667 VDD.n2168 VDD.n1777 6.3005
R1668 VDD.n2167 VDD.n2166 6.3005
R1669 VDD VDD.n1782 6.3005
R1670 VDD.n2162 VDD.n1786 6.3005
R1671 VDD.n2158 VDD.n1790 6.3005
R1672 VDD.n1923 VDD.n1922 6.3005
R1673 VDD.n1921 VDD.n1920 6.3005
R1674 VDD.n1912 VDD.n1911 6.3005
R1675 VDD.n1906 VDD.n1905 6.3005
R1676 VDD.n1910 VDD 6.3005
R1677 VDD.n1904 VDD.n1903 6.3005
R1678 VDD.n1895 VDD.n1894 6.3005
R1679 VDD.n2172 VDD.n2171 6.3005
R1680 VDD.n2173 VDD.n2172 6.3005
R1681 VDD.n2169 VDD 6.3005
R1682 VDD.n2192 VDD.n1729 6.3005
R1683 VDD.n1758 VDD.n1733 6.3005
R1684 VDD.n1755 VDD.n1736 6.3005
R1685 VDD VDD.n1737 6.3005
R1686 VDD.n1753 VDD.n1739 6.3005
R1687 VDD.n1749 VDD.n1744 6.3005
R1688 VDD.n1743 VDD.n1501 6.3005
R1689 VDD.n2217 VDD.n2216 6.3005
R1690 VDD VDD.n2208 6.3005
R1691 VDD.n2215 VDD.n2214 6.3005
R1692 VDD.n2207 VDD.n2206 6.3005
R1693 VDD VDD.n2197 6.3005
R1694 VDD.n2201 VDD.n2200 6.3005
R1695 VDD.n2196 VDD.n2195 6.3005
R1696 VDD.n1723 VDD.n1722 6.3005
R1697 VDD.n1547 VDD 6.3005
R1698 VDD.n1546 VDD.n1545 6.3005
R1699 VDD.n1548 VDD.n1535 6.3005
R1700 VDD.n1550 VDD.n1549 6.3005
R1701 VDD VDD.n1527 6.3005
R1702 VDD.n1553 VDD.n1526 6.3005
R1703 VDD.n1681 VDD.n1680 6.3005
R1704 VDD.n1678 VDD.n1677 6.3005
R1705 VDD.n1687 VDD.n1686 6.3005
R1706 VDD VDD.n1688 6.3005
R1707 VDD.n1605 VDD.n1567 6.3005
R1708 VDD VDD.n1648 6.3005
R1709 VDD.n1655 VDD.n1654 6.3005
R1710 VDD.n1657 VDD.n1656 6.3005
R1711 VDD.n1647 VDD.n1646 6.3005
R1712 VDD.n1641 VDD.n1640 6.3005
R1713 VDD VDD.n1637 6.3005
R1714 VDD.n1636 VDD.n1635 6.3005
R1715 VDD.n2474 VDD.n15 6.3005
R1716 VDD.n2479 VDD.n2 6.3005
R1717 VDD.n178 VDD.n168 6.24711
R1718 VDD.n551 VDD.n550 6.01865
R1719 VDD.n1282 VDD.n1281 6.01865
R1720 VDD.n364 VDD.n363 6.01865
R1721 VDD.n728 VDD.n727 6.01865
R1722 VDD.n1028 VDD.n1027 6.01865
R1723 VDD.n1208 VDD.n1207 6.01865
R1724 VDD.n238 VDD.n237 6.01865
R1725 VDD.n486 VDD.n485 6.01863
R1726 VDD.n2448 VDD.n2447 6.01863
R1727 VDD.n315 VDD.n314 6.01863
R1728 VDD.n787 VDD.n786 6.01863
R1729 VDD.n86 VDD.n85 6.01863
R1730 VDD.n2398 VDD.n2397 6.01863
R1731 VDD.n1261 VDD.n1260 6.01863
R1732 VDD.n1684 VDD.n1683 6.01863
R1733 VDD.n14 VDD.t1188 5.62158
R1734 VDD.n0 VDD.t27 5.62158
R1735 VDD.n28 VDD.t1182 5.62158
R1736 VDD.n8 VDD.t2126 5.56425
R1737 VDD.n21 VDD.t2112 5.56425
R1738 VDD.n35 VDD.t2131 5.56425
R1739 VDD.n505 VDD.t961 5.49501
R1740 VDD.t1219 VDD.n123 5.39424
R1741 VDD.t1556 VDD.n306 5.39424
R1742 VDD.t1500 VDD.n1319 5.39424
R1743 VDD.t1554 VDD.n748 5.39424
R1744 VDD.n714 VDD.t1581 5.39424
R1745 VDD.t1533 VDD.n620 5.39424
R1746 VDD.n1031 VDD.n376 5.39424
R1747 VDD.n1046 VDD.t1281 5.39424
R1748 VDD.n2452 VDD.t1289 5.39424
R1749 VDD.n139 VDD.n138 5.22436
R1750 VDD.n681 VDD.n680 5.22436
R1751 VDD.n405 VDD.n401 5.22436
R1752 VDD.n174 VDD.n170 5.22436
R1753 VDD.n1137 VDD.n1133 5.22436
R1754 VDD.n266 VDD.n265 5.22436
R1755 VDD.n502 VDD.n498 5.22436
R1756 VDD.n346 VDD.n345 5.20342
R1757 VDD.n756 VDD.n755 5.20342
R1758 VDD.n700 VDD.n699 5.20342
R1759 VDD.n1006 VDD.t2210 5.20342
R1760 VDD.n1074 VDD.t535 5.20342
R1761 VDD.n1093 VDD.t426 5.20342
R1762 VDD.n1180 VDD.t149 5.20342
R1763 VDD.n1154 VDD.t1692 5.20342
R1764 VDD.n228 VDD.n227 5.20342
R1765 VDD.n517 VDD.t198 5.20342
R1766 VDD.n1572 VDD.t2349 5.20242
R1767 VDD.n154 VDD.n152 5.20242
R1768 VDD.n286 VDD.n284 5.20242
R1769 VDD.n1327 VDD.n1325 5.20242
R1770 VDD.n652 VDD.n650 5.20242
R1771 VDD.n62 VDD.t1035 5.20242
R1772 VDD.n43 VDD.t177 5.20242
R1773 VDD.n114 VDD.n112 5.20242
R1774 VDD.n2372 VDD.t693 5.20242
R1775 VDD.n1235 VDD.t677 5.20242
R1776 VDD.n458 VDD.t159 5.20242
R1777 VDD.n439 VDD.t859 5.20242
R1778 VDD.n1801 VDD.t2350 5.20242
R1779 VDD.n1672 VDD.t826 5.20242
R1780 VDD.n1568 VDD.t979 5.17246
R1781 VDD.n585 VDD.t82 5.17246
R1782 VDD.n165 VDD.n164 5.17246
R1783 VDD.n281 VDD.n280 5.17246
R1784 VDD.n1341 VDD.n1340 5.17246
R1785 VDD.n1066 VDD.n1064 5.17246
R1786 VDD.n879 VDD.t2078 5.17246
R1787 VDD.n760 VDD.n758 5.17246
R1788 VDD.n695 VDD.n693 5.17246
R1789 VDD.n647 VDD.n646 5.17246
R1790 VDD.n392 VDD.t632 5.17246
R1791 VDD.n52 VDD.t577 5.17246
R1792 VDD.n40 VDD.t547 5.17246
R1793 VDD.n119 VDD.n118 5.17246
R1794 VDD.n2367 VDD.t72 5.17246
R1795 VDD.n1071 VDD.t101 5.17246
R1796 VDD.n1089 VDD.t948 5.17246
R1797 VDD.n1121 VDD.t183 5.17246
R1798 VDD.n1176 VDD.t488 5.17246
R1799 VDD.n1156 VDD.t1031 5.17246
R1800 VDD.n257 VDD.n255 5.17246
R1801 VDD.n513 VDD.t2328 5.17246
R1802 VDD.n454 VDD.t722 5.17246
R1803 VDD.n1803 VDD.t191 5.17246
R1804 VDD.n1669 VDD.t440 5.17246
R1805 VDD.n859 VDD.n858 5.155
R1806 VDD.n2053 VDD.n2052 5.155
R1807 VDD.n480 VDD.n479 5.107
R1808 VDD.n543 VDD.n542 5.107
R1809 VDD.n1276 VDD.n1275 5.107
R1810 VDD.n107 VDD.t569 5.107
R1811 VDD.n424 VDD.n423 5.107
R1812 VDD.n1334 VDD.t338 5.107
R1813 VDD.n319 VDD.t1067 5.107
R1814 VDD.n359 VDD.t711 5.107
R1815 VDD.n723 VDD.t465 5.107
R1816 VDD.n766 VDD.t470 5.107
R1817 VDD.n634 VDD.t1080 5.107
R1818 VDD.n391 VDD.n390 5.107
R1819 VDD.n81 VDD.n80 5.107
R1820 VDD.n149 VDD.t447 5.107
R1821 VDD.n2393 VDD.n2392 5.107
R1822 VDD.n1298 VDD.n1297 5.107
R1823 VDD.n1120 VDD.n1119 5.107
R1824 VDD.n1202 VDD.n1201 5.107
R1825 VDD.n1160 VDD.n1159 5.107
R1826 VDD.n242 VDD.t413 5.107
R1827 VDD.n571 VDD.n570 5.107
R1828 VDD.n1377 VDD.n1376 5.107
R1829 VDD.n1668 VDD.n1667 5.107
R1830 VDD.n1534 VDD.n1533 5.01686
R1831 VDD.n827 VDD.n826 5.01686
R1832 VDD.n1867 VDD.n1866 5.01686
R1833 VDD.n2205 VDD.n2204 5.01686
R1834 VDD.n1645 VDD.n1644 5.01686
R1835 VDD VDD.t2530 5.00492
R1836 VDD VDD.t747 5.00492
R1837 VDD VDD.t2591 5.00492
R1838 VDD VDD.t2642 5.00492
R1839 VDD VDD.t2524 5.00492
R1840 VDD.n1268 VDD.n1267 4.99544
R1841 VDD.n1781 VDD.n1780 4.97139
R1842 VDD VDD.t1156 4.94116
R1843 VDD.n278 VDD.n277 4.92985
R1844 VDD.n298 VDD.n297 4.92985
R1845 VDD.n1043 VDD.n1041 4.92985
R1846 VDD.n713 VDD.n711 4.92985
R1847 VDD.n692 VDD.n690 4.92985
R1848 VDD.n618 VDD.n617 4.92985
R1849 VDD.n1038 VDD.t1288 4.92985
R1850 VDD.n89 VDD.t1298 4.92985
R1851 VDD.n53 VDD.t1297 4.92985
R1852 VDD.n92 VDD.n91 4.92985
R1853 VDD.n122 VDD.n121 4.92985
R1854 VDD.n2406 VDD.t1882 4.92985
R1855 VDD.n1088 VDD.t1895 4.92985
R1856 VDD.n1107 VDD.t1861 4.92985
R1857 VDD.n1265 VDD.t1848 4.92985
R1858 VDD.n1194 VDD.t1880 4.92985
R1859 VDD.n1175 VDD.t1898 4.92985
R1860 VDD.n203 VDD.n201 4.92985
R1861 VDD.n1366 VDD.t1602 4.92985
R1862 VDD.n472 VDD.t1570 4.92985
R1863 VDD.n453 VDD.t1568 4.92985
R1864 VDD.n1555 VDD.t1343 4.92985
R1865 VDD.n842 VDD.t2098 4.75175
R1866 VDD.n1893 VDD.n1797 4.73288
R1867 VDD.n2466 VDD.n36 4.72058
R1868 VDD.n2463 VDD.t2103 4.71604
R1869 VDD.n1625 VDD.n1590 4.6676
R1870 VDD.n1691 VDD.n1521 4.6676
R1871 VDD.n814 VDD.n602 4.6676
R1872 VDD.n1854 VDD.n1819 4.6676
R1873 VDD.n2193 VDD.n1728 4.6676
R1874 VDD.n1721 VDD.t2618 4.65357
R1875 VDD.n840 VDD.t2638 4.65357
R1876 VDD.n1880 VDD.t757 4.65357
R1877 VDD.n2218 VDD.t2614 4.65357
R1878 VDD.n1658 VDD.t2511 4.65357
R1879 VDD.n2157 VDD.t2662 4.65233
R1880 VDD.n1621 VDD.n1594 4.65007
R1881 VDD.n1618 VDD.t2009 4.65007
R1882 VDD.n1616 VDD.n1600 4.65007
R1883 VDD.n1613 VDD.t481 4.65007
R1884 VDD.n1612 VDD.n1604 4.65007
R1885 VDD.n1609 VDD.t2499 4.65007
R1886 VDD.n1696 VDD.n1518 4.65007
R1887 VDD.n1699 VDD.t2705 4.65007
R1888 VDD.n1706 VDD.n1705 4.65007
R1889 VDD.n1711 VDD.t63 4.65007
R1890 VDD.n1712 VDD.n1515 4.65007
R1891 VDD.n1715 VDD.t2602 4.65007
R1892 VDD.n1536 VDD.t1045 4.65007
R1893 VDD.n1544 VDD.t2035 4.65007
R1894 VDD.n1540 VDD.n1539 4.65007
R1895 VDD.n1543 VDD.n1542 4.65007
R1896 VDD.n594 VDD.t800 4.65007
R1897 VDD.n835 VDD.t2028 4.65007
R1898 VDD.n831 VDD.n593 4.65007
R1899 VDD.n834 VDD.n833 4.65007
R1900 VDD.n820 VDD.n597 4.65007
R1901 VDD.n598 VDD.t609 4.65007
R1902 VDD.n815 VDD.n601 4.65007
R1903 VDD.n810 VDD.n606 4.65007
R1904 VDD.n807 VDD.t2033 4.65007
R1905 VDD.n805 VDD.n612 4.65007
R1906 VDD.n801 VDD.t917 4.65007
R1907 VDD.n800 VDD.n792 4.65007
R1908 VDD.n797 VDD.t2551 4.65007
R1909 VDD.n2308 VDD.n1387 4.65007
R1910 VDD.n2305 VDD.t2727 4.65007
R1911 VDD.n2302 VDD.n1397 4.65007
R1912 VDD.n2299 VDD.t1685 4.65007
R1913 VDD.n2298 VDD.n1401 4.65007
R1914 VDD.n2295 VDD.t1375 4.65007
R1915 VDD.n2292 VDD.n1411 4.65007
R1916 VDD.n2289 VDD.t245 4.65007
R1917 VDD.n2288 VDD.n1415 4.65007
R1918 VDD.n2285 VDD.t1972 4.65007
R1919 VDD.n1428 VDD.n1421 4.65007
R1920 VDD.n1434 VDD.t2167 4.65007
R1921 VDD.n1435 VDD.n1433 4.65007
R1922 VDD.n1438 VDD.t1333 4.65007
R1923 VDD.n1449 VDD.n1442 4.65007
R1924 VDD.n2277 VDD.t1401 4.65007
R1925 VDD.n2258 VDD.n2254 4.65007
R1926 VDD.n2259 VDD.t2410 4.65007
R1927 VDD.n2261 VDD.n2251 4.65007
R1928 VDD.n2245 VDD.t2484 4.65007
R1929 VDD.n2243 VDD.n2237 4.65007
R1930 VDD.n2242 VDD.t2093 4.65007
R1931 VDD.n2188 VDD.t37 4.65007
R1932 VDD.n1874 VDD.n1873 4.65007
R1933 VDD.n1875 VDD.t1815 4.65007
R1934 VDD.n1871 VDD.n1810 4.65007
R1935 VDD.n1811 VDD.t833 4.65007
R1936 VDD.n1860 VDD.n1814 4.65007
R1937 VDD.n1815 VDD.t11 4.65007
R1938 VDD.n1855 VDD.n1818 4.65007
R1939 VDD.n1850 VDD.n1823 4.65007
R1940 VDD.n1847 VDD.t1827 4.65007
R1941 VDD.n1845 VDD.n1829 4.65007
R1942 VDD.n1842 VDD.t1411 4.65007
R1943 VDD.n1841 VDD.n1833 4.65007
R1944 VDD.n1838 VDD.t739 4.65007
R1945 VDD.n2056 VDD.t1335 4.65007
R1946 VDD.n2071 VDD.n2041 4.65007
R1947 VDD.n2073 VDD.t2742 4.65007
R1948 VDD.n2079 VDD.n2033 4.65007
R1949 VDD.n2083 VDD.t1671 4.65007
R1950 VDD.n2082 VDD.n2081 4.65007
R1951 VDD.n2088 VDD.t1363 4.65007
R1952 VDD.n2095 VDD.n2094 4.65007
R1953 VDD.n2101 VDD.t230 4.65007
R1954 VDD.n2102 VDD.n2024 4.65007
R1955 VDD.n2104 VDD.t1962 4.65007
R1956 VDD.n2110 VDD.n2016 4.65007
R1957 VDD.n2114 VDD.t2192 4.65007
R1958 VDD.n2113 VDD.n2112 4.65007
R1959 VDD.n2119 VDD.t2459 4.65007
R1960 VDD.n2126 VDD.n2125 4.65007
R1961 VDD.n2132 VDD.t1390 4.65007
R1962 VDD.n1988 VDD.n1984 4.65007
R1963 VDD.n1989 VDD.t2429 4.65007
R1964 VDD.n1991 VDD.n1981 4.65007
R1965 VDD.n1975 VDD.t2472 4.65007
R1966 VDD.n1973 VDD.n1967 4.65007
R1967 VDD.n1972 VDD.t2077 4.65007
R1968 VDD.n1775 VDD.n1774 4.65007
R1969 VDD.n2165 VDD.t1085 4.65007
R1970 VDD.n2160 VDD.n1787 4.65007
R1971 VDD.n2161 VDD.t2538 4.65007
R1972 VDD.n2164 VDD.n1783 4.65007
R1973 VDD.n1915 VDD.n1791 4.65007
R1974 VDD.n1918 VDD.t1154 4.65007
R1975 VDD.n1908 VDD.n1907 4.65007
R1976 VDD.n1914 VDD.t2237 4.65007
R1977 VDD.n1898 VDD.n1794 4.65007
R1978 VDD.n1901 VDD.t2546 4.65007
R1979 VDD.n1891 VDD.n1889 4.65007
R1980 VDD.n2198 VDD.n1511 4.65007
R1981 VDD.n1759 VDD.n1732 4.65007
R1982 VDD.n1756 VDD.t2385 4.65007
R1983 VDD.n1754 VDD.n1738 4.65007
R1984 VDD.n1751 VDD.t2750 4.65007
R1985 VDD.n1750 VDD.n1742 4.65007
R1986 VDD.n1747 VDD.t2600 4.65007
R1987 VDD.n1508 VDD.t1802 4.65007
R1988 VDD.n2213 VDD.t2400 4.65007
R1989 VDD.n2209 VDD.n1507 4.65007
R1990 VDD.n2212 VDD.n2211 4.65007
R1991 VDD.n1552 VDD.n1528 4.65007
R1992 VDD.n1652 VDD.n1651 4.65007
R1993 VDD.n1653 VDD.t2001 4.65007
R1994 VDD.n1649 VDD.n1581 4.65007
R1995 VDD.n1582 VDD.t133 4.65007
R1996 VDD.n1638 VDD.n1585 4.65007
R1997 VDD.n1586 VDD.t118 4.65007
R1998 VDD.n1626 VDD.n1589 4.65007
R1999 VDD.n1622 VDD.t2365 4.64811
R2000 VDD.n1695 VDD.t2341 4.64811
R2001 VDD.n811 VDD.t2105 4.64811
R2002 VDD.n1851 VDD.t2147 4.64811
R2003 VDD.n1897 VDD.t1464 4.64811
R2004 VDD.n1760 VDD.t2221 4.64811
R2005 VDD.n1659 VDD.n1575 4.64487
R2006 VDD.n485 VDD.t1613 4.64447
R2007 VDD.n550 VDD.t1572 4.64447
R2008 VDD.n1281 VDD.t1890 4.64447
R2009 VDD.n2447 VDD.n102 4.64447
R2010 VDD.n428 VDD.t1213 4.64447
R2011 VDD.n271 VDD.n270 4.64447
R2012 VDD.n315 VDD.n291 4.64447
R2013 VDD.n363 VDD.n354 4.64447
R2014 VDD.n727 VDD.n718 4.64447
R2015 VDD.n685 VDD.n684 4.64447
R2016 VDD.n786 VDD.n629 4.64447
R2017 VDD.n1027 VDD.t1201 4.64447
R2018 VDD.n85 VDD.t1215 4.64447
R2019 VDD.n2429 VDD.n144 4.64447
R2020 VDD.n2397 VDD.t1903 4.64447
R2021 VDD.n1302 VDD.t1907 4.64447
R2022 VDD.n1260 VDD.t1905 4.64447
R2023 VDD.n1207 VDD.t1894 4.64447
R2024 VDD.n1140 VDD.t1909 4.64447
R2025 VDD.n238 VDD.n234 4.64447
R2026 VDD.n576 VDD.t1611 4.64447
R2027 VDD.n1683 VDD.t1345 4.64447
R2028 VDD.n310 VDD.t1139 4.61485
R2029 VDD.n293 VDD.n292 4.61485
R2030 VDD.n1344 VDD.t965 4.61485
R2031 VDD.n273 VDD.n272 4.61485
R2032 VDD.n348 VDD.t403 4.61485
R2033 VDD.n1050 VDD.n1049 4.61485
R2034 VDD.n717 VDD.n705 4.61485
R2035 VDD.n732 VDD.t545 4.61485
R2036 VDD.n687 VDD.n686 4.61485
R2037 VDD.n773 VDD.t986 4.61485
R2038 VDD.n654 VDD.t659 4.61485
R2039 VDD.n788 VDD.n627 4.61485
R2040 VDD.n385 VDD.t328 4.61485
R2041 VDD.n1011 VDD.n1010 4.61485
R2042 VDD.n87 VDD.t498 4.61485
R2043 VDD.n65 VDD.n59 4.61485
R2044 VDD.n417 VDD.t258 4.61485
R2045 VDD.n49 VDD.n48 4.61485
R2046 VDD.n2439 VDD.t1014 4.61485
R2047 VDD.n2449 VDD.n98 4.61485
R2048 VDD.n161 VDD.t379 4.61485
R2049 VDD.n2432 VDD.n129 4.61485
R2050 VDD.n2399 VDD.t783 4.61485
R2051 VDD.n2377 VDD.n2376 4.61485
R2052 VDD.n1308 VDD.n1076 4.61485
R2053 VDD.n1292 VDD.t639 4.61485
R2054 VDD.n1286 VDD.n1095 4.61485
R2055 VDD.n1270 VDD.t1704 4.61485
R2056 VDD.n1262 VDD.t135 4.61485
R2057 VDD.n1240 VDD.n1239 4.61485
R2058 VDD.n1212 VDD.n1182 4.61485
R2059 VDD.n1196 VDD.t815 4.61485
R2060 VDD.n1170 VDD.n1151 4.61485
R2061 VDD.n1218 VDD.t574 4.61485
R2062 VDD.n222 VDD.t647 4.61485
R2063 VDD.n236 VDD.n235 4.61485
R2064 VDD.n537 VDD.t592 4.61485
R2065 VDD.n558 VDD.n520 4.61485
R2066 VDD.n474 VDD.t302 4.61485
R2067 VDD.n490 VDD.n460 4.61485
R2068 VDD.n496 VDD.t1717 4.61485
R2069 VDD.n582 VDD.n441 4.61485
R2070 VDD.n1380 VDD.t211 4.61485
R2071 VDD.n1371 VDD.n1370 4.61485
R2072 VDD.n2309 VDD.t1786 4.61485
R2073 VDD.n2057 VDD.n2049 4.61485
R2074 VDD.n2063 VDD.t105 4.61485
R2075 VDD.n2062 VDD.n2061 4.61485
R2076 VDD.n2070 VDD.t1417 4.61485
R2077 VDD.n1662 VDD.t993 4.61485
R2078 VDD.n1675 VDD.n1674 4.61485
R2079 VDD.n866 VDD.t1056 4.58941
R2080 VDD.t1058 VDD.n2223 4.58941
R2081 VDD.n2221 VDD.t1062 4.58941
R2082 VDD.t1060 VDD.n2149 4.58941
R2083 VDD.n2154 VDD.t1053 4.58941
R2084 VDD.n335 VDD.n332 4.53072
R2085 VDD.n640 VDD.n637 4.53072
R2086 VDD.n395 VDD.t1752 4.53072
R2087 VDD.n2359 VDD.t2014 4.53072
R2088 VDD.n1124 VDD.t2454 4.53072
R2089 VDD.n249 VDD.n246 4.53072
R2090 VDD.n508 VDD.t956 4.53072
R2091 VDD.n136 VDD.n135 4.5005
R2092 VDD.n678 VDD.n677 4.5005
R2093 VDD.n1033 VDD.n380 4.5005
R2094 VDD.n1033 VDD.n1032 4.5005
R2095 VDD.n1032 VDD.n1031 4.5005
R2096 VDD.n404 VDD.n403 4.5005
R2097 VDD.n173 VDD.n172 4.5005
R2098 VDD.n2420 VDD.n178 4.5005
R2099 VDD.n2366 VDD.n178 4.5005
R2100 VDD.n1136 VDD.n1135 4.5005
R2101 VDD.n1129 VDD.n180 4.5005
R2102 VDD.n1226 VDD.n1129 4.5005
R2103 VDD.n263 VDD.n262 4.5005
R2104 VDD.n501 VDD.n500 4.5005
R2105 VDD.n379 VDD.n200 4.5005
R2106 VDD.n2183 VDD.n1763 4.5005
R2107 VDD.n2182 VDD.n2181 4.5005
R2108 VDD.n1887 VDD.n1886 4.5005
R2109 VDD.n2177 VDD.n1764 4.5005
R2110 VDD.n2177 VDD.n2176 4.5005
R2111 VDD.n2176 VDD.n2175 4.5005
R2112 VDD.n1798 VDD.n1767 4.5005
R2113 VDD.n2180 VDD.n2179 4.5005
R2114 VDD.n2156 VDD.n1923 4.28283
R2115 VDD.n14 VDD.t1194 4.2255
R2116 VDD.n8 VDD.t2140 4.2255
R2117 VDD.n0 VDD.t21 4.2255
R2118 VDD.n1568 VDD.t978 4.2255
R2119 VDD.n585 VDD.t81 4.2255
R2120 VDD.n165 VDD.n163 4.2255
R2121 VDD.n337 VDD.n336 4.2255
R2122 VDD.n142 VDD.n141 4.2255
R2123 VDD.n278 VDD.n276 4.2255
R2124 VDD.n281 VDD.n279 4.2255
R2125 VDD.n298 VDD.n296 4.2255
R2126 VDD.n1341 VDD.n1339 4.2255
R2127 VDD.n1066 VDD.n1065 4.2255
R2128 VDD.n1043 VDD.n1042 4.2255
R2129 VDD.n883 VDD.t2073 4.2255
R2130 VDD.n882 VDD.t2065 4.2255
R2131 VDD.n881 VDD.t2090 4.2255
R2132 VDD.n880 VDD.t2069 4.2255
R2133 VDD.n879 VDD.t2061 4.2255
R2134 VDD.t1056 VDD.n843 4.2255
R2135 VDD.n760 VDD.n759 4.2255
R2136 VDD.n713 VDD.n712 4.2255
R2137 VDD.n695 VDD.n694 4.2255
R2138 VDD.n692 VDD.n691 4.2255
R2139 VDD.n683 VDD.n674 4.2255
R2140 VDD.n641 VDD.n636 4.2255
R2141 VDD.n647 VDD.n645 4.2255
R2142 VDD.n618 VDD.n616 4.2255
R2143 VDD.n1038 VDD.t1287 4.2255
R2144 VDD.n392 VDD.t630 4.2255
R2145 VDD.n407 VDD.t2247 4.2255
R2146 VDD.n396 VDD.t203 4.2255
R2147 VDD.n89 VDD.t1206 4.2255
R2148 VDD.n52 VDD.t576 4.2255
R2149 VDD.n53 VDD.t1199 4.2255
R2150 VDD.n21 VDD.t2132 4.2255
R2151 VDD.n35 VDD.t2143 4.2255
R2152 VDD.n28 VDD.t1186 4.2255
R2153 VDD.n40 VDD.t548 4.2255
R2154 VDD.n92 VDD.n90 4.2255
R2155 VDD.n119 VDD.n117 4.2255
R2156 VDD.n122 VDD.n120 4.2255
R2157 VDD.n2406 VDD.t1923 4.2255
R2158 VDD.n2367 VDD.t70 4.2255
R2159 VDD.n2360 VDD.t1449 4.2255
R2160 VDD.n176 VDD.t623 4.2255
R2161 VDD.n1071 VDD.t103 4.2255
R2162 VDD.n1088 VDD.t1888 4.2255
R2163 VDD.n1089 VDD.t950 4.2255
R2164 VDD.n1107 VDD.t1860 4.2255
R2165 VDD.n1265 VDD.t1886 4.2255
R2166 VDD.n1121 VDD.t184 4.2255
R2167 VDD.n1125 VDD.t874 4.2255
R2168 VDD.n1139 VDD.t2448 4.2255
R2169 VDD.n1194 VDD.t1899 4.2255
R2170 VDD.n1176 VDD.t487 4.2255
R2171 VDD.n1175 VDD.t1892 4.2255
R2172 VDD.n1156 VDD.t1032 4.2255
R2173 VDD.n251 VDD.n250 4.2255
R2174 VDD.n269 VDD.n268 4.2255
R2175 VDD.n257 VDD.n256 4.2255
R2176 VDD.n203 VDD.n202 4.2255
R2177 VDD.n1366 VDD.t1508 4.2255
R2178 VDD.n513 VDD.t2326 4.2255
R2179 VDD.n504 VDD.t84 4.2255
R2180 VDD.n509 VDD.t1024 4.2255
R2181 VDD.n472 VDD.t1604 4.2255
R2182 VDD.n454 VDD.t721 4.2255
R2183 VDD.n453 VDD.t1603 4.2255
R2184 VDD.n2224 VDD.t1058 4.2255
R2185 VDD.n1500 VDD.t1062 4.2255
R2186 VDD.n1803 VDD.t192 4.2255
R2187 VDD.n2150 VDD.t1060 4.2255
R2188 VDD.t1053 VDD.n1924 4.2255
R2189 VDD.n1669 VDD.t439 4.2255
R2190 VDD.n1555 VDD.t1303 4.2255
R2191 VDD.n1690 VDD.n1689 4.12867
R2192 VDD.n851 VDD.n850 4.08391
R2193 VDD.n1482 VDD.n1481 4.08391
R2194 VDD.n1495 VDD.n1494 4.08391
R2195 VDD.n1945 VDD.n1944 4.08391
R2196 VDD.n1932 VDD.n1931 4.08391
R2197 VDD.n846 VDD.n845 4.07616
R2198 VDD.n1477 VDD.n1476 4.07616
R2199 VDD.n1490 VDD.n1489 4.07616
R2200 VDD.n1940 VDD.n1939 4.07616
R2201 VDD.n1927 VDD.n1926 4.07616
R2202 VDD.n1893 VDD.n1892 4.06552
R2203 VDD.n778 VDD.n777 3.77052
R2204 VDD.n1304 VDD.n1303 3.77052
R2205 VDD.n1220 VDD.n1219 3.77052
R2206 VDD.n1349 VDD.n1348 3.7705
R2207 VDD.n429 VDD.n418 3.7705
R2208 VDD.n578 VDD.n577 3.7705
R2209 VDD.n2431 VDD.n2430 3.7705
R2210 VDD.n335 VDD.n334 3.75093
R2211 VDD.n340 VDD.n339 3.75093
R2212 VDD.n640 VDD.n639 3.75093
R2213 VDD.n644 VDD.n643 3.75093
R2214 VDD.n395 VDD.n394 3.75093
R2215 VDD.n399 VDD.n398 3.75093
R2216 VDD.n2359 VDD.n2358 3.75093
R2217 VDD.n2363 VDD.n2362 3.75093
R2218 VDD.n1124 VDD.n1123 3.75093
R2219 VDD.n1128 VDD.n1127 3.75093
R2220 VDD.n249 VDD.n248 3.75093
R2221 VDD.n254 VDD.n253 3.75093
R2222 VDD.n508 VDD.n507 3.75093
R2223 VDD.n512 VDD.n511 3.75093
R2224 VDD VDD.n2225 3.73526
R2225 VDD VDD.n2151 3.73526
R2226 VDD.n869 VDD.n841 3.68288
R2227 VDD.n347 VDD.n346 3.60822
R2228 VDD.n757 VDD.n756 3.60822
R2229 VDD.n701 VDD.n700 3.60822
R2230 VDD.n229 VDD.n228 3.60822
R2231 VDD.n155 VDD.n154 3.60784
R2232 VDD.n287 VDD.n286 3.60784
R2233 VDD.n1328 VDD.n1327 3.60784
R2234 VDD.n653 VDD.n652 3.60784
R2235 VDD.n115 VDD.n114 3.60784
R2236 VDD.n1007 VDD.n1006 3.60762
R2237 VDD.n1075 VDD.n1074 3.60762
R2238 VDD.n1094 VDD.n1093 3.60762
R2239 VDD.n1181 VDD.n1180 3.60762
R2240 VDD.n1155 VDD.n1154 3.60762
R2241 VDD.n518 VDD.n517 3.60762
R2242 VDD.n1573 VDD.n1572 3.60724
R2243 VDD.n63 VDD.n62 3.60724
R2244 VDD.n44 VDD.n43 3.60724
R2245 VDD.n2373 VDD.n2372 3.60724
R2246 VDD.n1236 VDD.n1235 3.60724
R2247 VDD.n459 VDD.n458 3.60724
R2248 VDD.n440 VDD.n439 3.60724
R2249 VDD.n1802 VDD.n1801 3.60724
R2250 VDD.n1673 VDD.n1672 3.60724
R2251 VDD.n874 VDD.n871 3.54746
R2252 VDD.n435 VDD.n432 3.54746
R2253 VDD.n1396 VDD.n1393 3.54746
R2254 VDD.n1410 VDD.n1407 3.54746
R2255 VDD.n1426 VDD.n1423 3.54746
R2256 VDD.n1447 VDD.n1444 3.54746
R2257 VDD.n1460 VDD.n1459 3.54746
R2258 VDD.n2250 VDD.n2249 3.54746
R2259 VDD.n1466 VDD.n1465 3.54746
R2260 VDD.n2038 VDD.n2035 3.54746
R2261 VDD.n2093 VDD.n2090 3.54746
R2262 VDD.n2021 VDD.n2018 3.54746
R2263 VDD.n2124 VDD.n2121 3.54746
R2264 VDD.n2001 VDD.n2000 3.54746
R2265 VDD.n1980 VDD.n1979 3.54746
R2266 VDD.n1962 VDD.n1961 3.54746
R2267 VDD.n20 VDD.n19 3.5318
R2268 VDD.n13 VDD.n12 3.5318
R2269 VDD.n7 VDD.n6 3.5318
R2270 VDD.n1632 VDD.n1631 3.5318
R2271 VDD.n34 VDD.n33 3.5318
R2272 VDD.n27 VDD.n26 3.5318
R2273 VDD.n2176 VDD.n1771 3.49104
R2274 VDD VDD.n997 3.43071
R2275 VDD.n2263 VDD.n2245 3.4205
R2276 VDD.n2140 VDD.n1975 3.4205
R2277 VDD.n331 VDD.n330 3.30485
R2278 VDD.n303 VDD.n302 3.30485
R2279 VDD.n369 VDD.n366 3.30485
R2280 VDD.n710 VDD.n707 3.30485
R2281 VDD.n745 VDD.n742 3.30485
R2282 VDD.n625 VDD.n624 3.30485
R2283 VDD.n374 VDD.n371 3.30485
R2284 VDD.n72 VDD.n71 3.30485
R2285 VDD.n415 VDD.n414 3.30485
R2286 VDD.n97 VDD.n96 3.30485
R2287 VDD.n128 VDD.n127 3.30485
R2288 VDD.n2404 VDD.n2403 3.30485
R2289 VDD.n1086 VDD.n1083 3.30485
R2290 VDD.n1105 VDD.n1102 3.30485
R2291 VDD.n1112 VDD.n1111 3.30485
R2292 VDD.n1192 VDD.n1189 3.30485
R2293 VDD.n1148 VDD.n1145 3.30485
R2294 VDD.n210 VDD.n207 3.30485
R2295 VDD.n535 VDD.n532 3.30485
R2296 VDD.n470 VDD.n469 3.30485
R2297 VDD.n451 VDD.n450 3.30485
R2298 VDD.n1560 VDD.n1559 3.30485
R2299 VDD.n1031 VDD.t1229 3.23675
R2300 VDD.n2335 VDD.n2333 3.17341
R2301 VDD.n1224 VDD.n1223 3.1505
R2302 VDD.n1225 VDD.n1224 3.1505
R2303 VDD.n2174 VDD.n1771 3.1505
R2304 VDD.n2170 VDD.n1771 3.1505
R2305 VDD.n1886 VDD.n1885 3.10611
R2306 VDD.n1623 VDD.n1593 3.02507
R2307 VDD.n1619 VDD.n1597 3.02507
R2308 VDD.n1614 VDD.n1603 3.02507
R2309 VDD.n1610 VDD.n1608 3.02507
R2310 VDD.n1694 VDD.n1520 3.02507
R2311 VDD.n1700 VDD.n1698 3.02507
R2312 VDD.n1710 VDD.n1517 3.02507
R2313 VDD.n1716 VDD.n1714 3.02507
R2314 VDD.n1534 VDD.n1532 3.02507
R2315 VDD.n1541 VDD.n1538 3.02507
R2316 VDD.n1514 VDD.n1513 3.02507
R2317 VDD.n859 VDD.n857 3.02507
R2318 VDD.n827 VDD.n825 3.02507
R2319 VDD.n832 VDD.n592 3.02507
R2320 VDD.n590 VDD.n589 3.02507
R2321 VDD.n821 VDD.n596 3.02507
R2322 VDD.n816 VDD.n600 3.02507
R2323 VDD.n812 VDD.n605 3.02507
R2324 VDD.n808 VDD.n609 3.02507
R2325 VDD.n803 VDD.n615 3.02507
R2326 VDD.n798 VDD.n796 3.02507
R2327 VDD.n2307 VDD.n1389 3.02507
R2328 VDD.n2301 VDD.n1399 3.02507
R2329 VDD.n2297 VDD.n1403 3.02507
R2330 VDD.n2291 VDD.n1413 3.02507
R2331 VDD.n2287 VDD.n1417 3.02507
R2332 VDD.n1429 VDD.n1420 3.02507
R2333 VDD.n1436 VDD.n1432 3.02507
R2334 VDD.n1450 VDD.n1441 3.02507
R2335 VDD.n1454 VDD.n1453 3.02507
R2336 VDD.n2257 VDD.n2256 3.02507
R2337 VDD.n2260 VDD.n2253 3.02507
R2338 VDD.n2244 VDD.n2236 3.02507
R2339 VDD.n2241 VDD.n2239 3.02507
R2340 VDD.n1471 VDD.n1470 3.02507
R2341 VDD.n1807 VDD.n1806 3.02507
R2342 VDD.n1872 VDD.n1809 3.02507
R2343 VDD.n1867 VDD.n1865 3.02507
R2344 VDD.n1861 VDD.n1813 3.02507
R2345 VDD.n1856 VDD.n1817 3.02507
R2346 VDD.n1852 VDD.n1822 3.02507
R2347 VDD.n1848 VDD.n1826 3.02507
R2348 VDD.n1843 VDD.n1832 3.02507
R2349 VDD.n1839 VDD.n1837 3.02507
R2350 VDD.n2053 VDD.n2051 3.02507
R2351 VDD.n2072 VDD.n2040 3.02507
R2352 VDD.n2080 VDD.n2032 3.02507
R2353 VDD.n2030 VDD.n2029 3.02507
R2354 VDD.n2027 VDD.n2026 3.02507
R2355 VDD.n2103 VDD.n2023 3.02507
R2356 VDD.n2111 VDD.n2015 3.02507
R2357 VDD.n2013 VDD.n2012 3.02507
R2358 VDD.n2010 VDD.n2009 3.02507
R2359 VDD.n2006 VDD.n2005 3.02507
R2360 VDD.n1987 VDD.n1986 3.02507
R2361 VDD.n1990 VDD.n1983 3.02507
R2362 VDD.n1974 VDD.n1966 3.02507
R2363 VDD.n1971 VDD.n1969 3.02507
R2364 VDD.n1953 VDD.n1952 3.02507
R2365 VDD.n1776 VDD.n1773 3.02507
R2366 VDD.n1781 VDD.n1779 3.02507
R2367 VDD.n2159 VDD.n1789 3.02507
R2368 VDD.n2163 VDD.n1785 3.02507
R2369 VDD.n1919 VDD.n1917 3.02507
R2370 VDD.n1913 VDD.n1793 3.02507
R2371 VDD.n1902 VDD.n1900 3.02507
R2372 VDD.n1896 VDD.n1796 3.02507
R2373 VDD.n1770 VDD.n1769 3.02507
R2374 VDD.n2199 VDD.n1510 3.02507
R2375 VDD.n1727 VDD.n1726 3.02507
R2376 VDD.n2191 VDD.n1731 3.02507
R2377 VDD.n1757 VDD.n1735 3.02507
R2378 VDD.n1752 VDD.n1741 3.02507
R2379 VDD.n1748 VDD.n1746 3.02507
R2380 VDD.n2205 VDD.n2203 3.02507
R2381 VDD.n2210 VDD.n1506 3.02507
R2382 VDD.n1504 VDD.n1503 3.02507
R2383 VDD.n1551 VDD.n1530 3.02507
R2384 VDD.n1525 VDD.n1524 3.02507
R2385 VDD.n1578 VDD.n1577 3.02507
R2386 VDD.n1650 VDD.n1580 3.02507
R2387 VDD.n1645 VDD.n1643 3.02507
R2388 VDD.n1639 VDD.n1584 3.02507
R2389 VDD.n1627 VDD.n1588 3.02507
R2390 VDD.n997 VDD.n996 2.99957
R2391 VDD.n484 VDD.n476 2.98985
R2392 VDD.n480 VDD.n478 2.98985
R2393 VDD.n543 VDD.n541 2.98985
R2394 VDD.n549 VDD.n539 2.98985
R2395 VDD.n1276 VDD.n1274 2.98985
R2396 VDD.n1280 VDD.n1272 2.98985
R2397 VDD.n107 VDD.n106 2.98985
R2398 VDD.n2446 VDD.n104 2.98985
R2399 VDD.n427 VDD.n420 2.98985
R2400 VDD.n424 VDD.n422 2.98985
R2401 VDD.n1334 VDD.n1333 2.98985
R2402 VDD.n1331 VDD.n1330 2.98985
R2403 VDD.n319 VDD.n318 2.98985
R2404 VDD.n316 VDD.n290 2.98985
R2405 VDD.n311 VDD.n309 2.98985
R2406 VDD.n313 VDD.n295 2.98985
R2407 VDD.n1345 VDD.n1322 2.98985
R2408 VDD.n1347 VDD.n275 2.98985
R2409 VDD.n1054 VDD.n353 2.98985
R2410 VDD.n351 VDD.n350 2.98985
R2411 VDD.n362 VDD.n356 2.98985
R2412 VDD.n359 VDD.n358 2.98985
R2413 VDD.n726 VDD.n720 2.98985
R2414 VDD.n723 VDD.n722 2.98985
R2415 VDD.n763 VDD.n762 2.98985
R2416 VDD.n766 VDD.n765 2.98985
R2417 VDD.n729 VDD.n704 2.98985
R2418 VDD.n733 VDD.n731 2.98985
R2419 VDD.n776 VDD.n689 2.98985
R2420 VDD.n774 VDD.n751 2.98985
R2421 VDD.n634 VDD.n633 2.98985
R2422 VDD.n785 VDD.n631 2.98985
R2423 VDD.n657 VDD.n656 2.98985
R2424 VDD.n661 VDD.n660 2.98985
R2425 VDD.n391 VDD.n389 2.98985
R2426 VDD.n1026 VDD.n387 2.98985
R2427 VDD.n1016 VDD.n1015 2.98985
R2428 VDD.n383 VDD.n382 2.98985
R2429 VDD.n84 VDD.n77 2.98985
R2430 VDD.n81 VDD.n79 2.98985
R2431 VDD.n75 VDD.n74 2.98985
R2432 VDD.n66 VDD.n58 2.98985
R2433 VDD.n410 VDD.n409 2.98985
R2434 VDD.n50 VDD.n47 2.98985
R2435 VDD.n2440 VDD.n109 2.98985
R2436 VDD.n101 VDD.n100 2.98985
R2437 VDD.n160 VDD.n157 2.98985
R2438 VDD.n132 VDD.n131 2.98985
R2439 VDD.n149 VDD.n148 2.98985
R2440 VDD.n2428 VDD.n146 2.98985
R2441 VDD.n2396 VDD.n2389 2.98985
R2442 VDD.n2393 VDD.n2391 2.98985
R2443 VDD.n2386 VDD.n2385 2.98985
R2444 VDD.n2382 VDD.n2381 2.98985
R2445 VDD.n1298 VDD.n1296 2.98985
R2446 VDD.n1301 VDD.n1294 2.98985
R2447 VDD.n1307 VDD.n1078 2.98985
R2448 VDD.n1305 VDD.n1081 2.98985
R2449 VDD.n1285 VDD.n1097 2.98985
R2450 VDD.n1283 VDD.n1100 2.98985
R2451 VDD.n1259 VDD.n1116 2.98985
R2452 VDD.n1120 VDD.n1118 2.98985
R2453 VDD.n1248 VDD.n1247 2.98985
R2454 VDD.n1245 VDD.n1244 2.98985
R2455 VDD.n1202 VDD.n1200 2.98985
R2456 VDD.n1206 VDD.n1198 2.98985
R2457 VDD.n1211 VDD.n1184 2.98985
R2458 VDD.n1209 VDD.n1187 2.98985
R2459 VDD.n1171 VDD.n1150 2.98985
R2460 VDD.n1143 VDD.n1142 2.98985
R2461 VDD.n1160 VDD.n1158 2.98985
R2462 VDD.n1163 VDD.n1162 2.98985
R2463 VDD.n215 VDD.n214 2.98985
R2464 VDD.n219 VDD.n218 2.98985
R2465 VDD.n239 VDD.n233 2.98985
R2466 VDD.n242 VDD.n241 2.98985
R2467 VDD.n555 VDD.n524 2.98985
R2468 VDD.n553 VDD.n527 2.98985
R2469 VDD.n575 VDD.n567 2.98985
R2470 VDD.n571 VDD.n569 2.98985
R2471 VDD.n487 VDD.n465 2.98985
R2472 VDD.n489 VDD.n462 2.98985
R2473 VDD.n579 VDD.n446 2.98985
R2474 VDD.n581 VDD.n443 2.98985
R2475 VDD.n1377 VDD.n1375 2.98985
R2476 VDD.n1381 VDD.n1379 2.98985
R2477 VDD.n2312 VDD.n1373 2.98985
R2478 VDD.n2310 VDD.n1386 2.98985
R2479 VDD.n2058 VDD.n2048 2.98985
R2480 VDD.n2064 VDD.n2060 2.98985
R2481 VDD.n2046 VDD.n2045 2.98985
R2482 VDD.n2069 VDD.n2043 2.98985
R2483 VDD.n1682 VDD.n1664 2.98985
R2484 VDD.n1668 VDD.n1666 2.98985
R2485 VDD.n1685 VDD.n1566 2.98985
R2486 VDD.n1564 VDD.n1563 2.98985
R2487 VDD.n2464 VDD.n39 2.95711
R2488 VDD.n996 VDD.n995 2.94069
R2489 VDD.n868 VDD.n842 2.91309
R2490 VDD.n1572 VDD.t2337 2.84673
R2491 VDD.n154 VDD.n153 2.84673
R2492 VDD.n286 VDD.n285 2.84673
R2493 VDD.n1327 VDD.n1326 2.84673
R2494 VDD.n652 VDD.n651 2.84673
R2495 VDD.n62 VDD.t1034 2.84673
R2496 VDD.n43 VDD.t174 2.84673
R2497 VDD.n114 VDD.n113 2.84673
R2498 VDD.n2372 VDD.t689 2.84673
R2499 VDD.n1235 VDD.t673 2.84673
R2500 VDD.n458 VDD.t162 2.84673
R2501 VDD.n439 VDD.t860 2.84673
R2502 VDD.n1801 VDD.t2339 2.84673
R2503 VDD.n1672 VDD.t824 2.84673
R2504 VDD.n346 VDD.n344 2.84631
R2505 VDD.n756 VDD.n754 2.84631
R2506 VDD.n700 VDD.n698 2.84631
R2507 VDD.n1006 VDD.t2214 2.84631
R2508 VDD.n1074 VDD.t540 2.84631
R2509 VDD.n1093 VDD.t430 2.84631
R2510 VDD.n1180 VDD.t150 2.84631
R2511 VDD.n1154 VDD.t1697 2.84631
R2512 VDD.n228 VDD.n226 2.84631
R2513 VDD.n517 VDD.t196 2.84631
R2514 VDD.n868 VDD.n867 2.82929
R2515 VDD.n2262 VDD.n2261 2.63697
R2516 VDD.n1992 VDD.n1991 2.63697
R2517 VDD VDD.n165 2.61227
R2518 VDD VDD.n1341 2.61227
R2519 VDD VDD.n760 2.61227
R2520 VDD VDD.n1071 2.61227
R2521 VDD VDD.n1156 2.61227
R2522 VDD VDD.n1669 2.61227
R2523 VDD.n999 VDD.t1751 2.6092
R2524 VDD.n2365 VDD.t2015 2.6092
R2525 VDD.n1225 VDD.t2453 2.6092
R2526 VDD.n20 VDD.n17 2.6005
R2527 VDD.n13 VDD.n10 2.6005
R2528 VDD.n7 VDD.n4 2.6005
R2529 VDD.n1632 VDD.n1629 2.6005
R2530 VDD.n331 VDD.n328 2.6005
R2531 VDD.n303 VDD.n300 2.6005
R2532 VDD.n369 VDD.n368 2.6005
R2533 VDD.n874 VDD.n873 2.6005
R2534 VDD.n710 VDD.n709 2.6005
R2535 VDD.n745 VDD.n744 2.6005
R2536 VDD.n625 VDD.n622 2.6005
R2537 VDD.n374 VDD.n373 2.6005
R2538 VDD.n72 VDD.n69 2.6005
R2539 VDD.n415 VDD.n412 2.6005
R2540 VDD.n34 VDD.n31 2.6005
R2541 VDD.n27 VDD.n24 2.6005
R2542 VDD.n97 VDD.n94 2.6005
R2543 VDD.n128 VDD.n125 2.6005
R2544 VDD.n2404 VDD.n2401 2.6005
R2545 VDD.n1086 VDD.n1085 2.6005
R2546 VDD.n1105 VDD.n1104 2.6005
R2547 VDD.n1112 VDD.n1109 2.6005
R2548 VDD.n1192 VDD.n1191 2.6005
R2549 VDD.n1148 VDD.n1147 2.6005
R2550 VDD.n210 VDD.n209 2.6005
R2551 VDD.n535 VDD.n534 2.6005
R2552 VDD.n470 VDD.n467 2.6005
R2553 VDD.n451 VDD.n448 2.6005
R2554 VDD.n435 VDD.n434 2.6005
R2555 VDD.n1396 VDD.n1395 2.6005
R2556 VDD.n1410 VDD.n1409 2.6005
R2557 VDD.n1426 VDD.n1425 2.6005
R2558 VDD.n1447 VDD.n1446 2.6005
R2559 VDD.n1460 VDD.n1457 2.6005
R2560 VDD.n2250 VDD.n2247 2.6005
R2561 VDD.n1466 VDD.n1463 2.6005
R2562 VDD.n2038 VDD.n2037 2.6005
R2563 VDD.n2093 VDD.n2092 2.6005
R2564 VDD.n2021 VDD.n2020 2.6005
R2565 VDD.n2124 VDD.n2123 2.6005
R2566 VDD.n2001 VDD.n1998 2.6005
R2567 VDD.n1980 VDD.n1977 2.6005
R2568 VDD.n1962 VDD.n1959 2.6005
R2569 VDD.n1560 VDD.n1557 2.6005
R2570 VDD.n140 VDD.n133 2.58689
R2571 VDD.n682 VDD.n675 2.58689
R2572 VDD.n406 VDD.n400 2.58689
R2573 VDD.n175 VDD.n169 2.58689
R2574 VDD.n1138 VDD.n1132 2.58689
R2575 VDD.n267 VDD.n260 2.58689
R2576 VDD.n503 VDD.n497 2.58689
R2577 VDD.n855 VDD.n854 2.57852
R2578 VDD.n1486 VDD.n1485 2.57852
R2579 VDD.n1499 VDD.n1498 2.57852
R2580 VDD.n1949 VDD.n1948 2.57852
R2581 VDD.n1936 VDD.n1935 2.57852
R2582 VDD.n2243 VDD.n2242 2.44638
R2583 VDD.n1973 VDD.n1972 2.44638
R2584 VDD.n854 VDD.n852 2.39186
R2585 VDD.n1485 VDD.n1483 2.39186
R2586 VDD.n1498 VDD.n1496 2.39186
R2587 VDD.n1948 VDD.n1946 2.39186
R2588 VDD.n1935 VDD.n1933 2.39186
R2589 VDD.n892 VDD.n888 2.36621
R2590 VDD.n2333 VDD.n190 2.36511
R2591 VDD.n586 VDD.n585 2.32427
R2592 VDD.n984 VDD.n982 2.31745
R2593 VDD.n1035 VDD.n377 2.31316
R2594 VDD.n981 VDD.n190 2.30648
R2595 VDD.n2242 VDD.n2241 2.28756
R2596 VDD.n2244 VDD.n2243 2.28756
R2597 VDD.n2245 VDD.n2244 2.28756
R2598 VDD.n2261 VDD.n2260 2.28756
R2599 VDD.n2260 VDD.n2259 2.28756
R2600 VDD.n2258 VDD.n2257 2.28756
R2601 VDD.n1972 VDD.n1971 2.28756
R2602 VDD.n1974 VDD.n1973 2.28756
R2603 VDD.n1975 VDD.n1974 2.28756
R2604 VDD.n1991 VDD.n1990 2.28756
R2605 VDD.n1990 VDD.n1989 2.28756
R2606 VDD.n1988 VDD.n1987 2.28756
R2607 VDD.n969 VDD.n885 2.28191
R2608 VDD.n2157 VDD.n2156 2.28105
R2609 VDD.n1892 VDD.n1891 2.273
R2610 VDD.n997 VDD.n884 2.25729
R2611 VDD.n379 VDD.n378 2.25698
R2612 VDD.n2319 VDD.n2318 2.25213
R2613 VDD.n962 VDD.n961 2.25213
R2614 VDD.n893 VDD.n892 2.25213
R2615 VDD.n915 VDD.n914 2.25213
R2616 VDD.n2334 VDD.n187 2.25213
R2617 VDD.n975 VDD.n974 2.25213
R2618 VDD.n2323 VDD.n198 2.25176
R2619 VDD.n951 VDD.n948 2.25176
R2620 VDD.n904 VDD.n903 2.25176
R2621 VDD.n921 VDD.n918 2.25176
R2622 VDD.n2347 VDD.n2346 2.25176
R2623 VDD.n981 VDD.n978 2.25176
R2624 VDD.n1881 VDD.n1880 2.25151
R2625 VDD.n2219 VDD.n2218 2.2515
R2626 VDD.n2346 VDD.n2345 2.25144
R2627 VDD.n2186 VDD.n2185 2.25142
R2628 VDD.n384 VDD.n380 2.25122
R2629 VDD.n2323 VDD.n2322 2.25107
R2630 VDD.n1349 VDD.n271 2.25102
R2631 VDD.n778 VDD.n685 2.25102
R2632 VDD.n429 VDD.n428 2.25102
R2633 VDD.n2430 VDD.n2429 2.25102
R2634 VDD.n1303 VDD.n1302 2.25102
R2635 VDD.n1220 VDD.n1140 2.25102
R2636 VDD.n577 VDD.n576 2.25102
R2637 VDD.n986 VDD.n971 2.25088
R2638 VDD.n2330 VDD.n2329 2.2505
R2639 VDD.n2324 VDD.n199 2.2505
R2640 VDD.n197 VDD.n195 2.2505
R2641 VDD.n2328 VDD.n196 2.2505
R2642 VDD.n2327 VDD.n2326 2.2505
R2643 VDD.n958 VDD.n941 2.2505
R2644 VDD.n953 VDD.n952 2.2505
R2645 VDD.n959 VDD.n937 2.2505
R2646 VDD.n960 VDD.n959 2.2505
R2647 VDD.n949 VDD.n942 2.2505
R2648 VDD.n950 VDD.n946 2.2505
R2649 VDD.n898 VDD.n891 2.2505
R2650 VDD.n905 VDD.n901 2.2505
R2651 VDD.n897 VDD.n896 2.2505
R2652 VDD.n907 VDD.n899 2.2505
R2653 VDD.n891 VDD.n886 2.2505
R2654 VDD.n906 VDD.n900 2.2505
R2655 VDD.n933 VDD.n932 2.2505
R2656 VDD.n934 VDD.n916 2.2505
R2657 VDD.n931 VDD.n917 2.2505
R2658 VDD.n930 VDD.n929 2.2505
R2659 VDD.n2341 VDD.n186 2.2505
R2660 VDD.n2348 VDD.n2344 2.2505
R2661 VDD.n2339 VDD.n2338 2.2505
R2662 VDD.n2340 VDD.n2339 2.2505
R2663 VDD.n2350 VDD.n2342 2.2505
R2664 VDD.n2349 VDD.n2343 2.2505
R2665 VDD.n2338 VDD.n2337 2.2505
R2666 VDD.n2335 VDD.n2334 2.2505
R2667 VDD.n184 VDD.n182 2.2505
R2668 VDD.n186 VDD.n184 2.2505
R2669 VDD.n2336 VDD.n189 2.2505
R2670 VDD.n189 VDD.n188 2.2505
R2671 VDD.n921 VDD.n179 2.2505
R2672 VDD.n922 VDD.n919 2.2505
R2673 VDD.n924 VDD.n922 2.2505
R2674 VDD.n936 VDD.n935 2.2505
R2675 VDD.n935 VDD.n934 2.2505
R2676 VDD.n914 VDD.n910 2.2505
R2677 VDD.n923 VDD.n920 2.2505
R2678 VDD.n920 VDD.n917 2.2505
R2679 VDD.n933 VDD.n912 2.2505
R2680 VDD.n925 VDD.n912 2.2505
R2681 VDD.n926 VDD.n911 2.2505
R2682 VDD.n913 VDD.n911 2.2505
R2683 VDD.n929 VDD.n928 2.2505
R2684 VDD.n928 VDD.n927 2.2505
R2685 VDD.n2344 VDD.n183 2.2505
R2686 VDD.n2352 VDD.n2351 2.2505
R2687 VDD.n2351 VDD.n2350 2.2505
R2688 VDD.n2349 VDD.n185 2.2505
R2689 VDD.n2345 VDD.n185 2.2505
R2690 VDD.n992 VDD.n991 2.2505
R2691 VDD.n982 VDD.n979 2.2505
R2692 VDD.n993 VDD.n976 2.2505
R2693 VDD.n990 VDD.n977 2.2505
R2694 VDD.n989 VDD.n988 2.2505
R2695 VDD.n995 VDD.n994 2.2505
R2696 VDD.n994 VDD.n993 2.2505
R2697 VDD.n974 VDD.n970 2.2505
R2698 VDD.n983 VDD.n980 2.2505
R2699 VDD.n980 VDD.n977 2.2505
R2700 VDD.n985 VDD.n972 2.2505
R2701 VDD.n992 VDD.n972 2.2505
R2702 VDD.n973 VDD.n971 2.2505
R2703 VDD.n988 VDD.n987 2.2505
R2704 VDD.n987 VDD.n986 2.2505
R2705 VDD.n968 VDD.n886 2.2505
R2706 VDD.n903 VDD.n902 2.2505
R2707 VDD.n894 VDD.n885 2.2505
R2708 VDD.n906 VDD.n890 2.2505
R2709 VDD.n890 VDD.n887 2.2505
R2710 VDD.n901 VDD.n889 2.2505
R2711 VDD.n895 VDD.n888 2.2505
R2712 VDD.n896 VDD.n895 2.2505
R2713 VDD.n909 VDD.n908 2.2505
R2714 VDD.n908 VDD.n907 2.2505
R2715 VDD.n964 VDD.n937 2.2505
R2716 VDD.n953 VDD.n944 2.2505
R2717 VDD.n963 VDD.n962 2.2505
R2718 VDD.n943 VDD.n938 2.2505
R2719 VDD.n943 VDD.n942 2.2505
R2720 VDD.n957 VDD.n956 2.2505
R2721 VDD.n958 VDD.n957 2.2505
R2722 VDD.n948 VDD.n947 2.2505
R2723 VDD.n945 VDD.n939 2.2505
R2724 VDD.n940 VDD.n939 2.2505
R2725 VDD.n954 VDD.n946 2.2505
R2726 VDD.n955 VDD.n954 2.2505
R2727 VDD.n2318 VDD.n2317 2.2505
R2728 VDD.n2324 VDD.n191 2.2505
R2729 VDD.n2315 VDD.n193 2.2505
R2730 VDD.n195 VDD.n193 2.2505
R2731 VDD.n2316 VDD.n194 2.2505
R2732 VDD.n196 VDD.n194 2.2505
R2733 VDD.n2332 VDD.n2331 2.2505
R2734 VDD.n2331 VDD.n2330 2.2505
R2735 VDD.n2322 VDD.n2321 2.2505
R2736 VDD.n2321 VDD.n2320 2.2505
R2737 VDD.n2326 VDD.n2325 2.2505
R2738 VDD.n2325 VDD.n192 2.2505
R2739 VDD.n1762 VDD.n1761 2.2505
R2740 VDD.n2179 VDD.n2178 2.2505
R2741 VDD.n1890 VDD.n1888 2.2505
R2742 VDD.n1659 VDD.n1658 2.2505
R2743 VDD.n1575 VDD.n1568 2.21762
R2744 VDD.n2220 VDD.n2219 2.15367
R2745 VDD.n2156 VDD.n2155 2.12779
R2746 VDD.n2421 VDD.n168 2.1005
R2747 VDD.n2365 VDD.n168 2.1005
R2748 VDD.n1882 VDD.n1803 2.03935
R2749 VDD.n965 VDD.n936 1.96654
R2750 VDD.n2259 VDD.n2258 1.94874
R2751 VDD.n1989 VDD.n1988 1.94874
R2752 VDD.n1882 VDD.n1881 1.91888
R2753 VDD.n325 VDD.n281 1.88267
R2754 VDD.n1067 VDD.n1066 1.88267
R2755 VDD.n739 VDD.n695 1.88267
R2756 VDD.n672 VDD.n647 1.88267
R2757 VDD.n1002 VDD.n392 1.88267
R2758 VDD.n55 VDD.n52 1.88267
R2759 VDD.n2462 VDD.n40 1.88267
R2760 VDD.n2436 VDD.n119 1.88267
R2761 VDD.n2368 VDD.n2367 1.88267
R2762 VDD.n1289 VDD.n1089 1.88267
R2763 VDD.n1231 VDD.n1121 1.88267
R2764 VDD.n1215 VDD.n1176 1.88267
R2765 VDD.n258 VDD.n257 1.88267
R2766 VDD.n562 VDD.n513 1.88267
R2767 VDD.n493 VDD.n454 1.88267
R2768 VDD.n2355 VDD.n2354 1.80258
R2769 VDD.n966 VDD.n965 1.79408
R2770 VDD.n1313 VDD.t913 1.73963
R2771 VDD.n781 VDD.t1470 1.73963
R2772 VDD.n1352 VDD.t2710 1.73963
R2773 VDD.n1354 VDD.n245 1.65613
R2774 VDD.n17 VDD.t2116 1.6255
R2775 VDD.n17 VDD.n16 1.6255
R2776 VDD.n19 VDD.t2134 1.6255
R2777 VDD.n19 VDD.n18 1.6255
R2778 VDD.n10 VDD.t1195 1.6255
R2779 VDD.n10 VDD.n9 1.6255
R2780 VDD.n12 VDD.t1190 1.6255
R2781 VDD.n12 VDD.n11 1.6255
R2782 VDD.n4 VDD.t2135 1.6255
R2783 VDD.n4 VDD.n3 1.6255
R2784 VDD.n6 VDD.t2121 1.6255
R2785 VDD.n6 VDD.n5 1.6255
R2786 VDD.n1629 VDD.t28 1.6255
R2787 VDD.n1629 VDD.n1628 1.6255
R2788 VDD.n1631 VDD.t23 1.6255
R2789 VDD.n1631 VDD.n1630 1.6255
R2790 VDD.n1571 VDD.t2348 1.6255
R2791 VDD.n1571 VDD.n1570 1.6255
R2792 VDD.n1593 VDD.t2360 1.6255
R2793 VDD.n1593 VDD.n1592 1.6255
R2794 VDD.n1597 VDD.t1997 1.6255
R2795 VDD.n1597 VDD.n1596 1.6255
R2796 VDD.n1603 VDD.t483 1.6255
R2797 VDD.n1603 VDD.n1602 1.6255
R2798 VDD.n1608 VDD.t2506 1.6255
R2799 VDD.n1608 VDD.n1607 1.6255
R2800 VDD.n1520 VDD.t2333 1.6255
R2801 VDD.n1520 VDD.n1519 1.6255
R2802 VDD.n1698 VDD.t2700 1.6255
R2803 VDD.n1698 VDD.n1697 1.6255
R2804 VDD.n1517 VDD.t55 1.6255
R2805 VDD.n1517 VDD.n1516 1.6255
R2806 VDD.n1714 VDD.t2630 1.6255
R2807 VDD.n1714 VDD.n1713 1.6255
R2808 VDD.n1532 VDD.t1047 1.6255
R2809 VDD.n1532 VDD.n1531 1.6255
R2810 VDD.n1538 VDD.t2707 1.6255
R2811 VDD.n1538 VDD.n1537 1.6255
R2812 VDD.n1513 VDD.t2610 1.6255
R2813 VDD.n1513 VDD.n1512 1.6255
R2814 VDD.n476 VDD.t2625 1.6255
R2815 VDD.n476 VDD.n475 1.6255
R2816 VDD.n478 VDD.t1175 1.6255
R2817 VDD.n478 VDD.n477 1.6255
R2818 VDD.n541 VDD.t333 1.6255
R2819 VDD.n541 VDD.n540 1.6255
R2820 VDD.n539 VDD.t2476 1.6255
R2821 VDD.n539 VDD.n538 1.6255
R2822 VDD.n1274 VDD.t143 1.6255
R2823 VDD.n1274 VDD.n1273 1.6255
R2824 VDD.n1272 VDD.t2640 1.6255
R2825 VDD.n1272 VDD.n1271 1.6255
R2826 VDD.n151 VDD.t516 1.6255
R2827 VDD.n151 VDD.n150 1.6255
R2828 VDD.n106 VDD.t2598 1.6255
R2829 VDD.n106 VDD.n105 1.6255
R2830 VDD.n104 VDD.t1278 1.6255
R2831 VDD.n104 VDD.n103 1.6255
R2832 VDD.n420 VDD.t1329 1.6255
R2833 VDD.n420 VDD.n419 1.6255
R2834 VDD.n422 VDD.t1125 1.6255
R2835 VDD.n422 VDD.n421 1.6255
R2836 VDD.n334 VDD.t911 1.6255
R2837 VDD.n334 VDD.n333 1.6255
R2838 VDD.n339 VDD.t885 1.6255
R2839 VDD.n339 VDD.n338 1.6255
R2840 VDD.n328 VDD.t1548 1.6255
R2841 VDD.n328 VDD.n327 1.6255
R2842 VDD.n330 VDD.t1501 1.6255
R2843 VDD.n330 VDD.n329 1.6255
R2844 VDD.n1333 VDD.t1365 1.6255
R2845 VDD.n1333 VDD.n1332 1.6255
R2846 VDD.n1330 VDD.t1493 1.6255
R2847 VDD.n1330 VDD.n1329 1.6255
R2848 VDD.n318 VDD.t2651 1.6255
R2849 VDD.n318 VDD.n317 1.6255
R2850 VDD.n290 VDD.t1506 1.6255
R2851 VDD.n290 VDD.n289 1.6255
R2852 VDD.n283 VDD.t523 1.6255
R2853 VDD.n283 VDD.n282 1.6255
R2854 VDD.n309 VDD.t226 1.6255
R2855 VDD.n309 VDD.n308 1.6255
R2856 VDD.n295 VDD.t1436 1.6255
R2857 VDD.n295 VDD.n294 1.6255
R2858 VDD.n300 VDD.t1593 1.6255
R2859 VDD.n300 VDD.n299 1.6255
R2860 VDD.n302 VDD.t1557 1.6255
R2861 VDD.n302 VDD.n301 1.6255
R2862 VDD.n1324 VDD.t974 1.6255
R2863 VDD.n1324 VDD.n1323 1.6255
R2864 VDD.n1322 VDD.t315 1.6255
R2865 VDD.n1322 VDD.n1321 1.6255
R2866 VDD.n275 VDD.t599 1.6255
R2867 VDD.n275 VDD.n274 1.6255
R2868 VDD.n343 VDD.t354 1.6255
R2869 VDD.n343 VDD.n342 1.6255
R2870 VDD.n353 VDD.t561 1.6255
R2871 VDD.n353 VDD.n352 1.6255
R2872 VDD.n350 VDD.t931 1.6255
R2873 VDD.n350 VDD.n349 1.6255
R2874 VDD.n368 VDD.t1282 1.6255
R2875 VDD.n368 VDD.n367 1.6255
R2876 VDD.n366 VDD.t1285 1.6255
R2877 VDD.n366 VDD.n365 1.6255
R2878 VDD.n356 VDD.t1232 1.6255
R2879 VDD.n356 VDD.n355 1.6255
R2880 VDD.n358 VDD.t1936 1.6255
R2881 VDD.n358 VDD.n357 1.6255
R2882 VDD.n873 VDD.t1674 1.6255
R2883 VDD.n873 VDD.n872 1.6255
R2884 VDD.n871 VDD.t1665 1.6255
R2885 VDD.n871 VDD.n870 1.6255
R2886 VDD.n845 VDD.t1756 1.6255
R2887 VDD.n845 VDD.n844 1.6255
R2888 VDD.n854 VDD.t1760 1.6255
R2889 VDD.n854 VDD.n853 1.6255
R2890 VDD.n850 VDD.t1757 1.6255
R2891 VDD.n850 VDD.n849 1.6255
R2892 VDD.n848 VDD.t1759 1.6255
R2893 VDD.n848 VDD.n847 1.6255
R2894 VDD.n857 VDD.t2110 1.6255
R2895 VDD.n857 VDD.n856 1.6255
R2896 VDD.n825 VDD.t802 1.6255
R2897 VDD.n825 VDD.n824 1.6255
R2898 VDD.n592 VDD.t2026 1.6255
R2899 VDD.n592 VDD.n591 1.6255
R2900 VDD.n589 VDD.t2623 1.6255
R2901 VDD.n589 VDD.n588 1.6255
R2902 VDD.n596 VDD.t2616 1.6255
R2903 VDD.n596 VDD.n595 1.6255
R2904 VDD.n600 VDD.t614 1.6255
R2905 VDD.n600 VDD.n599 1.6255
R2906 VDD.n605 VDD.t2054 1.6255
R2907 VDD.n605 VDD.n604 1.6255
R2908 VDD.n609 VDD.t2021 1.6255
R2909 VDD.n609 VDD.n608 1.6255
R2910 VDD.n615 VDD.t915 1.6255
R2911 VDD.n615 VDD.n614 1.6255
R2912 VDD.n720 VDD.t1632 1.6255
R2913 VDD.n720 VDD.n719 1.6255
R2914 VDD.n722 VDD.t2667 1.6255
R2915 VDD.n722 VDD.n721 1.6255
R2916 VDD.n762 VDD.t1606 1.6255
R2917 VDD.n762 VDD.n761 1.6255
R2918 VDD.n765 VDD.t2283 1.6255
R2919 VDD.n765 VDD.n764 1.6255
R2920 VDD.n753 VDD.t850 1.6255
R2921 VDD.n753 VDD.n752 1.6255
R2922 VDD.n709 VDD.t1609 1.6255
R2923 VDD.n709 VDD.n708 1.6255
R2924 VDD.n707 VDD.t1582 1.6255
R2925 VDD.n707 VDD.n706 1.6255
R2926 VDD.n704 VDD.t584 1.6255
R2927 VDD.n704 VDD.n703 1.6255
R2928 VDD.n731 VDD.t2298 1.6255
R2929 VDD.n731 VDD.n730 1.6255
R2930 VDD.n697 VDD.t1099 1.6255
R2931 VDD.n697 VDD.n696 1.6255
R2932 VDD.n744 VDD.t1623 1.6255
R2933 VDD.n744 VDD.n743 1.6255
R2934 VDD.n742 VDD.t1555 1.6255
R2935 VDD.n742 VDD.n741 1.6255
R2936 VDD.n689 VDD.t307 1.6255
R2937 VDD.n689 VDD.n688 1.6255
R2938 VDD.n751 VDD.t724 1.6255
R2939 VDD.n751 VDD.n750 1.6255
R2940 VDD.n633 VDD.t2261 1.6255
R2941 VDD.n633 VDD.n632 1.6255
R2942 VDD.n631 VDD.t1510 1.6255
R2943 VDD.n631 VDD.n630 1.6255
R2944 VDD.n639 VDD.t1473 1.6255
R2945 VDD.n639 VDD.n638 1.6255
R2946 VDD.n643 VDD.t2317 1.6255
R2947 VDD.n643 VDD.n642 1.6255
R2948 VDD.n649 VDD.t389 1.6255
R2949 VDD.n649 VDD.n648 1.6255
R2950 VDD.n656 VDD.t4 1.6255
R2951 VDD.n656 VDD.n655 1.6255
R2952 VDD.n660 VDD.t1762 1.6255
R2953 VDD.n660 VDD.n659 1.6255
R2954 VDD.n622 VDD.t1583 1.6255
R2955 VDD.n622 VDD.n621 1.6255
R2956 VDD.n624 VDD.t1534 1.6255
R2957 VDD.n624 VDD.n623 1.6255
R2958 VDD.n796 VDD.t2681 1.6255
R2959 VDD.n796 VDD.n795 1.6255
R2960 VDD.n389 VDD.t1131 1.6255
R2961 VDD.n389 VDD.n388 1.6255
R2962 VDD.n387 VDD.t1305 1.6255
R2963 VDD.n387 VDD.n386 1.6255
R2964 VDD.n373 VDD.t1230 1.6255
R2965 VDD.n373 VDD.n372 1.6255
R2966 VDD.n371 VDD.t1244 1.6255
R2967 VDD.n371 VDD.n370 1.6255
R2968 VDD.n1015 VDD.t2207 1.6255
R2969 VDD.n1015 VDD.n1014 1.6255
R2970 VDD.n382 VDD.t2252 1.6255
R2971 VDD.n382 VDD.n381 1.6255
R2972 VDD.n1005 VDD.t2208 1.6255
R2973 VDD.n1005 VDD.n1004 1.6255
R2974 VDD.n394 VDD.t209 1.6255
R2975 VDD.n394 VDD.n393 1.6255
R2976 VDD.n398 VDD.t208 1.6255
R2977 VDD.n398 VDD.n397 1.6255
R2978 VDD.n77 VDD.t2556 1.6255
R2979 VDD.n77 VDD.n76 1.6255
R2980 VDD.n79 VDD.t397 1.6255
R2981 VDD.n79 VDD.n78 1.6255
R2982 VDD.n69 VDD.t1225 1.6255
R2983 VDD.n69 VDD.n68 1.6255
R2984 VDD.n71 VDD.t1265 1.6255
R2985 VDD.n71 VDD.n70 1.6255
R2986 VDD.n74 VDD.t2612 1.6255
R2987 VDD.n74 VDD.n73 1.6255
R2988 VDD.n58 VDD.t506 1.6255
R2989 VDD.n58 VDD.n57 1.6255
R2990 VDD.n61 VDD.t1036 1.6255
R2991 VDD.n61 VDD.n60 1.6255
R2992 VDD.n412 VDD.t1211 1.6255
R2993 VDD.n412 VDD.n411 1.6255
R2994 VDD.n414 VDD.t1264 1.6255
R2995 VDD.n414 VDD.n413 1.6255
R2996 VDD.n409 VDD.t273 1.6255
R2997 VDD.n409 VDD.n408 1.6255
R2998 VDD.n47 VDD.t170 1.6255
R2999 VDD.n47 VDD.n46 1.6255
R3000 VDD.n31 VDD.t2133 1.6255
R3001 VDD.n31 VDD.n30 1.6255
R3002 VDD.n33 VDD.t2114 1.6255
R3003 VDD.n33 VDD.n32 1.6255
R3004 VDD.n24 VDD.t1183 1.6255
R3005 VDD.n24 VDD.n23 1.6255
R3006 VDD.n26 VDD.t1177 1.6255
R3007 VDD.n26 VDD.n25 1.6255
R3008 VDD.n39 VDD.t788 1.6255
R3009 VDD.n39 VDD.n38 1.6255
R3010 VDD.n42 VDD.t172 1.6255
R3011 VDD.n42 VDD.n41 1.6255
R3012 VDD.n94 VDD.t1299 1.6255
R3013 VDD.n94 VDD.n93 1.6255
R3014 VDD.n96 VDD.t1290 1.6255
R3015 VDD.n96 VDD.n95 1.6255
R3016 VDD.n109 VDD.t2089 1.6255
R3017 VDD.n109 VDD.n108 1.6255
R3018 VDD.n100 VDD.t1103 1.6255
R3019 VDD.n100 VDD.n99 1.6255
R3020 VDD.n111 VDD.t284 1.6255
R3021 VDD.n111 VDD.n110 1.6255
R3022 VDD.n125 VDD.t1220 1.6255
R3023 VDD.n125 VDD.n124 1.6255
R3024 VDD.n127 VDD.t1271 1.6255
R3025 VDD.n127 VDD.n126 1.6255
R3026 VDD.n157 VDD.t701 1.6255
R3027 VDD.n157 VDD.n156 1.6255
R3028 VDD.n131 VDD.t374 1.6255
R3029 VDD.n131 VDD.n130 1.6255
R3030 VDD.n148 VDD.t1948 1.6255
R3031 VDD.n148 VDD.n147 1.6255
R3032 VDD.n146 VDD.t1276 1.6255
R3033 VDD.n146 VDD.n145 1.6255
R3034 VDD.n2389 VDD.t1958 1.6255
R3035 VDD.n2389 VDD.n2388 1.6255
R3036 VDD.n2391 VDD.t323 1.6255
R3037 VDD.n2391 VDD.n2390 1.6255
R3038 VDD.n2401 VDD.t1858 1.6255
R3039 VDD.n2401 VDD.n2400 1.6255
R3040 VDD.n2403 VDD.t1925 1.6255
R3041 VDD.n2403 VDD.n2402 1.6255
R3042 VDD.n2385 VDD.t625 1.6255
R3043 VDD.n2385 VDD.n2384 1.6255
R3044 VDD.n2381 VDD.t684 1.6255
R3045 VDD.n2381 VDD.n2380 1.6255
R3046 VDD.n2371 VDD.t694 1.6255
R3047 VDD.n2371 VDD.n2370 1.6255
R3048 VDD.n2358 VDD.t1455 1.6255
R3049 VDD.n2358 VDD.n2357 1.6255
R3050 VDD.n2362 VDD.t1454 1.6255
R3051 VDD.n2362 VDD.n2361 1.6255
R3052 VDD.n1296 VDD.t1699 1.6255
R3053 VDD.n1296 VDD.n1295 1.6255
R3054 VDD.n1294 VDD.t1960 1.6255
R3055 VDD.n1294 VDD.n1293 1.6255
R3056 VDD.n1073 VDD.t536 1.6255
R3057 VDD.n1073 VDD.n1072 1.6255
R3058 VDD.n1078 VDD.t186 1.6255
R3059 VDD.n1078 VDD.n1077 1.6255
R3060 VDD.n1081 VDD.t553 1.6255
R3061 VDD.n1081 VDD.n1080 1.6255
R3062 VDD.n1085 VDD.t1915 1.6255
R3063 VDD.n1085 VDD.n1084 1.6255
R3064 VDD.n1083 VDD.t1916 1.6255
R3065 VDD.n1083 VDD.n1082 1.6255
R3066 VDD.n1092 VDD.t424 1.6255
R3067 VDD.n1092 VDD.n1091 1.6255
R3068 VDD.n1097 VDD.t1709 1.6255
R3069 VDD.n1097 VDD.n1096 1.6255
R3070 VDD.n1100 VDD.t2190 1.6255
R3071 VDD.n1100 VDD.n1099 1.6255
R3072 VDD.n1104 VDD.t1919 1.6255
R3073 VDD.n1104 VDD.n1103 1.6255
R3074 VDD.n1102 VDD.t1922 1.6255
R3075 VDD.n1102 VDD.n1101 1.6255
R3076 VDD.n1116 VDD.t2723 1.6255
R3077 VDD.n1116 VDD.n1115 1.6255
R3078 VDD.n1118 VDD.t292 1.6255
R3079 VDD.n1118 VDD.n1117 1.6255
R3080 VDD.n1109 VDD.t1926 1.6255
R3081 VDD.n1109 VDD.n1108 1.6255
R3082 VDD.n1111 VDD.t1913 1.6255
R3083 VDD.n1111 VDD.n1110 1.6255
R3084 VDD.n1247 VDD.t2447 1.6255
R3085 VDD.n1247 VDD.n1246 1.6255
R3086 VDD.n1244 VDD.t706 1.6255
R3087 VDD.n1244 VDD.n1243 1.6255
R3088 VDD.n1234 VDD.t671 1.6255
R3089 VDD.n1234 VDD.n1233 1.6255
R3090 VDD.n1123 VDD.t875 1.6255
R3091 VDD.n1123 VDD.n1122 1.6255
R3092 VDD.n1127 VDD.t872 1.6255
R3093 VDD.n1127 VDD.n1126 1.6255
R3094 VDD.n1200 VDD.t1748 1.6255
R3095 VDD.n1200 VDD.n1199 1.6255
R3096 VDD.n1198 VDD.t2649 1.6255
R3097 VDD.n1198 VDD.n1197 1.6255
R3098 VDD.n1191 VDD.t1921 1.6255
R3099 VDD.n1191 VDD.n1190 1.6255
R3100 VDD.n1189 VDD.t1924 1.6255
R3101 VDD.n1189 VDD.n1188 1.6255
R3102 VDD.n1184 VDD.t120 1.6255
R3103 VDD.n1184 VDD.n1183 1.6255
R3104 VDD.n1187 VDD.t1683 1.6255
R3105 VDD.n1187 VDD.n1186 1.6255
R3106 VDD.n1179 VDD.t148 1.6255
R3107 VDD.n1179 VDD.n1178 1.6255
R3108 VDD.n1147 VDD.t1838 1.6255
R3109 VDD.n1147 VDD.n1146 1.6255
R3110 VDD.n1145 VDD.t1917 1.6255
R3111 VDD.n1145 VDD.n1144 1.6255
R3112 VDD.n1153 VDD.t1696 1.6255
R3113 VDD.n1153 VDD.n1152 1.6255
R3114 VDD.n1150 VDD.t1687 1.6255
R3115 VDD.n1150 VDD.n1149 1.6255
R3116 VDD.n1142 VDD.t841 1.6255
R3117 VDD.n1142 VDD.n1141 1.6255
R3118 VDD.n1158 VDD.t1646 1.6255
R3119 VDD.n1158 VDD.n1157 1.6255
R3120 VDD.n1162 VDD.t2725 1.6255
R3121 VDD.n1162 VDD.n1161 1.6255
R3122 VDD.n248 VDD.t2713 1.6255
R3123 VDD.n248 VDD.n247 1.6255
R3124 VDD.n253 VDD.t1784 1.6255
R3125 VDD.n253 VDD.n252 1.6255
R3126 VDD.n225 VDD.t346 1.6255
R3127 VDD.n225 VDD.n224 1.6255
R3128 VDD.n214 VDD.t2383 1.6255
R3129 VDD.n214 VDD.n213 1.6255
R3130 VDD.n218 VDD.t2019 1.6255
R3131 VDD.n218 VDD.n217 1.6255
R3132 VDD.n209 VDD.t1634 1.6255
R3133 VDD.n209 VDD.n208 1.6255
R3134 VDD.n207 VDD.t1590 1.6255
R3135 VDD.n207 VDD.n206 1.6255
R3136 VDD.n233 VDD.t1625 1.6255
R3137 VDD.n233 VDD.n232 1.6255
R3138 VDD.n241 VDD.t1356 1.6255
R3139 VDD.n241 VDD.n240 1.6255
R3140 VDD.n534 VDD.t1585 1.6255
R3141 VDD.n534 VDD.n533 1.6255
R3142 VDD.n532 VDD.t1518 1.6255
R3143 VDD.n532 VDD.n531 1.6255
R3144 VDD.n524 VDD.t594 1.6255
R3145 VDD.n524 VDD.n523 1.6255
R3146 VDD.n527 VDD.t86 1.6255
R3147 VDD.n527 VDD.n526 1.6255
R3148 VDD.n516 VDD.t194 1.6255
R3149 VDD.n516 VDD.n515 1.6255
R3150 VDD.n507 VDD.t1026 1.6255
R3151 VDD.n507 VDD.n506 1.6255
R3152 VDD.n511 VDD.t1019 1.6255
R3153 VDD.n511 VDD.n510 1.6255
R3154 VDD.n567 VDD.t2488 1.6255
R3155 VDD.n567 VDD.n566 1.6255
R3156 VDD.n569 VDD.t432 1.6255
R3157 VDD.n569 VDD.n568 1.6255
R3158 VDD.n467 VDD.t1527 1.6255
R3159 VDD.n467 VDD.n466 1.6255
R3160 VDD.n469 VDD.t1488 1.6255
R3161 VDD.n469 VDD.n468 1.6255
R3162 VDD.n465 VDD.t2440 1.6255
R3163 VDD.n465 VDD.n464 1.6255
R3164 VDD.n462 VDD.t155 1.6255
R3165 VDD.n462 VDD.n461 1.6255
R3166 VDD.n457 VDD.t161 1.6255
R3167 VDD.n457 VDD.n456 1.6255
R3168 VDD.n448 VDD.t1526 1.6255
R3169 VDD.n448 VDD.n447 1.6255
R3170 VDD.n450 VDD.t1486 1.6255
R3171 VDD.n450 VDD.n449 1.6255
R3172 VDD.n446 VDD.t652 1.6255
R3173 VDD.n446 VDD.n445 1.6255
R3174 VDD.n443 VDD.t654 1.6255
R3175 VDD.n443 VDD.n442 1.6255
R3176 VDD.n438 VDD.t858 1.6255
R3177 VDD.n438 VDD.n437 1.6255
R3178 VDD.n434 VDD.t2181 1.6255
R3179 VDD.n434 VDD.n433 1.6255
R3180 VDD.n432 VDD.t2177 1.6255
R3181 VDD.n432 VDD.n431 1.6255
R3182 VDD.n1375 VDD.t219 1.6255
R3183 VDD.n1375 VDD.n1374 1.6255
R3184 VDD.n1379 VDD.t2405 1.6255
R3185 VDD.n1379 VDD.n1378 1.6255
R3186 VDD.n1373 VDD.t679 1.6255
R3187 VDD.n1373 VDD.n1372 1.6255
R3188 VDD.n1386 VDD.t870 1.6255
R3189 VDD.n1386 VDD.n1385 1.6255
R3190 VDD.n1389 VDD.t2737 1.6255
R3191 VDD.n1389 VDD.n1388 1.6255
R3192 VDD.n1395 VDD.t670 1.6255
R3193 VDD.n1395 VDD.n1394 1.6255
R3194 VDD.n1393 VDD.t1669 1.6255
R3195 VDD.n1393 VDD.n1392 1.6255
R3196 VDD.n1399 VDD.t1655 1.6255
R3197 VDD.n1399 VDD.n1398 1.6255
R3198 VDD.n1403 VDD.t1358 1.6255
R3199 VDD.n1403 VDD.n1402 1.6255
R3200 VDD.n1409 VDD.t820 1.6255
R3201 VDD.n1409 VDD.n1408 1.6255
R3202 VDD.n1407 VDD.t241 1.6255
R3203 VDD.n1407 VDD.n1406 1.6255
R3204 VDD.n1413 VDD.t256 1.6255
R3205 VDD.n1413 VDD.n1412 1.6255
R3206 VDD.n1417 VDD.t1977 1.6255
R3207 VDD.n1417 VDD.n1416 1.6255
R3208 VDD.n1425 VDD.t266 1.6255
R3209 VDD.n1425 VDD.n1424 1.6255
R3210 VDD.n1423 VDD.t2188 1.6255
R3211 VDD.n1423 VDD.n1422 1.6255
R3212 VDD.n1420 VDD.t2180 1.6255
R3213 VDD.n1420 VDD.n1419 1.6255
R3214 VDD.n1432 VDD.t1340 1.6255
R3215 VDD.n1432 VDD.n1431 1.6255
R3216 VDD.n1446 VDD.t807 1.6255
R3217 VDD.n1446 VDD.n1445 1.6255
R3218 VDD.n1444 VDD.t1396 1.6255
R3219 VDD.n1444 VDD.n1443 1.6255
R3220 VDD.n1441 VDD.t1392 1.6255
R3221 VDD.n1441 VDD.n1440 1.6255
R3222 VDD.n1453 VDD.t2296 1.6255
R3223 VDD.n1453 VDD.n1452 1.6255
R3224 VDD.n1457 VDD.t607 1.6255
R3225 VDD.n1457 VDD.n1456 1.6255
R3226 VDD.n1459 VDD.t2309 1.6255
R3227 VDD.n1459 VDD.n1458 1.6255
R3228 VDD.n2256 VDD.t2281 1.6255
R3229 VDD.n2256 VDD.n2255 1.6255
R3230 VDD.n2253 VDD.t2423 1.6255
R3231 VDD.n2253 VDD.n2252 1.6255
R3232 VDD.n2247 VDD.t297 1.6255
R3233 VDD.n2247 VDD.n2246 1.6255
R3234 VDD.n2249 VDD.t2438 1.6255
R3235 VDD.n2249 VDD.n2248 1.6255
R3236 VDD.n2236 VDD.t2486 1.6255
R3237 VDD.n2236 VDD.n2235 1.6255
R3238 VDD.n2239 VDD.t2075 1.6255
R3239 VDD.n2239 VDD.n2238 1.6255
R3240 VDD.n1463 VDD.t1735 1.6255
R3241 VDD.n1463 VDD.n1462 1.6255
R3242 VDD.n1465 VDD.t2091 1.6255
R3243 VDD.n1465 VDD.n1464 1.6255
R3244 VDD.n1470 VDD.t1953 1.6255
R3245 VDD.n1470 VDD.n1469 1.6255
R3246 VDD.n1476 VDD.t773 1.6255
R3247 VDD.n1476 VDD.n1475 1.6255
R3248 VDD.n1485 VDD.t364 1.6255
R3249 VDD.n1485 VDD.n1484 1.6255
R3250 VDD.n1481 VDD.t772 1.6255
R3251 VDD.n1481 VDD.n1480 1.6255
R3252 VDD.n1479 VDD.t365 1.6255
R3253 VDD.n1479 VDD.n1478 1.6255
R3254 VDD.n1489 VDD.t1111 1.6255
R3255 VDD.n1489 VDD.n1488 1.6255
R3256 VDD.n1498 VDD.t1109 1.6255
R3257 VDD.n1498 VDD.n1497 1.6255
R3258 VDD.n1494 VDD.t1112 1.6255
R3259 VDD.n1494 VDD.n1493 1.6255
R3260 VDD.n1492 VDD.t1108 1.6255
R3261 VDD.n1492 VDD.n1491 1.6255
R3262 VDD.n1806 VDD.t729 1.6255
R3263 VDD.n1806 VDD.n1805 1.6255
R3264 VDD.n1809 VDD.t1819 1.6255
R3265 VDD.n1809 VDD.n1808 1.6255
R3266 VDD.n1865 VDD.t828 1.6255
R3267 VDD.n1865 VDD.n1864 1.6255
R3268 VDD.n1813 VDD.t749 1.6255
R3269 VDD.n1813 VDD.n1812 1.6255
R3270 VDD.n1817 VDD.t13 1.6255
R3271 VDD.n1817 VDD.n1816 1.6255
R3272 VDD.n1822 VDD.t2155 1.6255
R3273 VDD.n1822 VDD.n1821 1.6255
R3274 VDD.n1826 VDD.t1817 1.6255
R3275 VDD.n1826 VDD.n1825 1.6255
R3276 VDD.n1832 VDD.t1413 1.6255
R3277 VDD.n1832 VDD.n1831 1.6255
R3278 VDD.n1837 VDD.t737 1.6255
R3279 VDD.n1837 VDD.n1836 1.6255
R3280 VDD.n1800 VDD.t2342 1.6255
R3281 VDD.n1800 VDD.n1799 1.6255
R3282 VDD.n2051 VDD.t1342 1.6255
R3283 VDD.n2051 VDD.n2050 1.6255
R3284 VDD.n2048 VDD.t1725 1.6255
R3285 VDD.n2048 VDD.n2047 1.6255
R3286 VDD.n2060 VDD.t53 1.6255
R3287 VDD.n2060 VDD.n2059 1.6255
R3288 VDD.n2045 VDD.t1791 1.6255
R3289 VDD.n2045 VDD.n2044 1.6255
R3290 VDD.n2043 VDD.t935 1.6255
R3291 VDD.n2043 VDD.n2042 1.6255
R3292 VDD.n2040 VDD.t2729 1.6255
R3293 VDD.n2040 VDD.n2039 1.6255
R3294 VDD.n2037 VDD.t637 1.6255
R3295 VDD.n2037 VDD.n2036 1.6255
R3296 VDD.n2035 VDD.t1653 1.6255
R3297 VDD.n2035 VDD.n2034 1.6255
R3298 VDD.n2032 VDD.t1681 1.6255
R3299 VDD.n2032 VDD.n2031 1.6255
R3300 VDD.n2029 VDD.t1370 1.6255
R3301 VDD.n2029 VDD.n2028 1.6255
R3302 VDD.n2092 VDD.t310 1.6255
R3303 VDD.n2092 VDD.n2091 1.6255
R3304 VDD.n2090 VDD.t228 1.6255
R3305 VDD.n2090 VDD.n2089 1.6255
R3306 VDD.n2026 VDD.t243 1.6255
R3307 VDD.n2026 VDD.n2025 1.6255
R3308 VDD.n2023 VDD.t1970 1.6255
R3309 VDD.n2023 VDD.n2022 1.6255
R3310 VDD.n2020 VDD.t1727 1.6255
R3311 VDD.n2020 VDD.n2019 1.6255
R3312 VDD.n2018 VDD.t2178 1.6255
R3313 VDD.n2018 VDD.n2017 1.6255
R3314 VDD.n2015 VDD.t2162 1.6255
R3315 VDD.n2015 VDD.n2014 1.6255
R3316 VDD.n2012 VDD.t2461 1.6255
R3317 VDD.n2012 VDD.n2011 1.6255
R3318 VDD.n2123 VDD.t843 1.6255
R3319 VDD.n2123 VDD.n2122 1.6255
R3320 VDD.n2121 VDD.t1385 1.6255
R3321 VDD.n2121 VDD.n2120 1.6255
R3322 VDD.n2009 VDD.t1377 1.6255
R3323 VDD.n2009 VDD.n2008 1.6255
R3324 VDD.n2005 VDD.t2292 1.6255
R3325 VDD.n2005 VDD.n2004 1.6255
R3326 VDD.n1998 VDD.t579 1.6255
R3327 VDD.n1998 VDD.n1997 1.6255
R3328 VDD.n2000 VDD.t2302 1.6255
R3329 VDD.n2000 VDD.n1999 1.6255
R3330 VDD.n1986 VDD.t2271 1.6255
R3331 VDD.n1986 VDD.n1985 1.6255
R3332 VDD.n1983 VDD.t2418 1.6255
R3333 VDD.n1983 VDD.n1982 1.6255
R3334 VDD.n1977 VDD.t74 1.6255
R3335 VDD.n1977 VDD.n1976 1.6255
R3336 VDD.n1979 VDD.t2424 1.6255
R3337 VDD.n1979 VDD.n1978 1.6255
R3338 VDD.n1966 VDD.t2474 1.6255
R3339 VDD.n1966 VDD.n1965 1.6255
R3340 VDD.n1969 VDD.t2059 1.6255
R3341 VDD.n1969 VDD.n1968 1.6255
R3342 VDD.n1959 VDD.t991 1.6255
R3343 VDD.n1959 VDD.n1958 1.6255
R3344 VDD.n1961 VDD.t2079 1.6255
R3345 VDD.n1961 VDD.n1960 1.6255
R3346 VDD.n1952 VDD.t1938 1.6255
R3347 VDD.n1952 VDD.n1951 1.6255
R3348 VDD.n1939 VDD.t490 1.6255
R3349 VDD.n1939 VDD.n1938 1.6255
R3350 VDD.n1948 VDD.t1078 1.6255
R3351 VDD.n1948 VDD.n1947 1.6255
R3352 VDD.n1944 VDD.t491 1.6255
R3353 VDD.n1944 VDD.n1943 1.6255
R3354 VDD.n1942 VDD.t1077 1.6255
R3355 VDD.n1942 VDD.n1941 1.6255
R3356 VDD.n1926 VDD.t1797 1.6255
R3357 VDD.n1926 VDD.n1925 1.6255
R3358 VDD.n1935 VDD.t1133 1.6255
R3359 VDD.n1935 VDD.n1934 1.6255
R3360 VDD.n1931 VDD.t1796 1.6255
R3361 VDD.n1931 VDD.n1930 1.6255
R3362 VDD.n1929 VDD.t1134 1.6255
R3363 VDD.n1929 VDD.n1928 1.6255
R3364 VDD.n1773 VDD.t1161 1.6255
R3365 VDD.n1773 VDD.n1772 1.6255
R3366 VDD.n1779 VDD.t1093 1.6255
R3367 VDD.n1779 VDD.n1778 1.6255
R3368 VDD.n1789 VDD.t2593 1.6255
R3369 VDD.n1789 VDD.n1788 1.6255
R3370 VDD.n1785 VDD.t2575 1.6255
R3371 VDD.n1785 VDD.n1784 1.6255
R3372 VDD.n1917 VDD.t1152 1.6255
R3373 VDD.n1917 VDD.n1916 1.6255
R3374 VDD.n1793 VDD.t2245 1.6255
R3375 VDD.n1793 VDD.n1792 1.6255
R3376 VDD.n1900 VDD.t2589 1.6255
R3377 VDD.n1900 VDD.n1899 1.6255
R3378 VDD.n1796 VDD.t1466 1.6255
R3379 VDD.n1796 VDD.n1795 1.6255
R3380 VDD.n1769 VDD.t42 1.6255
R3381 VDD.n1769 VDD.n1768 1.6255
R3382 VDD.n1510 VDD.t2528 1.6255
R3383 VDD.n1510 VDD.n1509 1.6255
R3384 VDD.n1726 VDD.t2367 1.6255
R3385 VDD.n1726 VDD.n1725 1.6255
R3386 VDD.n1731 VDD.t2223 1.6255
R3387 VDD.n1731 VDD.n1730 1.6255
R3388 VDD.n1735 VDD.t2387 1.6255
R3389 VDD.n1735 VDD.n1734 1.6255
R3390 VDD.n1741 VDD.t1428 1.6255
R3391 VDD.n1741 VDD.n1740 1.6255
R3392 VDD.n1746 VDD.t2644 1.6255
R3393 VDD.n1746 VDD.n1745 1.6255
R3394 VDD.n2203 VDD.t1810 1.6255
R3395 VDD.n2203 VDD.n2202 1.6255
R3396 VDD.n1506 VDD.t2389 1.6255
R3397 VDD.n1506 VDD.n1505 1.6255
R3398 VDD.n1503 VDD.t2526 1.6255
R3399 VDD.n1503 VDD.n1502 1.6255
R3400 VDD.n1530 VDD.t2573 1.6255
R3401 VDD.n1530 VDD.n1529 1.6255
R3402 VDD.n1524 VDD.t1012 1.6255
R3403 VDD.n1524 VDD.n1523 1.6255
R3404 VDD.n1664 VDD.t2145 1.6255
R3405 VDD.n1664 VDD.n1663 1.6255
R3406 VDD.n1666 VDD.t699 1.6255
R3407 VDD.n1666 VDD.n1665 1.6255
R3408 VDD.n1671 VDD.t825 1.6255
R3409 VDD.n1671 VDD.n1670 1.6255
R3410 VDD.n1566 VDD.t2355 1.6255
R3411 VDD.n1566 VDD.n1565 1.6255
R3412 VDD.n1563 VDD.t943 1.6255
R3413 VDD.n1563 VDD.n1562 1.6255
R3414 VDD.n1557 VDD.t1301 1.6255
R3415 VDD.n1557 VDD.n1556 1.6255
R3416 VDD.n1559 VDD.t1312 1.6255
R3417 VDD.n1559 VDD.n1558 1.6255
R3418 VDD.n1577 VDD.t2504 1.6255
R3419 VDD.n1577 VDD.n1576 1.6255
R3420 VDD.n1580 VDD.t1999 1.6255
R3421 VDD.n1580 VDD.n1579 1.6255
R3422 VDD.n1643 VDD.t125 1.6255
R3423 VDD.n1643 VDD.n1642 1.6255
R3424 VDD.n1584 VDD.t2513 1.6255
R3425 VDD.n1584 VDD.n1583 1.6255
R3426 VDD.n1588 VDD.t113 1.6255
R3427 VDD.n1588 VDD.n1587 1.6255
R3428 VDD.n135 VDD.t716 1.59425
R3429 VDD.n677 VDD.t2689 1.59425
R3430 VDD.n403 VDD.n402 1.59425
R3431 VDD.n172 VDD.n171 1.59425
R3432 VDD.n1135 VDD.n1134 1.59425
R3433 VDD.n262 VDD.t460 1.59425
R3434 VDD.n500 VDD.n499 1.59425
R3435 VDD.n2185 VDD.n2184 1.5005
R3436 VDD.n1766 VDD.n1765 1.5005
R3437 VDD.n1661 VDD.n1660 1.4405
R3438 VDD.n2263 VDD.n2262 1.3505
R3439 VDD.n2140 VDD.n1992 1.3505
R3440 VDD.n2276 VDD.n1455 1.328
R3441 VDD.n2133 VDD.n2007 1.328
R3442 VDD.n2187 VDD.n2186 1.27445
R3443 VDD.n851 VDD.n848 1.23657
R3444 VDD.n1482 VDD.n1479 1.23657
R3445 VDD.n1495 VDD.n1492 1.23657
R3446 VDD.n1945 VDD.n1942 1.23657
R3447 VDD.n1932 VDD.n1929 1.23657
R3448 VDD.n1573 VDD.n1571 1.23637
R3449 VDD.n155 VDD.n151 1.23637
R3450 VDD.n287 VDD.n283 1.23637
R3451 VDD.n1328 VDD.n1324 1.23637
R3452 VDD.n653 VDD.n649 1.23637
R3453 VDD.n63 VDD.n61 1.23637
R3454 VDD.n44 VDD.n42 1.23637
R3455 VDD.n115 VDD.n111 1.23637
R3456 VDD.n2373 VDD.n2371 1.23637
R3457 VDD.n1236 VDD.n1234 1.23637
R3458 VDD.n459 VDD.n457 1.23637
R3459 VDD.n440 VDD.n438 1.23637
R3460 VDD.n1802 VDD.n1800 1.23637
R3461 VDD.n1673 VDD.n1671 1.23637
R3462 VDD.n347 VDD.n343 1.23591
R3463 VDD.n757 VDD.n753 1.23591
R3464 VDD.n701 VDD.n697 1.23591
R3465 VDD.n1007 VDD.n1005 1.23591
R3466 VDD.n1075 VDD.n1073 1.23591
R3467 VDD.n1094 VDD.n1092 1.23591
R3468 VDD.n1181 VDD.n1179 1.23591
R3469 VDD.n1155 VDD.n1153 1.23591
R3470 VDD.n229 VDD.n225 1.23591
R3471 VDD.n518 VDD.n516 1.23591
R3472 VDD.n2264 VDD 1.21734
R3473 VDD VDD.n2141 1.21734
R3474 VDD.n2319 VDD.n197 1.17585
R3475 VDD.n961 VDD.n960 1.17585
R3476 VDD.n897 VDD.n893 1.17585
R3477 VDD.n916 VDD.n915 1.17585
R3478 VDD.n2340 VDD.n187 1.17585
R3479 VDD.n976 VDD.n975 1.17585
R3480 VDD.n2327 VDD.n198 1.17044
R3481 VDD.n951 VDD.n950 1.17044
R3482 VDD.n904 VDD.n900 1.17044
R3483 VDD.n930 VDD.n918 1.17044
R3484 VDD.n2347 VDD.n2343 1.17044
R3485 VDD.n989 VDD.n978 1.17044
R3486 VDD.n947 VDD.n200 1.15088
R3487 VDD.n2271 VDD 1.13101
R3488 VDD VDD.n2137 1.13101
R3489 VDD.n996 VDD.n969 1.11767
R3490 VDD.n2354 VDD.n2353 1.08484
R3491 VDD.n2315 VDD.n2314 1.07484
R3492 VDD.n2268 VDD.n2267 1.05938
R3493 VDD.n2139 VDD.n2138 1.05938
R3494 VDD.n2356 VDD.n2355 0.985783
R3495 VDD.n1369 VDD.n200 0.98484
R3496 VDD VDD.n2230 0.97948
R3497 VDD.n2145 VDD 0.97948
R3498 VDD VDD.n2263 0.973969
R3499 VDD VDD.n2140 0.973969
R3500 VDD.n326 VDD.n325 0.969146
R3501 VDD.n740 VDD.n739 0.969146
R3502 VDD.n55 VDD.n54 0.969146
R3503 VDD.n2436 VDD.n2435 0.969146
R3504 VDD.n1290 VDD.n1289 0.969146
R3505 VDD.n1216 VDD.n1215 0.969146
R3506 VDD.n494 VDD.n493 0.969146
R3507 VDD VDD.n598 0.948722
R3508 VDD VDD.n1815 0.948722
R3509 VDD VDD.n1586 0.948722
R3510 VDD.n880 VDD.n879 0.947457
R3511 VDD.n881 VDD.n880 0.947457
R3512 VDD.n882 VDD.n881 0.947457
R3513 VDD.n883 VDD.n882 0.947457
R3514 VDD.n138 VDD.n137 0.938
R3515 VDD.n680 VDD.n679 0.938
R3516 VDD.n401 VDD.t2253 0.938
R3517 VDD.n170 VDD.t622 0.938
R3518 VDD.n1133 VDD.t2442 0.938
R3519 VDD.n265 VDD.n264 0.938
R3520 VDD.n498 VDD.t88 0.938
R3521 VDD.n2172 VDD.n1771 0.936986
R3522 VDD.n1909 VDD.n1906 0.923351
R3523 VDD.n142 VDD.n140 0.919433
R3524 VDD.n683 VDD.n682 0.919433
R3525 VDD.n407 VDD.n406 0.919433
R3526 VDD.n176 VDD.n175 0.919433
R3527 VDD.n1139 VDD.n1138 0.919433
R3528 VDD.n269 VDD.n267 0.919433
R3529 VDD.n504 VDD.n503 0.919433
R3530 VDD.n1617 VDD 0.90746
R3531 VDD VDD.n1704 0.90746
R3532 VDD.n806 VDD 0.90746
R3533 VDD.n1846 VDD 0.90746
R3534 VDD.n1755 VDD 0.90746
R3535 VDD VDD.n1633 0.894579
R3536 VDD.n2314 VDD.n1369 0.888236
R3537 VDD VDD.n1536 0.883046
R3538 VDD VDD.n594 0.883046
R3539 VDD VDD.n1811 0.883046
R3540 VDD VDD.n1508 0.883046
R3541 VDD VDD.n1582 0.883046
R3542 VDD.n2234 VDD.n1467 0.870194
R3543 VDD.n2275 VDD.n1461 0.870194
R3544 VDD.n2143 VDD.n2142 0.870194
R3545 VDD.n2135 VDD.n2134 0.870194
R3546 VDD.n852 VDD.n851 0.831962
R3547 VDD.n1483 VDD.n1482 0.831962
R3548 VDD.n1496 VDD.n1495 0.831962
R3549 VDD.n1946 VDD.n1945 0.831962
R3550 VDD.n1933 VDD.n1932 0.831962
R3551 VDD.n1067 VDD.n341 0.817542
R3552 VDD.n673 VDD.n672 0.817542
R3553 VDD.n1002 VDD.n1001 0.817542
R3554 VDD.n2368 VDD.n2364 0.817542
R3555 VDD.n1231 VDD.n1230 0.817542
R3556 VDD.n259 VDD.n258 0.817542
R3557 VDD.n563 VDD.n562 0.817542
R3558 VDD VDD.n298 0.792598
R3559 VDD VDD.n713 0.792598
R3560 VDD VDD.n89 0.792598
R3561 VDD VDD.n92 0.792598
R3562 VDD VDD.n1107 0.792598
R3563 VDD VDD.n1194 0.792598
R3564 VDD VDD.n472 0.792598
R3565 VDD.n875 VDD.n874 0.763264
R3566 VDD VDD.n435 0.750764
R3567 VDD.n780 VDD.n673 0.74033
R3568 VDD.n1351 VDD.n259 0.74033
R3569 VDD.n1001 VDD.n1000 0.739568
R3570 VDD.n564 VDD.n563 0.739568
R3571 VDD.n2165 VDD 0.731756
R3572 VDD.n325 VDD 0.7301
R3573 VDD VDD.n1067 0.7301
R3574 VDD.n739 VDD 0.7301
R3575 VDD.n672 VDD 0.7301
R3576 VDD VDD.n1002 0.7301
R3577 VDD VDD.n55 0.7301
R3578 VDD.n2462 VDD 0.7301
R3579 VDD VDD.n2436 0.7301
R3580 VDD VDD.n2368 0.7301
R3581 VDD.n1289 VDD 0.7301
R3582 VDD VDD.n1231 0.7301
R3583 VDD.n1215 VDD 0.7301
R3584 VDD.n258 VDD 0.7301
R3585 VDD.n562 VDD 0.7301
R3586 VDD.n493 VDD 0.7301
R3587 VDD.n2477 VDD.n2476 0.715763
R3588 VDD.n138 VDD.n133 0.688
R3589 VDD.n680 VDD.n675 0.688
R3590 VDD.n401 VDD.n400 0.688
R3591 VDD.n170 VDD.n169 0.688
R3592 VDD.n1133 VDD.n1132 0.688
R3593 VDD.n265 VDD.n260 0.688
R3594 VDD.n498 VDD.n497 0.688
R3595 VDD.n162 VDD.n161 0.652313
R3596 VDD.n310 VDD.n288 0.652313
R3597 VDD.n1344 VDD.n1343 0.652313
R3598 VDD.n773 VDD.n772 0.652313
R3599 VDD.n732 VDD.n702 0.652313
R3600 VDD.n65 VDD.n64 0.652313
R3601 VDD.n49 VDD.n45 0.652313
R3602 VDD.n2439 VDD.n2438 0.652313
R3603 VDD.n1309 VDD.n1308 0.652313
R3604 VDD.n1287 VDD.n1286 0.652313
R3605 VDD.n1213 VDD.n1212 0.652313
R3606 VDD.n1170 VDD.n1169 0.652313
R3607 VDD.n491 VDD.n490 0.652313
R3608 VDD.n583 VDD.n582 0.652313
R3609 VDD.n1676 VDD.n1675 0.652313
R3610 VDD.n1574 VDD.n1573 0.64106
R3611 VDD VDD.n2471 0.639914
R3612 VDD.n2295 VDD 0.630343
R3613 VDD VDD.n1438 0.630343
R3614 VDD VDD.n2088 0.630343
R3615 VDD.n2104 VDD 0.630343
R3616 VDD VDD.n2119 0.630343
R3617 VDD.n2305 VDD 0.624338
R3618 VDD.n2073 VDD 0.624338
R3619 VDD.n717 VDD.n716 0.579377
R3620 VDD.n746 VDD.n687 0.579377
R3621 VDD.n88 VDD.n87 0.579377
R3622 VDD.n417 VDD.n416 0.579377
R3623 VDD.n2450 VDD.n2449 0.579377
R3624 VDD.n2433 VDD.n2432 0.579377
R3625 VDD.n1196 VDD.n1195 0.579377
R3626 VDD.n1218 VDD.n1217 0.579377
R3627 VDD.n474 VDD.n473 0.579377
R3628 VDD.n496 VDD.n495 0.579377
R3629 VDD.n304 VDD.n293 0.579377
R3630 VDD.n1292 VDD.n1291 0.579377
R3631 VDD.n1270 VDD.n1269 0.579377
R3632 VDD.n1689 VDD.n1555 0.578376
R3633 VDD.n2467 VDD.n35 0.569616
R3634 VDD VDD.n869 0.566011
R3635 VDD VDD.n1882 0.565659
R3636 VDD.n2299 VDD.n2298 0.561058
R3637 VDD.n2083 VDD.n2082 0.561058
R3638 VDD.n802 VDD.n791 0.55925
R3639 VDD.n841 VDD.n587 0.555209
R3640 VDD.n337 VDD.n335 0.552239
R3641 VDD.n143 VDD.n142 0.552239
R3642 VDD.n779 VDD.n683 0.552239
R3643 VDD.n641 VDD.n640 0.552239
R3644 VDD.n430 VDD.n407 0.552239
R3645 VDD.n396 VDD.n395 0.552239
R3646 VDD.n2360 VDD.n2359 0.552239
R3647 VDD.n177 VDD.n176 0.552239
R3648 VDD.n1125 VDD.n1124 0.552239
R3649 VDD.n1221 VDD.n1139 0.552239
R3650 VDD.n251 VDD.n249 0.552239
R3651 VDD.n1350 VDD.n269 0.552239
R3652 VDD.n565 VDD.n504 0.552239
R3653 VDD.n509 VDD.n508 0.552239
R3654 VDD.n2419 VDD.n2364 0.550415
R3655 VDD.n1230 VDD.n1229 0.54889
R3656 VDD.n1044 VDD.n1043 0.537223
R3657 VDD.n619 VDD.n618 0.537223
R3658 VDD.n1039 VDD.n1038 0.537223
R3659 VDD.n2407 VDD.n2406 0.537223
R3660 VDD.n1266 VDD.n1265 0.537223
R3661 VDD.n204 VDD.n203 0.537223
R3662 VDD.n1367 VDD.n1366 0.537223
R3663 VDD.n2285 VDD.n181 0.530241
R3664 VDD.n2471 VDD.n2470 0.512079
R3665 VDD.n1633 VDD.n1 0.512079
R3666 VDD.n2478 VDD.n2477 0.512079
R3667 VDD.n2476 VDD.n2475 0.512079
R3668 VDD.n2473 VDD.n2472 0.510717
R3669 VDD.n1614 VDD.n1613 0.505435
R3670 VDD.n1711 VDD.n1710 0.505435
R3671 VDD.n1543 VDD.n1514 0.505435
R3672 VDD.n834 VDD.n590 0.505435
R3673 VDD.n1874 VDD.n1807 0.505435
R3674 VDD.n1843 VDD.n1842 0.505435
R3675 VDD.n1914 VDD.n1913 0.505435
R3676 VDD.n1752 VDD.n1751 0.505435
R3677 VDD.n2212 VDD.n1504 0.505435
R3678 VDD.n1652 VDD.n1578 0.505435
R3679 VDD.n1623 VDD.n1622 0.50509
R3680 VDD.n1695 VDD.n1694 0.50509
R3681 VDD.n812 VDD.n811 0.50509
R3682 VDD.n1852 VDD.n1851 0.50509
R3683 VDD.n1897 VDD.n1896 0.50509
R3684 VDD.n1885 VDD.n1802 0.499244
R3685 VDD.n311 VDD.n310 0.492652
R3686 VDD.n1345 VDD.n1344 0.492652
R3687 VDD.n733 VDD.n732 0.492652
R3688 VDD.n774 VDD.n773 0.492652
R3689 VDD.n66 VDD.n65 0.492652
R3690 VDD.n50 VDD.n49 0.492652
R3691 VDD.n2440 VDD.n2439 0.492652
R3692 VDD.n161 VDD.n160 0.492652
R3693 VDD.n1308 VDD.n1307 0.492652
R3694 VDD.n1286 VDD.n1285 0.492652
R3695 VDD.n1212 VDD.n1211 0.492652
R3696 VDD.n1171 VDD.n1170 0.492652
R3697 VDD.n490 VDD.n489 0.492652
R3698 VDD.n582 VDD.n581 0.492652
R3699 VDD.n1381 VDD.n1380 0.492652
R3700 VDD.n2310 VDD.n2309 0.492652
R3701 VDD.n2058 VDD.n2057 0.492652
R3702 VDD.n2064 VDD.n2063 0.492652
R3703 VDD.n2062 VDD.n2046 0.492652
R3704 VDD.n2070 VDD.n2069 0.492652
R3705 VDD.n1675 VDD.n1564 0.492652
R3706 VDD.n867 VDD.n843 0.485854
R3707 VDD.n1616 VDD 0.484396
R3708 VDD.n1706 VDD 0.484396
R3709 VDD.n805 VDD 0.484396
R3710 VDD.n1845 VDD 0.484396
R3711 VDD.n1908 VDD 0.484396
R3712 VDD.n1754 VDD 0.484396
R3713 VDD.n162 VDD.n155 0.48386
R3714 VDD.n288 VDD.n287 0.48386
R3715 VDD.n1343 VDD.n1328 0.48386
R3716 VDD.n670 VDD.n653 0.48386
R3717 VDD.n64 VDD.n63 0.48386
R3718 VDD.n45 VDD.n44 0.48386
R3719 VDD.n2438 VDD.n115 0.48386
R3720 VDD.n2374 VDD.n2373 0.48386
R3721 VDD.n1237 VDD.n1236 0.48386
R3722 VDD.n491 VDD.n459 0.48386
R3723 VDD.n583 VDD.n440 0.48386
R3724 VDD.n1676 VDD.n1673 0.48386
R3725 VDD.n1662 VDD.n1661 0.483752
R3726 VDD.n1063 VDD.n347 0.483349
R3727 VDD.n772 VDD.n757 0.483349
R3728 VDD.n702 VDD.n701 0.483349
R3729 VDD.n1008 VDD.n1007 0.483349
R3730 VDD.n1309 VDD.n1075 0.483349
R3731 VDD.n1287 VDD.n1094 0.483349
R3732 VDD.n1213 VDD.n1181 0.483349
R3733 VDD.n1169 VDD.n1155 0.483349
R3734 VDD.n230 VDD.n229 0.483349
R3735 VDD.n560 VDD.n518 0.483349
R3736 VDD VDD.n1721 0.48089
R3737 VDD.n840 VDD 0.48089
R3738 VDD.n1880 VDD 0.48089
R3739 VDD.n2218 VDD 0.48089
R3740 VDD.n1658 VDD 0.48089
R3741 VDD.n1625 VDD 0.466864
R3742 VDD VDD.n1691 0.466864
R3743 VDD.n814 VDD 0.466864
R3744 VDD.n1854 VDD 0.466864
R3745 VDD.n2193 VDD 0.466864
R3746 VDD.n2056 VDD 0.465572
R3747 VDD.n485 VDD.n484 0.463032
R3748 VDD.n550 VDD.n549 0.463032
R3749 VDD.n1281 VDD.n1280 0.463032
R3750 VDD.n2447 VDD.n2446 0.463032
R3751 VDD.n428 VDD.n427 0.463032
R3752 VDD.n1331 VDD.n271 0.463032
R3753 VDD.n316 VDD.n315 0.463032
R3754 VDD.n314 VDD.n313 0.463032
R3755 VDD.n1348 VDD.n1347 0.463032
R3756 VDD.n363 VDD.n362 0.463032
R3757 VDD.n727 VDD.n726 0.463032
R3758 VDD.n763 VDD.n685 0.463032
R3759 VDD.n729 VDD.n728 0.463032
R3760 VDD.n777 VDD.n776 0.463032
R3761 VDD.n786 VDD.n785 0.463032
R3762 VDD.n1027 VDD.n1026 0.463032
R3763 VDD.n85 VDD.n84 0.463032
R3764 VDD.n86 VDD.n75 0.463032
R3765 VDD.n418 VDD.n410 0.463032
R3766 VDD.n2448 VDD.n101 0.463032
R3767 VDD.n2431 VDD.n132 0.463032
R3768 VDD.n2429 VDD.n2428 0.463032
R3769 VDD.n2397 VDD.n2396 0.463032
R3770 VDD.n1302 VDD.n1301 0.463032
R3771 VDD.n1305 VDD.n1304 0.463032
R3772 VDD.n1283 VDD.n1282 0.463032
R3773 VDD.n1260 VDD.n1259 0.463032
R3774 VDD.n1207 VDD.n1206 0.463032
R3775 VDD.n1209 VDD.n1208 0.463032
R3776 VDD.n1219 VDD.n1143 0.463032
R3777 VDD.n1163 VDD.n1140 0.463032
R3778 VDD.n239 VDD.n238 0.463032
R3779 VDD.n576 VDD.n575 0.463032
R3780 VDD.n487 VDD.n486 0.463032
R3781 VDD.n579 VDD.n578 0.463032
R3782 VDD.n1683 VDD.n1682 0.463032
R3783 VDD.n1685 VDD.n1684 0.463032
R3784 VDD.n2473 VDD.n20 0.458326
R3785 VDD.n2476 VDD.n13 0.458326
R3786 VDD.n2478 VDD.n7 0.458326
R3787 VDD.n1633 VDD.n1632 0.458326
R3788 VDD.n2468 VDD.n34 0.458326
R3789 VDD.n2471 VDD.n27 0.458326
R3790 VDD.n1315 VDD.n341 0.456602
R3791 VDD.n2225 VDD.n2224 0.454602
R3792 VDD.n2151 VDD.n2150 0.454602
R3793 VDD.n2475 VDD.n14 0.45408
R3794 VDD.n1 VDD.n0 0.45408
R3795 VDD.n2470 VDD.n28 0.45408
R3796 VDD.n884 VDD.n883 0.453435
R3797 VDD.n2313 VDD.n1371 0.451639
R3798 VDD.n2293 VDD.n2292 0.450109
R3799 VDD.n1428 VDD.n1427 0.450109
R3800 VDD.n1449 VDD.n1448 0.450109
R3801 VDD.n2096 VDD.n2095 0.450109
R3802 VDD.n2110 VDD.n2109 0.450109
R3803 VDD.n2127 VDD.n2126 0.450109
R3804 VDD.n2477 VDD.n8 0.450011
R3805 VDD.n2303 VDD.n2302 0.446018
R3806 VDD.n2079 VDD.n2078 0.446018
R3807 VDD.n2472 VDD.n21 0.442185
R3808 VDD.n2309 VDD.n2308 0.436623
R3809 VDD.n2071 VDD.n2070 0.436623
R3810 VDD.n1317 VDD.n331 0.434848
R3811 VDD.n326 VDD.n278 0.434848
R3812 VDD.n304 VDD.n303 0.434848
R3813 VDD.n1048 VDD.n369 0.434848
R3814 VDD.n716 VDD.n710 0.434848
R3815 VDD.n740 VDD.n692 0.434848
R3816 VDD.n746 VDD.n745 0.434848
R3817 VDD.n789 VDD.n625 0.434848
R3818 VDD.n88 VDD.n72 0.434848
R3819 VDD.n54 VDD.n53 0.434848
R3820 VDD.n416 VDD.n415 0.434848
R3821 VDD.n2450 VDD.n97 0.434848
R3822 VDD.n2433 VDD.n128 0.434848
R3823 VDD.n2435 VDD.n122 0.434848
R3824 VDD.n2408 VDD.n2404 0.434848
R3825 VDD.n1291 VDD.n1086 0.434848
R3826 VDD.n1290 VDD.n1088 0.434848
R3827 VDD.n1269 VDD.n1105 0.434848
R3828 VDD.n1113 VDD.n1112 0.434848
R3829 VDD.n1195 VDD.n1192 0.434848
R3830 VDD.n1217 VDD.n1148 0.434848
R3831 VDD.n1216 VDD.n1175 0.434848
R3832 VDD.n211 VDD.n210 0.434848
R3833 VDD.n536 VDD.n535 0.434848
R3834 VDD.n473 VDD.n470 0.434848
R3835 VDD.n494 VDD.n453 0.434848
R3836 VDD.n495 VDD.n451 0.434848
R3837 VDD.n1561 VDD.n1560 0.434848
R3838 VDD VDD.n143 0.434483
R3839 VDD VDD.n779 0.434483
R3840 VDD VDD.n430 0.434483
R3841 VDD VDD.n1350 0.434483
R3842 VDD.n565 VDD 0.434483
R3843 VDD.n2057 VDD.n2056 0.421551
R3844 VDD.n2220 VDD.n1500 0.41984
R3845 VDD.n2155 VDD.n1924 0.41984
R3846 VDD.n1618 VDD 0.417987
R3847 VDD.n1609 VDD 0.417987
R3848 VDD.n1699 VDD 0.417987
R3849 VDD.n1715 VDD 0.417987
R3850 VDD.n1540 VDD 0.417987
R3851 VDD.n831 VDD 0.417987
R3852 VDD.n820 VDD 0.417987
R3853 VDD.n807 VDD 0.417987
R3854 VDD.n797 VDD 0.417987
R3855 VDD.n1871 VDD 0.417987
R3856 VDD.n1860 VDD 0.417987
R3857 VDD.n1847 VDD 0.417987
R3858 VDD.n1838 VDD 0.417987
R3859 VDD.n1918 VDD 0.417987
R3860 VDD.n1901 VDD 0.417987
R3861 VDD.n2198 VDD 0.417987
R3862 VDD.n1756 VDD 0.417987
R3863 VDD.n1747 VDD 0.417987
R3864 VDD.n2209 VDD 0.417987
R3865 VDD VDD.n1552 0.417987
R3866 VDD.n1649 VDD 0.417987
R3867 VDD.n1638 VDD 0.417987
R3868 VDD VDD.n788 0.412675
R3869 VDD VDD.n1050 0.412675
R3870 VDD VDD.n2399 0.412675
R3871 VDD VDD.n1262 0.412675
R3872 VDD.n236 VDD 0.412675
R3873 VDD.n537 VDD 0.412675
R3874 VDD.n375 VDD.n374 0.4055
R3875 VDD.n816 VDD.n815 0.401325
R3876 VDD.n1856 VDD.n1855 0.401325
R3877 VDD.n1627 VDD.n1626 0.401325
R3878 VDD.n1032 VDD.n377 0.399234
R3879 VDD VDD.n1893 0.398608
R3880 VDD.n2293 VDD.n1410 0.397674
R3881 VDD.n1427 VDD.n1426 0.397674
R3882 VDD.n1448 VDD.n1447 0.397674
R3883 VDD.n1461 VDD.n1460 0.397674
R3884 VDD.n1467 VDD.n1466 0.397674
R3885 VDD.n2096 VDD.n2093 0.397674
R3886 VDD.n2109 VDD.n2021 0.397674
R3887 VDD.n2127 VDD.n2124 0.397674
R3888 VDD.n2135 VDD.n2001 0.397674
R3889 VDD.n2143 VDD.n1962 0.397674
R3890 VDD VDD.n586 0.39672
R3891 VDD.n2303 VDD.n1396 0.395717
R3892 VDD.n2078 VDD.n2038 0.395717
R3893 VDD.n2189 VDD.n2188 0.393036
R3894 VDD.n2468 VDD.n2467 0.392474
R3895 VDD.n866 VDD.n865 0.392399
R3896 VDD.n2223 VDD.n1487 0.392399
R3897 VDD.n2222 VDD.n2221 0.392399
R3898 VDD.n2149 VDD.n2148 0.392399
R3899 VDD.n2154 VDD.n2153 0.392399
R3900 VDD.n2375 VDD.n2374 0.389831
R3901 VDD.n1238 VDD.n1237 0.389831
R3902 VDD.n1063 VDD.n1062 0.38879
R3903 VDD.n670 VDD.n669 0.38879
R3904 VDD.n1009 VDD.n1008 0.38879
R3905 VDD.n230 VDD.n223 0.38879
R3906 VDD.n560 VDD.n559 0.38879
R3907 VDD.n1575 VDD 0.385855
R3908 VDD VDD.n598 0.384624
R3909 VDD VDD.n1815 0.384624
R3910 VDD VDD.n842 0.382708
R3911 VDD.n385 VDD.n384 0.381864
R3912 VDD.n1380 VDD.n1371 0.381006
R3913 VDD.n2063 VDD.n2062 0.381006
R3914 VDD.n1619 VDD.n1618 0.370786
R3915 VDD.n1610 VDD.n1609 0.370786
R3916 VDD.n1700 VDD.n1699 0.370786
R3917 VDD.n1716 VDD.n1715 0.370786
R3918 VDD.n1541 VDD.n1540 0.370786
R3919 VDD.n832 VDD.n831 0.370786
R3920 VDD.n821 VDD.n820 0.370786
R3921 VDD.n808 VDD.n807 0.370786
R3922 VDD.n798 VDD.n797 0.370786
R3923 VDD.n1872 VDD.n1871 0.370786
R3924 VDD.n1861 VDD.n1860 0.370786
R3925 VDD.n1848 VDD.n1847 0.370786
R3926 VDD.n1839 VDD.n1838 0.370786
R3927 VDD.n1919 VDD.n1918 0.370786
R3928 VDD.n1902 VDD.n1901 0.370786
R3929 VDD.n2199 VDD.n2198 0.370786
R3930 VDD.n1757 VDD.n1756 0.370786
R3931 VDD.n1748 VDD.n1747 0.370786
R3932 VDD.n2210 VDD.n2209 0.370786
R3933 VDD.n1552 VDD.n1551 0.370786
R3934 VDD.n1650 VDD.n1649 0.370786
R3935 VDD.n1639 VDD.n1638 0.370786
R3936 VDD.n2464 VDD.n2463 0.368475
R3937 VDD.n2262 VDD.n2250 0.364413
R3938 VDD.n1992 VDD.n1980 0.364413
R3939 VDD VDD.n326 0.35825
R3940 VDD VDD.n740 0.35825
R3941 VDD.n54 VDD 0.35825
R3942 VDD.n2435 VDD 0.35825
R3943 VDD VDD.n1290 0.35825
R3944 VDD VDD.n1216 0.35825
R3945 VDD VDD.n494 0.35825
R3946 VDD.n1621 VDD 0.355357
R3947 VDD.n1612 VDD 0.355357
R3948 VDD VDD.n1696 0.355357
R3949 VDD VDD.n1712 0.355357
R3950 VDD VDD.n1544 0.355357
R3951 VDD VDD.n835 0.355357
R3952 VDD.n810 VDD 0.355357
R3953 VDD.n800 VDD 0.355357
R3954 VDD VDD.n1875 0.355357
R3955 VDD.n1850 VDD 0.355357
R3956 VDD.n1841 VDD 0.355357
R3957 VDD VDD.n1915 0.355357
R3958 VDD VDD.n1898 0.355357
R3959 VDD.n1759 VDD 0.355357
R3960 VDD.n1750 VDD 0.355357
R3961 VDD VDD.n2213 0.355357
R3962 VDD VDD.n1653 0.355357
R3963 VDD.n1536 VDD 0.352009
R3964 VDD VDD.n594 0.352009
R3965 VDD VDD.n1811 0.352009
R3966 VDD VDD.n1508 0.352009
R3967 VDD VDD.n1582 0.352009
R3968 VDD VDD.n1616 0.348937
R3969 VDD VDD.n1706 0.348937
R3970 VDD VDD.n805 0.348937
R3971 VDD VDD.n1845 0.348937
R3972 VDD VDD.n1754 0.348937
R3973 VDD VDD.n2164 0.345969
R3974 VDD.n1316 VDD.n273 0.342002
R3975 VDD.n2302 VDD.n2301 0.338587
R3976 VDD.n2292 VDD.n2291 0.338587
R3977 VDD.n1429 VDD.n1428 0.338587
R3978 VDD.n1450 VDD.n1449 0.338587
R3979 VDD.n2080 VDD.n2079 0.338587
R3980 VDD.n2095 VDD.n2027 0.338587
R3981 VDD.n2111 VDD.n2110 0.338587
R3982 VDD.n2126 VDD.n2010 0.338587
R3983 VDD.n1222 VDD.n1221 0.338381
R3984 VDD.n1316 VDD.n1315 0.337206
R3985 VDD.n2422 VDD.n177 0.336093
R3986 VDD.n2308 VDD.n2307 0.335672
R3987 VDD.n2298 VDD.n2297 0.335672
R3988 VDD.n2288 VDD.n2287 0.335672
R3989 VDD.n1436 VDD.n1435 0.335672
R3990 VDD.n2072 VDD.n2071 0.335672
R3991 VDD.n2082 VDD.n2030 0.335672
R3992 VDD.n2103 VDD.n2102 0.335672
R3993 VDD.n2113 VDD.n2013 0.335672
R3994 VDD.n1909 VDD.n1908 0.33125
R3995 VDD.n2164 VDD.n2163 0.327223
R3996 VDD.n2160 VDD.n2159 0.327223
R3997 VDD.n2470 VDD 0.326158
R3998 VDD VDD.n1 0.326158
R3999 VDD.n2475 VDD 0.326158
R4000 VDD VDD.n2299 0.3245
R4001 VDD VDD.n2289 0.3245
R4002 VDD.n1434 VDD 0.3245
R4003 VDD VDD.n2277 0.3245
R4004 VDD VDD.n2083 0.3245
R4005 VDD.n2101 VDD 0.3245
R4006 VDD VDD.n2114 0.3245
R4007 VDD.n2132 VDD 0.3245
R4008 VDD VDD.n2305 0.321707
R4009 VDD VDD.n2295 0.321707
R4010 VDD VDD.n2285 0.321707
R4011 VDD.n1438 VDD 0.321707
R4012 VDD VDD.n2073 0.321707
R4013 VDD.n2088 VDD 0.321707
R4014 VDD VDD.n2104 0.321707
R4015 VDD.n2119 VDD 0.321707
R4016 VDD.n1775 VDD 0.320891
R4017 VDD.n2189 VDD 0.320538
R4018 VDD VDD.n2161 0.313609
R4019 VDD VDD.n2157 0.31134
R4020 VDD VDD.n2165 0.308434
R4021 VDD.n802 VDD.n801 0.306734
R4022 VDD.n340 VDD.n337 0.305717
R4023 VDD.n644 VDD.n641 0.305717
R4024 VDD.n399 VDD.n396 0.305717
R4025 VDD.n2363 VDD.n2360 0.305717
R4026 VDD.n1128 VDD.n1125 0.305717
R4027 VDD.n254 VDD.n251 0.305717
R4028 VDD.n512 VDD.n509 0.305717
R4029 VDD.n1776 VDD.n1775 0.30425
R4030 VDD.n865 VDD.n855 0.290533
R4031 VDD.n1487 VDD.n1486 0.290533
R4032 VDD.n2222 VDD.n1499 0.290533
R4033 VDD.n2148 VDD.n1949 0.290533
R4034 VDD.n2153 VDD.n1936 0.290533
R4035 VDD.n865 VDD.n864 0.289867
R4036 VDD.n2229 VDD.n1487 0.289867
R4037 VDD.n2226 VDD.n2222 0.289867
R4038 VDD.n2148 VDD.n2147 0.289867
R4039 VDD.n2153 VDD.n2152 0.289867
R4040 VDD.n1435 VDD.n1434 0.288115
R4041 VDD.n2114 VDD.n2113 0.288115
R4042 VDD.n1622 VDD.n1621 0.287841
R4043 VDD.n1696 VDD.n1695 0.287841
R4044 VDD.n811 VDD.n810 0.287841
R4045 VDD.n1851 VDD.n1850 0.287841
R4046 VDD.n1898 VDD.n1897 0.287841
R4047 VDD.n1760 VDD.n1759 0.287841
R4048 VDD.n1315 VDD.n1314 0.284229
R4049 VDD.n2289 VDD.n2288 0.281855
R4050 VDD.n2102 VDD.n2101 0.281855
R4051 VDD.n1613 VDD.n1612 0.281308
R4052 VDD.n1712 VDD.n1711 0.281308
R4053 VDD.n801 VDD.n800 0.281308
R4054 VDD.n1842 VDD.n1841 0.281308
R4055 VDD.n1915 VDD.n1914 0.281308
R4056 VDD.n1751 VDD.n1750 0.281308
R4057 VDD.n1888 VDD.n1887 0.261586
R4058 VDD.n1892 VDD.n1888 0.261539
R4059 VDD.n1044 VDD 0.255875
R4060 VDD.n1039 VDD 0.255875
R4061 VDD VDD.n2407 0.255875
R4062 VDD VDD.n1266 0.255875
R4063 VDD VDD.n204 0.255875
R4064 VDD.n1053 VDD.n364 0.249097
R4065 VDD.n787 VDD.n628 0.249097
R4066 VDD.n1029 VDD.n1028 0.249097
R4067 VDD.n2398 VDD.n2387 0.249097
R4068 VDD.n1261 VDD.n1114 0.249097
R4069 VDD.n237 VDD.n212 0.249097
R4070 VDD.n552 VDD.n551 0.249097
R4071 VDD.n2191 VDD.n2190 0.248062
R4072 VDD.n483 VDD.n480 0.246576
R4073 VDD.n548 VDD.n543 0.246576
R4074 VDD.n1279 VDD.n1276 0.246576
R4075 VDD.n2445 VDD.n107 0.246576
R4076 VDD.n426 VDD.n424 0.246576
R4077 VDD.n1335 VDD.n1334 0.246576
R4078 VDD.n320 VDD.n319 0.246576
R4079 VDD.n312 VDD.n311 0.246576
R4080 VDD.n1346 VDD.n1345 0.246576
R4081 VDD.n1055 VDD.n351 0.246576
R4082 VDD.n361 VDD.n359 0.246576
R4083 VDD.n725 VDD.n723 0.246576
R4084 VDD.n767 VDD.n766 0.246576
R4085 VDD.n734 VDD.n733 0.246576
R4086 VDD.n775 VDD.n774 0.246576
R4087 VDD.n784 VDD.n634 0.246576
R4088 VDD.n662 VDD.n657 0.246576
R4089 VDD.n1025 VDD.n391 0.246576
R4090 VDD.n1017 VDD.n1016 0.246576
R4091 VDD.n83 VDD.n81 0.246576
R4092 VDD.n67 VDD.n66 0.246576
R4093 VDD.n51 VDD.n50 0.246576
R4094 VDD.n2441 VDD.n2440 0.246576
R4095 VDD.n160 VDD.n159 0.246576
R4096 VDD.n2427 VDD.n149 0.246576
R4097 VDD.n2395 VDD.n2393 0.246576
R4098 VDD.n2383 VDD.n2382 0.246576
R4099 VDD.n1300 VDD.n1298 0.246576
R4100 VDD.n1307 VDD.n1306 0.246576
R4101 VDD.n1285 VDD.n1284 0.246576
R4102 VDD.n1258 VDD.n1120 0.246576
R4103 VDD.n1249 VDD.n1245 0.246576
R4104 VDD.n1205 VDD.n1202 0.246576
R4105 VDD.n1211 VDD.n1210 0.246576
R4106 VDD.n1172 VDD.n1171 0.246576
R4107 VDD.n1164 VDD.n1160 0.246576
R4108 VDD.n219 VDD.n216 0.246576
R4109 VDD.n243 VDD.n242 0.246576
R4110 VDD.n555 VDD.n554 0.246576
R4111 VDD.n574 VDD.n571 0.246576
R4112 VDD.n489 VDD.n488 0.246576
R4113 VDD.n581 VDD.n580 0.246576
R4114 VDD.n1382 VDD.n1377 0.246576
R4115 VDD.n2312 VDD.n2311 0.246576
R4116 VDD.n2065 VDD.n2058 0.246576
R4117 VDD.n2068 VDD.n2046 0.246576
R4118 VDD.n1681 VDD.n1668 0.246576
R4119 VDD.n1686 VDD.n1564 0.246576
R4120 VDD.n484 VDD 0.245437
R4121 VDD.n549 VDD 0.245437
R4122 VDD.n1280 VDD 0.245437
R4123 VDD.n2446 VDD 0.245437
R4124 VDD.n427 VDD 0.245437
R4125 VDD VDD.n1331 0.245437
R4126 VDD VDD.n316 0.245437
R4127 VDD.n313 VDD 0.245437
R4128 VDD.n1347 VDD 0.245437
R4129 VDD VDD.n1054 0.245437
R4130 VDD.n362 VDD 0.245437
R4131 VDD.n726 VDD 0.245437
R4132 VDD VDD.n763 0.245437
R4133 VDD VDD.n729 0.245437
R4134 VDD.n776 VDD 0.245437
R4135 VDD.n785 VDD 0.245437
R4136 VDD VDD.n661 0.245437
R4137 VDD.n1026 VDD 0.245437
R4138 VDD VDD.n383 0.245437
R4139 VDD.n84 VDD 0.245437
R4140 VDD.n75 VDD 0.245437
R4141 VDD.n410 VDD 0.245437
R4142 VDD VDD.n101 0.245437
R4143 VDD VDD.n132 0.245437
R4144 VDD.n2428 VDD 0.245437
R4145 VDD.n2396 VDD 0.245437
R4146 VDD.n2386 VDD 0.245437
R4147 VDD.n1301 VDD 0.245437
R4148 VDD VDD.n1305 0.245437
R4149 VDD VDD.n1283 0.245437
R4150 VDD.n1259 VDD 0.245437
R4151 VDD VDD.n1248 0.245437
R4152 VDD.n1206 VDD 0.245437
R4153 VDD VDD.n1209 0.245437
R4154 VDD VDD.n1143 0.245437
R4155 VDD VDD.n1163 0.245437
R4156 VDD VDD.n215 0.245437
R4157 VDD VDD.n239 0.245437
R4158 VDD VDD.n553 0.245437
R4159 VDD.n575 VDD 0.245437
R4160 VDD VDD.n487 0.245437
R4161 VDD VDD.n579 0.245437
R4162 VDD VDD.n1381 0.245437
R4163 VDD VDD.n2310 0.245437
R4164 VDD VDD.n2064 0.245437
R4165 VDD.n2069 VDD 0.245437
R4166 VDD.n1682 VDD 0.245437
R4167 VDD VDD.n1685 0.245437
R4168 VDD.n902 VDD.n889 0.244844
R4169 VDD.n1544 VDD.n1543 0.243929
R4170 VDD.n835 VDD.n834 0.243929
R4171 VDD.n1875 VDD.n1874 0.243929
R4172 VDD.n2213 VDD.n2212 0.243929
R4173 VDD.n1653 VDD.n1652 0.243929
R4174 VDD.n2356 VDD.n179 0.240311
R4175 VDD.n2190 VDD.n1760 0.225771
R4176 VDD.n1059 VDD.n1058 0.225329
R4177 VDD.n666 VDD.n665 0.225329
R4178 VDD.n1013 VDD.n1012 0.225329
R4179 VDD.n2379 VDD.n2378 0.225329
R4180 VDD.n1242 VDD.n1241 0.225329
R4181 VDD.n221 VDD.n220 0.225329
R4182 VDD.n557 VDD.n556 0.225329
R4183 VDD.n1660 VDD.n1567 0.218719
R4184 VDD.n2469 VDD.n2468 0.217211
R4185 VDD.n2479 VDD.n2478 0.217211
R4186 VDD.n2474 VDD.n2473 0.217211
R4187 VDD.n1054 VDD.n1053 0.212555
R4188 VDD.n661 VDD.n628 0.212555
R4189 VDD.n1029 VDD.n383 0.212555
R4190 VDD.n2387 VDD.n2386 0.212555
R4191 VDD.n1248 VDD.n1114 0.212555
R4192 VDD.n215 VDD.n212 0.212555
R4193 VDD.n553 VDD.n552 0.212555
R4194 VDD.n1689 VDD 0.208873
R4195 VDD VDD.n1634 0.204624
R4196 VDD.n1690 VDD.n1554 0.202885
R4197 VDD.n803 VDD.n802 0.199201
R4198 VDD VDD.n2464 0.190753
R4199 VDD.n586 VDD 0.1901
R4200 VDD.n2221 VDD.n2220 0.189965
R4201 VDD.n2155 VDD.n2154 0.189965
R4202 VDD.n2294 VDD.n2293 0.189684
R4203 VDD.n1427 VDD.n1418 0.189684
R4204 VDD.n1448 VDD.n1439 0.189684
R4205 VDD.n2231 VDD.n1467 0.189684
R4206 VDD.n2272 VDD.n1461 0.189684
R4207 VDD.n2097 VDD.n2096 0.189684
R4208 VDD.n2109 VDD.n2108 0.189684
R4209 VDD.n2128 VDD.n2127 0.189684
R4210 VDD.n2144 VDD.n2143 0.189684
R4211 VDD.n2136 VDD.n2135 0.189684
R4212 VDD.n2304 VDD.n2303 0.187773
R4213 VDD.n2078 VDD.n2077 0.187773
R4214 VDD.n1634 VDD.n1586 0.1805
R4215 VDD.n2466 VDD.n2465 0.175943
R4216 VDD.n884 VDD.n878 0.174566
R4217 VDD.n2161 VDD.n2160 0.166887
R4218 VDD.n1890 VDD.n1767 0.1595
R4219 VDD.n1368 VDD.n1367 0.157922
R4220 VDD.n166 VDD.n162 0.1577
R4221 VDD.n324 VDD.n288 0.1577
R4222 VDD.n1343 VDD.n1342 0.1577
R4223 VDD.n1068 VDD.n1063 0.1577
R4224 VDD.n772 VDD.n771 0.1577
R4225 VDD.n738 VDD.n702 0.1577
R4226 VDD.n671 VDD.n670 0.1577
R4227 VDD.n1008 VDD.n1003 0.1577
R4228 VDD.n64 VDD.n56 0.1577
R4229 VDD.n2461 VDD.n45 0.1577
R4230 VDD.n2438 VDD.n2437 0.1577
R4231 VDD.n2374 VDD.n2369 0.1577
R4232 VDD.n1310 VDD.n1309 0.1577
R4233 VDD.n1288 VDD.n1287 0.1577
R4234 VDD.n1237 VDD.n1232 0.1577
R4235 VDD.n1214 VDD.n1213 0.1577
R4236 VDD.n1169 VDD.n1168 0.1577
R4237 VDD.n231 VDD.n230 0.1577
R4238 VDD.n561 VDD.n560 0.1577
R4239 VDD.n492 VDD.n491 0.1577
R4240 VDD.n584 VDD.n583 0.1577
R4241 VDD.n1677 VDD.n1676 0.1577
R4242 VDD.n341 VDD.n340 0.157022
R4243 VDD.n673 VDD.n644 0.157022
R4244 VDD.n1001 VDD.n399 0.157022
R4245 VDD.n2364 VDD.n2363 0.157022
R4246 VDD.n1230 VDD.n1128 0.157022
R4247 VDD.n259 VDD.n254 0.157022
R4248 VDD.n563 VDD.n512 0.157022
R4249 VDD.n1058 VDD.n351 0.155679
R4250 VDD.n665 VDD.n657 0.155679
R4251 VDD.n1016 VDD.n1013 0.155679
R4252 VDD.n2382 VDD.n2379 0.155679
R4253 VDD.n1245 VDD.n1242 0.155679
R4254 VDD.n220 VDD.n219 0.155679
R4255 VDD.n556 VDD.n555 0.155679
R4256 VDD.n2187 VDD.n1761 0.150448
R4257 VDD.n2183 VDD.n2182 0.1503
R4258 VDD.n2225 VDD.n2223 0.150192
R4259 VDD.n2151 VDD.n2149 0.150192
R4260 VDD.n1885 VDD.n1884 0.143178
R4261 VDD.n1062 VDD.n348 0.143147
R4262 VDD.n669 VDD.n654 0.143147
R4263 VDD.n1011 VDD.n1009 0.143147
R4264 VDD.n2377 VDD.n2375 0.143147
R4265 VDD.n1240 VDD.n1238 0.143147
R4266 VDD.n223 VDD.n222 0.143147
R4267 VDD.n559 VDD.n558 0.143147
R4268 VDD.n1317 VDD.n1316 0.14225
R4269 VDD.n2276 VDD 0.14101
R4270 VDD VDD.n2133 0.14101
R4271 VDD.n791 VDD 0.134375
R4272 VDD.n2181 VDD.n1763 0.132152
R4273 VDD VDD.n88 0.12875
R4274 VDD.n416 VDD 0.12875
R4275 VDD.n2408 VDD 0.12875
R4276 VDD.n1291 VDD 0.12875
R4277 VDD.n1195 VDD 0.12875
R4278 VDD.n1217 VDD 0.12875
R4279 VDD.n536 VDD 0.12875
R4280 VDD.n473 VDD 0.12875
R4281 VDD.n495 VDD 0.12875
R4282 VDD VDD.n1561 0.12875
R4283 VDD.n1891 VDD.n1890 0.128
R4284 VDD.n305 VDD.n304 0.127625
R4285 VDD.n1318 VDD.n1317 0.127625
R4286 VDD.n1048 VDD.n1047 0.127625
R4287 VDD.n716 VDD.n715 0.127625
R4288 VDD.n747 VDD.n746 0.127625
R4289 VDD.n790 VDD.n789 0.127625
R4290 VDD.n2451 VDD.n2450 0.127625
R4291 VDD.n2434 VDD.n2433 0.127625
R4292 VDD.n211 VDD.n205 0.127625
R4293 VDD.n867 VDD.n866 0.125816
R4294 VDD VDD.n375 0.124664
R4295 VDD.n1267 VDD 0.123125
R4296 VDD.n791 VDD.n619 0.122
R4297 VDD.n1268 VDD 0.122
R4298 VDD VDD.n1048 0.113
R4299 VDD.n789 VDD 0.113
R4300 VDD VDD.n2408 0.113
R4301 VDD VDD.n1113 0.113
R4302 VDD VDD.n211 0.113
R4303 VDD VDD.n536 0.113
R4304 VDD.n1059 VDD.n348 0.108884
R4305 VDD.n666 VDD.n654 0.108884
R4306 VDD.n1012 VDD.n1011 0.108884
R4307 VDD.n2378 VDD.n2377 0.108884
R4308 VDD.n1241 VDD.n1240 0.108884
R4309 VDD.n222 VDD.n221 0.108884
R4310 VDD.n558 VDD.n557 0.108884
R4311 VDD.n1455 VDD.n1454 0.1085
R4312 VDD.n2007 VDD.n2006 0.1085
R4313 VDD VDD.n181 0.100602
R4314 VDD.n2420 VDD.n2419 0.100415
R4315 VDD.n909 VDD.n889 0.100143
R4316 VDD.n2422 VDD 0.0988898
R4317 VDD.n966 VDD.n909 0.0985357
R4318 VDD.n1229 VDD.n180 0.0981271
R4319 VDD VDD.n1222 0.0966017
R4320 VDD.n1661 VDD.n1561 0.096125
R4321 VDD.n1223 VDD.n180 0.0935509
R4322 VDD.n1368 VDD 0.0918605
R4323 VDD.n2421 VDD.n2420 0.0897373
R4324 VDD.n140 VDD.n139 0.0859548
R4325 VDD.n682 VDD.n681 0.0859548
R4326 VDD.n406 VDD.n405 0.0859548
R4327 VDD.n175 VDD.n174 0.0859548
R4328 VDD.n1138 VDD.n1137 0.0859548
R4329 VDD.n267 VDD.n266 0.0859548
R4330 VDD.n503 VDD.n502 0.0859548
R4331 VDD.n2171 VDD.n1761 0.07625
R4332 VDD.n2472 VDD 0.07475
R4333 VDD.n2188 VDD.n2187 0.0745657
R4334 VDD.n1034 VDD.n375 0.0664514
R4335 VDD.n855 VDD.n846 0.0542576
R4336 VDD.n1486 VDD.n1477 0.0542576
R4337 VDD.n1499 VDD.n1490 0.0542576
R4338 VDD.n1949 VDD.n1940 0.0542576
R4339 VDD.n1936 VDD.n1927 0.0542576
R4340 VDD.n2330 VDD.n196 0.053063
R4341 VDD.n2331 VDD.n194 0.053063
R4342 VDD.n958 VDD.n942 0.053063
R4343 VDD.n957 VDD.n943 0.053063
R4344 VDD.n907 VDD.n891 0.053063
R4345 VDD.n908 VDD.n886 0.053063
R4346 VDD.n933 VDD.n917 0.053063
R4347 VDD.n920 VDD.n912 0.053063
R4348 VDD.n2350 VDD.n186 0.053063
R4349 VDD.n2351 VDD.n184 0.053063
R4350 VDD.n992 VDD.n977 0.053063
R4351 VDD.n980 VDD.n972 0.053063
R4352 VDD.n2320 VDD.n195 0.0526849
R4353 VDD.n2321 VDD.n193 0.0526849
R4354 VDD.n959 VDD.n940 0.0526849
R4355 VDD.n939 VDD.n937 0.0526849
R4356 VDD.n896 VDD.n894 0.0526849
R4357 VDD.n895 VDD.n885 0.0526849
R4358 VDD.n934 VDD.n913 0.0526849
R4359 VDD.n935 VDD.n911 0.0526849
R4360 VDD.n2339 VDD.n188 0.0526849
R4361 VDD.n2338 VDD.n189 0.0526849
R4362 VDD.n993 VDD.n973 0.0526849
R4363 VDD.n994 VDD.n971 0.0526849
R4364 VDD.n2329 VDD.n2328 0.050741
R4365 VDD.n949 VDD.n941 0.050741
R4366 VDD.n899 VDD.n898 0.050741
R4367 VDD.n932 VDD.n931 0.050741
R4368 VDD.n2342 VDD.n2341 0.050741
R4369 VDD.n991 VDD.n990 0.050741
R4370 VDD.n965 VDD.n964 0.0506887
R4371 VDD.n2326 VDD.n199 0.0470126
R4372 VDD.n2325 VDD.n2324 0.0470126
R4373 VDD.n952 VDD.n946 0.0470126
R4374 VDD.n954 VDD.n953 0.0470126
R4375 VDD.n906 VDD.n905 0.0470126
R4376 VDD.n901 VDD.n890 0.0470126
R4377 VDD.n929 VDD.n919 0.0470126
R4378 VDD.n928 VDD.n922 0.0470126
R4379 VDD.n2349 VDD.n2348 0.0470126
R4380 VDD.n2344 VDD.n185 0.0470126
R4381 VDD.n988 VDD.n979 0.0470126
R4382 VDD.n987 VDD.n982 0.0470126
R4383 VDD.n2263 VDD 0.0445816
R4384 VDD.n2140 VDD 0.0445816
R4385 VDD.n2194 VDD.n1727 0.0420385
R4386 VDD.n1554 VDD.n1525 0.0420385
R4387 VDD.n2313 VDD.n2312 0.0415127
R4388 VDD.n852 VDD.n846 0.0411256
R4389 VDD.n1483 VDD.n1477 0.0411256
R4390 VDD.n1496 VDD.n1490 0.0411256
R4391 VDD.n1946 VDD.n1940 0.0411256
R4392 VDD.n1933 VDD.n1927 0.0411256
R4393 VDD.n2230 VDD 0.0390714
R4394 VDD.n2145 VDD 0.0390714
R4395 VDD.n1472 VDD.n1471 0.0322647
R4396 VDD.n1954 VDD.n1953 0.0322647
R4397 VDD.n135 VDD.n133 0.03175
R4398 VDD.n677 VDD.n675 0.03175
R4399 VDD.n403 VDD.n400 0.03175
R4400 VDD.n172 VDD.n169 0.03175
R4401 VDD.n1135 VDD.n1132 0.03175
R4402 VDD.n262 VDD.n260 0.03175
R4403 VDD.n500 VDD.n497 0.03175
R4404 VDD.n1886 VDD.n1765 0.0316538
R4405 VDD.n2181 VDD.n2180 0.0316538
R4406 VDD.n2184 VDD.n2183 0.0316538
R4407 VDD.n902 VDD.n887 0.0302656
R4408 VDD.n314 VDD.n293 0.0301203
R4409 VDD.n1348 VDD.n273 0.0301203
R4410 VDD.n1050 VDD.n364 0.0301203
R4411 VDD.n728 VDD.n717 0.0301203
R4412 VDD.n777 VDD.n687 0.0301203
R4413 VDD.n788 VDD.n787 0.0301203
R4414 VDD.n1028 VDD.n385 0.0301203
R4415 VDD.n87 VDD.n86 0.0301203
R4416 VDD.n418 VDD.n417 0.0301203
R4417 VDD.n2449 VDD.n2448 0.0301203
R4418 VDD.n2432 VDD.n2431 0.0301203
R4419 VDD.n2399 VDD.n2398 0.0301203
R4420 VDD.n1304 VDD.n1292 0.0301203
R4421 VDD.n1282 VDD.n1270 0.0301203
R4422 VDD.n1262 VDD.n1261 0.0301203
R4423 VDD.n1208 VDD.n1196 0.0301203
R4424 VDD.n1219 VDD.n1218 0.0301203
R4425 VDD.n237 VDD.n236 0.0301203
R4426 VDD.n551 VDD.n537 0.0301203
R4427 VDD.n486 VDD.n474 0.0301203
R4428 VDD.n578 VDD.n496 0.0301203
R4429 VDD.n1684 VDD.n1662 0.0301203
R4430 VDD.n967 VDD.n887 0.0297969
R4431 VDD.n2185 VDD.n1763 0.0290882
R4432 VDD.n2337 VDD.n2336 0.0265377
R4433 VDD.n1034 VDD 0.0255962
R4434 VDD.n2195 VDD.n2194 0.0251429
R4435 VDD.n1554 VDD.n1553 0.0251429
R4436 VDD.n1474 VDD.n1472 0.0216225
R4437 VDD.n1955 VDD.n1954 0.0216225
R4438 VDD.n2345 VDD.n183 0.0212547
R4439 VDD.n925 VDD.n924 0.0208774
R4440 VDD.n956 VDD.n944 0.0208774
R4441 VDD.n1624 VDD.n1623 0.0203701
R4442 VDD.n1615 VDD.n1614 0.0203701
R4443 VDD.n1694 VDD.n1693 0.0203701
R4444 VDD.n1710 VDD.n1709 0.0203701
R4445 VDD.n1722 VDD.n1514 0.0203701
R4446 VDD.n860 VDD.n859 0.0203701
R4447 VDD.n839 VDD.n590 0.0203701
R4448 VDD.n813 VDD.n812 0.0203701
R4449 VDD.n804 VDD.n803 0.0203701
R4450 VDD.n1879 VDD.n1807 0.0203701
R4451 VDD.n1853 VDD.n1852 0.0203701
R4452 VDD.n1844 VDD.n1843 0.0203701
R4453 VDD.n2055 VDD.n2053 0.0203701
R4454 VDD.n1913 VDD.n1912 0.0203701
R4455 VDD.n1896 VDD.n1895 0.0203701
R4456 VDD.n2192 VDD.n2191 0.0203701
R4457 VDD.n1753 VDD.n1752 0.0203701
R4458 VDD.n2217 VDD.n1504 0.0203701
R4459 VDD.n1657 VDD.n1578 0.0203701
R4460 VDD.n1887 VDD.n1798 0.0202561
R4461 VDD.n2177 VDD.n1770 0.0185
R4462 VDD.n2179 VDD.n1764 0.018061
R4463 VDD.n2186 VDD.n1762 0.0164742
R4464 VDD.n817 VDD.n816 0.0162732
R4465 VDD.n1857 VDD.n1856 0.0162732
R4466 VDD.n1635 VDD.n1627 0.0162732
R4467 VDD.n2353 VDD.n182 0.0161604
R4468 VDD.n1620 VDD.n1619 0.0150714
R4469 VDD.n1611 VDD.n1610 0.0150714
R4470 VDD.n1701 VDD.n1700 0.0150714
R4471 VDD.n1717 VDD.n1716 0.0150714
R4472 VDD.n1545 VDD.n1541 0.0150714
R4473 VDD.n836 VDD.n832 0.0150714
R4474 VDD.n822 VDD.n821 0.0150714
R4475 VDD.n809 VDD.n808 0.0150714
R4476 VDD.n799 VDD.n798 0.0150714
R4477 VDD.n1876 VDD.n1872 0.0150714
R4478 VDD.n1862 VDD.n1861 0.0150714
R4479 VDD.n1849 VDD.n1848 0.0150714
R4480 VDD.n1840 VDD.n1839 0.0150714
R4481 VDD.n1920 VDD.n1919 0.0150714
R4482 VDD.n1903 VDD.n1902 0.0150714
R4483 VDD.n2200 VDD.n2199 0.0150714
R4484 VDD.n1758 VDD.n1757 0.0150714
R4485 VDD.n1749 VDD.n1748 0.0150714
R4486 VDD.n2214 VDD.n2210 0.0150714
R4487 VDD.n1551 VDD.n1550 0.0150714
R4488 VDD.n1654 VDD.n1650 0.0150714
R4489 VDD.n1640 VDD.n1639 0.0150714
R4490 VDD.n967 VDD.n888 0.0149643
R4491 VDD.n1535 VDD.n1534 0.014934
R4492 VDD.n828 VDD.n827 0.014934
R4493 VDD.n1868 VDD.n1867 0.014934
R4494 VDD.n2206 VDD.n2205 0.014934
R4495 VDD.n1646 VDD.n1645 0.014934
R4496 VDD.n2333 VDD.n2332 0.0144623
R4497 VDD.n2301 VDD.n2300 0.0138043
R4498 VDD.n2291 VDD.n2290 0.0138043
R4499 VDD.n1430 VDD.n1429 0.0138043
R4500 VDD.n2278 VDD.n1450 0.0138043
R4501 VDD.n2084 VDD.n2080 0.0138043
R4502 VDD.n2100 VDD.n2027 0.0138043
R4503 VDD.n2115 VDD.n2111 0.0138043
R4504 VDD.n2131 VDD.n2010 0.0138043
R4505 VDD.n2307 VDD.n2306 0.0136897
R4506 VDD.n2297 VDD.n2296 0.0136897
R4507 VDD.n2287 VDD.n2286 0.0136897
R4508 VDD.n1437 VDD.n1436 0.0136897
R4509 VDD.n2074 VDD.n2072 0.0136897
R4510 VDD.n2087 VDD.n2030 0.0136897
R4511 VDD.n2105 VDD.n2103 0.0136897
R4512 VDD.n2118 VDD.n2013 0.0136897
R4513 VDD.n384 VDD.n378 0.0135493
R4514 VDD.n2163 VDD.n2162 0.0133571
R4515 VDD.n2159 VDD.n2158 0.0133571
R4516 VDD.n2170 VDD.n1770 0.01325
R4517 VDD.n2166 VDD.n1781 0.0131446
R4518 VDD.n984 VDD.n983 0.0125755
R4519 VDD.n2182 VDD.n1764 0.0125732
R4520 VDD.n2178 VDD.n2177 0.0125
R4521 VDD.n1777 VDD.n1776 0.0124531
R4522 VDD.n1798 VDD.n1766 0.010378
R4523 VDD.n985 VDD.n984 0.00936793
R4524 VDD.n2178 VDD.n1767 0.008
R4525 VDD.n2171 VDD 0.008
R4526 VDD.n1269 VDD.n1268 0.00725
R4527 VDD.n2333 VDD.n191 0.00691509
R4528 VDD.n1267 VDD.n1113 0.006125
R4529 VDD VDD.n1033 0.00482692
R4530 VDD.n2353 VDD.n2352 0.00427358
R4531 VDD.n968 VDD.n967 0.00401562
R4532 VDD.n984 VDD.n190 0.00379268
R4533 VDD VDD.n1909 0.00292001
R4534 VDD VDD.n2469 0.00286842
R4535 VDD VDD.n2479 0.00286842
R4536 VDD VDD.n2474 0.00286842
R4537 VDD.n2321 VDD.n2318 0.00276891
R4538 VDD.n962 VDD.n939 0.00276891
R4539 VDD.n892 VDD.n885 0.00276891
R4540 VDD.n914 VDD.n911 0.00276891
R4541 VDD.n2334 VDD.n189 0.00276891
R4542 VDD.n974 VDD.n971 0.00276891
R4543 VDD.n969 VDD.n968 0.00214062
R4544 VDD.n2320 VDD.n2319 0.00213334
R4545 VDD.n961 VDD.n940 0.00213334
R4546 VDD.n894 VDD.n893 0.00213334
R4547 VDD.n915 VDD.n913 0.00213334
R4548 VDD.n188 VDD.n187 0.00213334
R4549 VDD.n975 VDD.n973 0.00213334
R4550 VDD.n967 VDD.n966 0.00210714
R4551 VDD.n1000 VDD 0.00202542
R4552 VDD VDD.n2421 0.00202542
R4553 VDD.n1223 VDD 0.00202542
R4554 VDD VDD.n564 0.00202542
R4555 VDD.n2324 VDD.n2323 0.00201261
R4556 VDD.n953 VDD.n948 0.00201261
R4557 VDD.n903 VDD.n901 0.00201261
R4558 VDD.n922 VDD.n921 0.00201261
R4559 VDD.n2346 VDD.n2344 0.00201261
R4560 VDD.n982 VDD.n981 0.00201261
R4561 VDD.n199 VDD.n198 0.00175581
R4562 VDD.n952 VDD.n951 0.00175581
R4563 VDD.n905 VDD.n904 0.00175581
R4564 VDD.n919 VDD.n918 0.00175581
R4565 VDD.n2348 VDD.n2347 0.00175581
R4566 VDD.n979 VDD.n978 0.00175581
R4567 VDD.n875 VDD 0.00175
R4568 VDD VDD.n1617 0.00173288
R4569 VDD.n1704 VDD 0.00173288
R4570 VDD.n1720 VDD 0.00173288
R4571 VDD VDD.n806 0.00173288
R4572 VDD VDD.n587 0.00173288
R4573 VDD VDD.n1846 0.00173288
R4574 VDD VDD.n1804 0.00173288
R4575 VDD.n1923 VDD 0.00173288
R4576 VDD.n1906 VDD 0.00173288
R4577 VDD VDD.n1755 0.00173288
R4578 VDD VDD.n1501 0.00173288
R4579 VDD VDD.n1567 0.00173288
R4580 VDD VDD.n1574 0.0017
R4581 VDD.n166 VDD 0.0017
R4582 VDD VDD.n324 0.0017
R4583 VDD.n1342 VDD 0.0017
R4584 VDD.n1068 VDD 0.0017
R4585 VDD.n771 VDD 0.0017
R4586 VDD VDD.n738 0.0017
R4587 VDD VDD.n671 0.0017
R4588 VDD.n1003 VDD 0.0017
R4589 VDD.n56 VDD 0.0017
R4590 VDD VDD.n2461 0.0017
R4591 VDD.n2437 VDD 0.0017
R4592 VDD.n2369 VDD 0.0017
R4593 VDD.n1310 VDD 0.0017
R4594 VDD VDD.n1288 0.0017
R4595 VDD.n1232 VDD 0.0017
R4596 VDD VDD.n1214 0.0017
R4597 VDD.n1168 VDD 0.0017
R4598 VDD VDD.n231 0.0017
R4599 VDD VDD.n561 0.0017
R4600 VDD VDD.n492 0.0017
R4601 VDD VDD.n584 0.0017
R4602 VDD.n1884 VDD 0.0017
R4603 VDD.n1677 VDD 0.0017
R4604 VDD VDD.n1624 0.00166883
R4605 VDD VDD.n1615 0.00166883
R4606 VDD.n1693 VDD 0.00166883
R4607 VDD.n1709 VDD 0.00166883
R4608 VDD.n1722 VDD 0.00166883
R4609 VDD.n860 VDD 0.00166883
R4610 VDD VDD.n839 0.00166883
R4611 VDD VDD.n813 0.00166883
R4612 VDD VDD.n804 0.00166883
R4613 VDD VDD.n1879 0.00166883
R4614 VDD VDD.n1853 0.00166883
R4615 VDD VDD.n1844 0.00166883
R4616 VDD VDD.n2055 0.00166883
R4617 VDD.n1912 VDD 0.00166883
R4618 VDD.n1895 VDD 0.00166883
R4619 VDD VDD.n2192 0.00166883
R4620 VDD VDD.n1753 0.00166883
R4621 VDD VDD.n2217 0.00166883
R4622 VDD VDD.n1657 0.00166883
R4623 VDD.n878 VDD 0.00165385
R4624 VDD.n2180 VDD.n1765 0.00165385
R4625 VDD.n2184 VDD.n1762 0.00165385
R4626 VDD VDD.n483 0.00163924
R4627 VDD VDD.n548 0.00163924
R4628 VDD VDD.n1279 0.00163924
R4629 VDD VDD.n2445 0.00163924
R4630 VDD VDD.n426 0.00163924
R4631 VDD.n1335 VDD 0.00163924
R4632 VDD.n320 VDD 0.00163924
R4633 VDD VDD.n312 0.00163924
R4634 VDD VDD.n1346 0.00163924
R4635 VDD.n1055 VDD 0.00163924
R4636 VDD VDD.n361 0.00163924
R4637 VDD.n864 VDD 0.00163924
R4638 VDD VDD.n725 0.00163924
R4639 VDD.n767 VDD 0.00163924
R4640 VDD.n734 VDD 0.00163924
R4641 VDD VDD.n775 0.00163924
R4642 VDD VDD.n784 0.00163924
R4643 VDD.n662 VDD 0.00163924
R4644 VDD VDD.n1025 0.00163924
R4645 VDD.n1017 VDD 0.00163924
R4646 VDD VDD.n83 0.00163924
R4647 VDD VDD.n67 0.00163924
R4648 VDD VDD.n51 0.00163924
R4649 VDD.n2465 VDD 0.00163924
R4650 VDD.n2441 VDD 0.00163924
R4651 VDD.n159 VDD 0.00163924
R4652 VDD VDD.n2427 0.00163924
R4653 VDD VDD.n2395 0.00163924
R4654 VDD VDD.n2383 0.00163924
R4655 VDD VDD.n1300 0.00163924
R4656 VDD.n1306 VDD 0.00163924
R4657 VDD.n1284 VDD 0.00163924
R4658 VDD VDD.n1258 0.00163924
R4659 VDD.n1249 VDD 0.00163924
R4660 VDD VDD.n1205 0.00163924
R4661 VDD.n1210 VDD 0.00163924
R4662 VDD.n1172 VDD 0.00163924
R4663 VDD.n1164 VDD 0.00163924
R4664 VDD.n216 VDD 0.00163924
R4665 VDD.n243 VDD 0.00163924
R4666 VDD.n554 VDD 0.00163924
R4667 VDD VDD.n574 0.00163924
R4668 VDD.n488 VDD 0.00163924
R4669 VDD.n580 VDD 0.00163924
R4670 VDD.n1382 VDD 0.00163924
R4671 VDD.n2311 VDD 0.00163924
R4672 VDD VDD.n2229 0.00163924
R4673 VDD.n2226 VDD 0.00163924
R4674 VDD.n2065 VDD 0.00163924
R4675 VDD VDD.n2068 0.00163924
R4676 VDD.n2147 VDD 0.00163924
R4677 VDD.n2152 VDD 0.00163924
R4678 VDD VDD.n1681 0.00163924
R4679 VDD.n1686 VDD 0.00163924
R4680 VDD.n2330 VDD.n195 0.00163445
R4681 VDD.n2331 VDD.n193 0.00163445
R4682 VDD.n959 VDD.n958 0.00163445
R4683 VDD.n957 VDD.n937 0.00163445
R4684 VDD.n896 VDD.n891 0.00163445
R4685 VDD.n895 VDD.n886 0.00163445
R4686 VDD.n934 VDD.n933 0.00163445
R4687 VDD.n935 VDD.n912 0.00163445
R4688 VDD.n2339 VDD.n186 0.00163445
R4689 VDD.n2338 VDD.n184 0.00163445
R4690 VDD.n993 VDD.n992 0.00163445
R4691 VDD.n994 VDD.n972 0.00163445
R4692 VDD.n2336 VDD.n2335 0.00163208
R4693 VDD.n305 VDD 0.001625
R4694 VDD.n1318 VDD 0.001625
R4695 VDD.n1047 VDD 0.001625
R4696 VDD.n715 VDD 0.001625
R4697 VDD.n747 VDD 0.001625
R4698 VDD VDD.n790 0.001625
R4699 VDD.n2451 VDD 0.001625
R4700 VDD VDD.n2434 0.001625
R4701 VDD.n205 VDD 0.001625
R4702 VDD.n2179 VDD.n1766 0.00159756
R4703 VDD.n2329 VDD.n197 0.00158434
R4704 VDD.n960 VDD.n941 0.00158434
R4705 VDD.n898 VDD.n897 0.00158434
R4706 VDD.n932 VDD.n916 0.00158434
R4707 VDD.n2341 VDD.n2340 0.00158434
R4708 VDD.n139 VDD.n136 0.00158434
R4709 VDD.n681 VDD.n678 0.00158434
R4710 VDD.n405 VDD.n404 0.00158434
R4711 VDD.n174 VDD.n173 0.00158434
R4712 VDD.n1137 VDD.n1136 0.00158434
R4713 VDD.n266 VDD.n263 0.00158434
R4714 VDD.n502 VDD.n501 0.00158434
R4715 VDD.n991 VDD.n976 0.00158434
R4716 VDD.n2195 VDD 0.00157143
R4717 VDD.n1553 VDD 0.00157143
R4718 VDD.n380 VDD.n379 0.00142783
R4719 VDD.n817 VDD 0.00142783
R4720 VDD.n1857 VDD 0.00142783
R4721 VDD.n1635 VDD 0.00142783
R4722 VDD VDD.n2294 0.00141837
R4723 VDD.n1418 VDD 0.00141837
R4724 VDD.n1439 VDD 0.00141837
R4725 VDD VDD.n1474 0.00141837
R4726 VDD.n2231 VDD 0.00141837
R4727 VDD VDD.n2234 0.00141837
R4728 VDD.n2264 VDD 0.00141837
R4729 VDD.n2267 VDD 0.00141837
R4730 VDD.n2268 VDD 0.00141837
R4731 VDD VDD.n2271 0.00141837
R4732 VDD.n2272 VDD 0.00141837
R4733 VDD VDD.n2275 0.00141837
R4734 VDD.n2097 VDD 0.00141837
R4735 VDD.n2108 VDD 0.00141837
R4736 VDD.n2128 VDD 0.00141837
R4737 VDD.n1955 VDD 0.00141837
R4738 VDD VDD.n2144 0.00141837
R4739 VDD.n2142 VDD 0.00141837
R4740 VDD.n2141 VDD 0.00141837
R4741 VDD VDD.n2139 0.00141837
R4742 VDD.n2138 VDD 0.00141837
R4743 VDD.n2137 VDD 0.00141837
R4744 VDD VDD.n2136 0.00141837
R4745 VDD.n2134 VDD 0.00141837
R4746 VDD VDD.n2304 0.00140909
R4747 VDD.n2077 VDD 0.00140909
R4748 VDD.n1033 VDD.n378 0.00136539
R4749 VDD VDD.n1620 0.00135714
R4750 VDD VDD.n1611 0.00135714
R4751 VDD.n1701 VDD 0.00135714
R4752 VDD.n1717 VDD 0.00135714
R4753 VDD.n1545 VDD 0.00135714
R4754 VDD.n836 VDD 0.00135714
R4755 VDD.n822 VDD 0.00135714
R4756 VDD VDD.n809 0.00135714
R4757 VDD VDD.n799 0.00135714
R4758 VDD.n1876 VDD 0.00135714
R4759 VDD.n1862 VDD 0.00135714
R4760 VDD VDD.n1849 0.00135714
R4761 VDD VDD.n1840 0.00135714
R4762 VDD.n1920 VDD 0.00135714
R4763 VDD.n1903 VDD 0.00135714
R4764 VDD.n2200 VDD 0.00135714
R4765 VDD VDD.n1758 0.00135714
R4766 VDD VDD.n1749 0.00135714
R4767 VDD.n2214 VDD 0.00135714
R4768 VDD.n1550 VDD 0.00135714
R4769 VDD.n1654 VDD 0.00135714
R4770 VDD.n1640 VDD 0.00135714
R4771 VDD VDD.n1535 0.00134906
R4772 VDD.n828 VDD 0.00134906
R4773 VDD.n1868 VDD 0.00134906
R4774 VDD.n2206 VDD 0.00134906
R4775 VDD.n1646 VDD 0.00134906
R4776 VDD.n2300 VDD 0.00128261
R4777 VDD.n2290 VDD 0.00128261
R4778 VDD VDD.n1430 0.00128261
R4779 VDD.n2278 VDD 0.00128261
R4780 VDD.n2084 VDD 0.00128261
R4781 VDD VDD.n2100 0.00128261
R4782 VDD.n2115 VDD 0.00128261
R4783 VDD VDD.n2131 0.00128261
R4784 VDD.n2306 VDD 0.00127586
R4785 VDD.n2296 VDD 0.00127586
R4786 VDD.n2286 VDD 0.00127586
R4787 VDD VDD.n1437 0.00127586
R4788 VDD.n2074 VDD 0.00127586
R4789 VDD VDD.n2087 0.00127586
R4790 VDD.n2105 VDD 0.00127586
R4791 VDD VDD.n2118 0.00127586
R4792 VDD.n1314 VDD 0.00126271
R4793 VDD.n780 VDD 0.00126271
R4794 VDD.n1351 VDD 0.00126271
R4795 VDD.n2162 VDD 0.0012563
R4796 VDD.n2158 VDD 0.0012563
R4797 VDD.n923 VDD.n910 0.00125472
R4798 VDD.n983 VDD.n970 0.00125472
R4799 VDD.n963 VDD.n938 0.00125472
R4800 VDD.n2317 VDD.n2316 0.00125472
R4801 VDD VDD.n2170 0.00125
R4802 VDD.n2166 VDD 0.0012438
R4803 VDD.n1777 VDD 0.00120312
R4804 VDD.n2337 VDD.n182 0.00106604
R4805 VDD.n924 VDD.n923 0.00106604
R4806 VDD.n926 VDD.n179 0.00106604
R4807 VDD.n2352 VDD.n183 0.00106604
R4808 VDD.n944 VDD.n938 0.00106604
R4809 VDD.n947 VDD.n945 0.00106604
R4810 VDD.n2316 VDD.n191 0.00106604
R4811 VDD.n2326 VDD.n196 0.000878151
R4812 VDD.n2325 VDD.n194 0.000878151
R4813 VDD.n946 VDD.n942 0.000878151
R4814 VDD.n954 VDD.n943 0.000878151
R4815 VDD.n907 VDD.n906 0.000878151
R4816 VDD.n908 VDD.n890 0.000878151
R4817 VDD.n929 VDD.n917 0.000878151
R4818 VDD.n928 VDD.n920 0.000878151
R4819 VDD.n2350 VDD.n2349 0.000878151
R4820 VDD.n2351 VDD.n185 0.000878151
R4821 VDD.n988 VDD.n977 0.000878151
R4822 VDD.n987 VDD.n980 0.000878151
R4823 VDD.n936 VDD.n910 0.000877358
R4824 VDD.n927 VDD.n925 0.000877358
R4825 VDD.n927 VDD.n926 0.000877358
R4826 VDD.n995 VDD.n970 0.000877358
R4827 VDD.n986 VDD.n985 0.000877358
R4828 VDD.n964 VDD.n963 0.000877358
R4829 VDD.n956 VDD.n955 0.000877358
R4830 VDD.n955 VDD.n945 0.000877358
R4831 VDD.n2317 VDD.n2315 0.000877358
R4832 VDD.n2332 VDD.n192 0.000877358
R4833 VDD.n2322 VDD.n192 0.000877358
R4834 VDD.n2328 VDD.n2327 0.000861446
R4835 VDD.n950 VDD.n949 0.000861446
R4836 VDD.n900 VDD.n899 0.000861446
R4837 VDD.n931 VDD.n930 0.000861446
R4838 VDD.n2343 VDD.n2342 0.000861446
R4839 VDD.n990 VDD.n989 0.000861446
R4840 CLK.t40 CLK.t9 47.8944
R4841 CLK.t28 CLK.t119 47.8944
R4842 CLK.t78 CLK.t126 47.8944
R4843 CLK.t13 CLK.t66 47.8944
R4844 CLK.t70 CLK.t107 47.8944
R4845 CLK.t8 CLK.t114 47.8944
R4846 CLK.t99 CLK.t22 47.8944
R4847 CLK.t27 CLK.t6 47.8944
R4848 CLK.t35 CLK.t23 47.8944
R4849 CLK.t87 CLK.t2 47.8944
R4850 CLK.t10 CLK.t74 47.8944
R4851 CLK.t24 CLK.t97 47.8944
R4852 CLK.t21 CLK.t112 44.058
R4853 CLK.t106 CLK.t61 44.058
R4854 CLK.t33 CLK.t125 44.058
R4855 CLK.t80 CLK.t63 44.058
R4856 CLK.t102 CLK.t92 44.058
R4857 CLK.t105 CLK.t94 44.058
R4858 CLK.t84 CLK.t45 44.058
R4859 CLK.t110 CLK.t118 44.058
R4860 CLK.n43 CLK.t108 38.8649
R4861 CLK.n34 CLK.t50 38.8649
R4862 CLK.n32 CLK.t116 38.8649
R4863 CLK.n31 CLK.t117 38.8649
R4864 CLK.n36 CLK.t30 38.8649
R4865 CLK.n38 CLK.t42 38.8649
R4866 CLK.n28 CLK.t39 38.8649
R4867 CLK.n5 CLK.t54 38.8649
R4868 CLK.n16 CLK.t90 38.7949
R4869 CLK.n15 CLK.t43 38.7949
R4870 CLK.n20 CLK.t3 38.7949
R4871 CLK.n19 CLK.t36 38.7949
R4872 CLK.n8 CLK.t29 38.7949
R4873 CLK.n9 CLK.t115 38.7949
R4874 CLK.n49 CLK.t58 38.7949
R4875 CLK.n50 CLK.t53 38.7949
R4876 CLK.n57 CLK.t51 38.7949
R4877 CLK.n56 CLK.t89 38.7949
R4878 CLK.n62 CLK.t77 38.7949
R4879 CLK.n61 CLK.t34 38.7949
R4880 CLK.n67 CLK.t81 38.7949
R4881 CLK.n66 CLK.t67 38.7949
R4882 CLK.n79 CLK.t12 38.7949
R4883 CLK.n78 CLK.t16 38.7949
R4884 CLK.n75 CLK.t113 38.7949
R4885 CLK.n74 CLK.t122 38.7949
R4886 CLK.n69 CLK.t25 38.7949
R4887 CLK.n70 CLK.t120 38.7949
R4888 CLK.n86 CLK.t65 38.7949
R4889 CLK.n87 CLK.t109 38.7949
R4890 CLK.n2 CLK.t101 38.7949
R4891 CLK.n1 CLK.t11 38.7949
R4892 CLK.n22 CLK.t59 36.2535
R4893 CLK.n59 CLK.t60 36.2535
R4894 CLK.n4 CLK.t17 36.2535
R4895 CLK.n73 CLK.t55 36.1638
R4896 CLK.n16 CLK.n15 31.4949
R4897 CLK.n20 CLK.n19 31.4949
R4898 CLK.n9 CLK.n8 31.4949
R4899 CLK.n50 CLK.n49 31.4949
R4900 CLK.n57 CLK.n56 31.4949
R4901 CLK.n62 CLK.n61 31.4949
R4902 CLK.n67 CLK.n66 31.4949
R4903 CLK.n79 CLK.n78 31.4949
R4904 CLK.n75 CLK.n74 31.4949
R4905 CLK.n70 CLK.n69 31.4949
R4906 CLK.n87 CLK.n86 31.4949
R4907 CLK.n2 CLK.n1 31.4949
R4908 CLK.t108 CLK.t21 28.6791
R4909 CLK.t50 CLK.t106 28.6791
R4910 CLK.t116 CLK.t33 28.6791
R4911 CLK.t117 CLK.t80 28.6791
R4912 CLK.t30 CLK.t102 28.6791
R4913 CLK.t42 CLK.t105 28.6791
R4914 CLK.t39 CLK.t84 28.6791
R4915 CLK.t54 CLK.t110 28.6791
R4916 CLK.n18 CLK.t62 26.9781
R4917 CLK.n18 CLK.t111 26.9781
R4918 CLK.n11 CLK.t103 26.9781
R4919 CLK.n11 CLK.t48 26.9781
R4920 CLK.n52 CLK.t72 26.9781
R4921 CLK.n52 CLK.t88 26.9781
R4922 CLK.n55 CLK.t95 26.9781
R4923 CLK.n55 CLK.t4 26.9781
R4924 CLK.n77 CLK.t75 26.9781
R4925 CLK.n77 CLK.t20 26.9781
R4926 CLK.n72 CLK.t79 26.9781
R4927 CLK.n72 CLK.t31 26.9781
R4928 CLK.n89 CLK.t91 26.9781
R4929 CLK.n89 CLK.t1 26.9781
R4930 CLK.n0 CLK.t71 26.9781
R4931 CLK.n0 CLK.t83 26.9781
R4932 CLK.n81 CLK.t19 20.269
R4933 CLK.n12 CLK.t93 20.2675
R4934 CLK.n53 CLK.t18 20.2675
R4935 CLK.n90 CLK.t15 20.2675
R4936 CLK.n17 CLK.t127 17.9416
R4937 CLK.n21 CLK.t121 17.9416
R4938 CLK.n10 CLK.t123 17.9416
R4939 CLK.n51 CLK.t100 17.9416
R4940 CLK.n58 CLK.t14 17.9416
R4941 CLK.n63 CLK.t38 17.9416
R4942 CLK.n68 CLK.t41 17.9416
R4943 CLK.n80 CLK.t68 17.9416
R4944 CLK.n71 CLK.t52 17.9416
R4945 CLK.n88 CLK.t96 17.9416
R4946 CLK.n3 CLK.t56 17.9416
R4947 CLK.n76 CLK.t86 17.6937
R4948 CLK.n41 CLK.n40 17.1932
R4949 CLK.n83 CLK 16.3788
R4950 CLK.n40 CLK.n39 14.7225
R4951 CLK.n84 CLK.n83 14.5859
R4952 CLK.n17 CLK.t40 11.957
R4953 CLK.n21 CLK.t28 11.957
R4954 CLK.n10 CLK.t78 11.957
R4955 CLK.n51 CLK.t13 11.957
R4956 CLK.n58 CLK.t70 11.957
R4957 CLK.n63 CLK.t8 11.957
R4958 CLK.n68 CLK.t99 11.957
R4959 CLK.n80 CLK.t27 11.957
R4960 CLK.n71 CLK.t87 11.957
R4961 CLK.n88 CLK.t10 11.957
R4962 CLK.n3 CLK.t24 11.957
R4963 CLK.n23 CLK 10.8825
R4964 CLK.n64 CLK 10.1333
R4965 CLK.n65 CLK.n64 9.77639
R4966 CLK.n48 CLK 9.69699
R4967 CLK.n27 CLK.n26 9.56219
R4968 CLK CLK.n47 9.4671
R4969 CLK.n76 CLK.t35 9.20812
R4970 CLK.n48 CLK.n27 8.87892
R4971 CLK.n60 CLK.n54 8.06233
R4972 CLK.n92 CLK.n91 8.06233
R4973 CLK.n92 CLK 7.82643
R4974 CLK.n43 CLK.t104 7.3005
R4975 CLK.n34 CLK.t44 7.3005
R4976 CLK.n32 CLK.t124 7.3005
R4977 CLK.n31 CLK.t0 7.3005
R4978 CLK.n36 CLK.t69 7.3005
R4979 CLK.n38 CLK.t82 7.3005
R4980 CLK.n28 CLK.t49 7.3005
R4981 CLK.n15 CLK.t85 7.3005
R4982 CLK.t127 CLK.n16 7.3005
R4983 CLK.n19 CLK.t76 7.3005
R4984 CLK.t121 CLK.n20 7.3005
R4985 CLK.t59 CLK.n18 7.3005
R4986 CLK.n8 CLK.t32 7.3005
R4987 CLK.t123 CLK.n9 7.3005
R4988 CLK.t93 CLK.n11 7.3005
R4989 CLK.n5 CLK.t57 7.3005
R4990 CLK.n49 CLK.t26 7.3005
R4991 CLK.t100 CLK.n50 7.3005
R4992 CLK.t18 CLK.n52 7.3005
R4993 CLK.n56 CLK.t5 7.3005
R4994 CLK.t14 CLK.n57 7.3005
R4995 CLK.t60 CLK.n55 7.3005
R4996 CLK.n61 CLK.t7 7.3005
R4997 CLK.t38 CLK.n62 7.3005
R4998 CLK.n66 CLK.t73 7.3005
R4999 CLK.t41 CLK.n67 7.3005
R5000 CLK.n78 CLK.t46 7.3005
R5001 CLK.t68 CLK.n79 7.3005
R5002 CLK.t19 CLK.n77 7.3005
R5003 CLK.n74 CLK.t64 7.3005
R5004 CLK.t86 CLK.n75 7.3005
R5005 CLK.n69 CLK.t98 7.3005
R5006 CLK.t52 CLK.n70 7.3005
R5007 CLK.t55 CLK.n72 7.3005
R5008 CLK.n86 CLK.t37 7.3005
R5009 CLK.t96 CLK.n87 7.3005
R5010 CLK.t15 CLK.n89 7.3005
R5011 CLK.n1 CLK.t47 7.3005
R5012 CLK.t56 CLK.n2 7.3005
R5013 CLK.t17 CLK.n0 7.3005
R5014 CLK.n42 CLK.n41 6.44858
R5015 CLK.n83 CLK.n82 6.20325
R5016 CLK CLK.n17 5.96162
R5017 CLK CLK.n63 5.96162
R5018 CLK CLK.n68 5.96162
R5019 CLK.n14 CLK.n13 5.77702
R5020 CLK.n22 CLK.n21 5.77618
R5021 CLK.n59 CLK.n58 5.77618
R5022 CLK.n81 CLK.n80 5.77618
R5023 CLK.n4 CLK.n3 5.77618
R5024 CLK.n12 CLK.n10 5.67753
R5025 CLK.n53 CLK.n51 5.67753
R5026 CLK.n73 CLK.n71 5.67753
R5027 CLK.n90 CLK.n88 5.67753
R5028 CLK CLK.n43 5.27587
R5029 CLK CLK.n34 5.27587
R5030 CLK CLK.n32 5.27587
R5031 CLK CLK.n31 5.27587
R5032 CLK CLK.n36 5.27587
R5033 CLK CLK.n38 5.27587
R5034 CLK CLK.n28 5.27587
R5035 CLK CLK.n5 5.27587
R5036 CLK.n82 CLK 4.72813
R5037 CLK CLK.n76 4.68152
R5038 CLK.n46 CLK.n45 4.5005
R5039 CLK.n14 CLK.n7 4.5005
R5040 CLK.n65 CLK.n48 4.17208
R5041 CLK.n33 CLK 4.13571
R5042 CLK.n40 CLK.n37 3.87524
R5043 CLK.n82 CLK 3.82364
R5044 CLK.n27 CLK.n6 3.77382
R5045 CLK.n35 CLK.n33 3.07781
R5046 CLK.n47 CLK.n29 2.63121
R5047 CLK.n44 CLK 2.58323
R5048 CLK.n47 CLK.n46 2.37292
R5049 CLK.n33 CLK 2.26896
R5050 CLK.n26 CLK.n25 2.251
R5051 CLK.n24 CLK.n7 2.24958
R5052 CLK.n42 CLK.n30 2.24324
R5053 CLK.n85 CLK.n65 1.87775
R5054 CLK.n35 CLK 1.52886
R5055 CLK.n24 CLK.n23 1.50904
R5056 CLK.n45 CLK.n44 1.5081
R5057 CLK CLK.n85 1.33289
R5058 CLK.n41 CLK.n35 1.23732
R5059 CLK.n85 CLK.n84 1.08658
R5060 CLK.n23 CLK 0.81937
R5061 CLK.n60 CLK 0.81937
R5062 CLK CLK.n92 0.81937
R5063 CLK.n64 CLK.n60 0.749691
R5064 CLK.n84 CLK 0.473978
R5065 CLK CLK.n73 0.187712
R5066 CLK CLK.n22 0.185948
R5067 CLK CLK.n59 0.185948
R5068 CLK CLK.n4 0.185948
R5069 CLK CLK.n81 0.183616
R5070 CLK.n37 CLK 0.183172
R5071 CLK CLK.n12 0.182986
R5072 CLK CLK.n53 0.182986
R5073 CLK CLK.n90 0.182986
R5074 CLK.n39 CLK 0.141537
R5075 CLK.n13 CLK 0.0449156
R5076 CLK.n54 CLK 0.0449156
R5077 CLK.n91 CLK 0.0449156
R5078 CLK.n13 CLK 0.0332273
R5079 CLK.n54 CLK 0.0332273
R5080 CLK.n91 CLK 0.0332273
R5081 CLK.n39 CLK 0.0329
R5082 CLK.n46 CLK.n30 0.0316538
R5083 CLK.n25 CLK.n14 0.0267025
R5084 CLK.n45 CLK.n42 0.017677
R5085 CLK.n29 CLK 0.0123421
R5086 CLK.n6 CLK 0.01175
R5087 CLK.n29 CLK 0.0111579
R5088 CLK.n6 CLK 0.010625
R5089 CLK.n26 CLK.n7 0.00645454
R5090 CLK.n37 CLK 0.00517532
R5091 CLK.n25 CLK.n24 0.0038463
R5092 CLK.n44 CLK.n30 0.00176987
R5093 VSS.n2960 VSS.n2959 7.02327e+06
R5094 VSS.t1189 VSS.t816 41809.4
R5095 VSS.t1137 VSS.t402 41809.4
R5096 VSS.t1132 VSS.t198 41809.4
R5097 VSS.t1443 VSS.t203 41809.4
R5098 VSS.n3737 VSS.t810 24773.8
R5099 VSS.n3738 VSS.n3737 21563.7
R5100 VSS.n1157 VSS.n1156 18483.1
R5101 VSS.n4244 VSS.n4243 13993.8
R5102 VSS.n5499 VSS.n5498 13611.1
R5103 VSS.n5436 VSS.n61 12047.2
R5104 VSS.n5017 VSS.n5016 12047.2
R5105 VSS.n1332 VSS.n1331 8086.33
R5106 VSS.n5499 VSS.n3 8008.43
R5107 VSS.n5496 VSS.n4 7098.75
R5108 VSS.t134 VSS.t1206 6847.71
R5109 VSS.t125 VSS.t1198 6847.71
R5110 VSS.t238 VSS.t829 6829.13
R5111 VSS.t839 VSS.t516 6829.13
R5112 VSS.n2928 VSS.n2927 5649.3
R5113 VSS.n5496 VSS.n5495 5241.73
R5114 VSS.n4338 VSS.n1723 4962.02
R5115 VSS.n4334 VSS.n4333 4922.24
R5116 VSS.n2497 VSS.t1526 4530.79
R5117 VSS.n2929 VSS.n2928 4291.67
R5118 VSS.n2495 VSS.n2494 3845.48
R5119 VSS.n42 VSS.n40 3818.95
R5120 VSS.n2931 VSS.n3 3720.83
R5121 VSS.n1645 VSS.n1643 3443.07
R5122 VSS.n5497 VSS.t1285 3046.22
R5123 VSS.n2959 VSS.t1368 3012.77
R5124 VSS.t1526 VSS.t1523 2881.77
R5125 VSS.t814 VSS.t1007 2827.3
R5126 VSS.n2780 VSS.t514 2685.77
R5127 VSS.t1231 VSS.t739 2456.82
R5128 VSS.t1347 VSS.t146 2368.09
R5129 VSS.t523 VSS.t497 2166.67
R5130 VSS.t1002 VSS.t1003 2166.67
R5131 VSS.t412 VSS.t348 2166.67
R5132 VSS.t187 VSS.t189 2166.67
R5133 VSS.t293 VSS.t200 2166.67
R5134 VSS.t685 VSS.t529 2166.67
R5135 VSS.t143 VSS.t100 2166.67
R5136 VSS.t267 VSS.t268 2166.67
R5137 VSS.t170 VSS.t1278 2166.67
R5138 VSS.t328 VSS.t109 2166.67
R5139 VSS.t309 VSS.t509 2166.67
R5140 VSS.t1383 VSS.t330 2166.67
R5141 VSS.t874 VSS.t703 2166.67
R5142 VSS.t299 VSS.t994 2166.67
R5143 VSS.t162 VSS.t518 2166.67
R5144 VSS.t1024 VSS.t340 2166.67
R5145 VSS.t304 VSS.t281 2166.67
R5146 VSS.t1006 VSS.t338 2166.67
R5147 VSS.t160 VSS.t92 2166.67
R5148 VSS.t306 VSS.t307 2166.67
R5149 VSS.t85 VSS.t359 2166.67
R5150 VSS.t425 VSS.t78 2166.67
R5151 VSS.t298 VSS.t1067 2072.98
R5152 VSS.n1333 VSS.n1332 1851.17
R5153 VSS.t810 VSS.t522 1791.59
R5154 VSS.n5382 VSS.t858 1779.25
R5155 VSS.n5126 VSS.t849 1779.25
R5156 VSS.n2821 VSS.n2820 1769.44
R5157 VSS.t629 VSS.t715 1701.21
R5158 VSS.t1162 VSS.t1472 1701.21
R5159 VSS.t595 VSS.t1500 1701.21
R5160 VSS.t1389 VSS.t576 1701.21
R5161 VSS.t603 VSS.t1174 1701.21
R5162 VSS.t387 VSS.t1051 1701.21
R5163 VSS.t716 VSS.t591 1699.79
R5164 VSS.t1498 VSS.t666 1699.79
R5165 VSS.t1173 VSS.t618 1699.79
R5166 VSS.t1047 VSS.t386 1699.79
R5167 VSS.n4154 VSS.t806 1584.15
R5168 VSS.t858 VSS.t855 1549.67
R5169 VSS.t849 VSS.t846 1549.67
R5170 VSS.n2932 VSS.n2931 1515.27
R5171 VSS.n1331 VSS.t1236 1506.44
R5172 VSS.t119 VSS.t120 1485.71
R5173 VSS.n1323 VSS.t1222 1374.84
R5174 VSS.t987 VSS.n5436 1374.11
R5175 VSS.n5017 VSS.t992 1374.11
R5176 VSS.n5498 VSS.n5497 1342.09
R5177 VSS.n23 VSS.t587 1317.42
R5178 VSS.n2844 VSS.t1159 1317.42
R5179 VSS.t1510 VSS.n2561 1317.42
R5180 VSS.n2452 VSS.t1392 1317.42
R5181 VSS.t1179 VSS.n1112 1317.42
R5182 VSS.t1042 VSS.n4027 1317.42
R5183 VSS.n1331 VSS.t1212 1272.89
R5184 VSS.t845 VSS.t1349 1205.23
R5185 VSS.t854 VSS.t1338 1205.23
R5186 VSS.t1360 VSS.n3 1183.66
R5187 VSS.n5495 VSS.t896 1183.26
R5188 VSS.n4555 VSS.t1001 1153.55
R5189 VSS.t413 VSS.n4555 1153.55
R5190 VSS.t188 VSS.n4468 1153.55
R5191 VSS.n4441 VSS.t294 1153.55
R5192 VSS.t686 VSS.n4441 1153.55
R5193 VSS.n4382 VSS.t142 1153.55
R5194 VSS.n4416 VSS.t266 1153.55
R5195 VSS.n4416 VSS.t171 1153.55
R5196 VSS.n4519 VSS.t329 1153.55
R5197 VSS.n4995 VSS.t310 1153.55
R5198 VSS.n4274 VSS.t1384 1153.55
R5199 VSS.t875 VSS.n4274 1153.55
R5200 VSS.t161 VSS.n1731 1153.55
R5201 VSS.n2925 VSS.t1025 1153.55
R5202 VSS.n2925 VSS.t303 1153.55
R5203 VSS.n4313 VSS.t1005 1153.55
R5204 VSS.n4226 VSS.t159 1153.55
R5205 VSS.t305 VSS.n4226 1153.55
R5206 VSS.t86 VSS.n4956 1153.55
R5207 VSS.n4956 VSS.t426 1153.55
R5208 VSS.n1323 VSS.t730 1151.13
R5209 VSS.n5497 VSS.n5496 1126.94
R5210 VSS.n4967 VSS.t107 1088.19
R5211 VSS.t882 VSS.t49 1088.19
R5212 VSS.t300 VSS.t115 1088.19
R5213 VSS.t463 VSS.t460 1088.19
R5214 VSS.t708 VSS.t1028 1088.19
R5215 VSS.t409 VSS.t1352 1088.19
R5216 VSS.t532 VSS.t370 1088.19
R5217 VSS.t1375 VSS.t1373 1083.33
R5218 VSS.t522 VSS.t1375 1083.33
R5219 VSS.t1263 VSS.t1266 1083.33
R5220 VSS.t1266 VSS.t1001 1083.33
R5221 VSS.t317 VSS.t319 1083.33
R5222 VSS.t319 VSS.t413 1083.33
R5223 VSS.t357 VSS.t188 1083.33
R5224 VSS.t354 VSS.t357 1083.33
R5225 VSS.t294 VSS.t484 1083.33
R5226 VSS.t484 VSS.t486 1083.33
R5227 VSS.t1196 VSS.t686 1083.33
R5228 VSS.t1201 VSS.t1196 1083.33
R5229 VSS.t147 VSS.t150 1083.33
R5230 VSS.t142 VSS.t147 1083.33
R5231 VSS.t556 VSS.t667 1083.33
R5232 VSS.t667 VSS.t266 1083.33
R5233 VSS.t1304 VSS.t1302 1083.33
R5234 VSS.t171 VSS.t1304 1083.33
R5235 VSS.t288 VSS.t291 1083.33
R5236 VSS.t329 VSS.t288 1083.33
R5237 VSS.t167 VSS.t310 1083.33
R5238 VSS.t164 VSS.t167 1083.33
R5239 VSS.t1384 VSS.t872 1083.33
R5240 VSS.t872 VSS.t1167 1083.33
R5241 VSS.t137 VSS.t875 1083.33
R5242 VSS.t139 VSS.t137 1083.33
R5243 VSS.t442 VSS.t439 1083.33
R5244 VSS.t439 VSS.t298 1083.33
R5245 VSS.t372 VSS.t161 1083.33
R5246 VSS.t374 VSS.t372 1083.33
R5247 VSS.t6 VSS.t1025 1083.33
R5248 VSS.t3 VSS.t6 1083.33
R5249 VSS.t303 VSS.t1345 1083.33
R5250 VSS.t1345 VSS.t1341 1083.33
R5251 VSS.t333 VSS.t336 1083.33
R5252 VSS.t1005 VSS.t333 1083.33
R5253 VSS.t1412 VSS.t1410 1083.33
R5254 VSS.t159 VSS.t1412 1083.33
R5255 VSS.t55 VSS.t57 1083.33
R5256 VSS.t57 VSS.t305 1083.33
R5257 VSS.t1429 VSS.t1426 1083.33
R5258 VSS.t1426 VSS.t86 1083.33
R5259 VSS.t975 VSS.t978 1083.33
R5260 VSS.t978 VSS.t426 1083.33
R5261 VSS.n4336 VSS.n4331 1067.69
R5262 VSS.n1330 VSS.t735 977.444
R5263 VSS.n1314 VSS.t18 976.221
R5264 VSS.n1322 VSS.t737 976.221
R5265 VSS.n2928 VSS.n2858 960.069
R5266 VSS.t1060 VSS.t87 932.271
R5267 VSS.t194 VSS.t758 932.271
R5268 VSS.t756 VSS.t295 932.271
R5269 VSS.t922 VSS.t205 932.271
R5270 VSS.t245 VSS.t924 932.271
R5271 VSS.t909 VSS.t172 932.271
R5272 VSS.t1063 VSS.t156 932.271
R5273 VSS.t1297 VSS.n23 927.644
R5274 VSS.t254 VSS.n2844 927.644
R5275 VSS.n2561 VSS.t40 927.644
R5276 VSS.t869 VSS.n2452 927.644
R5277 VSS.n1112 VSS.t479 927.644
R5278 VSS.n4027 VSS.t860 927.644
R5279 VSS.t87 VSS.t215 905.265
R5280 VSS.t537 VSS.t194 905.265
R5281 VSS.t295 VSS.t152 905.265
R5282 VSS.t205 VSS.t177 905.265
R5283 VSS.t192 VSS.t245 905.265
R5284 VSS.t172 VSS.t94 905.265
R5285 VSS.t156 VSS.t89 905.265
R5286 VSS.n5382 VSS.n5381 898.529
R5287 VSS.t1224 VSS.n1330 895.99
R5288 VSS.n1314 VSS.t1226 894.87
R5289 VSS.t1238 VSS.n1322 894.87
R5290 VSS.t732 VSS.t735 879.699
R5291 VSS.t1233 VSS.t1224 879.699
R5292 VSS.t1236 VSS.t1233 879.699
R5293 VSS.t730 VSS.t732 879.414
R5294 VSS.t15 VSS.t13 878.598
R5295 VSS.t18 VSS.t15 878.598
R5296 VSS.t1226 VSS.t1228 878.598
R5297 VSS.t1228 VSS.t1231 878.598
R5298 VSS.t739 VSS.t741 878.598
R5299 VSS.t741 VSS.t737 878.598
R5300 VSS.t1240 VSS.t1238 878.598
R5301 VSS.t1222 VSS.t1240 878.598
R5302 VSS.t1080 VSS.t1055 863.47
R5303 VSS.t1067 VSS.n4969 859.471
R5304 VSS.t400 VSS.t222 849.053
R5305 VSS.t641 VSS.n2585 831.183
R5306 VSS.n1332 VSS.t414 824.217
R5307 VSS.n1642 VSS.t1215 824.146
R5308 VSS.n4331 VSS.t52 797.835
R5309 VSS.t414 VSS.t416 773.981
R5310 VSS.t471 VSS.t470 768.221
R5311 VSS.t1373 VSS.n3736 767.361
R5312 VSS.n4526 VSS.t1263 767.361
R5313 VSS.n4556 VSS.t317 767.361
R5314 VSS.n4469 VSS.t354 767.361
R5315 VSS.t486 VSS.n1010 767.361
R5316 VSS.n4442 VSS.t1201 767.361
R5317 VSS.t150 VSS.n4381 767.361
R5318 VSS.n4403 VSS.t556 767.361
R5319 VSS.t1302 VSS.n4415 767.361
R5320 VSS.t291 VSS.n4518 767.361
R5321 VSS.n326 VSS.t164 767.361
R5322 VSS.t1167 VSS.n4263 767.361
R5323 VSS.n4275 VSS.t139 767.361
R5324 VSS.n4970 VSS.t442 767.361
R5325 VSS.n1732 VSS.t374 767.361
R5326 VSS.n2889 VSS.t3 767.361
R5327 VSS.t1341 VSS.n2924 767.361
R5328 VSS.t336 VSS.n4195 767.361
R5329 VSS.t1410 VSS.n4225 767.361
R5330 VSS.n4227 VSS.t55 767.361
R5331 VSS.n4957 VSS.t1429 767.361
R5332 VSS.n533 VSS.t975 767.361
R5333 VSS.t1404 VSS.t1401 742.857
R5334 VSS.t38 VSS.t35 739.726
R5335 VSS.t657 VSS.n1136 735.85
R5336 VSS.t284 VSS.n4354 733.75
R5337 VSS.t776 VSS.t744 728.448
R5338 VSS.n86 VSS.t471 725.543
R5339 VSS.t248 VSS.t445 713.264
R5340 VSS.t1401 VSS.n2465 694.71
R5341 VSS.t35 VSS.n36 691.782
R5342 VSS.n4361 VSS.t1204 689.797
R5343 VSS.t270 VSS.t224 687.824
R5344 VSS.t999 VSS.t278 687.824
R5345 VSS.t174 VSS.t512 687.824
R5346 VSS.t695 VSS.t102 677.587
R5347 VSS.n4335 VSS.n4332 676.828
R5348 VSS.n2585 VSS.t578 656.51
R5349 VSS.n36 VSS.t717 625.524
R5350 VSS.n2937 VSS.t1473 625.524
R5351 VSS.n2465 VSS.t594 625.524
R5352 VSS.t570 VSS.n1086 625.524
R5353 VSS.n4053 VSS.t380 625.524
R5354 VSS.n4543 VSS.t49 597.375
R5355 VSS.n4397 VSS.t300 597.375
R5356 VSS.t460 VSS.n4458 597.375
R5357 VSS.n4997 VSS.t708 597.375
R5358 VSS.n2916 VSS.t409 597.375
R5359 VSS.t370 VSS.n4311 597.375
R5360 VSS.t107 VSS.n4966 597.375
R5361 VSS.n5497 VSS.t571 592.4
R5362 VSS.t1090 VSS.n4954 587.324
R5363 VSS.t560 VSS.n2460 543.255
R5364 VSS.t638 VSS.n31 542.461
R5365 VSS.n2466 VSS.t1404 526.191
R5366 VSS.n37 VSS.t38 523.973
R5367 VSS.n2858 VSS.t1288 515.982
R5368 VSS.t1423 VSS.n4360 500.765
R5369 VSS.n4555 VSS.t1062 496.349
R5370 VSS.n4441 VSS.t747 496.349
R5371 VSS.n4274 VSS.t918 496.349
R5372 VSS.n2925 VSS.t919 496.349
R5373 VSS.n4956 VSS.t1066 496.349
R5374 VSS.n1299 VSS.t1219 490.904
R5375 VSS.n2933 VSS.n2932 482.353
R5376 VSS.n4336 VSS.n4335 472.248
R5377 VSS.t1062 VSS.t598 466.135
R5378 VSS.t550 VSS.t785 466.135
R5379 VSS.t747 VSS.t619 466.135
R5380 VSS.t918 VSS.t568 466.135
R5381 VSS.t615 VSS.t910 466.135
R5382 VSS.t584 VSS.t1066 466.135
R5383 VSS.t580 VSS.t728 449.122
R5384 VSS.t587 VSS.t713 449.122
R5385 VSS.t1152 VSS.t1486 449.122
R5386 VSS.t1159 VSS.t1490 449.122
R5387 VSS.t1511 VSS.t583 449.122
R5388 VSS.t636 VSS.t1510 449.122
R5389 VSS.t1393 VSS.t663 449.122
R5390 VSS.t1392 VSS.t596 449.122
R5391 VSS.t1183 VSS.t563 449.122
R5392 VSS.t632 VSS.t1179 449.122
R5393 VSS.t1044 VSS.t397 449.122
R5394 VSS.t395 VSS.t1042 449.122
R5395 VSS.t725 VSS.t644 448.745
R5396 VSS.t717 VSS.t634 448.745
R5397 VSS.t1475 VSS.t1156 448.745
R5398 VSS.t652 VSS.t1499 448.745
R5399 VSS.t1506 VSS.t578 448.745
R5400 VSS.t649 VSS.t1388 448.745
R5401 VSS.t594 VSS.t1399 448.745
R5402 VSS.t588 VSS.t1182 448.745
R5403 VSS.t1180 VSS.t570 448.745
R5404 VSS.t388 VSS.t1050 448.745
R5405 VSS.t380 VSS.t1040 448.745
R5406 VSS.n4554 VSS.t630 425.134
R5407 VSS.t558 VSS.n4423 425.134
R5408 VSS.n4233 VSS.t625 425.134
R5409 VSS.n548 VSS.t621 425.134
R5410 VSS.t1336 VSS.n5382 423.776
R5411 VSS.t1334 VSS.n5126 423.776
R5412 VSS.n4440 VSS.t612 422.976
R5413 VSS.n4273 VSS.t548 422.976
R5414 VSS.n2882 VSS.t609 422.976
R5415 VSS.t1288 VSS.n2857 421.623
R5416 VSS.t674 VSS.t977 418.253
R5417 VSS.t986 VSS.t180 418.253
R5418 VSS.n86 VSS.t865 415.048
R5419 VSS.t1321 VSS.t711 405.483
R5420 VSS.t424 VSS.t1333 405.483
R5421 VSS.t196 VSS.t1466 405.483
R5422 VSS.t144 VSS.t1409 405.483
R5423 VSS.t398 VSS.t1456 405.483
R5424 VSS.t1009 VSS.t1406 405.483
R5425 VSS.t182 VSS.t1316 405.483
R5426 VSS.t444 VSS.t1344 405.483
R5427 VSS.t806 VSS.n4153 397.815
R5428 VSS.t865 VSS.t1541 389.784
R5429 VSS.t222 VSS.t1547 389.784
R5430 VSS.t25 VSS.t145 388.274
R5431 VSS.t215 VSS.t47 384.026
R5432 VSS.t324 VSS.t537 384.026
R5433 VSS.t152 VSS.t97 384.026
R5434 VSS.t177 VSS.t227 384.026
R5435 VSS.t406 VSS.t192 384.026
R5436 VSS.t94 VSS.t500 384.026
R5437 VSS.t89 VSS.t105 384.026
R5438 VSS.t1212 VSS.n1303 370.296
R5439 VSS.n4153 VSS.t814 369.399
R5440 VSS.t1031 VSS.t654 365.745
R5441 VSS.t867 VSS.t627 365.209
R5442 VSS.n4244 VSS.t914 364.224
R5443 VSS.t927 VSS.n4244 364.224
R5444 VSS.t973 VSS.n347 355.769
R5445 VSS.n1303 VSS.t1191 343.846
R5446 VSS.t261 VSS.t1307 334.925
R5447 VSS.t489 VSS.t365 334.925
R5448 VSS.t210 VSS.t322 334.925
R5449 VSS.t243 VSS.t1170 334.925
R5450 VSS.t1496 VSS.t0 334.925
R5451 VSS.t467 VSS.t1431 334.925
R5452 VSS.t1434 VSS.t155 334.925
R5453 VSS.t155 VSS.t154 334.925
R5454 VSS.n4544 VSS.t630 330.18
R5455 VSS.n4424 VSS.t558 330.18
R5456 VSS.n4448 VSS.t612 330.18
R5457 VSS.n4292 VSS.t548 330.18
R5458 VSS.n2914 VSS.t609 330.18
R5459 VSS.t625 VSS.n4211 330.18
R5460 VSS.t621 VSS.n547 330.18
R5461 VSS.n4334 VSS.t218 329.661
R5462 VSS.n4868 VSS.n4867 321.615
R5463 VSS.n4351 VSS.t20 318.06
R5464 VSS.n4982 VSS.t535 316.466
R5465 VSS.n333 VSS.t273 316.466
R5466 VSS.n4479 VSS.t69 316.293
R5467 VSS.n4489 VSS.t879 316.293
R5468 VSS.n3736 VSS.t523 315.973
R5469 VSS.n4526 VSS.t1002 315.973
R5470 VSS.n4556 VSS.t412 315.973
R5471 VSS.n4469 VSS.t187 315.973
R5472 VSS.n1010 VSS.t293 315.973
R5473 VSS.n4442 VSS.t685 315.973
R5474 VSS.n4381 VSS.t143 315.973
R5475 VSS.n4403 VSS.t267 315.973
R5476 VSS.n4415 VSS.t170 315.973
R5477 VSS.n4518 VSS.t328 315.973
R5478 VSS.n326 VSS.t309 315.973
R5479 VSS.n4263 VSS.t1383 315.973
R5480 VSS.n4275 VSS.t874 315.973
R5481 VSS.n4970 VSS.t299 315.973
R5482 VSS.n1732 VSS.t162 315.973
R5483 VSS.n2889 VSS.t1024 315.973
R5484 VSS.n2924 VSS.t304 315.973
R5485 VSS.n4195 VSS.t1006 315.973
R5486 VSS.n4225 VSS.t160 315.973
R5487 VSS.n4227 VSS.t306 315.973
R5488 VSS.n4957 VSS.t85 315.973
R5489 VSS.n533 VSS.t425 315.973
R5490 VSS.n5381 VSS.n5380 313.151
R5491 VSS.t230 VSS.t674 311.447
R5492 VSS.t688 VSS.t401 311.447
R5493 VSS.t180 VSS.t405 311.447
R5494 VSS.t876 VSS.t270 311.033
R5495 VSS.t278 VSS.t276 311.033
R5496 VSS.t512 VSS.t427 311.033
R5497 VSS.n4954 VSS.n4953 309.228
R5498 VSS.t102 VSS.t697 304.029
R5499 VSS.n5476 VSS.t722 293.971
R5500 VSS.n2834 VSS.t1483 293.971
R5501 VSS.n2560 VSS.t573 293.971
R5502 VSS.n2442 VSS.t565 293.971
R5503 VSS.n1111 VSS.t553 293.971
R5504 VSS.n4026 VSS.t383 293.971
R5505 VSS.n29 VSS.t660 293.724
R5506 VSS.n2850 VSS.t1147 293.724
R5507 VSS.n2458 VSS.t1396 293.724
R5508 VSS.n1130 VSS.t1176 293.724
R5509 VSS.t1052 VSS.n2428 293.724
R5510 VSS.t664 VSS.n9 291.248
R5511 VSS.t1160 VSS.n2829 291.248
R5512 VSS.n2556 VSS.t1508 291.248
R5513 VSS.t1385 VSS.n2437 291.248
R5514 VSS.n1107 VSS.t1187 291.248
R5515 VSS.n4022 VSS.t1048 291.248
R5516 VSS.t718 VSS.n20 291.005
R5517 VSS.n2841 VSS.t1481 291.005
R5518 VSS.n2576 VSS.t592 291.005
R5519 VSS.n2449 VSS.t601 291.005
R5520 VSS.n1127 VSS.t546 291.005
R5521 VSS.n4041 VSS.t377 291.005
R5522 VSS.t416 VSS.n1299 283.077
R5523 VSS.n87 VSS.n86 275.279
R5524 VSS.n4338 VSS.t251 257.755
R5525 VSS.n4968 VSS.t1437 248.093
R5526 VSS.t449 VSS.t238 245.748
R5527 VSS.t1195 VSS.t134 245.748
R5528 VSS.t516 VSS.t45 245.748
R5529 VSS.t1211 VSS.t125 245.748
R5530 VSS.t401 VSS.n2497 242.237
R5531 VSS.n4555 VSS.t1069 238.666
R5532 VSS.n4567 VSS.t1057 238.666
R5533 VSS.t748 VSS.n4416 238.666
R5534 VSS.n4441 VSS.t750 238.666
R5535 VSS.n2928 VSS.t937 238.666
R5536 VSS.t901 VSS.n2925 238.666
R5537 VSS.n4226 VSS.t935 238.666
R5538 VSS.n4274 VSS.t940 238.666
R5539 VSS.n4956 VSS.t1071 238.666
R5540 VSS.t20 VSS.n4350 237.25
R5541 VSS.n2496 VSS.t452 234.696
R5542 VSS.t492 VSS.n41 234.352
R5543 VSS.n5037 VSS.t1115 231.411
R5544 VSS.n5430 VSS.t1105 231.411
R5545 VSS.t981 VSS.n4359 228.292
R5546 VSS.t1057 VSS.t1083 224.138
R5547 VSS.t753 VSS.t776 224.138
R5548 VSS.t744 VSS.t774 224.138
R5549 VSS.t937 VSS.t907 224.138
R5550 VSS.t914 VSS.t948 224.138
R5551 VSS.t899 VSS.t927 224.138
R5552 VSS.t1086 VSS.t1090 224.138
R5553 VSS.t1013 VSS.n4382 223.282
R5554 VSS.n4468 VSS.t472 223.282
R5555 VSS.n4995 VSS.t1518 223.282
R5556 VSS.t502 VSS.n4313 223.282
R5557 VSS.n4566 VSS.t1069 223.101
R5558 VSS.n4417 VSS.t748 223.101
R5559 VSS.n4435 VSS.t750 223.101
R5560 VSS.n2926 VSS.t901 223.101
R5561 VSS.n4238 VSS.t935 223.101
R5562 VSS.t940 VSS.n4245 223.101
R5563 VSS.t1071 VSS.n4955 223.101
R5564 VSS.t1539 VSS.t400 222.05
R5565 VSS.n4647 VSS.n4646 217.635
R5566 VSS.n2466 VSS.t119 216.667
R5567 VSS.n37 VSS.t72 215.754
R5568 VSS.n4360 VSS.t1347 215.561
R5569 VSS.n4337 VSS.n4336 215.53
R5570 VSS.n5060 VSS.t430 210.934
R5571 VSS.n5429 VSS.t163 210.934
R5572 VSS.t803 VSS.n5499 209.091
R5573 VSS.n1643 VSS.n1642 206.477
R5574 VSS.n347 VSS.t996 205.528
R5575 VSS.n2586 VSS.t641 204.15
R5576 VSS.t1541 VSS.n51 203.915
R5577 VSS.t1547 VSS.n2503 203.915
R5578 VSS.t789 VSS.t261 201.575
R5579 VSS.t1017 VSS.t791 201.575
R5580 VSS.t1016 VSS.t796 201.575
R5581 VSS.t1110 VSS.t475 201.575
R5582 VSS.t1112 VSS.t474 201.575
R5583 VSS.t365 VSS.t769 201.575
R5584 VSS.t1073 VSS.t210 201.575
R5585 VSS.t1134 VSS.t1165 201.575
R5586 VSS.t1142 VSS.t1166 201.575
R5587 VSS.t824 VSS.t1514 201.575
R5588 VSS.t821 VSS.t1520 201.575
R5589 VSS.t943 VSS.t243 201.575
R5590 VSS.t894 VSS.t1314 201.575
R5591 VSS.t895 VSS.t1330 201.575
R5592 VSS.t925 VSS.t1496 201.575
R5593 VSS.t921 VSS.t64 201.575
R5594 VSS.t1459 VSS.t506 201.575
R5595 VSS.t1463 VSS.t505 201.575
R5596 VSS.t1075 VSS.t467 201.575
R5597 VSS.t1544 VSS.t1439 201.575
R5598 VSS.t1550 VSS.t1433 201.575
R5599 VSS.t977 VSS.t233 200.305
R5600 VSS.t1290 VSS.t986 200.305
R5601 VSS.n2495 VSS.t455 200.148
R5602 VSS.t495 VSS.n42 199.855
R5603 VSS.t1115 VSS.t449 196.597
R5604 VSS.t826 VSS.t1010 196.597
R5605 VSS.t430 VSS.t1195 196.597
R5606 VSS.t45 VSS.t1105 196.597
R5607 VSS.t841 VSS.t521 196.597
R5608 VSS.t163 VSS.t1211 196.597
R5609 VSS.t793 VSS.t803 196.364
R5610 VSS.n5115 VSS.t818 194.549
R5611 VSS.n5099 VSS.t1126 194.549
R5612 VSS.t1139 VSS.n131 194.549
R5613 VSS.t1445 VSS.n5386 194.549
R5614 VSS.t996 VSS.t213 193.017
R5615 VSS.n2858 VSS.t1357 190.905
R5616 VSS.n2586 VSS.t571 189.569
R5617 VSS.t233 VSS.t327 189.478
R5618 VSS.t343 VSS.t1290 189.478
R5619 VSS.t327 VSS.n51 185.869
R5620 VSS.n2503 VSS.t343 185.869
R5621 VSS.n4332 VSS.t692 185.817
R5622 VSS.t455 VSS.n2470 182.276
R5623 VSS.n43 VSS.t495 182.011
R5624 VSS.n1137 VSS.t657 180.736
R5625 VSS.n4568 VSS.n4567 178.944
R5626 VSS.n4355 VSS.t1261 178.757
R5627 VSS.t1338 VSS.n5384 178.431
R5628 VSS.n5125 VSS.t1349 178.431
R5629 VSS.t1021 VSS.t764 176.522
R5630 VSS.t786 VSS.t1018 176.522
R5631 VSS.t476 VSS.t761 176.522
R5632 VSS.t778 VSS.t364 176.522
R5633 VSS.t1064 VSS.t186 176.522
R5634 VSS.t1163 VSS.t1095 176.522
R5635 VSS.t930 VSS.t1515 176.522
R5636 VSS.t967 VSS.t700 176.522
R5637 VSS.t954 VSS.t889 176.522
R5638 VSS.t1354 VSS.t959 176.522
R5639 VSS.t62 VSS.t933 176.522
R5640 VSS.t507 VSS.t911 176.522
R5641 VSS.n4352 VSS.t122 176.161
R5642 VSS.n90 VSS.t260 175.911
R5643 VSS.n2502 VSS.t404 175.911
R5644 VSS.n4395 VSS.t1020 175.405
R5645 VSS.n4459 VSS.t363 175.405
R5646 VSS.n4520 VSS.t185 175.405
R5647 VSS.n4996 VSS.t701 175.405
R5648 VSS.t1355 VSS.n1698 175.405
R5649 VSS.t63 VSS.n4312 175.405
R5650 VSS.n5114 VSS.t311 174.071
R5651 VSS.n5100 VSS.t158 174.071
R5652 VSS.n175 VSS.t51 174.071
R5653 VSS.n5385 VSS.t302 174.071
R5654 VSS.n24 VSS.n19 174.06
R5655 VSS.n2845 VSS.n2840 174.06
R5656 VSS.n2570 VSS.n2568 174.06
R5657 VSS.n2453 VSS.n2448 174.06
R5658 VSS.n1121 VSS.n1119 174.06
R5659 VSS.n4036 VSS.n4035 174.06
R5660 VSS.t47 VSS.n4543 170.679
R5661 VSS.n4397 VSS.t324 170.679
R5662 VSS.n4458 VSS.t97 170.679
R5663 VSS.n4997 VSS.t227 170.679
R5664 VSS.n2916 VSS.t406 170.679
R5665 VSS.n4311 VSS.t500 170.679
R5666 VSS.n4966 VSS.t105 170.679
R5667 VSS.n4352 VSS.t25 168.971
R5668 VSS.n1137 VSS.t623 167.826
R5669 VSS.n5437 VSS.t983 161.492
R5670 VSS.t1120 VSS.n5435 161.492
R5671 VSS.n5015 VSS.t989 161.492
R5672 VSS.n5018 VSS.t1102 161.492
R5673 VSS.n2533 VSS.n2532 155.786
R5674 VSS.n2958 VSS.n2957 155.786
R5675 VSS.n2551 VSS.n2550 155.786
R5676 VSS.n5494 VSS.n5493 155.786
R5677 VSS.n1102 VSS.n1101 155.786
R5678 VSS.n4017 VSS.n4016 155.786
R5679 VSS.t679 VSS.t1297 155.022
R5680 VSS.t1300 VSS.t682 155.022
R5681 VSS.t82 VSS.t254 155.022
R5682 VSS.t257 VSS.t80 155.022
R5683 VSS.t40 VSS.t541 155.022
R5684 VSS.t43 VSS.t544 155.022
R5685 VSS.t1036 VSS.t869 155.022
R5686 VSS.t1555 VSS.t1034 155.022
R5687 VSS.t479 VSS.t421 155.022
R5688 VSS.t482 VSS.t419 155.022
R5689 VSS.t860 VSS.t436 155.022
R5690 VSS.t863 VSS.t434 155.022
R5691 VSS.n95 VSS.t839 149.957
R5692 VSS.t829 VSS.n5036 149.957
R5693 VSS.t251 VSS.n4337 148.856
R5694 VSS.n4884 VSS.n4883 148.571
R5695 VSS.n11 VSS.t720 146.986
R5696 VSS.n2830 VSS.t1489 146.986
R5697 VSS.n2557 VSS.t647 146.986
R5698 VSS.n2438 VSS.t604 146.986
R5699 VSS.n1108 VSS.t605 146.986
R5700 VSS.n4023 VSS.t379 146.986
R5701 VSS.n27 VSS.t645 146.863
R5702 VSS.n2848 VSS.t1157 146.863
R5703 VSS.n2577 VSS.t1505 146.863
R5704 VSS.n2456 VSS.t1387 146.863
R5705 VSS.n1128 VSS.t1186 146.863
R5706 VSS.n4040 VSS.t1043 146.863
R5707 VSS.t1206 VSS.n5059 146.01
R5708 VSS.t1198 VSS.n5428 146.01
R5709 VSS.n2533 VSS.t1380 145.042
R5710 VSS.t73 VSS.n2958 145.042
R5711 VSS.n2550 VSS.t526 145.042
R5712 VSS.t30 VSS.n5494 145.042
R5713 VSS.n1101 VSS.t314 145.042
R5714 VSS.n4016 VSS.t10 145.042
R5715 VSS.n5475 VSS.t608 144.263
R5716 VSS.t1155 VSS.n2835 144.263
R5717 VSS.n2562 VSS.t1504 144.263
R5718 VSS.t1390 VSS.n2443 144.263
R5719 VSS.n1113 VSS.t1175 144.263
R5720 VSS.n4028 VSS.t1039 144.263
R5721 VSS.t721 VSS.n30 144.143
R5722 VSS.n2851 VSS.t1474 144.143
R5723 VSS.n2580 VSS.t648 144.143
R5724 VSS.t646 VSS.n2459 144.143
R5725 VSS.n1131 VSS.t577 144.143
R5726 VSS.t391 VSS.n4052 144.143
R5727 VSS.n5310 VSS.n5309 143
R5728 VSS.n2532 VSS.t1283 142.356
R5729 VSS.n2957 VSS.t1371 142.356
R5730 VSS.n2551 VSS.t1366 142.356
R5731 VSS.n5493 VSS.t887 142.356
R5732 VSS.n1102 VSS.t1220 142.356
R5733 VSS.n4017 VSS.t1246 142.356
R5734 VSS.t720 VSS.t580 138.82
R5735 VSS.t715 VSS.t664 138.82
R5736 VSS.t722 VSS.t629 138.82
R5737 VSS.t1489 VSS.t1152 138.82
R5738 VSS.t1472 VSS.t1160 138.82
R5739 VSS.t1483 VSS.t1162 138.82
R5740 VSS.t1490 VSS.t1155 138.82
R5741 VSS.t647 VSS.t1511 138.82
R5742 VSS.t1508 VSS.t595 138.82
R5743 VSS.t1500 VSS.t573 138.82
R5744 VSS.t1504 VSS.t636 138.82
R5745 VSS.t604 VSS.t1393 138.82
R5746 VSS.t576 VSS.t1385 138.82
R5747 VSS.t565 VSS.t1389 138.82
R5748 VSS.t596 VSS.t1390 138.82
R5749 VSS.t605 VSS.t1183 138.82
R5750 VSS.t1187 VSS.t603 138.82
R5751 VSS.t1174 VSS.t553 138.82
R5752 VSS.t1175 VSS.t632 138.82
R5753 VSS.t379 VSS.t1044 138.82
R5754 VSS.t1048 VSS.t387 138.82
R5755 VSS.t1051 VSS.t383 138.82
R5756 VSS.t1039 VSS.t395 138.82
R5757 VSS.t645 VSS.t725 138.703
R5758 VSS.t591 VSS.t718 138.703
R5759 VSS.t660 VSS.t716 138.703
R5760 VSS.t634 VSS.t721 138.703
R5761 VSS.t1157 VSS.t1475 138.703
R5762 VSS.t1481 VSS.t1158 138.703
R5763 VSS.t1147 VSS.t1492 138.703
R5764 VSS.t1474 VSS.t1150 138.703
R5765 VSS.t1505 VSS.t652 138.703
R5766 VSS.t592 VSS.t1498 138.703
R5767 VSS.t666 VSS.t1501 138.703
R5768 VSS.t648 VSS.t1506 138.703
R5769 VSS.t1387 VSS.t649 138.703
R5770 VSS.t601 VSS.t1391 138.703
R5771 VSS.t1396 VSS.t579 138.703
R5772 VSS.t1399 VSS.t646 138.703
R5773 VSS.t1186 VSS.t588 138.703
R5774 VSS.t546 VSS.t1173 138.703
R5775 VSS.t618 VSS.t1176 138.703
R5776 VSS.t577 VSS.t1180 138.703
R5777 VSS.t1043 VSS.t388 138.703
R5778 VSS.t377 VSS.t1047 138.703
R5779 VSS.t386 VSS.t1052 138.703
R5780 VSS.t1040 VSS.t391 138.703
R5781 VSS.n5383 VSS.t1336 137.011
R5782 VSS.n5127 VSS.t1334 137.011
R5783 VSS.t1380 VSS.t1285 136.983
R5784 VSS.t1283 VSS.t1378 136.983
R5785 VSS.t1368 VSS.t73 136.983
R5786 VSS.t1371 VSS.t76 136.983
R5787 VSS.t526 VSS.t1360 136.983
R5788 VSS.t1366 VSS.t524 136.983
R5789 VSS.t896 VSS.t30 136.983
R5790 VSS.t887 VSS.t28 136.983
R5791 VSS.t314 VSS.t1216 136.983
R5792 VSS.t1220 VSS.t312 136.983
R5793 VSS.t10 VSS.t1243 136.983
R5794 VSS.t1246 VSS.t8 136.983
R5795 VSS.n2497 VSS.n2496 136.084
R5796 VSS.n4544 VSS.t1060 135.957
R5797 VSS.n4424 VSS.t758 135.957
R5798 VSS.n4448 VSS.t756 135.957
R5799 VSS.n4292 VSS.t922 135.957
R5800 VSS.t924 VSS.n2914 135.957
R5801 VSS.n4211 VSS.t909 135.957
R5802 VSS.n547 VSS.t1063 135.957
R5803 VSS.n5058 VSS.t135 135.581
R5804 VSS.n5427 VSS.t129 135.581
R5805 VSS.n90 VSS.t230 135.537
R5806 VSS.t405 VSS.n2502 135.537
R5807 VSS.t697 VSS.n4373 135.124
R5808 VSS.n4799 VSS.n4798 134.333
R5809 VSS.t1307 VSS.t695 133.35
R5810 VSS.t791 VSS.t1016 133.35
R5811 VSS.t475 VSS.t1112 133.35
R5812 VSS.t224 VSS.t489 133.35
R5813 VSS.t322 VSS.t999 133.35
R5814 VSS.t1166 VSS.t1134 133.35
R5815 VSS.t1514 VSS.t821 133.35
R5816 VSS.t1170 VSS.t174 133.35
R5817 VSS.t1330 VSS.t894 133.35
R5818 VSS.t0 VSS.t248 133.35
R5819 VSS.t218 VSS.t60 133.35
R5820 VSS.t505 VSS.t1459 133.35
R5821 VSS.t1431 VSS.t973 133.35
R5822 VSS.t1433 VSS.t1544 133.35
R5823 VSS.t851 VSS.t284 130.901
R5824 VSS.n24 VSS.t679 130.544
R5825 VSS.n2845 VSS.t82 130.544
R5826 VSS.n2568 VSS.t541 130.544
R5827 VSS.n2453 VSS.t1036 130.544
R5828 VSS.n1119 VSS.t421 130.544
R5829 VSS.n4036 VSS.t436 130.544
R5830 VSS.n5436 VSS.t1120 129.061
R5831 VSS.t1102 VSS.n5017 129.061
R5832 VSS.t427 VSS.n4982 127.457
R5833 VSS.n4479 VSS.t876 127.398
R5834 VSS.t276 VSS.n4489 127.398
R5835 VSS.t1478 VSS.n2930 125.344
R5836 VSS.n4355 VSS.t851 125.272
R5837 VSS.t131 VSS.t1193 125.15
R5838 VSS.t126 VSS.t1209 125.15
R5839 VSS.t654 VSS.n2462 123.9
R5840 VSS.t627 VSS.n33 123.719
R5841 VSS.n5079 VSS.t1275 122.543
R5842 VSS.n242 VSS.t800 122.543
R5843 VSS.n265 VSS.t1129 122.543
R5844 VSS.n128 VSS.t1123 122.543
R5845 VSS.n139 VSS.t1269 122.543
R5846 VSS.n5388 VSS.t1440 122.543
R5847 VSS.n4359 VSS.t1022 116.843
R5848 VSS.n2930 VSS.t1487 116.391
R5849 VSS.n251 VSS.t1407 112.115
R5850 VSS.t1319 VSS.n5113 112.115
R5851 VSS.n274 VSS.t1461 112.115
R5852 VSS.n170 VSS.t1454 112.115
R5853 VSS.n160 VSS.t1418 112.115
R5854 VSS.n5387 VSS.t1312 112.115
R5855 VSS.t868 VSS.t1534 108.832
R5856 VSS.t346 VSS.t560 108.413
R5857 VSS.t1032 VSS.t638 108.254
R5858 VSS.t1487 VSS.n2929 102.962
R5859 VSS.n4376 VSS.t789 97.6866
R5860 VSS.t769 VSS.n4478 97.6866
R5861 VSS.n4490 VSS.t1073 97.6866
R5862 VSS.n4983 VSS.t943 97.6866
R5863 VSS.n4339 VSS.t925 97.6866
R5864 VSS.n1743 VSS.t921 97.6866
R5865 VSS.n348 VSS.t1075 97.6866
R5866 VSS.n1334 VSS.n1333 97.0154
R5867 VSS.n2405 VSS.n2404 94.1232
R5868 VSS.n346 VSS.n333 92.4513
R5869 VSS.t1536 VSS.t688 89.3971
R5870 VSS.t689 VSS.t1539 89.3971
R5871 VSS.n1158 VSS.n1157 81.2223
R5872 VSS.n5437 VSS.t675 80.7458
R5873 VSS.t1011 VSS.n5015 80.7458
R5874 VSS.n4382 VSS.t1021 80.4405
R5875 VSS.n4468 VSS.t364 80.4405
R5876 VSS.t186 VSS.n4519 80.4405
R5877 VSS.t700 VSS.n4995 80.4405
R5878 VSS.n1731 VSS.t1354 80.4405
R5879 VSS.n4313 VSS.t62 80.4405
R5880 VSS.n769 VSS.t367 75.9786
R5881 VSS.n4987 VSS.t240 75.9786
R5882 VSS.n1716 VSS.t1493 75.9786
R5883 VSS.n2470 VSS.t1031 75.0555
R5884 VSS.n43 VSS.t867 74.9456
R5885 VSS.n4388 VSS.t264 74.428
R5886 VSS.n4495 VSS.t208 74.428
R5887 VSS.n4320 VSS.t67 74.428
R5888 VSS.n344 VSS.t465 74.428
R5889 VSS.n4155 VSS.n4154 70.8693
R5890 VSS.t260 VSS.t983 69.2108
R5891 VSS.t675 VSS.t987 69.2108
R5892 VSS.t404 VSS.t989 69.2108
R5893 VSS.t992 VSS.t1011 69.2108
R5894 VSS.n18 VSS.t1300 67.9921
R5895 VSS.n2839 VSS.t257 67.9921
R5896 VSS.n2569 VSS.t43 67.9921
R5897 VSS.n2447 VSS.t1555 67.9921
R5898 VSS.n1120 VSS.t482 67.9921
R5899 VSS.n4034 VSS.t863 67.9921
R5900 VSS.t764 VSS.t1020 64.7994
R5901 VSS.t1018 VSS.t782 64.7994
R5902 VSS.t115 VSS.t786 64.7994
R5903 VSS.t761 VSS.t463 64.7994
R5904 VSS.t770 VSS.t476 64.7994
R5905 VSS.t363 VSS.t778 64.7994
R5906 VSS.t185 VSS.t1064 64.7994
R5907 VSS.t1076 VSS.t1163 64.7994
R5908 VSS.t1095 VSS.t882 64.7994
R5909 VSS.t1028 VSS.t930 64.7994
R5910 VSS.t1515 VSS.t944 64.7994
R5911 VSS.t701 VSS.t967 64.7994
R5912 VSS.t1352 VSS.t954 64.7994
R5913 VSS.t889 VSS.t964 64.7994
R5914 VSS.t959 VSS.t1355 64.7994
R5915 VSS.t933 VSS.t63 64.7994
R5916 VSS.t904 VSS.t507 64.7994
R5917 VSS.t911 VSS.t532 64.7994
R5918 VSS.n4968 VSS.n4967 62.5655
R5919 VSS.n1070 VSS.t790 62.0234
R5920 VSS.n4507 VSS.t1059 62.0234
R5921 VSS.n4316 VSS.t923 62.0234
R5922 VSS.n359 VSS.t1061 62.0234
R5923 VSS.n2504 VSS.t689 60.5595
R5924 VSS.n763 VSS.t757 60.4728
R5925 VSS.n304 VSS.t926 60.4728
R5926 VSS.n1708 VSS.t966 60.4728
R5927 VSS.n19 VSS.n18 59.8331
R5928 VSS.n2840 VSS.n2839 59.8331
R5929 VSS.n2570 VSS.n2569 59.8331
R5930 VSS.n2448 VSS.n2447 59.8331
R5931 VSS.n1121 VSS.n1120 59.8331
R5932 VSS.n4035 VSS.n4034 59.8331
R5933 VSS.t452 VSS.n2495 57.1852
R5934 VSS.n42 VSS.t492 57.1015
R5935 VSS.t445 VSS.n4338 53.2797
R5936 VSS.n5269 VSS.n5268 51.9102
R5937 VSS.n2498 VSS.t1536 46.1407
R5938 VSS.n2959 VSS.n2821 45.3916
R5939 VSS.t619 VSS.n4440 43.1612
R5940 VSS.t568 VSS.n4273 43.1612
R5941 VSS.n2882 VSS.t606 43.1612
R5942 VSS.t122 VSS.t1022 43.1421
R5943 VSS.t146 VSS.t981 43.1421
R5944 VSS.n4113 VSS.t111 41.8685
R5945 VSS.t598 VSS.n4554 41.0032
R5946 VSS.n4423 VSS.t550 41.0032
R5947 VSS.n4233 VSS.t615 41.0032
R5948 VSS.n548 VSS.t584 41.0032
R5949 VSS.n4373 VSS.t1261 38.004
R5950 VSS.t711 VSS.t1189 36.8625
R5951 VSS.t818 VSS.t1321 36.8625
R5952 VSS.n5115 VSS.n5114 36.8625
R5953 VSS.t311 VSS.t424 36.8625
R5954 VSS.t1333 VSS.t845 36.8625
R5955 VSS.t402 VSS.t196 36.8625
R5956 VSS.t1466 VSS.t1126 36.8625
R5957 VSS.n5100 VSS.n5099 36.8625
R5958 VSS.t158 VSS.t144 36.8625
R5959 VSS.t1409 VSS.t1274 36.8625
R5960 VSS.t198 VSS.t398 36.8625
R5961 VSS.t1456 VSS.t1139 36.8625
R5962 VSS.n175 VSS.n131 36.8625
R5963 VSS.t51 VSS.t1009 36.8625
R5964 VSS.t1406 VSS.t1265 36.8625
R5965 VSS.t203 VSS.t182 36.8625
R5966 VSS.t1316 VSS.t1445 36.8625
R5967 VSS.n5386 VSS.n5385 36.8625
R5968 VSS.t302 VSS.t444 36.8625
R5969 VSS.t1344 VSS.t854 36.8625
R5970 VSS.n4102 VSS.n4101 35.8284
R5971 VSS.n4376 VSS.t1017 35.6637
R5972 VSS.n4478 VSS.t474 35.6637
R5973 VSS.t1165 VSS.n4490 35.6637
R5974 VSS.t1520 VSS.n4983 35.6637
R5975 VSS.n4339 VSS.t895 35.6637
R5976 VSS.t506 VSS.n1743 35.6637
R5977 VSS.t1439 VSS.n348 35.6637
R5978 VSS.n4054 VSS.n4053 35.447
R5979 VSS.n5060 VSS.t1010 34.8146
R5980 VSS.t521 VSS.n5429 34.8146
R5981 VSS.n4758 VSS.n4757 34.6159
R5982 VSS.n3722 VSS.n3721 31.0162
R5983 VSS.n5384 VSS.n5383 28.677
R5984 VSS.n5127 VSS.n5125 28.677
R5985 VSS.n4064 VSS.n4063 28.2494
R5986 VSS.n1618 VSS.n1617 27.6079
R5987 VSS.n1136 VSS.n1086 27.4335
R5988 VSS.n4361 VSS.t1423 26.5311
R5989 VSS.n4335 VSS.n4334 26.1752
R5990 VSS.t213 VSS.n346 26.167
R5991 VSS.n4759 VSS.n4758 25.3911
R5992 VSS.n2462 VSS.t346 25.0188
R5993 VSS.n33 VSS.t1032 24.9822
R5994 VSS.t145 VSS.n4351 24.9752
R5995 VSS.n1614 VSS.n1613 24.5404
R5996 VSS.t1275 VSS.t1420 23.4662
R5997 VSS.t1407 VSS.t1259 23.4662
R5998 VSS.t800 VSS.t1309 23.4662
R5999 VSS.n5113 VSS.n242 23.4662
R6000 VSS.t816 VSS.t1319 23.4662
R6001 VSS.t1129 VSS.t1451 23.4662
R6002 VSS.t1461 VSS.t1137 23.4662
R6003 VSS.t1123 VSS.t1469 23.4662
R6004 VSS.t1454 VSS.t1132 23.4662
R6005 VSS.t1269 VSS.t1415 23.4662
R6006 VSS.t1418 VSS.t1272 23.4662
R6007 VSS.t1440 VSS.t1324 23.4662
R6008 VSS.n5388 VSS.n5387 23.4662
R6009 VSS.t1312 VSS.t1443 23.4662
R6010 VSS.n95 VSS.t1108 23.0706
R6011 VSS.n5036 VSS.t1118 23.0706
R6012 VSS.n41 VSS.t868 22.5772
R6013 VSS.n2496 VSS.t1030 22.5687
R6014 VSS.n4967 VSS.t457 22.2219
R6015 VSS.t1193 VSS.n5058 20.8589
R6016 VSS.t1209 VSS.n5427 20.8589
R6017 VSS.t472 VSS.n4467 20.1579
R6018 VSS.t1518 VSS.n4994 20.1579
R6019 VSS.n1706 VSS.t892 20.1579
R6020 VSS.n3739 VSS.n3738 20.1468
R6021 VSS.n3479 VSS.t352 19.3409
R6022 VSS.n4139 VSS.n4138 19.19
R6023 VSS.n4383 VSS.t1013 18.6074
R6024 VSS.n4505 VSS.t1529 18.6074
R6025 VSS.n4314 VSS.t502 18.6074
R6026 VSS.n357 VSS.t1434 18.6074
R6027 VSS.n3439 VSS.t220 18.1322
R6028 VSS.n4126 VSS.t885 17.4455
R6029 VSS.n4004 VSS.n4003 17.3263
R6030 VSS.n4885 VSS.n4884 16.9276
R6031 VSS.n2938 VSS.n2937 14.5494
R6032 VSS.n5037 VSS.t826 14.3357
R6033 VSS.n5430 VSS.t841 14.3357
R6034 VSS.n1513 VSS.n1508 14.3087
R6035 VSS.n2781 VSS.n2780 13.339
R6036 VSS.n983 VSS.n982 13.0165
R6037 VSS.n2465 VSS.t118 12.3882
R6038 VSS.n36 VSS.t71 12.3613
R6039 VSS.n5435 VSS.t831 11.5355
R6040 VSS.n5018 VSS.t836 11.5355
R6041 VSS.n11 VSS.n9 10.8883
R6042 VSS.n5476 VSS.n5475 10.8883
R6043 VSS.n2830 VSS.n2829 10.8883
R6044 VSS.n2835 VSS.n2834 10.8883
R6045 VSS.n2557 VSS.n2556 10.8883
R6046 VSS.n2562 VSS.n2560 10.8883
R6047 VSS.n2438 VSS.n2437 10.8883
R6048 VSS.n2443 VSS.n2442 10.8883
R6049 VSS.n1108 VSS.n1107 10.8883
R6050 VSS.n1113 VSS.n1111 10.8883
R6051 VSS.n4023 VSS.n4022 10.8883
R6052 VSS.n4028 VSS.n4026 10.8883
R6053 VSS.n27 VSS.n20 10.8792
R6054 VSS.n30 VSS.n29 10.8792
R6055 VSS.n2848 VSS.n2841 10.8792
R6056 VSS.n2851 VSS.n2850 10.8792
R6057 VSS.n2577 VSS.n2576 10.8792
R6058 VSS.n2580 VSS.n2579 10.8792
R6059 VSS.n2456 VSS.n2449 10.8792
R6060 VSS.n2459 VSS.n2458 10.8792
R6061 VSS.n1128 VSS.n1127 10.8792
R6062 VSS.n1131 VSS.n1130 10.8792
R6063 VSS.n4041 VSS.n4040 10.8792
R6064 VSS.n4052 VSS.n2428 10.8792
R6065 VSS.n1159 VSS.n1155 10.5005
R6066 VSS.n1512 VSS.n1510 10.5005
R6067 VSS.n889 VSS.n887 10.5005
R6068 VSS.n5059 VSS.t131 10.4297
R6069 VSS.n5428 VSS.t126 10.4297
R6070 VSS.n2822 VSS.n2609 9.95404
R6071 VSS.n554 VSS.n553 9.88396
R6072 VSS.n4082 VSS.t381 9.64646
R6073 VSS.n3745 VSS.t805 8.86487
R6074 VSS.n2590 VSS.n2589 8.84039
R6075 VSS VSS.n1078 8.3883
R6076 VSS.n4003 VSS.t799 8.05902
R6077 VSS.t1055 VSS.n4968 7.99558
R6078 VSS.n4366 VSS.n4365 7.78196
R6079 VSS.n3373 VSS.n3372 7.65609
R6080 VSS.n1746 VSS.n1069 6.91683
R6081 VSS.n4456 VSS.n298 6.88665
R6082 VSS.n5001 VSS.n5000 6.88175
R6083 VSS.n4186 VSS.n4185 6.85891
R6084 VSS.n3458 VSS.t33 6.85024
R6085 VSS.n991 VSS.n988 6.79475
R6086 VSS.n546 VSS.n224 6.75725
R6087 VSS.n4560 VSS.n4559 6.7505
R6088 VSS.n4562 VSS.n4561 6.7505
R6089 VSS.n4181 VSS.n4180 6.7505
R6090 VSS.n4392 VSS.n1058 6.7505
R6091 VSS.n990 VSS.n779 6.73295
R6092 VSS.n303 VSS.n302 6.73295
R6093 VSS.n4522 VSS.n4521 6.73247
R6094 VSS.n368 VSS.n367 6.73247
R6095 VSS.n4200 VSS.n4199 6.73137
R6096 VSS.n4394 VSS.n1039 6.73137
R6097 VSS.n4357 VSS.n4356 6.60306
R6098 VSS.n4538 VSS.n4537 6.23171
R6099 VSS.n4475 VSS.n4474 6.23171
R6100 VSS.n4445 VSS.n4444 6.23171
R6101 VSS.n4370 VSS.n1072 6.23171
R6102 VSS.n4406 VSS.n4405 6.23171
R6103 VSS.n330 VSS.n329 6.23171
R6104 VSS.n4278 VSS.n4277 6.23171
R6105 VSS.n2891 VSS.n2868 6.23171
R6106 VSS.n4328 VSS.n4327 6.23171
R6107 VSS.n4306 VSS.n4305 6.23171
R6108 VSS.n4961 VSS.n375 6.23171
R6109 VSS.n4224 VSS.n4204 6.23168
R6110 VSS.n4486 VSS.n754 6.23168
R6111 VSS.n4452 VSS.n4451 6.23168
R6112 VSS.n4409 VSS.n1033 6.23168
R6113 VSS.n4289 VSS.n4288 6.23168
R6114 VSS.n1735 VSS.n1734 6.23168
R6115 VSS.n4532 VSS.n4525 6.23168
R6116 VSS.n2922 VSS.n2921 6.23168
R6117 VSS.n532 VSS.n371 6.23168
R6118 VSS.n4976 VSS.n336 6.23168
R6119 VSS.t796 VSS.n4375 6.20279
R6120 VSS.n4497 VSS.t1142 6.20279
R6121 VSS.n4187 VSS.t1463 6.20279
R6122 VSS.n349 VSS.t1550 6.20279
R6123 VSS.n4304 VSS.n4303 6.02724
R6124 VSS.n4231 VSS.n4230 6.02724
R6125 VSS.n4326 VSS.n4325 6.02724
R6126 VSS.n1733 VSS.n1715 6.02724
R6127 VSS.n4530 VSS.n4529 6.02724
R6128 VSS.n2923 VSS.n2861 6.02724
R6129 VSS.n537 VSS.n536 6.02724
R6130 VSS.n749 VSS.n746 6.02724
R6131 VSS.n4515 VSS.n4514 6.02724
R6132 VSS.n4477 VSS.n4476 6.02724
R6133 VSS.n4450 VSS.n4449 6.02724
R6134 VSS.n4404 VSS.n1026 6.02724
R6135 VSS.n4447 VSS.n4446 6.02724
R6136 VSS.n4412 VSS.n4411 6.02724
R6137 VSS.n4378 VSS.n4377 6.02724
R6138 VSS.n328 VSS.n327 6.02724
R6139 VSS.n4291 VSS.n4254 6.02724
R6140 VSS.n4276 VSS.n4250 6.02724
R6141 VSS.n4974 VSS.n4973 6.02724
R6142 VSS.n2893 VSS.n2892 6.02724
R6143 VSS.n4959 VSS.n4958 6.02724
R6144 VSS.n4345 VSS.n4344 5.79501
R6145 VSS VSS.t121 5.6459
R6146 VSS VSS.t804 5.43302
R6147 VSS.n4430 VSS.n4429 5.41668
R6148 VSS VSS.t1367 5.39046
R6149 VSS VSS.t1247 5.39046
R6150 VSS VSS.t1221 5.39046
R6151 VSS.n2853 VSS.t1488 5.38269
R6152 VSS.n1302 VSS.t1192 5.38269
R6153 VSS VSS.t1262 5.36235
R6154 VSS.n366 VSS.t108 5.3339
R6155 VSS.n2917 VSS.n2871 5.3339
R6156 VSS.n750 VSS.t50 5.3339
R6157 VSS.n4396 VSS.t326 5.3339
R6158 VSS.n2856 VSS.t515 5.3339
R6159 VSS.n4330 VSS.t54 5.3339
R6160 VSS.n4310 VSS.t1356 5.3339
R6161 VSS.n4298 VSS.n4297 5.32067
R6162 VSS VSS.n1079 5.31891
R6163 VSS.n4031 VSS.n4030 5.30927
R6164 VSS.n1116 VSS.n1115 5.30927
R6165 VSS.n2565 VSS.n2564 5.30927
R6166 VSS.n2949 VSS.n2948 5.30927
R6167 VSS.n2524 VSS.n2523 5.30927
R6168 VSS.n4348 VSS.n4347 5.24868
R6169 VSS.n540 VSS.t1094 5.247
R6170 VSS.n5457 VSS.t1033 5.24132
R6171 VSS.n4132 VSS.t1363 5.23399
R6172 VSS.n2607 VSS.t498 5.23126
R6173 VSS.n4224 VSS.t308 5.23126
R6174 VSS.n4223 VSS.t173 5.23126
R6175 VSS.n1734 VSS.n1728 5.23126
R6176 VSS.n4525 VSS.t1004 5.23126
R6177 VSS.n2469 VSS.t347 5.23126
R6178 VSS.n34 VSS.t1008 5.23126
R6179 VSS.n2922 VSS.n2862 5.23126
R6180 VSS.n2864 VSS.n2863 5.23126
R6181 VSS.n532 VSS.t79 5.23126
R6182 VSS.n531 VSS.t1012 5.23126
R6183 VSS.n4537 VSS.t349 5.23126
R6184 VSS.n4531 VSS.t88 5.23126
R6185 VSS.n4536 VSS.t169 5.23126
R6186 VSS.n754 VSS.t110 5.23126
R6187 VSS.n4475 VSS.n4470 5.23126
R6188 VSS.n4451 VSS.n997 5.23126
R6189 VSS.n996 VSS.n995 5.23126
R6190 VSS.n4445 VSS.n4443 5.23126
R6191 VSS.n1007 VSS.n1006 5.23126
R6192 VSS.n1033 VSS.t1279 5.23126
R6193 VSS.n4410 VSS.t699 5.23126
R6194 VSS.n1073 VSS.t696 5.23126
R6195 VSS.n1072 VSS.t101 5.23126
R6196 VSS.n4400 VSS.t195 5.23126
R6197 VSS.n4405 VSS.t269 5.23126
R6198 VSS.n755 VSS.t1000 5.23126
R6199 VSS.n760 VSS.n759 5.23126
R6200 VSS.n329 VSS.n323 5.23126
R6201 VSS.n4288 VSS.n4287 5.23126
R6202 VSS.n4290 VSS.n4255 5.23126
R6203 VSS.n4277 VSS.n4258 5.23126
R6204 VSS.n4257 VSS.n4256 5.23126
R6205 VSS.n336 VSS.t995 5.23126
R6206 VSS.n4975 VSS.t974 5.23126
R6207 VSS.n322 VSS.n321 5.23126
R6208 VSS.n1727 VSS.n1726 5.23126
R6209 VSS.n2886 VSS.n2885 5.23126
R6210 VSS.n2891 VSS.n2890 5.23126
R6211 VSS.n1740 VSS.t219 5.23126
R6212 VSS.n4327 VSS.t339 5.23126
R6213 VSS.n4208 VSS.t729 5.23126
R6214 VSS.n4305 VSS.t93 5.23126
R6215 VSS.n4960 VSS.t157 5.23126
R6216 VSS.n375 VSS.t360 5.23126
R6217 VSS.n2610 VSS.t353 5.23126
R6218 VSS.n1015 VSS.n1014 5.21498
R6219 VSS.n4268 VSS.n4267 5.21498
R6220 VSS.n2875 VSS.n2874 5.21498
R6221 VSS.n4237 VSS.t920 5.21406
R6222 VSS.n4550 VSS.t1058 5.21406
R6223 VSS.n4418 VSS.t777 5.21406
R6224 VSS.n5085 VSS.t1320 5.20602
R6225 VSS.n263 VSS.t1462 5.20602
R6226 VSS.n275 VSS.t1138 5.20602
R6227 VSS.n5111 VSS.t817 5.20602
R6228 VSS.n5019 VSS.t1119 5.20602
R6229 VSS.n5034 VSS.t830 5.20602
R6230 VSS.n5451 VSS.t1535 5.20602
R6231 VSS.n5389 VSS.t1313 5.20602
R6232 VSS.n5405 VSS.t1455 5.20602
R6233 VSS.n151 VSS.t1444 5.20602
R6234 VSS.n172 VSS.t1133 5.20602
R6235 VSS.n69 VSS.t840 5.20602
R6236 VSS.n5433 VSS.t1109 5.20602
R6237 VSS.n2483 VSS.t1540 5.20602
R6238 VSS.n2458 VSS 5.20494
R6239 VSS VSS.n5476 5.20494
R6240 VSS.n29 VSS 5.20494
R6241 VSS.n2579 VSS 5.20494
R6242 VSS.n2560 VSS 5.20494
R6243 VSS.n4026 VSS 5.20494
R6244 VSS.n2850 VSS 5.20494
R6245 VSS.n2834 VSS 5.20494
R6246 VSS.n2442 VSS 5.20494
R6247 VSS.n1111 VSS 5.20494
R6248 VSS.n1130 VSS 5.20494
R6249 VSS VSS.n2428 5.20494
R6250 VSS.n3736 VSS 5.2005
R6251 VSS VSS.n4526 5.2005
R6252 VSS.n5114 VSS 5.2005
R6253 VSS VSS.n5115 5.2005
R6254 VSS.n5113 VSS.n5112 5.2005
R6255 VSS.n5080 VSS.n5079 5.2005
R6256 VSS.n5086 VSS.n242 5.2005
R6257 VSS.n252 VSS.n251 5.2005
R6258 VSS.n5099 VSS 5.2005
R6259 VSS VSS.n5100 5.2005
R6260 VSS VSS.n5037 5.2005
R6261 VSS.n5059 VSS.n5046 5.2005
R6262 VSS.n276 VSS.n274 5.2005
R6263 VSS.n266 VSS.n265 5.2005
R6264 VSS.n5058 VSS.n5057 5.2005
R6265 VSS VSS.n5060 5.2005
R6266 VSS VSS.n2466 5.2005
R6267 VSS VSS.n11 5.2005
R6268 VSS.n5479 VSS.n9 5.2005
R6269 VSS.n5475 VSS.n5474 5.2005
R6270 VSS VSS.n27 5.2005
R6271 VSS VSS.n24 5.2005
R6272 VSS.n5469 VSS.n19 5.2005
R6273 VSS.n5465 VSS.n30 5.2005
R6274 VSS.n5467 VSS.n20 5.2005
R6275 VSS VSS.n37 5.2005
R6276 VSS VSS.n5430 5.2005
R6277 VSS.n5429 VSS 5.2005
R6278 VSS.n5428 VSS.n118 5.2005
R6279 VSS.n171 VSS.n170 5.2005
R6280 VSS.n5406 VSS.n128 5.2005
R6281 VSS.n5427 VSS.n5426 5.2005
R6282 VSS VSS.n131 5.2005
R6283 VSS VSS.n175 5.2005
R6284 VSS.n5387 VSS.n145 5.2005
R6285 VSS.n140 VSS.n139 5.2005
R6286 VSS.n5390 VSS.n5388 5.2005
R6287 VSS.n161 VSS.n160 5.2005
R6288 VSS.n5385 VSS 5.2005
R6289 VSS.n5386 VSS 5.2005
R6290 VSS.n5383 VSS.n215 5.2005
R6291 VSS.n5384 VSS.n200 5.2005
R6292 VSS.n4153 VSS.n4152 5.2005
R6293 VSS.n2958 VSS 5.2005
R6294 VSS.n2957 VSS.n2956 5.2005
R6295 VSS VSS.n2830 5.2005
R6296 VSS.n2953 VSS.n2829 5.2005
R6297 VSS.n2950 VSS.n2835 5.2005
R6298 VSS.n2944 VSS.n2841 5.2005
R6299 VSS VSS.n2848 5.2005
R6300 VSS VSS.n2845 5.2005
R6301 VSS.n2946 VSS.n2840 5.2005
R6302 VSS.n2942 VSS.n2851 5.2005
R6303 VSS.n2930 VSS.n2853 5.2005
R6304 VSS.n2940 VSS.n2939 5.2005
R6305 VSS.n2939 VSS.n2938 5.2005
R6306 VSS.n2550 VSS 5.2005
R6307 VSS.n2552 VSS.n2551 5.2005
R6308 VSS VSS.n2557 5.2005
R6309 VSS.n2556 VSS.n2555 5.2005
R6310 VSS.n2563 VSS.n2562 5.2005
R6311 VSS.n2571 VSS.n2570 5.2005
R6312 VSS.n2581 VSS.n2580 5.2005
R6313 VSS.n2576 VSS.n2575 5.2005
R6314 VSS VSS.n2577 5.2005
R6315 VSS.n2568 VSS 5.2005
R6316 VSS.n2587 VSS.n2586 5.2005
R6317 VSS.n2585 VSS 5.2005
R6318 VSS.n5494 VSS 5.2005
R6319 VSS.n5493 VSS.n5492 5.2005
R6320 VSS.n5462 VSS.n33 5.2005
R6321 VSS VSS.n31 5.2005
R6322 VSS VSS.n43 5.2005
R6323 VSS.n5452 VSS.n48 5.2005
R6324 VSS.n88 VSS.n87 5.2005
R6325 VSS VSS.n51 5.2005
R6326 VSS.n5438 VSS.n5437 5.2005
R6327 VSS.n5435 VSS.n5434 5.2005
R6328 VSS.n91 VSS.n90 5.2005
R6329 VSS.n96 VSS.n95 5.2005
R6330 VSS.n5125 VSS.n5124 5.2005
R6331 VSS.n5128 VSS.n5127 5.2005
R6332 VSS VSS.n4556 5.2005
R6333 VSS.n4566 VSS 5.2005
R6334 VSS.n4566 VSS 5.2005
R6335 VSS.n4554 VSS.n4553 5.2005
R6336 VSS VSS.n4544 5.2005
R6337 VSS.n4544 VSS 5.2005
R6338 VSS.n4543 VSS.n750 5.2005
R6339 VSS.n4543 VSS.n4542 5.2005
R6340 VSS VSS.n4469 5.2005
R6341 VSS.n1010 VSS 5.2005
R6342 VSS VSS.n4442 5.2005
R6343 VSS.n4381 VSS 5.2005
R6344 VSS VSS.n4376 5.2005
R6345 VSS.n4385 VSS.n4384 5.2005
R6346 VSS.n4384 VSS.n4383 5.2005
R6347 VSS.n1071 VSS.n1070 5.2005
R6348 VSS.n4374 VSS.n1064 5.2005
R6349 VSS.n4375 VSS.n4374 5.2005
R6350 VSS.n4395 VSS 5.2005
R6351 VSS.n4398 VSS.n4397 5.2005
R6352 VSS.n4397 VSS.n4396 5.2005
R6353 VSS VSS.n4403 5.2005
R6354 VSS.n4415 VSS 5.2005
R6355 VSS.n4424 VSS 5.2005
R6356 VSS.n4423 VSS.n4422 5.2005
R6357 VSS VSS.n4424 5.2005
R6358 VSS.n4435 VSS 5.2005
R6359 VSS VSS.n4417 5.2005
R6360 VSS.n4417 VSS 5.2005
R6361 VSS VSS.n4435 5.2005
R6362 VSS.n4448 VSS 5.2005
R6363 VSS.n4440 VSS.n4439 5.2005
R6364 VSS VSS.n4448 5.2005
R6365 VSS.n775 VSS.n774 5.2005
R6366 VSS.n774 VSS.n773 5.2005
R6367 VSS.n4464 VSS.n764 5.2005
R6368 VSS.n764 VSS.n763 5.2005
R6369 VSS.n4466 VSS.n4465 5.2005
R6370 VSS.n4467 VSS.n4466 5.2005
R6371 VSS.n4506 VSS.n4504 5.2005
R6372 VSS.n4506 VSS.n4505 5.2005
R6373 VSS.n4509 VSS.n4508 5.2005
R6374 VSS.n4508 VSS.n4507 5.2005
R6375 VSS.n4499 VSS.n4498 5.2005
R6376 VSS.n4498 VSS.n4497 5.2005
R6377 VSS.n4518 VSS 5.2005
R6378 VSS VSS.n4520 5.2005
R6379 VSS VSS.n4490 5.2005
R6380 VSS.n4489 VSS.n4488 5.2005
R6381 VSS.n4480 VSS.n4479 5.2005
R6382 VSS.n4478 VSS 5.2005
R6383 VSS VSS.n4459 5.2005
R6384 VSS.n4458 VSS.n4457 5.2005
R6385 VSS VSS.n326 5.2005
R6386 VSS.n4263 VSS 5.2005
R6387 VSS VSS.n4275 5.2005
R6388 VSS VSS.n4292 5.2005
R6389 VSS.n4273 VSS.n4272 5.2005
R6390 VSS.n4292 VSS 5.2005
R6391 VSS.n4986 VSS.n4985 5.2005
R6392 VSS.n4985 VSS.n4984 5.2005
R6393 VSS.n4991 VSS.n305 5.2005
R6394 VSS.n305 VSS.n304 5.2005
R6395 VSS.n4993 VSS.n4992 5.2005
R6396 VSS.n4994 VSS.n4993 5.2005
R6397 VSS VSS.n4970 5.2005
R6398 VSS.n4983 VSS 5.2005
R6399 VSS.n4996 VSS 5.2005
R6400 VSS.n4997 VSS.n299 5.2005
R6401 VSS.n4998 VSS.n4997 5.2005
R6402 VSS.n2505 VSS.n2504 5.2005
R6403 VSS.n2499 VSS.n2498 5.2005
R6404 VSS.n2503 VSS 5.2005
R6405 VSS.n5015 VSS.n5014 5.2005
R6406 VSS.n5020 VSS.n5018 5.2005
R6407 VSS.n2502 VSS.n2501 5.2005
R6408 VSS.n5036 VSS.n5035 5.2005
R6409 VSS.n2514 VSS.n2462 5.2005
R6410 VSS VSS.n2460 5.2005
R6411 VSS VSS.n2470 5.2005
R6412 VSS.n2519 VSS.n2449 5.2005
R6413 VSS.n2521 VSS.n2448 5.2005
R6414 VSS.n2517 VSS.n2459 5.2005
R6415 VSS VSS.n2456 5.2005
R6416 VSS VSS.n2453 5.2005
R6417 VSS VSS.n2438 5.2005
R6418 VSS.n2528 VSS.n2437 5.2005
R6419 VSS.n2525 VSS.n2443 5.2005
R6420 VSS.n2532 VSS.n2531 5.2005
R6421 VSS VSS.n2533 5.2005
R6422 VSS VSS.n4339 5.2005
R6423 VSS.n1721 VSS.n1720 5.2005
R6424 VSS.n1722 VSS.n1721 5.2005
R6425 VSS.n1710 VSS.n1709 5.2005
R6426 VSS.n1709 VSS.n1708 5.2005
R6427 VSS.n1707 VSS.n1705 5.2005
R6428 VSS.n1707 VSS.n1706 5.2005
R6429 VSS.n4337 VSS.n1737 5.2005
R6430 VSS VSS.n1732 5.2005
R6431 VSS VSS.n1698 5.2005
R6432 VSS.n2917 VSS.n2916 5.2005
R6433 VSS.n2916 VSS.n2915 5.2005
R6434 VSS VSS.n2889 5.2005
R6435 VSS.n2924 VSS 5.2005
R6436 VSS.n2914 VSS 5.2005
R6437 VSS.n2883 VSS.n2882 5.2005
R6438 VSS.n2914 VSS 5.2005
R6439 VSS.n2926 VSS 5.2005
R6440 VSS.n2926 VSS 5.2005
R6441 VSS.n1101 VSS 5.2005
R6442 VSS.n1103 VSS.n1102 5.2005
R6443 VSS VSS.n1108 5.2005
R6444 VSS.n1107 VSS.n1106 5.2005
R6445 VSS.n1114 VSS.n1113 5.2005
R6446 VSS VSS.n1128 5.2005
R6447 VSS.n1119 VSS 5.2005
R6448 VSS.n1122 VSS.n1121 5.2005
R6449 VSS.n1132 VSS.n1131 5.2005
R6450 VSS.n1127 VSS.n1126 5.2005
R6451 VSS.n1303 VSS.n1302 5.2005
R6452 VSS.n1138 VSS.n1137 5.2005
R6453 VSS.n1136 VSS 5.2005
R6454 VSS.n2857 VSS.n2856 5.2005
R6455 VSS.n4331 VSS.n4330 5.2005
R6456 VSS.n4195 VSS 5.2005
R6457 VSS VSS.n1743 5.2005
R6458 VSS.n4315 VSS.n4194 5.2005
R6459 VSS.n4315 VSS.n4314 5.2005
R6460 VSS.n4318 VSS.n4317 5.2005
R6461 VSS.n4317 VSS.n4316 5.2005
R6462 VSS.n4189 VSS.n4188 5.2005
R6463 VSS.n4188 VSS.n4187 5.2005
R6464 VSS.n4312 VSS 5.2005
R6465 VSS.n4311 VSS.n4201 5.2005
R6466 VSS.n4311 VSS.n4310 5.2005
R6467 VSS.n4225 VSS 5.2005
R6468 VSS VSS.n4227 5.2005
R6469 VSS VSS.n4211 5.2005
R6470 VSS VSS.n4211 5.2005
R6471 VSS.n4234 VSS.n4233 5.2005
R6472 VSS VSS.n4238 5.2005
R6473 VSS VSS.n4245 5.2005
R6474 VSS VSS.n4245 5.2005
R6475 VSS.n4238 VSS 5.2005
R6476 VSS.n4982 VSS.n4981 5.2005
R6477 VSS.n4978 VSS.n333 5.2005
R6478 VSS.n358 VSS.n356 5.2005
R6479 VSS.n358 VSS.n357 5.2005
R6480 VSS.n361 VSS.n360 5.2005
R6481 VSS.n360 VSS.n359 5.2005
R6482 VSS.n351 VSS.n350 5.2005
R6483 VSS.n350 VSS.n349 5.2005
R6484 VSS.n348 VSS 5.2005
R6485 VSS.n4969 VSS 5.2005
R6486 VSS.n4966 VSS.n366 5.2005
R6487 VSS.n4966 VSS.n4965 5.2005
R6488 VSS VSS.n4957 5.2005
R6489 VSS VSS.n533 5.2005
R6490 VSS.n547 VSS 5.2005
R6491 VSS.n549 VSS.n548 5.2005
R6492 VSS.n547 VSS 5.2005
R6493 VSS.n4955 VSS 5.2005
R6494 VSS.n4955 VSS 5.2005
R6495 VSS VSS.n4355 5.2005
R6496 VSS.n4373 VSS.n4372 5.2005
R6497 VSS.n1299 VSS 5.2005
R6498 VSS VSS.n4361 5.2005
R6499 VSS.n4359 VSS 5.2005
R6500 VSS.n4353 VSS.n4352 5.2005
R6501 VSS VSS.n1314 5.2005
R6502 VSS.n1322 VSS 5.2005
R6503 VSS VSS.n1323 5.2005
R6504 VSS.n1330 VSS 5.2005
R6505 VSS.n4018 VSS.n4017 5.2005
R6506 VSS.n4016 VSS 5.2005
R6507 VSS.n4022 VSS.n4021 5.2005
R6508 VSS.n4029 VSS.n4028 5.2005
R6509 VSS VSS.n4023 5.2005
R6510 VSS.n4040 VSS 5.2005
R6511 VSS VSS.n4036 5.2005
R6512 VSS.n4105 VSS.n4104 5.2005
R6513 VSS VSS.n4102 5.2005
R6514 VSS.n4052 VSS.n4051 5.2005
R6515 VSS.n4042 VSS.n4041 5.2005
R6516 VSS.n4035 VSS.n4033 5.2005
R6517 VSS.n4108 VSS.n4107 5.2005
R6518 VSS.n5191 VSS.n5190 5.2005
R6519 VSS.n5183 VSS.n5182 5.2005
R6520 VSS.n1764 VSS.n1763 5.2005
R6521 VSS.n5214 VSS.n5213 5.2005
R6522 VSS.n5202 VSS.n5201 5.2005
R6523 VSS.n3454 VSS.n3453 5.2005
R6524 VSS VSS.n4004 5.2005
R6525 VSS VSS.n5500 5.2005
R6526 VSS.n4979 VSS.t536 5.18736
R6527 VSS.n1328 VSS.t1237 5.17491
R6528 VSS.n2822 VSS.t1372 5.17237
R6529 VSS.n2534 VSS.t1284 5.16935
R6530 VSS.n779 VSS.n778 5.16302
R6531 VSS.n303 VSS.n300 5.16302
R6532 VSS.n4343 VSS.n1697 5.16302
R6533 VSS.n4199 VSS.t912 5.1621
R6534 VSS.n4394 VSS.t787 5.1621
R6535 VSS.n4521 VSS.t1096 5.1621
R6536 VSS.n367 VSS.t1056 5.1621
R6537 VSS.n5000 VSS.n4999 5.1539
R6538 VSS.n2554 VSS.n2553 5.15366
R6539 VSS.n4020 VSS.n4019 5.15366
R6540 VSS.n2955 VSS.n2954 5.15366
R6541 VSS.n2530 VSS.n2529 5.15366
R6542 VSS.n1105 VSS.n1104 5.15366
R6543 VSS.n4032 VSS.n2595 5.14713
R6544 VSS.n2591 VSS.t435 5.14713
R6545 VSS.n4050 VSS.n2429 5.14713
R6546 VSS.n2424 VSS.t1041 5.14713
R6547 VSS.n4103 VSS.n2423 5.14713
R6548 VSS.n4106 VSS.t382 5.14713
R6549 VSS.n2526 VSS.n2441 5.14713
R6550 VSS.n2524 VSS.t597 5.14713
R6551 VSS.n295 VSS.t993 5.14713
R6552 VSS.n5006 VSS.n5004 5.14713
R6553 VSS.n2474 VSS.n2473 5.14713
R6554 VSS.n5077 VSS.n5075 5.14713
R6555 VSS.n5082 VSS.t1408 5.14713
R6556 VSS.n237 VSS.n235 5.14713
R6557 VSS.n232 VSS.t1335 5.14713
R6558 VSS.n5090 VSS.n5089 5.14713
R6559 VSS.n268 VSS.n264 5.14713
R6560 VSS.n271 VSS.n270 5.14713
R6561 VSS.n253 VSS.t1260 5.14713
R6562 VSS.n249 VSS.n247 5.14713
R6563 VSS.n244 VSS.n243 5.14713
R6564 VSS.n289 VSS.n287 5.14713
R6565 VSS.n284 VSS.t1194 5.14713
R6566 VSS.n5024 VSS.n5023 5.14713
R6567 VSS.n5053 VSS.t136 5.14713
R6568 VSS.n5050 VSS.n5047 5.14713
R6569 VSS.n5030 VSS.n5028 5.14713
R6570 VSS.n2522 VSS.n2446 5.14713
R6571 VSS.n2520 VSS.t1035 5.14713
R6572 VSS.n2518 VSS.n2450 5.14713
R6573 VSS.n2516 VSS.t1400 5.14713
R6574 VSS.n2515 VSS.n2461 5.14713
R6575 VSS.n2513 VSS.t655 5.14713
R6576 VSS.n2457 VSS.t602 5.14713
R6577 VSS.n2455 VSS.n2451 5.14713
R6578 VSS.n2454 VSS.t1556 5.14713
R6579 VSS.n2445 VSS.n2444 5.14713
R6580 VSS.n109 VSS.n107 5.14713
R6581 VSS.n104 VSS.t1210 5.14713
R6582 VSS.n4151 VSS.t815 5.14713
R6583 VSS.n4150 VSS.n2290 5.14713
R6584 VSS.n5470 VSS.n17 5.14713
R6585 VSS.n5468 VSS.t683 5.14713
R6586 VSS.n5466 VSS.n21 5.14713
R6587 VSS.n5464 VSS.t635 5.14713
R6588 VSS.n5463 VSS.n32 5.14713
R6589 VSS.n5461 VSS.t628 5.14713
R6590 VSS.n5486 VSS.n5483 5.14713
R6591 VSS.n5490 VSS.t29 5.14713
R6592 VSS.n5 VSS.t888 5.14713
R6593 VSS.n5485 VSS.n5484 5.14713
R6594 VSS.n14 VSS.n13 5.14713
R6595 VSS.n5473 VSS.t714 5.14713
R6596 VSS.n12 VSS.t665 5.14713
R6597 VSS.n8 VSS.n7 5.14713
R6598 VSS.n28 VSS.t719 5.14713
R6599 VSS.n26 VSS.n22 5.14713
R6600 VSS.n25 VSS.t1301 5.14713
R6601 VSS.n16 VSS.n15 5.14713
R6602 VSS.n5454 VSS.n47 5.14713
R6603 VSS.n5439 VSS.t988 5.14713
R6604 VSS.n59 VSS.n57 5.14713
R6605 VSS.n137 VSS.n135 5.14713
R6606 VSS.n142 VSS.t1419 5.14713
R6607 VSS.n190 VSS.n188 5.14713
R6608 VSS.n185 VSS.t1337 5.14713
R6609 VSS.n5394 VSS.n5393 5.14713
R6610 VSS.n5408 VSS.n127 5.14713
R6611 VSS.n202 VSS.t859 5.14713
R6612 VSS.n208 VSS.n206 5.14713
R6613 VSS.n153 VSS.n152 5.14713
R6614 VSS.n162 VSS.t1273 5.14713
R6615 VSS.n158 VSS.n156 5.14713
R6616 VSS.n124 VSS.n123 5.14713
R6617 VSS.n120 VSS.t130 5.14713
R6618 VSS.n5419 VSS.n5417 5.14713
R6619 VSS.n98 VSS.n94 5.14713
R6620 VSS.n71 VSS.n70 5.14713
R6621 VSS.n2540 VSS.n2539 5.14713
R6622 VSS.n2572 VSS.t545 5.14713
R6623 VSS.n2574 VSS.n2573 5.14713
R6624 VSS.n2582 VSS.t1507 5.14713
R6625 VSS.n2584 VSS.n2583 5.14713
R6626 VSS.n2588 VSS.t572 5.14713
R6627 VSS.n2578 VSS.t593 5.14713
R6628 VSS.n2537 VSS.n2536 5.14713
R6629 VSS.n2567 VSS.t44 5.14713
R6630 VSS.n2566 VSS.n2538 5.14713
R6631 VSS.n2542 VSS.n2541 5.14713
R6632 VSS.n2564 VSS.t637 5.14713
R6633 VSS.n2558 VSS.t1509 5.14713
R6634 VSS.n2545 VSS.n2544 5.14713
R6635 VSS.n2548 VSS.n2547 5.14713
R6636 VSS.n2553 VSS.t525 5.14713
R6637 VSS.n2549 VSS.n2546 5.14713
R6638 VSS.n2597 VSS.n2596 5.14713
R6639 VSS.n4030 VSS.t396 5.14713
R6640 VSS.n4024 VSS.t1049 5.14713
R6641 VSS.n2600 VSS.n2599 5.14713
R6642 VSS.n2603 VSS.n2602 5.14713
R6643 VSS.n4019 VSS.t9 5.14713
R6644 VSS.n4015 VSS.n2601 5.14713
R6645 VSS.n2900 VSS.n2899 5.14713
R6646 VSS.n2947 VSS.n2838 5.14713
R6647 VSS.n2945 VSS.t81 5.14713
R6648 VSS.n2943 VSS.n2842 5.14713
R6649 VSS.n2941 VSS.t1151 5.14713
R6650 VSS.n2849 VSS.t1482 5.14713
R6651 VSS.n2847 VSS.n2843 5.14713
R6652 VSS.n2846 VSS.t258 5.14713
R6653 VSS.n2837 VSS.n2836 5.14713
R6654 VSS.n2951 VSS.n2833 5.14713
R6655 VSS.n2949 VSS.t1491 5.14713
R6656 VSS.n2831 VSS.t1161 5.14713
R6657 VSS.n2828 VSS.n2827 5.14713
R6658 VSS.n2826 VSS.n2823 5.14713
R6659 VSS.n2955 VSS.t77 5.14713
R6660 VSS.n2825 VSS.n2824 5.14713
R6661 VSS.n5129 VSS.t850 5.14713
R6662 VSS.n229 VSS.n227 5.14713
R6663 VSS.n2439 VSS.t1386 5.14713
R6664 VSS.n2436 VSS.n2435 5.14713
R6665 VSS.n2434 VSS.n2433 5.14713
R6666 VSS.n2530 VSS.t1379 5.14713
R6667 VSS.n2432 VSS.n2431 5.14713
R6668 VSS.n1091 VSS.n1090 5.14713
R6669 VSS.n1123 VSS.t420 5.14713
R6670 VSS.n1125 VSS.n1124 5.14713
R6671 VSS.n1133 VSS.t1181 5.14713
R6672 VSS.n1135 VSS.n1134 5.14713
R6673 VSS.n1139 VSS.t624 5.14713
R6674 VSS.n1093 VSS.n1092 5.14713
R6675 VSS.n1115 VSS.t633 5.14713
R6676 VSS.n1109 VSS.t1188 5.14713
R6677 VSS.n1096 VSS.n1095 5.14713
R6678 VSS.n1099 VSS.n1098 5.14713
R6679 VSS.n1104 VSS.t313 5.14713
R6680 VSS.n1100 VSS.n1097 5.14713
R6681 VSS.n1129 VSS.t547 5.14713
R6682 VSS.n1088 VSS.n1087 5.14713
R6683 VSS.n1118 VSS.t483 5.14713
R6684 VSS.n1117 VSS.n1089 5.14713
R6685 VSS.n1301 VSS.n1300 5.14713
R6686 VSS.n4039 VSS.t378 5.14713
R6687 VSS.n4038 VSS.n2592 5.14713
R6688 VSS.n4037 VSS.t864 5.14713
R6689 VSS.n2594 VSS.n2593 5.14713
R6690 VSS.n2897 VSS.n2896 5.1454
R6691 VSS.n4431 VSS.n1019 5.1454
R6692 VSS.n4241 VSS.n4240 5.1454
R6693 VSS.n4428 VSS.t788 5.14447
R6694 VSS.n4239 VSS.t915 5.14447
R6695 VSS.n4358 VSS.t982 5.13735
R6696 VSS.n1075 VSS.n1074 5.13413
R6697 VSS.n554 VSS.t1089 5.13148
R6698 VSS.n553 VSS.t1091 5.12074
R6699 VSS.n4456 VSS.n4455 5.08183
R6700 VSS.n4482 VSS.n4481 5.07198
R6701 VSS.n4367 VSS.t285 5.07083
R6702 VSS.n4185 VSS.n4184 5.07083
R6703 VSS.n4522 VSS.t499 5.07083
R6704 VSS.n4200 VSS.t371 5.07083
R6705 VSS.n1039 VSS.t301 5.07083
R6706 VSS.n4483 VSS.t70 5.07083
R6707 VSS.n990 VSS.n989 5.07083
R6708 VSS.n4980 VSS.n332 5.07083
R6709 VSS.n302 VSS.n301 5.07083
R6710 VSS.n1696 VSS.n1695 5.07083
R6711 VSS.n368 VSS.t259 5.07083
R6712 VSS.n4109 VSS.t112 5.07083
R6713 VSS.n3448 VSS.t221 5.07083
R6714 VSS.n1313 VSS.t19 5.05713
R6715 VSS.n1316 VSS.t1232 5.05713
R6716 VSS.n1318 VSS.t738 5.05713
R6717 VSS.n1306 VSS.t1223 5.05713
R6718 VSS.n1325 VSS.t736 5.05713
R6719 VSS.n4364 VSS.t1205 4.92017
R6720 VSS.n2513 VSS.n2512 4.87494
R6721 VSS.n5461 VSS.n5460 4.86394
R6722 VSS.n5138 VSS.n5137 4.86308
R6723 VSS.n3455 VSS.n3454 4.83561
R6724 VSS.n99 VSS.n93 4.70151
R6725 VSS.n773 VSS.t1110 4.65222
R6726 VSS.n4984 VSS.t824 4.65222
R6727 VSS.t1314 VSS.n1722 4.65222
R6728 VSS.n2480 VSS.n2479 4.613
R6729 VSS.n2493 VSS.n2492 4.613
R6730 VSS.n84 VSS.n83 4.613
R6731 VSS.n78 VSS.n77 4.613
R6732 VSS.n1085 VSS.n1084 4.613
R6733 VSS.n5031 VSS.n5027 4.60595
R6734 VSS.n1705 VSS.n1704 4.60233
R6735 VSS.n4465 VSS.n766 4.60233
R6736 VSS.n4992 VSS.n307 4.60233
R6737 VSS.n4194 VSS.n4193 4.60133
R6738 VSS.n4504 VSS.n4503 4.60133
R6739 VSS.n356 VSS.n355 4.60133
R6740 VSS.n4341 VSS.n1712 4.56217
R6741 VSS.n364 VSS.n363 4.56217
R6742 VSS.n4323 VSS.n4322 4.56217
R6743 VSS.n4391 VSS.n4390 4.56217
R6744 VSS.n4462 VSS.n4461 4.56167
R6745 VSS.n4989 VSS.n313 4.56142
R6746 VSS.n4512 VSS.n4511 4.56117
R6747 VSS.n4013 VSS.n4011 4.50944
R6748 VSS.n4499 VSS.n4494 4.50733
R6749 VSS.n1064 VSS.n1063 4.50733
R6750 VSS.n351 VSS.n343 4.50733
R6751 VSS.n1720 VSS.n1719 4.50633
R6752 VSS.n775 VSS.n772 4.50633
R6753 VSS.n4986 VSS.n315 4.50633
R6754 VSS.n2934 VSS.n2852 4.5005
R6755 VSS.n2934 VSS.n2933 4.5005
R6756 VSS.n4390 VSS.n4389 4.5005
R6757 VSS.n4389 VSS.n4388 4.5005
R6758 VSS.n4462 VSS.n770 4.5005
R6759 VSS.n770 VSS.n769 4.5005
R6760 VSS.n4496 VSS.n4495 4.5005
R6761 VSS.n4989 VSS.n4988 4.5005
R6762 VSS.n4988 VSS.n4987 4.5005
R6763 VSS.n5444 VSS.n55 4.5005
R6764 VSS.n5003 VSS.n5002 4.5005
R6765 VSS.n1717 VSS.n1716 4.5005
R6766 VSS.n4322 VSS.n4321 4.5005
R6767 VSS.n4321 VSS.n4320 4.5005
R6768 VSS.n345 VSS.n344 4.5005
R6769 VSS.n4347 VSS.n4346 4.5005
R6770 VSS.n5181 VSS.n5180 4.5005
R6771 VSS.n1766 VSS.n1765 4.5005
R6772 VSS.n5204 VSS.n5203 4.5005
R6773 VSS.n5216 VSS.n5215 4.5005
R6774 VSS.n5193 VSS.n5192 4.5005
R6775 VSS.n2478 VSS.n2477 4.40426
R6776 VSS.n2491 VSS.n2490 4.40426
R6777 VSS.n82 VSS.n81 4.40426
R6778 VSS.n76 VSS.n75 4.40426
R6779 VSS.n1083 VSS.n1082 4.40426
R6780 VSS.n4364 VSS.n4363 4.30289
R6781 VSS.n2589 VSS.n2588 4.27175
R6782 VSS.n1069 VSS.n1068 4.12333
R6783 VSS.n3986 VSS.n3985 4.09657
R6784 VSS.n1313 VSS.n1312 4.07463
R6785 VSS.n2908 VSS.n2903 4.05733
R6786 VSS VSS.n3735 4.0484
R6787 VSS VSS.n4229 4.0484
R6788 VSS VSS.n1730 4.0484
R6789 VSS VSS.n4528 4.0484
R6790 VSS VSS.n2860 4.0484
R6791 VSS VSS.n535 4.0484
R6792 VSS VSS.n4517 4.0484
R6793 VSS VSS.n762 4.0484
R6794 VSS VSS.n999 4.0484
R6795 VSS VSS.n1009 4.0484
R6796 VSS VSS.n4414 4.0484
R6797 VSS VSS.n4380 4.0484
R6798 VSS VSS.n4402 4.0484
R6799 VSS VSS.n325 4.0484
R6800 VSS VSS.n4262 4.0484
R6801 VSS VSS.n4260 4.0484
R6802 VSS VSS.n4972 4.0484
R6803 VSS VSS.n2888 4.0484
R6804 VSS VSS.n1742 4.0484
R6805 VSS VSS.n4210 4.0484
R6806 VSS VSS.n377 4.0484
R6807 VSS.n4969 VSS.t1080 3.99804
R6808 VSS VSS.n2855 3.8414
R6809 VSS.n1711 VSS.n1702 3.83333
R6810 VSS.n4319 VSS.n4191 3.83333
R6811 VSS.n4186 VSS.n4183 3.83333
R6812 VSS.n4510 VSS.n4501 3.83333
R6813 VSS.n4463 VSS.n768 3.83333
R6814 VSS.n4387 VSS.n1066 3.83333
R6815 VSS.n4990 VSS.n309 3.83333
R6816 VSS.n362 VSS.n353 3.83333
R6817 VSS.n4344 VSS.n4343 3.79619
R6818 VSS.n4232 VSS.n4222 3.76876
R6819 VSS.n2510 VSS.n2472 3.76876
R6820 VSS.n2467 VSS.n2464 3.76876
R6821 VSS.n5458 VSS.n39 3.76876
R6822 VSS.n5456 VSS.n45 3.76876
R6823 VSS.n2913 VSS.n2895 3.76876
R6824 VSS.n545 VSS.n539 3.76876
R6825 VSS.n4563 VSS.n556 3.76876
R6826 VSS.n4545 VSS.n748 3.76876
R6827 VSS.n1002 VSS.n1001 3.76876
R6828 VSS.n1005 VSS.n1004 3.76876
R6829 VSS.n1029 VSS.n1028 3.76876
R6830 VSS.n1061 VSS.n1060 3.76876
R6831 VSS.n4425 VSS.n1025 3.76876
R6832 VSS.n4513 VSS.n4492 3.76876
R6833 VSS.n758 VSS.n757 3.76876
R6834 VSS.n4253 VSS.n4252 3.76876
R6835 VSS.n4293 VSS.n4249 3.76876
R6836 VSS.n341 VSS.n340 3.76876
R6837 VSS.n318 VSS.n317 3.76876
R6838 VSS.n4340 VSS.n1714 3.76876
R6839 VSS.n2884 VSS.n2873 3.76876
R6840 VSS.n4324 VSS.n1745 3.76876
R6841 VSS.n4302 VSS.n4213 3.76876
R6842 VSS.n530 VSS.n529 3.76876
R6843 VSS.n2606 VSS.n2605 3.76876
R6844 VSS.n1078 VSS.n1077 3.76485
R6845 VSS.n4006 VSS.n2608 3.75324
R6846 VSS.n4559 VSS.n4558 3.70003
R6847 VSS.n2 VSS.n1 3.66898
R6848 VSS.n4220 VSS.n4219 3.66898
R6849 VSS.n4460 VSS.n777 3.66898
R6850 VSS.n4548 VSS.n4547 3.66898
R6851 VSS.n2906 VSS.n2905 3.66898
R6852 VSS.n543 VSS.n542 3.66898
R6853 VSS.n526 VSS.n525 3.66898
R6854 VSS.n523 VSS.n522 3.66898
R6855 VSS.n4437 VSS.n1013 3.66898
R6856 VSS.n4434 VSS.n1018 3.66898
R6857 VSS.n1023 VSS.n1022 3.66898
R6858 VSS.n4420 VSS.n1032 3.66898
R6859 VSS.n4198 VSS.n4197 3.66898
R6860 VSS.n4393 VSS.n1041 3.66898
R6861 VSS.n753 VSS.n752 3.66898
R6862 VSS.n312 VSS.n311 3.66898
R6863 VSS.n4270 VSS.n4266 3.66898
R6864 VSS.n4300 VSS.n4216 3.66898
R6865 VSS.n4295 VSS.n4247 3.66898
R6866 VSS.n365 VSS.n338 3.66898
R6867 VSS.n4342 VSS.n1700 3.66898
R6868 VSS.n2880 VSS.n2878 3.66898
R6869 VSS.n241 VSS.n240 3.61615
R6870 VSS.n5071 VSS.n262 3.61615
R6871 VSS.n260 VSS.n259 3.61615
R6872 VSS.n5109 VSS.n5108 3.61615
R6873 VSS.n293 VSS.n292 3.61615
R6874 VSS.n282 VSS.n281 3.61615
R6875 VSS.n5448 VSS.n50 3.61615
R6876 VSS.n148 VSS.n147 3.61615
R6877 VSS.n5403 VSS.n130 3.61615
R6878 VSS.n183 VSS.n150 3.61615
R6879 VSS.n174 VSS.n168 3.61615
R6880 VSS.n102 VSS.n68 3.61615
R6881 VSS.n5431 VSS.n65 3.61615
R6882 VSS.n2486 VSS.n2485 3.61615
R6883 VSS.n4371 VSS.n4369 3.60833
R6884 VSS.n374 VSS.n373 3.60833
R6885 VSS.n2918 VSS.n2870 3.60833
R6886 VSS.n1736 VSS.n1725 3.60833
R6887 VSS.n4473 VSS.n4472 3.60833
R6888 VSS.n4535 VSS.n4534 3.60833
R6889 VSS.n4541 VSS.n4524 3.60833
R6890 VSS.n4207 VSS.n4206 3.60833
R6891 VSS.n4399 VSS.n1038 3.60833
R6892 VSS.n1036 VSS.n1035 3.60833
R6893 VSS.n4487 VSS.n4485 3.60833
R6894 VSS.n993 VSS.n783 3.60833
R6895 VSS.n4454 VSS.n781 3.60833
R6896 VSS.n331 VSS.n320 3.60833
R6897 VSS.n4977 VSS.n335 3.60833
R6898 VSS.n4281 VSS.n4280 3.60833
R6899 VSS.n4285 VSS.n4284 3.60833
R6900 VSS.n2867 VSS.n2866 3.60833
R6901 VSS.n4329 VSS.n1739 3.60833
R6902 VSS.n4309 VSS.n4203 3.60833
R6903 VSS.n4964 VSS.n370 3.60833
R6904 VSS.n2293 VSS.n2292 3.60833
R6905 VSS.n3452 VSS.n3450 3.60833
R6906 VSS.n1315 VSS.n1310 3.59463
R6907 VSS.n1317 VSS.n1308 3.59463
R6908 VSS.n1321 VSS.n1320 3.59463
R6909 VSS.n1324 VSS.n1305 3.59463
R6910 VSS.n1329 VSS.n1327 3.59463
R6911 VSS.t118 VSS.n2460 3.57455
R6912 VSS.t71 VSS.n31 3.56931
R6913 VSS.n1328 VSS.n1140 3.45115
R6914 VSS.n4049 VSS.n4048 3.39273
R6915 VSS.n2932 VSS.t1478 3.35794
R6916 VSS.n3751 VSS.t1250 3.22391
R6917 VSS.n5458 VSS.n5457 3.18833
R6918 VSS.n5472 VSS.n10 3.04115
R6919 VSS.n350 VSS.n345 3.01316
R6920 VSS.n360 VSS.n358 3.01316
R6921 VSS.n4317 VSS.n4315 3.01316
R6922 VSS.n1709 VSS.n1707 3.01316
R6923 VSS.n1721 VSS.n1717 3.01316
R6924 VSS.n4498 VSS.n4496 3.01316
R6925 VSS.n4508 VSS.n4506 3.01316
R6926 VSS.n4466 VSS.n764 3.01316
R6927 VSS.n4384 VSS.n1071 3.01316
R6928 VSS.n4993 VSS.n305 3.01316
R6929 VSS.n4357 VSS 2.96831
R6930 VSS.n4344 VSS.n1696 2.93836
R6931 VSS.n5472 VSS.n5471 2.9287
R6932 VSS.n2478 VSS.n2475 2.88323
R6933 VSS.n2491 VSS.n2488 2.88323
R6934 VSS.n82 VSS.n79 2.88323
R6935 VSS.n76 VSS.n73 2.88323
R6936 VSS.n1083 VSS.n1080 2.88323
R6937 VSS.n4046 VSS.n2590 2.77228
R6938 VSS.n5488 VSS.n5487 2.75971
R6939 VSS.n4180 VSS.n4179 2.73113
R6940 VSS.n5481 VSS.n5480 2.6759
R6941 VSS.n4169 VSS.n4166 2.62771
R6942 VSS.n2936 VSS 2.6005
R6943 VSS.n2936 VSS.n2935 2.6005
R6944 VSS.n5196 VSS.n5195 2.6005
R6945 VSS.n5277 VSS.n5276 2.6005
R6946 VSS.n5276 VSS.n5275 2.6005
R6947 VSS.n5274 VSS.n5273 2.6005
R6948 VSS.n5273 VSS.n5272 2.6005
R6949 VSS.n5271 VSS.n5270 2.6005
R6950 VSS.n5270 VSS.n5269 2.6005
R6951 VSS.n5267 VSS.n5266 2.6005
R6952 VSS.n5266 VSS.n5265 2.6005
R6953 VSS.n5264 VSS.n5263 2.6005
R6954 VSS.n5263 VSS.n5262 2.6005
R6955 VSS.n5261 VSS.n5260 2.6005
R6956 VSS.n5260 VSS.n5259 2.6005
R6957 VSS.n5258 VSS.n5257 2.6005
R6958 VSS.n5257 VSS.n5256 2.6005
R6959 VSS.n5255 VSS.n5254 2.6005
R6960 VSS.n5254 VSS.n5253 2.6005
R6961 VSS.n5252 VSS.n5251 2.6005
R6962 VSS.n5251 VSS.n5250 2.6005
R6963 VSS.n5249 VSS.n5248 2.6005
R6964 VSS.n5248 VSS.n5247 2.6005
R6965 VSS.n5246 VSS.n5245 2.6005
R6966 VSS.n5245 VSS.n5244 2.6005
R6967 VSS.n5243 VSS.n5242 2.6005
R6968 VSS.n5242 VSS.n5241 2.6005
R6969 VSS.n5240 VSS.n5239 2.6005
R6970 VSS.n5239 VSS.n5238 2.6005
R6971 VSS.n5237 VSS.n5236 2.6005
R6972 VSS.n5236 VSS.n5235 2.6005
R6973 VSS.n5234 VSS.n5233 2.6005
R6974 VSS.n5233 VSS.n5232 2.6005
R6975 VSS.n5231 VSS.n5230 2.6005
R6976 VSS.n5230 VSS.n5229 2.6005
R6977 VSS.n5228 VSS.n5227 2.6005
R6978 VSS.n5227 VSS.n5226 2.6005
R6979 VSS.n5225 VSS.n5224 2.6005
R6980 VSS.n5224 VSS.n5223 2.6005
R6981 VSS.n5219 VSS.n5218 2.6005
R6982 VSS.n5218 VSS.n5217 2.6005
R6983 VSS.n5207 VSS.n5206 2.6005
R6984 VSS.n5206 VSS.n5205 2.6005
R6985 VSS.n3759 VSS.n3758 2.6005
R6986 VSS.n3758 VSS.n3757 2.6005
R6987 VSS.n3756 VSS.n3755 2.6005
R6988 VSS.n3755 VSS.n3754 2.6005
R6989 VSS.n3753 VSS.n3752 2.6005
R6990 VSS.n3752 VSS.n3751 2.6005
R6991 VSS.n3750 VSS.n3749 2.6005
R6992 VSS.n3749 VSS.n3748 2.6005
R6993 VSS.n3747 VSS.n3746 2.6005
R6994 VSS.n3746 VSS.n3745 2.6005
R6995 VSS.n3744 VSS.n3743 2.6005
R6996 VSS.n3743 VSS.n3742 2.6005
R6997 VSS.n3741 VSS.n3740 2.6005
R6998 VSS.n3740 VSS.n3739 2.6005
R6999 VSS.n3733 VSS.n3732 2.6005
R7000 VSS.n3730 VSS.n3729 2.6005
R7001 VSS.n3728 VSS.n3727 2.6005
R7002 VSS.n3724 VSS.n3723 2.6005
R7003 VSS.n3723 VSS.n3722 2.6005
R7004 VSS.n3720 VSS.n3719 2.6005
R7005 VSS.n3719 VSS.n3718 2.6005
R7006 VSS.n3717 VSS.n3716 2.6005
R7007 VSS.n3716 VSS.n3715 2.6005
R7008 VSS.n3714 VSS.n3713 2.6005
R7009 VSS.n3713 VSS.n3712 2.6005
R7010 VSS.n3711 VSS.n3710 2.6005
R7011 VSS.n3710 VSS.n3709 2.6005
R7012 VSS.n3708 VSS.n3707 2.6005
R7013 VSS.n3707 VSS.n3706 2.6005
R7014 VSS.n3705 VSS.n3704 2.6005
R7015 VSS.n3704 VSS.n3703 2.6005
R7016 VSS.n3702 VSS.n3701 2.6005
R7017 VSS.n3701 VSS.n3700 2.6005
R7018 VSS.n3699 VSS.n3698 2.6005
R7019 VSS.n3698 VSS.n3697 2.6005
R7020 VSS.n3696 VSS.n3695 2.6005
R7021 VSS.n3695 VSS.n3694 2.6005
R7022 VSS.n3693 VSS.n3692 2.6005
R7023 VSS.n3692 VSS.n3691 2.6005
R7024 VSS.n3690 VSS.n3689 2.6005
R7025 VSS.n3689 VSS.n3688 2.6005
R7026 VSS.n3687 VSS.n3686 2.6005
R7027 VSS.n3686 VSS.n3685 2.6005
R7028 VSS.n3684 VSS.n3683 2.6005
R7029 VSS.n3683 VSS.n3682 2.6005
R7030 VSS.n3681 VSS.n3680 2.6005
R7031 VSS.n3680 VSS.n3679 2.6005
R7032 VSS.n3678 VSS.n3677 2.6005
R7033 VSS.n3677 VSS.n3676 2.6005
R7034 VSS.n3675 VSS.n3674 2.6005
R7035 VSS.n3674 VSS.n3673 2.6005
R7036 VSS.n3672 VSS.n3671 2.6005
R7037 VSS.n3671 VSS.n3670 2.6005
R7038 VSS.n3669 VSS.n3668 2.6005
R7039 VSS.n3668 VSS.n3667 2.6005
R7040 VSS.n3666 VSS.n3665 2.6005
R7041 VSS.n3665 VSS.n3664 2.6005
R7042 VSS.n3663 VSS.n3662 2.6005
R7043 VSS.n3662 VSS.n3661 2.6005
R7044 VSS.n3660 VSS.n3659 2.6005
R7045 VSS.n3659 VSS.n3658 2.6005
R7046 VSS.n3657 VSS.n3656 2.6005
R7047 VSS.n3656 VSS.n3655 2.6005
R7048 VSS.n3654 VSS.n3653 2.6005
R7049 VSS.n3653 VSS.n3652 2.6005
R7050 VSS.n3651 VSS.n3650 2.6005
R7051 VSS.n3650 VSS.n3649 2.6005
R7052 VSS.n3648 VSS.n3647 2.6005
R7053 VSS.n3647 VSS.n3646 2.6005
R7054 VSS.n3645 VSS.n3644 2.6005
R7055 VSS.n3644 VSS.n3643 2.6005
R7056 VSS.n3642 VSS.n3641 2.6005
R7057 VSS.n3641 VSS.n3640 2.6005
R7058 VSS.n3639 VSS.n3638 2.6005
R7059 VSS.n3638 VSS.n3637 2.6005
R7060 VSS.n3636 VSS.n3635 2.6005
R7061 VSS.n3635 VSS.n3634 2.6005
R7062 VSS.n3633 VSS.n3632 2.6005
R7063 VSS.n3632 VSS.n3631 2.6005
R7064 VSS.n3630 VSS.n3629 2.6005
R7065 VSS.n3629 VSS.n3628 2.6005
R7066 VSS.n3627 VSS.n3626 2.6005
R7067 VSS.n3626 VSS.n3625 2.6005
R7068 VSS.n3624 VSS.n3623 2.6005
R7069 VSS.n3623 VSS.n3622 2.6005
R7070 VSS.n3621 VSS.n3620 2.6005
R7071 VSS.n3620 VSS.n3619 2.6005
R7072 VSS.n3618 VSS.n3617 2.6005
R7073 VSS.n3617 VSS.n3616 2.6005
R7074 VSS.n3615 VSS.n3614 2.6005
R7075 VSS.n3614 VSS.n3613 2.6005
R7076 VSS.n3612 VSS.n3611 2.6005
R7077 VSS.n3611 VSS.n3610 2.6005
R7078 VSS.n3609 VSS.n3608 2.6005
R7079 VSS.n3608 VSS.n3607 2.6005
R7080 VSS.n3606 VSS.n3605 2.6005
R7081 VSS.n3605 VSS.n3604 2.6005
R7082 VSS.n3603 VSS.n3602 2.6005
R7083 VSS.n3602 VSS.n3601 2.6005
R7084 VSS.n3600 VSS.n3599 2.6005
R7085 VSS.n3599 VSS.n3598 2.6005
R7086 VSS.n3597 VSS.n3596 2.6005
R7087 VSS.n3596 VSS.n3595 2.6005
R7088 VSS.n3594 VSS.n3593 2.6005
R7089 VSS.n3593 VSS.n3592 2.6005
R7090 VSS.n3591 VSS.n3590 2.6005
R7091 VSS.n3590 VSS.n3589 2.6005
R7092 VSS.n3588 VSS.n3587 2.6005
R7093 VSS.n3587 VSS.n3586 2.6005
R7094 VSS.n3585 VSS.n3584 2.6005
R7095 VSS.n3584 VSS.n3583 2.6005
R7096 VSS.n3582 VSS.n3581 2.6005
R7097 VSS.n3581 VSS.n3580 2.6005
R7098 VSS.n3579 VSS.n3578 2.6005
R7099 VSS.n3578 VSS.n3577 2.6005
R7100 VSS.n3576 VSS.n3575 2.6005
R7101 VSS.n3575 VSS.n3574 2.6005
R7102 VSS.n3573 VSS.n3572 2.6005
R7103 VSS.n3572 VSS.n3571 2.6005
R7104 VSS.n3570 VSS.n3569 2.6005
R7105 VSS.n3569 VSS.n3568 2.6005
R7106 VSS.n3567 VSS.n3566 2.6005
R7107 VSS.n3566 VSS.n3565 2.6005
R7108 VSS.n3562 VSS.n3561 2.6005
R7109 VSS.n3561 VSS.n3560 2.6005
R7110 VSS.n3557 VSS.n3556 2.6005
R7111 VSS.n3556 VSS.n3555 2.6005
R7112 VSS.n3554 VSS.n3553 2.6005
R7113 VSS.n3553 VSS.n3552 2.6005
R7114 VSS.n3549 VSS.n3548 2.6005
R7115 VSS.n3548 VSS.n3547 2.6005
R7116 VSS.n3532 VSS.n3531 2.6005
R7117 VSS.n3531 VSS.n3530 2.6005
R7118 VSS.n3529 VSS.n3528 2.6005
R7119 VSS.n3528 VSS.n3527 2.6005
R7120 VSS.n3526 VSS.n3525 2.6005
R7121 VSS.n3525 VSS.n3524 2.6005
R7122 VSS.n3523 VSS.n3522 2.6005
R7123 VSS.n3522 VSS.n3521 2.6005
R7124 VSS.n2427 VSS.n2426 2.6005
R7125 VSS.n2426 VSS.n2425 2.6005
R7126 VSS.n4056 VSS.n4055 2.6005
R7127 VSS.n4055 VSS.n4054 2.6005
R7128 VSS.n4100 VSS.n4099 2.6005
R7129 VSS.n4101 VSS.n4100 2.6005
R7130 VSS.n4098 VSS.n4097 2.6005
R7131 VSS.n4097 VSS.n4096 2.6005
R7132 VSS.n4095 VSS.n4094 2.6005
R7133 VSS.n4094 VSS.n4093 2.6005
R7134 VSS.n4092 VSS.n4091 2.6005
R7135 VSS.n4091 VSS.n4090 2.6005
R7136 VSS.n4088 VSS.t392 2.6005
R7137 VSS.n4089 VSS.n4088 2.6005
R7138 VSS.n4087 VSS.n4086 2.6005
R7139 VSS.n4086 VSS.n4085 2.6005
R7140 VSS.n4084 VSS.n4083 2.6005
R7141 VSS.n4083 VSS.n4082 2.6005
R7142 VSS.n4081 VSS.n4080 2.6005
R7143 VSS.n4080 VSS.n4079 2.6005
R7144 VSS.n4078 VSS.n4077 2.6005
R7145 VSS.n4077 VSS.n4076 2.6005
R7146 VSS.n4075 VSS.n4074 2.6005
R7147 VSS.n4074 VSS.n4073 2.6005
R7148 VSS.n4072 VSS.n4071 2.6005
R7149 VSS.n4071 VSS.n4070 2.6005
R7150 VSS.n4069 VSS.n4068 2.6005
R7151 VSS.n4068 VSS.n4067 2.6005
R7152 VSS.n4066 VSS.n4065 2.6005
R7153 VSS.n4065 VSS.n4064 2.6005
R7154 VSS.n4062 VSS.n4061 2.6005
R7155 VSS.n4061 VSS.n4060 2.6005
R7156 VSS.n4059 VSS.n4058 2.6005
R7157 VSS.n4058 VSS.n4057 2.6005
R7158 VSS.n2422 VSS.n2421 2.6005
R7159 VSS.n2421 VSS.n2420 2.6005
R7160 VSS.n4112 VSS.n4111 2.6005
R7161 VSS.n4114 VSS.n4113 2.6005
R7162 VSS.n4119 VSS.n4118 2.6005
R7163 VSS.n4118 VSS.n4117 2.6005
R7164 VSS.n4122 VSS.n4121 2.6005
R7165 VSS.n4121 VSS.n4120 2.6005
R7166 VSS.n4125 VSS.n4124 2.6005
R7167 VSS.n4124 VSS.n4123 2.6005
R7168 VSS.n4128 VSS.n4127 2.6005
R7169 VSS.n4127 VSS.n4126 2.6005
R7170 VSS.n4131 VSS.n4130 2.6005
R7171 VSS.n4130 VSS.n4129 2.6005
R7172 VSS.n4134 VSS.n4133 2.6005
R7173 VSS.n4133 VSS.n4132 2.6005
R7174 VSS.n4137 VSS.n4136 2.6005
R7175 VSS.n4136 VSS.n4135 2.6005
R7176 VSS.n4141 VSS.n4140 2.6005
R7177 VSS.n4140 VSS.n4139 2.6005
R7178 VSS.n4145 VSS.n4144 2.6005
R7179 VSS.n2419 VSS.n2418 2.6005
R7180 VSS.n2417 VSS.n2416 2.6005
R7181 VSS.n2414 VSS.n2413 2.6005
R7182 VSS.n2412 VSS.n2411 2.6005
R7183 VSS.n2409 VSS.n2408 2.6005
R7184 VSS.n2407 VSS.n2406 2.6005
R7185 VSS.n2406 VSS.n2405 2.6005
R7186 VSS.n2403 VSS.n2402 2.6005
R7187 VSS.n2402 VSS.n2401 2.6005
R7188 VSS.n2400 VSS.n2399 2.6005
R7189 VSS.n2399 VSS.n2398 2.6005
R7190 VSS.n2397 VSS.n2396 2.6005
R7191 VSS.n2396 VSS.n2395 2.6005
R7192 VSS.n2394 VSS.n2393 2.6005
R7193 VSS.n2393 VSS.n2392 2.6005
R7194 VSS.n2387 VSS.n2386 2.6005
R7195 VSS.n2389 VSS.n2388 2.6005
R7196 VSS.n2385 VSS.n2384 2.6005
R7197 VSS.n2384 VSS.n2383 2.6005
R7198 VSS.n2382 VSS.n2381 2.6005
R7199 VSS.n2381 VSS.n2380 2.6005
R7200 VSS.n2379 VSS.n2378 2.6005
R7201 VSS.n2378 VSS.n2377 2.6005
R7202 VSS.n2376 VSS.n2375 2.6005
R7203 VSS.n2375 VSS.n2374 2.6005
R7204 VSS.n2373 VSS.n2372 2.6005
R7205 VSS.n2372 VSS.n2371 2.6005
R7206 VSS.n2370 VSS.n2369 2.6005
R7207 VSS.n2369 VSS.n2368 2.6005
R7208 VSS.n2367 VSS.n2366 2.6005
R7209 VSS.n2366 VSS.n2365 2.6005
R7210 VSS.n2364 VSS.n2363 2.6005
R7211 VSS.n2363 VSS.n2362 2.6005
R7212 VSS.n2360 VSS.n2359 2.6005
R7213 VSS.n2359 VSS.n2358 2.6005
R7214 VSS.n2357 VSS.n2356 2.6005
R7215 VSS.n2356 VSS.n2355 2.6005
R7216 VSS.n2354 VSS.n2353 2.6005
R7217 VSS.n2353 VSS.n2352 2.6005
R7218 VSS.n2351 VSS.n2350 2.6005
R7219 VSS.n2350 VSS.n2349 2.6005
R7220 VSS.n2348 VSS.n2347 2.6005
R7221 VSS.n2347 VSS.n2346 2.6005
R7222 VSS.n2345 VSS.n2344 2.6005
R7223 VSS.n2344 VSS.n2343 2.6005
R7224 VSS.n2342 VSS.n2341 2.6005
R7225 VSS.n2341 VSS.n2340 2.6005
R7226 VSS.n2338 VSS.n2337 2.6005
R7227 VSS.n2337 VSS.n2336 2.6005
R7228 VSS.n2335 VSS.n2334 2.6005
R7229 VSS.n2334 VSS.n2333 2.6005
R7230 VSS.n2332 VSS.n2331 2.6005
R7231 VSS.n2331 VSS.n2330 2.6005
R7232 VSS.n2329 VSS.n2328 2.6005
R7233 VSS.n2328 VSS.n2327 2.6005
R7234 VSS.n2326 VSS.n2325 2.6005
R7235 VSS.n2325 VSS.n2324 2.6005
R7236 VSS.n2323 VSS.n2322 2.6005
R7237 VSS.n2322 VSS.n2321 2.6005
R7238 VSS.n2316 VSS.n2315 2.6005
R7239 VSS.n2315 VSS.n2314 2.6005
R7240 VSS.n2307 VSS.n2306 2.6005
R7241 VSS.n2306 VSS.n2305 2.6005
R7242 VSS.n2304 VSS.n2303 2.6005
R7243 VSS.n2303 VSS.n2302 2.6005
R7244 VSS.n1753 VSS.n1752 2.6005
R7245 VSS.n1752 VSS.n1751 2.6005
R7246 VSS.n4169 VSS.n4168 2.6005
R7247 VSS.n4168 VSS.n4167 2.6005
R7248 VSS.n4166 VSS.n4165 2.6005
R7249 VSS.n4165 VSS.n4164 2.6005
R7250 VSS.n4163 VSS.n4162 2.6005
R7251 VSS.n4162 VSS.n4161 2.6005
R7252 VSS.n4160 VSS.n4159 2.6005
R7253 VSS.n4159 VSS.n4158 2.6005
R7254 VSS.n4157 VSS.n4156 2.6005
R7255 VSS.n4156 VSS.n4155 2.6005
R7256 VSS.n2289 VSS.n2288 2.6005
R7257 VSS.n2288 VSS.n2287 2.6005
R7258 VSS.n2286 VSS.n2285 2.6005
R7259 VSS.n2285 VSS.n2284 2.6005
R7260 VSS.n2283 VSS.n2282 2.6005
R7261 VSS.n2282 VSS.n2281 2.6005
R7262 VSS.n2280 VSS.n2279 2.6005
R7263 VSS.n2279 VSS.n2278 2.6005
R7264 VSS.n2277 VSS.n2276 2.6005
R7265 VSS.n2276 VSS.n2275 2.6005
R7266 VSS.n2274 VSS.n2273 2.6005
R7267 VSS.n2273 VSS.n2272 2.6005
R7268 VSS.n2271 VSS.n2270 2.6005
R7269 VSS.n2270 VSS.n2269 2.6005
R7270 VSS.n2268 VSS.n2267 2.6005
R7271 VSS.n2267 VSS.n2266 2.6005
R7272 VSS.n2265 VSS.n2264 2.6005
R7273 VSS.n2264 VSS.n2263 2.6005
R7274 VSS.n2262 VSS.n2261 2.6005
R7275 VSS.n2261 VSS.n2260 2.6005
R7276 VSS.n2259 VSS.n2258 2.6005
R7277 VSS.n2258 VSS.n2257 2.6005
R7278 VSS.n2256 VSS.n2255 2.6005
R7279 VSS.n2255 VSS.n2254 2.6005
R7280 VSS.n2253 VSS.n2252 2.6005
R7281 VSS.n2252 VSS.n2251 2.6005
R7282 VSS.n2250 VSS.n2249 2.6005
R7283 VSS.n2249 VSS.n2248 2.6005
R7284 VSS.n2247 VSS.n2246 2.6005
R7285 VSS.n2246 VSS.n2245 2.6005
R7286 VSS.n2244 VSS.n2243 2.6005
R7287 VSS.n2243 VSS.n2242 2.6005
R7288 VSS.n2241 VSS.n2240 2.6005
R7289 VSS.n2240 VSS.n2239 2.6005
R7290 VSS.n2238 VSS.n2237 2.6005
R7291 VSS.n2237 VSS.n2236 2.6005
R7292 VSS.n2235 VSS.n2234 2.6005
R7293 VSS.n2234 VSS.n2233 2.6005
R7294 VSS.n2232 VSS.n2231 2.6005
R7295 VSS.n2231 VSS.n2230 2.6005
R7296 VSS.n2229 VSS.n2228 2.6005
R7297 VSS.n2228 VSS.n2227 2.6005
R7298 VSS.n2226 VSS.n2225 2.6005
R7299 VSS.n2225 VSS.n2224 2.6005
R7300 VSS.n2223 VSS.n2222 2.6005
R7301 VSS.n2222 VSS.n2221 2.6005
R7302 VSS.n2220 VSS.n2219 2.6005
R7303 VSS.n2219 VSS.n2218 2.6005
R7304 VSS.n2217 VSS.n2216 2.6005
R7305 VSS.n2216 VSS.n2215 2.6005
R7306 VSS.n2214 VSS.n2213 2.6005
R7307 VSS.n2213 VSS.n2212 2.6005
R7308 VSS.n2211 VSS.n2210 2.6005
R7309 VSS.n2210 VSS.n2209 2.6005
R7310 VSS.n2208 VSS.n2207 2.6005
R7311 VSS.n2207 VSS.n2206 2.6005
R7312 VSS.n2205 VSS.n2204 2.6005
R7313 VSS.n2204 VSS.n2203 2.6005
R7314 VSS.n2202 VSS.n2201 2.6005
R7315 VSS.n2201 VSS.n2200 2.6005
R7316 VSS.n2199 VSS.n2198 2.6005
R7317 VSS.n2198 VSS.n2197 2.6005
R7318 VSS.n2196 VSS.n2195 2.6005
R7319 VSS.n2195 VSS.n2194 2.6005
R7320 VSS.n2193 VSS.n2192 2.6005
R7321 VSS.n2192 VSS.n2191 2.6005
R7322 VSS.n2190 VSS.n2189 2.6005
R7323 VSS.n2189 VSS.n2188 2.6005
R7324 VSS.n2187 VSS.n2186 2.6005
R7325 VSS.n2186 VSS.n2185 2.6005
R7326 VSS.n2184 VSS.n2183 2.6005
R7327 VSS.n2183 VSS.n2182 2.6005
R7328 VSS.n2181 VSS.n2180 2.6005
R7329 VSS.n2180 VSS.n2179 2.6005
R7330 VSS.n2178 VSS.n2177 2.6005
R7331 VSS.n2177 VSS.n2176 2.6005
R7332 VSS.n2175 VSS.n2174 2.6005
R7333 VSS.n2174 VSS.n2173 2.6005
R7334 VSS.n2172 VSS.n2171 2.6005
R7335 VSS.n2171 VSS.n2170 2.6005
R7336 VSS.n2169 VSS.n2168 2.6005
R7337 VSS.n2168 VSS.n2167 2.6005
R7338 VSS.n2166 VSS.n2165 2.6005
R7339 VSS.n2165 VSS.n2164 2.6005
R7340 VSS.n2163 VSS.n2162 2.6005
R7341 VSS.n2162 VSS.n2161 2.6005
R7342 VSS.n2160 VSS.n2159 2.6005
R7343 VSS.n2159 VSS.n2158 2.6005
R7344 VSS.n2157 VSS.n2156 2.6005
R7345 VSS.n2156 VSS.n2155 2.6005
R7346 VSS.n2154 VSS.n2153 2.6005
R7347 VSS.n2153 VSS.n2152 2.6005
R7348 VSS.n2151 VSS.n2150 2.6005
R7349 VSS.n2150 VSS.n2149 2.6005
R7350 VSS.n2148 VSS.n2147 2.6005
R7351 VSS.n2147 VSS.n2146 2.6005
R7352 VSS.n2145 VSS.n2144 2.6005
R7353 VSS.n2144 VSS.n2143 2.6005
R7354 VSS.n2142 VSS.n2141 2.6005
R7355 VSS.n2141 VSS.n2140 2.6005
R7356 VSS.n2139 VSS.n2138 2.6005
R7357 VSS.n2138 VSS.n2137 2.6005
R7358 VSS.n2136 VSS.n2135 2.6005
R7359 VSS.n2135 VSS.n2134 2.6005
R7360 VSS.n2133 VSS.n2132 2.6005
R7361 VSS.n2132 VSS.n2131 2.6005
R7362 VSS.n2130 VSS.n2129 2.6005
R7363 VSS.n2129 VSS.n2128 2.6005
R7364 VSS.n2127 VSS.n2126 2.6005
R7365 VSS.n2126 VSS.n2125 2.6005
R7366 VSS.n2124 VSS.n2123 2.6005
R7367 VSS.n2123 VSS.n2122 2.6005
R7368 VSS.n2121 VSS.n2120 2.6005
R7369 VSS.n2120 VSS.n2119 2.6005
R7370 VSS.n2118 VSS.n2117 2.6005
R7371 VSS.n2117 VSS.n2116 2.6005
R7372 VSS.n2115 VSS.n2114 2.6005
R7373 VSS.n2114 VSS.n2113 2.6005
R7374 VSS.n2112 VSS.n2111 2.6005
R7375 VSS.n2111 VSS.n2110 2.6005
R7376 VSS.n2109 VSS.n2108 2.6005
R7377 VSS.n2108 VSS.n2107 2.6005
R7378 VSS.n2106 VSS.n2105 2.6005
R7379 VSS.n2105 VSS.n2104 2.6005
R7380 VSS.n2103 VSS.n2102 2.6005
R7381 VSS.n2102 VSS.n2101 2.6005
R7382 VSS.n2100 VSS.n2099 2.6005
R7383 VSS.n2099 VSS.n2098 2.6005
R7384 VSS.n2097 VSS.n2096 2.6005
R7385 VSS.n2096 VSS.n2095 2.6005
R7386 VSS.n2094 VSS.n2093 2.6005
R7387 VSS.n2093 VSS.n2092 2.6005
R7388 VSS.n2091 VSS.n2090 2.6005
R7389 VSS.n2090 VSS.n2089 2.6005
R7390 VSS.n2088 VSS.n2087 2.6005
R7391 VSS.n2087 VSS.n2086 2.6005
R7392 VSS.n2085 VSS.n2084 2.6005
R7393 VSS.n2084 VSS.n2083 2.6005
R7394 VSS.n2082 VSS.n2081 2.6005
R7395 VSS.n2081 VSS.n2080 2.6005
R7396 VSS.n2079 VSS.n2078 2.6005
R7397 VSS.n2078 VSS.n2077 2.6005
R7398 VSS.n2076 VSS.n2075 2.6005
R7399 VSS.n2075 VSS.n2074 2.6005
R7400 VSS.n2067 VSS.n2066 2.6005
R7401 VSS.n2066 VSS.n2065 2.6005
R7402 VSS.n2064 VSS.n2063 2.6005
R7403 VSS.n2063 VSS.n2062 2.6005
R7404 VSS.n2055 VSS.n2054 2.6005
R7405 VSS.n2054 VSS.n2053 2.6005
R7406 VSS.n2046 VSS.n2045 2.6005
R7407 VSS.n2045 VSS.n2044 2.6005
R7408 VSS.n2040 VSS.n2039 2.6005
R7409 VSS.n2039 VSS.n2038 2.6005
R7410 VSS.n2037 VSS.n2036 2.6005
R7411 VSS.n2036 VSS.n2035 2.6005
R7412 VSS.n2034 VSS.n2033 2.6005
R7413 VSS.n2033 VSS.n2032 2.6005
R7414 VSS.n2031 VSS.n2030 2.6005
R7415 VSS.n2030 VSS.n2029 2.6005
R7416 VSS.n2028 VSS.n2027 2.6005
R7417 VSS.n2027 VSS.n2026 2.6005
R7418 VSS.n2025 VSS.n2024 2.6005
R7419 VSS.n2024 VSS.n2023 2.6005
R7420 VSS.n2022 VSS.n2021 2.6005
R7421 VSS.n2021 VSS.n2020 2.6005
R7422 VSS.n2019 VSS.n2018 2.6005
R7423 VSS.n2018 VSS.n2017 2.6005
R7424 VSS.n2016 VSS.n2015 2.6005
R7425 VSS.n2015 VSS.n2014 2.6005
R7426 VSS.n2013 VSS.n2012 2.6005
R7427 VSS.n2012 VSS.n2011 2.6005
R7428 VSS.n2010 VSS.n2009 2.6005
R7429 VSS.n2009 VSS.n2008 2.6005
R7430 VSS.n2007 VSS.n2006 2.6005
R7431 VSS.n2006 VSS.n2005 2.6005
R7432 VSS.n2004 VSS.n2003 2.6005
R7433 VSS.n2003 VSS.n2002 2.6005
R7434 VSS.n2001 VSS.n2000 2.6005
R7435 VSS.n2000 VSS.n1999 2.6005
R7436 VSS.n1998 VSS.n1997 2.6005
R7437 VSS.n1997 VSS.n1996 2.6005
R7438 VSS.n1995 VSS.n1994 2.6005
R7439 VSS.n1994 VSS.n1993 2.6005
R7440 VSS.n1992 VSS.n1991 2.6005
R7441 VSS.n1991 VSS.n1990 2.6005
R7442 VSS.n1989 VSS.n1988 2.6005
R7443 VSS.n1988 VSS.n1987 2.6005
R7444 VSS.n1986 VSS.n1985 2.6005
R7445 VSS.n1985 VSS.n1984 2.6005
R7446 VSS.n1983 VSS.n1982 2.6005
R7447 VSS.n1982 VSS.n1981 2.6005
R7448 VSS.n1980 VSS.n1979 2.6005
R7449 VSS.n1979 VSS.n1978 2.6005
R7450 VSS.n1977 VSS.n1976 2.6005
R7451 VSS.n1976 VSS.n1975 2.6005
R7452 VSS.n1974 VSS.n1973 2.6005
R7453 VSS.n1973 VSS.n1972 2.6005
R7454 VSS.n1971 VSS.n1970 2.6005
R7455 VSS.n1970 VSS.n1969 2.6005
R7456 VSS.n1968 VSS.n1967 2.6005
R7457 VSS.n1967 VSS.n1966 2.6005
R7458 VSS.n1965 VSS.n1964 2.6005
R7459 VSS.n1964 VSS.n1963 2.6005
R7460 VSS.n1962 VSS.n1961 2.6005
R7461 VSS.n1961 VSS.n1960 2.6005
R7462 VSS.n1959 VSS.n1958 2.6005
R7463 VSS.n1958 VSS.n1957 2.6005
R7464 VSS.n1956 VSS.n1955 2.6005
R7465 VSS.n1955 VSS.n1954 2.6005
R7466 VSS.n1953 VSS.n1952 2.6005
R7467 VSS.n1952 VSS.n1951 2.6005
R7468 VSS.n1950 VSS.n1949 2.6005
R7469 VSS.n1949 VSS.n1948 2.6005
R7470 VSS.n1947 VSS.n1946 2.6005
R7471 VSS.n1946 VSS.n1945 2.6005
R7472 VSS.n1944 VSS.n1943 2.6005
R7473 VSS.n1943 VSS.n1942 2.6005
R7474 VSS.n1941 VSS.n1940 2.6005
R7475 VSS.n1940 VSS.n1939 2.6005
R7476 VSS.n1938 VSS.n1937 2.6005
R7477 VSS.n1937 VSS.n1936 2.6005
R7478 VSS.n1935 VSS.n1934 2.6005
R7479 VSS.n1934 VSS.n1933 2.6005
R7480 VSS.n1932 VSS.n1931 2.6005
R7481 VSS.n1931 VSS.n1930 2.6005
R7482 VSS.n1929 VSS.n1928 2.6005
R7483 VSS.n1928 VSS.n1927 2.6005
R7484 VSS.n1926 VSS.n1925 2.6005
R7485 VSS.n1925 VSS.n1924 2.6005
R7486 VSS.n1923 VSS.n1922 2.6005
R7487 VSS.n1922 VSS.n1921 2.6005
R7488 VSS.n1920 VSS.n1919 2.6005
R7489 VSS.n1919 VSS.n1918 2.6005
R7490 VSS.n1917 VSS.n1916 2.6005
R7491 VSS.n1916 VSS.n1915 2.6005
R7492 VSS.n1914 VSS.n1913 2.6005
R7493 VSS.n1913 VSS.n1912 2.6005
R7494 VSS.n1911 VSS.n1910 2.6005
R7495 VSS.n1910 VSS.n1909 2.6005
R7496 VSS.n1908 VSS.n1907 2.6005
R7497 VSS.n1907 VSS.n1906 2.6005
R7498 VSS.n1905 VSS.n1904 2.6005
R7499 VSS.n1904 VSS.n1903 2.6005
R7500 VSS.n1902 VSS.n1901 2.6005
R7501 VSS.n1901 VSS.n1900 2.6005
R7502 VSS.n1899 VSS.n1898 2.6005
R7503 VSS.n1898 VSS.n1897 2.6005
R7504 VSS.n1896 VSS.n1895 2.6005
R7505 VSS.n1895 VSS.n1894 2.6005
R7506 VSS.n1893 VSS.n1892 2.6005
R7507 VSS.n1892 VSS.n1891 2.6005
R7508 VSS.n1890 VSS.n1889 2.6005
R7509 VSS.n1889 VSS.n1888 2.6005
R7510 VSS.n1887 VSS.n1886 2.6005
R7511 VSS.n1886 VSS.n1885 2.6005
R7512 VSS.n1884 VSS.n1883 2.6005
R7513 VSS.n1883 VSS.n1882 2.6005
R7514 VSS.n1881 VSS.n1880 2.6005
R7515 VSS.n1880 VSS.n1879 2.6005
R7516 VSS.n1878 VSS.n1877 2.6005
R7517 VSS.n1877 VSS.n1876 2.6005
R7518 VSS.n1875 VSS.n1874 2.6005
R7519 VSS.n1874 VSS.n1873 2.6005
R7520 VSS.n1872 VSS.n1871 2.6005
R7521 VSS.n1871 VSS.n1870 2.6005
R7522 VSS.n1869 VSS.n1868 2.6005
R7523 VSS.n1868 VSS.n1867 2.6005
R7524 VSS.n1866 VSS.n1865 2.6005
R7525 VSS.n1865 VSS.n1864 2.6005
R7526 VSS.n1863 VSS.n1862 2.6005
R7527 VSS.n1862 VSS.n1861 2.6005
R7528 VSS.n1860 VSS.n1859 2.6005
R7529 VSS.n1859 VSS.n1858 2.6005
R7530 VSS.n1857 VSS.n1856 2.6005
R7531 VSS.n1856 VSS.n1855 2.6005
R7532 VSS.n1854 VSS.n1853 2.6005
R7533 VSS.n1853 VSS.n1852 2.6005
R7534 VSS.n1851 VSS.n1850 2.6005
R7535 VSS.n1850 VSS.n1849 2.6005
R7536 VSS.n1848 VSS.n1847 2.6005
R7537 VSS.n1847 VSS.n1846 2.6005
R7538 VSS.n1845 VSS.n1844 2.6005
R7539 VSS.n1844 VSS.n1843 2.6005
R7540 VSS.n1842 VSS.n1841 2.6005
R7541 VSS.n1841 VSS.n1840 2.6005
R7542 VSS.n1839 VSS.n1838 2.6005
R7543 VSS.n1838 VSS.n1837 2.6005
R7544 VSS.n1836 VSS.n1835 2.6005
R7545 VSS.n1835 VSS.n1834 2.6005
R7546 VSS.n1833 VSS.n1832 2.6005
R7547 VSS.n1832 VSS.n1831 2.6005
R7548 VSS.n1830 VSS.n1829 2.6005
R7549 VSS.n1829 VSS.n1828 2.6005
R7550 VSS.n1827 VSS.n1826 2.6005
R7551 VSS.n1826 VSS.n1825 2.6005
R7552 VSS.n1824 VSS.n1823 2.6005
R7553 VSS.n1823 VSS.n1822 2.6005
R7554 VSS.n1821 VSS.n1820 2.6005
R7555 VSS.n1820 VSS.n1819 2.6005
R7556 VSS.n1818 VSS.n1817 2.6005
R7557 VSS.n1817 VSS.n1816 2.6005
R7558 VSS.n1815 VSS.n1814 2.6005
R7559 VSS.n1814 VSS.n1813 2.6005
R7560 VSS.n1812 VSS.n1811 2.6005
R7561 VSS.n1811 VSS.n1810 2.6005
R7562 VSS.n1809 VSS.n1808 2.6005
R7563 VSS.n1808 VSS.n1807 2.6005
R7564 VSS.n1806 VSS.n1805 2.6005
R7565 VSS.n1805 VSS.n1804 2.6005
R7566 VSS.n1803 VSS.n1802 2.6005
R7567 VSS.n1802 VSS.n1801 2.6005
R7568 VSS.n1800 VSS.n1799 2.6005
R7569 VSS.n1799 VSS.n1798 2.6005
R7570 VSS.n1797 VSS.n1796 2.6005
R7571 VSS.n1796 VSS.n1795 2.6005
R7572 VSS.n1794 VSS.n1793 2.6005
R7573 VSS.n1793 VSS.n1792 2.6005
R7574 VSS.n1791 VSS.n1790 2.6005
R7575 VSS.n1790 VSS.n1789 2.6005
R7576 VSS.n1788 VSS.n1787 2.6005
R7577 VSS.n1787 VSS.n1786 2.6005
R7578 VSS.n1785 VSS.n1784 2.6005
R7579 VSS.n1784 VSS.n1783 2.6005
R7580 VSS.n1782 VSS.n1781 2.6005
R7581 VSS.n1781 VSS.n1780 2.6005
R7582 VSS.n1779 VSS.n1778 2.6005
R7583 VSS.n1778 VSS.n1777 2.6005
R7584 VSS.n1776 VSS.n1775 2.6005
R7585 VSS.n1775 VSS.n1774 2.6005
R7586 VSS.n1773 VSS.n1772 2.6005
R7587 VSS.n1772 VSS.n1771 2.6005
R7588 VSS.n1769 VSS.n1768 2.6005
R7589 VSS.n1768 VSS.n1767 2.6005
R7590 VSS.n5175 VSS.n5174 2.6005
R7591 VSS.n5174 VSS.n5173 2.6005
R7592 VSS.n5186 VSS.n5185 2.6005
R7593 VSS.n5185 VSS.n5184 2.6005
R7594 VSS.n5195 VSS.n5194 2.6005
R7595 VSS.n3287 VSS.n3286 2.6005
R7596 VSS.n3286 VSS.n3285 2.6005
R7597 VSS.n3290 VSS.n3289 2.6005
R7598 VSS.n3289 VSS.n3288 2.6005
R7599 VSS.n3293 VSS.n3292 2.6005
R7600 VSS.n3292 VSS.n3291 2.6005
R7601 VSS.n3296 VSS.n3295 2.6005
R7602 VSS.n3295 VSS.n3294 2.6005
R7603 VSS.n3299 VSS.n3298 2.6005
R7604 VSS.n3298 VSS.n3297 2.6005
R7605 VSS.n3302 VSS.n3301 2.6005
R7606 VSS.n3301 VSS.n3300 2.6005
R7607 VSS.n3305 VSS.n3304 2.6005
R7608 VSS.n3304 VSS.n3303 2.6005
R7609 VSS.n3308 VSS.n3307 2.6005
R7610 VSS.n3307 VSS.n3306 2.6005
R7611 VSS.n3311 VSS.n3310 2.6005
R7612 VSS.n3310 VSS.n3309 2.6005
R7613 VSS.n3314 VSS.n3313 2.6005
R7614 VSS.n3313 VSS.n3312 2.6005
R7615 VSS.n3317 VSS.n3316 2.6005
R7616 VSS.n3316 VSS.n3315 2.6005
R7617 VSS.n3320 VSS.n3319 2.6005
R7618 VSS.n3319 VSS.n3318 2.6005
R7619 VSS.n3323 VSS.n3322 2.6005
R7620 VSS.n3322 VSS.n3321 2.6005
R7621 VSS.n3326 VSS.n3325 2.6005
R7622 VSS.n3325 VSS.n3324 2.6005
R7623 VSS.n3329 VSS.n3328 2.6005
R7624 VSS.n3328 VSS.n3327 2.6005
R7625 VSS.n3332 VSS.n3331 2.6005
R7626 VSS.n3331 VSS.n3330 2.6005
R7627 VSS.n3335 VSS.n3334 2.6005
R7628 VSS.n3334 VSS.n3333 2.6005
R7629 VSS.n3338 VSS.n3337 2.6005
R7630 VSS.n3337 VSS.n3336 2.6005
R7631 VSS.n3341 VSS.n3340 2.6005
R7632 VSS.n3340 VSS.n3339 2.6005
R7633 VSS.n3344 VSS.n3343 2.6005
R7634 VSS.n3343 VSS.n3342 2.6005
R7635 VSS.n3347 VSS.n3346 2.6005
R7636 VSS.n3346 VSS.n3345 2.6005
R7637 VSS.n3350 VSS.n3349 2.6005
R7638 VSS.n3349 VSS.n3348 2.6005
R7639 VSS.n3353 VSS.n3352 2.6005
R7640 VSS.n3352 VSS.n3351 2.6005
R7641 VSS.n3356 VSS.n3355 2.6005
R7642 VSS.n3355 VSS.n3354 2.6005
R7643 VSS.n3359 VSS.n3358 2.6005
R7644 VSS.n3358 VSS.n3357 2.6005
R7645 VSS.n3362 VSS.n3361 2.6005
R7646 VSS.n3361 VSS.n3360 2.6005
R7647 VSS.n3365 VSS.n3364 2.6005
R7648 VSS.n3364 VSS.n3363 2.6005
R7649 VSS.n3368 VSS.n3367 2.6005
R7650 VSS.n3367 VSS.n3366 2.6005
R7651 VSS.n3371 VSS.n3370 2.6005
R7652 VSS.n3370 VSS.n3369 2.6005
R7653 VSS.n3375 VSS.n3374 2.6005
R7654 VSS.n3374 VSS.n3373 2.6005
R7655 VSS.n3378 VSS.n3377 2.6005
R7656 VSS.n3377 VSS.n3376 2.6005
R7657 VSS.n3381 VSS.n3380 2.6005
R7658 VSS.n3380 VSS.n3379 2.6005
R7659 VSS.n3384 VSS.n3383 2.6005
R7660 VSS.n3383 VSS.n3382 2.6005
R7661 VSS.n3387 VSS.n3386 2.6005
R7662 VSS.n3386 VSS.n3385 2.6005
R7663 VSS.n3390 VSS.n3389 2.6005
R7664 VSS.n3389 VSS.n3388 2.6005
R7665 VSS.n3393 VSS.n3392 2.6005
R7666 VSS.n3392 VSS.n3391 2.6005
R7667 VSS.n3396 VSS.n3395 2.6005
R7668 VSS.n3395 VSS.n3394 2.6005
R7669 VSS.n3399 VSS.n3398 2.6005
R7670 VSS.n3398 VSS.n3397 2.6005
R7671 VSS.n3402 VSS.n3401 2.6005
R7672 VSS.n3401 VSS.n3400 2.6005
R7673 VSS.n3405 VSS.n3404 2.6005
R7674 VSS.n3404 VSS.n3403 2.6005
R7675 VSS.n3408 VSS.n3407 2.6005
R7676 VSS.n3407 VSS.n3406 2.6005
R7677 VSS.n3411 VSS.n3410 2.6005
R7678 VSS.n3410 VSS.n3409 2.6005
R7679 VSS.n3414 VSS.n3413 2.6005
R7680 VSS.n3413 VSS.n3412 2.6005
R7681 VSS.n3417 VSS.n3416 2.6005
R7682 VSS.n3416 VSS.n3415 2.6005
R7683 VSS.n3420 VSS.n3419 2.6005
R7684 VSS.n3419 VSS.n3418 2.6005
R7685 VSS.n3423 VSS.n3422 2.6005
R7686 VSS.n3422 VSS.n3421 2.6005
R7687 VSS.n3426 VSS.n3425 2.6005
R7688 VSS.n3425 VSS.n3424 2.6005
R7689 VSS.n3429 VSS.n3428 2.6005
R7690 VSS.n3428 VSS.n3427 2.6005
R7691 VSS.n3432 VSS.n3431 2.6005
R7692 VSS.n3431 VSS.n3430 2.6005
R7693 VSS.n3435 VSS.n3434 2.6005
R7694 VSS.n3434 VSS.n3433 2.6005
R7695 VSS.n3438 VSS.n3437 2.6005
R7696 VSS.n3437 VSS.n3436 2.6005
R7697 VSS.n3441 VSS.n3440 2.6005
R7698 VSS.n3440 VSS.n3439 2.6005
R7699 VSS.n3444 VSS.n3443 2.6005
R7700 VSS.n3443 VSS.n3442 2.6005
R7701 VSS.n3447 VSS.n3446 2.6005
R7702 VSS.n3446 VSS.n3445 2.6005
R7703 VSS.n3457 VSS.n3456 2.6005
R7704 VSS.n3456 VSS.n3455 2.6005
R7705 VSS.n3460 VSS.n3459 2.6005
R7706 VSS.n3459 VSS.n3458 2.6005
R7707 VSS.n3463 VSS.n3462 2.6005
R7708 VSS.n3462 VSS.n3461 2.6005
R7709 VSS.n3466 VSS.n3465 2.6005
R7710 VSS.n3465 VSS.n3464 2.6005
R7711 VSS.n3469 VSS.n3468 2.6005
R7712 VSS.n3468 VSS.n3467 2.6005
R7713 VSS.n3472 VSS.n3471 2.6005
R7714 VSS.n3471 VSS.n3470 2.6005
R7715 VSS.n3475 VSS.n3474 2.6005
R7716 VSS.n3474 VSS.n3473 2.6005
R7717 VSS.n3478 VSS.n3477 2.6005
R7718 VSS.n3477 VSS.n3476 2.6005
R7719 VSS.n3481 VSS.n3480 2.6005
R7720 VSS.n3480 VSS.n3479 2.6005
R7721 VSS.n3484 VSS.n3483 2.6005
R7722 VSS.n3483 VSS.n3482 2.6005
R7723 VSS.n3493 VSS.n3492 2.6005
R7724 VSS.n3492 VSS.n3491 2.6005
R7725 VSS.n3502 VSS.n3501 2.6005
R7726 VSS.n3501 VSS.n3500 2.6005
R7727 VSS.n4002 VSS.n4001 2.6005
R7728 VSS.n4003 VSS.n4002 2.6005
R7729 VSS.n4000 VSS.n3999 2.6005
R7730 VSS.n3999 VSS.n3998 2.6005
R7731 VSS.n5283 VSS.n5282 2.6005
R7732 VSS.n433 VSS.n432 2.6005
R7733 VSS.n432 VSS.n431 2.6005
R7734 VSS.n436 VSS.n435 2.6005
R7735 VSS.n435 VSS.n434 2.6005
R7736 VSS.n439 VSS.n438 2.6005
R7737 VSS.n438 VSS.n437 2.6005
R7738 VSS.n442 VSS.n441 2.6005
R7739 VSS.n441 VSS.n440 2.6005
R7740 VSS.n445 VSS.n444 2.6005
R7741 VSS.n444 VSS.n443 2.6005
R7742 VSS.n448 VSS.n447 2.6005
R7743 VSS.n447 VSS.n446 2.6005
R7744 VSS.n451 VSS.n450 2.6005
R7745 VSS.n450 VSS.n449 2.6005
R7746 VSS.n454 VSS.n453 2.6005
R7747 VSS.n453 VSS.n452 2.6005
R7748 VSS.n457 VSS.n456 2.6005
R7749 VSS.n456 VSS.n455 2.6005
R7750 VSS.n460 VSS.n459 2.6005
R7751 VSS.n459 VSS.n458 2.6005
R7752 VSS.n463 VSS.n462 2.6005
R7753 VSS.n462 VSS.n461 2.6005
R7754 VSS.n466 VSS.n465 2.6005
R7755 VSS.n465 VSS.n464 2.6005
R7756 VSS.n469 VSS.n468 2.6005
R7757 VSS.n468 VSS.n467 2.6005
R7758 VSS.n472 VSS.n471 2.6005
R7759 VSS.n471 VSS.n470 2.6005
R7760 VSS.n475 VSS.n474 2.6005
R7761 VSS.n474 VSS.n473 2.6005
R7762 VSS.n478 VSS.n477 2.6005
R7763 VSS.n477 VSS.n476 2.6005
R7764 VSS.n481 VSS.n480 2.6005
R7765 VSS.n480 VSS.n479 2.6005
R7766 VSS.n484 VSS.n483 2.6005
R7767 VSS.n483 VSS.n482 2.6005
R7768 VSS.n487 VSS.n486 2.6005
R7769 VSS.n486 VSS.n485 2.6005
R7770 VSS.n490 VSS.n489 2.6005
R7771 VSS.n489 VSS.n488 2.6005
R7772 VSS.n493 VSS.n492 2.6005
R7773 VSS.n492 VSS.n491 2.6005
R7774 VSS.n496 VSS.n495 2.6005
R7775 VSS.n495 VSS.n494 2.6005
R7776 VSS.n499 VSS.n498 2.6005
R7777 VSS.n498 VSS.n497 2.6005
R7778 VSS.n502 VSS.n501 2.6005
R7779 VSS.n501 VSS.n500 2.6005
R7780 VSS.n505 VSS.n504 2.6005
R7781 VSS.n504 VSS.n503 2.6005
R7782 VSS.n508 VSS.n507 2.6005
R7783 VSS.n507 VSS.n506 2.6005
R7784 VSS.n511 VSS.n510 2.6005
R7785 VSS.n510 VSS.n509 2.6005
R7786 VSS.n514 VSS.n513 2.6005
R7787 VSS.n513 VSS.n512 2.6005
R7788 VSS.n517 VSS.n516 2.6005
R7789 VSS.n516 VSS.n515 2.6005
R7790 VSS.n520 VSS.n519 2.6005
R7791 VSS.n519 VSS.n518 2.6005
R7792 VSS.n4570 VSS.n4569 2.6005
R7793 VSS.n4569 VSS.n4568 2.6005
R7794 VSS.n4573 VSS.n4572 2.6005
R7795 VSS.n4572 VSS.n4571 2.6005
R7796 VSS.n4576 VSS.n4575 2.6005
R7797 VSS.n4575 VSS.n4574 2.6005
R7798 VSS.n4579 VSS.n4578 2.6005
R7799 VSS.n4578 VSS.n4577 2.6005
R7800 VSS.n4582 VSS.n4581 2.6005
R7801 VSS.n4581 VSS.n4580 2.6005
R7802 VSS.n4585 VSS.n4584 2.6005
R7803 VSS.n4584 VSS.n4583 2.6005
R7804 VSS.n4588 VSS.n4587 2.6005
R7805 VSS.n4587 VSS.n4586 2.6005
R7806 VSS.n4591 VSS.n4590 2.6005
R7807 VSS.n4590 VSS.n4589 2.6005
R7808 VSS.n4594 VSS.n4593 2.6005
R7809 VSS.n4593 VSS.n4592 2.6005
R7810 VSS.n4597 VSS.n4596 2.6005
R7811 VSS.n4596 VSS.n4595 2.6005
R7812 VSS.n4600 VSS.n4599 2.6005
R7813 VSS.n4599 VSS.n4598 2.6005
R7814 VSS.n4603 VSS.n4602 2.6005
R7815 VSS.n4602 VSS.n4601 2.6005
R7816 VSS.n4606 VSS.n4605 2.6005
R7817 VSS.n4605 VSS.n4604 2.6005
R7818 VSS.n4609 VSS.n4608 2.6005
R7819 VSS.n4608 VSS.n4607 2.6005
R7820 VSS.n4612 VSS.n4611 2.6005
R7821 VSS.n4611 VSS.n4610 2.6005
R7822 VSS.n4615 VSS.n4614 2.6005
R7823 VSS.n4614 VSS.n4613 2.6005
R7824 VSS.n4618 VSS.n4617 2.6005
R7825 VSS.n4617 VSS.n4616 2.6005
R7826 VSS.n4621 VSS.n4620 2.6005
R7827 VSS.n4620 VSS.n4619 2.6005
R7828 VSS.n4624 VSS.n4623 2.6005
R7829 VSS.n4623 VSS.n4622 2.6005
R7830 VSS.n4627 VSS.n4626 2.6005
R7831 VSS.n4626 VSS.n4625 2.6005
R7832 VSS.n4630 VSS.n4629 2.6005
R7833 VSS.n4629 VSS.n4628 2.6005
R7834 VSS.n4633 VSS.n4632 2.6005
R7835 VSS.n4632 VSS.n4631 2.6005
R7836 VSS.n4636 VSS.n4635 2.6005
R7837 VSS.n4635 VSS.n4634 2.6005
R7838 VSS.n4639 VSS.n4638 2.6005
R7839 VSS.n4638 VSS.n4637 2.6005
R7840 VSS.n4642 VSS.n4641 2.6005
R7841 VSS.n4641 VSS.n4640 2.6005
R7842 VSS.n4645 VSS.n4644 2.6005
R7843 VSS.n4644 VSS.n4643 2.6005
R7844 VSS.n4649 VSS.n4648 2.6005
R7845 VSS.n4648 VSS.n4647 2.6005
R7846 VSS.n4652 VSS.n4651 2.6005
R7847 VSS.n4651 VSS.n4650 2.6005
R7848 VSS.n4655 VSS.n4654 2.6005
R7849 VSS.n4654 VSS.n4653 2.6005
R7850 VSS.n4658 VSS.n4657 2.6005
R7851 VSS.n4657 VSS.n4656 2.6005
R7852 VSS.n4661 VSS.n4660 2.6005
R7853 VSS.n4660 VSS.n4659 2.6005
R7854 VSS.n4664 VSS.n4663 2.6005
R7855 VSS.n4663 VSS.n4662 2.6005
R7856 VSS.n4667 VSS.n4666 2.6005
R7857 VSS.n4666 VSS.n4665 2.6005
R7858 VSS.n4670 VSS.n4669 2.6005
R7859 VSS.n4669 VSS.n4668 2.6005
R7860 VSS.n4673 VSS.n4672 2.6005
R7861 VSS.n4672 VSS.n4671 2.6005
R7862 VSS.n4676 VSS.n4675 2.6005
R7863 VSS.n4675 VSS.n4674 2.6005
R7864 VSS.n4679 VSS.n4678 2.6005
R7865 VSS.n4678 VSS.n4677 2.6005
R7866 VSS.n4681 VSS.n4680 2.6005
R7867 VSS.n4683 VSS.n4682 2.6005
R7868 VSS.n4685 VSS.n4684 2.6005
R7869 VSS.n4687 VSS.n4686 2.6005
R7870 VSS.n4689 VSS.n4688 2.6005
R7871 VSS.n4691 VSS.n4690 2.6005
R7872 VSS.n4693 VSS.n4692 2.6005
R7873 VSS.n4695 VSS.n4694 2.6005
R7874 VSS.n4697 VSS.n4696 2.6005
R7875 VSS.n4699 VSS.n4698 2.6005
R7876 VSS.n4701 VSS.n4700 2.6005
R7877 VSS.n4703 VSS.n4702 2.6005
R7878 VSS.n4705 VSS.n4704 2.6005
R7879 VSS.n4707 VSS.n4706 2.6005
R7880 VSS.n4709 VSS.n4708 2.6005
R7881 VSS.n4711 VSS.n4710 2.6005
R7882 VSS.n4713 VSS.n4712 2.6005
R7883 VSS.n4715 VSS.n4714 2.6005
R7884 VSS.n4717 VSS.n4716 2.6005
R7885 VSS.n4720 VSS.n4719 2.6005
R7886 VSS.n4722 VSS.n4721 2.6005
R7887 VSS.n4725 VSS.n4724 2.6005
R7888 VSS.n4727 VSS.n4726 2.6005
R7889 VSS.n4730 VSS.n4729 2.6005
R7890 VSS.n4732 VSS.n4731 2.6005
R7891 VSS.n4735 VSS.n4734 2.6005
R7892 VSS.n4737 VSS.n4736 2.6005
R7893 VSS.n4740 VSS.n4739 2.6005
R7894 VSS.n4742 VSS.n4741 2.6005
R7895 VSS.n4745 VSS.n4744 2.6005
R7896 VSS.n4747 VSS.n4746 2.6005
R7897 VSS.n4942 VSS.n4941 2.6005
R7898 VSS.n4940 VSS.n4939 2.6005
R7899 VSS.n4939 VSS.n4938 2.6005
R7900 VSS.n4937 VSS.n4936 2.6005
R7901 VSS.n4936 VSS.n4935 2.6005
R7902 VSS.n4934 VSS.n4933 2.6005
R7903 VSS.n4933 VSS.n4932 2.6005
R7904 VSS.n4931 VSS.n4930 2.6005
R7905 VSS.n4930 VSS.n4929 2.6005
R7906 VSS.n4928 VSS.n4927 2.6005
R7907 VSS.n4927 VSS.n4926 2.6005
R7908 VSS.n4925 VSS.n4924 2.6005
R7909 VSS.n4924 VSS.n4923 2.6005
R7910 VSS.n4922 VSS.n4921 2.6005
R7911 VSS.n4921 VSS.n4920 2.6005
R7912 VSS.n4919 VSS.n4918 2.6005
R7913 VSS.n4918 VSS.n4917 2.6005
R7914 VSS.n4916 VSS.n4915 2.6005
R7915 VSS.n4915 VSS.n4914 2.6005
R7916 VSS.n4913 VSS.n4912 2.6005
R7917 VSS.n4911 VSS.n4910 2.6005
R7918 VSS.n4908 VSS.n4907 2.6005
R7919 VSS.n4906 VSS.n4905 2.6005
R7920 VSS.n4903 VSS.n4902 2.6005
R7921 VSS.n4901 VSS.n4900 2.6005
R7922 VSS.n4898 VSS.n4897 2.6005
R7923 VSS.n4896 VSS.n4895 2.6005
R7924 VSS.n4893 VSS.n4892 2.6005
R7925 VSS.n4891 VSS.n4890 2.6005
R7926 VSS.n4887 VSS.n4886 2.6005
R7927 VSS.n4886 VSS.n4885 2.6005
R7928 VSS.n4882 VSS.n4881 2.6005
R7929 VSS.n4881 VSS.n4880 2.6005
R7930 VSS.n4879 VSS.n4878 2.6005
R7931 VSS.n4878 VSS.n4877 2.6005
R7932 VSS.n4876 VSS.n4875 2.6005
R7933 VSS.n4875 VSS.n4874 2.6005
R7934 VSS.n4873 VSS.n4872 2.6005
R7935 VSS.n4872 VSS.n4871 2.6005
R7936 VSS.n4870 VSS.n4869 2.6005
R7937 VSS.n4869 VSS.n4868 2.6005
R7938 VSS.n4866 VSS.n4865 2.6005
R7939 VSS.n4864 VSS.n4863 2.6005
R7940 VSS.n4862 VSS.n4861 2.6005
R7941 VSS.n4859 VSS.n4858 2.6005
R7942 VSS.n4857 VSS.n4856 2.6005
R7943 VSS.n4855 VSS.n4854 2.6005
R7944 VSS.n4853 VSS.n4852 2.6005
R7945 VSS.n4851 VSS.n4850 2.6005
R7946 VSS.n4849 VSS.n4848 2.6005
R7947 VSS.n4846 VSS.n4845 2.6005
R7948 VSS.n4844 VSS.n4843 2.6005
R7949 VSS.n4841 VSS.n4840 2.6005
R7950 VSS.n4839 VSS.n4838 2.6005
R7951 VSS.n4836 VSS.n4835 2.6005
R7952 VSS.n4834 VSS.n4833 2.6005
R7953 VSS.n4831 VSS.n4830 2.6005
R7954 VSS.n4829 VSS.n4828 2.6005
R7955 VSS.n4826 VSS.n4825 2.6005
R7956 VSS.n4824 VSS.n4823 2.6005
R7957 VSS.n4821 VSS.n4820 2.6005
R7958 VSS.n4819 VSS.n4818 2.6005
R7959 VSS.n4812 VSS.n4811 2.6005
R7960 VSS.n4810 VSS.n4809 2.6005
R7961 VSS.n4807 VSS.n4806 2.6005
R7962 VSS.n4805 VSS.n4804 2.6005
R7963 VSS.n4801 VSS.n4800 2.6005
R7964 VSS.n4800 VSS.n4799 2.6005
R7965 VSS.n4797 VSS.n4796 2.6005
R7966 VSS.n4796 VSS.n4795 2.6005
R7967 VSS.n4794 VSS.n4793 2.6005
R7968 VSS.n4793 VSS.n4792 2.6005
R7969 VSS.n4791 VSS.n4790 2.6005
R7970 VSS.n4790 VSS.n4789 2.6005
R7971 VSS.n4788 VSS.n4787 2.6005
R7972 VSS.n4787 VSS.n4786 2.6005
R7973 VSS.n4785 VSS.n4784 2.6005
R7974 VSS.n4784 VSS.n4783 2.6005
R7975 VSS.n4782 VSS.n4781 2.6005
R7976 VSS.n4780 VSS.n4779 2.6005
R7977 VSS.n4777 VSS.n4776 2.6005
R7978 VSS.n4775 VSS.n4774 2.6005
R7979 VSS.n4772 VSS.n4771 2.6005
R7980 VSS.n4770 VSS.n4769 2.6005
R7981 VSS.n4767 VSS.n4766 2.6005
R7982 VSS.n4765 VSS.n4764 2.6005
R7983 VSS.n4761 VSS.n4760 2.6005
R7984 VSS.n4760 VSS.n4759 2.6005
R7985 VSS.n4756 VSS.n4755 2.6005
R7986 VSS.n4755 VSS.n4754 2.6005
R7987 VSS.n4753 VSS.n4752 2.6005
R7988 VSS.n4752 VSS.n4751 2.6005
R7989 VSS.n4750 VSS.n4749 2.6005
R7990 VSS.n4749 VSS.n4748 2.6005
R7991 VSS.n218 VSS.n217 2.6005
R7992 VSS.n217 VSS.n216 2.6005
R7993 VSS.n5379 VSS.n5378 2.6005
R7994 VSS.n5380 VSS.n5379 2.6005
R7995 VSS.n5377 VSS.n5376 2.6005
R7996 VSS.n5375 VSS.n5374 2.6005
R7997 VSS.n5373 VSS.n5372 2.6005
R7998 VSS.n5370 VSS.n5369 2.6005
R7999 VSS.n5368 VSS.n5367 2.6005
R8000 VSS.n5366 VSS.n5365 2.6005
R8001 VSS.n5364 VSS.n5363 2.6005
R8002 VSS.n5362 VSS.n5361 2.6005
R8003 VSS.n5360 VSS.n5359 2.6005
R8004 VSS.n5357 VSS.n5356 2.6005
R8005 VSS.n5355 VSS.n5354 2.6005
R8006 VSS.n5352 VSS.n5351 2.6005
R8007 VSS.n5350 VSS.n5349 2.6005
R8008 VSS.n5347 VSS.n5346 2.6005
R8009 VSS.n5345 VSS.n5344 2.6005
R8010 VSS.n5342 VSS.n5341 2.6005
R8011 VSS.n5340 VSS.n5339 2.6005
R8012 VSS.n5337 VSS.n5336 2.6005
R8013 VSS.n5335 VSS.n5334 2.6005
R8014 VSS.n5332 VSS.n5331 2.6005
R8015 VSS.n5330 VSS.n5329 2.6005
R8016 VSS.n5323 VSS.n5322 2.6005
R8017 VSS.n5321 VSS.n5320 2.6005
R8018 VSS.n5318 VSS.n5317 2.6005
R8019 VSS.n5316 VSS.n5315 2.6005
R8020 VSS.n5312 VSS.n5311 2.6005
R8021 VSS.n5311 VSS.n5310 2.6005
R8022 VSS.n5308 VSS.n5307 2.6005
R8023 VSS.n5307 VSS.n5306 2.6005
R8024 VSS.n5305 VSS.n5304 2.6005
R8025 VSS.n5304 VSS.n5303 2.6005
R8026 VSS.n5302 VSS.n5301 2.6005
R8027 VSS.n5301 VSS.n5300 2.6005
R8028 VSS.n5299 VSS.n5298 2.6005
R8029 VSS.n5298 VSS.n5297 2.6005
R8030 VSS.n5296 VSS.n5295 2.6005
R8031 VSS.n5295 VSS.n5294 2.6005
R8032 VSS.n5293 VSS.n5292 2.6005
R8033 VSS.n5291 VSS.n5290 2.6005
R8034 VSS.n5288 VSS.n5287 2.6005
R8035 VSS.n5286 VSS.n5285 2.6005
R8036 VSS.n430 VSS.n429 2.6005
R8037 VSS.n429 VSS.n428 2.6005
R8038 VSS.n5281 VSS.n5280 2.6005
R8039 VSS.n427 VSS.n426 2.6005
R8040 VSS.n426 VSS.n425 2.6005
R8041 VSS.n3844 VSS.n3843 2.6005
R8042 VSS.n3846 VSS.n3845 2.6005
R8043 VSS.n3848 VSS.n3847 2.6005
R8044 VSS.n3850 VSS.n3849 2.6005
R8045 VSS.n3852 VSS.n3851 2.6005
R8046 VSS.n3854 VSS.n3853 2.6005
R8047 VSS.n3856 VSS.n3855 2.6005
R8048 VSS.n3858 VSS.n3857 2.6005
R8049 VSS.n3860 VSS.n3859 2.6005
R8050 VSS.n3862 VSS.n3861 2.6005
R8051 VSS.n3864 VSS.n3863 2.6005
R8052 VSS.n3866 VSS.n3865 2.6005
R8053 VSS.n3868 VSS.n3867 2.6005
R8054 VSS.n3870 VSS.n3869 2.6005
R8055 VSS.n3872 VSS.n3871 2.6005
R8056 VSS.n3874 VSS.n3873 2.6005
R8057 VSS.n3876 VSS.n3875 2.6005
R8058 VSS.n3878 VSS.n3877 2.6005
R8059 VSS.n3880 VSS.n3879 2.6005
R8060 VSS.n3882 VSS.n3881 2.6005
R8061 VSS.n3884 VSS.n3883 2.6005
R8062 VSS.n3886 VSS.n3885 2.6005
R8063 VSS.n3888 VSS.n3887 2.6005
R8064 VSS.n3890 VSS.n3889 2.6005
R8065 VSS.n3892 VSS.n3891 2.6005
R8066 VSS.n3894 VSS.n3893 2.6005
R8067 VSS.n3897 VSS.n3896 2.6005
R8068 VSS.n3899 VSS.n3898 2.6005
R8069 VSS.n3902 VSS.n3901 2.6005
R8070 VSS.n3904 VSS.n3903 2.6005
R8071 VSS.n3907 VSS.n3906 2.6005
R8072 VSS.n3909 VSS.n3908 2.6005
R8073 VSS.n3912 VSS.n3911 2.6005
R8074 VSS.n3916 VSS.n3915 2.6005
R8075 VSS.n3972 VSS.n3971 2.6005
R8076 VSS.n3976 VSS.n3975 2.6005
R8077 VSS.n1160 VSS.n1159 2.6005
R8078 VSS.n1159 VSS.n1158 2.6005
R8079 VSS.n1163 VSS.n1162 2.6005
R8080 VSS.n1162 VSS.n1161 2.6005
R8081 VSS.n1166 VSS.n1165 2.6005
R8082 VSS.n1165 VSS.n1164 2.6005
R8083 VSS.n1169 VSS.n1168 2.6005
R8084 VSS.n1168 VSS.n1167 2.6005
R8085 VSS.n1172 VSS.n1171 2.6005
R8086 VSS.n1171 VSS.n1170 2.6005
R8087 VSS.n1175 VSS.n1174 2.6005
R8088 VSS.n1174 VSS.n1173 2.6005
R8089 VSS.n1178 VSS.n1177 2.6005
R8090 VSS.n1177 VSS.n1176 2.6005
R8091 VSS.n1181 VSS.n1180 2.6005
R8092 VSS.n1180 VSS.n1179 2.6005
R8093 VSS.n1184 VSS.n1183 2.6005
R8094 VSS.n1183 VSS.n1182 2.6005
R8095 VSS.n1187 VSS.n1186 2.6005
R8096 VSS.n1186 VSS.n1185 2.6005
R8097 VSS.n1190 VSS.n1189 2.6005
R8098 VSS.n1189 VSS.n1188 2.6005
R8099 VSS.n1193 VSS.n1192 2.6005
R8100 VSS.n1192 VSS.n1191 2.6005
R8101 VSS.n1196 VSS.n1195 2.6005
R8102 VSS.n1195 VSS.n1194 2.6005
R8103 VSS.n1199 VSS.n1198 2.6005
R8104 VSS.n1198 VSS.n1197 2.6005
R8105 VSS.n1202 VSS.n1201 2.6005
R8106 VSS.n1201 VSS.n1200 2.6005
R8107 VSS.n1205 VSS.n1204 2.6005
R8108 VSS.n1204 VSS.n1203 2.6005
R8109 VSS.n1208 VSS.n1207 2.6005
R8110 VSS.n1207 VSS.n1206 2.6005
R8111 VSS.n1211 VSS.n1210 2.6005
R8112 VSS.n1210 VSS.n1209 2.6005
R8113 VSS.n1214 VSS.n1213 2.6005
R8114 VSS.n1213 VSS.n1212 2.6005
R8115 VSS.n1217 VSS.n1216 2.6005
R8116 VSS.n1216 VSS.n1215 2.6005
R8117 VSS.n1220 VSS.n1219 2.6005
R8118 VSS.n1219 VSS.n1218 2.6005
R8119 VSS.n1223 VSS.n1222 2.6005
R8120 VSS.n1222 VSS.n1221 2.6005
R8121 VSS.n1226 VSS.n1225 2.6005
R8122 VSS.n1225 VSS.n1224 2.6005
R8123 VSS.n1229 VSS.n1228 2.6005
R8124 VSS.n1228 VSS.n1227 2.6005
R8125 VSS.n1232 VSS.n1231 2.6005
R8126 VSS.n1231 VSS.n1230 2.6005
R8127 VSS.n1235 VSS.n1234 2.6005
R8128 VSS.n1234 VSS.n1233 2.6005
R8129 VSS.n1238 VSS.n1237 2.6005
R8130 VSS.n1237 VSS.n1236 2.6005
R8131 VSS.n1241 VSS.n1240 2.6005
R8132 VSS.n1240 VSS.n1239 2.6005
R8133 VSS.n1244 VSS.n1243 2.6005
R8134 VSS.n1243 VSS.n1242 2.6005
R8135 VSS.n1247 VSS.n1246 2.6005
R8136 VSS.n1246 VSS.n1245 2.6005
R8137 VSS.n1250 VSS.n1249 2.6005
R8138 VSS.n1249 VSS.n1248 2.6005
R8139 VSS.n1253 VSS.n1252 2.6005
R8140 VSS.n1252 VSS.n1251 2.6005
R8141 VSS.n1256 VSS.n1255 2.6005
R8142 VSS.n1255 VSS.n1254 2.6005
R8143 VSS.n1259 VSS.n1258 2.6005
R8144 VSS.n1258 VSS.n1257 2.6005
R8145 VSS.n1262 VSS.n1261 2.6005
R8146 VSS.n1261 VSS.n1260 2.6005
R8147 VSS.n1265 VSS.n1264 2.6005
R8148 VSS.n1264 VSS.n1263 2.6005
R8149 VSS.n1268 VSS.n1267 2.6005
R8150 VSS.n1267 VSS.n1266 2.6005
R8151 VSS.n1271 VSS.n1270 2.6005
R8152 VSS.n1270 VSS.n1269 2.6005
R8153 VSS.n1274 VSS.n1273 2.6005
R8154 VSS.n1273 VSS.n1272 2.6005
R8155 VSS.n1277 VSS.n1276 2.6005
R8156 VSS.n1276 VSS.n1275 2.6005
R8157 VSS.n1280 VSS.n1279 2.6005
R8158 VSS.n1279 VSS.n1278 2.6005
R8159 VSS.n1283 VSS.n1282 2.6005
R8160 VSS.n1282 VSS.n1281 2.6005
R8161 VSS.n1286 VSS.n1285 2.6005
R8162 VSS.n1285 VSS.n1284 2.6005
R8163 VSS.n1289 VSS.n1288 2.6005
R8164 VSS.n1288 VSS.n1287 2.6005
R8165 VSS.n1292 VSS.n1291 2.6005
R8166 VSS.n1291 VSS.n1290 2.6005
R8167 VSS.n1295 VSS.n1294 2.6005
R8168 VSS.n1294 VSS.n1293 2.6005
R8169 VSS.n1298 VSS.n1297 2.6005
R8170 VSS.n1297 VSS.n1296 2.6005
R8171 VSS.n1336 VSS.n1335 2.6005
R8172 VSS.n1335 VSS.n1334 2.6005
R8173 VSS.n1338 VSS.n1337 2.6005
R8174 VSS.n1341 VSS.n1340 2.6005
R8175 VSS.n1343 VSS.n1342 2.6005
R8176 VSS.n1346 VSS.n1345 2.6005
R8177 VSS.n1348 VSS.n1347 2.6005
R8178 VSS.n1351 VSS.n1350 2.6005
R8179 VSS.n1355 VSS.n1354 2.6005
R8180 VSS.n1359 VSS.n1358 2.6005
R8181 VSS.n1362 VSS.n1361 2.6005
R8182 VSS.n1682 VSS.n1681 2.6005
R8183 VSS.n1366 VSS.n1365 2.6005
R8184 VSS.n1368 VSS.n1367 2.6005
R8185 VSS.n1371 VSS.n1370 2.6005
R8186 VSS.n1373 VSS.n1372 2.6005
R8187 VSS.n1376 VSS.n1375 2.6005
R8188 VSS.n1378 VSS.n1377 2.6005
R8189 VSS.n1381 VSS.n1380 2.6005
R8190 VSS.n1383 VSS.n1382 2.6005
R8191 VSS.n1386 VSS.n1385 2.6005
R8192 VSS.n1677 VSS.n1676 2.6005
R8193 VSS.n1675 VSS.n1674 2.6005
R8194 VSS.n1674 VSS.n1673 2.6005
R8195 VSS.n1672 VSS.n1671 2.6005
R8196 VSS.n1671 VSS.n1670 2.6005
R8197 VSS.n1669 VSS.n1668 2.6005
R8198 VSS.n1668 VSS.n1667 2.6005
R8199 VSS.n1666 VSS.n1665 2.6005
R8200 VSS.n1665 VSS.n1664 2.6005
R8201 VSS.n1663 VSS.n1662 2.6005
R8202 VSS.n1662 VSS.n1661 2.6005
R8203 VSS.n1660 VSS.n1659 2.6005
R8204 VSS.n1659 VSS.n1658 2.6005
R8205 VSS.n1657 VSS.n1656 2.6005
R8206 VSS.n1656 VSS.n1655 2.6005
R8207 VSS.n1654 VSS.n1653 2.6005
R8208 VSS.n1653 VSS.n1652 2.6005
R8209 VSS.n1651 VSS.n1650 2.6005
R8210 VSS.n1650 VSS.n1649 2.6005
R8211 VSS.n1648 VSS.n1647 2.6005
R8212 VSS.n1641 VSS.n1640 2.6005
R8213 VSS.n1639 VSS.n1638 2.6005
R8214 VSS.n1636 VSS.n1635 2.6005
R8215 VSS.n1634 VSS.n1633 2.6005
R8216 VSS.n1631 VSS.n1630 2.6005
R8217 VSS.n1629 VSS.n1628 2.6005
R8218 VSS.n1626 VSS.n1625 2.6005
R8219 VSS.n1624 VSS.n1623 2.6005
R8220 VSS.n1622 VSS.n1621 2.6005
R8221 VSS.n1620 VSS.n1619 2.6005
R8222 VSS.n1619 VSS.n1618 2.6005
R8223 VSS.n1616 VSS.n1615 2.6005
R8224 VSS.n1615 VSS.n1614 2.6005
R8225 VSS.n1612 VSS.n1611 2.6005
R8226 VSS.n1611 VSS.n1610 2.6005
R8227 VSS.n1609 VSS.n1608 2.6005
R8228 VSS.n1608 VSS.n1607 2.6005
R8229 VSS.n1606 VSS.n1605 2.6005
R8230 VSS.n1605 VSS.n1604 2.6005
R8231 VSS.n1603 VSS.n1602 2.6005
R8232 VSS.n1602 VSS.n1601 2.6005
R8233 VSS.n1600 VSS.n1599 2.6005
R8234 VSS.n1599 VSS.n1598 2.6005
R8235 VSS.n1597 VSS.n1596 2.6005
R8236 VSS.n1596 VSS.n1595 2.6005
R8237 VSS.n1594 VSS.n1593 2.6005
R8238 VSS.n1593 VSS.n1592 2.6005
R8239 VSS.n1591 VSS.n1590 2.6005
R8240 VSS.n1590 VSS.n1589 2.6005
R8241 VSS.n1588 VSS.n1587 2.6005
R8242 VSS.n1587 VSS.n1586 2.6005
R8243 VSS.n1585 VSS.n1584 2.6005
R8244 VSS.n1584 VSS.n1583 2.6005
R8245 VSS.n1582 VSS.n1581 2.6005
R8246 VSS.n1581 VSS.n1580 2.6005
R8247 VSS.n1579 VSS.n1578 2.6005
R8248 VSS.n1578 VSS.n1577 2.6005
R8249 VSS.n1576 VSS.n1575 2.6005
R8250 VSS.n1575 VSS.n1574 2.6005
R8251 VSS.n1573 VSS.n1572 2.6005
R8252 VSS.n1572 VSS.n1571 2.6005
R8253 VSS.n1570 VSS.n1569 2.6005
R8254 VSS.n1569 VSS.n1568 2.6005
R8255 VSS.n1567 VSS.n1566 2.6005
R8256 VSS.n1566 VSS.n1565 2.6005
R8257 VSS.n1564 VSS.n1563 2.6005
R8258 VSS.n1563 VSS.n1562 2.6005
R8259 VSS.n1561 VSS.n1560 2.6005
R8260 VSS.n1560 VSS.n1559 2.6005
R8261 VSS.n1558 VSS.n1557 2.6005
R8262 VSS.n1557 VSS.n1556 2.6005
R8263 VSS.n1555 VSS.n1554 2.6005
R8264 VSS.n1554 VSS.n1553 2.6005
R8265 VSS.n1552 VSS.n1551 2.6005
R8266 VSS.n1551 VSS.n1550 2.6005
R8267 VSS.n1549 VSS.n1548 2.6005
R8268 VSS.n1548 VSS.n1547 2.6005
R8269 VSS.n1546 VSS.n1545 2.6005
R8270 VSS.n1545 VSS.n1544 2.6005
R8271 VSS.n1543 VSS.n1542 2.6005
R8272 VSS.n1542 VSS.n1541 2.6005
R8273 VSS.n1540 VSS.n1539 2.6005
R8274 VSS.n1539 VSS.n1538 2.6005
R8275 VSS.n1533 VSS.n1532 2.6005
R8276 VSS.n1532 VSS.n1531 2.6005
R8277 VSS.n1526 VSS.n1525 2.6005
R8278 VSS.n1525 VSS.n1524 2.6005
R8279 VSS.n1519 VSS.n1518 2.6005
R8280 VSS.n1518 VSS.n1517 2.6005
R8281 VSS.n1513 VSS.n1512 2.6005
R8282 VSS.n1512 VSS.n1511 2.6005
R8283 VSS.n1510 VSS.n1509 2.6005
R8284 VSS.n1507 VSS.n1506 2.6005
R8285 VSS.n1506 VSS.n1505 2.6005
R8286 VSS.n1504 VSS.n1503 2.6005
R8287 VSS.n1503 VSS.n1502 2.6005
R8288 VSS.n1501 VSS.n1500 2.6005
R8289 VSS.n1500 VSS.n1499 2.6005
R8290 VSS.n1498 VSS.n1497 2.6005
R8291 VSS.n1497 VSS.n1496 2.6005
R8292 VSS.n1495 VSS.n1494 2.6005
R8293 VSS.n1494 VSS.n1493 2.6005
R8294 VSS.n1492 VSS.n1491 2.6005
R8295 VSS.n1491 VSS.n1490 2.6005
R8296 VSS.n1489 VSS.n1488 2.6005
R8297 VSS.n1488 VSS.n1487 2.6005
R8298 VSS.n1486 VSS.n1485 2.6005
R8299 VSS.n1485 VSS.n1484 2.6005
R8300 VSS.n1483 VSS.n1482 2.6005
R8301 VSS.n1482 VSS.n1481 2.6005
R8302 VSS.n1480 VSS.n1479 2.6005
R8303 VSS.n1479 VSS.n1478 2.6005
R8304 VSS.n1477 VSS.n1476 2.6005
R8305 VSS.n1476 VSS.n1475 2.6005
R8306 VSS.n1474 VSS.n1473 2.6005
R8307 VSS.n1473 VSS.n1472 2.6005
R8308 VSS.n1471 VSS.n1470 2.6005
R8309 VSS.n1470 VSS.n1469 2.6005
R8310 VSS.n1468 VSS.n1467 2.6005
R8311 VSS.n1467 VSS.n1466 2.6005
R8312 VSS.n1465 VSS.n1464 2.6005
R8313 VSS.n1464 VSS.n1463 2.6005
R8314 VSS.n1462 VSS.n1461 2.6005
R8315 VSS.n1461 VSS.n1460 2.6005
R8316 VSS.n1459 VSS.n1458 2.6005
R8317 VSS.n1458 VSS.n1457 2.6005
R8318 VSS.n1456 VSS.n1455 2.6005
R8319 VSS.n1455 VSS.n1454 2.6005
R8320 VSS.n1453 VSS.n1452 2.6005
R8321 VSS.n1452 VSS.n1451 2.6005
R8322 VSS.n1450 VSS.n1449 2.6005
R8323 VSS.n1449 VSS.n1448 2.6005
R8324 VSS.n1447 VSS.n1446 2.6005
R8325 VSS.n1446 VSS.n1445 2.6005
R8326 VSS.n1444 VSS.n1443 2.6005
R8327 VSS.n1443 VSS.n1442 2.6005
R8328 VSS.n1441 VSS.n1440 2.6005
R8329 VSS.n1440 VSS.n1439 2.6005
R8330 VSS.n1438 VSS.n1437 2.6005
R8331 VSS.n1437 VSS.n1436 2.6005
R8332 VSS.n1435 VSS.n1434 2.6005
R8333 VSS.n1434 VSS.n1433 2.6005
R8334 VSS.n1432 VSS.n1431 2.6005
R8335 VSS.n1431 VSS.n1430 2.6005
R8336 VSS.n1429 VSS.n1428 2.6005
R8337 VSS.n1428 VSS.n1427 2.6005
R8338 VSS.n1426 VSS.n1425 2.6005
R8339 VSS.n1425 VSS.n1424 2.6005
R8340 VSS.n1423 VSS.n1422 2.6005
R8341 VSS.n1422 VSS.n1421 2.6005
R8342 VSS.n1420 VSS.n1419 2.6005
R8343 VSS.n1419 VSS.n1418 2.6005
R8344 VSS.n1417 VSS.n1416 2.6005
R8345 VSS.n1416 VSS.n1415 2.6005
R8346 VSS.n1414 VSS.n1413 2.6005
R8347 VSS.n1413 VSS.n1412 2.6005
R8348 VSS.n1411 VSS.n1410 2.6005
R8349 VSS.n1410 VSS.n1409 2.6005
R8350 VSS.n1408 VSS.n1407 2.6005
R8351 VSS.n1407 VSS.n1406 2.6005
R8352 VSS.n1405 VSS.n1404 2.6005
R8353 VSS.n1404 VSS.n1403 2.6005
R8354 VSS.n1402 VSS.n1401 2.6005
R8355 VSS.n1401 VSS.n1400 2.6005
R8356 VSS.n1399 VSS.n1398 2.6005
R8357 VSS.n1398 VSS.n1397 2.6005
R8358 VSS.n1396 VSS.n1395 2.6005
R8359 VSS.n1395 VSS.n1394 2.6005
R8360 VSS.n1393 VSS.n1392 2.6005
R8361 VSS.n1392 VSS.n1391 2.6005
R8362 VSS.n1390 VSS.n1389 2.6005
R8363 VSS.n1389 VSS.n1388 2.6005
R8364 VSS.n789 VSS.n788 2.6005
R8365 VSS.n788 VSS.n787 2.6005
R8366 VSS.n792 VSS.n791 2.6005
R8367 VSS.n791 VSS.n790 2.6005
R8368 VSS.n795 VSS.n794 2.6005
R8369 VSS.n794 VSS.n793 2.6005
R8370 VSS.n798 VSS.n797 2.6005
R8371 VSS.n797 VSS.n796 2.6005
R8372 VSS.n801 VSS.n800 2.6005
R8373 VSS.n800 VSS.n799 2.6005
R8374 VSS.n804 VSS.n803 2.6005
R8375 VSS.n803 VSS.n802 2.6005
R8376 VSS.n807 VSS.n806 2.6005
R8377 VSS.n806 VSS.n805 2.6005
R8378 VSS.n810 VSS.n809 2.6005
R8379 VSS.n809 VSS.n808 2.6005
R8380 VSS.n813 VSS.n812 2.6005
R8381 VSS.n812 VSS.n811 2.6005
R8382 VSS.n816 VSS.n815 2.6005
R8383 VSS.n815 VSS.n814 2.6005
R8384 VSS.n819 VSS.n818 2.6005
R8385 VSS.n818 VSS.n817 2.6005
R8386 VSS.n822 VSS.n821 2.6005
R8387 VSS.n821 VSS.n820 2.6005
R8388 VSS.n825 VSS.n824 2.6005
R8389 VSS.n824 VSS.n823 2.6005
R8390 VSS.n828 VSS.n827 2.6005
R8391 VSS.n827 VSS.n826 2.6005
R8392 VSS.n831 VSS.n830 2.6005
R8393 VSS.n830 VSS.n829 2.6005
R8394 VSS.n834 VSS.n833 2.6005
R8395 VSS.n833 VSS.n832 2.6005
R8396 VSS.n837 VSS.n836 2.6005
R8397 VSS.n836 VSS.n835 2.6005
R8398 VSS.n840 VSS.n839 2.6005
R8399 VSS.n839 VSS.n838 2.6005
R8400 VSS.n843 VSS.n842 2.6005
R8401 VSS.n842 VSS.n841 2.6005
R8402 VSS.n846 VSS.n845 2.6005
R8403 VSS.n845 VSS.n844 2.6005
R8404 VSS.n849 VSS.n848 2.6005
R8405 VSS.n848 VSS.n847 2.6005
R8406 VSS.n852 VSS.n851 2.6005
R8407 VSS.n851 VSS.n850 2.6005
R8408 VSS.n856 VSS.n855 2.6005
R8409 VSS.n855 VSS.n854 2.6005
R8410 VSS.n869 VSS.n868 2.6005
R8411 VSS.n868 VSS.n867 2.6005
R8412 VSS.n876 VSS.n875 2.6005
R8413 VSS.n875 VSS.n874 2.6005
R8414 VSS.n890 VSS.n889 2.6005
R8415 VSS.n889 VSS.n888 2.6005
R8416 VSS.n887 VSS.n886 2.6005
R8417 VSS.n981 VSS.n980 2.6005
R8418 VSS.n980 VSS.n979 2.6005
R8419 VSS.n978 VSS.n977 2.6005
R8420 VSS.n977 VSS.n976 2.6005
R8421 VSS.n975 VSS.n974 2.6005
R8422 VSS.n974 VSS.n973 2.6005
R8423 VSS.n972 VSS.n971 2.6005
R8424 VSS.n971 VSS.n970 2.6005
R8425 VSS.n969 VSS.n968 2.6005
R8426 VSS.n968 VSS.n967 2.6005
R8427 VSS.n966 VSS.n965 2.6005
R8428 VSS.n965 VSS.n964 2.6005
R8429 VSS.n963 VSS.n962 2.6005
R8430 VSS.n962 VSS.n961 2.6005
R8431 VSS.n960 VSS.n959 2.6005
R8432 VSS.n959 VSS.n958 2.6005
R8433 VSS.n957 VSS.n956 2.6005
R8434 VSS.n956 VSS.n955 2.6005
R8435 VSS.n954 VSS.n953 2.6005
R8436 VSS.n953 VSS.n952 2.6005
R8437 VSS.n951 VSS.n950 2.6005
R8438 VSS.n950 VSS.n949 2.6005
R8439 VSS.n948 VSS.n947 2.6005
R8440 VSS.n947 VSS.n946 2.6005
R8441 VSS.n945 VSS.n944 2.6005
R8442 VSS.n944 VSS.n943 2.6005
R8443 VSS.n942 VSS.n941 2.6005
R8444 VSS.n941 VSS.n940 2.6005
R8445 VSS.n939 VSS.n938 2.6005
R8446 VSS.n938 VSS.n937 2.6005
R8447 VSS.n936 VSS.n935 2.6005
R8448 VSS.n935 VSS.n934 2.6005
R8449 VSS.n933 VSS.n932 2.6005
R8450 VSS.n932 VSS.n931 2.6005
R8451 VSS.n930 VSS.n929 2.6005
R8452 VSS.n929 VSS.n928 2.6005
R8453 VSS.n927 VSS.n926 2.6005
R8454 VSS.n926 VSS.n925 2.6005
R8455 VSS.n924 VSS.n923 2.6005
R8456 VSS.n923 VSS.n922 2.6005
R8457 VSS.n921 VSS.n920 2.6005
R8458 VSS.n920 VSS.n919 2.6005
R8459 VSS.n918 VSS.n917 2.6005
R8460 VSS.n917 VSS.n916 2.6005
R8461 VSS.n915 VSS.n914 2.6005
R8462 VSS.n914 VSS.n913 2.6005
R8463 VSS.n912 VSS.n911 2.6005
R8464 VSS.n911 VSS.n910 2.6005
R8465 VSS.n909 VSS.n908 2.6005
R8466 VSS.n908 VSS.n907 2.6005
R8467 VSS.n906 VSS.n905 2.6005
R8468 VSS.n905 VSS.n904 2.6005
R8469 VSS.n903 VSS.n902 2.6005
R8470 VSS.n902 VSS.n901 2.6005
R8471 VSS.n900 VSS.n899 2.6005
R8472 VSS.n899 VSS.n898 2.6005
R8473 VSS.n897 VSS.n896 2.6005
R8474 VSS.n896 VSS.n895 2.6005
R8475 VSS.n894 VSS.n893 2.6005
R8476 VSS.n893 VSS.n892 2.6005
R8477 VSS.n586 VSS.n585 2.6005
R8478 VSS.n585 VSS.n584 2.6005
R8479 VSS.n589 VSS.n588 2.6005
R8480 VSS.n588 VSS.n587 2.6005
R8481 VSS.n592 VSS.n591 2.6005
R8482 VSS.n591 VSS.n590 2.6005
R8483 VSS.n595 VSS.n594 2.6005
R8484 VSS.n594 VSS.n593 2.6005
R8485 VSS.n598 VSS.n597 2.6005
R8486 VSS.n597 VSS.n596 2.6005
R8487 VSS.n601 VSS.n600 2.6005
R8488 VSS.n600 VSS.n599 2.6005
R8489 VSS.n604 VSS.n603 2.6005
R8490 VSS.n603 VSS.n602 2.6005
R8491 VSS.n607 VSS.n606 2.6005
R8492 VSS.n606 VSS.n605 2.6005
R8493 VSS.n610 VSS.n609 2.6005
R8494 VSS.n609 VSS.n608 2.6005
R8495 VSS.n613 VSS.n612 2.6005
R8496 VSS.n612 VSS.n611 2.6005
R8497 VSS.n616 VSS.n615 2.6005
R8498 VSS.n615 VSS.n614 2.6005
R8499 VSS.n619 VSS.n618 2.6005
R8500 VSS.n618 VSS.n617 2.6005
R8501 VSS.n622 VSS.n621 2.6005
R8502 VSS.n621 VSS.n620 2.6005
R8503 VSS.n625 VSS.n624 2.6005
R8504 VSS.n624 VSS.n623 2.6005
R8505 VSS.n628 VSS.n627 2.6005
R8506 VSS.n627 VSS.n626 2.6005
R8507 VSS.n631 VSS.n630 2.6005
R8508 VSS.n630 VSS.n629 2.6005
R8509 VSS.n634 VSS.n633 2.6005
R8510 VSS.n633 VSS.n632 2.6005
R8511 VSS.n637 VSS.n636 2.6005
R8512 VSS.n636 VSS.n635 2.6005
R8513 VSS.n640 VSS.n639 2.6005
R8514 VSS.n639 VSS.n638 2.6005
R8515 VSS.n643 VSS.n642 2.6005
R8516 VSS.n642 VSS.n641 2.6005
R8517 VSS.n646 VSS.n645 2.6005
R8518 VSS.n645 VSS.n644 2.6005
R8519 VSS.n649 VSS.n648 2.6005
R8520 VSS.n648 VSS.n647 2.6005
R8521 VSS.n652 VSS.n651 2.6005
R8522 VSS.n651 VSS.n650 2.6005
R8523 VSS.n655 VSS.n654 2.6005
R8524 VSS.n654 VSS.n653 2.6005
R8525 VSS.n658 VSS.n657 2.6005
R8526 VSS.n657 VSS.n656 2.6005
R8527 VSS.n661 VSS.n660 2.6005
R8528 VSS.n660 VSS.n659 2.6005
R8529 VSS.n664 VSS.n663 2.6005
R8530 VSS.n663 VSS.n662 2.6005
R8531 VSS.n667 VSS.n666 2.6005
R8532 VSS.n666 VSS.n665 2.6005
R8533 VSS.n670 VSS.n669 2.6005
R8534 VSS.n669 VSS.n668 2.6005
R8535 VSS.n673 VSS.n672 2.6005
R8536 VSS.n672 VSS.n671 2.6005
R8537 VSS.n676 VSS.n675 2.6005
R8538 VSS.n675 VSS.n674 2.6005
R8539 VSS.n679 VSS.n678 2.6005
R8540 VSS.n678 VSS.n677 2.6005
R8541 VSS.n682 VSS.n681 2.6005
R8542 VSS.n681 VSS.n680 2.6005
R8543 VSS.n685 VSS.n684 2.6005
R8544 VSS.n684 VSS.n683 2.6005
R8545 VSS.n688 VSS.n687 2.6005
R8546 VSS.n687 VSS.n686 2.6005
R8547 VSS.n691 VSS.n690 2.6005
R8548 VSS.n690 VSS.n689 2.6005
R8549 VSS.n694 VSS.n693 2.6005
R8550 VSS.n693 VSS.n692 2.6005
R8551 VSS.n697 VSS.n696 2.6005
R8552 VSS.n696 VSS.n695 2.6005
R8553 VSS.n700 VSS.n699 2.6005
R8554 VSS.n699 VSS.n698 2.6005
R8555 VSS.n703 VSS.n702 2.6005
R8556 VSS.n702 VSS.n701 2.6005
R8557 VSS.n706 VSS.n705 2.6005
R8558 VSS.n705 VSS.n704 2.6005
R8559 VSS.n709 VSS.n708 2.6005
R8560 VSS.n708 VSS.n707 2.6005
R8561 VSS.n712 VSS.n711 2.6005
R8562 VSS.n711 VSS.n710 2.6005
R8563 VSS.n715 VSS.n714 2.6005
R8564 VSS.n714 VSS.n713 2.6005
R8565 VSS.n718 VSS.n717 2.6005
R8566 VSS.n717 VSS.n716 2.6005
R8567 VSS.n721 VSS.n720 2.6005
R8568 VSS.n720 VSS.n719 2.6005
R8569 VSS.n724 VSS.n723 2.6005
R8570 VSS.n723 VSS.n722 2.6005
R8571 VSS.n727 VSS.n726 2.6005
R8572 VSS.n726 VSS.n725 2.6005
R8573 VSS.n563 VSS.n562 2.6005
R8574 VSS.n562 VSS.n561 2.6005
R8575 VSS.n569 VSS.n568 2.6005
R8576 VSS.n568 VSS.n567 2.6005
R8577 VSS.n579 VSS.n578 2.6005
R8578 VSS.n578 VSS.n577 2.6005
R8579 VSS.n740 VSS.n739 2.6005
R8580 VSS.n739 VSS.n738 2.6005
R8581 VSS.n380 VSS.n379 2.6005
R8582 VSS.n379 VSS.n378 2.6005
R8583 VSS.n383 VSS.n382 2.6005
R8584 VSS.n382 VSS.n381 2.6005
R8585 VSS.n386 VSS.n385 2.6005
R8586 VSS.n385 VSS.n384 2.6005
R8587 VSS.n389 VSS.n388 2.6005
R8588 VSS.n388 VSS.n387 2.6005
R8589 VSS.n392 VSS.n391 2.6005
R8590 VSS.n391 VSS.n390 2.6005
R8591 VSS.n395 VSS.n394 2.6005
R8592 VSS.n394 VSS.n393 2.6005
R8593 VSS.n398 VSS.n397 2.6005
R8594 VSS.n397 VSS.n396 2.6005
R8595 VSS.n401 VSS.n400 2.6005
R8596 VSS.n400 VSS.n399 2.6005
R8597 VSS.n404 VSS.n403 2.6005
R8598 VSS.n403 VSS.n402 2.6005
R8599 VSS.n407 VSS.n406 2.6005
R8600 VSS.n406 VSS.n405 2.6005
R8601 VSS.n410 VSS.n409 2.6005
R8602 VSS.n409 VSS.n408 2.6005
R8603 VSS.n412 VSS.n411 2.6005
R8604 VSS.n415 VSS.n414 2.6005
R8605 VSS.n417 VSS.n416 2.6005
R8606 VSS.n421 VSS.n420 2.6005
R8607 VSS.n424 VSS.n423 2.6005
R8608 VSS.n423 VSS.n422 2.6005
R8609 VSS.n3814 VSS.n3813 2.6005
R8610 VSS.n3813 VSS.n3812 2.6005
R8611 VSS.n3811 VSS.n3810 2.6005
R8612 VSS.n3810 VSS.n3809 2.6005
R8613 VSS.n3808 VSS.n3807 2.6005
R8614 VSS.n3807 VSS.n3806 2.6005
R8615 VSS.n3805 VSS.n3804 2.6005
R8616 VSS.n3804 VSS.n3803 2.6005
R8617 VSS.n3802 VSS.n3801 2.6005
R8618 VSS.n3801 VSS.n3800 2.6005
R8619 VSS.n3799 VSS.n3798 2.6005
R8620 VSS.n3798 VSS.n3797 2.6005
R8621 VSS.n3796 VSS.n3795 2.6005
R8622 VSS.n3795 VSS.n3794 2.6005
R8623 VSS.n3793 VSS.n3792 2.6005
R8624 VSS.n3792 VSS.n3791 2.6005
R8625 VSS.n3790 VSS.n3789 2.6005
R8626 VSS.n3789 VSS.n3788 2.6005
R8627 VSS.n3787 VSS.n3786 2.6005
R8628 VSS.n3786 VSS.n3785 2.6005
R8629 VSS.n3784 VSS.n3783 2.6005
R8630 VSS.n3783 VSS.n3782 2.6005
R8631 VSS.n3781 VSS.n3780 2.6005
R8632 VSS.n3780 VSS.n3779 2.6005
R8633 VSS.n3778 VSS.n3777 2.6005
R8634 VSS.n3777 VSS.n3776 2.6005
R8635 VSS.n2613 VSS.n2612 2.6005
R8636 VSS.n2612 VSS.n2611 2.6005
R8637 VSS.n2616 VSS.n2615 2.6005
R8638 VSS.n2615 VSS.n2614 2.6005
R8639 VSS.n2619 VSS.n2618 2.6005
R8640 VSS.n2618 VSS.n2617 2.6005
R8641 VSS.n2622 VSS.n2621 2.6005
R8642 VSS.n2621 VSS.n2620 2.6005
R8643 VSS.n2626 VSS.n2625 2.6005
R8644 VSS.n2625 VSS.n2624 2.6005
R8645 VSS.n2629 VSS.n2628 2.6005
R8646 VSS.n2628 VSS.n2627 2.6005
R8647 VSS.n2632 VSS.n2631 2.6005
R8648 VSS.n2631 VSS.n2630 2.6005
R8649 VSS.n2635 VSS.n2634 2.6005
R8650 VSS.n2634 VSS.n2633 2.6005
R8651 VSS.n2638 VSS.n2637 2.6005
R8652 VSS.n2637 VSS.n2636 2.6005
R8653 VSS.n2641 VSS.n2640 2.6005
R8654 VSS.n2640 VSS.n2639 2.6005
R8655 VSS.n2644 VSS.n2643 2.6005
R8656 VSS.n2643 VSS.n2642 2.6005
R8657 VSS.n2647 VSS.n2646 2.6005
R8658 VSS.n2646 VSS.n2645 2.6005
R8659 VSS.n2650 VSS.n2649 2.6005
R8660 VSS.n2649 VSS.n2648 2.6005
R8661 VSS.n2653 VSS.n2652 2.6005
R8662 VSS.n2652 VSS.n2651 2.6005
R8663 VSS.n2656 VSS.n2655 2.6005
R8664 VSS.n2655 VSS.n2654 2.6005
R8665 VSS.n2659 VSS.n2658 2.6005
R8666 VSS.n2658 VSS.n2657 2.6005
R8667 VSS.n2662 VSS.n2661 2.6005
R8668 VSS.n2661 VSS.n2660 2.6005
R8669 VSS.n2665 VSS.n2664 2.6005
R8670 VSS.n2664 VSS.n2663 2.6005
R8671 VSS.n2668 VSS.n2667 2.6005
R8672 VSS.n2667 VSS.n2666 2.6005
R8673 VSS.n2671 VSS.n2670 2.6005
R8674 VSS.n2670 VSS.n2669 2.6005
R8675 VSS.n2674 VSS.n2673 2.6005
R8676 VSS.n2673 VSS.n2672 2.6005
R8677 VSS.n2677 VSS.n2676 2.6005
R8678 VSS.n2676 VSS.n2675 2.6005
R8679 VSS.n2680 VSS.n2679 2.6005
R8680 VSS.n2679 VSS.n2678 2.6005
R8681 VSS.n2683 VSS.n2682 2.6005
R8682 VSS.n2682 VSS.n2681 2.6005
R8683 VSS.n2686 VSS.n2685 2.6005
R8684 VSS.n2685 VSS.n2684 2.6005
R8685 VSS.n2689 VSS.n2688 2.6005
R8686 VSS.n2688 VSS.n2687 2.6005
R8687 VSS.n2692 VSS.n2691 2.6005
R8688 VSS.n2691 VSS.n2690 2.6005
R8689 VSS.n2695 VSS.n2694 2.6005
R8690 VSS.n2694 VSS.n2693 2.6005
R8691 VSS.n2698 VSS.n2697 2.6005
R8692 VSS.n2697 VSS.n2696 2.6005
R8693 VSS.n2701 VSS.n2700 2.6005
R8694 VSS.n2700 VSS.n2699 2.6005
R8695 VSS.n2704 VSS.n2703 2.6005
R8696 VSS.n2703 VSS.n2702 2.6005
R8697 VSS.n2707 VSS.n2706 2.6005
R8698 VSS.n2706 VSS.n2705 2.6005
R8699 VSS.n2710 VSS.n2709 2.6005
R8700 VSS.n2709 VSS.n2708 2.6005
R8701 VSS.n2713 VSS.n2712 2.6005
R8702 VSS.n2712 VSS.n2711 2.6005
R8703 VSS.n2716 VSS.n2715 2.6005
R8704 VSS.n2715 VSS.n2714 2.6005
R8705 VSS.n2719 VSS.n2718 2.6005
R8706 VSS.n2718 VSS.n2717 2.6005
R8707 VSS.n2722 VSS.n2721 2.6005
R8708 VSS.n2721 VSS.n2720 2.6005
R8709 VSS.n2725 VSS.n2724 2.6005
R8710 VSS.n2724 VSS.n2723 2.6005
R8711 VSS.n2728 VSS.n2727 2.6005
R8712 VSS.n2727 VSS.n2726 2.6005
R8713 VSS.n2731 VSS.n2730 2.6005
R8714 VSS.n2730 VSS.n2729 2.6005
R8715 VSS.n2734 VSS.n2733 2.6005
R8716 VSS.n2733 VSS.n2732 2.6005
R8717 VSS.n2737 VSS.n2736 2.6005
R8718 VSS.n2736 VSS.n2735 2.6005
R8719 VSS.n2740 VSS.n2739 2.6005
R8720 VSS.n2739 VSS.n2738 2.6005
R8721 VSS.n2743 VSS.n2742 2.6005
R8722 VSS.n2742 VSS.n2741 2.6005
R8723 VSS.n2746 VSS.n2745 2.6005
R8724 VSS.n2745 VSS.n2744 2.6005
R8725 VSS.n2749 VSS.n2748 2.6005
R8726 VSS.n2748 VSS.n2747 2.6005
R8727 VSS.n2752 VSS.n2751 2.6005
R8728 VSS.n2751 VSS.n2750 2.6005
R8729 VSS.n2755 VSS.n2754 2.6005
R8730 VSS.n2754 VSS.n2753 2.6005
R8731 VSS.n2758 VSS.n2757 2.6005
R8732 VSS.n2757 VSS.n2756 2.6005
R8733 VSS.n2761 VSS.n2760 2.6005
R8734 VSS.n2760 VSS.n2759 2.6005
R8735 VSS.n2764 VSS.n2763 2.6005
R8736 VSS.n2763 VSS.n2762 2.6005
R8737 VSS.n2767 VSS.n2766 2.6005
R8738 VSS.n2766 VSS.n2765 2.6005
R8739 VSS.n2770 VSS.n2769 2.6005
R8740 VSS.n2769 VSS.n2768 2.6005
R8741 VSS.n2773 VSS.n2772 2.6005
R8742 VSS.n2772 VSS.n2771 2.6005
R8743 VSS.n2776 VSS.n2775 2.6005
R8744 VSS.n2775 VSS.n2774 2.6005
R8745 VSS.n2779 VSS.n2778 2.6005
R8746 VSS.n2778 VSS.n2777 2.6005
R8747 VSS.n2783 VSS.n2782 2.6005
R8748 VSS.n2782 VSS.n2781 2.6005
R8749 VSS.n2786 VSS.n2785 2.6005
R8750 VSS.n2785 VSS.n2784 2.6005
R8751 VSS.n2789 VSS.n2788 2.6005
R8752 VSS.n2788 VSS.n2787 2.6005
R8753 VSS.n2792 VSS.n2791 2.6005
R8754 VSS.n2791 VSS.n2790 2.6005
R8755 VSS.n2795 VSS.n2794 2.6005
R8756 VSS.n2794 VSS.n2793 2.6005
R8757 VSS.n2798 VSS.n2797 2.6005
R8758 VSS.n2797 VSS.n2796 2.6005
R8759 VSS.n2801 VSS.n2800 2.6005
R8760 VSS.n2800 VSS.n2799 2.6005
R8761 VSS.n2804 VSS.n2803 2.6005
R8762 VSS.n2803 VSS.n2802 2.6005
R8763 VSS.n2807 VSS.n2806 2.6005
R8764 VSS.n2806 VSS.n2805 2.6005
R8765 VSS.n2810 VSS.n2809 2.6005
R8766 VSS.n2809 VSS.n2808 2.6005
R8767 VSS.n2813 VSS.n2812 2.6005
R8768 VSS.n2812 VSS.n2811 2.6005
R8769 VSS.n2816 VSS.n2815 2.6005
R8770 VSS.n2815 VSS.n2814 2.6005
R8771 VSS.n2819 VSS.n2818 2.6005
R8772 VSS.n2818 VSS.n2817 2.6005
R8773 VSS.n2962 VSS.n2961 2.6005
R8774 VSS.n2961 VSS.n2960 2.6005
R8775 VSS.n2964 VSS.n2963 2.6005
R8776 VSS.n2966 VSS.n2965 2.6005
R8777 VSS.n2968 VSS.n2967 2.6005
R8778 VSS.n2970 VSS.n2969 2.6005
R8779 VSS.n2972 VSS.n2971 2.6005
R8780 VSS.n2975 VSS.n2974 2.6005
R8781 VSS.n2977 VSS.n2976 2.6005
R8782 VSS.n2980 VSS.n2979 2.6005
R8783 VSS.n2982 VSS.n2981 2.6005
R8784 VSS.n2985 VSS.n2984 2.6005
R8785 VSS.n2987 VSS.n2986 2.6005
R8786 VSS.n2990 VSS.n2989 2.6005
R8787 VSS.n2992 VSS.n2991 2.6005
R8788 VSS.n2995 VSS.n2994 2.6005
R8789 VSS.n2997 VSS.n2996 2.6005
R8790 VSS.n3000 VSS.n2999 2.6005
R8791 VSS.n3002 VSS.n3001 2.6005
R8792 VSS.n3008 VSS.n3007 2.6005
R8793 VSS.n3010 VSS.n3009 2.6005
R8794 VSS.n3013 VSS.n3012 2.6005
R8795 VSS.n3015 VSS.n3014 2.6005
R8796 VSS.n3018 VSS.n3017 2.6005
R8797 VSS.n3020 VSS.n3019 2.6005
R8798 VSS.n3024 VSS.n3023 2.6005
R8799 VSS.n3026 VSS.n3025 2.6005
R8800 VSS.n3028 VSS.n3027 2.6005
R8801 VSS.n3030 VSS.n3029 2.6005
R8802 VSS.n3032 VSS.n3031 2.6005
R8803 VSS.n3034 VSS.n3033 2.6005
R8804 VSS.n3036 VSS.n3035 2.6005
R8805 VSS.n3038 VSS.n3037 2.6005
R8806 VSS.n3040 VSS.n3039 2.6005
R8807 VSS.n3042 VSS.n3041 2.6005
R8808 VSS.n3044 VSS.n3043 2.6005
R8809 VSS.n3046 VSS.n3045 2.6005
R8810 VSS.n3048 VSS.n3047 2.6005
R8811 VSS.n3050 VSS.n3049 2.6005
R8812 VSS.n3052 VSS.n3051 2.6005
R8813 VSS.n3054 VSS.n3053 2.6005
R8814 VSS.n3057 VSS.n3056 2.6005
R8815 VSS.n3059 VSS.n3058 2.6005
R8816 VSS.n3062 VSS.n3061 2.6005
R8817 VSS.n3064 VSS.n3063 2.6005
R8818 VSS.n3067 VSS.n3066 2.6005
R8819 VSS.n3069 VSS.n3068 2.6005
R8820 VSS.n3072 VSS.n3071 2.6005
R8821 VSS.n3074 VSS.n3073 2.6005
R8822 VSS.n3077 VSS.n3076 2.6005
R8823 VSS.n3079 VSS.n3078 2.6005
R8824 VSS.n3082 VSS.n3081 2.6005
R8825 VSS.n3084 VSS.n3083 2.6005
R8826 VSS.n3095 VSS.n3094 2.6005
R8827 VSS.n3097 VSS.n3096 2.6005
R8828 VSS.n3817 VSS.n3816 2.6005
R8829 VSS.n3816 VSS.n3815 2.6005
R8830 VSS.n3221 VSS.n3220 2.6005
R8831 VSS.n3218 VSS.n3217 2.6005
R8832 VSS.n3216 VSS.n3215 2.6005
R8833 VSS.n3213 VSS.n3212 2.6005
R8834 VSS.n3211 VSS.n3210 2.6005
R8835 VSS.n3208 VSS.n3207 2.6005
R8836 VSS.n3206 VSS.n3205 2.6005
R8837 VSS.n3203 VSS.n3202 2.6005
R8838 VSS.n3201 VSS.n3200 2.6005
R8839 VSS.n3198 VSS.n3197 2.6005
R8840 VSS.n3196 VSS.n3195 2.6005
R8841 VSS.n3193 VSS.n3192 2.6005
R8842 VSS.n3191 VSS.n3190 2.6005
R8843 VSS.n3189 VSS.n3188 2.6005
R8844 VSS.n3187 VSS.n3186 2.6005
R8845 VSS.n3185 VSS.n3184 2.6005
R8846 VSS.n3183 VSS.n3182 2.6005
R8847 VSS.n3181 VSS.n3180 2.6005
R8848 VSS.n3179 VSS.n3178 2.6005
R8849 VSS.n3177 VSS.n3176 2.6005
R8850 VSS.n3175 VSS.n3174 2.6005
R8851 VSS.n3173 VSS.n3172 2.6005
R8852 VSS.n3171 VSS.n3170 2.6005
R8853 VSS.n3169 VSS.n3168 2.6005
R8854 VSS.n3167 VSS.n3166 2.6005
R8855 VSS.n3165 VSS.n3164 2.6005
R8856 VSS.n3163 VSS.n3162 2.6005
R8857 VSS.n3161 VSS.n3160 2.6005
R8858 VSS.n3159 VSS.n3158 2.6005
R8859 VSS.n3157 VSS.n3156 2.6005
R8860 VSS.n3155 VSS.n3154 2.6005
R8861 VSS.n3153 VSS.n3152 2.6005
R8862 VSS.n3151 VSS.n3150 2.6005
R8863 VSS.n3149 VSS.n3148 2.6005
R8864 VSS.n3147 VSS.n3146 2.6005
R8865 VSS.n3145 VSS.n3144 2.6005
R8866 VSS.n3143 VSS.n3142 2.6005
R8867 VSS.n3141 VSS.n3140 2.6005
R8868 VSS.n3139 VSS.n3138 2.6005
R8869 VSS.n3137 VSS.n3136 2.6005
R8870 VSS.n3135 VSS.n3134 2.6005
R8871 VSS.n3133 VSS.n3132 2.6005
R8872 VSS.n3131 VSS.n3130 2.6005
R8873 VSS.n3129 VSS.n3128 2.6005
R8874 VSS.n3127 VSS.n3126 2.6005
R8875 VSS.n3223 VSS.n3222 2.6005
R8876 VSS.n3284 VSS.n3283 2.6005
R8877 VSS.n2535 VSS.n2534 2.50768
R8878 VSS.n3757 VSS.t1248 2.41806
R8879 VSS.n35 VSS.n34 2.41121
R8880 VSS.n4013 VSS.n4012 2.39694
R8881 VSS.n2535 VSS.n2430 2.39323
R8882 VSS.n2908 VSS.n2907 2.38577
R8883 VSS.n5083 VSS.n5082 2.36606
R8884 VSS.n232 VSS.n231 2.36606
R8885 VSS.n284 VSS.n283 2.36606
R8886 VSS.n5053 VSS.n5052 2.36606
R8887 VSS.n104 VSS.n103 2.36606
R8888 VSS.n143 VSS.n142 2.36606
R8889 VSS.n185 VSS.n184 2.36606
R8890 VSS.n202 VSS.n201 2.36606
R8891 VSS.n120 VSS.n119 2.36606
R8892 VSS.n4358 VSS.n4357 2.36061
R8893 VSS.n2909 VSS.n2908 2.35343
R8894 VSS.n5482 VSS.n5481 2.31421
R8895 VSS.n1048 VSS.n1045 2.25899
R8896 VSS.n5169 VSS.n5142 2.25386
R8897 VSS.n2903 VSS.n2902 2.25315
R8898 VSS.n1688 VSS.n1687 2.25238
R8899 VSS.n3993 VSS.n3992 2.25176
R8900 VSS.n3543 VSS.n3534 2.25176
R8901 VSS.n3980 VSS.n3763 2.25176
R8902 VSS.n5123 VSS.n5122 2.2505
R8903 VSS.n255 VSS.n254 2.2505
R8904 VSS.n5045 VSS.n5044 2.2505
R8905 VSS.n5056 VSS.n5055 2.2505
R8906 VSS.n2512 VSS.n2511 2.2505
R8907 VSS.n117 VSS.n116 2.2505
R8908 VSS.n5489 VSS.n5488 2.2505
R8909 VSS.n5460 VSS.n5459 2.2505
R8910 VSS.n5441 VSS.n5440 2.2505
R8911 VSS.n199 VSS.n198 2.2505
R8912 VSS.n214 VSS.n213 2.2505
R8913 VSS.n164 VSS.n163 2.2505
R8914 VSS.n5425 VSS.n5424 2.2505
R8915 VSS.n4014 VSS.n4013 2.2505
R8916 VSS.n5131 VSS.n5130 2.2505
R8917 VSS.n730 VSS.n729 2.2505
R8918 VSS.n5168 VSS.n5167 2.2505
R8919 VSS.n744 VSS.n743 2.2505
R8920 VSS.n573 VSS.n572 2.2505
R8921 VSS.n734 VSS.n733 2.2505
R8922 VSS.n583 VSS.n582 2.2505
R8923 VSS.n2295 VSS.n2294 2.2505
R8924 VSS.n1051 VSS.n1050 2.2505
R8925 VSS.n1057 VSS.n1056 2.2505
R8926 VSS.n1054 VSS.n1053 2.2505
R8927 VSS.n1762 VSS.n1761 2.2505
R8928 VSS.n786 VSS.n785 2.2505
R8929 VSS.n860 VSS.n859 2.2505
R8930 VSS.n986 VSS.n985 2.2505
R8931 VSS.n873 VSS.n872 2.2505
R8932 VSS.n883 VSS.n882 2.2505
R8933 VSS.n5013 VSS.n5012 2.2505
R8934 VSS.n3545 VSS.n3544 2.2505
R8935 VSS.n3546 VSS.n3545 2.2505
R8936 VSS.n3511 VSS.n3510 2.2505
R8937 VSS.n3534 VSS.n3533 2.2505
R8938 VSS.n3519 VSS.n3518 2.2505
R8939 VSS.n3517 VSS.n3516 2.2505
R8940 VSS.n2590 VSS.n1694 2.2505
R8941 VSS.n4044 VSS.n4043 2.2505
R8942 VSS.n4174 VSS.n4173 2.2505
R8943 VSS.n4173 VSS.n4172 2.2505
R8944 VSS.n2312 VSS.n2311 2.2505
R8945 VSS.n2313 VSS.n2312 2.2505
R8946 VSS.n2320 VSS.n2295 2.2505
R8947 VSS.n2300 VSS.n2299 2.2505
R8948 VSS.n2301 VSS.n2300 2.2505
R8949 VSS.n2309 VSS.n2308 2.2505
R8950 VSS.n2310 VSS.n2309 2.2505
R8951 VSS.n4171 VSS.n4170 2.2505
R8952 VSS.n2318 VSS.n2317 2.2505
R8953 VSS.n2319 VSS.n2318 2.2505
R8954 VSS.n2297 VSS.n2296 2.2505
R8955 VSS.n2298 VSS.n2297 2.2505
R8956 VSS.n2043 VSS.n1762 2.2505
R8957 VSS.n2060 VSS.n2059 2.2505
R8958 VSS.n2061 VSS.n2060 2.2505
R8959 VSS.n2072 VSS.n2071 2.2505
R8960 VSS.n2073 VSS.n2072 2.2505
R8961 VSS.n2051 VSS.n2050 2.2505
R8962 VSS.n2052 VSS.n2051 2.2505
R8963 VSS.n2057 VSS.n2056 2.2505
R8964 VSS.n2058 VSS.n2057 2.2505
R8965 VSS.n2042 VSS.n2041 2.2505
R8966 VSS.n2069 VSS.n2068 2.2505
R8967 VSS.n2070 VSS.n2069 2.2505
R8968 VSS.n2048 VSS.n2047 2.2505
R8969 VSS.n2049 VSS.n2048 2.2505
R8970 VSS.n5162 VSS.n5161 2.2505
R8971 VSS.n5157 VSS.n5156 2.2505
R8972 VSS.n5151 VSS.n5150 2.2505
R8973 VSS.n5153 VSS.n5152 2.2505
R8974 VSS.n5165 VSS.n5164 2.2505
R8975 VSS.n5159 VSS.n5143 2.2505
R8976 VSS.n5147 VSS.n5146 2.2505
R8977 VSS.n3496 VSS.n3495 2.2505
R8978 VSS.n3504 VSS.n3503 2.2505
R8979 VSS.n3505 VSS.n3504 2.2505
R8980 VSS.n3997 VSS.n3996 2.2505
R8981 VSS.n3487 VSS.n3486 2.2505
R8982 VSS.n3499 VSS.n3498 2.2505
R8983 VSS.n3994 VSS.n3993 2.2505
R8984 VSS.n3490 VSS.n3489 2.2505
R8985 VSS.n3508 VSS.n3507 2.2505
R8986 VSS.n3996 VSS.n3995 2.2505
R8987 VSS.n3495 VSS.n3494 2.2505
R8988 VSS.n3486 VSS.n3485 2.2505
R8989 VSS.n3498 VSS.n3497 2.2505
R8990 VSS.n3489 VSS.n3488 2.2505
R8991 VSS.n3507 VSS.n3506 2.2505
R8992 VSS.n3771 VSS.n3770 2.2505
R8993 VSS.n3763 VSS.n3762 2.2505
R8994 VSS.n3979 VSS.n3978 2.2505
R8995 VSS.n3978 VSS.n3977 2.2505
R8996 VSS.n3765 VSS.n3764 2.2505
R8997 VSS.n3773 VSS.n3772 2.2505
R8998 VSS.n3767 VSS.n3766 2.2505
R8999 VSS.n3775 VSS.n3774 2.2505
R9000 VSS.n1687 VSS.n1686 2.2505
R9001 VSS.n1685 VSS.n1684 2.2505
R9002 VSS.n1684 VSS.n1683 2.2505
R9003 VSS.n1151 VSS.n1150 2.2505
R9004 VSS.n1149 VSS.n1148 2.2505
R9005 VSS.n1153 VSS.n1152 2.2505
R9006 VSS.n1514 VSS.n1387 2.2505
R9007 VSS.n1516 VSS.n1515 2.2505
R9008 VSS.n1530 VSS.n1529 2.2505
R9009 VSS.n1537 VSS.n1536 2.2505
R9010 VSS.n1523 VSS.n1522 2.2505
R9011 VSS.n1528 VSS.n1527 2.2505
R9012 VSS.n1535 VSS.n1534 2.2505
R9013 VSS.n1521 VSS.n1520 2.2505
R9014 VSS.n985 VSS.n984 2.2505
R9015 VSS.n984 VSS.n983 2.2505
R9016 VSS.n885 VSS.n884 2.2505
R9017 VSS.n866 VSS.n865 2.2505
R9018 VSS.n865 VSS.n864 2.2505
R9019 VSS.n879 VSS.n878 2.2505
R9020 VSS.n878 VSS.n877 2.2505
R9021 VSS.n872 VSS.n871 2.2505
R9022 VSS.n871 VSS.n870 2.2505
R9023 VSS.n859 VSS.n858 2.2505
R9024 VSS.n858 VSS.n857 2.2505
R9025 VSS.n882 VSS.n881 2.2505
R9026 VSS.n881 VSS.n880 2.2505
R9027 VSS.n743 VSS.n742 2.2505
R9028 VSS.n742 VSS.n741 2.2505
R9029 VSS.n576 VSS.n575 2.2505
R9030 VSS.n575 VSS.n574 2.2505
R9031 VSS.n566 VSS.n565 2.2505
R9032 VSS.n565 VSS.n564 2.2505
R9033 VSS.n736 VSS.n735 2.2505
R9034 VSS.n729 VSS.n728 2.2505
R9035 VSS.n572 VSS.n571 2.2505
R9036 VSS.n571 VSS.n570 2.2505
R9037 VSS.n733 VSS.n732 2.2505
R9038 VSS.n732 VSS.n731 2.2505
R9039 VSS.n582 VSS.n581 2.2505
R9040 VSS.n581 VSS.n580 2.2505
R9041 VSS.n4006 VSS.n4005 2.2505
R9042 VSS.n4008 VSS.n4007 2.2505
R9043 VSS.n4011 VSS.n4010 2.2505
R9044 VSS.n4461 VSS.n4460 2.17921
R9045 VSS.n313 VSS.n312 2.17921
R9046 VSS.n4342 VSS.n4341 2.17771
R9047 VSS.n4512 VSS.n753 2.17664
R9048 VSS.n365 VSS.n364 2.17664
R9049 VSS.n4150 VSS.n4149 2.10867
R9050 VSS.n2468 VSS.n2467 1.99937
R9051 VSS.n5185 VSS.n5183 1.97486
R9052 VSS.n4110 VSS.n4106 1.91985
R9053 VSS.n2936 VSS.n2934 1.90173
R9054 VSS.n4151 VSS.n35 1.83722
R9055 VSS.n4010 VSS.n4009 1.8127
R9056 VSS.n5195 VSS.n5191 1.79537
R9057 VSS.n5218 VSS.n5216 1.79537
R9058 VSS.n3924 VSS.n3922 1.74053
R9059 VSS.n3927 VSS.n3925 1.74053
R9060 VSS.n3930 VSS.n3928 1.74053
R9061 VSS.n3933 VSS.n3931 1.74053
R9062 VSS.n3936 VSS.n3934 1.74053
R9063 VSS.n3939 VSS.n3937 1.74053
R9064 VSS.n3942 VSS.n3940 1.74053
R9065 VSS.n3945 VSS.n3943 1.74053
R9066 VSS.n3948 VSS.n3946 1.74053
R9067 VSS.n3951 VSS.n3949 1.74053
R9068 VSS.n3954 VSS.n3952 1.74053
R9069 VSS.n3956 VSS.n3955 1.74053
R9070 VSS.n1369 VSS.n1366 1.74053
R9071 VSS.n1374 VSS.n1371 1.74053
R9072 VSS.n1379 VSS.n1376 1.74053
R9073 VSS.n1384 VSS.n1381 1.74053
R9074 VSS.n1678 VSS.n1386 1.74053
R9075 VSS.n1647 VSS.n1646 1.74053
R9076 VSS.n1638 VSS.n1637 1.74053
R9077 VSS.n1633 VSS.n1632 1.74053
R9078 VSS.n1628 VSS.n1627 1.74053
R9079 VSS.n3924 VSS.n3923 1.73995
R9080 VSS.n3927 VSS.n3926 1.73995
R9081 VSS.n3930 VSS.n3929 1.73995
R9082 VSS.n3933 VSS.n3932 1.73995
R9083 VSS.n3936 VSS.n3935 1.73995
R9084 VSS.n3939 VSS.n3938 1.73995
R9085 VSS.n3942 VSS.n3941 1.73995
R9086 VSS.n3945 VSS.n3944 1.73995
R9087 VSS.n3948 VSS.n3947 1.73995
R9088 VSS.n3951 VSS.n3950 1.73995
R9089 VSS.n3954 VSS.n3953 1.73995
R9090 VSS.n3896 VSS.n3895 1.73995
R9091 VSS.n3901 VSS.n3900 1.73995
R9092 VSS.n3906 VSS.n3905 1.73995
R9093 VSS.n3911 VSS.n3910 1.73995
R9094 VSS.n3971 VSS.n3970 1.73995
R9095 VSS.n1155 VSS.n1154 1.73995
R9096 VSS.n1340 VSS.n1339 1.73995
R9097 VSS.n1345 VSS.n1344 1.73995
R9098 VSS.n1350 VSS.n1349 1.73995
R9099 VSS.n1358 VSS.n1357 1.73995
R9100 VSS.n1681 VSS.n1680 1.73995
R9101 VSS.n1369 VSS.n1368 1.73995
R9102 VSS.n1374 VSS.n1373 1.73995
R9103 VSS.n1379 VSS.n1378 1.73995
R9104 VSS.n1384 VSS.n1383 1.73995
R9105 VSS.n1678 VSS.n1677 1.73995
R9106 VSS.n414 VSS.n413 1.73995
R9107 VSS.n420 VSS.n419 1.73995
R9108 VSS.n3921 VSS.n3919 1.72551
R9109 VSS.n3921 VSS.n3920 1.72493
R9110 VSS.n4115 VSS.n4112 1.65384
R9111 VSS.n4144 VSS.n4143 1.65384
R9112 VSS.n2416 VSS.n2415 1.65384
R9113 VSS.n2411 VSS.n2410 1.65384
R9114 VSS.n2390 VSS.n2387 1.65384
R9115 VSS.n4115 VSS.n4114 1.65327
R9116 VSS.n2390 VSS.n2389 1.65327
R9117 VSS.n4366 VSS.n1075 1.64468
R9118 VSS.n1768 VSS.n1766 1.61588
R9119 VSS.n4483 VSS.n4482 1.58545
R9120 VSS.n4323 VSS.n4181 1.54391
R9121 VSS.n2040 VSS.n2037 1.51729
R9122 VSS.n4392 VSS.n4391 1.5047
R9123 VSS.n5170 VSS.n5169 1.50064
R9124 VSS.n4046 VSS.n4045 1.4973
R9125 VSS.n4345 VSS.n1694 1.49567
R9126 VSS.n5285 VSS.n5284 1.49293
R9127 VSS.n5290 VSS.n5289 1.49293
R9128 VSS.n5320 VSS.n5319 1.49293
R9129 VSS.n4764 VSS.n4763 1.49293
R9130 VSS.n4769 VSS.n4768 1.49293
R9131 VSS.n4774 VSS.n4773 1.49293
R9132 VSS.n4779 VSS.n4778 1.49293
R9133 VSS.n4809 VSS.n4808 1.49293
R9134 VSS.n4890 VSS.n4889 1.49293
R9135 VSS.n4895 VSS.n4894 1.49293
R9136 VSS.n4900 VSS.n4899 1.49293
R9137 VSS.n4905 VSS.n4904 1.49293
R9138 VSS.n4910 VSS.n4909 1.49293
R9139 VSS.n5280 VSS.n5279 1.49293
R9140 VSS.n4719 VSS.n4718 1.4928
R9141 VSS.n4724 VSS.n4723 1.4928
R9142 VSS.n4729 VSS.n4728 1.4928
R9143 VSS.n4734 VSS.n4733 1.4928
R9144 VSS.n4739 VSS.n4738 1.4928
R9145 VSS.n4744 VSS.n4743 1.4928
R9146 VSS.n4943 VSS.n4942 1.4928
R9147 VSS.n4848 VSS.n4847 1.4928
R9148 VSS.n4843 VSS.n4842 1.4928
R9149 VSS.n4838 VSS.n4837 1.4928
R9150 VSS.n4833 VSS.n4832 1.4928
R9151 VSS.n4828 VSS.n4827 1.4928
R9152 VSS.n4823 VSS.n4822 1.4928
R9153 VSS.n4818 VSS.n4817 1.4928
R9154 VSS.n4804 VSS.n4803 1.4928
R9155 VSS.n5359 VSS.n5358 1.4928
R9156 VSS.n5354 VSS.n5353 1.4928
R9157 VSS.n5349 VSS.n5348 1.4928
R9158 VSS.n5344 VSS.n5343 1.4928
R9159 VSS.n5339 VSS.n5338 1.4928
R9160 VSS.n5334 VSS.n5333 1.4928
R9161 VSS.n5329 VSS.n5328 1.4928
R9162 VSS.n5315 VSS.n5314 1.4928
R9163 VSS.n3280 VSS.n3279 1.47425
R9164 VSS.n3280 VSS.n3278 1.47372
R9165 VSS.n3094 VSS.n3093 1.47372
R9166 VSS.n3081 VSS.n3080 1.47372
R9167 VSS.n3076 VSS.n3075 1.47372
R9168 VSS.n3071 VSS.n3070 1.47372
R9169 VSS.n3066 VSS.n3065 1.47372
R9170 VSS.n3061 VSS.n3060 1.47372
R9171 VSS.n3056 VSS.n3055 1.47372
R9172 VSS.n3023 VSS.n3022 1.47372
R9173 VSS.n3017 VSS.n3016 1.47372
R9174 VSS.n3012 VSS.n3011 1.47372
R9175 VSS.n3007 VSS.n3006 1.47372
R9176 VSS.n2999 VSS.n2998 1.47372
R9177 VSS.n2994 VSS.n2993 1.47372
R9178 VSS.n2989 VSS.n2988 1.47372
R9179 VSS.n2984 VSS.n2983 1.47372
R9180 VSS.n2979 VSS.n2978 1.47372
R9181 VSS.n2974 VSS.n2973 1.47372
R9182 VSS.n3277 VSS.n3275 1.47359
R9183 VSS.n3274 VSS.n3272 1.47359
R9184 VSS.n3271 VSS.n3269 1.47359
R9185 VSS.n3268 VSS.n3266 1.47359
R9186 VSS.n3265 VSS.n3263 1.47359
R9187 VSS.n3262 VSS.n3260 1.47359
R9188 VSS.n3259 VSS.n3257 1.47359
R9189 VSS.n3256 VSS.n3254 1.47359
R9190 VSS.n3253 VSS.n3251 1.47359
R9191 VSS.n3250 VSS.n3248 1.47359
R9192 VSS.n3247 VSS.n3245 1.47359
R9193 VSS.n3244 VSS.n3242 1.47359
R9194 VSS.n3195 VSS.n3194 1.47359
R9195 VSS.n3200 VSS.n3199 1.47359
R9196 VSS.n3205 VSS.n3204 1.47359
R9197 VSS.n3210 VSS.n3209 1.47359
R9198 VSS.n3215 VSS.n3214 1.47359
R9199 VSS.n3220 VSS.n3219 1.47359
R9200 VSS.n3283 VSS.n3282 1.47359
R9201 VSS.n3277 VSS.n3276 1.47359
R9202 VSS.n3274 VSS.n3273 1.47359
R9203 VSS.n3271 VSS.n3270 1.47359
R9204 VSS.n3241 VSS.n3240 1.47359
R9205 VSS.n3244 VSS.n3243 1.47359
R9206 VSS.n3247 VSS.n3246 1.47359
R9207 VSS.n3250 VSS.n3249 1.47359
R9208 VSS.n3253 VSS.n3252 1.47359
R9209 VSS.n3256 VSS.n3255 1.47359
R9210 VSS.n3259 VSS.n3258 1.47359
R9211 VSS.n3262 VSS.n3261 1.47359
R9212 VSS.n3265 VSS.n3264 1.47359
R9213 VSS.n3268 VSS.n3267 1.47359
R9214 VSS.n1 VSS.t811 1.463
R9215 VSS.n1 VSS.n0 1.463
R9216 VSS.n3735 VSS.t1374 1.463
R9217 VSS.n3735 VSS.n3734 1.463
R9218 VSS.n4369 VSS.t698 1.463
R9219 VSS.n4369 VSS.n4368 1.463
R9220 VSS.n373 VSS.t106 1.463
R9221 VSS.n373 VSS.n372 1.463
R9222 VSS.n4229 VSS.t56 1.463
R9223 VSS.n4229 VSS.n4228 1.463
R9224 VSS.n4219 VSS.t951 1.463
R9225 VSS.n4219 VSS.n4218 1.463
R9226 VSS.n4222 VSS.t1448 1.463
R9227 VSS.n4222 VSS.n4221 1.463
R9228 VSS.n2870 VSS.t193 1.463
R9229 VSS.n2870 VSS.n2869 1.463
R9230 VSS.n1704 VSS.t1353 1.463
R9231 VSS.n1704 VSS.n1703 1.463
R9232 VSS.n1702 VSS.t893 1.463
R9233 VSS.n1702 VSS.n1701 1.463
R9234 VSS.n1719 VSS.t1497 1.463
R9235 VSS.n1719 VSS.n1718 1.463
R9236 VSS.n1730 VSS.t373 1.463
R9237 VSS.n1730 VSS.n1729 1.463
R9238 VSS.n4193 VSS.t508 1.463
R9239 VSS.n4193 VSS.n4192 1.463
R9240 VSS.n4191 VSS.t68 1.463
R9241 VSS.n4191 VSS.n4190 1.463
R9242 VSS.n4183 VSS.t61 1.463
R9243 VSS.n4183 VSS.n4182 1.463
R9244 VSS.n1725 VSS.t446 1.463
R9245 VSS.n1725 VSS.n1724 1.463
R9246 VSS.n777 VSS.t771 1.463
R9247 VSS.n777 VSS.n776 1.463
R9248 VSS.n4472 VSS.t271 1.463
R9249 VSS.n4472 VSS.n4471 1.463
R9250 VSS.n4547 VSS.t1079 1.463
R9251 VSS.n4547 VSS.n4546 1.463
R9252 VSS.n4534 VSS.t48 1.463
R9253 VSS.n4534 VSS.n4533 1.463
R9254 VSS.n4528 VSS.t1264 1.463
R9255 VSS.n4528 VSS.n4527 1.463
R9256 VSS.n2477 VSS.t687 1.463
R9257 VSS.n2477 VSS.n2476 1.463
R9258 VSS.n2490 VSS.t181 1.463
R9259 VSS.n2490 VSS.n2489 1.463
R9260 VSS.n240 VSS.t1190 1.463
R9261 VSS.n240 VSS.n239 1.463
R9262 VSS.n262 VSS.t403 1.463
R9263 VSS.n262 VSS.n261 1.463
R9264 VSS.n259 VSS.t197 1.463
R9265 VSS.n259 VSS.n258 1.463
R9266 VSS.n5108 VSS.t712 1.463
R9267 VSS.n5108 VSS.n5107 1.463
R9268 VSS.n292 VSS.t239 1.463
R9269 VSS.n292 VSS.n291 1.463
R9270 VSS.n281 VSS.t450 1.463
R9271 VSS.n281 VSS.n280 1.463
R9272 VSS.n2472 VSS.t456 1.463
R9273 VSS.n2472 VSS.n2471 1.463
R9274 VSS.n2464 VSS.t1405 1.463
R9275 VSS.n2464 VSS.n2463 1.463
R9276 VSS.n81 VSS.t702 1.463
R9277 VSS.n81 VSS.n80 1.463
R9278 VSS.n39 VSS.t39 1.463
R9279 VSS.n39 VSS.n38 1.463
R9280 VSS.n45 VSS.t496 1.463
R9281 VSS.n45 VSS.n44 1.463
R9282 VSS.n50 VSS.t866 1.463
R9283 VSS.n50 VSS.n49 1.463
R9284 VSS.n75 VSS.t676 1.463
R9285 VSS.n75 VSS.n74 1.463
R9286 VSS.n147 VSS.t204 1.463
R9287 VSS.n147 VSS.n146 1.463
R9288 VSS.n130 VSS.t199 1.463
R9289 VSS.n130 VSS.n129 1.463
R9290 VSS.n150 VSS.t183 1.463
R9291 VSS.n150 VSS.n149 1.463
R9292 VSS.n168 VSS.t399 1.463
R9293 VSS.n168 VSS.n167 1.463
R9294 VSS.n68 VSS.t46 1.463
R9295 VSS.n68 VSS.n67 1.463
R9296 VSS.n65 VSS.t517 1.463
R9297 VSS.n65 VSS.n64 1.463
R9298 VSS.n2860 VSS.t1346 1.463
R9299 VSS.n2860 VSS.n2859 1.463
R9300 VSS.n2895 VSS.t607 1.463
R9301 VSS.n2895 VSS.n2894 1.463
R9302 VSS.n2905 VSS.t908 1.463
R9303 VSS.n2905 VSS.n2904 1.463
R9304 VSS.n542 VSS.t1074 1.463
R9305 VSS.n542 VSS.n541 1.463
R9306 VSS.n535 VSS.t976 1.463
R9307 VSS.n535 VSS.n534 1.463
R9308 VSS.n539 VSS.t622 1.463
R9309 VSS.n539 VSS.n538 1.463
R9310 VSS.n4558 VSS.t318 1.463
R9311 VSS.n4558 VSS.n4557 1.463
R9312 VSS.n525 VSS.t1072 1.463
R9313 VSS.n525 VSS.n524 1.463
R9314 VSS.n522 VSS.t1070 1.463
R9315 VSS.n522 VSS.n521 1.463
R9316 VSS.n556 VSS.t631 1.463
R9317 VSS.n556 VSS.n555 1.463
R9318 VSS.n4524 VSS.t540 1.463
R9319 VSS.n4524 VSS.n4523 1.463
R9320 VSS.n748 VSS.t1136 1.463
R9321 VSS.n748 VSS.n747 1.463
R9322 VSS.n4517 VSS.t292 1.463
R9323 VSS.n4517 VSS.n4516 1.463
R9324 VSS.n4494 VSS.t323 1.463
R9325 VSS.n4494 VSS.n4493 1.463
R9326 VSS.n4501 VSS.t209 1.463
R9327 VSS.n4501 VSS.n4500 1.463
R9328 VSS.n4503 VSS.t1164 1.463
R9329 VSS.n4503 VSS.n4502 1.463
R9330 VSS.n772 VSS.t366 1.463
R9331 VSS.n772 VSS.n771 1.463
R9332 VSS.n768 VSS.t473 1.463
R9333 VSS.n768 VSS.n767 1.463
R9334 VSS.n766 VSS.t464 1.463
R9335 VSS.n766 VSS.n765 1.463
R9336 VSS.n762 VSS.t358 1.463
R9337 VSS.n762 VSS.n761 1.463
R9338 VSS.n999 VSS.t485 1.463
R9339 VSS.n999 VSS.n998 1.463
R9340 VSS.n1001 VSS.t1099 1.463
R9341 VSS.n1001 VSS.n1000 1.463
R9342 VSS.n1013 VSS.t775 1.463
R9343 VSS.n1013 VSS.n1012 1.463
R9344 VSS.n1018 VSS.t781 1.463
R9345 VSS.n1018 VSS.n1017 1.463
R9346 VSS.n1009 VSS.t1197 1.463
R9347 VSS.n1009 VSS.n1008 1.463
R9348 VSS.n1004 VSS.t620 1.463
R9349 VSS.n1004 VSS.n1003 1.463
R9350 VSS.n1022 VSS.t766 1.463
R9351 VSS.n1022 VSS.n1021 1.463
R9352 VSS.n4414 VSS.t1303 1.463
R9353 VSS.n4414 VSS.n4413 1.463
R9354 VSS.n1032 VSS.t749 1.463
R9355 VSS.n1032 VSS.n1031 1.463
R9356 VSS.n1028 VSS.t809 1.463
R9357 VSS.n1028 VSS.n1027 1.463
R9358 VSS.n1066 VSS.t265 1.463
R9359 VSS.n1066 VSS.n1065 1.463
R9360 VSS.n1063 VSS.t1308 1.463
R9361 VSS.n1063 VSS.n1062 1.463
R9362 VSS.n1068 VSS.t1019 1.463
R9363 VSS.n1068 VSS.n1067 1.463
R9364 VSS.n4206 VSS.t501 1.463
R9365 VSS.n4206 VSS.n4205 1.463
R9366 VSS.n4197 VSS.t934 1.463
R9367 VSS.n4197 VSS.n4196 1.463
R9368 VSS.n1038 VSS.t451 1.463
R9369 VSS.n1038 VSS.n1037 1.463
R9370 VSS.n1041 VSS.t765 1.463
R9371 VSS.n1041 VSS.n1040 1.463
R9372 VSS.n1060 VSS.t792 1.463
R9373 VSS.n1060 VSS.n1059 1.463
R9374 VSS.n4380 VSS.t151 1.463
R9375 VSS.n4380 VSS.n4379 1.463
R9376 VSS.n1035 VSS.t325 1.463
R9377 VSS.n1035 VSS.n1034 1.463
R9378 VSS.n1025 VSS.t559 1.463
R9379 VSS.n1025 VSS.n1024 1.463
R9380 VSS.n4402 VSS.t557 1.463
R9381 VSS.n4402 VSS.n4401 1.463
R9382 VSS.n752 VSS.t1065 1.463
R9383 VSS.n752 VSS.n751 1.463
R9384 VSS.n4492 VSS.t1135 1.463
R9385 VSS.n4492 VSS.n4491 1.463
R9386 VSS.n4485 VSS.t277 1.463
R9387 VSS.n4485 VSS.n4484 1.463
R9388 VSS.n757 VSS.t1111 1.463
R9389 VSS.n757 VSS.n756 1.463
R9390 VSS.n783 VSS.t153 1.463
R9391 VSS.n783 VSS.n782 1.463
R9392 VSS.n781 VSS.t179 1.463
R9393 VSS.n781 VSS.n780 1.463
R9394 VSS.n311 VSS.t945 1.463
R9395 VSS.n311 VSS.n310 1.463
R9396 VSS.n325 VSS.t168 1.463
R9397 VSS.n325 VSS.n324 1.463
R9398 VSS.n4262 VSS.t873 1.463
R9399 VSS.n4262 VSS.n4261 1.463
R9400 VSS.n4266 VSS.t913 1.463
R9401 VSS.n4266 VSS.n4265 1.463
R9402 VSS.n4252 VSS.t844 1.463
R9403 VSS.n4252 VSS.n4251 1.463
R9404 VSS.n4260 VSS.t138 1.463
R9405 VSS.n4260 VSS.n4259 1.463
R9406 VSS.n4216 VSS.t936 1.463
R9407 VSS.n4216 VSS.n4215 1.463
R9408 VSS.n4247 VSS.t900 1.463
R9409 VSS.n4247 VSS.n4246 1.463
R9410 VSS.n4249 VSS.t569 1.463
R9411 VSS.n4249 VSS.n4248 1.463
R9412 VSS.n315 VSS.t244 1.463
R9413 VSS.n315 VSS.n314 1.463
R9414 VSS.n309 VSS.t1519 1.463
R9415 VSS.n309 VSS.n308 1.463
R9416 VSS.n307 VSS.t1029 1.463
R9417 VSS.n307 VSS.n306 1.463
R9418 VSS.n320 VSS.t513 1.463
R9419 VSS.n320 VSS.n319 1.463
R9420 VSS.n343 VSS.t1432 1.463
R9421 VSS.n343 VSS.n342 1.463
R9422 VSS.n353 VSS.t466 1.463
R9423 VSS.n353 VSS.n352 1.463
R9424 VSS.n355 VSS.t1438 1.463
R9425 VSS.n355 VSS.n354 1.463
R9426 VSS.n4972 VSS.t443 1.463
R9427 VSS.n4972 VSS.n4971 1.463
R9428 VSS.n338 VSS.t1068 1.463
R9429 VSS.n338 VSS.n337 1.463
R9430 VSS.n340 VSS.t1545 1.463
R9431 VSS.n340 VSS.n339 1.463
R9432 VSS.n335 VSS.t214 1.463
R9433 VSS.n335 VSS.n334 1.463
R9434 VSS.n317 VSS.t825 1.463
R9435 VSS.n317 VSS.n316 1.463
R9436 VSS.n4280 VSS.t272 1.463
R9437 VSS.n4280 VSS.n4279 1.463
R9438 VSS.n4284 VSS.t178 1.463
R9439 VSS.n4284 VSS.n4283 1.463
R9440 VSS.n2485 VSS.t223 1.463
R9441 VSS.n2485 VSS.n2484 1.463
R9442 VSS.n1700 VSS.t965 1.463
R9443 VSS.n1700 VSS.n1699 1.463
R9444 VSS.n1714 VSS.t1315 1.463
R9445 VSS.n1714 VSS.n1713 1.463
R9446 VSS.n2866 VSS.t684 1.463
R9447 VSS.n2866 VSS.n2865 1.463
R9448 VSS.n2878 VSS.t970 1.463
R9449 VSS.n2878 VSS.n2877 1.463
R9450 VSS.n2873 VSS.t1329 1.463
R9451 VSS.n2873 VSS.n2872 1.463
R9452 VSS.n2888 VSS.t7 1.463
R9453 VSS.n2888 VSS.n2887 1.463
R9454 VSS.n2855 VSS.t1289 1.463
R9455 VSS.n2855 VSS.n2854 1.463
R9456 VSS.n1739 VSS.t53 1.463
R9457 VSS.n1739 VSS.n1738 1.463
R9458 VSS.n1745 VSS.t1460 1.463
R9459 VSS.n1745 VSS.n1744 1.463
R9460 VSS.n1742 VSS.t337 1.463
R9461 VSS.n1742 VSS.n1741 1.463
R9462 VSS.n4203 VSS.t1282 1.463
R9463 VSS.n4203 VSS.n4202 1.463
R9464 VSS.n4213 VSS.t626 1.463
R9465 VSS.n4213 VSS.n4212 1.463
R9466 VSS.n4210 VSS.t1411 1.463
R9467 VSS.n4210 VSS.n4209 1.463
R9468 VSS.n370 VSS.t184 1.463
R9469 VSS.n370 VSS.n369 1.463
R9470 VSS.n529 VSS.t1546 1.463
R9471 VSS.n529 VSS.n528 1.463
R9472 VSS.n377 VSS.t1430 1.463
R9473 VSS.n377 VSS.n376 1.463
R9474 VSS.n4363 VSS.t1348 1.463
R9475 VSS.n4363 VSS.n4362 1.463
R9476 VSS.n1077 VSS.t415 1.463
R9477 VSS.n1077 VSS.n1076 1.463
R9478 VSS.n1082 VSS.t1023 1.463
R9479 VSS.n1082 VSS.n1081 1.463
R9480 VSS.n1312 VSS.t14 1.463
R9481 VSS.n1312 VSS.n1311 1.463
R9482 VSS.n1310 VSS.t1227 1.463
R9483 VSS.n1310 VSS.n1309 1.463
R9484 VSS.n1308 VSS.t740 1.463
R9485 VSS.n1308 VSS.n1307 1.463
R9486 VSS.n1320 VSS.t1239 1.463
R9487 VSS.n1320 VSS.n1319 1.463
R9488 VSS.n1305 VSS.t731 1.463
R9489 VSS.n1305 VSS.n1304 1.463
R9490 VSS.n1327 VSS.t1225 1.463
R9491 VSS.n1327 VSS.n1326 1.463
R9492 VSS.n2292 VSS.t886 1.463
R9493 VSS.n2292 VSS.n2291 1.463
R9494 VSS.n3450 VSS.t34 1.463
R9495 VSS.n3450 VSS.n3449 1.463
R9496 VSS.n2605 VSS.t1249 1.463
R9497 VSS.n2605 VSS.n2604 1.463
R9498 VSS.n5104 VSS.n5103 1.45973
R9499 VSS.n179 VSS.n178 1.45973
R9500 VSS.n89 VSS 1.4209
R9501 VSS.n2500 VSS 1.4209
R9502 VSS.n4432 VSS.n4431 1.41164
R9503 VSS.n4428 VSS.n4427 1.41164
R9504 VSS.n4239 VSS.n4214 1.41164
R9505 VSS.n4242 VSS.n4241 1.41164
R9506 VSS.n3732 VSS.n3731 1.39845
R9507 VSS.n3727 VSS.n3726 1.39845
R9508 VSS.n2624 VSS.n2623 1.38035
R9509 VSS.n204 VSS 1.34435
R9510 VSS VSS.n2487 1.34435
R9511 VSS.n5101 VSS 1.34261
R9512 VSS.n5061 VSS 1.34261
R9513 VSS.n176 VSS 1.34261
R9514 VSS.n121 VSS 1.34261
R9515 VSS.n5065 VSS.n5064 1.32493
R9516 VSS.n5414 VSS.n5413 1.32493
R9517 VSS.n5092 VSS.n5091 1.315
R9518 VSS.n5396 VSS.n5395 1.315
R9519 VSS.n4552 VSS.n4548 1.30108
R9520 VSS.n4434 VSS.n4433 1.30108
R9521 VSS.n4426 VSS.n1023 1.30108
R9522 VSS.n4301 VSS.n4300 1.30108
R9523 VSS.n4295 VSS.n4294 1.30108
R9524 VSS.n2881 VSS.n2880 1.30108
R9525 VSS.n4235 VSS.n4220 1.29958
R9526 VSS.n544 VSS.n543 1.29958
R9527 VSS.n4564 VSS.n523 1.29958
R9528 VSS.n4438 VSS.n4437 1.29958
R9529 VSS.n4421 VSS.n4420 1.29958
R9530 VSS.n4271 VSS.n4270 1.29958
R9531 VSS.n5139 VSS.n5138 1.27516
R9532 VSS.n249 VSS.n248 1.26641
R9533 VSS.n5050 VSS.n5049 1.26641
R9534 VSS.n209 VSS.n208 1.26641
R9535 VSS.n158 VSS.n157 1.26641
R9536 VSS.n5420 VSS.n5419 1.26641
R9537 VSS.n229 VSS.n228 1.26641
R9538 VSS.n5007 VSS.n5006 1.26641
R9539 VSS.n4349 VSS.n4348 1.26524
R9540 VSS.n4980 VSS.n4979 1.25337
R9541 VSS.n1301 VSS.n1140 1.25097
R9542 VSS.n5116 VSS 1.24292
R9543 VSS VSS.n5098 1.24292
R9544 VSS.n5038 VSS 1.24292
R9545 VSS VSS.n66 1.24292
R9546 VSS VSS.n5447 1.24292
R9547 VSS.n192 VSS 1.24292
R9548 VSS VSS.n5402 1.24292
R9549 VSS.n4861 VSS.n4860 1.23073
R9550 VSS.n5372 VSS.n5371 1.23073
R9551 VSS.n5077 VSS.n5076 1.22108
R9552 VSS.n238 VSS.n237 1.22108
R9553 VSS.n290 VSS.n289 1.22108
R9554 VSS.n110 VSS.n109 1.22108
R9555 VSS.n59 VSS.n58 1.22108
R9556 VSS.n137 VSS.n136 1.22108
R9557 VSS.n191 VSS.n190 1.22108
R9558 VSS.n3464 VSS.t431 1.20928
R9559 VSS.n4346 VSS.n4345 1.20218
R9560 VSS.n5473 VSS.n5472 1.19064
R9561 VSS.n4116 VSS.n4110 1.18807
R9562 VSS.n4176 VSS.n4175 1.18142
R9563 VSS.n3543 VSS.n3542 1.17635
R9564 VSS.n1689 VSS.n1688 1.1727
R9565 VSS.n3981 VSS.n3980 1.17251
R9566 VSS.n5142 VSS.n5141 1.171
R9567 VSS.n5206 VSS.n5204 1.16717
R9568 VSS.n3992 VSS.n3991 1.16534
R9569 VSS.n5002 VSS.n5001 1.15749
R9570 VSS.n1760 VSS.n1759 1.14506
R9571 VSS.n2589 VSS.n2535 1.12164
R9572 VSS.n2481 VSS.n2480 1.11939
R9573 VSS.n85 VSS.n84 1.11939
R9574 VSS.t782 VSS.n4395 1.11772
R9575 VSS.n4459 VSS.t770 1.11772
R9576 VSS.n4520 VSS.t1076 1.11772
R9577 VSS.t944 VSS.n4996 1.11772
R9578 VSS.t964 VSS.n1698 1.11772
R9579 VSS.n4312 VSS.t904 1.11772
R9580 VSS.n5001 VSS.n298 1.08721
R9581 VSS.n5206 VSS.n5202 1.07742
R9582 VSS.t1083 VSS.n4566 1.03818
R9583 VSS.n4417 VSS.t753 1.03818
R9584 VSS.n4435 VSS.t774 1.03818
R9585 VSS.t907 VSS.n2926 1.03818
R9586 VSS.t948 VSS.n4238 1.03818
R9587 VSS.n4245 VSS.t899 1.03818
R9588 VSS.n4955 VSS.t1086 1.03818
R9589 VSS.n3539 VSS.n1694 1.03581
R9590 VSS.n2913 VSS.n2912 1.03184
R9591 VSS.n545 VSS.n544 1.03184
R9592 VSS.n4433 VSS.n1005 1.03184
R9593 VSS.n4426 VSS.n4425 1.03184
R9594 VSS.n4302 VSS.n4301 1.03184
R9595 VSS.n4294 VSS.n4293 1.03184
R9596 VSS.n4237 VSS.n4236 1.01411
R9597 VSS.n552 VSS.n551 1.01411
R9598 VSS.n4551 VSS.n4550 1.01411
R9599 VSS.n1015 VSS.n1011 1.01411
R9600 VSS.n4418 VSS.n1030 1.01411
R9601 VSS.n4268 VSS.n4264 1.01411
R9602 VSS.n2876 VSS.n2875 1.01411
R9603 VSS.n4564 VSS.n4563 1.0114
R9604 VSS.n5138 VSS.n224 0.983736
R9605 VSS.n4561 VSS.n224 0.976784
R9606 VSS.n4348 VSS.n1139 0.936031
R9607 VSS.n4235 VSS 0.935416
R9608 VSS.n550 VSS 0.935416
R9609 VSS VSS.n4552 0.935416
R9610 VSS VSS.n4438 0.935416
R9611 VSS VSS.n4421 0.935416
R9612 VSS VSS.n4271 0.935416
R9613 VSS VSS.n2881 0.935416
R9614 VSS.n5002 VSS.n55 0.932808
R9615 VSS.n544 VSS.n540 0.92521
R9616 VSS.n4565 VSS.n4564 0.92521
R9617 VSS.n4816 VSS.n4815 0.914514
R9618 VSS.n5327 VSS.n5326 0.914514
R9619 VSS.n5500 VSS.t793 0.909591
R9620 VSS.n2520 VSS.n2519 0.881611
R9621 VSS.n5468 VSS.n5467 0.881611
R9622 VSS.n2575 VSS.n2572 0.881611
R9623 VSS.n2945 VSS.n2944 0.881611
R9624 VSS.n1126 VSS.n1123 0.881611
R9625 VSS.n4042 VSS.n2591 0.881611
R9626 VSS.n4146 VSS.n4145 0.880263
R9627 VSS.n4474 VSS.n4473 0.87647
R9628 VSS.n331 VSS.n330 0.87647
R9629 VSS.n1736 VSS.n1735 0.876262
R9630 VSS.n4371 VSS.n4370 0.87613
R9631 VSS.n4329 VSS.n4328 0.875129
R9632 VSS.n3452 VSS.n3451 0.875129
R9633 VSS.n4487 VSS.n4486 0.874923
R9634 VSS.n4977 VSS.n4976 0.874923
R9635 VSS.n2510 VSS.n2509 0.874807
R9636 VSS.n5456 VSS.n5455 0.874807
R9637 VSS.n5137 VSS 0.86396
R9638 VSS.n4007 VSS.n4006 0.845198
R9639 VSS.n4180 VSS.n1746 0.839031
R9640 VSS VSS.n2457 0.803833
R9641 VSS VSS.n2518 0.803833
R9642 VSS VSS.n28 0.803833
R9643 VSS VSS.n5466 0.803833
R9644 VSS VSS.n2578 0.803833
R9645 VSS VSS.n2574 0.803833
R9646 VSS VSS.n2849 0.803833
R9647 VSS VSS.n2943 0.803833
R9648 VSS VSS.n1129 0.803833
R9649 VSS VSS.n1125 0.803833
R9650 VSS.n4039 VSS 0.803833
R9651 VSS.n4432 VSS.n1016 0.803577
R9652 VSS.n4427 VSS.n1020 0.803577
R9653 VSS.n4299 VSS.n4214 0.803577
R9654 VSS.n4296 VSS.n4242 0.803577
R9655 VSS.n3726 VSS.n3725 0.802703
R9656 VSS.n2911 VSS.n2910 0.802588
R9657 VSS.n4236 VSS.n4217 0.788242
R9658 VSS.n551 VSS.n527 0.788242
R9659 VSS.n4551 VSS.n4549 0.788242
R9660 VSS.n4436 VSS.n1011 0.788242
R9661 VSS.n4419 VSS.n1030 0.788242
R9662 VSS.n4269 VSS.n4264 0.788242
R9663 VSS.n2879 VSS.n2876 0.788242
R9664 VSS.n2500 VSS.n2493 0.777239
R9665 VSS.n89 VSS.n78 0.777239
R9666 VSS.n4349 VSS.n1085 0.777239
R9667 VSS.n5026 VSS 0.77007
R9668 VSS.n92 VSS 0.77007
R9669 VSS.n2455 VSS.n2454 0.71601
R9670 VSS.n26 VSS.n25 0.71601
R9671 VSS.n2567 VSS.n2537 0.71601
R9672 VSS.n2847 VSS.n2846 0.71601
R9673 VSS.n1118 VSS.n1088 0.71601
R9674 VSS.n4038 VSS.n4037 0.71601
R9675 VSS.n4189 VSS.n4186 0.6745
R9676 VSS.n1317 VSS.n1316 0.671611
R9677 VSS.n4346 VSS.n1693 0.662178
R9678 VSS.n988 VSS.n987 0.656724
R9679 VSS.n2480 VSS.n2478 0.656358
R9680 VSS.n2493 VSS.n2491 0.656358
R9681 VSS.n84 VSS.n82 0.656358
R9682 VSS.n78 VSS.n76 0.656358
R9683 VSS.n1085 VSS.n1083 0.656358
R9684 VSS.n1768 VSS.n1764 0.628705
R9685 VSS.n5064 VSS.n5063 0.597038
R9686 VSS.n5415 VSS.n5414 0.597038
R9687 VSS.n4393 VSS.n4392 0.590319
R9688 VSS.n1058 VSS.n1057 0.584346
R9689 VSS VSS.n5478 0.582722
R9690 VSS VSS.n2543 0.582722
R9691 VSS VSS.n2598 0.582722
R9692 VSS VSS.n2952 0.582722
R9693 VSS VSS.n2527 0.582722
R9694 VSS VSS.n1094 0.582722
R9695 VSS.n4454 VSS.n4453 0.574328
R9696 VSS.n4286 VSS.n4285 0.574328
R9697 VSS.n2919 VSS.n2918 0.573536
R9698 VSS.n994 VSS.n993 0.573536
R9699 VSS.n4282 VSS.n4281 0.573536
R9700 VSS.n2920 VSS.n2867 0.573328
R9701 VSS.n4539 VSS.n4535 0.572195
R9702 VSS.n4407 VSS.n4399 0.572195
R9703 VSS.n4307 VSS.n4207 0.572195
R9704 VSS.n4962 VSS.n374 0.572195
R9705 VSS.n4541 VSS.n4540 0.571989
R9706 VSS.n4408 VSS.n1036 0.571989
R9707 VSS.n4309 VSS.n4308 0.571989
R9708 VSS.n4964 VSS.n4963 0.571989
R9709 VSS.n2501 VSS.n2500 0.568021
R9710 VSS.n91 VSS.n89 0.568021
R9711 VSS.n4353 VSS.n4349 0.568021
R9712 VSS.n3005 VSS.n3003 0.564944
R9713 VSS.n3005 VSS.n3004 0.564944
R9714 VSS.n3006 VSS.n3005 0.564944
R9715 VSS.n3022 VSS.n3021 0.564944
R9716 VSS.n3092 VSS.n3085 0.564944
R9717 VSS.n3092 VSS.n3086 0.564944
R9718 VSS.n3092 VSS.n3087 0.564944
R9719 VSS.n3092 VSS.n3088 0.564944
R9720 VSS.n3092 VSS.n3089 0.564944
R9721 VSS.n3092 VSS.n3090 0.564944
R9722 VSS.n3092 VSS.n3091 0.564944
R9723 VSS.n3093 VSS.n3092 0.564944
R9724 VSS.n3281 VSS.n3280 0.564944
R9725 VSS.n3281 VSS.n3277 0.564705
R9726 VSS.n3281 VSS.n3274 0.564705
R9727 VSS.n3281 VSS.n3271 0.564705
R9728 VSS.n3281 VSS.n3224 0.564705
R9729 VSS.n3281 VSS.n3225 0.564705
R9730 VSS.n3281 VSS.n3226 0.564705
R9731 VSS.n3281 VSS.n3227 0.564705
R9732 VSS.n3281 VSS.n3228 0.564705
R9733 VSS.n3281 VSS.n3229 0.564705
R9734 VSS.n3281 VSS.n3230 0.564705
R9735 VSS.n3281 VSS.n3231 0.564705
R9736 VSS.n3281 VSS.n3232 0.564705
R9737 VSS.n3281 VSS.n3233 0.564705
R9738 VSS.n3281 VSS.n3234 0.564705
R9739 VSS.n3281 VSS.n3235 0.564705
R9740 VSS.n3281 VSS.n3236 0.564705
R9741 VSS.n3281 VSS.n3237 0.564705
R9742 VSS.n3281 VSS.n3238 0.564705
R9743 VSS.n3281 VSS.n3239 0.564705
R9744 VSS.n3281 VSS.n3241 0.564705
R9745 VSS.n3281 VSS.n3244 0.564705
R9746 VSS.n3281 VSS.n3247 0.564705
R9747 VSS.n3281 VSS.n3250 0.564705
R9748 VSS.n3281 VSS.n3253 0.564705
R9749 VSS.n3281 VSS.n3256 0.564705
R9750 VSS.n3281 VSS.n3259 0.564705
R9751 VSS.n3281 VSS.n3262 0.564705
R9752 VSS.n3281 VSS.n3265 0.564705
R9753 VSS.n3281 VSS.n3268 0.564705
R9754 VSS.n3282 VSS.n3281 0.564705
R9755 VSS.n4147 VSS.n4146 0.561269
R9756 VSS.n4953 VSS.n4952 0.555337
R9757 VSS.n4889 VSS.n4888 0.555337
R9758 VSS.n4763 VSS.n4762 0.555337
R9759 VSS.n5279 VSS.n5278 0.555337
R9760 VSS.n4953 VSS.n4951 0.555098
R9761 VSS.n4953 VSS.n4950 0.555098
R9762 VSS.n4953 VSS.n4949 0.555098
R9763 VSS.n4953 VSS.n4948 0.555098
R9764 VSS.n4953 VSS.n4947 0.555098
R9765 VSS.n4953 VSS.n4946 0.555098
R9766 VSS.n4953 VSS.n4945 0.555098
R9767 VSS.n4953 VSS.n4944 0.555098
R9768 VSS.n4953 VSS.n4943 0.555098
R9769 VSS.n4816 VSS.n4814 0.555098
R9770 VSS.n4816 VSS.n4813 0.555098
R9771 VSS.n4817 VSS.n4816 0.555098
R9772 VSS.n4803 VSS.n4802 0.555098
R9773 VSS.n5327 VSS.n5325 0.555098
R9774 VSS.n5327 VSS.n5324 0.555098
R9775 VSS.n5328 VSS.n5327 0.555098
R9776 VSS.n5314 VSS.n5313 0.555098
R9777 VSS.n4198 VSS.n4181 0.554405
R9778 VSS.n5084 VSS.n241 0.50331
R9779 VSS.n5071 VSS.n5070 0.50331
R9780 VSS.n273 VSS.n260 0.50331
R9781 VSS.n5110 VSS.n5109 0.50331
R9782 VSS.n294 VSS.n293 0.50331
R9783 VSS.n5033 VSS.n282 0.50331
R9784 VSS.n5450 VSS.n5448 0.50331
R9785 VSS.n148 VSS.n144 0.50331
R9786 VSS.n5404 VSS.n5403 0.50331
R9787 VSS.n183 VSS.n182 0.50331
R9788 VSS.n174 VSS.n173 0.50331
R9789 VSS.n102 VSS.n101 0.50331
R9790 VSS.n5432 VSS.n5431 0.50331
R9791 VSS.n2486 VSS.n2482 0.50331
R9792 VSS.n4148 VSS.n4147 0.499494
R9793 VSS.n5486 VSS.n5485 0.487216
R9794 VSS.n2549 VSS.n2548 0.487216
R9795 VSS.n2826 VSS.n2825 0.487216
R9796 VSS.n1100 VSS.n1099 0.487216
R9797 VSS.n1316 VSS.n1315 0.4805
R9798 VSS.n1318 VSS.n1317 0.4805
R9799 VSS.n1321 VSS.n1306 0.4805
R9800 VSS.n1325 VSS.n1324 0.4805
R9801 VSS.n5137 VSS.n5136 0.480148
R9802 VSS.n4116 VSS.n4115 0.475159
R9803 VSS.n4143 VSS.n4142 0.475159
R9804 VSS.n2391 VSS.n2390 0.475159
R9805 VSS.n1754 VSS.n55 0.465605
R9806 VSS.n5477 VSS 0.457167
R9807 VSS VSS.n2559 0.457167
R9808 VSS VSS.n4025 0.457167
R9809 VSS VSS.n2832 0.457167
R9810 VSS VSS.n2440 0.457167
R9811 VSS VSS.n1110 0.457167
R9812 VSS.n2434 VSS.n2430 0.454994
R9813 VSS.n2912 VSS.n2911 0.4505
R9814 VSS.n4433 VSS.n4432 0.4505
R9815 VSS.n4427 VSS.n4426 0.4505
R9816 VSS.n4301 VSS.n4214 0.4505
R9817 VSS.n4294 VSS.n4242 0.4505
R9818 VSS.n5195 VSS.n5193 0.449218
R9819 VSS.n5218 VSS.n5214 0.449218
R9820 VSS.n5121 VSS.n233 0.445885
R9821 VSS.n5043 VSS.n285 0.445885
R9822 VSS.n115 VSS.n105 0.445885
R9823 VSS.n197 VSS.n186 0.445885
R9824 VSS.n5092 VSS.n5083 0.441269
R9825 VSS.n5396 VSS.n143 0.441269
R9826 VSS.n3969 VSS.n3921 0.439329
R9827 VSS.n1324 VSS 0.434944
R9828 VSS.n3969 VSS.n3924 0.431816
R9829 VSS.n3969 VSS.n3927 0.431816
R9830 VSS.n3969 VSS.n3930 0.431816
R9831 VSS.n3969 VSS.n3933 0.431816
R9832 VSS.n3969 VSS.n3936 0.431816
R9833 VSS.n3969 VSS.n3939 0.431816
R9834 VSS.n3969 VSS.n3942 0.431816
R9835 VSS.n3969 VSS.n3945 0.431816
R9836 VSS.n3969 VSS.n3948 0.431816
R9837 VSS.n3969 VSS.n3951 0.431816
R9838 VSS.n3969 VSS.n3954 0.431816
R9839 VSS.n3969 VSS.n3956 0.431816
R9840 VSS.n3969 VSS.n3957 0.431816
R9841 VSS.n3969 VSS.n3958 0.431816
R9842 VSS.n3969 VSS.n3959 0.431816
R9843 VSS.n3969 VSS.n3960 0.431816
R9844 VSS.n3969 VSS.n3961 0.431816
R9845 VSS.n3969 VSS.n3962 0.431816
R9846 VSS.n3969 VSS.n3963 0.431816
R9847 VSS.n3969 VSS.n3964 0.431816
R9848 VSS.n3969 VSS.n3965 0.431816
R9849 VSS.n3969 VSS.n3966 0.431816
R9850 VSS.n3969 VSS.n3967 0.431816
R9851 VSS.n3969 VSS.n3968 0.431816
R9852 VSS.n3970 VSS.n3969 0.431816
R9853 VSS.n1680 VSS.n1679 0.431816
R9854 VSS.n1679 VSS.n1369 0.431816
R9855 VSS.n1679 VSS.n1374 0.431816
R9856 VSS.n1679 VSS.n1379 0.431816
R9857 VSS.n1679 VSS.n1384 0.431816
R9858 VSS.n1679 VSS.n1678 0.431816
R9859 VSS.n1646 VSS.n1645 0.431816
R9860 VSS.n1645 VSS.n1644 0.431816
R9861 VSS.n419 VSS.n418 0.431816
R9862 VSS.n4146 VSS.n2293 0.413044
R9863 VSS.n5457 VSS 0.406011
R9864 VSS.n5120 VSS.n234 0.4055
R9865 VSS.n5096 VSS.n5095 0.4055
R9866 VSS.n5102 VSS.n257 0.4055
R9867 VSS.n5042 VSS.n286 0.4055
R9868 VSS.n5062 VSS.n279 0.4055
R9869 VSS.n114 VSS.n106 0.4055
R9870 VSS.n5445 VSS.n54 0.4055
R9871 VSS.n196 VSS.n187 0.4055
R9872 VSS.n5400 VSS.n5399 0.4055
R9873 VSS.n211 VSS.n205 0.4055
R9874 VSS.n177 VSS.n166 0.4055
R9875 VSS.n5422 VSS.n5416 0.4055
R9876 VSS.n5135 VSS.n5133 0.4055
R9877 VSS.n212 VSS.n203 0.403192
R9878 VSS.n5118 VSS.n5117 0.400885
R9879 VSS.n5093 VSS.n5073 0.400885
R9880 VSS.n5097 VSS.n5072 0.400885
R9881 VSS.n5040 VSS.n5039 0.400885
R9882 VSS.n112 VSS.n111 0.400885
R9883 VSS.n5446 VSS.n52 0.400885
R9884 VSS.n194 VSS.n193 0.400885
R9885 VSS.n5397 VSS.n133 0.400885
R9886 VSS.n5401 VSS.n132 0.400885
R9887 VSS.n4015 VSS.n4014 0.398328
R9888 VSS.n2511 VSS 0.395857
R9889 VSS.n5459 VSS 0.394786
R9890 VSS.n5103 VSS.n5102 0.388192
R9891 VSS.n5063 VSS.n5062 0.388192
R9892 VSS.n178 VSS.n177 0.388192
R9893 VSS.n5416 VSS.n5415 0.388192
R9894 VSS VSS.n2515 0.387167
R9895 VSS VSS.n5463 0.387167
R9896 VSS VSS.n2584 0.387167
R9897 VSS VSS.n1135 0.387167
R9898 VSS.n4103 VSS 0.387167
R9899 VSS.n4385 VSS.n1069 0.3805
R9900 VSS.n5068 VSS.n5067 0.37418
R9901 VSS.n5411 VSS.n5409 0.37418
R9902 VSS.n4149 VSS.n4148 0.367956
R9903 VSS.n1315 VSS 0.364944
R9904 VSS VSS.n1321 0.364944
R9905 VSS VSS.n1329 0.364944
R9906 VSS.n4560 VSS.n745 0.362755
R9907 VSS.n1329 VSS.n1328 0.362722
R9908 VSS.n5443 VSS.n5442 0.352423
R9909 VSS VSS.n2608 0.347643
R9910 VSS.n4230 VSS 0.347643
R9911 VSS VSS.n4231 0.347643
R9912 VSS.n1733 VSS 0.347643
R9913 VSS.n4529 VSS 0.347643
R9914 VSS VSS.n2923 0.347643
R9915 VSS VSS.n2861 0.347643
R9916 VSS.n536 VSS 0.347643
R9917 VSS VSS.n537 0.347643
R9918 VSS VSS.n746 0.347643
R9919 VSS.n4530 VSS 0.347643
R9920 VSS VSS.n749 0.347643
R9921 VSS VSS.n4515 0.347643
R9922 VSS.n4476 VSS 0.347643
R9923 VSS.n4450 VSS 0.347643
R9924 VSS.n4449 VSS 0.347643
R9925 VSS.n4446 VSS 0.347643
R9926 VSS VSS.n4447 0.347643
R9927 VSS VSS.n4412 0.347643
R9928 VSS.n4411 VSS 0.347643
R9929 VSS.n4377 VSS 0.347643
R9930 VSS VSS.n4378 0.347643
R9931 VSS VSS.n1026 0.347643
R9932 VSS.n4404 VSS 0.347643
R9933 VSS.n4514 VSS 0.347643
R9934 VSS VSS.n4477 0.347643
R9935 VSS.n328 VSS 0.347643
R9936 VSS VSS.n4254 0.347643
R9937 VSS VSS.n4291 0.347643
R9938 VSS.n4276 VSS 0.347643
R9939 VSS VSS.n4250 0.347643
R9940 VSS.n4973 VSS 0.347643
R9941 VSS.n4974 VSS 0.347643
R9942 VSS.n327 VSS 0.347643
R9943 VSS VSS.n1715 0.347643
R9944 VSS VSS.n2893 0.347643
R9945 VSS.n2892 VSS 0.347643
R9946 VSS.n4325 VSS 0.347643
R9947 VSS.n4326 VSS 0.347643
R9948 VSS.n4303 VSS 0.347643
R9949 VSS.n4304 VSS 0.347643
R9950 VSS.n4959 VSS 0.347643
R9951 VSS.n4958 VSS 0.347643
R9952 VSS.n4005 VSS 0.347643
R9953 VSS.n5477 VSS.n12 0.347167
R9954 VSS.n2559 VSS.n2558 0.347167
R9955 VSS.n4025 VSS.n4024 0.347167
R9956 VSS.n2832 VSS.n2831 0.347167
R9957 VSS.n2440 VSS.n2439 0.347167
R9958 VSS.n1110 VSS.n1109 0.347167
R9959 VSS.n2939 VSS.n2936 0.346179
R9960 VSS.n2516 VSS 0.338278
R9961 VSS.n5464 VSS 0.338278
R9962 VSS VSS.n2582 0.338278
R9963 VSS VSS.n1133 0.338278
R9964 VSS VSS.n2424 0.338278
R9965 VSS.n2941 VSS.n2940 0.333376
R9966 VSS.n5102 VSS.n5101 0.3305
R9967 VSS.n5062 VSS.n5061 0.3305
R9968 VSS.n205 VSS.n204 0.3305
R9969 VSS.n177 VSS.n176 0.3305
R9970 VSS.n5416 VSS.n121 0.3305
R9971 VSS.n5136 VSS.n5135 0.3305
R9972 VSS.n5009 VSS.n5003 0.330435
R9973 VSS.n5480 VSS.n5479 0.328278
R9974 VSS.n2555 VSS.n2554 0.328278
R9975 VSS.n4021 VSS.n4020 0.328278
R9976 VSS.n2954 VSS.n2953 0.328278
R9977 VSS.n2529 VSS.n2528 0.328278
R9978 VSS.n1106 VSS.n1105 0.328278
R9979 VSS.n2901 VSS.n2900 0.322918
R9980 VSS.n4540 VSS.n4539 0.320287
R9981 VSS.n4408 VSS.n4407 0.320287
R9982 VSS.n4453 VSS.n994 0.320287
R9983 VSS.n4286 VSS.n4282 0.320287
R9984 VSS.n2920 VSS.n2919 0.320287
R9985 VSS.n4308 VSS.n4307 0.320287
R9986 VSS.n4963 VSS.n4962 0.320287
R9987 VSS.n5088 VSS.n5087 0.30866
R9988 VSS.n278 VSS.n277 0.30866
R9989 VSS.n5106 VSS.n5105 0.30866
R9990 VSS.n5022 VSS.n5021 0.30866
R9991 VSS.n5392 VSS.n5391 0.30866
R9992 VSS.n181 VSS.n180 0.30866
R9993 VSS.n169 VSS.n122 0.30866
R9994 VSS.n63 VSS.n62 0.30866
R9995 VSS.n2507 VSS.n2506 0.30866
R9996 VSS.n2487 VSS.n297 0.303962
R9997 VSS.n2921 VSS.n2920 0.303434
R9998 VSS.n4963 VSS.n371 0.303434
R9999 VSS.n4539 VSS.n4538 0.303434
R10000 VSS.n4453 VSS.n4452 0.303434
R10001 VSS.n4444 VSS.n994 0.303434
R10002 VSS.n4407 VSS.n4406 0.303434
R10003 VSS.n4289 VSS.n4286 0.303434
R10004 VSS.n4282 VSS.n4278 0.303434
R10005 VSS.n2919 VSS.n2868 0.303434
R10006 VSS.n4307 VSS.n4306 0.303434
R10007 VSS.n4962 VSS.n4961 0.303434
R10008 VSS.n4308 VSS.n4204 0.303434
R10009 VSS.n4540 VSS.n4532 0.303434
R10010 VSS.n4409 VSS.n4408 0.303434
R10011 VSS.n179 VSS.n153 0.302175
R10012 VSS.n5104 VSS.n244 0.302175
R10013 VSS.n5091 VSS.n5090 0.299507
R10014 VSS.n5395 VSS.n5394 0.299507
R10015 VSS.n4561 VSS.n4560 0.296241
R10016 VSS.n2523 VSS.n2445 0.293141
R10017 VSS.n5471 VSS.n16 0.293141
R10018 VSS.n2566 VSS.n2565 0.293141
R10019 VSS.n2948 VSS.n2837 0.293141
R10020 VSS.n1117 VSS.n1116 0.293141
R10021 VSS.n4031 VSS.n2594 0.293141
R10022 VSS.n4006 VSS.n2609 0.284171
R10023 VSS.n4232 VSS 0.280143
R10024 VSS VSS.n2510 0.280143
R10025 VSS.n2467 VSS 0.280143
R10026 VSS VSS.n5458 0.280143
R10027 VSS VSS.n5456 0.280143
R10028 VSS VSS.n2913 0.280143
R10029 VSS.n4545 VSS 0.280143
R10030 VSS VSS.n1002 0.280143
R10031 VSS VSS.n1005 0.280143
R10032 VSS.n1029 VSS 0.280143
R10033 VSS VSS.n1061 0.280143
R10034 VSS.n4425 VSS 0.280143
R10035 VSS VSS.n4513 0.280143
R10036 VSS VSS.n758 0.280143
R10037 VSS VSS.n4253 0.280143
R10038 VSS.n4293 VSS 0.280143
R10039 VSS.n341 VSS 0.280143
R10040 VSS VSS.n318 0.280143
R10041 VSS.n4340 VSS 0.280143
R10042 VSS VSS.n2884 0.280143
R10043 VSS VSS.n4324 0.280143
R10044 VSS VSS.n4302 0.280143
R10045 VSS.n530 VSS 0.280143
R10046 VSS VSS.n2606 0.280143
R10047 VSS.n5085 VSS.n5084 0.27986
R10048 VSS.n5070 VSS.n263 0.27986
R10049 VSS.n5019 VSS.n294 0.27986
R10050 VSS.n5389 VSS.n144 0.27986
R10051 VSS.n5405 VSS.n5404 0.27986
R10052 VSS.n5433 VSS.n5432 0.27986
R10053 VSS.n297 VSS.n296 0.279618
R10054 VSS.n5068 VSS.n268 0.279241
R10055 VSS.n5409 VSS.n5408 0.279241
R10056 VSS.n275 VSS.n273 0.27914
R10057 VSS.n5111 VSS.n5110 0.27914
R10058 VSS.n5034 VSS.n5033 0.27914
R10059 VSS.n5451 VSS.n5450 0.27914
R10060 VSS.n182 VSS.n151 0.27914
R10061 VSS.n173 VSS.n172 0.27914
R10062 VSS.n101 VSS.n69 0.27914
R10063 VSS.n2483 VSS.n2482 0.27914
R10064 VSS.n4199 VSS 0.271428
R10065 VSS VSS.n4394 0.271428
R10066 VSS.n4521 VSS 0.271428
R10067 VSS.n367 VSS 0.271428
R10068 VSS VSS.n779 0.2705
R10069 VSS VSS.n303 0.2705
R10070 VSS.n4343 VSS 0.2705
R10071 VSS.n5185 VSS.n5181 0.269731
R10072 VSS.n4043 VSS 0.266056
R10073 VSS.n5066 VSS.n272 0.26546
R10074 VSS.n5412 VSS.n125 0.26546
R10075 VSS.n4185 VSS.n1737 0.263577
R10076 VSS.n4542 VSS.n4522 0.263577
R10077 VSS.n4201 VSS.n4200 0.263577
R10078 VSS.n4398 VSS.n1039 0.263577
R10079 VSS.n4488 VSS.n4483 0.263577
R10080 VSS.n4981 VSS.n4980 0.263577
R10081 VSS.n302 VSS.n299 0.263577
R10082 VSS.n2915 VSS.n1696 0.263577
R10083 VSS.n4965 VSS.n368 0.263577
R10084 VSS.n4372 VSS.n4367 0.263577
R10085 VSS.n3453 VSS.n3448 0.263577
R10086 VSS.n4010 VSS.n4008 0.263
R10087 VSS.n4482 VSS.n4480 0.262423
R10088 VSS.n4365 VSS 0.262029
R10089 VSS.n5093 VSS.n5092 0.26172
R10090 VSS.n5397 VSS.n5396 0.26172
R10091 VSS VSS.n1306 0.256056
R10092 VSS.n5135 VSS.n5134 0.25308
R10093 VSS.n1746 VSS.n1058 0.251199
R10094 VSS.n5121 VSS.n5120 0.250885
R10095 VSS.n257 VSS.n256 0.250885
R10096 VSS.n5043 VSS.n5042 0.250885
R10097 VSS.n5054 VSS.n279 0.250885
R10098 VSS.n115 VSS.n114 0.250885
R10099 VSS.n197 VSS.n196 0.250885
R10100 VSS.n212 VSS.n211 0.250885
R10101 VSS.n166 VSS.n165 0.250885
R10102 VSS.n5423 VSS.n5422 0.250885
R10103 VSS.n5133 VSS.n5132 0.250885
R10104 VSS.n5010 VSS.n5009 0.250885
R10105 VSS.n2523 VSS.n2522 0.249389
R10106 VSS.n5471 VSS.n5470 0.249389
R10107 VSS.n2565 VSS.n2540 0.249389
R10108 VSS.n2948 VSS.n2947 0.249389
R10109 VSS.n1116 VSS.n1091 0.249389
R10110 VSS.n4032 VSS.n4031 0.249389
R10111 VSS.n5096 VSS.n5093 0.248689
R10112 VSS.n5400 VSS.n5397 0.248689
R10113 VSS.n2457 VSS 0.243833
R10114 VSS.n2454 VSS 0.243833
R10115 VSS.n2522 VSS 0.243833
R10116 VSS.n2518 VSS 0.243833
R10117 VSS.n2515 VSS 0.243833
R10118 VSS VSS.n4150 0.243833
R10119 VSS VSS.n14 0.243833
R10120 VSS.n12 VSS 0.243833
R10121 VSS.n28 VSS 0.243833
R10122 VSS.n25 VSS 0.243833
R10123 VSS.n5470 VSS 0.243833
R10124 VSS.n5466 VSS 0.243833
R10125 VSS.n5463 VSS 0.243833
R10126 VSS.n2578 VSS 0.243833
R10127 VSS VSS.n2567 0.243833
R10128 VSS.n2540 VSS 0.243833
R10129 VSS.n2574 VSS 0.243833
R10130 VSS.n2584 VSS 0.243833
R10131 VSS.n2558 VSS 0.243833
R10132 VSS.n2542 VSS 0.243833
R10133 VSS.n2548 VSS 0.243833
R10134 VSS.n4024 VSS 0.243833
R10135 VSS.n2597 VSS 0.243833
R10136 VSS.n2900 VSS 0.243833
R10137 VSS.n2849 VSS 0.243833
R10138 VSS.n2846 VSS 0.243833
R10139 VSS.n2947 VSS 0.243833
R10140 VSS.n2943 VSS 0.243833
R10141 VSS.n2831 VSS 0.243833
R10142 VSS.n2951 VSS 0.243833
R10143 VSS VSS.n2826 0.243833
R10144 VSS.n2439 VSS 0.243833
R10145 VSS.n2526 VSS 0.243833
R10146 VSS VSS.n2434 0.243833
R10147 VSS.n1109 VSS 0.243833
R10148 VSS.n1093 VSS 0.243833
R10149 VSS.n1099 VSS 0.243833
R10150 VSS.n1129 VSS 0.243833
R10151 VSS VSS.n1118 0.243833
R10152 VSS.n1091 VSS 0.243833
R10153 VSS.n1125 VSS 0.243833
R10154 VSS.n1135 VSS 0.243833
R10155 VSS VSS.n1301 0.243833
R10156 VSS VSS.n4039 0.243833
R10157 VSS.n4037 VSS 0.243833
R10158 VSS VSS.n4032 0.243833
R10159 VSS VSS.n4050 0.243833
R10160 VSS VSS.n4103 0.243833
R10161 VSS.n5025 VSS.n5024 0.238749
R10162 VSS.n72 VSS.n71 0.238749
R10163 VSS VSS.n2455 0.237167
R10164 VSS VSS.n2445 0.237167
R10165 VSS.n5485 VSS 0.237167
R10166 VSS VSS.n8 0.237167
R10167 VSS VSS.n26 0.237167
R10168 VSS VSS.n16 0.237167
R10169 VSS VSS.n2537 0.237167
R10170 VSS VSS.n2566 0.237167
R10171 VSS VSS.n2545 0.237167
R10172 VSS VSS.n2549 0.237167
R10173 VSS VSS.n2600 0.237167
R10174 VSS VSS.n4015 0.237167
R10175 VSS VSS.n2847 0.237167
R10176 VSS VSS.n2837 0.237167
R10177 VSS VSS.n2828 0.237167
R10178 VSS.n2825 VSS 0.237167
R10179 VSS VSS.n2436 0.237167
R10180 VSS VSS.n2432 0.237167
R10181 VSS VSS.n1096 0.237167
R10182 VSS VSS.n1100 0.237167
R10183 VSS VSS.n1088 0.237167
R10184 VSS VSS.n1117 0.237167
R10185 VSS VSS.n4038 0.237167
R10186 VSS VSS.n2594 0.237167
R10187 VSS.n5027 VSS.n5026 0.236264
R10188 VSS.n2521 VSS.n2520 0.236056
R10189 VSS.n2517 VSS.n2516 0.236056
R10190 VSS.n2514 VSS.n2513 0.236056
R10191 VSS.n4152 VSS.n4151 0.236056
R10192 VSS.n5474 VSS.n5473 0.236056
R10193 VSS.n5469 VSS.n5468 0.236056
R10194 VSS.n5465 VSS.n5464 0.236056
R10195 VSS.n5462 VSS.n5461 0.236056
R10196 VSS.n2572 VSS.n2571 0.236056
R10197 VSS.n2582 VSS.n2581 0.236056
R10198 VSS.n2588 VSS.n2587 0.236056
R10199 VSS.n2564 VSS.n2563 0.236056
R10200 VSS.n2553 VSS.n2552 0.236056
R10201 VSS.n4030 VSS.n4029 0.236056
R10202 VSS.n4019 VSS.n4018 0.236056
R10203 VSS.n2946 VSS.n2945 0.236056
R10204 VSS.n2942 VSS.n2941 0.236056
R10205 VSS.n2950 VSS.n2949 0.236056
R10206 VSS.n2956 VSS.n2955 0.236056
R10207 VSS.n2525 VSS.n2524 0.236056
R10208 VSS.n2531 VSS.n2530 0.236056
R10209 VSS.n1115 VSS.n1114 0.236056
R10210 VSS.n1104 VSS.n1103 0.236056
R10211 VSS.n1123 VSS.n1122 0.236056
R10212 VSS.n1133 VSS.n1132 0.236056
R10213 VSS.n1139 VSS.n1138 0.236056
R10214 VSS.n4033 VSS.n2591 0.236056
R10215 VSS.n4051 VSS.n2424 0.236056
R10216 VSS.n4106 VSS.n4105 0.236056
R10217 VSS.n374 VSS 0.233577
R10218 VSS.n2918 VSS 0.233577
R10219 VSS VSS.n1736 0.233577
R10220 VSS.n4535 VSS 0.233577
R10221 VSS VSS.n4541 0.233577
R10222 VSS.n4207 VSS 0.233577
R10223 VSS.n4399 VSS 0.233577
R10224 VSS VSS.n1036 0.233577
R10225 VSS VSS.n4487 0.233577
R10226 VSS.n4473 VSS 0.233577
R10227 VSS.n993 VSS 0.233577
R10228 VSS VSS.n4454 0.233577
R10229 VSS VSS.n4977 0.233577
R10230 VSS VSS.n331 0.233577
R10231 VSS.n4281 VSS 0.233577
R10232 VSS.n4285 VSS 0.233577
R10233 VSS VSS.n2867 0.233577
R10234 VSS VSS.n4329 0.233577
R10235 VSS VSS.n4309 0.233577
R10236 VSS VSS.n4964 0.233577
R10237 VSS VSS.n4371 0.233577
R10238 VSS VSS.n3452 0.233577
R10239 VSS.n5031 VSS.n5030 0.233545
R10240 VSS.n99 VSS.n98 0.233545
R10241 VSS.n6 VSS 0.2305
R10242 VSS.n5097 VSS.n5096 0.229074
R10243 VSS.n5446 VSS.n5445 0.229074
R10244 VSS.n5401 VSS.n5400 0.229074
R10245 VSS VSS.n4358 0.2255
R10246 VSS.n2543 VSS.n2542 0.221611
R10247 VSS.n2598 VSS.n2597 0.221611
R10248 VSS.n2952 VSS.n2951 0.221611
R10249 VSS.n2527 VSS.n2526 0.221611
R10250 VSS.n2534 VSS 0.221611
R10251 VSS.n1094 VSS.n1093 0.221611
R10252 VSS VSS.n4237 0.219469
R10253 VSS.n552 VSS 0.219469
R10254 VSS.n4550 VSS 0.219469
R10255 VSS VSS.n4418 0.219469
R10256 VSS VSS.n2822 0.219089
R10257 VSS VSS.n1015 0.218541
R10258 VSS VSS.n4268 0.218541
R10259 VSS.n2875 VSS 0.218541
R10260 VSS.n5487 VSS 0.217167
R10261 VSS.n5026 VSS.n5025 0.214098
R10262 VSS.n92 VSS.n72 0.214098
R10263 VSS.n5478 VSS.n10 0.212722
R10264 VSS.n5008 VSS.n5007 0.208926
R10265 VSS.n248 VSS.n245 0.208926
R10266 VSS.n5049 VSS.n5048 0.208926
R10267 VSS.n210 VSS.n209 0.208926
R10268 VSS.n157 VSS.n154 0.208926
R10269 VSS.n5421 VSS.n5420 0.208926
R10270 VSS.n228 VSS.n225 0.208926
R10271 VSS.n4562 VSS 0.204256
R10272 VSS.n2508 VSS.n2481 0.20138
R10273 VSS.n85 VSS.n46 0.20138
R10274 VSS.n4223 VSS.n4204 0.199786
R10275 VSS.n2921 VSS.n2864 0.199786
R10276 VSS.n531 VSS.n371 0.199786
R10277 VSS.n4532 VSS.n4531 0.199786
R10278 VSS.n4538 VSS.n4536 0.199786
R10279 VSS.n4452 VSS.n996 0.199786
R10280 VSS.n4444 VSS.n1007 0.199786
R10281 VSS.n4410 VSS.n4409 0.199786
R10282 VSS.n4370 VSS.n1073 0.199786
R10283 VSS.n4406 VSS.n4400 0.199786
R10284 VSS.n4486 VSS.n755 0.199786
R10285 VSS.n4474 VSS.n760 0.199786
R10286 VSS.n4290 VSS.n4289 0.199786
R10287 VSS.n4278 VSS.n4257 0.199786
R10288 VSS.n4976 VSS.n4975 0.199786
R10289 VSS.n330 VSS.n322 0.199786
R10290 VSS.n1735 VSS.n1727 0.199786
R10291 VSS.n2886 VSS.n2868 0.199786
R10292 VSS.n4328 VSS.n1740 0.199786
R10293 VSS.n4306 VSS.n4208 0.199786
R10294 VSS.n4961 VSS.n4960 0.199786
R10295 VSS.n3451 VSS.n2610 0.199786
R10296 VSS.n4236 VSS.n4235 0.192
R10297 VSS.n4438 VSS.n1011 0.192
R10298 VSS.n4421 VSS.n1030 0.192
R10299 VSS.n4271 VSS.n4264 0.192
R10300 VSS.n551 VSS.n550 0.1905
R10301 VSS.n4552 VSS.n4551 0.1905
R10302 VSS.n2881 VSS.n2876 0.1905
R10303 VSS.n5014 VSS.n5013 0.189389
R10304 VSS.n5081 VSS.n5080 0.189389
R10305 VSS.n5124 VSS.n5123 0.189389
R10306 VSS.n254 VSS.n252 0.189389
R10307 VSS.n5046 VSS.n5045 0.189389
R10308 VSS.n5057 VSS.n5056 0.189389
R10309 VSS.n118 VSS.n117 0.189389
R10310 VSS.n5440 VSS.n5438 0.189389
R10311 VSS.n141 VSS.n140 0.189389
R10312 VSS.n200 VSS.n199 0.189389
R10313 VSS.n215 VSS.n214 0.189389
R10314 VSS.n163 VSS.n161 0.189389
R10315 VSS.n5426 VSS.n5425 0.189389
R10316 VSS.n5130 VSS.n5128 0.189389
R10317 VSS.n5117 VSS.n5116 0.18928
R10318 VSS.n5098 VSS.n5097 0.18928
R10319 VSS.n5039 VSS.n5038 0.18928
R10320 VSS.n111 VSS.n66 0.18928
R10321 VSS.n5447 VSS.n5446 0.18928
R10322 VSS.n193 VSS.n192 0.18928
R10323 VSS.n5402 VSS.n5401 0.18928
R10324 VSS.n4559 VSS 0.187098
R10325 VSS.n5274 VSS.n5271 0.182808
R10326 VSS VSS.n546 0.1805
R10327 VSS.n5000 VSS.n4998 0.1805
R10328 VSS.n5005 VSS 0.178278
R10329 VSS VSS.n5078 0.178278
R10330 VSS.n236 VSS 0.178278
R10331 VSS VSS.n250 0.178278
R10332 VSS.n288 VSS 0.178278
R10333 VSS VSS.n5051 0.178278
R10334 VSS.n108 VSS 0.178278
R10335 VSS VSS.n60 0.178278
R10336 VSS VSS.n138 0.178278
R10337 VSS.n189 VSS 0.178278
R10338 VSS.n207 VSS 0.178278
R10339 VSS VSS.n159 0.178278
R10340 VSS.n5418 VSS 0.178278
R10341 VSS VSS.n230 0.178278
R10342 VSS.n5086 VSS.n5085 0.177167
R10343 VSS.n266 VSS.n263 0.177167
R10344 VSS.n276 VSS.n275 0.177167
R10345 VSS.n5112 VSS.n5111 0.177167
R10346 VSS.n5020 VSS.n5019 0.177167
R10347 VSS.n5035 VSS.n5034 0.177167
R10348 VSS.n5452 VSS.n5451 0.177167
R10349 VSS.n5390 VSS.n5389 0.177167
R10350 VSS.n5406 VSS.n5405 0.177167
R10351 VSS.n151 VSS.n145 0.177167
R10352 VSS.n172 VSS.n171 0.177167
R10353 VSS.n96 VSS.n69 0.177167
R10354 VSS.n5434 VSS.n5433 0.177167
R10355 VSS.n2505 VSS.n2483 0.177167
R10356 VSS.n5460 VSS.n35 0.176722
R10357 VSS.n4008 VSS.n2606 0.175143
R10358 VSS.n540 VSS 0.175034
R10359 VSS VSS.n4565 0.175034
R10360 VSS.n4365 VSS.n4364 0.173341
R10361 VSS.n4429 VSS.n1020 0.170294
R10362 VSS.n5083 VSS.n5074 0.168962
R10363 VSS.n255 VSS.n246 0.168962
R10364 VSS.n5441 VSS.n56 0.168962
R10365 VSS.n143 VSS.n134 0.168962
R10366 VSS.n164 VSS.n155 0.168962
R10367 VSS.n5131 VSS.n226 0.168962
R10368 VSS.n5012 VSS.n5011 0.168962
R10369 VSS.n4297 VSS.n4296 0.168438
R10370 VSS.n424 VSS.n421 0.167808
R10371 VSS.n2509 VSS.n2474 0.166424
R10372 VSS.n5455 VSS.n5454 0.166424
R10373 VSS.n5492 VSS.n5491 0.166056
R10374 VSS.n5119 VSS.n5118 0.1655
R10375 VSS.n5041 VSS.n5040 0.1655
R10376 VSS.n113 VSS.n112 0.1655
R10377 VSS.n195 VSS.n194 0.1655
R10378 VSS VSS.n241 0.16488
R10379 VSS VSS.n5071 0.16488
R10380 VSS VSS.n260 0.16488
R10381 VSS.n5109 VSS 0.16488
R10382 VSS VSS.n293 0.16488
R10383 VSS VSS.n282 0.16488
R10384 VSS.n5448 VSS 0.16488
R10385 VSS VSS.n148 0.16488
R10386 VSS.n5403 VSS 0.16488
R10387 VSS VSS.n183 0.16488
R10388 VSS VSS.n174 0.16488
R10389 VSS VSS.n102 0.16488
R10390 VSS.n5431 VSS 0.16488
R10391 VSS VSS.n2486 0.16488
R10392 VSS.n4050 VSS.n4049 0.159389
R10393 VSS.n1712 VSS.n1711 0.1575
R10394 VSS.n4463 VSS.n4462 0.1575
R10395 VSS.n4990 VSS.n4989 0.1575
R10396 VSS.n4322 VSS.n4319 0.1565
R10397 VSS.n4511 VSS.n4510 0.1565
R10398 VSS.n4390 VSS.n4387 0.1565
R10399 VSS.n363 VSS.n362 0.1565
R10400 VSS.n5480 VSS.n8 0.155275
R10401 VSS.n2554 VSS.n2545 0.155275
R10402 VSS.n4020 VSS.n2600 0.155275
R10403 VSS.n2954 VSS.n2828 0.155275
R10404 VSS.n2529 VSS.n2436 0.155275
R10405 VSS.n1105 VSS.n1096 0.155275
R10406 VSS.n4391 VSS.n1061 0.154786
R10407 VSS.n4513 VSS.n4512 0.154786
R10408 VSS.n364 VSS.n341 0.154786
R10409 VSS.n4324 VSS.n4323 0.154786
R10410 VSS.n4461 VSS.n758 0.153714
R10411 VSS.n318 VSS.n313 0.153714
R10412 VSS.n4341 VSS.n4340 0.153714
R10413 VSS.n4299 VSS.n4298 0.152665
R10414 VSS.n5445 VSS.n5444 0.151747
R10415 VSS.n992 VSS.n991 0.1505
R10416 VSS.n2512 VSS.n2468 0.149389
R10417 VSS VSS.n1313 0.147167
R10418 VSS VSS.n1318 0.147167
R10419 VSS VSS.n1325 0.147167
R10420 VSS.n4979 VSS.n4978 0.147038
R10421 VSS VSS.n1078 0.144346
R10422 VSS.n93 VSS.n92 0.140703
R10423 VSS.n5032 VSS.n5031 0.138684
R10424 VSS.n100 VSS.n99 0.138684
R10425 VSS.n4367 VSS.n4366 0.137808
R10426 VSS.n3820 VSS.n3819 0.1355
R10427 VSS.n3821 VSS.n3820 0.1355
R10428 VSS.n3822 VSS.n3821 0.1355
R10429 VSS.n3823 VSS.n3822 0.1355
R10430 VSS.n3824 VSS.n3823 0.1355
R10431 VSS.n3825 VSS.n3824 0.1355
R10432 VSS.n3826 VSS.n3825 0.1355
R10433 VSS.n3827 VSS.n3826 0.1355
R10434 VSS.n3828 VSS.n3827 0.1355
R10435 VSS.n3829 VSS.n3828 0.1355
R10436 VSS.n3830 VSS.n3829 0.1355
R10437 VSS.n3831 VSS.n3830 0.1355
R10438 VSS.n3832 VSS.n3831 0.1355
R10439 VSS.n3833 VSS.n3832 0.1355
R10440 VSS.n3834 VSS.n3833 0.1355
R10441 VSS.n3835 VSS.n3834 0.1355
R10442 VSS.n3836 VSS.n3835 0.1355
R10443 VSS.n3837 VSS.n3836 0.1355
R10444 VSS.n3838 VSS.n3837 0.1355
R10445 VSS.n3839 VSS.n3838 0.1355
R10446 VSS.n3840 VSS.n3839 0.1355
R10447 VSS.n3841 VSS.n3840 0.1355
R10448 VSS.n3842 VSS.n3841 0.1355
R10449 VSS.n3844 VSS.n3842 0.1355
R10450 VSS.n3846 VSS.n3844 0.1355
R10451 VSS.n3848 VSS.n3846 0.1355
R10452 VSS.n3850 VSS.n3848 0.1355
R10453 VSS.n3852 VSS.n3850 0.1355
R10454 VSS.n3854 VSS.n3852 0.1355
R10455 VSS.n3856 VSS.n3854 0.1355
R10456 VSS.n3858 VSS.n3856 0.1355
R10457 VSS.n3860 VSS.n3858 0.1355
R10458 VSS.n3862 VSS.n3860 0.1355
R10459 VSS.n3864 VSS.n3862 0.1355
R10460 VSS.n3866 VSS.n3864 0.1355
R10461 VSS.n3868 VSS.n3866 0.1355
R10462 VSS.n3870 VSS.n3868 0.1355
R10463 VSS.n3872 VSS.n3870 0.1355
R10464 VSS.n3874 VSS.n3872 0.1355
R10465 VSS.n3876 VSS.n3874 0.1355
R10466 VSS.n3878 VSS.n3876 0.1355
R10467 VSS.n3880 VSS.n3878 0.1355
R10468 VSS.n3882 VSS.n3880 0.1355
R10469 VSS.n3884 VSS.n3882 0.1355
R10470 VSS.n3886 VSS.n3884 0.1355
R10471 VSS.n3888 VSS.n3886 0.1355
R10472 VSS.n3890 VSS.n3888 0.1355
R10473 VSS.n3892 VSS.n3890 0.1355
R10474 VSS.n3894 VSS.n3892 0.1355
R10475 VSS.n3897 VSS.n3894 0.1355
R10476 VSS.n3899 VSS.n3897 0.1355
R10477 VSS.n3902 VSS.n3899 0.1355
R10478 VSS.n3904 VSS.n3902 0.1355
R10479 VSS.n3907 VSS.n3904 0.1355
R10480 VSS.n3909 VSS.n3907 0.1355
R10481 VSS.n1163 VSS.n1160 0.1355
R10482 VSS.n1166 VSS.n1163 0.1355
R10483 VSS.n1169 VSS.n1166 0.1355
R10484 VSS.n1172 VSS.n1169 0.1355
R10485 VSS.n1175 VSS.n1172 0.1355
R10486 VSS.n1178 VSS.n1175 0.1355
R10487 VSS.n1181 VSS.n1178 0.1355
R10488 VSS.n1184 VSS.n1181 0.1355
R10489 VSS.n1187 VSS.n1184 0.1355
R10490 VSS.n1190 VSS.n1187 0.1355
R10491 VSS.n1193 VSS.n1190 0.1355
R10492 VSS.n1196 VSS.n1193 0.1355
R10493 VSS.n1199 VSS.n1196 0.1355
R10494 VSS.n1202 VSS.n1199 0.1355
R10495 VSS.n1205 VSS.n1202 0.1355
R10496 VSS.n1208 VSS.n1205 0.1355
R10497 VSS.n1211 VSS.n1208 0.1355
R10498 VSS.n1214 VSS.n1211 0.1355
R10499 VSS.n1217 VSS.n1214 0.1355
R10500 VSS.n1220 VSS.n1217 0.1355
R10501 VSS.n1223 VSS.n1220 0.1355
R10502 VSS.n1226 VSS.n1223 0.1355
R10503 VSS.n1229 VSS.n1226 0.1355
R10504 VSS.n1232 VSS.n1229 0.1355
R10505 VSS.n1235 VSS.n1232 0.1355
R10506 VSS.n1238 VSS.n1235 0.1355
R10507 VSS.n1241 VSS.n1238 0.1355
R10508 VSS.n1244 VSS.n1241 0.1355
R10509 VSS.n1247 VSS.n1244 0.1355
R10510 VSS.n1250 VSS.n1247 0.1355
R10511 VSS.n1253 VSS.n1250 0.1355
R10512 VSS.n1256 VSS.n1253 0.1355
R10513 VSS.n1259 VSS.n1256 0.1355
R10514 VSS.n1262 VSS.n1259 0.1355
R10515 VSS.n1265 VSS.n1262 0.1355
R10516 VSS.n1268 VSS.n1265 0.1355
R10517 VSS.n1271 VSS.n1268 0.1355
R10518 VSS.n1274 VSS.n1271 0.1355
R10519 VSS.n1277 VSS.n1274 0.1355
R10520 VSS.n1280 VSS.n1277 0.1355
R10521 VSS.n1283 VSS.n1280 0.1355
R10522 VSS.n1286 VSS.n1283 0.1355
R10523 VSS.n1289 VSS.n1286 0.1355
R10524 VSS.n1292 VSS.n1289 0.1355
R10525 VSS.n1295 VSS.n1292 0.1355
R10526 VSS.n1298 VSS.n1295 0.1355
R10527 VSS.n1336 VSS.n1298 0.1355
R10528 VSS.n1338 VSS.n1336 0.1355
R10529 VSS.n1341 VSS.n1338 0.1355
R10530 VSS.n1343 VSS.n1341 0.1355
R10531 VSS.n1346 VSS.n1343 0.1355
R10532 VSS.n1348 VSS.n1346 0.1355
R10533 VSS.n1676 VSS.n1675 0.1355
R10534 VSS.n1675 VSS.n1672 0.1355
R10535 VSS.n1672 VSS.n1669 0.1355
R10536 VSS.n1669 VSS.n1666 0.1355
R10537 VSS.n1666 VSS.n1663 0.1355
R10538 VSS.n1663 VSS.n1660 0.1355
R10539 VSS.n1660 VSS.n1657 0.1355
R10540 VSS.n1657 VSS.n1654 0.1355
R10541 VSS.n1654 VSS.n1651 0.1355
R10542 VSS.n1651 VSS.n1648 0.1355
R10543 VSS.n1648 VSS.n1641 0.1355
R10544 VSS.n1641 VSS.n1639 0.1355
R10545 VSS.n1639 VSS.n1636 0.1355
R10546 VSS.n1636 VSS.n1634 0.1355
R10547 VSS.n1634 VSS.n1631 0.1355
R10548 VSS.n1631 VSS.n1629 0.1355
R10549 VSS.n1629 VSS.n1626 0.1355
R10550 VSS.n1626 VSS.n1624 0.1355
R10551 VSS.n1624 VSS.n1622 0.1355
R10552 VSS.n1622 VSS.n1620 0.1355
R10553 VSS.n1620 VSS.n1616 0.1355
R10554 VSS.n1616 VSS.n1612 0.1355
R10555 VSS.n1612 VSS.n1609 0.1355
R10556 VSS.n1609 VSS.n1606 0.1355
R10557 VSS.n1606 VSS.n1603 0.1355
R10558 VSS.n1603 VSS.n1600 0.1355
R10559 VSS.n1600 VSS.n1597 0.1355
R10560 VSS.n1597 VSS.n1594 0.1355
R10561 VSS.n1594 VSS.n1591 0.1355
R10562 VSS.n1591 VSS.n1588 0.1355
R10563 VSS.n1588 VSS.n1585 0.1355
R10564 VSS.n1585 VSS.n1582 0.1355
R10565 VSS.n1582 VSS.n1579 0.1355
R10566 VSS.n1579 VSS.n1576 0.1355
R10567 VSS.n1576 VSS.n1573 0.1355
R10568 VSS.n1573 VSS.n1570 0.1355
R10569 VSS.n1570 VSS.n1567 0.1355
R10570 VSS.n1567 VSS.n1564 0.1355
R10571 VSS.n1564 VSS.n1561 0.1355
R10572 VSS.n1561 VSS.n1558 0.1355
R10573 VSS.n1558 VSS.n1555 0.1355
R10574 VSS.n1555 VSS.n1552 0.1355
R10575 VSS.n1552 VSS.n1549 0.1355
R10576 VSS.n1549 VSS.n1546 0.1355
R10577 VSS.n1546 VSS.n1543 0.1355
R10578 VSS.n1508 VSS.n1507 0.1355
R10579 VSS.n1507 VSS.n1504 0.1355
R10580 VSS.n1504 VSS.n1501 0.1355
R10581 VSS.n1501 VSS.n1498 0.1355
R10582 VSS.n1498 VSS.n1495 0.1355
R10583 VSS.n1495 VSS.n1492 0.1355
R10584 VSS.n1492 VSS.n1489 0.1355
R10585 VSS.n1489 VSS.n1486 0.1355
R10586 VSS.n1486 VSS.n1483 0.1355
R10587 VSS.n1483 VSS.n1480 0.1355
R10588 VSS.n1480 VSS.n1477 0.1355
R10589 VSS.n1477 VSS.n1474 0.1355
R10590 VSS.n1474 VSS.n1471 0.1355
R10591 VSS.n1471 VSS.n1468 0.1355
R10592 VSS.n1468 VSS.n1465 0.1355
R10593 VSS.n1465 VSS.n1462 0.1355
R10594 VSS.n1462 VSS.n1459 0.1355
R10595 VSS.n1459 VSS.n1456 0.1355
R10596 VSS.n1456 VSS.n1453 0.1355
R10597 VSS.n1453 VSS.n1450 0.1355
R10598 VSS.n1450 VSS.n1447 0.1355
R10599 VSS.n1447 VSS.n1444 0.1355
R10600 VSS.n1444 VSS.n1441 0.1355
R10601 VSS.n1441 VSS.n1438 0.1355
R10602 VSS.n1438 VSS.n1435 0.1355
R10603 VSS.n1435 VSS.n1432 0.1355
R10604 VSS.n1432 VSS.n1429 0.1355
R10605 VSS.n1429 VSS.n1426 0.1355
R10606 VSS.n1426 VSS.n1423 0.1355
R10607 VSS.n1423 VSS.n1420 0.1355
R10608 VSS.n1420 VSS.n1417 0.1355
R10609 VSS.n1417 VSS.n1414 0.1355
R10610 VSS.n1414 VSS.n1411 0.1355
R10611 VSS.n1411 VSS.n1408 0.1355
R10612 VSS.n1408 VSS.n1405 0.1355
R10613 VSS.n1405 VSS.n1402 0.1355
R10614 VSS.n1402 VSS.n1399 0.1355
R10615 VSS.n1399 VSS.n1396 0.1355
R10616 VSS.n1396 VSS.n1393 0.1355
R10617 VSS.n1393 VSS.n1390 0.1355
R10618 VSS.n792 VSS.n789 0.1355
R10619 VSS.n795 VSS.n792 0.1355
R10620 VSS.n798 VSS.n795 0.1355
R10621 VSS.n801 VSS.n798 0.1355
R10622 VSS.n804 VSS.n801 0.1355
R10623 VSS.n807 VSS.n804 0.1355
R10624 VSS.n810 VSS.n807 0.1355
R10625 VSS.n813 VSS.n810 0.1355
R10626 VSS.n816 VSS.n813 0.1355
R10627 VSS.n819 VSS.n816 0.1355
R10628 VSS.n822 VSS.n819 0.1355
R10629 VSS.n825 VSS.n822 0.1355
R10630 VSS.n828 VSS.n825 0.1355
R10631 VSS.n831 VSS.n828 0.1355
R10632 VSS.n834 VSS.n831 0.1355
R10633 VSS.n837 VSS.n834 0.1355
R10634 VSS.n840 VSS.n837 0.1355
R10635 VSS.n843 VSS.n840 0.1355
R10636 VSS.n846 VSS.n843 0.1355
R10637 VSS.n849 VSS.n846 0.1355
R10638 VSS.n982 VSS.n981 0.1355
R10639 VSS.n981 VSS.n978 0.1355
R10640 VSS.n978 VSS.n975 0.1355
R10641 VSS.n975 VSS.n972 0.1355
R10642 VSS.n972 VSS.n969 0.1355
R10643 VSS.n969 VSS.n966 0.1355
R10644 VSS.n966 VSS.n963 0.1355
R10645 VSS.n963 VSS.n960 0.1355
R10646 VSS.n960 VSS.n957 0.1355
R10647 VSS.n957 VSS.n954 0.1355
R10648 VSS.n954 VSS.n951 0.1355
R10649 VSS.n951 VSS.n948 0.1355
R10650 VSS.n948 VSS.n945 0.1355
R10651 VSS.n945 VSS.n942 0.1355
R10652 VSS.n942 VSS.n939 0.1355
R10653 VSS.n939 VSS.n936 0.1355
R10654 VSS.n936 VSS.n933 0.1355
R10655 VSS.n933 VSS.n930 0.1355
R10656 VSS.n930 VSS.n927 0.1355
R10657 VSS.n927 VSS.n924 0.1355
R10658 VSS.n924 VSS.n921 0.1355
R10659 VSS.n921 VSS.n918 0.1355
R10660 VSS.n918 VSS.n915 0.1355
R10661 VSS.n915 VSS.n912 0.1355
R10662 VSS.n912 VSS.n909 0.1355
R10663 VSS.n909 VSS.n906 0.1355
R10664 VSS.n906 VSS.n903 0.1355
R10665 VSS.n903 VSS.n900 0.1355
R10666 VSS.n900 VSS.n897 0.1355
R10667 VSS.n897 VSS.n894 0.1355
R10668 VSS.n589 VSS.n586 0.1355
R10669 VSS.n592 VSS.n589 0.1355
R10670 VSS.n595 VSS.n592 0.1355
R10671 VSS.n598 VSS.n595 0.1355
R10672 VSS.n601 VSS.n598 0.1355
R10673 VSS.n604 VSS.n601 0.1355
R10674 VSS.n607 VSS.n604 0.1355
R10675 VSS.n610 VSS.n607 0.1355
R10676 VSS.n613 VSS.n610 0.1355
R10677 VSS.n616 VSS.n613 0.1355
R10678 VSS.n619 VSS.n616 0.1355
R10679 VSS.n622 VSS.n619 0.1355
R10680 VSS.n625 VSS.n622 0.1355
R10681 VSS.n628 VSS.n625 0.1355
R10682 VSS.n631 VSS.n628 0.1355
R10683 VSS.n634 VSS.n631 0.1355
R10684 VSS.n637 VSS.n634 0.1355
R10685 VSS.n640 VSS.n637 0.1355
R10686 VSS.n643 VSS.n640 0.1355
R10687 VSS.n646 VSS.n643 0.1355
R10688 VSS.n649 VSS.n646 0.1355
R10689 VSS.n652 VSS.n649 0.1355
R10690 VSS.n655 VSS.n652 0.1355
R10691 VSS.n658 VSS.n655 0.1355
R10692 VSS.n661 VSS.n658 0.1355
R10693 VSS.n664 VSS.n661 0.1355
R10694 VSS.n667 VSS.n664 0.1355
R10695 VSS.n670 VSS.n667 0.1355
R10696 VSS.n673 VSS.n670 0.1355
R10697 VSS.n676 VSS.n673 0.1355
R10698 VSS.n679 VSS.n676 0.1355
R10699 VSS.n682 VSS.n679 0.1355
R10700 VSS.n685 VSS.n682 0.1355
R10701 VSS.n688 VSS.n685 0.1355
R10702 VSS.n691 VSS.n688 0.1355
R10703 VSS.n694 VSS.n691 0.1355
R10704 VSS.n697 VSS.n694 0.1355
R10705 VSS.n700 VSS.n697 0.1355
R10706 VSS.n703 VSS.n700 0.1355
R10707 VSS.n706 VSS.n703 0.1355
R10708 VSS.n709 VSS.n706 0.1355
R10709 VSS.n712 VSS.n709 0.1355
R10710 VSS.n715 VSS.n712 0.1355
R10711 VSS.n718 VSS.n715 0.1355
R10712 VSS.n721 VSS.n718 0.1355
R10713 VSS.n724 VSS.n721 0.1355
R10714 VSS.n383 VSS.n380 0.1355
R10715 VSS.n386 VSS.n383 0.1355
R10716 VSS.n389 VSS.n386 0.1355
R10717 VSS.n392 VSS.n389 0.1355
R10718 VSS.n395 VSS.n392 0.1355
R10719 VSS.n398 VSS.n395 0.1355
R10720 VSS.n401 VSS.n398 0.1355
R10721 VSS.n404 VSS.n401 0.1355
R10722 VSS.n407 VSS.n404 0.1355
R10723 VSS.n410 VSS.n407 0.1355
R10724 VSS.n412 VSS.n410 0.1355
R10725 VSS.n415 VSS.n412 0.1355
R10726 VSS.n417 VSS.n415 0.1355
R10727 VSS.n421 VSS.n417 0.1355
R10728 VSS.n2499 VSS.n2481 0.132897
R10729 VSS.n88 VSS.n85 0.132897
R10730 VSS.n4012 VSS 0.132722
R10731 VSS.n3819 VSS.n3818 0.132038
R10732 VSS.n5489 VSS.n5482 0.129738
R10733 VSS.n1351 VSS.n1348 0.126287
R10734 VSS.n988 VSS.n298 0.122388
R10735 VSS.n2419 VSS.n2417 0.117038
R10736 VSS.n2417 VSS.n2414 0.117038
R10737 VSS.n2414 VSS.n2412 0.117038
R10738 VSS.n2412 VSS.n2409 0.117038
R10739 VSS.n2409 VSS.n2407 0.117038
R10740 VSS.n2407 VSS.n2403 0.117038
R10741 VSS.n2403 VSS.n2400 0.117038
R10742 VSS.n2400 VSS.n2397 0.117038
R10743 VSS.n2397 VSS.n2394 0.117038
R10744 VSS.n4122 VSS.n4119 0.117038
R10745 VSS.n4125 VSS.n4122 0.117038
R10746 VSS.n4128 VSS.n4125 0.117038
R10747 VSS.n4131 VSS.n4128 0.117038
R10748 VSS.n4134 VSS.n4131 0.117038
R10749 VSS.n4137 VSS.n4134 0.117038
R10750 VSS.n4141 VSS.n4137 0.117038
R10751 VSS.n5228 VSS.n5225 0.117038
R10752 VSS.n5231 VSS.n5228 0.117038
R10753 VSS.n5234 VSS.n5231 0.117038
R10754 VSS.n5237 VSS.n5234 0.117038
R10755 VSS.n5240 VSS.n5237 0.117038
R10756 VSS.n5243 VSS.n5240 0.117038
R10757 VSS.n5246 VSS.n5243 0.117038
R10758 VSS.n5249 VSS.n5246 0.117038
R10759 VSS.n5252 VSS.n5249 0.117038
R10760 VSS.n5255 VSS.n5252 0.117038
R10761 VSS.n5258 VSS.n5255 0.117038
R10762 VSS.n5261 VSS.n5258 0.117038
R10763 VSS.n5264 VSS.n5261 0.117038
R10764 VSS.n5267 VSS.n5264 0.117038
R10765 VSS.n5271 VSS.n5267 0.117038
R10766 VSS.n5277 VSS.n5274 0.117038
R10767 VSS.n2385 VSS.n2382 0.117038
R10768 VSS.n2382 VSS.n2379 0.117038
R10769 VSS.n2379 VSS.n2376 0.117038
R10770 VSS.n2376 VSS.n2373 0.117038
R10771 VSS.n2373 VSS.n2370 0.117038
R10772 VSS.n2370 VSS.n2367 0.117038
R10773 VSS.n3529 VSS.n3526 0.117038
R10774 VSS.n3526 VSS.n3523 0.117038
R10775 VSS.n3523 VSS.n2427 0.117038
R10776 VSS.n4056 VSS.n2427 0.117038
R10777 VSS.n4099 VSS.n4056 0.117038
R10778 VSS.n4099 VSS.n4098 0.117038
R10779 VSS.n4098 VSS.n4095 0.117038
R10780 VSS.n4095 VSS.n4092 0.117038
R10781 VSS.n4092 VSS.n4089 0.117038
R10782 VSS.n4089 VSS.n4087 0.117038
R10783 VSS.n4087 VSS.n4084 0.117038
R10784 VSS.n4084 VSS.n4081 0.117038
R10785 VSS.n4081 VSS.n4078 0.117038
R10786 VSS.n4078 VSS.n4075 0.117038
R10787 VSS.n4075 VSS.n4072 0.117038
R10788 VSS.n4072 VSS.n4069 0.117038
R10789 VSS.n4069 VSS.n4066 0.117038
R10790 VSS.n4066 VSS.n4062 0.117038
R10791 VSS.n4062 VSS.n4059 0.117038
R10792 VSS.n4059 VSS.n2422 0.117038
R10793 VSS.n3759 VSS.n3756 0.117038
R10794 VSS.n3756 VSS.n3753 0.117038
R10795 VSS.n3753 VSS.n3750 0.117038
R10796 VSS.n3750 VSS.n3747 0.117038
R10797 VSS.n3747 VSS.n3744 0.117038
R10798 VSS.n3744 VSS.n3741 0.117038
R10799 VSS.n3741 VSS.n3733 0.117038
R10800 VSS.n3733 VSS.n3730 0.117038
R10801 VSS.n3730 VSS.n3728 0.117038
R10802 VSS.n3728 VSS.n3724 0.117038
R10803 VSS.n3724 VSS.n3720 0.117038
R10804 VSS.n3720 VSS.n3717 0.117038
R10805 VSS.n3717 VSS.n3714 0.117038
R10806 VSS.n3714 VSS.n3711 0.117038
R10807 VSS.n3711 VSS.n3708 0.117038
R10808 VSS.n3708 VSS.n3705 0.117038
R10809 VSS.n3705 VSS.n3702 0.117038
R10810 VSS.n3702 VSS.n3699 0.117038
R10811 VSS.n3699 VSS.n3696 0.117038
R10812 VSS.n3696 VSS.n3693 0.117038
R10813 VSS.n3693 VSS.n3690 0.117038
R10814 VSS.n3690 VSS.n3687 0.117038
R10815 VSS.n3687 VSS.n3684 0.117038
R10816 VSS.n3684 VSS.n3681 0.117038
R10817 VSS.n3681 VSS.n3678 0.117038
R10818 VSS.n3678 VSS.n3675 0.117038
R10819 VSS.n3675 VSS.n3672 0.117038
R10820 VSS.n3672 VSS.n3669 0.117038
R10821 VSS.n3669 VSS.n3666 0.117038
R10822 VSS.n3666 VSS.n3663 0.117038
R10823 VSS.n3663 VSS.n3660 0.117038
R10824 VSS.n3660 VSS.n3657 0.117038
R10825 VSS.n3657 VSS.n3654 0.117038
R10826 VSS.n3654 VSS.n3651 0.117038
R10827 VSS.n3651 VSS.n3648 0.117038
R10828 VSS.n3648 VSS.n3645 0.117038
R10829 VSS.n3645 VSS.n3642 0.117038
R10830 VSS.n3642 VSS.n3639 0.117038
R10831 VSS.n3639 VSS.n3636 0.117038
R10832 VSS.n3636 VSS.n3633 0.117038
R10833 VSS.n3633 VSS.n3630 0.117038
R10834 VSS.n3630 VSS.n3627 0.117038
R10835 VSS.n3627 VSS.n3624 0.117038
R10836 VSS.n3624 VSS.n3621 0.117038
R10837 VSS.n3621 VSS.n3618 0.117038
R10838 VSS.n3618 VSS.n3615 0.117038
R10839 VSS.n3615 VSS.n3612 0.117038
R10840 VSS.n3612 VSS.n3609 0.117038
R10841 VSS.n3609 VSS.n3606 0.117038
R10842 VSS.n3606 VSS.n3603 0.117038
R10843 VSS.n3603 VSS.n3600 0.117038
R10844 VSS.n3600 VSS.n3597 0.117038
R10845 VSS.n3597 VSS.n3594 0.117038
R10846 VSS.n3594 VSS.n3591 0.117038
R10847 VSS.n3591 VSS.n3588 0.117038
R10848 VSS.n3588 VSS.n3585 0.117038
R10849 VSS.n3585 VSS.n3582 0.117038
R10850 VSS.n3582 VSS.n3579 0.117038
R10851 VSS.n3579 VSS.n3576 0.117038
R10852 VSS.n3576 VSS.n3573 0.117038
R10853 VSS.n3573 VSS.n3570 0.117038
R10854 VSS.n2338 VSS.n2335 0.117038
R10855 VSS.n2335 VSS.n2332 0.117038
R10856 VSS.n2332 VSS.n2329 0.117038
R10857 VSS.n2329 VSS.n2326 0.117038
R10858 VSS.n4166 VSS.n4163 0.117038
R10859 VSS.n4163 VSS.n4160 0.117038
R10860 VSS.n4160 VSS.n4157 0.117038
R10861 VSS.n4157 VSS.n2289 0.117038
R10862 VSS.n2289 VSS.n2286 0.117038
R10863 VSS.n2286 VSS.n2283 0.117038
R10864 VSS.n2283 VSS.n2280 0.117038
R10865 VSS.n2280 VSS.n2277 0.117038
R10866 VSS.n2277 VSS.n2274 0.117038
R10867 VSS.n2274 VSS.n2271 0.117038
R10868 VSS.n2271 VSS.n2268 0.117038
R10869 VSS.n2268 VSS.n2265 0.117038
R10870 VSS.n2265 VSS.n2262 0.117038
R10871 VSS.n2262 VSS.n2259 0.117038
R10872 VSS.n2259 VSS.n2256 0.117038
R10873 VSS.n2256 VSS.n2253 0.117038
R10874 VSS.n2253 VSS.n2250 0.117038
R10875 VSS.n2250 VSS.n2247 0.117038
R10876 VSS.n2247 VSS.n2244 0.117038
R10877 VSS.n2244 VSS.n2241 0.117038
R10878 VSS.n2241 VSS.n2238 0.117038
R10879 VSS.n2238 VSS.n2235 0.117038
R10880 VSS.n2235 VSS.n2232 0.117038
R10881 VSS.n2232 VSS.n2229 0.117038
R10882 VSS.n2229 VSS.n2226 0.117038
R10883 VSS.n2226 VSS.n2223 0.117038
R10884 VSS.n2223 VSS.n2220 0.117038
R10885 VSS.n2220 VSS.n2217 0.117038
R10886 VSS.n2217 VSS.n2214 0.117038
R10887 VSS.n2214 VSS.n2211 0.117038
R10888 VSS.n2211 VSS.n2208 0.117038
R10889 VSS.n2208 VSS.n2205 0.117038
R10890 VSS.n2205 VSS.n2202 0.117038
R10891 VSS.n2202 VSS.n2199 0.117038
R10892 VSS.n2199 VSS.n2196 0.117038
R10893 VSS.n2196 VSS.n2193 0.117038
R10894 VSS.n2193 VSS.n2190 0.117038
R10895 VSS.n2190 VSS.n2187 0.117038
R10896 VSS.n2187 VSS.n2184 0.117038
R10897 VSS.n2184 VSS.n2181 0.117038
R10898 VSS.n2181 VSS.n2178 0.117038
R10899 VSS.n2178 VSS.n2175 0.117038
R10900 VSS.n2175 VSS.n2172 0.117038
R10901 VSS.n2172 VSS.n2169 0.117038
R10902 VSS.n2169 VSS.n2166 0.117038
R10903 VSS.n2166 VSS.n2163 0.117038
R10904 VSS.n2163 VSS.n2160 0.117038
R10905 VSS.n2160 VSS.n2157 0.117038
R10906 VSS.n2157 VSS.n2154 0.117038
R10907 VSS.n2154 VSS.n2151 0.117038
R10908 VSS.n2151 VSS.n2148 0.117038
R10909 VSS.n2148 VSS.n2145 0.117038
R10910 VSS.n2145 VSS.n2142 0.117038
R10911 VSS.n2142 VSS.n2139 0.117038
R10912 VSS.n2139 VSS.n2136 0.117038
R10913 VSS.n2136 VSS.n2133 0.117038
R10914 VSS.n2133 VSS.n2130 0.117038
R10915 VSS.n2130 VSS.n2127 0.117038
R10916 VSS.n2127 VSS.n2124 0.117038
R10917 VSS.n2124 VSS.n2121 0.117038
R10918 VSS.n2121 VSS.n2118 0.117038
R10919 VSS.n2118 VSS.n2115 0.117038
R10920 VSS.n2115 VSS.n2112 0.117038
R10921 VSS.n2112 VSS.n2109 0.117038
R10922 VSS.n2109 VSS.n2106 0.117038
R10923 VSS.n2106 VSS.n2103 0.117038
R10924 VSS.n2103 VSS.n2100 0.117038
R10925 VSS.n2100 VSS.n2097 0.117038
R10926 VSS.n2097 VSS.n2094 0.117038
R10927 VSS.n2094 VSS.n2091 0.117038
R10928 VSS.n2091 VSS.n2088 0.117038
R10929 VSS.n2088 VSS.n2085 0.117038
R10930 VSS.n2085 VSS.n2082 0.117038
R10931 VSS.n2082 VSS.n2079 0.117038
R10932 VSS.n2037 VSS.n2034 0.117038
R10933 VSS.n2034 VSS.n2031 0.117038
R10934 VSS.n2031 VSS.n2028 0.117038
R10935 VSS.n2028 VSS.n2025 0.117038
R10936 VSS.n2025 VSS.n2022 0.117038
R10937 VSS.n2022 VSS.n2019 0.117038
R10938 VSS.n2019 VSS.n2016 0.117038
R10939 VSS.n2016 VSS.n2013 0.117038
R10940 VSS.n2013 VSS.n2010 0.117038
R10941 VSS.n2010 VSS.n2007 0.117038
R10942 VSS.n2007 VSS.n2004 0.117038
R10943 VSS.n2004 VSS.n2001 0.117038
R10944 VSS.n2001 VSS.n1998 0.117038
R10945 VSS.n1998 VSS.n1995 0.117038
R10946 VSS.n1995 VSS.n1992 0.117038
R10947 VSS.n1992 VSS.n1989 0.117038
R10948 VSS.n1989 VSS.n1986 0.117038
R10949 VSS.n1986 VSS.n1983 0.117038
R10950 VSS.n1983 VSS.n1980 0.117038
R10951 VSS.n1980 VSS.n1977 0.117038
R10952 VSS.n1977 VSS.n1974 0.117038
R10953 VSS.n1974 VSS.n1971 0.117038
R10954 VSS.n1971 VSS.n1968 0.117038
R10955 VSS.n1968 VSS.n1965 0.117038
R10956 VSS.n1965 VSS.n1962 0.117038
R10957 VSS.n1962 VSS.n1959 0.117038
R10958 VSS.n1959 VSS.n1956 0.117038
R10959 VSS.n1956 VSS.n1953 0.117038
R10960 VSS.n1953 VSS.n1950 0.117038
R10961 VSS.n1950 VSS.n1947 0.117038
R10962 VSS.n1947 VSS.n1944 0.117038
R10963 VSS.n1944 VSS.n1941 0.117038
R10964 VSS.n1941 VSS.n1938 0.117038
R10965 VSS.n1938 VSS.n1935 0.117038
R10966 VSS.n1935 VSS.n1932 0.117038
R10967 VSS.n1932 VSS.n1929 0.117038
R10968 VSS.n1929 VSS.n1926 0.117038
R10969 VSS.n1926 VSS.n1923 0.117038
R10970 VSS.n1923 VSS.n1920 0.117038
R10971 VSS.n1920 VSS.n1917 0.117038
R10972 VSS.n1917 VSS.n1914 0.117038
R10973 VSS.n1914 VSS.n1911 0.117038
R10974 VSS.n1911 VSS.n1908 0.117038
R10975 VSS.n1908 VSS.n1905 0.117038
R10976 VSS.n1905 VSS.n1902 0.117038
R10977 VSS.n1902 VSS.n1899 0.117038
R10978 VSS.n1899 VSS.n1896 0.117038
R10979 VSS.n1896 VSS.n1893 0.117038
R10980 VSS.n1893 VSS.n1890 0.117038
R10981 VSS.n1890 VSS.n1887 0.117038
R10982 VSS.n1887 VSS.n1884 0.117038
R10983 VSS.n1884 VSS.n1881 0.117038
R10984 VSS.n1881 VSS.n1878 0.117038
R10985 VSS.n1878 VSS.n1875 0.117038
R10986 VSS.n1875 VSS.n1872 0.117038
R10987 VSS.n1872 VSS.n1869 0.117038
R10988 VSS.n1869 VSS.n1866 0.117038
R10989 VSS.n1866 VSS.n1863 0.117038
R10990 VSS.n1863 VSS.n1860 0.117038
R10991 VSS.n1860 VSS.n1857 0.117038
R10992 VSS.n1857 VSS.n1854 0.117038
R10993 VSS.n1854 VSS.n1851 0.117038
R10994 VSS.n1851 VSS.n1848 0.117038
R10995 VSS.n1848 VSS.n1845 0.117038
R10996 VSS.n1845 VSS.n1842 0.117038
R10997 VSS.n1842 VSS.n1839 0.117038
R10998 VSS.n1839 VSS.n1836 0.117038
R10999 VSS.n1836 VSS.n1833 0.117038
R11000 VSS.n1833 VSS.n1830 0.117038
R11001 VSS.n1830 VSS.n1827 0.117038
R11002 VSS.n1827 VSS.n1824 0.117038
R11003 VSS.n1824 VSS.n1821 0.117038
R11004 VSS.n1821 VSS.n1818 0.117038
R11005 VSS.n1818 VSS.n1815 0.117038
R11006 VSS.n1815 VSS.n1812 0.117038
R11007 VSS.n1812 VSS.n1809 0.117038
R11008 VSS.n1809 VSS.n1806 0.117038
R11009 VSS.n1806 VSS.n1803 0.117038
R11010 VSS.n1803 VSS.n1800 0.117038
R11011 VSS.n1800 VSS.n1797 0.117038
R11012 VSS.n1797 VSS.n1794 0.117038
R11013 VSS.n1794 VSS.n1791 0.117038
R11014 VSS.n1791 VSS.n1788 0.117038
R11015 VSS.n1788 VSS.n1785 0.117038
R11016 VSS.n1785 VSS.n1782 0.117038
R11017 VSS.n1782 VSS.n1779 0.117038
R11018 VSS.n1779 VSS.n1776 0.117038
R11019 VSS.n1776 VSS.n1773 0.117038
R11020 VSS.n3290 VSS.n3287 0.117038
R11021 VSS.n3293 VSS.n3290 0.117038
R11022 VSS.n3296 VSS.n3293 0.117038
R11023 VSS.n3299 VSS.n3296 0.117038
R11024 VSS.n3302 VSS.n3299 0.117038
R11025 VSS.n3305 VSS.n3302 0.117038
R11026 VSS.n3308 VSS.n3305 0.117038
R11027 VSS.n3311 VSS.n3308 0.117038
R11028 VSS.n3314 VSS.n3311 0.117038
R11029 VSS.n3317 VSS.n3314 0.117038
R11030 VSS.n3320 VSS.n3317 0.117038
R11031 VSS.n3323 VSS.n3320 0.117038
R11032 VSS.n3326 VSS.n3323 0.117038
R11033 VSS.n3329 VSS.n3326 0.117038
R11034 VSS.n3332 VSS.n3329 0.117038
R11035 VSS.n3335 VSS.n3332 0.117038
R11036 VSS.n3338 VSS.n3335 0.117038
R11037 VSS.n3341 VSS.n3338 0.117038
R11038 VSS.n3344 VSS.n3341 0.117038
R11039 VSS.n3347 VSS.n3344 0.117038
R11040 VSS.n3350 VSS.n3347 0.117038
R11041 VSS.n3353 VSS.n3350 0.117038
R11042 VSS.n3356 VSS.n3353 0.117038
R11043 VSS.n3359 VSS.n3356 0.117038
R11044 VSS.n3362 VSS.n3359 0.117038
R11045 VSS.n3365 VSS.n3362 0.117038
R11046 VSS.n3368 VSS.n3365 0.117038
R11047 VSS.n3371 VSS.n3368 0.117038
R11048 VSS.n3375 VSS.n3371 0.117038
R11049 VSS.n3378 VSS.n3375 0.117038
R11050 VSS.n3381 VSS.n3378 0.117038
R11051 VSS.n3384 VSS.n3381 0.117038
R11052 VSS.n3387 VSS.n3384 0.117038
R11053 VSS.n3390 VSS.n3387 0.117038
R11054 VSS.n3393 VSS.n3390 0.117038
R11055 VSS.n3396 VSS.n3393 0.117038
R11056 VSS.n3399 VSS.n3396 0.117038
R11057 VSS.n3402 VSS.n3399 0.117038
R11058 VSS.n3405 VSS.n3402 0.117038
R11059 VSS.n3408 VSS.n3405 0.117038
R11060 VSS.n3411 VSS.n3408 0.117038
R11061 VSS.n3414 VSS.n3411 0.117038
R11062 VSS.n3417 VSS.n3414 0.117038
R11063 VSS.n3420 VSS.n3417 0.117038
R11064 VSS.n3423 VSS.n3420 0.117038
R11065 VSS.n3426 VSS.n3423 0.117038
R11066 VSS.n3429 VSS.n3426 0.117038
R11067 VSS.n3432 VSS.n3429 0.117038
R11068 VSS.n3435 VSS.n3432 0.117038
R11069 VSS.n3438 VSS.n3435 0.117038
R11070 VSS.n3441 VSS.n3438 0.117038
R11071 VSS.n3444 VSS.n3441 0.117038
R11072 VSS.n3447 VSS.n3444 0.117038
R11073 VSS.n3457 VSS.n3447 0.117038
R11074 VSS.n3460 VSS.n3457 0.117038
R11075 VSS.n3463 VSS.n3460 0.117038
R11076 VSS.n3466 VSS.n3463 0.117038
R11077 VSS.n3469 VSS.n3466 0.117038
R11078 VSS.n3472 VSS.n3469 0.117038
R11079 VSS.n3475 VSS.n3472 0.117038
R11080 VSS.n3478 VSS.n3475 0.117038
R11081 VSS.n3481 VSS.n3478 0.117038
R11082 VSS VSS.n1020 0.116479
R11083 VSS VSS.n4299 0.116479
R11084 VSS.n4109 VSS.n4108 0.116432
R11085 VSS.n3818 VSS.n3817 0.116342
R11086 VSS.n4565 VSS.n554 0.116021
R11087 VSS.n2910 VSS 0.115552
R11088 VSS VSS.n1016 0.115552
R11089 VSS.n4296 VSS 0.115552
R11090 VSS.n4356 VSS.n1075 0.115394
R11091 VSS.n2367 VSS.n2364 0.113698
R11092 VSS.n852 VSS.n849 0.113655
R11093 VSS.n991 VSS.n990 0.113577
R11094 VSS.n5067 VSS.n269 0.112682
R11095 VSS.n5411 VSS.n5410 0.112682
R11096 VSS.n745 VSS.n557 0.109786
R11097 VSS.n5025 VSS.n5022 0.109456
R11098 VSS.n72 VSS.n63 0.109456
R11099 VSS.n4430 VSS.n1016 0.106273
R11100 VSS.n2391 VSS.n2385 0.1055
R11101 VSS VSS.n2293 0.103212
R11102 VSS.n2509 VSS.n2508 0.102619
R11103 VSS.n5455 VSS.n46 0.102619
R11104 VSS.n3532 VSS.n3529 0.10182
R11105 VSS.n546 VSS.n545 0.100143
R11106 VSS.n543 VSS 0.0997784
R11107 VSS VSS.n523 0.0997784
R11108 VSS VSS.n4434 0.0997784
R11109 VSS VSS.n1023 0.0997784
R11110 VSS VSS.n4198 0.0997784
R11111 VSS VSS.n4393 0.0997784
R11112 VSS VSS.n753 0.0997784
R11113 VSS.n4460 VSS 0.0997784
R11114 VSS.n4300 VSS 0.0997784
R11115 VSS VSS.n4295 0.0997784
R11116 VSS VSS.n365 0.0997784
R11117 VSS.n312 VSS 0.0997784
R11118 VSS VSS.n4342 0.0997784
R11119 VSS VSS.n2 0.0997784
R11120 VSS.n2079 VSS.n2076 0.0987744
R11121 VSS.n1773 VSS.n1770 0.0977902
R11122 VSS.n4234 VSS.n4232 0.0958571
R11123 VSS.n4553 VSS.n4545 0.0958571
R11124 VSS.n4422 VSS.n1029 0.0958571
R11125 VSS.n549 VSS.n530 0.0958571
R11126 VSS.n4220 VSS.n4217 0.0951392
R11127 VSS.n527 VSS.n526 0.0951392
R11128 VSS.n4549 VSS.n4548 0.0951392
R11129 VSS.n4420 VSS.n4419 0.0951392
R11130 VSS.n268 VSS.n267 0.0949444
R11131 VSS.n5030 VSS.n5029 0.0949444
R11132 VSS.n5454 VSS.n5453 0.0949444
R11133 VSS.n5408 VSS.n5407 0.0949444
R11134 VSS.n98 VSS.n97 0.0949444
R11135 VSS.n4439 VSS.n1002 0.0947857
R11136 VSS.n4272 VSS.n4253 0.0947857
R11137 VSS.n2884 VSS.n2883 0.0947857
R11138 VSS.n4437 VSS.n4436 0.0942113
R11139 VSS.n4270 VSS.n4269 0.0942113
R11140 VSS.n2880 VSS.n2879 0.0942113
R11141 VSS.n2909 VSS.n2897 0.0923557
R11142 VSS.n5069 VSS.n5068 0.0919876
R11143 VSS.n5449 VSS.n46 0.0919876
R11144 VSS.n5409 VSS.n126 0.0919876
R11145 VSS.n2508 VSS.n2507 0.0919876
R11146 VSS.n4457 VSS.n4456 0.0916538
R11147 VSS.n4116 VSS.n2422 0.0916538
R11148 VSS.n430 VSS.n427 0.0905
R11149 VSS.n433 VSS.n430 0.0905
R11150 VSS.n436 VSS.n433 0.0905
R11151 VSS.n439 VSS.n436 0.0905
R11152 VSS.n442 VSS.n439 0.0905
R11153 VSS.n445 VSS.n442 0.0905
R11154 VSS.n448 VSS.n445 0.0905
R11155 VSS.n451 VSS.n448 0.0905
R11156 VSS.n454 VSS.n451 0.0905
R11157 VSS.n457 VSS.n454 0.0905
R11158 VSS.n460 VSS.n457 0.0905
R11159 VSS.n463 VSS.n460 0.0905
R11160 VSS.n466 VSS.n463 0.0905
R11161 VSS.n469 VSS.n466 0.0905
R11162 VSS.n472 VSS.n469 0.0905
R11163 VSS.n475 VSS.n472 0.0905
R11164 VSS.n478 VSS.n475 0.0905
R11165 VSS.n481 VSS.n478 0.0905
R11166 VSS.n484 VSS.n481 0.0905
R11167 VSS.n487 VSS.n484 0.0905
R11168 VSS.n490 VSS.n487 0.0905
R11169 VSS.n493 VSS.n490 0.0905
R11170 VSS.n496 VSS.n493 0.0905
R11171 VSS.n499 VSS.n496 0.0905
R11172 VSS.n502 VSS.n499 0.0905
R11173 VSS.n505 VSS.n502 0.0905
R11174 VSS.n508 VSS.n505 0.0905
R11175 VSS.n511 VSS.n508 0.0905
R11176 VSS.n514 VSS.n511 0.0905
R11177 VSS.n517 VSS.n514 0.0905
R11178 VSS.n520 VSS.n517 0.0905
R11179 VSS.n4570 VSS.n520 0.0905
R11180 VSS.n4573 VSS.n4570 0.0905
R11181 VSS.n4576 VSS.n4573 0.0905
R11182 VSS.n4579 VSS.n4576 0.0905
R11183 VSS.n4582 VSS.n4579 0.0905
R11184 VSS.n4585 VSS.n4582 0.0905
R11185 VSS.n4588 VSS.n4585 0.0905
R11186 VSS.n4591 VSS.n4588 0.0905
R11187 VSS.n4594 VSS.n4591 0.0905
R11188 VSS.n4597 VSS.n4594 0.0905
R11189 VSS.n4600 VSS.n4597 0.0905
R11190 VSS.n4603 VSS.n4600 0.0905
R11191 VSS.n4606 VSS.n4603 0.0905
R11192 VSS.n4609 VSS.n4606 0.0905
R11193 VSS.n4612 VSS.n4609 0.0905
R11194 VSS.n4615 VSS.n4612 0.0905
R11195 VSS.n4618 VSS.n4615 0.0905
R11196 VSS.n4621 VSS.n4618 0.0905
R11197 VSS.n4624 VSS.n4621 0.0905
R11198 VSS.n4627 VSS.n4624 0.0905
R11199 VSS.n4630 VSS.n4627 0.0905
R11200 VSS.n4633 VSS.n4630 0.0905
R11201 VSS.n4636 VSS.n4633 0.0905
R11202 VSS.n4639 VSS.n4636 0.0905
R11203 VSS.n4642 VSS.n4639 0.0905
R11204 VSS.n4645 VSS.n4642 0.0905
R11205 VSS.n4649 VSS.n4645 0.0905
R11206 VSS.n4652 VSS.n4649 0.0905
R11207 VSS.n4655 VSS.n4652 0.0905
R11208 VSS.n4658 VSS.n4655 0.0905
R11209 VSS.n4661 VSS.n4658 0.0905
R11210 VSS.n4664 VSS.n4661 0.0905
R11211 VSS.n4667 VSS.n4664 0.0905
R11212 VSS.n4670 VSS.n4667 0.0905
R11213 VSS.n4673 VSS.n4670 0.0905
R11214 VSS.n4676 VSS.n4673 0.0905
R11215 VSS.n4679 VSS.n4676 0.0905
R11216 VSS.n4681 VSS.n4679 0.0905
R11217 VSS.n4683 VSS.n4681 0.0905
R11218 VSS.n4685 VSS.n4683 0.0905
R11219 VSS.n4687 VSS.n4685 0.0905
R11220 VSS.n4689 VSS.n4687 0.0905
R11221 VSS.n4691 VSS.n4689 0.0905
R11222 VSS.n4693 VSS.n4691 0.0905
R11223 VSS.n4695 VSS.n4693 0.0905
R11224 VSS.n4697 VSS.n4695 0.0905
R11225 VSS.n4699 VSS.n4697 0.0905
R11226 VSS.n4701 VSS.n4699 0.0905
R11227 VSS.n4703 VSS.n4701 0.0905
R11228 VSS.n4705 VSS.n4703 0.0905
R11229 VSS.n4707 VSS.n4705 0.0905
R11230 VSS.n4709 VSS.n4707 0.0905
R11231 VSS.n4711 VSS.n4709 0.0905
R11232 VSS.n4713 VSS.n4711 0.0905
R11233 VSS.n4715 VSS.n4713 0.0905
R11234 VSS.n4717 VSS.n4715 0.0905
R11235 VSS.n4720 VSS.n4717 0.0905
R11236 VSS.n4722 VSS.n4720 0.0905
R11237 VSS.n4725 VSS.n4722 0.0905
R11238 VSS.n4727 VSS.n4725 0.0905
R11239 VSS.n4730 VSS.n4727 0.0905
R11240 VSS.n4732 VSS.n4730 0.0905
R11241 VSS.n4735 VSS.n4732 0.0905
R11242 VSS.n4737 VSS.n4735 0.0905
R11243 VSS.n4740 VSS.n4737 0.0905
R11244 VSS.n4742 VSS.n4740 0.0905
R11245 VSS.n4745 VSS.n4742 0.0905
R11246 VSS.n4747 VSS.n4745 0.0905
R11247 VSS.n4941 VSS.n4747 0.0905
R11248 VSS.n4941 VSS.n4940 0.0905
R11249 VSS.n4940 VSS.n4937 0.0905
R11250 VSS.n4937 VSS.n4934 0.0905
R11251 VSS.n4934 VSS.n4931 0.0905
R11252 VSS.n4931 VSS.n4928 0.0905
R11253 VSS.n4928 VSS.n4925 0.0905
R11254 VSS.n4925 VSS.n4922 0.0905
R11255 VSS.n4922 VSS.n4919 0.0905
R11256 VSS.n4919 VSS.n4916 0.0905
R11257 VSS.n4916 VSS.n4913 0.0905
R11258 VSS.n4913 VSS.n4911 0.0905
R11259 VSS.n4911 VSS.n4908 0.0905
R11260 VSS.n4908 VSS.n4906 0.0905
R11261 VSS.n4906 VSS.n4903 0.0905
R11262 VSS.n4903 VSS.n4901 0.0905
R11263 VSS.n4901 VSS.n4898 0.0905
R11264 VSS.n4898 VSS.n4896 0.0905
R11265 VSS.n4896 VSS.n4893 0.0905
R11266 VSS.n4893 VSS.n4891 0.0905
R11267 VSS.n4891 VSS.n4887 0.0905
R11268 VSS.n4887 VSS.n4882 0.0905
R11269 VSS.n4882 VSS.n4879 0.0905
R11270 VSS.n4879 VSS.n4876 0.0905
R11271 VSS.n4876 VSS.n4873 0.0905
R11272 VSS.n4873 VSS.n4870 0.0905
R11273 VSS.n4870 VSS.n4866 0.0905
R11274 VSS.n4866 VSS.n4864 0.0905
R11275 VSS.n4864 VSS.n4862 0.0905
R11276 VSS.n4862 VSS.n4859 0.0905
R11277 VSS.n4859 VSS.n4857 0.0905
R11278 VSS.n4857 VSS.n4855 0.0905
R11279 VSS.n4855 VSS.n4853 0.0905
R11280 VSS.n4853 VSS.n4851 0.0905
R11281 VSS.n4851 VSS.n4849 0.0905
R11282 VSS.n4849 VSS.n4846 0.0905
R11283 VSS.n4846 VSS.n4844 0.0905
R11284 VSS.n4844 VSS.n4841 0.0905
R11285 VSS.n4841 VSS.n4839 0.0905
R11286 VSS.n4839 VSS.n4836 0.0905
R11287 VSS.n4836 VSS.n4834 0.0905
R11288 VSS.n4834 VSS.n4831 0.0905
R11289 VSS.n4831 VSS.n4829 0.0905
R11290 VSS.n4829 VSS.n4826 0.0905
R11291 VSS.n4826 VSS.n4824 0.0905
R11292 VSS.n4824 VSS.n4821 0.0905
R11293 VSS.n4821 VSS.n4819 0.0905
R11294 VSS.n4819 VSS.n4812 0.0905
R11295 VSS.n4812 VSS.n4810 0.0905
R11296 VSS.n4810 VSS.n4807 0.0905
R11297 VSS.n4807 VSS.n4805 0.0905
R11298 VSS.n4805 VSS.n4801 0.0905
R11299 VSS.n4801 VSS.n4797 0.0905
R11300 VSS.n4797 VSS.n4794 0.0905
R11301 VSS.n4794 VSS.n4791 0.0905
R11302 VSS.n4791 VSS.n4788 0.0905
R11303 VSS.n4788 VSS.n4785 0.0905
R11304 VSS.n4785 VSS.n4782 0.0905
R11305 VSS.n4782 VSS.n4780 0.0905
R11306 VSS.n4780 VSS.n4777 0.0905
R11307 VSS.n4777 VSS.n4775 0.0905
R11308 VSS.n4775 VSS.n4772 0.0905
R11309 VSS.n4772 VSS.n4770 0.0905
R11310 VSS.n4770 VSS.n4767 0.0905
R11311 VSS.n4767 VSS.n4765 0.0905
R11312 VSS.n4765 VSS.n4761 0.0905
R11313 VSS.n4761 VSS.n4756 0.0905
R11314 VSS.n4756 VSS.n4753 0.0905
R11315 VSS.n4753 VSS.n4750 0.0905
R11316 VSS.n4750 VSS.n218 0.0905
R11317 VSS.n5378 VSS.n218 0.0905
R11318 VSS.n5378 VSS.n5377 0.0905
R11319 VSS.n5377 VSS.n5375 0.0905
R11320 VSS.n5375 VSS.n5373 0.0905
R11321 VSS.n5373 VSS.n5370 0.0905
R11322 VSS.n5370 VSS.n5368 0.0905
R11323 VSS.n5368 VSS.n5366 0.0905
R11324 VSS.n5366 VSS.n5364 0.0905
R11325 VSS.n5364 VSS.n5362 0.0905
R11326 VSS.n5362 VSS.n5360 0.0905
R11327 VSS.n5360 VSS.n5357 0.0905
R11328 VSS.n5357 VSS.n5355 0.0905
R11329 VSS.n5355 VSS.n5352 0.0905
R11330 VSS.n5352 VSS.n5350 0.0905
R11331 VSS.n5350 VSS.n5347 0.0905
R11332 VSS.n5347 VSS.n5345 0.0905
R11333 VSS.n5345 VSS.n5342 0.0905
R11334 VSS.n5342 VSS.n5340 0.0905
R11335 VSS.n5340 VSS.n5337 0.0905
R11336 VSS.n5337 VSS.n5335 0.0905
R11337 VSS.n5335 VSS.n5332 0.0905
R11338 VSS.n5332 VSS.n5330 0.0905
R11339 VSS.n5330 VSS.n5323 0.0905
R11340 VSS.n5323 VSS.n5321 0.0905
R11341 VSS.n5321 VSS.n5318 0.0905
R11342 VSS.n5318 VSS.n5316 0.0905
R11343 VSS.n5316 VSS.n5312 0.0905
R11344 VSS.n5312 VSS.n5308 0.0905
R11345 VSS.n5308 VSS.n5305 0.0905
R11346 VSS.n5305 VSS.n5302 0.0905
R11347 VSS.n5302 VSS.n5299 0.0905
R11348 VSS.n5299 VSS.n5296 0.0905
R11349 VSS.n5296 VSS.n5293 0.0905
R11350 VSS.n5293 VSS.n5291 0.0905
R11351 VSS.n5291 VSS.n5288 0.0905
R11352 VSS.n5288 VSS.n5286 0.0905
R11353 VSS.n5286 VSS.n5283 0.0905
R11354 VSS.n5283 VSS.n5281 0.0905
R11355 VSS.n5118 VSS.n238 0.0898896
R11356 VSS.n5076 VSS.n5072 0.0898896
R11357 VSS.n5040 VSS.n290 0.0898896
R11358 VSS.n112 VSS.n110 0.0898896
R11359 VSS.n58 VSS.n52 0.0898896
R11360 VSS.n194 VSS.n191 0.0898896
R11361 VSS.n136 VSS.n132 0.0898896
R11362 VSS.n1543 VSS.n1540 0.0898504
R11363 VSS.n4014 VSS.n2603 0.0893889
R11364 VSS.n427 VSS.n424 0.0879615
R11365 VSS.n3817 VSS.n3814 0.0878267
R11366 VSS.n3814 VSS.n3811 0.0878267
R11367 VSS.n3811 VSS.n3808 0.0878267
R11368 VSS.n3808 VSS.n3805 0.0878267
R11369 VSS.n3805 VSS.n3802 0.0878267
R11370 VSS.n3802 VSS.n3799 0.0878267
R11371 VSS.n3799 VSS.n3796 0.0878267
R11372 VSS.n3796 VSS.n3793 0.0878267
R11373 VSS.n3793 VSS.n3790 0.0878267
R11374 VSS.n3790 VSS.n3787 0.0878267
R11375 VSS.n3787 VSS.n3784 0.0878267
R11376 VSS.n3784 VSS.n3781 0.0878267
R11377 VSS.n3781 VSS.n3778 0.0878267
R11378 VSS.n2616 VSS.n2613 0.0878267
R11379 VSS.n2619 VSS.n2616 0.0878267
R11380 VSS.n2622 VSS.n2619 0.0878267
R11381 VSS.n2626 VSS.n2622 0.0878267
R11382 VSS.n2629 VSS.n2626 0.0878267
R11383 VSS.n2632 VSS.n2629 0.0878267
R11384 VSS.n2635 VSS.n2632 0.0878267
R11385 VSS.n2638 VSS.n2635 0.0878267
R11386 VSS.n2641 VSS.n2638 0.0878267
R11387 VSS.n2644 VSS.n2641 0.0878267
R11388 VSS.n2647 VSS.n2644 0.0878267
R11389 VSS.n2650 VSS.n2647 0.0878267
R11390 VSS.n2653 VSS.n2650 0.0878267
R11391 VSS.n2656 VSS.n2653 0.0878267
R11392 VSS.n2659 VSS.n2656 0.0878267
R11393 VSS.n2662 VSS.n2659 0.0878267
R11394 VSS.n2665 VSS.n2662 0.0878267
R11395 VSS.n2668 VSS.n2665 0.0878267
R11396 VSS.n2671 VSS.n2668 0.0878267
R11397 VSS.n2674 VSS.n2671 0.0878267
R11398 VSS.n2677 VSS.n2674 0.0878267
R11399 VSS.n2680 VSS.n2677 0.0878267
R11400 VSS.n2683 VSS.n2680 0.0878267
R11401 VSS.n2686 VSS.n2683 0.0878267
R11402 VSS.n2689 VSS.n2686 0.0878267
R11403 VSS.n2692 VSS.n2689 0.0878267
R11404 VSS.n2695 VSS.n2692 0.0878267
R11405 VSS.n2698 VSS.n2695 0.0878267
R11406 VSS.n2701 VSS.n2698 0.0878267
R11407 VSS.n2704 VSS.n2701 0.0878267
R11408 VSS.n2707 VSS.n2704 0.0878267
R11409 VSS.n2710 VSS.n2707 0.0878267
R11410 VSS.n2713 VSS.n2710 0.0878267
R11411 VSS.n2716 VSS.n2713 0.0878267
R11412 VSS.n2719 VSS.n2716 0.0878267
R11413 VSS.n2722 VSS.n2719 0.0878267
R11414 VSS.n2725 VSS.n2722 0.0878267
R11415 VSS.n2728 VSS.n2725 0.0878267
R11416 VSS.n2731 VSS.n2728 0.0878267
R11417 VSS.n2734 VSS.n2731 0.0878267
R11418 VSS.n2737 VSS.n2734 0.0878267
R11419 VSS.n2740 VSS.n2737 0.0878267
R11420 VSS.n2743 VSS.n2740 0.0878267
R11421 VSS.n2746 VSS.n2743 0.0878267
R11422 VSS.n2749 VSS.n2746 0.0878267
R11423 VSS.n2752 VSS.n2749 0.0878267
R11424 VSS.n2755 VSS.n2752 0.0878267
R11425 VSS.n2758 VSS.n2755 0.0878267
R11426 VSS.n2761 VSS.n2758 0.0878267
R11427 VSS.n2764 VSS.n2761 0.0878267
R11428 VSS.n2767 VSS.n2764 0.0878267
R11429 VSS.n2770 VSS.n2767 0.0878267
R11430 VSS.n2773 VSS.n2770 0.0878267
R11431 VSS.n2776 VSS.n2773 0.0878267
R11432 VSS.n2779 VSS.n2776 0.0878267
R11433 VSS.n2783 VSS.n2779 0.0878267
R11434 VSS.n2786 VSS.n2783 0.0878267
R11435 VSS.n2789 VSS.n2786 0.0878267
R11436 VSS.n2792 VSS.n2789 0.0878267
R11437 VSS.n2795 VSS.n2792 0.0878267
R11438 VSS.n2798 VSS.n2795 0.0878267
R11439 VSS.n2801 VSS.n2798 0.0878267
R11440 VSS.n2804 VSS.n2801 0.0878267
R11441 VSS.n2807 VSS.n2804 0.0878267
R11442 VSS.n2810 VSS.n2807 0.0878267
R11443 VSS.n2813 VSS.n2810 0.0878267
R11444 VSS.n2816 VSS.n2813 0.0878267
R11445 VSS.n2819 VSS.n2816 0.0878267
R11446 VSS.n2962 VSS.n2819 0.0878267
R11447 VSS.n2964 VSS.n2962 0.0878267
R11448 VSS.n2966 VSS.n2964 0.0878267
R11449 VSS.n2968 VSS.n2966 0.0878267
R11450 VSS.n2970 VSS.n2968 0.0878267
R11451 VSS.n2972 VSS.n2970 0.0878267
R11452 VSS.n2975 VSS.n2972 0.0878267
R11453 VSS.n2977 VSS.n2975 0.0878267
R11454 VSS.n2980 VSS.n2977 0.0878267
R11455 VSS.n2982 VSS.n2980 0.0878267
R11456 VSS.n2985 VSS.n2982 0.0878267
R11457 VSS.n2987 VSS.n2985 0.0878267
R11458 VSS.n2990 VSS.n2987 0.0878267
R11459 VSS.n2992 VSS.n2990 0.0878267
R11460 VSS.n2995 VSS.n2992 0.0878267
R11461 VSS.n2997 VSS.n2995 0.0878267
R11462 VSS.n3000 VSS.n2997 0.0878267
R11463 VSS.n3002 VSS.n3000 0.0878267
R11464 VSS.n3008 VSS.n3002 0.0878267
R11465 VSS.n3010 VSS.n3008 0.0878267
R11466 VSS.n3013 VSS.n3010 0.0878267
R11467 VSS.n3015 VSS.n3013 0.0878267
R11468 VSS.n3018 VSS.n3015 0.0878267
R11469 VSS.n3020 VSS.n3018 0.0878267
R11470 VSS.n3024 VSS.n3020 0.0878267
R11471 VSS.n3026 VSS.n3024 0.0878267
R11472 VSS.n3028 VSS.n3026 0.0878267
R11473 VSS.n3030 VSS.n3028 0.0878267
R11474 VSS.n3032 VSS.n3030 0.0878267
R11475 VSS.n3034 VSS.n3032 0.0878267
R11476 VSS.n3036 VSS.n3034 0.0878267
R11477 VSS.n3038 VSS.n3036 0.0878267
R11478 VSS.n3040 VSS.n3038 0.0878267
R11479 VSS.n3042 VSS.n3040 0.0878267
R11480 VSS.n3044 VSS.n3042 0.0878267
R11481 VSS.n3046 VSS.n3044 0.0878267
R11482 VSS.n3048 VSS.n3046 0.0878267
R11483 VSS.n3050 VSS.n3048 0.0878267
R11484 VSS.n3052 VSS.n3050 0.0878267
R11485 VSS.n3054 VSS.n3052 0.0878267
R11486 VSS.n3057 VSS.n3054 0.0878267
R11487 VSS.n3059 VSS.n3057 0.0878267
R11488 VSS.n3062 VSS.n3059 0.0878267
R11489 VSS.n3064 VSS.n3062 0.0878267
R11490 VSS.n3067 VSS.n3064 0.0878267
R11491 VSS.n3069 VSS.n3067 0.0878267
R11492 VSS.n3072 VSS.n3069 0.0878267
R11493 VSS.n3074 VSS.n3072 0.0878267
R11494 VSS.n3077 VSS.n3074 0.0878267
R11495 VSS.n3079 VSS.n3077 0.0878267
R11496 VSS.n3082 VSS.n3079 0.0878267
R11497 VSS.n3084 VSS.n3082 0.0878267
R11498 VSS.n3095 VSS.n3084 0.0878267
R11499 VSS.n3097 VSS.n3095 0.0878267
R11500 VSS.n3098 VSS.n3097 0.0878267
R11501 VSS.n3099 VSS.n3098 0.0878267
R11502 VSS.n3100 VSS.n3099 0.0878267
R11503 VSS.n3101 VSS.n3100 0.0878267
R11504 VSS.n3102 VSS.n3101 0.0878267
R11505 VSS.n3103 VSS.n3102 0.0878267
R11506 VSS.n3104 VSS.n3103 0.0878267
R11507 VSS.n3105 VSS.n3104 0.0878267
R11508 VSS.n3109 VSS.n3108 0.0878267
R11509 VSS.n3110 VSS.n3109 0.0878267
R11510 VSS.n3111 VSS.n3110 0.0878267
R11511 VSS.n3112 VSS.n3111 0.0878267
R11512 VSS.n3113 VSS.n3112 0.0878267
R11513 VSS.n3114 VSS.n3113 0.0878267
R11514 VSS.n3115 VSS.n3114 0.0878267
R11515 VSS.n3116 VSS.n3115 0.0878267
R11516 VSS.n3117 VSS.n3116 0.0878267
R11517 VSS.n3118 VSS.n3117 0.0878267
R11518 VSS.n3119 VSS.n3118 0.0878267
R11519 VSS.n3120 VSS.n3119 0.0878267
R11520 VSS.n3121 VSS.n3120 0.0878267
R11521 VSS.n3122 VSS.n3121 0.0878267
R11522 VSS.n3123 VSS.n3122 0.0878267
R11523 VSS.n3124 VSS.n3123 0.0878267
R11524 VSS.n3125 VSS.n3124 0.0878267
R11525 VSS.n3127 VSS.n3125 0.0878267
R11526 VSS.n3129 VSS.n3127 0.0878267
R11527 VSS.n3131 VSS.n3129 0.0878267
R11528 VSS.n3133 VSS.n3131 0.0878267
R11529 VSS.n3135 VSS.n3133 0.0878267
R11530 VSS.n3137 VSS.n3135 0.0878267
R11531 VSS.n3139 VSS.n3137 0.0878267
R11532 VSS.n3141 VSS.n3139 0.0878267
R11533 VSS.n3143 VSS.n3141 0.0878267
R11534 VSS.n3145 VSS.n3143 0.0878267
R11535 VSS.n3147 VSS.n3145 0.0878267
R11536 VSS.n3149 VSS.n3147 0.0878267
R11537 VSS.n3151 VSS.n3149 0.0878267
R11538 VSS.n3153 VSS.n3151 0.0878267
R11539 VSS.n3155 VSS.n3153 0.0878267
R11540 VSS.n3157 VSS.n3155 0.0878267
R11541 VSS.n3159 VSS.n3157 0.0878267
R11542 VSS.n3161 VSS.n3159 0.0878267
R11543 VSS.n3163 VSS.n3161 0.0878267
R11544 VSS.n3165 VSS.n3163 0.0878267
R11545 VSS.n3167 VSS.n3165 0.0878267
R11546 VSS.n3169 VSS.n3167 0.0878267
R11547 VSS.n3171 VSS.n3169 0.0878267
R11548 VSS.n3173 VSS.n3171 0.0878267
R11549 VSS.n3175 VSS.n3173 0.0878267
R11550 VSS.n3177 VSS.n3175 0.0878267
R11551 VSS.n3179 VSS.n3177 0.0878267
R11552 VSS.n3181 VSS.n3179 0.0878267
R11553 VSS.n3183 VSS.n3181 0.0878267
R11554 VSS.n3185 VSS.n3183 0.0878267
R11555 VSS.n3187 VSS.n3185 0.0878267
R11556 VSS.n3189 VSS.n3187 0.0878267
R11557 VSS.n3191 VSS.n3189 0.0878267
R11558 VSS.n3193 VSS.n3191 0.0878267
R11559 VSS.n3196 VSS.n3193 0.0878267
R11560 VSS.n3198 VSS.n3196 0.0878267
R11561 VSS.n3201 VSS.n3198 0.0878267
R11562 VSS.n3203 VSS.n3201 0.0878267
R11563 VSS.n3206 VSS.n3203 0.0878267
R11564 VSS.n3208 VSS.n3206 0.0878267
R11565 VSS.n3211 VSS.n3208 0.0878267
R11566 VSS.n3213 VSS.n3211 0.0878267
R11567 VSS.n3216 VSS.n3213 0.0878267
R11568 VSS.n3218 VSS.n3216 0.0878267
R11569 VSS.n3221 VSS.n3218 0.0878267
R11570 VSS.n3223 VSS.n3221 0.0878267
R11571 VSS.n3284 VSS.n3223 0.0878267
R11572 VSS.n4009 VSS.n2 0.0830773
R11573 VSS.n2910 VSS.n2909 0.0812216
R11574 VSS.n5491 VSS.n6 0.0805
R11575 VSS.n5088 VSS.n5084 0.079343
R11576 VSS.n5070 VSS.n5069 0.079343
R11577 VSS.n278 VSS.n273 0.079343
R11578 VSS.n5110 VSS.n5106 0.079343
R11579 VSS.n5022 VSS.n294 0.079343
R11580 VSS.n5033 VSS.n5032 0.079343
R11581 VSS.n5450 VSS.n5449 0.079343
R11582 VSS.n5392 VSS.n144 0.079343
R11583 VSS.n5404 VSS.n126 0.079343
R11584 VSS.n182 VSS.n181 0.079343
R11585 VSS.n173 VSS.n122 0.079343
R11586 VSS.n101 VSS.n100 0.079343
R11587 VSS.n5432 VSS.n63 0.079343
R11588 VSS.n2507 VSS.n2482 0.079343
R11589 VSS.n3570 VSS.n3567 0.0767533
R11590 VSS.n5478 VSS.n5477 0.0746176
R11591 VSS.n2559 VSS.n2543 0.0746176
R11592 VSS.n4025 VSS.n2598 0.0746176
R11593 VSS.n2952 VSS.n2832 0.0746176
R11594 VSS.n2527 VSS.n2440 0.0746176
R11595 VSS.n1110 VSS.n1094 0.0746176
R11596 VSS.n553 VSS.n552 0.073799
R11597 VSS.n3287 VSS.n3284 0.0731923
R11598 VSS.n5091 VSS.n5088 0.0726642
R11599 VSS.n5395 VSS.n5392 0.0726642
R11600 VSS.n5065 VSS.n278 0.072617
R11601 VSS.n5413 VSS.n122 0.072617
R11602 VSS.n5491 VSS.n5490 0.0705
R11603 VSS.n4356 VSS 0.0703936
R11604 VSS.n727 VSS.n724 0.0695408
R11605 VSS.n5106 VSS.n5104 0.0694814
R11606 VSS.n181 VSS.n179 0.0694814
R11607 VSS.n2326 VSS.n2323 0.0688819
R11608 VSS.n2360 VSS.n2357 0.0688459
R11609 VSS.n2357 VSS.n2354 0.0688459
R11610 VSS.n2354 VSS.n2351 0.0688459
R11611 VSS.n2351 VSS.n2348 0.0688459
R11612 VSS.n2348 VSS.n2345 0.0688459
R11613 VSS.n2345 VSS.n2342 0.0688459
R11614 VSS.n2608 VSS.n2607 0.068
R11615 VSS.n4230 VSS.n4224 0.068
R11616 VSS.n4231 VSS.n4223 0.068
R11617 VSS.n1734 VSS.n1733 0.068
R11618 VSS.n4529 VSS.n4525 0.068
R11619 VSS.n2923 VSS.n2922 0.068
R11620 VSS.n2864 VSS.n2861 0.068
R11621 VSS.n536 VSS.n532 0.068
R11622 VSS.n537 VSS.n531 0.068
R11623 VSS.n4537 VSS.n746 0.068
R11624 VSS.n4531 VSS.n4530 0.068
R11625 VSS.n4536 VSS.n749 0.068
R11626 VSS.n4515 VSS.n754 0.068
R11627 VSS.n4476 VSS.n4475 0.068
R11628 VSS.n4451 VSS.n4450 0.068
R11629 VSS.n4449 VSS.n996 0.068
R11630 VSS.n4446 VSS.n4445 0.068
R11631 VSS.n4447 VSS.n1007 0.068
R11632 VSS.n4412 VSS.n1033 0.068
R11633 VSS.n4411 VSS.n4410 0.068
R11634 VSS.n4377 VSS.n1073 0.068
R11635 VSS.n4378 VSS.n1072 0.068
R11636 VSS.n4400 VSS.n1026 0.068
R11637 VSS.n4405 VSS.n4404 0.068
R11638 VSS.n4514 VSS.n755 0.068
R11639 VSS.n4477 VSS.n760 0.068
R11640 VSS.n329 VSS.n328 0.068
R11641 VSS.n4288 VSS.n4254 0.068
R11642 VSS.n4291 VSS.n4290 0.068
R11643 VSS.n4277 VSS.n4276 0.068
R11644 VSS.n4257 VSS.n4250 0.068
R11645 VSS.n4973 VSS.n336 0.068
R11646 VSS.n4975 VSS.n4974 0.068
R11647 VSS.n327 VSS.n322 0.068
R11648 VSS.n1727 VSS.n1715 0.068
R11649 VSS.n2893 VSS.n2886 0.068
R11650 VSS.n2892 VSS.n2891 0.068
R11651 VSS.n4325 VSS.n1740 0.068
R11652 VSS.n4327 VSS.n4326 0.068
R11653 VSS.n4303 VSS.n4208 0.068
R11654 VSS.n4305 VSS.n4304 0.068
R11655 VSS.n4960 VSS.n4959 0.068
R11656 VSS.n4958 VSS.n375 0.068
R11657 VSS.n4005 VSS.n2610 0.068
R11658 VSS.n2907 VSS 0.0673041
R11659 VSS.n4431 VSS.n4430 0.0673041
R11660 VSS.n860 VSS.n784 0.0665432
R11661 VSS.n5120 VSS.n5119 0.0662692
R11662 VSS.n5122 VSS.n5121 0.0662692
R11663 VSS.n5095 VSS.n5094 0.0662692
R11664 VSS.n257 VSS.n245 0.0662692
R11665 VSS.n256 VSS.n255 0.0662692
R11666 VSS.n5042 VSS.n5041 0.0662692
R11667 VSS.n5044 VSS.n5043 0.0662692
R11668 VSS.n5048 VSS.n279 0.0662692
R11669 VSS.n5055 VSS.n5054 0.0662692
R11670 VSS.n114 VSS.n113 0.0662692
R11671 VSS.n116 VSS.n115 0.0662692
R11672 VSS.n54 VSS.n53 0.0662692
R11673 VSS.n5442 VSS.n5441 0.0662692
R11674 VSS.n196 VSS.n195 0.0662692
R11675 VSS.n198 VSS.n197 0.0662692
R11676 VSS.n5399 VSS.n5398 0.0662692
R11677 VSS.n211 VSS.n210 0.0662692
R11678 VSS.n213 VSS.n212 0.0662692
R11679 VSS.n166 VSS.n154 0.0662692
R11680 VSS.n165 VSS.n164 0.0662692
R11681 VSS.n5422 VSS.n5421 0.0662692
R11682 VSS.n5424 VSS.n5423 0.0662692
R11683 VSS.n5133 VSS.n225 0.0662692
R11684 VSS.n5132 VSS.n5131 0.0662692
R11685 VSS.n5009 VSS.n5008 0.0662692
R11686 VSS.n5012 VSS.n5010 0.0662692
R11687 VSS.n5006 VSS.n5005 0.0660556
R11688 VSS.n5078 VSS.n5077 0.0660556
R11689 VSS.n237 VSS.n236 0.0660556
R11690 VSS.n250 VSS.n249 0.0660556
R11691 VSS.n289 VSS.n288 0.0660556
R11692 VSS.n5051 VSS.n5050 0.0660556
R11693 VSS.n109 VSS.n108 0.0660556
R11694 VSS.n60 VSS.n59 0.0660556
R11695 VSS.n138 VSS.n137 0.0660556
R11696 VSS.n190 VSS.n189 0.0660556
R11697 VSS.n208 VSS.n207 0.0660556
R11698 VSS.n159 VSS.n158 0.0660556
R11699 VSS.n5419 VSS.n5418 0.0660556
R11700 VSS.n230 VSS.n229 0.0660556
R11701 VSS.n4119 VSS.n4116 0.0639615
R11702 VSS.n5066 VSS.n5065 0.0635185
R11703 VSS.n5413 VSS.n5412 0.0635185
R11704 VSS.n4319 VSS.n4318 0.0625
R11705 VSS.n4510 VSS.n4509 0.0625
R11706 VSS.n4387 VSS.n4386 0.0625
R11707 VSS.n362 VSS.n361 0.0625
R11708 VSS.n1711 VSS.n1710 0.0615
R11709 VSS.n4464 VSS.n4463 0.0615
R11710 VSS.n4991 VSS.n4990 0.0615
R11711 VSS.n4178 VSS.n1750 0.0608
R11712 VSS.n863 VSS.n861 0.058921
R11713 VSS.n1048 VSS.n1043 0.0571038
R11714 VSS.n4347 VSS.n1140 0.0534048
R11715 VSS.n1151 VSS.n1149 0.053063
R11716 VSS.n3519 VSS.n3517 0.053063
R11717 VSS.n3773 VSS.n3771 0.053063
R11718 VSS.n560 VSS.n558 0.0527581
R11719 VSS.n1147 VSS.n1146 0.0526849
R11720 VSS.n1144 VSS.n1143 0.0526849
R11721 VSS.n3515 VSS.n3514 0.0526849
R11722 VSS.n3513 VSS.n3512 0.0526849
R11723 VSS.n3768 VSS.n3767 0.0526849
R11724 VSS.n4110 VSS.n4109 0.0503305
R11725 VSS.n2394 VSS.n2391 0.0501154
R11726 VSS.n5444 VSS.n5443 0.049129
R11727 VSS.n5013 VSS.n295 0.0471667
R11728 VSS.n5082 VSS.n5081 0.0471667
R11729 VSS.n5123 VSS.n232 0.0471667
R11730 VSS.n254 VSS.n253 0.0471667
R11731 VSS.n5045 VSS.n284 0.0471667
R11732 VSS.n5056 VSS.n5053 0.0471667
R11733 VSS.n117 VSS.n104 0.0471667
R11734 VSS.n5440 VSS.n5439 0.0471667
R11735 VSS.n142 VSS.n141 0.0471667
R11736 VSS.n199 VSS.n185 0.0471667
R11737 VSS.n214 VSS.n202 0.0471667
R11738 VSS.n163 VSS.n162 0.0471667
R11739 VSS.n5425 VSS.n120 0.0471667
R11740 VSS.n5130 VSS.n5129 0.0471667
R11741 VSS.n1685 VSS.n1153 0.0470126
R11742 VSS.n3545 VSS.n3509 0.0470126
R11743 VSS.n3544 VSS.n3520 0.0470126
R11744 VSS.n3979 VSS.n3775 0.0470126
R11745 VSS.n3540 VSS.n3536 0.0467273
R11746 VSS.n5281 VSS.n5277 0.0455
R11747 VSS.n2339 VSS.n2338 0.0436087
R11748 VSS.n222 VSS.n221 0.0434545
R11749 VSS.n3484 VSS.n3481 0.0428588
R11750 VSS.n272 VSS.n271 0.0427222
R11751 VSS.n125 VSS.n124 0.0427222
R11752 VSS.n3912 VSS.n3909 0.0425965
R11753 VSS.n5166 VSS.n5165 0.0422273
R11754 VSS.n3983 VSS.n3982 0.0417185
R11755 VSS.n5027 VSS 0.040834
R11756 VSS.n3994 VSS.n3759 0.0390371
R11757 VSS.n1691 VSS.n1690 0.0383151
R11758 VSS.n2364 VSS.n2361 0.037718
R11759 VSS.n3539 VSS.n3538 0.0367416
R11760 VSS.n3538 VSS.n3537 0.0361376
R11761 VSS.n1720 VSS.n1712 0.0345
R11762 VSS.n4322 VSS.n4189 0.0345
R11763 VSS.n4511 VSS.n4499 0.0345
R11764 VSS.n4462 VSS.n775 0.0345
R11765 VSS.n4390 VSS.n1064 0.0345
R11766 VSS.n4989 VSS.n4986 0.0345
R11767 VSS.n363 VSS.n351 0.0345
R11768 VSS.n5160 VSS.n5159 0.0336364
R11769 VSS.n1748 VSS.n1747 0.0330131
R11770 VSS.n2907 VSS.n2906 0.0329742
R11771 VSS.n5155 VSS.n5154 0.0328182
R11772 VSS.n2432 VSS.n2430 0.0327222
R11773 VSS.n4194 VSS 0.0325
R11774 VSS.n4504 VSS 0.0325
R11775 VSS VSS.n4385 0.0325
R11776 VSS.n356 VSS 0.0325
R11777 VSS.n5149 VSS.n5148 0.0324091
R11778 VSS.n5003 VSS.n297 0.03218
R11779 VSS.n2361 VSS.n2360 0.0316278
R11780 VSS.n1705 VSS 0.0315
R11781 VSS.n4465 VSS 0.0315
R11782 VSS.n4992 VSS 0.0315
R11783 VSS.n1047 VSS.n1046 0.0307655
R11784 VSS.n560 VSS.n559 0.0306935
R11785 VSS.n1043 VSS.n1042 0.0295733
R11786 VSS.n5225 VSS.n5222 0.0291851
R11787 VSS.n1362 VSS.n1360 0.0274767
R11788 VSS.n1356 VSS.n1355 0.0272442
R11789 VSS.n5487 VSS.n5486 0.0271667
R11790 VSS.n4001 VSS.n4000 0.0267717
R11791 VSS.n3557 VSS.n3554 0.0266207
R11792 VSS.n3505 VSS.n3502 0.0262514
R11793 VSS.n2342 VSS.n2339 0.0262143
R11794 VSS.n3107 VSS.n3105 0.0254505
R11795 VSS.n3562 VSS.n3559 0.0253276
R11796 VSS.n2307 VSS.n2304 0.0252684
R11797 VSS.n93 VSS 0.02496
R11798 VSS.n5490 VSS.n5489 0.0249444
R11799 VSS.n2067 VSS.n2064 0.0248048
R11800 VSS.n1519 VSS.n1516 0.0245
R11801 VSS.n4179 VSS.n1748 0.0240602
R11802 VSS.n5188 VSS.n5187 0.0234091
R11803 VSS.n5140 VSS.n5139 0.023
R11804 VSS.n1526 VSS.n1523 0.0229444
R11805 VSS.n5200 VSS.n5199 0.0225909
R11806 VSS.n5175 VSS.n5172 0.0221818
R11807 VSS.n5212 VSS.n5211 0.0221818
R11808 VSS.n1682 VSS.n1364 0.0221279
R11809 VSS.n2316 VSS.n2313 0.0220804
R11810 VSS.n3916 VSS.n3914 0.0220686
R11811 VSS.n3493 VSS.n3490 0.0213092
R11812 VSS.n1352 VSS.n1351 0.0209651
R11813 VSS.n4298 VSS.n4239 0.0209124
R11814 VSS.n2902 VSS.n2852 0.0207941
R11815 VSS.n4563 VSS.n4562 0.0207649
R11816 VSS.n5176 VSS.n5175 0.0205455
R11817 VSS.n2046 VSS.n2043 0.0204733
R11818 VSS.n4145 VSS.n4141 0.0201154
R11819 VSS.n3108 VSS.n3107 0.020104
R11820 VSS.n2852 VSS 0.0199118
R11821 VSS.n2511 VSS.n2469 0.0197857
R11822 VSS.n2058 VSS.n2055 0.0195107
R11823 VSS.n2076 VSS.n2073 0.0190294
R11824 VSS.n4145 VSS.n2419 0.0189615
R11825 VSS.n2298 VSS.n1753 0.0181567
R11826 VSS.n570 VSS.n569 0.018061
R11827 VSS.n1533 VSS.n1530 0.0173889
R11828 VSS.n3972 VSS.n3918 0.0173627
R11829 VSS.n5141 VSS.n5140 0.0172727
R11830 VSS.n4009 VSS 0.017201
R11831 VSS.n3550 VSS.n3549 0.0170517
R11832 VSS.n863 VSS.n862 0.0168158
R11833 VSS.n1691 VSS.n1141 0.0162531
R11834 VSS.n223 VSS.n222 0.0160455
R11835 VSS.n853 VSS.n852 0.0158061
R11836 VSS.n3549 VSS.n3546 0.0157586
R11837 VSS.n3496 VSS.n3493 0.0155867
R11838 VSS.n4047 VSS.n4046 0.015145
R11839 VSS.n2055 VSS.n2052 0.0149385
R11840 VSS.n5139 VSS.n223 0.0144091
R11841 VSS.n1535 VSS.n1533 0.0142778
R11842 VSS.n564 VSS.n563 0.0142195
R11843 VSS.n3567 VSS.n3564 0.0142069
R11844 VSS.n1759 VSS.n1758 0.0141364
R11845 VSS.n5067 VSS.n5066 0.0138884
R11846 VSS.n5412 VSS.n5411 0.0138884
R11847 VSS.n6 VSS.n5 0.0138333
R11848 VSS.n1048 VSS.n1047 0.0137168
R11849 VSS.n3991 VSS.n3990 0.013135
R11850 VSS.n4172 VSS.n1753 0.0130068
R11851 VSS.n3976 VSS.n3974 0.0128529
R11852 VSS.n2319 VSS.n2316 0.0127616
R11853 VSS.n3977 VSS.n3976 0.0122647
R11854 VSS.n5159 VSS.n5158 0.0119545
R11855 VSS.n4171 VSS.n4169 0.0117807
R11856 VSS.n580 VSS.n579 0.01175
R11857 VSS.n2323 VSS.n2320 0.0115354
R11858 VSS.n987 VSS.n860 0.0115072
R11859 VSS.n1540 VSS.n1537 0.0113889
R11860 VSS.n3563 VSS.n3562 0.0113621
R11861 VSS.n3541 VSS.n3540 0.0111364
R11862 VSS.n3502 VSS.n3499 0.0109046
R11863 VSS.n3973 VSS.n3972 0.0108922
R11864 VSS.n3762 VSS.n3761 0.0108922
R11865 VSS.n2903 VSS.n2898 0.0108124
R11866 VSS.n5087 VSS 0.0105
R11867 VSS.n267 VSS 0.0105
R11868 VSS.n277 VSS 0.0105
R11869 VSS.n5105 VSS 0.0105
R11870 VSS.n5021 VSS 0.0105
R11871 VSS.n5029 VSS 0.0105
R11872 VSS.n5453 VSS 0.0105
R11873 VSS.n5391 VSS 0.0105
R11874 VSS.n5407 VSS 0.0105
R11875 VSS.n180 VSS 0.0105
R11876 VSS VSS.n169 0.0105
R11877 VSS.n97 VSS 0.0105
R11878 VSS.n62 VSS 0.0105
R11879 VSS.n2506 VSS 0.0105
R11880 VSS.n3533 VSS.n3532 0.0103276
R11881 VSS.n4048 VSS.n4047 0.0101923
R11882 VSS.n1759 VSS.n1756 0.0101503
R11883 VSS.n2049 VSS.n2046 0.0101257
R11884 VSS.n3554 VSS.n3551 0.00981034
R11885 VSS.n5163 VSS.n5162 0.0095
R11886 VSS.n5178 VSS.n5177 0.0095
R11887 VSS.n5187 VSS.n5186 0.0095
R11888 VSS.n3991 VSS.n3988 0.00944168
R11889 VSS.n14 VSS.n10 0.00938889
R11890 VSS.n741 VSS.n740 0.0090061
R11891 VSS.n1528 VSS.n1526 0.00894444
R11892 VSS.n5157 VSS.n5155 0.00868182
R11893 VSS.n5196 VSS.n5189 0.00868182
R11894 VSS.n5199 VSS.n5198 0.00868182
R11895 VSS.n5220 VSS.n5219 0.00868182
R11896 VSS.n5165 VSS.n5163 0.00827273
R11897 VSS.n5177 VSS.n5176 0.00827273
R11898 VSS.n1692 VSS.n1691 0.00826224
R11899 VSS.n3107 VSS.n3106 0.00789726
R11900 VSS.n1769 VSS.n219 0.00786364
R11901 VSS.n857 VSS.n856 0.00784694
R11902 VSS.n5171 VSS.n5170 0.00781712
R11903 VSS.n1683 VSS.n1682 0.00747674
R11904 VSS.n2304 VSS.n2301 0.00736649
R11905 VSS.n728 VSS.n727 0.00681098
R11906 VSS.n5222 VSS.n5221 0.0065905
R11907 VSS.n5169 VSS.n5168 0.00622727
R11908 VSS.n4436 VSS 0.00606701
R11909 VSS.n4269 VSS 0.00606701
R11910 VSS.n2879 VSS 0.00606701
R11911 VSS.n3917 VSS.n3916 0.0059902
R11912 VSS.n4000 VSS.n3997 0.00596243
R11913 VSS.n573 VSS.n560 0.00594885
R11914 VSS.n1355 VSS.n1353 0.00584884
R11915 VSS.n1363 VSS.n1362 0.00584884
R11916 VSS.n5148 VSS.n5147 0.00581818
R11917 VSS.n5208 VSS.n5207 0.00581818
R11918 VSS.n5221 VSS.n5220 0.00581818
R11919 VSS.n5153 VSS.n5151 0.00540909
R11920 VSS.n5151 VSS.n5149 0.00540909
R11921 VSS.n5147 VSS.n5144 0.00540909
R11922 VSS.n221 VSS.n220 0.00540909
R11923 VSS.n5207 VSS.n5200 0.00540909
R11924 VSS.n5210 VSS.n5209 0.00540909
R11925 VSS.n5211 VSS.n5210 0.00540909
R11926 VSS.n3984 VSS.n3983 0.00516523
R11927 VSS VSS.n4217 0.00513918
R11928 VSS.n527 VSS 0.00513918
R11929 VSS.n4549 VSS 0.00513918
R11930 VSS.n4419 VSS 0.00513918
R11931 VSS.n4297 VSS.n4241 0.00513918
R11932 VSS.n2064 VSS.n2061 0.00507219
R11933 VSS.n2902 VSS.n2901 0.00491176
R11934 VSS.n2070 VSS.n2067 0.00483155
R11935 VSS.n5158 VSS.n5157 0.00459091
R11936 VSS.n5198 VSS.n5197 0.00459091
R11937 VSS.n4179 VSS.n4178 0.00448601
R11938 VSS.n3487 VSS.n3484 0.00440173
R11939 VSS.n3983 VSS.n3760 0.00436002
R11940 VSS.n2940 VSS 0.00402941
R11941 VSS.n891 VSS.n890 0.00396939
R11942 VSS.n2042 VSS.n2040 0.00386898
R11943 VSS.n2519 VSS 0.00383333
R11944 VSS.n5479 VSS 0.00383333
R11945 VSS.n5467 VSS 0.00383333
R11946 VSS.n2575 VSS 0.00383333
R11947 VSS.n2555 VSS 0.00383333
R11948 VSS.n4021 VSS 0.00383333
R11949 VSS.n2944 VSS 0.00383333
R11950 VSS.n2953 VSS 0.00383333
R11951 VSS.n2528 VSS 0.00383333
R11952 VSS.n1106 VSS 0.00383333
R11953 VSS.n1126 VSS 0.00383333
R11954 VSS VSS.n4042 0.00383333
R11955 VSS.n1521 VSS.n1519 0.00383333
R11956 VSS.n5168 VSS.n5166 0.00377273
R11957 VSS.n5162 VSS.n5160 0.00377273
R11958 VSS.n5172 VSS.n5171 0.00377273
R11959 VSS.n5179 VSS.n5178 0.00377273
R11960 VSS.n1710 VSS 0.0035
R11961 VSS VSS.n4464 0.0035
R11962 VSS VSS.n4991 0.0035
R11963 VSS.n5146 VSS.n5145 0.0034492
R11964 VSS.n987 VSS.n986 0.00343706
R11965 VSS.n1770 VSS.n1769 0.00336364
R11966 VSS.n4429 VSS.n4428 0.00328351
R11967 VSS.n873 VSS.n863 0.00322727
R11968 VSS.n5170 VSS.n219 0.00318129
R11969 VSS.n5154 VSS.n5153 0.00295455
R11970 VSS.n5209 VSS.n5208 0.00295455
R11971 VSS.n2310 VSS.n2307 0.00295232
R11972 VSS.n870 VSS.n869 0.00294898
R11973 VSS VSS.n366 0.00280769
R11974 VSS VSS.n2917 0.00280769
R11975 VSS.n1737 VSS 0.00280769
R11976 VSS VSS.n750 0.00280769
R11977 VSS.n4542 VSS 0.00280769
R11978 VSS VSS.n4201 0.00280769
R11979 VSS VSS.n4398 0.00280769
R11980 VSS.n4396 VSS 0.00280769
R11981 VSS.n4488 VSS 0.00280769
R11982 VSS.n4480 VSS 0.00280769
R11983 VSS VSS.n992 0.00280769
R11984 VSS.n4457 VSS 0.00280769
R11985 VSS.n4978 VSS 0.00280769
R11986 VSS.n4981 VSS 0.00280769
R11987 VSS VSS.n299 0.00280769
R11988 VSS.n4998 VSS 0.00280769
R11989 VSS.n2915 VSS 0.00280769
R11990 VSS.n2856 VSS 0.00280769
R11991 VSS.n4330 VSS 0.00280769
R11992 VSS.n4310 VSS 0.00280769
R11993 VSS.n4965 VSS 0.00280769
R11994 VSS.n4372 VSS 0.00280769
R11995 VSS.n3453 VSS 0.00280769
R11996 VSS.n733 VSS.n730 0.00276891
R11997 VSS.n1056 VSS.n1055 0.00276891
R11998 VSS.n859 VSS.n786 0.00276891
R11999 VSS.n1146 VSS.n1145 0.00276891
R12000 VSS.n1143 VSS.n1142 0.00276891
R12001 VSS.n3512 VSS.n3511 0.00276891
R12002 VSS.n3767 VSS.n3765 0.00276891
R12003 VSS.n4178 VSS.n4177 0.00275
R12004 VSS.n4439 VSS 0.00264286
R12005 VSS.n4272 VSS 0.00264286
R12006 VSS.n2883 VSS 0.00264286
R12007 VSS.n5197 VSS.n5196 0.00254545
R12008 VSS.n5219 VSS.n5212 0.00254545
R12009 VSS.n877 VSS.n876 0.00254082
R12010 VSS.n4318 VSS 0.0025
R12011 VSS.n4509 VSS 0.0025
R12012 VSS.n4386 VSS 0.0025
R12013 VSS.n361 VSS 0.0025
R12014 VSS.n3540 VSS.n3539 0.00238811
R12015 VSS.n1051 VSS.n1048 0.00217832
R12016 VSS.n1688 VSS.n1685 0.00213052
R12017 VSS.n3490 VSS.n3487 0.00206069
R12018 VSS.n3564 VSS.n3563 0.00205172
R12019 VSS.n743 VSS.n736 0.00201261
R12020 VSS.n1045 VSS.n1044 0.00201261
R12021 VSS.n985 VSS.n885 0.00201261
R12022 VSS.n2320 VSS.n2319 0.00197139
R12023 VSS.n2073 VSS.n2070 0.00194385
R12024 VSS.n1353 VSS.n1352 0.00189535
R12025 VSS.n1750 VSS.n1749 0.00185
R12026 VSS.n1537 VSS.n1535 0.00183333
R12027 VSS.n3980 VSS.n3979 0.00175579
R12028 VSS.n3544 VSS.n3543 0.00175577
R12029 VSS.n4175 VSS.n4174 0.00175575
R12030 VSS.n1761 VSS.n1760 0.00175281
R12031 VSS.n3536 VSS.n3535 0.00172727
R12032 VSS.n5186 VSS.n5179 0.00172727
R12033 VSS.n5189 VSS.n5188 0.00172727
R12034 VSS.n857 VSS.n853 0.00172449
R12035 VSS.n3914 VSS.n3913 0.00167647
R12036 VSS.n4045 VSS.n4044 0.00165385
R12037 VSS.n572 VSS.n566 0.00163445
R12038 VSS.n1050 VSS.n1049 0.00163445
R12039 VSS.n872 VSS.n866 0.00163445
R12040 VSS.n1148 VSS.n1147 0.00163445
R12041 VSS.n1149 VSS.n1144 0.00163445
R12042 VSS.n3516 VSS.n3515 0.00163445
R12043 VSS.n3517 VSS.n3513 0.00163445
R12044 VSS.n3771 VSS.n3768 0.00163445
R12045 VSS.n3770 VSS.n3769 0.00163445
R12046 VSS.n745 VSS.n744 0.00162735
R12047 VSS.n5014 VSS 0.00161111
R12048 VSS.n5080 VSS 0.00161111
R12049 VSS.n5124 VSS 0.00161111
R12050 VSS VSS.n5086 0.00161111
R12051 VSS VSS.n266 0.00161111
R12052 VSS VSS.n276 0.00161111
R12053 VSS.n252 VSS 0.00161111
R12054 VSS.n5112 VSS 0.00161111
R12055 VSS.n5046 VSS 0.00161111
R12056 VSS VSS.n5020 0.00161111
R12057 VSS.n5057 VSS 0.00161111
R12058 VSS.n5035 VSS 0.00161111
R12059 VSS VSS.n2521 0.00161111
R12060 VSS VSS.n2517 0.00161111
R12061 VSS VSS.n2514 0.00161111
R12062 VSS.n118 VSS 0.00161111
R12063 VSS.n4152 VSS 0.00161111
R12064 VSS.n5492 VSS 0.00161111
R12065 VSS.n5474 VSS 0.00161111
R12066 VSS VSS.n5469 0.00161111
R12067 VSS VSS.n5465 0.00161111
R12068 VSS VSS.n5462 0.00161111
R12069 VSS.n5438 VSS 0.00161111
R12070 VSS VSS.n5452 0.00161111
R12071 VSS.n140 VSS 0.00161111
R12072 VSS.n200 VSS 0.00161111
R12073 VSS VSS.n5390 0.00161111
R12074 VSS VSS.n5406 0.00161111
R12075 VSS.n215 VSS 0.00161111
R12076 VSS VSS.n145 0.00161111
R12077 VSS.n161 VSS 0.00161111
R12078 VSS.n171 VSS 0.00161111
R12079 VSS.n5426 VSS 0.00161111
R12080 VSS VSS.n96 0.00161111
R12081 VSS.n5434 VSS 0.00161111
R12082 VSS.n2571 VSS 0.00161111
R12083 VSS.n2581 VSS 0.00161111
R12084 VSS.n2587 VSS 0.00161111
R12085 VSS.n2563 VSS 0.00161111
R12086 VSS.n2552 VSS 0.00161111
R12087 VSS.n4029 VSS 0.00161111
R12088 VSS.n4018 VSS 0.00161111
R12089 VSS VSS.n2853 0.00161111
R12090 VSS VSS.n2946 0.00161111
R12091 VSS VSS.n2942 0.00161111
R12092 VSS VSS.n2950 0.00161111
R12093 VSS.n2956 VSS 0.00161111
R12094 VSS.n5128 VSS 0.00161111
R12095 VSS VSS.n2505 0.00161111
R12096 VSS VSS.n2525 0.00161111
R12097 VSS.n2531 VSS 0.00161111
R12098 VSS.n1114 VSS 0.00161111
R12099 VSS.n1103 VSS 0.00161111
R12100 VSS.n1122 VSS 0.00161111
R12101 VSS.n1132 VSS 0.00161111
R12102 VSS.n1138 VSS 0.00161111
R12103 VSS.n1302 VSS 0.00161111
R12104 VSS.n4033 VSS 0.00161111
R12105 VSS.n4051 VSS 0.00161111
R12106 VSS.n4105 VSS 0.00161111
R12107 VSS.n1514 VSS.n1513 0.00161111
R12108 VSS.n741 VSS.n737 0.00159756
R12109 VSS VSS.n4234 0.00157143
R12110 VSS.n4553 VSS 0.00157143
R12111 VSS.n4422 VSS 0.00157143
R12112 VSS VSS.n549 0.00157143
R12113 VSS.n986 VSS.n883 0.00154895
R12114 VSS.n3997 VSS.n3994 0.00154046
R12115 VSS.n4108 VSS 0.00151695
R12116 VSS.n4172 VSS.n4171 0.00148093
R12117 VSS.n2043 VSS.n2042 0.00146257
R12118 VSS.n1516 VSS.n1514 0.00138889
R12119 VSS.n1756 VSS.n1755 0.00133916
R12120 VSS.n1693 VSS.n1692 0.00133916
R12121 VSS.n983 VSS.n891 0.00131633
R12122 VSS.n3499 VSS.n3496 0.00128035
R12123 VSS.n3985 VSS.n3984 0.00127754
R12124 VSS.n3988 VSS.n3987 0.00127754
R12125 VSS.n3559 VSS.n3558 0.00127586
R12126 VSS.n2501 VSS 0.0012438
R12127 VSS VSS.n2499 0.0012438
R12128 VSS VSS.n88 0.0012438
R12129 VSS VSS.n91 0.0012438
R12130 VSS VSS.n4353 0.0012438
R12131 VSS.n2313 VSS.n2310 0.0012357
R12132 VSS.n2061 VSS.n2058 0.00122193
R12133 VSS.n1530 VSS.n1528 0.00116667
R12134 VSS.n3918 VSS.n3917 0.00108824
R12135 VSS.n744 VSS.n734 0.00106367
R12136 VSS.n3558 VSS.n3557 0.00101724
R12137 VSS.n1359 VSS.n1356 0.000965116
R12138 VSS.n4177 VSS.n4176 0.00095
R12139 VSS.n1054 VSS.n1051 0.00091958
R12140 VSS.n1057 VSS.n1054 0.00091958
R12141 VSS.n883 VSS.n873 0.00091958
R12142 VSS.n1755 VSS.n1754 0.00091958
R12143 VSS.n1758 VSS.n1757 0.00091958
R12144 VSS.n3542 VSS.n3541 0.000909091
R12145 VSS.n3987 VSS.n3986 0.000888769
R12146 VSS.n3990 VSS.n3989 0.000888769
R12147 VSS.n582 VSS.n576 0.000878151
R12148 VSS.n1053 VSS.n1052 0.000878151
R12149 VSS.n882 VSS.n879 0.000878151
R12150 VSS.n1153 VSS.n1151 0.000878151
R12151 VSS.n1690 VSS.n1689 0.000878151
R12152 VSS.n3520 VSS.n3519 0.000878151
R12153 VSS.n3775 VSS.n3773 0.000878151
R12154 VSS.n3982 VSS.n3981 0.000878151
R12155 VSS.n583 VSS.n573 0.000875783
R12156 VSS.n734 VSS.n583 0.000875783
R12157 VSS.n3508 VSS.n3505 0.000760116
R12158 VSS.n4001 VSS.n3508 0.000760116
R12159 VSS.n3551 VSS.n3550 0.000758621
R12160 VSS.n2301 VSS.n2298 0.000745232
R12161 VSS.n2052 VSS.n2049 0.000740642
R12162 VSS.n1360 VSS.n1359 0.000732558
R12163 VSS.n1364 VSS.n1363 0.000732558
R12164 VSS.n1523 VSS.n1521 0.000722222
R12165 VSS.n3913 VSS.n3912 0.000696078
R12166 VSS.n3974 VSS.n3973 0.000696078
R12167 7b_counter_0.MDFF_6.QB.n6 7b_counter_0.MDFF_6.QB.t8 53.2954
R12168 7b_counter_0.MDFF_6.QB.t9 7b_counter_0.MDFF_6.QB.t7 44.058
R12169 7b_counter_0.MDFF_6.QB.n0 7b_counter_0.MDFF_6.QB.t5 38.8649
R12170 7b_counter_0.MDFF_6.QB.t5 7b_counter_0.MDFF_6.QB.t9 28.6791
R12171 7b_counter_0.MDFF_6.QB 7b_counter_0.MDFF_6.QB.n7 19.3781
R12172 7b_counter_0.MDFF_6.QB.n7 7b_counter_0.MDFF_6.QB.t4 17.1425
R12173 7b_counter_0.MDFF_6.QB.n7 7b_counter_0.MDFF_6.QB.t10 14.405
R12174 7b_counter_0.MDFF_6.QB.n0 7b_counter_0.MDFF_6.QB.t6 7.3005
R12175 7b_counter_0.MDFF_6.QB.t10 7b_counter_0.MDFF_6.QB.n6 7.3005
R12176 7b_counter_0.MDFF_6.QB 7b_counter_0.MDFF_6.QB.n0 5.42109
R12177 7b_counter_0.MDFF_6.QB.n6 7b_counter_0.MDFF_6.QB.n5 4.51584
R12178 7b_counter_0.MDFF_6.QB.n5 7b_counter_0.MDFF_6.QB.n2 3.62007
R12179 7b_counter_0.MDFF_6.QB.n5 7b_counter_0.MDFF_6.QB.n4 3.15478
R12180 7b_counter_0.MDFF_6.QB.n4 7b_counter_0.MDFF_6.QB.t0 1.6255
R12181 7b_counter_0.MDFF_6.QB.n4 7b_counter_0.MDFF_6.QB.n3 1.6255
R12182 7b_counter_0.MDFF_6.QB.n2 7b_counter_0.MDFF_6.QB.t3 1.463
R12183 7b_counter_0.MDFF_6.QB.n2 7b_counter_0.MDFF_6.QB.n1 1.463
R12184 Q3.t15 Q3.t30 47.8944
R12185 Q3.t5 Q3.t21 47.8944
R12186 Q3.t14 Q3.t27 47.5387
R12187 Q3.t31 Q3.t19 47.5387
R12188 Q3.t28 Q3.t22 44.058
R12189 Q3.n24 Q3.n23 42.1039
R12190 Q3.n1 Q3.t8 38.8649
R12191 Q3.n11 Q3.t12 38.7949
R12192 Q3.n10 Q3.t7 38.7949
R12193 Q3.n4 Q3.t29 38.7949
R12194 Q3.n3 Q3.t25 38.7949
R12195 Q3.t3 Q3.t18 31.5469
R12196 Q3.t6 Q3.t16 31.5469
R12197 Q3.t26 Q3.t6 31.5469
R12198 Q3.t13 Q3.t26 31.5469
R12199 Q3.n11 Q3.n10 31.4949
R12200 Q3.n4 Q3.n3 31.4949
R12201 Q3.t18 Q3.t24 28.8094
R12202 Q3.t8 Q3.t28 28.6791
R12203 Q3.n30 Q3.n24 18.1935
R12204 Q3.n12 Q3.t4 17.9416
R12205 Q3.n5 Q3.t23 17.9416
R12206 Q3.n0 Q3.t13 16.3603
R12207 Q3.n14 Q3.t14 15.7085
R12208 Q3.n6 Q3.t31 15.7085
R12209 Q3.n0 Q3.t3 15.1871
R12210 Q3.n14 Q3.t17 13.4273
R12211 Q3.n6 Q3.t9 13.4273
R12212 Q3.n12 Q3.t15 11.957
R12213 Q3.n5 Q3.t5 11.957
R12214 Q3.n24 Q3.n2 9.75009
R12215 Q3.n1 Q3.t10 7.3005
R12216 Q3.n10 Q3.t20 7.3005
R12217 Q3.t4 Q3.n11 7.3005
R12218 Q3.n3 Q3.t11 7.3005
R12219 Q3.t23 Q3.n4 7.3005
R12220 Q3.n8 Q3.n7 7.10835
R12221 Q3 Q3.n0 6.7187
R12222 Q3 Q3.n12 5.94647
R12223 Q3 Q3.n5 5.94647
R12224 Q3.n28 Q3.n27 5.47387
R12225 Q3 Q3.n1 5.27587
R12226 Q3.n29 Q3.n25 4.65398
R12227 Q3.n28 Q3.n26 4.2255
R12228 Q3 Q3.n14 4.08021
R12229 Q3 Q3.n6 4.08021
R12230 Q3.n7 Q3 2.64035
R12231 Q3.n15 Q3 2.37798
R12232 Q3.n16 Q3.n15 2.2505
R12233 Q3.n23 Q3.n22 2.24343
R12234 Q3.n18 Q3.n17 1.49758
R12235 Q3.n13 Q3 0.473682
R12236 Q3.n7 Q3 0.472202
R12237 Q3.n29 Q3.n28 0.427022
R12238 Q3 Q3.n29 0.257096
R12239 Q3.n15 Q3.n13 0.229175
R12240 Q3 Q3.n31 0.184413
R12241 Q3.n19 Q3.n18 0.182545
R12242 Q3.n9 Q3.n8 0.030875
R12243 Q3.n30 Q3 0.0260556
R12244 Q3.n31 Q3 0.0238333
R12245 Q3.n23 Q3.n20 0.0172614
R12246 Q3.n20 Q3.n19 0.0161888
R12247 Q3.n2 Q3 0.0130316
R12248 Q3.n18 Q3.n9 0.012519
R12249 Q3.n2 Q3 0.00733544
R12250 Q3.n31 Q3.n30 0.00383333
R12251 Q3.n17 Q3.n16 0.00165385
R12252 Q3.n22 Q3.n21 0.00165385
R12253 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t15 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t14 47.8944
R12254 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n7 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t16 38.7949
R12255 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n8 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t17 38.7949
R12256 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n8 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n7 31.4949
R12257 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n9 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t13 17.9416
R12258 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n9 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t15 11.957
R12259 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n7 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t12 7.3005
R12260 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t13 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n8 7.3005
R12261 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n10 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN 5.93058
R12262 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n9 5.86474
R12263 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n2 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t1 5.68507
R12264 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n6 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t9 4.92604
R12265 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n15 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n12 3.6455
R12266 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n15 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n14 3.31072
R12267 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n5 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n4 3.1505
R12268 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n18 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n17 2.90572
R12269 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n2 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n1 2.6005
R12270 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n10 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN 1.88467
R12271 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n1 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t0 1.6255
R12272 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n1 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n0 1.6255
R12273 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n14 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t7 1.6255
R12274 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n14 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n13 1.6255
R12275 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n17 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t6 1.6255
R12276 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n17 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n16 1.6255
R12277 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n4 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t11 1.463
R12278 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n4 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n3 1.463
R12279 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n12 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t3 1.463
R12280 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n12 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n11 1.463
R12281 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n10 1.33598
R12282 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n6 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n5 1.15166
R12283 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n5 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n2 0.898543
R12284 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n18 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n15 0.4055
R12285 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n6 0.198522
R12286 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n18 0.178625
R12287 D2_4.t13 D2_4.t2 47.8944
R12288 D2_4.t4 D2_4.t21 47.8944
R12289 D2_4.t14 D2_4.t0 47.5387
R12290 D2_4.t5 D2_4.t18 47.5387
R12291 D2_4.t3 D2_4.t6 44.058
R12292 D2_4.t11 D2_4.t25 44.058
R12293 D2_4.n21 D2_4.t22 38.8649
R12294 D2_4.n18 D2_4.t24 38.8649
R12295 D2_4.n13 D2_4.t15 38.7949
R12296 D2_4.n12 D2_4.t16 38.7949
R12297 D2_4.n4 D2_4.t7 38.7949
R12298 D2_4.n3 D2_4.t9 38.7949
R12299 D2_4.n19 D2_4.n17 35.649
R12300 D2_4.n13 D2_4.n12 31.4949
R12301 D2_4.n4 D2_4.n3 31.4949
R12302 D2_4.t22 D2_4.t3 28.6791
R12303 D2_4.t24 D2_4.t11 28.6791
R12304 D2_4.n14 D2_4.t1 17.9416
R12305 D2_4.n5 D2_4.t19 17.9416
R12306 D2_4.n15 D2_4.t14 16.621
R12307 D2_4.n6 D2_4.t5 16.621
R12308 D2_4.n17 D2_4.n11 13.9752
R12309 D2_4.n15 D2_4.t17 12.5148
R12310 D2_4.n6 D2_4.t10 12.5148
R12311 D2_4.n14 D2_4.t13 11.957
R12312 D2_4.n5 D2_4.t4 11.957
R12313 D2_4.n20 D2_4.n19 8.296
R12314 D2_4.n21 D2_4.t23 7.3005
R12315 D2_4.n18 D2_4.t8 7.3005
R12316 D2_4.n12 D2_4.t20 7.3005
R12317 D2_4.t1 D2_4.n13 7.3005
R12318 D2_4.n3 D2_4.t12 7.3005
R12319 D2_4.t19 D2_4.n4 7.3005
R12320 D2_4 D2_4.n14 5.95286
R12321 D2_4 D2_4.n5 5.95286
R12322 D2_4 D2_4.n21 5.27587
R12323 D2_4 D2_4.n18 5.27587
R12324 D2_4 D2_4.n15 4.59246
R12325 D2_4 D2_4.n6 4.59246
R12326 D2_4.n2 D2_4.n1 4.5005
R12327 D2_4.n8 D2_4.n2 3.45961
R12328 D2_4.n19 D2_4 3.3199
R12329 D2_4.n17 D2_4.n16 2.62295
R12330 D2_4.n9 D2_4.n8 2.25138
R12331 D2_4.n11 D2_4.n1 2.24334
R12332 D2_4.n10 D2_4.n9 1.5081
R12333 D2_4.n7 D2_4 1.37202
R12334 D2_4.n16 D2_4 1.30354
R12335 D2_4.n16 D2_4 0.24123
R12336 D2_4.n7 D2_4 0.172752
R12337 D2_4.n8 D2_4.n7 0.167374
R12338 D2_4.n20 D2_4.n0 0.0468264
R12339 D2_4 D2_4.n20 0.0339615
R12340 D2_4.n10 D2_4.n2 0.0312595
R12341 D2_4.n11 D2_4.n10 0.0174666
R12342 D2_4.n0 D2_4 0.0108108
R12343 D2_4.n0 D2_4 0.00311992
R12344 D2_4.n9 D2_4.n1 0.00176987
R12345 p2_gen_magic_0.xnor_magic_3.OUT.t8 p2_gen_magic_0.xnor_magic_3.OUT.t6 28.8746
R12346 p2_gen_magic_0.xnor_magic_3.OUT.n1 p2_gen_magic_0.xnor_magic_3.OUT.t5 25.7891
R12347 p2_gen_magic_0.xnor_magic_3.OUT.t5 p2_gen_magic_0.xnor_magic_3.OUT.t4 23.4648
R12348 p2_gen_magic_0.xnor_magic_3.OUT.n5 p2_gen_magic_0.xnor_magic_3.OUT.n2 17.1813
R12349 p2_gen_magic_0.xnor_magic_3.OUT.n0 p2_gen_magic_0.xnor_magic_3.OUT.t7 17.1425
R12350 p2_gen_magic_0.xnor_magic_3.OUT.n0 p2_gen_magic_0.xnor_magic_3.OUT.t8 14.405
R12351 p2_gen_magic_0.xnor_magic_3.OUT.n5 p2_gen_magic_0.xnor_magic_3.OUT.n4 4.11507
R12352 p2_gen_magic_0.xnor_magic_3.OUT.n1 p2_gen_magic_0.xnor_magic_3.OUT.n0 3.62425
R12353 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_3.OUT.n5 3.61488
R12354 p2_gen_magic_0.xnor_magic_3.OUT.n2 p2_gen_magic_0.xnor_magic_3.OUT 2.33511
R12355 p2_gen_magic_0.xnor_magic_3.OUT.n4 p2_gen_magic_0.xnor_magic_3.OUT.t1 1.463
R12356 p2_gen_magic_0.xnor_magic_3.OUT.n4 p2_gen_magic_0.xnor_magic_3.OUT.n3 1.463
R12357 p2_gen_magic_0.xnor_magic_3.OUT.n2 p2_gen_magic_0.xnor_magic_3.OUT.n1 0.853219
R12358 P2.t13 P2.t8 47.8944
R12359 P2.t11 P2.t12 44.6331
R12360 P2.t6 P2.t11 43.4094
R12361 P2.n0 P2.t7 38.7949
R12362 P2.n1 P2.t14 38.7949
R12363 P2.t10 P2.t6 31.5469
R12364 P2.n1 P2.n0 31.4949
R12365 P2.n4 P2 24.839
R12366 P2.n2 P2.t9 17.9416
R12367 P2.n3 P2.t10 15.0567
R12368 P2.n3 P2.t16 13.6228
R12369 P2.n2 P2.t13 11.957
R12370 P2.n0 P2.t15 7.3005
R12371 P2.t9 P2.n1 7.3005
R12372 P2 P2.n2 5.86241
R12373 P2 P2.n3 4.2675
R12374 P2.n11 P2.n8 3.6455
R12375 P2.n11 P2.n10 3.31072
R12376 P2.n12 P2.n6 2.90572
R12377 P2.n6 P2.t4 1.6255
R12378 P2.n6 P2.n5 1.6255
R12379 P2.n10 P2.t3 1.6255
R12380 P2.n10 P2.n9 1.6255
R12381 P2.n8 P2.t1 1.463
R12382 P2.n8 P2.n7 1.463
R12383 P2.n13 P2 0.642239
R12384 P2.n4 P2 0.625183
R12385 P2.n12 P2.n11 0.4055
R12386 P2 P2.n4 0.382718
R12387 P2 P2.n12 0.178625
R12388 P2.n13 P2 0.12963
R12389 P2 P2.n13 0.112022
R12390 p3_gen_magic_0.xnor_magic_1.B.t6 p3_gen_magic_0.xnor_magic_1.B.t4 47.8944
R12391 p3_gen_magic_0.xnor_magic_1.B.t11 p3_gen_magic_0.xnor_magic_1.B.t9 47.5387
R12392 p3_gen_magic_0.xnor_magic_1.B.n1 p3_gen_magic_0.xnor_magic_1.B.t5 38.7949
R12393 p3_gen_magic_0.xnor_magic_1.B.n0 p3_gen_magic_0.xnor_magic_1.B.t3 38.7949
R12394 p3_gen_magic_0.xnor_magic_1.B.n1 p3_gen_magic_0.xnor_magic_1.B.n0 31.4949
R12395 p3_gen_magic_0.xnor_magic_1.B.n2 p3_gen_magic_0.xnor_magic_1.B.t10 17.9416
R12396 p3_gen_magic_0.xnor_magic_1.B.n3 p3_gen_magic_0.xnor_magic_1.B.t11 16.621
R12397 p3_gen_magic_0.xnor_magic_1.B.n3 p3_gen_magic_0.xnor_magic_1.B.t8 12.5148
R12398 p3_gen_magic_0.xnor_magic_1.B.n2 p3_gen_magic_0.xnor_magic_1.B.t6 11.957
R12399 p3_gen_magic_0.xnor_magic_1.B.n0 p3_gen_magic_0.xnor_magic_1.B.t7 7.3005
R12400 p3_gen_magic_0.xnor_magic_1.B.t10 p3_gen_magic_0.xnor_magic_1.B.n1 7.3005
R12401 p3_gen_magic_0.xnor_magic_1.B p3_gen_magic_0.xnor_magic_1.B.n2 5.95286
R12402 p3_gen_magic_0.xnor_magic_1.B p3_gen_magic_0.xnor_magic_1.B.n3 4.53752
R12403 D2_3.t6 D2_3.t21 47.8944
R12404 D2_3.t15 D2_3.t2 47.8944
R12405 D2_3.t4 D2_3.t18 47.5387
R12406 D2_3.t11 D2_3.t25 47.5387
R12407 D2_3.t22 D2_3.t14 44.058
R12408 D2_3.t10 D2_3.t3 44.058
R12409 D2_3.n1 D2_3.t13 38.8649
R12410 D2_3.n0 D2_3.t0 38.8649
R12411 D2_3.n16 D2_3.t7 38.7949
R12412 D2_3.n15 D2_3.t12 38.7949
R12413 D2_3.n6 D2_3.t19 38.7949
R12414 D2_3.n5 D2_3.t24 38.7949
R12415 D2_3.n16 D2_3.n15 31.4949
R12416 D2_3.n6 D2_3.n5 31.4949
R12417 D2_3.t13 D2_3.t22 28.6791
R12418 D2_3.t0 D2_3.t10 28.6791
R12419 D2_3.n24 D2_3.n23 23.7262
R12420 D2_3.n17 D2_3.t23 17.9416
R12421 D2_3.n7 D2_3.t5 17.9416
R12422 D2_3.n18 D2_3.t4 16.621
R12423 D2_3.n4 D2_3.t11 16.621
R12424 D2_3.n24 D2_3.n12 16.3468
R12425 D2_3.n18 D2_3.t8 12.5148
R12426 D2_3.n4 D2_3.t17 12.5148
R12427 D2_3.n17 D2_3.t6 11.957
R12428 D2_3.n7 D2_3.t15 11.957
R12429 D2_3.n25 D2_3 9.59299
R12430 D2_3.n15 D2_3.t9 7.3005
R12431 D2_3.t23 D2_3.n16 7.3005
R12432 D2_3.n5 D2_3.t20 7.3005
R12433 D2_3.t5 D2_3.n6 7.3005
R12434 D2_3.n1 D2_3.t16 7.3005
R12435 D2_3.n0 D2_3.t1 7.3005
R12436 D2_3 D2_3.n17 5.95286
R12437 D2_3 D2_3.n7 5.95286
R12438 D2_3.n25 D2_3.n24 5.52808
R12439 D2_3 D2_3.n1 5.27587
R12440 D2_3 D2_3.n0 5.27587
R12441 D2_3 D2_3.n18 4.59246
R12442 D2_3 D2_3.n4 4.59246
R12443 D2_3.n14 D2_3.n13 4.5005
R12444 D2_3.n3 D2_3.n2 4.5005
R12445 D2_3.n9 D2_3.n3 3.46105
R12446 D2_3.n20 D2_3.n14 3.45513
R12447 D2_3.n21 D2_3.n20 2.25138
R12448 D2_3.n10 D2_3.n9 2.25138
R12449 D2_3.n27 D2_3.n25 2.2505
R12450 D2_3.n23 D2_3.n13 2.24334
R12451 D2_3.n12 D2_3.n2 2.24334
R12452 D2_3.n22 D2_3.n21 1.5081
R12453 D2_3.n11 D2_3.n10 1.5081
R12454 D2_3.n19 D2_3 1.4092
R12455 D2_3.n8 D2_3 1.25659
R12456 D2_3.n20 D2_3.n19 0.143896
R12457 D2_3.n19 D2_3 0.135578
R12458 D2_3.n8 D2_3 0.133622
R12459 D2_3.n9 D2_3.n8 0.0563228
R12460 D2_3.n27 D2_3.n26 0.0468409
R12461 D2_3 D2_3.n27 0.0339615
R12462 D2_3.n22 D2_3.n14 0.0312595
R12463 D2_3.n11 D2_3.n3 0.0312595
R12464 D2_3.n23 D2_3.n22 0.0174666
R12465 D2_3.n12 D2_3.n11 0.0174666
R12466 D2_3.n26 D2_3 0.0108063
R12467 D2_3.n26 D2_3 0.00911964
R12468 D2_3.n21 D2_3.n13 0.00176987
R12469 D2_3.n10 D2_3.n2 0.00176987
R12470 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n2 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t10 130.41
R12471 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n0 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t7 35.3186
R12472 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n3 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t8 33.5023
R12473 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t4 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n3 33.5023
R12474 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n1 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t11 32.2349
R12475 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n0 31.632
R12476 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n5 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t6 19.0118
R12477 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n4 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t4 16.3786
R12478 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t6 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n2 13.2317
R12479 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n2 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n1 13.0005
R12480 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n4 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t5 11.3259
R12481 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n1 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t3 11.146
R12482 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n0 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t12 7.3005
R12483 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n3 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t9 7.3005
R12484 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n9 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n7 5.47387
R12485 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n10 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n6 4.65398
R12486 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n9 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n8 4.2255
R12487 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n5 3.63228
R12488 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n5 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n4 3.62977
R12489 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n10 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n9 0.427022
R12490 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n10 0.257096
R12491 7b_counter_0.MDFF_0.QB.n6 7b_counter_0.MDFF_0.QB.t10 53.0716
R12492 7b_counter_0.MDFF_0.QB.t7 7b_counter_0.MDFF_0.QB.t6 44.058
R12493 7b_counter_0.MDFF_0.QB.n0 7b_counter_0.MDFF_0.QB.t9 38.8649
R12494 7b_counter_0.MDFF_0.QB.t9 7b_counter_0.MDFF_0.QB.t7 28.6791
R12495 7b_counter_0.MDFF_0.QB 7b_counter_0.MDFF_0.QB.n7 19.3781
R12496 7b_counter_0.MDFF_0.QB.n7 7b_counter_0.MDFF_0.QB.t8 17.2076
R12497 7b_counter_0.MDFF_0.QB.n7 7b_counter_0.MDFF_0.QB.t5 14.3398
R12498 7b_counter_0.MDFF_0.QB.n0 7b_counter_0.MDFF_0.QB.t4 7.3005
R12499 7b_counter_0.MDFF_0.QB.t5 7b_counter_0.MDFF_0.QB.n6 7.3005
R12500 7b_counter_0.MDFF_0.QB 7b_counter_0.MDFF_0.QB.n0 5.42008
R12501 7b_counter_0.MDFF_0.QB.n6 7b_counter_0.MDFF_0.QB.n5 4.51584
R12502 7b_counter_0.MDFF_0.QB.n5 7b_counter_0.MDFF_0.QB.n2 3.62007
R12503 7b_counter_0.MDFF_0.QB.n5 7b_counter_0.MDFF_0.QB.n4 3.15478
R12504 7b_counter_0.MDFF_0.QB.n4 7b_counter_0.MDFF_0.QB.t3 1.6255
R12505 7b_counter_0.MDFF_0.QB.n4 7b_counter_0.MDFF_0.QB.n3 1.6255
R12506 7b_counter_0.MDFF_0.QB.n2 7b_counter_0.MDFF_0.QB.t0 1.463
R12507 7b_counter_0.MDFF_0.QB.n2 7b_counter_0.MDFF_0.QB.n1 1.463
R12508 p2_gen_magic_0.xnor_magic_1.OUT.t5 p2_gen_magic_0.xnor_magic_1.OUT.t8 44.058
R12509 p2_gen_magic_0.xnor_magic_1.OUT.n3 p2_gen_magic_0.xnor_magic_1.OUT.t7 38.8649
R12510 p2_gen_magic_0.xnor_magic_1.OUT.n4 p2_gen_magic_0.xnor_magic_1.OUT 36.2792
R12511 p2_gen_magic_0.xnor_magic_1.OUT.t7 p2_gen_magic_0.xnor_magic_1.OUT.t5 28.6791
R12512 p2_gen_magic_0.xnor_magic_1.OUT.n3 p2_gen_magic_0.xnor_magic_1.OUT.t6 7.3005
R12513 p2_gen_magic_0.xnor_magic_1.OUT p2_gen_magic_0.xnor_magic_1.OUT.n3 5.27587
R12514 p2_gen_magic_0.xnor_magic_1.OUT.n4 p2_gen_magic_0.xnor_magic_1.OUT.n2 4.11572
R12515 p2_gen_magic_0.xnor_magic_1.OUT p2_gen_magic_0.xnor_magic_1.OUT.n4 3.61488
R12516 p2_gen_magic_0.xnor_magic_1.OUT p2_gen_magic_0.xnor_magic_1.OUT.t1 3.11311
R12517 p2_gen_magic_0.xnor_magic_1.OUT.t1 p2_gen_magic_0.xnor_magic_1.OUT.n0 1.6255
R12518 p2_gen_magic_0.xnor_magic_1.OUT.n2 p2_gen_magic_0.xnor_magic_1.OUT.t0 1.463
R12519 p2_gen_magic_0.xnor_magic_1.OUT.n2 p2_gen_magic_0.xnor_magic_1.OUT.n1 1.463
R12520 Q2.t26 Q2.t18 47.8944
R12521 Q2.t7 Q2.t28 47.8944
R12522 Q2.t27 Q2.t19 47.5387
R12523 Q2.t8 Q2.t29 47.5387
R12524 Q2.t30 Q2.t20 44.058
R12525 Q2.n29 Q2.t12 38.8649
R12526 Q2.n7 Q2.t22 38.7949
R12527 Q2.n6 Q2.t23 38.7949
R12528 Q2.n15 Q2.t4 38.7949
R12529 Q2.n14 Q2.t5 38.7949
R12530 Q2.n28 Q2.n3 35.6043
R12531 Q2.t13 Q2.t21 31.5469
R12532 Q2.t6 Q2.t13 31.5469
R12533 Q2.t17 Q2.t6 31.5469
R12534 Q2.t10 Q2.t17 31.5469
R12535 Q2.n7 Q2.n6 31.4949
R12536 Q2.n15 Q2.n14 31.4949
R12537 Q2 Q2.n30 30.7641
R12538 Q2.t25 Q2.t31 28.8094
R12539 Q2.t12 Q2.t30 28.6791
R12540 Q2.n28 Q2.n27 28.6095
R12541 Q2.n11 Q2.n10 18.7921
R12542 Q2.n8 Q2.t14 17.9416
R12543 Q2.n16 Q2.t24 17.9416
R12544 Q2.n2 Q2.t10 15.9693
R12545 Q2.n9 Q2.t27 15.7085
R12546 Q2.n17 Q2.t8 15.7085
R12547 Q2.n2 Q2.t25 15.5782
R12548 Q2.n9 Q2.t3 13.4273
R12549 Q2.n17 Q2.t11 13.4273
R12550 Q2.n8 Q2.t26 11.957
R12551 Q2.n16 Q2.t7 11.957
R12552 Q2.n6 Q2.t9 7.3005
R12553 Q2.t14 Q2.n7 7.3005
R12554 Q2.n14 Q2.t16 7.3005
R12555 Q2.t24 Q2.n15 7.3005
R12556 Q2.n29 Q2.t15 7.3005
R12557 Q2.n23 Q2.n22 6.3692
R12558 Q2 Q2.n8 5.94647
R12559 Q2 Q2.n16 5.94647
R12560 Q2.n0 Q2.t0 5.47387
R12561 Q2 Q2.n29 5.27587
R12562 Q2.n1 Q2.t1 4.65398
R12563 Q2.n27 Q2.n26 4.5005
R12564 Q2.n11 Q2.n4 4.5005
R12565 Q2.n0 Q2.t2 4.2255
R12566 Q2.n3 Q2.n2 4.13791
R12567 Q2 Q2.n9 4.08021
R12568 Q2 Q2.n17 4.08021
R12569 Q2.n18 Q2.n13 3.28431
R12570 Q2.n10 Q2 2.48458
R12571 Q2.n18 Q2 2.40514
R12572 Q2.n3 Q2 2.32782
R12573 Q2.n20 Q2.n12 2.25826
R12574 Q2.n20 Q2.n19 2.25494
R12575 Q2.n21 Q2.n13 2.25218
R12576 Q2.n26 Q2.n5 2.2512
R12577 Q2.n25 Q2.n4 2.2507
R12578 Q2.n22 Q2.n21 2.24442
R12579 Q2 Q2.n28 1.96301
R12580 Q2.n24 Q2.n23 0.90303
R12581 Q2.n10 Q2 0.550045
R12582 Q2.n1 Q2.n0 0.427022
R12583 Q2.n19 Q2.n18 0.394756
R12584 Q2.n19 Q2 0.278682
R12585 Q2 Q2.n1 0.257096
R12586 Q2.n23 Q2.n5 0.217822
R12587 Q2.n30 Q2 0.18746
R12588 Q2.n24 Q2.n11 0.0324737
R12589 Q2.n27 Q2.n4 0.0316538
R12590 Q2.n5 Q2.n4 0.0165783
R12591 Q2.n22 Q2.n12 0.0151461
R12592 Q2.n13 Q2.n12 0.0142134
R12593 Q2.n30 Q2 0.00286842
R12594 Q2.n21 Q2.n20 0.00165385
R12595 Q2.n25 Q2.n24 0.00159203
R12596 Q2.n26 Q2.n25 0.00159203
R12597 D2_6.t11 D2_6.t1 47.8944
R12598 D2_6.t4 D2_6.t20 47.8944
R12599 D2_6.t25 D2_6.t19 47.5387
R12600 D2_6.t15 D2_6.t9 47.5387
R12601 D2_6.t24 D2_6.t16 44.058
R12602 D2_6.t3 D2_6.t2 44.058
R12603 D2_6.n20 D2_6.t12 38.8649
R12604 D2_6.n16 D2_6.t21 38.8649
R12605 D2_6.n12 D2_6.t8 38.7949
R12606 D2_6.n11 D2_6.t6 38.7949
R12607 D2_6.n3 D2_6.t0 38.7949
R12608 D2_6.n2 D2_6.t23 38.7949
R12609 D2_6.n18 D2_6.n10 34.6483
R12610 D2_6.n12 D2_6.n11 31.4949
R12611 D2_6.n3 D2_6.n2 31.4949
R12612 D2_6.t12 D2_6.t24 28.6791
R12613 D2_6.t21 D2_6.t3 28.6791
R12614 D2_6.n13 D2_6.t22 17.9416
R12615 D2_6.n4 D2_6.t14 17.9416
R12616 D2_6.n14 D2_6.t25 16.621
R12617 D2_6.n5 D2_6.t15 16.621
R12618 D2_6.n17 D2_6.n15 12.6238
R12619 D2_6.n14 D2_6.t17 12.5148
R12620 D2_6.n5 D2_6.t7 12.5148
R12621 D2_6.n13 D2_6.t11 11.957
R12622 D2_6.n4 D2_6.t4 11.957
R12623 D2_6.n20 D2_6.t10 7.3005
R12624 D2_6.n11 D2_6.t13 7.3005
R12625 D2_6.t22 D2_6.n12 7.3005
R12626 D2_6.n16 D2_6.t18 7.3005
R12627 D2_6.n2 D2_6.t5 7.3005
R12628 D2_6.t14 D2_6.n3 7.3005
R12629 D2_6 D2_6.n13 5.95286
R12630 D2_6 D2_6.n4 5.95286
R12631 D2_6.n18 D2_6.n17 5.61009
R12632 D2_6 D2_6.n20 5.27587
R12633 D2_6 D2_6.n16 5.27587
R12634 D2_6 D2_6.n14 4.59246
R12635 D2_6 D2_6.n5 4.59246
R12636 D2_6.n10 D2_6.n9 4.5005
R12637 D2_6.n8 D2_6.n7 3.45141
R12638 D2_6.n19 D2_6.n18 2.70648
R12639 D2_6.n7 D2_6.n1 2.25138
R12640 D2_6.n9 D2_6.n8 2.24334
R12641 D2_6.n17 D2_6 1.88904
R12642 D2_6.n1 D2_6.n0 1.5081
R12643 D2_6.n15 D2_6 1.36028
R12644 D2_6.n6 D2_6 1.34267
R12645 D2_6.n7 D2_6.n6 0.284443
R12646 D2_6.n6 D2_6 0.2021
R12647 D2_6.n15 D2_6 0.184491
R12648 D2_6.n19 D2_6 0.0740348
R12649 D2_6 D2_6.n19 0.0339615
R12650 D2_6.n10 D2_6.n0 0.0312595
R12651 D2_6.n8 D2_6.n0 0.0174666
R12652 D2_6.n9 D2_6.n1 0.00176987
R12653 D2_1.t18 D2_1.t11 144.929
R12654 D2_1.n19 D2_1.n18 58.5348
R12655 D2_1.t28 D2_1.t21 47.8944
R12656 D2_1.t29 D2_1.t16 47.8944
R12657 D2_1.t13 D2_1.t0 47.5387
R12658 D2_1.t34 D2_1.t19 44.058
R12659 D2_1.t20 D2_1.t9 44.058
R12660 D2_1.t3 D2_1.t30 44.058
R12661 D2_1.n1 D2_1.t4 38.8649
R12662 D2_1.n0 D2_1.t23 38.8649
R12663 D2_1.n8 D2_1.t27 38.7949
R12664 D2_1.n7 D2_1.t15 38.7949
R12665 D2_1.n3 D2_1.t26 38.7949
R12666 D2_1.n2 D2_1.t14 38.7949
R12667 D2_1.n14 D2_1.t24 32.714
R12668 D2_1.n8 D2_1.n7 31.4949
R12669 D2_1.n3 D2_1.n2 31.4949
R12670 D2_1.t4 D2_1.t20 28.6791
R12671 D2_1.t23 D2_1.t3 28.6791
R12672 D2_1.n18 D2_1.n17 25.7355
R12673 D2_1.n15 D2_1.n14 21.0471
R12674 D2_1.n9 D2_1.t5 17.9416
R12675 D2_1.n4 D2_1.t12 17.9416
R12676 D2_1.n5 D2_1.t13 16.621
R12677 D2_1.t24 D2_1 16.2341
R12678 D2_1.n11 D2_1.n10 15.8172
R12679 D2_1.n12 D2_1.n11 15.8172
R12680 D2_1.n17 D2_1 15.5683
R12681 D2_1.n13 D2_1.t18 14.7309
R12682 D2_1.n16 D2_1.t33 14.5353
R12683 D2_1.n13 D2_1.t34 13.9487
R12684 D2_1.n5 D2_1.t35 12.5148
R12685 D2_1.n9 D2_1.t28 11.957
R12686 D2_1.n4 D2_1.t29 11.957
R12687 D2_1.n17 D2_1 11.8316
R12688 D2_1.n10 D2_1.t1 11.7326
R12689 D2_1.n10 D2_1.t8 11.7326
R12690 D2_1.n11 D2_1.t7 11.7326
R12691 D2_1.n11 D2_1.t22 11.7326
R12692 D2_1.n12 D2_1.t2 11.7326
R12693 D2_1.t33 D2_1.n12 11.7326
R12694 D2_1.n15 D2_1.t17 11.6675
R12695 D2_1 D2_1.n13 9.83788
R12696 D2_1.n14 D2_1.t6 7.3005
R12697 D2_1.n7 D2_1.t32 7.3005
R12698 D2_1.t5 D2_1.n8 7.3005
R12699 D2_1.n2 D2_1.t31 7.3005
R12700 D2_1.t12 D2_1.n3 7.3005
R12701 D2_1.n1 D2_1.t10 7.3005
R12702 D2_1.n0 D2_1.t25 7.3005
R12703 D2_1.n21 D2_1.n19 6.74408
R12704 D2_1 D2_1.n9 5.95286
R12705 D2_1 D2_1.n4 5.95286
R12706 D2_1 D2_1.n1 5.27587
R12707 D2_1 D2_1.n0 5.27587
R12708 D2_1.n19 D2_1 5.07595
R12709 D2_1 D2_1.n5 4.59246
R12710 D2_1 D2_1.n16 4.19616
R12711 D2_1.n18 D2_1.n6 2.68069
R12712 D2_1.n16 D2_1.n15 2.47729
R12713 D2_1.n6 D2_1 1.3505
R12714 D2_1.n6 D2_1 0.194274
R12715 D2_1.n21 D2_1.n20 0.0468336
R12716 D2_1 D2_1.n21 0.0339615
R12717 D2_1.n20 D2_1 0.0115019
R12718 D2_1.n20 D2_1 0.00541341
R12719 a_29512_8496.t17 a_29512_8496.n3 39.6673
R12720 a_29512_8496.n3 a_29512_8496.t9 39.6673
R12721 a_29512_8496.n4 a_29512_8496.t13 39.3349
R12722 a_29512_8496.t11 a_29512_8496.n4 39.3349
R12723 a_29512_8496.t9 a_29512_8496.t14 31.0255
R12724 a_29512_8496.t10 a_29512_8496.t16 31.0255
R12725 a_29512_8496.t12 a_29512_8496.t11 29.1353
R12726 a_29512_8496.n5 a_29512_8496.t17 13.6103
R12727 a_29512_8496.n5 a_29512_8496.t12 12.9295
R12728 a_29512_8496.n3 a_29512_8496.t10 7.3005
R12729 a_29512_8496.n4 a_29512_8496.t15 7.3005
R12730 a_29512_8496.n6 a_29512_8496.n5 4.42281
R12731 a_29512_8496.n12 a_29512_8496.n11 4.2255
R12732 a_29512_8496.n8 a_29512_8496.n7 2.92502
R12733 a_29512_8496.n15 a_29512_8496.n14 2.90967
R12734 a_29512_8496.n14 a_29512_8496.n13 2.88695
R12735 a_29512_8496.n7 a_29512_8496.n2 2.86115
R12736 a_29512_8496.n17 a_29512_8496.n16 2.6005
R12737 a_29512_8496.n1 a_29512_8496.t3 1.6255
R12738 a_29512_8496.n1 a_29512_8496.n0 1.6255
R12739 a_29512_8496.n17 a_29512_8496.t8 1.6255
R12740 a_29512_8496.n18 a_29512_8496.n17 1.6255
R12741 a_29512_8496.n10 a_29512_8496.t7 1.463
R12742 a_29512_8496.n10 a_29512_8496.n9 1.463
R12743 a_29512_8496.n15 a_29512_8496.n10 1.42678
R12744 a_29512_8496.n8 a_29512_8496.n1 1.23627
R12745 a_29512_8496.n16 a_29512_8496.n8 0.901117
R12746 a_29512_8496.n14 a_29512_8496.n12 0.812613
R12747 a_29512_8496.n16 a_29512_8496.n15 0.801537
R12748 a_29512_8496.n7 a_29512_8496.n6 0.402865
R12749 7b_counter_0.MDFF_5.LD.t20 7b_counter_0.MDFF_5.LD.t28 165.293
R12750 7b_counter_0.MDFF_5.LD.t82 7b_counter_0.MDFF_5.LD.t70 144.929
R12751 7b_counter_0.MDFF_5.LD.t61 7b_counter_0.MDFF_5.LD.t21 144.929
R12752 7b_counter_0.MDFF_5.LD.t83 7b_counter_0.MDFF_5.LD.t60 144.929
R12753 7b_counter_0.MDFF_5.LD.t68 7b_counter_0.MDFF_5.LD.t72 144.929
R12754 7b_counter_0.MDFF_5.LD.t11 7b_counter_0.MDFF_5.LD.t17 144.929
R12755 7b_counter_0.MDFF_5.LD.t31 7b_counter_0.MDFF_5.LD.t43 44.058
R12756 7b_counter_0.MDFF_5.LD.t15 7b_counter_0.MDFF_5.LD.t16 44.058
R12757 7b_counter_0.MDFF_5.LD.t32 7b_counter_0.MDFF_5.LD.t34 44.058
R12758 7b_counter_0.MDFF_5.LD.t19 7b_counter_0.MDFF_5.LD.t41 44.058
R12759 7b_counter_0.MDFF_5.LD.t36 7b_counter_0.MDFF_5.LD.t69 44.058
R12760 7b_counter_0.MDFF_5.LD.t59 7b_counter_0.MDFF_5.LD.t67 44.058
R12761 7b_counter_0.MDFF_5.LD.n53 7b_counter_0.MDFF_5.LD.n52 36.1331
R12762 7b_counter_0.MDFF_5.LD.n34 7b_counter_0.MDFF_5.LD.t24 32.714
R12763 7b_counter_0.MDFF_5.LD.n16 7b_counter_0.MDFF_5.LD.t12 32.714
R12764 7b_counter_0.MDFF_5.LD.n26 7b_counter_0.MDFF_5.LD.t25 32.714
R12765 7b_counter_0.MDFF_5.LD.n1 7b_counter_0.MDFF_5.LD.t13 32.714
R12766 7b_counter_0.MDFF_5.LD.n11 7b_counter_0.MDFF_5.LD.t26 32.714
R12767 7b_counter_0.MDFF_5.LD.n60 7b_counter_0.MDFF_5.LD.t42 32.714
R12768 7b_counter_0.MDFF_5.LD.n35 7b_counter_0.MDFF_5.LD.n34 21.0471
R12769 7b_counter_0.MDFF_5.LD.n17 7b_counter_0.MDFF_5.LD.n16 21.0471
R12770 7b_counter_0.MDFF_5.LD.n27 7b_counter_0.MDFF_5.LD.n26 21.0471
R12771 7b_counter_0.MDFF_5.LD.n2 7b_counter_0.MDFF_5.LD.n1 21.0471
R12772 7b_counter_0.MDFF_5.LD.n12 7b_counter_0.MDFF_5.LD.n11 21.0471
R12773 7b_counter_0.MDFF_5.LD.n61 7b_counter_0.MDFF_5.LD.n60 21.0471
R12774 7b_counter_0.MDFF_5.LD.t24 7b_counter_0.MDFF_5.LD 16.2341
R12775 7b_counter_0.MDFF_5.LD.t25 7b_counter_0.MDFF_5.LD 16.2341
R12776 7b_counter_0.MDFF_5.LD.t26 7b_counter_0.MDFF_5.LD 16.2328
R12777 7b_counter_0.MDFF_5.LD.t42 7b_counter_0.MDFF_5.LD 16.2328
R12778 7b_counter_0.MDFF_5.LD.t12 7b_counter_0.MDFF_5.LD 16.1689
R12779 7b_counter_0.MDFF_5.LD.t13 7b_counter_0.MDFF_5.LD 16.1676
R12780 7b_counter_0.MDFF_5.LD.n31 7b_counter_0.MDFF_5.LD.n30 15.8172
R12781 7b_counter_0.MDFF_5.LD.n32 7b_counter_0.MDFF_5.LD.n31 15.8172
R12782 7b_counter_0.MDFF_5.LD.n19 7b_counter_0.MDFF_5.LD.n18 15.8172
R12783 7b_counter_0.MDFF_5.LD.n20 7b_counter_0.MDFF_5.LD.n19 15.8172
R12784 7b_counter_0.MDFF_5.LD.n23 7b_counter_0.MDFF_5.LD.n22 15.8172
R12785 7b_counter_0.MDFF_5.LD.n24 7b_counter_0.MDFF_5.LD.n23 15.8172
R12786 7b_counter_0.MDFF_5.LD.n4 7b_counter_0.MDFF_5.LD.n3 15.8172
R12787 7b_counter_0.MDFF_5.LD.n5 7b_counter_0.MDFF_5.LD.n4 15.8172
R12788 7b_counter_0.MDFF_5.LD.n8 7b_counter_0.MDFF_5.LD.n7 15.8172
R12789 7b_counter_0.MDFF_5.LD.n9 7b_counter_0.MDFF_5.LD.n8 15.8172
R12790 7b_counter_0.MDFF_5.LD.n57 7b_counter_0.MDFF_5.LD.n56 15.8172
R12791 7b_counter_0.MDFF_5.LD.n58 7b_counter_0.MDFF_5.LD.n57 15.8172
R12792 7b_counter_0.MDFF_5.LD.n15 7b_counter_0.MDFF_5.LD.t61 14.796
R12793 7b_counter_0.MDFF_5.LD.n0 7b_counter_0.MDFF_5.LD.t68 14.796
R12794 7b_counter_0.MDFF_5.LD.n33 7b_counter_0.MDFF_5.LD.t82 14.7309
R12795 7b_counter_0.MDFF_5.LD.n25 7b_counter_0.MDFF_5.LD.t83 14.7309
R12796 7b_counter_0.MDFF_5.LD.n10 7b_counter_0.MDFF_5.LD.t11 14.7309
R12797 7b_counter_0.MDFF_5.LD.n59 7b_counter_0.MDFF_5.LD.t20 14.7309
R12798 7b_counter_0.MDFF_5.LD.n36 7b_counter_0.MDFF_5.LD.t84 14.5353
R12799 7b_counter_0.MDFF_5.LD.n28 7b_counter_0.MDFF_5.LD.t85 14.5353
R12800 7b_counter_0.MDFF_5.LD.n13 7b_counter_0.MDFF_5.LD.t55 14.5353
R12801 7b_counter_0.MDFF_5.LD.n62 7b_counter_0.MDFF_5.LD.t56 14.5353
R12802 7b_counter_0.MDFF_5.LD.n21 7b_counter_0.MDFF_5.LD.t77 14.4701
R12803 7b_counter_0.MDFF_5.LD.n6 7b_counter_0.MDFF_5.LD.t45 14.4701
R12804 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n55 14.4277
R12805 7b_counter_0.MDFF_5.LD.n33 7b_counter_0.MDFF_5.LD.t31 13.9487
R12806 7b_counter_0.MDFF_5.LD.n25 7b_counter_0.MDFF_5.LD.t32 13.9487
R12807 7b_counter_0.MDFF_5.LD.n10 7b_counter_0.MDFF_5.LD.t36 13.9487
R12808 7b_counter_0.MDFF_5.LD.n59 7b_counter_0.MDFF_5.LD.t59 13.9487
R12809 7b_counter_0.MDFF_5.LD.n15 7b_counter_0.MDFF_5.LD.t15 13.8835
R12810 7b_counter_0.MDFF_5.LD.n0 7b_counter_0.MDFF_5.LD.t19 13.8835
R12811 7b_counter_0.MDFF_5.LD.n53 7b_counter_0.MDFF_5.LD 13.7929
R12812 7b_counter_0.MDFF_5.LD.n30 7b_counter_0.MDFF_5.LD.t27 11.7326
R12813 7b_counter_0.MDFF_5.LD.n30 7b_counter_0.MDFF_5.LD.t57 11.7326
R12814 7b_counter_0.MDFF_5.LD.n31 7b_counter_0.MDFF_5.LD.t48 11.7326
R12815 7b_counter_0.MDFF_5.LD.n31 7b_counter_0.MDFF_5.LD.t80 11.7326
R12816 7b_counter_0.MDFF_5.LD.n32 7b_counter_0.MDFF_5.LD.t9 11.7326
R12817 7b_counter_0.MDFF_5.LD.t84 7b_counter_0.MDFF_5.LD.n32 11.7326
R12818 7b_counter_0.MDFF_5.LD.n18 7b_counter_0.MDFF_5.LD.t47 11.7326
R12819 7b_counter_0.MDFF_5.LD.n18 7b_counter_0.MDFF_5.LD.t40 11.7326
R12820 7b_counter_0.MDFF_5.LD.n19 7b_counter_0.MDFF_5.LD.t53 11.7326
R12821 7b_counter_0.MDFF_5.LD.n19 7b_counter_0.MDFF_5.LD.t49 11.7326
R12822 7b_counter_0.MDFF_5.LD.n20 7b_counter_0.MDFF_5.LD.t76 11.7326
R12823 7b_counter_0.MDFF_5.LD.t77 7b_counter_0.MDFF_5.LD.n20 11.7326
R12824 7b_counter_0.MDFF_5.LD.n22 7b_counter_0.MDFF_5.LD.t38 11.7326
R12825 7b_counter_0.MDFF_5.LD.n22 7b_counter_0.MDFF_5.LD.t58 11.7326
R12826 7b_counter_0.MDFF_5.LD.n23 7b_counter_0.MDFF_5.LD.t81 11.7326
R12827 7b_counter_0.MDFF_5.LD.n23 7b_counter_0.MDFF_5.LD.t66 11.7326
R12828 7b_counter_0.MDFF_5.LD.n24 7b_counter_0.MDFF_5.LD.t18 11.7326
R12829 7b_counter_0.MDFF_5.LD.t85 7b_counter_0.MDFF_5.LD.n24 11.7326
R12830 7b_counter_0.MDFF_5.LD.n3 7b_counter_0.MDFF_5.LD.t51 11.7326
R12831 7b_counter_0.MDFF_5.LD.n3 7b_counter_0.MDFF_5.LD.t44 11.7326
R12832 7b_counter_0.MDFF_5.LD.n4 7b_counter_0.MDFF_5.LD.t75 11.7326
R12833 7b_counter_0.MDFF_5.LD.n4 7b_counter_0.MDFF_5.LD.t73 11.7326
R12834 7b_counter_0.MDFF_5.LD.n5 7b_counter_0.MDFF_5.LD.t39 11.7326
R12835 7b_counter_0.MDFF_5.LD.t45 7b_counter_0.MDFF_5.LD.n5 11.7326
R12836 7b_counter_0.MDFF_5.LD.n7 7b_counter_0.MDFF_5.LD.t50 11.7326
R12837 7b_counter_0.MDFF_5.LD.n7 7b_counter_0.MDFF_5.LD.t62 11.7326
R12838 7b_counter_0.MDFF_5.LD.n8 7b_counter_0.MDFF_5.LD.t86 11.7326
R12839 7b_counter_0.MDFF_5.LD.n8 7b_counter_0.MDFF_5.LD.t78 11.7326
R12840 7b_counter_0.MDFF_5.LD.n9 7b_counter_0.MDFF_5.LD.t71 11.7326
R12841 7b_counter_0.MDFF_5.LD.t55 7b_counter_0.MDFF_5.LD.n9 11.7326
R12842 7b_counter_0.MDFF_5.LD.n56 7b_counter_0.MDFF_5.LD.t46 11.7326
R12843 7b_counter_0.MDFF_5.LD.n56 7b_counter_0.MDFF_5.LD.t74 11.7326
R12844 7b_counter_0.MDFF_5.LD.n57 7b_counter_0.MDFF_5.LD.t35 11.7326
R12845 7b_counter_0.MDFF_5.LD.n57 7b_counter_0.MDFF_5.LD.t65 11.7326
R12846 7b_counter_0.MDFF_5.LD.n58 7b_counter_0.MDFF_5.LD.t79 11.7326
R12847 7b_counter_0.MDFF_5.LD.t56 7b_counter_0.MDFF_5.LD.n58 11.7326
R12848 7b_counter_0.MDFF_5.LD.n35 7b_counter_0.MDFF_5.LD.t63 11.6675
R12849 7b_counter_0.MDFF_5.LD.n17 7b_counter_0.MDFF_5.LD.t37 11.6675
R12850 7b_counter_0.MDFF_5.LD.n27 7b_counter_0.MDFF_5.LD.t64 11.6675
R12851 7b_counter_0.MDFF_5.LD.n2 7b_counter_0.MDFF_5.LD.t10 11.6675
R12852 7b_counter_0.MDFF_5.LD.n12 7b_counter_0.MDFF_5.LD.t22 11.6675
R12853 7b_counter_0.MDFF_5.LD.n61 7b_counter_0.MDFF_5.LD.t23 11.6675
R12854 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n33 9.83788
R12855 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n15 9.83788
R12856 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n25 9.83788
R12857 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n0 9.83788
R12858 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n10 9.83788
R12859 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n59 9.83788
R12860 7b_counter_0.MDFF_5.LD.n34 7b_counter_0.MDFF_5.LD.t54 7.3005
R12861 7b_counter_0.MDFF_5.LD.n16 7b_counter_0.MDFF_5.LD.t14 7.3005
R12862 7b_counter_0.MDFF_5.LD.n26 7b_counter_0.MDFF_5.LD.t30 7.3005
R12863 7b_counter_0.MDFF_5.LD.n1 7b_counter_0.MDFF_5.LD.t33 7.3005
R12864 7b_counter_0.MDFF_5.LD.n11 7b_counter_0.MDFF_5.LD.t52 7.3005
R12865 7b_counter_0.MDFF_5.LD.n60 7b_counter_0.MDFF_5.LD.t29 7.3005
R12866 7b_counter_0.MDFF_5.LD.n43 7b_counter_0.MDFF_5.LD.n37 4.2255
R12867 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n6 4.19721
R12868 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n13 4.19721
R12869 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n62 4.19721
R12870 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n36 4.19616
R12871 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n21 4.19616
R12872 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n28 4.19616
R12873 7b_counter_0.MDFF_5.LD.n51 7b_counter_0.MDFF_5.LD.n50 2.92992
R12874 7b_counter_0.MDFF_5.LD.n42 7b_counter_0.MDFF_5.LD.n41 2.90652
R12875 7b_counter_0.MDFF_5.LD.n42 7b_counter_0.MDFF_5.LD.n38 2.89193
R12876 7b_counter_0.MDFF_5.LD.n51 7b_counter_0.MDFF_5.LD.n44 2.85689
R12877 7b_counter_0.MDFF_5.LD.n49 7b_counter_0.MDFF_5.LD.n48 2.6005
R12878 7b_counter_0.MDFF_5.LD.n21 7b_counter_0.MDFF_5.LD.n17 2.54246
R12879 7b_counter_0.MDFF_5.LD.n6 7b_counter_0.MDFF_5.LD.n2 2.54246
R12880 7b_counter_0.MDFF_5.LD.n36 7b_counter_0.MDFF_5.LD.n35 2.47729
R12881 7b_counter_0.MDFF_5.LD.n28 7b_counter_0.MDFF_5.LD.n27 2.47729
R12882 7b_counter_0.MDFF_5.LD.n13 7b_counter_0.MDFF_5.LD.n12 2.47729
R12883 7b_counter_0.MDFF_5.LD.n62 7b_counter_0.MDFF_5.LD.n61 2.47729
R12884 7b_counter_0.MDFF_5.LD.n29 7b_counter_0.MDFF_5.LD 1.93071
R12885 7b_counter_0.MDFF_5.LD.n14 7b_counter_0.MDFF_5.LD 1.93071
R12886 7b_counter_0.MDFF_5.LD.n48 7b_counter_0.MDFF_5.LD.t4 1.6255
R12887 7b_counter_0.MDFF_5.LD.n48 7b_counter_0.MDFF_5.LD.n47 1.6255
R12888 7b_counter_0.MDFF_5.LD.n46 7b_counter_0.MDFF_5.LD.t7 1.6255
R12889 7b_counter_0.MDFF_5.LD.n46 7b_counter_0.MDFF_5.LD.n45 1.6255
R12890 7b_counter_0.MDFF_5.LD.n40 7b_counter_0.MDFF_5.LD.t0 1.463
R12891 7b_counter_0.MDFF_5.LD.n40 7b_counter_0.MDFF_5.LD.n39 1.463
R12892 7b_counter_0.MDFF_5.LD.n41 7b_counter_0.MDFF_5.LD.n40 1.43
R12893 7b_counter_0.MDFF_5.LD.n50 7b_counter_0.MDFF_5.LD.n46 1.23128
R12894 7b_counter_0.MDFF_5.LD.n54 7b_counter_0.MDFF_5.LD.n29 1.09582
R12895 7b_counter_0.MDFF_5.LD.n55 7b_counter_0.MDFF_5.LD.n14 1.09582
R12896 7b_counter_0.MDFF_5.LD.n50 7b_counter_0.MDFF_5.LD.n49 0.922675
R12897 7b_counter_0.MDFF_5.LD.n43 7b_counter_0.MDFF_5.LD.n42 0.789247
R12898 7b_counter_0.MDFF_5.LD.n54 7b_counter_0.MDFF_5.LD.n53 0.572499
R12899 7b_counter_0.MDFF_5.LD.n52 7b_counter_0.MDFF_5.LD.n51 0.456126
R12900 7b_counter_0.MDFF_5.LD.n52 7b_counter_0.MDFF_5.LD.n43 0.374196
R12901 7b_counter_0.MDFF_5.LD.n55 7b_counter_0.MDFF_5.LD.n54 0.26284
R12902 7b_counter_0.MDFF_5.LD.n29 7b_counter_0.MDFF_5.LD 0.181929
R12903 7b_counter_0.MDFF_5.LD.n14 7b_counter_0.MDFF_5.LD 0.1805
R12904 D2_2.t8 D2_2.t23 47.8944
R12905 D2_2.t16 D2_2.t3 47.8944
R12906 D2_2.t25 D2_2.t20 47.5387
R12907 D2_2.t9 D2_2.t1 47.5387
R12908 D2_2.t17 D2_2.t10 44.058
R12909 D2_2.t21 D2_2.t19 44.058
R12910 D2_2.n20 D2_2.t2 38.8649
R12911 D2_2.n0 D2_2.t12 38.8649
R12912 D2_2.n4 D2_2.t7 38.7949
R12913 D2_2.n3 D2_2.t5 38.7949
R12914 D2_2.n13 D2_2.t18 38.7949
R12915 D2_2.n12 D2_2.t15 38.7949
R12916 D2_2.n4 D2_2.n3 31.4949
R12917 D2_2.n13 D2_2.n12 31.4949
R12918 D2_2.t2 D2_2.t17 28.6791
R12919 D2_2.t12 D2_2.t21 28.6791
R12920 D2_2.n5 D2_2.t24 17.9416
R12921 D2_2.n14 D2_2.t6 17.9416
R12922 D2_2.n6 D2_2.t25 16.621
R12923 D2_2.n15 D2_2.t9 16.621
R12924 D2_2.n18 D2_2.n17 15.5756
R12925 D2_2.n6 D2_2.t4 12.5148
R12926 D2_2.n15 D2_2.t14 12.5148
R12927 D2_2.n5 D2_2.t8 11.957
R12928 D2_2.n14 D2_2.t16 11.957
R12929 D2_2.n17 D2_2.n11 9.32108
R12930 D2_2.n20 D2_2.t0 7.3005
R12931 D2_2.n3 D2_2.t13 7.3005
R12932 D2_2.t24 D2_2.n4 7.3005
R12933 D2_2.n12 D2_2.t22 7.3005
R12934 D2_2.t6 D2_2.n13 7.3005
R12935 D2_2.n0 D2_2.t11 7.3005
R12936 D2_2 D2_2.n5 5.95286
R12937 D2_2 D2_2.n14 5.95286
R12938 D2_2.n17 D2_2.n16 5.82172
R12939 D2_2.n19 D2_2.n18 5.72846
R12940 D2_2 D2_2.n20 5.27587
R12941 D2_2 D2_2.n0 5.27587
R12942 D2_2.n18 D2_2 4.76002
R12943 D2_2 D2_2.n6 4.59246
R12944 D2_2 D2_2.n15 4.59246
R12945 D2_2.n2 D2_2.n1 4.5005
R12946 D2_2.n8 D2_2.n2 3.49286
R12947 D2_2.n9 D2_2.n8 2.25138
R12948 D2_2.n11 D2_2.n1 2.24334
R12949 D2_2.n10 D2_2.n9 1.5081
R12950 D2_2.n16 D2_2 1.36924
R12951 D2_2.n7 D2_2 1.36028
R12952 D2_2.n8 D2_2.n7 0.204548
R12953 D2_2.n7 D2_2 0.184491
R12954 D2_2.n16 D2_2 0.108743
R12955 D2_2.n19 D2_2 0.0738303
R12956 D2_2 D2_2.n19 0.0339615
R12957 D2_2.n10 D2_2.n2 0.0312595
R12958 D2_2.n11 D2_2.n10 0.0174666
R12959 D2_2.n9 D2_2.n1 0.00176987
R12960 LD.t26 LD.t55 144.929
R12961 LD.t23 LD.t54 144.929
R12962 LD.t86 LD.t27 144.929
R12963 LD.t34 LD.t58 144.929
R12964 LD.t18 LD.t50 144.929
R12965 LD.t79 LD.t21 144.929
R12966 LD.n23 LD.n22 50.8638
R12967 LD.t59 LD.t33 44.058
R12968 LD.t63 LD.t39 44.058
R12969 LD.t47 LD.t15 44.058
R12970 LD.t61 LD.t36 44.058
R12971 LD.t62 LD.t35 44.058
R12972 LD.t43 LD.t14 44.058
R12973 LD.n35 LD.n34 32.8505
R12974 LD.n36 LD.n35 32.8505
R12975 LD.n59 LD.n58 32.8505
R12976 LD.n60 LD.n59 32.8505
R12977 LD.n4 LD.t60 32.714
R12978 LD.n25 LD.t41 32.714
R12979 LD.n32 LD.t51 32.714
R12980 LD.n43 LD.t46 32.714
R12981 LD.n48 LD.t32 32.714
R12982 LD.n56 LD.t45 32.714
R12983 LD.n5 LD.n4 21.0471
R12984 LD.n26 LD.n25 21.0471
R12985 LD.n33 LD.n32 21.0471
R12986 LD.n44 LD.n43 21.0471
R12987 LD.n49 LD.n48 21.0471
R12988 LD.n57 LD.n56 21.0471
R12989 LD.t60 LD 16.2341
R12990 LD.t46 LD 16.2341
R12991 LD.t41 LD 16.1689
R12992 LD.t51 LD 16.1689
R12993 LD.t32 LD 16.1689
R12994 LD.t45 LD 16.1689
R12995 LD.n1 LD.n0 15.8172
R12996 LD.n2 LD.n1 15.8172
R12997 LD.n28 LD.n27 15.8172
R12998 LD.n29 LD.n28 15.8172
R12999 LD.n40 LD.n39 15.8172
R13000 LD.n41 LD.n40 15.8172
R13001 LD.n51 LD.n50 15.8172
R13002 LD.n52 LD.n51 15.8172
R13003 LD.n38 LD 15.616
R13004 LD.n24 LD.t23 14.796
R13005 LD.n31 LD.t86 14.796
R13006 LD.n47 LD.t18 14.796
R13007 LD.n55 LD.t79 14.796
R13008 LD.n3 LD.t26 14.7309
R13009 LD.n42 LD.t34 14.7309
R13010 LD.n6 LD.t38 14.5353
R13011 LD.n45 LD.t17 14.5353
R13012 LD.n30 LD.t52 14.4701
R13013 LD.n37 LD.t37 14.4701
R13014 LD.n53 LD.t48 14.4701
R13015 LD.n61 LD.t28 14.4701
R13016 LD.n3 LD.t59 13.9487
R13017 LD.n42 LD.t61 13.9487
R13018 LD.n24 LD.t63 13.8835
R13019 LD.n31 LD.t47 13.8835
R13020 LD.n47 LD.t62 13.8835
R13021 LD.n55 LD.t43 13.8835
R13022 LD.n54 LD 13.8333
R13023 LD.n0 LD.t24 11.7326
R13024 LD.n0 LD.t84 11.7326
R13025 LD.n1 LD.t49 11.7326
R13026 LD.n1 LD.t30 11.7326
R13027 LD.n2 LD.t80 11.7326
R13028 LD.t38 LD.n2 11.7326
R13029 LD.n27 LD.t74 11.7326
R13030 LD.n27 LD.t13 11.7326
R13031 LD.n28 LD.t19 11.7326
R13032 LD.n28 LD.t57 11.7326
R13033 LD.n29 LD.t44 11.7326
R13034 LD.t52 LD.n29 11.7326
R13035 LD.n39 LD.t85 11.7326
R13036 LD.n39 LD.t68 11.7326
R13037 LD.n40 LD.t31 11.7326
R13038 LD.n40 LD.t11 11.7326
R13039 LD.n41 LD.t40 11.7326
R13040 LD.t17 LD.n41 11.7326
R13041 LD.n50 LD.t70 11.7326
R13042 LD.n50 LD.t69 11.7326
R13043 LD.n51 LD.t16 11.7326
R13044 LD.n51 LD.t12 11.7326
R13045 LD.n52 LD.t42 11.7326
R13046 LD.t48 LD.n52 11.7326
R13047 LD.n5 LD.t10 11.6675
R13048 LD.n26 LD.t9 11.6675
R13049 LD.n33 LD.t75 11.6675
R13050 LD.n44 LD.t72 11.6675
R13051 LD.n49 LD.t81 11.6675
R13052 LD.n57 LD.t71 11.6675
R13053 LD.n36 LD.t53 10.1684
R13054 LD.n34 LD.t77 10.1684
R13055 LD.n34 LD.t83 10.1684
R13056 LD.n35 LD.t65 10.1684
R13057 LD.n35 LD.t29 10.1684
R13058 LD.t37 LD.n36 10.1684
R13059 LD.n60 LD.t25 10.1684
R13060 LD.n58 LD.t76 10.1684
R13061 LD.n58 LD.t78 10.1684
R13062 LD.n59 LD.t20 10.1684
R13063 LD.n59 LD.t22 10.1684
R13064 LD.t28 LD.n60 10.1684
R13065 LD LD.n3 9.83788
R13066 LD LD.n24 9.83788
R13067 LD LD.n31 9.83788
R13068 LD LD.n42 9.83788
R13069 LD LD.n47 9.83788
R13070 LD LD.n55 9.83788
R13071 LD.n4 LD.t82 7.3005
R13072 LD.n25 LD.t64 7.3005
R13073 LD.n32 LD.t73 7.3005
R13074 LD.n43 LD.t67 7.3005
R13075 LD.n48 LD.t56 7.3005
R13076 LD.n56 LD.t66 7.3005
R13077 LD.n21 LD.n9 4.2255
R13078 LD LD.n6 4.19616
R13079 LD LD.n30 4.19616
R13080 LD LD.n37 4.19616
R13081 LD LD.n45 4.19616
R13082 LD LD.n53 4.19616
R13083 LD LD.n61 4.19616
R13084 LD.n46 LD 4.02178
R13085 LD.n15 LD.n8 2.93105
R13086 LD.n20 LD.n19 2.90828
R13087 LD.n20 LD.n10 2.8925
R13088 LD.n8 LD.n7 2.85689
R13089 LD.n18 LD.n17 2.6005
R13090 LD.n30 LD.n26 2.54246
R13091 LD.n37 LD.n33 2.54246
R13092 LD.n53 LD.n49 2.54246
R13093 LD.n61 LD.n57 2.54246
R13094 LD.n6 LD.n5 2.47729
R13095 LD.n45 LD.n44 2.47729
R13096 LD LD.n38 1.93071
R13097 LD LD.n62 1.93071
R13098 LD.n54 LD.n46 1.92305
R13099 LD.n62 LD.n54 1.78327
R13100 LD.n17 LD.t3 1.6255
R13101 LD.n17 LD.n16 1.6255
R13102 LD.n14 LD.t7 1.6255
R13103 LD.n14 LD.n13 1.6255
R13104 LD.n12 LD.t2 1.463
R13105 LD.n12 LD.n11 1.463
R13106 LD.n19 LD.n12 1.42943
R13107 LD.n15 LD.n14 1.23144
R13108 LD.n18 LD.n15 0.922765
R13109 LD.n19 LD.n18 0.789247
R13110 LD.n21 LD.n20 0.788516
R13111 LD LD.n23 0.643813
R13112 LD.n22 LD.n8 0.456126
R13113 LD.n22 LD.n21 0.374196
R13114 LD.n23 LD 0.193357
R13115 LD.n38 LD 0.181929
R13116 LD.n46 LD 0.181929
R13117 LD.n62 LD 0.181929
R13118 D2_7.t12 D2_7.t2 47.8944
R13119 D2_7.t18 D2_7.t8 47.8944
R13120 D2_7.t4 D2_7.t16 47.5387
R13121 D2_7.t10 D2_7.t25 47.5387
R13122 D2_7.t1 D2_7.t24 44.058
R13123 D2_7.t0 D2_7.t22 44.058
R13124 D2_7.n1 D2_7.t13 38.8649
R13125 D2_7.n0 D2_7.t15 38.8649
R13126 D2_7.n4 D2_7.t3 38.7949
R13127 D2_7.n3 D2_7.t6 38.7949
R13128 D2_7.n8 D2_7.t11 38.7949
R13129 D2_7.n7 D2_7.t14 38.7949
R13130 D2_7.n4 D2_7.n3 31.4949
R13131 D2_7.n8 D2_7.n7 31.4949
R13132 D2_7.t13 D2_7.t1 28.6791
R13133 D2_7.t15 D2_7.t0 28.6791
R13134 D2_7.n12 D2_7.n6 27.9087
R13135 D2_7.n13 D2_7.n12 20.4279
R13136 D2_7.n5 D2_7.t21 17.9416
R13137 D2_7.n9 D2_7.t7 17.9416
R13138 D2_7.n2 D2_7.t4 16.621
R13139 D2_7.n10 D2_7.t10 16.621
R13140 D2_7.n2 D2_7.t19 12.5148
R13141 D2_7.n10 D2_7.t5 12.5148
R13142 D2_7.n5 D2_7.t12 11.957
R13143 D2_7.n9 D2_7.t18 11.957
R13144 D2_7.n12 D2_7.n11 9.33041
R13145 D2_7.n13 D2_7 9.23901
R13146 D2_7.n3 D2_7.t9 7.3005
R13147 D2_7.t21 D2_7.n4 7.3005
R13148 D2_7.n7 D2_7.t17 7.3005
R13149 D2_7.t7 D2_7.n8 7.3005
R13150 D2_7.n1 D2_7.t20 7.3005
R13151 D2_7.n0 D2_7.t23 7.3005
R13152 D2_7 D2_7.n5 5.95286
R13153 D2_7 D2_7.n9 5.95286
R13154 D2_7 D2_7.n1 5.27587
R13155 D2_7 D2_7.n0 5.27587
R13156 D2_7 D2_7.n2 4.59246
R13157 D2_7 D2_7.n10 4.59246
R13158 D2_7.n14 D2_7.n13 1.56771
R13159 D2_7.n11 D2_7 1.3818
R13160 D2_7.n6 D2_7 1.31528
R13161 D2_7.n11 D2_7 0.16297
R13162 D2_7.n6 D2_7 0.137535
R13163 D2_7 D2_7.n14 0.113121
R13164 D2_7.n14 D2_7 0.00367207
R13165 mux_magic_0.IN2.t5 mux_magic_0.IN2.t8 47.8944
R13166 mux_magic_0.IN2.t6 mux_magic_0.IN2.t11 44.058
R13167 mux_magic_0.IN2.n0 mux_magic_0.IN2.t10 38.8649
R13168 mux_magic_0.IN2.n1 mux_magic_0.IN2.t7 38.7949
R13169 mux_magic_0.IN2.n2 mux_magic_0.IN2.t9 38.7949
R13170 mux_magic_0.IN2.n2 mux_magic_0.IN2.n1 31.4949
R13171 mux_magic_0.IN2.t10 mux_magic_0.IN2.t6 28.6791
R13172 mux_magic_0.IN2.n3 mux_magic_0.IN2.t12 17.9416
R13173 mux_magic_0.IN2.n3 mux_magic_0.IN2.t5 11.957
R13174 mux_magic_0.IN2.n4 mux_magic_0.IN2 8.98052
R13175 mux_magic_0.IN2.n1 mux_magic_0.IN2.t13 7.3005
R13176 mux_magic_0.IN2.t12 mux_magic_0.IN2.n2 7.3005
R13177 mux_magic_0.IN2.n0 mux_magic_0.IN2.t14 7.3005
R13178 mux_magic_0.IN2 mux_magic_0.IN2.n3 5.86241
R13179 mux_magic_0.IN2 mux_magic_0.IN2.n0 5.47416
R13180 mux_magic_0.IN2.t4 mux_magic_0.IN2.t3 3.31072
R13181 mux_magic_0.IN2.t3 mux_magic_0.IN2.n5 1.6255
R13182 mux_magic_0.IN2.n4 mux_magic_0.IN2 1.25072
R13183 mux_magic_0.IN2 mux_magic_0.IN2.n4 0.642239
R13184 mux_magic_0.IN2 mux_magic_0.IN2.t4 0.583625
R13185 7b_counter_0.DFF_magic_0.Q.t13 7b_counter_0.DFF_magic_0.Q.t16 47.8944
R13186 7b_counter_0.DFF_magic_0.Q.t10 7b_counter_0.DFF_magic_0.Q.t21 47.8944
R13187 7b_counter_0.DFF_magic_0.Q.n7 7b_counter_0.DFF_magic_0.Q.t11 38.7949
R13188 7b_counter_0.DFF_magic_0.Q.n8 7b_counter_0.DFF_magic_0.Q.t19 38.7949
R13189 7b_counter_0.DFF_magic_0.Q.n1 7b_counter_0.DFF_magic_0.Q.t18 38.7949
R13190 7b_counter_0.DFF_magic_0.Q.n0 7b_counter_0.DFF_magic_0.Q.t15 38.7949
R13191 7b_counter_0.DFF_magic_0.Q.n3 7b_counter_0.DFF_magic_0.Q.t7 31.9191
R13192 7b_counter_0.DFF_magic_0.Q.n8 7b_counter_0.DFF_magic_0.Q.n7 31.4949
R13193 7b_counter_0.DFF_magic_0.Q.n1 7b_counter_0.DFF_magic_0.Q.n0 31.4949
R13194 7b_counter_0.DFF_magic_0.Q.n4 7b_counter_0.DFF_magic_0.Q.t14 31.1267
R13195 7b_counter_0.DFF_magic_0.Q.n10 7b_counter_0.DFF_magic_0.Q.n6 19.1157
R13196 7b_counter_0.DFF_magic_0.Q.n9 7b_counter_0.DFF_magic_0.Q.t8 17.9416
R13197 7b_counter_0.DFF_magic_0.Q.n2 7b_counter_0.DFF_magic_0.Q.t6 17.9416
R13198 7b_counter_0.DFF_magic_0.Q.n9 7b_counter_0.DFF_magic_0.Q.t13 11.957
R13199 7b_counter_0.DFF_magic_0.Q.n2 7b_counter_0.DFF_magic_0.Q.t10 11.957
R13200 7b_counter_0.DFF_magic_0.Q.n4 7b_counter_0.DFF_magic_0.Q.t12 10.9505
R13201 7b_counter_0.DFF_magic_0.Q.n3 7b_counter_0.DFF_magic_0.Q.t20 10.3639
R13202 7b_counter_0.DFF_magic_0.Q.n5 7b_counter_0.DFF_magic_0.Q.n3 10.1032
R13203 7b_counter_0.DFF_magic_0.Q.n6 7b_counter_0.DFF_magic_0.Q 7.60603
R13204 7b_counter_0.DFF_magic_0.Q.n7 7b_counter_0.DFF_magic_0.Q.t9 7.3005
R13205 7b_counter_0.DFF_magic_0.Q.t8 7b_counter_0.DFF_magic_0.Q.n8 7.3005
R13206 7b_counter_0.DFF_magic_0.Q.n0 7b_counter_0.DFF_magic_0.Q.t17 7.3005
R13207 7b_counter_0.DFF_magic_0.Q.t6 7b_counter_0.DFF_magic_0.Q.n1 7.3005
R13208 7b_counter_0.DFF_magic_0.Q 7b_counter_0.DFF_magic_0.Q.n2 5.96162
R13209 7b_counter_0.DFF_magic_0.Q 7b_counter_0.DFF_magic_0.Q.n9 5.86241
R13210 7b_counter_0.DFF_magic_0.Q.n5 7b_counter_0.DFF_magic_0.Q.n4 4.75854
R13211 7b_counter_0.DFF_magic_0.Q 7b_counter_0.DFF_magic_0.Q.n5 4.22152
R13212 7b_counter_0.DFF_magic_0.Q.n15 7b_counter_0.DFF_magic_0.Q.n12 3.6455
R13213 7b_counter_0.DFF_magic_0.Q.n15 7b_counter_0.DFF_magic_0.Q.n14 3.31072
R13214 7b_counter_0.DFF_magic_0.Q.n18 7b_counter_0.DFF_magic_0.Q.n17 2.90572
R13215 7b_counter_0.DFF_magic_0.Q.n6 7b_counter_0.DFF_magic_0.Q 2.29941
R13216 7b_counter_0.DFF_magic_0.Q.n14 7b_counter_0.DFF_magic_0.Q.t3 1.6255
R13217 7b_counter_0.DFF_magic_0.Q.n14 7b_counter_0.DFF_magic_0.Q.n13 1.6255
R13218 7b_counter_0.DFF_magic_0.Q.n17 7b_counter_0.DFF_magic_0.Q.t5 1.6255
R13219 7b_counter_0.DFF_magic_0.Q.n17 7b_counter_0.DFF_magic_0.Q.n16 1.6255
R13220 7b_counter_0.DFF_magic_0.Q.n12 7b_counter_0.DFF_magic_0.Q.t1 1.463
R13221 7b_counter_0.DFF_magic_0.Q.n12 7b_counter_0.DFF_magic_0.Q.n11 1.463
R13222 7b_counter_0.DFF_magic_0.Q.n10 7b_counter_0.DFF_magic_0.Q 1.25072
R13223 7b_counter_0.DFF_magic_0.Q 7b_counter_0.DFF_magic_0.Q.n10 0.642239
R13224 7b_counter_0.DFF_magic_0.Q.n18 7b_counter_0.DFF_magic_0.Q.n15 0.4055
R13225 7b_counter_0.DFF_magic_0.Q 7b_counter_0.DFF_magic_0.Q.n18 0.178625
R13226 DFF_magic_0.D.t35 DFF_magic_0.D.n15 39.8579
R13227 DFF_magic_0.D.n15 DFF_magic_0.D.t26 39.8579
R13228 DFF_magic_0.D.t25 DFF_magic_0.D.n11 39.8579
R13229 DFF_magic_0.D.n11 DFF_magic_0.D.t13 39.8579
R13230 DFF_magic_0.D.t33 DFF_magic_0.D.n7 39.8579
R13231 DFF_magic_0.D.n7 DFF_magic_0.D.t29 39.8579
R13232 DFF_magic_0.D.n16 DFF_magic_0.D.t11 39.3349
R13233 DFF_magic_0.D.t23 DFF_magic_0.D.n16 39.3349
R13234 DFF_magic_0.D.n12 DFF_magic_0.D.t27 39.3349
R13235 DFF_magic_0.D.t9 DFF_magic_0.D.n12 39.3349
R13236 DFF_magic_0.D.n8 DFF_magic_0.D.t15 39.3349
R13237 DFF_magic_0.D.t19 DFF_magic_0.D.n8 39.3349
R13238 DFF_magic_0.D.t26 DFF_magic_0.D.t12 31.0255
R13239 DFF_magic_0.D.t34 DFF_magic_0.D.t22 31.0255
R13240 DFF_magic_0.D.t13 DFF_magic_0.D.t28 31.0255
R13241 DFF_magic_0.D.t14 DFF_magic_0.D.t31 31.0255
R13242 DFF_magic_0.D.t29 DFF_magic_0.D.t16 31.0255
R13243 DFF_magic_0.D.t32 DFF_magic_0.D.t18 31.0255
R13244 DFF_magic_0.D.t24 DFF_magic_0.D.t23 29.1353
R13245 DFF_magic_0.D.t10 DFF_magic_0.D.t9 29.1353
R13246 DFF_magic_0.D.t20 DFF_magic_0.D.t19 29.1353
R13247 DFF_magic_0.D.n10 DFF_magic_0.D 27.3045
R13248 DFF_magic_0.D.n17 DFF_magic_0.D.t35 13.5376
R13249 DFF_magic_0.D.n13 DFF_magic_0.D.t25 13.5376
R13250 DFF_magic_0.D.n9 DFF_magic_0.D.t33 13.5376
R13251 DFF_magic_0.D.n17 DFF_magic_0.D.t24 12.5549
R13252 DFF_magic_0.D.n13 DFF_magic_0.D.t10 12.5549
R13253 DFF_magic_0.D.n9 DFF_magic_0.D.t20 12.5549
R13254 DFF_magic_0.D.n15 DFF_magic_0.D.t34 7.3005
R13255 DFF_magic_0.D.n16 DFF_magic_0.D.t21 7.3005
R13256 DFF_magic_0.D.n11 DFF_magic_0.D.t14 7.3005
R13257 DFF_magic_0.D.n12 DFF_magic_0.D.t30 7.3005
R13258 DFF_magic_0.D.n7 DFF_magic_0.D.t32 7.3005
R13259 DFF_magic_0.D.n8 DFF_magic_0.D.t17 7.3005
R13260 DFF_magic_0.D.n10 DFF_magic_0.D.n9 5.73946
R13261 DFF_magic_0.D.n2 DFF_magic_0.D.t0 5.68507
R13262 DFF_magic_0.D.n14 DFF_magic_0.D.n13 5.6754
R13263 DFF_magic_0.D.n6 DFF_magic_0.D.t6 4.928
R13264 DFF_magic_0.D.n18 DFF_magic_0.D.n17 3.62559
R13265 DFF_magic_0.D DFF_magic_0.D.n18 3.5586
R13266 DFF_magic_0.D.n5 DFF_magic_0.D.n4 3.1505
R13267 DFF_magic_0.D.n2 DFF_magic_0.D.n1 2.6005
R13268 DFF_magic_0.D.n18 DFF_magic_0.D.n14 2.54453
R13269 DFF_magic_0.D.n14 DFF_magic_0.D.n10 2.36537
R13270 DFF_magic_0.D.n1 DFF_magic_0.D.t1 1.6255
R13271 DFF_magic_0.D.n1 DFF_magic_0.D.n0 1.6255
R13272 DFF_magic_0.D.n4 DFF_magic_0.D.t7 1.463
R13273 DFF_magic_0.D.n4 DFF_magic_0.D.n3 1.463
R13274 DFF_magic_0.D.n6 DFF_magic_0.D.n5 1.16072
R13275 DFF_magic_0.D.n5 DFF_magic_0.D.n2 0.898543
R13276 DFF_magic_0.D DFF_magic_0.D.n6 0.291602
R13277 Q1.t5 Q1.t23 47.8944
R13278 Q1.t24 Q1.t15 47.8944
R13279 Q1.t6 Q1.t28 47.5387
R13280 Q1.t25 Q1.t19 47.5387
R13281 Q1.t8 Q1.t26 44.058
R13282 Q1.n37 Q1.t16 38.8649
R13283 Q1.n13 Q1.t29 38.7949
R13284 Q1.n12 Q1.t30 38.7949
R13285 Q1.n20 Q1.t17 38.7949
R13286 Q1.n19 Q1.t20 38.7949
R13287 Q1.t7 Q1.t13 31.5469
R13288 Q1.t27 Q1.t7 31.5469
R13289 Q1.t10 Q1.t27 31.5469
R13290 Q1.t4 Q1.t10 31.5469
R13291 Q1.t18 Q1.t4 31.5469
R13292 Q1.n13 Q1.n12 31.4949
R13293 Q1.n20 Q1.n19 31.4949
R13294 Q1.n40 Q1.n38 28.7686
R13295 Q1.t16 Q1.t8 28.6791
R13296 Q1.n42 Q1.n36 21.8018
R13297 Q1.n14 Q1.t22 17.9416
R13298 Q1.n21 Q1.t11 17.9416
R13299 Q1.n31 Q1.t6 15.7085
R13300 Q1.n22 Q1.t25 15.7085
R13301 Q1.n6 Q1.t18 15.2523
R13302 Q1.n28 Q1.n27 14.3627
R13303 Q1.n6 Q1.t21 13.5576
R13304 Q1.n31 Q1.t9 13.4273
R13305 Q1.n22 Q1.t31 13.4273
R13306 Q1.n14 Q1.t5 11.957
R13307 Q1.n21 Q1.t24 11.957
R13308 Q1.n37 Q1.t12 7.3005
R13309 Q1.n12 Q1.t14 7.3005
R13310 Q1.t22 Q1.n13 7.3005
R13311 Q1.n19 Q1.t3 7.3005
R13312 Q1.t11 Q1.n20 7.3005
R13313 Q1 Q1.n14 5.94647
R13314 Q1 Q1.n21 5.94647
R13315 Q1.n3 Q1.n2 5.47387
R13316 Q1 Q1.n37 5.27587
R13317 Q1.n4 Q1.n0 4.65398
R13318 Q1.n18 Q1.n17 4.5005
R13319 Q1.n28 Q1.n15 4.5005
R13320 Q1.n41 Q1.n8 4.5005
R13321 Q1.n42 Q1.n41 4.5005
R13322 Q1.n39 Q1.n7 4.5005
R13323 Q1.n41 Q1.n9 4.5005
R13324 Q1.n3 Q1.n1 4.2255
R13325 Q1 Q1.n6 4.10124
R13326 Q1 Q1.n31 4.08021
R13327 Q1 Q1.n22 4.08021
R13328 Q1.n45 Q1.n44 3.38735
R13329 Q1.n23 Q1.n18 3.25748
R13330 Q1.n32 Q1 2.46385
R13331 Q1.n44 Q1.n43 2.33504
R13332 Q1.n23 Q1 2.3324
R13333 Q1.n30 Q1.n29 2.25926
R13334 Q1.n34 Q1.n10 2.25826
R13335 Q1.n40 Q1.n39 2.25825
R13336 Q1.n34 Q1.n33 2.25808
R13337 Q1.n35 Q1.n11 2.25252
R13338 Q1.n25 Q1.n24 2.25138
R13339 Q1.n32 Q1.n30 2.2505
R13340 Q1.n27 Q1.n17 2.24528
R13341 Q1.n36 Q1.n35 2.24475
R13342 Q1.n26 Q1.n25 1.5081
R13343 Q1.n16 Q1.n15 1.4988
R13344 Q1 Q1.n45 0.8075
R13345 Q1.n43 Q1.n8 0.626519
R13346 Q1.n24 Q1 0.46057
R13347 Q1.n45 Q1 0.454173
R13348 Q1.n4 Q1.n3 0.427022
R13349 Q1.n24 Q1.n23 0.260825
R13350 Q1.n33 Q1 0.259591
R13351 Q1 Q1.n4 0.257096
R13352 Q1.n33 Q1.n32 0.229763
R13353 Q1.n16 Q1.n11 0.212131
R13354 Q1.n38 Q1 0.18935
R13355 Q1.n5 Q1 0.186245
R13356 Q1.n44 Q1.n7 0.121611
R13357 Q1 Q1.n5 0.0995
R13358 Q1.n41 Q1.n7 0.0316111
R13359 Q1.n29 Q1.n28 0.0255515
R13360 Q1.n39 Q1.n8 0.0255515
R13361 Q1.n26 Q1.n18 0.0234245
R13362 Q1.n43 Q1.n42 0.0209124
R13363 Q1.n36 Q1.n10 0.0144188
R13364 Q1.n5 Q1 0.0139043
R13365 Q1.n11 Q1.n10 0.0135342
R13366 Q1.n27 Q1.n26 0.0132822
R13367 Q1.n29 Q1.n16 0.010624
R13368 Q1.n43 Q1.n9 0.00513918
R13369 Q1.n25 Q1.n17 0.00176987
R13370 Q1.n38 Q1 0.00166883
R13371 Q1.n30 Q1.n15 0.00165385
R13372 Q1.n35 Q1.n34 0.00165385
R13373 Q1.n41 Q1.n40 0.00161111
R13374 Q1.n39 Q1.n9 0.00142783
R13375 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n5 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t6 130.41
R13376 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n7 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t7 35.3186
R13377 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n2 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t5 33.5023
R13378 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t12 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n2 33.5023
R13379 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n4 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t11 32.2349
R13380 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n7 31.543
R13381 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n6 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t9 18.9789
R13382 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n3 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t12 16.3786
R13383 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t9 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n5 13.2317
R13384 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n5 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n4 13.0005
R13385 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n3 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t8 11.3259
R13386 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n4 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t10 11.146
R13387 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n2 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t4 7.3005
R13388 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n7 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t3 7.3005
R13389 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n0 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t0 5.47387
R13390 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n1 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t1 4.65398
R13391 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n0 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t2 4.2255
R13392 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n6 3.66281
R13393 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n6 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n3 3.63303
R13394 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n1 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n0 0.427022
R13395 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n1 0.257096
R13396 p3_gen_magic_0.P3.t15 p3_gen_magic_0.P3.t11 47.8944
R13397 p3_gen_magic_0.P3.t16 p3_gen_magic_0.P3.t12 44.6331
R13398 p3_gen_magic_0.P3.t7 p3_gen_magic_0.P3.t16 43.4094
R13399 p3_gen_magic_0.P3.n0 p3_gen_magic_0.P3.t10 38.7949
R13400 p3_gen_magic_0.P3.n1 p3_gen_magic_0.P3.t8 38.7949
R13401 p3_gen_magic_0.P3.t13 p3_gen_magic_0.P3.t7 31.5469
R13402 p3_gen_magic_0.P3.n1 p3_gen_magic_0.P3.n0 31.4949
R13403 p3_gen_magic_0.P3.n2 p3_gen_magic_0.P3.t14 17.9416
R13404 p3_gen_magic_0.P3.n3 p3_gen_magic_0.P3.t13 15.0567
R13405 p3_gen_magic_0.P3.n3 p3_gen_magic_0.P3.t6 13.6228
R13406 p3_gen_magic_0.P3.n2 p3_gen_magic_0.P3.t15 11.957
R13407 p3_gen_magic_0.P3.n0 p3_gen_magic_0.P3.t9 7.3005
R13408 p3_gen_magic_0.P3.t14 p3_gen_magic_0.P3.n1 7.3005
R13409 p3_gen_magic_0.P3 p3_gen_magic_0.P3.n2 5.86241
R13410 p3_gen_magic_0.P3 p3_gen_magic_0.P3.n3 4.2675
R13411 p3_gen_magic_0.P3.n9 p3_gen_magic_0.P3.n6 3.6455
R13412 p3_gen_magic_0.P3.n9 p3_gen_magic_0.P3.n8 3.31072
R13413 p3_gen_magic_0.P3.n12 p3_gen_magic_0.P3.n11 2.90572
R13414 p3_gen_magic_0.P3.n8 p3_gen_magic_0.P3.t3 1.6255
R13415 p3_gen_magic_0.P3.n8 p3_gen_magic_0.P3.n7 1.6255
R13416 p3_gen_magic_0.P3.n11 p3_gen_magic_0.P3.t5 1.6255
R13417 p3_gen_magic_0.P3.n11 p3_gen_magic_0.P3.n10 1.6255
R13418 p3_gen_magic_0.P3.n6 p3_gen_magic_0.P3.t1 1.463
R13419 p3_gen_magic_0.P3.n6 p3_gen_magic_0.P3.n5 1.463
R13420 p3_gen_magic_0.P3.n4 p3_gen_magic_0.P3 1.24289
R13421 p3_gen_magic_0.P3 p3_gen_magic_0.P3.n4 0.634257
R13422 p3_gen_magic_0.P3.n12 p3_gen_magic_0.P3.n9 0.4055
R13423 p3_gen_magic_0.P3 p3_gen_magic_0.P3.n12 0.178625
R13424 p3_gen_magic_0.P3.n4 p3_gen_magic_0.P3 0.1319
R13425 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t14 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t12 47.8944
R13426 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n7 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t13 38.7949
R13427 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n8 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t15 38.7949
R13428 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n8 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n7 31.4949
R13429 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n9 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t17 17.9416
R13430 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n9 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t14 11.957
R13431 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n7 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t16 7.3005
R13432 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t17 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n8 7.3005
R13433 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n10 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN 5.93058
R13434 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n9 5.86474
R13435 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n2 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t10 5.68507
R13436 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n6 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t0 4.92604
R13437 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n15 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n12 3.6455
R13438 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n15 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n14 3.31072
R13439 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n5 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n4 3.1505
R13440 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n18 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n17 2.90572
R13441 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n2 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n1 2.6005
R13442 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n10 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN 1.88467
R13443 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n1 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t11 1.6255
R13444 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n1 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n0 1.6255
R13445 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n14 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t6 1.6255
R13446 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n14 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n13 1.6255
R13447 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n17 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t7 1.6255
R13448 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n17 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n16 1.6255
R13449 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n4 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t2 1.463
R13450 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n4 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n3 1.463
R13451 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n12 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.t4 1.463
R13452 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n12 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n11 1.463
R13453 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n10 1.33598
R13454 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n6 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n5 1.15166
R13455 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n5 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n2 0.898543
R13456 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n18 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n15 0.4055
R13457 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n6 0.198522
R13458 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN.n18 0.178625
R13459 7b_counter_0.MDFF_4.LD.t62 7b_counter_0.MDFF_4.LD.t37 165.293
R13460 7b_counter_0.MDFF_4.LD.t89 7b_counter_0.MDFF_4.LD.t102 165.293
R13461 7b_counter_0.MDFF_4.LD.t31 7b_counter_0.MDFF_4.LD.t38 144.929
R13462 7b_counter_0.MDFF_4.LD.t63 7b_counter_0.MDFF_4.LD.t19 144.929
R13463 7b_counter_0.MDFF_4.LD.t20 7b_counter_0.MDFF_4.LD.t92 144.929
R13464 7b_counter_0.MDFF_4.LD.t66 7b_counter_0.MDFF_4.LD.t78 144.929
R13465 7b_counter_0.MDFF_4.LD.t119 7b_counter_0.MDFF_4.LD.t73 144.929
R13466 7b_counter_0.MDFF_4.LD.t34 7b_counter_0.MDFF_4.LD.t71 144.929
R13467 7b_counter_0.MDFF_4.LD.t70 7b_counter_0.MDFF_4.LD.t114 144.929
R13468 7b_counter_0.MDFF_4.LD.n60 7b_counter_0.MDFF_4.LD.t110 44.4466
R13469 7b_counter_0.MDFF_4.LD.t77 7b_counter_0.MDFF_4.LD.t117 44.058
R13470 7b_counter_0.MDFF_4.LD.t97 7b_counter_0.MDFF_4.LD.t118 44.058
R13471 7b_counter_0.MDFF_4.LD.t98 7b_counter_0.MDFF_4.LD.t100 44.058
R13472 7b_counter_0.MDFF_4.LD.t67 7b_counter_0.MDFF_4.LD.t72 44.058
R13473 7b_counter_0.MDFF_4.LD.t125 7b_counter_0.MDFF_4.LD.t21 44.058
R13474 7b_counter_0.MDFF_4.LD.t107 7b_counter_0.MDFF_4.LD.t30 44.058
R13475 7b_counter_0.MDFF_4.LD.t56 7b_counter_0.MDFF_4.LD.t88 44.058
R13476 7b_counter_0.MDFF_4.LD.t84 7b_counter_0.MDFF_4.LD.t121 44.058
R13477 7b_counter_0.MDFF_4.LD.t111 7b_counter_0.MDFF_4.LD.t33 44.058
R13478 7b_counter_0.MDFF_4.LD.n0 7b_counter_0.MDFF_4.LD 40.6939
R13479 7b_counter_0.MDFF_4.LD.n61 7b_counter_0.MDFF_4.LD.n60 34.2788
R13480 7b_counter_0.MDFF_4.LD.n64 7b_counter_0.MDFF_4.LD.n63 32.8505
R13481 7b_counter_0.MDFF_4.LD.n63 7b_counter_0.MDFF_4.LD.n62 32.8505
R13482 7b_counter_0.MDFF_4.LD.n28 7b_counter_0.MDFF_4.LD.t95 32.714
R13483 7b_counter_0.MDFF_4.LD.n35 7b_counter_0.MDFF_4.LD.t96 32.714
R13484 7b_counter_0.MDFF_4.LD.n39 7b_counter_0.MDFF_4.LD.t106 32.714
R13485 7b_counter_0.MDFF_4.LD.n49 7b_counter_0.MDFF_4.LD.t122 32.714
R13486 7b_counter_0.MDFF_4.LD.n56 7b_counter_0.MDFF_4.LD.t101 32.714
R13487 7b_counter_0.MDFF_4.LD.n11 7b_counter_0.MDFF_4.LD.t112 32.714
R13488 7b_counter_0.MDFF_4.LD.n18 7b_counter_0.MDFF_4.LD.t27 32.714
R13489 7b_counter_0.MDFF_4.LD.n7 7b_counter_0.MDFF_4.LD.t11 32.714
R13490 7b_counter_0.MDFF_4.LD.n29 7b_counter_0.MDFF_4.LD.n28 21.0471
R13491 7b_counter_0.MDFF_4.LD.n36 7b_counter_0.MDFF_4.LD.n35 21.0471
R13492 7b_counter_0.MDFF_4.LD.n40 7b_counter_0.MDFF_4.LD.n39 21.0471
R13493 7b_counter_0.MDFF_4.LD.n50 7b_counter_0.MDFF_4.LD.n49 21.0471
R13494 7b_counter_0.MDFF_4.LD.n57 7b_counter_0.MDFF_4.LD.n56 21.0471
R13495 7b_counter_0.MDFF_4.LD.n12 7b_counter_0.MDFF_4.LD.n11 21.0471
R13496 7b_counter_0.MDFF_4.LD.n19 7b_counter_0.MDFF_4.LD.n18 21.0471
R13497 7b_counter_0.MDFF_4.LD.n8 7b_counter_0.MDFF_4.LD.n7 21.0471
R13498 7b_counter_0.MDFF_4.LD.n0 7b_counter_0.MDFF_4.LD.n1 20.2647
R13499 7b_counter_0.MDFF_4.LD.t95 7b_counter_0.MDFF_4.LD 16.2341
R13500 7b_counter_0.MDFF_4.LD.t96 7b_counter_0.MDFF_4.LD 16.2341
R13501 7b_counter_0.MDFF_4.LD.t122 7b_counter_0.MDFF_4.LD 16.2328
R13502 7b_counter_0.MDFF_4.LD.t101 7b_counter_0.MDFF_4.LD 16.2328
R13503 7b_counter_0.MDFF_4.LD.t11 7b_counter_0.MDFF_4.LD 16.2328
R13504 7b_counter_0.MDFF_4.LD.t106 7b_counter_0.MDFF_4.LD 16.1689
R13505 7b_counter_0.MDFF_4.LD.t110 7b_counter_0.MDFF_4.LD 16.1676
R13506 7b_counter_0.MDFF_4.LD.t112 7b_counter_0.MDFF_4.LD 16.1676
R13507 7b_counter_0.MDFF_4.LD.t27 7b_counter_0.MDFF_4.LD 16.1676
R13508 7b_counter_0.MDFF_4.LD.n25 7b_counter_0.MDFF_4.LD.n24 15.8172
R13509 7b_counter_0.MDFF_4.LD.n26 7b_counter_0.MDFF_4.LD.n25 15.8172
R13510 7b_counter_0.MDFF_4.LD.n32 7b_counter_0.MDFF_4.LD.n31 15.8172
R13511 7b_counter_0.MDFF_4.LD.n33 7b_counter_0.MDFF_4.LD.n32 15.8172
R13512 7b_counter_0.MDFF_4.LD.n42 7b_counter_0.MDFF_4.LD.n41 15.8172
R13513 7b_counter_0.MDFF_4.LD.n43 7b_counter_0.MDFF_4.LD.n42 15.8172
R13514 7b_counter_0.MDFF_4.LD.n46 7b_counter_0.MDFF_4.LD.n45 15.8172
R13515 7b_counter_0.MDFF_4.LD.n47 7b_counter_0.MDFF_4.LD.n46 15.8172
R13516 7b_counter_0.MDFF_4.LD.n53 7b_counter_0.MDFF_4.LD.n52 15.8172
R13517 7b_counter_0.MDFF_4.LD.n54 7b_counter_0.MDFF_4.LD.n53 15.8172
R13518 7b_counter_0.MDFF_4.LD.n14 7b_counter_0.MDFF_4.LD.n13 15.8172
R13519 7b_counter_0.MDFF_4.LD.n15 7b_counter_0.MDFF_4.LD.n14 15.8172
R13520 7b_counter_0.MDFF_4.LD.n21 7b_counter_0.MDFF_4.LD.n20 15.8172
R13521 7b_counter_0.MDFF_4.LD.n22 7b_counter_0.MDFF_4.LD.n21 15.8172
R13522 7b_counter_0.MDFF_4.LD.n4 7b_counter_0.MDFF_4.LD.n3 15.8172
R13523 7b_counter_0.MDFF_4.LD.n5 7b_counter_0.MDFF_4.LD.n4 15.8172
R13524 7b_counter_0.MDFF_4.LD.n59 7b_counter_0.MDFF_4.LD.t31 14.796
R13525 7b_counter_0.MDFF_4.LD.n38 7b_counter_0.MDFF_4.LD.t20 14.796
R13526 7b_counter_0.MDFF_4.LD.n10 7b_counter_0.MDFF_4.LD.t119 14.796
R13527 7b_counter_0.MDFF_4.LD.n17 7b_counter_0.MDFF_4.LD.t34 14.796
R13528 7b_counter_0.MDFF_4.LD.n27 7b_counter_0.MDFF_4.LD.t62 14.7309
R13529 7b_counter_0.MDFF_4.LD.n34 7b_counter_0.MDFF_4.LD.t63 14.7309
R13530 7b_counter_0.MDFF_4.LD.n48 7b_counter_0.MDFF_4.LD.t89 14.7309
R13531 7b_counter_0.MDFF_4.LD.n55 7b_counter_0.MDFF_4.LD.t66 14.7309
R13532 7b_counter_0.MDFF_4.LD.n6 7b_counter_0.MDFF_4.LD.t70 14.7309
R13533 7b_counter_0.MDFF_4.LD.n30 7b_counter_0.MDFF_4.LD.t64 14.5353
R13534 7b_counter_0.MDFF_4.LD.n37 7b_counter_0.MDFF_4.LD.t65 14.5353
R13535 7b_counter_0.MDFF_4.LD.n51 7b_counter_0.MDFF_4.LD.t15 14.5353
R13536 7b_counter_0.MDFF_4.LD.n58 7b_counter_0.MDFF_4.LD.t14 14.5353
R13537 7b_counter_0.MDFF_4.LD.n9 7b_counter_0.MDFF_4.LD.t22 14.5353
R13538 7b_counter_0.MDFF_4.LD.n65 7b_counter_0.MDFF_4.LD.t39 14.4701
R13539 7b_counter_0.MDFF_4.LD.n44 7b_counter_0.MDFF_4.LD.t85 14.4701
R13540 7b_counter_0.MDFF_4.LD.n16 7b_counter_0.MDFF_4.LD.t47 14.4701
R13541 7b_counter_0.MDFF_4.LD.n23 7b_counter_0.MDFF_4.LD.t46 14.4701
R13542 7b_counter_0.MDFF_4.LD.n27 7b_counter_0.MDFF_4.LD.t97 13.9487
R13543 7b_counter_0.MDFF_4.LD.n34 7b_counter_0.MDFF_4.LD.t98 13.9487
R13544 7b_counter_0.MDFF_4.LD.n48 7b_counter_0.MDFF_4.LD.t125 13.9487
R13545 7b_counter_0.MDFF_4.LD.n55 7b_counter_0.MDFF_4.LD.t107 13.9487
R13546 7b_counter_0.MDFF_4.LD.n6 7b_counter_0.MDFF_4.LD.t111 13.9487
R13547 7b_counter_0.MDFF_4.LD.n59 7b_counter_0.MDFF_4.LD.t77 13.8835
R13548 7b_counter_0.MDFF_4.LD.n38 7b_counter_0.MDFF_4.LD.t67 13.8835
R13549 7b_counter_0.MDFF_4.LD.n10 7b_counter_0.MDFF_4.LD.t56 13.8835
R13550 7b_counter_0.MDFF_4.LD.n17 7b_counter_0.MDFF_4.LD.t84 13.8835
R13551 7b_counter_0.MDFF_4.LD.n24 7b_counter_0.MDFF_4.LD.t44 11.7326
R13552 7b_counter_0.MDFF_4.LD.n24 7b_counter_0.MDFF_4.LD.t16 11.7326
R13553 7b_counter_0.MDFF_4.LD.n25 7b_counter_0.MDFF_4.LD.t83 11.7326
R13554 7b_counter_0.MDFF_4.LD.n25 7b_counter_0.MDFF_4.LD.t61 11.7326
R13555 7b_counter_0.MDFF_4.LD.n26 7b_counter_0.MDFF_4.LD.t86 11.7326
R13556 7b_counter_0.MDFF_4.LD.t64 7b_counter_0.MDFF_4.LD.n26 11.7326
R13557 7b_counter_0.MDFF_4.LD.n31 7b_counter_0.MDFF_4.LD.t45 11.7326
R13558 7b_counter_0.MDFF_4.LD.n31 7b_counter_0.MDFF_4.LD.t17 11.7326
R13559 7b_counter_0.MDFF_4.LD.n32 7b_counter_0.MDFF_4.LD.t55 11.7326
R13560 7b_counter_0.MDFF_4.LD.n32 7b_counter_0.MDFF_4.LD.t29 11.7326
R13561 7b_counter_0.MDFF_4.LD.n33 7b_counter_0.MDFF_4.LD.t87 11.7326
R13562 7b_counter_0.MDFF_4.LD.t65 7b_counter_0.MDFF_4.LD.n33 11.7326
R13563 7b_counter_0.MDFF_4.LD.n41 7b_counter_0.MDFF_4.LD.t40 11.7326
R13564 7b_counter_0.MDFF_4.LD.n41 7b_counter_0.MDFF_4.LD.t76 11.7326
R13565 7b_counter_0.MDFF_4.LD.n42 7b_counter_0.MDFF_4.LD.t53 11.7326
R13566 7b_counter_0.MDFF_4.LD.n42 7b_counter_0.MDFF_4.LD.t59 11.7326
R13567 7b_counter_0.MDFF_4.LD.n43 7b_counter_0.MDFF_4.LD.t32 11.7326
R13568 7b_counter_0.MDFF_4.LD.t85 7b_counter_0.MDFF_4.LD.n43 11.7326
R13569 7b_counter_0.MDFF_4.LD.n45 7b_counter_0.MDFF_4.LD.t68 11.7326
R13570 7b_counter_0.MDFF_4.LD.n45 7b_counter_0.MDFF_4.LD.t41 11.7326
R13571 7b_counter_0.MDFF_4.LD.n46 7b_counter_0.MDFF_4.LD.t54 11.7326
R13572 7b_counter_0.MDFF_4.LD.n46 7b_counter_0.MDFF_4.LD.t28 11.7326
R13573 7b_counter_0.MDFF_4.LD.n47 7b_counter_0.MDFF_4.LD.t43 11.7326
R13574 7b_counter_0.MDFF_4.LD.t15 7b_counter_0.MDFF_4.LD.n47 11.7326
R13575 7b_counter_0.MDFF_4.LD.n52 7b_counter_0.MDFF_4.LD.t51 11.7326
R13576 7b_counter_0.MDFF_4.LD.n52 7b_counter_0.MDFF_4.LD.t23 11.7326
R13577 7b_counter_0.MDFF_4.LD.n53 7b_counter_0.MDFF_4.LD.t81 11.7326
R13578 7b_counter_0.MDFF_4.LD.n53 7b_counter_0.MDFF_4.LD.t58 11.7326
R13579 7b_counter_0.MDFF_4.LD.n54 7b_counter_0.MDFF_4.LD.t42 11.7326
R13580 7b_counter_0.MDFF_4.LD.t14 7b_counter_0.MDFF_4.LD.n54 11.7326
R13581 7b_counter_0.MDFF_4.LD.n13 7b_counter_0.MDFF_4.LD.t52 11.7326
R13582 7b_counter_0.MDFF_4.LD.n13 7b_counter_0.MDFF_4.LD.t90 11.7326
R13583 7b_counter_0.MDFF_4.LD.n14 7b_counter_0.MDFF_4.LD.t57 11.7326
R13584 7b_counter_0.MDFF_4.LD.n14 7b_counter_0.MDFF_4.LD.t115 11.7326
R13585 7b_counter_0.MDFF_4.LD.n15 7b_counter_0.MDFF_4.LD.t18 11.7326
R13586 7b_counter_0.MDFF_4.LD.t47 7b_counter_0.MDFF_4.LD.n15 11.7326
R13587 7b_counter_0.MDFF_4.LD.n20 7b_counter_0.MDFF_4.LD.t80 11.7326
R13588 7b_counter_0.MDFF_4.LD.n20 7b_counter_0.MDFF_4.LD.t69 11.7326
R13589 7b_counter_0.MDFF_4.LD.n21 7b_counter_0.MDFF_4.LD.t74 11.7326
R13590 7b_counter_0.MDFF_4.LD.n21 7b_counter_0.MDFF_4.LD.t91 11.7326
R13591 7b_counter_0.MDFF_4.LD.n22 7b_counter_0.MDFF_4.LD.t120 11.7326
R13592 7b_counter_0.MDFF_4.LD.t46 7b_counter_0.MDFF_4.LD.n22 11.7326
R13593 7b_counter_0.MDFF_4.LD.n3 7b_counter_0.MDFF_4.LD.t82 11.7326
R13594 7b_counter_0.MDFF_4.LD.n3 7b_counter_0.MDFF_4.LD.t60 11.7326
R13595 7b_counter_0.MDFF_4.LD.n4 7b_counter_0.MDFF_4.LD.t75 11.7326
R13596 7b_counter_0.MDFF_4.LD.n4 7b_counter_0.MDFF_4.LD.t48 11.7326
R13597 7b_counter_0.MDFF_4.LD.n5 7b_counter_0.MDFF_4.LD.t49 11.7326
R13598 7b_counter_0.MDFF_4.LD.t22 7b_counter_0.MDFF_4.LD.n5 11.7326
R13599 7b_counter_0.MDFF_4.LD.n29 7b_counter_0.MDFF_4.LD.t24 11.6675
R13600 7b_counter_0.MDFF_4.LD.n36 7b_counter_0.MDFF_4.LD.t26 11.6675
R13601 7b_counter_0.MDFF_4.LD.n40 7b_counter_0.MDFF_4.LD.t35 11.6675
R13602 7b_counter_0.MDFF_4.LD.n50 7b_counter_0.MDFF_4.LD.t94 11.6675
R13603 7b_counter_0.MDFF_4.LD.n57 7b_counter_0.MDFF_4.LD.t93 11.6675
R13604 7b_counter_0.MDFF_4.LD.n12 7b_counter_0.MDFF_4.LD.t109 11.6675
R13605 7b_counter_0.MDFF_4.LD.n19 7b_counter_0.MDFF_4.LD.t108 11.6675
R13606 7b_counter_0.MDFF_4.LD.n8 7b_counter_0.MDFF_4.LD.t99 11.6675
R13607 7b_counter_0.MDFF_4.LD.n61 7b_counter_0.MDFF_4.LD.t104 10.1684
R13608 7b_counter_0.MDFF_4.LD.n60 7b_counter_0.MDFF_4.LD.t25 10.1684
R13609 7b_counter_0.MDFF_4.LD.n64 7b_counter_0.MDFF_4.LD.t36 10.1684
R13610 7b_counter_0.MDFF_4.LD.n63 7b_counter_0.MDFF_4.LD.t123 10.1684
R13611 7b_counter_0.MDFF_4.LD.n63 7b_counter_0.MDFF_4.LD.t79 10.1684
R13612 7b_counter_0.MDFF_4.LD.n62 7b_counter_0.MDFF_4.LD.t9 10.1684
R13613 7b_counter_0.MDFF_4.LD.n62 7b_counter_0.MDFF_4.LD.t50 10.1684
R13614 7b_counter_0.MDFF_4.LD.t39 7b_counter_0.MDFF_4.LD.n64 10.1684
R13615 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n59 9.83788
R13616 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n27 9.83788
R13617 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n34 9.83788
R13618 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n38 9.83788
R13619 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n48 9.83788
R13620 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n55 9.83788
R13621 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n10 9.83788
R13622 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n17 9.83788
R13623 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n6 9.83788
R13624 7b_counter_0.MDFF_4.LD.n28 7b_counter_0.MDFF_4.LD.t12 7.3005
R13625 7b_counter_0.MDFF_4.LD.n35 7b_counter_0.MDFF_4.LD.t105 7.3005
R13626 7b_counter_0.MDFF_4.LD.n39 7b_counter_0.MDFF_4.LD.t113 7.3005
R13627 7b_counter_0.MDFF_4.LD.n49 7b_counter_0.MDFF_4.LD.t103 7.3005
R13628 7b_counter_0.MDFF_4.LD.n56 7b_counter_0.MDFF_4.LD.t10 7.3005
R13629 7b_counter_0.MDFF_4.LD.n11 7b_counter_0.MDFF_4.LD.t116 7.3005
R13630 7b_counter_0.MDFF_4.LD.n18 7b_counter_0.MDFF_4.LD.t13 7.3005
R13631 7b_counter_0.MDFF_4.LD.n7 7b_counter_0.MDFF_4.LD.t124 7.3005
R13632 7b_counter_0.MDFF_4.LD.n1 7b_counter_0.MDFF_4.LD.n66 4.2255
R13633 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n65 4.19721
R13634 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n51 4.19721
R13635 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n58 4.19721
R13636 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n16 4.19721
R13637 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n23 4.19721
R13638 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n9 4.19721
R13639 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n30 4.19616
R13640 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n37 4.19616
R13641 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n44 4.19616
R13642 7b_counter_0.MDFF_4.LD.n2 7b_counter_0.MDFF_4.LD 3.73837
R13643 7b_counter_0.MDFF_4.LD.n2 7b_counter_0.MDFF_4.LD 3.73837
R13644 7b_counter_0.MDFF_4.LD.n79 7b_counter_0.MDFF_4.LD.n78 2.92988
R13645 7b_counter_0.MDFF_4.LD.n71 7b_counter_0.MDFF_4.LD.n70 2.90652
R13646 7b_counter_0.MDFF_4.LD.n71 7b_counter_0.MDFF_4.LD.n67 2.89193
R13647 7b_counter_0.MDFF_4.LD.n79 7b_counter_0.MDFF_4.LD.n72 2.85715
R13648 7b_counter_0.MDFF_4.LD.n77 7b_counter_0.MDFF_4.LD.n76 2.6005
R13649 7b_counter_0.MDFF_4.LD.n44 7b_counter_0.MDFF_4.LD.n40 2.54246
R13650 7b_counter_0.MDFF_4.LD.n16 7b_counter_0.MDFF_4.LD.n12 2.54246
R13651 7b_counter_0.MDFF_4.LD.n23 7b_counter_0.MDFF_4.LD.n19 2.54246
R13652 7b_counter_0.MDFF_4.LD.n30 7b_counter_0.MDFF_4.LD.n29 2.47729
R13653 7b_counter_0.MDFF_4.LD.n37 7b_counter_0.MDFF_4.LD.n36 2.47729
R13654 7b_counter_0.MDFF_4.LD.n51 7b_counter_0.MDFF_4.LD.n50 2.47729
R13655 7b_counter_0.MDFF_4.LD.n58 7b_counter_0.MDFF_4.LD.n57 2.47729
R13656 7b_counter_0.MDFF_4.LD.n9 7b_counter_0.MDFF_4.LD.n8 2.47729
R13657 7b_counter_0.MDFF_4.LD.n76 7b_counter_0.MDFF_4.LD.t4 1.6255
R13658 7b_counter_0.MDFF_4.LD.n76 7b_counter_0.MDFF_4.LD.n75 1.6255
R13659 7b_counter_0.MDFF_4.LD.n74 7b_counter_0.MDFF_4.LD.t8 1.6255
R13660 7b_counter_0.MDFF_4.LD.n74 7b_counter_0.MDFF_4.LD.n73 1.6255
R13661 7b_counter_0.MDFF_4.LD.n69 7b_counter_0.MDFF_4.LD.t3 1.463
R13662 7b_counter_0.MDFF_4.LD.n69 7b_counter_0.MDFF_4.LD.n68 1.463
R13663 7b_counter_0.MDFF_4.LD.n70 7b_counter_0.MDFF_4.LD.n69 1.43
R13664 7b_counter_0.MDFF_4.LD.n0 7b_counter_0.MDFF_4.LD 1.23561
R13665 7b_counter_0.MDFF_4.LD.n78 7b_counter_0.MDFF_4.LD.n74 1.23154
R13666 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n0 1.17946
R13667 7b_counter_0.MDFF_4.LD.n65 7b_counter_0.MDFF_4.LD.n61 1.04336
R13668 7b_counter_0.MDFF_4.LD.n78 7b_counter_0.MDFF_4.LD.n77 0.922667
R13669 7b_counter_0.MDFF_4.LD.n1 7b_counter_0.MDFF_4.LD.n79 0.829813
R13670 7b_counter_0.MDFF_4.LD.n1 7b_counter_0.MDFF_4.LD.n71 0.789247
R13671 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n2 0.601715
R13672 7b_counter_0.MDFF_4.LD.n2 7b_counter_0.MDFF_4.LD 0.465333
R13673 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n2 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t3 130.41
R13674 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n0 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t8 35.3186
R13675 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n3 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t5 33.5023
R13676 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t12 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n3 33.5023
R13677 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n1 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t4 32.2349
R13678 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n0 31.632
R13679 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n5 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t11 19.0118
R13680 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n4 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t12 16.3786
R13681 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t11 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n2 13.2317
R13682 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n2 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n1 13.0005
R13683 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n4 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t7 11.3259
R13684 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n1 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t6 11.146
R13685 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n0 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t9 7.3005
R13686 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n3 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t10 7.3005
R13687 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n8 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n6 5.47387
R13688 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n10 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n9 4.65398
R13689 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n8 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n7 4.2255
R13690 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n5 3.63228
R13691 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n5 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n4 3.62977
R13692 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n10 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n8 0.427022
R13693 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n10 0.257096
R13694 p3_gen_magic_0.3_inp_AND_magic_0.C.t6 p3_gen_magic_0.3_inp_AND_magic_0.C.t3 28.8746
R13695 p3_gen_magic_0.3_inp_AND_magic_0.C.n1 p3_gen_magic_0.3_inp_AND_magic_0.C.t4 25.7894
R13696 p3_gen_magic_0.3_inp_AND_magic_0.C.t4 p3_gen_magic_0.3_inp_AND_magic_0.C.t5 23.4648
R13697 p3_gen_magic_0.3_inp_AND_magic_0.C.n0 p3_gen_magic_0.3_inp_AND_magic_0.C.t7 17.1425
R13698 p3_gen_magic_0.3_inp_AND_magic_0.C.n0 p3_gen_magic_0.3_inp_AND_magic_0.C.t6 14.405
R13699 p3_gen_magic_0.3_inp_AND_magic_0.C.n1 p3_gen_magic_0.3_inp_AND_magic_0.C.n0 3.62425
R13700 p3_gen_magic_0.3_inp_AND_magic_0.C p3_gen_magic_0.3_inp_AND_magic_0.C.t1 3.46108
R13701 p3_gen_magic_0.3_inp_AND_magic_0.C p3_gen_magic_0.3_inp_AND_magic_0.C.n1 3.11402
R13702 p3_gen_magic_0.3_inp_AND_magic_0.C.t1 p3_gen_magic_0.3_inp_AND_magic_0.C.n2 1.6255
R13703 D2_5.t5 D2_5.t23 47.8944
R13704 D2_5.t10 D2_5.t6 47.8944
R13705 D2_5.t16 D2_5.t13 47.5387
R13706 D2_5.t2 D2_5.t20 47.5387
R13707 D2_5.t4 D2_5.t25 44.058
R13708 D2_5.t3 D2_5.t24 44.058
R13709 D2_5.n24 D2_5.t14 38.8649
R13710 D2_5.n0 D2_5.t15 38.8649
R13711 D2_5.n4 D2_5.t22 38.7949
R13712 D2_5.n3 D2_5.t1 38.7949
R13713 D2_5.n15 D2_5.t7 38.7949
R13714 D2_5.n14 D2_5.t9 38.7949
R13715 D2_5.n4 D2_5.n3 31.4949
R13716 D2_5.n15 D2_5.n14 31.4949
R13717 D2_5.t14 D2_5.t4 28.6791
R13718 D2_5.t15 D2_5.t3 28.6791
R13719 D2_5.n5 D2_5.t12 17.9416
R13720 D2_5.n16 D2_5.t19 17.9416
R13721 D2_5.n6 D2_5.t16 16.621
R13722 D2_5.n17 D2_5.t2 16.621
R13723 D2_5.n23 D2_5.n11 14.0832
R13724 D2_5.n25 D2_5.n23 13.4988
R13725 D2_5.n6 D2_5.t11 12.5148
R13726 D2_5.n17 D2_5.t18 12.5148
R13727 D2_5.n5 D2_5.t5 11.957
R13728 D2_5.n16 D2_5.t10 11.957
R13729 D2_5.n23 D2_5.n22 9.97869
R13730 D2_5.n3 D2_5.t8 7.3005
R13731 D2_5.t12 D2_5.n4 7.3005
R13732 D2_5.n14 D2_5.t17 7.3005
R13733 D2_5.t19 D2_5.n15 7.3005
R13734 D2_5.n24 D2_5.t21 7.3005
R13735 D2_5.n0 D2_5.t0 7.3005
R13736 D2_5 D2_5.n5 5.95286
R13737 D2_5 D2_5.n16 5.95286
R13738 D2_5.n26 D2_5.n25 5.86456
R13739 D2_5.n25 D2_5 5.66695
R13740 D2_5 D2_5.n24 5.27587
R13741 D2_5 D2_5.n0 5.27587
R13742 D2_5 D2_5.n6 4.59246
R13743 D2_5 D2_5.n17 4.59246
R13744 D2_5.n2 D2_5.n1 4.5005
R13745 D2_5.n19 D2_5.n13 3.38419
R13746 D2_5.n8 D2_5.n2 3.23516
R13747 D2_5.n9 D2_5.n8 2.60829
R13748 D2_5.n20 D2_5.n12 2.25826
R13749 D2_5.n22 D2_5.n21 2.25258
R13750 D2_5.n20 D2_5.n19 2.2505
R13751 D2_5.n21 D2_5.n13 2.24482
R13752 D2_5.n11 D2_5.n1 2.2437
R13753 D2_5.n10 D2_5.n9 1.5081
R13754 D2_5.n7 D2_5 1.4268
R13755 D2_5.n18 D2_5 1.35441
R13756 D2_5.n19 D2_5.n18 0.255095
R13757 D2_5.n18 D2_5 0.190361
R13758 D2_5.n8 D2_5.n7 0.137704
R13759 D2_5.n7 D2_5 0.11797
R13760 D2_5.n26 D2_5 0.0740494
R13761 D2_5 D2_5.n26 0.0339615
R13762 D2_5.n10 D2_5.n2 0.0297771
R13763 D2_5.n11 D2_5.n10 0.0166754
R13764 D2_5.n13 D2_5.n12 0.0142823
R13765 D2_5.n22 D2_5.n12 0.0134067
R13766 D2_5.n9 D2_5.n1 0.00176987
R13767 D2_5.n21 D2_5.n20 0.00165385
R13768 divide_by_2_1.tg_magic_3.CLK.t5 divide_by_2_1.tg_magic_3.CLK.t14 47.8944
R13769 divide_by_2_1.tg_magic_3.CLK.t4 divide_by_2_1.tg_magic_3.CLK.t3 47.8944
R13770 divide_by_2_1.tg_magic_3.CLK.n4 divide_by_2_1.tg_magic_3.CLK.t20 38.7949
R13771 divide_by_2_1.tg_magic_3.CLK.n5 divide_by_2_1.tg_magic_3.CLK.t18 38.7949
R13772 divide_by_2_1.tg_magic_3.CLK.n2 divide_by_2_1.tg_magic_3.CLK.t16 38.7949
R13773 divide_by_2_1.tg_magic_3.CLK.n1 divide_by_2_1.tg_magic_3.CLK.t11 38.7949
R13774 divide_by_2_1.tg_magic_3.CLK divide_by_2_1.tg_magic_3.CLK.t9 36.2535
R13775 divide_by_2_1.tg_magic_3.CLK divide_by_2_1.tg_magic_3.CLK.t7 36.1638
R13776 divide_by_2_1.tg_magic_3.CLK.n5 divide_by_2_1.tg_magic_3.CLK.n4 31.4949
R13777 divide_by_2_1.tg_magic_3.CLK.n2 divide_by_2_1.tg_magic_3.CLK.n1 31.4949
R13778 divide_by_2_1.tg_magic_3.CLK.n7 divide_by_2_1.tg_magic_3.CLK.t12 26.9781
R13779 divide_by_2_1.tg_magic_3.CLK.n7 divide_by_2_1.tg_magic_3.CLK.t19 26.9781
R13780 divide_by_2_1.tg_magic_3.CLK.n0 divide_by_2_1.tg_magic_3.CLK.t10 26.9781
R13781 divide_by_2_1.tg_magic_3.CLK.n0 divide_by_2_1.tg_magic_3.CLK.t8 26.9781
R13782 divide_by_2_1.tg_magic_3.CLK.n6 divide_by_2_1.tg_magic_3.CLK.t13 17.9416
R13783 divide_by_2_1.tg_magic_3.CLK.n3 divide_by_2_1.tg_magic_3.CLK.t17 17.9416
R13784 divide_by_2_1.tg_magic_3.CLK.n6 divide_by_2_1.tg_magic_3.CLK.t5 11.957
R13785 divide_by_2_1.tg_magic_3.CLK.n3 divide_by_2_1.tg_magic_3.CLK.t4 11.957
R13786 divide_by_2_1.tg_magic_3.CLK.n4 divide_by_2_1.tg_magic_3.CLK.t6 7.3005
R13787 divide_by_2_1.tg_magic_3.CLK.t13 divide_by_2_1.tg_magic_3.CLK.n5 7.3005
R13788 divide_by_2_1.tg_magic_3.CLK.t7 divide_by_2_1.tg_magic_3.CLK.n7 7.3005
R13789 divide_by_2_1.tg_magic_3.CLK.n1 divide_by_2_1.tg_magic_3.CLK.t15 7.3005
R13790 divide_by_2_1.tg_magic_3.CLK.t17 divide_by_2_1.tg_magic_3.CLK.n2 7.3005
R13791 divide_by_2_1.tg_magic_3.CLK.t9 divide_by_2_1.tg_magic_3.CLK.n0 7.3005
R13792 divide_by_2_1.tg_magic_3.CLK divide_by_2_1.tg_magic_3.CLK.n6 5.99387
R13793 divide_by_2_1.tg_magic_3.CLK divide_by_2_1.tg_magic_3.CLK.n3 5.77618
R13794 Q6.t15 Q6.t4 48.3065
R13795 Q6.n5 Q6 48.0285
R13796 Q6.t5 Q6.t29 47.8944
R13797 Q6.t24 Q6.t19 47.8944
R13798 Q6.t7 Q6.t21 47.5387
R13799 Q6.t27 Q6.t13 47.5387
R13800 Q6.t22 Q6.t20 44.058
R13801 Q6.n3 Q6.t12 38.8649
R13802 Q6.n18 Q6.t6 38.7949
R13803 Q6.n17 Q6.t10 38.7949
R13804 Q6.n9 Q6.t23 38.7949
R13805 Q6.n8 Q6.t26 38.7949
R13806 Q6.t4 Q6.t25 31.5469
R13807 Q6.t11 Q6.t15 31.5469
R13808 Q6.n18 Q6.n17 31.4949
R13809 Q6.n9 Q6.n8 31.4949
R13810 Q6.t12 Q6.t22 28.6791
R13811 Q6 Q6.n2 20.7556
R13812 Q6.n2 Q6.t11 18.2505
R13813 Q6.n19 Q6.t16 17.9416
R13814 Q6.n10 Q6.t9 17.9416
R13815 Q6.n5 Q6.n4 16.591
R13816 Q6.n20 Q6.t7 15.7085
R13817 Q6.n6 Q6.t27 15.7085
R13818 Q6 Q6.n22 14.6026
R13819 Q6.n22 Q6.n16 13.7743
R13820 Q6.n20 Q6.t28 13.4273
R13821 Q6.n6 Q6.t17 13.4273
R13822 Q6.n19 Q6.t5 11.957
R13823 Q6.n10 Q6.t24 11.957
R13824 Q6.n2 Q6.t8 11.4067
R13825 Q6.n3 Q6.t18 7.3005
R13826 Q6.n17 Q6.t14 7.3005
R13827 Q6.t16 Q6.n18 7.3005
R13828 Q6.n8 Q6.t3 7.3005
R13829 Q6.t9 Q6.n9 7.3005
R13830 Q6 Q6.n19 5.94647
R13831 Q6 Q6.n10 5.94647
R13832 Q6.n0 Q6.t0 5.47387
R13833 Q6 Q6.n3 5.27587
R13834 Q6.n1 Q6.t2 4.65398
R13835 Q6.n0 Q6.t1 4.2255
R13836 Q6 Q6.n20 4.08021
R13837 Q6 Q6.n6 4.08021
R13838 Q6.n12 Q6.n11 3.21398
R13839 Q6.n7 Q6 2.31011
R13840 Q6.n21 Q6 1.96503
R13841 Q6.n22 Q6.n21 1.95297
R13842 Q6 Q6.n5 1.88133
R13843 Q6.n15 Q6.n14 1.5081
R13844 Q6.n21 Q6 1.15959
R13845 Q6.n11 Q6 0.540318
R13846 Q6.n1 Q6.n0 0.427022
R13847 Q6 Q6.n1 0.257096
R13848 Q6.n11 Q6.n7 0.222553
R13849 Q6.n15 Q6.n12 0.0312595
R13850 Q6.n16 Q6.n15 0.0174666
R13851 Q6.n4 Q6 0.010625
R13852 Q6.n4 Q6 0.0095
R13853 Q6.n14 Q6.n13 0.00176987
R13854 divide_by_2_0.tg_magic_3.CLK.t13 divide_by_2_0.tg_magic_3.CLK.t19 47.8944
R13855 divide_by_2_0.tg_magic_3.CLK.t9 divide_by_2_0.tg_magic_3.CLK.t22 47.8944
R13856 divide_by_2_0.tg_magic_3.CLK.n5 divide_by_2_0.tg_magic_3.CLK.t17 38.7949
R13857 divide_by_2_0.tg_magic_3.CLK.n6 divide_by_2_0.tg_magic_3.CLK.t5 38.7949
R13858 divide_by_2_0.tg_magic_3.CLK.n3 divide_by_2_0.tg_magic_3.CLK.t6 38.7949
R13859 divide_by_2_0.tg_magic_3.CLK.n2 divide_by_2_0.tg_magic_3.CLK.t18 38.7949
R13860 divide_by_2_0.tg_magic_3.CLK divide_by_2_0.tg_magic_3.CLK.t12 36.2535
R13861 divide_by_2_0.tg_magic_3.CLK divide_by_2_0.tg_magic_3.CLK.t7 36.1638
R13862 divide_by_2_0.tg_magic_3.CLK.n6 divide_by_2_0.tg_magic_3.CLK.n5 31.4949
R13863 divide_by_2_0.tg_magic_3.CLK.n3 divide_by_2_0.tg_magic_3.CLK.n2 31.4949
R13864 divide_by_2_0.tg_magic_3.CLK.n8 divide_by_2_0.tg_magic_3.CLK.t10 26.9781
R13865 divide_by_2_0.tg_magic_3.CLK.n8 divide_by_2_0.tg_magic_3.CLK.t21 26.9781
R13866 divide_by_2_0.tg_magic_3.CLK.n1 divide_by_2_0.tg_magic_3.CLK.t15 26.9781
R13867 divide_by_2_0.tg_magic_3.CLK.n1 divide_by_2_0.tg_magic_3.CLK.t20 26.9781
R13868 divide_by_2_0.tg_magic_3.CLK.n7 divide_by_2_0.tg_magic_3.CLK.t8 17.9416
R13869 divide_by_2_0.tg_magic_3.CLK.n4 divide_by_2_0.tg_magic_3.CLK.t14 17.9416
R13870 divide_by_2_0.tg_magic_3.CLK.t2 divide_by_2_0.tg_magic_3.CLK 16.117
R13871 divide_by_2_0.tg_magic_3.CLK.n7 divide_by_2_0.tg_magic_3.CLK.t13 11.957
R13872 divide_by_2_0.tg_magic_3.CLK.n4 divide_by_2_0.tg_magic_3.CLK.t9 11.957
R13873 divide_by_2_0.tg_magic_3.CLK.n5 divide_by_2_0.tg_magic_3.CLK.t16 7.3005
R13874 divide_by_2_0.tg_magic_3.CLK.t8 divide_by_2_0.tg_magic_3.CLK.n6 7.3005
R13875 divide_by_2_0.tg_magic_3.CLK.t7 divide_by_2_0.tg_magic_3.CLK.n8 7.3005
R13876 divide_by_2_0.tg_magic_3.CLK.n2 divide_by_2_0.tg_magic_3.CLK.t11 7.3005
R13877 divide_by_2_0.tg_magic_3.CLK.t14 divide_by_2_0.tg_magic_3.CLK.n3 7.3005
R13878 divide_by_2_0.tg_magic_3.CLK.t12 divide_by_2_0.tg_magic_3.CLK.n1 7.3005
R13879 divide_by_2_0.tg_magic_3.CLK divide_by_2_0.tg_magic_3.CLK.n7 5.99387
R13880 divide_by_2_0.tg_magic_3.CLK divide_by_2_0.tg_magic_3.CLK.n4 5.77618
R13881 divide_by_2_0.tg_magic_3.CLK.t2 divide_by_2_0.tg_magic_3.CLK.t3 2.90572
R13882 divide_by_2_0.tg_magic_3.CLK.t3 divide_by_2_0.tg_magic_3.CLK.n0 1.6255
R13883 divide_by_2_0.tg_magic_3.CLK.t2 divide_by_2_0.tg_magic_3.CLK 1.31541
R13884 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t17 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t6 47.8944
R13885 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t23 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t19 47.8944
R13886 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n13 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t9 38.7949
R13887 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n14 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t22 38.7949
R13888 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n10 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t21 38.7949
R13889 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n9 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t14 38.7949
R13890 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n12 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t7 36.2535
R13891 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n17 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t12 36.1638
R13892 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n14 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n13 31.4949
R13893 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n10 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n9 31.4949
R13894 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n16 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t16 26.9781
R13895 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n16 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t10 26.9781
R13896 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n8 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t15 26.9781
R13897 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n8 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t8 26.9781
R13898 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n15 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t11 17.9416
R13899 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n11 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t20 17.9416
R13900 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n18 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK 16.117
R13901 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n15 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t17 11.957
R13902 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n11 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t23 11.957
R13903 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n13 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t18 7.3005
R13904 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t11 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n14 7.3005
R13905 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t12 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n16 7.3005
R13906 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n9 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t13 7.3005
R13907 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t20 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n10 7.3005
R13908 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t7 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n8 7.3005
R13909 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n12 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n11 5.77618
R13910 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n17 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n15 5.67753
R13911 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n4 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n1 3.6455
R13912 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n4 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n3 3.31072
R13913 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n7 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n6 2.90572
R13914 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n3 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t3 1.6255
R13915 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n3 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n2 1.6255
R13916 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n6 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t4 1.6255
R13917 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n6 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n5 1.6255
R13918 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n1 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t0 1.463
R13919 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n1 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n0 1.463
R13920 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n18 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK 0.717689
R13921 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n7 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n4 0.4055
R13922 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n17 0.187712
R13923 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n12 0.185948
R13924 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n7 0.179883
R13925 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n18 0.104263
R13926 Q7.t17 Q7.t19 48.5227
R13927 Q7.t7 Q7.t4 47.8944
R13928 Q7.t25 Q7.t21 47.8944
R13929 Q7.t6 Q7.t20 47.5387
R13930 Q7.t24 Q7.t12 47.5387
R13931 Q7.n5 Q7.t23 38.7949
R13932 Q7.n4 Q7.t22 38.7949
R13933 Q7.n15 Q7.t14 38.7949
R13934 Q7.n14 Q7.t13 38.7949
R13935 Q7.n29 Q7.n28 36.5454
R13936 Q7.n29 Q7.n1 34.6595
R13937 Q7.t19 Q7.t11 31.5469
R13938 Q7.n5 Q7.n4 31.4949
R13939 Q7.n15 Q7.n14 31.4949
R13940 Q7.t11 Q7.t10 29.6567
R13941 Q7.n6 Q7.t18 17.9416
R13942 Q7.n16 Q7.t8 17.9416
R13943 Q7.n0 Q7.t17 16.7514
R13944 Q7.n7 Q7.t6 15.7085
R13945 Q7.n13 Q7.t24 15.7085
R13946 Q7.n0 Q7.t9 14.796
R13947 Q7.n7 Q7.t3 13.4273
R13948 Q7.n13 Q7.t16 13.4273
R13949 Q7.n6 Q7.t7 11.957
R13950 Q7.n16 Q7.t25 11.957
R13951 Q7.n4 Q7.t15 7.3005
R13952 Q7.t18 Q7.n5 7.3005
R13953 Q7.n14 Q7.t5 7.3005
R13954 Q7.t8 Q7.n15 7.3005
R13955 Q7 Q7.n6 5.94647
R13956 Q7 Q7.n16 5.94647
R13957 Q7.n22 Q7.n21 5.85774
R13958 Q7.n33 Q7.n31 5.47387
R13959 Q7.n1 Q7.n0 4.97066
R13960 Q7.n35 Q7.n34 4.65398
R13961 Q7.n22 Q7.n9 4.5005
R13962 Q7.n3 Q7.n2 4.5005
R13963 Q7.n18 Q7.n17 4.47899
R13964 Q7.n33 Q7.n32 4.2255
R13965 Q7 Q7.n7 4.08021
R13966 Q7 Q7.n13 4.08021
R13967 Q7.n21 Q7.n20 3.15993
R13968 Q7.n8 Q7 3.0464
R13969 Q7.n17 Q7 2.86847
R13970 Q7.n30 Q7.n29 2.66587
R13971 Q7.n26 Q7.n25 2.51888
R13972 Q7.n21 Q7.n11 2.50168
R13973 Q7.n1 Q7 2.3623
R13974 Q7.n12 Q7.n11 2.25826
R13975 Q7.n19 Q7.n18 2.25218
R13976 Q7.n25 Q7.n24 2.25172
R13977 Q7.n20 Q7.n19 2.24442
R13978 Q7.n10 Q7.n9 2.24334
R13979 Q7.n28 Q7.n2 2.24334
R13980 Q7.n27 Q7.n26 1.5081
R13981 Q7.n24 Q7.n23 1.50776
R13982 Q7.n35 Q7.n33 0.427022
R13983 Q7 Q7.n35 0.257096
R13984 Q7.n10 Q7.n3 0.24236
R13985 Q7.n17 Q7 0.169666
R13986 Q7.n25 Q7.n8 0.133791
R13987 Q7.n8 Q7 0.0782273
R13988 Q7.n23 Q7.n22 0.0312595
R13989 Q7.n27 Q7.n3 0.0312595
R13990 Q7.n30 Q7 0.030875
R13991 Q7 Q7.n30 0.023
R13992 Q7.n23 Q7.n10 0.0174666
R13993 Q7.n28 Q7.n27 0.0174666
R13994 Q7.n20 Q7.n12 0.0151461
R13995 Q7.n18 Q7.n12 0.0142134
R13996 Q7.n24 Q7.n9 0.00243627
R13997 Q7.n26 Q7.n2 0.00176987
R13998 Q7.n19 Q7.n11 0.00165385
R13999 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n3 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t5 130.41
R14000 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n7 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t12 35.3186
R14001 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n4 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t6 33.5023
R14002 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t8 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n4 33.5023
R14003 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n2 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t10 32.2349
R14004 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n7 31.543
R14005 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n6 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t9 19.0138
R14006 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n5 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t8 16.3421
R14007 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t9 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n3 13.2317
R14008 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n3 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n2 13.0005
R14009 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n5 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t4 11.3624
R14010 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n2 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t3 11.146
R14011 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n4 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t7 7.3005
R14012 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n7 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t11 7.3005
R14013 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n0 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t0 5.47387
R14014 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n1 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t2 4.65398
R14015 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n0 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t1 4.2255
R14016 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n6 3.63214
R14017 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n6 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n5 3.62977
R14018 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n1 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n0 0.427022
R14019 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n1 0.257096
R14020 7b_counter_0.MDFF_4.QB.n5 7b_counter_0.MDFF_4.QB.t9 53.2571
R14021 7b_counter_0.MDFF_4.QB.t4 7b_counter_0.MDFF_4.QB.t6 44.058
R14022 7b_counter_0.MDFF_4.QB.n7 7b_counter_0.MDFF_4.QB.t8 38.8649
R14023 7b_counter_0.MDFF_4.QB.t8 7b_counter_0.MDFF_4.QB.t4 28.6791
R14024 7b_counter_0.MDFF_4.QB 7b_counter_0.MDFF_4.QB.n6 19.3781
R14025 7b_counter_0.MDFF_4.QB.n6 7b_counter_0.MDFF_4.QB.t10 17.1425
R14026 7b_counter_0.MDFF_4.QB.n6 7b_counter_0.MDFF_4.QB.t7 14.405
R14027 7b_counter_0.MDFF_4.QB.n7 7b_counter_0.MDFF_4.QB.t5 7.3005
R14028 7b_counter_0.MDFF_4.QB.t7 7b_counter_0.MDFF_4.QB.n5 7.3005
R14029 7b_counter_0.MDFF_4.QB 7b_counter_0.MDFF_4.QB.n7 5.4273
R14030 7b_counter_0.MDFF_4.QB.n5 7b_counter_0.MDFF_4.QB.n4 4.57931
R14031 7b_counter_0.MDFF_4.QB.n4 7b_counter_0.MDFF_4.QB.n1 3.62007
R14032 7b_counter_0.MDFF_4.QB.n4 7b_counter_0.MDFF_4.QB.n3 3.15478
R14033 7b_counter_0.MDFF_4.QB.n3 7b_counter_0.MDFF_4.QB.t1 1.6255
R14034 7b_counter_0.MDFF_4.QB.n3 7b_counter_0.MDFF_4.QB.n2 1.6255
R14035 7b_counter_0.MDFF_4.QB.n1 7b_counter_0.MDFF_4.QB.t3 1.463
R14036 7b_counter_0.MDFF_4.QB.n1 7b_counter_0.MDFF_4.QB.n0 1.463
R14037 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t20 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t22 47.8944
R14038 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t17 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t15 47.8944
R14039 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n13 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t12 38.7949
R14040 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n14 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t19 38.7949
R14041 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n10 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t10 38.7949
R14042 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n9 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t23 38.7949
R14043 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n12 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t21 36.2535
R14044 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n17 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t14 36.1638
R14045 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n14 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n13 31.4949
R14046 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n10 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n9 31.4949
R14047 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n16 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t16 26.9781
R14048 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n16 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t13 26.9781
R14049 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n8 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t7 26.9781
R14050 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n8 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t18 26.9781
R14051 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n15 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t6 17.9416
R14052 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n11 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t11 17.9416
R14053 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n18 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 16.117
R14054 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n15 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t20 11.957
R14055 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n11 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t17 11.957
R14056 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n13 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t8 7.3005
R14057 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t6 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n14 7.3005
R14058 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t14 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n16 7.3005
R14059 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n9 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t9 7.3005
R14060 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t11 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n10 7.3005
R14061 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t21 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n8 7.3005
R14062 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n12 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n11 5.77618
R14063 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n17 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n15 5.67753
R14064 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n4 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n1 3.6455
R14065 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n4 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n3 3.31072
R14066 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n7 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n6 2.90572
R14067 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n3 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t2 1.6255
R14068 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n3 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n2 1.6255
R14069 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n6 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t5 1.6255
R14070 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n6 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n5 1.6255
R14071 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n1 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t1 1.463
R14072 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n1 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n0 1.463
R14073 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n18 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 0.717689
R14074 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n7 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n4 0.4055
R14075 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n17 0.187712
R14076 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n12 0.185948
R14077 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n7 0.179883
R14078 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n18 0.104263
R14079 Q4.t22 Q4.t21 48.3065
R14080 Q4.t20 Q4.t16 47.8944
R14081 Q4.t29 Q4.t25 47.8944
R14082 Q4.t12 Q4.t7 47.5387
R14083 Q4.t23 Q4.t18 47.5387
R14084 Q4.t27 Q4.t4 44.058
R14085 Q4.n23 Q4.n22 42.2373
R14086 Q4.n21 Q4.t3 38.8649
R14087 Q4.n8 Q4.t19 38.7949
R14088 Q4.n7 Q4.t10 38.7949
R14089 Q4.n16 Q4.t28 38.7949
R14090 Q4.n15 Q4.t24 38.7949
R14091 Q4.t21 Q4.t13 31.5469
R14092 Q4.t14 Q4.t22 31.5469
R14093 Q4.n8 Q4.n7 31.4949
R14094 Q4.n16 Q4.n15 31.4949
R14095 Q4.t3 Q4.t27 28.6791
R14096 Q4.n20 Q4.n14 19.7703
R14097 Q4.n0 Q4.t14 18.2505
R14098 Q4.n1 Q4.n0 18.0612
R14099 Q4.n9 Q4.t5 17.9416
R14100 Q4.n17 Q4.t15 17.9416
R14101 Q4.n23 Q4.n20 17.379
R14102 Q4.n6 Q4.t12 15.7085
R14103 Q4.n18 Q4.t23 15.7085
R14104 Q4.n20 Q4.n19 14.7053
R14105 Q4 Q4.n1 14.0114
R14106 Q4.n6 Q4.t6 13.4273
R14107 Q4.n18 Q4.t17 13.4273
R14108 Q4.n9 Q4.t20 11.957
R14109 Q4.n17 Q4.t29 11.957
R14110 Q4.n0 Q4.t11 11.4067
R14111 Q4.n21 Q4.t9 7.3005
R14112 Q4.n7 Q4.t26 7.3005
R14113 Q4.t5 Q4.n8 7.3005
R14114 Q4.n15 Q4.t8 7.3005
R14115 Q4.t15 Q4.n16 7.3005
R14116 Q4 Q4.n9 5.94647
R14117 Q4 Q4.n17 5.94647
R14118 Q4.n2 Q4.t0 5.47387
R14119 Q4 Q4.n21 5.27587
R14120 Q4.n3 Q4.t1 4.65398
R14121 Q4.n14 Q4.n13 4.5005
R14122 Q4.n2 Q4.t2 4.2255
R14123 Q4 Q4.n6 4.08021
R14124 Q4 Q4.n18 4.08021
R14125 Q4.n12 Q4.n11 3.28355
R14126 Q4.n19 Q4 3.06276
R14127 Q4.n24 Q4.n23 2.54473
R14128 Q4.n11 Q4 2.3422
R14129 Q4.n10 Q4.n5 2.25138
R14130 Q4.n13 Q4.n12 2.24334
R14131 Q4.n5 Q4.n4 1.5081
R14132 Q4.n10 Q4 0.466518
R14133 Q4.n3 Q4.n2 0.427022
R14134 Q4.n24 Q4 0.291564
R14135 Q4.n11 Q4.n10 0.279201
R14136 Q4 Q4.n3 0.257096
R14137 Q4.n22 Q4 0.167977
R14138 Q4.n1 Q4 0.103054
R14139 Q4.n24 Q4 0.0713511
R14140 Q4.n19 Q4 0.0618636
R14141 Q4.n14 Q4.n4 0.0312595
R14142 Q4.n12 Q4.n4 0.0174666
R14143 Q4.n22 Q4 0.0156948
R14144 Q4 Q4.n24 0.00915385
R14145 Q4.n13 Q4.n5 0.00176987
R14146 OR_magic_2.A.t11 OR_magic_2.A.t16 47.8944
R14147 OR_magic_2.A.t6 OR_magic_2.A.t19 44.6331
R14148 OR_magic_2.A.t18 OR_magic_2.A.t15 44.6331
R14149 OR_magic_2.A.n1 OR_magic_2.A.t14 38.7949
R14150 OR_magic_2.A.n2 OR_magic_2.A.t17 38.7949
R14151 OR_magic_2.A.t10 OR_magic_2.A.t20 31.5469
R14152 OR_magic_2.A.t13 OR_magic_2.A.t21 31.5469
R14153 OR_magic_2.A.n2 OR_magic_2.A.n1 31.4949
R14154 OR_magic_2.A.t20 OR_magic_2.A.t9 28.6791
R14155 OR_magic_2.A.t21 OR_magic_2.A.t12 28.6791
R14156 OR_magic_2.A.n4 OR_magic_2.A 22.1185
R14157 OR_magic_2.A.n5 OR_magic_2.A.t6 19.4237
R14158 OR_magic_2.A.n0 OR_magic_2.A.t18 19.4237
R14159 OR_magic_2.A.n3 OR_magic_2.A.t7 17.9416
R14160 OR_magic_2.A.n6 OR_magic_2.A 13.8488
R14161 OR_magic_2.A.n5 OR_magic_2.A.t10 12.1237
R14162 OR_magic_2.A.n0 OR_magic_2.A.t13 12.1237
R14163 OR_magic_2.A.n3 OR_magic_2.A.t11 11.957
R14164 OR_magic_2.A.n1 OR_magic_2.A.t8 7.3005
R14165 OR_magic_2.A.t7 OR_magic_2.A.n2 7.3005
R14166 OR_magic_2.A OR_magic_2.A.n3 5.86241
R14167 OR_magic_2.A OR_magic_2.A.n5 4.23754
R14168 OR_magic_2.A OR_magic_2.A.n0 4.22853
R14169 OR_magic_2.A.n11 OR_magic_2.A.n8 3.6455
R14170 OR_magic_2.A.n11 OR_magic_2.A.n10 3.31072
R14171 OR_magic_2.A.n14 OR_magic_2.A.n13 2.90572
R14172 OR_magic_2.A.n10 OR_magic_2.A.t4 1.6255
R14173 OR_magic_2.A.n10 OR_magic_2.A.n9 1.6255
R14174 OR_magic_2.A.n13 OR_magic_2.A.t2 1.6255
R14175 OR_magic_2.A.n13 OR_magic_2.A.n12 1.6255
R14176 OR_magic_2.A.n8 OR_magic_2.A.t1 1.463
R14177 OR_magic_2.A.n8 OR_magic_2.A.n7 1.463
R14178 OR_magic_2.A.n6 OR_magic_2.A 1.25072
R14179 OR_magic_2.A OR_magic_2.A.n4 1.08637
R14180 OR_magic_2.A OR_magic_2.A.n6 0.642239
R14181 OR_magic_2.A.n4 OR_magic_2.A 0.594783
R14182 OR_magic_2.A.n14 OR_magic_2.A.n11 0.4055
R14183 OR_magic_2.A OR_magic_2.A.n14 0.178625
R14184 p2_gen_magic_0.3_inp_AND_magic_0.C.t3 p2_gen_magic_0.3_inp_AND_magic_0.C.t5 28.8746
R14185 p2_gen_magic_0.3_inp_AND_magic_0.C.n1 p2_gen_magic_0.3_inp_AND_magic_0.C.t7 25.7894
R14186 p2_gen_magic_0.3_inp_AND_magic_0.C.t7 p2_gen_magic_0.3_inp_AND_magic_0.C.t6 23.4648
R14187 p2_gen_magic_0.3_inp_AND_magic_0.C.n0 p2_gen_magic_0.3_inp_AND_magic_0.C.t4 17.1425
R14188 p2_gen_magic_0.3_inp_AND_magic_0.C.n0 p2_gen_magic_0.3_inp_AND_magic_0.C.t3 14.405
R14189 p2_gen_magic_0.3_inp_AND_magic_0.C.n1 p2_gen_magic_0.3_inp_AND_magic_0.C.n0 3.62425
R14190 p2_gen_magic_0.3_inp_AND_magic_0.C p2_gen_magic_0.3_inp_AND_magic_0.C.t1 3.46108
R14191 p2_gen_magic_0.3_inp_AND_magic_0.C p2_gen_magic_0.3_inp_AND_magic_0.C.n1 3.11402
R14192 p2_gen_magic_0.3_inp_AND_magic_0.C.t1 p2_gen_magic_0.3_inp_AND_magic_0.C.n2 1.6255
R14193 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n7 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t6 11.8647
R14194 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n2 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t10 5.68507
R14195 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n11 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n10 5.47974
R14196 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n6 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t0 4.928
R14197 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n12 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n8 4.77528
R14198 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n13 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t7 4.52027
R14199 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n11 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n9 4.2255
R14200 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t7 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n7 4.2255
R14201 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n5 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n4 3.1505
R14202 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n2 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n1 2.6005
R14203 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n1 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t8 1.6255
R14204 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n1 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n0 1.6255
R14205 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n4 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t1 1.463
R14206 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n4 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n3 1.463
R14207 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n6 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n5 1.16072
R14208 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n5 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n2 0.898543
R14209 p3_gen_magic_0.3_inp_AND_magic_0.VOUT p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n14 0.5135
R14210 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n14 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n13 0.3875
R14211 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n12 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n11 0.305717
R14212 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n14 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n7 0.299848
R14213 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n13 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n12 0.244879
R14214 p3_gen_magic_0.3_inp_AND_magic_0.VOUT p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n6 0.23682
R14215 OR_magic_1.VOUT.t14 OR_magic_1.VOUT.t16 47.8944
R14216 OR_magic_1.VOUT.t25 OR_magic_1.VOUT.t18 47.8944
R14217 OR_magic_1.VOUT.t23 OR_magic_1.VOUT.t15 47.8944
R14218 OR_magic_1.VOUT.n4 OR_magic_1.VOUT.t4 38.7949
R14219 OR_magic_1.VOUT.n5 OR_magic_1.VOUT.t20 38.7949
R14220 OR_magic_1.VOUT.n10 OR_magic_1.VOUT.t21 38.7949
R14221 OR_magic_1.VOUT.n9 OR_magic_1.VOUT.t9 38.7949
R14222 OR_magic_1.VOUT.n1 OR_magic_1.VOUT.t11 38.7949
R14223 OR_magic_1.VOUT.n0 OR_magic_1.VOUT.t5 38.7949
R14224 OR_magic_1.VOUT.n12 OR_magic_1.VOUT.t24 36.2535
R14225 OR_magic_1.VOUT.n5 OR_magic_1.VOUT.n4 31.4949
R14226 OR_magic_1.VOUT.n10 OR_magic_1.VOUT.n9 31.4949
R14227 OR_magic_1.VOUT.n1 OR_magic_1.VOUT.n0 31.4949
R14228 OR_magic_1.VOUT.n7 OR_magic_1.VOUT.t10 26.9781
R14229 OR_magic_1.VOUT.n7 OR_magic_1.VOUT.t26 26.9781
R14230 OR_magic_1.VOUT.n8 OR_magic_1.VOUT.t6 26.9781
R14231 OR_magic_1.VOUT.n8 OR_magic_1.VOUT.t22 26.9781
R14232 OR_magic_1.VOUT.n3 OR_magic_1.VOUT.t12 20.2675
R14233 OR_magic_1.VOUT.n6 OR_magic_1.VOUT.t8 17.9416
R14234 OR_magic_1.VOUT.n11 OR_magic_1.VOUT.t19 17.9416
R14235 OR_magic_1.VOUT.n2 OR_magic_1.VOUT.t17 17.9416
R14236 OR_magic_1.VOUT.n6 OR_magic_1.VOUT.t14 11.957
R14237 OR_magic_1.VOUT.n11 OR_magic_1.VOUT.t25 11.957
R14238 OR_magic_1.VOUT.n2 OR_magic_1.VOUT.t23 11.957
R14239 OR_magic_1.VOUT.n13 OR_magic_1.VOUT 8.06233
R14240 OR_magic_1.VOUT.n14 OR_magic_1.VOUT.n13 7.58578
R14241 OR_magic_1.VOUT.n4 OR_magic_1.VOUT.t3 7.3005
R14242 OR_magic_1.VOUT.t8 OR_magic_1.VOUT.n5 7.3005
R14243 OR_magic_1.VOUT.t12 OR_magic_1.VOUT.n7 7.3005
R14244 OR_magic_1.VOUT.n9 OR_magic_1.VOUT.t13 7.3005
R14245 OR_magic_1.VOUT.t19 OR_magic_1.VOUT.n10 7.3005
R14246 OR_magic_1.VOUT.t24 OR_magic_1.VOUT.n8 7.3005
R14247 OR_magic_1.VOUT.n0 OR_magic_1.VOUT.t7 7.3005
R14248 OR_magic_1.VOUT.t17 OR_magic_1.VOUT.n1 7.3005
R14249 OR_magic_1.VOUT OR_magic_1.VOUT.n2 5.96162
R14250 OR_magic_1.VOUT.n12 OR_magic_1.VOUT.n11 5.77618
R14251 OR_magic_1.VOUT.n3 OR_magic_1.VOUT.n6 5.67753
R14252 OR_magic_1.VOUT.n16 OR_magic_1.VOUT.n15 4.2255
R14253 OR_magic_1.VOUT.n14 OR_magic_1.VOUT 3.20528
R14254 OR_magic_1.VOUT OR_magic_1.VOUT.n14 2.28497
R14255 OR_magic_1.VOUT.n13 OR_magic_1.VOUT 0.81937
R14256 OR_magic_1.VOUT.n17 OR_magic_1.VOUT.n16 0.427022
R14257 OR_magic_1.VOUT OR_magic_1.VOUT.n12 0.315078
R14258 OR_magic_1.VOUT OR_magic_1.VOUT.n17 0.257096
R14259 OR_magic_1.VOUT OR_magic_1.VOUT.n3 0.227402
R14260 divide_by_2_0.tg_magic_1.IN.t12 divide_by_2_0.tg_magic_1.IN.t16 47.8944
R14261 divide_by_2_0.tg_magic_1.IN.n7 divide_by_2_0.tg_magic_1.IN.t15 38.7949
R14262 divide_by_2_0.tg_magic_1.IN.n8 divide_by_2_0.tg_magic_1.IN.t14 38.7949
R14263 divide_by_2_0.tg_magic_1.IN.n8 divide_by_2_0.tg_magic_1.IN.n7 31.4949
R14264 divide_by_2_0.tg_magic_1.IN.n9 divide_by_2_0.tg_magic_1.IN.t17 17.9416
R14265 divide_by_2_0.tg_magic_1.IN.n9 divide_by_2_0.tg_magic_1.IN.t12 11.957
R14266 divide_by_2_0.tg_magic_1.IN.n7 divide_by_2_0.tg_magic_1.IN.t13 7.3005
R14267 divide_by_2_0.tg_magic_1.IN.t17 divide_by_2_0.tg_magic_1.IN.n8 7.3005
R14268 divide_by_2_0.tg_magic_1.IN.n10 divide_by_2_0.tg_magic_1.IN 5.93058
R14269 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_1.IN.n9 5.86474
R14270 divide_by_2_0.tg_magic_1.IN.n2 divide_by_2_0.tg_magic_1.IN.t11 5.68507
R14271 divide_by_2_0.tg_magic_1.IN.n6 divide_by_2_0.tg_magic_1.IN.t1 4.92604
R14272 divide_by_2_0.tg_magic_1.IN.n17 divide_by_2_0.tg_magic_1.IN.n14 3.6455
R14273 divide_by_2_0.tg_magic_1.IN.n17 divide_by_2_0.tg_magic_1.IN.n16 3.31072
R14274 divide_by_2_0.tg_magic_1.IN.n5 divide_by_2_0.tg_magic_1.IN.n4 3.1505
R14275 divide_by_2_0.tg_magic_1.IN.n18 divide_by_2_0.tg_magic_1.IN.n12 2.90572
R14276 divide_by_2_0.tg_magic_1.IN.n2 divide_by_2_0.tg_magic_1.IN.n1 2.6005
R14277 divide_by_2_0.tg_magic_1.IN.n10 divide_by_2_0.tg_magic_1.IN 1.88467
R14278 divide_by_2_0.tg_magic_1.IN.n1 divide_by_2_0.tg_magic_1.IN.t10 1.6255
R14279 divide_by_2_0.tg_magic_1.IN.n1 divide_by_2_0.tg_magic_1.IN.n0 1.6255
R14280 divide_by_2_0.tg_magic_1.IN.n12 divide_by_2_0.tg_magic_1.IN.t6 1.6255
R14281 divide_by_2_0.tg_magic_1.IN.n12 divide_by_2_0.tg_magic_1.IN.n11 1.6255
R14282 divide_by_2_0.tg_magic_1.IN.n16 divide_by_2_0.tg_magic_1.IN.t8 1.6255
R14283 divide_by_2_0.tg_magic_1.IN.n16 divide_by_2_0.tg_magic_1.IN.n15 1.6255
R14284 divide_by_2_0.tg_magic_1.IN.n4 divide_by_2_0.tg_magic_1.IN.t2 1.463
R14285 divide_by_2_0.tg_magic_1.IN.n4 divide_by_2_0.tg_magic_1.IN.n3 1.463
R14286 divide_by_2_0.tg_magic_1.IN.n14 divide_by_2_0.tg_magic_1.IN.t4 1.463
R14287 divide_by_2_0.tg_magic_1.IN.n14 divide_by_2_0.tg_magic_1.IN.n13 1.463
R14288 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_1.IN.n10 1.33598
R14289 divide_by_2_0.tg_magic_1.IN.n6 divide_by_2_0.tg_magic_1.IN.n5 1.15166
R14290 divide_by_2_0.tg_magic_1.IN.n5 divide_by_2_0.tg_magic_1.IN.n2 0.898543
R14291 divide_by_2_0.tg_magic_1.IN.n18 divide_by_2_0.tg_magic_1.IN.n17 0.4055
R14292 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_1.IN.n6 0.198522
R14293 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_1.IN.n18 0.178625
R14294 divide_by_2_0.tg_magic_3.IN.t20 divide_by_2_0.tg_magic_3.IN.t22 47.8944
R14295 divide_by_2_0.tg_magic_3.IN.n8 divide_by_2_0.tg_magic_3.IN.t18 38.7949
R14296 divide_by_2_0.tg_magic_3.IN.n7 divide_by_2_0.tg_magic_3.IN.t23 38.7949
R14297 divide_by_2_0.tg_magic_3.IN.n8 divide_by_2_0.tg_magic_3.IN.n7 31.4949
R14298 divide_by_2_0.tg_magic_3.IN.n9 divide_by_2_0.tg_magic_3.IN.t21 17.9416
R14299 divide_by_2_0.tg_magic_3.IN.n9 divide_by_2_0.tg_magic_3.IN.t20 11.957
R14300 divide_by_2_0.tg_magic_3.IN.n7 divide_by_2_0.tg_magic_3.IN.t19 7.3005
R14301 divide_by_2_0.tg_magic_3.IN.t21 divide_by_2_0.tg_magic_3.IN.n8 7.3005
R14302 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_3.IN.n9 5.96162
R14303 divide_by_2_0.tg_magic_3.IN.n2 divide_by_2_0.tg_magic_3.IN.t1 5.68507
R14304 divide_by_2_0.tg_magic_3.IN.n25 divide_by_2_0.tg_magic_3.IN.n24 4.96909
R14305 divide_by_2_0.tg_magic_3.IN.n16 divide_by_2_0.tg_magic_3.IN.t13 4.96909
R14306 divide_by_2_0.tg_magic_3.IN.n6 divide_by_2_0.tg_magic_3.IN.t10 4.928
R14307 divide_by_2_0.tg_magic_3.IN.n14 divide_by_2_0.tg_magic_3.IN.n11 3.97619
R14308 divide_by_2_0.tg_magic_3.IN.n21 divide_by_2_0.tg_magic_3.IN.n20 3.97568
R14309 divide_by_2_0.tg_magic_3.IN.n5 divide_by_2_0.tg_magic_3.IN.n4 3.1505
R14310 divide_by_2_0.tg_magic_3.IN.n15 divide_by_2_0.tg_magic_3.IN.t15 2.87015
R14311 divide_by_2_0.tg_magic_3.IN.n23 divide_by_2_0.tg_magic_3.IN.n22 2.86969
R14312 divide_by_2_0.tg_magic_3.IN.n23 divide_by_2_0.tg_magic_3.IN.n21 2.86627
R14313 divide_by_2_0.tg_magic_3.IN.n15 divide_by_2_0.tg_magic_3.IN.n14 2.86528
R14314 divide_by_2_0.tg_magic_3.IN.n2 divide_by_2_0.tg_magic_3.IN.n1 2.6005
R14315 divide_by_2_0.tg_magic_3.IN.n18 divide_by_2_0.tg_magic_3.IN.t6 1.6255
R14316 divide_by_2_0.tg_magic_3.IN.n18 divide_by_2_0.tg_magic_3.IN.n17 1.6255
R14317 divide_by_2_0.tg_magic_3.IN.n13 divide_by_2_0.tg_magic_3.IN.t17 1.6255
R14318 divide_by_2_0.tg_magic_3.IN.n13 divide_by_2_0.tg_magic_3.IN.n12 1.6255
R14319 divide_by_2_0.tg_magic_3.IN.n1 divide_by_2_0.tg_magic_3.IN.t0 1.6255
R14320 divide_by_2_0.tg_magic_3.IN.n1 divide_by_2_0.tg_magic_3.IN.n0 1.6255
R14321 divide_by_2_0.tg_magic_3.IN.n4 divide_by_2_0.tg_magic_3.IN.t9 1.463
R14322 divide_by_2_0.tg_magic_3.IN.n4 divide_by_2_0.tg_magic_3.IN.n3 1.463
R14323 divide_by_2_0.tg_magic_3.IN.n20 divide_by_2_0.tg_magic_3.IN.t3 1.463
R14324 divide_by_2_0.tg_magic_3.IN.n20 divide_by_2_0.tg_magic_3.IN.n19 1.463
R14325 divide_by_2_0.tg_magic_3.IN.n11 divide_by_2_0.tg_magic_3.IN.t12 1.463
R14326 divide_by_2_0.tg_magic_3.IN.n11 divide_by_2_0.tg_magic_3.IN.n10 1.463
R14327 divide_by_2_0.tg_magic_3.IN.n14 divide_by_2_0.tg_magic_3.IN.n13 1.24557
R14328 divide_by_2_0.tg_magic_3.IN.n21 divide_by_2_0.tg_magic_3.IN.n18 1.24556
R14329 divide_by_2_0.tg_magic_3.IN.n6 divide_by_2_0.tg_magic_3.IN.n5 1.16072
R14330 divide_by_2_0.tg_magic_3.IN.n5 divide_by_2_0.tg_magic_3.IN.n2 0.898543
R14331 divide_by_2_0.tg_magic_3.IN.n16 divide_by_2_0.tg_magic_3.IN.n15 0.380457
R14332 divide_by_2_0.tg_magic_3.IN.n25 divide_by_2_0.tg_magic_3.IN.n23 0.379952
R14333 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_3.IN.n25 0.274825
R14334 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_3.IN.n6 0.260717
R14335 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_3.IN.n16 0.199452
R14336 a_27567_8496.t17 a_27567_8496.n0 39.6673
R14337 a_27567_8496.n0 a_27567_8496.t15 39.6673
R14338 a_27567_8496.n1 a_27567_8496.t9 39.3349
R14339 a_27567_8496.t13 a_27567_8496.n1 39.3349
R14340 a_27567_8496.t15 a_27567_8496.t10 31.0255
R14341 a_27567_8496.t16 a_27567_8496.t12 31.0255
R14342 a_27567_8496.t14 a_27567_8496.t13 29.1353
R14343 a_27567_8496.n2 a_27567_8496.t17 13.6103
R14344 a_27567_8496.n2 a_27567_8496.t14 12.9295
R14345 a_27567_8496.n0 a_27567_8496.t16 7.3005
R14346 a_27567_8496.n1 a_27567_8496.t11 7.3005
R14347 a_27567_8496.n8 a_27567_8496.n2 4.42281
R14348 a_27567_8496.n18 a_27567_8496.n17 4.2255
R14349 a_27567_8496.n7 a_27567_8496.n6 2.92496
R14350 a_27567_8496.n16 a_27567_8496.n15 2.9101
R14351 a_27567_8496.n16 a_27567_8496.n9 2.88638
R14352 a_27567_8496.n7 a_27567_8496.n3 2.86141
R14353 a_27567_8496.n12 a_27567_8496.n11 2.6005
R14354 a_27567_8496.n11 a_27567_8496.t7 1.6255
R14355 a_27567_8496.n11 a_27567_8496.n10 1.6255
R14356 a_27567_8496.n5 a_27567_8496.t4 1.6255
R14357 a_27567_8496.n5 a_27567_8496.n4 1.6255
R14358 a_27567_8496.n14 a_27567_8496.t1 1.463
R14359 a_27567_8496.n14 a_27567_8496.n13 1.463
R14360 a_27567_8496.n15 a_27567_8496.n14 1.42734
R14361 a_27567_8496.n6 a_27567_8496.n5 1.23607
R14362 a_27567_8496.n17 a_27567_8496.n16 0.813345
R14363 a_27567_8496.n15 a_27567_8496.n12 0.800806
R14364 a_27567_8496.n8 a_27567_8496.n7 0.402859
R14365 a_27567_8496.n17 a_27567_8496.n8 0.395717
R14366 a_31440_8496.t9 a_31440_8496.n0 39.6673
R14367 a_31440_8496.n0 a_31440_8496.t16 39.6673
R14368 a_31440_8496.n1 a_31440_8496.t10 39.3349
R14369 a_31440_8496.t14 a_31440_8496.n1 39.3349
R14370 a_31440_8496.t16 a_31440_8496.t11 31.0255
R14371 a_31440_8496.t17 a_31440_8496.t13 31.0255
R14372 a_31440_8496.t15 a_31440_8496.t14 29.1353
R14373 a_31440_8496.n2 a_31440_8496.t9 13.6103
R14374 a_31440_8496.n2 a_31440_8496.t15 12.9295
R14375 a_31440_8496.n0 a_31440_8496.t17 7.3005
R14376 a_31440_8496.n1 a_31440_8496.t12 7.3005
R14377 a_31440_8496.n8 a_31440_8496.n2 4.42281
R14378 a_31440_8496.n18 a_31440_8496.n17 4.2255
R14379 a_31440_8496.n7 a_31440_8496.n6 2.92496
R14380 a_31440_8496.n16 a_31440_8496.n15 2.9101
R14381 a_31440_8496.n16 a_31440_8496.n9 2.88638
R14382 a_31440_8496.n7 a_31440_8496.n3 2.86141
R14383 a_31440_8496.n12 a_31440_8496.n11 2.6005
R14384 a_31440_8496.n11 a_31440_8496.t7 1.6255
R14385 a_31440_8496.n11 a_31440_8496.n10 1.6255
R14386 a_31440_8496.n5 a_31440_8496.t4 1.6255
R14387 a_31440_8496.n5 a_31440_8496.n4 1.6255
R14388 a_31440_8496.n14 a_31440_8496.t1 1.463
R14389 a_31440_8496.n14 a_31440_8496.n13 1.463
R14390 a_31440_8496.n15 a_31440_8496.n14 1.42734
R14391 a_31440_8496.n6 a_31440_8496.n5 1.23607
R14392 a_31440_8496.n17 a_31440_8496.n16 0.813345
R14393 a_31440_8496.n15 a_31440_8496.n12 0.800806
R14394 a_31440_8496.n8 a_31440_8496.n7 0.402859
R14395 a_31440_8496.n17 a_31440_8496.n8 0.395717
R14396 p3_gen_magic_0.xnor_magic_5.OUT.t6 p3_gen_magic_0.xnor_magic_5.OUT.t8 144.929
R14397 p3_gen_magic_0.xnor_magic_5.OUT.t5 p3_gen_magic_0.xnor_magic_5.OUT.t7 44.058
R14398 p3_gen_magic_0.xnor_magic_5.OUT.n4 p3_gen_magic_0.xnor_magic_5.OUT 22.3661
R14399 p3_gen_magic_0.xnor_magic_5.OUT.n3 p3_gen_magic_0.xnor_magic_5.OUT.t6 14.796
R14400 p3_gen_magic_0.xnor_magic_5.OUT.n3 p3_gen_magic_0.xnor_magic_5.OUT.t5 13.8835
R14401 p3_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_5.OUT.n3 9.82332
R14402 p3_gen_magic_0.xnor_magic_5.OUT.n4 p3_gen_magic_0.xnor_magic_5.OUT.n2 4.11572
R14403 p3_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_5.OUT.n4 3.61488
R14404 p3_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_5.OUT.t0 2.96833
R14405 p3_gen_magic_0.xnor_magic_5.OUT.t0 p3_gen_magic_0.xnor_magic_5.OUT.n0 1.6255
R14406 p3_gen_magic_0.xnor_magic_5.OUT.n2 p3_gen_magic_0.xnor_magic_5.OUT.t4 1.463
R14407 p3_gen_magic_0.xnor_magic_5.OUT.n2 p3_gen_magic_0.xnor_magic_5.OUT.n1 1.463
R14408 divide_by_2_1.tg_magic_3.IN.t23 divide_by_2_1.tg_magic_3.IN.t20 47.8944
R14409 divide_by_2_1.tg_magic_3.IN.n1 divide_by_2_1.tg_magic_3.IN.t22 38.7949
R14410 divide_by_2_1.tg_magic_3.IN.n0 divide_by_2_1.tg_magic_3.IN.t18 38.7949
R14411 divide_by_2_1.tg_magic_3.IN.n1 divide_by_2_1.tg_magic_3.IN.n0 31.4949
R14412 divide_by_2_1.tg_magic_3.IN.n2 divide_by_2_1.tg_magic_3.IN.t21 17.9416
R14413 divide_by_2_1.tg_magic_3.IN.n2 divide_by_2_1.tg_magic_3.IN.t23 11.957
R14414 divide_by_2_1.tg_magic_3.IN.n0 divide_by_2_1.tg_magic_3.IN.t19 7.3005
R14415 divide_by_2_1.tg_magic_3.IN.t21 divide_by_2_1.tg_magic_3.IN.n1 7.3005
R14416 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_3.IN.n2 5.96162
R14417 divide_by_2_1.tg_magic_3.IN.n5 divide_by_2_1.tg_magic_3.IN.t15 5.68507
R14418 divide_by_2_1.tg_magic_3.IN.n25 divide_by_2_1.tg_magic_3.IN.t13 4.96909
R14419 divide_by_2_1.tg_magic_3.IN.n18 divide_by_2_1.tg_magic_3.IN.n17 4.96909
R14420 divide_by_2_1.tg_magic_3.IN.n9 divide_by_2_1.tg_magic_3.IN.t9 4.928
R14421 divide_by_2_1.tg_magic_3.IN.n23 divide_by_2_1.tg_magic_3.IN.n20 3.97619
R14422 divide_by_2_1.tg_magic_3.IN.n14 divide_by_2_1.tg_magic_3.IN.n13 3.97568
R14423 divide_by_2_1.tg_magic_3.IN.n8 divide_by_2_1.tg_magic_3.IN.n7 3.1505
R14424 divide_by_2_1.tg_magic_3.IN.n24 divide_by_2_1.tg_magic_3.IN.t2 2.87015
R14425 divide_by_2_1.tg_magic_3.IN.n16 divide_by_2_1.tg_magic_3.IN.n15 2.86969
R14426 divide_by_2_1.tg_magic_3.IN.n16 divide_by_2_1.tg_magic_3.IN.n14 2.86627
R14427 divide_by_2_1.tg_magic_3.IN.n24 divide_by_2_1.tg_magic_3.IN.n23 2.86504
R14428 divide_by_2_1.tg_magic_3.IN.n5 divide_by_2_1.tg_magic_3.IN.n4 2.6005
R14429 divide_by_2_1.tg_magic_3.IN.n4 divide_by_2_1.tg_magic_3.IN.t17 1.6255
R14430 divide_by_2_1.tg_magic_3.IN.n4 divide_by_2_1.tg_magic_3.IN.n3 1.6255
R14431 divide_by_2_1.tg_magic_3.IN.n11 divide_by_2_1.tg_magic_3.IN.t3 1.6255
R14432 divide_by_2_1.tg_magic_3.IN.n11 divide_by_2_1.tg_magic_3.IN.n10 1.6255
R14433 divide_by_2_1.tg_magic_3.IN.n22 divide_by_2_1.tg_magic_3.IN.t0 1.6255
R14434 divide_by_2_1.tg_magic_3.IN.n22 divide_by_2_1.tg_magic_3.IN.n21 1.6255
R14435 divide_by_2_1.tg_magic_3.IN.n7 divide_by_2_1.tg_magic_3.IN.t11 1.463
R14436 divide_by_2_1.tg_magic_3.IN.n7 divide_by_2_1.tg_magic_3.IN.n6 1.463
R14437 divide_by_2_1.tg_magic_3.IN.n13 divide_by_2_1.tg_magic_3.IN.t6 1.463
R14438 divide_by_2_1.tg_magic_3.IN.n13 divide_by_2_1.tg_magic_3.IN.n12 1.463
R14439 divide_by_2_1.tg_magic_3.IN.n20 divide_by_2_1.tg_magic_3.IN.t12 1.463
R14440 divide_by_2_1.tg_magic_3.IN.n20 divide_by_2_1.tg_magic_3.IN.n19 1.463
R14441 divide_by_2_1.tg_magic_3.IN.n23 divide_by_2_1.tg_magic_3.IN.n22 1.24557
R14442 divide_by_2_1.tg_magic_3.IN.n14 divide_by_2_1.tg_magic_3.IN.n11 1.24556
R14443 divide_by_2_1.tg_magic_3.IN.n9 divide_by_2_1.tg_magic_3.IN.n8 1.16072
R14444 divide_by_2_1.tg_magic_3.IN.n8 divide_by_2_1.tg_magic_3.IN.n5 0.898543
R14445 divide_by_2_1.tg_magic_3.IN.n25 divide_by_2_1.tg_magic_3.IN.n24 0.380457
R14446 divide_by_2_1.tg_magic_3.IN.n18 divide_by_2_1.tg_magic_3.IN.n16 0.379952
R14447 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_3.IN.n18 0.274825
R14448 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_3.IN.n9 0.260717
R14449 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_3.IN.n25 0.199452
R14450 mux_magic_0.IN1.t8 mux_magic_0.IN1.t11 47.8944
R14451 mux_magic_0.IN1.t7 mux_magic_0.IN1.t6 44.058
R14452 mux_magic_0.IN1.n0 mux_magic_0.IN1.t12 38.8649
R14453 mux_magic_0.IN1.n1 mux_magic_0.IN1.t14 38.7949
R14454 mux_magic_0.IN1.n2 mux_magic_0.IN1.t13 38.7949
R14455 mux_magic_0.IN1.n2 mux_magic_0.IN1.n1 31.4949
R14456 mux_magic_0.IN1.t12 mux_magic_0.IN1.t7 28.6791
R14457 mux_magic_0.IN1.n3 mux_magic_0.IN1.t10 17.9416
R14458 mux_magic_0.IN1.n4 mux_magic_0.IN1 17.0637
R14459 mux_magic_0.IN1.n3 mux_magic_0.IN1.t8 11.957
R14460 mux_magic_0.IN1.n0 mux_magic_0.IN1.t15 7.3005
R14461 mux_magic_0.IN1.n1 mux_magic_0.IN1.t9 7.3005
R14462 mux_magic_0.IN1.t10 mux_magic_0.IN1.n2 7.3005
R14463 mux_magic_0.IN1 mux_magic_0.IN1.n3 5.86241
R14464 mux_magic_0.IN1 mux_magic_0.IN1.n0 5.27587
R14465 mux_magic_0.IN1.n9 mux_magic_0.IN1.n6 3.6455
R14466 mux_magic_0.IN1.n9 mux_magic_0.IN1.n8 3.31072
R14467 mux_magic_0.IN1.n12 mux_magic_0.IN1.n11 2.90572
R14468 mux_magic_0.IN1.n8 mux_magic_0.IN1.t3 1.6255
R14469 mux_magic_0.IN1.n8 mux_magic_0.IN1.n7 1.6255
R14470 mux_magic_0.IN1.n11 mux_magic_0.IN1.t5 1.6255
R14471 mux_magic_0.IN1.n11 mux_magic_0.IN1.n10 1.6255
R14472 mux_magic_0.IN1.n6 mux_magic_0.IN1.t1 1.463
R14473 mux_magic_0.IN1.n6 mux_magic_0.IN1.n5 1.463
R14474 mux_magic_0.IN1 mux_magic_0.IN1.n4 1.08637
R14475 mux_magic_0.IN1.n4 mux_magic_0.IN1 0.594783
R14476 mux_magic_0.IN1.n12 mux_magic_0.IN1.n9 0.4055
R14477 mux_magic_0.IN1 mux_magic_0.IN1.n12 0.178625
R14478 p3_gen_magic_0.xnor_magic_3.OUT.t6 p3_gen_magic_0.xnor_magic_3.OUT.t5 28.8746
R14479 p3_gen_magic_0.xnor_magic_3.OUT.n2 p3_gen_magic_0.xnor_magic_3.OUT.t7 25.7891
R14480 p3_gen_magic_0.xnor_magic_3.OUT.t7 p3_gen_magic_0.xnor_magic_3.OUT.t8 23.4648
R14481 p3_gen_magic_0.xnor_magic_3.OUT.n6 p3_gen_magic_0.xnor_magic_3.OUT.n3 17.1813
R14482 p3_gen_magic_0.xnor_magic_3.OUT.n1 p3_gen_magic_0.xnor_magic_3.OUT.t9 17.1425
R14483 p3_gen_magic_0.xnor_magic_3.OUT.n1 p3_gen_magic_0.xnor_magic_3.OUT.t6 14.405
R14484 p3_gen_magic_0.xnor_magic_3.OUT.n6 p3_gen_magic_0.xnor_magic_3.OUT.n5 4.11507
R14485 p3_gen_magic_0.xnor_magic_3.OUT.n2 p3_gen_magic_0.xnor_magic_3.OUT.n1 3.62425
R14486 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_3.OUT.n6 3.61488
R14487 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_3.OUT.t1 3.11311
R14488 p3_gen_magic_0.xnor_magic_3.OUT.n3 p3_gen_magic_0.xnor_magic_3.OUT 2.33511
R14489 p3_gen_magic_0.xnor_magic_3.OUT.t1 p3_gen_magic_0.xnor_magic_3.OUT.n0 1.6255
R14490 p3_gen_magic_0.xnor_magic_3.OUT.n5 p3_gen_magic_0.xnor_magic_3.OUT.t3 1.463
R14491 p3_gen_magic_0.xnor_magic_3.OUT.n5 p3_gen_magic_0.xnor_magic_3.OUT.n4 1.463
R14492 p3_gen_magic_0.xnor_magic_3.OUT.n3 p3_gen_magic_0.xnor_magic_3.OUT.n2 0.853219
R14493 divide_by_2_1.tg_magic_1.IN.t14 divide_by_2_1.tg_magic_1.IN.t16 47.8944
R14494 divide_by_2_1.tg_magic_1.IN.n7 divide_by_2_1.tg_magic_1.IN.t13 38.7949
R14495 divide_by_2_1.tg_magic_1.IN.n8 divide_by_2_1.tg_magic_1.IN.t17 38.7949
R14496 divide_by_2_1.tg_magic_1.IN.n8 divide_by_2_1.tg_magic_1.IN.n7 31.4949
R14497 divide_by_2_1.tg_magic_1.IN.n9 divide_by_2_1.tg_magic_1.IN.t15 17.9416
R14498 divide_by_2_1.tg_magic_1.IN.n9 divide_by_2_1.tg_magic_1.IN.t14 11.957
R14499 divide_by_2_1.tg_magic_1.IN.n7 divide_by_2_1.tg_magic_1.IN.t12 7.3005
R14500 divide_by_2_1.tg_magic_1.IN.t15 divide_by_2_1.tg_magic_1.IN.n8 7.3005
R14501 divide_by_2_1.tg_magic_1.IN.n10 divide_by_2_1.tg_magic_1.IN 5.93058
R14502 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_1.IN.n9 5.86474
R14503 divide_by_2_1.tg_magic_1.IN.n2 divide_by_2_1.tg_magic_1.IN.t6 5.68507
R14504 divide_by_2_1.tg_magic_1.IN.n6 divide_by_2_1.tg_magic_1.IN.t11 4.92604
R14505 divide_by_2_1.tg_magic_1.IN.n17 divide_by_2_1.tg_magic_1.IN.n14 3.6455
R14506 divide_by_2_1.tg_magic_1.IN.n17 divide_by_2_1.tg_magic_1.IN.n16 3.31072
R14507 divide_by_2_1.tg_magic_1.IN.n5 divide_by_2_1.tg_magic_1.IN.n4 3.1505
R14508 divide_by_2_1.tg_magic_1.IN.n18 divide_by_2_1.tg_magic_1.IN.n12 2.90572
R14509 divide_by_2_1.tg_magic_1.IN.n2 divide_by_2_1.tg_magic_1.IN.n1 2.6005
R14510 divide_by_2_1.tg_magic_1.IN.n10 divide_by_2_1.tg_magic_1.IN 1.88467
R14511 divide_by_2_1.tg_magic_1.IN.n1 divide_by_2_1.tg_magic_1.IN.t8 1.6255
R14512 divide_by_2_1.tg_magic_1.IN.n1 divide_by_2_1.tg_magic_1.IN.n0 1.6255
R14513 divide_by_2_1.tg_magic_1.IN.n12 divide_by_2_1.tg_magic_1.IN.t3 1.6255
R14514 divide_by_2_1.tg_magic_1.IN.n12 divide_by_2_1.tg_magic_1.IN.n11 1.6255
R14515 divide_by_2_1.tg_magic_1.IN.n16 divide_by_2_1.tg_magic_1.IN.t4 1.6255
R14516 divide_by_2_1.tg_magic_1.IN.n16 divide_by_2_1.tg_magic_1.IN.n15 1.6255
R14517 divide_by_2_1.tg_magic_1.IN.n4 divide_by_2_1.tg_magic_1.IN.t10 1.463
R14518 divide_by_2_1.tg_magic_1.IN.n4 divide_by_2_1.tg_magic_1.IN.n3 1.463
R14519 divide_by_2_1.tg_magic_1.IN.n14 divide_by_2_1.tg_magic_1.IN.t1 1.463
R14520 divide_by_2_1.tg_magic_1.IN.n14 divide_by_2_1.tg_magic_1.IN.n13 1.463
R14521 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_1.IN.n10 1.33598
R14522 divide_by_2_1.tg_magic_1.IN.n6 divide_by_2_1.tg_magic_1.IN.n5 1.15166
R14523 divide_by_2_1.tg_magic_1.IN.n5 divide_by_2_1.tg_magic_1.IN.n2 0.898543
R14524 divide_by_2_1.tg_magic_1.IN.n18 divide_by_2_1.tg_magic_1.IN.n17 0.4055
R14525 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_1.IN.n6 0.198522
R14526 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_1.IN.n18 0.178625
R14527 Q5.t4 Q5.t14 48.5227
R14528 Q5.t13 Q5.t9 47.8944
R14529 Q5.t23 Q5.t17 47.8944
R14530 Q5.t16 Q5.t10 47.5387
R14531 Q5.t24 Q5.t19 47.5387
R14532 Q5.t15 Q5.t7 44.058
R14533 Q5.n33 Q5.n16 39.7927
R14534 Q5.n0 Q5.t28 38.8649
R14535 Q5.n13 Q5.t11 38.7949
R14536 Q5.n12 Q5.t12 38.7949
R14537 Q5.n23 Q5.t21 38.7949
R14538 Q5.n22 Q5.t22 38.7949
R14539 Q5.n37 Q5 34.8562
R14540 Q5.t14 Q5.t5 31.5469
R14541 Q5.n13 Q5.n12 31.4949
R14542 Q5.n23 Q5.n22 31.4949
R14543 Q5.t5 Q5.t3 29.6567
R14544 Q5.t28 Q5.t15 28.6791
R14545 Q5.n7 Q5.n1 23.6541
R14546 Q5.n14 Q5.t25 17.9416
R14547 Q5.n24 Q5.t6 17.9416
R14548 Q5.n9 Q5.t4 16.7514
R14549 Q5.n15 Q5.t16 15.7085
R14550 Q5.n21 Q5.t24 15.7085
R14551 Q5.n9 Q5.t27 14.796
R14552 Q5.n15 Q5.t8 13.4273
R14553 Q5.n21 Q5.t18 13.4273
R14554 Q5.n14 Q5.t13 11.957
R14555 Q5.n24 Q5.t23 11.957
R14556 Q5 Q5.n9 7.34862
R14557 Q5.n0 Q5.t26 7.3005
R14558 Q5.n12 Q5.t20 7.3005
R14559 Q5.t25 Q5.n13 7.3005
R14560 Q5.n22 Q5.t29 7.3005
R14561 Q5.t6 Q5.n23 7.3005
R14562 Q5.n37 Q5.n36 6.32392
R14563 Q5 Q5.n14 5.94647
R14564 Q5 Q5.n24 5.94647
R14565 Q5.n30 Q5.n29 5.62253
R14566 Q5.n4 Q5.n2 5.47387
R14567 Q5 Q5.n0 5.27587
R14568 Q5.n6 Q5.n5 4.65398
R14569 Q5.n20 Q5.n19 4.5005
R14570 Q5.n30 Q5.n17 4.5005
R14571 Q5.n11 Q5.n10 4.5005
R14572 Q5.n4 Q5.n3 4.2255
R14573 Q5 Q5.n15 4.08021
R14574 Q5 Q5.n21 4.08021
R14575 Q5.n25 Q5.n20 3.4766
R14576 Q5.n34 Q5.n33 2.47039
R14577 Q5.n33 Q5.n32 2.46133
R14578 Q5.n27 Q5.n26 2.25138
R14579 Q5.n29 Q5.n19 2.24334
R14580 Q5.n18 Q5.n17 2.24334
R14581 Q5.n36 Q5.n10 2.24334
R14582 Q5.n16 Q5 1.96503
R14583 Q5.n26 Q5 1.90207
R14584 Q5.n28 Q5.n27 1.5081
R14585 Q5.n35 Q5.n34 1.5081
R14586 Q5.n32 Q5.n31 1.50776
R14587 Q5 Q5.n37 1.43232
R14588 Q5.n16 Q5 1.15959
R14589 Q5.n25 Q5 0.702722
R14590 Q5.n18 Q5.n11 0.49553
R14591 Q5.n26 Q5.n25 0.47224
R14592 Q5.n6 Q5.n4 0.427022
R14593 Q5 Q5.n6 0.257096
R14594 Q5 Q5.n8 0.113409
R14595 Q5.n28 Q5.n20 0.0312595
R14596 Q5.n31 Q5.n30 0.0312595
R14597 Q5.n35 Q5.n11 0.0312595
R14598 Q5.n7 Q5 0.02675
R14599 Q5.n8 Q5 0.02425
R14600 Q5.n1 Q5 0.0182778
R14601 Q5.n29 Q5.n28 0.0174666
R14602 Q5.n31 Q5.n18 0.0174666
R14603 Q5.n36 Q5.n35 0.0174666
R14604 Q5.n8 Q5.n7 0.00925
R14605 Q5.n32 Q5.n17 0.00243627
R14606 Q5.n34 Q5.n10 0.00176987
R14607 Q5.n27 Q5.n19 0.00176987
R14608 Q5.n1 Q5 0.00161111
R14609 DFF_magic_0.tg_magic_3.CLK.t18 DFF_magic_0.tg_magic_3.CLK.t16 47.8944
R14610 DFF_magic_0.tg_magic_3.CLK.t15 DFF_magic_0.tg_magic_3.CLK.t11 47.8944
R14611 DFF_magic_0.tg_magic_3.CLK.n13 DFF_magic_0.tg_magic_3.CLK.t20 38.7949
R14612 DFF_magic_0.tg_magic_3.CLK.n14 DFF_magic_0.tg_magic_3.CLK.t23 38.7949
R14613 DFF_magic_0.tg_magic_3.CLK.n10 DFF_magic_0.tg_magic_3.CLK.t22 38.7949
R14614 DFF_magic_0.tg_magic_3.CLK.n9 DFF_magic_0.tg_magic_3.CLK.t19 38.7949
R14615 DFF_magic_0.tg_magic_3.CLK.n12 DFF_magic_0.tg_magic_3.CLK.t14 36.2535
R14616 DFF_magic_0.tg_magic_3.CLK.n17 DFF_magic_0.tg_magic_3.CLK.t13 36.1638
R14617 DFF_magic_0.tg_magic_3.CLK.n14 DFF_magic_0.tg_magic_3.CLK.n13 31.4949
R14618 DFF_magic_0.tg_magic_3.CLK.n10 DFF_magic_0.tg_magic_3.CLK.n9 31.4949
R14619 DFF_magic_0.tg_magic_3.CLK.n16 DFF_magic_0.tg_magic_3.CLK.t17 26.9781
R14620 DFF_magic_0.tg_magic_3.CLK.n16 DFF_magic_0.tg_magic_3.CLK.t10 26.9781
R14621 DFF_magic_0.tg_magic_3.CLK.n8 DFF_magic_0.tg_magic_3.CLK.t6 26.9781
R14622 DFF_magic_0.tg_magic_3.CLK.n8 DFF_magic_0.tg_magic_3.CLK.t9 26.9781
R14623 DFF_magic_0.tg_magic_3.CLK.n15 DFF_magic_0.tg_magic_3.CLK.t12 17.9416
R14624 DFF_magic_0.tg_magic_3.CLK.n11 DFF_magic_0.tg_magic_3.CLK.t7 17.9416
R14625 DFF_magic_0.tg_magic_3.CLK.n18 DFF_magic_0.tg_magic_3.CLK 16.117
R14626 DFF_magic_0.tg_magic_3.CLK.n15 DFF_magic_0.tg_magic_3.CLK.t18 11.957
R14627 DFF_magic_0.tg_magic_3.CLK.n11 DFF_magic_0.tg_magic_3.CLK.t15 11.957
R14628 DFF_magic_0.tg_magic_3.CLK.n13 DFF_magic_0.tg_magic_3.CLK.t8 7.3005
R14629 DFF_magic_0.tg_magic_3.CLK.t12 DFF_magic_0.tg_magic_3.CLK.n14 7.3005
R14630 DFF_magic_0.tg_magic_3.CLK.t13 DFF_magic_0.tg_magic_3.CLK.n16 7.3005
R14631 DFF_magic_0.tg_magic_3.CLK.n9 DFF_magic_0.tg_magic_3.CLK.t21 7.3005
R14632 DFF_magic_0.tg_magic_3.CLK.t7 DFF_magic_0.tg_magic_3.CLK.n10 7.3005
R14633 DFF_magic_0.tg_magic_3.CLK.t14 DFF_magic_0.tg_magic_3.CLK.n8 7.3005
R14634 DFF_magic_0.tg_magic_3.CLK.n12 DFF_magic_0.tg_magic_3.CLK.n11 5.77618
R14635 DFF_magic_0.tg_magic_3.CLK.n17 DFF_magic_0.tg_magic_3.CLK.n15 5.67753
R14636 DFF_magic_0.tg_magic_3.CLK.n6 DFF_magic_0.tg_magic_3.CLK.n3 3.6455
R14637 DFF_magic_0.tg_magic_3.CLK.n6 DFF_magic_0.tg_magic_3.CLK.n5 3.31072
R14638 DFF_magic_0.tg_magic_3.CLK.n7 DFF_magic_0.tg_magic_3.CLK.n1 2.90572
R14639 DFF_magic_0.tg_magic_3.CLK.n1 DFF_magic_0.tg_magic_3.CLK.t4 1.6255
R14640 DFF_magic_0.tg_magic_3.CLK.n1 DFF_magic_0.tg_magic_3.CLK.n0 1.6255
R14641 DFF_magic_0.tg_magic_3.CLK.n5 DFF_magic_0.tg_magic_3.CLK.t5 1.6255
R14642 DFF_magic_0.tg_magic_3.CLK.n5 DFF_magic_0.tg_magic_3.CLK.n4 1.6255
R14643 DFF_magic_0.tg_magic_3.CLK.n3 DFF_magic_0.tg_magic_3.CLK.t1 1.463
R14644 DFF_magic_0.tg_magic_3.CLK.n3 DFF_magic_0.tg_magic_3.CLK.n2 1.463
R14645 DFF_magic_0.tg_magic_3.CLK.n18 DFF_magic_0.tg_magic_3.CLK 0.717689
R14646 DFF_magic_0.tg_magic_3.CLK.n7 DFF_magic_0.tg_magic_3.CLK.n6 0.4055
R14647 DFF_magic_0.tg_magic_3.CLK DFF_magic_0.tg_magic_3.CLK.n17 0.187712
R14648 DFF_magic_0.tg_magic_3.CLK DFF_magic_0.tg_magic_3.CLK.n12 0.185948
R14649 DFF_magic_0.tg_magic_3.CLK DFF_magic_0.tg_magic_3.CLK.n7 0.179883
R14650 DFF_magic_0.tg_magic_3.CLK DFF_magic_0.tg_magic_3.CLK.n18 0.104263
R14651 7b_counter_0.MDFF_7.QB.n5 7b_counter_0.MDFF_7.QB.t4 53.0329
R14652 7b_counter_0.MDFF_7.QB.t5 7b_counter_0.MDFF_7.QB.t6 44.058
R14653 7b_counter_0.MDFF_7.QB.n7 7b_counter_0.MDFF_7.QB.t8 38.8649
R14654 7b_counter_0.MDFF_7.QB.t8 7b_counter_0.MDFF_7.QB.t5 28.6791
R14655 7b_counter_0.MDFF_7.QB 7b_counter_0.MDFF_7.QB.n6 19.3781
R14656 7b_counter_0.MDFF_7.QB.n6 7b_counter_0.MDFF_7.QB.t10 17.2076
R14657 7b_counter_0.MDFF_7.QB.n6 7b_counter_0.MDFF_7.QB.t7 14.3398
R14658 7b_counter_0.MDFF_7.QB.n7 7b_counter_0.MDFF_7.QB.t9 7.3005
R14659 7b_counter_0.MDFF_7.QB.t7 7b_counter_0.MDFF_7.QB.n5 7.3005
R14660 7b_counter_0.MDFF_7.QB 7b_counter_0.MDFF_7.QB.n7 5.4249
R14661 7b_counter_0.MDFF_7.QB.n5 7b_counter_0.MDFF_7.QB.n4 4.57931
R14662 7b_counter_0.MDFF_7.QB.n4 7b_counter_0.MDFF_7.QB.n1 3.62007
R14663 7b_counter_0.MDFF_7.QB.n4 7b_counter_0.MDFF_7.QB.n3 3.15478
R14664 7b_counter_0.MDFF_7.QB.n3 7b_counter_0.MDFF_7.QB.t2 1.6255
R14665 7b_counter_0.MDFF_7.QB.n3 7b_counter_0.MDFF_7.QB.n2 1.6255
R14666 7b_counter_0.MDFF_7.QB.n1 7b_counter_0.MDFF_7.QB.t1 1.463
R14667 7b_counter_0.MDFF_7.QB.n1 7b_counter_0.MDFF_7.QB.n0 1.463
R14668 DFF_magic_0.tg_magic_1.IN.t14 DFF_magic_0.tg_magic_1.IN.t15 47.8944
R14669 DFF_magic_0.tg_magic_1.IN.n7 DFF_magic_0.tg_magic_1.IN.t17 38.7949
R14670 DFF_magic_0.tg_magic_1.IN.n8 DFF_magic_0.tg_magic_1.IN.t16 38.7949
R14671 DFF_magic_0.tg_magic_1.IN.n8 DFF_magic_0.tg_magic_1.IN.n7 31.4949
R14672 DFF_magic_0.tg_magic_1.IN.n9 DFF_magic_0.tg_magic_1.IN.t12 17.9416
R14673 DFF_magic_0.tg_magic_1.IN.n9 DFF_magic_0.tg_magic_1.IN.t14 11.957
R14674 DFF_magic_0.tg_magic_1.IN.n7 DFF_magic_0.tg_magic_1.IN.t13 7.3005
R14675 DFF_magic_0.tg_magic_1.IN.t12 DFF_magic_0.tg_magic_1.IN.n8 7.3005
R14676 DFF_magic_0.tg_magic_1.IN.n10 DFF_magic_0.tg_magic_1.IN 5.93058
R14677 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_1.IN.n9 5.86474
R14678 DFF_magic_0.tg_magic_1.IN.n2 DFF_magic_0.tg_magic_1.IN.t9 5.68507
R14679 DFF_magic_0.tg_magic_1.IN.n6 DFF_magic_0.tg_magic_1.IN.t7 4.92604
R14680 DFF_magic_0.tg_magic_1.IN.n17 DFF_magic_0.tg_magic_1.IN.n14 3.6455
R14681 DFF_magic_0.tg_magic_1.IN.n17 DFF_magic_0.tg_magic_1.IN.n16 3.31072
R14682 DFF_magic_0.tg_magic_1.IN.n5 DFF_magic_0.tg_magic_1.IN.n4 3.1505
R14683 DFF_magic_0.tg_magic_1.IN.n18 DFF_magic_0.tg_magic_1.IN.n12 2.90572
R14684 DFF_magic_0.tg_magic_1.IN.n2 DFF_magic_0.tg_magic_1.IN.n1 2.6005
R14685 DFF_magic_0.tg_magic_1.IN.n10 DFF_magic_0.tg_magic_1.IN 1.88467
R14686 DFF_magic_0.tg_magic_1.IN.n1 DFF_magic_0.tg_magic_1.IN.t11 1.6255
R14687 DFF_magic_0.tg_magic_1.IN.n1 DFF_magic_0.tg_magic_1.IN.n0 1.6255
R14688 DFF_magic_0.tg_magic_1.IN.n12 DFF_magic_0.tg_magic_1.IN.t2 1.6255
R14689 DFF_magic_0.tg_magic_1.IN.n12 DFF_magic_0.tg_magic_1.IN.n11 1.6255
R14690 DFF_magic_0.tg_magic_1.IN.n16 DFF_magic_0.tg_magic_1.IN.t5 1.6255
R14691 DFF_magic_0.tg_magic_1.IN.n16 DFF_magic_0.tg_magic_1.IN.n15 1.6255
R14692 DFF_magic_0.tg_magic_1.IN.n4 DFF_magic_0.tg_magic_1.IN.t6 1.463
R14693 DFF_magic_0.tg_magic_1.IN.n4 DFF_magic_0.tg_magic_1.IN.n3 1.463
R14694 DFF_magic_0.tg_magic_1.IN.n14 DFF_magic_0.tg_magic_1.IN.t0 1.463
R14695 DFF_magic_0.tg_magic_1.IN.n14 DFF_magic_0.tg_magic_1.IN.n13 1.463
R14696 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_1.IN.n10 1.33598
R14697 DFF_magic_0.tg_magic_1.IN.n6 DFF_magic_0.tg_magic_1.IN.n5 1.15166
R14698 DFF_magic_0.tg_magic_1.IN.n5 DFF_magic_0.tg_magic_1.IN.n2 0.898543
R14699 DFF_magic_0.tg_magic_1.IN.n18 DFF_magic_0.tg_magic_1.IN.n17 0.4055
R14700 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_1.IN.n6 0.198522
R14701 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_1.IN.n18 0.178625
R14702 p3_gen_magic_0.xnor_magic_1.OUT.t7 p3_gen_magic_0.xnor_magic_1.OUT.t6 44.058
R14703 p3_gen_magic_0.xnor_magic_1.OUT.n2 p3_gen_magic_0.xnor_magic_1.OUT.t5 38.8649
R14704 p3_gen_magic_0.xnor_magic_1.OUT.n3 p3_gen_magic_0.xnor_magic_1.OUT 31.5208
R14705 p3_gen_magic_0.xnor_magic_1.OUT.t5 p3_gen_magic_0.xnor_magic_1.OUT.t7 28.6791
R14706 p3_gen_magic_0.xnor_magic_1.OUT.n2 p3_gen_magic_0.xnor_magic_1.OUT.t4 7.3005
R14707 p3_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_1.OUT.n2 5.27587
R14708 p3_gen_magic_0.xnor_magic_1.OUT.n3 p3_gen_magic_0.xnor_magic_1.OUT.n1 4.11572
R14709 p3_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_1.OUT.n3 3.61488
R14710 p3_gen_magic_0.xnor_magic_1.OUT.n1 p3_gen_magic_0.xnor_magic_1.OUT.t1 1.463
R14711 p3_gen_magic_0.xnor_magic_1.OUT.n1 p3_gen_magic_0.xnor_magic_1.OUT.n0 1.463
R14712 7b_counter_0.MDFF_1.QB.n6 7b_counter_0.MDFF_1.QB.t10 53.2954
R14713 7b_counter_0.MDFF_1.QB.t5 7b_counter_0.MDFF_1.QB.t7 44.058
R14714 7b_counter_0.MDFF_1.QB.n0 7b_counter_0.MDFF_1.QB.t8 38.8649
R14715 7b_counter_0.MDFF_1.QB.t8 7b_counter_0.MDFF_1.QB.t5 28.6791
R14716 7b_counter_0.MDFF_1.QB 7b_counter_0.MDFF_1.QB.n7 19.3781
R14717 7b_counter_0.MDFF_1.QB.n7 7b_counter_0.MDFF_1.QB.t4 17.1425
R14718 7b_counter_0.MDFF_1.QB.n7 7b_counter_0.MDFF_1.QB.t6 14.405
R14719 7b_counter_0.MDFF_1.QB.n0 7b_counter_0.MDFF_1.QB.t9 7.3005
R14720 7b_counter_0.MDFF_1.QB.t6 7b_counter_0.MDFF_1.QB.n6 7.3005
R14721 7b_counter_0.MDFF_1.QB 7b_counter_0.MDFF_1.QB.n0 5.42776
R14722 7b_counter_0.MDFF_1.QB.n6 7b_counter_0.MDFF_1.QB.n5 4.51584
R14723 7b_counter_0.MDFF_1.QB.n5 7b_counter_0.MDFF_1.QB.n2 3.62007
R14724 7b_counter_0.MDFF_1.QB.n5 7b_counter_0.MDFF_1.QB.n4 3.15478
R14725 7b_counter_0.MDFF_1.QB.n4 7b_counter_0.MDFF_1.QB.t1 1.6255
R14726 7b_counter_0.MDFF_1.QB.n4 7b_counter_0.MDFF_1.QB.n3 1.6255
R14727 7b_counter_0.MDFF_1.QB.n2 7b_counter_0.MDFF_1.QB.t3 1.463
R14728 7b_counter_0.MDFF_1.QB.n2 7b_counter_0.MDFF_1.QB.n1 1.463
R14729 OR_magic_2.VOUT.t9 OR_magic_2.VOUT.t21 47.8944
R14730 OR_magic_2.VOUT.t17 OR_magic_2.VOUT.t3 47.8944
R14731 OR_magic_2.VOUT.t22 OR_magic_2.VOUT.t10 47.8944
R14732 OR_magic_2.VOUT.n1 OR_magic_2.VOUT.t25 38.7949
R14733 OR_magic_2.VOUT.n0 OR_magic_2.VOUT.t24 38.7949
R14734 OR_magic_2.VOUT.n4 OR_magic_2.VOUT.t12 38.7949
R14735 OR_magic_2.VOUT.n5 OR_magic_2.VOUT.t5 38.7949
R14736 OR_magic_2.VOUT.n10 OR_magic_2.VOUT.t18 38.7949
R14737 OR_magic_2.VOUT.n9 OR_magic_2.VOUT.t13 38.7949
R14738 OR_magic_2.VOUT.n12 OR_magic_2.VOUT.t6 36.2535
R14739 OR_magic_2.VOUT.n1 OR_magic_2.VOUT.n0 31.4949
R14740 OR_magic_2.VOUT.n5 OR_magic_2.VOUT.n4 31.4949
R14741 OR_magic_2.VOUT.n10 OR_magic_2.VOUT.n9 31.4949
R14742 OR_magic_2.VOUT.n7 OR_magic_2.VOUT.t8 26.9781
R14743 OR_magic_2.VOUT.n7 OR_magic_2.VOUT.t14 26.9781
R14744 OR_magic_2.VOUT.n8 OR_magic_2.VOUT.t16 26.9781
R14745 OR_magic_2.VOUT.n8 OR_magic_2.VOUT.t26 26.9781
R14746 OR_magic_2.VOUT.n3 OR_magic_2.VOUT.t20 20.2675
R14747 OR_magic_2.VOUT.n2 OR_magic_2.VOUT.t15 17.9416
R14748 OR_magic_2.VOUT.n6 OR_magic_2.VOUT.t11 17.9416
R14749 OR_magic_2.VOUT.n11 OR_magic_2.VOUT.t7 17.9416
R14750 OR_magic_2.VOUT.n2 OR_magic_2.VOUT.t9 11.957
R14751 OR_magic_2.VOUT.n6 OR_magic_2.VOUT.t17 11.957
R14752 OR_magic_2.VOUT.n11 OR_magic_2.VOUT.t22 11.957
R14753 OR_magic_2.VOUT.n14 OR_magic_2.VOUT.n13 10.5271
R14754 OR_magic_2.VOUT.n13 OR_magic_2.VOUT 8.06233
R14755 OR_magic_2.VOUT.n0 OR_magic_2.VOUT.t4 7.3005
R14756 OR_magic_2.VOUT.t15 OR_magic_2.VOUT.n1 7.3005
R14757 OR_magic_2.VOUT.n4 OR_magic_2.VOUT.t23 7.3005
R14758 OR_magic_2.VOUT.t11 OR_magic_2.VOUT.n5 7.3005
R14759 OR_magic_2.VOUT.t20 OR_magic_2.VOUT.n7 7.3005
R14760 OR_magic_2.VOUT.n9 OR_magic_2.VOUT.t19 7.3005
R14761 OR_magic_2.VOUT.t7 OR_magic_2.VOUT.n10 7.3005
R14762 OR_magic_2.VOUT.t6 OR_magic_2.VOUT.n8 7.3005
R14763 OR_magic_2.VOUT OR_magic_2.VOUT.n2 5.96162
R14764 OR_magic_2.VOUT.n12 OR_magic_2.VOUT.n11 5.77618
R14765 OR_magic_2.VOUT.n3 OR_magic_2.VOUT.n6 5.67753
R14766 OR_magic_2.VOUT OR_magic_2.VOUT.n14 1.45773
R14767 OR_magic_2.VOUT.n13 OR_magic_2.VOUT 0.81937
R14768 OR_magic_2.VOUT.n14 OR_magic_2.VOUT 0.35463
R14769 OR_magic_2.VOUT OR_magic_2.VOUT.n12 0.315078
R14770 OR_magic_2.VOUT OR_magic_2.VOUT.n3 0.227402
R14771 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t15 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t17 47.8944
R14772 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n7 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t13 38.7949
R14773 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n8 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t16 38.7949
R14774 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n8 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n7 31.4949
R14775 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n9 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t12 17.9416
R14776 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n9 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t15 11.957
R14777 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n7 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t14 7.3005
R14778 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t12 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n8 7.3005
R14779 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n10 7b_counter_0.DFF_magic_0.tg_magic_1.IN 5.93058
R14780 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n9 5.86474
R14781 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n2 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t9 5.68507
R14782 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n6 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t7 4.92604
R14783 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n15 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n12 3.6455
R14784 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n15 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n14 3.31072
R14785 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n5 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n4 3.1505
R14786 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n18 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n17 2.90572
R14787 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n2 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n1 2.6005
R14788 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n10 7b_counter_0.DFF_magic_0.tg_magic_1.IN 1.88467
R14789 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n1 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t11 1.6255
R14790 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n1 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n0 1.6255
R14791 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n14 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t2 1.6255
R14792 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n14 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n13 1.6255
R14793 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n17 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t5 1.6255
R14794 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n17 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n16 1.6255
R14795 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n4 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t6 1.463
R14796 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n4 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n3 1.463
R14797 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n12 7b_counter_0.DFF_magic_0.tg_magic_1.IN.t1 1.463
R14798 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n12 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n11 1.463
R14799 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n10 1.33598
R14800 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n6 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n5 1.15166
R14801 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n5 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n2 0.898543
R14802 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n18 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n15 0.4055
R14803 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n6 0.198522
R14804 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_1.IN.n18 0.178625
R14805 OUT1.n11 OUT1.n10 5.47387
R14806 OUT1.n12 OUT1.n8 4.65398
R14807 OUT1.n11 OUT1.n9 4.2255
R14808 OUT1 OUT1.n7 3.93486
R14809 OUT1.n7 OUT1.n1 2.2505
R14810 OUT1.n7 OUT1.n6 2.2505
R14811 OUT1.n3 OUT1.n2 1.49801
R14812 OUT1.n6 OUT1.n5 1.498
R14813 OUT1.n4 OUT1.n0 1.13034
R14814 OUT1.n5 OUT1.n4 1.12833
R14815 OUT1.n12 OUT1.n11 0.427022
R14816 OUT1 OUT1.n12 0.257096
R14817 OUT1.n5 OUT1.n3 0.0109978
R14818 OUT1.n6 OUT1.n2 0.00995968
R14819 OUT1.n4 OUT1.n1 0.00808653
R14820 OUT1.n3 OUT1.n0 0.0079912
R14821 OUT1.n7 OUT1.n0 0.0079912
R14822 OUT1.n2 OUT1.n1 0.00547984
R14823 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n7 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.t6 11.8647
R14824 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n2 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.t3 5.68507
R14825 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n11 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n10 5.47974
R14826 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n6 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.t0 4.928
R14827 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n12 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n8 4.77528
R14828 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n13 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.t7 4.52027
R14829 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n11 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n9 4.2255
R14830 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.t7 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n7 4.2255
R14831 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n5 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n4 3.1505
R14832 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n2 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n1 2.6005
R14833 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n1 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.t5 1.6255
R14834 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n1 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n0 1.6255
R14835 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n4 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.t1 1.463
R14836 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n4 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n3 1.463
R14837 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n6 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n5 1.16072
R14838 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n5 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n2 0.898543
R14839 p2_gen_magic_0.3_inp_AND_magic_0.VOUT p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n14 0.5135
R14840 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n14 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n13 0.3875
R14841 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n12 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n11 0.305717
R14842 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n14 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n7 0.299848
R14843 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n13 p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n12 0.244879
R14844 p2_gen_magic_0.3_inp_AND_magic_0.VOUT p2_gen_magic_0.3_inp_AND_magic_0.VOUT.n6 0.235505
R14845 7b_counter_0.MDFF_5.QB.n5 7b_counter_0.MDFF_5.QB.t10 53.2571
R14846 7b_counter_0.MDFF_5.QB.t4 7b_counter_0.MDFF_5.QB.t8 44.058
R14847 7b_counter_0.MDFF_5.QB.n7 7b_counter_0.MDFF_5.QB.t7 38.8649
R14848 7b_counter_0.MDFF_5.QB.t7 7b_counter_0.MDFF_5.QB.t4 28.6791
R14849 7b_counter_0.MDFF_5.QB 7b_counter_0.MDFF_5.QB.n6 19.3781
R14850 7b_counter_0.MDFF_5.QB.n6 7b_counter_0.MDFF_5.QB.t9 17.1425
R14851 7b_counter_0.MDFF_5.QB.n6 7b_counter_0.MDFF_5.QB.t6 14.405
R14852 7b_counter_0.MDFF_5.QB.n7 7b_counter_0.MDFF_5.QB.t5 7.3005
R14853 7b_counter_0.MDFF_5.QB.t6 7b_counter_0.MDFF_5.QB.n5 7.3005
R14854 7b_counter_0.MDFF_5.QB 7b_counter_0.MDFF_5.QB.n7 5.4273
R14855 7b_counter_0.MDFF_5.QB.n5 7b_counter_0.MDFF_5.QB.n4 4.57931
R14856 7b_counter_0.MDFF_5.QB.n4 7b_counter_0.MDFF_5.QB.n1 3.62007
R14857 7b_counter_0.MDFF_5.QB.n4 7b_counter_0.MDFF_5.QB.n3 3.15478
R14858 7b_counter_0.MDFF_5.QB.n3 7b_counter_0.MDFF_5.QB.t1 1.6255
R14859 7b_counter_0.MDFF_5.QB.n3 7b_counter_0.MDFF_5.QB.n2 1.6255
R14860 7b_counter_0.MDFF_5.QB.n1 7b_counter_0.MDFF_5.QB.t3 1.463
R14861 7b_counter_0.MDFF_5.QB.n1 7b_counter_0.MDFF_5.QB.n0 1.463
R14862 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n3 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t10 130.41
R14863 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n7 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t7 35.3186
R14864 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n4 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t4 33.5023
R14865 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t11 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n4 33.5023
R14866 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n2 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t5 32.2349
R14867 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n7 31.543
R14868 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n6 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t3 19.0138
R14869 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n5 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t11 16.3421
R14870 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t3 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n3 13.2317
R14871 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n3 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n2 13.0005
R14872 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n5 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t9 11.3624
R14873 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n2 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t8 11.146
R14874 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n4 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t12 7.3005
R14875 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n7 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t6 7.3005
R14876 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n0 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t0 5.47387
R14877 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n1 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t1 4.65398
R14878 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n0 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t2 4.2255
R14879 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n6 3.63214
R14880 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n6 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n5 3.62977
R14881 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n1 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n0 0.427022
R14882 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n1 0.257096
C0 7b_counter_0.MDFF_5.tspc2_magic_0.Q 7b_counter_0.MDFF_5.LD 0.12f
C1 a_26126_1124# CLK 0.0622f
C2 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A Q1 2.58e-19
C3 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A VDD 1.37f
C4 a_5036_n8579# VDD 0.476f
C5 a_5054_n1526# D2_3 0.229f
C6 7b_counter_0.MDFF_6.tspc2_magic_0.Q VDD 1.18f
C7 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A 0.00618f
C8 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B 0.0069f
C9 a_30365_3514# P2 0.477f
C10 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B 0.00112f
C11 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 2.27e-20
C12 p3_gen_magic_0.xnor_magic_4.OUT a_11708_n6613# 0.0456f
C13 a_2749_10148# a_2749_8740# 0.475f
C14 a_1209_6275# a_1209_4557# 0.00776f
C15 Q1 D2_4 0.0738f
C16 7b_counter_0.MDFF_7.tspc2_magic_0.CLK D2_4 0.249f
C17 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A CLK 0.00307f
C18 7b_counter_0.MDFF_6.tspc2_magic_0.Q D2_1 0.169f
C19 a_13353_n2115# p2_gen_magic_0.3_inp_AND_magic_0.VOUT 0.115f
C20 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_12174_n4081# 0.0815f
C21 7b_counter_0.3_inp_AND_magic_0.A Q1 1.15e-19
C22 7b_counter_0.3_inp_AND_magic_0.A 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 2.83e-20
C23 a_5185_7469# Q6 2.54e-19
C24 a_12387_8536# a_12931_8580# 0.298f
C25 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 7b_counter_0.DFF_magic_0.tg_magic_2.IN 0.694f
C26 a_12174_n7648# a_12174_n8095# 0.0139f
C27 a_27234_552# DFF_magic_0.tg_magic_3.OUT 0.00293f
C28 a_14556_n3644# Q4 0.0188f
C29 a_27234_1746# Q3 4.62e-19
C30 a_23560_3728# Q3 0.00422f
C31 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.3_inp_AND_magic_0.A 0.91f
C32 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.3_inp_AND_magic_0.B 0.00468f
C33 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_6.OUT 5.45e-19
C34 7b_counter_0.3_inp_AND_magic_0.C Q4 0.0696f
C35 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_19841_8580# 6.68e-20
C36 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_12387_5769# 1.37e-19
C37 a_12387_1746# a_12931_2253# 0.298f
C38 a_1559_n6471# a_1975_n6471# 0.00222f
C39 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN 0.654f
C40 a_17405_684# Q1 0.00119f
C41 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT 0.246f
C42 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B Q5 0.0215f
C43 7b_counter_0.MDFF_6.tspc2_magic_0.Q LD 7.02e-19
C44 p2_gen_magic_0.3_inp_AND_magic_0.C p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 1.07e-19
C45 a_4235_3947# D2_5 0.0338f
C46 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A Q3 2.33e-19
C47 Q1 Q2 0.505f
C48 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A a_1409_6275# 0.0292f
C49 7b_counter_0.MDFF_7.tspc2_magic_0.D a_23560_3728# 0.0379f
C50 a_5036_n8095# Q5 5.75e-19
C51 p2_gen_magic_0.xnor_magic_3.OUT D2_7 0.0475f
C52 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_9412_739# 1.29e-19
C53 a_30365_3514# VDD 1.16f
C54 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 4.89e-20
C55 a_1209_1059# a_1559_n1042# 6.47e-20
C56 a_23802_2253# VDD 0.0879f
C57 a_9212_739# D2_6 0.0646f
C58 a_1409_3363# VDD 0.0124f
C59 a_11191_684# p2_gen_magic_0.xnor_magic_0.OUT 2.52e-20
C60 a_5036_n7648# Q6 0.315f
C61 7b_counter_0.3_inp_AND_magic_0.VOUT D2_4 0.0316f
C62 a_23793_5904# VDD 1.08f
C63 7b_counter_0.3_inp_AND_magic_0.VOUT 7b_counter_0.3_inp_AND_magic_0.A 0.00143f
C64 a_12931_8580# VDD 0.0124f
C65 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B D2_4 0.0113f
C66 a_1209_7469# a_2749_5900# 1.14e-19
C67 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_1209_8579# 4.8e-20
C68 mux_magic_0.AND2_magic_0.A mux_magic_0.OR_magic_0.A 0.00108f
C69 a_1559_n1973# a_1975_n1973# 0.00222f
C70 a_19841_3363# a_19152_1223# 3.03e-19
C71 a_17405_7309# 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 2.4e-20
C72 a_2749_684# VDD 1.55f
C73 a_11279_1124# VDD 0.936f
C74 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT VDD 1.07f
C75 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 0.162f
C76 divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT VDD 1.09f
C77 p3_gen_magic_0.3_inp_AND_magic_0.C p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.00142f
C78 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B VDD 1.2f
C79 7b_counter_0.MDFF_4.LD a_12387_3319# 0.195f
C80 a_2749_7308# CLK 0.0106f
C81 7b_counter_0.MDFF_4.LD a_27234_1746# 0.195f
C82 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B Q4 0.00109f
C83 7b_counter_0.MDFF_4.LD a_23560_3728# 0.00691f
C84 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B 0.00112f
C85 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 0.00315f
C86 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_1 5.89e-19
C87 7b_counter_0.3_inp_AND_magic_0.VOUT Q2 3.64e-20
C88 7b_counter_0.MDFF_4.LD 7b_counter_0.DFF_magic_0.tg_magic_0.IN 5.63e-20
C89 a_1409_3363# LD 0.0292f
C90 a_7303_3480# Q7 0.0391f
C91 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A a_20041_3363# 5.46e-20
C92 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B D2_1 0.0061f
C93 a_16065_4557# CLK 0.00454f
C94 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A 0.00618f
C95 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_11279_6341# 0.00904f
C96 p3_gen_magic_0.3_inp_AND_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK 0.244f
C97 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT D2_3 0.00103f
C98 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A 1.1e-20
C99 a_21381_3524# Q5 0.00555f
C100 a_5036_n8095# Q2 6.69e-21
C101 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN VDD 1.18f
C102 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT a_8939_n3150# 0.00157f
C103 a_2749_684# LD 0.00267f
C104 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT a_12174_n8095# 0.0834f
C105 a_6725_7308# Q2 4.35e-19
C106 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A 0.443f
C107 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A Q1 0.00809f
C108 7b_counter_0.DFF_magic_0.D 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 0.846f
C109 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A D2_5 4.23e-19
C110 7b_counter_0.MDFF_4.tspc2_magic_0.CLK VDD 2.18f
C111 a_27234_3319# D2_4 0.241f
C112 a_9212_739# D2_2 9.14e-19
C113 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN D2_1 0.00752f
C114 a_12387_4513# Q1 8.5e-19
C115 a_5185_2253# a_6725_2092# 0.00114f
C116 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A a_20041_3363# 1.77e-19
C117 a_1541_n8579# VDD 0.415f
C118 a_30365_4922# P2 0.173f
C119 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A 3.81e-19
C120 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A 0.00108f
C121 p3_gen_magic_0.3_inp_AND_magic_0.C Q4 0.161f
C122 p3_gen_magic_0.xnor_magic_4.OUT a_11492_n6613# 0.104f
C123 7b_counter_0.DFF_magic_0.Q 7b_counter_0.MDFF_5.LD 0.169f
C124 7b_counter_0.MDFF_4.tspc2_magic_0.Q Q6 2.13e-19
C125 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A Q1 0.00434f
C126 a_15865_7470# 7b_counter_0.MDFF_6.tspc2_magic_0.D 7.57e-20
C127 a_12174_n3150# a_12174_n3597# 0.0139f
C128 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A a_15865_3363# 1.03e-19
C129 p3_gen_magic_0.AND2_magic_1.A a_12590_n7648# 0.0629f
C130 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A Q1 0.0462f
C131 a_12174_n3597# Q4 0.0843f
C132 a_23802_2253# Q3 4.83e-19
C133 a_23793_5904# Q3 0.00192f
C134 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 0.412f
C135 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A a_8411_3319# 1.03e-19
C136 p2_gen_magic_0.xnor_magic_1.OUT Q5 0.00362f
C137 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B a_17405_4932# 0.173f
C138 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_15865_1059# 1.37e-19
C139 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT a_5452_n7648# 6.1e-19
C140 OR_magic_2.VOUT divide_by_2_0.tg_magic_3.IN 0.619f
C141 p3_gen_magic_0.xnor_magic_3.OUT a_11292_n6613# 0.483f
C142 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_5.OUT 5.37e-19
C143 a_2749_684# Q3 3.98e-19
C144 7b_counter_0.MDFF_3.tspc2_magic_0.Q CLK 0.0529f
C145 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B Q2 8.2e-19
C146 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A a_1209_6275# 0.251f
C147 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8643_n1526# 0.0827f
C148 a_15865_1059# Q4 6.05e-19
C149 p3_gen_magic_0.3_inp_AND_magic_0.VOUT VDD 2.16f
C150 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B 0.00594f
C151 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B VDD 1.2f
C152 a_30365_4922# VDD 1.59f
C153 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK a_16386_n8142# 0.016f
C154 a_19152_1223# VDD 0.759f
C155 a_8411_3319# VDD 0.982f
C156 p2_gen_magic_0.xnor_magic_1.OUT D2_4 0.248f
C157 p3_gen_magic_0.3_inp_AND_magic_0.VOUT D2_1 0.00935f
C158 a_21504_5904# VDD 1.11f
C159 7b_counter_0.DFF_magic_0.Q 7b_counter_0.3_inp_AND_magic_0.B 0.00209f
C160 p2_gen_magic_0.xnor_magic_4.OUT a_5036_n3597# 0.00929f
C161 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_6 0.127f
C162 a_23985_7877# VDD 1.21f
C163 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A a_1409_4557# 9.27e-19
C164 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 0.179f
C165 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_5 0.0103f
C166 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A a_16065_4557# 9.27e-19
C167 a_6725_5900# a_5185_6275# 7.98e-19
C168 OR_magic_2.A a_30365_3514# 0.0435f
C169 p3_gen_magic_0.xnor_magic_4.OUT a_5054_n5540# 0.297f
C170 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_3.IN 0.797f
C171 a_6725_2092# VDD 0.943f
C172 7b_counter_0.MDFF_5.LD D2_4 0.103f
C173 7b_counter_0.MDFF_4.LD a_30365_3514# 4.86e-20
C174 a_16065_7470# VDD 0.0191f
C175 7b_counter_0.MDFF_4.tspc2_magic_0.CLK Q3 4.75e-19
C176 a_1409_2253# Q4 0.002f
C177 7b_counter_0.MDFF_4.LD a_23802_2253# 0.0279f
C178 7b_counter_0.MDFF_5.LD 7b_counter_0.3_inp_AND_magic_0.A 8.74e-20
C179 p2_gen_magic_0.AND2_magic_1.A a_11292_n6613# 1.68e-19
C180 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A a_11279_3480# 2.4e-20
C181 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_20171_1669# 5.37e-19
C182 p2_gen_magic_0.xnor_magic_1.OUT Q2 0.0181f
C183 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT 0.00275f
C184 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A Q7 0.0252f
C185 a_16065_7470# D2_1 0.168f
C186 mux_magic_0.IN1 divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT 0.004f
C187 a_23985_7877# LD 0.0102f
C188 a_13353_n6613# p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK 9.82e-21
C189 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A 0.00108f
C190 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_1209_6275# 1.63e-20
C191 a_5054_n1042# D2_3 0.0088f
C192 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT a_12174_n3597# 0.0834f
C193 p3_gen_magic_0.xnor_magic_1.B Q4 0.00258f
C194 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 0.00325f
C195 a_8713_1625# D2_3 2.66e-19
C196 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.xnor_magic_5.OUT 0.00433f
C197 7b_counter_0.3_inp_AND_magic_0.B Q5 8.09e-19
C198 a_13769_n6613# VDD 0.0206f
C199 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A a_1559_n1042# 6.06e-20
C200 p2_gen_magic_0.3_inp_AND_magic_0.B Q4 0.0509f
C201 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A a_21381_3524# 2.4e-20
C202 a_15865_4557# Q1 8.5e-19
C203 7b_counter_0.MDFF_5.LD Q2 3.8f
C204 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B 0.00121f
C205 a_17405_4932# VDD 1.55f
C206 a_9689_6886# D2_6 0.00514f
C207 7b_counter_0.MDFF_6.tspc2_magic_0.D a_19152_6440# 0.037f
C208 a_24536_3947# D2_4 0.00993f
C209 divide_by_2_1.tg_magic_2.IN VDD 1.22f
C210 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A a_12931_4557# 0.0292f
C211 7b_counter_0.MDFF_5.tspc2_magic_0.Q a_8411_4513# 1.1e-19
C212 a_8643_n5540# Q1 0.0138f
C213 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_2 0.926f
C214 a_16386_n8142# VDD 0.0248f
C215 DFF_magic_0.tg_magic_2.OUT P2 0.0139f
C216 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A Q7 0.0843f
C217 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A VDD 1.23f
C218 p2_gen_magic_0.AND2_magic_1.A a_12590_n3150# 0.0629f
C219 a_16386_n8142# D2_1 0.00483f
C220 7b_counter_0.3_inp_AND_magic_0.B D2_4 0.00634f
C221 a_19841_8580# Q1 0.00342f
C222 a_15865_9774# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A 0.128f
C223 a_23352_n6798# CLK 2.13e-20
C224 7b_counter_0.3_inp_AND_magic_0.A 7b_counter_0.3_inp_AND_magic_0.B 0.254f
C225 a_17405_3524# Q1 0.017f
C226 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 0.0847f
C227 a_8939_n7648# a_8523_n8095# 0.013f
C228 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A a_21381_3524# 0.0334f
C229 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B Q3 0.0177f
C230 a_19152_1223# Q3 8.01e-20
C231 7b_counter_0.MDFF_4.tspc2_magic_0.Q a_8955_3363# 0.017f
C232 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A a_1409_8579# 7.81e-19
C233 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT a_5452_n3150# 6.1e-19
C234 a_21504_5904# Q3 0.191f
C235 7b_counter_0.MDFF_3.tspc2_magic_0.Q 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 6.87e-19
C236 a_23985_7877# Q3 0.00167f
C237 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A Q1 0.00647f
C238 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B Q6 0.00143f
C239 a_1559_n6024# a_1975_n6471# 0.013f
C240 Q7 D2_6 0.0788f
C241 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_27234_3319# 0.125f
C242 OR_magic_2.VOUT a_23352_n6798# 0.12f
C243 a_4235_9163# CLK 0.00818f
C244 a_1409_4557# D2_5 0.00471f
C245 7b_counter_0.3_inp_AND_magic_0.B Q2 0.176f
C246 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.3_inp_AND_magic_0.A 0.0111f
C247 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A LD 0.00221f
C248 a_13353_n6613# VDD 1.23f
C249 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT a_5054_n5540# 7.56e-21
C250 a_9689_6886# D2_2 3.14e-21
C251 p3_gen_magic_0.xnor_magic_5.OUT VDD 2.24f
C252 7b_counter_0.3_inp_AND_magic_0.VOUT a_24401_7877# 0.192f
C253 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A a_11191_4932# 1.51e-21
C254 DFF_magic_0.tg_magic_2.OUT VDD 1.23f
C255 a_26126_3480# VDD 0.943f
C256 a_18891_1669# VDD 0.969f
C257 a_5054_n5540# Q6 0.0445f
C258 mux_magic_0.AND2_magic_0.A mux_magic_0.IN2 0.0162f
C259 a_13353_n6613# D2_1 0.0078f
C260 a_1541_n3150# D2_4 0.0409f
C261 p2_gen_magic_0.xnor_magic_5.OUT D2_3 0.132f
C262 OR_magic_1.VOUT divide_by_2_1.tg_magic_3.CLK 0.566f
C263 divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT VDD 1.09f
C264 a_19152_5956# VDD 0.721f
C265 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.AND2_magic_1.A 2.36e-19
C266 p3_gen_magic_0.3_inp_AND_magic_0.B p3_gen_magic_0.AND2_magic_1.A 0.00771f
C267 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_5.tspc2_magic_0.D 0.00171f
C268 p3_gen_magic_0.xnor_magic_5.OUT D2_1 0.00389f
C269 DFF_magic_0.tg_magic_2.OUT D2_1 0.00225f
C270 a_2749_2092# D2_4 0.00422f
C271 a_1559_n1526# a_1975_n1973# 0.013f
C272 OR_magic_2.A a_30365_4922# 0.297f
C273 a_23560_3728# a_23802_2253# 5.39e-19
C274 divide_by_2_1.tg_magic_1.IN a_34156_n889# 5.83e-20
C275 7b_counter_0.MDFF_6.tspc2_magic_0.CLK Q6 2.96e-19
C276 a_5185_1059# D2_3 0.00246f
C277 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B 0.00561f
C278 a_23793_5904# a_23560_3728# 4.74e-19
C279 a_12931_7470# VDD 0.00388f
C280 7b_counter_0.MDFF_4.LD a_30365_4922# 0.0254f
C281 7b_counter_0.MDFF_4.tspc2_magic_0.D a_12387_552# 1.63e-20
C282 DFF_magic_0.D a_27778_3363# 0.00228f
C283 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_5515_3947# 0.112f
C284 7b_counter_0.MDFF_4.LD a_19152_1223# 0.00678f
C285 a_17405_7309# 7b_counter_0.MDFF_6.tspc2_magic_0.D 0.123f
C286 a_9212_5956# a_9689_6886# 0.153f
C287 7b_counter_0.MDFF_4.LD a_8411_3319# 0.195f
C288 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_19307_1669# 0.00409f
C289 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A a_23258_552# 0.251f
C290 7b_counter_0.MDFF_5.LD a_8955_8580# 0.0279f
C291 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A a_11191_4932# 3.58e-20
C292 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A VDD 1.3f
C293 a_15865_9774# Q7 7.52e-19
C294 7b_counter_0.MDFF_7.tspc2_magic_0.Q a_23258_1746# 0.0276f
C295 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1975_n6471# 6.1e-19
C296 D2_2 Q7 0.0683f
C297 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A P2 5.23e-20
C298 p2_gen_magic_0.3_inp_AND_magic_0.C p2_gen_magic_0.xnor_magic_6.OUT 0.0267f
C299 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 0.0847f
C300 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A a_1409_1059# 9.27e-19
C301 7b_counter_0.DFF_magic_0.D DFF_magic_0.D 0.00552f
C302 a_13553_n6613# VDD 0.0178f
C303 a_11279_3480# Q1 0.00512f
C304 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B D2_7 0.00401f
C305 a_8825_6886# D2_6 4.84e-19
C306 a_7303_8697# Q2 0.161f
C307 7b_counter_0.MDFF_4.tspc2_magic_0.D p2_gen_magic_0.xnor_magic_3.OUT 2.45e-19
C308 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN 0.164f
C309 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A CLK 0.00118f
C310 7b_counter_0.MDFF_6.tspc2_magic_0.D a_18891_6886# 0.278f
C311 p2_gen_magic_0.xnor_magic_0.OUT a_11292_n2115# 0.379f
C312 7b_counter_0.DFF_magic_0.Q 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 0.0315f
C313 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.xnor_magic_3.OUT 0.88f
C314 a_27234_4513# VDD 0.975f
C315 a_11279_1124# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A 0.0334f
C316 a_23672_3947# D2_4 6.09e-19
C317 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A D2_3 0.0293f
C318 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A Q7 0.096f
C319 a_14756_n8142# VDD 0.0541f
C320 p3_gen_magic_0.xnor_magic_6.OUT D2_6 0.375f
C321 a_5054_n1973# a_5036_n3150# 0.0732f
C322 a_8643_n1973# p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT 7.47e-19
C323 p3_gen_magic_0.AND2_magic_1.A D2_5 0.191f
C324 a_8713_6842# Q6 1.07e-20
C325 7b_counter_0.MDFF_0.tspc2_magic_0.D D2_5 0.00383f
C326 a_19841_4557# a_19841_3363# 0.00638f
C327 a_14756_n3644# D2_3 0.0266f
C328 a_17405_4932# a_15865_3363# 1.14e-19
C329 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_12387_3319# 1.08e-19
C330 a_27234_4513# a_27778_4557# 0.297f
C331 p3_gen_magic_0.xnor_magic_4.OUT a_8643_n6471# 7.33e-19
C332 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_0.OUT 7.63e-21
C333 a_8939_n3150# a_8523_n3597# 0.013f
C334 a_5185_7469# VDD 1.02f
C335 mux_magic_0.IN1 divide_by_2_1.tg_magic_2.IN 0.303f
C336 p3_gen_magic_0.xnor_magic_1.OUT Q4 4.22e-19
C337 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A Q7 0.0126f
C338 a_2749_3524# a_2749_2092# 0.00112f
C339 a_5054_n6024# p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT 7.12e-21
C340 a_8955_9774# D2_2 0.00581f
C341 a_23352_n6798# p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN 0.00396f
C342 a_12931_4557# Q1 6.2e-19
C343 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A VDD 1.3f
C344 7b_counter_0.MDFF_4.LD a_17405_4932# 0.00267f
C345 a_12174_n7648# a_12590_n7648# 0.00222f
C346 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A Q7 0.0249f
C347 a_9689_6886# CLK 0.00191f
C348 p2_gen_magic_0.3_inp_AND_magic_0.C VDD 2.55f
C349 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A CLK 0.0296f
C350 Q5 D2_5 1.15f
C351 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B D2_6 0.0068f
C352 a_19841_9774# Q1 1.63e-20
C353 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT Q4 1.93e-19
C354 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A a_2749_3524# 0.0334f
C355 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A 0.0037f
C356 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A DFF_magic_0.tg_magic_3.OUT 0.0012f
C357 a_19152_6440# Q7 4.12e-19
C358 a_1559_n6024# a_1559_n6471# 0.0142f
C359 7b_counter_0.MDFF_1.tspc2_magic_0.Q Q5 0.476f
C360 a_1957_n3150# Q7 0.00335f
C361 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN D2_6 0.0101f
C362 p2_gen_magic_0.3_inp_AND_magic_0.C D2_1 0.00476f
C363 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT a_1957_n7648# 6.1e-19
C364 7b_counter_0.MDFF_5.tspc2_magic_0.D D2_6 0.0792f
C365 7b_counter_0.MDFF_7.tspc2_magic_0.D a_26126_3480# 0.123f
C366 a_5185_7469# LD 0.195f
C367 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A a_17405_8741# 0.0334f
C368 a_8825_6886# D2_2 4.39e-19
C369 a_5036_n7648# VDD 0.0434f
C370 7b_counter_0.3_inp_AND_magic_0.VOUT a_24185_7877# 1.9e-20
C371 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT Q5 0.00576f
C372 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK a_16186_n8142# 0.00336f
C373 a_11191_684# VDD 1.55f
C374 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A Q3 5.49e-20
C375 a_24259_4877# VDD 0.728f
C376 D2_5 D2_4 0.0802f
C377 D2_6 D2_3 0.66f
C378 a_5036_n3150# D2_3 1.85e-19
C379 a_16065_6276# VDD 0.0609f
C380 7b_counter_0.DFF_magic_0.tg_magic_3.CLK D2_4 0.0288f
C381 p3_gen_magic_0.xnor_magic_6.OUT D2_2 5.59e-20
C382 7b_counter_0.MDFF_1.tspc2_magic_0.Q D2_4 0.00648f
C383 a_8411_4513# a_7215_4932# 7.98e-19
C384 a_1209_4557# a_1409_4557# 0.297f
C385 p2_gen_magic_0.3_inp_AND_magic_0.A Q5 7.55e-20
C386 CLK Q7 0.864f
C387 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A a_8955_9774# 0.0292f
C388 7b_counter_0.3_inp_AND_magic_0.A 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 2.7e-20
C389 a_1559_n1526# a_1559_n1973# 0.0142f
C390 a_8411_4513# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A 0.128f
C391 a_16065_6276# D2_1 0.00452f
C392 a_27234_1746# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B 0.125f
C393 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_5.OUT 5.24e-19
C394 OR_magic_2.A DFF_magic_0.tg_magic_2.OUT 0.318f
C395 a_15865_7470# D2_3 0.002f
C396 p3_gen_magic_0.xnor_magic_1.B p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 0.00195f
C397 DFF_magic_0.tg_magic_0.IN DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 4.89e-20
C398 a_9212_5956# a_8825_6886# 0.00652f
C399 7b_counter_0.MDFF_4.LD a_18891_1669# 1.61e-20
C400 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_4651_3947# 0.0618f
C401 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A a_6725_5900# 3.58e-20
C402 p3_gen_magic_0.xnor_magic_4.OUT Q1 0.34f
C403 7b_counter_0.MDFF_5.LD a_19841_8580# 0.195f
C404 Q2 D2_5 0.0947f
C405 D2_7 Q5 0.42f
C406 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B D2_2 0.023f
C407 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1559_n6471# 0.102f
C408 a_11279_8697# Q7 0.00668f
C409 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_3.OUT 2.35e-19
C410 p2_gen_magic_0.3_inp_AND_magic_0.A D2_4 0.00729f
C411 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.xnor_magic_5.OUT 5.85e-19
C412 a_11292_n6613# Q4 4.98e-19
C413 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A a_1209_9773# 0.25f
C414 7b_counter_0.MDFF_5.tspc2_magic_0.D D2_2 0.0123f
C415 divide_by_2_0.tg_magic_2.IN VDD 1.23f
C416 7b_counter_0.MDFF_4.tspc2_magic_0.Q 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 0.255f
C417 7b_counter_0.MDFF_5.LD a_17405_10149# 0.0332f
C418 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A a_1209_1059# 0.128f
C419 a_27234_4513# 7b_counter_0.MDFF_7.tspc2_magic_0.D 1.63e-20
C420 p3_gen_magic_0.3_inp_AND_magic_0.A p3_gen_magic_0.3_inp_AND_magic_0.B 0.318f
C421 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B Q6 6.05e-19
C422 a_8643_n6024# D2_6 7.09e-20
C423 a_11708_n6613# VDD 0.0137f
C424 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT a_12590_n7648# 0.00157f
C425 a_11191_4932# Q1 0.00215f
C426 7b_counter_0.3_inp_AND_magic_0.C Q7 1.73e-19
C427 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A Q3 0.00169f
C428 a_1409_7469# D2_7 0.0346f
C429 a_8955_9774# CLK 4.55e-19
C430 a_19841_4557# VDD 0.988f
C431 p2_gen_magic_0.3_inp_AND_magic_0.C Q3 0.197f
C432 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT D2_7 0.0248f
C433 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A 0.401f
C434 D2_2 D2_3 0.0996f
C435 D2_7 D2_4 0.937f
C436 divide_by_2_1.tg_magic_1.IN mux_magic_0.OR_magic_0.B 9.17e-20
C437 DFF_magic_0.tg_magic_3.CLK DFF_magic_0.tg_magic_3.OUT 0.528f
C438 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT a_23352_n5390# 1.09e-19
C439 p2_gen_magic_0.xnor_magic_6.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 2.61e-19
C440 7b_counter_0.MDFF_0.tspc2_magic_0.Q Q4 0.00136f
C441 a_8523_n7648# D2_6 0.0571f
C442 a_16186_n8142# VDD 0.895f
C443 a_8643_n1526# D2_6 0.0168f
C444 7b_counter_0.MDFF_4.tspc2_magic_0.Q VDD 1.23f
C445 a_2749_3524# D2_5 0.0422f
C446 a_23207_5815# Q1 0.00574f
C447 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A CLK 0.0197f
C448 7b_counter_0.3_inp_AND_magic_0.B a_24401_7877# 0.0502f
C449 a_2749_5900# Q6 0.0148f
C450 p3_gen_magic_0.xnor_magic_0.OUT D2_6 0.0156f
C451 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT Q5 0.0014f
C452 7b_counter_0.MDFF_5.tspc2_magic_0.D a_9212_5956# 0.278f
C453 a_12174_n3150# a_12590_n3150# 0.00222f
C454 a_16186_n8142# D2_1 0.00993f
C455 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 0.00186f
C456 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_4496_4393# 0.00119f
C457 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B a_7303_3480# 0.412f
C458 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_20041_8580# 0.00741f
C459 a_22150_1124# VDD 1.02f
C460 7b_counter_0.MDFF_4.LD a_27234_4513# 3.96e-19
C461 a_16065_3363# Q2 0.002f
C462 7b_counter_0.3_inp_AND_magic_0.VOUT DFF_magic_0.D 2.51e-20
C463 a_8825_6886# CLK 0.00221f
C464 a_12590_n3150# Q4 0.0034f
C465 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_14756_n8142# 7.91e-19
C466 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.0032f
C467 a_23258_552# CLK 0.0437f
C468 p3_gen_magic_0.xnor_magic_4.OUT a_5036_n8095# 0.0164f
C469 Q2 D2_7 2.13f
C470 7b_counter_0.MDFF_1.tspc2_magic_0.D a_19307_1669# 0.00451f
C471 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_21504_5904# 0.0222f
C472 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_15865_8580# 1.08e-19
C473 a_21381_10149# a_19841_8580# 1.14e-19
C474 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_11279_1124# 0.0183f
C475 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A a_2749_4932# 0.397f
C476 a_1209_4557# 7b_counter_0.MDFF_0.tspc2_magic_0.D 1.63e-20
C477 a_17405_2092# 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 2.4e-20
C478 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B a_19152_739# 1.29e-19
C479 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_1.tspc2_magic_0.Q 0.252f
C480 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_4 0.00688f
C481 a_1409_9773# CLK 4.61e-19
C482 mux_magic_0.IN2 OR_magic_2.VOUT 3.1e-19
C483 a_8411_8536# a_8713_6842# 3.03e-19
C484 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B Q7 0.027f
C485 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B a_19841_3363# 0.125f
C486 a_8643_n6024# D2_2 0.237f
C487 p3_gen_magic_0.3_inp_AND_magic_0.A D2_5 0.06f
C488 a_12387_552# Q4 0.00131f
C489 7b_counter_0.MDFF_3.QB a_5185_7469# 2.1e-19
C490 7b_counter_0.MDFF_7.tspc2_magic_0.D a_24259_4877# 0.103f
C491 a_2749_7308# a_1209_6275# 7.16e-20
C492 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A 8.54e-19
C493 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT a_11292_n6613# 3.07e-20
C494 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT VDD 1.17f
C495 a_1957_n7648# VDD 0.0018f
C496 7b_counter_0.MDFF_4.LD p2_gen_magic_0.3_inp_AND_magic_0.C 9.66e-19
C497 7b_counter_0.MDFF_0.tspc2_magic_0.CLK Q7 0.0465f
C498 a_32616_n1264# a_32616_n2458# 0.00638f
C499 a_1409_1059# VDD 0.0559f
C500 a_24059_4877# VDD 0.976f
C501 a_19152_6440# D2_3 0.0264f
C502 a_15865_6276# VDD 0.988f
C503 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A a_27778_2253# 1.77e-19
C504 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT D2_1 8.45e-19
C505 a_12387_6963# 7b_counter_0.MDFF_5.tspc2_magic_0.D 7.57e-20
C506 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A a_6725_7308# 0.0334f
C507 a_8523_n7648# D2_2 1.85e-19
C508 a_8643_n1526# D2_2 0.229f
C509 a_1541_n8095# D2_7 1.21e-19
C510 p2_gen_magic_0.xnor_magic_3.OUT a_12174_n3150# 4.14e-19
C511 p2_gen_magic_0.xnor_magic_0.OUT Q1 0.147f
C512 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_5.OUT 4.35e-20
C513 a_20171_6886# Q6 9.64e-20
C514 Q1 Q6 0.427f
C515 7b_counter_0.MDFF_1.tspc2_magic_0.Q 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A 0.00118f
C516 p3_gen_magic_0.xnor_magic_0.OUT D2_2 0.148f
C517 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN CLK 0.0167f
C518 a_4496_4393# a_5515_3947# 0.0292f
C519 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT Q2 0.00596f
C520 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A D2_2 0.0021f
C521 a_15865_6276# D2_1 2.51e-19
C522 a_30365_4922# a_30365_3514# 0.475f
C523 7b_counter_0.MDFF_5.tspc2_magic_0.D CLK 0.00375f
C524 p2_gen_magic_0.xnor_magic_3.OUT Q4 0.0254f
C525 a_26126_3480# a_23560_3728# 6.34e-20
C526 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A a_17405_4932# 3.58e-20
C527 a_19841_4557# Q3 4.89e-20
C528 DFF_magic_0.D a_27234_3319# 7.25e-19
C529 a_8643_n1973# Q5 6.4e-19
C530 a_12931_3363# Q5 0.0664f
C531 a_1409_1059# LD 0.00428f
C532 CLK D2_3 1.61f
C533 a_11191_10149# Q7 0.00975f
C534 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B CLK 3.4e-19
C535 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT D2_6 0.116f
C536 7b_counter_0.MDFF_1.tspc2_magic_0.D Q5 0.0029f
C537 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT VDD 1.18f
C538 7b_counter_0.MDFF_7.tspc2_magic_0.Q Q5 0.148f
C539 p2_gen_magic_0.3_inp_AND_magic_0.VOUT D2_6 0.188f
C540 a_5185_6275# a_5385_6275# 0.297f
C541 7b_counter_0.MDFF_5.LD a_19841_9774# 0.00256f
C542 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT a_12590_n3150# 0.00157f
C543 divide_by_2_0.tg_magic_3.CLK divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT 1.37f
C544 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT D2_3 3.68e-19
C545 DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT CLK 2.41e-19
C546 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A VDD 1.28f
C547 a_11492_n6613# VDD 0.0143f
C548 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT D2_5 0.055f
C549 a_22150_1124# Q3 0.0214f
C550 a_1209_7469# D2_7 0.0192f
C551 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT VDD 1.17f
C552 a_4496_9609# CLK 0.0471f
C553 7b_counter_0.3_inp_AND_magic_0.VOUT Q6 1.06e-20
C554 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_1.OUT 3.33e-19
C555 divide_by_2_1.tg_magic_3.CLK P2 6.12e-20
C556 p3_gen_magic_0.3_inp_AND_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN 0.0147f
C557 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A D2_1 0.00966f
C558 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A a_7215_10149# 3.58e-20
C559 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B Q6 0.0854f
C560 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A 0.00108f
C561 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT Q4 0.00409f
C562 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT D2_1 0.00721f
C563 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A CLK 0.0126f
C564 7b_counter_0.MDFF_1.tspc2_magic_0.D D2_4 0.0179f
C565 a_12174_n7648# D2_5 0.0813f
C566 a_14556_n8142# VDD 0.937f
C567 a_12931_9774# Q7 0.0263f
C568 7b_counter_0.MDFF_7.tspc2_magic_0.Q D2_4 0.361f
C569 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A 0.00108f
C570 a_22991_5815# Q1 0.201f
C571 7b_counter_0.MDFF_3.tspc2_magic_0.D CLK 0.00841f
C572 7b_counter_0.3_inp_AND_magic_0.B a_24185_7877# 0.111f
C573 a_5036_n8095# Q6 0.0818f
C574 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_4.OUT 1.56e-19
C575 a_6725_7308# Q6 0.251f
C576 a_14556_n3644# D2_3 0.0261f
C577 DFF_magic_0.D DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 0.0258f
C578 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_8411_3319# 4.65e-19
C579 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B a_8411_8536# 0.125f
C580 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_14756_n3644# 0.00251f
C581 p3_gen_magic_0.xnor_magic_5.OUT a_5036_n8579# 0.423f
C582 7b_counter_0.DFF_magic_0.tg_magic_0.IN a_27234_4513# 2.82e-20
C583 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A LD 0.409f
C584 a_17405_2092# VDD 0.936f
C585 7b_counter_0.MDFF_4.LD a_19841_4557# 3.96e-19
C586 a_1409_1059# Q3 5.91e-20
C587 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT LD 1.36e-19
C588 a_24059_4877# Q3 0.00209f
C589 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.0215f
C590 a_26038_684# CLK 0.00646f
C591 a_23802_1059# D2_4 0.0308f
C592 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B VDD 1.21f
C593 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.AND2_magic_1.A 2.36e-19
C594 a_17405_8741# D2_3 0.00152f
C595 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 2.64e-19
C596 a_16065_9774# a_15865_8580# 0.00308f
C597 7b_counter_0.MDFF_1.tspc2_magic_0.D a_17405_684# 1.08e-19
C598 a_17405_7309# D2_3 0.0295f
C599 a_12387_1746# D2_6 0.241f
C600 a_1209_4557# a_2749_3524# 7.16e-20
C601 a_16065_1059# D2_3 0.00452f
C602 7b_counter_0.MDFF_5.tspc2_magic_0.Q 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B 4.47e-20
C603 divide_by_2_1.tg_magic_2.IN divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT 0.258f
C604 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.tspc2_magic_0.Q 0.12f
C605 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A 0.00108f
C606 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 0.516f
C607 7b_counter_0.MDFF_7.tspc2_magic_0.Q Q2 2.54e-20
C608 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT DFF_magic_0.tg_magic_1.IN 4.63e-20
C609 divide_by_2_1.tg_magic_1.IN mux_magic_0.OR_magic_0.A 0.00251f
C610 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_17405_4932# 4.22e-19
C611 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_9412_5956# 1.29e-19
C612 a_7215_10149# CLK 0.002f
C613 a_19841_9774# a_21381_10149# 7.98e-19
C614 divide_by_2_1.tg_magic_3.CLK VDD 4.15f
C615 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT D2_7 0.0098f
C616 7b_counter_0.MDFF_7.tspc2_magic_0.D a_24059_4877# 0.278f
C617 a_8643_n5540# D2_5 0.00158f
C618 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A CLK 0.00612f
C619 a_1409_2253# Q7 0.00875f
C620 a_5054_n1042# a_5054_n1526# 0.0335f
C621 a_8643_n1526# p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 1.86e-20
C622 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT 0.165f
C623 7b_counter_0.MDFF_5.LD DFF_magic_0.D 0.465f
C624 a_5054_n5540# VDD 0.497f
C625 OR_magic_1.VOUT divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT 1.31f
C626 p2_gen_magic_0.3_inp_AND_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 0.226f
C627 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT D2_6 0.00148f
C628 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B 0.178f
C629 p3_gen_magic_0.xnor_magic_3.OUT Q5 5.14e-19
C630 divide_by_2_1.tg_magic_3.CLK D2_1 0.00101f
C631 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_0.OUT 1.06e-20
C632 mux_magic_0.AND2_magic_0.A a_32616_n2458# 1.03e-19
C633 a_1209_1059# VDD 0.971f
C634 a_20041_4557# VDD 0.101f
C635 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK p2_gen_magic_0.xnor_magic_1.OUT 0.00316f
C636 a_18891_6886# D2_3 0.0424f
C637 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A VDD 1.24f
C638 a_12931_6276# VDD 0.0542f
C639 a_12931_2253# D2_6 0.172f
C640 p3_gen_magic_0.3_inp_AND_magic_0.C p3_gen_magic_0.xnor_magic_6.OUT 0.029f
C641 a_15865_2253# CLK 3.82e-19
C642 p3_gen_magic_0.xnor_magic_1.B Q7 0.0242f
C643 a_11292_n2115# p2_gen_magic_0.xnor_magic_6.OUT 0.0227f
C644 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A D2_3 0.00135f
C645 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B Q1 0.00733f
C646 a_21381_3524# Q6 2e-20
C647 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN 6.95e-19
C648 a_4496_4393# a_4651_3947# 0.235f
C649 a_12174_n4081# D2_2 0.00121f
C650 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_17405_3524# 1.23e-19
C651 p2_gen_magic_0.3_inp_AND_magic_0.C p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.00145f
C652 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN a_16386_n8142# 3.05e-19
C653 7b_counter_0.MDFF_6.tspc2_magic_0.CLK VDD 2.17f
C654 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A Q4 0.00101f
C655 7b_counter_0.MDFF_5.LD a_23207_5815# 1.42e-19
C656 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A Q1 0.287f
C657 a_24259_4877# a_23560_3728# 0.0141f
C658 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A a_27778_4557# 9.27e-19
C659 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A D2_2 0.0182f
C660 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q3 0.586f
C661 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT 9.92e-19
C662 a_8955_3363# Q1 0.0118f
C663 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B D2_6 0.00268f
C664 p3_gen_magic_0.xnor_magic_3.OUT D2_4 0.216f
C665 7b_counter_0.MDFF_6.tspc2_magic_0.CLK D2_1 0.123f
C666 a_1209_1059# LD 0.00288f
C667 a_12387_1746# D2_2 0.00207f
C668 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT D2_5 0.134f
C669 7b_counter_0.MDFF_4.LD a_15865_6276# 0.0015f
C670 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1559_n6024# 0.0629f
C671 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A a_11191_684# 0.397f
C672 a_9689_1669# Q5 0.0016f
C673 a_13353_n2115# D2_6 0.00532f
C674 a_8713_6842# 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 8.41e-19
C675 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT D2_4 0.163f
C676 a_1409_7469# 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A 0.00103f
C677 a_9059_n6471# VDD 0.0018f
C678 a_23258_1746# Q4 1.26e-19
C679 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_1.OUT 0.00194f
C680 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_19152_5956# 1.29e-19
C681 a_12387_9730# 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A 0.128f
C682 a_11292_n2115# VDD 1.22f
C683 divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT divide_by_2_1.tg_magic_1.IN 4.63e-20
C684 p2_gen_magic_0.xnor_magic_1.OUT Q6 0.0359f
C685 p3_gen_magic_0.xnor_magic_3.OUT Q2 0.289f
C686 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 0.469f
C687 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 0.00576f
C688 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B Q3 0.00777f
C689 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_5515_3947# 5.37e-19
C690 p3_gen_magic_0.3_inp_AND_magic_0.VOUT a_13769_n6613# 0.192f
C691 p3_gen_magic_0.3_inp_AND_magic_0.C D2_3 0.0256f
C692 a_1541_n4081# p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT 8.45e-21
C693 a_8713_6842# VDD 0.757f
C694 a_12174_n8095# VDD 0.181f
C695 a_8713_1625# a_9412_739# 0.0141f
C696 a_15865_2253# a_16065_1059# 0.00308f
C697 a_8939_n7648# D2_5 0.00143f
C698 a_20041_8580# a_20171_6886# 0.00565f
C699 a_11279_1124# 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A 2.4e-20
C700 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 4e-20
C701 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A VDD 1.23f
C702 a_26038_4932# D2_4 0.0163f
C703 7b_counter_0.3_inp_AND_magic_0.B a_23207_5815# 0.0474f
C704 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT CLK 0.413f
C705 a_20041_8580# Q1 0.00357f
C706 a_2749_8740# CLK 0.0161f
C707 p2_gen_magic_0.3_inp_AND_magic_0.VOUT CLK 0.0415f
C708 a_8523_n4081# D2_6 0.00786f
C709 p2_gen_magic_0.xnor_magic_5.OUT a_5036_n4081# 0.414f
C710 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT Q2 0.00334f
C711 7b_counter_0.MDFF_5.LD Q6 0.157f
C712 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT 0.157f
C713 a_9412_5956# D2_6 0.0395f
C714 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_3.QB 0.367f
C715 a_15865_8580# Q1 0.0154f
C716 divide_by_2_0.tg_magic_3.CLK divide_by_2_0.tg_magic_2.IN 0.694f
C717 DFF_magic_0.tg_magic_2.IN CLK 0.00111f
C718 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A Q2 0.0938f
C719 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_14556_n8142# 0.00817f
C720 a_1209_1059# Q3 8.82e-19
C721 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT 0.0205f
C722 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT a_8939_n7648# 6.1e-19
C723 7b_counter_0.MDFF_4.tspc2_magic_0.D Q5 0.00385f
C724 p2_gen_magic_0.xnor_magic_4.OUT Q5 0.147f
C725 a_15865_1059# D2_3 2.51e-19
C726 p3_gen_magic_0.xnor_magic_1.B p3_gen_magic_0.xnor_magic_6.OUT 0.0537f
C727 a_1209_4557# a_2749_4932# 7.98e-19
C728 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1559_n5540# 0.057f
C729 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT Q4 0.00578f
C730 a_16065_2253# a_16065_1059# 0.0206f
C731 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_20171_1669# 0.112f
C732 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A VDD 1.31f
C733 7b_counter_0.MDFF_5.tspc2_magic_0.D a_11191_5901# 1.08e-19
C734 a_12387_6963# 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 1.03e-19
C735 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN VDD 1.18f
C736 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A a_23802_2253# 1.77e-19
C737 a_4496_4393# Q7 0.0576f
C738 a_27778_3363# VDD 0.0124f
C739 p2_gen_magic_0.xnor_magic_0.OUT a_11708_n2115# 0.0247f
C740 a_12387_9730# CLK 6.58e-19
C741 a_1559_n1042# D2_7 0.0172f
C742 a_1209_2253# Q7 0.0429f
C743 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A CLK 0.0666f
C744 a_13353_n6613# p3_gen_magic_0.3_inp_AND_magic_0.VOUT 0.115f
C745 7b_counter_0.MDFF_4.tspc2_magic_0.D D2_4 0.00204f
C746 VDD OUT1 0.345f
C747 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q7 0.0364f
C748 p2_gen_magic_0.xnor_magic_4.OUT D2_4 0.00295f
C749 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.0636f
C750 a_12387_5769# VDD 0.975f
C751 a_27778_4557# a_27778_3363# 0.0206f
C752 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT a_8523_n8579# 0.057f
C753 a_19841_3363# a_20041_3363# 0.296f
C754 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_4235_3947# 6.31e-20
C755 divide_by_2_1.tg_magic_3.CLK mux_magic_0.IN1 0.104f
C756 OR_magic_2.A divide_by_2_1.tg_magic_3.CLK 0.00209f
C757 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.xnor_magic_1.B 3.86e-19
C758 7b_counter_0.DFF_magic_0.D VDD 1.61f
C759 a_12387_9730# a_11279_8697# 7.16e-20
C760 7b_counter_0.3_inp_AND_magic_0.B Q6 0.0615f
C761 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.3_inp_AND_magic_0.A 0.91f
C762 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.3_inp_AND_magic_0.B 0.00468f
C763 divide_by_2_0.tg_magic_3.OUT VDD 1.15f
C764 a_16065_9774# VDD 0.0609f
C765 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A Q1 0.00239f
C766 a_18891_1669# a_19152_1223# 0.299f
C767 7b_counter_0.MDFF_5.LD a_22991_5815# 1.46e-19
C768 7b_counter_0.MDFF_3.tspc2_magic_0.CLK Q2 0.00281f
C769 a_24059_4877# a_23560_3728# 0.299f
C770 a_11292_n2115# Q3 0.0121f
C771 a_19841_3363# Q1 0.0309f
C772 a_21381_10149# Q6 0.0563f
C773 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_19841_4557# 1.1e-19
C774 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_9059_n6471# 6.1e-19
C775 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5470_n1973# 6.1e-19
C776 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT 0.156f
C777 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT CLK 0.313f
C778 divide_by_2_0.tg_magic_3.OUT D2_1 0.0297f
C779 7b_counter_0.MDFF_4.LD a_20041_4557# 1.1e-19
C780 a_22062_684# a_23258_552# 7.98e-19
C781 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A 1.1e-20
C782 a_12174_n8095# a_12174_n8579# 0.0335f
C783 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A a_1209_3363# 0.00184f
C784 p2_gen_magic_0.xnor_magic_4.OUT Q2 0.133f
C785 DFF_magic_0.D DFF_magic_0.tg_magic_1.IN 0.0675f
C786 a_1209_1059# p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT 0.0021f
C787 a_11279_1124# a_11191_684# 0.475f
C788 p2_gen_magic_0.3_inp_AND_magic_0.B D2_3 0.158f
C789 a_8825_1669# Q5 0.00166f
C790 p3_gen_magic_0.xnor_magic_1.OUT Q7 0.153f
C791 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B VDD 1.2f
C792 a_1409_9773# a_1209_8579# 0.00289f
C793 7b_counter_0.DFF_magic_0.D LD 0.0811f
C794 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 7b_counter_0.MDFF_4.LD 3.09e-20
C795 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B a_7215_4932# 4.85e-19
C796 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B Q1 0.0133f
C797 a_8643_n6471# VDD 0.0014f
C798 a_1209_7469# 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A 1.03e-19
C799 7b_counter_0.DFF_magic_0.D a_24003_10051# 0.461f
C800 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT CLK 0.33f
C801 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B Q2 8.23e-19
C802 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 0.00576f
C803 a_9212_5956# a_9412_5956# 0.651f
C804 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B D2_1 3.46e-19
C805 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A VDD 1.28f
C806 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A a_5385_6275# 0.0292f
C807 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT VDD 1.17f
C808 a_1541_n3150# Q6 0.00192f
C809 a_13769_n2115# p2_gen_magic_0.xnor_magic_6.OUT 0.00231f
C810 a_4235_3947# a_5515_3947# 0.00652f
C811 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_4651_3947# 0.00409f
C812 a_13353_n6613# a_13769_n6613# 0.278f
C813 p3_gen_magic_0.3_inp_AND_magic_0.VOUT a_13553_n6613# 1.9e-20
C814 p2_gen_magic_0.AND2_magic_1.A p3_gen_magic_0.3_inp_AND_magic_0.A 3.88e-20
C815 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A D2_1 0.00116f
C816 a_8411_9730# 7b_counter_0.MDFF_5.LD 3.96e-19
C817 a_15865_2253# a_15865_1059# 0.00638f
C818 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT D2_1 0.0833f
C819 a_8523_n8095# VDD 0.181f
C820 a_2749_5900# VDD 1.55f
C821 a_11279_6341# VDD 0.921f
C822 7b_counter_0.3_inp_AND_magic_0.B a_22991_5815# 0.0366f
C823 a_2749_10148# CLK 0.002f
C824 p3_gen_magic_0.xnor_magic_4.OUT D2_5 0.139f
C825 a_1541_n3597# D2_4 5.31e-19
C826 a_13353_n2115# CLK 0.00102f
C827 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B 0.178f
C828 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B LD 6.07e-19
C829 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_11191_684# 0.00215f
C830 p2_gen_magic_0.xnor_magic_6.OUT Q1 0.123f
C831 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B 0.00298f
C832 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A a_12931_3363# 1.77e-19
C833 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B 0.0069f
C834 a_7303_8697# Q6 6.49e-19
C835 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A Q6 0.02f
C836 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_14556_n3644# 0.00818f
C837 a_12387_8536# Q1 0.0151f
C838 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A 2.42e-19
C839 p3_gen_magic_0.xnor_magic_5.OUT a_16386_n8142# 0.0292f
C840 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A LD 0.413f
C841 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT a_8939_n3150# 6.1e-19
C842 a_5385_2253# 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A 5.46e-20
C843 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_12174_n8095# 0.0629f
C844 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A 0.412f
C845 7b_counter_0.DFF_magic_0.D 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 0.244f
C846 p3_gen_magic_0.xnor_magic_3.OUT a_12174_n7648# 4.14e-19
C847 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B Q2 1.74e-19
C848 DFF_magic_0.D 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 0.382f
C849 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A 0.00113f
C850 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A Q1 0.00412f
C851 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_19307_1669# 0.0618f
C852 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A D2_4 0.00176f
C853 a_2749_5900# LD 0.00267f
C854 a_13769_n2115# VDD 0.0181f
C855 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_1209_7469# 1.08e-19
C856 a_1541_n3597# Q2 0.00139f
C857 a_5185_2253# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B 0.125f
C858 p2_gen_magic_0.xnor_magic_0.OUT a_11492_n2115# 0.0655f
C859 a_20041_3363# VDD 0.0856f
C860 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN D2_4 0.00451f
C861 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_26038_4932# 0.173f
C862 7b_counter_0.MDFF_5.LD a_8411_8536# 0.195f
C863 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 1.32f
C864 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT a_8523_n4081# 0.057f
C865 a_13553_n6613# a_13769_n6613# 0.326f
C866 a_20171_6886# VDD 0.075f
C867 7b_counter_0.MDFF_7.tspc2_magic_0.CLK VDD 2.25f
C868 VDD Q1 6.51f
C869 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.00246f
C870 a_1209_3363# D2_5 0.241f
C871 7b_counter_0.MDFF_3.tspc2_magic_0.D a_1209_8579# 7.57e-20
C872 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A 0.412f
C873 p3_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_6.OUT 0.0543f
C874 a_12387_9730# a_11191_10149# 7.98e-19
C875 p3_gen_magic_0.xnor_magic_4.OUT D2_7 0.00894f
C876 7b_counter_0.MDFF_4.LD a_27778_3363# 0.0293f
C877 a_20171_6886# D2_1 4.39e-19
C878 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN a_16186_n8142# 1.97e-20
C879 Q1 D2_1 1.89f
C880 a_5515_9163# VDD 0.0859f
C881 7b_counter_0.MDFF_5.LD a_20041_8580# 0.0279f
C882 mux_magic_0.IN1 OUT1 0.0791f
C883 a_5054_n1973# a_5036_n3597# 6.43e-20
C884 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B a_21381_10149# 0.173f
C885 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A Q3 0.00623f
C886 a_9412_739# D2_6 0.0123f
C887 a_21381_3524# a_19841_3363# 0.00114f
C888 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q3 7.95e-19
C889 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_8643_n6471# 0.102f
C890 a_23793_5904# a_24059_4877# 2.1e-21
C891 a_12174_n3597# a_12174_n4081# 0.0335f
C892 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5054_n1973# 0.102f
C893 7b_counter_0.MDFF_4.tspc2_magic_0.Q 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 0.00507f
C894 7b_counter_0.MDFF_5.LD a_15865_8580# 0.196f
C895 p3_gen_magic_0.AND2_magic_1.A Q4 0.464f
C896 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B Q7 7.61e-19
C897 7b_counter_0.MDFF_0.tspc2_magic_0.Q Q7 0.0796f
C898 7b_counter_0.MDFF_4.LD a_12387_5769# 0.0015f
C899 a_14756_n8142# a_16386_n8142# 0.00333f
C900 OR_magic_1.VOUT divide_by_2_1.tg_magic_0.IN 0.61f
C901 LD Q1 0.00377f
C902 a_1541_n7648# Q7 0.303f
C903 a_12387_9730# a_12931_9774# 0.297f
C904 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT D2_6 0.03f
C905 a_5185_1059# a_5385_1059# 0.297f
C906 7b_counter_0.MDFF_1.tspc2_magic_0.CLK Q5 0.00519f
C907 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT D2_5 0.0482f
C908 a_16065_7470# a_16065_6276# 0.0206f
C909 7b_counter_0.3_inp_AND_magic_0.VOUT VDD 2.57f
C910 a_5515_9163# LD 8.29e-19
C911 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN 0.971f
C912 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 0.228f
C913 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A a_5185_6275# 0.251f
C914 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B a_2749_7308# 0.412f
C915 Q6 D2_5 1.17f
C916 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 0.179f
C917 Q4 Q5 5.12f
C918 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B D2_6 0.00229f
C919 divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.IN 0.29f
C920 DFF_magic_0.D a_27234_552# 2.25e-19
C921 a_13553_n2115# p2_gen_magic_0.xnor_magic_6.OUT 0.0114f
C922 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 5.72e-19
C923 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B VDD 1.2f
C924 a_13353_n6613# a_13553_n6613# 0.519f
C925 a_4235_3947# a_4651_3947# 0.153f
C926 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD 1.1f
C927 a_8411_9730# a_7303_8697# 7.16e-20
C928 a_12931_4557# a_12931_3363# 0.0206f
C929 DFF_magic_0.tg_magic_3.CLK D2_4 2.41e-19
C930 a_5036_n8095# VDD 0.236f
C931 a_1209_3363# D2_7 0.0119f
C932 a_6725_7308# VDD 0.941f
C933 7b_counter_0.DFF_magic_0.tg_magic_3.CLK OR_magic_1.VOUT 1.81e-19
C934 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B CLK 0.0751f
C935 7b_counter_0.MDFF_3.QB 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B 0.00176f
C936 a_5036_n3597# D2_3 4.88e-20
C937 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT D2_1 0.0152f
C938 p2_gen_magic_0.xnor_magic_5.OUT a_16386_n3644# 0.0292f
C939 7b_counter_0.MDFF_1.tspc2_magic_0.CLK D2_4 0.026f
C940 p2_gen_magic_0.3_inp_AND_magic_0.B p2_gen_magic_0.3_inp_AND_magic_0.VOUT 0.0177f
C941 a_8523_n3150# Q1 0.0609f
C942 a_27234_4513# a_26126_3480# 7.16e-20
C943 a_8411_4513# Q6 5.01e-20
C944 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_3 0.978f
C945 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_12174_n3597# 0.0629f
C946 a_9412_739# D2_2 1.68e-20
C947 a_11191_5901# 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 3.58e-20
C948 p3_gen_magic_0.xnor_magic_5.OUT a_14756_n8142# 0.0285f
C949 7b_counter_0.3_inp_AND_magic_0.VOUT LD 0.164f
C950 Q4 D2_4 0.742f
C951 a_2749_2092# 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A 2.07e-19
C952 7b_counter_0.3_inp_AND_magic_0.A Q4 0.0414f
C953 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.3_inp_AND_magic_0.A 0.00121f
C954 7b_counter_0.3_inp_AND_magic_0.VOUT a_24003_10051# 0.187f
C955 7b_counter_0.MDFF_4.tspc2_magic_0.Q a_8411_3319# 0.0276f
C956 a_11292_n6613# p3_gen_magic_0.xnor_magic_6.OUT 0.0227f
C957 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A a_11292_n2115# 2.09e-19
C958 Q1 Q3 0.187f
C959 7b_counter_0.MDFF_7.tspc2_magic_0.CLK Q3 0.0665f
C960 divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT VDD 1.08f
C961 a_26126_1124# D2_4 0.024f
C962 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_17405_684# 0.00215f
C963 p2_gen_magic_0.xnor_magic_3.OUT Q7 0.0898f
C964 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A D2_7 0.00485f
C965 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT Q1 0.0171f
C966 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT D2_2 0.0548f
C967 a_13553_n2115# VDD 0.0169f
C968 a_22150_1124# a_19152_1223# 0.0013f
C969 7b_counter_0.MDFF_6.tspc2_magic_0.Q 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 0.00643f
C970 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A a_2749_2092# 0.0334f
C971 a_5185_2253# a_5385_2253# 0.296f
C972 a_27234_3319# VDD 0.87f
C973 p2_gen_magic_0.xnor_magic_0.OUT a_9059_n1973# 0.0762f
C974 divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT D2_1 0.00175f
C975 7b_counter_0.MDFF_4.tspc2_magic_0.Q a_6725_2092# 0.00134f
C976 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT D2_7 0.0591f
C977 7b_counter_0.MDFF_5.LD a_20041_9774# 0.00109f
C978 a_7303_8697# a_8411_8536# 0.00114f
C979 D2_7 Q6 1f
C980 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 7b_counter_0.MDFF_7.tspc2_magic_0.D 0.423f
C981 Q2 Q4 0.0294f
C982 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK 1.07f
C983 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B D2_2 0.0641f
C984 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A 0.00112f
C985 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A a_12387_3319# 1.03e-19
C986 p2_gen_magic_0.xnor_magic_1.OUT p2_gen_magic_0.xnor_magic_6.OUT 0.0806f
C987 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B VDD 1.2f
C988 a_27778_4557# a_27234_3319# 0.00308f
C989 a_19307_6886# VDD 0.00407f
C990 a_21381_3524# VDD 0.949f
C991 a_2749_8740# a_1209_8579# 0.00114f
C992 a_5036_n7648# p3_gen_magic_0.xnor_magic_5.OUT 0.0924f
C993 p3_gen_magic_0.xnor_magic_1.OUT a_8523_n7648# 4.75e-19
C994 mux_magic_0.AND2_magic_0.A a_32616_n1264# 0.212f
C995 7b_counter_0.MDFF_4.LD a_20041_3363# 0.0279f
C996 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B D2_1 0.00542f
C997 a_19307_6886# D2_1 9.21e-20
C998 a_4651_9163# VDD 0.0501f
C999 7b_counter_0.3_inp_AND_magic_0.VOUT Q3 1.6e-21
C1000 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A p2_gen_magic_0.3_inp_AND_magic_0.C 3.74e-19
C1001 a_24259_4877# a_26126_3480# 1.39e-20
C1002 a_15865_3363# Q1 0.0212f
C1003 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A Q2 0.0282f
C1004 a_11292_n6613# D2_3 0.018f
C1005 a_14756_n3644# a_16386_n3644# 0.00333f
C1006 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B Q3 2.94e-19
C1007 divide_by_2_1.tg_magic_3.CLK divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT 1.37f
C1008 a_1409_8579# D2_7 0.193f
C1009 7b_counter_0.MDFF_5.LD a_12387_8536# 0.195f
C1010 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.26f
C1011 a_4235_3947# Q7 0.0116f
C1012 a_27778_2253# 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 0.00103f
C1013 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT a_5054_n5540# 8.17e-21
C1014 a_1209_4557# a_1209_3363# 0.00638f
C1015 a_8523_n8095# a_8523_n8579# 0.0335f
C1016 a_16186_n8142# a_16386_n8142# 0.299f
C1017 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 0.0847f
C1018 7b_counter_0.MDFF_4.LD Q1 0.192f
C1019 DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD 1.09f
C1020 a_2749_684# a_1209_1059# 7.98e-19
C1021 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT Q6 0.0207f
C1022 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B LD 6.05e-19
C1023 a_8939_n3150# Q5 3.02e-20
C1024 a_8713_1625# D2_6 0.0258f
C1025 a_21381_8741# Q1 0.127f
C1026 p2_gen_magic_0.3_inp_AND_magic_0.B p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT 2.64e-19
C1027 a_16065_9774# a_16065_8580# 0.0206f
C1028 a_17405_5901# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B 4.22e-19
C1029 7b_counter_0.MDFF_3.QB a_5515_9163# 0.167f
C1030 a_11191_684# 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A 3.58e-20
C1031 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_1.tspc2_magic_0.CLK 0.00315f
C1032 p2_gen_magic_0.xnor_magic_1.OUT VDD 6.8f
C1033 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B D2_3 5.05e-19
C1034 a_11708_n2115# p2_gen_magic_0.xnor_magic_6.OUT 0.00656f
C1035 a_4496_4877# a_4651_3947# 0.00164f
C1036 a_5385_2253# VDD 0.109f
C1037 divide_by_2_0.tg_magic_3.CLK divide_by_2_0.tg_magic_3.OUT 0.53f
C1038 p2_gen_magic_0.xnor_magic_1.OUT D2_1 0.529f
C1039 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B 0.00594f
C1040 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT VDD 1.15f
C1041 a_12590_n7648# VDD 0.0018f
C1042 divide_by_2_0.tg_magic_2.IN divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT 0.258f
C1043 a_1559_n1526# a_1957_n3150# 3.01e-19
C1044 p3_gen_magic_0.3_inp_AND_magic_0.A Q4 0.0115f
C1045 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1975_n6471# 0.00157f
C1046 a_16386_n3644# D2_6 7.6e-19
C1047 7b_counter_0.MDFF_5.LD VDD 21.1f
C1048 p2_gen_magic_0.xnor_magic_5.OUT a_14756_n3644# 0.0285f
C1049 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT D2_1 0.0591f
C1050 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A D2_5 0.0946f
C1051 7b_counter_0.MDFF_1.tspc2_magic_0.CLK 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A 0.0037f
C1052 a_1559_n6471# p3_gen_magic_0.xnor_magic_1.B 0.00101f
C1053 p2_gen_magic_0.3_inp_AND_magic_0.B a_13353_n2115# 0.381f
C1054 a_1209_4557# Q6 0.0254f
C1055 p3_gen_magic_0.xnor_magic_5.OUT a_16186_n8142# 0.2f
C1056 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A Q4 4.99e-19
C1057 7b_counter_0.MDFF_5.LD D2_1 0.59f
C1058 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT 0.00385f
C1059 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 7.81e-19
C1060 7b_counter_0.3_inp_AND_magic_0.VOUT a_21381_8741# 4.62e-22
C1061 p2_gen_magic_0.xnor_magic_0.OUT a_8643_n1042# 0.297f
C1062 a_22062_684# p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT 1.69e-19
C1063 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B CLK 0.00238f
C1064 a_5385_2253# LD 0.0279f
C1065 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A Q4 0.00222f
C1066 7b_counter_0.MDFF_7.tspc2_magic_0.D a_27234_3319# 7.57e-20
C1067 a_21381_3524# Q3 0.148f
C1068 a_12387_552# D2_3 4.13e-19
C1069 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A D2_5 0.00285f
C1070 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B p2_gen_magic_0.xnor_magic_3.OUT 3.48e-20
C1071 a_27778_1059# VDD 0.0559f
C1072 p3_gen_magic_0.xnor_magic_0.OUT a_11292_n6613# 0.379f
C1073 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.xnor_magic_3.OUT 0.88f
C1074 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A Q7 0.00332f
C1075 a_11708_n2115# VDD 0.0137f
C1076 a_17405_2092# a_19152_1223# 7.92e-19
C1077 DFF_magic_0.tg_magic_0.IN DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.26f
C1078 a_16065_4557# Q2 0.12f
C1079 7b_counter_0.MDFF_5.LD LD 0.809f
C1080 a_24536_3947# VDD 0.00498f
C1081 p2_gen_magic_0.xnor_magic_0.OUT a_8643_n1973# 0.291f
C1082 7b_counter_0.MDFF_5.LD a_24003_10051# 0.221f
C1083 a_21504_5904# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B 5.98e-19
C1084 mux_magic_0.IN1 divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT 6.54e-20
C1085 OR_magic_1.VOUT divide_by_2_1.tg_magic_3.OUT 0.413f
C1086 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B 0.00112f
C1087 p2_gen_magic_0.xnor_magic_5.OUT D2_6 6.3e-19
C1088 a_5036_n3150# p2_gen_magic_0.xnor_magic_5.OUT 0.0924f
C1089 a_26038_684# DFF_magic_0.tg_magic_3.OUT 8.55e-20
C1090 p2_gen_magic_0.xnor_magic_3.OUT D2_3 0.0812f
C1091 a_17405_5901# VDD 1.55f
C1092 7b_counter_0.3_inp_AND_magic_0.B VDD 0.697f
C1093 a_2749_10148# a_1209_8579# 1.14e-19
C1094 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 0.00594f
C1095 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q4 3.03e-19
C1096 7b_counter_0.MDFF_4.LD a_27234_3319# 0.195f
C1097 a_21381_10149# VDD 1.56f
C1098 p2_gen_magic_0.xnor_magic_1.OUT Q3 0.00147f
C1099 a_24059_4877# a_26126_3480# 0.00212f
C1100 a_12387_3319# Q1 0.0213f
C1101 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B D2_6 0.00814f
C1102 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_27234_1746# 1.08e-19
C1103 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_23560_3728# 0.51f
C1104 a_16186_n3644# a_16386_n3644# 0.299f
C1105 a_8523_n3597# a_8523_n4081# 0.0335f
C1106 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p3_gen_magic_0.3_inp_AND_magic_0.A 1.5e-19
C1107 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 2.82e-19
C1108 a_12174_n7648# Q4 0.304f
C1109 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.P3 3.85e-19
C1110 a_14556_n8142# a_16386_n8142# 0.00107f
C1111 a_16065_8580# Q1 0.0502f
C1112 a_16186_n8142# a_14756_n8142# 3.21e-19
C1113 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT Q5 0.00376f
C1114 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A D2_7 0.00417f
C1115 7b_counter_0.MDFF_3.QB 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B 0.00258f
C1116 7b_counter_0.3_inp_AND_magic_0.B LD 0.01f
C1117 a_9212_739# Q5 0.00772f
C1118 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_21504_5904# 1.75e-21
C1119 7b_counter_0.MDFF_5.LD Q3 5.6e-19
C1120 7b_counter_0.MDFF_5.tspc2_magic_0.Q a_9689_6886# 1.18e-19
C1121 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A Q1 0.00436f
C1122 a_24003_10051# 7b_counter_0.3_inp_AND_magic_0.B 2.42e-20
C1123 p3_gen_magic_0.P3 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 4.95e-19
C1124 7b_counter_0.MDFF_3.QB a_4651_9163# 9.15e-20
C1125 a_1541_n3150# VDD 0.0151f
C1126 a_15865_4557# 7b_counter_0.MDFF_1.tspc2_magic_0.CLK 1.63e-20
C1127 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_5.OUT 0.0158f
C1128 7b_counter_0.MDFF_3.tspc2_magic_0.Q Q2 0.405f
C1129 a_1209_7469# a_2749_7308# 0.00114f
C1130 OR_magic_2.A DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 7.58e-20
C1131 a_11492_n2115# p2_gen_magic_0.xnor_magic_6.OUT 0.00991f
C1132 a_2749_2092# VDD 0.935f
C1133 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 8.78e-21
C1134 p2_gen_magic_0.xnor_magic_5.OUT D2_2 0.0653f
C1135 p3_gen_magic_0.xnor_magic_1.B p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT 0.00129f
C1136 a_1541_n3150# D2_1 0.0573f
C1137 7b_counter_0.MDFF_4.LD DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 0.00268f
C1138 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT D2_4 1.59e-20
C1139 a_27778_1059# Q3 0.146f
C1140 a_12387_1746# a_12931_1059# 0.00308f
C1141 divide_by_2_1.tg_magic_3.CLK divide_by_2_1.tg_magic_2.IN 0.679f
C1142 DFF_magic_0.tg_magic_1.IN P2 0.00193f
C1143 a_9212_739# D2_4 2.51e-20
C1144 a_22150_1124# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A 0.0334f
C1145 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_19841_3363# 0.0276f
C1146 a_7303_8697# VDD 0.941f
C1147 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A VDD 1.23f
C1148 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1559_n6471# 0.0115f
C1149 p2_gen_magic_0.xnor_magic_5.OUT a_16186_n3644# 0.2f
C1150 a_24536_3947# Q3 9.92e-19
C1151 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_3.OUT 2.3e-19
C1152 p3_gen_magic_0.xnor_magic_3.OUT Q6 0.0389f
C1153 divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT VDD 1.08f
C1154 p3_gen_magic_0.xnor_magic_5.OUT a_14556_n8142# 0.0515f
C1155 a_17405_3524# 7b_counter_0.MDFF_1.tspc2_magic_0.CLK 0.121f
C1156 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B D2_2 0.0662f
C1157 7b_counter_0.MDFF_5.tspc2_magic_0.Q Q7 0.198f
C1158 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_12590_n7648# 6.1e-19
C1159 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A a_2749_684# 3.58e-20
C1160 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A Q1 0.00526f
C1161 a_2749_2092# LD 0.00115f
C1162 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_20171_6886# 5.37e-19
C1163 a_23258_1746# a_23258_552# 0.00638f
C1164 7b_counter_0.MDFF_6.tspc2_magic_0.Q Q1 0.458f
C1165 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 0.00709f
C1166 7b_counter_0.MDFF_7.tspc2_magic_0.D a_24536_3947# 0.00451f
C1167 7b_counter_0.3_inp_AND_magic_0.B Q3 0.283f
C1168 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT Q2 7.53e-21
C1169 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT D2_7 0.0299f
C1170 a_5185_2253# D2_5 0.233f
C1171 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT Q6 0.00788f
C1172 a_12931_2253# a_12931_1059# 0.0206f
C1173 OR_magic_2.VOUT a_23352_n5390# 2.68e-19
C1174 p3_gen_magic_0.P3 VDD 2.63f
C1175 DFF_magic_0.tg_magic_3.CLK DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 1.31f
C1176 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_4.LD 0.0352f
C1177 a_1209_9773# D2_7 0.0239f
C1178 a_17405_2092# a_18891_1669# 0.00212f
C1179 a_11492_n2115# VDD 0.0143f
C1180 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A LD 0.00115f
C1181 a_16386_n3644# CLK 2.19e-20
C1182 a_23672_3947# VDD 0.0794f
C1183 p3_gen_magic_0.3_inp_AND_magic_0.B VDD 0.802f
C1184 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A Q6 0.31f
C1185 p3_gen_magic_0.P3 D2_1 0.14f
C1186 7b_counter_0.MDFF_5.LD 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 0.00217f
C1187 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q5 3.37e-19
C1188 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_9212_5956# 4.79e-21
C1189 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT Q4 0.647f
C1190 DFF_magic_0.tg_magic_1.IN VDD 2.02f
C1191 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A 0.00108f
C1192 p3_gen_magic_0.3_inp_AND_magic_0.B D2_1 0.00265f
C1193 p2_gen_magic_0.xnor_magic_6.OUT D2_5 0.0684f
C1194 a_27234_3319# a_27234_1746# 0.00329f
C1195 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A D2_3 0.00203f
C1196 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.AND2_magic_1.A 3.88e-19
C1197 7b_counter_0.MDFF_4.LD a_27778_1059# 0.00428f
C1198 DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK 1.31f
C1199 7b_counter_0.DFF_magic_0.tg_magic_3.CLK P2 0.00249f
C1200 7b_counter_0.MDFF_5.tspc2_magic_0.Q a_8955_9774# 0.12f
C1201 a_1559_n1042# Q4 6.32e-20
C1202 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B a_22062_684# 0.173f
C1203 a_26126_1124# DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 5.8e-22
C1204 divide_by_2_1.tg_magic_0.IN VDD 1.18f
C1205 a_1541_n3150# Q3 0.00207f
C1206 a_24059_4877# a_24259_4877# 0.651f
C1207 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT D2_4 0.758f
C1208 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A a_26126_3480# 0.0334f
C1209 7b_counter_0.MDFF_0.tspc2_magic_0.D a_4651_3947# 0.00451f
C1210 a_19152_5956# a_20041_4557# 3.41e-19
C1211 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_23802_2253# 0.00751f
C1212 a_21381_3524# a_23560_3728# 0.0013f
C1213 a_16186_n3644# a_14756_n3644# 3.21e-19
C1214 a_14556_n3644# a_16386_n3644# 0.00107f
C1215 a_15865_6276# a_16065_6276# 0.297f
C1216 a_23793_5904# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 0.00108f
C1217 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A 0.00108f
C1218 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 0.0037f
C1219 a_12931_8580# Q1 0.00653f
C1220 a_5036_n8095# a_5036_n8579# 0.0335f
C1221 a_14556_n8142# a_14756_n8142# 0.299f
C1222 p2_gen_magic_0.xnor_magic_5.OUT CLK 0.00324f
C1223 7b_counter_0.DFF_magic_0.D a_23985_7877# 1.7e-19
C1224 p2_gen_magic_0.3_inp_AND_magic_0.A p2_gen_magic_0.xnor_magic_6.OUT 0.0397f
C1225 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_19152_5956# 0.347f
C1226 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B Q7 0.00749f
C1227 7b_counter_0.MDFF_5.tspc2_magic_0.Q a_8825_6886# 5.37e-19
C1228 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.3_inp_AND_magic_0.VOUT 1.75e-19
C1229 a_11279_1124# Q1 0.0103f
C1230 7b_counter_0.MDFF_3.tspc2_magic_0.CLK Q6 0.00347f
C1231 a_8411_4513# 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 0.251f
C1232 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT Q5 1.56e-19
C1233 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A 0.178f
C1234 a_12387_6963# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B 0.125f
C1235 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_5.OUT 0.0155f
C1236 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN 6.95e-19
C1237 VDD D2_5 4.74f
C1238 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q2 0.497f
C1239 a_15865_4557# a_16065_4557# 0.297f
C1240 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B Q1 1.46e-19
C1241 a_4235_9163# Q2 1.57e-20
C1242 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 0.00105f
C1243 7b_counter_0.MDFF_1.tspc2_magic_0.Q VDD 1.16f
C1244 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.xnor_magic_4.OUT 0.356f
C1245 a_21381_10149# a_21381_8741# 0.475f
C1246 7b_counter_0.DFF_magic_0.tg_magic_3.CLK VDD 4.27f
C1247 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B CLK 0.00565f
C1248 a_11191_5901# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B 4.22e-19
C1249 p2_gen_magic_0.xnor_magic_4.OUT Q6 0.0101f
C1250 D2_2 D2_6 3.11f
C1251 D2_1 D2_5 1.74f
C1252 p2_gen_magic_0.xnor_magic_6.OUT D2_7 0.00173f
C1253 a_12387_1746# a_12387_552# 0.00638f
C1254 DFF_magic_0.D 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A 2.04e-19
C1255 p2_gen_magic_0.xnor_magic_3.OUT a_1975_n1973# 0.0629f
C1256 7b_counter_0.DFF_magic_0.tg_magic_3.CLK a_27778_4557# 0.022f
C1257 a_16186_n3644# D2_6 9.83e-19
C1258 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A Q7 9.01e-19
C1259 a_8411_4513# VDD 0.984f
C1260 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B Q6 3.81e-19
C1261 a_23672_3947# Q3 9.07e-19
C1262 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT VDD 1.04f
C1263 p2_gen_magic_0.xnor_magic_5.OUT a_14556_n3644# 0.0484f
C1264 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT D2_6 0.0442f
C1265 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_4 3.32e-19
C1266 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B 7b_counter_0.MDFF_0.tspc2_magic_0.Q 4.45e-20
C1267 a_1559_n6024# p3_gen_magic_0.xnor_magic_1.B 5.31e-19
C1268 a_27234_4513# 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A 0.128f
C1269 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_12590_n3150# 6.1e-19
C1270 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_3 6.5e-19
C1271 7b_counter_0.MDFF_4.tspc2_magic_0.CLK Q1 0.0461f
C1272 LD D2_5 0.847f
C1273 DFF_magic_0.tg_magic_1.IN Q3 2.59e-20
C1274 a_6725_684# Q7 8.78e-19
C1275 p2_gen_magic_0.3_inp_AND_magic_0.A VDD 1.33f
C1276 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1541_n3150# 9.19e-19
C1277 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_19307_6886# 1.08e-19
C1278 a_9212_5956# D2_6 0.0554f
C1279 a_20171_1669# D2_3 4.39e-19
C1280 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.OUT 0.00933f
C1281 7b_counter_0.MDFF_6.tspc2_magic_0.D 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 2.05e-19
C1282 7b_counter_0.MDFF_5.LD a_16065_8580# 0.0292f
C1283 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A D2_6 0.00297f
C1284 a_9059_n1973# VDD 0.0018f
C1285 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT CLK 0.0124f
C1286 7b_counter_0.MDFF_3.QB a_7303_8697# 0.00363f
C1287 a_16065_3363# VDD 0.0191f
C1288 VDD D2_7 5.81f
C1289 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN 0.0617f
C1290 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A D2_6 0.0603f
C1291 a_1559_n6471# a_1541_n7648# 0.0128f
C1292 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B Q6 0.0522f
C1293 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A a_12931_7470# 1.77e-19
C1294 a_27234_1746# a_27778_1059# 0.00308f
C1295 7b_counter_0.MDFF_0.tspc2_magic_0.D Q7 0.0106f
C1296 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8523_n3597# 1.63e-19
C1297 a_5470_n6471# D2_4 0.00551f
C1298 a_11492_n6613# a_11708_n6613# 0.326f
C1299 D2_7 D2_1 0.661f
C1300 divide_by_2_0.tg_magic_0.IN VDD 1.18f
C1301 OR_magic_2.A p3_gen_magic_0.P3 0.218f
C1302 a_8523_n3150# D2_5 6.39e-20
C1303 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A Q2 7.6e-19
C1304 a_20041_3363# a_19152_1223# 5.39e-19
C1305 a_23560_3728# a_24536_3947# 0.235f
C1306 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A D2_4 5.7e-19
C1307 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A CLK 7.36e-19
C1308 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A CLK 0.0294f
C1309 p3_gen_magic_0.3_inp_AND_magic_0.B p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT 2.64e-19
C1310 7b_counter_0.MDFF_1.tspc2_magic_0.D 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 8.78e-21
C1311 7b_counter_0.MDFF_4.LD a_23672_3947# 8.29e-19
C1312 OR_magic_2.A DFF_magic_0.tg_magic_1.IN 0.00104f
C1313 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 1.31f
C1314 a_12174_n8579# D2_5 0.00786f
C1315 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.B 4e-19
C1316 Q3 D2_5 0.044f
C1317 Q7 Q5 0.946f
C1318 a_27234_552# VDD 0.971f
C1319 a_1559_n5540# D2_4 0.00786f
C1320 LD D2_7 1.05f
C1321 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN Q4 0.00811f
C1322 7b_counter_0.MDFF_4.LD DFF_magic_0.tg_magic_1.IN 8.9e-20
C1323 a_2749_3524# a_4651_3947# 2.12e-20
C1324 a_19152_1223# Q1 0.0395f
C1325 a_12387_6963# D2_6 3.28e-20
C1326 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_5 0.0258f
C1327 a_8411_3319# Q1 0.0202f
C1328 a_5036_n3597# a_5036_n4081# 0.0335f
C1329 a_14556_n3644# a_14756_n3644# 0.299f
C1330 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5054_n1526# 0.0628f
C1331 a_5470_n6471# Q2 2.48e-20
C1332 a_8643_n1526# p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT 2.26e-20
C1333 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A a_17405_8741# 2.07e-19
C1334 a_21504_5904# Q1 0.0483f
C1335 a_7215_4932# Q7 0.0197f
C1336 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT VDD 1.07f
C1337 CLK D2_6 0.66f
C1338 DFF_magic_0.D DFF_magic_0.tg_magic_3.CLK 0.539f
C1339 a_14556_n8142# a_16186_n8142# 3.4e-19
C1340 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A Q7 0.0173f
C1341 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_0.OUT 3.68e-20
C1342 a_9689_6886# Q2 0.0301f
C1343 p3_gen_magic_0.xnor_magic_4.OUT Q4 0.00134f
C1344 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 1.19e-19
C1345 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_6.tspc2_magic_0.Q 0.125f
C1346 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_1 6.11e-19
C1347 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A D2_2 0.00179f
C1348 a_6725_2092# Q1 0.0171f
C1349 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A a_2749_5900# 0.397f
C1350 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q7 0.495f
C1351 a_11292_n2115# p2_gen_magic_0.3_inp_AND_magic_0.C 2.07e-19
C1352 p2_gen_magic_0.xnor_magic_3.OUT a_13353_n2115# 0.00201f
C1353 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT D2_6 0.0558f
C1354 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.153f
C1355 a_5385_7469# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A 1.77e-19
C1356 DFF_magic_0.tg_magic_0.IN CLK 0.61f
C1357 a_5470_n1973# Q2 2.48e-20
C1358 Q7 D2_4 0.0373f
C1359 a_1559_n5540# Q2 0.0143f
C1360 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A D2_2 0.0881f
C1361 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 4.02e-20
C1362 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT 0.00385f
C1363 divide_by_2_1.tg_magic_3.OUT P2 3.4e-19
C1364 p2_gen_magic_0.3_inp_AND_magic_0.A Q3 0.00409f
C1365 a_11279_8697# D2_6 0.0127f
C1366 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.3_inp_AND_magic_0.C 7.01e-19
C1367 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A 7b_counter_0.MDFF_5.tspc2_magic_0.Q 0.00118f
C1368 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT D2_5 0.974f
C1369 p2_gen_magic_0.xnor_magic_3.OUT a_1559_n1973# 0.0924f
C1370 a_11191_684# a_11292_n2115# 8.67e-20
C1371 a_1209_4557# VDD 0.975f
C1372 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1559_n6024# 0.0834f
C1373 7b_counter_0.DFF_magic_0.tg_magic_3.CLK OR_magic_2.A 1.13e-19
C1374 a_19841_4557# a_20041_4557# 0.297f
C1375 D2_7 Q3 1.15f
C1376 Q2 Q7 1.94f
C1377 7b_counter_0.3_inp_AND_magic_0.VOUT a_23985_7877# 0.117f
C1378 a_23207_5815# Q4 0.0204f
C1379 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_1.tspc2_magic_0.Q 0.114f
C1380 a_17405_4932# Q1 0.00215f
C1381 p3_gen_magic_0.xnor_magic_6.OUT p3_gen_magic_0.AND2_magic_1.A 0.238f
C1382 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK Q4 0.274f
C1383 7b_counter_0.MDFF_4.LD 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 0.0408f
C1384 a_12387_6963# D2_2 0.248f
C1385 a_8643_n1042# VDD 0.376f
C1386 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A a_1409_4557# 0.0292f
C1387 a_5185_6275# a_4496_4393# 2.33e-20
C1388 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_1.OUT 0.00181f
C1389 a_5054_n6471# Q5 0.579f
C1390 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 1.84e-19
C1391 CLK D2_2 0.54f
C1392 a_15865_9774# CLK 0.223f
C1393 7b_counter_0.MDFF_6.tspc2_magic_0.Q 7b_counter_0.3_inp_AND_magic_0.B 0.00247f
C1394 a_19307_1669# D2_3 0.00746f
C1395 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B a_6725_2092# 0.409f
C1396 a_1541_n4081# p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT 7.56e-21
C1397 divide_by_2_1.tg_magic_3.OUT VDD 1.15f
C1398 7b_counter_0.MDFF_5.LD a_12931_8580# 0.0293f
C1399 7b_counter_0.MDFF_4.LD a_8411_4513# 3.96e-19
C1400 a_8643_n1973# VDD 0.0014f
C1401 a_27234_552# Q3 0.25f
C1402 a_16186_n3644# CLK 0.00253f
C1403 a_1209_4557# LD 0.0019f
C1404 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A D2_4 0.0157f
C1405 a_5054_n1973# Q5 0.0456f
C1406 a_12931_3363# VDD 0.0124f
C1407 p3_gen_magic_0.xnor_magic_6.OUT Q5 0.146f
C1408 a_6725_684# D2_3 2.92e-20
C1409 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT CLK 0.00519f
C1410 p2_gen_magic_0.3_inp_AND_magic_0.B a_16386_n3644# 6.81e-19
C1411 divide_by_2_1.tg_magic_3.OUT D2_1 9.28e-21
C1412 a_1541_n8095# Q7 0.0805f
C1413 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 0.00754f
C1414 a_15865_7470# a_17405_7309# 0.00114f
C1415 7b_counter_0.MDFF_1.tspc2_magic_0.D VDD 1.38f
C1416 a_2749_3524# Q7 0.0209f
C1417 a_5054_n6471# D2_4 0.00867f
C1418 7b_counter_0.MDFF_7.tspc2_magic_0.Q VDD 1.21f
C1419 a_11279_8697# D2_2 0.0364f
C1420 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 0.0041f
C1421 a_5452_n3150# D2_5 0.00278f
C1422 a_15865_3363# a_16065_3363# 0.298f
C1423 divide_by_2_0.tg_magic_3.CLK divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT 0.0636f
C1424 p2_gen_magic_0.xnor_magic_0.OUT a_12174_n3150# 0.00199f
C1425 a_23258_552# D2_4 0.031f
C1426 a_9212_5956# CLK 0.00355f
C1427 a_23560_3728# a_23672_3947# 0.0292f
C1428 a_19152_739# CLK 4.53e-22
C1429 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT 0.0214f
C1430 a_8955_3363# a_8825_1669# 0.00565f
C1431 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B Q5 0.00237f
C1432 p2_gen_magic_0.xnor_magic_0.OUT Q4 0.0278f
C1433 7b_counter_0.MDFF_4.LD a_16065_3363# 0.0293f
C1434 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN 0.848f
C1435 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A CLK 0.00612f
C1436 a_23802_1059# VDD 0.0979f
C1437 Q6 Q4 0.266f
C1438 a_1209_1059# a_1409_1059# 0.297f
C1439 7b_counter_0.MDFF_3.QB D2_7 0.299f
C1440 p3_gen_magic_0.P3 divide_by_2_0.tg_magic_3.CLK 5.98e-20
C1441 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_9689_6886# 0.0618f
C1442 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A a_24059_4877# 3.22e-21
C1443 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A CLK 0.00246f
C1444 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_11191_5901# 0.173f
C1445 a_18891_1669# Q1 0.00561f
C1446 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT Q4 0.00132f
C1447 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_7 0.151f
C1448 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_26126_3480# 0.019f
C1449 a_14556_n3644# a_16186_n3644# 3.4e-19
C1450 a_5054_n6471# Q2 0.302f
C1451 a_19152_5956# Q1 1.39e-19
C1452 a_15865_9774# a_17405_8741# 7.16e-20
C1453 a_1209_9773# 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 1.37e-19
C1454 a_8825_6886# Q2 0.00202f
C1455 a_8713_6842# 7b_counter_0.MDFF_4.tspc2_magic_0.Q 0.00119f
C1456 p2_gen_magic_0.3_inp_AND_magic_0.B p2_gen_magic_0.xnor_magic_5.OUT 0.049f
C1457 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_15865_6276# 1.37e-19
C1458 Q5 D2_3 0.625f
C1459 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A a_11279_8697# 0.0334f
C1460 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B D2_4 0.014f
C1461 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT a_8523_n8579# 0.0846f
C1462 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B Q5 0.00222f
C1463 7b_counter_0.MDFF_4.LD a_27234_552# 0.00396f
C1464 a_5054_n1973# Q2 0.302f
C1465 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A a_11279_8697# 2.07e-19
C1466 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_17405_5901# 0.173f
C1467 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A a_21381_4932# 3.58e-20
C1468 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_0.tspc2_magic_0.D 8.78e-21
C1469 a_1409_9773# Q2 6.99e-19
C1470 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A Q7 0.00247f
C1471 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT VDD 1.09f
C1472 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A Q1 0.00239f
C1473 a_12387_6963# CLK 0.0316f
C1474 a_8643_n1973# a_8523_n3150# 0.186f
C1475 p3_gen_magic_0.3_inp_AND_magic_0.C D2_6 0.06f
C1476 a_11191_10149# D2_6 0.00522f
C1477 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.3_inp_AND_magic_0.VOUT 4.16e-20
C1478 a_5452_n3150# D2_7 0.00371f
C1479 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_9059_n6471# 0.00157f
C1480 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5470_n1973# 0.00157f
C1481 a_7303_3480# a_4496_4393# 0.00153f
C1482 7b_counter_0.MDFF_5.tspc2_magic_0.CLK Q7 0.00459f
C1483 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK 1.34f
C1484 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT D2_1 0.00732f
C1485 p2_gen_magic_0.xnor_magic_3.OUT a_5054_n1526# 1.65e-19
C1486 D2_3 D2_4 1.59f
C1487 p3_gen_magic_0.xnor_magic_3.OUT VDD 2.84f
C1488 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B D2_4 0.0139f
C1489 p2_gen_magic_0.xnor_magic_6.OUT p2_gen_magic_0.AND2_magic_1.A 0.241f
C1490 p3_gen_magic_0.3_inp_AND_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT 0.702f
C1491 a_22991_5815# Q4 0.00728f
C1492 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 7b_counter_0.DFF_magic_0.tg_magic_0.IN 0.164f
C1493 a_27234_4513# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 1.37e-19
C1494 p3_gen_magic_0.xnor_magic_5.OUT a_5036_n8095# 0.368f
C1495 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A a_21381_4932# 0.397f
C1496 7b_counter_0.MDFF_5.tspc2_magic_0.D Q2 0.103f
C1497 p3_gen_magic_0.xnor_magic_3.OUT D2_1 1.59f
C1498 7b_counter_0.MDFF_1.tspc2_magic_0.D Q3 2.79e-19
C1499 divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT VDD 1.08f
C1500 7b_counter_0.MDFF_7.tspc2_magic_0.Q Q3 0.479f
C1501 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.AND2_magic_1.A 3.88e-19
C1502 a_8643_n6024# Q5 6.51e-20
C1503 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 5.4e-19
C1504 a_11279_8697# CLK 0.0159f
C1505 p2_gen_magic_0.3_inp_AND_magic_0.C a_13769_n2115# 0.0441f
C1506 a_2749_2092# a_2749_684# 0.475f
C1507 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A a_1409_3363# 1.77e-19
C1508 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT VDD 1.03f
C1509 a_17405_7309# a_19152_6440# 6.34e-20
C1510 a_15865_1059# D2_6 4.11e-19
C1511 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B a_17405_684# 0.173f
C1512 divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT D2_1 0.00124f
C1513 Q2 D2_3 0.0512f
C1514 7b_counter_0.MDFF_5.LD a_23985_7877# 8.82e-20
C1515 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A VDD 1.31f
C1516 a_32816_n1264# VDD 0.0559f
C1517 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT D2_1 1.1f
C1518 a_8523_n7648# Q5 0.319f
C1519 a_14556_n3644# CLK 0.00444f
C1520 a_8643_n1526# Q5 6.51e-20
C1521 p2_gen_magic_0.3_inp_AND_magic_0.B a_14756_n3644# 0.00227f
C1522 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A a_17405_10149# 0.397f
C1523 7b_counter_0.3_inp_AND_magic_0.C CLK 0.0743f
C1524 a_1559_n6024# a_1541_n7648# 0.00121f
C1525 p3_gen_magic_0.xnor_magic_0.OUT Q5 4.41e-20
C1526 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A D2_1 6.27e-20
C1527 a_32816_n1264# D2_1 0.00329f
C1528 a_2749_7308# Q6 0.00926f
C1529 a_9689_1669# VDD 0.00407f
C1530 a_2749_4932# Q7 0.00254f
C1531 a_26038_4932# VDD 1.56f
C1532 7b_counter_0.MDFF_5.LD a_16065_7470# 0.0293f
C1533 a_4496_9609# Q2 0.00123f
C1534 p2_gen_magic_0.AND2_magic_1.A VDD 1.4f
C1535 a_18891_6886# a_19152_6440# 0.299f
C1536 a_11191_5901# D2_6 0.00491f
C1537 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5054_n1042# 0.0846f
C1538 p3_gen_magic_0.3_inp_AND_magic_0.A p3_gen_magic_0.xnor_magic_6.OUT 0.0397f
C1539 p2_gen_magic_0.xnor_magic_0.OUT a_8939_n3150# 1.73e-19
C1540 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.xnor_magic_6.OUT 0.0308f
C1541 a_23672_3947# a_23802_2253# 0.00565f
C1542 a_26126_3480# a_27234_3319# 0.00114f
C1543 7b_counter_0.MDFF_3.tspc2_magic_0.Q 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A 0.00118f
C1544 a_8955_8580# a_8825_6886# 0.00565f
C1545 a_8955_4557# D2_6 0.00606f
C1546 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A Q2 0.0972f
C1547 p2_gen_magic_0.AND2_magic_1.A D2_1 2.23e-19
C1548 7b_counter_0.MDFF_4.LD a_12931_3363# 0.0292f
C1549 a_5185_6275# 7b_counter_0.MDFF_0.tspc2_magic_0.Q 1.11e-19
C1550 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A LD 0.412f
C1551 7b_counter_0.MDFF_3.tspc2_magic_0.D Q2 0.0011f
C1552 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 2.63e-19
C1553 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_8825_6886# 0.112f
C1554 a_11191_684# Q1 0.00119f
C1555 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_1.tspc2_magic_0.D 0.00121f
C1556 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B a_12387_8536# 0.125f
C1557 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_7.tspc2_magic_0.Q 0.111f
C1558 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_24259_4877# 0.35f
C1559 a_19307_6886# a_19152_5956# 0.00164f
C1560 7b_counter_0.3_inp_AND_magic_0.B a_21504_5904# 0.898f
C1561 p3_gen_magic_0.xnor_magic_1.B D2_6 0.0483f
C1562 7b_counter_0.3_inp_AND_magic_0.B a_23985_7877# 0.322f
C1563 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT a_8523_n4081# 0.0846f
C1564 a_27234_1746# a_27234_552# 0.00638f
C1565 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_20041_4557# 0.00103f
C1566 7b_counter_0.MDFF_3.tspc2_magic_0.CLK VDD 2.44f
C1567 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A Q4 0.00146f
C1568 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A a_11191_10149# 0.397f
C1569 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B a_4235_3947# 7.16e-19
C1570 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A CLK 0.00225f
C1571 a_15865_2253# D2_4 0.00225f
C1572 p3_gen_magic_0.xnor_magic_3.OUT Q3 0.145f
C1573 divide_by_2_0.tg_magic_3.CLK divide_by_2_0.tg_magic_0.IN 0.164f
C1574 7b_counter_0.MDFF_4.LD a_23802_1059# 1.1e-19
C1575 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 0.00956f
C1576 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A D2_3 0.188f
C1577 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B CLK 0.00118f
C1578 a_5185_7469# a_6725_7308# 0.00114f
C1579 7b_counter_0.MDFF_3.tspc2_magic_0.CLK D2_1 0.0423f
C1580 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.00246f
C1581 a_19841_8580# Q7 0.0011f
C1582 7b_counter_0.MDFF_4.tspc2_magic_0.D VDD 1.38f
C1583 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1541_n7648# 9.19e-19
C1584 p2_gen_magic_0.xnor_magic_4.OUT VDD 1.5f
C1585 DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT DFF_magic_0.tg_magic_2.OUT 0.156f
C1586 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A a_2749_3524# 2.4e-20
C1587 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A Q2 0.00278f
C1588 divide_by_2_1.tg_magic_0.IN divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT 4.89e-20
C1589 p3_gen_magic_0.3_inp_AND_magic_0.A D2_3 0.02f
C1590 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A Q4 0.0022f
C1591 p2_gen_magic_0.xnor_magic_1.OUT a_13353_n6613# 1.57e-19
C1592 a_11191_5901# D2_2 0.0429f
C1593 a_17405_8741# a_17405_7309# 0.00112f
C1594 a_27234_4513# a_27234_3319# 0.00638f
C1595 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8643_n6471# 0.00638f
C1596 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5054_n1973# 0.00941f
C1597 a_15865_2253# a_17405_684# 1.14e-19
C1598 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B VDD 1.2f
C1599 a_22062_684# 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 3.58e-20
C1600 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN CLK 0.595f
C1601 p2_gen_magic_0.xnor_magic_3.OUT a_1559_n1526# 0.368f
C1602 a_1409_3363# D2_5 0.171f
C1603 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A a_16065_3363# 0.00103f
C1604 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A D2_3 0.00213f
C1605 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 7b_counter_0.MDFF_5.tspc2_magic_0.D 0.414f
C1606 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A a_1409_1059# 0.0292f
C1607 7b_counter_0.MDFF_3.tspc2_magic_0.CLK LD 0.087f
C1608 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A a_12931_9774# 9.27e-19
C1609 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A 0.178f
C1610 p2_gen_magic_0.xnor_magic_5.OUT a_5036_n3597# 0.368f
C1611 a_23258_1746# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B 0.125f
C1612 a_8523_n3597# D2_6 0.231f
C1613 a_5036_n8579# D2_7 0.0381f
C1614 7b_counter_0.MDFF_3.tspc2_magic_0.Q Q6 0.155f
C1615 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_5385_1059# 0.12f
C1616 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B D2_1 3.46e-19
C1617 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT Q5 4.95e-19
C1618 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.xnor_magic_5.OUT 5.78e-19
C1619 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8523_n8095# 1.63e-19
C1620 p3_gen_magic_0.xnor_magic_6.OUT a_12174_n7648# 0.144f
C1621 a_19841_4557# Q1 0.0143f
C1622 a_5036_n7648# a_5036_n8095# 0.0142f
C1623 a_2749_684# D2_5 0.00292f
C1624 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_5 0.0913f
C1625 p2_gen_magic_0.3_inp_AND_magic_0.C a_13553_n2115# 0.00138f
C1626 a_11191_10149# CLK 0.002f
C1627 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A a_12931_6276# 9.27e-19
C1628 p3_gen_magic_0.3_inp_AND_magic_0.C CLK 0.687f
C1629 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 0.193f
C1630 a_17405_7309# a_18891_6886# 0.00212f
C1631 a_32816_n2458# VDD 0.0124f
C1632 a_1559_n1042# Q7 0.0489f
C1633 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_5054_n1042# 6.8e-20
C1634 7b_counter_0.MDFF_4.tspc2_magic_0.Q Q1 0.153f
C1635 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A a_4496_4393# 2.58e-19
C1636 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B LD 6.07e-19
C1637 a_34156_n2297# VDD 0.926f
C1638 a_32816_n2458# D2_1 0.0324f
C1639 7b_counter_0.MDFF_7.tspc2_magic_0.D a_26038_4932# 1.08e-19
C1640 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT D2_4 0.0143f
C1641 a_8643_n6471# p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 0.0016f
C1642 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B VDD 1.21f
C1643 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_7303_3480# 0.00134f
C1644 p2_gen_magic_0.3_inp_AND_magic_0.B a_16186_n3644# 0.0437f
C1645 p2_gen_magic_0.3_inp_AND_magic_0.VOUT D2_4 0.00249f
C1646 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.0032f
C1647 a_8825_1669# VDD 0.075f
C1648 a_11191_10149# a_11279_8697# 0.475f
C1649 a_1975_n6471# D2_4 0.00157f
C1650 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT Q6 0.593f
C1651 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT D2_3 0.0531f
C1652 p3_gen_magic_0.3_inp_AND_magic_0.B p3_gen_magic_0.3_inp_AND_magic_0.VOUT 0.0231f
C1653 7b_counter_0.MDFF_5.LD a_12931_7470# 0.0248f
C1654 a_1541_n3597# VDD 0.181f
C1655 mux_magic_0.IN1 a_32816_n1264# 0.12f
C1656 a_12931_9774# CLK 0.00494f
C1657 a_12387_3319# a_12931_3363# 0.298f
C1658 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT a_8523_n8095# 0.0834f
C1659 a_26126_3480# a_24536_3947# 2.12e-20
C1660 a_15865_1059# CLK 1.92e-19
C1661 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.3_inp_AND_magic_0.A 0.00121f
C1662 a_5515_3947# Q6 0.00144f
C1663 a_1409_3363# D2_7 0.00916f
C1664 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A a_27778_3363# 1.77e-19
C1665 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT 0.00142f
C1666 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT 0.00888f
C1667 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 1.41f
C1668 a_1541_n3597# D2_1 0.231f
C1669 a_12387_1746# Q5 3.88e-19
C1670 a_8523_n3597# D2_2 3.13e-19
C1671 a_1975_n1973# D2_4 0.00157f
C1672 7b_counter_0.MDFF_7.tspc2_magic_0.Q a_23560_3728# 0.013f
C1673 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q1 0.615f
C1674 7b_counter_0.MDFF_4.tspc2_magic_0.D Q3 4.06e-19
C1675 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_19841_3363# 4.65e-19
C1676 p2_gen_magic_0.xnor_magic_4.OUT Q3 0.00283f
C1677 a_12387_6963# a_11191_5901# 1.14e-19
C1678 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_24059_4877# 0.654f
C1679 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A Q4 6.96e-19
C1680 p2_gen_magic_0.xnor_magic_5.OUT a_11292_n6613# 7.66e-21
C1681 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_7 1.14f
C1682 a_1975_n6471# Q2 7.44e-19
C1683 a_12387_5769# a_12931_6276# 0.297f
C1684 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A VDD 1.23f
C1685 7b_counter_0.MDFF_4.tspc2_magic_0.Q 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B 4.45e-20
C1686 a_19841_3363# Q4 2.73e-20
C1687 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A a_8955_8580# 1.77e-19
C1688 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN VDD 2.02f
C1689 DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.153f
C1690 p2_gen_magic_0.3_inp_AND_magic_0.C p2_gen_magic_0.xnor_magic_1.OUT 0.0215f
C1691 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B a_4496_4877# 1.29e-19
C1692 a_15865_2253# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A 0.00184f
C1693 a_12387_1746# D2_4 0.00225f
C1694 p2_gen_magic_0.xnor_magic_3.OUT a_5054_n1042# 0.128f
C1695 divide_by_2_0.tg_magic_1.IN VDD 2.02f
C1696 a_1409_2253# CLK 0.12f
C1697 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_6.OUT 0.0173f
C1698 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A 0.00619f
C1699 a_12387_9730# Q2 9.61e-19
C1700 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A a_2749_4932# 3.58e-20
C1701 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A VDD 1.24f
C1702 p3_gen_magic_0.3_inp_AND_magic_0.B a_13769_n6613# 0.109f
C1703 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A Q2 0.0507f
C1704 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT Q1 2.49e-19
C1705 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK Q4 0.0114f
C1706 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A a_4235_9163# 3.22e-21
C1707 p3_gen_magic_0.xnor_magic_1.OUT D2_6 2.34f
C1708 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT D2_4 6.16e-19
C1709 a_1975_n6471# a_1541_n8095# 3.04e-19
C1710 a_19841_9774# Q7 0.0527f
C1711 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B Q5 4.93e-19
C1712 a_15865_1059# a_16065_1059# 0.297f
C1713 DFF_magic_0.tg_magic_3.CLK P2 0.655f
C1714 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 0.00312f
C1715 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 0.00322f
C1716 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A D2_1 0.00213f
C1717 7b_counter_0.MDFF_3.QB 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 0.0751f
C1718 p3_gen_magic_0.xnor_magic_4.OUT a_5470_n6471# 0.0761f
C1719 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A a_1209_1059# 0.251f
C1720 p2_gen_magic_0.3_inp_AND_magic_0.B CLK 1.01e-19
C1721 7b_counter_0.DFF_magic_0.tg_magic_3.CLK a_30365_4922# 4.31e-19
C1722 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_19152_1223# 0.0129f
C1723 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q6 0.0158f
C1724 a_16065_2253# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A 1.77e-19
C1725 a_19841_8580# D2_3 0.00302f
C1726 p2_gen_magic_0.xnor_magic_6.OUT a_12174_n3150# 0.144f
C1727 a_5036_n3150# a_5036_n3597# 0.0142f
C1728 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_5185_1059# 0.223f
C1729 a_1541_n8579# D2_7 0.0628f
C1730 p3_gen_magic_0.3_inp_AND_magic_0.B a_16386_n8142# 6.81e-19
C1731 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B a_7215_4932# 0.173f
C1732 a_17405_3524# D2_3 0.00646f
C1733 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5036_n3150# 5.22e-19
C1734 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD 1.08f
C1735 a_13353_n2115# Q5 7.55e-20
C1736 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A 0.178f
C1737 a_19841_4557# a_21381_3524# 7.16e-20
C1738 p3_gen_magic_0.xnor_magic_6.OUT a_8939_n7648# 0.0629f
C1739 Q4 P2 0.315f
C1740 p2_gen_magic_0.xnor_magic_6.OUT Q4 0.386f
C1741 a_1559_n6471# Q5 0.582f
C1742 p3_gen_magic_0.xnor_magic_0.OUT a_12174_n7648# 0.00199f
C1743 a_1541_n3597# Q3 6.69e-21
C1744 DFF_magic_0.D 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 0.0111f
C1745 a_8411_4513# a_8411_3319# 0.00638f
C1746 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A a_12387_5769# 0.128f
C1747 a_12931_1059# D2_6 0.00452f
C1748 divide_by_2_0.tg_magic_3.CLK divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT 1.31f
C1749 7b_counter_0.MDFF_5.LD a_16065_6276# 0.00329f
C1750 a_8643_n5540# a_8643_n6024# 0.0335f
C1751 a_34156_n889# VDD 1.55f
C1752 a_5385_7469# VDD 0.109f
C1753 a_13353_n2115# D2_4 0.00384f
C1754 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A p2_gen_magic_0.3_inp_AND_magic_0.VOUT 1e-19
C1755 p2_gen_magic_0.3_inp_AND_magic_0.B a_14556_n3644# 0.127f
C1756 a_17405_2092# Q1 0.0106f
C1757 a_21381_3524# a_22150_1124# 7.9e-19
C1758 mux_magic_0.IN1 a_32816_n2458# 0.002f
C1759 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B 9.4e-20
C1760 a_8523_n4081# Q5 2.81e-19
C1761 DFF_magic_0.tg_magic_3.CLK VDD 4.17f
C1762 a_1559_n6471# p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT 0.00274f
C1763 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B Q1 0.075f
C1764 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT a_8523_n3597# 0.0834f
C1765 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A Q3 0.0143f
C1766 a_8643_n6471# a_9059_n6471# 5.82e-19
C1767 p3_gen_magic_0.3_inp_AND_magic_0.B a_13353_n6613# 0.381f
C1768 a_1559_n6471# D2_4 0.0571f
C1769 7b_counter_0.MDFF_1.tspc2_magic_0.CLK VDD 2.18f
C1770 p3_gen_magic_0.3_inp_AND_magic_0.B p3_gen_magic_0.xnor_magic_5.OUT 0.049f
C1771 a_12174_n3150# VDD 0.0014f
C1772 a_1209_8579# CLK 0.0201f
C1773 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.141f
C1774 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN Q3 0.0653f
C1775 a_24259_4877# a_24536_3947# 0.00164f
C1776 a_22062_684# CLK 0.0278f
C1777 a_4651_3947# Q6 6.8e-19
C1778 divide_by_2_0.tg_magic_3.CLK divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT 1.84e-19
C1779 p3_gen_magic_0.xnor_magic_0.OUT a_8643_n5540# 0.297f
C1780 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_2.OUT 1.09f
C1781 VDD Q4 13f
C1782 a_9059_n6471# a_8523_n8095# 1.25e-19
C1783 a_1559_n1973# D2_4 0.101f
C1784 7b_counter_0.MDFF_7.tspc2_magic_0.Q a_23802_2253# 0.017f
C1785 a_5054_n5540# Q1 5.54e-20
C1786 a_5385_7469# LD 0.0279f
C1787 D2_1 Q4 0.135f
C1788 7b_counter_0.MDFF_4.LD a_8825_1669# 8.29e-19
C1789 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A Q6 3.37e-19
C1790 a_5185_1059# p2_gen_magic_0.xnor_magic_3.OUT 1.7e-19
C1791 a_20041_4557# Q1 0.00191f
C1792 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A a_5385_1059# 8.53e-19
C1793 a_26126_1124# VDD 0.929f
C1794 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A 0.0037f
C1795 a_1559_n6471# Q2 5.68e-19
C1796 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A Q7 0.033f
C1797 a_1409_6275# CLK 0.00449f
C1798 OR_magic_1.VOUT divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT 0.00519f
C1799 a_11279_6341# a_8713_6842# 6.34e-20
C1800 a_11279_6341# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A 0.0294f
C1801 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1541_n3597# 6.14e-19
C1802 a_23207_5815# Q7 2.68e-19
C1803 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_6.OUT 0.0153f
C1804 a_12387_9730# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 1.63e-20
C1805 a_26038_684# DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 1.9e-19
C1806 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A VDD 1.38f
C1807 7b_counter_0.MDFF_6.tspc2_magic_0.CLK Q1 0.0867f
C1808 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_20171_6886# 0.112f
C1809 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_8643_n1042# 3.46e-20
C1810 a_1209_2253# CLK 0.223f
C1811 LD Q4 1.93f
C1812 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B 0.00691f
C1813 a_5470_n6471# Q6 0.00199f
C1814 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A D2_1 0.0157f
C1815 a_1209_3363# Q7 0.0097f
C1816 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 0.00178f
C1817 p3_gen_magic_0.3_inp_AND_magic_0.B a_13553_n6613# 0.163f
C1818 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A 0.00305f
C1819 a_13353_n6613# D2_5 0.0257f
C1820 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 2.76e-19
C1821 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p3_gen_magic_0.3_inp_AND_magic_0.A 9.87e-20
C1822 a_1559_n6471# a_1541_n8095# 5.02e-19
C1823 p3_gen_magic_0.xnor_magic_5.OUT D2_5 0.00104f
C1824 a_5470_n1973# Q6 8.88e-19
C1825 p3_gen_magic_0.xnor_magic_4.OUT a_5054_n6471# 0.3f
C1826 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_18891_1669# 1.94e-20
C1827 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT Q5 0.013f
C1828 p3_gen_magic_0.3_inp_AND_magic_0.B a_14756_n8142# 0.00777f
C1829 DFF_magic_0.D 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A 0.00788f
C1830 p2_gen_magic_0.xnor_magic_6.OUT a_8939_n3150# 0.0629f
C1831 a_9059_n6471# Q1 6.09e-19
C1832 7b_counter_0.DFF_magic_0.tg_magic_1.IN CLK 0.839f
C1833 DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_0.IN 0.85f
C1834 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B Q5 3.04e-19
C1835 a_8523_n7648# a_8939_n7648# 0.00222f
C1836 DFF_magic_0.tg_magic_3.CLK Q3 0.0168f
C1837 a_11292_n6613# D2_2 0.00277f
C1838 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A D2_7 0.00176f
C1839 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A 0.00113f
C1840 a_19841_9774# D2_3 0.00296f
C1841 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.xnor_magic_6.OUT 0.0308f
C1842 p3_gen_magic_0.xnor_magic_0.OUT a_8939_n7648# 1.73e-19
C1843 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT VDD 1.17f
C1844 p3_gen_magic_0.3_inp_AND_magic_0.C p3_gen_magic_0.xnor_magic_1.B 0.0107f
C1845 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_5.OUT 5.24e-19
C1846 7b_counter_0.MDFF_1.tspc2_magic_0.CLK Q3 4.27e-19
C1847 a_11279_6341# a_12387_5769# 7.16e-20
C1848 a_12387_552# D2_6 3.07e-19
C1849 7b_counter_0.MDFF_5.LD a_15865_6276# 3.96e-19
C1850 7b_counter_0.DFF_magic_0.tg_magic_2.IN 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.258f
C1851 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 0.00749f
C1852 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT D2_1 4.8e-19
C1853 a_12174_n8579# Q4 0.0369f
C1854 Q3 Q4 0.493f
C1855 Q7 Q6 6.56f
C1856 divide_by_2_1.tg_magic_3.CLK divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT 0.0636f
C1857 a_5054_n1526# Q5 0.00816f
C1858 a_2749_7308# VDD 0.935f
C1859 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B D2_4 0.0218f
C1860 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_3.OUT 2.35e-19
C1861 a_5036_n4081# Q5 1.88e-19
C1862 a_26126_1124# Q3 0.0118f
C1863 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B a_21381_3524# 0.412f
C1864 a_5054_n6024# D2_4 0.104f
C1865 a_13553_n6613# D2_5 0.00409f
C1866 a_8939_n3150# VDD 0.0018f
C1867 a_16065_4557# VDD 0.0609f
C1868 p3_gen_magic_0.xnor_magic_5.OUT D2_7 0.308f
C1869 p2_gen_magic_0.xnor_magic_3.OUT D2_6 0.0434f
C1870 a_24059_4877# a_24536_3947# 0.153f
C1871 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A Q1 0.00426f
C1872 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_0.tspc2_magic_0.D 0.00171f
C1873 a_21381_4932# Q6 4.02e-19
C1874 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A a_27234_3319# 0.00184f
C1875 7b_counter_0.DFF_magic_0.tg_magic_3.CLK a_27234_4513# 0.0157f
C1876 7b_counter_0.MDFF_1.tspc2_magic_0.D a_19152_1223# 0.0384f
C1877 a_8643_n6471# a_8523_n8095# 3.68e-19
C1878 OR_magic_2.A DFF_magic_0.tg_magic_3.CLK 0.0312f
C1879 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A p2_gen_magic_0.3_inp_AND_magic_0.A 0.00113f
C1880 a_14756_n8142# D2_5 0.00324f
C1881 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_15865_3363# 1.08e-19
C1882 7b_counter_0.MDFF_3.QB a_5385_7469# 2.44e-20
C1883 a_2749_7308# LD 0.00115f
C1884 p3_gen_magic_0.xnor_magic_4.OUT D2_3 0.172f
C1885 divide_by_2_0.tg_magic_0.IN divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT 4.89e-20
C1886 7b_counter_0.MDFF_4.LD DFF_magic_0.tg_magic_3.CLK 0.00535f
C1887 mux_magic_0.OR_magic_0.B VDD 1.19f
C1888 a_1209_2253# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B 0.125f
C1889 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A a_5185_1059# 0.128f
C1890 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A a_4235_3947# 6.32e-20
C1891 a_17405_5901# a_15865_6276# 7.98e-19
C1892 a_5054_n6024# Q2 0.0805f
C1893 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_4496_4393# 0.51f
C1894 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_1.tspc2_magic_0.CLK 0.086f
C1895 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT Q4 0.0442f
C1896 a_12387_552# D2_2 0.00341f
C1897 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_1209_2253# 1.08e-19
C1898 a_11279_1124# a_9689_1669# 2.12e-20
C1899 a_6725_7308# a_8713_6842# 0.00152f
C1900 a_22991_5815# Q7 4.31e-19
C1901 7b_counter_0.MDFF_4.LD Q4 3.33f
C1902 a_16065_9774# Q1 5.64e-20
C1903 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_19307_6886# 0.0618f
C1904 a_27234_1746# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A 0.00184f
C1905 divide_by_2_0.tg_magic_3.IN VDD 2.5f
C1906 a_5054_n1526# Q2 0.0805f
C1907 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_9412_5956# 0.35f
C1908 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT Q4 1.93e-19
C1909 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT D2_6 0.00199f
C1910 a_5054_n6471# Q6 0.0341f
C1911 p3_gen_magic_0.3_inp_AND_magic_0.B a_11708_n6613# 0.00272f
C1912 7b_counter_0.MDFF_4.LD a_26126_1124# 0.00115f
C1913 divide_by_2_0.tg_magic_3.IN D2_1 1.19f
C1914 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A a_1409_9773# 9.27e-19
C1915 p2_gen_magic_0.xnor_magic_3.OUT D2_2 0.19f
C1916 a_5054_n1973# p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 0.00271f
C1917 a_5036_n7648# D2_5 0.00377f
C1918 p3_gen_magic_0.xnor_magic_4.OUT a_8643_n6024# 2.24e-19
C1919 a_5054_n1973# Q6 0.00892f
C1920 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 0.00177f
C1921 7b_counter_0.MDFF_3.tspc2_magic_0.Q VDD 1.39f
C1922 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK D2_3 0.00402f
C1923 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_9689_1669# 0.0618f
C1924 a_8523_n3150# a_8939_n3150# 0.00222f
C1925 p2_gen_magic_0.3_inp_AND_magic_0.A p2_gen_magic_0.3_inp_AND_magic_0.C 0.0449f
C1926 a_8643_n6471# Q1 0.302f
C1927 p3_gen_magic_0.3_inp_AND_magic_0.B a_16186_n8142# 0.0437f
C1928 7b_counter_0.3_inp_AND_magic_0.VOUT 7b_counter_0.DFF_magic_0.D 0.785f
C1929 7b_counter_0.MDFF_3.tspc2_magic_0.Q D2_1 0.00109f
C1930 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_5.OUT 4.35e-20
C1931 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.3_inp_AND_magic_0.VOUT 1.75e-19
C1932 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q5 8.52e-19
C1933 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 5.61e-19
C1934 a_5185_7469# D2_7 0.223f
C1935 a_8411_9730# Q7 0.0241f
C1936 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B CLK 0.00118f
C1937 divide_by_2_0.tg_magic_3.CLK divide_by_2_0.tg_magic_1.IN 0.0617f
C1938 a_11279_1124# 7b_counter_0.MDFF_4.tspc2_magic_0.D 0.123f
C1939 a_1559_n6024# Q5 7.45e-19
C1940 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT 0.0086f
C1941 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B p2_gen_magic_0.xnor_magic_0.OUT 0.00107f
C1942 a_8523_n8095# Q1 1.86e-20
C1943 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.xnor_magic_4.OUT 0.354f
C1944 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A a_15865_8580# 0.00184f
C1945 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B Q5 0.00368f
C1946 7b_counter_0.MDFF_5.LD a_12931_6276# 0.00242f
C1947 DFF_magic_0.tg_magic_3.OUT CLK 0.441f
C1948 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B Q7 0.0779f
C1949 7b_counter_0.MDFF_3.tspc2_magic_0.Q LD 0.12f
C1950 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 0.089f
C1951 a_1409_9773# a_1409_8579# 0.0142f
C1952 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A a_6725_5900# 0.397f
C1953 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN 4.63e-20
C1954 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A a_1209_3363# 1.03e-19
C1955 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A Q7 0.0249f
C1956 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT 0.229f
C1957 a_27234_3319# a_27778_3363# 0.298f
C1958 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT VDD 1.48f
C1959 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT D2_4 3.24e-19
C1960 a_1559_n6024# p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT 6.69e-21
C1961 a_9212_739# VDD 0.969f
C1962 7b_counter_0.3_inp_AND_magic_0.B 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B 2.65e-20
C1963 a_1559_n6024# D2_4 0.239f
C1964 a_11708_n6613# D2_5 0.0189f
C1965 p2_gen_magic_0.xnor_magic_0.OUT D2_3 1.73e-19
C1966 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A Q7 3.39e-19
C1967 p3_gen_magic_0.3_inp_AND_magic_0.C p3_gen_magic_0.xnor_magic_1.OUT 0.0176f
C1968 a_5515_3947# VDD 0.0859f
C1969 a_5036_n7648# D2_7 0.0578f
C1970 Q6 D2_3 0.0989f
C1971 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1541_n3150# 4.77e-19
C1972 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B a_2749_3524# 0.412f
C1973 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 7b_counter_0.MDFF_4.tspc2_magic_0.D 0.399f
C1974 a_24059_4877# a_23672_3947# 0.00652f
C1975 7b_counter_0.MDFF_4.tspc2_magic_0.CLK p2_gen_magic_0.xnor_magic_4.OUT 9.91e-20
C1976 a_23258_1746# 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 1.03e-19
C1977 a_20041_3363# Q1 0.0131f
C1978 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_19841_4557# 0.223f
C1979 a_8411_9730# a_8955_9774# 0.297f
C1980 p2_gen_magic_0.AND2_magic_1.A p3_gen_magic_0.3_inp_AND_magic_0.VOUT 1.34e-19
C1981 a_8411_8536# Q7 5.24e-19
C1982 7b_counter_0.MDFF_1.tspc2_magic_0.D a_18891_1669# 0.278f
C1983 a_1559_n1526# D2_4 0.231f
C1984 a_16065_4557# a_15865_3363# 0.00308f
C1985 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A Q7 0.031f
C1986 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B a_17405_8741# 0.412f
C1987 a_4496_9609# Q6 3.63e-19
C1988 a_1209_2253# a_1409_2253# 0.298f
C1989 a_20171_6886# Q1 0.00228f
C1990 a_1559_n6024# Q2 0.00423f
C1991 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT Q5 0.00211f
C1992 7b_counter_0.MDFF_4.LD a_16065_4557# 0.00357f
C1993 a_23560_3728# Q4 0.00344f
C1994 a_12590_n7648# a_12174_n8095# 0.013f
C1995 a_5515_3947# LD 8.29e-19
C1996 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A Q6 0.0155f
C1997 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_22150_1124# 6.72e-19
C1998 7b_counter_0.MDFF_5.LD a_8713_6842# 0.00664f
C1999 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_17405_5901# 0.00215f
C2000 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A 1.1e-20
C2001 mux_magic_0.IN1 mux_magic_0.OR_magic_0.B 1.06e-19
C2002 a_8411_4513# 7b_counter_0.MDFF_4.tspc2_magic_0.Q 0.223f
C2003 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5036_n7648# 5.22e-19
C2004 a_23352_n6798# VDD 0.976f
C2005 a_27234_1746# a_26126_1124# 0.00114f
C2006 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A Q4 0.00101f
C2007 a_1541_n4081# Q2 0.00271f
C2008 7b_counter_0.MDFF_6.tspc2_magic_0.D VDD 1.39f
C2009 p3_gen_magic_0.3_inp_AND_magic_0.B a_11492_n6613# 7.27e-19
C2010 a_6725_5900# Q6 0.0264f
C2011 a_11292_n2115# a_11708_n2115# 0.278f
C2012 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT Q4 0.0201f
C2013 a_23352_n6798# D2_1 0.0239f
C2014 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_4 0.981f
C2015 7b_counter_0.DFF_magic_0.tg_magic_2.IN CLK 0.0147f
C2016 mux_magic_0.OR_magic_0.A VDD 1.23f
C2017 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT D2_5 0.106f
C2018 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5054_n1526# 0.0821f
C2019 7b_counter_0.MDFF_6.tspc2_magic_0.D D2_1 0.00827f
C2020 OR_magic_2.A divide_by_2_0.tg_magic_3.IN 0.00136f
C2021 p2_gen_magic_0.xnor_magic_0.OUT a_8643_n1526# 0.415f
C2022 a_1409_1059# D2_5 0.00121f
C2023 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT VDD 1.36f
C2024 a_4235_9163# VDD 1.06f
C2025 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_8825_1669# 0.112f
C2026 7b_counter_0.3_inp_AND_magic_0.VOUT Q1 1.62e-19
C2027 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A 1.19e-19
C2028 p3_gen_magic_0.3_inp_AND_magic_0.B a_14556_n8142# 0.127f
C2029 mux_magic_0.OR_magic_0.A D2_1 1.1e-20
C2030 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 7b_counter_0.MDFF_0.tspc2_magic_0.Q 0.0189f
C2031 a_2749_2092# a_1209_1059# 7.16e-20
C2032 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A Q6 3.37e-19
C2033 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A 0.00108f
C2034 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT D2_1 8.59e-19
C2035 a_4235_9163# D2_1 0.0021f
C2036 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT Q7 0.00572f
C2037 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_6 1.13f
C2038 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B Q1 0.0124f
C2039 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT CLK 2.41e-19
C2040 a_5054_n1042# Q5 0.00879f
C2041 a_11292_n6613# p3_gen_magic_0.3_inp_AND_magic_0.C 2.07e-19
C2042 p3_gen_magic_0.xnor_magic_3.OUT a_13353_n6613# 0.00201f
C2043 a_8713_1625# Q5 0.00762f
C2044 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT Q2 0.0585f
C2045 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_1.tspc2_magic_0.CLK 8.78e-21
C2046 p3_gen_magic_0.xnor_magic_4.OUT a_5452_n7648# 7.38e-19
C2047 p3_gen_magic_0.xnor_magic_1.B p3_gen_magic_0.xnor_magic_1.OUT 0.458f
C2048 7b_counter_0.MDFF_5.LD a_12387_5769# 3.96e-19
C2049 a_7303_3480# Q5 0.00756f
C2050 7b_counter_0.DFF_magic_0.D 7b_counter_0.MDFF_5.LD 0.0518f
C2051 7b_counter_0.MDFF_3.QB 7b_counter_0.MDFF_3.tspc2_magic_0.Q 0.292f
C2052 7b_counter_0.MDFF_7.tspc2_magic_0.Q 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A 0.00118f
C2053 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A 0.178f
C2054 a_4235_9163# LD 2.62e-21
C2055 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT 0.54f
C2056 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT D2_5 0.0536f
C2057 7b_counter_0.MDFF_5.tspc2_magic_0.Q D2_6 0.0433f
C2058 a_13553_n2115# a_13769_n2115# 0.326f
C2059 7b_counter_0.MDFF_5.LD a_16065_9774# 0.0341f
C2060 p2_gen_magic_0.3_inp_AND_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK 0.429f
C2061 a_7215_4932# a_7303_3480# 0.475f
C2062 a_5054_n1042# D2_4 1.31e-19
C2063 a_8713_1625# D2_4 7.9e-19
C2064 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A a_7303_3480# 0.0334f
C2065 a_11492_n6613# D2_5 0.0289f
C2066 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A D2_5 0.00477f
C2067 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A a_23802_1059# 9.27e-19
C2068 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN 0.965f
C2069 a_4651_3947# VDD 0.0502f
C2070 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT VDD 1.03f
C2071 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1541_n8095# 5.59e-19
C2072 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_1.OUT 0.24f
C2073 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 0.00894f
C2074 a_27778_2253# CLK 0.196f
C2075 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B a_2749_4932# 0.173f
C2076 a_1409_1059# D2_7 0.0195f
C2077 a_6725_684# a_5185_1059# 7.98e-19
C2078 p2_gen_magic_0.AND2_magic_1.A a_13353_n6613# 3.76e-20
C2079 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_27234_3319# 4.8e-20
C2080 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 0.0213f
C2081 a_20041_9774# Q7 0.0329f
C2082 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B p2_gen_magic_0.xnor_magic_3.OUT 1.55e-19
C2083 a_14556_n8142# D2_5 0.00162f
C2084 a_26038_4932# a_26126_3480# 0.475f
C2085 divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT VDD 1.09f
C2086 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A VDD 1.23f
C2087 a_5185_2253# Q7 0.012f
C2088 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_2 0.0114f
C2089 a_21381_4932# a_19841_3363# 1.14e-19
C2090 p3_gen_magic_0.xnor_magic_3.OUT a_13553_n6613# 3.87e-19
C2091 a_5054_n1042# Q2 0.00355f
C2092 divide_by_2_1.tg_magic_3.CLK divide_by_2_1.tg_magic_0.IN 0.164f
C2093 a_12590_n3150# a_12174_n3597# 0.013f
C2094 a_19307_6886# a_20171_6886# 0.00862f
C2095 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A a_2749_8740# 0.0334f
C2096 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.26f
C2097 a_19307_6886# Q1 0.0148f
C2098 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A D2_1 0.0145f
C2099 a_21381_3524# Q1 0.11f
C2100 a_6725_2092# a_8825_1669# 1.19e-20
C2101 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A 9.4e-20
C2102 a_23793_5904# Q4 0.356f
C2103 p2_gen_magic_0.xnor_magic_5.OUT Q5 0.0322f
C2104 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 0.00618f
C2105 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A 0.178f
C2106 a_5470_n6471# VDD 0.00291f
C2107 7b_counter_0.MDFF_5.tspc2_magic_0.Q D2_2 0.418f
C2108 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT D2_7 0.00376f
C2109 a_12387_8536# Q7 4.58e-19
C2110 a_9689_6886# VDD 0.00407f
C2111 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A LD 5.51e-19
C2112 a_4651_9163# a_5515_9163# 0.00862f
C2113 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A VDD 1.29f
C2114 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A D2_7 0.088f
C2115 a_11292_n2115# a_11492_n2115# 0.519f
C2116 a_5054_n5540# D2_5 0.0385f
C2117 a_1209_9773# a_1409_9773# 0.297f
C2118 a_5185_1059# Q5 0.0151f
C2119 a_8411_9730# a_7215_10149# 7.98e-19
C2120 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT D2_7 9.85e-19
C2121 a_20041_8580# D2_3 8.6e-19
C2122 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT 0.469f
C2123 a_5470_n1973# VDD 0.00361f
C2124 a_8411_9730# 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A 0.128f
C2125 OR_magic_2.A a_23352_n6798# 0.0334f
C2126 a_1559_n5540# VDD 0.414f
C2127 a_1209_1059# D2_5 0.00166f
C2128 7b_counter_0.DFF_magic_0.Q 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 4.95e-19
C2129 a_23258_1746# CLK 0.0567f
C2130 a_4496_10093# VDD 0.763f
C2131 a_5452_n7648# Q6 0.00158f
C2132 p2_gen_magic_0.xnor_magic_5.OUT D2_4 0.00761f
C2133 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_20041_4557# 0.12f
C2134 p2_gen_magic_0.xnor_magic_1.OUT Q1 0.0108f
C2135 a_27234_4513# a_26038_4932# 7.98e-19
C2136 p2_gen_magic_0.xnor_magic_3.OUT a_12174_n3597# 2.99e-20
C2137 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_8523_n3150# 3.55e-19
C2138 a_12387_9730# Q6 3.77e-19
C2139 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_4235_3947# 0.654f
C2140 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A 0.0042f
C2141 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_6.tspc2_magic_0.D 0.00851f
C2142 a_4496_10093# D2_1 0.00321f
C2143 mux_magic_0.IN1 mux_magic_0.OR_magic_0.A 0.00129f
C2144 divide_by_2_0.tg_magic_3.CLK divide_by_2_0.tg_magic_3.IN 0.951f
C2145 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_1.OUT 9.88e-19
C2146 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A a_16065_4557# 0.0292f
C2147 7b_counter_0.MDFF_4.tspc2_magic_0.CLK Q4 0.00162f
C2148 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 7b_counter_0.MDFF_1.tspc2_magic_0.Q 0.00105f
C2149 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT Q3 5.29e-19
C2150 a_5185_1059# D2_4 7.56e-19
C2151 p3_gen_magic_0.3_inp_AND_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.00569f
C2152 p3_gen_magic_0.xnor_magic_1.B a_1541_n7648# 0.0839f
C2153 VDD Q7 8.54f
C2154 7b_counter_0.MDFF_5.LD a_20171_6886# 8.29e-19
C2155 7b_counter_0.MDFF_5.tspc2_magic_0.Q 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A 0.255f
C2156 7b_counter_0.MDFF_5.LD Q1 0.206f
C2157 7b_counter_0.MDFF_4.tspc2_magic_0.D 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A 8.78e-21
C2158 p2_gen_magic_0.xnor_magic_5.OUT Q2 1.22e-20
C2159 7b_counter_0.MDFF_3.QB a_4235_9163# 0.0278f
C2160 a_16065_7470# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A 1.77e-19
C2161 D2_1 Q7 0.343f
C2162 a_13353_n2115# p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK 1.16e-20
C2163 a_7215_10149# a_8411_8536# 1.14e-19
C2164 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_0.tspc2_magic_0.D 2.05e-19
C2165 p2_gen_magic_0.3_inp_AND_magic_0.C p2_gen_magic_0.AND2_magic_1.A 0.00428f
C2166 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT 0.195f
C2167 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A a_8411_8536# 0.00184f
C2168 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT 0.153f
C2169 a_9059_n6471# D2_5 0.00231f
C2170 a_1209_6275# a_1409_6275# 0.297f
C2171 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B Q2 0.0496f
C2172 a_21381_4932# VDD 1.56f
C2173 mux_magic_0.IN2 P2 4.03e-19
C2174 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 0.0214f
C2175 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT a_1541_n3150# 0.0088f
C2176 a_20171_1669# CLK 0.002f
C2177 a_1209_1059# D2_7 0.0168f
C2178 LD Q7 0.164f
C2179 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A D2_3 0.103f
C2180 a_2749_2092# 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A 2.4e-20
C2181 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_24536_3947# 0.0618f
C2182 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A a_17405_4932# 1.51e-21
C2183 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B a_7303_8697# 0.412f
C2184 a_19841_3363# D2_3 0.223f
C2185 a_12174_n8095# D2_5 0.24f
C2186 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_5185_7469# 4.65e-19
C2187 p3_gen_magic_0.AND2_magic_1.A D2_6 0.0933f
C2188 7b_counter_0.MDFF_7.tspc2_magic_0.Q a_24059_4877# 1.94e-20
C2189 a_8955_9774# VDD 0.0935f
C2190 7b_counter_0.MDFF_5.tspc2_magic_0.Q CLK 0.0701f
C2191 7b_counter_0.3_inp_AND_magic_0.VOUT 7b_counter_0.MDFF_5.LD 0.102f
C2192 p3_gen_magic_0.xnor_magic_3.OUT a_11708_n6613# 0.0446f
C2193 p3_gen_magic_0.3_inp_AND_magic_0.VOUT Q4 0.195f
C2194 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_19152_1223# 0.51f
C2195 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A Q3 0.352f
C2196 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A 0.178f
C2197 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A a_2749_10148# 0.397f
C2198 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B Q6 0.0104f
C2199 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN 0.659f
C2200 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 3.8e-19
C2201 a_1209_9773# 7b_counter_0.MDFF_3.tspc2_magic_0.D 1.63e-20
C2202 a_19152_1223# Q4 2.83e-19
C2203 7b_counter_0.3_inp_AND_magic_0.B Q1 0.0584f
C2204 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A a_9212_739# 3.22e-21
C2205 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A VDD 1.29f
C2206 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A a_15865_9774# 0.251f
C2207 a_1559_n5540# Q3 2.81e-19
C2208 a_21504_5904# Q4 0.00237f
C2209 a_20041_9774# D2_3 0.00138f
C2210 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A Q2 0.00108f
C2211 a_2749_5900# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A 1.52e-21
C2212 a_8713_6842# a_8411_4513# 1.73e-19
C2213 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.3_inp_AND_magic_0.B 0.0103f
C2214 a_11292_n2115# p2_gen_magic_0.3_inp_AND_magic_0.A 0.116f
C2215 a_23985_7877# Q4 7.55e-20
C2216 p2_gen_magic_0.xnor_magic_0.OUT a_13353_n2115# 1.73e-20
C2217 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5054_n1042# 0.0582f
C2218 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B D2_3 0.00564f
C2219 a_5036_n3150# Q5 3.01e-19
C2220 Q5 D2_6 1.57f
C2221 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A D2_4 0.103f
C2222 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B 0.00112f
C2223 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B a_26126_1124# 0.412f
C2224 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5054_n5540# 0.0846f
C2225 7b_counter_0.MDFF_5.tspc2_magic_0.Q a_11279_8697# 0.00137f
C2226 a_5054_n6471# VDD 0.0269f
C2227 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.0032f
C2228 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT a_16386_n8142# 2.74e-19
C2229 a_1559_n6471# Q6 7.08e-19
C2230 mux_magic_0.IN2 VDD 2.01f
C2231 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A a_27778_4557# 0.0292f
C2232 a_8825_6886# VDD 0.075f
C2233 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT 0.0171f
C2234 a_23258_552# VDD 0.994f
C2235 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A D2_6 0.00222f
C2236 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.3_inp_AND_magic_0.A 2.07e-20
C2237 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_4496_4393# 0.0116f
C2238 mux_magic_0.IN2 D2_1 0.276f
C2239 a_1559_n1042# a_1559_n1526# 0.0335f
C2240 p3_gen_magic_0.xnor_magic_6.OUT VDD 1.38f
C2241 Q3 Q7 0.922f
C2242 a_5054_n1973# VDD 0.0325f
C2243 a_19307_1669# a_19152_739# 0.00164f
C2244 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT 0.0032f
C2245 7b_counter_0.MDFF_4.tspc2_magic_0.D a_11191_684# 1.08e-19
C2246 D2_6 D2_4 1.09f
C2247 p3_gen_magic_0.xnor_magic_4.OUT a_5054_n6024# 0.415f
C2248 a_1409_9773# VDD 0.0523f
C2249 a_11191_684# p2_gen_magic_0.xnor_magic_4.OUT 1.34e-19
C2250 p2_gen_magic_0.xnor_magic_6.OUT D2_3 0.14f
C2251 7b_counter_0.MDFF_5.tspc2_magic_0.D 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 2.05e-19
C2252 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_4496_4877# 0.35f
C2253 OR_magic_2.A 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 2.72e-20
C2254 7b_counter_0.3_inp_AND_magic_0.VOUT 7b_counter_0.3_inp_AND_magic_0.B 0.00395f
C2255 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT a_5036_n8579# 0.057f
C2256 a_13769_n6613# Q4 0.00917f
C2257 a_1409_9773# D2_1 0.0175f
C2258 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 0.413f
C2259 DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT P2 0.00143f
C2260 7b_counter_0.DFF_magic_0.D 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 0.589f
C2261 a_12387_9730# 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A 0.251f
C2262 a_5185_7469# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B 0.125f
C2263 a_1409_4557# CLK 7.14e-19
C2264 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 0.00956f
C2265 7b_counter_0.MDFF_4.tspc2_magic_0.Q a_9689_1669# 0.00409f
C2266 a_16065_7470# 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 0.00103f
C2267 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1541_n7648# 0.00283f
C2268 divide_by_2_0.tg_magic_3.CLK a_23352_n6798# 1.85e-19
C2269 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B VDD 1.2f
C2270 a_21381_4932# Q3 0.0012f
C2271 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_5.OUT 0.00982f
C2272 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B CLK 0.0105f
C2273 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN VDD 2.03f
C2274 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B a_11279_3480# 0.412f
C2275 7b_counter_0.MDFF_5.tspc2_magic_0.D VDD 1.39f
C2276 a_17405_2092# 7b_counter_0.MDFF_1.tspc2_magic_0.D 0.123f
C2277 D2_2 Q5 0.123f
C2278 a_5036_n3150# Q2 0.00136f
C2279 Q2 D2_6 0.25f
C2280 7b_counter_0.MDFF_3.QB a_4496_10093# 3.52e-19
C2281 a_1409_9773# LD 0.00391f
C2282 a_15865_2253# 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 1.03e-19
C2283 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B 7b_counter_0.MDFF_7.tspc2_magic_0.Q 1.17e-20
C2284 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN D2_1 0.0532f
C2285 divide_by_2_1.tg_magic_3.CLK divide_by_2_1.tg_magic_3.OUT 0.537f
C2286 a_7303_8697# a_5515_9163# 1.36e-20
C2287 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B 0.00234f
C2288 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT Q5 3.73e-19
C2289 a_8643_n6471# D2_5 0.0634f
C2290 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_5.OUT 9.88e-19
C2291 VDD D2_3 5.78f
C2292 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B VDD 1.2f
C2293 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A D2_5 0.0126f
C2294 a_15865_7470# Q2 5.69e-19
C2295 7b_counter_0.MDFF_3.QB Q7 5.73e-19
C2296 a_19307_1669# CLK 0.00196f
C2297 a_1541_n7648# p3_gen_magic_0.xnor_magic_1.OUT 0.0925f
C2298 D2_2 D2_4 0.0841f
C2299 DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD 1.09f
C2300 D2_1 D2_3 2.17f
C2301 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A CLK 0.307f
C2302 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT Q7 0.0256f
C2303 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_23672_3947# 0.112f
C2304 DFF_magic_0.tg_magic_3.CLK DFF_magic_0.tg_magic_2.OUT 0.469f
C2305 7b_counter_0.MDFF_0.tspc2_magic_0.Q p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 0.00168f
C2306 a_21381_8741# Q7 0.0519f
C2307 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A a_5385_6275# 9.27e-19
C2308 a_16065_2253# 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 0.00103f
C2309 a_8523_n8095# D2_5 0.00185f
C2310 a_4496_9609# VDD 1.07f
C2311 a_23258_552# Q3 3.93e-19
C2312 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_18891_1669# 0.654f
C2313 7b_counter_0.MDFF_7.tspc2_magic_0.D 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A 8.78e-21
C2314 p3_gen_magic_0.xnor_magic_3.OUT a_11492_n6613# 0.00138f
C2315 a_13353_n6613# Q4 0.0219f
C2316 a_8643_n6471# p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT 7.47e-19
C2317 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT D2_4 0.00344f
C2318 p3_gen_magic_0.xnor_magic_5.OUT Q4 0.0641f
C2319 a_1209_9773# a_2749_8740# 7.16e-20
C2320 a_4496_9609# D2_1 0.00131f
C2321 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A VDD 1.29f
C2322 a_18891_1669# Q4 7.16e-21
C2323 7b_counter_0.DFF_magic_0.Q CLK 1.33f
C2324 LD D2_3 0.0167f
C2325 a_11279_1124# a_9212_739# 0.00212f
C2326 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT Q6 0.00618f
C2327 7b_counter_0.MDFF_3.tspc2_magic_0.D VDD 1.4f
C2328 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_0.IN 0.85f
C2329 a_15865_9774# Q2 9.61e-19
C2330 Q2 D2_2 0.257f
C2331 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT a_8523_n8095# 0.0629f
C2332 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A D2_1 6.27e-20
C2333 a_7303_8697# a_6725_7308# 1.62e-19
C2334 a_19152_739# D2_4 0.0131f
C2335 a_8643_n6024# VDD 0.181f
C2336 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A a_16065_8580# 1.77e-19
C2337 7b_counter_0.MDFF_3.tspc2_magic_0.D D2_1 0.00592f
C2338 a_17405_684# p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 1.78e-19
C2339 a_26126_3480# a_26126_1124# 0.00112f
C2340 a_5054_n6024# Q6 0.0335f
C2341 a_4496_9609# LD 0.00751f
C2342 a_6725_5900# VDD 1.55f
C2343 a_26038_684# VDD 1.55f
C2344 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A OR_magic_2.A 1.39e-19
C2345 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B Q3 2.69e-19
C2346 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_20041_3363# 0.017f
C2347 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A D2_7 0.0996f
C2348 a_4235_3947# a_4496_4393# 0.299f
C2349 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A 0.405f
C2350 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A Q4 0.00146f
C2351 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.P3 6.97e-20
C2352 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B a_1209_3363# 0.125f
C2353 a_8523_n7648# VDD 0.0014f
C2354 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT D2_7 0.00494f
C2355 a_8643_n1526# VDD 0.181f
C2356 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A LD 0.412f
C2357 a_5054_n1526# p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 6.69e-21
C2358 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A a_17405_8741# 2.4e-20
C2359 a_12387_552# a_12931_1059# 0.297f
C2360 7b_counter_0.MDFF_3.tspc2_magic_0.D LD 8.18e-19
C2361 a_5054_n1526# Q6 1.77e-20
C2362 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A Q2 7.6e-19
C2363 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A D2_6 5.77e-19
C2364 a_7215_10149# VDD 1.55f
C2365 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_2.IN 6.95e-19
C2366 p3_gen_magic_0.xnor_magic_0.OUT VDD 0.632f
C2367 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT Q5 3.72e-19
C2368 mux_magic_0.IN1 mux_magic_0.IN2 0.0039f
C2369 a_9212_5956# Q2 0.0979f
C2370 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT a_5036_n4081# 0.057f
C2371 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_1.IN 1.16f
C2372 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_9212_739# 0.654f
C2373 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A VDD 1.23f
C2374 a_27234_1746# 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 1.03e-19
C2375 OR_magic_2.A mux_magic_0.IN2 0.0108f
C2376 Q1 D2_5 0.214f
C2377 7b_counter_0.DFF_magic_0.Q 7b_counter_0.3_inp_AND_magic_0.C 0.003f
C2378 CLK Q5 0.219f
C2379 a_5036_n4081# Q6 0.015f
C2380 7b_counter_0.MDFF_1.tspc2_magic_0.Q Q1 0.0862f
C2381 a_13553_n6613# Q4 0.00458f
C2382 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A Q2 7.6e-19
C2383 p3_gen_magic_0.xnor_magic_0.OUT D2_1 0.00576f
C2384 7b_counter_0.MDFF_4.LD a_23258_552# 0.00147f
C2385 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A a_16065_6276# 9.27e-19
C2386 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 0.0338f
C2387 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_6.OUT 0.0372f
C2388 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT Q5 0.513f
C2389 a_5385_6275# Q6 1.77e-19
C2390 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A D2_1 3.01e-19
C2391 7b_counter_0.MDFF_4.tspc2_magic_0.Q a_8825_1669# 5.37e-19
C2392 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A a_2749_7308# 0.0334f
C2393 a_5185_7469# a_5385_7469# 0.296f
C2394 Q3 D2_3 1.98f
C2395 p3_gen_magic_0.xnor_magic_3.OUT a_5054_n5540# 0.128f
C2396 7b_counter_0.MDFF_5.tspc2_magic_0.CLK D2_6 0.503f
C2397 a_15865_2253# VDD 0.884f
C2398 p2_gen_magic_0.3_inp_AND_magic_0.A a_13769_n2115# 0.0247f
C2399 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B Q3 2.23e-19
C2400 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A Q2 0.00109f
C2401 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_3 0.00277f
C2402 a_1409_7469# CLK 0.125f
C2403 7b_counter_0.MDFF_5.LD 7b_counter_0.3_inp_AND_magic_0.B 8.74e-20
C2404 a_8411_4513# Q1 8.5e-19
C2405 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_6.tspc2_magic_0.D 0.00171f
C2406 a_14756_n8142# Q4 0.0349f
C2407 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B a_11191_4932# 0.173f
C2408 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT D2_4 1.13e-19
C2409 7b_counter_0.MDFF_3.QB a_1409_9773# 0.122f
C2410 CLK D2_4 0.923f
C2411 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A LD 5.51e-19
C2412 7b_counter_0.3_inp_AND_magic_0.A CLK 2.69e-19
C2413 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A a_12931_3363# 0.00103f
C2414 7b_counter_0.MDFF_5.LD a_21381_10149# 0.00606f
C2415 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_2.IN 6.95e-19
C2416 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B Q6 0.0137f
C2417 a_12387_4513# D2_2 0.013f
C2418 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A Q4 5.53e-19
C2419 p3_gen_magic_0.3_inp_AND_magic_0.A D2_2 1.35e-20
C2420 7b_counter_0.3_inp_AND_magic_0.C Q5 0.297f
C2421 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5036_n3150# 0.0028f
C2422 p2_gen_magic_0.3_inp_AND_magic_0.C Q4 0.309f
C2423 a_1541_n3150# p2_gen_magic_0.xnor_magic_1.OUT 0.0924f
C2424 a_16065_2253# VDD 0.0179f
C2425 DFF_magic_0.tg_magic_2.IN P2 0.00821f
C2426 a_12387_6963# Q2 0.0938f
C2427 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B D2_5 0.00145f
C2428 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_5.tspc2_magic_0.D 0.00851f
C2429 a_9059_n1973# Q1 0.00128f
C2430 a_23258_1746# a_22062_684# 1.14e-19
C2431 a_21381_3524# a_23672_3947# 6.59e-21
C2432 a_16065_3363# Q1 0.0108f
C2433 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A a_19841_8580# 1.03e-19
C2434 CLK Q2 0.39f
C2435 a_8955_8580# D2_2 0.125f
C2436 a_16065_1059# Q5 8.32e-19
C2437 divide_by_2_1.tg_magic_0.IN divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT 0.26f
C2438 a_5036_n8095# D2_5 5.71e-19
C2439 a_15865_3363# D2_3 4e-19
C2440 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A a_5185_6275# 0.128f
C2441 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A a_26038_4932# 0.397f
C2442 a_26038_684# Q3 0.0113f
C2443 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_8643_n6024# 0.0629f
C2444 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 0.00238f
C2445 a_5515_9163# D2_7 4.39e-19
C2446 a_12387_9730# a_12387_8536# 0.00638f
C2447 7b_counter_0.3_inp_AND_magic_0.C D2_4 0.0288f
C2448 7b_counter_0.MDFF_4.LD D2_3 0.872f
C2449 7b_counter_0.MDFF_5.tspc2_magic_0.CLK D2_2 0.0552f
C2450 a_1209_9773# a_2749_10148# 7.98e-19
C2451 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B 9.09e-19
C2452 p3_gen_magic_0.xnor_magic_6.OUT a_8523_n8579# 0.462f
C2453 7b_counter_0.3_inp_AND_magic_0.A 7b_counter_0.3_inp_AND_magic_0.C 0.229f
C2454 OR_magic_2.A DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.00128f
C2455 a_1559_n6471# p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT 7.35e-19
C2456 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT a_8523_n3597# 0.0629f
C2457 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT VDD 1.17f
C2458 a_2749_8740# VDD 0.941f
C2459 p2_gen_magic_0.3_inp_AND_magic_0.VOUT VDD 2.04f
C2460 p3_gen_magic_0.xnor_magic_3.OUT a_12174_n8095# 2.99e-20
C2461 7b_counter_0.MDFF_0.tspc2_magic_0.D 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 0.423f
C2462 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_8523_n7648# 3.55e-19
C2463 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_27234_552# 1.63e-20
C2464 a_16065_1059# D2_4 0.0041f
C2465 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 0.228f
C2466 a_19152_6440# 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 9.17e-19
C2467 a_1975_n6471# VDD 0.0018f
C2468 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT a_16186_n8142# 8.71e-20
C2469 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.141f
C2470 a_2749_8740# D2_1 0.00218f
C2471 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 0.229f
C2472 DFF_magic_0.tg_magic_2.IN VDD 1.23f
C2473 7b_counter_0.MDFF_3.QB a_4496_9609# 0.111f
C2474 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B Q5 2.92e-19
C2475 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT Q1 0.0149f
C2476 7b_counter_0.MDFF_0.tspc2_magic_0.Q p2_gen_magic_0.xnor_magic_3.OUT 1.7e-19
C2477 7b_counter_0.3_inp_AND_magic_0.C Q2 0.0812f
C2478 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.3_inp_AND_magic_0.B 2.27e-19
C2479 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_9212_5956# 0.654f
C2480 a_4496_4877# a_4496_4393# 0.0141f
C2481 7b_counter_0.MDFF_6.tspc2_magic_0.Q Q7 0.185f
C2482 a_5452_n7648# VDD 0.0042f
C2483 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A a_8955_8580# 5.46e-20
C2484 a_1975_n1973# VDD 0.0018f
C2485 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT P2 0.312f
C2486 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A a_16065_6276# 0.0292f
C2487 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT 0.265f
C2488 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_11279_3480# 1e-20
C2489 7b_counter_0.MDFF_3.QB 7b_counter_0.MDFF_3.tspc2_magic_0.D 0.00346f
C2490 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.153f
C2491 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT 0.153f
C2492 a_12174_n4081# VDD 0.379f
C2493 a_12387_9730# VDD 0.97f
C2494 a_5036_n8095# D2_7 0.244f
C2495 p3_gen_magic_0.3_inp_AND_magic_0.C p3_gen_magic_0.AND2_magic_1.A 0.00445f
C2496 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1541_n3597# 1.73e-19
C2497 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 0.00315f
C2498 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_6.OUT 0.0371f
C2499 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A VDD 1.3f
C2500 7b_counter_0.MDFF_4.tspc2_magic_0.CLK p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.00152f
C2501 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A CLK 1.75e-19
C2502 a_11708_n6613# Q4 2.92e-19
C2503 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A a_15865_6276# 0.128f
C2504 7b_counter_0.MDFF_4.LD a_26038_684# 0.00267f
C2505 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B D2_4 0.0125f
C2506 a_12387_9730# D2_1 3.33e-19
C2507 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.154f
C2508 a_5185_6275# Q6 5.24e-19
C2509 a_12387_4513# CLK 0.0162f
C2510 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A D2_6 1.41e-19
C2511 a_12387_1746# VDD 0.871f
C2512 p2_gen_magic_0.3_inp_AND_magic_0.A a_13553_n2115# 0.0655f
C2513 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.OUT 0.163f
C2514 7b_counter_0.MDFF_0.tspc2_magic_0.CLK D2_4 5.78e-19
C2515 mux_magic_0.IN2 divide_by_2_0.tg_magic_3.CLK 0.0281f
C2516 a_12387_552# p2_gen_magic_0.xnor_magic_3.OUT 5.56e-20
C2517 a_1209_7469# CLK 0.24f
C2518 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT D2_6 0.00117f
C2519 7b_counter_0.MDFF_3.QB a_7215_10149# 1.88e-20
C2520 a_12387_9730# LD 6.64e-19
C2521 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A CLK 3.05e-19
C2522 a_15865_3363# a_15865_2253# 0.00329f
C2523 a_4235_3947# 7b_counter_0.MDFF_0.tspc2_magic_0.Q 1.94e-20
C2524 a_11492_n2115# a_11708_n2115# 0.326f
C2525 a_8955_8580# CLK 0.00991f
C2526 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A Q2 0.00118f
C2527 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_12387_6963# 4.8e-20
C2528 a_8643_n1042# Q1 0.00125f
C2529 a_13353_n2115# p2_gen_magic_0.xnor_magic_6.OUT 0.0385f
C2530 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A CLK 2.5e-20
C2531 divide_by_2_1.tg_magic_3.CLK a_34156_n2297# 1.79e-19
C2532 a_23672_3947# a_24536_3947# 0.00862f
C2533 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B Q2 2.56e-19
C2534 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT VDD 1.24f
C2535 a_8643_n5540# D2_2 0.0167f
C2536 a_22150_1124# Q4 0.126f
C2537 7b_counter_0.MDFF_4.LD a_15865_2253# 0.195f
C2538 p2_gen_magic_0.xnor_magic_1.OUT D2_5 0.295f
C2539 a_23793_5904# Q7 2.05e-20
C2540 a_32616_n2458# P2 3.9e-19
C2541 a_12931_2253# VDD 0.0124f
C2542 7b_counter_0.MDFF_5.tspc2_magic_0.CLK CLK 0.0381f
C2543 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT 4e-20
C2544 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT Q3 0.138f
C2545 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT VDD 1.04f
C2546 p2_gen_magic_0.xnor_magic_4.OUT a_11292_n2115# 0.315f
C2547 p2_gen_magic_0.3_inp_AND_magic_0.VOUT Q3 0.0207f
C2548 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_5.OUT 0.243f
C2549 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A 0.178f
C2550 a_5385_2253# D2_5 0.122f
C2551 a_8643_n1973# Q1 0.319f
C2552 a_2749_684# Q7 0.00982f
C2553 a_12931_3363# Q1 0.0111f
C2554 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B D2_7 0.00813f
C2555 a_1975_n6471# Q3 2.48e-20
C2556 a_15865_1059# Q5 0.00287f
C2557 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT VDD 1.36f
C2558 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT D2_1 4.91e-19
C2559 a_12590_n7648# D2_5 0.0046f
C2560 a_8939_n7648# D2_6 0.00157f
C2561 7b_counter_0.MDFF_1.tspc2_magic_0.D Q1 0.00608f
C2562 7b_counter_0.MDFF_7.tspc2_magic_0.Q Q1 0.00308f
C2563 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B CLK 0.00333f
C2564 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B VDD 1.2f
C2565 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK a_16386_n3644# 0.0171f
C2566 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 7b_counter_0.MDFF_7.tspc2_magic_0.Q 0.00349f
C2567 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_4.OUT 7.63e-21
C2568 p2_gen_magic_0.xnor_magic_6.OUT a_8523_n4081# 0.462f
C2569 a_4651_9163# D2_7 0.00739f
C2570 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT D2_1 0.0792f
C2571 a_5385_1059# Q6 0.0361f
C2572 a_11279_8697# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 0.121f
C2573 a_15865_9774# a_17405_10149# 7.98e-19
C2574 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A a_19841_9774# 0.251f
C2575 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A D2_2 0.0372f
C2576 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_3.OUT 2.31e-19
C2577 7b_counter_0.MDFF_4.LD a_16065_2253# 0.0292f
C2578 a_1409_1059# Q4 0.121f
C2579 a_1975_n1973# Q3 2.06e-19
C2580 a_24059_4877# Q4 3.69e-19
C2581 a_2749_10148# VDD 1.55f
C2582 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A D2_3 3.7e-19
C2583 a_13353_n2115# VDD 1.23f
C2584 a_2749_3524# 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 0.019f
C2585 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A a_16065_1059# 9.27e-19
C2586 a_15865_1059# D2_4 0.0257f
C2587 p3_gen_magic_0.xnor_magic_1.B p3_gen_magic_0.AND2_magic_1.A 0.00142f
C2588 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT D2_3 3.26e-20
C2589 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A a_19841_8580# 0.00184f
C2590 a_1559_n6471# VDD 0.0151f
C2591 a_5054_n1042# Q6 0.00443f
C2592 a_18891_6886# 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 6.3e-20
C2593 a_11279_3480# D2_6 0.00616f
C2594 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_5185_7469# 0.0276f
C2595 a_2749_10148# D2_1 0.00324f
C2596 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT 0.0214f
C2597 a_32616_n2458# VDD 0.87f
C2598 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A 0.00112f
C2599 7b_counter_0.MDFF_0.tspc2_magic_0.Q 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A 0.00118f
C2600 p2_gen_magic_0.xnor_magic_1.OUT D2_7 0.0652f
C2601 a_7303_3480# Q6 0.141f
C2602 a_1541_n8579# Q7 2.81e-19
C2603 a_32616_n2458# D2_1 0.196f
C2604 7b_counter_0.MDFF_4.LD p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT 6.76e-19
C2605 a_1559_n1973# VDD 0.0151f
C2606 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A a_8955_4557# 9.27e-19
C2607 7b_counter_0.MDFF_4.LD p2_gen_magic_0.3_inp_AND_magic_0.VOUT 6.67e-20
C2608 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A a_15865_6276# 0.251f
C2609 a_17405_684# a_15865_1059# 7.98e-19
C2610 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_11191_4932# 4.22e-19
C2611 OR_magic_2.A DFF_magic_0.tg_magic_2.IN 0.305f
C2612 p3_gen_magic_0.xnor_magic_1.B Q5 0.0461f
C2613 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A a_2749_5900# 3.58e-20
C2614 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK p2_gen_magic_0.xnor_magic_5.OUT 0.005f
C2615 a_8523_n4081# VDD 0.414f
C2616 a_27234_1746# a_26038_684# 1.14e-19
C2617 a_19841_8580# a_19152_6440# 3.03e-19
C2618 7b_counter_0.DFF_magic_0.tg_magic_3.OUT CLK 0.439f
C2619 a_1559_n1973# D2_1 3.7e-19
C2620 7b_counter_0.MDFF_6.tspc2_magic_0.D a_19152_5956# 0.103f
C2621 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A 0.00112f
C2622 p2_gen_magic_0.3_inp_AND_magic_0.B Q5 7.55e-20
C2623 a_15865_4557# CLK 3.56e-19
C2624 a_9412_5956# VDD 0.721f
C2625 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT Q3 0.0915f
C2626 OR_magic_1.VOUT a_32616_n1264# 4.36e-19
C2627 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q4 0.00229f
C2628 7b_counter_0.MDFF_6.tspc2_magic_0.Q D2_3 0.0116f
C2629 p2_gen_magic_0.3_inp_AND_magic_0.A a_11708_n2115# 0.192f
C2630 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A 0.0037f
C2631 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_1.B 0.105f
C2632 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT 0.153f
C2633 a_14556_n8142# Q4 0.0335f
C2634 p3_gen_magic_0.xnor_magic_3.OUT Q1 0.298f
C2635 p3_gen_magic_0.xnor_magic_1.B D2_4 0.00131f
C2636 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 2.82e-19
C2637 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT a_8643_n5540# 8.92e-20
C2638 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1975_n1973# 6.1e-19
C2639 a_11191_5901# Q2 0.0437f
C2640 a_5054_n1973# p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT 5.8e-19
C2641 a_11279_3480# D2_2 0.124f
C2642 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_17405_2092# 0.019f
C2643 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 0.00177f
C2644 DFF_magic_0.D 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 8.02e-19
C2645 p2_gen_magic_0.3_inp_AND_magic_0.B D2_4 0.00225f
C2646 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B P2 7.78e-21
C2647 divide_by_2_1.tg_magic_3.CLK a_34156_n889# 7.92e-19
C2648 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_2.IN 0.965f
C2649 a_17405_3524# CLK 0.0436f
C2650 a_8523_n3597# Q5 0.0805f
C2651 a_8411_3319# Q7 0.00415f
C2652 p3_gen_magic_0.3_inp_AND_magic_0.A p3_gen_magic_0.3_inp_AND_magic_0.C 0.0449f
C2653 7b_counter_0.MDFF_4.LD a_12387_1746# 0.195f
C2654 a_21504_5904# Q7 0.467f
C2655 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_5.OUT 0.243f
C2656 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A CLK 0.00189f
C2657 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B Q4 0.00563f
C2658 p2_gen_magic_0.xnor_magic_5.OUT Q6 0.297f
C2659 a_34156_n2297# OUT1 0.128f
C2660 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A p2_gen_magic_0.xnor_magic_3.OUT 1.55e-19
C2661 a_13353_n2115# Q3 0.00786f
C2662 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT a_5036_n7648# 0.0115f
C2663 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_11279_1124# 0.412f
C2664 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN D2_6 6.72e-19
C2665 a_2749_2092# D2_5 0.0562f
C2666 a_27234_552# a_27778_1059# 0.297f
C2667 a_6725_2092# Q7 0.00432f
C2668 a_1559_n6471# Q3 0.303f
C2669 a_12931_4557# D2_2 0.0012f
C2670 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT CLK 0.00519f
C2671 7b_counter_0.3_inp_AND_magic_0.C a_24401_7877# 0.0446f
C2672 7b_counter_0.MDFF_4.LD p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT 6.94e-19
C2673 a_9689_1669# Q1 0.00188f
C2674 a_21381_3524# 7b_counter_0.MDFF_7.tspc2_magic_0.Q 6.46e-19
C2675 p3_gen_magic_0.xnor_magic_4.OUT D2_6 3.57e-20
C2676 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_26038_4932# 0.00215f
C2677 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A D2_5 0.00213f
C2678 a_5185_1059# Q6 0.0584f
C2679 7b_counter_0.MDFF_0.tspc2_magic_0.D a_4496_4393# 0.0384f
C2680 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A 0.00108f
C2681 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT VDD 1.07f
C2682 7b_counter_0.MDFF_4.LD a_12931_2253# 0.0292f
C2683 a_1209_1059# Q4 0.23f
C2684 a_1559_n6024# p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT 7.02e-19
C2685 a_1559_n1973# Q3 0.305f
C2686 7b_counter_0.DFF_magic_0.tg_magic_2.OUT CLK 0.365f
C2687 OR_magic_2.A p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT 0.00271f
C2688 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B VDD 1.24f
C2689 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_3 1.35e-19
C2690 a_2749_4932# 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 0.00215f
C2691 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN 0.287f
C2692 7b_counter_0.DFF_magic_0.Q 7b_counter_0.DFF_magic_0.tg_magic_1.IN 8.34e-19
C2693 a_22062_684# D2_4 0.0213f
C2694 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A a_15865_1059# 0.128f
C2695 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B D2_3 0.0261f
C2696 p3_gen_magic_0.xnor_magic_1.B a_1541_n8095# 0.302f
C2697 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A a_5385_1059# 0.0292f
C2698 a_11191_4932# D2_6 0.00117f
C2699 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B 0.00594f
C2700 a_5054_n6024# VDD 0.221f
C2701 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN 0.29f
C2702 a_8523_n4081# p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 8.96e-20
C2703 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A a_1409_3363# 0.00103f
C2704 a_15865_4557# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A 0.128f
C2705 p3_gen_magic_0.3_inp_AND_magic_0.B D2_5 0.0317f
C2706 a_17405_10149# a_17405_8741# 0.475f
C2707 a_19841_9774# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A 0.128f
C2708 a_1541_n3150# D2_7 0.00164f
C2709 a_8955_3363# a_8713_1625# 5.39e-19
C2710 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A Q6 4.74e-19
C2711 a_5054_n1526# VDD 0.233f
C2712 a_1409_7469# a_1409_6275# 0.0206f
C2713 7b_counter_0.MDFF_4.LD a_13353_n2115# 9.73e-19
C2714 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q5 0.011f
C2715 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A a_5054_n1042# 7.09e-20
C2716 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK D2_6 0.211f
C2717 a_1209_8579# Q2 0.00318f
C2718 a_5036_n4081# VDD 0.494f
C2719 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A Q7 0.00107f
C2720 7b_counter_0.MDFF_4.tspc2_magic_0.D Q1 0.00374f
C2721 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_5515_9163# 0.112f
C2722 7b_counter_0.MDFF_4.tspc2_magic_0.CLK D2_3 6.8e-19
C2723 p2_gen_magic_0.xnor_magic_4.OUT Q1 0.367f
C2724 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT a_1541_n3597# 0.0834f
C2725 p3_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.AND2_magic_1.A 0.00117f
C2726 a_5385_6275# VDD 0.115f
C2727 OR_magic_1.VOUT mux_magic_0.AND2_magic_0.A 0.00134f
C2728 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.153f
C2729 p3_gen_magic_0.xnor_magic_4.OUT D2_2 0.163f
C2730 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_1.IN 0.316f
C2731 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5036_n7648# 1.55e-19
C2732 p2_gen_magic_0.3_inp_AND_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.00627f
C2733 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A a_17405_3524# 0.0334f
C2734 7b_counter_0.MDFF_4.tspc2_magic_0.Q a_9212_739# 1.94e-20
C2735 a_11292_n2115# Q4 0.0208f
C2736 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_11191_5901# 8.42e-19
C2737 p2_gen_magic_0.3_inp_AND_magic_0.A a_11492_n2115# 1.9e-20
C2738 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B Q1 7.94e-19
C2739 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT 0.0331f
C2740 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT 0.00888f
C2741 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT D2_4 0.0731f
C2742 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A Q6 0.00669f
C2743 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK 1.31f
C2744 a_12174_n8095# Q4 0.0876f
C2745 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1559_n1973# 0.102f
C2746 divide_by_2_0.tg_magic_0.IN divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT 0.26f
C2747 p3_gen_magic_0.xnor_magic_1.OUT Q5 0.077f
C2748 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B VDD 1.2f
C2749 a_11191_4932# D2_2 0.0425f
C2750 a_4496_4877# a_4235_3947# 0.651f
C2751 a_12387_3319# a_12387_1746# 0.00329f
C2752 a_12931_4557# CLK 0.00968f
C2753 a_5385_6275# LD 1.1e-19
C2754 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_6.OUT 6.31e-19
C2755 a_5036_n3597# Q5 2.14e-20
C2756 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT Q5 0.135f
C2757 p2_gen_magic_0.xnor_magic_0.OUT D2_6 0.201f
C2758 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT a_5036_n3150# 0.0115f
C2759 a_26038_4932# a_27234_3319# 1.14e-19
C2760 Q6 D2_6 0.068f
C2761 7b_counter_0.MDFF_7.tspc2_magic_0.Q a_24536_3947# 0.00409f
C2762 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B Q3 0.00469f
C2763 a_5036_n3150# Q6 0.328f
C2764 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q2 0.0673f
C2765 a_12387_1746# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A 0.00184f
C2766 p3_gen_magic_0.3_inp_AND_magic_0.VOUT D2_3 0.0073f
C2767 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_1.OUT 0.277f
C2768 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT D2_6 0.059f
C2769 a_13769_n6613# p3_gen_magic_0.xnor_magic_6.OUT 0.00231f
C2770 a_12931_1059# Q5 4.49e-19
C2771 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN Q4 0.0131f
C2772 a_19152_1223# D2_3 2.21e-19
C2773 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B LD 0.00121f
C2774 a_9412_739# VDD 0.721f
C2775 7b_counter_0.3_inp_AND_magic_0.C a_24185_7877# 0.00138f
C2776 a_8825_1669# Q1 0.00654f
C2777 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK a_16186_n3644# 0.00677f
C2778 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 1.31f
C2779 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_5 0.00704f
C2780 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_3.OUT 0.0201f
C2781 a_2749_3524# a_4496_4393# 7.92e-19
C2782 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B 9.4e-20
C2783 divide_by_2_1.tg_magic_3.CLK mux_magic_0.OR_magic_0.B 9.26e-19
C2784 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_4 3.32e-19
C2785 a_27234_552# DFF_magic_0.tg_magic_1.IN 7.13e-21
C2786 a_1209_8579# a_1209_7469# 0.00329f
C2787 p2_gen_magic_0.3_inp_AND_magic_0.A D2_5 0.00656f
C2788 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 3.44e-20
C2789 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A a_12931_2253# 1.77e-19
C2790 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1541_n8095# 1.73e-19
C2791 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT VDD 1.17f
C2792 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN CLK 0.00111f
C2793 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_1.OUT 0.124f
C2794 a_12931_1059# D2_4 0.00381f
C2795 a_1209_4557# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A 0.128f
C2796 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A a_5185_1059# 0.251f
C2797 a_1559_n6024# VDD 0.181f
C2798 a_5036_n3597# Q2 6.69e-21
C2799 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B VDD 1.2f
C2800 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A a_26126_3480# 2.4e-20
C2801 D2_7 D2_5 0.556f
C2802 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT Q2 0.00596f
C2803 p2_gen_magic_0.xnor_magic_0.OUT D2_2 0.218f
C2804 a_15865_9774# Q6 3.77e-19
C2805 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 0.00594f
C2806 D2_2 Q6 0.059f
C2807 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B 9.09e-19
C2808 a_1559_n1526# VDD 0.181f
C2809 a_1209_7469# a_1409_6275# 0.00308f
C2810 a_13769_n6613# D2_3 0.00184f
C2811 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_4.OUT 5.37e-20
C2812 DFF_magic_0.D CLK 0.957f
C2813 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B a_26038_684# 0.173f
C2814 a_1541_n4081# VDD 0.412f
C2815 a_5185_7469# Q7 0.0357f
C2816 p2_gen_magic_0.xnor_magic_1.OUT p2_gen_magic_0.AND2_magic_1.A 0.0115f
C2817 a_17405_4932# D2_3 0.00247f
C2818 a_1559_n1526# D2_1 5.31e-19
C2819 a_13353_n6613# p3_gen_magic_0.xnor_magic_6.OUT 0.0385f
C2820 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_4651_9163# 0.0618f
C2821 mux_magic_0.IN2 divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT 4.95e-19
C2822 7b_counter_0.MDFF_6.tspc2_magic_0.D a_15865_6276# 1.63e-20
C2823 a_5185_6275# VDD 1.02f
C2824 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B a_6725_7308# 0.412f
C2825 p3_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_6.OUT 0.982f
C2826 p3_gen_magic_0.xnor_magic_1.OUT a_1541_n8095# 0.371f
C2827 a_1541_n4081# D2_1 0.0982f
C2828 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A Q1 1.35e-19
C2829 a_16186_n3644# p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 7.26e-20
C2830 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A Q4 0.295f
C2831 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A CLK 6.07e-20
C2832 a_11191_5901# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A 1.51e-21
C2833 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A Q6 0.0273f
C2834 7b_counter_0.MDFF_0.tspc2_magic_0.Q Q5 6.39e-19
C2835 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_5 0.0858f
C2836 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 1.84e-19
C2837 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK CLK 0.566f
C2838 a_1541_n7648# Q5 0.685f
C2839 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A Q6 3.37e-19
C2840 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT VDD 1.03f
C2841 a_1209_3363# CLK 0.0023f
C2842 a_27234_4513# 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A 0.251f
C2843 a_5185_6275# LD 3.96e-19
C2844 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8523_n3150# 0.00261f
C2845 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A Q6 4.53e-19
C2846 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_1 4.67e-19
C2847 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A a_20041_8580# 5.46e-20
C2848 7b_counter_0.MDFF_7.tspc2_magic_0.Q a_23672_3947# 5.37e-19
C2849 7b_counter_0.MDFF_0.tspc2_magic_0.Q D2_4 8.18e-19
C2850 a_19152_6440# Q6 4.92e-19
C2851 a_12387_1746# a_11279_1124# 0.00114f
C2852 a_13353_n6613# D2_3 0.018f
C2853 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_20041_3363# 0.00751f
C2854 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q3 0.00106f
C2855 p3_gen_magic_0.xnor_magic_1.B p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 0.00123f
C2856 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT a_1541_n7648# 0.0115f
C2857 a_13553_n6613# p3_gen_magic_0.xnor_magic_6.OUT 0.0114f
C2858 a_1541_n7648# D2_4 2.58e-19
C2859 a_1559_n6024# Q3 0.0805f
C2860 a_12387_552# Q5 0.00287f
C2861 a_8955_3363# D2_6 0.125f
C2862 a_13769_n2115# Q4 0.00722f
C2863 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_0.IN 0.85f
C2864 a_18891_1669# D2_3 0.0335f
C2865 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B a_18891_1669# 7.16e-19
C2866 a_5385_1059# VDD 0.109f
C2867 7b_counter_0.3_inp_AND_magic_0.C a_23207_5815# 0.656f
C2868 a_19152_5956# D2_3 0.0594f
C2869 a_1209_4557# D2_5 2.51e-19
C2870 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A CLK 0.0061f
C2871 7b_counter_0.DFF_magic_0.Q 7b_counter_0.DFF_magic_0.tg_magic_2.IN 0.289f
C2872 a_5515_9163# a_5385_7469# 0.00565f
C2873 DFF_magic_0.tg_magic_2.OUT DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.153f
C2874 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A a_7303_3480# 2.4e-20
C2875 7b_counter_0.MDFF_1.tspc2_magic_0.CLK Q1 0.0455f
C2876 p3_gen_magic_0.xnor_magic_6.OUT a_14756_n8142# 0.12f
C2877 a_1559_n1526# Q3 0.0805f
C2878 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B Q2 8.23e-19
C2879 CLK Q6 0.131f
C2880 Q1 Q4 0.0513f
C2881 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A a_23258_552# 0.128f
C2882 7b_counter_0.MDFF_7.tspc2_magic_0.CLK Q4 0.0011f
C2883 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_7 6.27e-21
C2884 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B 0.0047f
C2885 a_5054_n1042# VDD 0.497f
C2886 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT a_1541_n3150# 0.102f
C2887 a_8713_1625# VDD 0.757f
C2888 DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT P2 0.00143f
C2889 p2_gen_magic_0.xnor_magic_3.OUT Q5 0.097f
C2890 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 1.42e-19
C2891 a_12387_552# D2_4 0.0258f
C2892 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT CLK 1.33f
C2893 a_23352_n5390# VDD 1.56f
C2894 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_12387_1746# 4.8e-20
C2895 OR_magic_1.VOUT CLK 0.0154f
C2896 a_8411_9730# D2_2 0.018f
C2897 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A D2_3 0.00233f
C2898 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK 2.19e-20
C2899 a_7303_3480# VDD 0.929f
C2900 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_26126_1124# 0.121f
C2901 a_5385_1059# LD 1.1e-19
C2902 p2_gen_magic_0.xnor_magic_4.OUT a_11708_n2115# 0.0456f
C2903 a_23352_n5390# D2_1 0.0113f
C2904 a_1209_7469# a_1209_6275# 0.00638f
C2905 a_32616_n1264# VDD 0.97f
C2906 a_5185_2253# a_5185_1059# 0.00638f
C2907 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A Q1 9.62e-19
C2908 a_13553_n6613# D2_3 8.12e-19
C2909 a_1409_8579# CLK 0.0097f
C2910 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5036_n3597# 6.98e-21
C2911 divide_by_2_1.tg_magic_3.CLK mux_magic_0.OR_magic_0.A 0.00129f
C2912 p2_gen_magic_0.xnor_magic_5.OUT p2_gen_magic_0.xnor_magic_6.OUT 0.981f
C2913 p2_gen_magic_0.xnor_magic_1.OUT a_1541_n3597# 0.368f
C2914 a_16386_n3644# VDD 0.0248f
C2915 p2_gen_magic_0.xnor_magic_3.OUT D2_4 0.193f
C2916 7b_counter_0.MDFF_0.tspc2_magic_0.D a_4235_3947# 0.278f
C2917 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A D2_2 5.7e-19
C2918 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT Q3 0.00576f
C2919 a_2749_7308# a_2749_5900# 0.475f
C2920 a_32616_n1264# D2_1 3.96e-19
C2921 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 0.0207f
C2922 7b_counter_0.3_inp_AND_magic_0.C Q6 2.08e-22
C2923 a_19841_4557# a_21381_4932# 7.98e-19
C2924 a_1541_n7648# a_1541_n8095# 0.00457f
C2925 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.3_inp_AND_magic_0.B 0.0103f
C2926 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5054_n5540# 0.0558f
C2927 a_11292_n6613# p3_gen_magic_0.3_inp_AND_magic_0.A 0.116f
C2928 p3_gen_magic_0.xnor_magic_0.OUT a_13353_n6613# 1.73e-20
C2929 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B 0.0047f
C2930 a_16386_n3644# D2_1 0.0231f
C2931 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN 0.0107f
C2932 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_3.IN 0.779f
C2933 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_1.IN 0.316f
C2934 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 7b_counter_0.MDFF_6.tspc2_magic_0.D 0.412f
C2935 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B Q4 0.00109f
C2936 DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD 1.08f
C2937 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B 0.178f
C2938 a_8411_8536# D2_2 0.298f
C2939 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A a_20041_9774# 0.0292f
C2940 a_15865_8580# a_15865_7470# 0.00329f
C2941 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_1209_3363# 4.8e-20
C2942 a_8411_9730# 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A 0.251f
C2943 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1559_n1526# 0.0629f
C2944 p2_gen_magic_0.xnor_magic_3.OUT Q2 0.863f
C2945 a_8643_n1973# a_9059_n1973# 5.82e-19
C2946 p2_gen_magic_0.3_inp_AND_magic_0.C D2_3 0.295f
C2947 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_11191_684# 0.173f
C2948 a_1957_n7648# Q7 2.48e-20
C2949 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A a_6725_684# 0.397f
C2950 a_1409_1059# Q7 0.01f
C2951 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A 0.00108f
C2952 mux_magic_0.IN2 divide_by_2_0.tg_magic_2.IN 0.289f
C2953 a_4496_9609# a_5185_7469# 3.03e-19
C2954 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT a_5036_n8579# 0.0846f
C2955 p2_gen_magic_0.xnor_magic_5.OUT VDD 1.98f
C2956 a_18891_6886# Q6 3.53e-20
C2957 p2_gen_magic_0.AND2_magic_1.A p3_gen_magic_0.3_inp_AND_magic_0.B 2.73e-20
C2958 p2_gen_magic_0.xnor_magic_5.OUT D2_1 1.51f
C2959 a_8713_1625# Q3 8.58e-20
C2960 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A D2_6 0.00237f
C2961 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B 7b_counter_0.MDFF_3.tspc2_magic_0.Q 4.47e-20
C2962 a_15865_9774# a_15865_8580# 0.00638f
C2963 a_11708_n6613# p3_gen_magic_0.xnor_magic_6.OUT 0.00656f
C2964 a_5036_n7648# D2_3 1.85e-19
C2965 a_13553_n2115# Q4 0.00847f
C2966 mux_magic_0.AND2_magic_0.A P2 0.00993f
C2967 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT P2 1.48e-19
C2968 7b_counter_0.3_inp_AND_magic_0.C a_22991_5815# 0.0191f
C2969 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B VDD 1.2f
C2970 a_5185_1059# VDD 0.994f
C2971 a_8411_9730# CLK 6.58e-19
C2972 p2_gen_magic_0.xnor_magic_6.OUT a_14756_n3644# 0.12f
C2973 p3_gen_magic_0.xnor_magic_3.OUT D2_5 0.125f
C2974 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A a_27778_1059# 9.27e-19
C2975 divide_by_2_1.tg_magic_3.CLK divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT 1.31f
C2976 7b_counter_0.MDFF_0.tspc2_magic_0.CLK Q6 0.0233f
C2977 a_16065_4557# Q1 6.2e-19
C2978 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A a_8411_8536# 1.03e-19
C2979 a_8939_n3150# Q1 0.00635f
C2980 a_5185_7469# a_6725_5900# 1.14e-19
C2981 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A 1.1e-20
C2982 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A a_20041_8580# 1.77e-19
C2983 a_21381_3524# Q4 0.00462f
C2984 a_22150_1124# a_23258_552# 7.16e-20
C2985 a_15865_1059# p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK 0.0033f
C2986 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B a_8411_3319# 0.125f
C2987 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 1.09f
C2988 a_27778_2253# D2_4 0.0401f
C2989 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_1.OUT 1.62e-19
C2990 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A Q5 0.0236f
C2991 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.149f
C2992 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A CLK 0.0214f
C2993 DFF_magic_0.tg_magic_3.CLK DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 1.84e-19
C2994 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK D2_6 0.294f
C2995 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q7 0.117f
C2996 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A D2_5 1.39e-19
C2997 a_5185_1059# LD 3.96e-19
C2998 p2_gen_magic_0.xnor_magic_4.OUT a_11492_n2115# 0.104f
C2999 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A VDD 1.32f
C3000 mux_magic_0.AND2_magic_0.A VDD 1.3f
C3001 a_20041_8580# a_19152_6440# 5.39e-19
C3002 OR_magic_2.A a_23352_n5390# 0.38f
C3003 DFF_magic_0.tg_magic_2.OUT DFF_magic_0.tg_magic_2.IN 0.965f
C3004 a_11708_n6613# D2_3 0.00184f
C3005 a_19307_1669# a_20171_1669# 0.00862f
C3006 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A D2_1 0.016f
C3007 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD 1.1f
C3008 a_8411_8536# CLK 0.0192f
C3009 7b_counter_0.MDFF_4.LD a_8713_1625# 0.00664f
C3010 a_14756_n3644# VDD 0.0501f
C3011 a_1541_n3150# a_1541_n3597# 0.0142f
C3012 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B a_12387_3319# 0.125f
C3013 p2_gen_magic_0.xnor_magic_6.OUT D2_6 0.217f
C3014 p2_gen_magic_0.AND2_magic_1.A D2_5 0.27f
C3015 7b_counter_0.MDFF_0.tspc2_magic_0.D a_4496_4877# 0.103f
C3016 a_2749_3524# a_4235_3947# 0.00212f
C3017 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A a_11279_8697# 2.4e-20
C3018 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A D2_4 0.00666f
C3019 mux_magic_0.AND2_magic_0.A D2_1 0.402f
C3020 a_19841_4557# D2_3 5.4e-19
C3021 a_11292_n2115# p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.011f
C3022 p3_gen_magic_0.xnor_magic_1.OUT a_8939_n7648# 6.88e-19
C3023 p3_gen_magic_0.xnor_magic_5.OUT a_5452_n7648# 0.0629f
C3024 p3_gen_magic_0.xnor_magic_3.OUT D2_7 0.37f
C3025 p2_gen_magic_0.xnor_magic_1.OUT Q4 0.185f
C3026 divide_by_2_0.tg_magic_3.OUT a_23352_n6798# 1.86e-20
C3027 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A a_17405_5901# 0.397f
C3028 mux_magic_0.IN1 a_32616_n1264# 0.391f
C3029 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B Q7 0.00721f
C3030 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A VDD 1.4f
C3031 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A LD 7.66e-19
C3032 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A D2_6 0.107f
C3033 OR_magic_1.VOUT divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT 1.33f
C3034 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A VDD 1.33f
C3035 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 1.59e-20
C3036 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT Q4 8.15e-19
C3037 a_12590_n7648# Q4 0.00106f
C3038 a_5054_n1526# p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT 7.12e-21
C3039 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT D2_7 0.0374f
C3040 a_23258_1746# D2_4 0.224f
C3041 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_5515_9163# 5.37e-19
C3042 a_15865_8580# CLK 0.247f
C3043 a_5185_1059# Q3 2.83e-19
C3044 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 5.61e-19
C3045 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT a_5036_n4081# 0.0846f
C3046 OR_magic_2.A DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 7.82e-19
C3047 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A D2_7 0.106f
C3048 a_1209_1059# Q7 0.0442f
C3049 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B a_21381_4932# 0.173f
C3050 VDD D2_6 6.14f
C3051 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 0.0285f
C3052 a_5036_n3150# VDD 0.0414f
C3053 p2_gen_magic_0.xnor_magic_4.OUT D2_5 0.0974f
C3054 a_16186_n3644# p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK 2.71e-20
C3055 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A LD 0.4f
C3056 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_6.OUT 0.246f
C3057 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT Q5 0.00576f
C3058 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 0.0338f
C3059 a_11292_n6613# p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 0.00128f
C3060 a_12931_7470# 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 5.46e-20
C3061 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A a_20041_9774# 8.53e-19
C3062 D2_1 D2_6 0.257f
C3063 DFF_magic_0.tg_magic_0.IN VDD 1.18f
C3064 p2_gen_magic_0.xnor_magic_6.OUT D2_2 0.2f
C3065 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT D2_3 6.64e-19
C3066 a_11492_n6613# p3_gen_magic_0.xnor_magic_6.OUT 0.00991f
C3067 a_12387_8536# D2_2 0.0119f
C3068 a_20171_1669# Q5 5.94e-20
C3069 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 0.402f
C3070 a_11708_n2115# Q4 0.00854f
C3071 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A a_1409_9773# 0.0285f
C3072 a_8713_6842# a_9689_6886# 0.235f
C3073 p3_gen_magic_0.xnor_magic_0.OUT a_11708_n6613# 0.0247f
C3074 a_12387_1746# 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A 1.03e-19
C3075 a_15865_7470# VDD 0.884f
C3076 a_9212_739# Q1 0.00797f
C3077 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B a_17405_10149# 0.173f
C3078 a_15865_6276# D2_3 0.00228f
C3079 p2_gen_magic_0.3_inp_AND_magic_0.C p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT 0.00958f
C3080 a_1209_9773# CLK 6.34e-19
C3081 p2_gen_magic_0.3_inp_AND_magic_0.C p2_gen_magic_0.3_inp_AND_magic_0.VOUT 0.792f
C3082 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT 5.61e-19
C3083 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A D2_2 0.00272f
C3084 p3_gen_magic_0.xnor_magic_6.OUT a_14556_n8142# 0.228f
C3085 LD D2_6 0.0169f
C3086 a_15865_7470# D2_1 0.237f
C3087 p3_gen_magic_0.xnor_magic_1.B Q6 0.0388f
C3088 7b_counter_0.MDFF_7.tspc2_magic_0.Q a_23802_1059# 0.12f
C3089 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A 9.4e-20
C3090 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.3_inp_AND_magic_0.B 9.01e-19
C3091 7b_counter_0.3_inp_AND_magic_0.B Q4 0.00157f
C3092 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.3_inp_AND_magic_0.A 0.00329f
C3093 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_1.OUT 0.00178f
C3094 a_20171_1669# D2_4 0.00149f
C3095 a_17405_8741# a_15865_8580# 0.00114f
C3096 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A CLK 0.00322f
C3097 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A 0.00315f
C3098 7b_counter_0.MDFF_3.tspc2_magic_0.CLK D2_7 0.0658f
C3099 a_19841_3363# CLK 0.00133f
C3100 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT DFF_magic_0.tg_magic_3.OUT 0.163f
C3101 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B 0.00121f
C3102 a_12931_2253# 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A 0.00103f
C3103 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A a_12387_8536# 0.00184f
C3104 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A a_16065_9774# 9.27e-19
C3105 a_15865_9774# VDD 0.983f
C3106 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A 0.178f
C3107 a_11279_1124# a_9412_739# 1.39e-20
C3108 VDD D2_2 4.21f
C3109 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A 0.00108f
C3110 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8643_n6024# 0.0827f
C3111 a_8713_6842# Q7 0.00548f
C3112 p2_gen_magic_0.xnor_magic_4.OUT D2_7 0.334f
C3113 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A Q3 0.0809f
C3114 a_9212_5956# 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 6.3e-20
C3115 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A a_17405_5901# 3.58e-20
C3116 a_11492_n6613# D2_3 8.12e-19
C3117 a_15865_9774# D2_1 0.00337f
C3118 D2_2 D2_1 0.117f
C3119 a_8523_n3150# D2_6 0.121f
C3120 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD 1.1f
C3121 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A a_11191_10149# 3.58e-20
C3122 a_16186_n3644# VDD 0.882f
C3123 p2_gen_magic_0.xnor_magic_5.OUT a_5452_n3150# 0.0629f
C3124 a_2749_3524# a_4496_4877# 1.39e-20
C3125 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B CLK 0.00638f
C3126 p2_gen_magic_0.xnor_magic_0.OUT a_8523_n3597# 0.0118f
C3127 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8523_n7648# 1.55e-19
C3128 7b_counter_0.MDFF_6.tspc2_magic_0.D Q1 3.55e-19
C3129 a_5036_n7648# a_5452_n7648# 0.00222f
C3130 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT a_5036_n8095# 0.0834f
C3131 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A a_1209_8579# 0.00184f
C3132 DFF_magic_0.D 7b_counter_0.DFF_magic_0.tg_magic_1.IN 0.0132f
C3133 mux_magic_0.IN1 mux_magic_0.AND2_magic_0.A 0.479f
C3134 a_16186_n3644# D2_1 0.018f
C3135 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK CLK 0.847f
C3136 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 0.228f
C3137 OR_magic_2.A mux_magic_0.AND2_magic_0.A 0.00321f
C3138 Q3 D2_6 0.28f
C3139 7b_counter_0.MDFF_5.tspc2_magic_0.Q Q2 0.29f
C3140 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A VDD 1.22f
C3141 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT OR_magic_2.A 0.00636f
C3142 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A a_13353_n2115# 1.33e-19
C3143 a_15865_9774# LD 6.64e-19
C3144 a_9212_5956# VDD 0.969f
C3145 a_1209_3363# a_1209_2253# 0.00329f
C3146 LD D2_2 0.0153f
C3147 a_19152_739# VDD 0.721f
C3148 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_6 1.86e-19
C3149 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A a_21381_8741# 2.4e-20
C3150 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_9412_739# 0.35f
C3151 7b_counter_0.MDFF_4.LD 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.00313f
C3152 a_12387_8536# a_12387_6963# 0.00329f
C3153 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A VDD 1.23f
C3154 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT CLK 1.31f
C3155 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT P2 6.97e-20
C3156 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A a_12931_9774# 0.0292f
C3157 a_8643_n6024# p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 1.86e-20
C3158 a_17405_2092# D2_3 0.0419f
C3159 CLK P2 0.153f
C3160 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_3.tspc2_magic_0.D 8.78e-21
C3161 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A a_16065_1059# 0.0292f
C3162 p2_gen_magic_0.xnor_magic_6.OUT CLK 9.29e-19
C3163 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B a_17405_2092# 0.412f
C3164 a_4235_9163# a_5515_9163# 0.00652f
C3165 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_4651_9163# 0.00409f
C3166 a_12387_8536# CLK 0.243f
C3167 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A VDD 1.32f
C3168 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B D2_3 0.00118f
C3169 a_12387_1746# a_11191_684# 1.14e-19
C3170 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A D2_1 3.01e-19
C3171 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_6.OUT 0.233f
C3172 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B D2_7 0.00118f
C3173 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A D2_1 4.06e-19
C3174 a_19152_6440# VDD 0.76f
C3175 a_1957_n3150# VDD 0.0018f
C3176 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 0.402f
C3177 p2_gen_magic_0.xnor_magic_3.OUT a_1559_n1042# 0.454f
C3178 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A LD 5.51e-19
C3179 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT a_8523_n7648# 0.0115f
C3180 a_1409_6275# Q6 0.13f
C3181 a_1209_8579# a_1409_8579# 0.298f
C3182 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 1.42e-19
C3183 DFF_magic_0.tg_magic_3.CLK DFF_magic_0.tg_magic_1.IN 0.0617f
C3184 a_19152_6440# D2_1 4.14e-19
C3185 a_1957_n3150# D2_1 0.00157f
C3186 a_4496_4393# Q6 0.0379f
C3187 a_1541_n3597# D2_7 0.00213f
C3188 a_8523_n3150# D2_2 5.07e-19
C3189 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A LD 5.51e-19
C3190 a_17405_7309# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B 1e-20
C3191 a_5054_n5540# D2_3 0.011f
C3192 a_11279_8697# a_12387_8536# 0.00114f
C3193 a_11492_n2115# Q4 0.00957f
C3194 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT D2_6 6.9e-19
C3195 p3_gen_magic_0.xnor_magic_0.OUT a_11492_n6613# 0.0655f
C3196 a_8713_6842# a_8825_6886# 0.0292f
C3197 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A LD 7.66e-19
C3198 a_12387_6963# VDD 0.87f
C3199 p3_gen_magic_0.3_inp_AND_magic_0.B Q4 0.0907f
C3200 a_11279_6341# a_9689_6886# 2.12e-20
C3201 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT a_1559_n5540# 7.56e-21
C3202 p2_gen_magic_0.xnor_magic_6.OUT a_14556_n3644# 0.228f
C3203 p2_gen_magic_0.3_inp_AND_magic_0.C a_13353_n2115# 0.556f
C3204 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 7b_counter_0.DFF_magic_0.tg_magic_2.IN 0.965f
C3205 7b_counter_0.MDFF_4.LD D2_6 1.12f
C3206 D2_2 Q3 0.109f
C3207 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT Q1 0.00991f
C3208 a_6725_684# Q5 0.0185f
C3209 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD 1.09f
C3210 p3_gen_magic_0.xnor_magic_6.OUT a_12174_n8095# 0.0235f
C3211 VDD CLK 39.2f
C3212 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5036_n8095# 9.93e-20
C3213 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_2 0.998f
C3214 7b_counter_0.MDFF_6.tspc2_magic_0.CLK D2_3 0.493f
C3215 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B Q7 0.0376f
C3216 p2_gen_magic_0.xnor_magic_4.OUT a_8643_n1042# 0.384f
C3217 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A a_27778_3363# 0.00103f
C3218 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT Q3 0.0247f
C3219 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT VDD 1.17f
C3220 CLK D2_1 1.82f
C3221 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A Q1 0.00225f
C3222 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_11292_n2115# 1.28e-19
C3223 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_5.OUT 0.149f
C3224 a_19307_1669# D2_4 6.91e-19
C3225 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_5.OUT 0.00989f
C3226 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A Q7 0.0212f
C3227 p3_gen_magic_0.xnor_magic_4.OUT a_11292_n6613# 0.315f
C3228 OR_magic_2.VOUT VDD 7.52f
C3229 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B 0.178f
C3230 a_27778_4557# CLK 3.73e-20
C3231 OR_magic_1.VOUT divide_by_2_1.tg_magic_1.IN 0.682f
C3232 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q7 0.675f
C3233 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT D2_1 4.09e-19
C3234 p2_gen_magic_0.xnor_magic_4.OUT a_8643_n1973# 7.33e-19
C3235 a_6725_684# D2_4 0.00736f
C3236 a_11279_8697# VDD 0.929f
C3237 a_1409_2253# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A 1.77e-19
C3238 OR_magic_2.VOUT D2_1 0.126f
C3239 7b_counter_0.MDFF_5.tspc2_magic_0.Q a_8955_8580# 0.017f
C3240 a_2749_5900# Q7 0.00294f
C3241 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A a_27234_552# 0.128f
C3242 LD CLK 0.634f
C3243 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_0.IN 0.287f
C3244 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_5185_2253# 4.65e-19
C3245 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_3.OUT 2.4e-19
C3246 p3_gen_magic_0.xnor_magic_1.OUT Q6 4.67e-19
C3247 7b_counter_0.MDFF_5.tspc2_magic_0.D a_8713_6842# 0.0368f
C3248 7b_counter_0.DFF_magic_0.Q D2_4 0.113f
C3249 a_14556_n3644# VDD 0.955f
C3250 a_5036_n3150# a_5452_n3150# 0.00222f
C3251 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT a_5036_n3597# 0.0828f
C3252 a_12174_n3150# D2_5 0.0576f
C3253 7b_counter_0.DFF_magic_0.Q 7b_counter_0.3_inp_AND_magic_0.A 0.00206f
C3254 a_11292_n2115# D2_3 1.74e-19
C3255 a_15865_2253# a_17405_2092# 0.00114f
C3256 7b_counter_0.3_inp_AND_magic_0.C VDD 1.46f
C3257 7b_counter_0.MDFF_5.tspc2_magic_0.Q 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 0.00482f
C3258 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A Q2 0.00108f
C3259 7b_counter_0.MDFF_1.tspc2_magic_0.Q 7b_counter_0.MDFF_1.tspc2_magic_0.CLK 0.00351f
C3260 7b_counter_0.MDFF_6.tspc2_magic_0.D a_19307_6886# 0.00451f
C3261 a_5036_n3597# Q6 0.0836f
C3262 a_11279_1124# a_8713_1625# 6.34e-20
C3263 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 8.78e-21
C3264 Q4 D2_5 0.298f
C3265 a_5515_3947# a_5385_2253# 0.00565f
C3266 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT Q6 0.00395f
C3267 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN 5.37e-19
C3268 a_14556_n3644# D2_1 6.98e-19
C3269 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B a_2749_3524# 1.01e-20
C3270 a_8523_n8579# D2_6 0.0172f
C3271 7b_counter_0.MDFF_4.LD D2_2 0.0327f
C3272 a_17405_8741# VDD 0.929f
C3273 a_17405_7309# VDD 0.936f
C3274 a_16065_1059# VDD 0.0609f
C3275 7b_counter_0.DFF_magic_0.tg_magic_0.IN 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 4.89e-20
C3276 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B a_4235_9163# 7.16e-19
C3277 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A Q5 8.66e-19
C3278 7b_counter_0.DFF_magic_0.Q Q2 1.69e-19
C3279 a_17405_8741# D2_1 0.0352f
C3280 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.258f
C3281 a_17405_7309# D2_1 0.0464f
C3282 7b_counter_0.MDFF_4.LD p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 5.15e-19
C3283 DFF_magic_0.D DFF_magic_0.tg_magic_3.OUT 0.822f
C3284 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A a_2749_8740# 2.4e-20
C3285 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A a_15865_1059# 0.251f
C3286 a_4235_9163# a_4651_9163# 0.153f
C3287 7b_counter_0.3_inp_AND_magic_0.C LD 0.0551f
C3288 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q5 0.24f
C3289 p3_gen_magic_0.3_inp_AND_magic_0.C p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK 0.00927f
C3290 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT Q4 0.0133f
C3291 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A a_7215_4932# 0.397f
C3292 Q5 D2_4 0.587f
C3293 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT CLK 0.00733f
C3294 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT a_8523_n3150# 0.00463f
C3295 a_8643_n6024# a_9059_n6471# 0.0115f
C3296 7b_counter_0.3_inp_AND_magic_0.A Q5 0.256f
C3297 a_5385_7469# D2_7 0.119f
C3298 p2_gen_magic_0.3_inp_AND_magic_0.A Q4 0.0404f
C3299 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT Q3 0.0249f
C3300 a_18891_6886# VDD 0.97f
C3301 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_8713_1625# 0.51f
C3302 Q1 Q7 0.168f
C3303 CLK Q3 0.832f
C3304 a_1209_6275# Q6 0.266f
C3305 7b_counter_0.MDFF_5.tspc2_magic_0.D a_12387_5769# 1.63e-20
C3306 a_1209_7469# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B 0.125f
C3307 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A VDD 1.24f
C3308 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A a_21381_8741# 0.0334f
C3309 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B VDD 1.2f
C3310 a_18891_6886# D2_1 0.0289f
C3311 p2_gen_magic_0.xnor_magic_6.OUT p3_gen_magic_0.3_inp_AND_magic_0.C 1.04e-19
C3312 a_5515_9163# Q7 2.48e-19
C3313 a_11191_10149# a_12387_8536# 1.14e-19
C3314 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.B 0.933f
C3315 a_5470_n6471# a_5036_n8095# 1.26e-19
C3316 a_12387_3319# D2_6 4e-19
C3317 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 2.76e-19
C3318 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1975_n1973# 0.00157f
C3319 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT a_8643_n5540# 9.33e-20
C3320 7b_counter_0.MDFF_0.tspc2_magic_0.CLK VDD 2.44f
C3321 p3_gen_magic_0.xnor_magic_0.OUT a_9059_n6471# 0.0762f
C3322 7b_counter_0.MDFF_7.tspc2_magic_0.D CLK 1.54e-19
C3323 Q2 Q5 0.61f
C3324 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A 0.178f
C3325 D2_7 Q4 0.32f
C3326 p2_gen_magic_0.xnor_magic_6.OUT a_12174_n3597# 0.0235f
C3327 7b_counter_0.3_inp_AND_magic_0.A D2_4 0.013f
C3328 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_6.tspc2_magic_0.Q 0.255f
C3329 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT 3.44e-20
C3330 a_21381_4932# Q1 0.0505f
C3331 p3_gen_magic_0.xnor_magic_6.OUT a_8523_n8095# 0.368f
C3332 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN VDD 1.25f
C3333 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A D2_6 0.00229f
C3334 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_5.OUT 0.146f
C3335 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT D2_5 0.139f
C3336 a_2749_3524# 7b_counter_0.MDFF_0.tspc2_magic_0.D 0.123f
C3337 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A 8.78e-21
C3338 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B LD 0.0047f
C3339 a_17405_684# D2_4 0.0167f
C3340 7b_counter_0.3_inp_AND_magic_0.C Q3 0.262f
C3341 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_7303_8697# 0.001f
C3342 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT D2_6 0.0457f
C3343 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN D2_1 0.046f
C3344 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT a_5036_n7648# 0.102f
C3345 a_12931_9774# a_12387_8536# 0.00308f
C3346 a_15865_3363# CLK 0.242f
C3347 Q2 D2_4 0.616f
C3348 OR_magic_2.A CLK 0.516f
C3349 7b_counter_0.MDFF_0.tspc2_magic_0.CLK LD 0.0847f
C3350 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B Q7 0.00698f
C3351 7b_counter_0.3_inp_AND_magic_0.A Q2 0.001f
C3352 a_1209_2253# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A 0.00184f
C3353 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.258f
C3354 a_11191_10149# VDD 1.55f
C3355 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B Q6 3.81e-19
C3356 p3_gen_magic_0.3_inp_AND_magic_0.C VDD 2.51f
C3357 7b_counter_0.MDFF_0.tspc2_magic_0.Q Q6 0.289f
C3358 a_1541_n8095# Q5 7.64e-19
C3359 7b_counter_0.MDFF_4.LD p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 5.14e-19
C3360 7b_counter_0.MDFF_4.LD CLK 1.5f
C3361 a_8411_3319# a_8713_1625# 3.03e-19
C3362 a_6725_7308# Q7 0.165f
C3363 7b_counter_0.MDFF_3.QB CLK 0.00694f
C3364 DFF_magic_0.D 7b_counter_0.DFF_magic_0.tg_magic_2.IN 0.011f
C3365 a_26126_1124# a_27234_552# 7.16e-20
C3366 7b_counter_0.MDFF_4.tspc2_magic_0.D a_9689_1669# 0.00451f
C3367 a_1541_n7648# Q6 0.00128f
C3368 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK 1.34f
C3369 p3_gen_magic_0.3_inp_AND_magic_0.C D2_1 0.281f
C3370 a_11279_6341# 7b_counter_0.MDFF_5.tspc2_magic_0.D 0.123f
C3371 OR_magic_2.A OR_magic_2.VOUT 0.00267f
C3372 a_12174_n3597# VDD 0.181f
C3373 a_8939_n3150# D2_5 7.68e-20
C3374 divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT VDD 1.09f
C3375 p2_gen_magic_0.3_inp_AND_magic_0.A p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 3.27e-20
C3376 a_12387_3319# D2_2 0.0108f
C3377 a_7303_3480# a_8411_3319# 0.00114f
C3378 7b_counter_0.MDFF_6.tspc2_magic_0.D a_17405_5901# 1.08e-19
C3379 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.xnor_magic_1.B 2.99e-20
C3380 a_1209_9773# a_1209_8579# 0.00638f
C3381 a_6725_2092# a_8713_1625# 0.00153f
C3382 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B a_2749_4932# 4.23e-19
C3383 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT a_1541_n8095# 0.0828f
C3384 a_8523_n4081# p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 9.33e-20
C3385 a_1541_n8095# D2_4 5.31e-19
C3386 a_12931_9774# VDD 0.0559f
C3387 p3_gen_magic_0.xnor_magic_6.OUT Q1 1.36e-19
C3388 a_15865_1059# VDD 0.984f
C3389 a_7303_3480# a_6725_2092# 1.63e-19
C3390 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B a_4496_10093# 1.29e-19
C3391 a_12387_4513# Q5 0.223f
C3392 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A D2_2 0.0148f
C3393 a_32816_n1264# a_32816_n2458# 0.0206f
C3394 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B Q3 2.49e-19
C3395 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A a_8955_4557# 0.0292f
C3396 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A a_12931_6276# 0.0292f
C3397 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A a_2749_10148# 3.58e-20
C3398 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 2.31e-19
C3399 a_4496_10093# a_4651_9163# 0.00164f
C3400 p2_gen_magic_0.3_inp_AND_magic_0.B p2_gen_magic_0.xnor_magic_6.OUT 0.197f
C3401 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 6.36e-20
C3402 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A Q5 0.00211f
C3403 a_23802_2253# 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 5.46e-20
C3404 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A 0.0224f
C3405 a_21381_8741# 7b_counter_0.3_inp_AND_magic_0.C 7.58e-20
C3406 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT a_1541_n3597# 0.0629f
C3407 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B Q1 0.00937f
C3408 a_8643_n6024# a_8643_n6471# 0.0137f
C3409 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT a_16186_n3644# 8.76e-20
C3410 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A Q5 5.18e-19
C3411 a_2749_7308# D2_7 0.0363f
C3412 a_11191_5901# VDD 1.55f
C3413 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 1.37f
C3414 a_21381_3524# Q7 0.00105f
C3415 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT divide_by_2_0.tg_magic_1.IN 4.63e-20
C3416 7b_counter_0.MDFF_4.LD a_16065_1059# 0.00329f
C3417 a_13769_n2115# D2_3 0.00843f
C3418 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.xnor_magic_3.OUT 0.0455f
C3419 a_20041_3363# D2_3 0.119f
C3420 p2_gen_magic_0.xnor_magic_3.OUT Q6 0.0455f
C3421 a_1209_7469# a_1409_7469# 0.298f
C3422 a_8955_4557# VDD 0.0935f
C3423 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.3_inp_AND_magic_0.VOUT 1.99e-23
C3424 a_16065_4557# a_16065_3363# 0.0206f
C3425 a_1409_2253# VDD 0.0124f
C3426 a_4651_9163# Q7 1.15e-19
C3427 DFF_magic_0.D a_27778_2253# 0.00228f
C3428 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B a_7215_10149# 0.173f
C3429 a_8643_n6471# a_8523_n7648# 0.186f
C3430 a_5054_n6471# a_5036_n8095# 2.84e-19
C3431 a_8825_1669# a_9689_1669# 0.00862f
C3432 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A 0.178f
C3433 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1559_n1973# 0.0115f
C3434 7b_counter_0.MDFF_1.tspc2_magic_0.CLK 7b_counter_0.MDFF_1.tspc2_magic_0.D 0.423f
C3435 p3_gen_magic_0.xnor_magic_0.OUT a_8643_n6471# 0.291f
C3436 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A D2_4 0.0202f
C3437 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B a_22150_1124# 0.412f
C3438 a_6725_7308# a_8825_6886# 1.36e-20
C3439 a_20171_6886# D2_3 4.33e-19
C3440 p2_gen_magic_0.xnor_magic_6.OUT a_8523_n3597# 0.368f
C3441 Q1 D2_3 1.19f
C3442 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A a_15865_3363# 0.00184f
C3443 p3_gen_magic_0.xnor_magic_1.B VDD 6.52f
C3444 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B Q1 0.00936f
C3445 7b_counter_0.MDFF_1.tspc2_magic_0.D Q4 7.41e-19
C3446 a_21381_4932# a_21381_3524# 0.475f
C3447 7b_counter_0.MDFF_7.tspc2_magic_0.Q Q4 0.207f
C3448 a_12174_n7648# p3_gen_magic_0.AND2_magic_1.A 0.0924f
C3449 a_8523_n7648# a_8523_n8095# 0.0142f
C3450 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT 0.229f
C3451 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A 0.00221f
C3452 p2_gen_magic_0.3_inp_AND_magic_0.B VDD 0.777f
C3453 a_11279_1124# D2_6 0.0425f
C3454 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT a_5036_n3150# 0.102f
C3455 p3_gen_magic_0.xnor_magic_0.OUT a_8523_n8095# 0.0118f
C3456 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q5 0.00231f
C3457 p3_gen_magic_0.xnor_magic_1.B D2_1 0.331f
C3458 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN 0.85f
C3459 7b_counter_0.DFF_magic_0.Q 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 0.00455f
C3460 a_2749_4932# 7b_counter_0.MDFF_0.tspc2_magic_0.D 1.08e-19
C3461 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A a_27234_3319# 1.03e-19
C3462 p2_gen_magic_0.3_inp_AND_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN 0.0142f
C3463 a_1409_2253# LD 0.0292f
C3464 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A a_17405_684# 0.397f
C3465 p2_gen_magic_0.xnor_magic_1.OUT Q7 0.188f
C3466 p3_gen_magic_0.P3 a_23352_n6798# 0.33f
C3467 7b_counter_0.MDFF_7.tspc2_magic_0.Q a_26126_1124# 1.23e-19
C3468 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.OUT 0.134f
C3469 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 0.00108f
C3470 a_12387_3319# CLK 0.259f
C3471 a_27234_1746# CLK 0.269f
C3472 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A a_27778_1059# 0.0292f
C3473 a_23560_3728# CLK 0.00196f
C3474 OR_magic_1.VOUT divide_by_2_1.tg_magic_3.IN 0.619f
C3475 OR_magic_2.A p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN 1.49e-19
C3476 a_5385_2253# Q7 0.00461f
C3477 a_4496_4393# a_5185_2253# 3.03e-19
C3478 a_8955_8580# Q2 5.02e-19
C3479 a_5185_7469# a_5185_6275# 0.00638f
C3480 a_4496_9609# a_5515_9163# 0.0292f
C3481 7b_counter_0.MDFF_6.tspc2_magic_0.Q 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A 0.00118f
C3482 7b_counter_0.DFF_magic_0.tg_magic_0.IN CLK 0.622f
C3483 a_4235_3947# Q6 0.0127f
C3484 a_6725_2092# a_5185_1059# 7.16e-20
C3485 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B D2_4 0.03f
C3486 a_16065_8580# CLK 0.136f
C3487 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 0.233f
C3488 a_15865_1059# Q3 2.13e-19
C3489 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A a_17405_10149# 3.58e-20
C3490 a_15865_7470# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B 0.125f
C3491 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_0.IN 0.0105f
C3492 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT D2_4 0.00131f
C3493 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN D2_6 0.1f
C3494 7b_counter_0.MDFF_5.tspc2_magic_0.CLK Q2 0.237f
C3495 7b_counter_0.MDFF_5.LD Q7 2.37f
C3496 a_8523_n3597# VDD 0.181f
C3497 a_8643_n6024# Q1 0.0849f
C3498 a_5515_3947# D2_5 4.39e-19
C3499 7b_counter_0.MDFF_4.tspc2_magic_0.CLK D2_6 0.262f
C3500 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B D2_3 4.21e-19
C3501 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK 1.31f
C3502 7b_counter_0.MDFF_0.tspc2_magic_0.Q 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A 0.255f
C3503 7b_counter_0.MDFF_3.tspc2_magic_0.Q D2_7 0.17f
C3504 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A 0.00894f
C3505 a_5036_n8095# D2_3 3.01e-19
C3506 a_12931_8580# D2_2 0.0401f
C3507 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_19152_6440# 0.0127f
C3508 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT a_30365_4922# 2.63e-19
C3509 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 0.0082f
C3510 a_8643_n1526# Q1 0.0808f
C3511 a_1209_8579# VDD 0.87f
C3512 a_8523_n7648# Q1 0.00802f
C3513 OR_magic_2.VOUT divide_by_2_0.tg_magic_3.CLK 0.569f
C3514 a_22062_684# VDD 1.59f
C3515 divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT mux_magic_0.IN1 6.97e-20
C3516 a_11279_1124# D2_2 0.044f
C3517 p3_gen_magic_0.xnor_magic_0.OUT Q1 0.143f
C3518 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q2 0.506f
C3519 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A a_12387_5769# 0.251f
C3520 a_24401_7877# Q5 4.38e-20
C3521 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_4.OUT 4.49e-20
C3522 p3_gen_magic_0.xnor_magic_3.OUT Q4 0.00214f
C3523 DFF_magic_0.tg_magic_2.OUT DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 3.44e-20
C3524 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 9.4e-20
C3525 7b_counter_0.DFF_magic_0.tg_magic_3.OUT D2_4 0.00958f
C3526 a_11292_n2115# a_13353_n2115# 6.01e-20
C3527 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.xnor_magic_1.OUT 0.00267f
C3528 7b_counter_0.MDFF_5.LD a_8955_9774# 1.1e-19
C3529 a_15865_2253# Q1 0.0156f
C3530 7b_counter_0.DFF_magic_0.Q 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 0.316f
C3531 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN 0.0105f
C3532 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A CLK 0.0234f
C3533 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p3_gen_magic_0.AND2_magic_1.A 0.25f
C3534 a_1409_6275# VDD 0.0559f
C3535 7b_counter_0.MDFF_4.LD a_15865_1059# 0.00147f
C3536 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT D2_7 0.153f
C3537 7b_counter_0.3_inp_AND_magic_0.B Q7 0.251f
C3538 a_13553_n2115# D2_3 0.00245f
C3539 a_1209_8579# LD 0.195f
C3540 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A 0.00108f
C3541 p2_gen_magic_0.3_inp_AND_magic_0.B Q3 0.00261f
C3542 a_4496_4393# VDD 1.07f
C3543 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A Q6 0.108f
C3544 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B a_15865_8580# 0.125f
C3545 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A a_12931_8580# 1.77e-19
C3546 p3_gen_magic_0.3_inp_AND_magic_0.VOUT D2_6 0.341f
C3547 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A Q5 0.00339f
C3548 p2_gen_magic_0.xnor_magic_5.OUT a_13353_n6613# 7.66e-21
C3549 a_1209_2253# VDD 0.87f
C3550 7b_counter_0.MDFF_4.tspc2_magic_0.Q p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 2.14e-20
C3551 a_21381_10149# Q7 0.0162f
C3552 a_24401_7877# D2_4 0.00564f
C3553 7b_counter_0.MDFF_4.tspc2_magic_0.CLK D2_2 0.222f
C3554 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT D2_5 4.98e-19
C3555 7b_counter_0.3_inp_AND_magic_0.A a_24401_7877# 0.0247f
C3556 a_8411_3319# D2_6 0.27f
C3557 a_6725_7308# a_6725_5900# 0.475f
C3558 a_19307_6886# D2_3 0.00338f
C3559 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT VDD 1.18f
C3560 a_8523_n3150# a_8523_n3597# 0.0142f
C3561 a_12174_n3150# p2_gen_magic_0.AND2_magic_1.A 0.0924f
C3562 7b_counter_0.MDFF_5.LD a_8825_6886# 8.29e-19
C3563 a_15865_4557# Q2 0.228f
C3564 a_16065_2253# Q1 0.00496f
C3565 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A p2_gen_magic_0.xnor_magic_3.OUT 2.11e-19
C3566 p3_gen_magic_0.xnor_magic_6.OUT a_12590_n7648# 0.00294f
C3567 a_1409_6275# LD 0.00387f
C3568 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT D2_1 4.54e-19
C3569 p2_gen_magic_0.AND2_magic_1.A Q4 0.173f
C3570 7b_counter_0.MDFF_4.LD a_8955_4557# 1.1e-19
C3571 divide_by_2_1.tg_magic_1.IN VDD 2.02f
C3572 a_2749_4932# a_2749_3524# 0.475f
C3573 a_4496_4393# LD 0.00664f
C3574 p2_gen_magic_0.3_inp_AND_magic_0.VOUT a_13769_n2115# 0.192f
C3575 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_8955_8580# 0.00751f
C3576 7b_counter_0.DFF_magic_0.tg_magic_1.IN VDD 2.03f
C3577 a_1209_2253# LD 0.195f
C3578 a_1541_n3150# Q7 0.344f
C3579 a_8713_6842# a_9412_5956# 0.0134f
C3580 a_11279_6341# 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 2.4e-20
C3581 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A p2_gen_magic_0.xnor_magic_3.OUT 1.55e-19
C3582 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT a_1541_n7648# 0.102f
C3583 p3_gen_magic_0.xnor_magic_1.B p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT 0.00129f
C3584 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_5385_7469# 0.00751f
C3585 a_30365_3514# CLK 0.0166f
C3586 a_23802_2253# CLK 0.0674f
C3587 a_1409_3363# CLK 7.14e-19
C3588 a_2749_2092# Q7 0.014f
C3589 a_19841_8580# Q2 1.92e-20
C3590 a_8939_n7648# Q5 2.48e-20
C3591 a_4496_9609# a_4651_9163# 0.235f
C3592 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_17405_8741# 0.00137f
C3593 a_4496_4877# Q6 0.0125f
C3594 a_12931_8580# CLK 0.13f
C3595 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_3.tspc2_magic_0.D 0.00171f
C3596 a_5054_n5540# a_5054_n6024# 0.0335f
C3597 p2_gen_magic_0.3_inp_AND_magic_0.C a_16386_n3644# 0.00263f
C3598 a_22062_684# Q3 0.0012f
C3599 a_1559_n6024# a_1957_n7648# 3.01e-19
C3600 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_3.OUT 7.86e-20
C3601 p3_gen_magic_0.xnor_magic_1.OUT VDD 1.62f
C3602 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN 0.321f
C3603 a_1559_n1042# D2_4 0.00889f
C3604 a_15865_7470# a_16065_7470# 0.298f
C3605 p2_gen_magic_0.xnor_magic_1.OUT D2_3 0.0611f
C3606 a_7303_8697# Q7 0.0498f
C3607 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A Q7 0.00783f
C3608 a_32616_n2458# OUT1 7.57e-20
C3609 a_5036_n3597# VDD 0.237f
C3610 7b_counter_0.MDFF_3.tspc2_magic_0.D a_4651_9163# 0.00451f
C3611 p3_gen_magic_0.xnor_magic_1.OUT D2_1 0.00238f
C3612 a_4651_3947# D2_5 0.00739f
C3613 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT VDD 1.07f
C3614 a_4235_9163# D2_7 0.0335f
C3615 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 0.00813f
C3616 DFF_magic_0.tg_magic_2.OUT mux_magic_0.AND2_magic_0.A 1.68e-20
C3617 7b_counter_0.MDFF_4.tspc2_magic_0.D Q4 0.00144f
C3618 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT 0.0182f
C3619 p2_gen_magic_0.xnor_magic_4.OUT Q4 0.0106f
C3620 a_16386_n8142# D2_6 0.0103f
C3621 a_11279_3480# Q5 0.0328f
C3622 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A 0.00108f
C3623 7b_counter_0.MDFF_5.LD D2_3 0.272f
C3624 a_12931_1059# VDD 0.0559f
C3625 a_12387_9730# Q1 0.223f
C3626 a_1559_n1042# Q2 2.48e-19
C3627 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_5185_2253# 0.0276f
C3628 7b_counter_0.3_inp_AND_magic_0.C a_23793_5904# 0.0541f
C3629 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN CLK 0.00105f
C3630 a_24185_7877# Q5 2.88e-19
C3631 a_34156_n889# a_34156_n2297# 0.475f
C3632 p2_gen_magic_0.3_inp_AND_magic_0.C p2_gen_magic_0.xnor_magic_5.OUT 0.007f
C3633 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p2_gen_magic_0.AND2_magic_1.A 0.25f
C3634 a_19152_1223# a_19152_739# 0.0141f
C3635 7b_counter_0.MDFF_5.tspc2_magic_0.Q Q6 0.0266f
C3636 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q3 0.502f
C3637 a_2749_7308# 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A 2.4e-20
C3638 a_12387_1746# Q1 0.0156f
C3639 a_12931_4557# Q5 0.12f
C3640 a_1209_6275# VDD 0.975f
C3641 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 0.0206f
C3642 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.IN 0.29f
C3643 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_1.IN 4.63e-20
C3644 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A a_17405_3524# 2.07e-19
C3645 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_9059_n1973# 6.1e-19
C3646 a_1409_4557# a_1209_3363# 0.00308f
C3647 7b_counter_0.MDFF_4.tspc2_magic_0.Q a_8713_1625# 0.0125f
C3648 a_24185_7877# D2_4 0.0032f
C3649 a_5470_n1973# D2_5 0.00214f
C3650 p3_gen_magic_0.xnor_magic_5.OUT D2_6 0.465f
C3651 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT D2_4 0.00361f
C3652 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_17405_7309# 0.412f
C3653 DFF_magic_0.tg_magic_3.OUT P2 3.51e-19
C3654 7b_counter_0.3_inp_AND_magic_0.A a_24185_7877# 0.0655f
C3655 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1559_n1526# 0.0824f
C3656 a_1559_n1973# p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT 1.81e-19
C3657 a_12387_4513# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A 0.128f
C3658 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_0.OUT 1.56e-19
C3659 a_11292_n6613# VDD 1.22f
C3660 a_17405_5901# D2_3 0.0164f
C3661 p2_gen_magic_0.xnor_magic_6.OUT a_12590_n3150# 0.00294f
C3662 a_12931_2253# Q1 0.00496f
C3663 DFF_magic_0.tg_magic_2.OUT DFF_magic_0.tg_magic_0.IN 0.0105f
C3664 p3_gen_magic_0.xnor_magic_1.OUT Q3 1.22e-20
C3665 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A 0.00108f
C3666 a_5452_n7648# a_5036_n8095# 0.013f
C3667 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT 0.195f
C3668 a_1209_6275# LD 0.00288f
C3669 a_11292_n6613# D2_1 0.0124f
C3670 7b_counter_0.DFF_magic_0.Q DFF_magic_0.D 0.849f
C3671 p3_gen_magic_0.3_inp_AND_magic_0.A p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 3.27e-20
C3672 p3_gen_magic_0.3_inp_AND_magic_0.VOUT CLK 0.329f
C3673 a_13353_n2115# a_13769_n2115# 0.278f
C3674 p2_gen_magic_0.3_inp_AND_magic_0.VOUT a_13553_n2115# 1.9e-20
C3675 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_18891_6886# 7.16e-19
C3676 Q7 D2_5 0.831f
C3677 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT Q3 5.29e-19
C3678 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A 7b_counter_0.MDFF_5.LD 1.1e-20
C3679 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B a_2749_684# 0.173f
C3680 a_11279_6341# a_9412_5956# 1.39e-20
C3681 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B CLK 0.0351f
C3682 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_2749_7308# 0.121f
C3683 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B Q1 0.00344f
C3684 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A D2_6 0.0622f
C3685 a_30365_4922# CLK 0.0127f
C3686 a_19152_1223# CLK 0.00834f
C3687 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B VDD 1.2f
C3688 7b_counter_0.MDFF_0.tspc2_magic_0.Q VDD 1.35f
C3689 divide_by_2_1.tg_magic_1.IN mux_magic_0.IN1 0.00449f
C3690 a_1409_4557# Q6 0.00399f
C3691 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B a_2749_8740# 0.412f
C3692 p2_gen_magic_0.3_inp_AND_magic_0.C a_14756_n3644# 0.00112f
C3693 a_1541_n7648# VDD 0.014f
C3694 p3_gen_magic_0.xnor_magic_4.OUT Q5 0.478f
C3695 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B D2_1 0.0224f
C3696 DFF_magic_0.tg_magic_3.OUT VDD 1.15f
C3697 a_5185_7469# 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A 1.03e-19
C3698 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B Q6 0.0123f
C3699 a_19841_9774# Q2 9.61e-19
C3700 a_8411_4513# Q7 0.00531f
C3701 7b_counter_0.MDFF_4.LD 7b_counter_0.DFF_magic_0.tg_magic_1.IN 0.00645f
C3702 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN Q4 0.00524f
C3703 a_12590_n3150# VDD 0.0018f
C3704 a_2749_8740# a_4651_9163# 2.12e-20
C3705 a_5470_n1973# D2_7 6.9e-19
C3706 p3_gen_magic_0.3_inp_AND_magic_0.B p3_gen_magic_0.xnor_magic_6.OUT 0.198f
C3707 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_6.OUT 0.0529f
C3708 a_26126_1124# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A 0.0334f
C3709 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 0.00108f
C3710 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 0.229f
C3711 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.OUT 1.91e-19
C3712 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B LD 6.07e-19
C3713 a_14756_n8142# D2_6 0.0139f
C3714 7b_counter_0.MDFF_0.tspc2_magic_0.Q LD 0.12f
C3715 a_12387_552# VDD 0.973f
C3716 p3_gen_magic_0.xnor_magic_4.OUT D2_4 0.207f
C3717 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A a_27234_552# 0.251f
C3718 a_8523_n4081# Q1 0.0072f
C3719 7b_counter_0.MDFF_0.tspc2_magic_0.D a_1209_3363# 7.57e-20
C3720 a_8411_9730# 7b_counter_0.MDFF_5.tspc2_magic_0.Q 0.223f
C3721 7b_counter_0.DFF_magic_0.tg_magic_2.IN P2 2.12e-19
C3722 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5470_n6471# 6.1e-19
C3723 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT 0.156f
C3724 a_12387_4513# a_11279_3480# 7.16e-20
C3725 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A Q6 4.53e-19
C3726 7b_counter_0.3_inp_AND_magic_0.C a_23985_7877# 0.615f
C3727 a_23207_5815# Q5 4.56e-20
C3728 D2_7 Q7 0.777f
C3729 a_12931_7470# D2_2 0.164f
C3730 p2_gen_magic_0.3_inp_AND_magic_0.C D2_6 0.0188f
C3731 DFF_magic_0.D D2_4 0.0401f
C3732 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK Q5 4.95e-19
C3733 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A 0.0175f
C3734 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_8643_n1042# 0.0802f
C3735 a_6725_684# Q6 0.0175f
C3736 a_18891_1669# a_19152_739# 0.651f
C3737 a_7303_8697# a_4496_9609# 0.00152f
C3738 a_5054_n6471# D2_5 0.0789f
C3739 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT a_12174_n7648# 0.00915f
C3740 a_12931_9774# a_12931_8580# 0.0206f
C3741 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 0.00108f
C3742 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT P2 4.95e-19
C3743 7b_counter_0.MDFF_4.LD a_12931_1059# 0.00329f
C3744 a_11292_n6613# p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.0109f
C3745 p2_gen_magic_0.xnor_magic_3.OUT VDD 2.86f
C3746 7b_counter_0.DFF_magic_0.Q Q6 1.47e-19
C3747 a_15865_4557# a_17405_3524# 7.16e-20
C3748 p3_gen_magic_0.xnor_magic_4.OUT Q2 0.128f
C3749 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A 0.00108f
C3750 p3_gen_magic_0.3_inp_AND_magic_0.B D2_3 0.00751f
C3751 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_8643_n1973# 0.102f
C3752 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A CLK 0.00433f
C3753 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 7b_counter_0.MDFF_3.tspc2_magic_0.Q 0.0189f
C3754 a_12387_4513# a_12931_4557# 0.297f
C3755 p2_gen_magic_0.xnor_magic_3.OUT D2_1 0.0282f
C3756 a_5054_n1973# D2_5 0.0756f
C3757 p3_gen_magic_0.xnor_magic_6.OUT D2_5 0.135f
C3758 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 1.56e-20
C3759 a_9212_739# a_9689_1669# 0.153f
C3760 7b_counter_0.3_inp_AND_magic_0.A a_23207_5815# 2.57e-19
C3761 divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.OUT 0.163f
C3762 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK D2_4 0.00166f
C3763 7b_counter_0.MDFF_0.tspc2_magic_0.Q Q3 3.07e-19
C3764 a_19152_6440# a_19152_5956# 0.0141f
C3765 7b_counter_0.MDFF_0.tspc2_magic_0.D Q6 0.0177f
C3766 7b_counter_0.MDFF_5.tspc2_magic_0.Q a_8411_8536# 0.0276f
C3767 a_5452_n3150# a_5036_n3597# 0.013f
C3768 7b_counter_0.DFF_magic_0.tg_magic_2.IN VDD 1.23f
C3769 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.0032f
C3770 p3_gen_magic_0.xnor_magic_1.OUT a_8523_n8579# 0.01f
C3771 mux_magic_0.OR_magic_0.B a_34156_n2297# 0.412f
C3772 a_1541_n7648# Q3 1.88e-19
C3773 DFF_magic_0.tg_magic_3.OUT Q3 3.73e-19
C3774 a_12174_n3150# Q4 0.368f
C3775 p2_gen_magic_0.xnor_magic_3.OUT LD 2.3e-19
C3776 divide_by_2_1.tg_magic_3.IN VDD 2.79f
C3777 7b_counter_0.MDFF_1.tspc2_magic_0.CLK Q4 8.64e-19
C3778 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A Q2 6.29e-19
C3779 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_6.OUT 0.2f
C3780 p2_gen_magic_0.xnor_magic_0.OUT Q5 1.2e-19
C3781 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 0.0277f
C3782 a_13353_n6613# CLK 0.00103f
C3783 a_13353_n2115# a_13553_n2115# 0.519f
C3784 a_23207_5815# Q2 0.271f
C3785 a_12387_9730# 7b_counter_0.MDFF_5.LD 0.00288f
C3786 a_7215_10149# a_7303_8697# 0.475f
C3787 a_15865_7470# a_16065_6276# 0.00308f
C3788 Q6 Q5 0.353f
C3789 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A a_7303_8697# 0.0334f
C3790 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD 1.09f
C3791 a_5185_2253# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A 0.00184f
C3792 DFF_magic_0.tg_magic_2.OUT CLK 0.287f
C3793 a_18891_1669# CLK 0.00484f
C3794 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 0.401f
C3795 a_26126_3480# CLK 9.95e-19
C3796 a_4235_3947# VDD 1.06f
C3797 a_5054_n6471# D2_7 1.85e-19
C3798 a_7215_4932# Q6 0.00283f
C3799 p2_gen_magic_0.3_inp_AND_magic_0.C a_16186_n3644# 0.126f
C3800 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B a_2749_10148# 0.173f
C3801 a_12387_552# Q3 2.57e-19
C3802 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A Q6 0.00755f
C3803 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_0.IN 0.287f
C3804 7b_counter_0.MDFF_4.tspc2_magic_0.D a_9212_739# 0.278f
C3805 a_1409_7469# Q6 0.002f
C3806 a_12387_6963# a_12931_7470# 0.293f
C3807 D2_5 D2_3 3.47f
C3808 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT D2_4 0.00486f
C3809 a_1209_4557# Q7 9.91e-19
C3810 p3_gen_magic_0.3_inp_AND_magic_0.C p3_gen_magic_0.3_inp_AND_magic_0.VOUT 0.793f
C3811 mux_magic_0.OR_magic_0.A a_32816_n1264# 9.27e-19
C3812 p2_gen_magic_0.xnor_magic_0.OUT D2_4 0.00405f
C3813 a_2749_5900# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B 4.23e-19
C3814 divide_by_2_1.tg_magic_3.CLK a_32616_n1264# 0.00207f
C3815 OR_magic_2.VOUT divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT 2.41e-19
C3816 p3_gen_magic_0.xnor_magic_6.OUT D2_7 0.00181f
C3817 a_5054_n1973# D2_7 0.496f
C3818 7b_counter_0.MDFF_1.tspc2_magic_0.Q D2_3 0.284f
C3819 Q6 D2_4 1.67f
C3820 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_1.OUT 0.00179f
C3821 a_22150_1124# 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 2.4e-20
C3822 a_11191_684# D2_2 0.0153f
C3823 a_12931_7470# CLK 0.0106f
C3824 a_1409_9773# D2_7 0.0103f
C3825 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.3_inp_AND_magic_0.A 0.00329f
C3826 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.3_inp_AND_magic_0.B 9.01e-19
C3827 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A a_17405_4932# 0.397f
C3828 OR_magic_2.A DFF_magic_0.tg_magic_3.OUT 0.00798f
C3829 a_16186_n8142# D2_6 0.0188f
C3830 7b_counter_0.MDFF_4.tspc2_magic_0.Q D2_6 0.41f
C3831 p2_gen_magic_0.xnor_magic_3.OUT Q3 1.29f
C3832 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A Q2 7.57e-19
C3833 a_27778_2253# VDD 0.0124f
C3834 7b_counter_0.MDFF_4.LD DFF_magic_0.tg_magic_3.OUT 0.00114f
C3835 a_2749_3524# a_1209_3363# 0.00114f
C3836 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5054_n6471# 0.102f
C3837 a_12387_4513# a_11191_4932# 7.98e-19
C3838 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT Q2 0.00151f
C3839 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT 0.00172f
C3840 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A D2_5 0.0167f
C3841 Q2 Q6 1.38f
C3842 p2_gen_magic_0.3_inp_AND_magic_0.A D2_3 0.0097f
C3843 a_22991_5815# Q5 2.42e-20
C3844 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.153f
C3845 a_27234_4513# CLK 3.94e-19
C3846 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT a_12174_n3150# 0.00871f
C3847 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_1.IN 1.16f
C3848 p3_gen_magic_0.xnor_magic_1.B a_1541_n8579# 0.0698f
C3849 a_17405_7309# a_19152_5956# 1.39e-20
C3850 a_8643_n6024# D2_5 0.00419f
C3851 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT a_5036_n8095# 0.0629f
C3852 7b_counter_0.MDFF_4.LD a_12387_552# 3.96e-19
C3853 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT Q4 0.646f
C3854 7b_counter_0.DFF_magic_0.Q 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B 2.36e-20
C3855 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A VDD 1.22f
C3856 p3_gen_magic_0.3_inp_AND_magic_0.C a_13769_n6613# 0.0441f
C3857 a_11708_n6613# D2_2 1.63e-20
C3858 D2_7 D2_3 0.0121f
C3859 a_24185_7877# a_24401_7877# 0.326f
C3860 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_4235_9163# 0.654f
C3861 a_5185_7469# CLK 2.95e-19
C3862 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A a_12931_1059# 9.27e-19
C3863 a_9212_739# a_8825_1669# 0.00652f
C3864 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A a_6725_684# 3.58e-20
C3865 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT D2_6 2.08e-19
C3866 a_8523_n7648# D2_5 0.0136f
C3867 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A a_11279_3480# 0.0334f
C3868 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A CLK 0.0742f
C3869 7b_counter_0.3_inp_AND_magic_0.A a_22991_5815# 8.94e-20
C3870 a_1541_n8095# Q6 1.35e-19
C3871 p2_gen_magic_0.3_inp_AND_magic_0.C CLK 0.67f
C3872 p3_gen_magic_0.xnor_magic_0.OUT D2_5 0.172f
C3873 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK 3.24e-20
C3874 a_1559_n1526# p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT 6.69e-21
C3875 a_8643_n6024# p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT 2.26e-20
C3876 a_18891_6886# a_19152_5956# 0.651f
C3877 a_11279_6341# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B 1e-20
C3878 a_2749_3524# Q6 0.0105f
C3879 p3_gen_magic_0.3_inp_AND_magic_0.C a_16386_n8142# 0.00263f
C3880 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT a_1541_n4081# 0.057f
C3881 mux_magic_0.OR_magic_0.B a_34156_n889# 0.173f
C3882 7b_counter_0.MDFF_4.tspc2_magic_0.Q D2_2 5.09e-20
C3883 a_4496_9609# D2_7 5.51e-20
C3884 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_6.OUT 0.176f
C3885 a_23258_1746# VDD 0.998f
C3886 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A LD 1.1e-20
C3887 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT 0.156f
C3888 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A D2_7 0.0869f
C3889 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT a_8523_n7648# 0.102f
C3890 p3_gen_magic_0.xnor_magic_3.OUT a_1559_n5540# 0.454f
C3891 a_19841_9774# a_19841_8580# 0.00638f
C3892 a_22991_5815# Q2 0.175f
C3893 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A a_12931_4557# 9.27e-19
C3894 7b_counter_0.MDFF_3.tspc2_magic_0.D D2_7 0.00366f
C3895 a_1209_2253# a_2749_684# 1.14e-19
C3896 7b_counter_0.DFF_magic_0.tg_magic_2.IN OR_magic_2.A 2.97e-20
C3897 a_15865_7470# a_15865_6276# 0.00638f
C3898 a_9412_739# Q1 0.00312f
C3899 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT 0.0188f
C3900 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_3 0.983f
C3901 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A a_15865_8580# 1.03e-19
C3902 a_4496_4877# VDD 0.762f
C3903 divide_by_2_1.tg_magic_3.IN mux_magic_0.IN1 0.321f
C3904 7b_counter_0.MDFF_4.LD 7b_counter_0.DFF_magic_0.tg_magic_2.IN 0.0113f
C3905 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT D2_6 0.0812f
C3906 a_8955_3363# Q5 3.88e-19
C3907 mux_magic_0.OR_magic_0.A a_32816_n2458# 1.77e-19
C3908 a_9212_5956# 7b_counter_0.MDFF_4.tspc2_magic_0.Q 6.28e-20
C3909 p2_gen_magic_0.3_inp_AND_magic_0.C a_14556_n3644# 5.23e-19
C3910 a_27778_2253# Q3 0.002f
C3911 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT a_1559_n5540# 8.17e-21
C3912 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 3.44e-20
C3913 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A Q5 5.99e-19
C3914 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q1 0.64f
C3915 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_2.IN 6.95e-19
C3916 a_1209_7469# Q6 0.00139f
C3917 a_8643_n1526# a_9059_n1973# 0.0115f
C3918 mux_magic_0.OR_magic_0.A a_34156_n2297# 0.0334f
C3919 p3_gen_magic_0.xnor_magic_3.OUT Q7 6.24e-19
C3920 p3_gen_magic_0.3_inp_AND_magic_0.C a_13353_n6613# 0.556f
C3921 divide_by_2_1.tg_magic_3.CLK mux_magic_0.AND2_magic_0.A 0.00159f
C3922 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A a_8955_3363# 1.77e-19
C3923 7b_counter_0.MDFF_7.tspc2_magic_0.Q a_23258_552# 0.223f
C3924 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT D2_2 0.0788f
C3925 p3_gen_magic_0.3_inp_AND_magic_0.C p3_gen_magic_0.xnor_magic_5.OUT 0.007f
C3926 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT 0.0032f
C3927 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.101f
C3928 a_19152_6440# a_19841_4557# 1.73e-19
C3929 DFF_magic_0.D 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 0.0196f
C3930 p3_gen_magic_0.xnor_magic_4.OUT a_8643_n5540# 0.384f
C3931 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_5385_7469# 0.017f
C3932 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT VDD 1.04f
C3933 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B Q1 0.00762f
C3934 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A Q6 0.0039f
C3935 a_14556_n8142# D2_6 0.0635f
C3936 a_32616_n1264# OUT1 1.63e-20
C3937 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A Q5 2.57e-19
C3938 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT Q7 0.00753f
C3939 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_1 4.19e-19
C3940 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A Q3 2.56e-19
C3941 a_8411_9730# Q2 0.00105f
C3942 a_26038_684# a_27234_552# 7.98e-19
C3943 a_23258_552# a_23802_1059# 0.297f
C3944 7b_counter_0.MDFF_5.tspc2_magic_0.CLK Q6 1.99e-20
C3945 a_20171_1669# VDD 0.075f
C3946 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 0.00315f
C3947 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A D2_4 0.00103f
C3948 a_2749_4932# a_1209_3363# 1.14e-19
C3949 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B Q2 0.00107f
C3950 7b_counter_0.MDFF_5.tspc2_magic_0.Q VDD 1.22f
C3951 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A 0.178f
C3952 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT a_5036_n3597# 0.0629f
C3953 OR_magic_2.VOUT divide_by_2_0.tg_magic_2.IN 0.00111f
C3954 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A D2_4 0.0121f
C3955 p3_gen_magic_0.xnor_magic_1.B a_16386_n8142# 7.65e-19
C3956 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A Q2 0.00108f
C3957 7b_counter_0.MDFF_5.tspc2_magic_0.Q D2_1 3.67e-19
C3958 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 0.0357f
C3959 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT 0.00535f
C3960 7b_counter_0.MDFF_4.LD a_27778_2253# 0.0293f
C3961 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q6 0.212f
C3962 a_23258_1746# Q3 1.56e-19
C3963 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A a_1209_4557# 0.251f
C3964 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A Q2 3.98e-20
C3965 a_11492_n6613# D2_2 2.63e-20
C3966 p3_gen_magic_0.3_inp_AND_magic_0.C a_13553_n6613# 0.00138f
C3967 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_4496_10093# 0.35f
C3968 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A a_12387_552# 0.128f
C3969 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A a_11191_4932# 0.397f
C3970 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.P3 0.312f
C3971 7b_counter_0.MDFF_1.tspc2_magic_0.D D2_3 0.00366f
C3972 a_1559_n1973# a_1541_n3150# 0.191f
C3973 a_22150_1124# CLK 0.095f
C3974 p2_gen_magic_0.xnor_magic_4.OUT a_5470_n1973# 0.0761f
C3975 a_8411_8536# Q2 0.0026f
C3976 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_1.tspc2_magic_0.D 0.00171f
C3977 7b_counter_0.MDFF_5.tspc2_magic_0.Q LD 7.02e-19
C3978 DFF_magic_0.D DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 0.301f
C3979 a_12174_n4081# D2_5 0.0272f
C3980 p2_gen_magic_0.xnor_magic_1.OUT a_5036_n4081# 2.1e-19
C3981 a_2749_4932# Q6 0.0164f
C3982 p2_gen_magic_0.3_inp_AND_magic_0.A p2_gen_magic_0.3_inp_AND_magic_0.VOUT 3.5e-19
C3983 p3_gen_magic_0.3_inp_AND_magic_0.C a_14756_n8142# 0.00228f
C3984 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A Q2 2.21e-19
C3985 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT Q5 0.00718f
C3986 p3_gen_magic_0.xnor_magic_1.OUT a_1541_n8579# 0.338f
C3987 a_9212_739# Q4 1.76e-20
C3988 a_5185_2253# a_6725_684# 1.14e-19
C3989 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT a_8523_n3150# 0.102f
C3990 7b_counter_0.MDFF_3.tspc2_magic_0.CLK Q7 0.0208f
C3991 DFF_magic_0.D 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 0.0903f
C3992 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_6.OUT 0.0529f
C3993 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A p2_gen_magic_0.xnor_magic_3.OUT 0.00109f
C3994 mux_magic_0.IN2 divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT 7.64e-20
C3995 p3_gen_magic_0.xnor_magic_1.B p3_gen_magic_0.xnor_magic_5.OUT 0.851f
C3996 a_2749_8740# D2_7 0.0422f
C3997 a_6725_7308# a_5185_6275# 7.16e-20
C3998 a_1409_1059# CLK 0.00449f
C3999 a_8643_n1042# a_8643_n1526# 0.0335f
C4000 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT 0.0154f
C4001 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A a_26038_4932# 3.58e-20
C4002 a_24059_4877# CLK 0.00118f
C4003 a_1409_4557# VDD 0.0559f
C4004 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A Q5 0.00312f
C4005 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT D2_4 2.45e-19
C4006 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 0.00212f
C4007 a_17405_2092# p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 6.42e-22
C4008 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.00222f
C4009 a_19841_3363# Q5 6.21e-20
C4010 a_32816_n1264# mux_magic_0.IN2 0.00449f
C4011 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_15865_7470# 4.8e-20
C4012 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B VDD 1.2f
C4013 7b_counter_0.MDFF_4.LD a_23258_1746# 0.195f
C4014 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B Q7 0.0132f
C4015 a_5054_n1042# Q1 8.14e-20
C4016 a_8713_1625# Q1 0.0602f
C4017 a_9059_n6471# D2_6 1.05e-19
C4018 mux_magic_0.OR_magic_0.A a_34156_n889# 0.397f
C4019 a_8643_n1526# a_8643_n1973# 0.0137f
C4020 a_5452_n7648# D2_7 0.00236f
C4021 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT D2_5 1.01f
C4022 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1957_n3150# 6.85e-21
C4023 a_17405_2092# a_19152_739# 1.39e-20
C4024 a_19841_8580# Q6 1.23e-19
C4025 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_2749_7308# 0.00137f
C4026 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A D2_4 0.0236f
C4027 a_12931_6276# D2_2 0.0035f
C4028 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A p2_gen_magic_0.3_inp_AND_magic_0.B 3.97e-19
C4029 a_5185_2253# Q5 0.00146f
C4030 mux_magic_0.AND2_magic_0.A OUT1 8.78e-21
C4031 a_1409_4557# LD 0.00329f
C4032 a_8713_6842# D2_6 0.0511f
C4033 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A D2_6 2.27e-19
C4034 a_1209_9773# Q2 9.57e-19
C4035 a_11191_4932# a_11279_3480# 0.475f
C4036 a_19307_1669# VDD 0.00407f
C4037 p3_gen_magic_0.xnor_magic_3.OUT D2_3 0.135f
C4038 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A VDD 1.38f
C4039 a_15865_9774# 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 1.63e-20
C4040 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B LD 0.0047f
C4041 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A a_1409_6275# 9.27e-19
C4042 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B 0.00112f
C4043 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A 0.00112f
C4044 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A CLK 0.00315f
C4045 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 8.78e-21
C4046 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 0.00108f
C4047 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A a_17405_684# 3.58e-20
C4048 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B Q7 0.0311f
C4049 a_15865_2253# 7b_counter_0.MDFF_1.tspc2_magic_0.D 7.57e-20
C4050 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A D2_1 4.06e-19
C4051 a_6725_684# VDD 1.55f
C4052 a_13353_n2115# D2_5 4.86e-20
C4053 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_11279_6341# 0.409f
C4054 p2_gen_magic_0.3_inp_AND_magic_0.A p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT 0.00302f
C4055 a_27234_1746# a_27778_2253# 0.298f
C4056 p2_gen_magic_0.xnor_magic_6.OUT Q5 0.15f
C4057 a_8411_8536# a_8955_8580# 0.296f
C4058 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_2.IN 6.95e-19
C4059 a_17405_7309# a_15865_6276# 7.16e-20
C4060 7b_counter_0.MDFF_6.tspc2_magic_0.D 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 8.78e-21
C4061 7b_counter_0.DFF_magic_0.Q VDD 6.53f
C4062 a_1541_n3597# Q7 0.0832f
C4063 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT a_1541_n8095# 0.0627f
C4064 7b_counter_0.MDFF_4.LD a_20171_1669# 8.29e-19
C4065 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN D2_6 0.109f
C4066 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_8411_8536# 4.65e-19
C4067 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A LD 7.66e-19
C4068 a_9059_n6471# D2_2 0.00157f
C4069 a_11279_1124# a_12387_552# 7.16e-20
C4070 a_11292_n2115# D2_2 0.038f
C4071 p3_gen_magic_0.AND2_magic_1.A VDD 1.4f
C4072 p2_gen_magic_0.xnor_magic_4.OUT a_5054_n1973# 0.299f
C4073 a_17405_2092# CLK 2.46e-19
C4074 7b_counter_0.MDFF_0.tspc2_magic_0.D VDD 1.41f
C4075 a_8523_n4081# D2_5 0.00782f
C4076 p2_gen_magic_0.AND2_magic_1.A D2_3 0.109f
C4077 p2_gen_magic_0.xnor_magic_1.OUT a_1541_n4081# 0.332f
C4078 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 0.00168f
C4079 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B CLK 1.23e-19
C4080 a_12387_5769# D2_6 2.15e-20
C4081 p2_gen_magic_0.3_inp_AND_magic_0.B p2_gen_magic_0.3_inp_AND_magic_0.C 1.29f
C4082 p2_gen_magic_0.3_inp_AND_magic_0.A a_13353_n2115# 0.467f
C4083 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A a_7215_4932# 3.58e-20
C4084 a_8713_6842# D2_2 1.65e-19
C4085 p2_gen_magic_0.xnor_magic_5.OUT Q1 0.0303f
C4086 p3_gen_magic_0.3_inp_AND_magic_0.C a_16186_n8142# 0.126f
C4087 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 0.00108f
C4088 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A D2_2 0.0403f
C4089 7b_counter_0.DFF_magic_0.Q LD 0.406f
C4090 p3_gen_magic_0.xnor_magic_1.OUT a_16386_n8142# 0.132f
C4091 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A 0.00896f
C4092 7b_counter_0.DFF_magic_0.Q a_24003_10051# 0.09f
C4093 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_19152_6440# 0.509f
C4094 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT Q4 1.93e-19
C4095 divide_by_2_1.tg_magic_3.CLK CLK 0.00249f
C4096 VDD Q5 20.7f
C4097 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_4.tspc2_magic_0.D 0.00171f
C4098 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B p2_gen_magic_0.xnor_magic_4.OUT 1.05e-19
C4099 a_2749_10148# D2_7 2.25e-19
C4100 a_12387_6963# a_12931_6276# 0.00152f
C4101 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.xnor_magic_3.OUT 0.0455f
C4102 mux_magic_0.IN2 a_32816_n2458# 0.12f
C4103 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_12387_552# 1.37e-19
C4104 D2_1 Q5 0.43f
C4105 7b_counter_0.MDFF_0.tspc2_magic_0.D LD 0.00852f
C4106 a_7215_4932# VDD 1.55f
C4107 7b_counter_0.MDFF_1.tspc2_magic_0.D p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT 0.00126f
C4108 a_23560_3728# a_23258_1746# 3.03e-19
C4109 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A VDD 1.24f
C4110 a_1559_n6471# D2_7 4.09e-19
C4111 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A CLK 0.00127f
C4112 a_12931_6276# CLK 0.00519f
C4113 a_8713_6842# a_9212_5956# 0.299f
C4114 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT 2.82e-19
C4115 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A D2_2 0.00397f
C4116 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A a_19841_3363# 1.03e-19
C4117 a_1409_7469# VDD 0.0124f
C4118 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT VDD 1.17f
C4119 a_8643_n6471# D2_6 1.85e-19
C4120 VDD D2_4 7.59f
C4121 7b_counter_0.MDFF_4.tspc2_magic_0.D D2_3 5.71e-19
C4122 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A 0.00112f
C4123 p2_gen_magic_0.xnor_magic_4.OUT D2_3 0.159f
C4124 LD Q5 0.135f
C4125 7b_counter_0.3_inp_AND_magic_0.A VDD 0.464f
C4126 a_1559_n1973# D2_7 0.00377f
C4127 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT 0.153f
C4128 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN 0.694f
C4129 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A a_22062_684# 0.397f
C4130 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN a_16186_n3644# 2.1e-20
C4131 7b_counter_0.DFF_magic_0.Q 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 0.00184f
C4132 7b_counter_0.MDFF_4.tspc2_magic_0.CLK p2_gen_magic_0.xnor_magic_3.OUT 2.45e-19
C4133 p3_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_5.OUT 1.34f
C4134 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B a_19841_8580# 0.125f
C4135 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B 0.178f
C4136 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_4496_9609# 0.51f
C4137 D2_1 D2_4 0.773f
C4138 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 0.00108f
C4139 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A Q1 8.6e-19
C4140 a_12387_5769# D2_2 0.013f
C4141 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B 9.4e-20
C4142 a_27778_4557# D2_4 0.00452f
C4143 a_8523_n8095# D2_6 0.24f
C4144 a_11279_6341# D2_6 0.0229f
C4145 a_19841_9774# Q6 4.57e-19
C4146 a_17405_684# VDD 1.55f
C4147 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A a_19841_3363# 0.00184f
C4148 a_15865_9774# a_16065_9774# 0.297f
C4149 a_1409_7469# LD 0.0292f
C4150 7b_counter_0.MDFF_3.tspc2_magic_0.D 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 0.423f
C4151 7b_counter_0.MDFF_4.tspc2_magic_0.Q a_8955_4557# 0.12f
C4152 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A a_1209_6275# 0.128f
C4153 VDD Q2 9.49f
C4154 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_5 0.00449f
C4155 p3_gen_magic_0.AND2_magic_1.A a_12174_n8579# 0.613f
C4156 LD D2_4 0.112f
C4157 a_26126_1124# 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 2.4e-20
C4158 a_5385_7469# Q7 0.0146f
C4159 7b_counter_0.3_inp_AND_magic_0.A LD 0.005f
C4160 a_24003_10051# D2_4 0.00342f
C4161 mux_magic_0.OR_magic_0.A mux_magic_0.OR_magic_0.B 0.178f
C4162 Q2 D2_1 1.21f
C4163 7b_counter_0.MDFF_1.tspc2_magic_0.Q 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B 1.17e-20
C4164 a_12387_6963# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A 0.00184f
C4165 a_8523_n3150# Q5 0.303f
C4166 a_24003_10051# 7b_counter_0.3_inp_AND_magic_0.A 2.55e-20
C4167 p3_gen_magic_0.xnor_magic_1.B a_16186_n8142# 0.0015f
C4168 a_5054_n6024# D2_5 0.04f
C4169 a_8713_6842# CLK 0.0391f
C4170 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 0.00315f
C4171 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B D2_2 0.00258f
C4172 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A CLK 0.00486f
C4173 a_13769_n2115# D2_6 5.08e-20
C4174 a_17405_8741# 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 0.121f
C4175 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_17405_7309# 0.019f
C4176 a_8643_n6471# D2_2 0.0541f
C4177 Q3 Q5 1.46f
C4178 Q7 Q4 0.0457f
C4179 LD Q2 11.2f
C4180 a_1559_n1526# a_1541_n3150# 0.00121f
C4181 a_1541_n8095# VDD 0.18f
C4182 a_5054_n1526# D2_5 0.0503f
C4183 p2_gen_magic_0.xnor_magic_4.OUT a_8643_n1526# 2.24e-19
C4184 a_2749_3524# VDD 0.941f
C4185 a_24003_10051# Q2 9.92e-20
C4186 a_19841_8580# a_20041_8580# 0.296f
C4187 a_18891_6886# a_20041_4557# 7.7e-19
C4188 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_4.OUT 1.59e-21
C4189 p3_gen_magic_0.xnor_magic_3.OUT a_1975_n6471# 0.0629f
C4190 a_5036_n4081# D2_5 0.05f
C4191 p2_gen_magic_0.xnor_magic_1.OUT a_16386_n3644# 0.132f
C4192 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A a_12931_1059# 0.0292f
C4193 Q1 D2_6 0.897f
C4194 p3_gen_magic_0.3_inp_AND_magic_0.C a_14556_n8142# 5.36e-19
C4195 7b_counter_0.DFF_magic_0.Q 7b_counter_0.MDFF_4.LD 1.05f
C4196 a_8523_n8095# D2_2 3.13e-19
C4197 a_11279_6341# D2_2 0.132f
C4198 p3_gen_magic_0.xnor_magic_4.OUT Q6 0.121f
C4199 a_1409_2253# a_1409_1059# 0.0206f
C4200 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT D2_4 0.00273f
C4201 p3_gen_magic_0.xnor_magic_1.OUT a_14756_n8142# 1.75e-19
C4202 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q3 0.00144f
C4203 7b_counter_0.DFF_magic_0.Q 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 0.00191f
C4204 a_11292_n6613# a_13353_n6613# 6.01e-20
C4205 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p3_gen_magic_0.AND2_magic_1.A 0.212f
C4206 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A CLK 0.0864f
C4207 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_18891_6886# 0.654f
C4208 a_21381_4932# Q4 0.00304f
C4209 Q3 D2_4 2.86f
C4210 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN CLK 0.61f
C4211 a_27778_3363# CLK 0.00209f
C4212 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_7 1.01f
C4213 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_1209_1059# 1.63e-20
C4214 7b_counter_0.3_inp_AND_magic_0.A Q3 0.0113f
C4215 a_4235_9163# 7b_counter_0.MDFF_3.tspc2_magic_0.Q 1.94e-20
C4216 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_12387_8536# 1.08e-19
C4217 a_17405_10149# a_15865_8580# 1.14e-19
C4218 p3_gen_magic_0.xnor_magic_1.B a_1957_n7648# 0.00157f
C4219 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A VDD 1.33f
C4220 a_12387_6963# a_12387_5769# 0.00638f
C4221 a_15865_7470# Q1 3.82e-19
C4222 a_12387_4513# VDD 0.975f
C4223 DFF_magic_0.D OR_magic_1.VOUT 0.00188f
C4224 a_23258_1746# a_23802_2253# 0.296f
C4225 p3_gen_magic_0.3_inp_AND_magic_0.A VDD 1.34f
C4226 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B D2_5 0.0063f
C4227 a_5054_n6024# D2_7 6.69e-21
C4228 a_12387_5769# CLK 0.0162f
C4229 7b_counter_0.MDFF_7.tspc2_magic_0.D D2_4 0.0841f
C4230 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A Q6 0.0232f
C4231 a_11279_6341# a_9212_5956# 8.2e-19
C4232 a_6725_7308# 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A 2.4e-20
C4233 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 0.00753f
C4234 7b_counter_0.DFF_magic_0.D CLK 0.678f
C4235 a_1209_7469# VDD 0.87f
C4236 7b_counter_0.3_inp_AND_magic_0.A 7b_counter_0.MDFF_7.tspc2_magic_0.D 3.94e-20
C4237 divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT mux_magic_0.AND2_magic_0.A 4.32e-20
C4238 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B a_6725_5900# 0.173f
C4239 7b_counter_0.MDFF_4.LD Q5 2.49f
C4240 p3_gen_magic_0.3_inp_AND_magic_0.A D2_1 0.0042f
C4241 a_23207_5815# Q6 3.27e-21
C4242 Q2 Q3 2.44f
C4243 a_16065_9774# CLK 0.124f
C4244 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A VDD 1.23f
C4245 p2_gen_magic_0.xnor_magic_1.OUT p2_gen_magic_0.xnor_magic_5.OUT 1.31f
C4246 a_8955_8580# VDD 0.0856f
C4247 a_5054_n1526# D2_7 1.66e-20
C4248 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A VDD 1.24f
C4249 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT a_1957_n3150# 0.00157f
C4250 a_22150_1124# a_22062_684# 0.475f
C4251 a_17405_2092# a_15865_1059# 7.16e-20
C4252 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A D2_3 0.0145f
C4253 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT Q5 0.00101f
C4254 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 5.61e-19
C4255 divide_by_2_1.tg_magic_3.CLK divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT 1.84e-19
C4256 a_5036_n4081# D2_7 0.00786f
C4257 a_15865_9774# Q1 3.56e-19
C4258 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT 0.00535f
C4259 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 0.00123f
C4260 a_1209_3363# Q6 0.0021f
C4261 Q1 D2_2 0.723f
C4262 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A 1.1e-20
C4263 p3_gen_magic_0.xnor_magic_1.B p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 0.00123f
C4264 7b_counter_0.MDFF_5.tspc2_magic_0.CLK VDD 2.16f
C4265 a_23258_552# Q4 5.53e-20
C4266 OR_magic_2.VOUT divide_by_2_0.tg_magic_3.OUT 0.413f
C4267 p2_gen_magic_0.AND2_magic_1.A a_12174_n4081# 0.613f
C4268 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B CLK 0.0127f
C4269 a_1209_7469# LD 0.195f
C4270 7b_counter_0.MDFF_4.LD D2_4 0.812f
C4271 a_2749_8740# 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 0.019f
C4272 p3_gen_magic_0.xnor_magic_6.OUT Q4 0.228f
C4273 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_3.OUT 3.29e-20
C4274 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5054_n6024# 0.0628f
C4275 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A a_26038_684# 0.397f
C4276 a_1541_n8095# Q3 6.69e-21
C4277 a_2749_7308# Q7 0.0104f
C4278 7b_counter_0.DFF_magic_0.D 7b_counter_0.3_inp_AND_magic_0.C 0.152f
C4279 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A CLK 0.0147f
C4280 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_4 1.17f
C4281 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B VDD 1.21f
C4282 a_12387_6963# a_11279_6341# 0.00114f
C4283 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_2.IN 0.965f
C4284 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A Q1 3.35e-19
C4285 p3_gen_magic_0.xnor_magic_1.B a_14556_n8142# 0.00128f
C4286 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT VDD 1.49f
C4287 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B a_17405_3524# 0.412f
C4288 a_2749_5900# CLK 0.00119f
C4289 a_11279_6341# CLK 0.0096f
C4290 a_5036_n4081# p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 8.45e-21
C4291 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B Q4 0.00109f
C4292 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT Q6 0.631f
C4293 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A a_16065_8580# 0.00103f
C4294 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A Q1 0.00118f
C4295 a_8523_n8579# Q5 2.81e-19
C4296 7b_counter_0.MDFF_4.LD Q2 0.204f
C4297 a_22991_5815# a_23207_5815# 0.914f
C4298 7b_counter_0.MDFF_3.QB Q2 2.59f
C4299 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A Q3 8.78e-21
C4300 a_12174_n7648# VDD 0.0014f
C4301 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT Q2 0.0231f
C4302 a_21381_8741# Q2 5.13e-19
C4303 a_2749_4932# VDD 1.55f
C4304 a_9212_739# p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 5.26e-20
C4305 p3_gen_magic_0.xnor_magic_3.OUT a_1559_n6471# 0.0924f
C4306 a_12174_n3150# D2_3 6.39e-19
C4307 p2_gen_magic_0.xnor_magic_1.OUT a_14756_n3644# 0.00254f
C4308 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A a_12387_552# 0.251f
C4309 7b_counter_0.MDFF_1.tspc2_magic_0.CLK D2_3 0.0697f
C4310 a_19152_6440# a_20171_6886# 0.0292f
C4311 a_19152_6440# Q1 0.0126f
C4312 7b_counter_0.MDFF_1.tspc2_magic_0.CLK 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B 0.00594f
C4313 DFF_magic_0.tg_magic_3.CLK DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 1.37f
C4314 a_11279_8697# a_11279_6341# 0.00112f
C4315 a_4651_3947# a_5515_3947# 0.00862f
C4316 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.AND2_magic_1.A 0.212f
C4317 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A a_1409_8579# 1.77e-19
C4318 p3_gen_magic_0.xnor_magic_1.OUT a_16186_n8142# 0.254f
C4319 a_1209_2253# a_1409_1059# 0.00308f
C4320 a_4496_9609# a_5385_7469# 5.39e-19
C4321 Q4 D2_3 0.556f
C4322 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A 0.421f
C4323 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B Q4 5.49e-19
C4324 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A Q3 1.93e-19
C4325 7b_counter_0.DFF_magic_0.tg_magic_3.OUT VDD 1.15f
C4326 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1957_n7648# 1.46e-20
C4327 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A a_1209_8579# 1.03e-19
C4328 a_20041_3363# CLK 3.99e-19
C4329 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A a_6725_2092# 0.0334f
C4330 a_12387_1746# 7b_counter_0.MDFF_4.tspc2_magic_0.D 7.57e-20
C4331 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A Q3 0.00376f
C4332 a_15865_4557# VDD 0.988f
C4333 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_9059_n1973# 0.00157f
C4334 p3_gen_magic_0.P3 a_23352_n5390# 0.175f
C4335 a_32816_n1264# a_32616_n2458# 0.00308f
C4336 a_8643_n5540# VDD 0.376f
C4337 7b_counter_0.MDFF_7.tspc2_magic_0.CLK CLK 0.0421f
C4338 Q1 CLK 1.17f
C4339 a_1559_n1973# p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT 7.35e-19
C4340 a_12387_3319# Q5 0.0418f
C4341 a_23560_3728# Q5 7.87e-19
C4342 a_24401_7877# VDD 0.0231f
C4343 7b_counter_0.MDFF_3.tspc2_magic_0.Q Q7 0.101f
C4344 a_22991_5815# Q6 2.82e-19
C4345 a_5515_9163# CLK 0.00291f
C4346 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT Q1 0.265f
C4347 p2_gen_magic_0.xnor_magic_1.OUT D2_6 0.00505f
C4348 a_19841_8580# VDD 0.982f
C4349 7b_counter_0.DFF_magic_0.tg_magic_3.OUT LD 0.0186f
C4350 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 0.4f
C4351 a_1409_4557# a_1409_3363# 0.0206f
C4352 a_1559_n1526# D2_7 0.0159f
C4353 p3_gen_magic_0.3_inp_AND_magic_0.A p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT 0.00302f
C4354 a_17405_3524# VDD 0.929f
C4355 p3_gen_magic_0.xnor_magic_1.OUT a_1957_n7648# 0.0636f
C4356 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A Q5 0.00225f
C4357 7b_counter_0.MDFF_4.LD a_12387_4513# 0.00288f
C4358 a_1541_n4081# D2_7 0.00265f
C4359 a_19841_8580# D2_1 0.223f
C4360 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q3 0.00122f
C4361 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT D2_6 0.0827f
C4362 a_17405_10149# VDD 1.55f
C4363 a_1975_n1973# a_1541_n3597# 3.04e-19
C4364 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A VDD 1.23f
C4365 a_27234_1746# D2_4 0.0119f
C4366 a_23560_3728# D2_4 0.0195f
C4367 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A a_11191_5901# 0.397f
C4368 a_5385_1059# D2_5 0.00754f
C4369 7b_counter_0.MDFF_5.LD D2_6 0.0923f
C4370 a_11292_n6613# a_11708_n6613# 0.278f
C4371 7b_counter_0.DFF_magic_0.tg_magic_0.IN D2_4 0.00267f
C4372 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A 8.78e-21
C4373 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN 0.316f
C4374 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A a_21381_10149# 3.58e-20
C4375 a_2749_10148# 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 0.00215f
C4376 7b_counter_0.MDFF_7.tspc2_magic_0.D 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B 0.00171f
C4377 mux_magic_0.OR_magic_0.B mux_magic_0.IN2 0.00118f
C4378 a_17405_10149# D2_1 0.0161f
C4379 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A 8.54e-19
C4380 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT VDD 1.17f
C4381 7b_counter_0.3_inp_AND_magic_0.C Q1 0.0446f
C4382 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD 1.09f
C4383 a_26126_1124# a_26038_684# 0.475f
C4384 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A 1.1e-20
C4385 p3_gen_magic_0.xnor_magic_0.OUT Q4 0.00945f
C4386 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 5.61e-19
C4387 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT D2_3 2.9e-19
C4388 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A D2_4 0.0203f
C4389 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.3_inp_AND_magic_0.C 0.00798f
C4390 a_11292_n2115# p2_gen_magic_0.3_inp_AND_magic_0.B 0.00234f
C4391 a_5054_n1042# D2_5 0.0504f
C4392 a_19152_1223# a_20171_1669# 0.0292f
C4393 a_11191_684# a_12387_552# 7.98e-19
C4394 a_8411_9730# Q6 3.77e-19
C4395 a_17405_8741# Q1 0.0436f
C4396 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_15865_2253# 4.8e-20
C4397 a_1559_n1042# VDD 0.415f
C4398 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_7 8.88e-19
C4399 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK 0.00408f
C4400 7b_counter_0.MDFF_5.LD a_15865_7470# 0.195f
C4401 a_17405_7309# Q1 1.7e-19
C4402 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 7b_counter_0.MDFF_4.LD 3.09e-20
C4403 7b_counter_0.DFF_magic_0.tg_magic_2.OUT VDD 1.21f
C4404 a_5515_3947# Q7 0.00491f
C4405 mux_magic_0.IN2 divide_by_2_0.tg_magic_3.IN 0.324f
C4406 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 0.157f
C4407 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_1.OUT 0.0623f
C4408 a_6725_7308# CLK 9.8e-20
C4409 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A Q5 6.14e-19
C4410 a_5036_n8579# Q5 1.88e-19
C4411 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B Q6 0.0539f
C4412 a_19841_9774# a_20041_9774# 0.297f
C4413 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.3_inp_AND_magic_0.B 7.68e-21
C4414 p2_gen_magic_0.xnor_magic_1.OUT D2_2 0.00537f
C4415 a_8939_n7648# VDD 0.0018f
C4416 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5470_n6471# 0.00157f
C4417 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A a_11279_3480# 2.07e-19
C4418 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A Q6 4.53e-19
C4419 p3_gen_magic_0.xnor_magic_3.OUT a_5054_n6024# 1.65e-19
C4420 p2_gen_magic_0.xnor_magic_1.OUT a_16186_n3644# 0.256f
C4421 a_18891_6886# Q1 0.00247f
C4422 7b_counter_0.3_inp_AND_magic_0.VOUT 7b_counter_0.3_inp_AND_magic_0.C 0.407f
C4423 a_11191_5901# a_12387_5769# 7.98e-19
C4424 a_19152_6440# a_19307_6886# 0.235f
C4425 a_18891_6886# a_20171_6886# 0.00652f
C4426 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8643_n1042# 0.0528f
C4427 a_8411_4513# a_7303_3480# 7.16e-20
C4428 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A Q6 0.0438f
C4429 7b_counter_0.MDFF_5.LD a_15865_9774# 0.0336f
C4430 p3_gen_magic_0.xnor_magic_1.OUT a_14556_n8142# 0.0203f
C4431 a_1209_2253# a_1209_1059# 0.00638f
C4432 a_24401_7877# Q3 7.62e-20
C4433 7b_counter_0.MDFF_5.LD D2_2 0.504f
C4434 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A Q1 0.00645f
C4435 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_8643_n5540# 0.0802f
C4436 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B 0.00506f
C4437 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 0.00677f
C4438 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_12174_n7648# 0.102f
C4439 a_27234_3319# CLK 0.00757f
C4440 divide_by_2_1.tg_magic_3.CLK divide_by_2_1.tg_magic_1.IN 0.0617f
C4441 a_4496_10093# a_4235_9163# 0.651f
C4442 a_11279_3480# VDD 0.929f
C4443 a_32616_n2458# a_32816_n2458# 0.298f
C4444 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8643_n1973# 0.00941f
C4445 a_15865_7470# a_17405_5901# 1.14e-19
C4446 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT 1.09f
C4447 a_34156_n2297# a_32616_n2458# 0.00114f
C4448 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B CLK 0.0127f
C4449 a_21381_3524# CLK 0.00325f
C4450 a_5054_n6471# p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 0.00172f
C4451 a_15865_4557# a_15865_3363# 0.00638f
C4452 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A 0.00157f
C4453 a_24185_7877# VDD 0.021f
C4454 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A Q2 0.335f
C4455 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD 1.09f
C4456 a_11708_n2115# D2_2 0.0064f
C4457 a_23793_5904# Q5 0.531f
C4458 7b_counter_0.MDFF_6.tspc2_magic_0.Q Q2 0.001f
C4459 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT a_12174_n8579# 0.0542f
C4460 DFF_magic_0.tg_magic_3.CLK DFF_magic_0.tg_magic_2.IN 0.694f
C4461 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT Q4 0.0237f
C4462 7b_counter_0.MDFF_4.LD 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 1.64e-20
C4463 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5452_n3150# 7.77e-21
C4464 a_4651_9163# CLK 0.00289f
C4465 a_12387_4513# a_12387_3319# 0.00638f
C4466 p2_gen_magic_0.xnor_magic_1.OUT a_1957_n3150# 0.0629f
C4467 p2_gen_magic_0.xnor_magic_5.OUT D2_5 1.1f
C4468 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT Q3 0.00347f
C4469 p2_gen_magic_0.3_inp_AND_magic_0.VOUT Q4 0.139f
C4470 7b_counter_0.MDFF_4.LD a_15865_4557# 0.00288f
C4471 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A 0.00221f
C4472 a_12931_4557# VDD 0.0559f
C4473 a_11279_1124# Q5 5.93e-19
C4474 a_1541_n7648# a_1957_n7648# 0.00222f
C4475 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT Q5 0.0148f
C4476 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN P2 0.29f
C4477 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 4e-20
C4478 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.LD 0.4f
C4479 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK 2.39e-20
C4480 a_1409_2253# 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A 0.00103f
C4481 a_1559_n1042# Q3 0.00132f
C4482 a_1559_n1973# a_1541_n3597# 5.1e-19
C4483 a_19841_9774# VDD 0.959f
C4484 a_23802_2253# D2_4 0.119f
C4485 DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK 1.33f
C4486 a_11279_6341# a_11191_5901# 0.473f
C4487 a_5185_1059# D2_5 0.0195f
C4488 a_23793_5904# D2_4 0.00663f
C4489 a_11292_n6613# a_11492_n6613# 0.519f
C4490 7b_counter_0.MDFF_5.LD a_19152_6440# 0.00691f
C4491 a_17405_3524# a_15865_3363# 0.00114f
C4492 7b_counter_0.3_inp_AND_magic_0.A a_23793_5904# 0.896f
C4493 a_1209_9773# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A 0.128f
C4494 p2_gen_magic_0.xnor_magic_1.OUT CLK 0.151f
C4495 a_2749_684# D2_4 0.00871f
C4496 7b_counter_0.MDFF_4.LD a_17405_3524# 0.00115f
C4497 a_12174_n4081# Q4 0.00175f
C4498 a_11279_1124# D2_4 0.00853f
C4499 DFF_magic_0.D P2 0.627f
C4500 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_9212_739# 7.16e-19
C4501 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT Q6 0.0205f
C4502 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_4496_9609# 0.0125f
C4503 a_21381_8741# a_19841_8580# 0.00114f
C4504 a_19152_1223# a_19307_1669# 0.235f
C4505 a_18891_1669# a_20171_1669# 0.00652f
C4506 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_1.OUT 0.00178f
C4507 a_12931_9774# Q1 0.12f
C4508 7b_counter_0.MDFF_5.LD a_12387_6963# 0.195f
C4509 7b_counter_0.MDFF_4.tspc2_magic_0.CLK Q5 0.307f
C4510 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A 0.00221f
C4511 a_17405_7309# a_19307_6886# 2.12e-20
C4512 a_4651_3947# Q7 0.00361f
C4513 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT CLK 0.229f
C4514 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 0.0214f
C4515 a_19841_9774# LD 6.64e-19
C4516 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A a_21381_10149# 0.397f
C4517 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN VDD 1.25f
C4518 7b_counter_0.MDFF_5.LD CLK 0.929f
C4519 a_1541_n8579# Q5 0.00425f
C4520 p3_gen_magic_0.3_inp_AND_magic_0.B D2_6 0.0452f
C4521 p2_gen_magic_0.xnor_magic_5.OUT D2_7 0.136f
C4522 7b_counter_0.MDFF_4.LD DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 8.64e-19
C4523 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5054_n6471# 0.00265f
C4524 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A Q7 6.76e-19
C4525 p2_gen_magic_0.xnor_magic_4.OUT a_5054_n1526# 0.415f
C4526 a_23258_1746# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A 0.00184f
C4527 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK P2 0.0281f
C4528 p3_gen_magic_0.xnor_magic_3.OUT a_1559_n6024# 0.368f
C4529 p3_gen_magic_0.xnor_magic_4.OUT VDD 1.47f
C4530 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 0.00325f
C4531 p2_gen_magic_0.xnor_magic_1.OUT a_14556_n3644# 0.0229f
C4532 a_14756_n3644# D2_5 0.00137f
C4533 a_18891_6886# a_19307_6886# 0.153f
C4534 a_6725_2092# a_6725_684# 0.475f
C4535 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 1.37f
C4536 7b_counter_0.DFF_magic_0.Q a_23985_7877# 0.00115f
C4537 7b_counter_0.MDFF_4.tspc2_magic_0.CLK D2_4 0.00126f
C4538 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT Q4 0.00236f
C4539 7b_counter_0.MDFF_4.LD 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 0.00112f
C4540 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_0.IN 0.287f
C4541 7b_counter_0.3_inp_AND_magic_0.B a_19152_6440# 8.75e-21
C4542 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_12174_n3150# 0.102f
C4543 a_8411_9730# a_8411_8536# 0.00638f
C4544 a_27778_1059# CLK 0.00664f
C4545 a_24185_7877# Q3 1.32e-19
C4546 7b_counter_0.MDFF_5.LD a_11279_8697# 0.00115f
C4547 a_8955_4557# Q1 6.2e-19
C4548 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT a_1541_n8579# 0.057f
C4549 p3_gen_magic_0.xnor_magic_4.OUT D2_1 0.00287f
C4550 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1559_n1042# 0.0846f
C4551 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 0.156f
C4552 DFF_magic_0.D VDD 8.74f
C4553 a_9689_1669# a_9412_739# 0.00164f
C4554 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT Q4 0.0252f
C4555 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A 0.178f
C4556 a_24536_3947# CLK 1.41e-20
C4557 p2_gen_magic_0.3_inp_AND_magic_0.B a_13769_n2115# 0.109f
C4558 a_11191_4932# VDD 1.55f
C4559 a_2749_8740# a_2749_7308# 0.00112f
C4560 a_5185_2253# Q6 0.00164f
C4561 7b_counter_0.MDFF_5.LD 7b_counter_0.3_inp_AND_magic_0.C 0.00111f
C4562 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 1.59e-20
C4563 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A VDD 1.24f
C4564 a_34156_n889# a_32616_n2458# 1.14e-19
C4565 a_1559_n1526# p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT 7.02e-19
C4566 a_19152_1223# Q5 8.58e-19
C4567 a_8411_3319# Q5 7.02e-19
C4568 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT a_12174_n4081# 0.0542f
C4569 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK 0.043f
C4570 a_23207_5815# VDD 0.185f
C4571 7b_counter_0.MDFF_5.LD a_17405_8741# 0.0139f
C4572 a_11492_n2115# D2_2 0.00891f
C4573 a_1559_n5540# Q7 1.35e-19
C4574 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT a_1541_n4081# 0.0832f
C4575 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_0.IN 0.85f
C4576 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK VDD 4.25f
C4577 a_23985_7877# Q5 5.61e-19
C4578 D2_5 D2_6 0.029f
C4579 DFF_magic_0.D LD 0.478f
C4580 a_1541_n3150# a_1957_n3150# 0.00222f
C4581 a_13353_n2115# Q4 0.0198f
C4582 a_5036_n3150# D2_5 0.0786f
C4583 7b_counter_0.MDFF_6.tspc2_magic_0.D D2_3 0.0977f
C4584 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.xnor_magic_6.OUT 0.149f
C4585 7b_counter_0.MDFF_4.LD a_11279_3480# 0.00115f
C4586 a_7215_4932# a_8411_3319# 1.14e-19
C4587 a_1209_3363# VDD 0.87f
C4588 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A a_8411_3319# 0.00184f
C4589 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT 0.244f
C4590 a_6725_2092# Q5 0.156f
C4591 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT 0.156f
C4592 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A a_7303_8697# 2.4e-20
C4593 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B D2_4 0.00379f
C4594 a_1209_2253# 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A 1.03e-19
C4595 OR_magic_1.VOUT P2 0.0146f
C4596 a_19152_1223# D2_4 0.0429f
C4597 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A LD 1.1e-20
C4598 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT D2_3 0.047f
C4599 7b_counter_0.MDFF_4.tspc2_magic_0.D a_9412_739# 0.103f
C4600 a_8411_4513# D2_6 0.0187f
C4601 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A Q6 8.78e-21
C4602 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_6 1.01f
C4603 a_23985_7877# D2_4 0.0117f
C4604 a_8523_n3597# Q1 0.022f
C4605 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A D2_7 0.0168f
C4606 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_5385_2253# 0.00751f
C4607 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT 0.00322f
C4608 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT 0.00312f
C4609 7b_counter_0.3_inp_AND_magic_0.B 7b_counter_0.3_inp_AND_magic_0.C 0.347f
C4610 7b_counter_0.3_inp_AND_magic_0.A a_23985_7877# 0.383f
C4611 a_1541_n8095# a_1541_n8579# 0.0335f
C4612 p3_gen_magic_0.AND2_magic_1.A a_16386_n8142# 3.84e-19
C4613 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A a_12387_3319# 0.00184f
C4614 7b_counter_0.MDFF_4.LD a_12931_4557# 0.00428f
C4615 a_6725_2092# D2_4 0.00548f
C4616 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A VDD 1.23f
C4617 a_1209_3363# LD 0.195f
C4618 a_4235_9163# a_4496_9609# 0.299f
C4619 a_18891_1669# a_19307_1669# 0.153f
C4620 a_5054_n6471# a_5470_n6471# 5.82e-19
C4621 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 0.16f
C4622 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 0.0213f
C4623 DFF_magic_0.D 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 0.00183f
C4624 a_17405_7309# a_17405_5901# 0.475f
C4625 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.101f
C4626 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT VDD 1.48f
C4627 p2_gen_magic_0.xnor_magic_0.OUT VDD 0.632f
C4628 a_21381_4932# Q7 0.00278f
C4629 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A D2_1 0.00542f
C4630 a_9059_n1973# D2_6 0.00115f
C4631 VDD Q6 9.42f
C4632 DFF_magic_0.D Q3 0.32f
C4633 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A 0.00112f
C4634 a_19841_9774# a_21381_8741# 7.16e-20
C4635 a_8825_6886# a_9689_6886# 0.00862f
C4636 a_7303_8697# CLK 0.0164f
C4637 a_23985_7877# Q2 4.76e-19
C4638 7b_counter_0.MDFF_3.tspc2_magic_0.D a_4235_9163# 0.278f
C4639 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.3_inp_AND_magic_0.C 0.236f
C4640 D2_2 D2_5 0.297f
C4641 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT D2_1 0.00981f
C4642 a_5036_n3150# D2_7 0.642f
C4643 a_12387_4513# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 1.63e-20
C4644 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A a_15865_4557# 0.251f
C4645 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD 1.09f
C4646 D2_1 Q6 2.17f
C4647 OR_magic_1.VOUT VDD 7.84f
C4648 a_8955_9774# Q7 0.0263f
C4649 a_23258_1746# a_22150_1124# 0.00114f
C4650 a_1209_1059# p2_gen_magic_0.xnor_magic_3.OUT 1.7e-19
C4651 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A LD 5.6e-19
C4652 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT D2_1 0.0166f
C4653 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 7b_counter_0.DFF_magic_0.tg_magic_0.IN 0.0105f
C4654 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_3 3.57e-19
C4655 p3_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.AND2_magic_1.A 0.426f
C4656 p3_gen_magic_0.xnor_magic_1.OUT a_8523_n8095# 0.00376f
C4657 a_5054_n1973# a_5470_n1973# 5.82e-19
C4658 a_23207_5815# Q3 0.187f
C4659 7b_counter_0.MDFF_5.LD a_11191_10149# 0.00267f
C4660 OR_magic_2.VOUT divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT 1.31f
C4661 a_17405_5901# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A 1.51e-21
C4662 p3_gen_magic_0.P3 CLK 0.234f
C4663 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_2 0.00101f
C4664 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK Q3 0.0676f
C4665 a_1409_8579# VDD 0.0124f
C4666 LD Q6 1.55f
C4667 a_1409_7469# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A 1.77e-19
C4668 a_23672_3947# CLK 1.38e-20
C4669 p2_gen_magic_0.3_inp_AND_magic_0.B a_13553_n2115# 0.163f
C4670 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_19841_8580# 0.0276f
C4671 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A a_17405_3524# 2.4e-20
C4672 divide_by_2_1.tg_magic_3.CLK divide_by_2_1.tg_magic_3.IN 0.951f
C4673 p2_gen_magic_0.3_inp_AND_magic_0.A D2_2 0.00592f
C4674 DFF_magic_0.tg_magic_1.IN CLK 0.682f
C4675 a_8825_6886# Q7 0.0019f
C4676 p3_gen_magic_0.P3 OR_magic_2.VOUT 0.00359f
C4677 7b_counter_0.MDFF_5.tspc2_magic_0.D a_9689_6886# 0.00451f
C4678 p3_gen_magic_0.xnor_magic_5.OUT Q5 0.0296f
C4679 DFF_magic_0.D OR_magic_2.A 0.394f
C4680 a_18891_1669# Q5 3.37e-20
C4681 a_8713_1625# a_9689_1669# 0.235f
C4682 7b_counter_0.MDFF_5.LD a_12931_9774# 0.00428f
C4683 a_22991_5815# VDD 1.1f
C4684 a_11279_3480# a_12387_3319# 0.00114f
C4685 a_9059_n1973# D2_2 0.00157f
C4686 DFF_magic_0.D 7b_counter_0.MDFF_4.LD 1.05f
C4687 p3_gen_magic_0.3_inp_AND_magic_0.A p3_gen_magic_0.3_inp_AND_magic_0.VOUT 3.5e-19
C4688 a_5470_n6471# D2_3 0.00157f
C4689 a_1409_8579# LD 0.0292f
C4690 a_32616_n1264# a_32816_n1264# 0.297f
C4691 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B Q4 0.00246f
C4692 a_5185_2253# 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A 1.03e-19
C4693 p2_gen_magic_0.xnor_magic_0.OUT a_8523_n3150# 0.0374f
C4694 7b_counter_0.MDFF_4.LD a_11191_4932# 0.00267f
C4695 DFF_magic_0.D 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 0.0258f
C4696 a_19152_6440# 7b_counter_0.MDFF_1.tspc2_magic_0.Q 0.00119f
C4697 p2_gen_magic_0.xnor_magic_3.OUT a_11292_n2115# 0.483f
C4698 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT a_5452_n7648# 0.00157f
C4699 a_22150_1124# a_20171_1669# 6.59e-21
C4700 a_5470_n1973# D2_3 0.00157f
C4701 a_2749_5900# a_1209_6275# 7.98e-19
C4702 p2_gen_magic_0.xnor_magic_0.OUT Q3 0.00577f
C4703 a_18891_1669# D2_4 0.0163f
C4704 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_8643_n1526# 0.0629f
C4705 7b_counter_0.DFF_magic_0.tg_magic_0.IN 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.26f
C4706 a_26126_3480# D2_4 0.0852f
C4707 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A a_12387_8536# 1.03e-19
C4708 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B a_2749_2092# 0.412f
C4709 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A Q5 0.00312f
C4710 Q3 Q6 0.0406f
C4711 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_3.OUT 7.64e-21
C4712 p2_gen_magic_0.AND2_magic_1.A a_16386_n3644# 3.84e-19
C4713 a_1541_n3597# a_1541_n4081# 0.0335f
C4714 a_12931_4557# a_12387_3319# 0.00308f
C4715 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 1.61e-19
C4716 mux_magic_0.OR_magic_0.B a_32616_n2458# 0.125f
C4717 7b_counter_0.MDFF_4.LD p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK 6.76e-19
C4718 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_2749_2092# 0.121f
C4719 p3_gen_magic_0.AND2_magic_1.A a_14756_n8142# 0.0292f
C4720 a_21504_5904# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A 3.96e-19
C4721 CLK D2_5 2.04f
C4722 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT Q1 0.0189f
C4723 a_8643_n1042# D2_6 0.0186f
C4724 p2_gen_magic_0.3_inp_AND_magic_0.B p2_gen_magic_0.xnor_magic_1.OUT 0.0406f
C4725 7b_counter_0.MDFF_1.tspc2_magic_0.Q CLK 0.247f
C4726 7b_counter_0.DFF_magic_0.tg_magic_3.CLK CLK 0.635f
C4727 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A a_8955_3363# 5.46e-20
C4728 a_8411_9730# VDD 0.972f
C4729 7b_counter_0.MDFF_7.tspc2_magic_0.Q 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 0.25f
C4730 a_4496_10093# a_4496_9609# 0.0141f
C4731 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT D2_5 0.0567f
C4732 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B a_1209_8579# 0.125f
C4733 p2_gen_magic_0.xnor_magic_4.OUT a_5054_n1042# 0.297f
C4734 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_5.OUT 5.37e-19
C4735 7b_counter_0.MDFF_4.tspc2_magic_0.D a_8713_1625# 0.0379f
C4736 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 0.0037f
C4737 p3_gen_magic_0.xnor_magic_5.OUT Q2 1.22e-20
C4738 Q7 D2_3 0.0599f
C4739 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A D2_4 0.0293f
C4740 a_8411_9730# D2_1 3.33e-19
C4741 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_17405_3524# 1e-20
C4742 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B VDD 1.2f
C4743 a_8643_n1973# D2_6 0.0124f
C4744 p3_gen_magic_0.3_inp_AND_magic_0.A a_13769_n6613# 0.0247f
C4745 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B 0.00112f
C4746 7b_counter_0.MDFF_3.tspc2_magic_0.D a_4496_10093# 0.103f
C4747 a_2749_8740# a_4235_9163# 0.00212f
C4748 a_1957_n3150# D2_7 6.21e-19
C4749 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A a_23802_1059# 0.0292f
C4750 a_26038_684# 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 3.58e-20
C4751 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B D2_1 0.00118f
C4752 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A VDD 1.32f
C4753 a_8955_3363# VDD 0.0856f
C4754 a_4496_9609# Q7 5.19e-19
C4755 7b_counter_0.MDFF_3.QB 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A 0.00362f
C4756 a_14556_n3644# D2_5 5.98e-19
C4757 p2_gen_magic_0.xnor_magic_5.OUT p2_gen_magic_0.AND2_magic_1.A 0.425f
C4758 a_8411_9730# LD 6.64e-19
C4759 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A D2_1 4.06e-19
C4760 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A VDD 1.39f
C4761 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A Q5 1.03e-21
C4762 a_27234_4513# D2_4 0.00447f
C4763 a_12931_7470# Q2 0.073f
C4764 p2_gen_magic_0.3_inp_AND_magic_0.C Q5 7.55e-20
C4765 a_22991_5815# Q3 0.032f
C4766 7b_counter_0.3_inp_AND_magic_0.C 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 5.03e-20
C4767 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT 5.61e-19
C4768 p3_gen_magic_0.P3 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN 0.289f
C4769 OR_magic_1.VOUT mux_magic_0.IN1 0.00723f
C4770 7b_counter_0.MDFF_3.QB Q6 0.124f
C4771 OR_magic_2.A OR_magic_1.VOUT 0.0582f
C4772 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B LD 6.96e-19
C4773 a_8411_8536# VDD 0.982f
C4774 a_16065_3363# CLK 0.172f
C4775 a_1209_7469# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A 0.00184f
C4776 p2_gen_magic_0.3_inp_AND_magic_0.B a_11708_n2115# 0.00272f
C4777 a_21381_8741# Q6 0.153f
C4778 7b_counter_0.MDFF_4.LD OR_magic_1.VOUT 0.003f
C4779 CLK D2_7 0.69f
C4780 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A VDD 1.23f
C4781 a_8643_n1042# D2_2 0.00867f
C4782 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A LD 7.66e-19
C4783 a_6725_5900# Q7 0.0153f
C4784 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT D2_7 0.00173f
C4785 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A D2_4 0.0208f
C4786 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 4.89e-20
C4787 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_19841_9774# 0.223f
C4788 a_5036_n7648# Q5 0.69f
C4789 divide_by_2_1.tg_magic_3.IN OUT1 2.8e-19
C4790 DFF_magic_0.D a_27234_1746# 6.41e-19
C4791 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A LD 0.4f
C4792 p2_gen_magic_0.3_inp_AND_magic_0.C D2_4 0.00218f
C4793 a_8713_1625# a_8825_1669# 0.0292f
C4794 a_24259_4877# Q5 8.26e-19
C4795 a_11191_4932# a_12387_3319# 1.14e-19
C4796 a_8643_n1973# D2_2 0.0542f
C4797 a_20041_8580# VDD 0.0856f
C4798 a_5054_n6471# D2_3 0.0541f
C4799 a_12931_3363# D2_2 0.0012f
C4800 p3_gen_magic_0.3_inp_AND_magic_0.B p3_gen_magic_0.3_inp_AND_magic_0.C 1.3f
C4801 p3_gen_magic_0.3_inp_AND_magic_0.A a_13353_n6613# 0.467f
C4802 a_7215_10149# Q7 0.0266f
C4803 7b_counter_0.MDFF_3.QB a_1409_8579# 0.0013f
C4804 a_27234_552# CLK 0.00729f
C4805 mux_magic_0.AND2_magic_0.A a_32816_n1264# 0.0291f
C4806 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A Q7 0.0248f
C4807 a_32616_n1264# a_34156_n2297# 7.16e-20
C4808 OR_magic_2.VOUT divide_by_2_0.tg_magic_0.IN 0.61f
C4809 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT a_5452_n3150# 0.00157f
C4810 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.xnor_magic_5.OUT 1.36e-19
C4811 a_15865_8580# VDD 0.884f
C4812 a_18891_6886# 7b_counter_0.MDFF_1.tspc2_magic_0.Q 9.59e-20
C4813 a_20041_8580# D2_1 0.119f
C4814 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q4 1.89e-19
C4815 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A p2_gen_magic_0.xnor_magic_3.OUT 2.5e-19
C4816 a_5452_n3150# Q6 7.91e-19
C4817 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A LD 0.00221f
C4818 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT 3.27e-21
C4819 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B Q1 0.0052f
C4820 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B D2_5 0.0166f
C4821 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT a_23352_n6798# 1.08e-20
C4822 a_5054_n1973# D2_3 0.0541f
C4823 a_11279_3480# a_11279_1124# 0.00112f
C4824 a_15865_8580# D2_1 0.0028f
C4825 a_4496_4393# a_5385_2253# 5.39e-19
C4826 a_11191_684# D2_4 0.0144f
C4827 a_24259_4877# D2_4 0.00761f
C4828 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A a_18891_1669# 3.22e-21
C4829 7b_counter_0.MDFF_0.tspc2_magic_0.CLK D2_5 0.11f
C4830 a_23985_7877# a_24401_7877# 0.278f
C4831 p3_gen_magic_0.xnor_magic_3.OUT D2_6 5.14e-19
C4832 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT 2.83e-19
C4833 p2_gen_magic_0.AND2_magic_1.A a_14756_n3644# 0.0292f
C4834 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT VDD 1.03f
C4835 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B D2_3 4.21e-19
C4836 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B 0.00112f
C4837 a_1209_9773# VDD 0.97f
C4838 7b_counter_0.MDFF_1.tspc2_magic_0.D a_19152_739# 0.103f
C4839 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A Q3 3.45e-19
C4840 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A a_8955_9774# 9.27e-19
C4841 a_5036_n7648# Q2 1.88e-19
C4842 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.0636f
C4843 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A a_2749_4932# 1.52e-21
C4844 a_2749_7308# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B 1.01e-20
C4845 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 3.69e-19
C4846 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 0.00317f
C4847 a_11279_3480# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 0.121f
C4848 a_1209_9773# D2_1 0.00992f
C4849 a_15865_4557# a_17405_4932# 7.98e-19
C4850 p3_gen_magic_0.3_inp_AND_magic_0.A a_13553_n6613# 0.0655f
C4851 a_1209_4557# CLK 0.00168f
C4852 p3_gen_magic_0.3_inp_AND_magic_0.C D2_5 0.00693f
C4853 a_2749_8740# a_4496_10093# 1.39e-20
C4854 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_26126_3480# 0.412f
C4855 7b_counter_0.MDFF_4.tspc2_magic_0.Q Q5 0.428f
C4856 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A VDD 1.38f
C4857 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A Q3 0.0014f
C4858 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A a_16065_3363# 1.77e-19
C4859 a_19841_3363# VDD 0.982f
C4860 a_9689_1669# D2_6 0.0117f
C4861 mux_magic_0.OR_magic_0.A a_32616_n2458# 0.00184f
C4862 7b_counter_0.MDFF_5.LD 7b_counter_0.DFF_magic_0.tg_magic_1.IN 0.0153f
C4863 a_12174_n3597# D2_5 0.243f
C4864 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B D2_3 0.0061f
C4865 p2_gen_magic_0.xnor_magic_1.OUT a_5036_n3597# 1.79e-22
C4866 a_1209_9773# LD 0.00106f
C4867 a_22150_1124# Q5 0.00127f
C4868 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A 7b_counter_0.MDFF_4.tspc2_magic_0.Q 0.00118f
C4869 p2_gen_magic_0.xnor_magic_3.OUT Q1 0.144f
C4870 a_8523_n7648# p3_gen_magic_0.xnor_magic_6.OUT 0.102f
C4871 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A 0.00315f
C4872 p3_gen_magic_0.xnor_magic_3.OUT D2_2 0.0785f
C4873 a_17405_4932# a_17405_3524# 0.475f
C4874 a_20041_9774# VDD 0.0877f
C4875 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.xnor_magic_6.OUT 0.149f
C4876 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B VDD 1.2f
C4877 7b_counter_0.MDFF_4.tspc2_magic_0.Q D2_4 4.33e-19
C4878 a_12931_3363# CLK 0.125f
C4879 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B a_21381_8741# 0.409f
C4880 p2_gen_magic_0.3_inp_AND_magic_0.B a_11492_n2115# 7.27e-19
C4881 7b_counter_0.MDFF_4.LD a_8955_3363# 0.0279f
C4882 a_5185_2253# VDD 1.02f
C4883 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 0.0213f
C4884 a_8643_n1973# p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 1.81e-19
C4885 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK VDD 3.52f
C4886 7b_counter_0.MDFF_1.tspc2_magic_0.D CLK 0.0012f
C4887 7b_counter_0.MDFF_7.tspc2_magic_0.Q CLK 0.0706f
C4888 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_5385_6275# 0.12f
C4889 a_22150_1124# D2_4 0.0128f
C4890 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q5 7.94e-22
C4891 DFF_magic_0.D a_30365_3514# 0.00374f
C4892 a_1957_n7648# Q5 0.0012f
C4893 mux_magic_0.AND2_magic_0.A a_32816_n2458# 0.00103f
C4894 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK D2_1 0.17f
C4895 a_24059_4877# Q5 0.00197f
C4896 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_4.OUT 4.68e-21
C4897 a_5054_n6024# p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 6.69e-21
C4898 a_1975_n1973# Q7 0.0055f
C4899 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8939_n3150# 5.84e-19
C4900 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD 1.09f
C4901 a_12387_9730# Q7 0.0228f
C4902 a_32616_n1264# a_34156_n889# 7.98e-19
C4903 p2_gen_magic_0.xnor_magic_6.OUT VDD 1.34f
C4904 7b_counter_0.MDFF_4.tspc2_magic_0.D D2_6 0.0439f
C4905 VDD P2 4.85f
C4906 mux_magic_0.AND2_magic_0.A a_34156_n2297# 2.4e-20
C4907 a_23802_1059# CLK 0.0052f
C4908 p2_gen_magic_0.xnor_magic_4.OUT D2_6 0.0424f
C4909 7b_counter_0.MDFF_5.tspc2_magic_0.Q a_8713_6842# 0.0129f
C4910 p2_gen_magic_0.xnor_magic_4.OUT a_5036_n3150# 0.0349f
C4911 a_12387_8536# VDD 0.871f
C4912 a_8713_1625# Q4 0.00113f
C4913 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT D2_1 0.0171f
C4914 7b_counter_0.MDFF_3.tspc2_magic_0.D a_4496_9609# 0.0384f
C4915 a_5185_2253# LD 0.195f
C4916 a_17405_2092# a_19307_1669# 2.12e-20
C4917 D2_1 P2 0.53f
C4918 a_1409_2253# D2_5 0.0784f
C4919 p2_gen_magic_0.xnor_magic_6.OUT D2_1 6.7e-19
C4920 p2_gen_magic_0.AND2_magic_1.A D2_2 0.00215f
C4921 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B p2_gen_magic_0.xnor_magic_3.OUT 1.55e-19
C4922 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT a_1957_n7648# 0.00157f
C4923 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B D2_6 0.00902f
C4924 a_5036_n8579# Q6 3.19e-19
C4925 a_24059_4877# D2_4 0.0541f
C4926 a_23985_7877# a_24185_7877# 0.519f
C4927 7b_counter_0.MDFF_6.tspc2_magic_0.Q Q6 0.197f
C4928 p3_gen_magic_0.xnor_magic_0.OUT D2_3 0.0073f
C4929 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A VDD 1.33f
C4930 a_1209_2253# a_2749_2092# 0.00114f
C4931 p2_gen_magic_0.xnor_magic_1.OUT a_11292_n6613# 1.57e-19
C4932 a_1209_3363# a_1409_3363# 0.298f
C4933 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT Q5 0.502f
C4934 p3_gen_magic_0.xnor_magic_1.B D2_5 0.00258f
C4935 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A Q3 0.00154f
C4936 a_8411_4513# a_8955_4557# 0.297f
C4937 p3_gen_magic_0.AND2_magic_1.A a_14556_n8142# 0.203f
C4938 a_19841_3363# Q3 1.54e-19
C4939 a_16386_n3644# Q4 0.0114f
C4940 p2_gen_magic_0.3_inp_AND_magic_0.B D2_5 6.85e-21
C4941 DFF_magic_0.tg_magic_3.CLK DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.0636f
C4942 a_15865_2253# D2_3 0.246f
C4943 a_15865_2253# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B 0.125f
C4944 a_1209_4557# 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 1.37e-19
C4945 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q5 0.00236f
C4946 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT a_1957_n3150# 6.1e-19
C4947 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_5.OUT 0.0149f
C4948 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A a_19841_4557# 0.251f
C4949 DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 4e-20
C4950 p3_gen_magic_0.xnor_magic_1.B p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT 0.00129f
C4951 p3_gen_magic_0.3_inp_AND_magic_0.A a_11708_n6613# 0.192f
C4952 OR_magic_2.VOUT divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT 0.00519f
C4953 p2_gen_magic_0.xnor_magic_3.OUT a_13553_n2115# 3.87e-19
C4954 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_24259_4877# 1.29e-19
C4955 VDD D2_1 8.91f
C4956 7b_counter_0.MDFF_4.tspc2_magic_0.D D2_2 0.139f
C4957 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_5385_2253# 0.017f
C4958 p2_gen_magic_0.xnor_magic_4.OUT D2_2 0.244f
C4959 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 8.78e-21
C4960 a_27778_4557# VDD 0.0579f
C4961 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5054_n6024# 0.0766f
C4962 a_8825_1669# D2_6 7.98e-19
C4963 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_3.OUT 2.3e-19
C4964 p3_gen_magic_0.xnor_magic_0.OUT a_8643_n6024# 0.415f
C4965 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B Q7 0.0259f
C4966 a_1409_2253# D2_7 0.00916f
C4967 a_16065_2253# D2_3 0.175f
C4968 7b_counter_0.MDFF_3.QB a_1209_9773# 0.231f
C4969 a_8523_n3597# D2_5 0.00322f
C4970 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT D2_4 0.049f
C4971 p2_gen_magic_0.3_inp_AND_magic_0.A p2_gen_magic_0.3_inp_AND_magic_0.B 0.318f
C4972 a_8523_n3150# p2_gen_magic_0.xnor_magic_6.OUT 0.0924f
C4973 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B 0.0303f
C4974 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B D2_2 0.00443f
C4975 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A Q1 0.0071f
C4976 VDD LD 20f
C4977 a_1957_n7648# a_1541_n8095# 0.013f
C4978 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B Q5 4.71e-19
C4979 a_30365_3514# OR_magic_1.VOUT 0.127f
C4980 a_19841_4557# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A 0.128f
C4981 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT 3.44e-20
C4982 p2_gen_magic_0.xnor_magic_5.OUT Q4 0.074f
C4983 a_9689_6886# a_9412_5956# 0.00164f
C4984 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A CLK 0.026f
C4985 p3_gen_magic_0.xnor_magic_1.B D2_7 0.24f
C4986 OR_magic_2.VOUT divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT 1.33f
C4987 a_24003_10051# VDD 0.0331f
C4988 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 0.0206f
C4989 p3_gen_magic_0.xnor_magic_0.OUT a_8523_n7648# 0.0374f
C4990 a_9212_739# a_9412_739# 0.651f
C4991 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 0.41f
C4992 Q3 P2 0.0165f
C4993 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT Q6 0.00782f
C4994 a_5036_n4081# p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 7.56e-21
C4995 LD D2_1 0.917f
C4996 a_1559_n6471# Q7 9.27e-19
C4997 7b_counter_0.MDFF_4.LD a_19841_3363# 0.195f
C4998 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A a_7215_10149# 0.397f
C4999 p2_gen_magic_0.xnor_magic_6.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 2.29e-19
C5000 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A Q2 0.111f
C5001 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_5185_6275# 0.223f
C5002 DFF_magic_0.D 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B 2.35e-19
C5003 a_5185_1059# Q4 0.00131f
C5004 DFF_magic_0.D a_30365_4922# 0.016f
C5005 a_17405_2092# D2_4 0.0108f
C5006 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q2 0.0142f
C5007 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT D2_3 4.44e-19
C5008 OR_magic_1.VOUT divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT 2.41e-19
C5009 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B a_15865_3363# 0.125f
C5010 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN D2_6 0.0267f
C5011 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 7b_counter_0.MDFF_4.tspc2_magic_0.Q 6.86e-19
C5012 p2_gen_magic_0.3_inp_AND_magic_0.VOUT D2_3 0.126f
C5013 a_1209_1059# Q5 2.91e-19
C5014 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT 1.05e-19
C5015 a_1559_n1973# Q7 0.042f
C5016 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_23258_1746# 4.65e-19
C5017 DFF_magic_0.D a_23985_7877# 1.36e-20
C5018 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B 0.0047f
C5019 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A 0.178f
C5020 a_24003_10051# LD 0.024f
C5021 a_8523_n3150# VDD 0.0014f
C5022 mux_magic_0.AND2_magic_0.A a_34156_n889# 3.58e-20
C5023 p3_gen_magic_0.3_inp_AND_magic_0.B p3_gen_magic_0.xnor_magic_1.OUT 0.0464f
C5024 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_0.IN 0.287f
C5025 a_9059_n1973# a_8523_n3597# 1.25e-19
C5026 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT 4e-20
C5027 a_4496_4393# D2_5 5.51e-20
C5028 a_2749_8740# a_4496_9609# 7.92e-19
C5029 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B 9.4e-20
C5030 a_17405_2092# a_17405_684# 0.475f
C5031 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD 1.09f
C5032 a_1209_2253# D2_5 0.049f
C5033 7b_counter_0.MDFF_5.tspc2_magic_0.D 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 8.78e-21
C5034 a_5054_n5540# D2_4 0.0212f
C5035 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A 0.178f
C5036 a_12387_1746# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B 0.125f
C5037 DFF_magic_0.tg_magic_2.IN DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.258f
C5038 a_12174_n8579# VDD 0.382f
C5039 VDD Q3 9.3f
C5040 mux_magic_0.IN1 P2 0.0475f
C5041 a_1541_n8579# Q6 1.74e-19
C5042 OR_magic_2.A P2 0.921f
C5043 7b_counter_0.MDFF_3.tspc2_magic_0.CLK CLK 0.048f
C5044 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A D2_4 0.0173f
C5045 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT VDD 1.03f
C5046 a_2749_8740# 7b_counter_0.MDFF_3.tspc2_magic_0.D 0.123f
C5047 p2_gen_magic_0.AND2_magic_1.A a_14556_n3644# 0.203f
C5048 D2_1 Q3 0.153f
C5049 7b_counter_0.MDFF_4.LD P2 0.00181f
C5050 a_1209_8579# D2_7 0.422f
C5051 a_15865_7470# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A 0.00184f
C5052 a_5385_7469# 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A 5.46e-20
C5053 a_20041_3363# a_20171_1669# 0.00565f
C5054 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT D2_6 0.0431f
C5055 p3_gen_magic_0.AND2_magic_1.A a_12174_n8095# 0.368f
C5056 a_15865_8580# a_16065_8580# 0.298f
C5057 a_14756_n3644# Q4 0.00317f
C5058 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_1 9.14e-19
C5059 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT Q1 0.0983f
C5060 7b_counter_0.MDFF_7.tspc2_magic_0.D VDD 1.39f
C5061 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_5.OUT 0.0155f
C5062 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A DFF_magic_0.tg_magic_3.CLK 7.43e-20
C5063 7b_counter_0.MDFF_1.tspc2_magic_0.D a_15865_1059# 1.63e-20
C5064 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT LD 0.00146f
C5065 a_5054_n5540# Q2 0.00454f
C5066 a_15865_2253# a_16065_2253# 0.298f
C5067 a_11292_n2115# Q5 7.55e-20
C5068 a_5054_n6024# a_5470_n6471# 0.0115f
C5069 a_1209_1059# Q2 2.43e-19
C5070 7b_counter_0.DFF_magic_0.tg_magic_3.CLK 7b_counter_0.DFF_magic_0.tg_magic_1.IN 0.0617f
C5071 a_20171_1669# Q1 0.00233f
C5072 LD Q3 0.0105f
C5073 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 0.4f
C5074 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B CLK 0.0139f
C5075 a_12931_6276# Q2 0.0298f
C5076 mux_magic_0.IN2 a_32616_n2458# 0.223f
C5077 p3_gen_magic_0.3_inp_AND_magic_0.A a_11492_n6613# 1.9e-20
C5078 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A Q4 8.78e-21
C5079 p2_gen_magic_0.xnor_magic_3.OUT a_11708_n2115# 0.0446f
C5080 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_24059_4877# 7.16e-19
C5081 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_2749_2092# 0.00137f
C5082 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN 4.63e-20
C5083 p3_gen_magic_0.xnor_magic_1.OUT D2_5 3.68e-19
C5084 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A a_16065_9774# 0.0292f
C5085 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT 0.96f
C5086 a_15865_3363# VDD 0.884f
C5087 mux_magic_0.IN1 VDD 6.48f
C5088 OR_magic_2.A VDD 5.4f
C5089 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT VDD 1.04f
C5090 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT a_27234_4513# 0.00721f
C5091 a_1209_2253# D2_7 0.0119f
C5092 a_5036_n3597# D2_5 0.0501f
C5093 a_26126_1124# 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 2.07e-19
C5094 p3_gen_magic_0.3_inp_AND_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 0.214f
C5095 a_8411_3319# Q6 1.47e-19
C5096 a_11292_n2115# D2_4 0.00766f
C5097 a_1957_n3150# a_1541_n3597# 0.013f
C5098 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT D2_3 0.0185f
C5099 7b_counter_0.MDFF_4.LD VDD 31f
C5100 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B a_11279_8697# 0.412f
C5101 DFF_magic_0.tg_magic_3.CLK DFF_magic_0.tg_magic_0.IN 0.164f
C5102 a_21504_5904# Q6 0.287f
C5103 7b_counter_0.DFF_magic_0.Q 7b_counter_0.DFF_magic_0.D 1.28f
C5104 mux_magic_0.IN1 D2_1 0.0522f
C5105 OR_magic_2.A D2_1 0.256f
C5106 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_5 0.0448f
C5107 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B a_2749_5900# 0.173f
C5108 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_20041_8580# 0.017f
C5109 a_5054_n1526# a_5470_n1973# 0.0115f
C5110 7b_counter_0.MDFF_3.QB VDD 5.29f
C5111 Q4 D2_6 3.19f
C5112 a_11292_n6613# p3_gen_magic_0.3_inp_AND_magic_0.B 0.00234f
C5113 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT D2_7 0.0459f
C5114 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.3_inp_AND_magic_0.C 0.00798f
C5115 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT VDD 1.04f
C5116 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD 1.08f
C5117 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.xnor_magic_5.OUT 1.38e-19
C5118 a_21381_8741# VDD 0.944f
C5119 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.OUT 0.0108f
C5120 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A a_12931_8580# 0.00103f
C5121 7b_counter_0.MDFF_3.QB D2_1 0.0532f
C5122 a_6725_2092# Q6 0.0744f
C5123 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B CLK 7.16e-20
C5124 7b_counter_0.MDFF_4.LD a_27778_4557# 0.00329f
C5125 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A Q5 0.273f
C5126 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_1 5.05e-21
C5127 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A a_17405_2092# 0.0334f
C5128 DFF_magic_0.D DFF_magic_0.tg_magic_2.OUT 0.0613f
C5129 a_13353_n2115# D2_3 0.0227f
C5130 a_8713_1625# a_9212_739# 0.299f
C5131 7b_counter_0.MDFF_3.QB LD 0.051f
C5132 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A a_20041_4557# 0.0292f
C5133 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.0211f
C5134 a_8713_6842# Q2 0.00818f
C5135 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B 0.178f
C5136 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT LD 1.39e-19
C5137 a_15865_6276# a_15865_4557# 0.00775f
C5138 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A Q2 0.053f
C5139 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8643_n5540# 0.0528f
C5140 a_21381_8741# LD 1.6e-20
C5141 a_5452_n3150# VDD 0.00519f
C5142 p3_gen_magic_0.xnor_magic_1.OUT D2_7 1.68f
C5143 a_5385_6275# Q7 0.00931f
C5144 7b_counter_0.MDFF_5.tspc2_magic_0.Q a_6725_7308# 0.00135f
C5145 a_27778_3363# D2_4 0.168f
C5146 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 4.28e-19
C5147 a_8643_n1973# a_8523_n3597# 3.68e-19
C5148 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A a_2749_684# 0.397f
C5149 a_7303_3480# a_5515_3947# 1.19e-20
C5150 a_12174_n3150# D2_2 3e-19
C5151 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A CLK 0.016f
C5152 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 0.00849f
C5153 a_5385_2253# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A 1.77e-19
C5154 7b_counter_0.MDFF_5.tspc2_magic_0.D a_9412_5956# 0.103f
C5155 a_5036_n3597# D2_7 0.243f
C5156 p2_gen_magic_0.AND2_magic_1.A p3_gen_magic_0.3_inp_AND_magic_0.C 5.66e-19
C5157 DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_1.IN 0.316f
C5158 a_15865_7470# 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 1.03e-19
C5159 a_8523_n8579# VDD 0.417f
C5160 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A 0.00112f
C5161 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_7 0.00216f
C5162 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 0.229f
C5163 a_27778_2253# a_27778_1059# 0.0206f
C5164 D2_2 Q4 0.472f
C5165 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN CLK 0.691f
C5166 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_8955_3363# 0.00751f
C5167 a_2749_10148# 7b_counter_0.MDFF_3.tspc2_magic_0.D 1.08e-19
C5168 a_11292_n6613# D2_5 0.0483f
C5169 OR_magic_1.VOUT divide_by_2_1.tg_magic_2.IN 0.00111f
C5170 p2_gen_magic_0.AND2_magic_1.A a_12174_n3597# 0.368f
C5171 p2_gen_magic_0.3_inp_AND_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT 0.708f
C5172 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A a_20041_4557# 9.27e-19
C5173 a_6725_5900# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B 4.85e-19
C5174 a_5054_n6471# p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT 5.8e-19
C5175 7b_counter_0.DFF_magic_0.D D2_4 0.0615f
C5176 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A Q6 0.0219f
C5177 a_2749_7308# 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A 2.07e-19
C5178 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B Q7 0.0163f
C5179 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A Q2 0.00117f
C5180 a_16186_n3644# Q4 0.0575f
C5181 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_12174_n8579# 0.0815f
C5182 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT Q4 8.46e-19
C5183 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT D2_6 2.34e-19
C5184 a_8643_n6471# Q5 3.78e-19
C5185 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A Q5 3.49e-19
C5186 7b_counter_0.MDFF_4.LD Q3 0.948f
C5187 a_23352_n5390# a_23352_n6798# 0.475f
C5188 a_5054_n6024# a_5054_n6471# 0.0137f
C5189 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_6.OUT 5.45e-19
C5190 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_19152_739# 0.35f
C5191 OR_magic_2.VOUT divide_by_2_0.tg_magic_1.IN 0.682f
C5192 a_19307_1669# Q1 0.00209f
C5193 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A Q1 0.00274f
C5194 7b_counter_0.MDFF_0.tspc2_magic_0.Q D2_5 0.214f
C5195 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT Q3 0.0062f
C5196 a_12387_5769# Q2 0.0294f
C5197 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_20041_9774# 0.12f
C5198 a_8523_n8095# Q5 0.0805f
C5199 p2_gen_magic_0.xnor_magic_3.OUT a_11492_n2115# 0.00138f
C5200 a_1209_6275# D2_7 0.00117f
C5201 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A 0.178f
C5202 a_6725_684# Q1 0.0075f
C5203 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK 1.83e-19
C5204 7b_counter_0.MDFF_4.tspc2_magic_0.Q a_11279_3480# 0.00137f
C5205 a_12387_3319# VDD 0.871f
C5206 a_27234_1746# VDD 0.87f
C5207 a_1559_n5540# a_1559_n6024# 0.0335f
C5208 p3_gen_magic_0.xnor_magic_5.OUT Q6 0.158f
C5209 a_23560_3728# VDD 0.774f
C5210 a_8939_n3150# D2_6 0.00157f
C5211 7b_counter_0.DFF_magic_0.tg_magic_0.IN VDD 1.18f
C5212 a_12590_n3150# D2_5 0.00223f
C5213 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT D2_4 1.42e-19
C5214 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A a_4235_3947# 3.22e-21
C5215 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B a_11191_10149# 0.173f
C5216 a_16065_8580# VDD 0.0173f
C5217 a_19152_5956# Q6 1.13e-20
C5218 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8939_n7648# 1.05e-19
C5219 a_32616_n1264# mux_magic_0.OR_magic_0.A 0.128f
C5220 a_5054_n1526# a_5054_n1973# 0.0137f
C5221 a_5185_7469# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A 0.00184f
C5222 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_1.OUT 0.00179f
C5223 a_8411_3319# a_8955_3363# 0.296f
C5224 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_1.IN 0.316f
C5225 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A VDD 1.23f
C5226 p3_gen_magic_0.xnor_magic_4.OUT a_5036_n7648# 0.0354f
C5227 divide_by_2_0.tg_magic_3.CLK VDD 4.16f
C5228 a_8955_8580# a_8713_6842# 5.39e-19
C5229 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B Q2 0.00493f
C5230 a_1559_n6024# Q7 5.03e-21
C5231 7b_counter_0.MDFF_4.LD a_15865_3363# 0.195f
C5232 a_5385_7469# CLK 0.00127f
C5233 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD 1.08f
C5234 7b_counter_0.MDFF_4.LD OR_magic_2.A 1.04f
C5235 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT D2_2 0.0174f
C5236 DFF_magic_0.tg_magic_3.CLK CLK 0.569f
C5237 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_3 1.35e-19
C5238 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A a_17405_7309# 0.0334f
C5239 a_11492_n6613# p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 5.63e-20
C5240 divide_by_2_0.tg_magic_3.CLK D2_1 0.0281f
C5241 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A Q2 0.0987f
C5242 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_8713_6842# 0.509f
C5243 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q2 0.00962f
C5244 a_12387_4513# 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A 0.251f
C5245 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A 0.00114f
C5246 7b_counter_0.MDFF_1.tspc2_magic_0.CLK CLK 0.119f
C5247 p2_gen_magic_0.3_inp_AND_magic_0.C p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK 0.0189f
C5248 p2_gen_magic_0.3_inp_AND_magic_0.B p2_gen_magic_0.AND2_magic_1.A 0.00753f
C5249 a_17405_3524# a_17405_2092# 0.00112f
C5250 a_1559_n1526# Q7 0.0526f
C5251 a_6725_2092# 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A 2.4e-20
C5252 7b_counter_0.MDFF_3.tspc2_magic_0.Q 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A 0.255f
C5253 7b_counter_0.MDFF_4.LD 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 6.05e-21
C5254 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT Q4 8.43e-19
C5255 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A 2.8e-19
C5256 CLK Q4 1.39f
C5257 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B a_6725_684# 0.173f
C5258 Q1 Q5 0.828f
C5259 a_5054_n6024# D2_3 0.231f
C5260 7b_counter_0.MDFF_7.tspc2_magic_0.CLK Q5 0.0124f
C5261 7b_counter_0.DFF_magic_0.Q 7b_counter_0.3_inp_AND_magic_0.VOUT 0.0989f
C5262 a_1541_n4081# Q7 0.00277f
C5263 a_11279_6341# Q2 0.129f
C5264 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT a_1541_n8579# 0.0846f
C5265 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_0.IN 0.0105f
C5266 a_1541_n7648# D2_7 4.29e-19
C5267 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1559_n1042# 0.057f
C5268 p2_gen_magic_0.xnor_magic_3.OUT D2_5 0.0413f
C5269 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT a_8939_n7648# 0.00157f
C5270 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1559_n5540# 0.0846f
C5271 a_5185_6275# Q7 0.0385f
C5272 a_12387_5769# a_12387_4513# 0.00775f
C5273 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A a_18891_6886# 3.22e-21
C5274 a_12387_552# p2_gen_magic_0.3_inp_AND_magic_0.A 5.12e-20
.ends

