* NGSPICE file created from mux_4x1_ibr_flat.ext - technology: gf180mcuC

.subckt mux_4x1_ibr_flat I1 I2 I3 S1 S0 OUT VDD VSS I0
X0 VDD S1.t0 mux_2x1_ibr_2.nand2_ibr_1.IN2 VDD.t19 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1 mux_2x1_ibr_1.nand2_ibr_2.IN2 S0.t0 VSS.t19 VSS.t18 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2 mux_2x1_ibr_2.I1 mux_2x1_ibr_1.nand2_ibr_1.IN2 VDD.t45 VDD.t44 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3 mux_2x1_ibr_1.nand2_ibr_2.OUT I2.t0 a_733_712# VSS.t5 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X4 VDD I2.t1 mux_2x1_ibr_1.nand2_ibr_2.OUT VDD.t4 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X5 mux_2x1_ibr_2.I0 mux_2x1_ibr_0.nand2_ibr_1.IN2 VDD.t43 VDD.t42 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X6 mux_2x1_ibr_2.nand2_ibr_2.IN2 S1.t1 VDD.t18 VDD.t17 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X7 mux_2x1_ibr_0.nand2_ibr_1.IN2 S0.t1 a_n956_1312# VSS.t17 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X8 VDD mux_2x1_ibr_2.nand2_ibr_2.OUT OUT.t1 VDD.t9 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X9 a_1859_712# mux_2x1_ibr_2.nand2_ibr_2.IN2 VSS.t11 VSS.t10 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X10 mux_2x1_ibr_2.nand2_ibr_2.OUT mux_2x1_ibr_2.nand2_ibr_2.IN2 VDD.t28 VDD.t27 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X11 OUT mux_2x1_ibr_2.nand2_ibr_1.IN2 VDD.t50 VDD.t49 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X12 a_n393_712# mux_2x1_ibr_0.nand2_ibr_2.IN2 VSS.t21 VSS.t20 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X13 mux_2x1_ibr_0.nand2_ibr_2.OUT mux_2x1_ibr_0.nand2_ibr_2.IN2 VDD.t38 VDD.t37 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X14 mux_2x1_ibr_2.nand2_ibr_1.IN2 mux_2x1_ibr_2.I1 VDD.t30 VDD.t29 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X15 mux_2x1_ibr_1.nand2_ibr_1.IN2 S0.t2 a_170_1312# VSS.t16 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X16 mux_2x1_ibr_2.I1 mux_2x1_ibr_1.nand2_ibr_2.OUT a_733_1312# VSS.t5 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X17 mux_2x1_ibr_0.nand2_ibr_2.IN2 S0.t3 VDD.t3 VDD.t2 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X18 mux_2x1_ibr_0.nand2_ibr_1.IN2 I1.t0 VDD.t23 VDD.t22 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X19 VDD mux_2x1_ibr_0.nand2_ibr_2.OUT mux_2x1_ibr_2.I0 VDD.t14 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X20 a_170_1312# I3.t0 VSS.t4 VSS.t3 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X21 mux_2x1_ibr_2.nand2_ibr_2.OUT mux_2x1_ibr_2.I0 a_1859_712# VSS.t2 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X22 VDD mux_2x1_ibr_2.I0 mux_2x1_ibr_2.nand2_ibr_2.OUT VDD.t31 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X23 mux_2x1_ibr_2.nand2_ibr_2.IN2 S1.t2 VSS.t9 VSS.t8 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X24 mux_2x1_ibr_2.nand2_ibr_1.IN2 S1.t3 a_1296_1312# VSS.t7 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X25 a_733_1312# mux_2x1_ibr_1.nand2_ibr_1.IN2 VSS.t25 VSS.t0 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X26 VDD S0.t4 mux_2x1_ibr_0.nand2_ibr_1.IN2 VDD.t34 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X27 a_n393_1312# mux_2x1_ibr_0.nand2_ibr_1.IN2 VSS.t24 VSS.t20 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X28 mux_2x1_ibr_0.nand2_ibr_2.IN2 S0.t5 VSS.t15 VSS.t14 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X29 a_733_712# mux_2x1_ibr_1.nand2_ibr_2.IN2 VSS.t1 VSS.t0 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X30 mux_2x1_ibr_1.nand2_ibr_2.OUT mux_2x1_ibr_1.nand2_ibr_2.IN2 VDD.t8 VDD.t7 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X31 OUT mux_2x1_ibr_2.nand2_ibr_2.OUT a_1859_1312# VSS.t2 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X32 a_1859_1312# mux_2x1_ibr_2.nand2_ibr_1.IN2 VSS.t26 VSS.t10 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X33 mux_2x1_ibr_1.nand2_ibr_2.IN2 S0.t6 VDD.t1 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X34 VDD mux_2x1_ibr_1.nand2_ibr_2.OUT mux_2x1_ibr_2.I1 VDD.t39 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X35 a_1296_1312# mux_2x1_ibr_2.I1 VSS.t13 VSS.t12 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X36 VDD S0.t7 mux_2x1_ibr_1.nand2_ibr_1.IN2 VDD.t46 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X37 VDD I0.t0 mux_2x1_ibr_0.nand2_ibr_2.OUT VDD.t24 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X38 mux_2x1_ibr_1.nand2_ibr_1.IN2 I3.t1 VDD.t13 VDD.t12 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X39 mux_2x1_ibr_0.nand2_ibr_2.OUT I0.t1 a_n393_712# VSS.t6 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X40 a_n956_1312# I1.t1 VSS.t23 VSS.t22 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X41 mux_2x1_ibr_2.I0 mux_2x1_ibr_0.nand2_ibr_2.OUT a_n393_1312# VSS.t6 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
R0 S1.n4 S1.t3 31.528
R1 S1.n1 S1.t1 25.7638
R2 S1.n4 S1.t0 15.3826
R3 S1.n1 S1.t2 13.2969
R4 S1.n5 S1.n4 7.62076
R5 S1.n7 S1.n6 4.54699
R6 S1.n3 S1 4.52833
R7 S1.n2 S1.n1 2.11815
R8 S1.n6 S1.n3 1.33848
R9 S1.n2 S1.n0 1.1266
R10 S1.n6 S1.n5 1.12145
R11 S1 S1.n7 0.0780197
R12 S1.n7 S1 0.0359098
R13 S1.n3 S1.n0 0.0344967
R14 S1.n0 S1 0.0125466
R15 S1.n5 S1 0.00197541
R16 S1 S1.n2 0.00142783
R17 VDD.t49 VDD.t19 763.259
R18 VDD.t39 VDD.t29 763.259
R19 VDD.t14 VDD.t12 763.259
R20 VDD.t34 VDD.t42 763.259
R21 VDD.n10 VDD.t27 386.348
R22 VDD.n36 VDD.t7 386.348
R23 VDD.n42 VDD.t37 386.348
R24 VDD.n10 VDD.t17 362.409
R25 VDD.n36 VDD.t0 362.409
R26 VDD.n42 VDD.t2 362.409
R27 VDD.n43 VDD.n42 319.75
R28 VDD.n37 VDD.n36 319.75
R29 VDD.n14 VDD.n10 319.75
R30 VDD.n19 VDD.t9 193.183
R31 VDD.n27 VDD.t19 193.183
R32 VDD.n28 VDD.t39 193.183
R33 VDD.n2 VDD.t46 193.183
R34 VDD.n4 VDD.t14 193.183
R35 VDD.n48 VDD.t34 193.183
R36 VDD.n9 VDD.t31 193.183
R37 VDD.n35 VDD.t4 193.183
R38 VDD.n41 VDD.t24 193.183
R39 VDD.n19 VDD.t49 109.849
R40 VDD.t29 VDD.n27 109.849
R41 VDD.n28 VDD.t44 109.849
R42 VDD.t12 VDD.n2 109.849
R43 VDD.t42 VDD.n4 109.849
R44 VDD.n48 VDD.t22 109.849
R45 VDD.t27 VDD.n9 109.849
R46 VDD.t7 VDD.n35 109.849
R47 VDD.t37 VDD.n41 109.849
R48 VDD.n15 VDD 11.7877
R49 VDD.n41 VDD.n40 6.3005
R50 VDD.n35 VDD.n34 6.3005
R51 VDD.n9 VDD.n8 6.3005
R52 VDD.n20 VDD.n19 6.3005
R53 VDD.n27 VDD.n26 6.3005
R54 VDD.n29 VDD.n28 6.3005
R55 VDD.n55 VDD.n2 6.3005
R56 VDD.n52 VDD.n4 6.3005
R57 VDD.n49 VDD.n48 6.3005
R58 VDD VDD.n18 5.23855
R59 VDD VDD.n7 5.23796
R60 VDD.n49 VDD.t23 5.21701
R61 VDD.n43 VDD.t3 5.19258
R62 VDD.n38 VDD.t1 5.14703
R63 VDD.n13 VDD.t18 5.14703
R64 VDD.n54 VDD.t13 5.13746
R65 VDD.n25 VDD.t30 5.13746
R66 VDD.n50 VDD.n47 5.13287
R67 VDD.n53 VDD.n3 5.13287
R68 VDD.n1 VDD.n0 5.13287
R69 VDD.n24 VDD.n23 5.13287
R70 VDD.n22 VDD.n6 5.13287
R71 VDD.n39 VDD.n5 5.13287
R72 VDD.n12 VDD.n11 5.13287
R73 VDD.n46 VDD.t43 3.91303
R74 VDD.n31 VDD.t45 3.91303
R75 VDD.n17 VDD.t50 3.91303
R76 VDD.n46 VDD.n45 3.87623
R77 VDD.n32 VDD.n31 3.87623
R78 VDD.n17 VDD.n16 3.87523
R79 VDD.n16 VDD.t28 3.51093
R80 VDD.n45 VDD.t38 3.51093
R81 VDD.n32 VDD.t8 3.51093
R82 VDD.n13 VDD.n12 0.852084
R83 VDD.n44 VDD 0.31523
R84 VDD.n33 VDD 0.31523
R85 VDD.n45 VDD.n44 0.272927
R86 VDD.n33 VDD.n32 0.272927
R87 VDD.n16 VDD.n15 0.272927
R88 VDD.n51 VDD.n46 0.22389
R89 VDD.n31 VDD.n30 0.22389
R90 VDD.n21 VDD.n17 0.22389
R91 VDD.n39 VDD.n38 0.197419
R92 VDD.n22 VDD.n21 0.141016
R93 VDD.n25 VDD.n24 0.141016
R94 VDD.n30 VDD.n1 0.141016
R95 VDD.n54 VDD.n53 0.141016
R96 VDD.n51 VDD.n50 0.141016
R97 VDD VDD.n22 0.106177
R98 VDD.n24 VDD 0.106177
R99 VDD VDD.n1 0.106177
R100 VDD.n53 VDD 0.106177
R101 VDD.n50 VDD 0.106177
R102 VDD VDD.n39 0.105597
R103 VDD.n12 VDD 0.105597
R104 VDD.n44 VDD.n40 0.0800484
R105 VDD.n34 VDD.n33 0.0800484
R106 VDD.n15 VDD.n8 0.0800484
R107 VDD.n21 VDD.n20 0.0800484
R108 VDD.n26 VDD.n25 0.0800484
R109 VDD.n30 VDD.n29 0.0800484
R110 VDD.n52 VDD.n51 0.0800484
R111 VDD VDD.n54 0.0788871
R112 VDD.n38 VDD.n37 0.0460556
R113 VDD.n14 VDD.n13 0.0460556
R114 VDD.n40 VDD 0.00166129
R115 VDD.n34 VDD 0.00166129
R116 VDD.n8 VDD 0.00166129
R117 VDD.n20 VDD 0.00166129
R118 VDD.n26 VDD 0.00166129
R119 VDD.n29 VDD 0.00166129
R120 VDD VDD.n55 0.00166129
R121 VDD.n55 VDD 0.00166129
R122 VDD VDD.n52 0.00166129
R123 VDD VDD.n49 0.00166129
R124 VDD VDD.n43 0.00105556
R125 VDD.n37 VDD 0.00105556
R126 VDD VDD.n14 0.00105556
R127 S0.n3 S0.t1 31.528
R128 S0.n0 S0.t2 31.528
R129 S0.n7 S0.t3 25.7638
R130 S0.n14 S0.t6 25.7638
R131 S0.n3 S0.t4 15.3826
R132 S0.n0 S0.t7 15.3826
R133 S0.n7 S0.t5 13.2969
R134 S0.n14 S0.t0 13.2969
R135 S0.n1 S0.n0 7.6289
R136 S0.n4 S0.n3 7.62076
R137 S0.n2 S0 4.53443
R138 S0.n9 S0 4.52833
R139 S0 S0.n13 4.52833
R140 S0.n12 S0.n11 2.19776
R141 S0.n8 S0.n7 2.11815
R142 S0.n15 S0.n14 2.11815
R143 S0.n5 S0.n4 1.5005
R144 S0.n10 S0.n9 1.31042
R145 S0.n13 S0.n12 1.28387
R146 S0.n8 S0.n6 1.1266
R147 S0.n16 S0.n15 1.1266
R148 S0.n12 S0.n1 0.948428
R149 S0.n1 S0 0.108522
R150 S0.n2 S0 0.0780742
R151 S0.n4 S0.n2 0.0373852
R152 S0.n11 S0.n10 0.0359098
R153 S0.n9 S0.n6 0.0344967
R154 S0.n16 S0.n13 0.0344967
R155 S0.n6 S0 0.0125466
R156 S0 S0.n16 0.0125466
R157 S0.n5 S0 0.00345082
R158 S0.n11 S0.n5 0.00197541
R159 S0 S0.n8 0.00142783
R160 S0.n15 S0 0.00142783
R161 VSS.t7 VSS.t10 1483.3
R162 VSS.t12 VSS.t5 1483.3
R163 VSS.t16 VSS.t0 1483.3
R164 VSS.t6 VSS.t3 1483.3
R165 VSS.t17 VSS.t20 1483.3
R166 VSS.n5 VSS.t2 353.341
R167 VSS.n11 VSS.t5 353.341
R168 VSS.n15 VSS.t6 353.341
R169 VSS.t10 VSS.n5 235.561
R170 VSS.n7 VSS.t12 235.561
R171 VSS.t0 VSS.n11 235.561
R172 VSS.t3 VSS.n14 235.561
R173 VSS.t20 VSS.n15 235.561
R174 VSS.n17 VSS.t22 235.561
R175 VSS.n16 VSS.t15 9.34566
R176 VSS.n2 VSS.t9 9.34566
R177 VSS.n0 VSS.t19 9.34566
R178 VSS VSS.t23 7.24801
R179 VSS.n21 VSS.t24 7.19156
R180 VSS.n21 VSS.t21 7.19156
R181 VSS.n4 VSS.t26 7.19156
R182 VSS.n4 VSS.t11 7.19156
R183 VSS.n9 VSS.t13 7.19156
R184 VSS.n10 VSS.t25 7.19156
R185 VSS.n10 VSS.t1 7.19156
R186 VSS.n22 VSS.t4 7.19156
R187 VSS.t8 VSS.t7 3.68113
R188 VSS.t18 VSS.t16 3.68113
R189 VSS.t14 VSS.t17 3.68113
R190 VSS.n13 VSS.n12 3.37613
R191 VSS.n8 VSS.n6 3.37613
R192 VSS.n19 VSS.n18 3.37613
R193 VSS VSS.n15 2.6035
R194 VSS.n11 VSS 2.6035
R195 VSS.n5 VSS 2.60269
R196 VSS.n18 VSS 2.6005
R197 VSS.n18 VSS.n17 2.6005
R198 VSS.n20 VSS.n19 2.6005
R199 VSS.n19 VSS.t14 2.6005
R200 VSS VSS.n8 2.6005
R201 VSS.n8 VSS.n7 2.6005
R202 VSS.n6 VSS.n3 2.6005
R203 VSS.n6 VSS.t8 2.6005
R204 VSS VSS.n13 2.6005
R205 VSS.n14 VSS.n13 2.6005
R206 VSS.n12 VSS.n1 2.6005
R207 VSS.n12 VSS.t18 2.6005
R208 VSS.n22 VSS 0.171522
R209 VSS VSS.n9 0.171522
R210 VSS.n21 VSS 0.113253
R211 VSS.n4 VSS 0.113253
R212 VSS.n10 VSS 0.113253
R213 VSS VSS.n21 0.0595367
R214 VSS VSS.n4 0.0595367
R215 VSS VSS.n10 0.0595367
R216 VSS.n9 VSS 0.0569474
R217 VSS VSS.n22 0.0569474
R218 VSS.n16 VSS 0.0340526
R219 VSS VSS.n2 0.0340526
R220 VSS VSS.n0 0.0340526
R221 VSS VSS.n20 0.0182632
R222 VSS VSS.n3 0.0182632
R223 VSS VSS.n1 0.0182632
R224 VSS VSS.n16 0.00405263
R225 VSS VSS.n2 0.00405263
R226 VSS.n0 VSS 0.00247368
R227 VSS.n20 VSS 0.000894737
R228 VSS.n3 VSS 0.000894737
R229 VSS.n1 VSS 0.000894737
R230 I2.n0 I2.t0 31.528
R231 I2.n0 I2.t1 15.3826
R232 I2.n1 I2.n0 8.74076
R233 I2 I2.n1 0.00507627
R234 I2.n1 I2 0.00202542
R235 OUT OUT.n2 7.15141
R236 OUT.n3 OUT.n1 3.2163
R237 OUT.n1 OUT.t1 2.2755
R238 OUT.n1 OUT.n0 2.2755
R239 OUT OUT.n3 0.035398
R240 OUT.n3 OUT 0.0119545
R241 I1.n0 I1.t0 30.9379
R242 I1.n0 I1.t1 21.6422
R243 I1 I1.n0 4.005
R244 I3.n0 I3.t1 30.9379
R245 I3.n0 I3.t0 21.6422
R246 I3 I3.n0 4.0005
R247 I0.n0 I0.t1 31.528
R248 I0.n0 I0.t0 15.3826
R249 I0 I0.n0 8.74076
C0 mux_2x1_ibr_1.nand2_ibr_1.IN2 I3 0.0959f
C1 S0 S1 0.00205f
C2 a_n393_712# mux_2x1_ibr_2.I0 1.5e-19
C3 mux_2x1_ibr_1.nand2_ibr_2.OUT mux_2x1_ibr_2.nand2_ibr_2.IN2 0.0112f
C4 a_733_1312# VDD 0.00444f
C5 mux_2x1_ibr_2.I0 mux_2x1_ibr_2.nand2_ibr_2.IN2 0.0646f
C6 VDD a_1859_712# 0.00444f
C7 mux_2x1_ibr_2.nand2_ibr_2.OUT a_1859_1312# 0.00949f
C8 VDD a_n393_1312# 0.00444f
C9 mux_2x1_ibr_2.I1 mux_2x1_ibr_2.nand2_ibr_1.IN2 0.11f
C10 a_1296_1312# mux_2x1_ibr_2.nand2_ibr_1.IN2 0.069f
C11 a_733_712# mux_2x1_ibr_1.nand2_ibr_2.OUT 0.0964f
C12 a_170_1312# mux_2x1_ibr_2.I0 0.00211f
C13 S0 mux_2x1_ibr_0.nand2_ibr_2.IN2 0.138f
C14 mux_2x1_ibr_2.nand2_ibr_2.IN2 S1 0.136f
C15 a_733_712# mux_2x1_ibr_2.I0 8.2e-19
C16 mux_2x1_ibr_1.nand2_ibr_2.IN2 a_733_712# 0.00372f
C17 VDD I1 0.146f
C18 S0 a_n393_712# 6.89e-19
C19 I2 mux_2x1_ibr_2.nand2_ibr_2.IN2 0.0036f
C20 VDD mux_2x1_ibr_1.nand2_ibr_2.OUT 0.666f
C21 I0 VDD 0.254f
C22 a_n956_1312# mux_2x1_ibr_0.nand2_ibr_1.IN2 0.069f
C23 a_733_1312# mux_2x1_ibr_1.nand2_ibr_1.IN2 0.00372f
C24 mux_2x1_ibr_2.nand2_ibr_2.OUT mux_2x1_ibr_2.nand2_ibr_1.IN2 0.053f
C25 a_n393_712# mux_2x1_ibr_0.nand2_ibr_2.IN2 0.00372f
C26 a_733_712# S1 2.15e-19
C27 VDD mux_2x1_ibr_2.I0 1.29f
C28 a_733_1312# mux_2x1_ibr_2.I1 0.069f
C29 VDD mux_2x1_ibr_1.nand2_ibr_2.IN2 0.402f
C30 mux_2x1_ibr_0.nand2_ibr_2.OUT a_n393_1312# 0.00949f
C31 I2 a_733_712# 0.00293f
C32 mux_2x1_ibr_2.nand2_ibr_1.IN2 a_1859_1312# 0.00372f
C33 S0 a_170_1312# 0.0151f
C34 S0 a_733_712# 2.62e-19
C35 VDD S1 0.595f
C36 mux_2x1_ibr_2.I0 OUT 5.19e-19
C37 I0 mux_2x1_ibr_0.nand2_ibr_2.OUT 0.202f
C38 I2 VDD 0.255f
C39 mux_2x1_ibr_1.nand2_ibr_2.OUT mux_2x1_ibr_1.nand2_ibr_1.IN2 0.053f
C40 mux_2x1_ibr_0.nand2_ibr_2.OUT mux_2x1_ibr_2.I0 0.63f
C41 mux_2x1_ibr_2.nand2_ibr_2.OUT a_1859_712# 0.0964f
C42 S0 VDD 1.57f
C43 mux_2x1_ibr_0.nand2_ibr_2.OUT mux_2x1_ibr_1.nand2_ibr_2.IN2 0.0112f
C44 mux_2x1_ibr_2.I1 mux_2x1_ibr_1.nand2_ibr_2.OUT 0.328f
C45 a_1296_1312# mux_2x1_ibr_1.nand2_ibr_2.OUT 9.43e-19
C46 S1 OUT 0.00946f
C47 mux_2x1_ibr_2.I0 mux_2x1_ibr_1.nand2_ibr_1.IN2 0.0169f
C48 mux_2x1_ibr_1.nand2_ibr_2.IN2 mux_2x1_ibr_1.nand2_ibr_1.IN2 0.00212f
C49 VDD mux_2x1_ibr_0.nand2_ibr_2.IN2 0.401f
C50 a_n393_1312# mux_2x1_ibr_0.nand2_ibr_1.IN2 0.00372f
C51 mux_2x1_ibr_2.I1 mux_2x1_ibr_2.I0 0.00147f
C52 a_1296_1312# mux_2x1_ibr_2.I0 1.04e-19
C53 VDD a_n393_712# 0.00444f
C54 S0 OUT 6.5e-20
C55 S1 mux_2x1_ibr_1.nand2_ibr_1.IN2 4.51e-21
C56 mux_2x1_ibr_0.nand2_ibr_1.IN2 I1 0.0959f
C57 VDD mux_2x1_ibr_2.nand2_ibr_2.IN2 0.402f
C58 mux_2x1_ibr_2.I1 S1 0.0593f
C59 a_1296_1312# S1 0.0144f
C60 S0 mux_2x1_ibr_0.nand2_ibr_2.OUT 0.0522f
C61 mux_2x1_ibr_2.nand2_ibr_2.OUT mux_2x1_ibr_2.I0 0.25f
C62 mux_2x1_ibr_0.nand2_ibr_1.IN2 mux_2x1_ibr_2.I0 0.109f
C63 S0 mux_2x1_ibr_1.nand2_ibr_1.IN2 0.378f
C64 I2 mux_2x1_ibr_2.I1 1.36e-19
C65 VDD a_170_1312# 3.14e-19
C66 mux_2x1_ibr_0.nand2_ibr_2.OUT mux_2x1_ibr_0.nand2_ibr_2.IN2 0.12f
C67 VDD a_733_712# 0.00444f
C68 S0 mux_2x1_ibr_2.I1 0.0109f
C69 mux_2x1_ibr_2.I0 a_1859_1312# 2.44e-19
C70 mux_2x1_ibr_0.nand2_ibr_2.OUT a_n393_712# 0.0964f
C71 mux_2x1_ibr_2.nand2_ibr_2.OUT S1 4.46e-19
C72 a_n956_1312# I1 0.00347f
C73 mux_2x1_ibr_2.I0 I3 0.0454f
C74 mux_2x1_ibr_2.nand2_ibr_1.IN2 mux_2x1_ibr_1.nand2_ibr_2.OUT 0.0106f
C75 S0 mux_2x1_ibr_0.nand2_ibr_1.IN2 0.368f
C76 mux_2x1_ibr_2.I0 mux_2x1_ibr_2.nand2_ibr_1.IN2 0.00155f
C77 a_170_1312# mux_2x1_ibr_1.nand2_ibr_1.IN2 0.069f
C78 mux_2x1_ibr_0.nand2_ibr_1.IN2 mux_2x1_ibr_0.nand2_ibr_2.IN2 0.00212f
C79 VDD OUT 0.234f
C80 mux_2x1_ibr_2.nand2_ibr_1.IN2 S1 0.341f
C81 mux_2x1_ibr_2.nand2_ibr_2.OUT mux_2x1_ibr_2.nand2_ibr_2.IN2 0.12f
C82 mux_2x1_ibr_0.nand2_ibr_2.OUT VDD 0.662f
C83 a_733_1312# mux_2x1_ibr_1.nand2_ibr_2.OUT 0.00949f
C84 S0 I3 0.0665f
C85 VDD mux_2x1_ibr_1.nand2_ibr_1.IN2 0.46f
C86 S0 a_n956_1312# 0.0144f
C87 a_733_1312# mux_2x1_ibr_2.I0 2.44e-19
C88 VDD mux_2x1_ibr_2.I1 0.423f
C89 VDD a_1296_1312# 3.14e-19
C90 S0 mux_2x1_ibr_2.nand2_ibr_1.IN2 4.45e-19
C91 mux_2x1_ibr_2.I0 a_1859_712# 0.00375f
C92 a_n393_1312# mux_2x1_ibr_2.I0 0.069f
C93 S1 a_1859_712# 2.62e-19
C94 mux_2x1_ibr_2.nand2_ibr_2.OUT VDD 0.634f
C95 mux_2x1_ibr_0.nand2_ibr_2.OUT mux_2x1_ibr_1.nand2_ibr_1.IN2 0.0102f
C96 VDD mux_2x1_ibr_0.nand2_ibr_1.IN2 0.456f
C97 mux_2x1_ibr_2.nand2_ibr_1.IN2 mux_2x1_ibr_2.nand2_ibr_2.IN2 0.00212f
C98 a_170_1312# I3 0.00347f
C99 mux_2x1_ibr_2.I0 mux_2x1_ibr_1.nand2_ibr_2.OUT 0.0242f
C100 I0 mux_2x1_ibr_2.I0 0.0148f
C101 I0 mux_2x1_ibr_1.nand2_ibr_2.IN2 0.0036f
C102 mux_2x1_ibr_1.nand2_ibr_2.IN2 mux_2x1_ibr_1.nand2_ibr_2.OUT 0.12f
C103 VDD a_1859_1312# 0.00444f
C104 mux_2x1_ibr_2.I1 mux_2x1_ibr_1.nand2_ibr_1.IN2 0.109f
C105 mux_2x1_ibr_1.nand2_ibr_2.IN2 mux_2x1_ibr_2.I0 0.019f
C106 S0 a_n393_1312# 9.5e-19
C107 mux_2x1_ibr_2.nand2_ibr_2.OUT OUT 0.303f
C108 mux_2x1_ibr_2.I1 a_1296_1312# 0.00372f
C109 mux_2x1_ibr_1.nand2_ibr_2.OUT S1 0.108f
C110 VDD I3 0.153f
C111 mux_2x1_ibr_2.I0 S1 0.0157f
C112 a_1859_1312# OUT 0.069f
C113 a_n956_1312# VDD 3.14e-19
C114 mux_2x1_ibr_0.nand2_ibr_2.OUT mux_2x1_ibr_0.nand2_ibr_1.IN2 0.053f
C115 S0 I1 0.0576f
C116 mux_2x1_ibr_1.nand2_ibr_2.IN2 S1 3.65e-19
C117 I2 mux_2x1_ibr_1.nand2_ibr_2.OUT 0.202f
C118 VDD mux_2x1_ibr_2.nand2_ibr_1.IN2 0.461f
C119 S0 mux_2x1_ibr_1.nand2_ibr_2.OUT 0.00113f
C120 S0 I0 0.00438f
C121 mux_2x1_ibr_2.nand2_ibr_2.IN2 a_1859_712# 0.00372f
C122 I2 mux_2x1_ibr_2.I0 0.0101f
C123 I2 mux_2x1_ibr_1.nand2_ibr_2.IN2 0.0473f
C124 I0 mux_2x1_ibr_0.nand2_ibr_2.IN2 0.0473f
C125 S0 mux_2x1_ibr_2.I0 0.198f
C126 S0 mux_2x1_ibr_1.nand2_ibr_2.IN2 0.136f
C127 mux_2x1_ibr_2.I0 mux_2x1_ibr_0.nand2_ibr_2.IN2 0.0048f
C128 I0 a_n393_712# 0.00293f
C129 mux_2x1_ibr_0.nand2_ibr_2.OUT I3 0.0174f
C130 I2 S1 0.00408f
C131 mux_2x1_ibr_2.nand2_ibr_1.IN2 OUT 0.109f
C132 a_1859_712# VSS 0.0676f
C133 mux_2x1_ibr_2.nand2_ibr_2.IN2 VSS 0.422f
C134 a_733_712# VSS 0.0676f
C135 I2 VSS 0.232f
C136 mux_2x1_ibr_1.nand2_ibr_2.IN2 VSS 0.422f
C137 a_n393_712# VSS 0.0676f
C138 I0 VSS 0.232f
C139 mux_2x1_ibr_0.nand2_ibr_2.IN2 VSS 0.437f
C140 a_1859_1312# VSS 0.0676f
C141 a_1296_1312# VSS 0.0676f
C142 a_733_1312# VSS 0.0676f
C143 a_170_1312# VSS 0.0676f
C144 a_n393_1312# VSS 0.0676f
C145 a_n956_1312# VSS 0.0678f
C146 OUT VSS 0.14f
C147 mux_2x1_ibr_2.I0 VSS 1.1f
C148 mux_2x1_ibr_2.nand2_ibr_2.OUT VSS 0.651f
C149 mux_2x1_ibr_2.nand2_ibr_1.IN2 VSS 0.412f
C150 S1 VSS 0.702f
C151 mux_2x1_ibr_2.I1 VSS 0.416f
C152 mux_2x1_ibr_1.nand2_ibr_2.OUT VSS 0.489f
C153 mux_2x1_ibr_1.nand2_ibr_1.IN2 VSS 0.412f
C154 I3 VSS 0.257f
C155 mux_2x1_ibr_0.nand2_ibr_2.OUT VSS 0.437f
C156 mux_2x1_ibr_0.nand2_ibr_1.IN2 VSS 0.435f
C157 S0 VSS 1.75f
C158 I1 VSS 0.292f
C159 VDD VSS 12.3f
.ends

