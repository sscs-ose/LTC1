magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -932 -1968 16833 52982
use M2_M1_CDNS_6903358316533  M2_M1_CDNS_6903358316533_0
timestamp 1713338890
transform 1 0 14795 0 1 35896
box -38 -686 38 686
use M2_M1_CDNS_6903358316533  M2_M1_CDNS_6903358316533_1
timestamp 1713338890
transform 1 0 14795 0 1 50296
box -38 -686 38 686
use M3_M2_CDNS_6903358316534  M3_M2_CDNS_6903358316534_0
timestamp 1713338890
transform 1 0 14795 0 1 35896
box -38 -686 38 686
use M3_M2_CDNS_6903358316534  M3_M2_CDNS_6903358316534_1
timestamp 1713338890
transform 1 0 14795 0 1 50296
box -38 -686 38 686
use M3_M2_CDNS_69033583165370  M3_M2_CDNS_69033583165370_0
timestamp 1713338890
transform 1 0 1602 0 1 10296
box -534 -658 534 658
use M3_M2_CDNS_69033583165370  M3_M2_CDNS_69033583165370_1
timestamp 1713338890
transform 1 0 6892 0 1 11896
box -534 -658 534 658
use M3_M2_CDNS_69033583165370  M3_M2_CDNS_69033583165370_2
timestamp 1713338890
transform 1 0 8086 0 1 10296
box -534 -658 534 658
use M3_M2_CDNS_69033583165370  M3_M2_CDNS_69033583165370_3
timestamp 1713338890
transform 1 0 13376 0 1 11896
box -534 -658 534 658
use M3_M2_CDNS_69033583165370  M3_M2_CDNS_69033583165370_4
timestamp 1713338890
transform 1 0 6892 0 1 26296
box -534 -658 534 658
use M3_M2_CDNS_69033583165370  M3_M2_CDNS_69033583165370_5
timestamp 1713338890
transform 1 0 8086 0 1 27896
box -534 -658 534 658
use M3_M2_CDNS_69033583165370  M3_M2_CDNS_69033583165370_6
timestamp 1713338890
transform 1 0 13376 0 1 26296
box -534 -658 534 658
use M3_M2_CDNS_69033583165370  M3_M2_CDNS_69033583165370_7
timestamp 1713338890
transform 1 0 8086 0 1 40696
box -534 -658 534 658
use M3_M2_CDNS_69033583165370  M3_M2_CDNS_69033583165370_8
timestamp 1713338890
transform 1 0 8086 0 1 39096
box -534 -658 534 658
use M3_M2_CDNS_69033583165370  M3_M2_CDNS_69033583165370_9
timestamp 1713338890
transform 1 0 8086 0 1 42296
box -534 -658 534 658
use M3_M2_CDNS_69033583165370  M3_M2_CDNS_69033583165370_10
timestamp 1713338890
transform 1 0 13376 0 1 43896
box -534 -658 534 658
use M3_M2_CDNS_69033583165371  M3_M2_CDNS_69033583165371_0
timestamp 1713338890
transform 1 0 6892 0 1 4696
box -534 -1464 534 1464
use M3_M2_CDNS_69033583165371  M3_M2_CDNS_69033583165371_1
timestamp 1713338890
transform 1 0 6892 0 1 1496
box -534 -1464 534 1464
use M3_M2_CDNS_69033583165371  M3_M2_CDNS_69033583165371_2
timestamp 1713338890
transform 1 0 13376 0 1 4696
box -534 -1464 534 1464
use M3_M2_CDNS_69033583165371  M3_M2_CDNS_69033583165371_3
timestamp 1713338890
transform 1 0 13376 0 1 1496
box -534 -1464 534 1464
use M3_M2_CDNS_69033583165371  M3_M2_CDNS_69033583165371_4
timestamp 1713338890
transform 1 0 6892 0 1 7896
box -534 -1464 534 1464
use M3_M2_CDNS_69033583165371  M3_M2_CDNS_69033583165371_5
timestamp 1713338890
transform 1 0 13376 0 1 7896
box -534 -1464 534 1464
use M3_M2_CDNS_69033583165371  M3_M2_CDNS_69033583165371_6
timestamp 1713338890
transform 1 0 1602 0 1 17496
box -534 -1464 534 1464
use M3_M2_CDNS_69033583165371  M3_M2_CDNS_69033583165371_7
timestamp 1713338890
transform 1 0 1602 0 1 14296
box -534 -1464 534 1464
use M3_M2_CDNS_69033583165371  M3_M2_CDNS_69033583165371_8
timestamp 1713338890
transform 1 0 8086 0 1 17496
box -534 -1464 534 1464
use M3_M2_CDNS_69033583165371  M3_M2_CDNS_69033583165371_9
timestamp 1713338890
transform 1 0 8086 0 1 14296
box -534 -1464 534 1464
use M3_M2_CDNS_69033583165371  M3_M2_CDNS_69033583165371_10
timestamp 1713338890
transform 1 0 1602 0 1 20696
box -534 -1464 534 1464
use M3_M2_CDNS_69033583165371  M3_M2_CDNS_69033583165371_11
timestamp 1713338890
transform 1 0 8086 0 1 20696
box -534 -1464 534 1464
use M3_M2_CDNS_69033583165371  M3_M2_CDNS_69033583165371_12
timestamp 1713338890
transform 1 0 1602 0 1 23896
box -534 -1464 534 1464
use M3_M2_CDNS_69033583165371  M3_M2_CDNS_69033583165371_13
timestamp 1713338890
transform 1 0 8086 0 1 23896
box -534 -1464 534 1464
use M3_M2_CDNS_69033583165371  M3_M2_CDNS_69033583165371_14
timestamp 1713338890
transform 1 0 6892 0 1 33496
box -534 -1464 534 1464
use M3_M2_CDNS_69033583165371  M3_M2_CDNS_69033583165371_15
timestamp 1713338890
transform 1 0 8086 0 1 30296
box -534 -1464 534 1464
use M3_M2_CDNS_69033583165371  M3_M2_CDNS_69033583165371_16
timestamp 1713338890
transform 1 0 13376 0 1 33496
box -534 -1464 534 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_0
timestamp 1713338890
transform 1 0 3403 0 1 4696
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_1
timestamp 1713338890
transform 1 0 3403 0 1 1496
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_2
timestamp 1713338890
transform 1 0 9647 0 1 1496
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_3
timestamp 1713338890
transform 1 0 9647 0 1 4696
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_4
timestamp 1713338890
transform 1 0 3403 0 1 7896
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_5
timestamp 1713338890
transform 1 0 9647 0 1 7896
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_6
timestamp 1713338890
transform 1 0 5331 0 1 14296
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_7
timestamp 1713338890
transform 1 0 5331 0 1 17496
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_8
timestamp 1713338890
transform 1 0 11575 0 1 17496
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_9
timestamp 1713338890
transform 1 0 11575 0 1 14296
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_10
timestamp 1713338890
transform 1 0 5331 0 1 20696
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_11
timestamp 1713338890
transform 1 0 11575 0 1 20696
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_12
timestamp 1713338890
transform 1 0 5331 0 1 23896
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_13
timestamp 1713338890
transform 1 0 11575 0 1 23896
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_14
timestamp 1713338890
transform 1 0 5331 0 1 30296
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_15
timestamp 1713338890
transform 1 0 9647 0 1 33496
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165372  M3_M2_CDNS_69033583165372_16
timestamp 1713338890
transform 1 0 11575 0 1 30296
box -906 -1464 906 1464
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_0
timestamp 1713338890
transform 1 0 3403 0 1 11896
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_1
timestamp 1713338890
transform 1 0 5331 0 1 10296
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_2
timestamp 1713338890
transform 1 0 9647 0 1 11896
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_3
timestamp 1713338890
transform 1 0 11575 0 1 10296
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_4
timestamp 1713338890
transform 1 0 3403 0 1 26296
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_5
timestamp 1713338890
transform 1 0 5331 0 1 27896
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_6
timestamp 1713338890
transform 1 0 9647 0 1 26296
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_7
timestamp 1713338890
transform 1 0 11575 0 1 27896
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_8
timestamp 1713338890
transform 1 0 11575 0 1 40696
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_9
timestamp 1713338890
transform 1 0 11575 0 1 39096
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_10
timestamp 1713338890
transform 1 0 9647 0 1 43896
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_11
timestamp 1713338890
transform 1 0 11575 0 1 42296
box -906 -658 906 658
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_0
timestamp 1713338890
transform 1 0 1527 0 1 28088
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_1
timestamp 1713338890
transform 1 0 4622 0 1 40831
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_2
timestamp 1713338890
transform 1 0 4498 0 1 40955
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_3
timestamp 1713338890
transform 1 0 5118 0 1 40335
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_4
timestamp 1713338890
transform 1 0 4994 0 1 40459
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_5
timestamp 1713338890
transform 1 0 4870 0 1 40583
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_6
timestamp 1713338890
transform 1 0 5614 0 1 39839
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_7
timestamp 1713338890
transform 1 0 5490 0 1 39963
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_8
timestamp 1713338890
transform 1 0 5366 0 1 40087
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_9
timestamp 1713338890
transform 1 0 5242 0 1 40211
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_10
timestamp 1713338890
transform 1 0 5986 0 1 39467
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_11
timestamp 1713338890
transform 1 0 5862 0 1 39591
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_12
timestamp 1713338890
transform 1 0 5738 0 1 39715
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_13
timestamp 1713338890
transform 1 0 6110 0 1 39343
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_14
timestamp 1713338890
transform 1 0 4746 0 1 40707
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_15
timestamp 1713338890
transform 1 0 4498 0 1 43190
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_16
timestamp 1713338890
transform 1 0 4622 0 1 43066
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_17
timestamp 1713338890
transform 1 0 4622 0 1 45365
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_18
timestamp 1713338890
transform 1 0 4870 0 1 42818
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_19
timestamp 1713338890
transform 1 0 4746 0 1 42942
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_20
timestamp 1713338890
transform 1 0 5118 0 1 42570
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_21
timestamp 1713338890
transform 1 0 4994 0 1 42694
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_22
timestamp 1713338890
transform 1 0 5242 0 1 42446
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_23
timestamp 1713338890
transform 1 0 5366 0 1 42322
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_24
timestamp 1713338890
transform 1 0 5490 0 1 42198
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_25
timestamp 1713338890
transform 1 0 5614 0 1 42074
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_26
timestamp 1713338890
transform 1 0 5738 0 1 41950
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_27
timestamp 1713338890
transform 1 0 5862 0 1 41826
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_28
timestamp 1713338890
transform 1 0 5986 0 1 41702
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_29
timestamp 1713338890
transform 1 0 6110 0 1 41578
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_30
timestamp 1713338890
transform 1 0 5366 0 1 44621
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_31
timestamp 1713338890
transform 1 0 5614 0 1 44373
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_32
timestamp 1713338890
transform 1 0 5490 0 1 44497
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_33
timestamp 1713338890
transform 1 0 5738 0 1 44249
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_34
timestamp 1713338890
transform 1 0 5862 0 1 44125
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_35
timestamp 1713338890
transform 1 0 5986 0 1 44001
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_36
timestamp 1713338890
transform 1 0 6110 0 1 43877
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_37
timestamp 1713338890
transform 1 0 4870 0 1 45117
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_38
timestamp 1713338890
transform 1 0 4746 0 1 45241
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_39
timestamp 1713338890
transform 1 0 5118 0 1 44869
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_40
timestamp 1713338890
transform 1 0 4994 0 1 44993
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_41
timestamp 1713338890
transform 1 0 5242 0 1 44745
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_42
timestamp 1713338890
transform 1 0 6918 0 1 45340
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_43
timestamp 1713338890
transform 1 0 7290 0 1 44968
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_44
timestamp 1713338890
transform 1 0 7042 0 1 45216
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_45
timestamp 1713338890
transform 1 0 7166 0 1 45092
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_46
timestamp 1713338890
transform 1 0 4498 0 1 45489
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_47
timestamp 1713338890
transform 1 0 6422 0 1 45836
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_48
timestamp 1713338890
transform 1 0 6794 0 1 45464
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_49
timestamp 1713338890
transform 1 0 6546 0 1 45712
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_50
timestamp 1713338890
transform 1 0 6670 0 1 45588
box -38 -844 38 844
use M3_M2_CDNS_69033583165375  M3_M2_CDNS_69033583165375_0
timestamp 1713338890
transform 1 0 1899 0 1 27891
box -38 -658 38 658
use M3_M2_CDNS_69033583165375  M3_M2_CDNS_69033583165375_1
timestamp 1713338890
transform 1 0 2023 0 1 27889
box -38 -658 38 658
use M3_M2_CDNS_69033583165376  M3_M2_CDNS_69033583165376_0
timestamp 1713338890
transform 1 0 1651 0 1 28036
box -38 -782 38 782
use M3_M2_CDNS_69033583165377  M3_M2_CDNS_69033583165377_0
timestamp 1713338890
transform 1 0 1775 0 1 27943
box -38 -720 38 720
use M3_M2_CDNS_69033583165378  M3_M2_CDNS_69033583165378_0
timestamp 1713338890
transform 1 0 3671 0 1 33925
box -38 -1898 38 1898
use M3_M2_CDNS_69033583165379  M3_M2_CDNS_69033583165379_0
timestamp 1713338890
transform 1 0 3547 0 1 33996
box -38 -1960 38 1960
use M3_M2_CDNS_69033583165380  M3_M2_CDNS_69033583165380_0
timestamp 1713338890
transform 1 0 1555 0 1 31382
box -38 -2022 38 2022
use M3_M2_CDNS_69033583165380  M3_M2_CDNS_69033583165380_1
timestamp 1713338890
transform 1 0 1803 0 1 31134
box -38 -2022 38 2022
use M3_M2_CDNS_69033583165380  M3_M2_CDNS_69033583165380_2
timestamp 1713338890
transform 1 0 1679 0 1 31258
box -38 -2022 38 2022
use M3_M2_CDNS_69033583165380  M3_M2_CDNS_69033583165380_3
timestamp 1713338890
transform 1 0 1431 0 1 31506
box -38 -2022 38 2022
use M3_M2_CDNS_69033583165380  M3_M2_CDNS_69033583165380_4
timestamp 1713338890
transform 1 0 1307 0 1 31630
box -38 -2022 38 2022
use M3_M2_CDNS_69033583165380  M3_M2_CDNS_69033583165380_5
timestamp 1713338890
transform 1 0 2051 0 1 30886
box -38 -2022 38 2022
use M3_M2_CDNS_69033583165380  M3_M2_CDNS_69033583165380_6
timestamp 1713338890
transform 1 0 1927 0 1 31010
box -38 -2022 38 2022
use M3_M2_CDNS_69033583165380  M3_M2_CDNS_69033583165380_7
timestamp 1713338890
transform 1 0 1183 0 1 31754
box -38 -2022 38 2022
use M3_M2_CDNS_69033583165380  M3_M2_CDNS_69033583165380_8
timestamp 1713338890
transform 1 0 3299 0 1 34244
box -38 -2022 38 2022
use M3_M2_CDNS_69033583165380  M3_M2_CDNS_69033583165380_9
timestamp 1713338890
transform 1 0 3423 0 1 34120
box -38 -2022 38 2022
use M3_M2_CDNS_69033583165380  M3_M2_CDNS_69033583165380_10
timestamp 1713338890
transform 1 0 3175 0 1 34368
box -38 -2022 38 2022
use M3_M2_CDNS_69033583165380  M3_M2_CDNS_69033583165380_11
timestamp 1713338890
transform 1 0 2803 0 1 34740
box -38 -2022 38 2022
use M3_M2_CDNS_69033583165380  M3_M2_CDNS_69033583165380_12
timestamp 1713338890
transform 1 0 2679 0 1 34864
box -38 -2022 38 2022
use M3_M2_CDNS_69033583165380  M3_M2_CDNS_69033583165380_13
timestamp 1713338890
transform 1 0 2555 0 1 34988
box -38 -2022 38 2022
use M3_M2_CDNS_69033583165380  M3_M2_CDNS_69033583165380_14
timestamp 1713338890
transform 1 0 3051 0 1 34492
box -38 -2022 38 2022
use M3_M2_CDNS_69033583165380  M3_M2_CDNS_69033583165380_15
timestamp 1713338890
transform 1 0 2927 0 1 34616
box -38 -2022 38 2022
use M3_M2_CDNS_69033583165381  M3_M2_CDNS_69033583165381_0
timestamp 1713338890
transform 1 0 1155 0 1 28411
box -38 -906 38 906
use M3_M2_CDNS_69033583165381  M3_M2_CDNS_69033583165381_1
timestamp 1713338890
transform 1 0 1279 0 1 28287
box -38 -906 38 906
use M3_M2_CDNS_69033583165381  M3_M2_CDNS_69033583165381_2
timestamp 1713338890
transform 1 0 1403 0 1 28163
box -38 -906 38 906
use M3_M2_CDNS_69033583165381  M3_M2_CDNS_69033583165381_3
timestamp 1713338890
transform 1 0 1132 0 1 44359
box -38 -906 38 906
use M3_M2_CDNS_69033583165381  M3_M2_CDNS_69033583165381_4
timestamp 1713338890
transform 1 0 2000 0 1 43491
box -38 -906 38 906
use M3_M2_CDNS_69033583165381  M3_M2_CDNS_69033583165381_5
timestamp 1713338890
transform 1 0 1504 0 1 43987
box -38 -906 38 906
use M3_M2_CDNS_69033583165381  M3_M2_CDNS_69033583165381_6
timestamp 1713338890
transform 1 0 1628 0 1 43863
box -38 -906 38 906
use M3_M2_CDNS_69033583165381  M3_M2_CDNS_69033583165381_7
timestamp 1713338890
transform 1 0 1752 0 1 43739
box -38 -906 38 906
use M3_M2_CDNS_69033583165381  M3_M2_CDNS_69033583165381_8
timestamp 1713338890
transform 1 0 1876 0 1 43615
box -38 -906 38 906
use M3_M2_CDNS_69033583165381  M3_M2_CDNS_69033583165381_9
timestamp 1713338890
transform 1 0 1256 0 1 44235
box -38 -906 38 906
use M3_M2_CDNS_69033583165381  M3_M2_CDNS_69033583165381_10
timestamp 1713338890
transform 1 0 1380 0 1 44111
box -38 -906 38 906
use M3_M2_CDNS_69033583165382  M3_M2_CDNS_69033583165382_0
timestamp 1713338890
transform 1 0 4167 0 1 33715
box -38 -1712 38 1712
use M3_M2_CDNS_69033583165383  M3_M2_CDNS_69033583165383_0
timestamp 1713338890
transform 1 0 4043 0 1 33771
box -38 -1774 38 1774
use M3_M2_CDNS_69033583165383  M3_M2_CDNS_69033583165383_1
timestamp 1713338890
transform 1 0 3919 0 1 33842
box -38 -1774 38 1774
use M3_M2_CDNS_69033583165384  M3_M2_CDNS_69033583165384_0
timestamp 1713338890
transform 1 0 3795 0 1 33884
box -38 -1836 38 1836
<< end >>
