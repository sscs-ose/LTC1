magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2541 -2045 2541 2045
<< psubdiff >>
rect -541 23 541 45
rect -541 -23 -519 23
rect -473 -23 -395 23
rect -349 -23 -271 23
rect -225 -23 -147 23
rect -101 -23 -23 23
rect 23 -23 101 23
rect 147 -23 225 23
rect 271 -23 349 23
rect 395 -23 473 23
rect 519 -23 541 23
rect -541 -45 541 -23
<< psubdiffcont >>
rect -519 -23 -473 23
rect -395 -23 -349 23
rect -271 -23 -225 23
rect -147 -23 -101 23
rect -23 -23 23 23
rect 101 -23 147 23
rect 225 -23 271 23
rect 349 -23 395 23
rect 473 -23 519 23
<< metal1 >>
rect -530 23 530 34
rect -530 -23 -519 23
rect -473 -23 -395 23
rect -349 -23 -271 23
rect -225 -23 -147 23
rect -101 -23 -23 23
rect 23 -23 101 23
rect 147 -23 225 23
rect 271 -23 349 23
rect 395 -23 473 23
rect 519 -23 530 23
rect -530 -34 530 -23
<< end >>
