* NGSPICE file created from Mux2x1_flat.ext - technology: gf180mcuC

.subckt pex_Mux2x1 VDD VSS A B SEL OUT
X0 a_672_1152# B.t0 VSS.t1 VSS.t0 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X1 a_268_215# A.t0 VSS.t5 VSS.t4 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X2 AND_0.B SEL.t0 VDD.t12 VDD.t11 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X3 VDD SEL.t1 AND_1.Inverter_0.IN VDD.t8 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X4 OR_0.Inverter_0.IN OR_0.B VSS.t12 VSS.t11 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X5 AND_0.Inverter_0.IN AND_0.B a_672_1152# VSS.t13 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X6 AND_0.B SEL.t2 VSS.t3 VSS.t2 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X7 a_1557_553# OR_0.A OR_0.Inverter_0.IN VDD.t23 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X8 OR_0.Inverter_0.IN OR_0.A VSS.t17 VSS.t16 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X9 OR_0.A AND_0.Inverter_0.IN VDD.t21 VDD.t20 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X10 OUT OR_0.Inverter_0.IN VDD.t7 VDD.t6 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X11 a_1557_553# OR_0.B VDD.t17 VDD.t16 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X12 AND_0.Inverter_0.IN B.t1 VDD.t1 VDD.t0 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X13 OR_0.B AND_1.Inverter_0.IN VDD.t3 VDD.t2 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X14 AND_1.Inverter_0.IN SEL.t3 a_268_215# VSS.t10 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X15 AND_1.Inverter_0.IN A.t1 VDD.t5 VDD.t4 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X16 OR_0.A AND_0.Inverter_0.IN VSS.t15 VSS.t14 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X17 OUT OR_0.Inverter_0.IN VSS.t9 VSS.t8 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X18 VDD OR_0.B a_1557_553# VDD.t13 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X19 VDD AND_0.B AND_0.Inverter_0.IN VDD.t0 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X20 OR_0.B AND_1.Inverter_0.IN VSS.t7 VSS.t6 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X21 OR_0.Inverter_0.IN OR_0.A a_1557_553# VDD.t22 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
R0 B.n0 B.t0 31.938
R1 B.n1 B.n0 29.9741
R2 B.n0 B.t1 12.2541
R3 B B.n1 3.09278
R4 B B.n2 2.264
R5 B.n1 B 0.00183811
R6 VSS.t4 VSS.n22 11315.1
R7 VSS.n7 VSS.t11 3284.06
R8 VSS.n1 VSS.t16 2649.77
R9 VSS.n17 VSS.n16 1755.05
R10 VSS.n6 VSS.t16 1537.16
R11 VSS.t10 VSS.n8 1475.28
R12 VSS.t0 VSS.n13 1462.13
R13 VSS.t11 VSS.n6 1420.05
R14 VSS.n18 VSS.t13 1410.64
R15 VSS.n18 VSS.t0 1382.98
R16 VSS.n22 VSS.n13 1071.17
R17 VSS VSS.n1 934.77
R18 VSS.n15 VSS.t14 603.342
R19 VSS.n7 VSS.t6 498.764
R20 VSS.n1 VSS.t8 426.344
R21 VSS.n13 VSS.t2 414.541
R22 VSS.n8 VSS.n7 80.4465
R23 VSS.n23 VSS.t4 80.3376
R24 VSS.n16 VSS.n15 72.402
R25 VSS.n9 VSS.t10 58.4275
R26 VSS.n19 VSS.n17 56.8118
R27 VSS.n10 VSS.n0 38.0173
R28 VSS VSS.t3 9.03788
R29 VSS.n3 VSS.t17 9.0005
R30 VSS.n5 VSS.t12 9.0005
R31 VSS.n14 VSS.t15 8.96939
R32 VSS.n2 VSS.t9 8.96939
R33 VSS.n4 VSS.t7 8.96939
R34 VSS.n25 VSS.t5 6.77303
R35 VSS.n20 VSS.t1 6.71411
R36 VSS.n22 VSS 5.2005
R37 VSS.n6 VSS 5.2005
R38 VSS.n11 VSS.n10 5.2005
R39 VSS.n10 VSS.n9 5.2005
R40 VSS.n25 VSS.n24 5.2005
R41 VSS.n24 VSS.n23 5.2005
R42 VSS.n21 VSS.n12 5.03032
R43 VSS.n27 VSS.n26 4.5005
R44 VSS VSS.n19 2.6005
R45 VSS.n19 VSS.n18 2.6005
R46 VSS.n17 VSS 2.6005
R47 VSS VSS.n0 2.6005
R48 VSS VSS.n29 2.6005
R49 VSS.n29 VSS.n28 2.6005
R50 VSS.n29 VSS.n27 0.671733
R51 VSS.n3 VSS.n2 0.445721
R52 VSS.n5 VSS 0.42093
R53 VSS VSS.n14 0.400161
R54 VSS VSS.n5 0.221916
R55 VSS.n20 VSS 0.214059
R56 VSS VSS.n21 0.197853
R57 VSS.n12 VSS.n11 0.122874
R58 VSS VSS.n25 0.122874
R59 VSS.n11 VSS 0.109277
R60 VSS.n4 VSS 0.10359
R61 VSS VSS.n3 0.100854
R62 VSS.n21 VSS.n20 0.0897373
R63 VSS VSS.n14 0.0689956
R64 VSS.n2 VSS 0.0689956
R65 VSS VSS.n4 0.0582612
R66 VSS VSS.n12 0.00503237
R67 A A.n0 32.7191
R68 A.n0 A.t0 31.938
R69 A.n0 A.t1 12.2541
R70 SEL.n2 SEL.n1 33.2812
R71 SEL.n1 SEL.t1 31.5469
R72 SEL.n0 SEL.t2 19.0247
R73 SEL.n0 SEL.t0 17.3935
R74 SEL.n1 SEL.t3 12.6451
R75 SEL.n3 SEL.n2 5.99599
R76 SEL.n3 SEL.n0 4.08939
R77 SEL.n2 SEL 0.0705334
R78 SEL SEL.n3 0.0638333
R79 VDD.t23 VDD.n5 826.923
R80 VDD.t16 VDD.n12 596.154
R81 VDD.n13 VDD.t22 448.719
R82 VDD.t8 VDD.n11 443.255
R83 VDD.n12 VDD.t8 432.548
R84 VDD.n11 VDD.t4 421.842
R85 VDD.n13 VDD.t13 414.531
R86 VDD.t22 VDD.t23 341.88
R87 VDD.t13 VDD.t16 341.88
R88 VDD.n12 VDD 315.707
R89 VDD.n18 VDD 315.707
R90 VDD.n18 VDD.t20 116.338
R91 VDD.n12 VDD.t2 116.338
R92 VDD.n19 VDD.n18 100.001
R93 VDD.n19 VDD.n1 71.9005
R94 VDD.n5 VDD.t6 36.3253
R95 VDD.t0 VDD.t11 26.4005
R96 VDD.n18 VDD.t0 11.2005
R97 VDD VDD.t5 6.7809
R98 VDD.n6 VDD.t17 6.61028
R99 VDD.n3 VDD.n2 6.61028
R100 VDD.n9 VDD.n7 6.57115
R101 VDD.n0 VDD.t1 6.57115
R102 VDD.n16 VDD.n15 6.57115
R103 VDD VDD.t12 6.44123
R104 VDD.n4 VDD.t7 6.40636
R105 VDD.n8 VDD.t3 6.40636
R106 VDD.n17 VDD.t21 6.40636
R107 VDD VDD.n13 6.30198
R108 VDD.n5 VDD 6.3005
R109 VDD.n11 VDD.n10 6.3005
R110 VDD VDD.n19 6.3005
R111 VDD VDD.n14 0.919595
R112 VDD.n14 VDD.n4 0.501259
R113 VDD.n6 VDD.n3 0.291409
R114 VDD VDD.n6 0.284603
R115 VDD.n10 VDD.n9 0.219398
R116 VDD.n16 VDD.n1 0.219398
R117 VDD VDD.n0 0.210246
R118 VDD.n0 VDD 0.18379
R119 VDD.n9 VDD.n8 0.145855
R120 VDD.n17 VDD.n16 0.145855
R121 VDD.n14 VDD.n3 0.0595909
R122 VDD.n8 VDD 0.0353691
R123 VDD VDD.n17 0.0353691
R124 VDD VDD.n4 0.0319151
R125 VDD.n14 VDD 0.00713934
R126 VDD.n10 VDD 0.00202542
R127 VDD.n1 VDD 0.00202542
R128 OUT.n2 OUT.n1 9.02722
R129 OUT.n2 OUT.n0 6.48941
R130 OUT OUT.n2 0.130713
C0 a_1557_553# A 5.22e-21
C1 SEL A 0.148f
C2 a_268_215# VDD 0.00253f
C3 a_1557_553# VDD 0.899f
C4 SEL AND_0.B 0.108f
C5 B a_672_1152# 8.64e-19
C6 AND_1.Inverter_0.IN A 0.00979f
C7 SEL VDD 0.547f
C8 VDD OR_0.Inverter_0.IN 0.305f
C9 OR_0.B OR_0.A 0.335f
C10 AND_1.Inverter_0.IN AND_0.B 0.0024f
C11 SEL AND_0.Inverter_0.IN 0.00162f
C12 a_672_1152# OR_0.A 0.00337f
C13 AND_1.Inverter_0.IN VDD 0.582f
C14 OUT VDD 0.125f
C15 B A 0.00236f
C16 B AND_0.B 0.191f
C17 OR_0.A A 1.16e-20
C18 B VDD 0.443f
C19 B AND_0.Inverter_0.IN 0.0126f
C20 OR_0.A AND_0.B 0.00664f
C21 SEL a_268_215# 0.155f
C22 OR_0.A VDD 0.938f
C23 a_1557_553# OR_0.Inverter_0.IN 0.162f
C24 OR_0.A AND_0.Inverter_0.IN 0.162f
C25 AND_1.Inverter_0.IN a_268_215# 0.0608f
C26 AND_1.Inverter_0.IN a_1557_553# 7.88e-20
C27 SEL OR_0.Inverter_0.IN 2.23e-22
C28 AND_1.Inverter_0.IN SEL 0.128f
C29 AND_1.Inverter_0.IN OR_0.Inverter_0.IN 1.3e-19
C30 OUT OR_0.Inverter_0.IN 0.116f
C31 OR_0.B A 1.57e-20
C32 a_268_215# B 2.56e-19
C33 a_672_1152# AND_0.B 0.155f
C34 SEL B 0.0965f
C35 OR_0.B VDD 0.418f
C36 a_1557_553# OR_0.A 0.2f
C37 OR_0.B AND_0.Inverter_0.IN 7.69e-20
C38 a_672_1152# VDD 0.00253f
C39 AND_1.Inverter_0.IN B 6.91e-19
C40 a_672_1152# AND_0.Inverter_0.IN 0.0608f
C41 SEL OR_0.A 0.015f
C42 OR_0.A OR_0.Inverter_0.IN 0.261f
C43 AND_1.Inverter_0.IN OR_0.A 0.00447f
C44 A AND_0.B 1.12e-19
C45 OUT OR_0.A 3.24e-19
C46 A VDD 0.251f
C47 VDD AND_0.B 0.374f
C48 AND_0.Inverter_0.IN AND_0.B 0.129f
C49 OR_0.B a_268_215# 4.07e-20
C50 B OR_0.A 0.00142f
C51 OR_0.B a_1557_553# 0.0243f
C52 AND_0.Inverter_0.IN VDD 0.582f
C53 OR_0.B SEL 0.00118f
C54 OR_0.B OR_0.Inverter_0.IN 0.0441f
C55 SEL a_672_1152# 0.00164f
C56 OR_0.B AND_1.Inverter_0.IN 0.12f
C57 AND_1.Inverter_0.IN a_672_1152# 5.44e-20
C58 a_268_215# A 8.64e-19
C59 a_268_215# VSS 0.214f
C60 OUT VSS 0.188f
C61 OR_0.Inverter_0.IN VSS 0.762f
C62 a_1557_553# VSS 0.132f
C63 AND_1.Inverter_0.IN VSS 0.448f
C64 OR_0.B VSS 0.611f
C65 A VSS 0.359f
C66 a_672_1152# VSS 0.188f
C67 OR_0.A VSS 0.769f
C68 AND_0.Inverter_0.IN VSS 0.408f
C69 AND_0.B VSS 0.536f
C70 B VSS 0.418f
C71 SEL VSS 1.14f
C72 VDD VSS 9.46f
.ends

