magic
tech gf180mcuC
magscale 1 10
timestamp 1693459011
<< nwell >>
rect -264 -386 264 386
<< nsubdiff >>
rect -240 290 240 362
rect -240 -290 -168 290
rect 168 -290 240 290
rect -240 -362 240 -290
<< polysilicon >>
rect -80 189 80 202
rect -80 143 -67 189
rect 67 143 80 189
rect -80 100 80 143
rect -80 -143 80 -100
rect -80 -189 -67 -143
rect 67 -189 80 -143
rect -80 -202 80 -189
<< polycontact >>
rect -67 143 67 189
rect -67 -189 67 -143
<< ppolyres >>
rect -80 -100 80 100
<< metal1 >>
rect -78 143 -67 189
rect 67 143 78 189
rect -78 -189 -67 -143
rect 67 -189 78 -143
<< properties >>
string FIXED_BBOX -204 -326 204 326
string gencell ppolyf_u
string library gf180mcu
string parameters w 0.80 l 1.00 m 1 nx 1 wmin 0.80 lmin 1.00 rho 315 val 431.506 dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0
<< end >>
