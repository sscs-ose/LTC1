* NGSPICE file created from Local_Enc_flat.ext - technology: gf180mcuC

.subckt Local_Enc_flat VDD VSS Q QB Ci Ri Ri-1
X0 a_305_1140# Ci.t0 VSS.t21 VSS.t20 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X1 NAND_6.A Ri.t0 VDD.t16 VDD.t15 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X2 VDD NAND_6.A NAND_5.A VDD.t26 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X3 NAND_1.B Ri-1.t0 VDD.t11 VDD.t10 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X4 Q NAND_8.A a_1879_1140# VSS.t25 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X5 a_305_2111# Ri-1.t1 VSS.t6 VSS.t5 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X6 a_1879_1140# QB.t3 VSS.t9 VSS.t8 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X7 a_1068_164# NAND_6.B VSS.t16 VSS.t15 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X8 VDD Q.t3 QB.t2 VDD.t29 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X9 a_305_165# Ri.t1 VSS.t11 VSS.t10 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X10 VDD NAND_5.A NAND_8.A VDD.t19 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X11 NAND_5.A NAND_6.A a_1068_164# VSS.t17 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X12 QB NAND_4.B VDD.t6 VDD.t5 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X13 QB Q.t4 a_1879_2111# VSS.t18 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X14 VDD Ci.t1 NAND_6.B VDD.t34 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X15 a_1879_2111# NAND_4.B VSS.t4 VSS.t3 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X16 NAND_8.A NAND_5.B VDD.t18 VDD.t17 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X17 VDD Ri.t2 NAND_6.A VDD.t12 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X18 NAND_4.B NAND_8.A VDD.t44 VDD.t43 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X19 VDD NAND_8.A NAND_4.B VDD.t40 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X20 NAND_8.A NAND_5.A a_1068_1140# VSS.t14 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X21 NAND_6.B Ci.t2 VDD.t33 VDD.t32 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X22 NAND_6.B Ci.t3 a_305_1140# VSS.t19 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X23 a_1068_1140# NAND_5.B VSS.t13 VSS.t12 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X24 NAND_6.A Ri.t3 a_305_165# VSS.t26 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X25 a_1879_164# NAND_8.A VSS.t24 VSS.t23 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X26 VDD NAND_1.B NAND_5.B VDD.t2 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X27 VDD Ri-1.t2 NAND_1.B VDD.t7 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X28 NAND_5.B NAND_1.B VDD.t1 VDD.t0 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X29 VDD NAND_8.A Q.t2 VDD.t37 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X30 NAND_5.B NAND_1.B a_1068_2111# VSS.t2 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X31 NAND_4.B NAND_8.A a_1879_164# VSS.t22 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X32 NAND_1.B Ri-1.t3 a_305_2111# VSS.t7 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X33 a_1068_2111# NAND_1.B VSS.t1 VSS.t0 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X34 Q QB.t4 VDD.t23 VDD.t22 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X35 NAND_5.A NAND_6.B VDD.t25 VDD.t24 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
R0 Ci.n0 Ci.t1 28.2228
R1 Ci.n1 Ci.t0 26.9784
R2 Ci.n1 Ci.t2 14.7248
R3 Ci.n0 Ci.t3 14.4701
R4 Ci Ci.n0 4.53357
R5 Ci Ci.n1 4.18544
R6 VSS.t18 VSS.n4 9953.06
R7 VSS.n8 VSS.n7 6710.53
R8 VSS.t20 VSS.n16 2739.78
R9 VSS.t23 VSS.n20 2616.05
R10 VSS.n20 VSS.t17 2608.02
R11 VSS.n27 VSS.t15 2421.48
R12 VSS.t26 VSS.n27 2409.48
R13 VSS.n7 VSS.t3 2298.26
R14 VSS.t8 VSS.n8 2273.61
R15 VSS.n4 VSS.t25 2148.07
R16 VSS.n2 VSS.t0 2129.07
R17 VSS.t7 VSS.n2 2122.02
R18 VSS.n15 VSS.t12 2106.22
R19 VSS.t19 VSS.n15 2102.28
R20 VSS.n21 VSS.t22 682.1
R21 VSS.n26 VSS.t17 682.1
R22 VSS.n28 VSS.t26 680.419
R23 VSS.n21 VSS.t23 601.852
R24 VSS.t15 VSS.n26 601.852
R25 VSS.n28 VSS.t10 600.37
R26 VSS.n6 VSS.t18 599.241
R27 VSS.n1 VSS.t2 599.241
R28 VSS.n3 VSS.t7 599.241
R29 VSS.n17 VSS.t19 594.087
R30 VSS.n14 VSS.t14 592.812
R31 VSS.t3 VSS.n6 528.742
R32 VSS.t0 VSS.n1 528.742
R33 VSS.n3 VSS.t5 528.742
R34 VSS.n17 VSS.t20 524.194
R35 VSS.n9 VSS.t8 523.069
R36 VSS.t12 VSS.n14 523.069
R37 VSS.n11 VSS.t9 6.65541
R38 VSS.n12 VSS.t13 6.65541
R39 VSS.n19 VSS.t21 6.65541
R40 VSS.n32 VSS.t6 6.65541
R41 VSS.n30 VSS.t11 6.65541
R42 VSS.n24 VSS.t16 6.65541
R43 VSS.n23 VSS.t24 6.65541
R44 VSS.n0 VSS.t4 6.65541
R45 VSS.n34 VSS.t1 6.65541
R46 VSS.n22 VSS.n21 5.2005
R47 VSS.n26 VSS.n25 5.2005
R48 VSS.n29 VSS.n28 5.2005
R49 VSS.n10 VSS.n9 5.2005
R50 VSS.n14 VSS.n13 5.2005
R51 VSS.n18 VSS.n17 5.2005
R52 VSS.n33 VSS.n3 5.2005
R53 VSS.n6 VSS.n5 5.2005
R54 VSS.n35 VSS.n1 5.2005
R55 VSS.n32 VSS.n31 3.81335
R56 VSS.n31 VSS.n30 3.80502
R57 VSS.n31 VSS.n19 2.53474
R58 VSS VSS.n11 0.684889
R59 VSS VSS.n23 0.684889
R60 VSS VSS.n0 0.684889
R61 VSS.n12 VSS 0.620412
R62 VSS.n34 VSS 0.620412
R63 VSS.n24 VSS 0.620412
R64 VSS.n11 VSS.n10 0.142847
R65 VSS.n13 VSS.n12 0.142847
R66 VSS.n19 VSS.n18 0.142847
R67 VSS.n33 VSS.n32 0.142847
R68 VSS.n30 VSS.n29 0.142847
R69 VSS.n25 VSS.n24 0.142847
R70 VSS.n23 VSS.n22 0.142847
R71 VSS.n5 VSS.n0 0.142847
R72 VSS VSS.n34 0.130908
R73 VSS.n35 VSS 0.0124388
R74 VSS.n10 VSS 0.00141837
R75 VSS.n13 VSS 0.00141837
R76 VSS.n18 VSS 0.00141837
R77 VSS VSS.n33 0.00141837
R78 VSS.n29 VSS 0.00141837
R79 VSS.n25 VSS 0.00141837
R80 VSS.n22 VSS 0.00141837
R81 VSS.n5 VSS 0.00141837
R82 VSS VSS.n35 0.00141837
R83 Ri.n0 Ri.t2 28.2228
R84 Ri.n1 Ri.t1 26.9784
R85 Ri.n1 Ri.t0 14.7248
R86 Ri.n0 Ri.t3 14.4701
R87 Ri Ri.n0 4.53357
R88 Ri Ri.n1 4.18544
R89 VDD.n6 VDD.t2 178.431
R90 VDD.n9 VDD.t7 178.431
R91 VDD.n21 VDD.t34 178.431
R92 VDD.n17 VDD.t19 178.431
R93 VDD.n13 VDD.t37 178.431
R94 VDD.n35 VDD.t12 178.431
R95 VDD.n31 VDD.t26 178.431
R96 VDD.n27 VDD.t40 178.431
R97 VDD.n2 VDD.t29 178.431
R98 VDD.n6 VDD.t0 135.294
R99 VDD.n9 VDD.t10 135.294
R100 VDD.n21 VDD.t32 135.294
R101 VDD.n17 VDD.t17 135.294
R102 VDD.n13 VDD.t22 135.294
R103 VDD.n35 VDD.t15 135.294
R104 VDD.n31 VDD.t24 135.294
R105 VDD.n27 VDD.t43 135.294
R106 VDD.n2 VDD.t5 135.294
R107 VDD.n14 VDD.n12 6.69527
R108 VDD.n28 VDD.n26 6.69527
R109 VDD.n3 VDD.n1 6.69527
R110 VDD.n16 VDD.n11 6.59267
R111 VDD.n20 VDD.n10 6.59267
R112 VDD.n30 VDD.n25 6.59267
R113 VDD.n34 VDD.n24 6.59267
R114 VDD.n41 VDD.n8 6.59267
R115 VDD.n5 VDD.n0 6.59267
R116 VDD.n15 VDD.t23 6.55815
R117 VDD.n19 VDD.t18 6.55815
R118 VDD.n23 VDD.t33 6.55815
R119 VDD.n29 VDD.t44 6.55815
R120 VDD.n33 VDD.t25 6.55815
R121 VDD.n37 VDD.t16 6.55815
R122 VDD.n39 VDD.t11 6.55815
R123 VDD.n4 VDD.t6 6.55815
R124 VDD.n42 VDD.t1 6.55815
R125 VDD.n14 VDD.n13 6.3005
R126 VDD.n18 VDD.n17 6.3005
R127 VDD.n22 VDD.n21 6.3005
R128 VDD.n28 VDD.n27 6.3005
R129 VDD.n32 VDD.n31 6.3005
R130 VDD.n36 VDD.n35 6.3005
R131 VDD.n40 VDD.n9 6.3005
R132 VDD.n3 VDD.n2 6.3005
R133 VDD.n7 VDD.n6 6.3005
R134 VDD.n39 VDD.n38 3.9851
R135 VDD.n38 VDD.n37 3.87957
R136 VDD.n38 VDD.n23 2.58214
R137 VDD.n16 VDD.n15 0.339604
R138 VDD.n30 VDD.n29 0.339604
R139 VDD.n5 VDD.n4 0.339604
R140 VDD.n20 VDD.n19 0.302039
R141 VDD.n34 VDD.n33 0.302039
R142 VDD.n42 VDD.n41 0.302039
R143 VDD.n18 VDD.n16 0.1031
R144 VDD.n22 VDD.n20 0.1031
R145 VDD.n32 VDD.n30 0.1031
R146 VDD.n36 VDD.n34 0.1031
R147 VDD.n41 VDD.n40 0.1031
R148 VDD.n7 VDD.n5 0.1031
R149 VDD.n15 VDD 0.0893
R150 VDD.n19 VDD 0.0893
R151 VDD.n23 VDD 0.0893
R152 VDD.n29 VDD 0.0893
R153 VDD.n33 VDD 0.0893
R154 VDD.n37 VDD 0.0893
R155 VDD VDD.n39 0.0893
R156 VDD.n4 VDD 0.0893
R157 VDD VDD.n42 0.0839
R158 VDD VDD.n14 0.0017
R159 VDD VDD.n18 0.0017
R160 VDD VDD.n22 0.0017
R161 VDD VDD.n28 0.0017
R162 VDD VDD.n32 0.0017
R163 VDD VDD.n36 0.0017
R164 VDD.n40 VDD 0.0017
R165 VDD VDD.n3 0.0017
R166 VDD VDD.n7 0.0017
R167 Ri-1.n0 Ri-1.t2 28.2228
R168 Ri-1.n1 Ri-1.t1 26.9784
R169 Ri-1.n1 Ri-1.t0 14.7248
R170 Ri-1.n0 Ri-1.t3 14.4701
R171 Ri-1 Ri-1.n0 4.53357
R172 Ri-1 Ri-1.n1 4.18544
R173 Q.n1 Q.t3 28.2228
R174 Q.n1 Q.t4 14.4701
R175 Q.n5 Q.n0 6.8765
R176 Q.n4 Q 6.04981
R177 Q Q.n1 4.53357
R178 Q.n3 Q.t2 3.6405
R179 Q.n3 Q.n2 3.6405
R180 Q.n4 Q.n3 2.6005
R181 Q.n5 Q.n4 0.484465
R182 Q Q.n5 0.17463
R183 QB.n0 QB.t3 26.9784
R184 QB.n0 QB.t4 14.7248
R185 QB.n1 QB 10.3144
R186 QB.n5 QB.n2 6.8765
R187 QB QB.n0 4.18544
R188 QB.n4 QB.t2 3.6405
R189 QB.n4 QB.n3 3.6405
R190 QB.n5 QB.n4 3.08447
R191 QB QB.n1 0.241152
R192 QB QB.n5 0.17463
R193 QB.n1 QB 0.112881
C0 VDD Q 0.585f
C1 NAND_1.B a_1068_2111# 0.0852f
C2 NAND_5.A Q 2.28e-19
C3 Ri a_1879_164# 3.42e-22
C4 Ri VDD 0.36f
C5 Ri NAND_5.A 9e-19
C6 Q a_1068_2111# 6.06e-19
C7 Ri a_1068_164# 1.61e-21
C8 VDD NAND_5.B 0.864f
C9 NAND_5.A NAND_5.B 0.316f
C10 NAND_5.B a_1068_2111# 0.0469f
C11 VDD Ri-1 0.382f
C12 VDD NAND_6.B 0.618f
C13 VDD a_305_2111# 8.42e-19
C14 NAND_6.B NAND_5.A 0.232f
C15 QB Ci 5.92e-19
C16 NAND_6.B a_1068_164# 0.00403f
C17 QB a_1879_2111# 0.0423f
C18 NAND_4.B NAND_6.A 1.31e-19
C19 NAND_8.A NAND_6.A 0.0124f
C20 NAND_1.B QB 1.31e-19
C21 a_1068_1140# NAND_5.B 0.0043f
C22 a_305_1140# NAND_5.A 2.15e-19
C23 QB Q 0.302f
C24 a_1068_1140# NAND_6.B 2.79e-20
C25 a_1879_1140# QB 0.00549f
C26 NAND_5.B QB 0.00682f
C27 a_1879_2111# Q 0.0961f
C28 Ri Ci 0.00475f
C29 VDD NAND_6.A 0.358f
C30 NAND_8.A NAND_4.B 0.345f
C31 NAND_5.A NAND_6.A 0.216f
C32 NAND_6.A a_1068_164# 0.0812f
C33 NAND_5.B Ci 0.0105f
C34 NAND_1.B Q 0.004f
C35 NAND_6.B QB 4.6e-19
C36 NAND_5.B a_1879_2111# 6.99e-20
C37 Ri-1 Ci 0.00479f
C38 NAND_6.B Ci 0.235f
C39 NAND_1.B NAND_5.B 0.344f
C40 Ci a_305_2111# 5.76e-20
C41 NAND_4.B a_1879_164# 0.0419f
C42 a_1879_1140# Q 0.043f
C43 NAND_5.B Q 0.0478f
C44 NAND_8.A a_1879_164# 0.0852f
C45 NAND_1.B Ri-1 0.24f
C46 VDD NAND_4.B 0.673f
C47 a_1068_1140# NAND_6.A 5.69e-20
C48 NAND_1.B NAND_6.B 1.35e-19
C49 NAND_1.B a_305_2111# 0.0419f
C50 NAND_5.A NAND_4.B 0.00496f
C51 NAND_8.A VDD 0.864f
C52 NAND_8.A NAND_5.A 0.333f
C53 a_305_1140# Ci 0.0852f
C54 Ri a_305_165# 0.0852f
C55 Ri NAND_6.B 0.0132f
C56 Ri-1 NAND_5.B 0.00958f
C57 NAND_6.B NAND_5.B 0.0342f
C58 NAND_5.B a_305_2111# 0.00175f
C59 NAND_5.A a_1879_164# 1.88e-20
C60 NAND_6.A Ci 1.17e-19
C61 a_1068_1140# NAND_8.A 0.045f
C62 VDD NAND_5.A 0.503f
C63 NAND_6.B Ri-1 1.18e-19
C64 Ri-1 a_305_2111# 0.0852f
C65 NAND_5.A a_1068_164# 0.0451f
C66 a_305_1140# Ri 5.71e-20
C67 NAND_5.A a_1068_2111# 5.76e-20
C68 NAND_4.B QB 0.453f
C69 NAND_8.A QB 0.427f
C70 a_305_1140# NAND_6.B 0.0444f
C71 Ri NAND_6.A 0.233f
C72 NAND_8.A Ci 8.19e-19
C73 a_1068_1140# NAND_5.A 0.0874f
C74 NAND_4.B a_1879_2111# 0.00495f
C75 NAND_8.A a_1879_2111# 5.76e-20
C76 NAND_6.A a_305_165# 0.0419f
C77 NAND_1.B NAND_4.B 0.00819f
C78 NAND_8.A NAND_1.B 1.18e-19
C79 a_1879_164# QB 3.34e-19
C80 NAND_6.B NAND_6.A 0.429f
C81 VDD QB 0.625f
C82 NAND_4.B Q 0.601f
C83 NAND_5.A QB 0.00927f
C84 NAND_8.A Q 0.201f
C85 Ri NAND_4.B 2.34e-22
C86 VDD Ci 0.372f
C87 Ri NAND_8.A 5.07e-19
C88 NAND_5.A Ci 0.00321f
C89 a_1879_1140# NAND_4.B 0.00331f
C90 NAND_4.B NAND_5.B 0.026f
C91 a_1879_1140# NAND_8.A 0.0821f
C92 NAND_8.A NAND_5.B 0.0646f
C93 NAND_1.B VDD 0.628f
C94 NAND_1.B NAND_5.A 0.00251f
C95 NAND_4.B Ri-1 1.08e-19
C96 NAND_6.B NAND_4.B 2.09e-20
C97 a_1879_164# Q 1.23e-19
C98 NAND_8.A NAND_6.B 0.00405f
C99 a_1879_164# VSS 0.0983f
C100 a_1068_164# VSS 0.0986f
C101 a_305_165# VSS 0.0998f
C102 NAND_6.A VSS 0.56f
C103 Ri VSS 0.622f
C104 a_1879_1140# VSS 0.0983f
C105 a_1068_1140# VSS 0.0983f
C106 a_305_1140# VSS 0.0997f
C107 NAND_6.B VSS 0.682f
C108 NAND_8.A VSS 1.43f
C109 NAND_5.A VSS 0.707f
C110 Ci VSS 0.609f
C111 a_1879_2111# VSS 0.0983f
C112 a_1068_2111# VSS 0.0983f
C113 a_305_2111# VSS 0.0983f
C114 QB VSS 0.903f
C115 NAND_5.B VSS 0.697f
C116 Q VSS 0.76f
C117 NAND_4.B VSS 0.764f
C118 NAND_1.B VSS 0.754f
C119 Ri-1 VSS 0.591f
C120 VDD VSS 13.9f
.ends

