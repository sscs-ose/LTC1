magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1451 -1046 1451 1046
<< metal1 >>
rect -451 40 451 46
rect -451 14 -445 40
rect -419 14 -391 40
rect -365 14 -337 40
rect -311 14 -283 40
rect -257 14 -229 40
rect -203 14 -175 40
rect -149 14 -121 40
rect -95 14 -67 40
rect -41 14 -13 40
rect 13 14 41 40
rect 67 14 95 40
rect 121 14 149 40
rect 175 14 203 40
rect 229 14 257 40
rect 283 14 311 40
rect 337 14 365 40
rect 391 14 419 40
rect 445 14 451 40
rect -451 -14 451 14
rect -451 -40 -445 -14
rect -419 -40 -391 -14
rect -365 -40 -337 -14
rect -311 -40 -283 -14
rect -257 -40 -229 -14
rect -203 -40 -175 -14
rect -149 -40 -121 -14
rect -95 -40 -67 -14
rect -41 -40 -13 -14
rect 13 -40 41 -14
rect 67 -40 95 -14
rect 121 -40 149 -14
rect 175 -40 203 -14
rect 229 -40 257 -14
rect 283 -40 311 -14
rect 337 -40 365 -14
rect 391 -40 419 -14
rect 445 -40 451 -14
rect -451 -46 451 -40
<< via1 >>
rect -445 14 -419 40
rect -391 14 -365 40
rect -337 14 -311 40
rect -283 14 -257 40
rect -229 14 -203 40
rect -175 14 -149 40
rect -121 14 -95 40
rect -67 14 -41 40
rect -13 14 13 40
rect 41 14 67 40
rect 95 14 121 40
rect 149 14 175 40
rect 203 14 229 40
rect 257 14 283 40
rect 311 14 337 40
rect 365 14 391 40
rect 419 14 445 40
rect -445 -40 -419 -14
rect -391 -40 -365 -14
rect -337 -40 -311 -14
rect -283 -40 -257 -14
rect -229 -40 -203 -14
rect -175 -40 -149 -14
rect -121 -40 -95 -14
rect -67 -40 -41 -14
rect -13 -40 13 -14
rect 41 -40 67 -14
rect 95 -40 121 -14
rect 149 -40 175 -14
rect 203 -40 229 -14
rect 257 -40 283 -14
rect 311 -40 337 -14
rect 365 -40 391 -14
rect 419 -40 445 -14
<< metal2 >>
rect -451 40 451 46
rect -451 14 -445 40
rect -419 14 -391 40
rect -365 14 -337 40
rect -311 14 -283 40
rect -257 14 -229 40
rect -203 14 -175 40
rect -149 14 -121 40
rect -95 14 -67 40
rect -41 14 -13 40
rect 13 14 41 40
rect 67 14 95 40
rect 121 14 149 40
rect 175 14 203 40
rect 229 14 257 40
rect 283 14 311 40
rect 337 14 365 40
rect 391 14 419 40
rect 445 14 451 40
rect -451 -14 451 14
rect -451 -40 -445 -14
rect -419 -40 -391 -14
rect -365 -40 -337 -14
rect -311 -40 -283 -14
rect -257 -40 -229 -14
rect -203 -40 -175 -14
rect -149 -40 -121 -14
rect -95 -40 -67 -14
rect -41 -40 -13 -14
rect 13 -40 41 -14
rect 67 -40 95 -14
rect 121 -40 149 -14
rect 175 -40 203 -14
rect 229 -40 257 -14
rect 283 -40 311 -14
rect 337 -40 365 -14
rect 391 -40 419 -14
rect 445 -40 451 -14
rect -451 -46 451 -40
<< end >>
