* NGSPICE file created from CLK_div_2_mag_flat.ext - technology: gf180mcuC

.subckt CLK_div_2_mag_flat VDD Vdiv2 CLK RST VSS
X0 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_1.OUT a_1288_1433# VSS.t11 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1 a_1852_1433# JK_FF_mag_0.nand3_mag_1.IN1 VSS.t21 VSS.t20 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2 VDD RST.t0 JK_FF_mag_0.nand3_mag_1.OUT VDD.t31 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X3 a_1288_1433# JK_FF_mag_0.nand3_mag_0.OUT VSS.t1 VSS.t0 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X4 Vdiv2 JK_FF_mag_0.QB a_2416_1433# VSS.t7 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X5 VDD JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_4.IN2 VDD.t7 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X6 Vdiv2 JK_FF_mag_0.nand2_mag_1.IN2 VDD.t47 VDD.t46 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X7 a_718_292# CLK.t0 a_558_292# VSS.t26 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X8 a_2006_336# JK_FF_mag_0.nand3_mag_1.OUT VSS.t10 VSS.t9 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X9 a_1282_292# JK_FF_mag_0.nand3_mag_2.OUT VSS.t3 VSS.t2 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X10 JK_FF_mag_0.nand2_mag_3.IN1 CLK.t1 VSS.t23 VSS.t22 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X11 JK_FF_mag_0.nand3_mag_2.OUT Vdiv2.t3 VDD.t49 VDD.t48 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X12 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand2_mag_3.IN1 a_2006_336# VSS.t5 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X13 a_2416_1433# JK_FF_mag_0.nand2_mag_1.IN2 VSS.t25 VSS.t24 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X14 a_1442_292# RST.t1 a_1282_292# VSS.t12 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X15 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 VDD.t42 VDD.t41 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X16 VDD JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_1.IN2 VDD.t4 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X17 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.QB VDD.t14 VDD.t13 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X18 JK_FF_mag_0.nand3_mag_2.OUT Vdiv2.t4 a_718_292# VSS.t14 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X19 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.QB a_724_1389# VSS.t6 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X20 JK_FF_mag_0.QB JK_FF_mag_0.nand2_mag_4.IN2 VDD.t38 VDD.t37 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X21 JK_FF_mag_0.nand3_mag_2.OUT VDD.t26 VDD.t28 VDD.t27 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X22 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand2_mag_3.IN1 a_1852_1433# VSS.t4 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X23 VDD JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 VDD.t20 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X24 VDD Vdiv2.t5 JK_FF_mag_0.QB VDD.t43 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X25 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 a_1442_292# VSS.t19 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X26 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand3_mag_1.IN1 VDD.t40 VDD.t39 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X27 VDD JK_FF_mag_0.QB Vdiv2.t1 VDD.t10 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X28 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_0.OUT VDD.t1 VDD.t0 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X29 VDD CLK.t2 JK_FF_mag_0.nand3_mag_2.OUT VDD.t15 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X30 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_2.OUT VDD.t3 VDD.t2 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X31 a_2570_336# JK_FF_mag_0.nand2_mag_4.IN2 VSS.t18 VSS.t17 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X32 VDD CLK.t3 JK_FF_mag_0.nand3_mag_0.OUT VDD.t34 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X33 JK_FF_mag_0.nand2_mag_3.IN1 CLK.t4 VDD.t30 VDD.t29 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X34 JK_FF_mag_0.nand3_mag_0.OUT VDD.t23 VDD.t25 VDD.t24 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X35 a_724_1389# CLK.t5 a_564_1389# VSS.t13 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X36 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand3_mag_1.OUT VDD.t19 VDD.t18 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X37 a_564_1389# VDD.t50 VSS.t28 VSS.t27 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X38 a_558_292# VDD.t51 VSS.t16 VSS.t15 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X39 JK_FF_mag_0.QB Vdiv2.t6 a_2570_336# VSS.t8 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
R0 VSS.t8 VSS.n13 9652.01
R1 VSS.n24 VSS.t15 5796.73
R2 VSS.t24 VSS.t4 2307.56
R3 VSS.t11 VSS.t20 2307.56
R4 VSS.t0 VSS.t6 2307.56
R5 VSS.t22 VSS.t27 2307.56
R6 VSS.n13 VSS.t7 2244.73
R7 VSS.t5 VSS.t17 2221.66
R8 VSS.t14 VSS.t2 2221.66
R9 VSS.t6 VSS.t13 913.885
R10 VSS.t12 VSS.t19 879.865
R11 VSS.t26 VSS.t14 879.865
R12 VSS.n7 VSS.t4 548.331
R13 VSS.n8 VSS.t11 548.331
R14 VSS.n12 VSS.t13 548.331
R15 VSS.n16 VSS.t8 527.919
R16 VSS.n17 VSS.t5 527.919
R17 VSS.n22 VSS.t12 527.919
R18 VSS.n23 VSS.t26 527.919
R19 VSS.n25 VSS.n24 376.978
R20 VSS.n2 VSS.t24 365.555
R21 VSS.t20 VSS.n7 365.555
R22 VSS.n8 VSS.t0 365.555
R23 VSS.t27 VSS.n12 365.555
R24 VSS.t17 VSS.n16 351.947
R25 VSS.n17 VSS.t9 351.947
R26 VSS.t2 VSS.n22 351.947
R27 VSS.t15 VSS.n23 351.947
R28 VSS.n25 VSS.t22 34.2711
R29 VSS.n26 VSS.t23 9.3736
R30 VSS.n14 VSS.t18 7.19156
R31 VSS.n19 VSS.t10 7.19156
R32 VSS.n4 VSS.t25 7.19156
R33 VSS.n5 VSS.t21 7.19156
R34 VSS.n10 VSS.t1 7.19156
R35 VSS.n20 VSS.t3 5.91399
R36 VSS.n28 VSS.t16 5.91399
R37 VSS.n1 VSS.t28 5.91399
R38 VSS.n26 VSS.n25 5.2005
R39 VSS.n12 VSS.n11 5.2005
R40 VSS.n9 VSS.n8 5.2005
R41 VSS.n7 VSS.n6 5.2005
R42 VSS.n3 VSS.n2 5.2005
R43 VSS.n23 VSS.n0 5.2005
R44 VSS.n22 VSS.n21 5.2005
R45 VSS.n18 VSS.n17 5.2005
R46 VSS.n16 VSS.n15 5.2005
R47 VSS.n28 VSS.n27 0.961338
R48 VSS VSS.n4 0.343161
R49 VSS.n5 VSS 0.343161
R50 VSS.n21 VSS.n19 0.295924
R51 VSS.n11 VSS 0.289491
R52 VSS.n14 VSS 0.211517
R53 VSS VSS.n10 0.191234
R54 VSS VSS.n0 0.168805
R55 VSS.n27 VSS 0.137685
R56 VSS.n20 VSS 0.127619
R57 VSS.n4 VSS.n3 0.118573
R58 VSS.n6 VSS.n5 0.118573
R59 VSS.n10 VSS.n9 0.118573
R60 VSS VSS.n1 0.115271
R61 VSS.n27 VSS.n1 0.10206
R62 VSS.n15 VSS.n14 0.0732119
R63 VSS.n19 VSS.n18 0.0732119
R64 VSS VSS.n20 0.071178
R65 VSS VSS.n28 0.071178
R66 VSS.n3 VSS 0.00545413
R67 VSS.n6 VSS 0.00545413
R68 VSS.n9 VSS 0.00545413
R69 VSS.n11 VSS 0.00380275
R70 VSS.n15 VSS 0.00355085
R71 VSS.n18 VSS 0.00355085
R72 VSS.n21 VSS 0.0025339
R73 VSS VSS.n0 0.0025339
R74 VSS VSS.n26 0.00219811
R75 RST.n0 RST.t1 36.935
R76 RST.n0 RST.t0 18.1962
R77 RST.n1 RST.n0 2.12207
R78 RST.n3 RST 1.63657
R79 RST.n6 RST.n5 1.5005
R80 RST.n4 RST.n3 1.12901
R81 RST RST.n7 0.0379319
R82 RST.n7 RST.n6 0.0361897
R83 RST.n5 RST.n2 0.0145153
R84 RST.n6 RST.n1 0.0067069
R85 RST.n5 RST.n4 0.00523684
R86 VDD.t4 VDD.t46 765.152
R87 VDD.t39 VDD.t20 765.152
R88 VDD.t13 VDD.t0 765.152
R89 VDD.t7 VDD.t37 765.152
R90 VDD.t41 VDD.t18 765.152
R91 VDD.t48 VDD.t2 765.152
R92 VDD VDD.n47 429.187
R93 VDD.t34 VDD.t13 303.031
R94 VDD.t31 VDD.t41 303.031
R95 VDD.t15 VDD.t48 303.031
R96 VDD.n33 VDD.t10 193.183
R97 VDD.n34 VDD.t4 193.183
R98 VDD.n43 VDD.t20 193.183
R99 VDD.n44 VDD.t34 193.183
R100 VDD.n5 VDD.t43 193.183
R101 VDD.n7 VDD.t7 193.183
R102 VDD.n10 VDD.t31 193.183
R103 VDD.n13 VDD.t15 193.183
R104 VDD.t46 VDD.n33 109.849
R105 VDD.n34 VDD.t39 109.849
R106 VDD.t0 VDD.n43 109.849
R107 VDD.n44 VDD.t24 109.849
R108 VDD.t37 VDD.n5 109.849
R109 VDD.t18 VDD.n7 109.849
R110 VDD.t2 VDD.n10 109.849
R111 VDD.n13 VDD.t27 109.849
R112 VDD.n47 VDD.t29 59.702
R113 VDD.n14 VDD.t23 30.9379
R114 VDD.n16 VDD.t26 30.9379
R115 VDD.n14 VDD.t50 24.5101
R116 VDD.n16 VDD.t51 24.5101
R117 VDD.n19 VDD.n13 6.3005
R118 VDD.n22 VDD.n10 6.3005
R119 VDD.n25 VDD.n7 6.3005
R120 VDD.n28 VDD.n5 6.3005
R121 VDD.n33 VDD.n32 6.3005
R122 VDD.n35 VDD.n34 6.3005
R123 VDD.n43 VDD.n42 6.3005
R124 VDD.n45 VDD.n44 6.3005
R125 VDD VDD.t30 5.13604
R126 VDD.n18 VDD.t28 5.13287
R127 VDD.n21 VDD.t3 5.13287
R128 VDD.n24 VDD.t19 5.13287
R129 VDD.n26 VDD.n6 5.13287
R130 VDD.n27 VDD.t38 5.13287
R131 VDD.n29 VDD.n4 5.13287
R132 VDD.n46 VDD.t25 5.11708
R133 VDD.n41 VDD.t1 5.11708
R134 VDD.n37 VDD.n0 5.11708
R135 VDD.n36 VDD.t40 5.11708
R136 VDD.n2 VDD.n1 5.11708
R137 VDD.n31 VDD.t47 5.11708
R138 VDD.n30 VDD.n3 5.11708
R139 VDD VDD.n16 4.08487
R140 VDD.n15 VDD.n14 4.07684
R141 VDD.n17 VDD.n15 3.00126
R142 VDD.n17 VDD 2.87711
R143 VDD.n20 VDD.n12 2.85787
R144 VDD.n23 VDD.n9 2.85787
R145 VDD.n40 VDD.n39 2.84208
R146 VDD.n18 VDD.n17 2.28069
R147 VDD.n39 VDD.t14 2.2755
R148 VDD.n39 VDD.n38 2.2755
R149 VDD.n12 VDD.t49 2.2755
R150 VDD.n12 VDD.n11 2.2755
R151 VDD.n9 VDD.t42 2.2755
R152 VDD.n9 VDD.n8 2.2755
R153 VDD.n30 VDD.n29 1.1341
R154 VDD.n24 VDD.n23 0.233919
R155 VDD.n21 VDD.n20 0.233919
R156 VDD VDD.n46 0.165331
R157 VDD.n27 VDD.n26 0.141016
R158 VDD.n31 VDD.n2 0.12286
R159 VDD.n37 VDD.n36 0.12286
R160 VDD.n29 VDD.n28 0.107339
R161 VDD.n26 VDD.n25 0.107339
R162 VDD.n23 VDD 0.106177
R163 VDD.n20 VDD 0.106177
R164 VDD VDD.n40 0.0975787
R165 VDD.n32 VDD.n30 0.0935337
R166 VDD.n35 VDD.n2 0.0935337
R167 VDD.n42 VDD.n37 0.0935337
R168 VDD.n40 VDD 0.0925225
R169 VDD.n22 VDD.n21 0.080629
R170 VDD.n19 VDD.n18 0.080629
R171 VDD VDD.n27 0.0794677
R172 VDD VDD.n24 0.0794677
R173 VDD.n46 VDD.n45 0.0702753
R174 VDD VDD.n31 0.069264
R175 VDD.n36 VDD 0.069264
R176 VDD VDD.n41 0.069264
R177 VDD.n41 VDD 0.0510618
R178 VDD.n15 VDD 0.003875
R179 VDD.n28 VDD 0.00166129
R180 VDD.n25 VDD 0.00166129
R181 VDD VDD.n22 0.00166129
R182 VDD VDD.n19 0.00166129
R183 VDD.n32 VDD 0.00151124
R184 VDD VDD.n35 0.00151124
R185 VDD.n42 VDD 0.00151124
R186 VDD.n45 VDD 0.00151124
R187 Vdiv2.n4 Vdiv2.t4 36.935
R188 Vdiv2.n6 Vdiv2.t6 31.528
R189 Vdiv2.n4 Vdiv2.t3 18.1962
R190 Vdiv2.n6 Vdiv2.t5 15.3826
R191 Vdiv2.n3 Vdiv2.n0 7.09905
R192 Vdiv2.n7 Vdiv2.n6 6.86134
R193 Vdiv2.n8 Vdiv2.n5 5.01116
R194 Vdiv2.n3 Vdiv2.n2 3.25085
R195 Vdiv2.n10 Vdiv2.n9 2.33232
R196 Vdiv2.n2 Vdiv2.t1 2.2755
R197 Vdiv2.n2 Vdiv2.n1 2.2755
R198 Vdiv2.n5 Vdiv2.n4 2.13398
R199 Vdiv2.n9 Vdiv2.n8 1.35708
R200 Vdiv2.n8 Vdiv2.n7 1.12056
R201 Vdiv2.n9 Vdiv2 0.41675
R202 Vdiv2.n10 Vdiv2.n3 0.0919062
R203 Vdiv2.n7 Vdiv2 0.0857632
R204 Vdiv2.n5 Vdiv2 0.0810725
R205 Vdiv2 Vdiv2.n10 0.073625
R206 CLK.n10 CLK.t5 36.935
R207 CLK.n3 CLK.t0 36.935
R208 CLK.n0 CLK.t4 25.5361
R209 CLK.n10 CLK.t3 18.1962
R210 CLK.n3 CLK.t2 18.1962
R211 CLK.n0 CLK.t1 14.0734
R212 CLK.n13 CLK.n12 2.25107
R213 CLK.n16 CLK.n15 2.24235
R214 CLK.n4 CLK.n3 2.12175
R215 CLK.n11 CLK.n10 2.12075
R216 CLK.n8 CLK.n7 1.74297
R217 CLK.n7 CLK.n5 1.49778
R218 CLK.n1 CLK.n0 1.42775
R219 CLK.n15 CLK.n13 0.97145
R220 CLK CLK.n17 0.1605
R221 CLK.n9 CLK 0.0473512
R222 CLK.n2 CLK 0.0473512
R223 CLK.n12 CLK.n9 0.0361897
R224 CLK.n5 CLK.n2 0.0361897
R225 CLK.n17 CLK.n16 0.03175
R226 CLK.n15 CLK.n14 0.0246174
R227 CLK.n7 CLK.n6 0.0131772
R228 CLK.n13 CLK.n8 0.0122182
R229 CLK.n12 CLK.n11 0.00515517
R230 CLK.n5 CLK.n4 0.00515517
R231 CLK.n16 CLK.n1 0.00175
C0 CLK a_1288_1433# 6.43e-21
C1 m2_n31_595# m1_n31_595# 0.021f
C2 VDD JK_FF_mag_0.nand3_mag_1.IN1 0.656f
C3 RST JK_FF_mag_0.nand2_mag_4.IN2 2.17e-19
C4 JK_FF_mag_0.nand2_mag_3.IN1 a_724_1389# 0.00119f
C5 a_1282_292# JK_FF_mag_0.nand3_mag_1.OUT 0.0203f
C6 JK_FF_mag_0.nand2_mag_3.IN1 a_1288_1433# 1.43e-19
C7 Vdiv2 JK_FF_mag_0.nand3_mag_1.IN1 0.00335f
C8 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C9 JK_FF_mag_0.nand2_mag_1.IN2 CLK 1.48e-20
C10 VDD Vdiv2 1.06f
C11 JK_FF_mag_0.nand3_mag_0.OUT VDD 0.758f
C12 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.QB 0.103f
C13 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C14 JK_FF_mag_0.nand2_mag_3.IN1 a_1852_1433# 0.011f
C15 RST JK_FF_mag_0.nand3_mag_1.OUT 0.253f
C16 VDD a_564_1389# 0.00492f
C17 JK_FF_mag_0.nand3_mag_0.OUT Vdiv2 7.24e-19
C18 a_1282_292# JK_FF_mag_0.nand3_mag_2.OUT 9.1e-19
C19 a_1288_1433# JK_FF_mag_0.nand3_mag_1.IN1 0.0697f
C20 JK_FF_mag_0.nand3_mag_0.OUT a_564_1389# 0.0203f
C21 a_1288_1433# VDD 3.18e-19
C22 CLK JK_FF_mag_0.QB 0.307f
C23 a_1442_292# JK_FF_mag_0.QB 0.00696f
C24 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand3_mag_1.IN1 0.109f
C25 a_1852_1433# JK_FF_mag_0.nand3_mag_1.IN1 0.0059f
C26 RST JK_FF_mag_0.nand3_mag_2.OUT 0.0816f
C27 a_724_1389# Vdiv2 2.79e-20
C28 JK_FF_mag_0.nand3_mag_0.OUT a_724_1389# 0.0732f
C29 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.QB 0.28f
C30 JK_FF_mag_0.nand3_mag_0.OUT a_1288_1433# 0.00378f
C31 JK_FF_mag_0.nand2_mag_1.IN2 VDD 0.402f
C32 a_1852_1433# VDD 3.18e-19
C33 a_1282_292# a_1442_292# 0.0504f
C34 a_724_1389# a_564_1389# 0.0504f
C35 JK_FF_mag_0.QB a_2570_336# 0.0811f
C36 a_558_292# RST 0.00188f
C37 JK_FF_mag_0.nand2_mag_1.IN2 Vdiv2 0.107f
C38 RST CLK 0.0415f
C39 RST a_1442_292# 0.00153f
C40 JK_FF_mag_0.nand2_mag_3.IN1 a_2416_1433# 0.00118f
C41 JK_FF_mag_0.QB JK_FF_mag_0.nand3_mag_1.IN1 0.0386f
C42 JK_FF_mag_0.nand2_mag_3.IN1 RST 0.00463f
C43 JK_FF_mag_0.QB VDD 0.907f
C44 a_718_292# RST 0.00188f
C45 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.QB 0.343f
C46 JK_FF_mag_0.QB Vdiv2 1.94f
C47 a_1282_292# VDD 2.21e-19
C48 JK_FF_mag_0.nand2_mag_1.IN2 a_1852_1433# 0.069f
C49 RST JK_FF_mag_0.nand3_mag_1.IN1 0.152f
C50 a_2416_1433# VDD 3.6e-19
C51 a_1282_292# Vdiv2 0.0102f
C52 RST VDD 0.32f
C53 a_2416_1433# Vdiv2 0.069f
C54 JK_FF_mag_0.QB a_724_1389# 0.00392f
C55 JK_FF_mag_0.QB a_1288_1433# 3e-19
C56 JK_FF_mag_0.nand3_mag_0.OUT RST 0.00531f
C57 RST Vdiv2 0.0427f
C58 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.QB 0.0592f
C59 RST a_564_1389# 9.23e-19
C60 a_1852_1433# JK_FF_mag_0.QB 2.96e-19
C61 m2_n31_595# CLK 6.19e-19
C62 RST a_724_1389# 7.69e-19
C63 RST a_1288_1433# 3.11e-19
C64 JK_FF_mag_0.nand2_mag_4.IN2 a_2006_336# 0.069f
C65 JK_FF_mag_0.nand2_mag_1.IN2 a_2416_1433# 0.00372f
C66 m1_n31_595# CLK 2.36e-20
C67 JK_FF_mag_0.nand3_mag_1.OUT a_2006_336# 0.00378f
C68 a_1282_292# JK_FF_mag_0.QB 0.00695f
C69 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand3_mag_1.OUT 0.122f
C70 a_2416_1433# JK_FF_mag_0.QB 0.0114f
C71 m2_n31_595# VDD 0.0194f
C72 RST JK_FF_mag_0.QB 0.0996f
C73 m1_n31_595# VDD 6.13e-19
C74 a_1282_292# RST 0.0017f
C75 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C76 JK_FF_mag_0.nand2_mag_3.IN1 a_2006_336# 0.0036f
C77 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C78 a_558_292# JK_FF_mag_0.nand3_mag_1.OUT 1.17e-20
C79 JK_FF_mag_0.nand2_mag_4.IN2 a_2570_336# 0.00372f
C80 CLK JK_FF_mag_0.nand3_mag_1.OUT 6.64e-19
C81 a_1442_292# JK_FF_mag_0.nand3_mag_1.OUT 0.0733f
C82 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand3_mag_1.OUT 0.16f
C83 a_2006_336# VDD 3.14e-19
C84 a_558_292# JK_FF_mag_0.nand3_mag_2.OUT 0.0202f
C85 a_718_292# JK_FF_mag_0.nand3_mag_1.OUT 1.5e-20
C86 a_2006_336# Vdiv2 0.00859f
C87 JK_FF_mag_0.nand2_mag_4.IN2 VDD 0.391f
C88 JK_FF_mag_0.nand3_mag_2.OUT CLK 0.235f
C89 JK_FF_mag_0.nand3_mag_2.OUT a_1442_292# 2.88e-20
C90 JK_FF_mag_0.nand2_mag_4.IN2 Vdiv2 0.0635f
C91 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand3_mag_2.OUT 0.00118f
C92 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C93 m2_n31_595# RST 0.0301f
C94 a_558_292# CLK 0.00117f
C95 JK_FF_mag_0.nand3_mag_1.OUT VDD 0.995f
C96 a_718_292# JK_FF_mag_0.nand3_mag_2.OUT 0.0731f
C97 m1_n31_595# RST 7.56e-19
C98 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C99 JK_FF_mag_0.nand3_mag_1.OUT Vdiv2 0.0343f
C100 JK_FF_mag_0.nand2_mag_3.IN1 CLK 0.406f
C101 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.nand3_mag_1.IN1 0.00165f
C102 a_558_292# a_718_292# 0.0504f
C103 JK_FF_mag_0.nand3_mag_2.OUT VDD 0.747f
C104 a_718_292# CLK 0.00164f
C105 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C106 JK_FF_mag_0.nand3_mag_1.OUT a_1288_1433# 0.0202f
C107 JK_FF_mag_0.nand3_mag_2.OUT Vdiv2 0.338f
C108 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C109 JK_FF_mag_0.nand2_mag_3.IN1 a_718_292# 1.46e-19
C110 CLK JK_FF_mag_0.nand3_mag_1.IN1 9.71e-20
C111 a_558_292# VDD 0.00108f
C112 a_1442_292# JK_FF_mag_0.nand3_mag_1.IN1 8.64e-19
C113 JK_FF_mag_0.QB a_2006_336# 0.00964f
C114 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand3_mag_1.OUT 0.00975f
C115 a_1852_1433# JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C116 CLK VDD 1.05f
C117 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand3_mag_1.IN1 0.233f
C118 a_558_292# Vdiv2 0.00335f
C119 JK_FF_mag_0.QB JK_FF_mag_0.nand2_mag_4.IN2 0.199f
C120 JK_FF_mag_0.nand2_mag_3.IN1 VDD 1.21f
C121 CLK Vdiv2 0.149f
C122 JK_FF_mag_0.nand3_mag_0.OUT CLK 0.267f
C123 a_1442_292# Vdiv2 0.0101f
C124 VDD a_2570_336# 3.14e-19
C125 CLK a_564_1389# 0.0101f
C126 JK_FF_mag_0.nand2_mag_3.IN1 Vdiv2 0.0168f
C127 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand3_mag_0.OUT 0.0889f
C128 Vdiv2 a_2570_336# 0.0157f
C129 JK_FF_mag_0.QB JK_FF_mag_0.nand3_mag_1.OUT 0.25f
C130 a_718_292# Vdiv2 0.00789f
C131 a_2416_1433# JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C132 CLK a_724_1389# 0.00939f
C133 m2_n31_595# VSS 0.0654f $ **FLOATING
C134 m1_n31_595# VSS 0.15f $ **FLOATING
C135 a_2570_336# VSS 0.0675f
C136 a_2006_336# VSS 0.0676f
C137 a_1442_292# VSS 0.0343f
C138 a_1282_292# VSS 0.0881f
C139 a_718_292# VSS 0.0343f
C140 a_558_292# VSS 0.0881f
C141 JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.416f
C142 RST VSS 0.595f
C143 JK_FF_mag_0.nand3_mag_2.OUT VSS 0.54f
C144 a_2416_1433# VSS 0.0676f
C145 a_1852_1433# VSS 0.0676f
C146 a_1288_1433# VSS 0.0676f
C147 a_724_1389# VSS 0.0343f
C148 a_564_1389# VSS 0.0881f
C149 Vdiv2 VSS 1.64f
C150 JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C151 JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.958f
C152 JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.725f
C153 JK_FF_mag_0.nand3_mag_1.OUT VSS 0.81f
C154 JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C155 JK_FF_mag_0.QB VSS 0.918f
C156 CLK VSS 0.926f
C157 VDD VSS 13.4f
.ends

