magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2045 -2045 2045 2045
<< psubdiff >>
rect -45 23 45 45
rect -45 -23 -23 23
rect 23 -23 45 23
rect -45 -45 45 -23
<< psubdiffcont >>
rect -23 -23 23 23
<< metal1 >>
rect -34 23 34 34
rect -34 -23 -23 23
rect 23 -23 34 23
rect -34 -34 34 -23
<< end >>
