magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1382 -1019 986 1019
<< metal3 >>
rect -382 14 -14 19
rect -382 -14 -377 14
rect -349 -14 -311 14
rect -283 -14 -245 14
rect -217 -14 -179 14
rect -151 -14 -113 14
rect -85 -14 -47 14
rect -19 -14 -14 14
rect -382 -19 -14 -14
<< via3 >>
rect -377 -14 -349 14
rect -311 -14 -283 14
rect -245 -14 -217 14
rect -179 -14 -151 14
rect -113 -14 -85 14
rect -47 -14 -19 14
<< metal4 >>
rect -382 14 -14 19
rect -382 -14 -377 14
rect -349 -14 -311 14
rect -283 -14 -245 14
rect -217 -14 -179 14
rect -151 -14 -113 14
rect -85 -14 -47 14
rect -19 -14 -14 14
rect -382 -19 -14 -14
<< end >>
