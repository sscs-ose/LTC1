* NGSPICE file created from Tr_Gate_flat.ext - technology: gf180mcuC

.subckt Tr_Gate_flat VSS OUT IN CLK VDD
X0 IN a_105_n678.t6 OUT.t3 VDD.t0 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X1 IN CLK.t0 OUT.t7 VSS.t3 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X2 OUT a_105_n678.t7 IN.t2 VDD.t5 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X3 VDD CLK.t2 a_105_n678.t4 VDD.t3 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X4 VSS CLK.t3 a_105_n678.t1 VSS.t3 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X5 VDD CLK.t5 a_105_n678.t0 VDD.t0 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X6 OUT a_105_n678.t8 IN.t1 VDD.t4 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X7 OUT CLK.t6 IN.t5 VSS.t1 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X8 IN CLK.t7 OUT.t6 VSS.t0 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X9 IN a_105_n678.t9 OUT.t2 VDD.t3 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X10 IN CLK.t9 OUT.t4 VSS.t0 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
R0 a_105_n678.n0 a_105_n678.t7 29.2961
R1 a_105_n678.n1 a_105_n678.n0 21.9292
R2 a_105_n678.n2 a_105_n678.n1 18.1271
R3 a_105_n678.n2 a_105_n678.t6 11.1695
R4 a_105_n678.n0 a_105_n678.t9 6.1325
R5 a_105_n678.n1 a_105_n678.t8 6.1325
R6 a_105_n678.n6 a_105_n678.n5 4.93252
R7 a_105_n678.n6 a_105_n678.t1 4.70348
R8 a_105_n678.n8 a_105_n678.n2 4.6311
R9 a_105_n678.n10 a_105_n678.n8 2.85093
R10 a_105_n678.n4 a_105_n678.t4 2.16717
R11 a_105_n678.n4 a_105_n678.n3 2.16717
R12 a_105_n678.t0 a_105_n678.n10 2.16717
R13 a_105_n678.n10 a_105_n678.n9 2.16717
R14 a_105_n678.n7 a_105_n678.n6 1.58582
R15 a_105_n678.n7 a_105_n678.n4 1.24371
R16 a_105_n678.n8 a_105_n678.n7 0.971051
R17 OUT.n6 OUT.t7 6.74332
R18 OUT.n7 OUT.t6 5.1005
R19 OUT.n4 OUT.n1 3.57508
R20 OUT.n6 OUT.n5 3.40011
R21 OUT.n8 OUT.t4 3.00158
R22 OUT OUT.n9 2.58112
R23 OUT.n3 OUT.t3 2.16717
R24 OUT.n3 OUT.n2 2.16717
R25 OUT.n1 OUT.t2 2.16717
R26 OUT.n1 OUT.n0 2.16717
R27 OUT.n9 OUT.n8 1.84821
R28 OUT.n4 OUT.n3 1.25233
R29 OUT.n9 OUT.n4 1.12554
R30 OUT.n8 OUT.n7 0.445613
R31 OUT.n7 OUT.n6 0.11326
R32 IN.n2 IN.t2 5.81586
R33 IN.n10 IN.n7 5.10148
R34 IN.n6 IN.n5 5.10116
R35 IN.n4 IN.n3 5.08021
R36 IN.n10 IN.n9 4.66166
R37 IN.n2 IN.n1 2.85093
R38 IN IN.n11 2.36593
R39 IN.n1 IN.t1 2.16717
R40 IN.n1 IN.n0 2.16717
R41 IN.n9 IN.t5 1.9505
R42 IN.n9 IN.n8 1.9505
R43 IN.n4 IN.n2 0.644196
R44 IN.n6 IN.n4 0.450839
R45 IN.n11 IN.n10 0.358498
R46 IN.n11 IN.n6 0.229792
R47 VDD.n10 VDD.t3 104.945
R48 VDD.n10 VDD.t4 100.909
R49 VDD.n6 VDD.t0 84.7634
R50 VDD.n8 VDD.t5 49.4444
R51 VDD.n7 VDD.n6 6.3005
R52 VDD.n2 VDD.t9 5.77744
R53 VDD.n4 VDD.n3 5.07264
R54 VDD.n12 VDD.n8 3.68253
R55 VDD.n12 VDD.n11 3.1505
R56 VDD.n11 VDD.n10 3.1505
R57 VDD.n2 VDD.n1 2.87637
R58 VDD.n1 VDD.t6 2.16717
R59 VDD.n1 VDD.n0 2.16717
R60 VDD.n4 VDD.n2 0.6395
R61 VDD VDD.n7 0.173395
R62 VDD.n7 VDD.n5 0.1355
R63 VDD.n5 VDD.n4 0.0893158
R64 VDD.n11 VDD.n9 0.0833947
R65 VDD VDD.n12 0.00128947
R66 CLK.n3 CLK.t7 45.6363
R67 CLK.n0 CLK.t5 29.6446
R68 CLK.t1 CLK.n1 29.6446
R69 CLK.n2 CLK.t8 24.6117
R70 CLK.n1 CLK.n0 22.2047
R71 CLK.t7 CLK.t9 22.1925
R72 CLK.n4 CLK.n3 20.9314
R73 CLK CLK.t1 18.5191
R74 CLK.n2 CLK.t3 6.1325
R75 CLK.n0 CLK.t4 6.1325
R76 CLK.n1 CLK.t2 6.1325
R77 CLK.n3 CLK.t6 6.1325
R78 CLK.n4 CLK.t0 6.1325
R79 CLK.n5 CLK.n4 5.38991
R80 CLK.n5 CLK.n2 4.83094
R81 CLK CLK.n5 0.658318
R82 VSS.n12 VSS.t1 292.541
R83 VSS.n15 VSS.t3 189.34
R84 VSS.n2 VSS.t0 108.201
R85 VSS.n7 VSS.n6 5.2005
R86 VSS.n6 VSS.n5 5.2005
R87 VSS.n10 VSS.n9 5.2005
R88 VSS.n9 VSS.n8 5.2005
R89 VSS.n4 VSS.n1 4.88525
R90 VSS.n4 VSS.n3 4.5005
R91 VSS.n3 VSS.n2 4.5005
R92 VSS VSS.n15 3.34763
R93 VSS.n14 VSS.n13 2.6005
R94 VSS.n13 VSS.n12 2.6005
R95 VSS.n1 VSS.t2 2.02837
R96 VSS.n1 VSS.n0 1.80405
R97 VSS.n13 VSS.n11 0.512695
R98 VSS.n14 VSS.n10 0.151571
R99 VSS.n7 VSS.n4 0.028625
R100 VSS.n10 VSS.n7 0.0101429
R101 VSS VSS.n14 0.00532143
C0 IN VDD 0.108f
C1 IN OUT 1.19f
C2 CLK IN 0.487f
C3 OUT VDD 0.0834f
C4 CLK VDD 1f
C5 CLK OUT 0.385f
.ends

