magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1184 -1283 1184 1283
<< metal1 >>
rect -184 277 184 283
rect -184 251 -178 277
rect -152 251 -112 277
rect -86 251 -46 277
rect -20 251 20 277
rect 46 251 86 277
rect 112 251 152 277
rect 178 251 184 277
rect -184 211 184 251
rect -184 185 -178 211
rect -152 185 -112 211
rect -86 185 -46 211
rect -20 185 20 211
rect 46 185 86 211
rect 112 185 152 211
rect 178 185 184 211
rect -184 145 184 185
rect -184 119 -178 145
rect -152 119 -112 145
rect -86 119 -46 145
rect -20 119 20 145
rect 46 119 86 145
rect 112 119 152 145
rect 178 119 184 145
rect -184 79 184 119
rect -184 53 -178 79
rect -152 53 -112 79
rect -86 53 -46 79
rect -20 53 20 79
rect 46 53 86 79
rect 112 53 152 79
rect 178 53 184 79
rect -184 13 184 53
rect -184 -13 -178 13
rect -152 -13 -112 13
rect -86 -13 -46 13
rect -20 -13 20 13
rect 46 -13 86 13
rect 112 -13 152 13
rect 178 -13 184 13
rect -184 -53 184 -13
rect -184 -79 -178 -53
rect -152 -79 -112 -53
rect -86 -79 -46 -53
rect -20 -79 20 -53
rect 46 -79 86 -53
rect 112 -79 152 -53
rect 178 -79 184 -53
rect -184 -119 184 -79
rect -184 -145 -178 -119
rect -152 -145 -112 -119
rect -86 -145 -46 -119
rect -20 -145 20 -119
rect 46 -145 86 -119
rect 112 -145 152 -119
rect 178 -145 184 -119
rect -184 -185 184 -145
rect -184 -211 -178 -185
rect -152 -211 -112 -185
rect -86 -211 -46 -185
rect -20 -211 20 -185
rect 46 -211 86 -185
rect 112 -211 152 -185
rect 178 -211 184 -185
rect -184 -251 184 -211
rect -184 -277 -178 -251
rect -152 -277 -112 -251
rect -86 -277 -46 -251
rect -20 -277 20 -251
rect 46 -277 86 -251
rect 112 -277 152 -251
rect 178 -277 184 -251
rect -184 -283 184 -277
<< via1 >>
rect -178 251 -152 277
rect -112 251 -86 277
rect -46 251 -20 277
rect 20 251 46 277
rect 86 251 112 277
rect 152 251 178 277
rect -178 185 -152 211
rect -112 185 -86 211
rect -46 185 -20 211
rect 20 185 46 211
rect 86 185 112 211
rect 152 185 178 211
rect -178 119 -152 145
rect -112 119 -86 145
rect -46 119 -20 145
rect 20 119 46 145
rect 86 119 112 145
rect 152 119 178 145
rect -178 53 -152 79
rect -112 53 -86 79
rect -46 53 -20 79
rect 20 53 46 79
rect 86 53 112 79
rect 152 53 178 79
rect -178 -13 -152 13
rect -112 -13 -86 13
rect -46 -13 -20 13
rect 20 -13 46 13
rect 86 -13 112 13
rect 152 -13 178 13
rect -178 -79 -152 -53
rect -112 -79 -86 -53
rect -46 -79 -20 -53
rect 20 -79 46 -53
rect 86 -79 112 -53
rect 152 -79 178 -53
rect -178 -145 -152 -119
rect -112 -145 -86 -119
rect -46 -145 -20 -119
rect 20 -145 46 -119
rect 86 -145 112 -119
rect 152 -145 178 -119
rect -178 -211 -152 -185
rect -112 -211 -86 -185
rect -46 -211 -20 -185
rect 20 -211 46 -185
rect 86 -211 112 -185
rect 152 -211 178 -185
rect -178 -277 -152 -251
rect -112 -277 -86 -251
rect -46 -277 -20 -251
rect 20 -277 46 -251
rect 86 -277 112 -251
rect 152 -277 178 -251
<< metal2 >>
rect -184 277 184 283
rect -184 251 -178 277
rect -152 251 -112 277
rect -86 251 -46 277
rect -20 251 20 277
rect 46 251 86 277
rect 112 251 152 277
rect 178 251 184 277
rect -184 211 184 251
rect -184 185 -178 211
rect -152 185 -112 211
rect -86 185 -46 211
rect -20 185 20 211
rect 46 185 86 211
rect 112 185 152 211
rect 178 185 184 211
rect -184 145 184 185
rect -184 119 -178 145
rect -152 119 -112 145
rect -86 119 -46 145
rect -20 119 20 145
rect 46 119 86 145
rect 112 119 152 145
rect 178 119 184 145
rect -184 79 184 119
rect -184 53 -178 79
rect -152 53 -112 79
rect -86 53 -46 79
rect -20 53 20 79
rect 46 53 86 79
rect 112 53 152 79
rect 178 53 184 79
rect -184 13 184 53
rect -184 -13 -178 13
rect -152 -13 -112 13
rect -86 -13 -46 13
rect -20 -13 20 13
rect 46 -13 86 13
rect 112 -13 152 13
rect 178 -13 184 13
rect -184 -53 184 -13
rect -184 -79 -178 -53
rect -152 -79 -112 -53
rect -86 -79 -46 -53
rect -20 -79 20 -53
rect 46 -79 86 -53
rect 112 -79 152 -53
rect 178 -79 184 -53
rect -184 -119 184 -79
rect -184 -145 -178 -119
rect -152 -145 -112 -119
rect -86 -145 -46 -119
rect -20 -145 20 -119
rect 46 -145 86 -119
rect 112 -145 152 -119
rect 178 -145 184 -119
rect -184 -185 184 -145
rect -184 -211 -178 -185
rect -152 -211 -112 -185
rect -86 -211 -46 -185
rect -20 -211 20 -185
rect 46 -211 86 -185
rect 112 -211 152 -185
rect 178 -211 184 -185
rect -184 -251 184 -211
rect -184 -277 -178 -251
rect -152 -277 -112 -251
rect -86 -277 -46 -251
rect -20 -277 20 -251
rect 46 -277 86 -251
rect 112 -277 152 -251
rect 178 -277 184 -251
rect -184 -283 184 -277
<< end >>
