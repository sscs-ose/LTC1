magic
tech gf180mcuC
magscale 1 10
timestamp 1699956126
<< pwell >>
rect -162 -368 162 368
<< nmos >>
rect -50 -300 50 300
<< ndiff >>
rect -138 287 -50 300
rect -138 -287 -125 287
rect -79 -287 -50 287
rect -138 -300 -50 -287
rect 50 287 138 300
rect 50 -287 79 287
rect 125 -287 138 287
rect 50 -300 138 -287
<< ndiffc >>
rect -125 -287 -79 287
rect 79 -287 125 287
<< polysilicon >>
rect -50 300 50 344
rect -50 -344 50 -300
<< metal1 >>
rect -125 287 -79 298
rect -125 -298 -79 -287
rect 79 287 125 298
rect 79 -298 125 -287
<< properties >>
string gencell nfet_03v3
string library gf180mcu
string parameters w 3 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
