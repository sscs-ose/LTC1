magic
tech gf180mcuC
magscale 1 10
timestamp 1694754755
<< nwell >>
rect 493 -2440 10701 2440
<< nsubdiff >>
rect 543 2377 10651 2394
rect 543 2327 560 2377
rect 606 2331 658 2377
rect 704 2331 756 2377
rect 802 2331 854 2377
rect 900 2331 952 2377
rect 998 2331 1050 2377
rect 1096 2331 1148 2377
rect 1194 2331 1246 2377
rect 1292 2331 1344 2377
rect 1390 2331 1442 2377
rect 1488 2331 1540 2377
rect 1586 2331 1638 2377
rect 1684 2331 1736 2377
rect 1782 2331 1834 2377
rect 1880 2331 1932 2377
rect 1978 2331 2030 2377
rect 2076 2331 2128 2377
rect 2174 2331 2226 2377
rect 2272 2331 2324 2377
rect 2370 2331 2422 2377
rect 2468 2331 2520 2377
rect 2566 2331 2618 2377
rect 2664 2331 2716 2377
rect 2762 2331 2814 2377
rect 2860 2331 2912 2377
rect 2958 2331 3010 2377
rect 3056 2331 3108 2377
rect 3154 2331 3206 2377
rect 3252 2331 3304 2377
rect 3350 2331 3402 2377
rect 3448 2331 3500 2377
rect 3546 2331 3598 2377
rect 3644 2331 3696 2377
rect 3742 2331 3794 2377
rect 3840 2331 3892 2377
rect 3938 2331 3990 2377
rect 4036 2331 4088 2377
rect 4134 2331 4186 2377
rect 4232 2331 4284 2377
rect 4330 2331 4382 2377
rect 4428 2331 4480 2377
rect 4526 2331 4578 2377
rect 4624 2331 4676 2377
rect 4722 2331 4774 2377
rect 4820 2331 4872 2377
rect 4918 2331 4970 2377
rect 5016 2331 5068 2377
rect 5114 2331 5166 2377
rect 5212 2331 5264 2377
rect 5310 2331 5362 2377
rect 5408 2331 5460 2377
rect 5506 2331 5558 2377
rect 5604 2331 5656 2377
rect 5702 2331 5754 2377
rect 5800 2331 5852 2377
rect 5898 2331 5950 2377
rect 5996 2331 6048 2377
rect 6094 2331 6146 2377
rect 6192 2331 6244 2377
rect 6290 2331 6342 2377
rect 6388 2331 6440 2377
rect 6486 2331 6538 2377
rect 6584 2331 6636 2377
rect 6682 2331 6734 2377
rect 6780 2331 6832 2377
rect 6878 2331 6930 2377
rect 6976 2331 7028 2377
rect 7074 2331 7126 2377
rect 7172 2331 7224 2377
rect 7270 2331 7322 2377
rect 7368 2331 7420 2377
rect 7466 2331 7518 2377
rect 7564 2331 7616 2377
rect 7662 2331 7714 2377
rect 7760 2331 7812 2377
rect 7858 2331 7910 2377
rect 7956 2331 8008 2377
rect 8054 2331 8106 2377
rect 8152 2331 8204 2377
rect 8250 2331 8302 2377
rect 8348 2331 8400 2377
rect 8446 2331 8498 2377
rect 8544 2331 8596 2377
rect 8642 2331 8694 2377
rect 8740 2331 8792 2377
rect 8838 2331 8890 2377
rect 8936 2331 8988 2377
rect 9034 2331 9086 2377
rect 9132 2331 9184 2377
rect 9230 2331 9282 2377
rect 9328 2331 9380 2377
rect 9426 2331 9478 2377
rect 9524 2331 9576 2377
rect 9622 2331 9674 2377
rect 9720 2331 9772 2377
rect 9818 2331 9870 2377
rect 9916 2331 9968 2377
rect 10014 2331 10066 2377
rect 10112 2331 10164 2377
rect 10210 2331 10262 2377
rect 10308 2331 10360 2377
rect 10406 2331 10458 2377
rect 10504 2331 10588 2377
rect 606 2327 10588 2331
rect 10634 2327 10651 2377
rect 543 2314 10651 2327
rect 543 2275 623 2314
rect 543 2229 560 2275
rect 606 2229 623 2275
rect 10571 2275 10651 2314
rect 543 2177 623 2229
rect 543 2131 560 2177
rect 606 2131 623 2177
rect 543 2079 623 2131
rect 543 2033 560 2079
rect 606 2033 623 2079
rect 543 1981 623 2033
rect 543 1935 560 1981
rect 606 1935 623 1981
rect 543 1883 623 1935
rect 543 1837 560 1883
rect 606 1837 623 1883
rect 543 1785 623 1837
rect 543 1739 560 1785
rect 606 1739 623 1785
rect 543 1687 623 1739
rect 543 1641 560 1687
rect 606 1641 623 1687
rect 543 1589 623 1641
rect 543 1543 560 1589
rect 606 1543 623 1589
rect 543 1491 623 1543
rect 543 1445 560 1491
rect 606 1445 623 1491
rect 543 1393 623 1445
rect 543 1347 560 1393
rect 606 1347 623 1393
rect 543 1295 623 1347
rect 543 1249 560 1295
rect 606 1249 623 1295
rect 543 1197 623 1249
rect 543 1151 560 1197
rect 606 1151 623 1197
rect 543 1099 623 1151
rect 543 1053 560 1099
rect 606 1053 623 1099
rect 543 1001 623 1053
rect 543 955 560 1001
rect 606 955 623 1001
rect 543 903 623 955
rect 543 857 560 903
rect 606 857 623 903
rect 543 805 623 857
rect 543 759 560 805
rect 606 759 623 805
rect 543 707 623 759
rect 543 661 560 707
rect 606 661 623 707
rect 543 609 623 661
rect 543 563 560 609
rect 606 563 623 609
rect 543 511 623 563
rect 543 465 560 511
rect 606 465 623 511
rect 543 413 623 465
rect 543 367 560 413
rect 606 367 623 413
rect 543 315 623 367
rect 543 269 560 315
rect 606 269 623 315
rect 543 217 623 269
rect 717 2186 10477 2258
rect 717 1606 789 2186
rect 10405 1606 10477 2186
rect 717 1534 10477 1606
rect 717 954 789 1534
rect 10405 954 10477 1534
rect 717 882 10477 954
rect 717 302 789 882
rect 10405 302 10477 882
rect 717 230 10477 302
rect 10571 2229 10588 2275
rect 10634 2229 10651 2275
rect 10571 2177 10651 2229
rect 10571 2131 10588 2177
rect 10634 2131 10651 2177
rect 10571 2079 10651 2131
rect 10571 2033 10588 2079
rect 10634 2033 10651 2079
rect 10571 1981 10651 2033
rect 10571 1935 10588 1981
rect 10634 1935 10651 1981
rect 10571 1883 10651 1935
rect 10571 1837 10588 1883
rect 10634 1837 10651 1883
rect 10571 1785 10651 1837
rect 10571 1739 10588 1785
rect 10634 1739 10651 1785
rect 10571 1687 10651 1739
rect 10571 1641 10588 1687
rect 10634 1641 10651 1687
rect 10571 1589 10651 1641
rect 10571 1543 10588 1589
rect 10634 1543 10651 1589
rect 10571 1491 10651 1543
rect 10571 1445 10588 1491
rect 10634 1445 10651 1491
rect 10571 1393 10651 1445
rect 10571 1347 10588 1393
rect 10634 1347 10651 1393
rect 10571 1295 10651 1347
rect 10571 1249 10588 1295
rect 10634 1249 10651 1295
rect 10571 1197 10651 1249
rect 10571 1151 10588 1197
rect 10634 1151 10651 1197
rect 10571 1099 10651 1151
rect 10571 1053 10588 1099
rect 10634 1053 10651 1099
rect 10571 1001 10651 1053
rect 10571 955 10588 1001
rect 10634 955 10651 1001
rect 10571 903 10651 955
rect 10571 857 10588 903
rect 10634 857 10651 903
rect 10571 805 10651 857
rect 10571 759 10588 805
rect 10634 759 10651 805
rect 10571 707 10651 759
rect 10571 661 10588 707
rect 10634 661 10651 707
rect 10571 609 10651 661
rect 10571 563 10588 609
rect 10634 563 10651 609
rect 10571 511 10651 563
rect 10571 465 10588 511
rect 10634 465 10651 511
rect 10571 413 10651 465
rect 10571 367 10588 413
rect 10634 367 10651 413
rect 10571 315 10651 367
rect 10571 269 10588 315
rect 10634 269 10651 315
rect 543 171 560 217
rect 606 171 623 217
rect 543 136 623 171
rect 10571 217 10651 269
rect 10571 171 10588 217
rect 10634 171 10651 217
rect 10571 136 10651 171
rect 543 119 10651 136
rect 543 73 560 119
rect 606 73 658 119
rect 704 73 756 119
rect 802 73 854 119
rect 900 73 952 119
rect 998 73 1050 119
rect 1096 73 1148 119
rect 1194 73 1246 119
rect 1292 73 1344 119
rect 1390 73 1442 119
rect 1488 73 1540 119
rect 1586 73 1638 119
rect 1684 73 1736 119
rect 1782 73 1834 119
rect 1880 73 1932 119
rect 1978 73 2030 119
rect 2076 73 2128 119
rect 2174 73 2226 119
rect 2272 73 2324 119
rect 2370 73 2422 119
rect 2468 73 2520 119
rect 2566 73 2618 119
rect 2664 73 2716 119
rect 2762 73 2814 119
rect 2860 73 2912 119
rect 2958 73 3010 119
rect 3056 73 3108 119
rect 3154 73 3206 119
rect 3252 73 3304 119
rect 3350 73 3402 119
rect 3448 73 3500 119
rect 3546 73 3598 119
rect 3644 73 3696 119
rect 3742 73 3794 119
rect 3840 73 3892 119
rect 3938 73 3990 119
rect 4036 73 4088 119
rect 4134 73 4186 119
rect 4232 73 4284 119
rect 4330 73 4382 119
rect 4428 73 4480 119
rect 4526 73 4578 119
rect 4624 73 4676 119
rect 4722 73 4774 119
rect 4820 73 4872 119
rect 4918 73 4970 119
rect 5016 73 5068 119
rect 5114 73 5166 119
rect 5212 73 5264 119
rect 5310 73 5362 119
rect 5408 73 5460 119
rect 5506 73 5558 119
rect 5604 73 5656 119
rect 5702 73 5754 119
rect 5800 73 5852 119
rect 5898 73 5950 119
rect 5996 73 6048 119
rect 6094 73 6146 119
rect 6192 73 6244 119
rect 6290 73 6342 119
rect 6388 73 6440 119
rect 6486 73 6538 119
rect 6584 73 6636 119
rect 6682 73 6734 119
rect 6780 73 6832 119
rect 6878 73 6930 119
rect 6976 73 7028 119
rect 7074 73 7126 119
rect 7172 73 7224 119
rect 7270 73 7322 119
rect 7368 73 7420 119
rect 7466 73 7518 119
rect 7564 73 7616 119
rect 7662 73 7714 119
rect 7760 73 7812 119
rect 7858 73 7910 119
rect 7956 73 8008 119
rect 8054 73 8106 119
rect 8152 73 8204 119
rect 8250 73 8302 119
rect 8348 73 8400 119
rect 8446 73 8498 119
rect 8544 73 8596 119
rect 8642 73 8694 119
rect 8740 73 8792 119
rect 8838 73 8890 119
rect 8936 73 8988 119
rect 9034 73 9086 119
rect 9132 73 9184 119
rect 9230 73 9282 119
rect 9328 73 9380 119
rect 9426 73 9478 119
rect 9524 73 9576 119
rect 9622 73 9674 119
rect 9720 73 9772 119
rect 9818 73 9870 119
rect 9916 73 9968 119
rect 10014 73 10066 119
rect 10112 73 10164 119
rect 10210 73 10262 119
rect 10308 73 10360 119
rect 10406 73 10458 119
rect 10504 73 10588 119
rect 10634 73 10651 119
rect 543 56 10651 73
rect 543 -73 10651 -56
rect 543 -119 560 -73
rect 606 -119 658 -73
rect 704 -119 756 -73
rect 802 -119 854 -73
rect 900 -119 952 -73
rect 998 -119 1050 -73
rect 1096 -119 1148 -73
rect 1194 -119 1246 -73
rect 1292 -119 1344 -73
rect 1390 -119 1442 -73
rect 1488 -119 1540 -73
rect 1586 -119 1638 -73
rect 1684 -119 1736 -73
rect 1782 -119 1834 -73
rect 1880 -119 1932 -73
rect 1978 -119 2030 -73
rect 2076 -119 2128 -73
rect 2174 -119 2226 -73
rect 2272 -119 2324 -73
rect 2370 -119 2422 -73
rect 2468 -119 2520 -73
rect 2566 -119 2618 -73
rect 2664 -119 2716 -73
rect 2762 -119 2814 -73
rect 2860 -119 2912 -73
rect 2958 -119 3010 -73
rect 3056 -119 3108 -73
rect 3154 -119 3206 -73
rect 3252 -119 3304 -73
rect 3350 -119 3402 -73
rect 3448 -119 3500 -73
rect 3546 -119 3598 -73
rect 3644 -119 3696 -73
rect 3742 -119 3794 -73
rect 3840 -119 3892 -73
rect 3938 -119 3990 -73
rect 4036 -119 4088 -73
rect 4134 -119 4186 -73
rect 4232 -119 4284 -73
rect 4330 -119 4382 -73
rect 4428 -119 4480 -73
rect 4526 -119 4578 -73
rect 4624 -119 4676 -73
rect 4722 -119 4774 -73
rect 4820 -119 4872 -73
rect 4918 -119 4970 -73
rect 5016 -119 5068 -73
rect 5114 -119 5166 -73
rect 5212 -119 5264 -73
rect 5310 -119 5362 -73
rect 5408 -119 5460 -73
rect 5506 -119 5558 -73
rect 5604 -119 5656 -73
rect 5702 -119 5754 -73
rect 5800 -119 5852 -73
rect 5898 -119 5950 -73
rect 5996 -119 6048 -73
rect 6094 -119 6146 -73
rect 6192 -119 6244 -73
rect 6290 -119 6342 -73
rect 6388 -119 6440 -73
rect 6486 -119 6538 -73
rect 6584 -119 6636 -73
rect 6682 -119 6734 -73
rect 6780 -119 6832 -73
rect 6878 -119 6930 -73
rect 6976 -119 7028 -73
rect 7074 -119 7126 -73
rect 7172 -119 7224 -73
rect 7270 -119 7322 -73
rect 7368 -119 7420 -73
rect 7466 -119 7518 -73
rect 7564 -119 7616 -73
rect 7662 -119 7714 -73
rect 7760 -119 7812 -73
rect 7858 -119 7910 -73
rect 7956 -119 8008 -73
rect 8054 -119 8106 -73
rect 8152 -119 8204 -73
rect 8250 -119 8302 -73
rect 8348 -119 8400 -73
rect 8446 -119 8498 -73
rect 8544 -119 8596 -73
rect 8642 -119 8694 -73
rect 8740 -119 8792 -73
rect 8838 -119 8890 -73
rect 8936 -119 8988 -73
rect 9034 -119 9086 -73
rect 9132 -119 9184 -73
rect 9230 -119 9282 -73
rect 9328 -119 9380 -73
rect 9426 -119 9478 -73
rect 9524 -119 9576 -73
rect 9622 -119 9674 -73
rect 9720 -119 9772 -73
rect 9818 -119 9870 -73
rect 9916 -119 9968 -73
rect 10014 -119 10066 -73
rect 10112 -119 10164 -73
rect 10210 -119 10262 -73
rect 10308 -119 10360 -73
rect 10406 -119 10458 -73
rect 10504 -119 10588 -73
rect 10634 -119 10651 -73
rect 543 -136 10651 -119
rect 543 -171 623 -136
rect 543 -217 560 -171
rect 606 -217 623 -171
rect 543 -269 623 -217
rect 10571 -171 10651 -136
rect 10571 -217 10588 -171
rect 10634 -217 10651 -171
rect 543 -315 560 -269
rect 606 -315 623 -269
rect 543 -367 623 -315
rect 543 -413 560 -367
rect 606 -413 623 -367
rect 543 -465 623 -413
rect 543 -511 560 -465
rect 606 -511 623 -465
rect 543 -563 623 -511
rect 543 -609 560 -563
rect 606 -609 623 -563
rect 543 -661 623 -609
rect 543 -707 560 -661
rect 606 -707 623 -661
rect 543 -759 623 -707
rect 543 -805 560 -759
rect 606 -805 623 -759
rect 543 -857 623 -805
rect 543 -903 560 -857
rect 606 -903 623 -857
rect 543 -955 623 -903
rect 543 -1001 560 -955
rect 606 -1001 623 -955
rect 543 -1053 623 -1001
rect 543 -1099 560 -1053
rect 606 -1099 623 -1053
rect 543 -1151 623 -1099
rect 543 -1197 560 -1151
rect 606 -1197 623 -1151
rect 543 -1249 623 -1197
rect 543 -1295 560 -1249
rect 606 -1295 623 -1249
rect 543 -1347 623 -1295
rect 543 -1393 560 -1347
rect 606 -1393 623 -1347
rect 543 -1445 623 -1393
rect 543 -1491 560 -1445
rect 606 -1491 623 -1445
rect 543 -1543 623 -1491
rect 543 -1589 560 -1543
rect 606 -1589 623 -1543
rect 543 -1641 623 -1589
rect 543 -1687 560 -1641
rect 606 -1687 623 -1641
rect 543 -1739 623 -1687
rect 543 -1785 560 -1739
rect 606 -1785 623 -1739
rect 543 -1837 623 -1785
rect 543 -1883 560 -1837
rect 606 -1883 623 -1837
rect 543 -1935 623 -1883
rect 543 -1981 560 -1935
rect 606 -1981 623 -1935
rect 543 -2033 623 -1981
rect 543 -2079 560 -2033
rect 606 -2079 623 -2033
rect 543 -2131 623 -2079
rect 543 -2177 560 -2131
rect 606 -2177 623 -2131
rect 543 -2229 623 -2177
rect 543 -2275 560 -2229
rect 606 -2275 623 -2229
rect 717 -302 10477 -230
rect 717 -882 789 -302
rect 10405 -882 10477 -302
rect 717 -954 10477 -882
rect 717 -1534 789 -954
rect 10405 -1534 10477 -954
rect 717 -1606 10477 -1534
rect 717 -2186 789 -1606
rect 10405 -2186 10477 -1606
rect 717 -2258 10477 -2186
rect 10571 -269 10651 -217
rect 10571 -315 10588 -269
rect 10634 -315 10651 -269
rect 10571 -367 10651 -315
rect 10571 -413 10588 -367
rect 10634 -413 10651 -367
rect 10571 -465 10651 -413
rect 10571 -511 10588 -465
rect 10634 -511 10651 -465
rect 10571 -563 10651 -511
rect 10571 -609 10588 -563
rect 10634 -609 10651 -563
rect 10571 -661 10651 -609
rect 10571 -707 10588 -661
rect 10634 -707 10651 -661
rect 10571 -759 10651 -707
rect 10571 -805 10588 -759
rect 10634 -805 10651 -759
rect 10571 -857 10651 -805
rect 10571 -903 10588 -857
rect 10634 -903 10651 -857
rect 10571 -955 10651 -903
rect 10571 -1001 10588 -955
rect 10634 -1001 10651 -955
rect 10571 -1053 10651 -1001
rect 10571 -1099 10588 -1053
rect 10634 -1099 10651 -1053
rect 10571 -1151 10651 -1099
rect 10571 -1197 10588 -1151
rect 10634 -1197 10651 -1151
rect 10571 -1249 10651 -1197
rect 10571 -1295 10588 -1249
rect 10634 -1295 10651 -1249
rect 10571 -1347 10651 -1295
rect 10571 -1393 10588 -1347
rect 10634 -1393 10651 -1347
rect 10571 -1445 10651 -1393
rect 10571 -1491 10588 -1445
rect 10634 -1491 10651 -1445
rect 10571 -1543 10651 -1491
rect 10571 -1589 10588 -1543
rect 10634 -1589 10651 -1543
rect 10571 -1641 10651 -1589
rect 10571 -1687 10588 -1641
rect 10634 -1687 10651 -1641
rect 10571 -1739 10651 -1687
rect 10571 -1785 10588 -1739
rect 10634 -1785 10651 -1739
rect 10571 -1837 10651 -1785
rect 10571 -1883 10588 -1837
rect 10634 -1883 10651 -1837
rect 10571 -1935 10651 -1883
rect 10571 -1981 10588 -1935
rect 10634 -1981 10651 -1935
rect 10571 -2033 10651 -1981
rect 10571 -2079 10588 -2033
rect 10634 -2079 10651 -2033
rect 10571 -2131 10651 -2079
rect 10571 -2177 10588 -2131
rect 10634 -2177 10651 -2131
rect 10571 -2229 10651 -2177
rect 543 -2314 623 -2275
rect 10571 -2275 10588 -2229
rect 10634 -2275 10651 -2229
rect 10571 -2314 10651 -2275
rect 543 -2327 10651 -2314
rect 543 -2377 560 -2327
rect 606 -2331 10588 -2327
rect 606 -2377 658 -2331
rect 704 -2377 756 -2331
rect 802 -2377 854 -2331
rect 900 -2377 952 -2331
rect 998 -2377 1050 -2331
rect 1096 -2377 1148 -2331
rect 1194 -2377 1246 -2331
rect 1292 -2377 1344 -2331
rect 1390 -2377 1442 -2331
rect 1488 -2377 1540 -2331
rect 1586 -2377 1638 -2331
rect 1684 -2377 1736 -2331
rect 1782 -2377 1834 -2331
rect 1880 -2377 1932 -2331
rect 1978 -2377 2030 -2331
rect 2076 -2377 2128 -2331
rect 2174 -2377 2226 -2331
rect 2272 -2377 2324 -2331
rect 2370 -2377 2422 -2331
rect 2468 -2377 2520 -2331
rect 2566 -2377 2618 -2331
rect 2664 -2377 2716 -2331
rect 2762 -2377 2814 -2331
rect 2860 -2377 2912 -2331
rect 2958 -2377 3010 -2331
rect 3056 -2377 3108 -2331
rect 3154 -2377 3206 -2331
rect 3252 -2377 3304 -2331
rect 3350 -2377 3402 -2331
rect 3448 -2377 3500 -2331
rect 3546 -2377 3598 -2331
rect 3644 -2377 3696 -2331
rect 3742 -2377 3794 -2331
rect 3840 -2377 3892 -2331
rect 3938 -2377 3990 -2331
rect 4036 -2377 4088 -2331
rect 4134 -2377 4186 -2331
rect 4232 -2377 4284 -2331
rect 4330 -2377 4382 -2331
rect 4428 -2377 4480 -2331
rect 4526 -2377 4578 -2331
rect 4624 -2377 4676 -2331
rect 4722 -2377 4774 -2331
rect 4820 -2377 4872 -2331
rect 4918 -2377 4970 -2331
rect 5016 -2377 5068 -2331
rect 5114 -2377 5166 -2331
rect 5212 -2377 5264 -2331
rect 5310 -2377 5362 -2331
rect 5408 -2377 5460 -2331
rect 5506 -2377 5558 -2331
rect 5604 -2377 5656 -2331
rect 5702 -2377 5754 -2331
rect 5800 -2377 5852 -2331
rect 5898 -2377 5950 -2331
rect 5996 -2377 6048 -2331
rect 6094 -2377 6146 -2331
rect 6192 -2377 6244 -2331
rect 6290 -2377 6342 -2331
rect 6388 -2377 6440 -2331
rect 6486 -2377 6538 -2331
rect 6584 -2377 6636 -2331
rect 6682 -2377 6734 -2331
rect 6780 -2377 6832 -2331
rect 6878 -2377 6930 -2331
rect 6976 -2377 7028 -2331
rect 7074 -2377 7126 -2331
rect 7172 -2377 7224 -2331
rect 7270 -2377 7322 -2331
rect 7368 -2377 7420 -2331
rect 7466 -2377 7518 -2331
rect 7564 -2377 7616 -2331
rect 7662 -2377 7714 -2331
rect 7760 -2377 7812 -2331
rect 7858 -2377 7910 -2331
rect 7956 -2377 8008 -2331
rect 8054 -2377 8106 -2331
rect 8152 -2377 8204 -2331
rect 8250 -2377 8302 -2331
rect 8348 -2377 8400 -2331
rect 8446 -2377 8498 -2331
rect 8544 -2377 8596 -2331
rect 8642 -2377 8694 -2331
rect 8740 -2377 8792 -2331
rect 8838 -2377 8890 -2331
rect 8936 -2377 8988 -2331
rect 9034 -2377 9086 -2331
rect 9132 -2377 9184 -2331
rect 9230 -2377 9282 -2331
rect 9328 -2377 9380 -2331
rect 9426 -2377 9478 -2331
rect 9524 -2377 9576 -2331
rect 9622 -2377 9674 -2331
rect 9720 -2377 9772 -2331
rect 9818 -2377 9870 -2331
rect 9916 -2377 9968 -2331
rect 10014 -2377 10066 -2331
rect 10112 -2377 10164 -2331
rect 10210 -2377 10262 -2331
rect 10308 -2377 10360 -2331
rect 10406 -2377 10458 -2331
rect 10504 -2377 10588 -2331
rect 10634 -2377 10651 -2327
rect 543 -2394 10651 -2377
<< nsubdiffcont >>
rect 560 2327 606 2377
rect 658 2331 704 2377
rect 756 2331 802 2377
rect 854 2331 900 2377
rect 952 2331 998 2377
rect 1050 2331 1096 2377
rect 1148 2331 1194 2377
rect 1246 2331 1292 2377
rect 1344 2331 1390 2377
rect 1442 2331 1488 2377
rect 1540 2331 1586 2377
rect 1638 2331 1684 2377
rect 1736 2331 1782 2377
rect 1834 2331 1880 2377
rect 1932 2331 1978 2377
rect 2030 2331 2076 2377
rect 2128 2331 2174 2377
rect 2226 2331 2272 2377
rect 2324 2331 2370 2377
rect 2422 2331 2468 2377
rect 2520 2331 2566 2377
rect 2618 2331 2664 2377
rect 2716 2331 2762 2377
rect 2814 2331 2860 2377
rect 2912 2331 2958 2377
rect 3010 2331 3056 2377
rect 3108 2331 3154 2377
rect 3206 2331 3252 2377
rect 3304 2331 3350 2377
rect 3402 2331 3448 2377
rect 3500 2331 3546 2377
rect 3598 2331 3644 2377
rect 3696 2331 3742 2377
rect 3794 2331 3840 2377
rect 3892 2331 3938 2377
rect 3990 2331 4036 2377
rect 4088 2331 4134 2377
rect 4186 2331 4232 2377
rect 4284 2331 4330 2377
rect 4382 2331 4428 2377
rect 4480 2331 4526 2377
rect 4578 2331 4624 2377
rect 4676 2331 4722 2377
rect 4774 2331 4820 2377
rect 4872 2331 4918 2377
rect 4970 2331 5016 2377
rect 5068 2331 5114 2377
rect 5166 2331 5212 2377
rect 5264 2331 5310 2377
rect 5362 2331 5408 2377
rect 5460 2331 5506 2377
rect 5558 2331 5604 2377
rect 5656 2331 5702 2377
rect 5754 2331 5800 2377
rect 5852 2331 5898 2377
rect 5950 2331 5996 2377
rect 6048 2331 6094 2377
rect 6146 2331 6192 2377
rect 6244 2331 6290 2377
rect 6342 2331 6388 2377
rect 6440 2331 6486 2377
rect 6538 2331 6584 2377
rect 6636 2331 6682 2377
rect 6734 2331 6780 2377
rect 6832 2331 6878 2377
rect 6930 2331 6976 2377
rect 7028 2331 7074 2377
rect 7126 2331 7172 2377
rect 7224 2331 7270 2377
rect 7322 2331 7368 2377
rect 7420 2331 7466 2377
rect 7518 2331 7564 2377
rect 7616 2331 7662 2377
rect 7714 2331 7760 2377
rect 7812 2331 7858 2377
rect 7910 2331 7956 2377
rect 8008 2331 8054 2377
rect 8106 2331 8152 2377
rect 8204 2331 8250 2377
rect 8302 2331 8348 2377
rect 8400 2331 8446 2377
rect 8498 2331 8544 2377
rect 8596 2331 8642 2377
rect 8694 2331 8740 2377
rect 8792 2331 8838 2377
rect 8890 2331 8936 2377
rect 8988 2331 9034 2377
rect 9086 2331 9132 2377
rect 9184 2331 9230 2377
rect 9282 2331 9328 2377
rect 9380 2331 9426 2377
rect 9478 2331 9524 2377
rect 9576 2331 9622 2377
rect 9674 2331 9720 2377
rect 9772 2331 9818 2377
rect 9870 2331 9916 2377
rect 9968 2331 10014 2377
rect 10066 2331 10112 2377
rect 10164 2331 10210 2377
rect 10262 2331 10308 2377
rect 10360 2331 10406 2377
rect 10458 2331 10504 2377
rect 10588 2327 10634 2377
rect 560 2229 606 2275
rect 560 2131 606 2177
rect 560 2033 606 2079
rect 560 1935 606 1981
rect 560 1837 606 1883
rect 560 1739 606 1785
rect 560 1641 606 1687
rect 560 1543 606 1589
rect 560 1445 606 1491
rect 560 1347 606 1393
rect 560 1249 606 1295
rect 560 1151 606 1197
rect 560 1053 606 1099
rect 560 955 606 1001
rect 560 857 606 903
rect 560 759 606 805
rect 560 661 606 707
rect 560 563 606 609
rect 560 465 606 511
rect 560 367 606 413
rect 560 269 606 315
rect 10588 2229 10634 2275
rect 10588 2131 10634 2177
rect 10588 2033 10634 2079
rect 10588 1935 10634 1981
rect 10588 1837 10634 1883
rect 10588 1739 10634 1785
rect 10588 1641 10634 1687
rect 10588 1543 10634 1589
rect 10588 1445 10634 1491
rect 10588 1347 10634 1393
rect 10588 1249 10634 1295
rect 10588 1151 10634 1197
rect 10588 1053 10634 1099
rect 10588 955 10634 1001
rect 10588 857 10634 903
rect 10588 759 10634 805
rect 10588 661 10634 707
rect 10588 563 10634 609
rect 10588 465 10634 511
rect 10588 367 10634 413
rect 10588 269 10634 315
rect 560 171 606 217
rect 10588 171 10634 217
rect 560 73 606 119
rect 658 73 704 119
rect 756 73 802 119
rect 854 73 900 119
rect 952 73 998 119
rect 1050 73 1096 119
rect 1148 73 1194 119
rect 1246 73 1292 119
rect 1344 73 1390 119
rect 1442 73 1488 119
rect 1540 73 1586 119
rect 1638 73 1684 119
rect 1736 73 1782 119
rect 1834 73 1880 119
rect 1932 73 1978 119
rect 2030 73 2076 119
rect 2128 73 2174 119
rect 2226 73 2272 119
rect 2324 73 2370 119
rect 2422 73 2468 119
rect 2520 73 2566 119
rect 2618 73 2664 119
rect 2716 73 2762 119
rect 2814 73 2860 119
rect 2912 73 2958 119
rect 3010 73 3056 119
rect 3108 73 3154 119
rect 3206 73 3252 119
rect 3304 73 3350 119
rect 3402 73 3448 119
rect 3500 73 3546 119
rect 3598 73 3644 119
rect 3696 73 3742 119
rect 3794 73 3840 119
rect 3892 73 3938 119
rect 3990 73 4036 119
rect 4088 73 4134 119
rect 4186 73 4232 119
rect 4284 73 4330 119
rect 4382 73 4428 119
rect 4480 73 4526 119
rect 4578 73 4624 119
rect 4676 73 4722 119
rect 4774 73 4820 119
rect 4872 73 4918 119
rect 4970 73 5016 119
rect 5068 73 5114 119
rect 5166 73 5212 119
rect 5264 73 5310 119
rect 5362 73 5408 119
rect 5460 73 5506 119
rect 5558 73 5604 119
rect 5656 73 5702 119
rect 5754 73 5800 119
rect 5852 73 5898 119
rect 5950 73 5996 119
rect 6048 73 6094 119
rect 6146 73 6192 119
rect 6244 73 6290 119
rect 6342 73 6388 119
rect 6440 73 6486 119
rect 6538 73 6584 119
rect 6636 73 6682 119
rect 6734 73 6780 119
rect 6832 73 6878 119
rect 6930 73 6976 119
rect 7028 73 7074 119
rect 7126 73 7172 119
rect 7224 73 7270 119
rect 7322 73 7368 119
rect 7420 73 7466 119
rect 7518 73 7564 119
rect 7616 73 7662 119
rect 7714 73 7760 119
rect 7812 73 7858 119
rect 7910 73 7956 119
rect 8008 73 8054 119
rect 8106 73 8152 119
rect 8204 73 8250 119
rect 8302 73 8348 119
rect 8400 73 8446 119
rect 8498 73 8544 119
rect 8596 73 8642 119
rect 8694 73 8740 119
rect 8792 73 8838 119
rect 8890 73 8936 119
rect 8988 73 9034 119
rect 9086 73 9132 119
rect 9184 73 9230 119
rect 9282 73 9328 119
rect 9380 73 9426 119
rect 9478 73 9524 119
rect 9576 73 9622 119
rect 9674 73 9720 119
rect 9772 73 9818 119
rect 9870 73 9916 119
rect 9968 73 10014 119
rect 10066 73 10112 119
rect 10164 73 10210 119
rect 10262 73 10308 119
rect 10360 73 10406 119
rect 10458 73 10504 119
rect 10588 73 10634 119
rect 560 -119 606 -73
rect 658 -119 704 -73
rect 756 -119 802 -73
rect 854 -119 900 -73
rect 952 -119 998 -73
rect 1050 -119 1096 -73
rect 1148 -119 1194 -73
rect 1246 -119 1292 -73
rect 1344 -119 1390 -73
rect 1442 -119 1488 -73
rect 1540 -119 1586 -73
rect 1638 -119 1684 -73
rect 1736 -119 1782 -73
rect 1834 -119 1880 -73
rect 1932 -119 1978 -73
rect 2030 -119 2076 -73
rect 2128 -119 2174 -73
rect 2226 -119 2272 -73
rect 2324 -119 2370 -73
rect 2422 -119 2468 -73
rect 2520 -119 2566 -73
rect 2618 -119 2664 -73
rect 2716 -119 2762 -73
rect 2814 -119 2860 -73
rect 2912 -119 2958 -73
rect 3010 -119 3056 -73
rect 3108 -119 3154 -73
rect 3206 -119 3252 -73
rect 3304 -119 3350 -73
rect 3402 -119 3448 -73
rect 3500 -119 3546 -73
rect 3598 -119 3644 -73
rect 3696 -119 3742 -73
rect 3794 -119 3840 -73
rect 3892 -119 3938 -73
rect 3990 -119 4036 -73
rect 4088 -119 4134 -73
rect 4186 -119 4232 -73
rect 4284 -119 4330 -73
rect 4382 -119 4428 -73
rect 4480 -119 4526 -73
rect 4578 -119 4624 -73
rect 4676 -119 4722 -73
rect 4774 -119 4820 -73
rect 4872 -119 4918 -73
rect 4970 -119 5016 -73
rect 5068 -119 5114 -73
rect 5166 -119 5212 -73
rect 5264 -119 5310 -73
rect 5362 -119 5408 -73
rect 5460 -119 5506 -73
rect 5558 -119 5604 -73
rect 5656 -119 5702 -73
rect 5754 -119 5800 -73
rect 5852 -119 5898 -73
rect 5950 -119 5996 -73
rect 6048 -119 6094 -73
rect 6146 -119 6192 -73
rect 6244 -119 6290 -73
rect 6342 -119 6388 -73
rect 6440 -119 6486 -73
rect 6538 -119 6584 -73
rect 6636 -119 6682 -73
rect 6734 -119 6780 -73
rect 6832 -119 6878 -73
rect 6930 -119 6976 -73
rect 7028 -119 7074 -73
rect 7126 -119 7172 -73
rect 7224 -119 7270 -73
rect 7322 -119 7368 -73
rect 7420 -119 7466 -73
rect 7518 -119 7564 -73
rect 7616 -119 7662 -73
rect 7714 -119 7760 -73
rect 7812 -119 7858 -73
rect 7910 -119 7956 -73
rect 8008 -119 8054 -73
rect 8106 -119 8152 -73
rect 8204 -119 8250 -73
rect 8302 -119 8348 -73
rect 8400 -119 8446 -73
rect 8498 -119 8544 -73
rect 8596 -119 8642 -73
rect 8694 -119 8740 -73
rect 8792 -119 8838 -73
rect 8890 -119 8936 -73
rect 8988 -119 9034 -73
rect 9086 -119 9132 -73
rect 9184 -119 9230 -73
rect 9282 -119 9328 -73
rect 9380 -119 9426 -73
rect 9478 -119 9524 -73
rect 9576 -119 9622 -73
rect 9674 -119 9720 -73
rect 9772 -119 9818 -73
rect 9870 -119 9916 -73
rect 9968 -119 10014 -73
rect 10066 -119 10112 -73
rect 10164 -119 10210 -73
rect 10262 -119 10308 -73
rect 10360 -119 10406 -73
rect 10458 -119 10504 -73
rect 10588 -119 10634 -73
rect 560 -217 606 -171
rect 10588 -217 10634 -171
rect 560 -315 606 -269
rect 560 -413 606 -367
rect 560 -511 606 -465
rect 560 -609 606 -563
rect 560 -707 606 -661
rect 560 -805 606 -759
rect 560 -903 606 -857
rect 560 -1001 606 -955
rect 560 -1099 606 -1053
rect 560 -1197 606 -1151
rect 560 -1295 606 -1249
rect 560 -1393 606 -1347
rect 560 -1491 606 -1445
rect 560 -1589 606 -1543
rect 560 -1687 606 -1641
rect 560 -1785 606 -1739
rect 560 -1883 606 -1837
rect 560 -1981 606 -1935
rect 560 -2079 606 -2033
rect 560 -2177 606 -2131
rect 560 -2275 606 -2229
rect 10588 -315 10634 -269
rect 10588 -413 10634 -367
rect 10588 -511 10634 -465
rect 10588 -609 10634 -563
rect 10588 -707 10634 -661
rect 10588 -805 10634 -759
rect 10588 -903 10634 -857
rect 10588 -1001 10634 -955
rect 10588 -1099 10634 -1053
rect 10588 -1197 10634 -1151
rect 10588 -1295 10634 -1249
rect 10588 -1393 10634 -1347
rect 10588 -1491 10634 -1445
rect 10588 -1589 10634 -1543
rect 10588 -1687 10634 -1641
rect 10588 -1785 10634 -1739
rect 10588 -1883 10634 -1837
rect 10588 -1981 10634 -1935
rect 10588 -2079 10634 -2033
rect 10588 -2177 10634 -2131
rect 10588 -2275 10634 -2229
rect 560 -2377 606 -2327
rect 658 -2377 704 -2331
rect 756 -2377 802 -2331
rect 854 -2377 900 -2331
rect 952 -2377 998 -2331
rect 1050 -2377 1096 -2331
rect 1148 -2377 1194 -2331
rect 1246 -2377 1292 -2331
rect 1344 -2377 1390 -2331
rect 1442 -2377 1488 -2331
rect 1540 -2377 1586 -2331
rect 1638 -2377 1684 -2331
rect 1736 -2377 1782 -2331
rect 1834 -2377 1880 -2331
rect 1932 -2377 1978 -2331
rect 2030 -2377 2076 -2331
rect 2128 -2377 2174 -2331
rect 2226 -2377 2272 -2331
rect 2324 -2377 2370 -2331
rect 2422 -2377 2468 -2331
rect 2520 -2377 2566 -2331
rect 2618 -2377 2664 -2331
rect 2716 -2377 2762 -2331
rect 2814 -2377 2860 -2331
rect 2912 -2377 2958 -2331
rect 3010 -2377 3056 -2331
rect 3108 -2377 3154 -2331
rect 3206 -2377 3252 -2331
rect 3304 -2377 3350 -2331
rect 3402 -2377 3448 -2331
rect 3500 -2377 3546 -2331
rect 3598 -2377 3644 -2331
rect 3696 -2377 3742 -2331
rect 3794 -2377 3840 -2331
rect 3892 -2377 3938 -2331
rect 3990 -2377 4036 -2331
rect 4088 -2377 4134 -2331
rect 4186 -2377 4232 -2331
rect 4284 -2377 4330 -2331
rect 4382 -2377 4428 -2331
rect 4480 -2377 4526 -2331
rect 4578 -2377 4624 -2331
rect 4676 -2377 4722 -2331
rect 4774 -2377 4820 -2331
rect 4872 -2377 4918 -2331
rect 4970 -2377 5016 -2331
rect 5068 -2377 5114 -2331
rect 5166 -2377 5212 -2331
rect 5264 -2377 5310 -2331
rect 5362 -2377 5408 -2331
rect 5460 -2377 5506 -2331
rect 5558 -2377 5604 -2331
rect 5656 -2377 5702 -2331
rect 5754 -2377 5800 -2331
rect 5852 -2377 5898 -2331
rect 5950 -2377 5996 -2331
rect 6048 -2377 6094 -2331
rect 6146 -2377 6192 -2331
rect 6244 -2377 6290 -2331
rect 6342 -2377 6388 -2331
rect 6440 -2377 6486 -2331
rect 6538 -2377 6584 -2331
rect 6636 -2377 6682 -2331
rect 6734 -2377 6780 -2331
rect 6832 -2377 6878 -2331
rect 6930 -2377 6976 -2331
rect 7028 -2377 7074 -2331
rect 7126 -2377 7172 -2331
rect 7224 -2377 7270 -2331
rect 7322 -2377 7368 -2331
rect 7420 -2377 7466 -2331
rect 7518 -2377 7564 -2331
rect 7616 -2377 7662 -2331
rect 7714 -2377 7760 -2331
rect 7812 -2377 7858 -2331
rect 7910 -2377 7956 -2331
rect 8008 -2377 8054 -2331
rect 8106 -2377 8152 -2331
rect 8204 -2377 8250 -2331
rect 8302 -2377 8348 -2331
rect 8400 -2377 8446 -2331
rect 8498 -2377 8544 -2331
rect 8596 -2377 8642 -2331
rect 8694 -2377 8740 -2331
rect 8792 -2377 8838 -2331
rect 8890 -2377 8936 -2331
rect 8988 -2377 9034 -2331
rect 9086 -2377 9132 -2331
rect 9184 -2377 9230 -2331
rect 9282 -2377 9328 -2331
rect 9380 -2377 9426 -2331
rect 9478 -2377 9524 -2331
rect 9576 -2377 9622 -2331
rect 9674 -2377 9720 -2331
rect 9772 -2377 9818 -2331
rect 9870 -2377 9916 -2331
rect 9968 -2377 10014 -2331
rect 10066 -2377 10112 -2331
rect 10164 -2377 10210 -2331
rect 10262 -2377 10308 -2331
rect 10360 -2377 10406 -2331
rect 10458 -2377 10504 -2331
rect 10588 -2377 10634 -2327
<< polysilicon >>
rect 877 2085 1077 2098
rect 877 2039 890 2085
rect 1064 2039 1077 2085
rect 877 1996 1077 2039
rect 877 1753 1077 1796
rect 877 1707 890 1753
rect 1064 1707 1077 1753
rect 877 1694 1077 1707
rect 1157 2085 1357 2098
rect 1157 2039 1170 2085
rect 1344 2039 1357 2085
rect 1157 1996 1357 2039
rect 1157 1753 1357 1796
rect 1157 1707 1170 1753
rect 1344 1707 1357 1753
rect 1157 1694 1357 1707
rect 1437 2085 1637 2098
rect 1437 2039 1450 2085
rect 1624 2039 1637 2085
rect 1437 1996 1637 2039
rect 1437 1753 1637 1796
rect 1437 1707 1450 1753
rect 1624 1707 1637 1753
rect 1437 1694 1637 1707
rect 1717 2085 1917 2098
rect 1717 2039 1730 2085
rect 1904 2039 1917 2085
rect 1717 1996 1917 2039
rect 1717 1753 1917 1796
rect 1717 1707 1730 1753
rect 1904 1707 1917 1753
rect 1717 1694 1917 1707
rect 1997 2085 2197 2098
rect 1997 2039 2010 2085
rect 2184 2039 2197 2085
rect 1997 1996 2197 2039
rect 1997 1753 2197 1796
rect 1997 1707 2010 1753
rect 2184 1707 2197 1753
rect 1997 1694 2197 1707
rect 2277 2085 2477 2098
rect 2277 2039 2290 2085
rect 2464 2039 2477 2085
rect 2277 1996 2477 2039
rect 2277 1753 2477 1796
rect 2277 1707 2290 1753
rect 2464 1707 2477 1753
rect 2277 1694 2477 1707
rect 2557 2085 2757 2098
rect 2557 2039 2570 2085
rect 2744 2039 2757 2085
rect 2557 1996 2757 2039
rect 2557 1753 2757 1796
rect 2557 1707 2570 1753
rect 2744 1707 2757 1753
rect 2557 1694 2757 1707
rect 2837 2085 3037 2098
rect 2837 2039 2850 2085
rect 3024 2039 3037 2085
rect 2837 1996 3037 2039
rect 2837 1753 3037 1796
rect 2837 1707 2850 1753
rect 3024 1707 3037 1753
rect 2837 1694 3037 1707
rect 3117 2085 3317 2098
rect 3117 2039 3130 2085
rect 3304 2039 3317 2085
rect 3117 1996 3317 2039
rect 3117 1753 3317 1796
rect 3117 1707 3130 1753
rect 3304 1707 3317 1753
rect 3117 1694 3317 1707
rect 3397 2085 3597 2098
rect 3397 2039 3410 2085
rect 3584 2039 3597 2085
rect 3397 1996 3597 2039
rect 3397 1753 3597 1796
rect 3397 1707 3410 1753
rect 3584 1707 3597 1753
rect 3397 1694 3597 1707
rect 3677 2085 3877 2098
rect 3677 2039 3690 2085
rect 3864 2039 3877 2085
rect 3677 1996 3877 2039
rect 3677 1753 3877 1796
rect 3677 1707 3690 1753
rect 3864 1707 3877 1753
rect 3677 1694 3877 1707
rect 3957 2085 4157 2098
rect 3957 2039 3970 2085
rect 4144 2039 4157 2085
rect 3957 1996 4157 2039
rect 3957 1753 4157 1796
rect 3957 1707 3970 1753
rect 4144 1707 4157 1753
rect 3957 1694 4157 1707
rect 4237 2085 4437 2098
rect 4237 2039 4250 2085
rect 4424 2039 4437 2085
rect 4237 1996 4437 2039
rect 4237 1753 4437 1796
rect 4237 1707 4250 1753
rect 4424 1707 4437 1753
rect 4237 1694 4437 1707
rect 4517 2085 4717 2098
rect 4517 2039 4530 2085
rect 4704 2039 4717 2085
rect 4517 1996 4717 2039
rect 4517 1753 4717 1796
rect 4517 1707 4530 1753
rect 4704 1707 4717 1753
rect 4517 1694 4717 1707
rect 4797 2085 4997 2098
rect 4797 2039 4810 2085
rect 4984 2039 4997 2085
rect 4797 1996 4997 2039
rect 4797 1753 4997 1796
rect 4797 1707 4810 1753
rect 4984 1707 4997 1753
rect 4797 1694 4997 1707
rect 5077 2085 5277 2098
rect 5077 2039 5090 2085
rect 5264 2039 5277 2085
rect 5077 1996 5277 2039
rect 5077 1753 5277 1796
rect 5077 1707 5090 1753
rect 5264 1707 5277 1753
rect 5077 1694 5277 1707
rect 5357 2085 5557 2098
rect 5357 2039 5370 2085
rect 5544 2039 5557 2085
rect 5357 1996 5557 2039
rect 5357 1753 5557 1796
rect 5357 1707 5370 1753
rect 5544 1707 5557 1753
rect 5357 1694 5557 1707
rect 5637 2085 5837 2098
rect 5637 2039 5650 2085
rect 5824 2039 5837 2085
rect 5637 1996 5837 2039
rect 5637 1753 5837 1796
rect 5637 1707 5650 1753
rect 5824 1707 5837 1753
rect 5637 1694 5837 1707
rect 5917 2085 6117 2098
rect 5917 2039 5930 2085
rect 6104 2039 6117 2085
rect 5917 1996 6117 2039
rect 5917 1753 6117 1796
rect 5917 1707 5930 1753
rect 6104 1707 6117 1753
rect 5917 1694 6117 1707
rect 6197 2085 6397 2098
rect 6197 2039 6210 2085
rect 6384 2039 6397 2085
rect 6197 1996 6397 2039
rect 6197 1753 6397 1796
rect 6197 1707 6210 1753
rect 6384 1707 6397 1753
rect 6197 1694 6397 1707
rect 6477 2085 6677 2098
rect 6477 2039 6490 2085
rect 6664 2039 6677 2085
rect 6477 1996 6677 2039
rect 6477 1753 6677 1796
rect 6477 1707 6490 1753
rect 6664 1707 6677 1753
rect 6477 1694 6677 1707
rect 6757 2085 6957 2098
rect 6757 2039 6770 2085
rect 6944 2039 6957 2085
rect 6757 1996 6957 2039
rect 6757 1753 6957 1796
rect 6757 1707 6770 1753
rect 6944 1707 6957 1753
rect 6757 1694 6957 1707
rect 7037 2085 7237 2098
rect 7037 2039 7050 2085
rect 7224 2039 7237 2085
rect 7037 1996 7237 2039
rect 7037 1753 7237 1796
rect 7037 1707 7050 1753
rect 7224 1707 7237 1753
rect 7037 1694 7237 1707
rect 7317 2085 7517 2098
rect 7317 2039 7330 2085
rect 7504 2039 7517 2085
rect 7317 1996 7517 2039
rect 7317 1753 7517 1796
rect 7317 1707 7330 1753
rect 7504 1707 7517 1753
rect 7317 1694 7517 1707
rect 7597 2085 7797 2098
rect 7597 2039 7610 2085
rect 7784 2039 7797 2085
rect 7597 1996 7797 2039
rect 7597 1753 7797 1796
rect 7597 1707 7610 1753
rect 7784 1707 7797 1753
rect 7597 1694 7797 1707
rect 7877 2085 8077 2098
rect 7877 2039 7890 2085
rect 8064 2039 8077 2085
rect 7877 1996 8077 2039
rect 7877 1753 8077 1796
rect 7877 1707 7890 1753
rect 8064 1707 8077 1753
rect 7877 1694 8077 1707
rect 8157 2085 8357 2098
rect 8157 2039 8170 2085
rect 8344 2039 8357 2085
rect 8157 1996 8357 2039
rect 8157 1753 8357 1796
rect 8157 1707 8170 1753
rect 8344 1707 8357 1753
rect 8157 1694 8357 1707
rect 8437 2085 8637 2098
rect 8437 2039 8450 2085
rect 8624 2039 8637 2085
rect 8437 1996 8637 2039
rect 8437 1753 8637 1796
rect 8437 1707 8450 1753
rect 8624 1707 8637 1753
rect 8437 1694 8637 1707
rect 8717 2085 8917 2098
rect 8717 2039 8730 2085
rect 8904 2039 8917 2085
rect 8717 1996 8917 2039
rect 8717 1753 8917 1796
rect 8717 1707 8730 1753
rect 8904 1707 8917 1753
rect 8717 1694 8917 1707
rect 8997 2085 9197 2098
rect 8997 2039 9010 2085
rect 9184 2039 9197 2085
rect 8997 1996 9197 2039
rect 8997 1753 9197 1796
rect 8997 1707 9010 1753
rect 9184 1707 9197 1753
rect 8997 1694 9197 1707
rect 9277 2085 9477 2098
rect 9277 2039 9290 2085
rect 9464 2039 9477 2085
rect 9277 1996 9477 2039
rect 9277 1753 9477 1796
rect 9277 1707 9290 1753
rect 9464 1707 9477 1753
rect 9277 1694 9477 1707
rect 9557 2085 9757 2098
rect 9557 2039 9570 2085
rect 9744 2039 9757 2085
rect 9557 1996 9757 2039
rect 9557 1753 9757 1796
rect 9557 1707 9570 1753
rect 9744 1707 9757 1753
rect 9557 1694 9757 1707
rect 9837 2085 10037 2098
rect 9837 2039 9850 2085
rect 10024 2039 10037 2085
rect 9837 1996 10037 2039
rect 9837 1753 10037 1796
rect 9837 1707 9850 1753
rect 10024 1707 10037 1753
rect 9837 1694 10037 1707
rect 10117 2085 10317 2098
rect 10117 2039 10130 2085
rect 10304 2039 10317 2085
rect 10117 1996 10317 2039
rect 10117 1753 10317 1796
rect 10117 1707 10130 1753
rect 10304 1707 10317 1753
rect 10117 1694 10317 1707
rect 877 1433 1077 1446
rect 877 1387 890 1433
rect 1064 1387 1077 1433
rect 877 1344 1077 1387
rect 877 1101 1077 1144
rect 877 1055 890 1101
rect 1064 1055 1077 1101
rect 877 1042 1077 1055
rect 1157 1433 1357 1446
rect 1157 1387 1170 1433
rect 1344 1387 1357 1433
rect 1157 1344 1357 1387
rect 1157 1101 1357 1144
rect 1157 1055 1170 1101
rect 1344 1055 1357 1101
rect 1157 1042 1357 1055
rect 1437 1433 1637 1446
rect 1437 1387 1450 1433
rect 1624 1387 1637 1433
rect 1437 1344 1637 1387
rect 1437 1101 1637 1144
rect 1437 1055 1450 1101
rect 1624 1055 1637 1101
rect 1437 1042 1637 1055
rect 1717 1433 1917 1446
rect 1717 1387 1730 1433
rect 1904 1387 1917 1433
rect 1717 1344 1917 1387
rect 1717 1101 1917 1144
rect 1717 1055 1730 1101
rect 1904 1055 1917 1101
rect 1717 1042 1917 1055
rect 1997 1433 2197 1446
rect 1997 1387 2010 1433
rect 2184 1387 2197 1433
rect 1997 1344 2197 1387
rect 1997 1101 2197 1144
rect 1997 1055 2010 1101
rect 2184 1055 2197 1101
rect 1997 1042 2197 1055
rect 2277 1433 2477 1446
rect 2277 1387 2290 1433
rect 2464 1387 2477 1433
rect 2277 1344 2477 1387
rect 2277 1101 2477 1144
rect 2277 1055 2290 1101
rect 2464 1055 2477 1101
rect 2277 1042 2477 1055
rect 2557 1433 2757 1446
rect 2557 1387 2570 1433
rect 2744 1387 2757 1433
rect 2557 1344 2757 1387
rect 2557 1101 2757 1144
rect 2557 1055 2570 1101
rect 2744 1055 2757 1101
rect 2557 1042 2757 1055
rect 2837 1433 3037 1446
rect 2837 1387 2850 1433
rect 3024 1387 3037 1433
rect 2837 1344 3037 1387
rect 2837 1101 3037 1144
rect 2837 1055 2850 1101
rect 3024 1055 3037 1101
rect 2837 1042 3037 1055
rect 3117 1433 3317 1446
rect 3117 1387 3130 1433
rect 3304 1387 3317 1433
rect 3117 1344 3317 1387
rect 3117 1101 3317 1144
rect 3117 1055 3130 1101
rect 3304 1055 3317 1101
rect 3117 1042 3317 1055
rect 3397 1433 3597 1446
rect 3397 1387 3410 1433
rect 3584 1387 3597 1433
rect 3397 1344 3597 1387
rect 3397 1101 3597 1144
rect 3397 1055 3410 1101
rect 3584 1055 3597 1101
rect 3397 1042 3597 1055
rect 3677 1433 3877 1446
rect 3677 1387 3690 1433
rect 3864 1387 3877 1433
rect 3677 1344 3877 1387
rect 3677 1101 3877 1144
rect 3677 1055 3690 1101
rect 3864 1055 3877 1101
rect 3677 1042 3877 1055
rect 3957 1433 4157 1446
rect 3957 1387 3970 1433
rect 4144 1387 4157 1433
rect 3957 1344 4157 1387
rect 3957 1101 4157 1144
rect 3957 1055 3970 1101
rect 4144 1055 4157 1101
rect 3957 1042 4157 1055
rect 4237 1433 4437 1446
rect 4237 1387 4250 1433
rect 4424 1387 4437 1433
rect 4237 1344 4437 1387
rect 4237 1101 4437 1144
rect 4237 1055 4250 1101
rect 4424 1055 4437 1101
rect 4237 1042 4437 1055
rect 4517 1433 4717 1446
rect 4517 1387 4530 1433
rect 4704 1387 4717 1433
rect 4517 1344 4717 1387
rect 4517 1101 4717 1144
rect 4517 1055 4530 1101
rect 4704 1055 4717 1101
rect 4517 1042 4717 1055
rect 4797 1433 4997 1446
rect 4797 1387 4810 1433
rect 4984 1387 4997 1433
rect 4797 1344 4997 1387
rect 4797 1101 4997 1144
rect 4797 1055 4810 1101
rect 4984 1055 4997 1101
rect 4797 1042 4997 1055
rect 5077 1433 5277 1446
rect 5077 1387 5090 1433
rect 5264 1387 5277 1433
rect 5077 1344 5277 1387
rect 5077 1101 5277 1144
rect 5077 1055 5090 1101
rect 5264 1055 5277 1101
rect 5077 1042 5277 1055
rect 5357 1433 5557 1446
rect 5357 1387 5370 1433
rect 5544 1387 5557 1433
rect 5357 1344 5557 1387
rect 5357 1101 5557 1144
rect 5357 1055 5370 1101
rect 5544 1055 5557 1101
rect 5357 1042 5557 1055
rect 5637 1433 5837 1446
rect 5637 1387 5650 1433
rect 5824 1387 5837 1433
rect 5637 1344 5837 1387
rect 5637 1101 5837 1144
rect 5637 1055 5650 1101
rect 5824 1055 5837 1101
rect 5637 1042 5837 1055
rect 5917 1433 6117 1446
rect 5917 1387 5930 1433
rect 6104 1387 6117 1433
rect 5917 1344 6117 1387
rect 5917 1101 6117 1144
rect 5917 1055 5930 1101
rect 6104 1055 6117 1101
rect 5917 1042 6117 1055
rect 6197 1433 6397 1446
rect 6197 1387 6210 1433
rect 6384 1387 6397 1433
rect 6197 1344 6397 1387
rect 6197 1101 6397 1144
rect 6197 1055 6210 1101
rect 6384 1055 6397 1101
rect 6197 1042 6397 1055
rect 6477 1433 6677 1446
rect 6477 1387 6490 1433
rect 6664 1387 6677 1433
rect 6477 1344 6677 1387
rect 6477 1101 6677 1144
rect 6477 1055 6490 1101
rect 6664 1055 6677 1101
rect 6477 1042 6677 1055
rect 6757 1433 6957 1446
rect 6757 1387 6770 1433
rect 6944 1387 6957 1433
rect 6757 1344 6957 1387
rect 6757 1101 6957 1144
rect 6757 1055 6770 1101
rect 6944 1055 6957 1101
rect 6757 1042 6957 1055
rect 7037 1433 7237 1446
rect 7037 1387 7050 1433
rect 7224 1387 7237 1433
rect 7037 1344 7237 1387
rect 7037 1101 7237 1144
rect 7037 1055 7050 1101
rect 7224 1055 7237 1101
rect 7037 1042 7237 1055
rect 7317 1433 7517 1446
rect 7317 1387 7330 1433
rect 7504 1387 7517 1433
rect 7317 1344 7517 1387
rect 7317 1101 7517 1144
rect 7317 1055 7330 1101
rect 7504 1055 7517 1101
rect 7317 1042 7517 1055
rect 7597 1433 7797 1446
rect 7597 1387 7610 1433
rect 7784 1387 7797 1433
rect 7597 1344 7797 1387
rect 7597 1101 7797 1144
rect 7597 1055 7610 1101
rect 7784 1055 7797 1101
rect 7597 1042 7797 1055
rect 7877 1433 8077 1446
rect 7877 1387 7890 1433
rect 8064 1387 8077 1433
rect 7877 1344 8077 1387
rect 7877 1101 8077 1144
rect 7877 1055 7890 1101
rect 8064 1055 8077 1101
rect 7877 1042 8077 1055
rect 8157 1433 8357 1446
rect 8157 1387 8170 1433
rect 8344 1387 8357 1433
rect 8157 1344 8357 1387
rect 8157 1101 8357 1144
rect 8157 1055 8170 1101
rect 8344 1055 8357 1101
rect 8157 1042 8357 1055
rect 8437 1433 8637 1446
rect 8437 1387 8450 1433
rect 8624 1387 8637 1433
rect 8437 1344 8637 1387
rect 8437 1101 8637 1144
rect 8437 1055 8450 1101
rect 8624 1055 8637 1101
rect 8437 1042 8637 1055
rect 8717 1433 8917 1446
rect 8717 1387 8730 1433
rect 8904 1387 8917 1433
rect 8717 1344 8917 1387
rect 8717 1101 8917 1144
rect 8717 1055 8730 1101
rect 8904 1055 8917 1101
rect 8717 1042 8917 1055
rect 8997 1433 9197 1446
rect 8997 1387 9010 1433
rect 9184 1387 9197 1433
rect 8997 1344 9197 1387
rect 8997 1101 9197 1144
rect 8997 1055 9010 1101
rect 9184 1055 9197 1101
rect 8997 1042 9197 1055
rect 9277 1433 9477 1446
rect 9277 1387 9290 1433
rect 9464 1387 9477 1433
rect 9277 1344 9477 1387
rect 9277 1101 9477 1144
rect 9277 1055 9290 1101
rect 9464 1055 9477 1101
rect 9277 1042 9477 1055
rect 9557 1433 9757 1446
rect 9557 1387 9570 1433
rect 9744 1387 9757 1433
rect 9557 1344 9757 1387
rect 9557 1101 9757 1144
rect 9557 1055 9570 1101
rect 9744 1055 9757 1101
rect 9557 1042 9757 1055
rect 9837 1433 10037 1446
rect 9837 1387 9850 1433
rect 10024 1387 10037 1433
rect 9837 1344 10037 1387
rect 9837 1101 10037 1144
rect 9837 1055 9850 1101
rect 10024 1055 10037 1101
rect 9837 1042 10037 1055
rect 10117 1433 10317 1446
rect 10117 1387 10130 1433
rect 10304 1387 10317 1433
rect 10117 1344 10317 1387
rect 10117 1101 10317 1144
rect 10117 1055 10130 1101
rect 10304 1055 10317 1101
rect 10117 1042 10317 1055
rect 877 781 1077 794
rect 877 735 890 781
rect 1064 735 1077 781
rect 877 692 1077 735
rect 877 449 1077 492
rect 877 403 890 449
rect 1064 403 1077 449
rect 877 390 1077 403
rect 1157 781 1357 794
rect 1157 735 1170 781
rect 1344 735 1357 781
rect 1157 692 1357 735
rect 1157 449 1357 492
rect 1157 403 1170 449
rect 1344 403 1357 449
rect 1157 390 1357 403
rect 1437 781 1637 794
rect 1437 735 1450 781
rect 1624 735 1637 781
rect 1437 692 1637 735
rect 1437 449 1637 492
rect 1437 403 1450 449
rect 1624 403 1637 449
rect 1437 390 1637 403
rect 1717 781 1917 794
rect 1717 735 1730 781
rect 1904 735 1917 781
rect 1717 692 1917 735
rect 1717 449 1917 492
rect 1717 403 1730 449
rect 1904 403 1917 449
rect 1717 390 1917 403
rect 1997 781 2197 794
rect 1997 735 2010 781
rect 2184 735 2197 781
rect 1997 692 2197 735
rect 1997 449 2197 492
rect 1997 403 2010 449
rect 2184 403 2197 449
rect 1997 390 2197 403
rect 2277 781 2477 794
rect 2277 735 2290 781
rect 2464 735 2477 781
rect 2277 692 2477 735
rect 2277 449 2477 492
rect 2277 403 2290 449
rect 2464 403 2477 449
rect 2277 390 2477 403
rect 2557 781 2757 794
rect 2557 735 2570 781
rect 2744 735 2757 781
rect 2557 692 2757 735
rect 2557 449 2757 492
rect 2557 403 2570 449
rect 2744 403 2757 449
rect 2557 390 2757 403
rect 2837 781 3037 794
rect 2837 735 2850 781
rect 3024 735 3037 781
rect 2837 692 3037 735
rect 2837 449 3037 492
rect 2837 403 2850 449
rect 3024 403 3037 449
rect 2837 390 3037 403
rect 3117 781 3317 794
rect 3117 735 3130 781
rect 3304 735 3317 781
rect 3117 692 3317 735
rect 3117 449 3317 492
rect 3117 403 3130 449
rect 3304 403 3317 449
rect 3117 390 3317 403
rect 3397 781 3597 794
rect 3397 735 3410 781
rect 3584 735 3597 781
rect 3397 692 3597 735
rect 3397 449 3597 492
rect 3397 403 3410 449
rect 3584 403 3597 449
rect 3397 390 3597 403
rect 3677 781 3877 794
rect 3677 735 3690 781
rect 3864 735 3877 781
rect 3677 692 3877 735
rect 3677 449 3877 492
rect 3677 403 3690 449
rect 3864 403 3877 449
rect 3677 390 3877 403
rect 3957 781 4157 794
rect 3957 735 3970 781
rect 4144 735 4157 781
rect 3957 692 4157 735
rect 3957 449 4157 492
rect 3957 403 3970 449
rect 4144 403 4157 449
rect 3957 390 4157 403
rect 4237 781 4437 794
rect 4237 735 4250 781
rect 4424 735 4437 781
rect 4237 692 4437 735
rect 4237 449 4437 492
rect 4237 403 4250 449
rect 4424 403 4437 449
rect 4237 390 4437 403
rect 4517 781 4717 794
rect 4517 735 4530 781
rect 4704 735 4717 781
rect 4517 692 4717 735
rect 4517 449 4717 492
rect 4517 403 4530 449
rect 4704 403 4717 449
rect 4517 390 4717 403
rect 4797 781 4997 794
rect 4797 735 4810 781
rect 4984 735 4997 781
rect 4797 692 4997 735
rect 4797 449 4997 492
rect 4797 403 4810 449
rect 4984 403 4997 449
rect 4797 390 4997 403
rect 5077 781 5277 794
rect 5077 735 5090 781
rect 5264 735 5277 781
rect 5077 692 5277 735
rect 5077 449 5277 492
rect 5077 403 5090 449
rect 5264 403 5277 449
rect 5077 390 5277 403
rect 5357 781 5557 794
rect 5357 735 5370 781
rect 5544 735 5557 781
rect 5357 692 5557 735
rect 5357 449 5557 492
rect 5357 403 5370 449
rect 5544 403 5557 449
rect 5357 390 5557 403
rect 5637 781 5837 794
rect 5637 735 5650 781
rect 5824 735 5837 781
rect 5637 692 5837 735
rect 5637 449 5837 492
rect 5637 403 5650 449
rect 5824 403 5837 449
rect 5637 390 5837 403
rect 5917 781 6117 794
rect 5917 735 5930 781
rect 6104 735 6117 781
rect 5917 692 6117 735
rect 5917 449 6117 492
rect 5917 403 5930 449
rect 6104 403 6117 449
rect 5917 390 6117 403
rect 6197 781 6397 794
rect 6197 735 6210 781
rect 6384 735 6397 781
rect 6197 692 6397 735
rect 6197 449 6397 492
rect 6197 403 6210 449
rect 6384 403 6397 449
rect 6197 390 6397 403
rect 6477 781 6677 794
rect 6477 735 6490 781
rect 6664 735 6677 781
rect 6477 692 6677 735
rect 6477 449 6677 492
rect 6477 403 6490 449
rect 6664 403 6677 449
rect 6477 390 6677 403
rect 6757 781 6957 794
rect 6757 735 6770 781
rect 6944 735 6957 781
rect 6757 692 6957 735
rect 6757 449 6957 492
rect 6757 403 6770 449
rect 6944 403 6957 449
rect 6757 390 6957 403
rect 7037 781 7237 794
rect 7037 735 7050 781
rect 7224 735 7237 781
rect 7037 692 7237 735
rect 7037 449 7237 492
rect 7037 403 7050 449
rect 7224 403 7237 449
rect 7037 390 7237 403
rect 7317 781 7517 794
rect 7317 735 7330 781
rect 7504 735 7517 781
rect 7317 692 7517 735
rect 7317 449 7517 492
rect 7317 403 7330 449
rect 7504 403 7517 449
rect 7317 390 7517 403
rect 7597 781 7797 794
rect 7597 735 7610 781
rect 7784 735 7797 781
rect 7597 692 7797 735
rect 7597 449 7797 492
rect 7597 403 7610 449
rect 7784 403 7797 449
rect 7597 390 7797 403
rect 7877 781 8077 794
rect 7877 735 7890 781
rect 8064 735 8077 781
rect 7877 692 8077 735
rect 7877 449 8077 492
rect 7877 403 7890 449
rect 8064 403 8077 449
rect 7877 390 8077 403
rect 8157 781 8357 794
rect 8157 735 8170 781
rect 8344 735 8357 781
rect 8157 692 8357 735
rect 8157 449 8357 492
rect 8157 403 8170 449
rect 8344 403 8357 449
rect 8157 390 8357 403
rect 8437 781 8637 794
rect 8437 735 8450 781
rect 8624 735 8637 781
rect 8437 692 8637 735
rect 8437 449 8637 492
rect 8437 403 8450 449
rect 8624 403 8637 449
rect 8437 390 8637 403
rect 8717 781 8917 794
rect 8717 735 8730 781
rect 8904 735 8917 781
rect 8717 692 8917 735
rect 8717 449 8917 492
rect 8717 403 8730 449
rect 8904 403 8917 449
rect 8717 390 8917 403
rect 8997 781 9197 794
rect 8997 735 9010 781
rect 9184 735 9197 781
rect 8997 692 9197 735
rect 8997 449 9197 492
rect 8997 403 9010 449
rect 9184 403 9197 449
rect 8997 390 9197 403
rect 9277 781 9477 794
rect 9277 735 9290 781
rect 9464 735 9477 781
rect 9277 692 9477 735
rect 9277 449 9477 492
rect 9277 403 9290 449
rect 9464 403 9477 449
rect 9277 390 9477 403
rect 9557 781 9757 794
rect 9557 735 9570 781
rect 9744 735 9757 781
rect 9557 692 9757 735
rect 9557 449 9757 492
rect 9557 403 9570 449
rect 9744 403 9757 449
rect 9557 390 9757 403
rect 9837 781 10037 794
rect 9837 735 9850 781
rect 10024 735 10037 781
rect 9837 692 10037 735
rect 9837 449 10037 492
rect 9837 403 9850 449
rect 10024 403 10037 449
rect 9837 390 10037 403
rect 10117 781 10317 794
rect 10117 735 10130 781
rect 10304 735 10317 781
rect 10117 692 10317 735
rect 10117 449 10317 492
rect 10117 403 10130 449
rect 10304 403 10317 449
rect 10117 390 10317 403
rect 877 -403 1077 -390
rect 877 -449 890 -403
rect 1064 -449 1077 -403
rect 877 -492 1077 -449
rect 877 -735 1077 -692
rect 877 -781 890 -735
rect 1064 -781 1077 -735
rect 877 -794 1077 -781
rect 1157 -403 1357 -390
rect 1157 -449 1170 -403
rect 1344 -449 1357 -403
rect 1157 -492 1357 -449
rect 1157 -735 1357 -692
rect 1157 -781 1170 -735
rect 1344 -781 1357 -735
rect 1157 -794 1357 -781
rect 1437 -403 1637 -390
rect 1437 -449 1450 -403
rect 1624 -449 1637 -403
rect 1437 -492 1637 -449
rect 1437 -735 1637 -692
rect 1437 -781 1450 -735
rect 1624 -781 1637 -735
rect 1437 -794 1637 -781
rect 1717 -403 1917 -390
rect 1717 -449 1730 -403
rect 1904 -449 1917 -403
rect 1717 -492 1917 -449
rect 1717 -735 1917 -692
rect 1717 -781 1730 -735
rect 1904 -781 1917 -735
rect 1717 -794 1917 -781
rect 1997 -403 2197 -390
rect 1997 -449 2010 -403
rect 2184 -449 2197 -403
rect 1997 -492 2197 -449
rect 1997 -735 2197 -692
rect 1997 -781 2010 -735
rect 2184 -781 2197 -735
rect 1997 -794 2197 -781
rect 2277 -403 2477 -390
rect 2277 -449 2290 -403
rect 2464 -449 2477 -403
rect 2277 -492 2477 -449
rect 2277 -735 2477 -692
rect 2277 -781 2290 -735
rect 2464 -781 2477 -735
rect 2277 -794 2477 -781
rect 2557 -403 2757 -390
rect 2557 -449 2570 -403
rect 2744 -449 2757 -403
rect 2557 -492 2757 -449
rect 2557 -735 2757 -692
rect 2557 -781 2570 -735
rect 2744 -781 2757 -735
rect 2557 -794 2757 -781
rect 2837 -403 3037 -390
rect 2837 -449 2850 -403
rect 3024 -449 3037 -403
rect 2837 -492 3037 -449
rect 2837 -735 3037 -692
rect 2837 -781 2850 -735
rect 3024 -781 3037 -735
rect 2837 -794 3037 -781
rect 3117 -403 3317 -390
rect 3117 -449 3130 -403
rect 3304 -449 3317 -403
rect 3117 -492 3317 -449
rect 3117 -735 3317 -692
rect 3117 -781 3130 -735
rect 3304 -781 3317 -735
rect 3117 -794 3317 -781
rect 3397 -403 3597 -390
rect 3397 -449 3410 -403
rect 3584 -449 3597 -403
rect 3397 -492 3597 -449
rect 3397 -735 3597 -692
rect 3397 -781 3410 -735
rect 3584 -781 3597 -735
rect 3397 -794 3597 -781
rect 3677 -403 3877 -390
rect 3677 -449 3690 -403
rect 3864 -449 3877 -403
rect 3677 -492 3877 -449
rect 3677 -735 3877 -692
rect 3677 -781 3690 -735
rect 3864 -781 3877 -735
rect 3677 -794 3877 -781
rect 3957 -403 4157 -390
rect 3957 -449 3970 -403
rect 4144 -449 4157 -403
rect 3957 -492 4157 -449
rect 3957 -735 4157 -692
rect 3957 -781 3970 -735
rect 4144 -781 4157 -735
rect 3957 -794 4157 -781
rect 4237 -403 4437 -390
rect 4237 -449 4250 -403
rect 4424 -449 4437 -403
rect 4237 -492 4437 -449
rect 4237 -735 4437 -692
rect 4237 -781 4250 -735
rect 4424 -781 4437 -735
rect 4237 -794 4437 -781
rect 4517 -403 4717 -390
rect 4517 -449 4530 -403
rect 4704 -449 4717 -403
rect 4517 -492 4717 -449
rect 4517 -735 4717 -692
rect 4517 -781 4530 -735
rect 4704 -781 4717 -735
rect 4517 -794 4717 -781
rect 4797 -403 4997 -390
rect 4797 -449 4810 -403
rect 4984 -449 4997 -403
rect 4797 -492 4997 -449
rect 4797 -735 4997 -692
rect 4797 -781 4810 -735
rect 4984 -781 4997 -735
rect 4797 -794 4997 -781
rect 5077 -403 5277 -390
rect 5077 -449 5090 -403
rect 5264 -449 5277 -403
rect 5077 -492 5277 -449
rect 5077 -735 5277 -692
rect 5077 -781 5090 -735
rect 5264 -781 5277 -735
rect 5077 -794 5277 -781
rect 5357 -403 5557 -390
rect 5357 -449 5370 -403
rect 5544 -449 5557 -403
rect 5357 -492 5557 -449
rect 5357 -735 5557 -692
rect 5357 -781 5370 -735
rect 5544 -781 5557 -735
rect 5357 -794 5557 -781
rect 5637 -403 5837 -390
rect 5637 -449 5650 -403
rect 5824 -449 5837 -403
rect 5637 -492 5837 -449
rect 5637 -735 5837 -692
rect 5637 -781 5650 -735
rect 5824 -781 5837 -735
rect 5637 -794 5837 -781
rect 5917 -403 6117 -390
rect 5917 -449 5930 -403
rect 6104 -449 6117 -403
rect 5917 -492 6117 -449
rect 5917 -735 6117 -692
rect 5917 -781 5930 -735
rect 6104 -781 6117 -735
rect 5917 -794 6117 -781
rect 6197 -403 6397 -390
rect 6197 -449 6210 -403
rect 6384 -449 6397 -403
rect 6197 -492 6397 -449
rect 6197 -735 6397 -692
rect 6197 -781 6210 -735
rect 6384 -781 6397 -735
rect 6197 -794 6397 -781
rect 6477 -403 6677 -390
rect 6477 -449 6490 -403
rect 6664 -449 6677 -403
rect 6477 -492 6677 -449
rect 6477 -735 6677 -692
rect 6477 -781 6490 -735
rect 6664 -781 6677 -735
rect 6477 -794 6677 -781
rect 6757 -403 6957 -390
rect 6757 -449 6770 -403
rect 6944 -449 6957 -403
rect 6757 -492 6957 -449
rect 6757 -735 6957 -692
rect 6757 -781 6770 -735
rect 6944 -781 6957 -735
rect 6757 -794 6957 -781
rect 7037 -403 7237 -390
rect 7037 -449 7050 -403
rect 7224 -449 7237 -403
rect 7037 -492 7237 -449
rect 7037 -735 7237 -692
rect 7037 -781 7050 -735
rect 7224 -781 7237 -735
rect 7037 -794 7237 -781
rect 7317 -403 7517 -390
rect 7317 -449 7330 -403
rect 7504 -449 7517 -403
rect 7317 -492 7517 -449
rect 7317 -735 7517 -692
rect 7317 -781 7330 -735
rect 7504 -781 7517 -735
rect 7317 -794 7517 -781
rect 7597 -403 7797 -390
rect 7597 -449 7610 -403
rect 7784 -449 7797 -403
rect 7597 -492 7797 -449
rect 7597 -735 7797 -692
rect 7597 -781 7610 -735
rect 7784 -781 7797 -735
rect 7597 -794 7797 -781
rect 7877 -403 8077 -390
rect 7877 -449 7890 -403
rect 8064 -449 8077 -403
rect 7877 -492 8077 -449
rect 7877 -735 8077 -692
rect 7877 -781 7890 -735
rect 8064 -781 8077 -735
rect 7877 -794 8077 -781
rect 8157 -403 8357 -390
rect 8157 -449 8170 -403
rect 8344 -449 8357 -403
rect 8157 -492 8357 -449
rect 8157 -735 8357 -692
rect 8157 -781 8170 -735
rect 8344 -781 8357 -735
rect 8157 -794 8357 -781
rect 8437 -403 8637 -390
rect 8437 -449 8450 -403
rect 8624 -449 8637 -403
rect 8437 -492 8637 -449
rect 8437 -735 8637 -692
rect 8437 -781 8450 -735
rect 8624 -781 8637 -735
rect 8437 -794 8637 -781
rect 8717 -403 8917 -390
rect 8717 -449 8730 -403
rect 8904 -449 8917 -403
rect 8717 -492 8917 -449
rect 8717 -735 8917 -692
rect 8717 -781 8730 -735
rect 8904 -781 8917 -735
rect 8717 -794 8917 -781
rect 8997 -403 9197 -390
rect 8997 -449 9010 -403
rect 9184 -449 9197 -403
rect 8997 -492 9197 -449
rect 8997 -735 9197 -692
rect 8997 -781 9010 -735
rect 9184 -781 9197 -735
rect 8997 -794 9197 -781
rect 9277 -403 9477 -390
rect 9277 -449 9290 -403
rect 9464 -449 9477 -403
rect 9277 -492 9477 -449
rect 9277 -735 9477 -692
rect 9277 -781 9290 -735
rect 9464 -781 9477 -735
rect 9277 -794 9477 -781
rect 9557 -403 9757 -390
rect 9557 -449 9570 -403
rect 9744 -449 9757 -403
rect 9557 -492 9757 -449
rect 9557 -735 9757 -692
rect 9557 -781 9570 -735
rect 9744 -781 9757 -735
rect 9557 -794 9757 -781
rect 9837 -403 10037 -390
rect 9837 -449 9850 -403
rect 10024 -449 10037 -403
rect 9837 -492 10037 -449
rect 9837 -735 10037 -692
rect 9837 -781 9850 -735
rect 10024 -781 10037 -735
rect 9837 -794 10037 -781
rect 10117 -403 10317 -390
rect 10117 -449 10130 -403
rect 10304 -449 10317 -403
rect 10117 -492 10317 -449
rect 10117 -735 10317 -692
rect 10117 -781 10130 -735
rect 10304 -781 10317 -735
rect 10117 -794 10317 -781
rect 877 -1055 1077 -1042
rect 877 -1101 890 -1055
rect 1064 -1101 1077 -1055
rect 877 -1144 1077 -1101
rect 877 -1387 1077 -1344
rect 877 -1433 890 -1387
rect 1064 -1433 1077 -1387
rect 877 -1446 1077 -1433
rect 1157 -1055 1357 -1042
rect 1157 -1101 1170 -1055
rect 1344 -1101 1357 -1055
rect 1157 -1144 1357 -1101
rect 1157 -1387 1357 -1344
rect 1157 -1433 1170 -1387
rect 1344 -1433 1357 -1387
rect 1157 -1446 1357 -1433
rect 1437 -1055 1637 -1042
rect 1437 -1101 1450 -1055
rect 1624 -1101 1637 -1055
rect 1437 -1144 1637 -1101
rect 1437 -1387 1637 -1344
rect 1437 -1433 1450 -1387
rect 1624 -1433 1637 -1387
rect 1437 -1446 1637 -1433
rect 1717 -1055 1917 -1042
rect 1717 -1101 1730 -1055
rect 1904 -1101 1917 -1055
rect 1717 -1144 1917 -1101
rect 1717 -1387 1917 -1344
rect 1717 -1433 1730 -1387
rect 1904 -1433 1917 -1387
rect 1717 -1446 1917 -1433
rect 1997 -1055 2197 -1042
rect 1997 -1101 2010 -1055
rect 2184 -1101 2197 -1055
rect 1997 -1144 2197 -1101
rect 1997 -1387 2197 -1344
rect 1997 -1433 2010 -1387
rect 2184 -1433 2197 -1387
rect 1997 -1446 2197 -1433
rect 2277 -1055 2477 -1042
rect 2277 -1101 2290 -1055
rect 2464 -1101 2477 -1055
rect 2277 -1144 2477 -1101
rect 2277 -1387 2477 -1344
rect 2277 -1433 2290 -1387
rect 2464 -1433 2477 -1387
rect 2277 -1446 2477 -1433
rect 2557 -1055 2757 -1042
rect 2557 -1101 2570 -1055
rect 2744 -1101 2757 -1055
rect 2557 -1144 2757 -1101
rect 2557 -1387 2757 -1344
rect 2557 -1433 2570 -1387
rect 2744 -1433 2757 -1387
rect 2557 -1446 2757 -1433
rect 2837 -1055 3037 -1042
rect 2837 -1101 2850 -1055
rect 3024 -1101 3037 -1055
rect 2837 -1144 3037 -1101
rect 2837 -1387 3037 -1344
rect 2837 -1433 2850 -1387
rect 3024 -1433 3037 -1387
rect 2837 -1446 3037 -1433
rect 3117 -1055 3317 -1042
rect 3117 -1101 3130 -1055
rect 3304 -1101 3317 -1055
rect 3117 -1144 3317 -1101
rect 3117 -1387 3317 -1344
rect 3117 -1433 3130 -1387
rect 3304 -1433 3317 -1387
rect 3117 -1446 3317 -1433
rect 3397 -1055 3597 -1042
rect 3397 -1101 3410 -1055
rect 3584 -1101 3597 -1055
rect 3397 -1144 3597 -1101
rect 3397 -1387 3597 -1344
rect 3397 -1433 3410 -1387
rect 3584 -1433 3597 -1387
rect 3397 -1446 3597 -1433
rect 3677 -1055 3877 -1042
rect 3677 -1101 3690 -1055
rect 3864 -1101 3877 -1055
rect 3677 -1144 3877 -1101
rect 3677 -1387 3877 -1344
rect 3677 -1433 3690 -1387
rect 3864 -1433 3877 -1387
rect 3677 -1446 3877 -1433
rect 3957 -1055 4157 -1042
rect 3957 -1101 3970 -1055
rect 4144 -1101 4157 -1055
rect 3957 -1144 4157 -1101
rect 3957 -1387 4157 -1344
rect 3957 -1433 3970 -1387
rect 4144 -1433 4157 -1387
rect 3957 -1446 4157 -1433
rect 4237 -1055 4437 -1042
rect 4237 -1101 4250 -1055
rect 4424 -1101 4437 -1055
rect 4237 -1144 4437 -1101
rect 4237 -1387 4437 -1344
rect 4237 -1433 4250 -1387
rect 4424 -1433 4437 -1387
rect 4237 -1446 4437 -1433
rect 4517 -1055 4717 -1042
rect 4517 -1101 4530 -1055
rect 4704 -1101 4717 -1055
rect 4517 -1144 4717 -1101
rect 4517 -1387 4717 -1344
rect 4517 -1433 4530 -1387
rect 4704 -1433 4717 -1387
rect 4517 -1446 4717 -1433
rect 4797 -1055 4997 -1042
rect 4797 -1101 4810 -1055
rect 4984 -1101 4997 -1055
rect 4797 -1144 4997 -1101
rect 4797 -1387 4997 -1344
rect 4797 -1433 4810 -1387
rect 4984 -1433 4997 -1387
rect 4797 -1446 4997 -1433
rect 5077 -1055 5277 -1042
rect 5077 -1101 5090 -1055
rect 5264 -1101 5277 -1055
rect 5077 -1144 5277 -1101
rect 5077 -1387 5277 -1344
rect 5077 -1433 5090 -1387
rect 5264 -1433 5277 -1387
rect 5077 -1446 5277 -1433
rect 5357 -1055 5557 -1042
rect 5357 -1101 5370 -1055
rect 5544 -1101 5557 -1055
rect 5357 -1144 5557 -1101
rect 5357 -1387 5557 -1344
rect 5357 -1433 5370 -1387
rect 5544 -1433 5557 -1387
rect 5357 -1446 5557 -1433
rect 5637 -1055 5837 -1042
rect 5637 -1101 5650 -1055
rect 5824 -1101 5837 -1055
rect 5637 -1144 5837 -1101
rect 5637 -1387 5837 -1344
rect 5637 -1433 5650 -1387
rect 5824 -1433 5837 -1387
rect 5637 -1446 5837 -1433
rect 5917 -1055 6117 -1042
rect 5917 -1101 5930 -1055
rect 6104 -1101 6117 -1055
rect 5917 -1144 6117 -1101
rect 5917 -1387 6117 -1344
rect 5917 -1433 5930 -1387
rect 6104 -1433 6117 -1387
rect 5917 -1446 6117 -1433
rect 6197 -1055 6397 -1042
rect 6197 -1101 6210 -1055
rect 6384 -1101 6397 -1055
rect 6197 -1144 6397 -1101
rect 6197 -1387 6397 -1344
rect 6197 -1433 6210 -1387
rect 6384 -1433 6397 -1387
rect 6197 -1446 6397 -1433
rect 6477 -1055 6677 -1042
rect 6477 -1101 6490 -1055
rect 6664 -1101 6677 -1055
rect 6477 -1144 6677 -1101
rect 6477 -1387 6677 -1344
rect 6477 -1433 6490 -1387
rect 6664 -1433 6677 -1387
rect 6477 -1446 6677 -1433
rect 6757 -1055 6957 -1042
rect 6757 -1101 6770 -1055
rect 6944 -1101 6957 -1055
rect 6757 -1144 6957 -1101
rect 6757 -1387 6957 -1344
rect 6757 -1433 6770 -1387
rect 6944 -1433 6957 -1387
rect 6757 -1446 6957 -1433
rect 7037 -1055 7237 -1042
rect 7037 -1101 7050 -1055
rect 7224 -1101 7237 -1055
rect 7037 -1144 7237 -1101
rect 7037 -1387 7237 -1344
rect 7037 -1433 7050 -1387
rect 7224 -1433 7237 -1387
rect 7037 -1446 7237 -1433
rect 7317 -1055 7517 -1042
rect 7317 -1101 7330 -1055
rect 7504 -1101 7517 -1055
rect 7317 -1144 7517 -1101
rect 7317 -1387 7517 -1344
rect 7317 -1433 7330 -1387
rect 7504 -1433 7517 -1387
rect 7317 -1446 7517 -1433
rect 7597 -1055 7797 -1042
rect 7597 -1101 7610 -1055
rect 7784 -1101 7797 -1055
rect 7597 -1144 7797 -1101
rect 7597 -1387 7797 -1344
rect 7597 -1433 7610 -1387
rect 7784 -1433 7797 -1387
rect 7597 -1446 7797 -1433
rect 7877 -1055 8077 -1042
rect 7877 -1101 7890 -1055
rect 8064 -1101 8077 -1055
rect 7877 -1144 8077 -1101
rect 7877 -1387 8077 -1344
rect 7877 -1433 7890 -1387
rect 8064 -1433 8077 -1387
rect 7877 -1446 8077 -1433
rect 8157 -1055 8357 -1042
rect 8157 -1101 8170 -1055
rect 8344 -1101 8357 -1055
rect 8157 -1144 8357 -1101
rect 8157 -1387 8357 -1344
rect 8157 -1433 8170 -1387
rect 8344 -1433 8357 -1387
rect 8157 -1446 8357 -1433
rect 8437 -1055 8637 -1042
rect 8437 -1101 8450 -1055
rect 8624 -1101 8637 -1055
rect 8437 -1144 8637 -1101
rect 8437 -1387 8637 -1344
rect 8437 -1433 8450 -1387
rect 8624 -1433 8637 -1387
rect 8437 -1446 8637 -1433
rect 8717 -1055 8917 -1042
rect 8717 -1101 8730 -1055
rect 8904 -1101 8917 -1055
rect 8717 -1144 8917 -1101
rect 8717 -1387 8917 -1344
rect 8717 -1433 8730 -1387
rect 8904 -1433 8917 -1387
rect 8717 -1446 8917 -1433
rect 8997 -1055 9197 -1042
rect 8997 -1101 9010 -1055
rect 9184 -1101 9197 -1055
rect 8997 -1144 9197 -1101
rect 8997 -1387 9197 -1344
rect 8997 -1433 9010 -1387
rect 9184 -1433 9197 -1387
rect 8997 -1446 9197 -1433
rect 9277 -1055 9477 -1042
rect 9277 -1101 9290 -1055
rect 9464 -1101 9477 -1055
rect 9277 -1144 9477 -1101
rect 9277 -1387 9477 -1344
rect 9277 -1433 9290 -1387
rect 9464 -1433 9477 -1387
rect 9277 -1446 9477 -1433
rect 9557 -1055 9757 -1042
rect 9557 -1101 9570 -1055
rect 9744 -1101 9757 -1055
rect 9557 -1144 9757 -1101
rect 9557 -1387 9757 -1344
rect 9557 -1433 9570 -1387
rect 9744 -1433 9757 -1387
rect 9557 -1446 9757 -1433
rect 9837 -1055 10037 -1042
rect 9837 -1101 9850 -1055
rect 10024 -1101 10037 -1055
rect 9837 -1144 10037 -1101
rect 9837 -1387 10037 -1344
rect 9837 -1433 9850 -1387
rect 10024 -1433 10037 -1387
rect 9837 -1446 10037 -1433
rect 10117 -1055 10317 -1042
rect 10117 -1101 10130 -1055
rect 10304 -1101 10317 -1055
rect 10117 -1144 10317 -1101
rect 10117 -1387 10317 -1344
rect 10117 -1433 10130 -1387
rect 10304 -1433 10317 -1387
rect 10117 -1446 10317 -1433
rect 877 -1707 1077 -1694
rect 877 -1753 890 -1707
rect 1064 -1753 1077 -1707
rect 877 -1796 1077 -1753
rect 877 -2039 1077 -1996
rect 877 -2085 890 -2039
rect 1064 -2085 1077 -2039
rect 877 -2098 1077 -2085
rect 1157 -1707 1357 -1694
rect 1157 -1753 1170 -1707
rect 1344 -1753 1357 -1707
rect 1157 -1796 1357 -1753
rect 1157 -2039 1357 -1996
rect 1157 -2085 1170 -2039
rect 1344 -2085 1357 -2039
rect 1157 -2098 1357 -2085
rect 1437 -1707 1637 -1694
rect 1437 -1753 1450 -1707
rect 1624 -1753 1637 -1707
rect 1437 -1796 1637 -1753
rect 1437 -2039 1637 -1996
rect 1437 -2085 1450 -2039
rect 1624 -2085 1637 -2039
rect 1437 -2098 1637 -2085
rect 1717 -1707 1917 -1694
rect 1717 -1753 1730 -1707
rect 1904 -1753 1917 -1707
rect 1717 -1796 1917 -1753
rect 1717 -2039 1917 -1996
rect 1717 -2085 1730 -2039
rect 1904 -2085 1917 -2039
rect 1717 -2098 1917 -2085
rect 1997 -1707 2197 -1694
rect 1997 -1753 2010 -1707
rect 2184 -1753 2197 -1707
rect 1997 -1796 2197 -1753
rect 1997 -2039 2197 -1996
rect 1997 -2085 2010 -2039
rect 2184 -2085 2197 -2039
rect 1997 -2098 2197 -2085
rect 2277 -1707 2477 -1694
rect 2277 -1753 2290 -1707
rect 2464 -1753 2477 -1707
rect 2277 -1796 2477 -1753
rect 2277 -2039 2477 -1996
rect 2277 -2085 2290 -2039
rect 2464 -2085 2477 -2039
rect 2277 -2098 2477 -2085
rect 2557 -1707 2757 -1694
rect 2557 -1753 2570 -1707
rect 2744 -1753 2757 -1707
rect 2557 -1796 2757 -1753
rect 2557 -2039 2757 -1996
rect 2557 -2085 2570 -2039
rect 2744 -2085 2757 -2039
rect 2557 -2098 2757 -2085
rect 2837 -1707 3037 -1694
rect 2837 -1753 2850 -1707
rect 3024 -1753 3037 -1707
rect 2837 -1796 3037 -1753
rect 2837 -2039 3037 -1996
rect 2837 -2085 2850 -2039
rect 3024 -2085 3037 -2039
rect 2837 -2098 3037 -2085
rect 3117 -1707 3317 -1694
rect 3117 -1753 3130 -1707
rect 3304 -1753 3317 -1707
rect 3117 -1796 3317 -1753
rect 3117 -2039 3317 -1996
rect 3117 -2085 3130 -2039
rect 3304 -2085 3317 -2039
rect 3117 -2098 3317 -2085
rect 3397 -1707 3597 -1694
rect 3397 -1753 3410 -1707
rect 3584 -1753 3597 -1707
rect 3397 -1796 3597 -1753
rect 3397 -2039 3597 -1996
rect 3397 -2085 3410 -2039
rect 3584 -2085 3597 -2039
rect 3397 -2098 3597 -2085
rect 3677 -1707 3877 -1694
rect 3677 -1753 3690 -1707
rect 3864 -1753 3877 -1707
rect 3677 -1796 3877 -1753
rect 3677 -2039 3877 -1996
rect 3677 -2085 3690 -2039
rect 3864 -2085 3877 -2039
rect 3677 -2098 3877 -2085
rect 3957 -1707 4157 -1694
rect 3957 -1753 3970 -1707
rect 4144 -1753 4157 -1707
rect 3957 -1796 4157 -1753
rect 3957 -2039 4157 -1996
rect 3957 -2085 3970 -2039
rect 4144 -2085 4157 -2039
rect 3957 -2098 4157 -2085
rect 4237 -1707 4437 -1694
rect 4237 -1753 4250 -1707
rect 4424 -1753 4437 -1707
rect 4237 -1796 4437 -1753
rect 4237 -2039 4437 -1996
rect 4237 -2085 4250 -2039
rect 4424 -2085 4437 -2039
rect 4237 -2098 4437 -2085
rect 4517 -1707 4717 -1694
rect 4517 -1753 4530 -1707
rect 4704 -1753 4717 -1707
rect 4517 -1796 4717 -1753
rect 4517 -2039 4717 -1996
rect 4517 -2085 4530 -2039
rect 4704 -2085 4717 -2039
rect 4517 -2098 4717 -2085
rect 4797 -1707 4997 -1694
rect 4797 -1753 4810 -1707
rect 4984 -1753 4997 -1707
rect 4797 -1796 4997 -1753
rect 4797 -2039 4997 -1996
rect 4797 -2085 4810 -2039
rect 4984 -2085 4997 -2039
rect 4797 -2098 4997 -2085
rect 5077 -1707 5277 -1694
rect 5077 -1753 5090 -1707
rect 5264 -1753 5277 -1707
rect 5077 -1796 5277 -1753
rect 5077 -2039 5277 -1996
rect 5077 -2085 5090 -2039
rect 5264 -2085 5277 -2039
rect 5077 -2098 5277 -2085
rect 5357 -1707 5557 -1694
rect 5357 -1753 5370 -1707
rect 5544 -1753 5557 -1707
rect 5357 -1796 5557 -1753
rect 5357 -2039 5557 -1996
rect 5357 -2085 5370 -2039
rect 5544 -2085 5557 -2039
rect 5357 -2098 5557 -2085
rect 5637 -1707 5837 -1694
rect 5637 -1753 5650 -1707
rect 5824 -1753 5837 -1707
rect 5637 -1796 5837 -1753
rect 5637 -2039 5837 -1996
rect 5637 -2085 5650 -2039
rect 5824 -2085 5837 -2039
rect 5637 -2098 5837 -2085
rect 5917 -1707 6117 -1694
rect 5917 -1753 5930 -1707
rect 6104 -1753 6117 -1707
rect 5917 -1796 6117 -1753
rect 5917 -2039 6117 -1996
rect 5917 -2085 5930 -2039
rect 6104 -2085 6117 -2039
rect 5917 -2098 6117 -2085
rect 6197 -1707 6397 -1694
rect 6197 -1753 6210 -1707
rect 6384 -1753 6397 -1707
rect 6197 -1796 6397 -1753
rect 6197 -2039 6397 -1996
rect 6197 -2085 6210 -2039
rect 6384 -2085 6397 -2039
rect 6197 -2098 6397 -2085
rect 6477 -1707 6677 -1694
rect 6477 -1753 6490 -1707
rect 6664 -1753 6677 -1707
rect 6477 -1796 6677 -1753
rect 6477 -2039 6677 -1996
rect 6477 -2085 6490 -2039
rect 6664 -2085 6677 -2039
rect 6477 -2098 6677 -2085
rect 6757 -1707 6957 -1694
rect 6757 -1753 6770 -1707
rect 6944 -1753 6957 -1707
rect 6757 -1796 6957 -1753
rect 6757 -2039 6957 -1996
rect 6757 -2085 6770 -2039
rect 6944 -2085 6957 -2039
rect 6757 -2098 6957 -2085
rect 7037 -1707 7237 -1694
rect 7037 -1753 7050 -1707
rect 7224 -1753 7237 -1707
rect 7037 -1796 7237 -1753
rect 7037 -2039 7237 -1996
rect 7037 -2085 7050 -2039
rect 7224 -2085 7237 -2039
rect 7037 -2098 7237 -2085
rect 7317 -1707 7517 -1694
rect 7317 -1753 7330 -1707
rect 7504 -1753 7517 -1707
rect 7317 -1796 7517 -1753
rect 7317 -2039 7517 -1996
rect 7317 -2085 7330 -2039
rect 7504 -2085 7517 -2039
rect 7317 -2098 7517 -2085
rect 7597 -1707 7797 -1694
rect 7597 -1753 7610 -1707
rect 7784 -1753 7797 -1707
rect 7597 -1796 7797 -1753
rect 7597 -2039 7797 -1996
rect 7597 -2085 7610 -2039
rect 7784 -2085 7797 -2039
rect 7597 -2098 7797 -2085
rect 7877 -1707 8077 -1694
rect 7877 -1753 7890 -1707
rect 8064 -1753 8077 -1707
rect 7877 -1796 8077 -1753
rect 7877 -2039 8077 -1996
rect 7877 -2085 7890 -2039
rect 8064 -2085 8077 -2039
rect 7877 -2098 8077 -2085
rect 8157 -1707 8357 -1694
rect 8157 -1753 8170 -1707
rect 8344 -1753 8357 -1707
rect 8157 -1796 8357 -1753
rect 8157 -2039 8357 -1996
rect 8157 -2085 8170 -2039
rect 8344 -2085 8357 -2039
rect 8157 -2098 8357 -2085
rect 8437 -1707 8637 -1694
rect 8437 -1753 8450 -1707
rect 8624 -1753 8637 -1707
rect 8437 -1796 8637 -1753
rect 8437 -2039 8637 -1996
rect 8437 -2085 8450 -2039
rect 8624 -2085 8637 -2039
rect 8437 -2098 8637 -2085
rect 8717 -1707 8917 -1694
rect 8717 -1753 8730 -1707
rect 8904 -1753 8917 -1707
rect 8717 -1796 8917 -1753
rect 8717 -2039 8917 -1996
rect 8717 -2085 8730 -2039
rect 8904 -2085 8917 -2039
rect 8717 -2098 8917 -2085
rect 8997 -1707 9197 -1694
rect 8997 -1753 9010 -1707
rect 9184 -1753 9197 -1707
rect 8997 -1796 9197 -1753
rect 8997 -2039 9197 -1996
rect 8997 -2085 9010 -2039
rect 9184 -2085 9197 -2039
rect 8997 -2098 9197 -2085
rect 9277 -1707 9477 -1694
rect 9277 -1753 9290 -1707
rect 9464 -1753 9477 -1707
rect 9277 -1796 9477 -1753
rect 9277 -2039 9477 -1996
rect 9277 -2085 9290 -2039
rect 9464 -2085 9477 -2039
rect 9277 -2098 9477 -2085
rect 9557 -1707 9757 -1694
rect 9557 -1753 9570 -1707
rect 9744 -1753 9757 -1707
rect 9557 -1796 9757 -1753
rect 9557 -2039 9757 -1996
rect 9557 -2085 9570 -2039
rect 9744 -2085 9757 -2039
rect 9557 -2098 9757 -2085
rect 9837 -1707 10037 -1694
rect 9837 -1753 9850 -1707
rect 10024 -1753 10037 -1707
rect 9837 -1796 10037 -1753
rect 9837 -2039 10037 -1996
rect 9837 -2085 9850 -2039
rect 10024 -2085 10037 -2039
rect 9837 -2098 10037 -2085
rect 10117 -1707 10317 -1694
rect 10117 -1753 10130 -1707
rect 10304 -1753 10317 -1707
rect 10117 -1796 10317 -1753
rect 10117 -2039 10317 -1996
rect 10117 -2085 10130 -2039
rect 10304 -2085 10317 -2039
rect 10117 -2098 10317 -2085
<< polycontact >>
rect 890 2039 1064 2085
rect 890 1707 1064 1753
rect 1170 2039 1344 2085
rect 1170 1707 1344 1753
rect 1450 2039 1624 2085
rect 1450 1707 1624 1753
rect 1730 2039 1904 2085
rect 1730 1707 1904 1753
rect 2010 2039 2184 2085
rect 2010 1707 2184 1753
rect 2290 2039 2464 2085
rect 2290 1707 2464 1753
rect 2570 2039 2744 2085
rect 2570 1707 2744 1753
rect 2850 2039 3024 2085
rect 2850 1707 3024 1753
rect 3130 2039 3304 2085
rect 3130 1707 3304 1753
rect 3410 2039 3584 2085
rect 3410 1707 3584 1753
rect 3690 2039 3864 2085
rect 3690 1707 3864 1753
rect 3970 2039 4144 2085
rect 3970 1707 4144 1753
rect 4250 2039 4424 2085
rect 4250 1707 4424 1753
rect 4530 2039 4704 2085
rect 4530 1707 4704 1753
rect 4810 2039 4984 2085
rect 4810 1707 4984 1753
rect 5090 2039 5264 2085
rect 5090 1707 5264 1753
rect 5370 2039 5544 2085
rect 5370 1707 5544 1753
rect 5650 2039 5824 2085
rect 5650 1707 5824 1753
rect 5930 2039 6104 2085
rect 5930 1707 6104 1753
rect 6210 2039 6384 2085
rect 6210 1707 6384 1753
rect 6490 2039 6664 2085
rect 6490 1707 6664 1753
rect 6770 2039 6944 2085
rect 6770 1707 6944 1753
rect 7050 2039 7224 2085
rect 7050 1707 7224 1753
rect 7330 2039 7504 2085
rect 7330 1707 7504 1753
rect 7610 2039 7784 2085
rect 7610 1707 7784 1753
rect 7890 2039 8064 2085
rect 7890 1707 8064 1753
rect 8170 2039 8344 2085
rect 8170 1707 8344 1753
rect 8450 2039 8624 2085
rect 8450 1707 8624 1753
rect 8730 2039 8904 2085
rect 8730 1707 8904 1753
rect 9010 2039 9184 2085
rect 9010 1707 9184 1753
rect 9290 2039 9464 2085
rect 9290 1707 9464 1753
rect 9570 2039 9744 2085
rect 9570 1707 9744 1753
rect 9850 2039 10024 2085
rect 9850 1707 10024 1753
rect 10130 2039 10304 2085
rect 10130 1707 10304 1753
rect 890 1387 1064 1433
rect 890 1055 1064 1101
rect 1170 1387 1344 1433
rect 1170 1055 1344 1101
rect 1450 1387 1624 1433
rect 1450 1055 1624 1101
rect 1730 1387 1904 1433
rect 1730 1055 1904 1101
rect 2010 1387 2184 1433
rect 2010 1055 2184 1101
rect 2290 1387 2464 1433
rect 2290 1055 2464 1101
rect 2570 1387 2744 1433
rect 2570 1055 2744 1101
rect 2850 1387 3024 1433
rect 2850 1055 3024 1101
rect 3130 1387 3304 1433
rect 3130 1055 3304 1101
rect 3410 1387 3584 1433
rect 3410 1055 3584 1101
rect 3690 1387 3864 1433
rect 3690 1055 3864 1101
rect 3970 1387 4144 1433
rect 3970 1055 4144 1101
rect 4250 1387 4424 1433
rect 4250 1055 4424 1101
rect 4530 1387 4704 1433
rect 4530 1055 4704 1101
rect 4810 1387 4984 1433
rect 4810 1055 4984 1101
rect 5090 1387 5264 1433
rect 5090 1055 5264 1101
rect 5370 1387 5544 1433
rect 5370 1055 5544 1101
rect 5650 1387 5824 1433
rect 5650 1055 5824 1101
rect 5930 1387 6104 1433
rect 5930 1055 6104 1101
rect 6210 1387 6384 1433
rect 6210 1055 6384 1101
rect 6490 1387 6664 1433
rect 6490 1055 6664 1101
rect 6770 1387 6944 1433
rect 6770 1055 6944 1101
rect 7050 1387 7224 1433
rect 7050 1055 7224 1101
rect 7330 1387 7504 1433
rect 7330 1055 7504 1101
rect 7610 1387 7784 1433
rect 7610 1055 7784 1101
rect 7890 1387 8064 1433
rect 7890 1055 8064 1101
rect 8170 1387 8344 1433
rect 8170 1055 8344 1101
rect 8450 1387 8624 1433
rect 8450 1055 8624 1101
rect 8730 1387 8904 1433
rect 8730 1055 8904 1101
rect 9010 1387 9184 1433
rect 9010 1055 9184 1101
rect 9290 1387 9464 1433
rect 9290 1055 9464 1101
rect 9570 1387 9744 1433
rect 9570 1055 9744 1101
rect 9850 1387 10024 1433
rect 9850 1055 10024 1101
rect 10130 1387 10304 1433
rect 10130 1055 10304 1101
rect 890 735 1064 781
rect 890 403 1064 449
rect 1170 735 1344 781
rect 1170 403 1344 449
rect 1450 735 1624 781
rect 1450 403 1624 449
rect 1730 735 1904 781
rect 1730 403 1904 449
rect 2010 735 2184 781
rect 2010 403 2184 449
rect 2290 735 2464 781
rect 2290 403 2464 449
rect 2570 735 2744 781
rect 2570 403 2744 449
rect 2850 735 3024 781
rect 2850 403 3024 449
rect 3130 735 3304 781
rect 3130 403 3304 449
rect 3410 735 3584 781
rect 3410 403 3584 449
rect 3690 735 3864 781
rect 3690 403 3864 449
rect 3970 735 4144 781
rect 3970 403 4144 449
rect 4250 735 4424 781
rect 4250 403 4424 449
rect 4530 735 4704 781
rect 4530 403 4704 449
rect 4810 735 4984 781
rect 4810 403 4984 449
rect 5090 735 5264 781
rect 5090 403 5264 449
rect 5370 735 5544 781
rect 5370 403 5544 449
rect 5650 735 5824 781
rect 5650 403 5824 449
rect 5930 735 6104 781
rect 5930 403 6104 449
rect 6210 735 6384 781
rect 6210 403 6384 449
rect 6490 735 6664 781
rect 6490 403 6664 449
rect 6770 735 6944 781
rect 6770 403 6944 449
rect 7050 735 7224 781
rect 7050 403 7224 449
rect 7330 735 7504 781
rect 7330 403 7504 449
rect 7610 735 7784 781
rect 7610 403 7784 449
rect 7890 735 8064 781
rect 7890 403 8064 449
rect 8170 735 8344 781
rect 8170 403 8344 449
rect 8450 735 8624 781
rect 8450 403 8624 449
rect 8730 735 8904 781
rect 8730 403 8904 449
rect 9010 735 9184 781
rect 9010 403 9184 449
rect 9290 735 9464 781
rect 9290 403 9464 449
rect 9570 735 9744 781
rect 9570 403 9744 449
rect 9850 735 10024 781
rect 9850 403 10024 449
rect 10130 735 10304 781
rect 10130 403 10304 449
rect 890 -449 1064 -403
rect 890 -781 1064 -735
rect 1170 -449 1344 -403
rect 1170 -781 1344 -735
rect 1450 -449 1624 -403
rect 1450 -781 1624 -735
rect 1730 -449 1904 -403
rect 1730 -781 1904 -735
rect 2010 -449 2184 -403
rect 2010 -781 2184 -735
rect 2290 -449 2464 -403
rect 2290 -781 2464 -735
rect 2570 -449 2744 -403
rect 2570 -781 2744 -735
rect 2850 -449 3024 -403
rect 2850 -781 3024 -735
rect 3130 -449 3304 -403
rect 3130 -781 3304 -735
rect 3410 -449 3584 -403
rect 3410 -781 3584 -735
rect 3690 -449 3864 -403
rect 3690 -781 3864 -735
rect 3970 -449 4144 -403
rect 3970 -781 4144 -735
rect 4250 -449 4424 -403
rect 4250 -781 4424 -735
rect 4530 -449 4704 -403
rect 4530 -781 4704 -735
rect 4810 -449 4984 -403
rect 4810 -781 4984 -735
rect 5090 -449 5264 -403
rect 5090 -781 5264 -735
rect 5370 -449 5544 -403
rect 5370 -781 5544 -735
rect 5650 -449 5824 -403
rect 5650 -781 5824 -735
rect 5930 -449 6104 -403
rect 5930 -781 6104 -735
rect 6210 -449 6384 -403
rect 6210 -781 6384 -735
rect 6490 -449 6664 -403
rect 6490 -781 6664 -735
rect 6770 -449 6944 -403
rect 6770 -781 6944 -735
rect 7050 -449 7224 -403
rect 7050 -781 7224 -735
rect 7330 -449 7504 -403
rect 7330 -781 7504 -735
rect 7610 -449 7784 -403
rect 7610 -781 7784 -735
rect 7890 -449 8064 -403
rect 7890 -781 8064 -735
rect 8170 -449 8344 -403
rect 8170 -781 8344 -735
rect 8450 -449 8624 -403
rect 8450 -781 8624 -735
rect 8730 -449 8904 -403
rect 8730 -781 8904 -735
rect 9010 -449 9184 -403
rect 9010 -781 9184 -735
rect 9290 -449 9464 -403
rect 9290 -781 9464 -735
rect 9570 -449 9744 -403
rect 9570 -781 9744 -735
rect 9850 -449 10024 -403
rect 9850 -781 10024 -735
rect 10130 -449 10304 -403
rect 10130 -781 10304 -735
rect 890 -1101 1064 -1055
rect 890 -1433 1064 -1387
rect 1170 -1101 1344 -1055
rect 1170 -1433 1344 -1387
rect 1450 -1101 1624 -1055
rect 1450 -1433 1624 -1387
rect 1730 -1101 1904 -1055
rect 1730 -1433 1904 -1387
rect 2010 -1101 2184 -1055
rect 2010 -1433 2184 -1387
rect 2290 -1101 2464 -1055
rect 2290 -1433 2464 -1387
rect 2570 -1101 2744 -1055
rect 2570 -1433 2744 -1387
rect 2850 -1101 3024 -1055
rect 2850 -1433 3024 -1387
rect 3130 -1101 3304 -1055
rect 3130 -1433 3304 -1387
rect 3410 -1101 3584 -1055
rect 3410 -1433 3584 -1387
rect 3690 -1101 3864 -1055
rect 3690 -1433 3864 -1387
rect 3970 -1101 4144 -1055
rect 3970 -1433 4144 -1387
rect 4250 -1101 4424 -1055
rect 4250 -1433 4424 -1387
rect 4530 -1101 4704 -1055
rect 4530 -1433 4704 -1387
rect 4810 -1101 4984 -1055
rect 4810 -1433 4984 -1387
rect 5090 -1101 5264 -1055
rect 5090 -1433 5264 -1387
rect 5370 -1101 5544 -1055
rect 5370 -1433 5544 -1387
rect 5650 -1101 5824 -1055
rect 5650 -1433 5824 -1387
rect 5930 -1101 6104 -1055
rect 5930 -1433 6104 -1387
rect 6210 -1101 6384 -1055
rect 6210 -1433 6384 -1387
rect 6490 -1101 6664 -1055
rect 6490 -1433 6664 -1387
rect 6770 -1101 6944 -1055
rect 6770 -1433 6944 -1387
rect 7050 -1101 7224 -1055
rect 7050 -1433 7224 -1387
rect 7330 -1101 7504 -1055
rect 7330 -1433 7504 -1387
rect 7610 -1101 7784 -1055
rect 7610 -1433 7784 -1387
rect 7890 -1101 8064 -1055
rect 7890 -1433 8064 -1387
rect 8170 -1101 8344 -1055
rect 8170 -1433 8344 -1387
rect 8450 -1101 8624 -1055
rect 8450 -1433 8624 -1387
rect 8730 -1101 8904 -1055
rect 8730 -1433 8904 -1387
rect 9010 -1101 9184 -1055
rect 9010 -1433 9184 -1387
rect 9290 -1101 9464 -1055
rect 9290 -1433 9464 -1387
rect 9570 -1101 9744 -1055
rect 9570 -1433 9744 -1387
rect 9850 -1101 10024 -1055
rect 9850 -1433 10024 -1387
rect 10130 -1101 10304 -1055
rect 10130 -1433 10304 -1387
rect 890 -1753 1064 -1707
rect 890 -2085 1064 -2039
rect 1170 -1753 1344 -1707
rect 1170 -2085 1344 -2039
rect 1450 -1753 1624 -1707
rect 1450 -2085 1624 -2039
rect 1730 -1753 1904 -1707
rect 1730 -2085 1904 -2039
rect 2010 -1753 2184 -1707
rect 2010 -2085 2184 -2039
rect 2290 -1753 2464 -1707
rect 2290 -2085 2464 -2039
rect 2570 -1753 2744 -1707
rect 2570 -2085 2744 -2039
rect 2850 -1753 3024 -1707
rect 2850 -2085 3024 -2039
rect 3130 -1753 3304 -1707
rect 3130 -2085 3304 -2039
rect 3410 -1753 3584 -1707
rect 3410 -2085 3584 -2039
rect 3690 -1753 3864 -1707
rect 3690 -2085 3864 -2039
rect 3970 -1753 4144 -1707
rect 3970 -2085 4144 -2039
rect 4250 -1753 4424 -1707
rect 4250 -2085 4424 -2039
rect 4530 -1753 4704 -1707
rect 4530 -2085 4704 -2039
rect 4810 -1753 4984 -1707
rect 4810 -2085 4984 -2039
rect 5090 -1753 5264 -1707
rect 5090 -2085 5264 -2039
rect 5370 -1753 5544 -1707
rect 5370 -2085 5544 -2039
rect 5650 -1753 5824 -1707
rect 5650 -2085 5824 -2039
rect 5930 -1753 6104 -1707
rect 5930 -2085 6104 -2039
rect 6210 -1753 6384 -1707
rect 6210 -2085 6384 -2039
rect 6490 -1753 6664 -1707
rect 6490 -2085 6664 -2039
rect 6770 -1753 6944 -1707
rect 6770 -2085 6944 -2039
rect 7050 -1753 7224 -1707
rect 7050 -2085 7224 -2039
rect 7330 -1753 7504 -1707
rect 7330 -2085 7504 -2039
rect 7610 -1753 7784 -1707
rect 7610 -2085 7784 -2039
rect 7890 -1753 8064 -1707
rect 7890 -2085 8064 -2039
rect 8170 -1753 8344 -1707
rect 8170 -2085 8344 -2039
rect 8450 -1753 8624 -1707
rect 8450 -2085 8624 -2039
rect 8730 -1753 8904 -1707
rect 8730 -2085 8904 -2039
rect 9010 -1753 9184 -1707
rect 9010 -2085 9184 -2039
rect 9290 -1753 9464 -1707
rect 9290 -2085 9464 -2039
rect 9570 -1753 9744 -1707
rect 9570 -2085 9744 -2039
rect 9850 -1753 10024 -1707
rect 9850 -2085 10024 -2039
rect 10130 -1753 10304 -1707
rect 10130 -2085 10304 -2039
<< ppolyres >>
rect 877 1796 1077 1996
rect 1157 1796 1357 1996
rect 1437 1796 1637 1996
rect 1717 1796 1917 1996
rect 1997 1796 2197 1996
rect 2277 1796 2477 1996
rect 2557 1796 2757 1996
rect 2837 1796 3037 1996
rect 3117 1796 3317 1996
rect 3397 1796 3597 1996
rect 3677 1796 3877 1996
rect 3957 1796 4157 1996
rect 4237 1796 4437 1996
rect 4517 1796 4717 1996
rect 4797 1796 4997 1996
rect 5077 1796 5277 1996
rect 5357 1796 5557 1996
rect 5637 1796 5837 1996
rect 5917 1796 6117 1996
rect 6197 1796 6397 1996
rect 6477 1796 6677 1996
rect 6757 1796 6957 1996
rect 7037 1796 7237 1996
rect 7317 1796 7517 1996
rect 7597 1796 7797 1996
rect 7877 1796 8077 1996
rect 8157 1796 8357 1996
rect 8437 1796 8637 1996
rect 8717 1796 8917 1996
rect 8997 1796 9197 1996
rect 9277 1796 9477 1996
rect 9557 1796 9757 1996
rect 9837 1796 10037 1996
rect 10117 1796 10317 1996
rect 877 1144 1077 1344
rect 1157 1144 1357 1344
rect 1437 1144 1637 1344
rect 1717 1144 1917 1344
rect 1997 1144 2197 1344
rect 2277 1144 2477 1344
rect 2557 1144 2757 1344
rect 2837 1144 3037 1344
rect 3117 1144 3317 1344
rect 3397 1144 3597 1344
rect 3677 1144 3877 1344
rect 3957 1144 4157 1344
rect 4237 1144 4437 1344
rect 4517 1144 4717 1344
rect 4797 1144 4997 1344
rect 5077 1144 5277 1344
rect 5357 1144 5557 1344
rect 5637 1144 5837 1344
rect 5917 1144 6117 1344
rect 6197 1144 6397 1344
rect 6477 1144 6677 1344
rect 6757 1144 6957 1344
rect 7037 1144 7237 1344
rect 7317 1144 7517 1344
rect 7597 1144 7797 1344
rect 7877 1144 8077 1344
rect 8157 1144 8357 1344
rect 8437 1144 8637 1344
rect 8717 1144 8917 1344
rect 8997 1144 9197 1344
rect 9277 1144 9477 1344
rect 9557 1144 9757 1344
rect 9837 1144 10037 1344
rect 10117 1144 10317 1344
rect 877 492 1077 692
rect 1157 492 1357 692
rect 1437 492 1637 692
rect 1717 492 1917 692
rect 1997 492 2197 692
rect 2277 492 2477 692
rect 2557 492 2757 692
rect 2837 492 3037 692
rect 3117 492 3317 692
rect 3397 492 3597 692
rect 3677 492 3877 692
rect 3957 492 4157 692
rect 4237 492 4437 692
rect 4517 492 4717 692
rect 4797 492 4997 692
rect 5077 492 5277 692
rect 5357 492 5557 692
rect 5637 492 5837 692
rect 5917 492 6117 692
rect 6197 492 6397 692
rect 6477 492 6677 692
rect 6757 492 6957 692
rect 7037 492 7237 692
rect 7317 492 7517 692
rect 7597 492 7797 692
rect 7877 492 8077 692
rect 8157 492 8357 692
rect 8437 492 8637 692
rect 8717 492 8917 692
rect 8997 492 9197 692
rect 9277 492 9477 692
rect 9557 492 9757 692
rect 9837 492 10037 692
rect 10117 492 10317 692
rect 877 -692 1077 -492
rect 1157 -692 1357 -492
rect 1437 -692 1637 -492
rect 1717 -692 1917 -492
rect 1997 -692 2197 -492
rect 2277 -692 2477 -492
rect 2557 -692 2757 -492
rect 2837 -692 3037 -492
rect 3117 -692 3317 -492
rect 3397 -692 3597 -492
rect 3677 -692 3877 -492
rect 3957 -692 4157 -492
rect 4237 -692 4437 -492
rect 4517 -692 4717 -492
rect 4797 -692 4997 -492
rect 5077 -692 5277 -492
rect 5357 -692 5557 -492
rect 5637 -692 5837 -492
rect 5917 -692 6117 -492
rect 6197 -692 6397 -492
rect 6477 -692 6677 -492
rect 6757 -692 6957 -492
rect 7037 -692 7237 -492
rect 7317 -692 7517 -492
rect 7597 -692 7797 -492
rect 7877 -692 8077 -492
rect 8157 -692 8357 -492
rect 8437 -692 8637 -492
rect 8717 -692 8917 -492
rect 8997 -692 9197 -492
rect 9277 -692 9477 -492
rect 9557 -692 9757 -492
rect 9837 -692 10037 -492
rect 10117 -692 10317 -492
rect 877 -1344 1077 -1144
rect 1157 -1344 1357 -1144
rect 1437 -1344 1637 -1144
rect 1717 -1344 1917 -1144
rect 1997 -1344 2197 -1144
rect 2277 -1344 2477 -1144
rect 2557 -1344 2757 -1144
rect 2837 -1344 3037 -1144
rect 3117 -1344 3317 -1144
rect 3397 -1344 3597 -1144
rect 3677 -1344 3877 -1144
rect 3957 -1344 4157 -1144
rect 4237 -1344 4437 -1144
rect 4517 -1344 4717 -1144
rect 4797 -1344 4997 -1144
rect 5077 -1344 5277 -1144
rect 5357 -1344 5557 -1144
rect 5637 -1344 5837 -1144
rect 5917 -1344 6117 -1144
rect 6197 -1344 6397 -1144
rect 6477 -1344 6677 -1144
rect 6757 -1344 6957 -1144
rect 7037 -1344 7237 -1144
rect 7317 -1344 7517 -1144
rect 7597 -1344 7797 -1144
rect 7877 -1344 8077 -1144
rect 8157 -1344 8357 -1144
rect 8437 -1344 8637 -1144
rect 8717 -1344 8917 -1144
rect 8997 -1344 9197 -1144
rect 9277 -1344 9477 -1144
rect 9557 -1344 9757 -1144
rect 9837 -1344 10037 -1144
rect 10117 -1344 10317 -1144
rect 877 -1996 1077 -1796
rect 1157 -1996 1357 -1796
rect 1437 -1996 1637 -1796
rect 1717 -1996 1917 -1796
rect 1997 -1996 2197 -1796
rect 2277 -1996 2477 -1796
rect 2557 -1996 2757 -1796
rect 2837 -1996 3037 -1796
rect 3117 -1996 3317 -1796
rect 3397 -1996 3597 -1796
rect 3677 -1996 3877 -1796
rect 3957 -1996 4157 -1796
rect 4237 -1996 4437 -1796
rect 4517 -1996 4717 -1796
rect 4797 -1996 4997 -1796
rect 5077 -1996 5277 -1796
rect 5357 -1996 5557 -1796
rect 5637 -1996 5837 -1796
rect 5917 -1996 6117 -1796
rect 6197 -1996 6397 -1796
rect 6477 -1996 6677 -1796
rect 6757 -1996 6957 -1796
rect 7037 -1996 7237 -1796
rect 7317 -1996 7517 -1796
rect 7597 -1996 7797 -1796
rect 7877 -1996 8077 -1796
rect 8157 -1996 8357 -1796
rect 8437 -1996 8637 -1796
rect 8717 -1996 8917 -1796
rect 8997 -1996 9197 -1796
rect 9277 -1996 9477 -1796
rect 9557 -1996 9757 -1796
rect 9837 -1996 10037 -1796
rect 10117 -1996 10317 -1796
<< metal1 >>
rect 543 2377 10651 2394
rect 543 2327 560 2377
rect 606 2331 658 2377
rect 704 2331 756 2377
rect 802 2331 854 2377
rect 900 2331 952 2377
rect 998 2331 1050 2377
rect 1096 2331 1148 2377
rect 1194 2331 1246 2377
rect 1292 2331 1344 2377
rect 1390 2331 1442 2377
rect 1488 2331 1540 2377
rect 1586 2331 1638 2377
rect 1684 2331 1736 2377
rect 1782 2331 1834 2377
rect 1880 2331 1932 2377
rect 1978 2331 2030 2377
rect 2076 2331 2128 2377
rect 2174 2331 2226 2377
rect 2272 2331 2324 2377
rect 2370 2331 2422 2377
rect 2468 2331 2520 2377
rect 2566 2331 2618 2377
rect 2664 2331 2716 2377
rect 2762 2331 2814 2377
rect 2860 2331 2912 2377
rect 2958 2331 3010 2377
rect 3056 2331 3108 2377
rect 3154 2331 3206 2377
rect 3252 2331 3304 2377
rect 3350 2331 3402 2377
rect 3448 2331 3500 2377
rect 3546 2331 3598 2377
rect 3644 2331 3696 2377
rect 3742 2331 3794 2377
rect 3840 2331 3892 2377
rect 3938 2331 3990 2377
rect 4036 2331 4088 2377
rect 4134 2331 4186 2377
rect 4232 2331 4284 2377
rect 4330 2331 4382 2377
rect 4428 2331 4480 2377
rect 4526 2331 4578 2377
rect 4624 2331 4676 2377
rect 4722 2331 4774 2377
rect 4820 2331 4872 2377
rect 4918 2331 4970 2377
rect 5016 2331 5068 2377
rect 5114 2331 5166 2377
rect 5212 2331 5264 2377
rect 5310 2331 5362 2377
rect 5408 2331 5460 2377
rect 5506 2331 5558 2377
rect 5604 2331 5656 2377
rect 5702 2331 5754 2377
rect 5800 2331 5852 2377
rect 5898 2331 5950 2377
rect 5996 2331 6048 2377
rect 6094 2331 6146 2377
rect 6192 2331 6244 2377
rect 6290 2331 6342 2377
rect 6388 2331 6440 2377
rect 6486 2331 6538 2377
rect 6584 2331 6636 2377
rect 6682 2331 6734 2377
rect 6780 2331 6832 2377
rect 6878 2331 6930 2377
rect 6976 2331 7028 2377
rect 7074 2331 7126 2377
rect 7172 2331 7224 2377
rect 7270 2331 7322 2377
rect 7368 2331 7420 2377
rect 7466 2331 7518 2377
rect 7564 2331 7616 2377
rect 7662 2331 7714 2377
rect 7760 2331 7812 2377
rect 7858 2331 7910 2377
rect 7956 2331 8008 2377
rect 8054 2331 8106 2377
rect 8152 2331 8204 2377
rect 8250 2331 8302 2377
rect 8348 2331 8400 2377
rect 8446 2331 8498 2377
rect 8544 2331 8596 2377
rect 8642 2331 8694 2377
rect 8740 2331 8792 2377
rect 8838 2331 8890 2377
rect 8936 2331 8988 2377
rect 9034 2331 9086 2377
rect 9132 2331 9184 2377
rect 9230 2331 9282 2377
rect 9328 2331 9380 2377
rect 9426 2331 9478 2377
rect 9524 2331 9576 2377
rect 9622 2331 9674 2377
rect 9720 2331 9772 2377
rect 9818 2331 9870 2377
rect 9916 2331 9968 2377
rect 10014 2331 10066 2377
rect 10112 2331 10164 2377
rect 10210 2331 10262 2377
rect 10308 2331 10360 2377
rect 10406 2331 10458 2377
rect 10504 2331 10588 2377
rect 606 2327 10588 2331
rect 10634 2327 10651 2377
rect 543 2314 10651 2327
rect 543 2275 623 2314
rect 543 2229 560 2275
rect 606 2229 623 2275
rect 543 2177 623 2229
rect 543 2131 560 2177
rect 606 2131 623 2177
rect 543 2079 623 2131
rect 951 2085 1020 2314
rect 10571 2275 10651 2314
rect 10571 2229 10588 2275
rect 10634 2229 10651 2275
rect 3036 2191 3226 2195
rect 3036 2182 3048 2191
rect 2138 2136 3048 2182
rect 2138 2085 2184 2136
rect 3036 2135 3048 2136
rect 3104 2135 3158 2191
rect 3214 2135 3226 2191
rect 3036 2131 3226 2135
rect 3488 2191 3678 2195
rect 3488 2135 3500 2191
rect 3556 2135 3610 2191
rect 3666 2182 3678 2191
rect 7516 2191 7706 2195
rect 7516 2182 7528 2191
rect 3666 2136 4576 2182
rect 3666 2135 3678 2136
rect 3488 2131 3678 2135
rect 2277 2085 2477 2089
rect 2634 2085 2684 2087
rect 4030 2085 4080 2087
rect 4237 2085 4437 2089
rect 4530 2085 4576 2136
rect 6618 2136 7528 2182
rect 6618 2085 6664 2136
rect 7516 2135 7528 2136
rect 7584 2135 7638 2191
rect 7694 2135 7706 2191
rect 7516 2131 7706 2135
rect 7968 2191 8158 2195
rect 7968 2135 7980 2191
rect 8036 2135 8090 2191
rect 8146 2182 8158 2191
rect 8146 2136 9056 2182
rect 8146 2135 8158 2136
rect 7968 2131 8158 2135
rect 6757 2085 6957 2089
rect 7114 2085 7164 2087
rect 8510 2085 8560 2087
rect 8717 2085 8917 2089
rect 9010 2085 9056 2136
rect 10571 2177 10651 2229
rect 10571 2131 10588 2177
rect 10634 2131 10651 2177
rect 10571 2091 10651 2131
rect 10302 2085 10651 2091
rect 543 2033 560 2079
rect 606 2033 623 2079
rect 879 2039 890 2085
rect 1064 2039 1075 2085
rect 1159 2039 1170 2085
rect 1344 2039 1450 2085
rect 1624 2039 1646 2085
rect 1719 2039 1730 2085
rect 1904 2039 1915 2085
rect 1999 2039 2010 2085
rect 2184 2039 2195 2085
rect 2277 2039 2290 2085
rect 2464 2039 2477 2085
rect 2559 2039 2570 2085
rect 2744 2039 2755 2085
rect 2839 2039 2850 2085
rect 3024 2039 3130 2085
rect 3304 2039 3315 2085
rect 3399 2039 3410 2085
rect 3584 2039 3690 2085
rect 3864 2039 3875 2085
rect 3959 2039 3970 2085
rect 4144 2039 4155 2085
rect 4237 2039 4250 2085
rect 4424 2039 4437 2085
rect 4519 2039 4530 2085
rect 4704 2039 4715 2085
rect 4799 2039 4810 2085
rect 4984 2039 4995 2085
rect 5068 2039 5090 2085
rect 5264 2039 5370 2085
rect 5544 2039 5555 2085
rect 5639 2039 5650 2085
rect 5824 2039 5930 2085
rect 6104 2039 6126 2085
rect 6199 2039 6210 2085
rect 6384 2039 6395 2085
rect 6479 2039 6490 2085
rect 6664 2039 6675 2085
rect 6757 2039 6770 2085
rect 6944 2039 6957 2085
rect 7039 2039 7050 2085
rect 7224 2039 7235 2085
rect 7319 2039 7330 2085
rect 7504 2039 7610 2085
rect 7784 2039 7795 2085
rect 7879 2039 7890 2085
rect 8064 2039 8170 2085
rect 8344 2039 8355 2085
rect 8439 2039 8450 2085
rect 8624 2039 8635 2085
rect 8717 2039 8730 2085
rect 8904 2039 8917 2085
rect 8999 2039 9010 2085
rect 9184 2039 9195 2085
rect 9279 2039 9290 2085
rect 9464 2039 9475 2085
rect 9548 2039 9570 2085
rect 9744 2039 9850 2085
rect 10024 2039 10035 2085
rect 10119 2039 10130 2085
rect 10304 2079 10651 2085
rect 10304 2039 10588 2079
rect 543 1981 623 2033
rect 543 1935 560 1981
rect 606 1935 623 1981
rect 543 1883 623 1935
rect 543 1837 560 1883
rect 606 1837 623 1883
rect 543 1785 623 1837
rect 543 1739 560 1785
rect 606 1739 623 1785
rect 951 1753 1020 2039
rect 1170 1753 1251 2039
rect 1774 1887 1831 2039
rect 2277 2024 2291 2039
rect 2347 2024 2401 2039
rect 2457 2024 2477 2039
rect 2277 2012 2477 2024
rect 2634 1983 2684 2039
rect 4030 1983 4080 2039
rect 4237 2024 4257 2039
rect 4313 2024 4367 2039
rect 4423 2024 4437 2039
rect 4237 2012 4437 2024
rect 2634 1933 4080 1983
rect 4883 1887 4940 2039
rect 1774 1830 4940 1887
rect 6254 1887 6311 2039
rect 6757 2024 6771 2039
rect 6827 2024 6881 2039
rect 6937 2024 6957 2039
rect 6757 2012 6957 2024
rect 7114 1983 7164 2039
rect 8510 1983 8560 2039
rect 8717 2024 8737 2039
rect 8793 2024 8847 2039
rect 8903 2024 8917 2039
rect 8717 2012 8917 2024
rect 7114 1933 8560 1983
rect 9363 1887 9420 2039
rect 10302 2034 10588 2039
rect 6254 1830 9420 1887
rect 10571 2033 10588 2034
rect 10634 2033 10651 2079
rect 10571 1981 10651 2033
rect 10571 1935 10588 1981
rect 10634 1935 10651 1981
rect 10571 1883 10651 1935
rect 10571 1837 10588 1883
rect 10634 1837 10651 1883
rect 10571 1785 10651 1837
rect 1437 1765 1637 1779
rect 543 1687 623 1739
rect 879 1707 890 1753
rect 1064 1707 1075 1753
rect 1159 1707 1170 1753
rect 1344 1707 1355 1753
rect 1437 1709 1449 1765
rect 1505 1753 1557 1765
rect 1613 1753 1637 1765
rect 1997 1772 2197 1780
rect 1437 1707 1450 1709
rect 1624 1707 1637 1753
rect 1719 1707 1730 1753
rect 1904 1707 1915 1753
rect 1997 1707 2010 1772
rect 2066 1753 2120 1772
rect 2176 1753 2197 1772
rect 2184 1707 2197 1753
rect 543 1641 560 1687
rect 606 1641 623 1687
rect 543 1589 623 1641
rect 543 1543 560 1589
rect 606 1543 623 1589
rect 915 1646 1112 1651
rect 915 1590 931 1646
rect 987 1590 1041 1646
rect 1097 1641 1112 1646
rect 1170 1641 1216 1707
rect 1437 1702 1637 1707
rect 1097 1595 1216 1641
rect 1097 1590 1112 1595
rect 915 1585 1112 1590
rect 543 1491 623 1543
rect 346 1431 412 1446
rect 346 1375 351 1431
rect 407 1375 412 1431
rect 346 1321 412 1375
rect 346 1265 351 1321
rect 407 1265 412 1321
rect 346 1249 412 1265
rect 543 1445 560 1491
rect 606 1445 623 1491
rect 543 1442 623 1445
rect 1296 1579 1611 1583
rect 1296 1523 1433 1579
rect 1489 1523 1543 1579
rect 1599 1523 1611 1579
rect 1296 1517 1611 1523
rect 1737 1536 1783 1707
rect 1997 1703 2197 1707
rect 2277 1769 2477 1780
rect 2277 1753 2291 1769
rect 2347 1753 2401 1769
rect 2457 1753 2477 1769
rect 2837 1766 3037 1780
rect 2277 1707 2290 1753
rect 2464 1707 2477 1753
rect 2559 1707 2570 1753
rect 2744 1707 2755 1753
rect 2837 1710 2849 1766
rect 2905 1753 2959 1766
rect 3015 1753 3037 1766
rect 3677 1766 3877 1780
rect 3677 1753 3699 1766
rect 3755 1753 3809 1766
rect 2837 1707 2850 1710
rect 3024 1707 3037 1753
rect 3119 1707 3130 1753
rect 3304 1707 3410 1753
rect 3584 1707 3595 1753
rect 3677 1707 3690 1753
rect 3865 1710 3877 1766
rect 4237 1769 4437 1780
rect 4237 1753 4257 1769
rect 4313 1753 4367 1769
rect 4423 1753 4437 1769
rect 3864 1707 3877 1710
rect 3959 1707 3970 1753
rect 4144 1707 4155 1753
rect 4237 1707 4250 1753
rect 4424 1707 4437 1753
rect 2277 1703 2477 1707
rect 1832 1645 2024 1647
rect 2570 1645 2620 1707
rect 2837 1703 3037 1707
rect 3677 1703 3877 1707
rect 1832 1644 2620 1645
rect 1832 1588 1844 1644
rect 1900 1588 1954 1644
rect 2010 1599 2620 1644
rect 4094 1645 4144 1707
rect 4237 1703 4437 1707
rect 4517 1772 4717 1780
rect 4517 1753 4538 1772
rect 4594 1753 4648 1772
rect 4517 1707 4530 1753
rect 4704 1707 4717 1772
rect 5077 1765 5277 1779
rect 5077 1753 5101 1765
rect 5157 1753 5209 1765
rect 4799 1707 4810 1753
rect 4984 1707 4995 1753
rect 5077 1707 5090 1753
rect 5265 1709 5277 1765
rect 5917 1765 6117 1779
rect 5264 1707 5277 1709
rect 5359 1707 5370 1753
rect 5544 1707 5555 1753
rect 5639 1707 5650 1753
rect 5824 1707 5835 1753
rect 5917 1709 5929 1765
rect 5985 1753 6037 1765
rect 6093 1753 6117 1765
rect 6477 1772 6677 1780
rect 5917 1707 5930 1709
rect 6104 1707 6117 1753
rect 6199 1707 6210 1753
rect 6384 1707 6395 1753
rect 6477 1707 6490 1772
rect 6546 1753 6600 1772
rect 6656 1753 6677 1772
rect 6664 1707 6677 1753
rect 4517 1703 4717 1707
rect 4690 1645 4882 1647
rect 4094 1644 4882 1645
rect 4094 1599 4704 1644
rect 2010 1588 2024 1599
rect 1832 1585 2024 1588
rect 4690 1588 4704 1599
rect 4760 1588 4814 1644
rect 4870 1588 4882 1644
rect 4690 1585 4882 1588
rect 4931 1536 4977 1707
rect 5077 1702 5277 1707
rect 5498 1661 5544 1707
rect 5650 1661 5696 1707
rect 5917 1702 6117 1707
rect 5466 1615 5696 1661
rect 543 1433 930 1442
rect 1296 1433 1344 1517
rect 1737 1490 2620 1536
rect 1437 1433 1637 1435
rect 543 1393 890 1433
rect 543 1347 560 1393
rect 606 1387 890 1393
rect 1064 1387 1075 1433
rect 1159 1387 1170 1433
rect 1344 1387 1355 1433
rect 1437 1387 1450 1433
rect 1624 1387 1637 1433
rect 606 1376 930 1387
rect 606 1347 623 1376
rect 1437 1367 1452 1387
rect 1508 1367 1562 1387
rect 1618 1367 1637 1387
rect 1437 1357 1637 1367
rect 1717 1433 1917 1437
rect 2073 1433 2123 1434
rect 2357 1433 2407 1434
rect 2570 1433 2620 1490
rect 4094 1490 4977 1536
rect 5101 1578 5418 1583
rect 5101 1522 5113 1578
rect 5169 1522 5223 1578
rect 5279 1522 5418 1578
rect 5101 1517 5418 1522
rect 2837 1433 3037 1436
rect 1717 1387 1730 1433
rect 1904 1387 1917 1433
rect 1999 1387 2010 1433
rect 2184 1387 2195 1433
rect 2279 1387 2290 1433
rect 2464 1387 2475 1433
rect 2559 1387 2570 1433
rect 2744 1387 2755 1433
rect 2837 1387 2850 1433
rect 3024 1387 3037 1433
rect 1717 1373 1732 1387
rect 1788 1373 1842 1387
rect 1898 1373 1917 1387
rect 1717 1360 1917 1373
rect 543 1295 623 1347
rect 543 1249 560 1295
rect 606 1249 623 1295
rect 678 1311 875 1315
rect 2073 1311 2123 1387
rect 678 1310 2123 1311
rect 678 1254 691 1310
rect 747 1254 801 1310
rect 857 1261 2123 1310
rect 2357 1309 2407 1387
rect 2837 1366 2851 1387
rect 2907 1366 2961 1387
rect 3017 1366 3037 1387
rect 2837 1356 3037 1366
rect 3117 1433 3317 1437
rect 3117 1368 3130 1433
rect 3304 1387 3317 1433
rect 3186 1368 3240 1387
rect 3296 1368 3317 1387
rect 3117 1360 3317 1368
rect 3397 1433 3597 1437
rect 3397 1387 3410 1433
rect 3397 1368 3418 1387
rect 3474 1368 3528 1387
rect 3584 1368 3597 1433
rect 3397 1360 3597 1368
rect 3677 1433 3877 1436
rect 4094 1433 4144 1490
rect 4307 1433 4357 1434
rect 4591 1433 4641 1434
rect 4797 1433 4997 1437
rect 3677 1387 3690 1433
rect 3864 1387 3877 1433
rect 3959 1387 3970 1433
rect 4144 1387 4155 1433
rect 4239 1387 4250 1433
rect 4424 1387 4435 1433
rect 4519 1387 4530 1433
rect 4704 1387 4715 1433
rect 4797 1387 4810 1433
rect 4984 1387 4997 1433
rect 3677 1366 3697 1387
rect 3753 1366 3807 1387
rect 3863 1366 3877 1387
rect 3677 1356 3877 1366
rect 4307 1309 4357 1387
rect 857 1254 875 1261
rect 2357 1259 4357 1309
rect 4591 1311 4641 1387
rect 4797 1373 4816 1387
rect 4872 1373 4926 1387
rect 4982 1373 4997 1387
rect 4797 1360 4997 1373
rect 5077 1433 5277 1435
rect 5370 1433 5418 1517
rect 5776 1579 6091 1583
rect 5776 1523 5913 1579
rect 5969 1523 6023 1579
rect 6079 1523 6091 1579
rect 5776 1517 6091 1523
rect 6217 1536 6263 1707
rect 6477 1703 6677 1707
rect 6757 1769 6957 1780
rect 6757 1753 6771 1769
rect 6827 1753 6881 1769
rect 6937 1753 6957 1769
rect 7317 1766 7517 1780
rect 6757 1707 6770 1753
rect 6944 1707 6957 1753
rect 7039 1707 7050 1753
rect 7224 1707 7235 1753
rect 7317 1710 7329 1766
rect 7385 1753 7439 1766
rect 7495 1753 7517 1766
rect 8157 1766 8357 1780
rect 8157 1753 8179 1766
rect 8235 1753 8289 1766
rect 7317 1707 7330 1710
rect 7504 1707 7517 1753
rect 7599 1707 7610 1753
rect 7784 1707 7890 1753
rect 8064 1707 8075 1753
rect 8157 1707 8170 1753
rect 8345 1710 8357 1766
rect 8717 1769 8917 1780
rect 8717 1753 8737 1769
rect 8793 1753 8847 1769
rect 8903 1753 8917 1769
rect 8344 1707 8357 1710
rect 8439 1707 8450 1753
rect 8624 1707 8635 1753
rect 8717 1707 8730 1753
rect 8904 1707 8917 1753
rect 6757 1703 6957 1707
rect 6312 1645 6504 1647
rect 7050 1645 7100 1707
rect 7317 1703 7517 1707
rect 8157 1703 8357 1707
rect 6312 1644 7100 1645
rect 6312 1588 6324 1644
rect 6380 1588 6434 1644
rect 6490 1599 7100 1644
rect 8574 1645 8624 1707
rect 8717 1703 8917 1707
rect 8997 1772 9197 1780
rect 8997 1753 9018 1772
rect 9074 1753 9128 1772
rect 8997 1707 9010 1753
rect 9184 1707 9197 1772
rect 9557 1765 9757 1779
rect 10571 1765 10588 1785
rect 9557 1753 9581 1765
rect 9637 1753 9689 1765
rect 9279 1707 9290 1753
rect 9464 1707 9475 1753
rect 9557 1707 9570 1753
rect 9745 1709 9757 1765
rect 10302 1753 10588 1765
rect 9744 1707 9757 1709
rect 9839 1707 9850 1753
rect 10024 1707 10035 1753
rect 10119 1707 10130 1753
rect 10304 1739 10588 1753
rect 10634 1739 10651 1785
rect 10304 1708 10651 1739
rect 10304 1707 10315 1708
rect 8997 1703 9197 1707
rect 9170 1645 9362 1647
rect 8574 1644 9362 1645
rect 8574 1599 9184 1644
rect 6490 1588 6504 1599
rect 6312 1585 6504 1588
rect 9170 1588 9184 1599
rect 9240 1588 9294 1644
rect 9350 1588 9362 1644
rect 9170 1585 9362 1588
rect 9411 1536 9457 1707
rect 9557 1702 9757 1707
rect 9978 1641 10024 1707
rect 10571 1687 10651 1708
rect 10282 1646 10479 1651
rect 10282 1641 10295 1646
rect 9978 1595 10295 1641
rect 10282 1590 10295 1595
rect 10353 1590 10405 1646
rect 10463 1590 10479 1646
rect 10282 1585 10479 1590
rect 10571 1641 10588 1687
rect 10634 1641 10651 1687
rect 10571 1589 10651 1641
rect 5776 1433 5824 1517
rect 6217 1490 7100 1536
rect 5917 1433 6117 1435
rect 5077 1387 5090 1433
rect 5264 1387 5277 1433
rect 5359 1387 5370 1433
rect 5544 1387 5555 1433
rect 5639 1387 5650 1433
rect 5824 1387 5835 1433
rect 5917 1387 5930 1433
rect 6104 1387 6117 1433
rect 5077 1367 5096 1387
rect 5152 1367 5206 1387
rect 5262 1367 5277 1387
rect 5077 1357 5277 1367
rect 5917 1367 5932 1387
rect 5988 1367 6042 1387
rect 6098 1367 6117 1387
rect 5917 1357 6117 1367
rect 6197 1433 6397 1437
rect 6553 1433 6603 1434
rect 6837 1433 6887 1434
rect 7050 1433 7100 1490
rect 8574 1490 9457 1536
rect 9581 1578 9898 1583
rect 9581 1522 9593 1578
rect 9649 1522 9703 1578
rect 9759 1522 9898 1578
rect 9581 1517 9898 1522
rect 7317 1433 7517 1436
rect 6197 1387 6210 1433
rect 6384 1387 6397 1433
rect 6479 1387 6490 1433
rect 6664 1387 6675 1433
rect 6759 1387 6770 1433
rect 6944 1387 6955 1433
rect 7039 1387 7050 1433
rect 7224 1387 7235 1433
rect 7317 1387 7330 1433
rect 7504 1387 7517 1433
rect 6197 1373 6212 1387
rect 6268 1373 6322 1387
rect 6378 1373 6397 1387
rect 6197 1360 6397 1373
rect 6553 1311 6603 1387
rect 4591 1261 6603 1311
rect 6837 1309 6887 1387
rect 7317 1366 7331 1387
rect 7387 1366 7441 1387
rect 7497 1366 7517 1387
rect 7317 1356 7517 1366
rect 7597 1433 7797 1437
rect 7597 1368 7610 1433
rect 7784 1387 7797 1433
rect 7666 1368 7720 1387
rect 7776 1368 7797 1387
rect 7597 1360 7797 1368
rect 7877 1433 8077 1437
rect 7877 1387 7890 1433
rect 7877 1368 7898 1387
rect 7954 1368 8008 1387
rect 8064 1368 8077 1433
rect 7877 1360 8077 1368
rect 8157 1433 8357 1436
rect 8574 1433 8624 1490
rect 8787 1433 8837 1434
rect 9071 1433 9121 1434
rect 9277 1433 9477 1437
rect 8157 1387 8170 1433
rect 8344 1387 8357 1433
rect 8439 1387 8450 1433
rect 8624 1387 8635 1433
rect 8719 1387 8730 1433
rect 8904 1387 8915 1433
rect 8999 1387 9010 1433
rect 9184 1387 9195 1433
rect 9277 1387 9290 1433
rect 9464 1387 9477 1433
rect 8157 1366 8177 1387
rect 8233 1366 8287 1387
rect 8343 1366 8357 1387
rect 8157 1356 8357 1366
rect 8787 1309 8837 1387
rect 6837 1259 8837 1309
rect 9071 1311 9121 1387
rect 9277 1373 9296 1387
rect 9352 1373 9406 1387
rect 9462 1373 9477 1387
rect 9277 1360 9477 1373
rect 9557 1433 9757 1435
rect 9850 1433 9898 1517
rect 10571 1543 10588 1589
rect 10634 1543 10651 1589
rect 10571 1491 10651 1543
rect 10571 1445 10588 1491
rect 10634 1445 10651 1491
rect 10571 1442 10651 1445
rect 10300 1433 10651 1442
rect 9557 1387 9570 1433
rect 9744 1387 9757 1433
rect 9839 1387 9850 1433
rect 10024 1387 10035 1433
rect 10119 1387 10130 1433
rect 10304 1393 10651 1433
rect 10304 1387 10588 1393
rect 9557 1367 9576 1387
rect 9632 1367 9686 1387
rect 9742 1367 9757 1387
rect 10300 1385 10588 1387
rect 9557 1357 9757 1367
rect 10571 1347 10588 1385
rect 10634 1347 10651 1393
rect 10067 1311 10264 1315
rect 9071 1310 10264 1311
rect 9071 1261 10085 1310
rect 678 1249 875 1254
rect 236 1126 302 1141
rect 236 1070 241 1126
rect 297 1070 302 1126
rect 114 1004 180 1019
rect 114 948 119 1004
rect 175 948 180 1004
rect 114 894 180 948
rect 114 838 119 894
rect 175 838 180 894
rect 114 832 180 838
rect 113 822 180 832
rect 236 1016 302 1070
rect 236 960 241 1016
rect 297 960 302 1016
rect 236 944 302 960
rect 0 412 66 427
rect 0 356 5 412
rect 61 356 66 412
rect 0 302 66 356
rect 0 246 5 302
rect 61 246 66 302
rect 0 232 66 246
rect 0 230 65 232
rect 2 -230 65 230
rect 0 -232 65 -230
rect 0 -246 66 -232
rect 0 -302 5 -246
rect 61 -302 66 -246
rect 0 -356 66 -302
rect 0 -412 5 -356
rect 61 -412 66 -356
rect 0 -427 66 -412
rect 113 -822 176 822
rect 113 -832 180 -822
rect 114 -838 180 -832
rect 114 -894 119 -838
rect 175 -894 180 -838
rect 114 -948 180 -894
rect 114 -1004 119 -948
rect 175 -1004 180 -948
rect 114 -1019 180 -1004
rect 236 -944 299 944
rect 236 -960 302 -944
rect 236 -1016 241 -960
rect 297 -1016 302 -960
rect 236 -1070 302 -1016
rect 236 -1126 241 -1070
rect 297 -1126 302 -1070
rect 236 -1141 302 -1126
rect 348 -1249 411 1249
rect 543 1197 623 1249
rect 543 1151 560 1197
rect 606 1151 623 1197
rect 543 1122 623 1151
rect 543 1101 931 1122
rect 1437 1117 1637 1127
rect 543 1099 890 1101
rect 543 1053 560 1099
rect 606 1056 890 1099
rect 606 1053 623 1056
rect 879 1055 890 1056
rect 1064 1055 1075 1101
rect 1159 1055 1170 1101
rect 1344 1055 1355 1101
rect 1437 1055 1450 1117
rect 1506 1101 1560 1117
rect 1616 1101 1637 1117
rect 1624 1055 1637 1101
rect 543 1001 623 1053
rect 543 955 560 1001
rect 606 955 623 1001
rect 543 903 623 955
rect 669 1005 866 1010
rect 669 949 682 1005
rect 738 949 792 1005
rect 848 1002 866 1005
rect 1170 1002 1216 1055
rect 1437 1050 1637 1055
rect 1717 1118 1917 1128
rect 1717 1055 1730 1118
rect 1786 1101 1840 1118
rect 1896 1101 1917 1118
rect 2837 1116 3037 1128
rect 2569 1101 2619 1102
rect 2837 1101 2852 1116
rect 2908 1101 2962 1116
rect 3018 1101 3037 1116
rect 1904 1055 1917 1101
rect 1999 1055 2010 1101
rect 2184 1055 2290 1101
rect 2464 1055 2475 1101
rect 2559 1055 2570 1101
rect 2744 1055 2755 1101
rect 2837 1055 2850 1101
rect 3024 1055 3037 1101
rect 3119 1116 3316 1121
rect 3119 1101 3135 1116
rect 3191 1101 3245 1116
rect 3301 1101 3316 1116
rect 3399 1116 3596 1121
rect 3399 1101 3415 1116
rect 3471 1101 3525 1116
rect 3581 1101 3596 1116
rect 3119 1055 3130 1101
rect 3304 1055 3410 1101
rect 3584 1055 3596 1101
rect 3677 1116 3877 1128
rect 3677 1101 3696 1116
rect 3752 1101 3806 1116
rect 3862 1101 3877 1116
rect 4797 1118 4997 1128
rect 4095 1101 4145 1102
rect 4797 1101 4818 1118
rect 4874 1101 4928 1118
rect 3677 1055 3690 1101
rect 3864 1055 3877 1101
rect 3959 1055 3970 1101
rect 4144 1055 4155 1101
rect 4239 1055 4250 1101
rect 4424 1055 4530 1101
rect 4704 1055 4715 1101
rect 4797 1055 4810 1101
rect 4984 1055 4997 1118
rect 1717 1051 1917 1055
rect 848 956 1216 1002
rect 2569 999 2619 1055
rect 2837 1050 3037 1055
rect 3677 1050 3877 1055
rect 848 949 866 956
rect 669 944 866 949
rect 1736 953 2619 999
rect 4095 999 4145 1055
rect 4797 1051 4997 1055
rect 5077 1117 5277 1127
rect 5077 1101 5098 1117
rect 5154 1101 5208 1117
rect 5077 1055 5090 1101
rect 5264 1055 5277 1117
rect 5917 1117 6117 1127
rect 5359 1055 5370 1101
rect 5544 1055 5555 1101
rect 5639 1055 5650 1101
rect 5824 1055 5835 1101
rect 5917 1055 5930 1117
rect 5986 1101 6040 1117
rect 6096 1101 6117 1117
rect 6104 1055 6117 1101
rect 5077 1050 5277 1055
rect 5498 1009 5544 1055
rect 5650 1009 5696 1055
rect 5917 1050 6117 1055
rect 6197 1118 6397 1128
rect 6197 1055 6210 1118
rect 6266 1101 6320 1118
rect 6376 1101 6397 1118
rect 7317 1116 7517 1128
rect 7049 1101 7099 1102
rect 7317 1101 7332 1116
rect 7388 1101 7442 1116
rect 7498 1101 7517 1116
rect 8157 1116 8357 1128
rect 8157 1101 8176 1116
rect 8232 1101 8286 1116
rect 8342 1101 8357 1116
rect 9277 1118 9477 1128
rect 8575 1101 8625 1102
rect 9277 1101 9298 1118
rect 9354 1101 9408 1118
rect 6384 1055 6397 1101
rect 6479 1055 6490 1101
rect 6664 1055 6770 1101
rect 6944 1055 6955 1101
rect 7039 1055 7050 1101
rect 7224 1055 7235 1101
rect 7317 1055 7330 1101
rect 7504 1055 7517 1101
rect 7599 1055 7610 1101
rect 7784 1055 7890 1101
rect 8064 1055 8075 1101
rect 8157 1055 8170 1101
rect 8344 1055 8357 1101
rect 8439 1055 8450 1101
rect 8624 1055 8635 1101
rect 8719 1055 8730 1101
rect 8904 1055 9010 1101
rect 9184 1055 9195 1101
rect 9277 1055 9290 1101
rect 9464 1055 9477 1118
rect 6197 1051 6397 1055
rect 4095 953 4978 999
rect 5466 963 5696 1009
rect 7049 999 7099 1055
rect 7317 1050 7517 1055
rect 8157 1050 8357 1055
rect 543 857 560 903
rect 606 857 623 903
rect 543 805 623 857
rect 932 888 1129 893
rect 932 832 948 888
rect 1004 832 1058 888
rect 1114 873 1129 888
rect 1114 832 1216 873
rect 932 827 1216 832
rect 543 759 560 805
rect 606 782 623 805
rect 606 781 895 782
rect 1170 781 1216 827
rect 1437 781 1637 785
rect 1736 781 1782 953
rect 1831 889 1911 894
rect 1831 833 1843 889
rect 1899 883 1911 889
rect 4803 889 4883 894
rect 4803 883 4815 889
rect 1899 837 2620 883
rect 1899 833 1911 837
rect 1831 827 1911 833
rect 1997 781 2197 785
rect 606 759 890 781
rect 543 735 890 759
rect 1064 735 1075 781
rect 1159 735 1170 781
rect 1344 735 1355 781
rect 543 707 623 735
rect 1437 719 1450 781
rect 1624 735 1637 781
rect 1719 735 1730 781
rect 1904 735 1915 781
rect 1997 735 2010 781
rect 2184 735 2197 781
rect 1506 719 1560 735
rect 1616 719 1637 735
rect 1437 708 1637 719
rect 1997 718 2011 735
rect 2067 718 2121 735
rect 2177 718 2197 735
rect 1997 708 2197 718
rect 2277 781 2477 785
rect 2570 781 2620 837
rect 4094 837 4815 883
rect 4094 781 4144 837
rect 4803 833 4815 837
rect 4871 833 4883 889
rect 4803 827 4883 833
rect 4237 781 4437 785
rect 2277 735 2290 781
rect 2464 735 2477 781
rect 2559 735 2570 781
rect 2744 735 2755 781
rect 2839 735 2850 781
rect 3024 735 3130 781
rect 3304 735 3315 781
rect 3399 735 3410 781
rect 3584 735 3690 781
rect 3864 735 3875 781
rect 3959 735 3970 781
rect 4144 735 4155 781
rect 4237 735 4250 781
rect 4424 735 4437 781
rect 2277 719 2292 735
rect 2348 719 2402 735
rect 2458 719 2477 735
rect 2277 708 2477 719
rect 4237 719 4256 735
rect 4312 719 4366 735
rect 4422 719 4437 735
rect 4237 708 4437 719
rect 4517 781 4717 785
rect 4932 781 4978 953
rect 6216 953 7099 999
rect 8575 999 8625 1055
rect 9277 1051 9477 1055
rect 9557 1117 9757 1127
rect 9557 1101 9578 1117
rect 9634 1101 9688 1117
rect 9557 1055 9570 1101
rect 9744 1055 9757 1117
rect 9850 1101 9908 1261
rect 10067 1254 10085 1261
rect 10141 1254 10195 1310
rect 10251 1254 10264 1310
rect 10067 1249 10264 1254
rect 10571 1295 10651 1347
rect 10571 1249 10588 1295
rect 10634 1249 10651 1295
rect 10571 1197 10651 1249
rect 10571 1151 10588 1197
rect 10634 1151 10651 1197
rect 10571 1104 10651 1151
rect 10299 1101 10651 1104
rect 9839 1055 9850 1101
rect 10024 1055 10035 1101
rect 10119 1055 10130 1101
rect 10304 1099 10651 1101
rect 10304 1055 10588 1099
rect 9557 1050 9757 1055
rect 10299 1053 10588 1055
rect 10634 1053 10651 1099
rect 10299 1047 10651 1053
rect 10571 1001 10651 1047
rect 8575 953 9458 999
rect 5466 827 5696 873
rect 5077 781 5277 785
rect 5498 781 5544 827
rect 5650 781 5696 827
rect 5917 781 6117 785
rect 6216 781 6262 953
rect 6311 889 6391 894
rect 6311 833 6323 889
rect 6379 883 6391 889
rect 9283 889 9363 894
rect 9283 883 9295 889
rect 6379 837 7100 883
rect 6379 833 6391 837
rect 6311 827 6391 833
rect 6477 781 6677 785
rect 4517 735 4530 781
rect 4704 735 4717 781
rect 4799 735 4810 781
rect 4984 735 4995 781
rect 5077 735 5090 781
rect 4517 718 4537 735
rect 4593 718 4647 735
rect 4703 718 4717 735
rect 4517 708 4717 718
rect 5077 719 5098 735
rect 5154 719 5208 735
rect 5264 719 5277 781
rect 5359 735 5370 781
rect 5544 735 5555 781
rect 5639 735 5650 781
rect 5824 735 5835 781
rect 5077 708 5277 719
rect 5917 719 5930 781
rect 6104 735 6117 781
rect 6199 735 6210 781
rect 6384 735 6395 781
rect 6477 735 6490 781
rect 6664 735 6677 781
rect 5986 719 6040 735
rect 6096 719 6117 735
rect 5917 708 6117 719
rect 6477 718 6491 735
rect 6547 718 6601 735
rect 6657 718 6677 735
rect 6477 708 6677 718
rect 6757 781 6957 785
rect 7050 781 7100 837
rect 8574 837 9295 883
rect 8574 781 8624 837
rect 9283 833 9295 837
rect 9351 833 9363 889
rect 9283 827 9363 833
rect 8717 781 8917 785
rect 6757 735 6770 781
rect 6944 735 6957 781
rect 7039 735 7050 781
rect 7224 735 7235 781
rect 7319 735 7330 781
rect 7504 735 7610 781
rect 7784 735 7795 781
rect 7879 735 7890 781
rect 8064 735 8170 781
rect 8344 735 8355 781
rect 8439 735 8450 781
rect 8624 735 8635 781
rect 8717 735 8730 781
rect 8904 735 8917 781
rect 6757 719 6772 735
rect 6828 719 6882 735
rect 6938 719 6957 735
rect 6757 708 6957 719
rect 8717 719 8736 735
rect 8792 719 8846 735
rect 8902 719 8917 735
rect 8717 708 8917 719
rect 8997 781 9197 785
rect 9412 781 9458 953
rect 10571 955 10588 1001
rect 10634 955 10651 1001
rect 10571 903 10651 955
rect 10066 888 10263 893
rect 10066 874 10084 888
rect 10024 873 10084 874
rect 9978 832 10084 873
rect 10140 832 10194 888
rect 10250 832 10263 888
rect 9978 827 10263 832
rect 10571 857 10588 903
rect 10634 857 10651 903
rect 9557 781 9757 785
rect 9978 781 10024 827
rect 10571 805 10651 857
rect 10571 786 10588 805
rect 8997 735 9010 781
rect 9184 735 9197 781
rect 9279 735 9290 781
rect 9464 735 9475 781
rect 9557 735 9570 781
rect 8997 718 9017 735
rect 9073 718 9127 735
rect 9183 718 9197 735
rect 8997 708 9197 718
rect 9557 719 9578 735
rect 9634 719 9688 735
rect 9744 719 9757 781
rect 9839 735 9850 781
rect 10024 735 10035 781
rect 10119 735 10130 781
rect 10304 759 10588 786
rect 10634 759 10651 805
rect 10304 729 10651 759
rect 9557 708 9757 719
rect 543 661 560 707
rect 606 661 623 707
rect 10571 707 10651 729
rect 543 609 623 661
rect 543 563 560 609
rect 606 563 623 609
rect 670 664 867 669
rect 670 608 683 664
rect 739 608 793 664
rect 849 662 867 664
rect 10315 664 10517 669
rect 10315 662 10333 664
rect 849 612 2620 662
rect 849 608 867 612
rect 670 603 867 608
rect 543 511 623 563
rect 543 465 560 511
rect 606 465 623 511
rect 543 456 623 465
rect 1439 472 1636 477
rect 543 449 909 456
rect 1439 449 1452 472
rect 1508 449 1562 472
rect 1618 449 1636 472
rect 1997 474 2194 479
rect 543 413 890 449
rect 543 367 560 413
rect 606 403 890 413
rect 1064 403 1075 449
rect 1159 403 1170 449
rect 1344 403 1450 449
rect 1624 411 1636 449
rect 1624 403 1635 411
rect 1719 403 1730 449
rect 1904 403 1915 449
rect 1997 413 2010 474
rect 2066 449 2120 474
rect 2176 449 2194 474
rect 2570 449 2620 612
rect 4094 612 7100 662
rect 2837 461 3037 476
rect 1999 403 2010 413
rect 2184 403 2195 449
rect 2279 403 2290 449
rect 2464 403 2475 449
rect 2559 403 2570 449
rect 2744 403 2755 449
rect 2837 405 2849 461
rect 2905 449 2959 461
rect 3015 449 3037 461
rect 3677 461 3877 476
rect 3677 449 3699 461
rect 3755 449 3809 461
rect 2837 403 2850 405
rect 3024 403 3037 449
rect 3119 403 3130 449
rect 3304 403 3410 449
rect 3584 403 3595 449
rect 3677 403 3690 449
rect 3865 405 3877 461
rect 4094 449 4144 612
rect 4915 501 6279 551
rect 4915 475 4984 501
rect 4914 449 4984 475
rect 6210 475 6279 501
rect 6210 449 6280 475
rect 7050 449 7100 612
rect 8574 612 10333 662
rect 7317 461 7517 476
rect 3864 403 3877 405
rect 3959 403 3970 449
rect 4144 403 4155 449
rect 4239 403 4250 449
rect 4424 403 4435 449
rect 4519 403 4530 449
rect 4704 403 4715 449
rect 4799 403 4810 449
rect 4984 403 4995 449
rect 5079 403 5090 449
rect 5264 403 5370 449
rect 5544 403 5555 449
rect 5639 403 5650 449
rect 5824 403 5930 449
rect 6104 403 6115 449
rect 6199 403 6210 449
rect 6384 403 6395 449
rect 6479 403 6490 449
rect 6664 403 6675 449
rect 6759 403 6770 449
rect 6944 403 6955 449
rect 7039 403 7050 449
rect 7224 403 7235 449
rect 7317 405 7329 461
rect 7385 449 7439 461
rect 7495 449 7517 461
rect 8157 461 8357 476
rect 8157 449 8179 461
rect 8235 449 8289 461
rect 7317 403 7330 405
rect 7504 403 7517 449
rect 7599 403 7610 449
rect 7784 403 7890 449
rect 8064 403 8075 449
rect 8157 403 8170 449
rect 8345 405 8357 461
rect 8574 449 8624 612
rect 10315 608 10333 612
rect 10389 608 10443 664
rect 10499 608 10517 664
rect 10315 603 10517 608
rect 10571 661 10588 707
rect 10634 661 10651 707
rect 10571 609 10651 661
rect 10065 561 10262 566
rect 10065 551 10083 561
rect 9395 505 10083 551
rect 10139 505 10193 561
rect 10249 505 10262 561
rect 9395 501 10262 505
rect 9395 475 9464 501
rect 10065 500 10262 501
rect 10571 563 10588 609
rect 10634 563 10651 609
rect 10571 511 10651 563
rect 9394 449 9464 475
rect 10571 465 10588 511
rect 10634 465 10651 511
rect 10571 456 10651 465
rect 10292 449 10651 456
rect 8344 403 8357 405
rect 8439 403 8450 449
rect 8624 403 8635 449
rect 8719 403 8730 449
rect 8904 403 8915 449
rect 8999 403 9010 449
rect 9184 403 9195 449
rect 9279 403 9290 449
rect 9464 403 9475 449
rect 9559 403 9570 449
rect 9744 403 9850 449
rect 10024 403 10035 449
rect 10119 403 10130 449
rect 10304 413 10651 449
rect 10304 403 10588 413
rect 606 399 909 403
rect 606 367 623 399
rect 543 315 623 367
rect 543 269 560 315
rect 606 269 623 315
rect 543 217 623 269
rect 674 291 871 296
rect 674 235 687 291
rect 743 235 797 291
rect 853 289 871 291
rect 1814 289 1904 403
rect 2011 289 2064 403
rect 853 236 2064 289
rect 853 235 871 236
rect 674 230 871 235
rect 2011 229 2064 236
rect 2409 284 2462 403
rect 2837 399 3037 403
rect 3677 399 3877 403
rect 4252 284 4305 403
rect 2409 231 4305 284
rect 4650 289 4703 403
rect 6491 289 6544 403
rect 4650 236 6544 289
rect 4650 229 4703 236
rect 6491 229 6544 236
rect 6889 284 6942 403
rect 7317 399 7517 403
rect 8157 399 8357 403
rect 8732 284 8785 403
rect 6889 231 8785 284
rect 9130 289 9183 403
rect 10292 399 10588 403
rect 10571 367 10588 399
rect 10634 367 10651 413
rect 10571 315 10651 367
rect 10295 291 10492 296
rect 10295 289 10313 291
rect 9130 236 10313 289
rect 9130 229 9183 236
rect 10295 235 10313 236
rect 10369 235 10423 291
rect 10479 235 10492 291
rect 10295 230 10492 235
rect 10571 269 10588 315
rect 10634 269 10651 315
rect 543 171 560 217
rect 606 171 623 217
rect 543 136 623 171
rect 10571 217 10651 269
rect 10571 171 10588 217
rect 10634 171 10651 217
rect 10571 136 10651 171
rect 543 119 10651 136
rect 543 73 560 119
rect 606 73 658 119
rect 704 73 756 119
rect 802 73 854 119
rect 900 73 952 119
rect 998 73 1050 119
rect 1096 73 1148 119
rect 1194 73 1246 119
rect 1292 73 1344 119
rect 1390 73 1442 119
rect 1488 73 1540 119
rect 1586 73 1638 119
rect 1684 73 1736 119
rect 1782 73 1834 119
rect 1880 73 1932 119
rect 1978 73 2030 119
rect 2076 73 2128 119
rect 2174 73 2226 119
rect 2272 73 2324 119
rect 2370 73 2422 119
rect 2468 73 2520 119
rect 2566 73 2618 119
rect 2664 73 2716 119
rect 2762 73 2814 119
rect 2860 73 2912 119
rect 2958 73 3010 119
rect 3056 73 3108 119
rect 3154 73 3206 119
rect 3252 73 3304 119
rect 3350 73 3402 119
rect 3448 73 3500 119
rect 3546 73 3598 119
rect 3644 73 3696 119
rect 3742 73 3794 119
rect 3840 73 3892 119
rect 3938 73 3990 119
rect 4036 73 4088 119
rect 4134 73 4186 119
rect 4232 73 4284 119
rect 4330 73 4382 119
rect 4428 73 4480 119
rect 4526 73 4578 119
rect 4624 73 4676 119
rect 4722 73 4774 119
rect 4820 73 4872 119
rect 4918 73 4970 119
rect 5016 73 5068 119
rect 5114 73 5166 119
rect 5212 73 5264 119
rect 5310 73 5362 119
rect 5408 73 5460 119
rect 5506 73 5558 119
rect 5604 73 5656 119
rect 5702 73 5754 119
rect 5800 73 5852 119
rect 5898 73 5950 119
rect 5996 73 6048 119
rect 6094 73 6146 119
rect 6192 73 6244 119
rect 6290 73 6342 119
rect 6388 73 6440 119
rect 6486 73 6538 119
rect 6584 73 6636 119
rect 6682 73 6734 119
rect 6780 73 6832 119
rect 6878 73 6930 119
rect 6976 73 7028 119
rect 7074 73 7126 119
rect 7172 73 7224 119
rect 7270 73 7322 119
rect 7368 73 7420 119
rect 7466 73 7518 119
rect 7564 73 7616 119
rect 7662 73 7714 119
rect 7760 73 7812 119
rect 7858 73 7910 119
rect 7956 73 8008 119
rect 8054 73 8106 119
rect 8152 73 8204 119
rect 8250 73 8302 119
rect 8348 73 8400 119
rect 8446 73 8498 119
rect 8544 73 8596 119
rect 8642 73 8694 119
rect 8740 73 8792 119
rect 8838 73 8890 119
rect 8936 73 8988 119
rect 9034 73 9086 119
rect 9132 73 9184 119
rect 9230 73 9282 119
rect 9328 73 9380 119
rect 9426 73 9478 119
rect 9524 73 9576 119
rect 9622 73 9674 119
rect 9720 73 9772 119
rect 9818 73 9870 119
rect 9916 73 9968 119
rect 10014 73 10066 119
rect 10112 73 10164 119
rect 10210 73 10262 119
rect 10308 73 10360 119
rect 10406 73 10458 119
rect 10504 73 10588 119
rect 10634 73 10651 119
rect 543 56 10651 73
rect 10704 1324 10767 1339
rect 10704 1268 10709 1324
rect 10765 1268 10767 1324
rect 10704 1214 10767 1268
rect 10704 1158 10709 1214
rect 10765 1158 10767 1214
rect 582 -56 10497 56
rect 543 -73 10651 -56
rect 543 -119 560 -73
rect 606 -119 658 -73
rect 704 -119 756 -73
rect 802 -119 854 -73
rect 900 -119 952 -73
rect 998 -119 1050 -73
rect 1096 -119 1148 -73
rect 1194 -119 1246 -73
rect 1292 -119 1344 -73
rect 1390 -119 1442 -73
rect 1488 -119 1540 -73
rect 1586 -119 1638 -73
rect 1684 -119 1736 -73
rect 1782 -119 1834 -73
rect 1880 -119 1932 -73
rect 1978 -119 2030 -73
rect 2076 -119 2128 -73
rect 2174 -119 2226 -73
rect 2272 -119 2324 -73
rect 2370 -119 2422 -73
rect 2468 -119 2520 -73
rect 2566 -119 2618 -73
rect 2664 -119 2716 -73
rect 2762 -119 2814 -73
rect 2860 -119 2912 -73
rect 2958 -119 3010 -73
rect 3056 -119 3108 -73
rect 3154 -119 3206 -73
rect 3252 -119 3304 -73
rect 3350 -119 3402 -73
rect 3448 -119 3500 -73
rect 3546 -119 3598 -73
rect 3644 -119 3696 -73
rect 3742 -119 3794 -73
rect 3840 -119 3892 -73
rect 3938 -119 3990 -73
rect 4036 -119 4088 -73
rect 4134 -119 4186 -73
rect 4232 -119 4284 -73
rect 4330 -119 4382 -73
rect 4428 -119 4480 -73
rect 4526 -119 4578 -73
rect 4624 -119 4676 -73
rect 4722 -119 4774 -73
rect 4820 -119 4872 -73
rect 4918 -119 4970 -73
rect 5016 -119 5068 -73
rect 5114 -119 5166 -73
rect 5212 -119 5264 -73
rect 5310 -119 5362 -73
rect 5408 -119 5460 -73
rect 5506 -119 5558 -73
rect 5604 -119 5656 -73
rect 5702 -119 5754 -73
rect 5800 -119 5852 -73
rect 5898 -119 5950 -73
rect 5996 -119 6048 -73
rect 6094 -119 6146 -73
rect 6192 -119 6244 -73
rect 6290 -119 6342 -73
rect 6388 -119 6440 -73
rect 6486 -119 6538 -73
rect 6584 -119 6636 -73
rect 6682 -119 6734 -73
rect 6780 -119 6832 -73
rect 6878 -119 6930 -73
rect 6976 -119 7028 -73
rect 7074 -119 7126 -73
rect 7172 -119 7224 -73
rect 7270 -119 7322 -73
rect 7368 -119 7420 -73
rect 7466 -119 7518 -73
rect 7564 -119 7616 -73
rect 7662 -119 7714 -73
rect 7760 -119 7812 -73
rect 7858 -119 7910 -73
rect 7956 -119 8008 -73
rect 8054 -119 8106 -73
rect 8152 -119 8204 -73
rect 8250 -119 8302 -73
rect 8348 -119 8400 -73
rect 8446 -119 8498 -73
rect 8544 -119 8596 -73
rect 8642 -119 8694 -73
rect 8740 -119 8792 -73
rect 8838 -119 8890 -73
rect 8936 -119 8988 -73
rect 9034 -119 9086 -73
rect 9132 -119 9184 -73
rect 9230 -119 9282 -73
rect 9328 -119 9380 -73
rect 9426 -119 9478 -73
rect 9524 -119 9576 -73
rect 9622 -119 9674 -73
rect 9720 -119 9772 -73
rect 9818 -119 9870 -73
rect 9916 -119 9968 -73
rect 10014 -119 10066 -73
rect 10112 -119 10164 -73
rect 10210 -119 10262 -73
rect 10308 -119 10360 -73
rect 10406 -119 10458 -73
rect 10504 -119 10588 -73
rect 10634 -119 10651 -73
rect 543 -136 10651 -119
rect 543 -171 623 -136
rect 543 -217 560 -171
rect 606 -217 623 -171
rect 543 -269 623 -217
rect 10571 -171 10651 -136
rect 10571 -217 10588 -171
rect 10634 -217 10651 -171
rect 543 -315 560 -269
rect 606 -315 623 -269
rect 674 -235 871 -230
rect 674 -291 687 -235
rect 743 -291 797 -235
rect 853 -236 871 -235
rect 2011 -236 2064 -229
rect 853 -289 2064 -236
rect 853 -291 871 -289
rect 674 -296 871 -291
rect 543 -367 623 -315
rect 543 -413 560 -367
rect 606 -399 623 -367
rect 606 -403 909 -399
rect 1814 -403 1904 -289
rect 2011 -403 2064 -289
rect 2409 -284 4305 -231
rect 2409 -403 2462 -284
rect 2837 -403 3037 -399
rect 3677 -403 3877 -399
rect 4252 -403 4305 -284
rect 4650 -236 4703 -229
rect 6491 -236 6544 -229
rect 4650 -289 6544 -236
rect 4650 -403 4703 -289
rect 6491 -403 6544 -289
rect 6889 -284 8785 -231
rect 6889 -403 6942 -284
rect 7317 -403 7517 -399
rect 8157 -403 8357 -399
rect 8732 -403 8785 -284
rect 9130 -236 9183 -229
rect 10295 -235 10492 -230
rect 10295 -236 10313 -235
rect 9130 -289 10313 -236
rect 9130 -403 9183 -289
rect 10295 -291 10313 -289
rect 10369 -291 10423 -235
rect 10479 -291 10492 -235
rect 10295 -296 10492 -291
rect 10571 -269 10651 -217
rect 10571 -315 10588 -269
rect 10634 -315 10651 -269
rect 10571 -367 10651 -315
rect 10571 -399 10588 -367
rect 10292 -403 10588 -399
rect 606 -413 890 -403
rect 543 -449 890 -413
rect 1064 -449 1075 -403
rect 1159 -449 1170 -403
rect 1344 -449 1450 -403
rect 1624 -411 1635 -403
rect 1624 -449 1636 -411
rect 1719 -449 1730 -403
rect 1904 -449 1915 -403
rect 1999 -413 2010 -403
rect 543 -456 909 -449
rect 543 -465 623 -456
rect 543 -511 560 -465
rect 606 -511 623 -465
rect 1439 -472 1452 -449
rect 1508 -472 1562 -449
rect 1618 -472 1636 -449
rect 1439 -477 1636 -472
rect 1997 -474 2010 -413
rect 2184 -449 2195 -403
rect 2279 -449 2290 -403
rect 2464 -449 2475 -403
rect 2559 -449 2570 -403
rect 2744 -449 2755 -403
rect 2837 -405 2850 -403
rect 2066 -474 2120 -449
rect 2176 -474 2194 -449
rect 1997 -479 2194 -474
rect 543 -563 623 -511
rect 543 -609 560 -563
rect 606 -609 623 -563
rect 543 -661 623 -609
rect 543 -707 560 -661
rect 606 -707 623 -661
rect 670 -608 867 -603
rect 670 -664 683 -608
rect 739 -664 793 -608
rect 849 -612 867 -608
rect 2570 -612 2620 -449
rect 2837 -461 2849 -405
rect 3024 -449 3037 -403
rect 3119 -449 3130 -403
rect 3304 -449 3410 -403
rect 3584 -449 3595 -403
rect 3677 -449 3690 -403
rect 3864 -405 3877 -403
rect 2905 -461 2959 -449
rect 3015 -461 3037 -449
rect 2837 -476 3037 -461
rect 3677 -461 3699 -449
rect 3755 -461 3809 -449
rect 3865 -461 3877 -405
rect 3959 -449 3970 -403
rect 4144 -449 4155 -403
rect 4239 -449 4250 -403
rect 4424 -449 4435 -403
rect 4519 -449 4530 -403
rect 4704 -449 4715 -403
rect 4799 -449 4810 -403
rect 4984 -449 4995 -403
rect 5079 -449 5090 -403
rect 5264 -449 5370 -403
rect 5544 -449 5555 -403
rect 5639 -449 5650 -403
rect 5824 -449 5930 -403
rect 6104 -449 6115 -403
rect 6199 -449 6210 -403
rect 6384 -449 6395 -403
rect 6479 -449 6490 -403
rect 6664 -449 6675 -403
rect 6759 -449 6770 -403
rect 6944 -449 6955 -403
rect 7039 -449 7050 -403
rect 7224 -449 7235 -403
rect 7317 -405 7330 -403
rect 3677 -476 3877 -461
rect 849 -662 2620 -612
rect 4094 -612 4144 -449
rect 4914 -475 4984 -449
rect 4915 -501 4984 -475
rect 6210 -475 6280 -449
rect 6210 -501 6279 -475
rect 4915 -551 6279 -501
rect 7050 -612 7100 -449
rect 7317 -461 7329 -405
rect 7504 -449 7517 -403
rect 7599 -449 7610 -403
rect 7784 -449 7890 -403
rect 8064 -449 8075 -403
rect 8157 -449 8170 -403
rect 8344 -405 8357 -403
rect 7385 -461 7439 -449
rect 7495 -461 7517 -449
rect 7317 -476 7517 -461
rect 8157 -461 8179 -449
rect 8235 -461 8289 -449
rect 8345 -461 8357 -405
rect 8439 -449 8450 -403
rect 8624 -449 8635 -403
rect 8719 -449 8730 -403
rect 8904 -449 8915 -403
rect 8999 -449 9010 -403
rect 9184 -449 9195 -403
rect 9279 -449 9290 -403
rect 9464 -449 9475 -403
rect 9559 -449 9570 -403
rect 9744 -449 9850 -403
rect 10024 -449 10035 -403
rect 10119 -449 10130 -403
rect 10304 -413 10588 -403
rect 10634 -413 10651 -367
rect 10304 -449 10651 -413
rect 8157 -476 8357 -461
rect 4094 -662 7100 -612
rect 8574 -612 8624 -449
rect 9394 -475 9464 -449
rect 10292 -456 10651 -449
rect 9395 -501 9464 -475
rect 10571 -465 10651 -456
rect 10065 -501 10262 -500
rect 9395 -505 10262 -501
rect 9395 -551 10083 -505
rect 10065 -561 10083 -551
rect 10139 -561 10193 -505
rect 10249 -561 10262 -505
rect 10065 -566 10262 -561
rect 10571 -511 10588 -465
rect 10634 -511 10651 -465
rect 10571 -563 10651 -511
rect 10315 -608 10517 -603
rect 10315 -612 10333 -608
rect 8574 -662 10333 -612
rect 849 -664 867 -662
rect 670 -669 867 -664
rect 10315 -664 10333 -662
rect 10389 -664 10443 -608
rect 10499 -664 10517 -608
rect 10315 -669 10517 -664
rect 10571 -609 10588 -563
rect 10634 -609 10651 -563
rect 10571 -661 10651 -609
rect 543 -735 623 -707
rect 10571 -707 10588 -661
rect 10634 -707 10651 -661
rect 1437 -719 1637 -708
rect 543 -759 890 -735
rect 543 -805 560 -759
rect 606 -781 890 -759
rect 1064 -781 1075 -735
rect 1159 -781 1170 -735
rect 1344 -781 1355 -735
rect 1437 -781 1450 -719
rect 1506 -735 1560 -719
rect 1616 -735 1637 -719
rect 1997 -718 2197 -708
rect 1997 -735 2011 -718
rect 2067 -735 2121 -718
rect 2177 -735 2197 -718
rect 1624 -781 1637 -735
rect 1719 -781 1730 -735
rect 1904 -781 1915 -735
rect 1997 -781 2010 -735
rect 2184 -781 2197 -735
rect 606 -782 895 -781
rect 606 -805 623 -782
rect 543 -857 623 -805
rect 1170 -827 1216 -781
rect 1437 -785 1637 -781
rect 543 -903 560 -857
rect 606 -903 623 -857
rect 932 -832 1216 -827
rect 932 -888 948 -832
rect 1004 -888 1058 -832
rect 1114 -873 1216 -832
rect 1114 -888 1129 -873
rect 932 -893 1129 -888
rect 543 -955 623 -903
rect 543 -1001 560 -955
rect 606 -1001 623 -955
rect 543 -1053 623 -1001
rect 669 -949 866 -944
rect 669 -1005 682 -949
rect 738 -1005 792 -949
rect 848 -956 866 -949
rect 1736 -953 1782 -781
rect 1997 -785 2197 -781
rect 2277 -719 2477 -708
rect 2277 -735 2292 -719
rect 2348 -735 2402 -719
rect 2458 -735 2477 -719
rect 4237 -719 4437 -708
rect 4237 -735 4256 -719
rect 4312 -735 4366 -719
rect 4422 -735 4437 -719
rect 2277 -781 2290 -735
rect 2464 -781 2477 -735
rect 2559 -781 2570 -735
rect 2744 -781 2755 -735
rect 2839 -781 2850 -735
rect 3024 -781 3130 -735
rect 3304 -781 3315 -735
rect 3399 -781 3410 -735
rect 3584 -781 3690 -735
rect 3864 -781 3875 -735
rect 3959 -781 3970 -735
rect 4144 -781 4155 -735
rect 4237 -781 4250 -735
rect 4424 -781 4437 -735
rect 2277 -785 2477 -781
rect 1831 -833 1911 -827
rect 1831 -889 1843 -833
rect 1899 -837 1911 -833
rect 2570 -837 2620 -781
rect 1899 -883 2620 -837
rect 4094 -837 4144 -781
rect 4237 -785 4437 -781
rect 4517 -718 4717 -708
rect 4517 -735 4537 -718
rect 4593 -735 4647 -718
rect 4703 -735 4717 -718
rect 5077 -719 5277 -708
rect 5077 -735 5098 -719
rect 5154 -735 5208 -719
rect 4517 -781 4530 -735
rect 4704 -781 4717 -735
rect 4799 -781 4810 -735
rect 4984 -781 4995 -735
rect 5077 -781 5090 -735
rect 5264 -781 5277 -719
rect 5917 -719 6117 -708
rect 5359 -781 5370 -735
rect 5544 -781 5555 -735
rect 5639 -781 5650 -735
rect 5824 -781 5835 -735
rect 5917 -781 5930 -719
rect 5986 -735 6040 -719
rect 6096 -735 6117 -719
rect 6477 -718 6677 -708
rect 6477 -735 6491 -718
rect 6547 -735 6601 -718
rect 6657 -735 6677 -718
rect 6104 -781 6117 -735
rect 6199 -781 6210 -735
rect 6384 -781 6395 -735
rect 6477 -781 6490 -735
rect 6664 -781 6677 -735
rect 4517 -785 4717 -781
rect 4803 -833 4883 -827
rect 4803 -837 4815 -833
rect 4094 -883 4815 -837
rect 1899 -889 1911 -883
rect 1831 -894 1911 -889
rect 4803 -889 4815 -883
rect 4871 -889 4883 -833
rect 4803 -894 4883 -889
rect 4932 -953 4978 -781
rect 5077 -785 5277 -781
rect 5498 -827 5544 -781
rect 5650 -827 5696 -781
rect 5917 -785 6117 -781
rect 5466 -873 5696 -827
rect 848 -1002 1216 -956
rect 1736 -999 2619 -953
rect 848 -1005 866 -1002
rect 669 -1010 866 -1005
rect 543 -1099 560 -1053
rect 606 -1056 623 -1053
rect 1170 -1055 1216 -1002
rect 1437 -1055 1637 -1050
rect 879 -1056 890 -1055
rect 606 -1099 890 -1056
rect 543 -1101 890 -1099
rect 1064 -1101 1075 -1055
rect 1159 -1101 1170 -1055
rect 1344 -1101 1355 -1055
rect 543 -1122 931 -1101
rect 1437 -1117 1450 -1055
rect 1624 -1101 1637 -1055
rect 1506 -1117 1560 -1101
rect 1616 -1117 1637 -1101
rect 543 -1151 623 -1122
rect 1437 -1127 1637 -1117
rect 1717 -1055 1917 -1051
rect 2569 -1055 2619 -999
rect 4095 -999 4978 -953
rect 6216 -953 6262 -781
rect 6477 -785 6677 -781
rect 6757 -719 6957 -708
rect 6757 -735 6772 -719
rect 6828 -735 6882 -719
rect 6938 -735 6957 -719
rect 8717 -719 8917 -708
rect 8717 -735 8736 -719
rect 8792 -735 8846 -719
rect 8902 -735 8917 -719
rect 6757 -781 6770 -735
rect 6944 -781 6957 -735
rect 7039 -781 7050 -735
rect 7224 -781 7235 -735
rect 7319 -781 7330 -735
rect 7504 -781 7610 -735
rect 7784 -781 7795 -735
rect 7879 -781 7890 -735
rect 8064 -781 8170 -735
rect 8344 -781 8355 -735
rect 8439 -781 8450 -735
rect 8624 -781 8635 -735
rect 8717 -781 8730 -735
rect 8904 -781 8917 -735
rect 6757 -785 6957 -781
rect 6311 -833 6391 -827
rect 6311 -889 6323 -833
rect 6379 -837 6391 -833
rect 7050 -837 7100 -781
rect 6379 -883 7100 -837
rect 8574 -837 8624 -781
rect 8717 -785 8917 -781
rect 8997 -718 9197 -708
rect 8997 -735 9017 -718
rect 9073 -735 9127 -718
rect 9183 -735 9197 -718
rect 9557 -719 9757 -708
rect 9557 -735 9578 -719
rect 9634 -735 9688 -719
rect 8997 -781 9010 -735
rect 9184 -781 9197 -735
rect 9279 -781 9290 -735
rect 9464 -781 9475 -735
rect 9557 -781 9570 -735
rect 9744 -781 9757 -719
rect 10571 -729 10651 -707
rect 9839 -781 9850 -735
rect 10024 -781 10035 -735
rect 10119 -781 10130 -735
rect 10304 -759 10651 -729
rect 8997 -785 9197 -781
rect 9283 -833 9363 -827
rect 9283 -837 9295 -833
rect 8574 -883 9295 -837
rect 6379 -889 6391 -883
rect 6311 -894 6391 -889
rect 9283 -889 9295 -883
rect 9351 -889 9363 -833
rect 9283 -894 9363 -889
rect 9412 -953 9458 -781
rect 9557 -785 9757 -781
rect 9978 -827 10024 -781
rect 10304 -786 10588 -759
rect 10571 -805 10588 -786
rect 10634 -805 10651 -759
rect 9978 -832 10263 -827
rect 9978 -873 10084 -832
rect 10024 -874 10084 -873
rect 10066 -888 10084 -874
rect 10140 -888 10194 -832
rect 10250 -888 10263 -832
rect 10066 -893 10263 -888
rect 10571 -857 10651 -805
rect 2837 -1055 3037 -1050
rect 3677 -1055 3877 -1050
rect 4095 -1055 4145 -999
rect 5466 -1009 5696 -963
rect 6216 -999 7099 -953
rect 4797 -1055 4997 -1051
rect 1717 -1118 1730 -1055
rect 1904 -1101 1917 -1055
rect 1999 -1101 2010 -1055
rect 2184 -1101 2290 -1055
rect 2464 -1101 2475 -1055
rect 2559 -1101 2570 -1055
rect 2744 -1101 2755 -1055
rect 2837 -1101 2850 -1055
rect 3024 -1101 3037 -1055
rect 1786 -1118 1840 -1101
rect 1896 -1118 1917 -1101
rect 2569 -1102 2619 -1101
rect 1717 -1128 1917 -1118
rect 2837 -1116 2852 -1101
rect 2908 -1116 2962 -1101
rect 3018 -1116 3037 -1101
rect 2837 -1128 3037 -1116
rect 3119 -1101 3130 -1055
rect 3304 -1101 3410 -1055
rect 3584 -1101 3596 -1055
rect 3119 -1116 3135 -1101
rect 3191 -1116 3245 -1101
rect 3301 -1116 3316 -1101
rect 3119 -1121 3316 -1116
rect 3399 -1116 3415 -1101
rect 3471 -1116 3525 -1101
rect 3581 -1116 3596 -1101
rect 3399 -1121 3596 -1116
rect 3677 -1101 3690 -1055
rect 3864 -1101 3877 -1055
rect 3959 -1101 3970 -1055
rect 4144 -1101 4155 -1055
rect 4239 -1101 4250 -1055
rect 4424 -1101 4530 -1055
rect 4704 -1101 4715 -1055
rect 4797 -1101 4810 -1055
rect 3677 -1116 3696 -1101
rect 3752 -1116 3806 -1101
rect 3862 -1116 3877 -1101
rect 4095 -1102 4145 -1101
rect 3677 -1128 3877 -1116
rect 4797 -1118 4818 -1101
rect 4874 -1118 4928 -1101
rect 4984 -1118 4997 -1055
rect 4797 -1128 4997 -1118
rect 5077 -1055 5277 -1050
rect 5498 -1055 5544 -1009
rect 5650 -1055 5696 -1009
rect 5917 -1055 6117 -1050
rect 5077 -1101 5090 -1055
rect 5077 -1117 5098 -1101
rect 5154 -1117 5208 -1101
rect 5264 -1117 5277 -1055
rect 5359 -1101 5370 -1055
rect 5544 -1101 5555 -1055
rect 5639 -1101 5650 -1055
rect 5824 -1101 5835 -1055
rect 5077 -1127 5277 -1117
rect 5917 -1117 5930 -1055
rect 6104 -1101 6117 -1055
rect 5986 -1117 6040 -1101
rect 6096 -1117 6117 -1101
rect 5917 -1127 6117 -1117
rect 6197 -1055 6397 -1051
rect 7049 -1055 7099 -999
rect 8575 -999 9458 -953
rect 10571 -903 10588 -857
rect 10634 -903 10651 -857
rect 10571 -955 10651 -903
rect 7317 -1055 7517 -1050
rect 8157 -1055 8357 -1050
rect 8575 -1055 8625 -999
rect 10571 -1001 10588 -955
rect 10634 -1001 10651 -955
rect 10571 -1047 10651 -1001
rect 9277 -1055 9477 -1051
rect 6197 -1118 6210 -1055
rect 6384 -1101 6397 -1055
rect 6479 -1101 6490 -1055
rect 6664 -1101 6770 -1055
rect 6944 -1101 6955 -1055
rect 7039 -1101 7050 -1055
rect 7224 -1101 7235 -1055
rect 7317 -1101 7330 -1055
rect 7504 -1101 7517 -1055
rect 7599 -1101 7610 -1055
rect 7784 -1101 7890 -1055
rect 8064 -1101 8075 -1055
rect 8157 -1101 8170 -1055
rect 8344 -1101 8357 -1055
rect 8439 -1101 8450 -1055
rect 8624 -1101 8635 -1055
rect 8719 -1101 8730 -1055
rect 8904 -1101 9010 -1055
rect 9184 -1101 9195 -1055
rect 9277 -1101 9290 -1055
rect 6266 -1118 6320 -1101
rect 6376 -1118 6397 -1101
rect 7049 -1102 7099 -1101
rect 6197 -1128 6397 -1118
rect 7317 -1116 7332 -1101
rect 7388 -1116 7442 -1101
rect 7498 -1116 7517 -1101
rect 7317 -1128 7517 -1116
rect 8157 -1116 8176 -1101
rect 8232 -1116 8286 -1101
rect 8342 -1116 8357 -1101
rect 8575 -1102 8625 -1101
rect 8157 -1128 8357 -1116
rect 9277 -1118 9298 -1101
rect 9354 -1118 9408 -1101
rect 9464 -1118 9477 -1055
rect 9277 -1128 9477 -1118
rect 9557 -1055 9757 -1050
rect 10299 -1053 10651 -1047
rect 10299 -1055 10588 -1053
rect 9557 -1101 9570 -1055
rect 9557 -1117 9578 -1101
rect 9634 -1117 9688 -1101
rect 9744 -1117 9757 -1055
rect 9839 -1101 9850 -1055
rect 10024 -1101 10035 -1055
rect 10119 -1101 10130 -1055
rect 10304 -1099 10588 -1055
rect 10634 -1099 10651 -1053
rect 10304 -1101 10651 -1099
rect 9557 -1127 9757 -1117
rect 543 -1197 560 -1151
rect 606 -1197 623 -1151
rect 543 -1249 623 -1197
rect 346 -1265 412 -1249
rect 346 -1321 351 -1265
rect 407 -1321 412 -1265
rect 346 -1375 412 -1321
rect 346 -1431 351 -1375
rect 407 -1431 412 -1375
rect 346 -1446 412 -1431
rect 543 -1295 560 -1249
rect 606 -1295 623 -1249
rect 543 -1347 623 -1295
rect 678 -1254 875 -1249
rect 678 -1310 691 -1254
rect 747 -1310 801 -1254
rect 857 -1261 875 -1254
rect 857 -1310 2123 -1261
rect 678 -1311 2123 -1310
rect 678 -1315 875 -1311
rect 543 -1393 560 -1347
rect 606 -1376 623 -1347
rect 1437 -1367 1637 -1357
rect 606 -1387 930 -1376
rect 1437 -1387 1452 -1367
rect 1508 -1387 1562 -1367
rect 1618 -1387 1637 -1367
rect 606 -1393 890 -1387
rect 543 -1433 890 -1393
rect 1064 -1433 1075 -1387
rect 1159 -1433 1170 -1387
rect 1344 -1433 1355 -1387
rect 1437 -1433 1450 -1387
rect 1624 -1433 1637 -1387
rect 543 -1442 930 -1433
rect 543 -1445 623 -1442
rect 543 -1491 560 -1445
rect 606 -1491 623 -1445
rect 543 -1543 623 -1491
rect 543 -1589 560 -1543
rect 606 -1589 623 -1543
rect 1296 -1517 1344 -1433
rect 1437 -1435 1637 -1433
rect 1717 -1373 1917 -1360
rect 1717 -1387 1732 -1373
rect 1788 -1387 1842 -1373
rect 1898 -1387 1917 -1373
rect 2073 -1387 2123 -1311
rect 2357 -1309 4357 -1259
rect 2357 -1387 2407 -1309
rect 2837 -1366 3037 -1356
rect 2837 -1387 2851 -1366
rect 2907 -1387 2961 -1366
rect 3017 -1387 3037 -1366
rect 1717 -1433 1730 -1387
rect 1904 -1433 1917 -1387
rect 1999 -1433 2010 -1387
rect 2184 -1433 2195 -1387
rect 2279 -1433 2290 -1387
rect 2464 -1433 2475 -1387
rect 2559 -1433 2570 -1387
rect 2744 -1433 2755 -1387
rect 2837 -1433 2850 -1387
rect 3024 -1433 3037 -1387
rect 1717 -1437 1917 -1433
rect 2073 -1434 2123 -1433
rect 2357 -1434 2407 -1433
rect 2570 -1490 2620 -1433
rect 2837 -1436 3037 -1433
rect 3117 -1368 3317 -1360
rect 3117 -1433 3130 -1368
rect 3186 -1387 3240 -1368
rect 3296 -1387 3317 -1368
rect 3304 -1433 3317 -1387
rect 3117 -1437 3317 -1433
rect 3397 -1368 3597 -1360
rect 3397 -1387 3418 -1368
rect 3474 -1387 3528 -1368
rect 3397 -1433 3410 -1387
rect 3584 -1433 3597 -1368
rect 3397 -1437 3597 -1433
rect 3677 -1366 3877 -1356
rect 3677 -1387 3697 -1366
rect 3753 -1387 3807 -1366
rect 3863 -1387 3877 -1366
rect 4307 -1387 4357 -1309
rect 4591 -1311 6603 -1261
rect 4591 -1387 4641 -1311
rect 4797 -1373 4997 -1360
rect 4797 -1387 4816 -1373
rect 4872 -1387 4926 -1373
rect 4982 -1387 4997 -1373
rect 3677 -1433 3690 -1387
rect 3864 -1433 3877 -1387
rect 3959 -1433 3970 -1387
rect 4144 -1433 4155 -1387
rect 4239 -1433 4250 -1387
rect 4424 -1433 4435 -1387
rect 4519 -1433 4530 -1387
rect 4704 -1433 4715 -1387
rect 4797 -1433 4810 -1387
rect 4984 -1433 4997 -1387
rect 3677 -1436 3877 -1433
rect 1296 -1523 1611 -1517
rect 1296 -1579 1433 -1523
rect 1489 -1579 1543 -1523
rect 1599 -1579 1611 -1523
rect 1296 -1583 1611 -1579
rect 1737 -1536 2620 -1490
rect 4094 -1490 4144 -1433
rect 4307 -1434 4357 -1433
rect 4591 -1434 4641 -1433
rect 4797 -1437 4997 -1433
rect 5077 -1367 5277 -1357
rect 5077 -1387 5096 -1367
rect 5152 -1387 5206 -1367
rect 5262 -1387 5277 -1367
rect 5917 -1367 6117 -1357
rect 5917 -1387 5932 -1367
rect 5988 -1387 6042 -1367
rect 6098 -1387 6117 -1367
rect 5077 -1433 5090 -1387
rect 5264 -1433 5277 -1387
rect 5359 -1433 5370 -1387
rect 5544 -1433 5555 -1387
rect 5639 -1433 5650 -1387
rect 5824 -1433 5835 -1387
rect 5917 -1433 5930 -1387
rect 6104 -1433 6117 -1387
rect 5077 -1435 5277 -1433
rect 4094 -1536 4977 -1490
rect 5370 -1517 5418 -1433
rect 543 -1641 623 -1589
rect 543 -1687 560 -1641
rect 606 -1687 623 -1641
rect 915 -1590 1112 -1585
rect 915 -1646 931 -1590
rect 987 -1646 1041 -1590
rect 1097 -1595 1112 -1590
rect 1097 -1641 1216 -1595
rect 1097 -1646 1112 -1641
rect 915 -1651 1112 -1646
rect 543 -1739 623 -1687
rect 1170 -1707 1216 -1641
rect 1437 -1707 1637 -1702
rect 1737 -1707 1783 -1536
rect 1832 -1588 2024 -1585
rect 1832 -1644 1844 -1588
rect 1900 -1644 1954 -1588
rect 2010 -1599 2024 -1588
rect 4690 -1588 4882 -1585
rect 4690 -1599 4704 -1588
rect 2010 -1644 2620 -1599
rect 1832 -1645 2620 -1644
rect 1832 -1647 2024 -1645
rect 1997 -1707 2197 -1703
rect 543 -1785 560 -1739
rect 606 -1785 623 -1739
rect 879 -1753 890 -1707
rect 1064 -1753 1075 -1707
rect 1159 -1753 1170 -1707
rect 1344 -1753 1355 -1707
rect 1437 -1709 1450 -1707
rect 543 -1837 623 -1785
rect 543 -1883 560 -1837
rect 606 -1883 623 -1837
rect 543 -1935 623 -1883
rect 543 -1981 560 -1935
rect 606 -1981 623 -1935
rect 543 -2033 623 -1981
rect 543 -2079 560 -2033
rect 606 -2079 623 -2033
rect 951 -2039 1020 -1753
rect 1170 -2039 1251 -1753
rect 1437 -1765 1449 -1709
rect 1624 -1753 1637 -1707
rect 1719 -1753 1730 -1707
rect 1904 -1753 1915 -1707
rect 1505 -1765 1557 -1753
rect 1613 -1765 1637 -1753
rect 1437 -1779 1637 -1765
rect 1997 -1772 2010 -1707
rect 2184 -1753 2197 -1707
rect 2066 -1772 2120 -1753
rect 2176 -1772 2197 -1753
rect 1997 -1780 2197 -1772
rect 2277 -1707 2477 -1703
rect 2570 -1707 2620 -1645
rect 4094 -1644 4704 -1599
rect 4760 -1644 4814 -1588
rect 4870 -1644 4882 -1588
rect 4094 -1645 4882 -1644
rect 2837 -1707 3037 -1703
rect 3677 -1707 3877 -1703
rect 4094 -1707 4144 -1645
rect 4690 -1647 4882 -1645
rect 4237 -1707 4437 -1703
rect 2277 -1753 2290 -1707
rect 2464 -1753 2477 -1707
rect 2559 -1753 2570 -1707
rect 2744 -1753 2755 -1707
rect 2837 -1710 2850 -1707
rect 2277 -1769 2291 -1753
rect 2347 -1769 2401 -1753
rect 2457 -1769 2477 -1753
rect 2277 -1780 2477 -1769
rect 2837 -1766 2849 -1710
rect 3024 -1753 3037 -1707
rect 3119 -1753 3130 -1707
rect 3304 -1753 3410 -1707
rect 3584 -1753 3595 -1707
rect 3677 -1753 3690 -1707
rect 3864 -1710 3877 -1707
rect 2905 -1766 2959 -1753
rect 3015 -1766 3037 -1753
rect 2837 -1780 3037 -1766
rect 3677 -1766 3699 -1753
rect 3755 -1766 3809 -1753
rect 3865 -1766 3877 -1710
rect 3959 -1753 3970 -1707
rect 4144 -1753 4155 -1707
rect 4237 -1753 4250 -1707
rect 4424 -1753 4437 -1707
rect 3677 -1780 3877 -1766
rect 4237 -1769 4257 -1753
rect 4313 -1769 4367 -1753
rect 4423 -1769 4437 -1753
rect 4237 -1780 4437 -1769
rect 4517 -1707 4717 -1703
rect 4931 -1707 4977 -1536
rect 5101 -1522 5418 -1517
rect 5101 -1578 5113 -1522
rect 5169 -1578 5223 -1522
rect 5279 -1578 5418 -1522
rect 5101 -1583 5418 -1578
rect 5776 -1517 5824 -1433
rect 5917 -1435 6117 -1433
rect 6197 -1373 6397 -1360
rect 6197 -1387 6212 -1373
rect 6268 -1387 6322 -1373
rect 6378 -1387 6397 -1373
rect 6553 -1387 6603 -1311
rect 6837 -1309 8837 -1259
rect 9850 -1261 9908 -1101
rect 10299 -1104 10651 -1101
rect 10571 -1151 10651 -1104
rect 10571 -1197 10588 -1151
rect 10634 -1197 10651 -1151
rect 10571 -1249 10651 -1197
rect 10067 -1254 10264 -1249
rect 10067 -1261 10085 -1254
rect 6837 -1387 6887 -1309
rect 7317 -1366 7517 -1356
rect 7317 -1387 7331 -1366
rect 7387 -1387 7441 -1366
rect 7497 -1387 7517 -1366
rect 6197 -1433 6210 -1387
rect 6384 -1433 6397 -1387
rect 6479 -1433 6490 -1387
rect 6664 -1433 6675 -1387
rect 6759 -1433 6770 -1387
rect 6944 -1433 6955 -1387
rect 7039 -1433 7050 -1387
rect 7224 -1433 7235 -1387
rect 7317 -1433 7330 -1387
rect 7504 -1433 7517 -1387
rect 6197 -1437 6397 -1433
rect 6553 -1434 6603 -1433
rect 6837 -1434 6887 -1433
rect 7050 -1490 7100 -1433
rect 7317 -1436 7517 -1433
rect 7597 -1368 7797 -1360
rect 7597 -1433 7610 -1368
rect 7666 -1387 7720 -1368
rect 7776 -1387 7797 -1368
rect 7784 -1433 7797 -1387
rect 7597 -1437 7797 -1433
rect 7877 -1368 8077 -1360
rect 7877 -1387 7898 -1368
rect 7954 -1387 8008 -1368
rect 7877 -1433 7890 -1387
rect 8064 -1433 8077 -1368
rect 7877 -1437 8077 -1433
rect 8157 -1366 8357 -1356
rect 8157 -1387 8177 -1366
rect 8233 -1387 8287 -1366
rect 8343 -1387 8357 -1366
rect 8787 -1387 8837 -1309
rect 9071 -1310 10085 -1261
rect 10141 -1310 10195 -1254
rect 10251 -1310 10264 -1254
rect 9071 -1311 10264 -1310
rect 9071 -1387 9121 -1311
rect 10067 -1315 10264 -1311
rect 10571 -1295 10588 -1249
rect 10634 -1295 10651 -1249
rect 10571 -1347 10651 -1295
rect 10704 -1158 10767 1158
rect 10813 785 10879 800
rect 10813 729 10818 785
rect 10874 729 10879 785
rect 10813 675 10879 729
rect 10813 619 10818 675
rect 10874 619 10879 675
rect 10813 603 10879 619
rect 10813 -603 10876 603
rect 10942 583 11005 598
rect 10942 527 10947 583
rect 11003 527 11005 583
rect 10942 473 11005 527
rect 10942 417 10947 473
rect 11003 417 11005 473
rect 10942 -417 11005 417
rect 11063 412 11127 427
rect 11063 356 11066 412
rect 11122 356 11127 412
rect 11063 302 11127 356
rect 11063 296 11066 302
rect 11061 246 11066 296
rect 11122 246 11127 302
rect 11061 230 11127 246
rect 11061 -230 11124 230
rect 11061 -246 11127 -230
rect 11061 -296 11066 -246
rect 10942 -473 10947 -417
rect 11003 -473 11005 -417
rect 11063 -302 11066 -296
rect 11122 -302 11127 -246
rect 11063 -356 11127 -302
rect 11063 -412 11066 -356
rect 11122 -412 11127 -356
rect 11063 -427 11127 -412
rect 10942 -527 11005 -473
rect 10942 -583 10947 -527
rect 11003 -583 11005 -527
rect 10942 -598 11005 -583
rect 10813 -619 10879 -603
rect 10813 -675 10818 -619
rect 10874 -675 10879 -619
rect 10813 -729 10879 -675
rect 10813 -785 10818 -729
rect 10874 -785 10879 -729
rect 10813 -800 10879 -785
rect 10704 -1214 10709 -1158
rect 10765 -1214 10767 -1158
rect 10704 -1268 10767 -1214
rect 10704 -1324 10709 -1268
rect 10765 -1324 10767 -1268
rect 10704 -1339 10767 -1324
rect 9277 -1373 9477 -1360
rect 9277 -1387 9296 -1373
rect 9352 -1387 9406 -1373
rect 9462 -1387 9477 -1373
rect 8157 -1433 8170 -1387
rect 8344 -1433 8357 -1387
rect 8439 -1433 8450 -1387
rect 8624 -1433 8635 -1387
rect 8719 -1433 8730 -1387
rect 8904 -1433 8915 -1387
rect 8999 -1433 9010 -1387
rect 9184 -1433 9195 -1387
rect 9277 -1433 9290 -1387
rect 9464 -1433 9477 -1387
rect 8157 -1436 8357 -1433
rect 5776 -1523 6091 -1517
rect 5776 -1579 5913 -1523
rect 5969 -1579 6023 -1523
rect 6079 -1579 6091 -1523
rect 5776 -1583 6091 -1579
rect 6217 -1536 7100 -1490
rect 8574 -1490 8624 -1433
rect 8787 -1434 8837 -1433
rect 9071 -1434 9121 -1433
rect 9277 -1437 9477 -1433
rect 9557 -1367 9757 -1357
rect 9557 -1387 9576 -1367
rect 9632 -1387 9686 -1367
rect 9742 -1387 9757 -1367
rect 10571 -1385 10588 -1347
rect 10300 -1387 10588 -1385
rect 9557 -1433 9570 -1387
rect 9744 -1433 9757 -1387
rect 9839 -1433 9850 -1387
rect 10024 -1433 10035 -1387
rect 10119 -1433 10130 -1387
rect 10304 -1393 10588 -1387
rect 10634 -1393 10651 -1347
rect 10304 -1433 10651 -1393
rect 9557 -1435 9757 -1433
rect 8574 -1536 9457 -1490
rect 9850 -1517 9898 -1433
rect 10300 -1442 10651 -1433
rect 5466 -1661 5696 -1615
rect 5077 -1707 5277 -1702
rect 5498 -1707 5544 -1661
rect 5650 -1707 5696 -1661
rect 5917 -1707 6117 -1702
rect 6217 -1707 6263 -1536
rect 6312 -1588 6504 -1585
rect 6312 -1644 6324 -1588
rect 6380 -1644 6434 -1588
rect 6490 -1599 6504 -1588
rect 9170 -1588 9362 -1585
rect 9170 -1599 9184 -1588
rect 6490 -1644 7100 -1599
rect 6312 -1645 7100 -1644
rect 6312 -1647 6504 -1645
rect 6477 -1707 6677 -1703
rect 4517 -1753 4530 -1707
rect 4517 -1772 4538 -1753
rect 4594 -1772 4648 -1753
rect 4704 -1772 4717 -1707
rect 4799 -1753 4810 -1707
rect 4984 -1753 4995 -1707
rect 5077 -1753 5090 -1707
rect 5264 -1709 5277 -1707
rect 4517 -1780 4717 -1772
rect 5077 -1765 5101 -1753
rect 5157 -1765 5209 -1753
rect 5265 -1765 5277 -1709
rect 5359 -1753 5370 -1707
rect 5544 -1753 5555 -1707
rect 5639 -1753 5650 -1707
rect 5824 -1753 5835 -1707
rect 5917 -1709 5930 -1707
rect 5077 -1779 5277 -1765
rect 5917 -1765 5929 -1709
rect 6104 -1753 6117 -1707
rect 6199 -1753 6210 -1707
rect 6384 -1753 6395 -1707
rect 5985 -1765 6037 -1753
rect 6093 -1765 6117 -1753
rect 5917 -1779 6117 -1765
rect 6477 -1772 6490 -1707
rect 6664 -1753 6677 -1707
rect 6546 -1772 6600 -1753
rect 6656 -1772 6677 -1753
rect 6477 -1780 6677 -1772
rect 6757 -1707 6957 -1703
rect 7050 -1707 7100 -1645
rect 8574 -1644 9184 -1599
rect 9240 -1644 9294 -1588
rect 9350 -1644 9362 -1588
rect 8574 -1645 9362 -1644
rect 7317 -1707 7517 -1703
rect 8157 -1707 8357 -1703
rect 8574 -1707 8624 -1645
rect 9170 -1647 9362 -1645
rect 8717 -1707 8917 -1703
rect 6757 -1753 6770 -1707
rect 6944 -1753 6957 -1707
rect 7039 -1753 7050 -1707
rect 7224 -1753 7235 -1707
rect 7317 -1710 7330 -1707
rect 6757 -1769 6771 -1753
rect 6827 -1769 6881 -1753
rect 6937 -1769 6957 -1753
rect 6757 -1780 6957 -1769
rect 7317 -1766 7329 -1710
rect 7504 -1753 7517 -1707
rect 7599 -1753 7610 -1707
rect 7784 -1753 7890 -1707
rect 8064 -1753 8075 -1707
rect 8157 -1753 8170 -1707
rect 8344 -1710 8357 -1707
rect 7385 -1766 7439 -1753
rect 7495 -1766 7517 -1753
rect 7317 -1780 7517 -1766
rect 8157 -1766 8179 -1753
rect 8235 -1766 8289 -1753
rect 8345 -1766 8357 -1710
rect 8439 -1753 8450 -1707
rect 8624 -1753 8635 -1707
rect 8717 -1753 8730 -1707
rect 8904 -1753 8917 -1707
rect 8157 -1780 8357 -1766
rect 8717 -1769 8737 -1753
rect 8793 -1769 8847 -1753
rect 8903 -1769 8917 -1753
rect 8717 -1780 8917 -1769
rect 8997 -1707 9197 -1703
rect 9411 -1707 9457 -1536
rect 9581 -1522 9898 -1517
rect 9581 -1578 9593 -1522
rect 9649 -1578 9703 -1522
rect 9759 -1578 9898 -1522
rect 9581 -1583 9898 -1578
rect 10571 -1445 10651 -1442
rect 10571 -1491 10588 -1445
rect 10634 -1491 10651 -1445
rect 10571 -1543 10651 -1491
rect 10282 -1590 10479 -1585
rect 10282 -1595 10295 -1590
rect 9978 -1641 10295 -1595
rect 9557 -1707 9757 -1702
rect 9978 -1707 10024 -1641
rect 10282 -1646 10295 -1641
rect 10353 -1646 10405 -1590
rect 10463 -1646 10479 -1590
rect 10282 -1651 10479 -1646
rect 10571 -1589 10588 -1543
rect 10634 -1589 10651 -1543
rect 10571 -1641 10651 -1589
rect 10571 -1687 10588 -1641
rect 10634 -1687 10651 -1641
rect 8997 -1753 9010 -1707
rect 8997 -1772 9018 -1753
rect 9074 -1772 9128 -1753
rect 9184 -1772 9197 -1707
rect 9279 -1753 9290 -1707
rect 9464 -1753 9475 -1707
rect 9557 -1753 9570 -1707
rect 9744 -1709 9757 -1707
rect 8997 -1780 9197 -1772
rect 9557 -1765 9581 -1753
rect 9637 -1765 9689 -1753
rect 9745 -1765 9757 -1709
rect 9839 -1753 9850 -1707
rect 10024 -1753 10035 -1707
rect 10119 -1753 10130 -1707
rect 10304 -1708 10315 -1707
rect 10571 -1708 10651 -1687
rect 10304 -1739 10651 -1708
rect 10304 -1753 10588 -1739
rect 10302 -1765 10588 -1753
rect 9557 -1779 9757 -1765
rect 10571 -1785 10588 -1765
rect 10634 -1785 10651 -1739
rect 1774 -1887 4940 -1830
rect 1774 -2039 1831 -1887
rect 2634 -1983 4080 -1933
rect 2277 -2024 2477 -2012
rect 2277 -2039 2291 -2024
rect 2347 -2039 2401 -2024
rect 2457 -2039 2477 -2024
rect 2634 -2039 2684 -1983
rect 4030 -2039 4080 -1983
rect 4237 -2024 4437 -2012
rect 4237 -2039 4257 -2024
rect 4313 -2039 4367 -2024
rect 4423 -2039 4437 -2024
rect 4883 -2039 4940 -1887
rect 6254 -1887 9420 -1830
rect 6254 -2039 6311 -1887
rect 7114 -1983 8560 -1933
rect 6757 -2024 6957 -2012
rect 6757 -2039 6771 -2024
rect 6827 -2039 6881 -2024
rect 6937 -2039 6957 -2024
rect 7114 -2039 7164 -1983
rect 8510 -2039 8560 -1983
rect 8717 -2024 8917 -2012
rect 8717 -2039 8737 -2024
rect 8793 -2039 8847 -2024
rect 8903 -2039 8917 -2024
rect 9363 -2039 9420 -1887
rect 10571 -1837 10651 -1785
rect 10571 -1883 10588 -1837
rect 10634 -1883 10651 -1837
rect 10571 -1935 10651 -1883
rect 10571 -1981 10588 -1935
rect 10634 -1981 10651 -1935
rect 10571 -2033 10651 -1981
rect 10571 -2034 10588 -2033
rect 10302 -2039 10588 -2034
rect 543 -2131 623 -2079
rect 879 -2085 890 -2039
rect 1064 -2085 1075 -2039
rect 1159 -2085 1170 -2039
rect 1344 -2085 1450 -2039
rect 1624 -2085 1646 -2039
rect 1719 -2085 1730 -2039
rect 1904 -2085 1915 -2039
rect 1999 -2085 2010 -2039
rect 2184 -2085 2195 -2039
rect 2277 -2085 2290 -2039
rect 2464 -2085 2477 -2039
rect 2559 -2085 2570 -2039
rect 2744 -2085 2755 -2039
rect 2839 -2085 2850 -2039
rect 3024 -2085 3130 -2039
rect 3304 -2085 3315 -2039
rect 3399 -2085 3410 -2039
rect 3584 -2085 3690 -2039
rect 3864 -2085 3875 -2039
rect 3959 -2085 3970 -2039
rect 4144 -2085 4155 -2039
rect 4237 -2085 4250 -2039
rect 4424 -2085 4437 -2039
rect 4519 -2085 4530 -2039
rect 4704 -2085 4715 -2039
rect 4799 -2085 4810 -2039
rect 4984 -2085 4995 -2039
rect 5068 -2085 5090 -2039
rect 5264 -2085 5370 -2039
rect 5544 -2085 5555 -2039
rect 5639 -2085 5650 -2039
rect 5824 -2085 5930 -2039
rect 6104 -2085 6126 -2039
rect 6199 -2085 6210 -2039
rect 6384 -2085 6395 -2039
rect 6479 -2085 6490 -2039
rect 6664 -2085 6675 -2039
rect 6757 -2085 6770 -2039
rect 6944 -2085 6957 -2039
rect 7039 -2085 7050 -2039
rect 7224 -2085 7235 -2039
rect 7319 -2085 7330 -2039
rect 7504 -2085 7610 -2039
rect 7784 -2085 7795 -2039
rect 7879 -2085 7890 -2039
rect 8064 -2085 8170 -2039
rect 8344 -2085 8355 -2039
rect 8439 -2085 8450 -2039
rect 8624 -2085 8635 -2039
rect 8717 -2085 8730 -2039
rect 8904 -2085 8917 -2039
rect 8999 -2085 9010 -2039
rect 9184 -2085 9195 -2039
rect 9279 -2085 9290 -2039
rect 9464 -2085 9475 -2039
rect 9548 -2085 9570 -2039
rect 9744 -2085 9850 -2039
rect 10024 -2085 10035 -2039
rect 10119 -2085 10130 -2039
rect 10304 -2079 10588 -2039
rect 10634 -2079 10651 -2033
rect 10304 -2085 10651 -2079
rect 543 -2177 560 -2131
rect 606 -2177 623 -2131
rect 543 -2229 623 -2177
rect 543 -2275 560 -2229
rect 606 -2275 623 -2229
rect 543 -2314 623 -2275
rect 951 -2314 1020 -2085
rect 2138 -2136 2184 -2085
rect 2277 -2089 2477 -2085
rect 2634 -2087 2684 -2085
rect 4030 -2087 4080 -2085
rect 4237 -2089 4437 -2085
rect 3036 -2135 3226 -2131
rect 3036 -2136 3048 -2135
rect 2138 -2182 3048 -2136
rect 3036 -2191 3048 -2182
rect 3104 -2191 3158 -2135
rect 3214 -2191 3226 -2135
rect 3036 -2195 3226 -2191
rect 3488 -2135 3678 -2131
rect 3488 -2191 3500 -2135
rect 3556 -2191 3610 -2135
rect 3666 -2136 3678 -2135
rect 4530 -2136 4576 -2085
rect 3666 -2182 4576 -2136
rect 6618 -2136 6664 -2085
rect 6757 -2089 6957 -2085
rect 7114 -2087 7164 -2085
rect 8510 -2087 8560 -2085
rect 8717 -2089 8917 -2085
rect 7516 -2135 7706 -2131
rect 7516 -2136 7528 -2135
rect 6618 -2182 7528 -2136
rect 3666 -2191 3678 -2182
rect 3488 -2195 3678 -2191
rect 7516 -2191 7528 -2182
rect 7584 -2191 7638 -2135
rect 7694 -2191 7706 -2135
rect 7516 -2195 7706 -2191
rect 7968 -2135 8158 -2131
rect 7968 -2191 7980 -2135
rect 8036 -2191 8090 -2135
rect 8146 -2136 8158 -2135
rect 9010 -2136 9056 -2085
rect 10302 -2091 10651 -2085
rect 8146 -2182 9056 -2136
rect 10571 -2131 10651 -2091
rect 10571 -2177 10588 -2131
rect 10634 -2177 10651 -2131
rect 8146 -2191 8158 -2182
rect 7968 -2195 8158 -2191
rect 10571 -2229 10651 -2177
rect 10571 -2275 10588 -2229
rect 10634 -2275 10651 -2229
rect 10571 -2314 10651 -2275
rect 543 -2327 10651 -2314
rect 543 -2377 560 -2327
rect 606 -2331 10588 -2327
rect 606 -2377 658 -2331
rect 704 -2377 756 -2331
rect 802 -2377 854 -2331
rect 900 -2377 952 -2331
rect 998 -2377 1050 -2331
rect 1096 -2377 1148 -2331
rect 1194 -2377 1246 -2331
rect 1292 -2377 1344 -2331
rect 1390 -2377 1442 -2331
rect 1488 -2377 1540 -2331
rect 1586 -2377 1638 -2331
rect 1684 -2377 1736 -2331
rect 1782 -2377 1834 -2331
rect 1880 -2377 1932 -2331
rect 1978 -2377 2030 -2331
rect 2076 -2377 2128 -2331
rect 2174 -2377 2226 -2331
rect 2272 -2377 2324 -2331
rect 2370 -2377 2422 -2331
rect 2468 -2377 2520 -2331
rect 2566 -2377 2618 -2331
rect 2664 -2377 2716 -2331
rect 2762 -2377 2814 -2331
rect 2860 -2377 2912 -2331
rect 2958 -2377 3010 -2331
rect 3056 -2377 3108 -2331
rect 3154 -2377 3206 -2331
rect 3252 -2377 3304 -2331
rect 3350 -2377 3402 -2331
rect 3448 -2377 3500 -2331
rect 3546 -2377 3598 -2331
rect 3644 -2377 3696 -2331
rect 3742 -2377 3794 -2331
rect 3840 -2377 3892 -2331
rect 3938 -2377 3990 -2331
rect 4036 -2377 4088 -2331
rect 4134 -2377 4186 -2331
rect 4232 -2377 4284 -2331
rect 4330 -2377 4382 -2331
rect 4428 -2377 4480 -2331
rect 4526 -2377 4578 -2331
rect 4624 -2377 4676 -2331
rect 4722 -2377 4774 -2331
rect 4820 -2377 4872 -2331
rect 4918 -2377 4970 -2331
rect 5016 -2377 5068 -2331
rect 5114 -2377 5166 -2331
rect 5212 -2377 5264 -2331
rect 5310 -2377 5362 -2331
rect 5408 -2377 5460 -2331
rect 5506 -2377 5558 -2331
rect 5604 -2377 5656 -2331
rect 5702 -2377 5754 -2331
rect 5800 -2377 5852 -2331
rect 5898 -2377 5950 -2331
rect 5996 -2377 6048 -2331
rect 6094 -2377 6146 -2331
rect 6192 -2377 6244 -2331
rect 6290 -2377 6342 -2331
rect 6388 -2377 6440 -2331
rect 6486 -2377 6538 -2331
rect 6584 -2377 6636 -2331
rect 6682 -2377 6734 -2331
rect 6780 -2377 6832 -2331
rect 6878 -2377 6930 -2331
rect 6976 -2377 7028 -2331
rect 7074 -2377 7126 -2331
rect 7172 -2377 7224 -2331
rect 7270 -2377 7322 -2331
rect 7368 -2377 7420 -2331
rect 7466 -2377 7518 -2331
rect 7564 -2377 7616 -2331
rect 7662 -2377 7714 -2331
rect 7760 -2377 7812 -2331
rect 7858 -2377 7910 -2331
rect 7956 -2377 8008 -2331
rect 8054 -2377 8106 -2331
rect 8152 -2377 8204 -2331
rect 8250 -2377 8302 -2331
rect 8348 -2377 8400 -2331
rect 8446 -2377 8498 -2331
rect 8544 -2377 8596 -2331
rect 8642 -2377 8694 -2331
rect 8740 -2377 8792 -2331
rect 8838 -2377 8890 -2331
rect 8936 -2377 8988 -2331
rect 9034 -2377 9086 -2331
rect 9132 -2377 9184 -2331
rect 9230 -2377 9282 -2331
rect 9328 -2377 9380 -2331
rect 9426 -2377 9478 -2331
rect 9524 -2377 9576 -2331
rect 9622 -2377 9674 -2331
rect 9720 -2377 9772 -2331
rect 9818 -2377 9870 -2331
rect 9916 -2377 9968 -2331
rect 10014 -2377 10066 -2331
rect 10112 -2377 10164 -2331
rect 10210 -2377 10262 -2331
rect 10308 -2377 10360 -2331
rect 10406 -2377 10458 -2331
rect 10504 -2377 10588 -2331
rect 10634 -2377 10651 -2327
rect 543 -2394 10651 -2377
<< via1 >>
rect 3048 2135 3104 2191
rect 3158 2135 3214 2191
rect 3500 2135 3556 2191
rect 3610 2135 3666 2191
rect 7528 2135 7584 2191
rect 7638 2135 7694 2191
rect 7980 2135 8036 2191
rect 8090 2135 8146 2191
rect 2291 2039 2347 2080
rect 2401 2039 2457 2080
rect 4257 2039 4313 2080
rect 4367 2039 4423 2080
rect 6771 2039 6827 2080
rect 6881 2039 6937 2080
rect 8737 2039 8793 2080
rect 8847 2039 8903 2080
rect 2291 2024 2347 2039
rect 2401 2024 2457 2039
rect 4257 2024 4313 2039
rect 4367 2024 4423 2039
rect 6771 2024 6827 2039
rect 6881 2024 6937 2039
rect 8737 2024 8793 2039
rect 8847 2024 8903 2039
rect 1449 1753 1505 1765
rect 1557 1753 1613 1765
rect 1449 1709 1450 1753
rect 1450 1709 1505 1753
rect 1557 1709 1613 1753
rect 2010 1753 2066 1772
rect 2120 1753 2176 1772
rect 2010 1716 2066 1753
rect 2120 1716 2176 1753
rect 931 1590 987 1646
rect 1041 1590 1097 1646
rect 351 1375 407 1431
rect 351 1265 407 1321
rect 1433 1523 1489 1579
rect 1543 1523 1599 1579
rect 2291 1753 2347 1769
rect 2401 1753 2457 1769
rect 2291 1713 2347 1753
rect 2401 1713 2457 1753
rect 2849 1753 2905 1766
rect 2959 1753 3015 1766
rect 3699 1753 3755 1766
rect 3809 1753 3865 1766
rect 2849 1710 2850 1753
rect 2850 1710 2905 1753
rect 2959 1710 3015 1753
rect 3699 1710 3755 1753
rect 3809 1710 3864 1753
rect 3864 1710 3865 1753
rect 4257 1753 4313 1769
rect 4367 1753 4423 1769
rect 4257 1713 4313 1753
rect 4367 1713 4423 1753
rect 1844 1588 1900 1644
rect 1954 1588 2010 1644
rect 4538 1753 4594 1772
rect 4648 1753 4704 1772
rect 4538 1716 4594 1753
rect 4648 1716 4704 1753
rect 5101 1753 5157 1765
rect 5209 1753 5265 1765
rect 5101 1709 5157 1753
rect 5209 1709 5264 1753
rect 5264 1709 5265 1753
rect 5929 1753 5985 1765
rect 6037 1753 6093 1765
rect 5929 1709 5930 1753
rect 5930 1709 5985 1753
rect 6037 1709 6093 1753
rect 6490 1753 6546 1772
rect 6600 1753 6656 1772
rect 6490 1716 6546 1753
rect 6600 1716 6656 1753
rect 4704 1588 4760 1644
rect 4814 1588 4870 1644
rect 1452 1387 1508 1423
rect 1562 1387 1618 1423
rect 1452 1367 1508 1387
rect 1562 1367 1618 1387
rect 5113 1522 5169 1578
rect 5223 1522 5279 1578
rect 1732 1387 1788 1429
rect 1842 1387 1898 1429
rect 2851 1387 2907 1422
rect 2961 1387 3017 1422
rect 1732 1373 1788 1387
rect 1842 1373 1898 1387
rect 691 1254 747 1310
rect 801 1254 857 1310
rect 2851 1366 2907 1387
rect 2961 1366 3017 1387
rect 3130 1387 3186 1424
rect 3240 1387 3296 1424
rect 3130 1368 3186 1387
rect 3240 1368 3296 1387
rect 3418 1387 3474 1424
rect 3528 1387 3584 1424
rect 3418 1368 3474 1387
rect 3528 1368 3584 1387
rect 3697 1387 3753 1422
rect 3807 1387 3863 1422
rect 4816 1387 4872 1429
rect 4926 1387 4982 1429
rect 3697 1366 3753 1387
rect 3807 1366 3863 1387
rect 4816 1373 4872 1387
rect 4926 1373 4982 1387
rect 5913 1523 5969 1579
rect 6023 1523 6079 1579
rect 6771 1753 6827 1769
rect 6881 1753 6937 1769
rect 6771 1713 6827 1753
rect 6881 1713 6937 1753
rect 7329 1753 7385 1766
rect 7439 1753 7495 1766
rect 8179 1753 8235 1766
rect 8289 1753 8345 1766
rect 7329 1710 7330 1753
rect 7330 1710 7385 1753
rect 7439 1710 7495 1753
rect 8179 1710 8235 1753
rect 8289 1710 8344 1753
rect 8344 1710 8345 1753
rect 8737 1753 8793 1769
rect 8847 1753 8903 1769
rect 8737 1713 8793 1753
rect 8847 1713 8903 1753
rect 6324 1588 6380 1644
rect 6434 1588 6490 1644
rect 9018 1753 9074 1772
rect 9128 1753 9184 1772
rect 9018 1716 9074 1753
rect 9128 1716 9184 1753
rect 9581 1753 9637 1765
rect 9689 1753 9745 1765
rect 9581 1709 9637 1753
rect 9689 1709 9744 1753
rect 9744 1709 9745 1753
rect 9184 1588 9240 1644
rect 9294 1588 9350 1644
rect 10295 1590 10353 1646
rect 10405 1590 10463 1646
rect 5096 1387 5152 1423
rect 5206 1387 5262 1423
rect 5932 1387 5988 1423
rect 6042 1387 6098 1423
rect 5096 1367 5152 1387
rect 5206 1367 5262 1387
rect 5932 1367 5988 1387
rect 6042 1367 6098 1387
rect 9593 1522 9649 1578
rect 9703 1522 9759 1578
rect 6212 1387 6268 1429
rect 6322 1387 6378 1429
rect 7331 1387 7387 1422
rect 7441 1387 7497 1422
rect 6212 1373 6268 1387
rect 6322 1373 6378 1387
rect 7331 1366 7387 1387
rect 7441 1366 7497 1387
rect 7610 1387 7666 1424
rect 7720 1387 7776 1424
rect 7610 1368 7666 1387
rect 7720 1368 7776 1387
rect 7898 1387 7954 1424
rect 8008 1387 8064 1424
rect 7898 1368 7954 1387
rect 8008 1368 8064 1387
rect 8177 1387 8233 1422
rect 8287 1387 8343 1422
rect 9296 1387 9352 1429
rect 9406 1387 9462 1429
rect 8177 1366 8233 1387
rect 8287 1366 8343 1387
rect 9296 1373 9352 1387
rect 9406 1373 9462 1387
rect 9576 1387 9632 1423
rect 9686 1387 9742 1423
rect 9576 1367 9632 1387
rect 9686 1367 9742 1387
rect 241 1070 297 1126
rect 119 948 175 1004
rect 119 838 175 894
rect 241 960 297 1016
rect 5 356 61 412
rect 5 246 61 302
rect 5 -302 61 -246
rect 5 -412 61 -356
rect 119 -894 175 -838
rect 119 -1004 175 -948
rect 241 -1016 297 -960
rect 241 -1126 297 -1070
rect 1450 1101 1506 1117
rect 1560 1101 1616 1117
rect 1450 1061 1506 1101
rect 1560 1061 1616 1101
rect 682 949 738 1005
rect 792 949 848 1005
rect 1730 1101 1786 1118
rect 1840 1101 1896 1118
rect 2852 1101 2908 1116
rect 2962 1101 3018 1116
rect 1730 1062 1786 1101
rect 1840 1062 1896 1101
rect 2852 1060 2908 1101
rect 2962 1060 3018 1101
rect 3135 1101 3191 1116
rect 3245 1101 3301 1116
rect 3415 1101 3471 1116
rect 3525 1101 3581 1116
rect 3135 1060 3191 1101
rect 3245 1060 3301 1101
rect 3415 1060 3471 1101
rect 3525 1060 3581 1101
rect 3696 1101 3752 1116
rect 3806 1101 3862 1116
rect 4818 1101 4874 1118
rect 4928 1101 4984 1118
rect 3696 1060 3752 1101
rect 3806 1060 3862 1101
rect 4818 1062 4874 1101
rect 4928 1062 4984 1101
rect 5098 1101 5154 1117
rect 5208 1101 5264 1117
rect 5098 1061 5154 1101
rect 5208 1061 5264 1101
rect 5930 1101 5986 1117
rect 6040 1101 6096 1117
rect 5930 1061 5986 1101
rect 6040 1061 6096 1101
rect 6210 1101 6266 1118
rect 6320 1101 6376 1118
rect 7332 1101 7388 1116
rect 7442 1101 7498 1116
rect 8176 1101 8232 1116
rect 8286 1101 8342 1116
rect 9298 1101 9354 1118
rect 9408 1101 9464 1118
rect 6210 1062 6266 1101
rect 6320 1062 6376 1101
rect 7332 1060 7388 1101
rect 7442 1060 7498 1101
rect 8176 1060 8232 1101
rect 8286 1060 8342 1101
rect 9298 1062 9354 1101
rect 9408 1062 9464 1101
rect 948 832 1004 888
rect 1058 832 1114 888
rect 1843 833 1899 889
rect 1450 735 1506 775
rect 1560 735 1616 775
rect 2011 735 2067 774
rect 2121 735 2177 774
rect 1450 719 1506 735
rect 1560 719 1616 735
rect 2011 718 2067 735
rect 2121 718 2177 735
rect 4815 833 4871 889
rect 2292 735 2348 775
rect 2402 735 2458 775
rect 4256 735 4312 775
rect 4366 735 4422 775
rect 2292 719 2348 735
rect 2402 719 2458 735
rect 4256 719 4312 735
rect 4366 719 4422 735
rect 9578 1101 9634 1117
rect 9688 1101 9744 1117
rect 9578 1061 9634 1101
rect 9688 1061 9744 1101
rect 10085 1254 10141 1310
rect 10195 1254 10251 1310
rect 6323 833 6379 889
rect 4537 735 4593 774
rect 4647 735 4703 774
rect 5098 735 5154 775
rect 5208 735 5264 775
rect 4537 718 4593 735
rect 4647 718 4703 735
rect 5098 719 5154 735
rect 5208 719 5264 735
rect 5930 735 5986 775
rect 6040 735 6096 775
rect 6491 735 6547 774
rect 6601 735 6657 774
rect 5930 719 5986 735
rect 6040 719 6096 735
rect 6491 718 6547 735
rect 6601 718 6657 735
rect 9295 833 9351 889
rect 6772 735 6828 775
rect 6882 735 6938 775
rect 8736 735 8792 775
rect 8846 735 8902 775
rect 6772 719 6828 735
rect 6882 719 6938 735
rect 8736 719 8792 735
rect 8846 719 8902 735
rect 10084 832 10140 888
rect 10194 832 10250 888
rect 9017 735 9073 774
rect 9127 735 9183 774
rect 9578 735 9634 775
rect 9688 735 9744 775
rect 9017 718 9073 735
rect 9127 718 9183 735
rect 9578 719 9634 735
rect 9688 719 9744 735
rect 683 608 739 664
rect 793 608 849 664
rect 1452 449 1508 472
rect 1562 449 1618 472
rect 1452 416 1508 449
rect 1562 416 1618 449
rect 2010 449 2066 474
rect 2120 449 2176 474
rect 2010 418 2066 449
rect 2120 418 2176 449
rect 2849 449 2905 461
rect 2959 449 3015 461
rect 3699 449 3755 461
rect 3809 449 3865 461
rect 2849 405 2850 449
rect 2850 405 2905 449
rect 2959 405 3015 449
rect 3699 405 3755 449
rect 3809 405 3864 449
rect 3864 405 3865 449
rect 7329 449 7385 461
rect 7439 449 7495 461
rect 8179 449 8235 461
rect 8289 449 8345 461
rect 7329 405 7330 449
rect 7330 405 7385 449
rect 7439 405 7495 449
rect 8179 405 8235 449
rect 8289 405 8344 449
rect 8344 405 8345 449
rect 10333 608 10389 664
rect 10443 608 10499 664
rect 10083 505 10139 561
rect 10193 505 10249 561
rect 687 235 743 291
rect 797 235 853 291
rect 10313 235 10369 291
rect 10423 235 10479 291
rect 10709 1268 10765 1324
rect 10709 1158 10765 1214
rect 687 -291 743 -235
rect 797 -291 853 -235
rect 10313 -291 10369 -235
rect 10423 -291 10479 -235
rect 1452 -449 1508 -416
rect 1562 -449 1618 -416
rect 1452 -472 1508 -449
rect 1562 -472 1618 -449
rect 2010 -449 2066 -418
rect 2120 -449 2176 -418
rect 2010 -474 2066 -449
rect 2120 -474 2176 -449
rect 683 -664 739 -608
rect 793 -664 849 -608
rect 2849 -449 2850 -405
rect 2850 -449 2905 -405
rect 2959 -449 3015 -405
rect 3699 -449 3755 -405
rect 3809 -449 3864 -405
rect 3864 -449 3865 -405
rect 2849 -461 2905 -449
rect 2959 -461 3015 -449
rect 3699 -461 3755 -449
rect 3809 -461 3865 -449
rect 7329 -449 7330 -405
rect 7330 -449 7385 -405
rect 7439 -449 7495 -405
rect 8179 -449 8235 -405
rect 8289 -449 8344 -405
rect 8344 -449 8345 -405
rect 7329 -461 7385 -449
rect 7439 -461 7495 -449
rect 8179 -461 8235 -449
rect 8289 -461 8345 -449
rect 10083 -561 10139 -505
rect 10193 -561 10249 -505
rect 10333 -664 10389 -608
rect 10443 -664 10499 -608
rect 1450 -735 1506 -719
rect 1560 -735 1616 -719
rect 2011 -735 2067 -718
rect 2121 -735 2177 -718
rect 1450 -775 1506 -735
rect 1560 -775 1616 -735
rect 2011 -774 2067 -735
rect 2121 -774 2177 -735
rect 948 -888 1004 -832
rect 1058 -888 1114 -832
rect 682 -1005 738 -949
rect 792 -1005 848 -949
rect 2292 -735 2348 -719
rect 2402 -735 2458 -719
rect 4256 -735 4312 -719
rect 4366 -735 4422 -719
rect 2292 -775 2348 -735
rect 2402 -775 2458 -735
rect 4256 -775 4312 -735
rect 4366 -775 4422 -735
rect 1843 -889 1899 -833
rect 4537 -735 4593 -718
rect 4647 -735 4703 -718
rect 5098 -735 5154 -719
rect 5208 -735 5264 -719
rect 4537 -774 4593 -735
rect 4647 -774 4703 -735
rect 5098 -775 5154 -735
rect 5208 -775 5264 -735
rect 5930 -735 5986 -719
rect 6040 -735 6096 -719
rect 6491 -735 6547 -718
rect 6601 -735 6657 -718
rect 5930 -775 5986 -735
rect 6040 -775 6096 -735
rect 6491 -774 6547 -735
rect 6601 -774 6657 -735
rect 4815 -889 4871 -833
rect 1450 -1101 1506 -1061
rect 1560 -1101 1616 -1061
rect 1450 -1117 1506 -1101
rect 1560 -1117 1616 -1101
rect 6772 -735 6828 -719
rect 6882 -735 6938 -719
rect 8736 -735 8792 -719
rect 8846 -735 8902 -719
rect 6772 -775 6828 -735
rect 6882 -775 6938 -735
rect 8736 -775 8792 -735
rect 8846 -775 8902 -735
rect 6323 -889 6379 -833
rect 9017 -735 9073 -718
rect 9127 -735 9183 -718
rect 9578 -735 9634 -719
rect 9688 -735 9744 -719
rect 9017 -774 9073 -735
rect 9127 -774 9183 -735
rect 9578 -775 9634 -735
rect 9688 -775 9744 -735
rect 9295 -889 9351 -833
rect 10084 -888 10140 -832
rect 10194 -888 10250 -832
rect 1730 -1101 1786 -1062
rect 1840 -1101 1896 -1062
rect 2852 -1101 2908 -1060
rect 2962 -1101 3018 -1060
rect 1730 -1118 1786 -1101
rect 1840 -1118 1896 -1101
rect 2852 -1116 2908 -1101
rect 2962 -1116 3018 -1101
rect 3135 -1101 3191 -1060
rect 3245 -1101 3301 -1060
rect 3415 -1101 3471 -1060
rect 3525 -1101 3581 -1060
rect 3135 -1116 3191 -1101
rect 3245 -1116 3301 -1101
rect 3415 -1116 3471 -1101
rect 3525 -1116 3581 -1101
rect 3696 -1101 3752 -1060
rect 3806 -1101 3862 -1060
rect 4818 -1101 4874 -1062
rect 4928 -1101 4984 -1062
rect 3696 -1116 3752 -1101
rect 3806 -1116 3862 -1101
rect 4818 -1118 4874 -1101
rect 4928 -1118 4984 -1101
rect 5098 -1101 5154 -1061
rect 5208 -1101 5264 -1061
rect 5098 -1117 5154 -1101
rect 5208 -1117 5264 -1101
rect 5930 -1101 5986 -1061
rect 6040 -1101 6096 -1061
rect 5930 -1117 5986 -1101
rect 6040 -1117 6096 -1101
rect 6210 -1101 6266 -1062
rect 6320 -1101 6376 -1062
rect 7332 -1101 7388 -1060
rect 7442 -1101 7498 -1060
rect 8176 -1101 8232 -1060
rect 8286 -1101 8342 -1060
rect 9298 -1101 9354 -1062
rect 9408 -1101 9464 -1062
rect 6210 -1118 6266 -1101
rect 6320 -1118 6376 -1101
rect 7332 -1116 7388 -1101
rect 7442 -1116 7498 -1101
rect 8176 -1116 8232 -1101
rect 8286 -1116 8342 -1101
rect 9298 -1118 9354 -1101
rect 9408 -1118 9464 -1101
rect 9578 -1101 9634 -1061
rect 9688 -1101 9744 -1061
rect 9578 -1117 9634 -1101
rect 9688 -1117 9744 -1101
rect 351 -1321 407 -1265
rect 351 -1431 407 -1375
rect 691 -1310 747 -1254
rect 801 -1310 857 -1254
rect 1452 -1387 1508 -1367
rect 1562 -1387 1618 -1367
rect 1452 -1423 1508 -1387
rect 1562 -1423 1618 -1387
rect 1732 -1387 1788 -1373
rect 1842 -1387 1898 -1373
rect 2851 -1387 2907 -1366
rect 2961 -1387 3017 -1366
rect 1732 -1429 1788 -1387
rect 1842 -1429 1898 -1387
rect 2851 -1422 2907 -1387
rect 2961 -1422 3017 -1387
rect 3130 -1387 3186 -1368
rect 3240 -1387 3296 -1368
rect 3130 -1424 3186 -1387
rect 3240 -1424 3296 -1387
rect 3418 -1387 3474 -1368
rect 3528 -1387 3584 -1368
rect 3418 -1424 3474 -1387
rect 3528 -1424 3584 -1387
rect 3697 -1387 3753 -1366
rect 3807 -1387 3863 -1366
rect 4816 -1387 4872 -1373
rect 4926 -1387 4982 -1373
rect 3697 -1422 3753 -1387
rect 3807 -1422 3863 -1387
rect 4816 -1429 4872 -1387
rect 4926 -1429 4982 -1387
rect 1433 -1579 1489 -1523
rect 1543 -1579 1599 -1523
rect 5096 -1387 5152 -1367
rect 5206 -1387 5262 -1367
rect 5932 -1387 5988 -1367
rect 6042 -1387 6098 -1367
rect 5096 -1423 5152 -1387
rect 5206 -1423 5262 -1387
rect 5932 -1423 5988 -1387
rect 6042 -1423 6098 -1387
rect 931 -1646 987 -1590
rect 1041 -1646 1097 -1590
rect 1844 -1644 1900 -1588
rect 1954 -1644 2010 -1588
rect 1449 -1753 1450 -1709
rect 1450 -1753 1505 -1709
rect 1557 -1753 1613 -1709
rect 1449 -1765 1505 -1753
rect 1557 -1765 1613 -1753
rect 2010 -1753 2066 -1716
rect 2120 -1753 2176 -1716
rect 2010 -1772 2066 -1753
rect 2120 -1772 2176 -1753
rect 4704 -1644 4760 -1588
rect 4814 -1644 4870 -1588
rect 2291 -1753 2347 -1713
rect 2401 -1753 2457 -1713
rect 2291 -1769 2347 -1753
rect 2401 -1769 2457 -1753
rect 2849 -1753 2850 -1710
rect 2850 -1753 2905 -1710
rect 2959 -1753 3015 -1710
rect 3699 -1753 3755 -1710
rect 3809 -1753 3864 -1710
rect 3864 -1753 3865 -1710
rect 2849 -1766 2905 -1753
rect 2959 -1766 3015 -1753
rect 3699 -1766 3755 -1753
rect 3809 -1766 3865 -1753
rect 4257 -1753 4313 -1713
rect 4367 -1753 4423 -1713
rect 4257 -1769 4313 -1753
rect 4367 -1769 4423 -1753
rect 5113 -1578 5169 -1522
rect 5223 -1578 5279 -1522
rect 6212 -1387 6268 -1373
rect 6322 -1387 6378 -1373
rect 7331 -1387 7387 -1366
rect 7441 -1387 7497 -1366
rect 6212 -1429 6268 -1387
rect 6322 -1429 6378 -1387
rect 7331 -1422 7387 -1387
rect 7441 -1422 7497 -1387
rect 7610 -1387 7666 -1368
rect 7720 -1387 7776 -1368
rect 7610 -1424 7666 -1387
rect 7720 -1424 7776 -1387
rect 7898 -1387 7954 -1368
rect 8008 -1387 8064 -1368
rect 7898 -1424 7954 -1387
rect 8008 -1424 8064 -1387
rect 8177 -1387 8233 -1366
rect 8287 -1387 8343 -1366
rect 10085 -1310 10141 -1254
rect 10195 -1310 10251 -1254
rect 10818 729 10874 785
rect 10818 619 10874 675
rect 10947 527 11003 583
rect 10947 417 11003 473
rect 11066 356 11122 412
rect 11066 246 11122 302
rect 10947 -473 11003 -417
rect 11066 -302 11122 -246
rect 11066 -412 11122 -356
rect 10947 -583 11003 -527
rect 10818 -675 10874 -619
rect 10818 -785 10874 -729
rect 10709 -1214 10765 -1158
rect 10709 -1324 10765 -1268
rect 9296 -1387 9352 -1373
rect 9406 -1387 9462 -1373
rect 8177 -1422 8233 -1387
rect 8287 -1422 8343 -1387
rect 9296 -1429 9352 -1387
rect 9406 -1429 9462 -1387
rect 5913 -1579 5969 -1523
rect 6023 -1579 6079 -1523
rect 9576 -1387 9632 -1367
rect 9686 -1387 9742 -1367
rect 9576 -1423 9632 -1387
rect 9686 -1423 9742 -1387
rect 6324 -1644 6380 -1588
rect 6434 -1644 6490 -1588
rect 4538 -1753 4594 -1716
rect 4648 -1753 4704 -1716
rect 4538 -1772 4594 -1753
rect 4648 -1772 4704 -1753
rect 5101 -1753 5157 -1709
rect 5209 -1753 5264 -1709
rect 5264 -1753 5265 -1709
rect 5101 -1765 5157 -1753
rect 5209 -1765 5265 -1753
rect 5929 -1753 5930 -1709
rect 5930 -1753 5985 -1709
rect 6037 -1753 6093 -1709
rect 5929 -1765 5985 -1753
rect 6037 -1765 6093 -1753
rect 6490 -1753 6546 -1716
rect 6600 -1753 6656 -1716
rect 6490 -1772 6546 -1753
rect 6600 -1772 6656 -1753
rect 9184 -1644 9240 -1588
rect 9294 -1644 9350 -1588
rect 6771 -1753 6827 -1713
rect 6881 -1753 6937 -1713
rect 6771 -1769 6827 -1753
rect 6881 -1769 6937 -1753
rect 7329 -1753 7330 -1710
rect 7330 -1753 7385 -1710
rect 7439 -1753 7495 -1710
rect 8179 -1753 8235 -1710
rect 8289 -1753 8344 -1710
rect 8344 -1753 8345 -1710
rect 7329 -1766 7385 -1753
rect 7439 -1766 7495 -1753
rect 8179 -1766 8235 -1753
rect 8289 -1766 8345 -1753
rect 8737 -1753 8793 -1713
rect 8847 -1753 8903 -1713
rect 8737 -1769 8793 -1753
rect 8847 -1769 8903 -1753
rect 9593 -1578 9649 -1522
rect 9703 -1578 9759 -1522
rect 10295 -1646 10353 -1590
rect 10405 -1646 10463 -1590
rect 9018 -1753 9074 -1716
rect 9128 -1753 9184 -1716
rect 9018 -1772 9074 -1753
rect 9128 -1772 9184 -1753
rect 9581 -1753 9637 -1709
rect 9689 -1753 9744 -1709
rect 9744 -1753 9745 -1709
rect 9581 -1765 9637 -1753
rect 9689 -1765 9745 -1753
rect 2291 -2039 2347 -2024
rect 2401 -2039 2457 -2024
rect 4257 -2039 4313 -2024
rect 4367 -2039 4423 -2024
rect 6771 -2039 6827 -2024
rect 6881 -2039 6937 -2024
rect 8737 -2039 8793 -2024
rect 8847 -2039 8903 -2024
rect 2291 -2080 2347 -2039
rect 2401 -2080 2457 -2039
rect 4257 -2080 4313 -2039
rect 4367 -2080 4423 -2039
rect 6771 -2080 6827 -2039
rect 6881 -2080 6937 -2039
rect 8737 -2080 8793 -2039
rect 8847 -2080 8903 -2039
rect 3048 -2191 3104 -2135
rect 3158 -2191 3214 -2135
rect 3500 -2191 3556 -2135
rect 3610 -2191 3666 -2135
rect 7528 -2191 7584 -2135
rect 7638 -2191 7694 -2135
rect 7980 -2191 8036 -2135
rect 8090 -2191 8146 -2135
<< metal2 >>
rect 3036 2191 3226 2195
rect 3036 2135 3048 2191
rect 3104 2135 3158 2191
rect 3214 2135 3226 2191
rect 3036 2131 3226 2135
rect 3488 2191 3678 2195
rect 3488 2135 3500 2191
rect 3556 2135 3610 2191
rect 3666 2135 3678 2191
rect 3488 2131 3678 2135
rect 7516 2191 7706 2195
rect 7516 2135 7528 2191
rect 7584 2135 7638 2191
rect 7694 2135 7706 2191
rect 7516 2131 7706 2135
rect 7968 2191 8158 2195
rect 7968 2135 7980 2191
rect 8036 2135 8090 2191
rect 8146 2135 8158 2191
rect 7968 2131 8158 2135
rect 2291 2089 2347 2090
rect 2277 2080 2477 2089
rect 2277 2024 2291 2080
rect 2347 2024 2401 2080
rect 2457 2024 2477 2080
rect 2277 2012 2477 2024
rect 2010 1780 2066 1782
rect 1437 1770 1637 1779
rect 1185 1765 1637 1770
rect 1185 1709 1449 1765
rect 1505 1709 1557 1765
rect 1613 1709 1637 1765
rect 1185 1704 1637 1709
rect 915 1646 1112 1651
rect 915 1590 931 1646
rect 987 1590 1041 1646
rect 1097 1590 1112 1646
rect 915 1585 1112 1590
rect 346 1431 412 1446
rect 346 1375 351 1431
rect 407 1375 412 1431
rect 346 1321 412 1375
rect 346 1265 351 1321
rect 407 1315 412 1321
rect 407 1310 875 1315
rect 407 1265 691 1310
rect 346 1254 691 1265
rect 747 1254 801 1310
rect 857 1254 875 1310
rect 346 1249 875 1254
rect 236 1126 302 1141
rect 236 1070 241 1126
rect 297 1070 302 1126
rect 114 1004 180 1019
rect 114 948 119 1004
rect 175 948 180 1004
rect 114 894 180 948
rect 236 1016 302 1070
rect 236 960 241 1016
rect 297 1010 302 1016
rect 297 1005 866 1010
rect 297 960 682 1005
rect 236 949 682 960
rect 738 949 792 1005
rect 848 949 866 1005
rect 236 944 866 949
rect 114 838 119 894
rect 175 888 180 894
rect 1012 893 1078 1585
rect 932 888 1129 893
rect 175 838 948 888
rect 114 832 948 838
rect 1004 832 1058 888
rect 1114 832 1129 888
rect 114 827 1129 832
rect 114 822 932 827
rect 670 664 867 669
rect 670 608 683 664
rect 739 608 793 664
rect 849 608 867 664
rect 670 603 867 608
rect 0 412 66 427
rect 0 356 5 412
rect 61 356 66 412
rect 0 302 66 356
rect 0 246 5 302
rect 61 296 66 302
rect 1185 355 1251 1704
rect 1437 1702 1637 1704
rect 1997 1772 2197 1780
rect 1997 1716 2010 1772
rect 2066 1716 2120 1772
rect 2176 1716 2197 1772
rect 1997 1703 2197 1716
rect 2277 1769 2477 1780
rect 2277 1713 2291 1769
rect 2347 1713 2401 1769
rect 2457 1713 2477 1769
rect 2277 1703 2477 1713
rect 2837 1766 3037 1780
rect 2837 1710 2849 1766
rect 2905 1710 2959 1766
rect 3015 1710 3037 1766
rect 2837 1703 3037 1710
rect 1447 1699 1503 1702
rect 1832 1644 2024 1647
rect 1832 1588 1844 1644
rect 1900 1588 1954 1644
rect 2010 1588 2024 1644
rect 1832 1585 2024 1588
rect 1421 1579 1611 1583
rect 1421 1523 1433 1579
rect 1489 1523 1543 1579
rect 1599 1523 1611 1579
rect 1421 1518 1611 1523
rect 1433 1517 1611 1518
rect 1838 1437 1904 1585
rect 1437 1423 1637 1435
rect 1437 1367 1452 1423
rect 1508 1367 1562 1423
rect 1618 1367 1637 1423
rect 1437 1357 1637 1367
rect 1717 1429 1917 1437
rect 1717 1373 1732 1429
rect 1788 1373 1842 1429
rect 1898 1373 1917 1429
rect 1717 1360 1917 1373
rect 2394 1379 2466 1703
rect 3124 1437 3190 2131
rect 3524 1437 3590 2131
rect 4367 2089 4423 2090
rect 6771 2089 6827 2090
rect 4237 2080 4437 2089
rect 4237 2024 4257 2080
rect 4313 2024 4367 2080
rect 4423 2024 4437 2080
rect 4237 2012 4437 2024
rect 6757 2080 6957 2089
rect 6757 2024 6771 2080
rect 6827 2024 6881 2080
rect 6937 2024 6957 2080
rect 6757 2012 6957 2024
rect 4648 1780 4704 1782
rect 6490 1780 6546 1782
rect 3677 1766 3877 1780
rect 3677 1710 3699 1766
rect 3755 1710 3809 1766
rect 3865 1710 3877 1766
rect 3677 1703 3877 1710
rect 4237 1769 4437 1780
rect 4237 1713 4257 1769
rect 4313 1713 4367 1769
rect 4423 1713 4437 1769
rect 4237 1703 4437 1713
rect 4517 1772 4717 1780
rect 4517 1716 4538 1772
rect 4594 1716 4648 1772
rect 4704 1716 4717 1772
rect 4517 1703 4717 1716
rect 5077 1770 5277 1779
rect 5917 1770 6117 1779
rect 5077 1765 5529 1770
rect 5077 1709 5101 1765
rect 5157 1709 5209 1765
rect 5265 1709 5529 1765
rect 5077 1704 5529 1709
rect 2837 1422 3037 1436
rect 2837 1379 2851 1422
rect 2394 1366 2851 1379
rect 2907 1366 2961 1422
rect 3017 1366 3037 1422
rect 2394 1356 3037 1366
rect 3117 1424 3317 1437
rect 3117 1368 3130 1424
rect 3186 1368 3240 1424
rect 3296 1368 3317 1424
rect 3117 1360 3317 1368
rect 3397 1424 3597 1437
rect 3397 1368 3418 1424
rect 3474 1368 3528 1424
rect 3584 1368 3597 1424
rect 3397 1360 3597 1368
rect 3677 1422 3877 1436
rect 3677 1366 3697 1422
rect 3753 1366 3807 1422
rect 3863 1379 3877 1422
rect 4248 1379 4320 1703
rect 5077 1702 5277 1704
rect 5211 1699 5267 1702
rect 4690 1644 4882 1647
rect 4690 1588 4704 1644
rect 4760 1588 4814 1644
rect 4870 1588 4882 1644
rect 4690 1585 4882 1588
rect 4810 1437 4876 1585
rect 5101 1578 5291 1583
rect 5101 1522 5113 1578
rect 5169 1522 5223 1578
rect 5279 1522 5291 1578
rect 5101 1517 5291 1522
rect 3863 1366 4320 1379
rect 3130 1358 3257 1360
rect 2394 1307 2952 1356
rect 1437 1117 1637 1127
rect 1437 1061 1450 1117
rect 1506 1061 1560 1117
rect 1616 1061 1637 1117
rect 1437 1050 1637 1061
rect 1717 1118 1917 1128
rect 1717 1062 1730 1118
rect 1786 1062 1840 1118
rect 1896 1062 1917 1118
rect 1717 1051 1917 1062
rect 2837 1116 3037 1128
rect 3181 1121 3257 1358
rect 3472 1358 3584 1360
rect 3472 1121 3548 1358
rect 3677 1356 4320 1366
rect 4797 1429 4997 1437
rect 4797 1373 4816 1429
rect 4872 1373 4926 1429
rect 4982 1373 4997 1429
rect 4797 1360 4997 1373
rect 5077 1423 5277 1435
rect 5077 1367 5096 1423
rect 5152 1367 5206 1423
rect 5262 1367 5277 1423
rect 5077 1357 5277 1367
rect 3762 1307 4320 1356
rect 2837 1060 2852 1116
rect 2908 1060 2962 1116
rect 3018 1060 3037 1116
rect 1838 894 1904 1051
rect 2837 1050 3037 1060
rect 3119 1116 3316 1121
rect 3119 1060 3135 1116
rect 3191 1060 3245 1116
rect 3301 1060 3316 1116
rect 3119 1055 3316 1060
rect 3399 1116 3596 1121
rect 3399 1060 3415 1116
rect 3471 1060 3525 1116
rect 3581 1060 3596 1116
rect 3399 1055 3596 1060
rect 3677 1116 3877 1128
rect 3677 1060 3696 1116
rect 3752 1060 3806 1116
rect 3862 1060 3877 1116
rect 3677 1050 3877 1060
rect 4797 1118 4997 1128
rect 4797 1062 4818 1118
rect 4874 1062 4928 1118
rect 4984 1062 4997 1118
rect 4797 1051 4997 1062
rect 5077 1117 5277 1127
rect 5077 1061 5098 1117
rect 5154 1061 5208 1117
rect 5264 1061 5277 1117
rect 2854 928 2922 1050
rect 1831 889 1911 894
rect 1831 833 1843 889
rect 1899 833 1911 889
rect 1831 827 1911 833
rect 2359 860 2922 928
rect 3792 928 3860 1050
rect 3792 860 4355 928
rect 4810 894 4876 1051
rect 5077 1050 5277 1061
rect 2359 785 2427 860
rect 4287 785 4355 860
rect 4803 889 4883 894
rect 4803 833 4815 889
rect 4871 833 4883 889
rect 4803 827 4883 833
rect 1437 775 1637 785
rect 1437 719 1450 775
rect 1506 719 1560 775
rect 1616 719 1637 775
rect 1437 708 1637 719
rect 1997 774 2197 785
rect 1997 718 2011 774
rect 2067 718 2121 774
rect 2177 718 2197 774
rect 1997 708 2197 718
rect 2277 775 2477 785
rect 2277 719 2292 775
rect 2348 719 2402 775
rect 2458 719 2477 775
rect 2277 708 2477 719
rect 4237 775 4437 785
rect 4237 719 4256 775
rect 4312 719 4366 775
rect 4422 719 4437 775
rect 4237 708 4437 719
rect 4517 774 4717 785
rect 4517 718 4537 774
rect 4593 718 4647 774
rect 4703 718 4717 774
rect 4517 708 4717 718
rect 5077 775 5277 785
rect 5077 719 5098 775
rect 5154 719 5208 775
rect 5264 719 5277 775
rect 5077 708 5277 719
rect 2059 479 2129 708
rect 1439 472 1636 477
rect 1439 416 1452 472
rect 1508 416 1562 472
rect 1618 416 1636 472
rect 1439 411 1636 416
rect 1997 474 2194 479
rect 1997 418 2010 474
rect 2066 418 2120 474
rect 2176 418 2194 474
rect 1997 413 2194 418
rect 2837 461 3037 476
rect 2837 405 2849 461
rect 2905 405 2959 461
rect 3015 405 3037 461
rect 2837 399 3037 405
rect 3677 461 3877 476
rect 3677 405 3699 461
rect 3755 405 3809 461
rect 3865 405 3877 461
rect 3677 399 3877 405
rect 2837 395 2905 399
rect 3809 395 3877 399
rect 2837 355 2903 395
rect 61 291 871 296
rect 61 246 687 291
rect 0 235 687 246
rect 743 235 797 291
rect 853 235 871 291
rect 1185 289 2903 355
rect 3811 355 3877 395
rect 5463 355 5529 1704
rect 3811 289 5529 355
rect 5665 1765 6117 1770
rect 5665 1709 5929 1765
rect 5985 1709 6037 1765
rect 6093 1709 6117 1765
rect 5665 1704 6117 1709
rect 5665 355 5731 1704
rect 5917 1702 6117 1704
rect 6477 1772 6677 1780
rect 6477 1716 6490 1772
rect 6546 1716 6600 1772
rect 6656 1716 6677 1772
rect 6477 1703 6677 1716
rect 6757 1769 6957 1780
rect 6757 1713 6771 1769
rect 6827 1713 6881 1769
rect 6937 1713 6957 1769
rect 6757 1703 6957 1713
rect 7317 1766 7517 1780
rect 7317 1710 7329 1766
rect 7385 1710 7439 1766
rect 7495 1710 7517 1766
rect 7317 1703 7517 1710
rect 5927 1699 5983 1702
rect 6312 1644 6504 1647
rect 6312 1588 6324 1644
rect 6380 1588 6434 1644
rect 6490 1588 6504 1644
rect 6312 1585 6504 1588
rect 5901 1579 6091 1583
rect 5901 1523 5913 1579
rect 5969 1523 6023 1579
rect 6079 1523 6091 1579
rect 5901 1518 6091 1523
rect 5913 1517 6091 1518
rect 6318 1437 6384 1585
rect 5917 1423 6117 1435
rect 5917 1367 5932 1423
rect 5988 1367 6042 1423
rect 6098 1367 6117 1423
rect 5917 1357 6117 1367
rect 6197 1429 6397 1437
rect 6197 1373 6212 1429
rect 6268 1373 6322 1429
rect 6378 1373 6397 1429
rect 6197 1360 6397 1373
rect 6874 1379 6946 1703
rect 7604 1437 7670 2131
rect 8004 1437 8070 2131
rect 8847 2089 8903 2090
rect 8717 2080 8917 2089
rect 8717 2024 8737 2080
rect 8793 2024 8847 2080
rect 8903 2024 8917 2080
rect 8717 2012 8917 2024
rect 9128 1780 9184 1782
rect 8157 1766 8357 1780
rect 8157 1710 8179 1766
rect 8235 1710 8289 1766
rect 8345 1710 8357 1766
rect 8157 1703 8357 1710
rect 8717 1769 8917 1780
rect 8717 1713 8737 1769
rect 8793 1713 8847 1769
rect 8903 1713 8917 1769
rect 8717 1703 8917 1713
rect 8997 1772 9197 1780
rect 8997 1716 9018 1772
rect 9074 1716 9128 1772
rect 9184 1716 9197 1772
rect 8997 1703 9197 1716
rect 9557 1770 9757 1779
rect 9557 1765 10009 1770
rect 9557 1709 9581 1765
rect 9637 1709 9689 1765
rect 9745 1709 10009 1765
rect 9557 1704 10009 1709
rect 7317 1422 7517 1436
rect 7317 1379 7331 1422
rect 6874 1366 7331 1379
rect 7387 1366 7441 1422
rect 7497 1366 7517 1422
rect 6874 1356 7517 1366
rect 7597 1424 7797 1437
rect 7597 1368 7610 1424
rect 7666 1368 7720 1424
rect 7776 1368 7797 1424
rect 7597 1360 7797 1368
rect 7877 1424 8077 1437
rect 7877 1368 7898 1424
rect 7954 1368 8008 1424
rect 8064 1368 8077 1424
rect 7877 1360 8077 1368
rect 8157 1422 8357 1436
rect 8157 1366 8177 1422
rect 8233 1366 8287 1422
rect 8343 1379 8357 1422
rect 8728 1379 8800 1703
rect 9557 1702 9757 1704
rect 9691 1699 9747 1702
rect 9170 1644 9362 1647
rect 9170 1588 9184 1644
rect 9240 1588 9294 1644
rect 9350 1588 9362 1644
rect 9170 1585 9362 1588
rect 9290 1437 9356 1585
rect 9581 1578 9771 1583
rect 9581 1522 9593 1578
rect 9649 1522 9703 1578
rect 9759 1522 9771 1578
rect 9581 1517 9771 1522
rect 8343 1366 8800 1379
rect 7610 1358 7666 1360
rect 8008 1358 8064 1360
rect 8157 1356 8800 1366
rect 9277 1429 9477 1437
rect 9277 1373 9296 1429
rect 9352 1373 9406 1429
rect 9462 1373 9477 1429
rect 9277 1360 9477 1373
rect 9557 1423 9757 1435
rect 9557 1367 9576 1423
rect 9632 1367 9686 1423
rect 9742 1367 9757 1423
rect 9557 1357 9757 1367
rect 6874 1307 7432 1356
rect 8242 1307 8800 1356
rect 5917 1117 6117 1127
rect 5917 1061 5930 1117
rect 5986 1061 6040 1117
rect 6096 1061 6117 1117
rect 5917 1050 6117 1061
rect 6197 1118 6397 1128
rect 6197 1062 6210 1118
rect 6266 1062 6320 1118
rect 6376 1062 6397 1118
rect 6197 1051 6397 1062
rect 7317 1116 7517 1128
rect 7317 1060 7332 1116
rect 7388 1060 7442 1116
rect 7498 1060 7517 1116
rect 6318 894 6384 1051
rect 7317 1050 7517 1060
rect 8157 1116 8357 1128
rect 8157 1060 8176 1116
rect 8232 1060 8286 1116
rect 8342 1060 8357 1116
rect 8157 1050 8357 1060
rect 9277 1118 9477 1128
rect 9277 1062 9298 1118
rect 9354 1062 9408 1118
rect 9464 1062 9477 1118
rect 9277 1051 9477 1062
rect 9557 1117 9757 1127
rect 9557 1061 9578 1117
rect 9634 1061 9688 1117
rect 9744 1061 9757 1117
rect 7334 928 7402 1050
rect 6311 889 6391 894
rect 6311 833 6323 889
rect 6379 833 6391 889
rect 6311 827 6391 833
rect 6839 860 7402 928
rect 8272 928 8340 1050
rect 8272 860 8835 928
rect 9290 894 9356 1051
rect 9557 1050 9757 1061
rect 6839 785 6907 860
rect 8767 785 8835 860
rect 9283 889 9363 894
rect 9283 833 9295 889
rect 9351 833 9363 889
rect 9283 827 9363 833
rect 5917 775 6117 785
rect 5917 719 5930 775
rect 5986 719 6040 775
rect 6096 719 6117 775
rect 5917 708 6117 719
rect 6477 774 6677 785
rect 6477 718 6491 774
rect 6547 718 6601 774
rect 6657 718 6677 774
rect 6477 708 6677 718
rect 6757 775 6957 785
rect 6757 719 6772 775
rect 6828 719 6882 775
rect 6938 719 6957 775
rect 6757 708 6957 719
rect 8717 775 8917 785
rect 8717 719 8736 775
rect 8792 719 8846 775
rect 8902 719 8917 775
rect 8717 708 8917 719
rect 8997 774 9197 785
rect 8997 718 9017 774
rect 9073 718 9127 774
rect 9183 718 9197 774
rect 8997 708 9197 718
rect 9557 775 9757 785
rect 9557 719 9578 775
rect 9634 719 9688 775
rect 9744 719 9757 775
rect 9557 708 9757 719
rect 7317 461 7517 476
rect 7317 405 7329 461
rect 7385 405 7439 461
rect 7495 405 7517 461
rect 7317 399 7517 405
rect 8157 461 8357 476
rect 8157 405 8179 461
rect 8235 405 8289 461
rect 8345 405 8357 461
rect 8157 399 8357 405
rect 7317 395 7385 399
rect 8289 395 8357 399
rect 7317 355 7383 395
rect 5665 289 7383 355
rect 8291 355 8357 395
rect 9943 355 10009 1704
rect 10282 1646 10479 1651
rect 10282 1590 10295 1646
rect 10353 1590 10405 1646
rect 10463 1590 10479 1646
rect 10282 1585 10479 1590
rect 10704 1324 10767 1339
rect 10704 1315 10709 1324
rect 10067 1310 10709 1315
rect 10067 1254 10085 1310
rect 10141 1254 10195 1310
rect 10251 1268 10709 1310
rect 10765 1315 10767 1324
rect 10765 1268 10893 1315
rect 10251 1254 10893 1268
rect 10067 1249 10893 1254
rect 10704 1214 10767 1249
rect 10704 1158 10709 1214
rect 10765 1158 10767 1214
rect 10704 1141 10767 1158
rect 10066 888 10263 893
rect 10066 832 10084 888
rect 10140 832 10194 888
rect 10250 832 10263 888
rect 10066 827 10263 832
rect 10137 566 10203 827
rect 10813 785 10879 800
rect 10813 729 10818 785
rect 10874 729 10879 785
rect 10813 675 10879 729
rect 10813 669 10818 675
rect 10315 664 10818 669
rect 10315 608 10333 664
rect 10389 608 10443 664
rect 10499 619 10818 664
rect 10874 619 10879 675
rect 10499 608 10879 619
rect 10315 603 10879 608
rect 10942 583 11005 598
rect 10065 561 10262 566
rect 10065 505 10083 561
rect 10139 505 10193 561
rect 10249 505 10262 561
rect 10065 500 10262 505
rect 10196 467 10262 500
rect 10942 527 10947 583
rect 11003 527 11005 583
rect 10942 473 11005 527
rect 10942 467 10947 473
rect 10196 417 10947 467
rect 11003 417 11005 473
rect 10196 401 11005 417
rect 11063 412 11127 427
rect 8291 289 10009 355
rect 11063 356 11066 412
rect 11122 356 11127 412
rect 11063 302 11127 356
rect 11063 296 11066 302
rect 10295 291 11066 296
rect 0 230 871 235
rect 10295 235 10313 291
rect 10369 235 10423 291
rect 10479 246 11066 291
rect 11122 246 11127 302
rect 10479 235 11127 246
rect 10295 230 11127 235
rect 0 -235 871 -230
rect 0 -246 687 -235
rect 0 -302 5 -246
rect 61 -291 687 -246
rect 743 -291 797 -235
rect 853 -291 871 -235
rect 10295 -235 11127 -230
rect 61 -296 871 -291
rect 61 -302 66 -296
rect 0 -356 66 -302
rect 0 -412 5 -356
rect 61 -412 66 -356
rect 0 -427 66 -412
rect 1185 -355 2903 -289
rect 670 -608 867 -603
rect 670 -664 683 -608
rect 739 -664 793 -608
rect 849 -664 867 -608
rect 670 -669 867 -664
rect 114 -827 932 -822
rect 114 -832 1129 -827
rect 114 -838 948 -832
rect 114 -894 119 -838
rect 175 -888 948 -838
rect 1004 -888 1058 -832
rect 1114 -888 1129 -832
rect 175 -894 180 -888
rect 932 -893 1129 -888
rect 114 -948 180 -894
rect 114 -1004 119 -948
rect 175 -1004 180 -948
rect 114 -1019 180 -1004
rect 236 -949 866 -944
rect 236 -960 682 -949
rect 236 -1016 241 -960
rect 297 -1005 682 -960
rect 738 -1005 792 -949
rect 848 -1005 866 -949
rect 297 -1010 866 -1005
rect 297 -1016 302 -1010
rect 236 -1070 302 -1016
rect 236 -1126 241 -1070
rect 297 -1126 302 -1070
rect 236 -1141 302 -1126
rect 346 -1254 875 -1249
rect 346 -1265 691 -1254
rect 346 -1321 351 -1265
rect 407 -1310 691 -1265
rect 747 -1310 801 -1254
rect 857 -1310 875 -1254
rect 407 -1315 875 -1310
rect 407 -1321 412 -1315
rect 346 -1375 412 -1321
rect 346 -1431 351 -1375
rect 407 -1431 412 -1375
rect 346 -1446 412 -1431
rect 1012 -1585 1078 -893
rect 915 -1590 1112 -1585
rect 915 -1646 931 -1590
rect 987 -1646 1041 -1590
rect 1097 -1646 1112 -1590
rect 915 -1651 1112 -1646
rect 1185 -1704 1251 -355
rect 2837 -395 2903 -355
rect 3811 -355 5529 -289
rect 3811 -395 3877 -355
rect 2837 -399 2905 -395
rect 3809 -399 3877 -395
rect 2837 -405 3037 -399
rect 1439 -416 1636 -411
rect 1439 -472 1452 -416
rect 1508 -472 1562 -416
rect 1618 -472 1636 -416
rect 1439 -477 1636 -472
rect 1997 -418 2194 -413
rect 1997 -474 2010 -418
rect 2066 -474 2120 -418
rect 2176 -474 2194 -418
rect 1997 -479 2194 -474
rect 2837 -461 2849 -405
rect 2905 -461 2959 -405
rect 3015 -461 3037 -405
rect 2837 -476 3037 -461
rect 3677 -405 3877 -399
rect 3677 -461 3699 -405
rect 3755 -461 3809 -405
rect 3865 -461 3877 -405
rect 3677 -476 3877 -461
rect 2059 -708 2129 -479
rect 1437 -719 1637 -708
rect 1437 -775 1450 -719
rect 1506 -775 1560 -719
rect 1616 -775 1637 -719
rect 1437 -785 1637 -775
rect 1997 -718 2197 -708
rect 1997 -774 2011 -718
rect 2067 -774 2121 -718
rect 2177 -774 2197 -718
rect 1997 -785 2197 -774
rect 2277 -719 2477 -708
rect 2277 -775 2292 -719
rect 2348 -775 2402 -719
rect 2458 -775 2477 -719
rect 2277 -785 2477 -775
rect 4237 -719 4437 -708
rect 4237 -775 4256 -719
rect 4312 -775 4366 -719
rect 4422 -775 4437 -719
rect 4237 -785 4437 -775
rect 4517 -718 4717 -708
rect 4517 -774 4537 -718
rect 4593 -774 4647 -718
rect 4703 -774 4717 -718
rect 4517 -785 4717 -774
rect 5077 -719 5277 -708
rect 5077 -775 5098 -719
rect 5154 -775 5208 -719
rect 5264 -775 5277 -719
rect 5077 -785 5277 -775
rect 1831 -833 1911 -827
rect 1831 -889 1843 -833
rect 1899 -889 1911 -833
rect 1831 -894 1911 -889
rect 2359 -860 2427 -785
rect 4287 -860 4355 -785
rect 1437 -1061 1637 -1050
rect 1838 -1051 1904 -894
rect 2359 -928 2922 -860
rect 2854 -1050 2922 -928
rect 3792 -928 4355 -860
rect 4803 -833 4883 -827
rect 4803 -889 4815 -833
rect 4871 -889 4883 -833
rect 4803 -894 4883 -889
rect 3792 -1050 3860 -928
rect 1437 -1117 1450 -1061
rect 1506 -1117 1560 -1061
rect 1616 -1117 1637 -1061
rect 1437 -1127 1637 -1117
rect 1717 -1062 1917 -1051
rect 1717 -1118 1730 -1062
rect 1786 -1118 1840 -1062
rect 1896 -1118 1917 -1062
rect 1717 -1128 1917 -1118
rect 2837 -1060 3037 -1050
rect 2837 -1116 2852 -1060
rect 2908 -1116 2962 -1060
rect 3018 -1116 3037 -1060
rect 2837 -1128 3037 -1116
rect 3119 -1060 3316 -1055
rect 3119 -1116 3135 -1060
rect 3191 -1116 3245 -1060
rect 3301 -1116 3316 -1060
rect 3119 -1121 3316 -1116
rect 3399 -1060 3596 -1055
rect 3399 -1116 3415 -1060
rect 3471 -1116 3525 -1060
rect 3581 -1116 3596 -1060
rect 3399 -1121 3596 -1116
rect 3677 -1060 3877 -1050
rect 4810 -1051 4876 -894
rect 3677 -1116 3696 -1060
rect 3752 -1116 3806 -1060
rect 3862 -1116 3877 -1060
rect 2394 -1356 2952 -1307
rect 1437 -1367 1637 -1357
rect 1437 -1423 1452 -1367
rect 1508 -1423 1562 -1367
rect 1618 -1423 1637 -1367
rect 1437 -1435 1637 -1423
rect 1717 -1373 1917 -1360
rect 1717 -1429 1732 -1373
rect 1788 -1429 1842 -1373
rect 1898 -1429 1917 -1373
rect 1717 -1437 1917 -1429
rect 2394 -1366 3037 -1356
rect 3181 -1358 3257 -1121
rect 3130 -1360 3257 -1358
rect 3472 -1358 3548 -1121
rect 3677 -1128 3877 -1116
rect 4797 -1062 4997 -1051
rect 4797 -1118 4818 -1062
rect 4874 -1118 4928 -1062
rect 4984 -1118 4997 -1062
rect 4797 -1128 4997 -1118
rect 5077 -1061 5277 -1050
rect 5077 -1117 5098 -1061
rect 5154 -1117 5208 -1061
rect 5264 -1117 5277 -1061
rect 5077 -1127 5277 -1117
rect 3762 -1356 4320 -1307
rect 3472 -1360 3584 -1358
rect 2394 -1379 2851 -1366
rect 1433 -1518 1611 -1517
rect 1421 -1523 1611 -1518
rect 1421 -1579 1433 -1523
rect 1489 -1579 1543 -1523
rect 1599 -1579 1611 -1523
rect 1421 -1583 1611 -1579
rect 1838 -1585 1904 -1437
rect 1832 -1588 2024 -1585
rect 1832 -1644 1844 -1588
rect 1900 -1644 1954 -1588
rect 2010 -1644 2024 -1588
rect 1832 -1647 2024 -1644
rect 1447 -1702 1503 -1699
rect 1437 -1704 1637 -1702
rect 2394 -1703 2466 -1379
rect 2837 -1422 2851 -1379
rect 2907 -1422 2961 -1366
rect 3017 -1422 3037 -1366
rect 2837 -1436 3037 -1422
rect 3117 -1368 3317 -1360
rect 3117 -1424 3130 -1368
rect 3186 -1424 3240 -1368
rect 3296 -1424 3317 -1368
rect 3117 -1437 3317 -1424
rect 3397 -1368 3597 -1360
rect 3397 -1424 3418 -1368
rect 3474 -1424 3528 -1368
rect 3584 -1424 3597 -1368
rect 3397 -1437 3597 -1424
rect 3677 -1366 4320 -1356
rect 3677 -1422 3697 -1366
rect 3753 -1422 3807 -1366
rect 3863 -1379 4320 -1366
rect 3863 -1422 3877 -1379
rect 3677 -1436 3877 -1422
rect 1185 -1709 1637 -1704
rect 1185 -1765 1449 -1709
rect 1505 -1765 1557 -1709
rect 1613 -1765 1637 -1709
rect 1185 -1770 1637 -1765
rect 1437 -1779 1637 -1770
rect 1997 -1716 2197 -1703
rect 1997 -1772 2010 -1716
rect 2066 -1772 2120 -1716
rect 2176 -1772 2197 -1716
rect 1997 -1780 2197 -1772
rect 2277 -1713 2477 -1703
rect 2277 -1769 2291 -1713
rect 2347 -1769 2401 -1713
rect 2457 -1769 2477 -1713
rect 2277 -1780 2477 -1769
rect 2837 -1710 3037 -1703
rect 2837 -1766 2849 -1710
rect 2905 -1766 2959 -1710
rect 3015 -1766 3037 -1710
rect 2837 -1780 3037 -1766
rect 2010 -1782 2066 -1780
rect 2277 -2024 2477 -2012
rect 2277 -2080 2291 -2024
rect 2347 -2080 2401 -2024
rect 2457 -2080 2477 -2024
rect 2277 -2089 2477 -2080
rect 2291 -2090 2347 -2089
rect 3124 -2131 3190 -1437
rect 3524 -2131 3590 -1437
rect 4248 -1703 4320 -1379
rect 4797 -1373 4997 -1360
rect 4797 -1429 4816 -1373
rect 4872 -1429 4926 -1373
rect 4982 -1429 4997 -1373
rect 4797 -1437 4997 -1429
rect 5077 -1367 5277 -1357
rect 5077 -1423 5096 -1367
rect 5152 -1423 5206 -1367
rect 5262 -1423 5277 -1367
rect 5077 -1435 5277 -1423
rect 4810 -1585 4876 -1437
rect 5101 -1522 5291 -1517
rect 5101 -1578 5113 -1522
rect 5169 -1578 5223 -1522
rect 5279 -1578 5291 -1522
rect 5101 -1583 5291 -1578
rect 4690 -1588 4882 -1585
rect 4690 -1644 4704 -1588
rect 4760 -1644 4814 -1588
rect 4870 -1644 4882 -1588
rect 4690 -1647 4882 -1644
rect 5211 -1702 5267 -1699
rect 3677 -1710 3877 -1703
rect 3677 -1766 3699 -1710
rect 3755 -1766 3809 -1710
rect 3865 -1766 3877 -1710
rect 3677 -1780 3877 -1766
rect 4237 -1713 4437 -1703
rect 4237 -1769 4257 -1713
rect 4313 -1769 4367 -1713
rect 4423 -1769 4437 -1713
rect 4237 -1780 4437 -1769
rect 4517 -1716 4717 -1703
rect 4517 -1772 4538 -1716
rect 4594 -1772 4648 -1716
rect 4704 -1772 4717 -1716
rect 4517 -1780 4717 -1772
rect 5077 -1704 5277 -1702
rect 5463 -1704 5529 -355
rect 5077 -1709 5529 -1704
rect 5077 -1765 5101 -1709
rect 5157 -1765 5209 -1709
rect 5265 -1765 5529 -1709
rect 5077 -1770 5529 -1765
rect 5665 -355 7383 -289
rect 5665 -1704 5731 -355
rect 7317 -395 7383 -355
rect 8291 -355 10009 -289
rect 10295 -291 10313 -235
rect 10369 -291 10423 -235
rect 10479 -246 11127 -235
rect 10479 -291 11066 -246
rect 10295 -296 11066 -291
rect 8291 -395 8357 -355
rect 7317 -399 7385 -395
rect 8289 -399 8357 -395
rect 7317 -405 7517 -399
rect 7317 -461 7329 -405
rect 7385 -461 7439 -405
rect 7495 -461 7517 -405
rect 7317 -476 7517 -461
rect 8157 -405 8357 -399
rect 8157 -461 8179 -405
rect 8235 -461 8289 -405
rect 8345 -461 8357 -405
rect 8157 -476 8357 -461
rect 5917 -719 6117 -708
rect 5917 -775 5930 -719
rect 5986 -775 6040 -719
rect 6096 -775 6117 -719
rect 5917 -785 6117 -775
rect 6477 -718 6677 -708
rect 6477 -774 6491 -718
rect 6547 -774 6601 -718
rect 6657 -774 6677 -718
rect 6477 -785 6677 -774
rect 6757 -719 6957 -708
rect 6757 -775 6772 -719
rect 6828 -775 6882 -719
rect 6938 -775 6957 -719
rect 6757 -785 6957 -775
rect 8717 -719 8917 -708
rect 8717 -775 8736 -719
rect 8792 -775 8846 -719
rect 8902 -775 8917 -719
rect 8717 -785 8917 -775
rect 8997 -718 9197 -708
rect 8997 -774 9017 -718
rect 9073 -774 9127 -718
rect 9183 -774 9197 -718
rect 8997 -785 9197 -774
rect 9557 -719 9757 -708
rect 9557 -775 9578 -719
rect 9634 -775 9688 -719
rect 9744 -775 9757 -719
rect 9557 -785 9757 -775
rect 6311 -833 6391 -827
rect 6311 -889 6323 -833
rect 6379 -889 6391 -833
rect 6311 -894 6391 -889
rect 6839 -860 6907 -785
rect 8767 -860 8835 -785
rect 5917 -1061 6117 -1050
rect 6318 -1051 6384 -894
rect 6839 -928 7402 -860
rect 7334 -1050 7402 -928
rect 8272 -928 8835 -860
rect 9283 -833 9363 -827
rect 9283 -889 9295 -833
rect 9351 -889 9363 -833
rect 9283 -894 9363 -889
rect 8272 -1050 8340 -928
rect 5917 -1117 5930 -1061
rect 5986 -1117 6040 -1061
rect 6096 -1117 6117 -1061
rect 5917 -1127 6117 -1117
rect 6197 -1062 6397 -1051
rect 6197 -1118 6210 -1062
rect 6266 -1118 6320 -1062
rect 6376 -1118 6397 -1062
rect 6197 -1128 6397 -1118
rect 7317 -1060 7517 -1050
rect 7317 -1116 7332 -1060
rect 7388 -1116 7442 -1060
rect 7498 -1116 7517 -1060
rect 7317 -1128 7517 -1116
rect 8157 -1060 8357 -1050
rect 9290 -1051 9356 -894
rect 8157 -1116 8176 -1060
rect 8232 -1116 8286 -1060
rect 8342 -1116 8357 -1060
rect 8157 -1128 8357 -1116
rect 9277 -1062 9477 -1051
rect 9277 -1118 9298 -1062
rect 9354 -1118 9408 -1062
rect 9464 -1118 9477 -1062
rect 9277 -1128 9477 -1118
rect 9557 -1061 9757 -1050
rect 9557 -1117 9578 -1061
rect 9634 -1117 9688 -1061
rect 9744 -1117 9757 -1061
rect 9557 -1127 9757 -1117
rect 6874 -1356 7432 -1307
rect 8242 -1356 8800 -1307
rect 5917 -1367 6117 -1357
rect 5917 -1423 5932 -1367
rect 5988 -1423 6042 -1367
rect 6098 -1423 6117 -1367
rect 5917 -1435 6117 -1423
rect 6197 -1373 6397 -1360
rect 6197 -1429 6212 -1373
rect 6268 -1429 6322 -1373
rect 6378 -1429 6397 -1373
rect 6197 -1437 6397 -1429
rect 6874 -1366 7517 -1356
rect 7610 -1360 7666 -1358
rect 8008 -1360 8064 -1358
rect 6874 -1379 7331 -1366
rect 5913 -1518 6091 -1517
rect 5901 -1523 6091 -1518
rect 5901 -1579 5913 -1523
rect 5969 -1579 6023 -1523
rect 6079 -1579 6091 -1523
rect 5901 -1583 6091 -1579
rect 6318 -1585 6384 -1437
rect 6312 -1588 6504 -1585
rect 6312 -1644 6324 -1588
rect 6380 -1644 6434 -1588
rect 6490 -1644 6504 -1588
rect 6312 -1647 6504 -1644
rect 5927 -1702 5983 -1699
rect 5917 -1704 6117 -1702
rect 6874 -1703 6946 -1379
rect 7317 -1422 7331 -1379
rect 7387 -1422 7441 -1366
rect 7497 -1422 7517 -1366
rect 7317 -1436 7517 -1422
rect 7597 -1368 7797 -1360
rect 7597 -1424 7610 -1368
rect 7666 -1424 7720 -1368
rect 7776 -1424 7797 -1368
rect 7597 -1437 7797 -1424
rect 7877 -1368 8077 -1360
rect 7877 -1424 7898 -1368
rect 7954 -1424 8008 -1368
rect 8064 -1424 8077 -1368
rect 7877 -1437 8077 -1424
rect 8157 -1366 8800 -1356
rect 8157 -1422 8177 -1366
rect 8233 -1422 8287 -1366
rect 8343 -1379 8800 -1366
rect 8343 -1422 8357 -1379
rect 8157 -1436 8357 -1422
rect 5665 -1709 6117 -1704
rect 5665 -1765 5929 -1709
rect 5985 -1765 6037 -1709
rect 6093 -1765 6117 -1709
rect 5665 -1770 6117 -1765
rect 5077 -1779 5277 -1770
rect 5917 -1779 6117 -1770
rect 6477 -1716 6677 -1703
rect 6477 -1772 6490 -1716
rect 6546 -1772 6600 -1716
rect 6656 -1772 6677 -1716
rect 6477 -1780 6677 -1772
rect 6757 -1713 6957 -1703
rect 6757 -1769 6771 -1713
rect 6827 -1769 6881 -1713
rect 6937 -1769 6957 -1713
rect 6757 -1780 6957 -1769
rect 7317 -1710 7517 -1703
rect 7317 -1766 7329 -1710
rect 7385 -1766 7439 -1710
rect 7495 -1766 7517 -1710
rect 7317 -1780 7517 -1766
rect 4648 -1782 4704 -1780
rect 6490 -1782 6546 -1780
rect 4237 -2024 4437 -2012
rect 4237 -2080 4257 -2024
rect 4313 -2080 4367 -2024
rect 4423 -2080 4437 -2024
rect 4237 -2089 4437 -2080
rect 6757 -2024 6957 -2012
rect 6757 -2080 6771 -2024
rect 6827 -2080 6881 -2024
rect 6937 -2080 6957 -2024
rect 6757 -2089 6957 -2080
rect 4367 -2090 4423 -2089
rect 6771 -2090 6827 -2089
rect 7604 -2131 7670 -1437
rect 8004 -2131 8070 -1437
rect 8728 -1703 8800 -1379
rect 9277 -1373 9477 -1360
rect 9277 -1429 9296 -1373
rect 9352 -1429 9406 -1373
rect 9462 -1429 9477 -1373
rect 9277 -1437 9477 -1429
rect 9557 -1367 9757 -1357
rect 9557 -1423 9576 -1367
rect 9632 -1423 9686 -1367
rect 9742 -1423 9757 -1367
rect 9557 -1435 9757 -1423
rect 9290 -1585 9356 -1437
rect 9581 -1522 9771 -1517
rect 9581 -1578 9593 -1522
rect 9649 -1578 9703 -1522
rect 9759 -1578 9771 -1522
rect 9581 -1583 9771 -1578
rect 9170 -1588 9362 -1585
rect 9170 -1644 9184 -1588
rect 9240 -1644 9294 -1588
rect 9350 -1644 9362 -1588
rect 9170 -1647 9362 -1644
rect 9691 -1702 9747 -1699
rect 8157 -1710 8357 -1703
rect 8157 -1766 8179 -1710
rect 8235 -1766 8289 -1710
rect 8345 -1766 8357 -1710
rect 8157 -1780 8357 -1766
rect 8717 -1713 8917 -1703
rect 8717 -1769 8737 -1713
rect 8793 -1769 8847 -1713
rect 8903 -1769 8917 -1713
rect 8717 -1780 8917 -1769
rect 8997 -1716 9197 -1703
rect 8997 -1772 9018 -1716
rect 9074 -1772 9128 -1716
rect 9184 -1772 9197 -1716
rect 8997 -1780 9197 -1772
rect 9557 -1704 9757 -1702
rect 9943 -1704 10009 -355
rect 11063 -302 11066 -296
rect 11122 -302 11127 -246
rect 11063 -356 11127 -302
rect 10196 -417 11005 -401
rect 10196 -467 10947 -417
rect 10196 -500 10262 -467
rect 10065 -505 10262 -500
rect 10065 -561 10083 -505
rect 10139 -561 10193 -505
rect 10249 -561 10262 -505
rect 10065 -566 10262 -561
rect 10942 -473 10947 -467
rect 11003 -473 11005 -417
rect 11063 -412 11066 -356
rect 11122 -412 11127 -356
rect 11063 -427 11127 -412
rect 10942 -527 11005 -473
rect 10137 -827 10203 -566
rect 10942 -583 10947 -527
rect 11003 -583 11005 -527
rect 10942 -598 11005 -583
rect 10315 -608 10879 -603
rect 10315 -664 10333 -608
rect 10389 -664 10443 -608
rect 10499 -619 10879 -608
rect 10499 -664 10818 -619
rect 10315 -669 10818 -664
rect 10813 -675 10818 -669
rect 10874 -675 10879 -619
rect 10813 -729 10879 -675
rect 10813 -785 10818 -729
rect 10874 -785 10879 -729
rect 10813 -800 10879 -785
rect 10066 -832 10263 -827
rect 10066 -888 10084 -832
rect 10140 -888 10194 -832
rect 10250 -888 10263 -832
rect 10066 -893 10263 -888
rect 10704 -1158 10767 -1141
rect 10704 -1214 10709 -1158
rect 10765 -1214 10767 -1158
rect 10704 -1249 10767 -1214
rect 10067 -1254 10893 -1249
rect 10067 -1310 10085 -1254
rect 10141 -1310 10195 -1254
rect 10251 -1268 10893 -1254
rect 10251 -1310 10709 -1268
rect 10067 -1315 10709 -1310
rect 10704 -1324 10709 -1315
rect 10765 -1315 10893 -1268
rect 10765 -1324 10767 -1315
rect 10704 -1339 10767 -1324
rect 10282 -1590 10479 -1585
rect 10282 -1646 10295 -1590
rect 10353 -1646 10405 -1590
rect 10463 -1646 10479 -1590
rect 10282 -1651 10479 -1646
rect 9557 -1709 10009 -1704
rect 9557 -1765 9581 -1709
rect 9637 -1765 9689 -1709
rect 9745 -1765 10009 -1709
rect 9557 -1770 10009 -1765
rect 9557 -1779 9757 -1770
rect 9128 -1782 9184 -1780
rect 8717 -2024 8917 -2012
rect 8717 -2080 8737 -2024
rect 8793 -2080 8847 -2024
rect 8903 -2080 8917 -2024
rect 8717 -2089 8917 -2080
rect 8847 -2090 8903 -2089
rect 3036 -2135 3226 -2131
rect 3036 -2191 3048 -2135
rect 3104 -2191 3158 -2135
rect 3214 -2191 3226 -2135
rect 3036 -2195 3226 -2191
rect 3488 -2135 3678 -2131
rect 3488 -2191 3500 -2135
rect 3556 -2191 3610 -2135
rect 3666 -2191 3678 -2135
rect 3488 -2195 3678 -2191
rect 7516 -2135 7706 -2131
rect 7516 -2191 7528 -2135
rect 7584 -2191 7638 -2135
rect 7694 -2191 7706 -2135
rect 7516 -2195 7706 -2191
rect 7968 -2135 8158 -2131
rect 7968 -2191 7980 -2135
rect 8036 -2191 8090 -2135
rect 8146 -2191 8158 -2135
rect 7968 -2195 8158 -2191
<< via2 >>
rect 2291 2024 2347 2080
rect 2401 2024 2457 2080
rect 691 1254 747 1310
rect 801 1254 857 1310
rect 683 608 739 664
rect 793 608 849 664
rect 2010 1716 2066 1772
rect 2120 1716 2176 1772
rect 2849 1710 2905 1766
rect 2959 1710 3015 1766
rect 1433 1523 1489 1579
rect 1543 1523 1599 1579
rect 1452 1367 1508 1423
rect 1562 1367 1618 1423
rect 4257 2024 4313 2080
rect 4367 2024 4423 2080
rect 6771 2024 6827 2080
rect 6881 2024 6937 2080
rect 3699 1710 3755 1766
rect 3809 1710 3865 1766
rect 4538 1716 4594 1772
rect 4648 1716 4704 1772
rect 5113 1522 5169 1578
rect 5223 1522 5279 1578
rect 1450 1061 1506 1117
rect 1560 1061 1616 1117
rect 5096 1367 5152 1423
rect 5206 1367 5262 1423
rect 5098 1061 5154 1117
rect 5208 1061 5264 1117
rect 1450 719 1506 775
rect 1560 719 1616 775
rect 2011 718 2067 774
rect 2121 718 2177 774
rect 4537 718 4593 774
rect 4647 718 4703 774
rect 5098 719 5154 775
rect 5208 719 5264 775
rect 1452 416 1508 472
rect 1562 416 1618 472
rect 2010 418 2066 474
rect 2120 418 2176 474
rect 6490 1716 6546 1772
rect 6600 1716 6656 1772
rect 7329 1710 7385 1766
rect 7439 1710 7495 1766
rect 5913 1523 5969 1579
rect 6023 1523 6079 1579
rect 5932 1367 5988 1423
rect 6042 1367 6098 1423
rect 8737 2024 8793 2080
rect 8847 2024 8903 2080
rect 8179 1710 8235 1766
rect 8289 1710 8345 1766
rect 9018 1716 9074 1772
rect 9128 1716 9184 1772
rect 9593 1522 9649 1578
rect 9703 1522 9759 1578
rect 9576 1367 9632 1423
rect 9686 1367 9742 1423
rect 5930 1061 5986 1117
rect 6040 1061 6096 1117
rect 9578 1061 9634 1117
rect 9688 1061 9744 1117
rect 5930 719 5986 775
rect 6040 719 6096 775
rect 6491 718 6547 774
rect 6601 718 6657 774
rect 9017 718 9073 774
rect 9127 718 9183 774
rect 9578 719 9634 775
rect 9688 719 9744 775
rect 10295 1590 10351 1646
rect 10405 1590 10461 1646
rect 10333 608 10389 664
rect 10443 608 10499 664
rect 683 -664 739 -608
rect 793 -664 849 -608
rect 691 -1310 747 -1254
rect 801 -1310 857 -1254
rect 1452 -472 1508 -416
rect 1562 -472 1618 -416
rect 2010 -474 2066 -418
rect 2120 -474 2176 -418
rect 1450 -775 1506 -719
rect 1560 -775 1616 -719
rect 2011 -774 2067 -718
rect 2121 -774 2177 -718
rect 4537 -774 4593 -718
rect 4647 -774 4703 -718
rect 5098 -775 5154 -719
rect 5208 -775 5264 -719
rect 1450 -1117 1506 -1061
rect 1560 -1117 1616 -1061
rect 1452 -1423 1508 -1367
rect 1562 -1423 1618 -1367
rect 5098 -1117 5154 -1061
rect 5208 -1117 5264 -1061
rect 1433 -1579 1489 -1523
rect 1543 -1579 1599 -1523
rect 2010 -1772 2066 -1716
rect 2120 -1772 2176 -1716
rect 2849 -1766 2905 -1710
rect 2959 -1766 3015 -1710
rect 2291 -2080 2347 -2024
rect 2401 -2080 2457 -2024
rect 5096 -1423 5152 -1367
rect 5206 -1423 5262 -1367
rect 5113 -1578 5169 -1522
rect 5223 -1578 5279 -1522
rect 3699 -1766 3755 -1710
rect 3809 -1766 3865 -1710
rect 4538 -1772 4594 -1716
rect 4648 -1772 4704 -1716
rect 5930 -775 5986 -719
rect 6040 -775 6096 -719
rect 6491 -774 6547 -718
rect 6601 -774 6657 -718
rect 9017 -774 9073 -718
rect 9127 -774 9183 -718
rect 9578 -775 9634 -719
rect 9688 -775 9744 -719
rect 5930 -1117 5986 -1061
rect 6040 -1117 6096 -1061
rect 9578 -1117 9634 -1061
rect 9688 -1117 9744 -1061
rect 5932 -1423 5988 -1367
rect 6042 -1423 6098 -1367
rect 5913 -1579 5969 -1523
rect 6023 -1579 6079 -1523
rect 6490 -1772 6546 -1716
rect 6600 -1772 6656 -1716
rect 7329 -1766 7385 -1710
rect 7439 -1766 7495 -1710
rect 4257 -2080 4313 -2024
rect 4367 -2080 4423 -2024
rect 6771 -2080 6827 -2024
rect 6881 -2080 6937 -2024
rect 9576 -1423 9632 -1367
rect 9686 -1423 9742 -1367
rect 9593 -1578 9649 -1522
rect 9703 -1578 9759 -1522
rect 8179 -1766 8235 -1710
rect 8289 -1766 8345 -1710
rect 9018 -1772 9074 -1716
rect 9128 -1772 9184 -1716
rect 10333 -664 10389 -608
rect 10443 -664 10499 -608
rect 10295 -1646 10351 -1590
rect 10405 -1646 10461 -1590
rect 8737 -2080 8793 -2024
rect 8847 -2080 8903 -2024
<< metal3 >>
rect 2277 2080 2477 2089
rect 2277 2024 2291 2080
rect 2347 2024 2401 2080
rect 2457 2024 2477 2080
rect 2277 2012 2477 2024
rect 4237 2080 4437 2089
rect 4237 2024 4257 2080
rect 4313 2024 4367 2080
rect 4423 2024 4437 2080
rect 4237 2012 4437 2024
rect 6757 2080 6957 2089
rect 6757 2024 6771 2080
rect 6827 2024 6881 2080
rect 6937 2024 6957 2080
rect 6757 2012 6957 2024
rect 8717 2080 8917 2089
rect 8717 2024 8737 2080
rect 8793 2024 8847 2080
rect 8903 2024 8917 2080
rect 8717 2012 8917 2024
rect 1997 1772 2197 1780
rect 1997 1716 2010 1772
rect 2066 1716 2120 1772
rect 2176 1716 2197 1772
rect 1997 1703 2197 1716
rect 2042 1583 2108 1703
rect 1295 1579 2108 1583
rect 1295 1523 1433 1579
rect 1489 1523 1543 1579
rect 1599 1523 2108 1579
rect 1295 1517 2108 1523
rect 1437 1423 1637 1435
rect 1437 1367 1452 1423
rect 1508 1367 1562 1423
rect 1618 1389 1637 1423
rect 1618 1367 1639 1389
rect 1437 1357 1639 1367
rect 1514 1347 1639 1357
rect 2290 1347 2354 2012
rect 2837 1766 3037 1780
rect 2837 1710 2849 1766
rect 2905 1710 2959 1766
rect 3015 1710 3037 1766
rect 2837 1703 3037 1710
rect 3677 1766 3877 1780
rect 3677 1710 3699 1766
rect 3755 1710 3809 1766
rect 3865 1710 3877 1766
rect 3677 1703 3877 1710
rect 678 1310 875 1315
rect 678 1254 691 1310
rect 747 1254 801 1310
rect 857 1254 875 1310
rect 678 1249 875 1254
rect 1514 1283 2354 1347
rect 742 669 808 1249
rect 1514 1127 1598 1283
rect 1437 1117 1637 1127
rect 1437 1061 1450 1117
rect 1506 1061 1560 1117
rect 1616 1061 1637 1117
rect 1437 1050 1637 1061
rect 1564 965 1637 1050
rect 1564 892 2096 965
rect 2023 785 2096 892
rect 1437 775 1637 785
rect 1437 719 1450 775
rect 1506 719 1560 775
rect 1616 719 1637 775
rect 1437 708 1637 719
rect 1997 774 2197 785
rect 1997 718 2011 774
rect 2067 718 2121 774
rect 2177 718 2197 774
rect 1997 708 2197 718
rect 670 664 867 669
rect 670 608 683 664
rect 739 608 793 664
rect 849 608 867 664
rect 670 603 867 608
rect 1536 652 1637 708
rect 2934 652 3000 1703
rect 1536 586 3000 652
rect 3714 652 3780 1703
rect 4360 1347 4424 2012
rect 4517 1772 4717 1780
rect 4517 1716 4538 1772
rect 4594 1716 4648 1772
rect 4704 1716 4717 1772
rect 4517 1703 4717 1716
rect 6477 1772 6677 1780
rect 6477 1716 6490 1772
rect 6546 1716 6600 1772
rect 6656 1716 6677 1772
rect 6477 1703 6677 1716
rect 4606 1583 4672 1703
rect 6522 1583 6588 1703
rect 4606 1578 5291 1583
rect 4606 1522 5113 1578
rect 5169 1522 5223 1578
rect 5279 1522 5291 1578
rect 4606 1517 5291 1522
rect 5775 1579 6588 1583
rect 5775 1523 5913 1579
rect 5969 1523 6023 1579
rect 6079 1523 6588 1579
rect 5775 1517 6588 1523
rect 5077 1423 5277 1435
rect 5077 1367 5096 1423
rect 5152 1367 5206 1423
rect 5262 1367 5277 1423
rect 5077 1357 5277 1367
rect 5917 1423 6117 1435
rect 5917 1367 5932 1423
rect 5988 1367 6042 1423
rect 6098 1367 6117 1423
rect 5917 1357 6117 1367
rect 5077 1347 5189 1357
rect 4360 1283 5189 1347
rect 6002 1347 6117 1357
rect 6770 1347 6834 2012
rect 7317 1766 7517 1780
rect 7317 1710 7329 1766
rect 7385 1710 7439 1766
rect 7495 1710 7517 1766
rect 7317 1703 7517 1710
rect 8157 1766 8357 1780
rect 8157 1710 8179 1766
rect 8235 1710 8289 1766
rect 8345 1710 8357 1766
rect 8157 1703 8357 1710
rect 6002 1283 6834 1347
rect 5077 1117 5277 1127
rect 5077 1061 5098 1117
rect 5154 1061 5208 1117
rect 5264 1061 5277 1117
rect 5077 1050 5277 1061
rect 5917 1117 6117 1127
rect 5917 1061 5930 1117
rect 5986 1061 6040 1117
rect 6096 1061 6117 1117
rect 5917 1050 6117 1061
rect 5077 965 5150 1050
rect 4618 892 5150 965
rect 6044 965 6117 1050
rect 6044 892 6576 965
rect 4618 785 4691 892
rect 6503 785 6576 892
rect 4517 774 4717 785
rect 4517 718 4537 774
rect 4593 718 4647 774
rect 4703 718 4717 774
rect 4517 708 4717 718
rect 5077 775 5277 785
rect 5077 719 5098 775
rect 5154 719 5208 775
rect 5264 719 5277 775
rect 5077 708 5277 719
rect 5917 775 6117 785
rect 5917 719 5930 775
rect 5986 719 6040 775
rect 6096 719 6117 775
rect 5917 708 6117 719
rect 6477 774 6677 785
rect 6477 718 6491 774
rect 6547 718 6601 774
rect 6657 718 6677 774
rect 6477 708 6677 718
rect 5077 652 5178 708
rect 3714 586 5178 652
rect 6016 652 6117 708
rect 7414 652 7480 1703
rect 6016 586 7480 652
rect 8194 652 8260 1703
rect 8840 1347 8904 2012
rect 8997 1772 9197 1780
rect 8997 1716 9018 1772
rect 9074 1716 9128 1772
rect 9184 1716 9197 1772
rect 8997 1703 9197 1716
rect 9086 1583 9152 1703
rect 10282 1646 10479 1651
rect 10282 1590 10295 1646
rect 10351 1590 10405 1646
rect 10461 1590 10479 1646
rect 10282 1585 10479 1590
rect 9086 1578 9771 1583
rect 9086 1522 9593 1578
rect 9649 1522 9703 1578
rect 9759 1522 9771 1578
rect 9086 1517 9771 1522
rect 9557 1423 9757 1435
rect 9557 1367 9576 1423
rect 9632 1367 9686 1423
rect 9742 1367 9757 1423
rect 9557 1357 9757 1367
rect 9557 1347 9669 1357
rect 8840 1283 9669 1347
rect 9557 1117 9757 1127
rect 9557 1061 9578 1117
rect 9634 1061 9688 1117
rect 9744 1061 9757 1117
rect 9557 1050 9757 1061
rect 9557 965 9630 1050
rect 9098 892 9630 965
rect 9098 785 9171 892
rect 8997 774 9197 785
rect 8997 718 9017 774
rect 9073 718 9127 774
rect 9183 718 9197 774
rect 8997 708 9197 718
rect 9557 775 9757 785
rect 9557 719 9578 775
rect 9634 719 9688 775
rect 9744 719 9757 775
rect 9557 708 9757 719
rect 9557 652 9658 708
rect 10383 669 10449 1585
rect 8194 586 9658 652
rect 10320 664 10517 669
rect 10320 608 10333 664
rect 10389 608 10443 664
rect 10499 608 10517 664
rect 10320 603 10517 608
rect 1536 477 1637 586
rect 1439 472 1637 477
rect 1439 416 1452 472
rect 1508 416 1562 472
rect 1618 448 1637 472
rect 1997 474 2194 479
rect 1618 416 1636 448
rect 1439 411 1636 416
rect 1997 418 2010 474
rect 2066 418 2120 474
rect 2176 418 2194 474
rect 1997 413 2194 418
rect 1439 -416 1636 -411
rect 1439 -472 1452 -416
rect 1508 -472 1562 -416
rect 1618 -448 1636 -416
rect 1997 -418 2194 -413
rect 1618 -472 1637 -448
rect 1439 -477 1637 -472
rect 1536 -586 1637 -477
rect 1997 -474 2010 -418
rect 2066 -474 2120 -418
rect 2176 -474 2194 -418
rect 1997 -479 2194 -474
rect 670 -608 867 -603
rect 670 -664 683 -608
rect 739 -664 793 -608
rect 849 -664 867 -608
rect 670 -669 867 -664
rect 1536 -652 3000 -586
rect 742 -1249 808 -669
rect 1536 -708 1637 -652
rect 1437 -719 1637 -708
rect 1437 -775 1450 -719
rect 1506 -775 1560 -719
rect 1616 -775 1637 -719
rect 1437 -785 1637 -775
rect 1997 -718 2197 -708
rect 1997 -774 2011 -718
rect 2067 -774 2121 -718
rect 2177 -774 2197 -718
rect 1997 -785 2197 -774
rect 2023 -892 2096 -785
rect 1564 -965 2096 -892
rect 1564 -1050 1637 -965
rect 1437 -1061 1637 -1050
rect 1437 -1117 1450 -1061
rect 1506 -1117 1560 -1061
rect 1616 -1117 1637 -1061
rect 1437 -1127 1637 -1117
rect 678 -1254 875 -1249
rect 678 -1310 691 -1254
rect 747 -1310 801 -1254
rect 857 -1310 875 -1254
rect 678 -1315 875 -1310
rect 1514 -1283 1598 -1127
rect 1514 -1347 2354 -1283
rect 1514 -1357 1639 -1347
rect 1437 -1367 1639 -1357
rect 1437 -1423 1452 -1367
rect 1508 -1423 1562 -1367
rect 1618 -1389 1639 -1367
rect 1618 -1423 1637 -1389
rect 1437 -1435 1637 -1423
rect 1295 -1523 2108 -1517
rect 1295 -1579 1433 -1523
rect 1489 -1579 1543 -1523
rect 1599 -1579 2108 -1523
rect 1295 -1583 2108 -1579
rect 2042 -1703 2108 -1583
rect 1997 -1716 2197 -1703
rect 1997 -1772 2010 -1716
rect 2066 -1772 2120 -1716
rect 2176 -1772 2197 -1716
rect 1997 -1780 2197 -1772
rect 2290 -2012 2354 -1347
rect 2934 -1703 3000 -652
rect 3714 -652 5178 -586
rect 3714 -1703 3780 -652
rect 5077 -708 5178 -652
rect 6016 -652 7480 -586
rect 6016 -708 6117 -652
rect 4517 -718 4717 -708
rect 4517 -774 4537 -718
rect 4593 -774 4647 -718
rect 4703 -774 4717 -718
rect 4517 -785 4717 -774
rect 5077 -719 5277 -708
rect 5077 -775 5098 -719
rect 5154 -775 5208 -719
rect 5264 -775 5277 -719
rect 5077 -785 5277 -775
rect 5917 -719 6117 -708
rect 5917 -775 5930 -719
rect 5986 -775 6040 -719
rect 6096 -775 6117 -719
rect 5917 -785 6117 -775
rect 6477 -718 6677 -708
rect 6477 -774 6491 -718
rect 6547 -774 6601 -718
rect 6657 -774 6677 -718
rect 6477 -785 6677 -774
rect 4618 -892 4691 -785
rect 6503 -892 6576 -785
rect 4618 -965 5150 -892
rect 5077 -1050 5150 -965
rect 6044 -965 6576 -892
rect 6044 -1050 6117 -965
rect 5077 -1061 5277 -1050
rect 5077 -1117 5098 -1061
rect 5154 -1117 5208 -1061
rect 5264 -1117 5277 -1061
rect 5077 -1127 5277 -1117
rect 5917 -1061 6117 -1050
rect 5917 -1117 5930 -1061
rect 5986 -1117 6040 -1061
rect 6096 -1117 6117 -1061
rect 5917 -1127 6117 -1117
rect 4360 -1347 5189 -1283
rect 2837 -1710 3037 -1703
rect 2837 -1766 2849 -1710
rect 2905 -1766 2959 -1710
rect 3015 -1766 3037 -1710
rect 2837 -1780 3037 -1766
rect 3677 -1710 3877 -1703
rect 3677 -1766 3699 -1710
rect 3755 -1766 3809 -1710
rect 3865 -1766 3877 -1710
rect 3677 -1780 3877 -1766
rect 4360 -2012 4424 -1347
rect 5077 -1357 5189 -1347
rect 6002 -1347 6834 -1283
rect 6002 -1357 6117 -1347
rect 5077 -1367 5277 -1357
rect 5077 -1423 5096 -1367
rect 5152 -1423 5206 -1367
rect 5262 -1423 5277 -1367
rect 5077 -1435 5277 -1423
rect 5917 -1367 6117 -1357
rect 5917 -1423 5932 -1367
rect 5988 -1423 6042 -1367
rect 6098 -1423 6117 -1367
rect 5917 -1435 6117 -1423
rect 4606 -1522 5291 -1517
rect 4606 -1578 5113 -1522
rect 5169 -1578 5223 -1522
rect 5279 -1578 5291 -1522
rect 4606 -1583 5291 -1578
rect 5775 -1523 6588 -1517
rect 5775 -1579 5913 -1523
rect 5969 -1579 6023 -1523
rect 6079 -1579 6588 -1523
rect 5775 -1583 6588 -1579
rect 4606 -1703 4672 -1583
rect 6522 -1703 6588 -1583
rect 4517 -1716 4717 -1703
rect 4517 -1772 4538 -1716
rect 4594 -1772 4648 -1716
rect 4704 -1772 4717 -1716
rect 4517 -1780 4717 -1772
rect 6477 -1716 6677 -1703
rect 6477 -1772 6490 -1716
rect 6546 -1772 6600 -1716
rect 6656 -1772 6677 -1716
rect 6477 -1780 6677 -1772
rect 6770 -2012 6834 -1347
rect 7414 -1703 7480 -652
rect 8194 -652 9658 -586
rect 8194 -1703 8260 -652
rect 9557 -708 9658 -652
rect 10320 -608 10517 -603
rect 10320 -664 10333 -608
rect 10389 -664 10443 -608
rect 10499 -664 10517 -608
rect 10320 -669 10517 -664
rect 8997 -718 9197 -708
rect 8997 -774 9017 -718
rect 9073 -774 9127 -718
rect 9183 -774 9197 -718
rect 8997 -785 9197 -774
rect 9557 -719 9757 -708
rect 9557 -775 9578 -719
rect 9634 -775 9688 -719
rect 9744 -775 9757 -719
rect 9557 -785 9757 -775
rect 9098 -892 9171 -785
rect 9098 -965 9630 -892
rect 9557 -1050 9630 -965
rect 9557 -1061 9757 -1050
rect 9557 -1117 9578 -1061
rect 9634 -1117 9688 -1061
rect 9744 -1117 9757 -1061
rect 9557 -1127 9757 -1117
rect 8840 -1347 9669 -1283
rect 7317 -1710 7517 -1703
rect 7317 -1766 7329 -1710
rect 7385 -1766 7439 -1710
rect 7495 -1766 7517 -1710
rect 7317 -1780 7517 -1766
rect 8157 -1710 8357 -1703
rect 8157 -1766 8179 -1710
rect 8235 -1766 8289 -1710
rect 8345 -1766 8357 -1710
rect 8157 -1780 8357 -1766
rect 8840 -2012 8904 -1347
rect 9557 -1357 9669 -1347
rect 9557 -1367 9757 -1357
rect 9557 -1423 9576 -1367
rect 9632 -1423 9686 -1367
rect 9742 -1423 9757 -1367
rect 9557 -1435 9757 -1423
rect 9086 -1522 9771 -1517
rect 9086 -1578 9593 -1522
rect 9649 -1578 9703 -1522
rect 9759 -1578 9771 -1522
rect 9086 -1583 9771 -1578
rect 9086 -1703 9152 -1583
rect 10383 -1585 10449 -669
rect 10282 -1590 10479 -1585
rect 10282 -1646 10295 -1590
rect 10351 -1646 10405 -1590
rect 10461 -1646 10479 -1590
rect 10282 -1651 10479 -1646
rect 8997 -1716 9197 -1703
rect 8997 -1772 9018 -1716
rect 9074 -1772 9128 -1716
rect 9184 -1772 9197 -1716
rect 8997 -1780 9197 -1772
rect 2277 -2024 2477 -2012
rect 2277 -2080 2291 -2024
rect 2347 -2080 2401 -2024
rect 2457 -2080 2477 -2024
rect 2277 -2089 2477 -2080
rect 4237 -2024 4437 -2012
rect 4237 -2080 4257 -2024
rect 4313 -2080 4367 -2024
rect 4423 -2080 4437 -2024
rect 4237 -2089 4437 -2080
rect 6757 -2024 6957 -2012
rect 6757 -2080 6771 -2024
rect 6827 -2080 6881 -2024
rect 6937 -2080 6957 -2024
rect 6757 -2089 6957 -2080
rect 8717 -2024 8917 -2012
rect 8717 -2080 8737 -2024
rect 8793 -2080 8847 -2024
rect 8903 -2080 8917 -2024
rect 8717 -2089 8917 -2080
<< labels >>
flabel metal1 4375 0 4384 9 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel metal1 257 743 257 743 0 FreeSans 1600 0 0 0 A
port 3 nsew
flabel metal1 381 686 381 686 0 FreeSans 1600 0 0 0 C
port 5 nsew
flabel metal1 140 454 140 454 0 FreeSans 1600 0 0 0 E
port 7 nsew
flabel metal1 32 -46 32 -46 0 FreeSans 1600 0 0 0 G
port 9 nsew
flabel metal1 10741 970 10741 970 0 FreeSans 1600 0 0 0 B
port 11 nsew
flabel metal1 10848 530 10848 530 0 FreeSans 1600 0 0 0 D
port 13 nsew
flabel metal1 10942 -417 11005 417 0 FreeSans 1600 0 0 0 F
port 14 nsew
flabel metal1 11103 -145 11103 -145 0 FreeSans 1600 0 0 0 H
port 15 nsew
flabel metal2 396 -856 396 -856 0 FreeSans 800 0 0 0 pag_res_magic_0.E
flabel metal2 10704 -622 10704 -622 0 FreeSans 800 0 0 0 pag_res_magic_0.D
flabel metal2 10695 -427 10695 -427 0 FreeSans 800 0 0 0 pag_res_magic_0.F
flabel metal2 10708 -257 10708 -257 0 FreeSans 800 0 0 0 pag_res_magic_0.H
flabel via1 375 -1273 375 -1273 0 FreeSans 800 0 0 0 pag_res_magic_0.C
flabel metal2 362 -261 362 -261 0 FreeSans 800 0 0 0 pag_res_magic_0.G
flabel metal2 10874 -1273 10874 -1273 0 FreeSans 800 0 0 0 pag_res_magic_0.B
flabel metal2 344 -969 344 -969 0 FreeSans 800 0 0 0 pag_res_magic_0.A
flabel metal1 5237 -2348 5237 -2348 0 FreeSans 1280 0 0 0 pag_res_magic_0.VDD
flabel metal2 396 856 396 856 0 FreeSans 800 0 0 0 pag_res_magic_1.E
flabel metal2 10704 622 10704 622 0 FreeSans 800 0 0 0 pag_res_magic_1.D
flabel metal2 10695 427 10695 427 0 FreeSans 800 0 0 0 pag_res_magic_1.F
flabel metal2 10708 257 10708 257 0 FreeSans 800 0 0 0 pag_res_magic_1.H
flabel via1 375 1273 375 1273 0 FreeSans 800 0 0 0 pag_res_magic_1.C
flabel metal2 362 261 362 261 0 FreeSans 800 0 0 0 pag_res_magic_1.G
flabel metal2 10874 1273 10874 1273 0 FreeSans 800 0 0 0 pag_res_magic_1.B
flabel metal2 344 969 344 969 0 FreeSans 800 0 0 0 pag_res_magic_1.A
flabel metal1 5237 2348 5237 2348 0 FreeSans 1280 0 0 0 pag_res_magic_1.VDD
<< end >>
