magic
tech gf180mcuC
magscale 1 10
timestamp 1692946346
<< pwell >>
rect 114 269 195 310
rect 3095 69 3144 170
rect 4933 20 4979 81
rect 1854 -190 1933 -149
rect 5124 -189 5202 -109
rect 520 -405 620 -365
rect 1132 -405 1232 -365
rect 1336 -405 1436 -365
rect 1948 -405 2048 -365
rect 2152 -405 2252 -365
rect 2764 -405 2864 -365
rect 2968 -405 3068 -365
rect 3580 -405 3680 -365
rect 3784 -404 3884 -364
rect 326 -446 405 -405
rect 530 -445 609 -405
rect 1142 -445 1221 -405
rect 1346 -445 1425 -405
rect 1958 -445 2037 -405
rect 2162 -445 2241 -405
rect 2774 -446 2853 -405
rect 2978 -446 3057 -405
rect 3590 -446 3669 -405
rect 3794 -445 3873 -404
rect 4396 -405 4496 -365
rect 4600 -405 4700 -365
rect 4406 -446 4485 -405
rect 5212 -406 5312 -366
rect 5416 -406 5516 -366
rect 6028 -406 6128 -366
rect 4609 -447 4688 -406
rect 5228 -408 5306 -406
rect 6232 -407 6332 -367
rect 5222 -448 5306 -408
rect 5425 -448 5507 -410
rect 6038 -448 6119 -410
rect 6243 -448 6324 -410
<< ndiff >>
rect 3095 69 3144 170
<< polysilicon >>
rect 84 306 210 345
rect 84 255 100 306
rect 151 290 210 306
rect 724 343 824 356
rect 724 290 744 343
rect 792 290 824 343
rect 151 255 212 290
rect 84 242 212 255
rect 86 241 212 242
rect 112 188 212 241
rect 724 190 824 290
rect 928 346 1028 360
rect 928 285 947 346
rect 1010 285 1028 346
rect 928 190 1028 285
rect 1540 348 1640 361
rect 1540 285 1558 348
rect 1617 285 1640 348
rect 1540 190 1640 285
rect 1744 347 1844 361
rect 1744 287 1764 347
rect 1826 287 1844 347
rect 1744 190 1844 287
rect 2356 349 2456 365
rect 2356 286 2372 349
rect 2440 286 2456 349
rect 2356 190 2456 286
rect 2560 349 2660 366
rect 2560 285 2577 349
rect 2640 285 2660 349
rect 2560 190 2660 285
rect 3172 350 3272 364
rect 3172 286 3188 350
rect 3256 286 3272 350
rect 3172 190 3272 286
rect 3376 352 3476 365
rect 3376 283 3389 352
rect 3461 283 3476 352
rect 3376 190 3476 283
rect 3988 350 4088 365
rect 3988 284 4004 350
rect 4069 284 4088 350
rect 3988 190 4088 284
rect 4192 349 4292 365
rect 4192 284 4207 349
rect 4274 284 4292 349
rect 4192 190 4292 284
rect 4804 341 4904 354
rect 4804 286 4825 341
rect 4883 286 4904 341
rect 4804 190 4904 286
rect 5008 340 5105 355
rect 5008 285 5030 340
rect 5088 290 5105 340
rect 5620 349 5720 362
rect 5831 353 5918 361
rect 5620 294 5643 349
rect 5701 294 5720 349
rect 5088 285 5108 290
rect 5008 232 5108 285
rect 5008 188 5105 232
rect 5620 190 5720 294
rect 5824 347 5924 353
rect 5824 293 5846 347
rect 5904 293 5924 347
rect 5824 190 5924 293
rect 6456 340 6537 356
rect 6456 291 6472 340
rect 6518 291 6537 340
rect 6456 290 6537 291
rect 6436 280 6537 290
rect 6436 232 6536 280
rect 316 26 393 68
rect 316 -31 416 24
rect 520 -31 620 24
rect 1132 -31 1232 24
rect 1336 -31 1436 24
rect 1948 -31 2048 24
rect 2152 -31 2252 24
rect 2764 -31 2864 24
rect 2968 -31 3068 24
rect 3580 -31 3680 25
rect 3784 -31 3884 24
rect 4396 -31 4496 25
rect 4600 -31 4700 27
rect 5212 -31 5312 24
rect 5416 -31 5516 27
rect 6028 -31 6128 27
rect 6232 -31 6332 29
rect 112 -85 6536 -31
rect 62 -99 6536 -85
rect 62 -150 76 -99
rect 127 -108 6536 -99
rect 127 -150 212 -108
rect 62 -164 212 -150
rect 112 -173 212 -164
rect 724 -173 824 -108
rect 928 -173 1028 -108
rect 1540 -173 1640 -108
rect 1744 -173 1844 -108
rect 2356 -173 2456 -108
rect 2560 -173 2660 -108
rect 3172 -173 3272 -108
rect 3376 -173 3476 -108
rect 3988 -173 4088 -108
rect 4192 -173 4292 -108
rect 4804 -173 4904 -108
rect 5008 -173 5108 -108
rect 5620 -173 5720 -108
rect 5824 -173 5924 -108
rect 6436 -173 6536 -108
rect 318 -379 416 -326
rect 318 -381 341 -379
rect 316 -430 341 -381
rect 392 -430 416 -379
rect 316 -447 416 -430
rect 520 -378 620 -365
rect 520 -430 545 -378
rect 596 -430 620 -378
rect 520 -447 620 -430
rect 1132 -378 1232 -365
rect 1132 -430 1157 -378
rect 1208 -430 1232 -378
rect 1132 -447 1232 -430
rect 1336 -378 1436 -365
rect 1336 -430 1361 -378
rect 1412 -430 1436 -378
rect 1336 -447 1436 -430
rect 1948 -378 2048 -365
rect 1948 -430 1973 -378
rect 2024 -430 2048 -378
rect 1948 -447 2048 -430
rect 2152 -378 2252 -365
rect 2152 -430 2177 -378
rect 2228 -430 2252 -378
rect 2152 -447 2252 -430
rect 2764 -379 2864 -365
rect 2764 -430 2789 -379
rect 2840 -430 2864 -379
rect 2764 -447 2864 -430
rect 2968 -379 3068 -365
rect 2968 -430 2993 -379
rect 3044 -430 3068 -379
rect 2968 -447 3068 -430
rect 3580 -379 3680 -365
rect 3580 -430 3605 -379
rect 3656 -430 3680 -379
rect 3580 -447 3680 -430
rect 3784 -378 3884 -364
rect 3784 -429 3809 -378
rect 3860 -429 3884 -378
rect 3784 -446 3884 -429
rect 4396 -379 4496 -365
rect 4396 -430 4421 -379
rect 4472 -430 4496 -379
rect 4396 -447 4496 -430
rect 4600 -379 4700 -365
rect 4600 -430 4625 -379
rect 4676 -430 4700 -379
rect 4600 -447 4700 -430
rect 5212 -380 5312 -366
rect 5212 -431 5237 -380
rect 5288 -431 5312 -380
rect 5212 -448 5312 -431
rect 5416 -380 5516 -366
rect 5416 -431 5441 -380
rect 5492 -431 5516 -380
rect 5416 -448 5516 -431
rect 6028 -380 6128 -366
rect 6028 -431 6053 -380
rect 6104 -431 6128 -380
rect 6028 -448 6128 -431
rect 6232 -381 6332 -367
rect 6232 -432 6257 -381
rect 6308 -432 6332 -381
rect 6232 -449 6332 -432
<< polycontact >>
rect 100 255 151 306
rect 744 290 792 343
rect 947 285 1010 346
rect 1558 285 1617 348
rect 1764 287 1826 347
rect 2372 286 2440 349
rect 2577 285 2640 349
rect 3188 286 3256 350
rect 3389 283 3461 352
rect 4004 284 4069 350
rect 4207 284 4274 349
rect 4825 286 4883 341
rect 5030 285 5088 340
rect 5643 294 5701 349
rect 5846 293 5904 347
rect 6472 291 6518 340
rect 76 -150 127 -99
rect 341 -430 392 -379
rect 545 -430 596 -378
rect 1157 -430 1208 -378
rect 1361 -430 1412 -378
rect 1973 -430 2024 -378
rect 2177 -430 2228 -378
rect 2789 -430 2840 -379
rect 2993 -430 3044 -379
rect 3605 -430 3656 -379
rect 3809 -429 3860 -378
rect 4421 -430 4472 -379
rect 4625 -430 4676 -379
rect 5237 -431 5288 -380
rect 5441 -431 5492 -380
rect 6053 -431 6104 -380
rect 6257 -432 6308 -381
<< metal1 >>
rect 0 435 6682 515
rect 114 335 195 348
rect 114 320 125 335
rect 86 306 125 320
rect 86 255 100 306
rect 179 281 195 335
rect 151 269 195 281
rect 151 255 166 269
rect 86 241 166 255
rect 224 191 301 202
rect 224 137 237 191
rect 291 137 301 191
rect 445 186 491 435
rect 732 345 811 356
rect 732 290 741 345
rect 797 290 811 345
rect 732 277 811 290
rect 934 346 1025 360
rect 934 285 947 346
rect 1010 285 1025 346
rect 934 273 1025 285
rect 634 194 711 209
rect 224 128 301 137
rect 634 140 645 194
rect 699 140 711 194
rect 634 128 711 140
rect 1041 195 1118 207
rect 1041 141 1053 195
rect 1107 141 1118 195
rect 1261 186 1307 435
rect 1546 348 1634 360
rect 1546 285 1558 348
rect 1617 285 1634 348
rect 1546 272 1634 285
rect 1752 347 1839 361
rect 1752 287 1764 347
rect 1826 287 1839 347
rect 1752 275 1839 287
rect 1450 195 1527 207
rect 1041 133 1118 141
rect 1450 141 1461 195
rect 1515 141 1527 195
rect 1450 133 1527 141
rect 1858 193 1935 205
rect 1858 139 1869 193
rect 1923 139 1935 193
rect 2077 186 2123 435
rect 2357 349 2455 364
rect 2357 286 2372 349
rect 2440 286 2455 349
rect 2357 273 2455 286
rect 2565 349 2656 366
rect 2565 285 2577 349
rect 2640 285 2656 349
rect 2565 272 2656 285
rect 2265 195 2342 206
rect 37 22 83 85
rect 238 69 289 128
rect 646 69 697 128
rect 853 22 899 72
rect 1054 69 1105 133
rect 1462 69 1513 133
rect 1858 131 1935 139
rect 2265 141 2276 195
rect 2330 141 2342 195
rect 2265 132 2342 141
rect 2671 193 2748 204
rect 2671 139 2683 193
rect 2737 139 2748 193
rect 2893 186 2939 435
rect 3174 350 3270 364
rect 3174 286 3188 350
rect 3256 286 3270 350
rect 3174 273 3270 286
rect 3377 352 3473 364
rect 3377 283 3389 352
rect 3461 283 3473 352
rect 3377 270 3473 283
rect 3082 198 3159 208
rect 1669 22 1715 72
rect 1870 69 1921 131
rect 2278 69 2329 132
rect 2671 130 2748 139
rect 3082 144 3093 198
rect 3147 144 3159 198
rect 3082 134 3159 144
rect 3488 193 3565 202
rect 3488 139 3500 193
rect 3554 139 3565 193
rect 3709 186 3755 435
rect 3991 350 4085 364
rect 3991 284 4004 350
rect 4069 284 4085 350
rect 3991 270 4085 284
rect 4192 349 4290 365
rect 4192 284 4207 349
rect 4274 284 4290 349
rect 4192 270 4290 284
rect 3896 197 3973 208
rect 2485 22 2531 72
rect 2686 69 2736 130
rect 3095 69 3144 134
rect 3488 128 3565 139
rect 3896 143 3908 197
rect 3962 143 3973 197
rect 3896 135 3973 143
rect 4305 202 4382 214
rect 4305 148 4316 202
rect 4370 148 4382 202
rect 4525 186 4571 435
rect 4814 341 4897 353
rect 4814 286 4825 341
rect 4883 286 4897 341
rect 4814 274 4897 286
rect 5017 340 5100 353
rect 5017 285 5030 340
rect 5088 285 5100 340
rect 5017 274 5100 285
rect 4712 200 4789 211
rect 4305 140 4382 148
rect 4712 146 4724 200
rect 4778 146 4789 200
rect 3301 22 3347 70
rect 3502 69 3552 128
rect 3910 69 3960 135
rect 4117 22 4163 80
rect 4318 69 4368 140
rect 4712 137 4789 146
rect 5122 183 5199 193
rect 5341 186 5387 435
rect 5628 349 5715 360
rect 5628 294 5643 349
rect 5701 294 5715 349
rect 5628 282 5715 294
rect 5831 347 5918 361
rect 5831 293 5846 347
rect 5904 293 5918 347
rect 5831 284 5918 293
rect 5529 216 5606 227
rect 4726 69 4776 137
rect 5122 129 5131 183
rect 5185 129 5199 183
rect 5529 162 5540 216
rect 5594 162 5606 216
rect 5529 153 5606 162
rect 5936 214 6013 227
rect 5936 160 5948 214
rect 6002 160 6013 214
rect 6157 186 6203 435
rect 6456 344 6537 356
rect 6456 288 6468 344
rect 6524 288 6537 344
rect 6456 280 6537 288
rect 6346 219 6423 231
rect 5122 119 5199 129
rect 4933 22 4979 81
rect 5134 69 5184 119
rect 5542 69 5592 153
rect 5936 150 6013 160
rect 6346 165 6356 219
rect 6410 165 6423 219
rect 6346 157 6423 165
rect 6355 156 6411 157
rect 5749 22 5795 80
rect 5950 69 6000 150
rect 6358 69 6408 156
rect 6565 22 6611 70
rect 37 -24 6611 22
rect 62 -99 140 -85
rect 62 -150 76 -99
rect 127 -150 140 -99
rect 62 -164 140 -150
rect 226 -124 307 -111
rect 226 -178 237 -124
rect 291 -178 307 -124
rect 226 -190 307 -178
rect 37 -519 83 -335
rect 238 -336 289 -190
rect 445 -219 491 -24
rect 631 -123 710 -110
rect 631 -179 644 -123
rect 700 -179 710 -123
rect 631 -189 710 -179
rect 1035 -123 1114 -110
rect 1035 -179 1047 -123
rect 1103 -179 1114 -123
rect 1035 -189 1114 -179
rect 646 -336 697 -189
rect 326 -367 404 -365
rect 530 -366 608 -365
rect 326 -379 405 -367
rect 326 -380 341 -379
rect 326 -434 337 -380
rect 392 -430 405 -379
rect 391 -434 405 -430
rect 326 -446 405 -434
rect 530 -378 609 -366
rect 530 -379 545 -378
rect 530 -433 541 -379
rect 596 -430 609 -378
rect 595 -433 609 -430
rect 530 -445 609 -433
rect 853 -519 899 -335
rect 1054 -336 1105 -189
rect 1261 -219 1307 -24
rect 1451 -123 1530 -111
rect 1451 -179 1463 -123
rect 1519 -179 1530 -123
rect 1451 -190 1530 -179
rect 1854 -123 1933 -111
rect 1854 -179 1866 -123
rect 1922 -179 1933 -123
rect 1854 -190 1933 -179
rect 1462 -336 1513 -190
rect 1142 -366 1220 -365
rect 1346 -366 1424 -365
rect 1142 -378 1221 -366
rect 1142 -379 1157 -378
rect 1142 -433 1153 -379
rect 1208 -430 1221 -378
rect 1207 -433 1221 -430
rect 1142 -445 1221 -433
rect 1346 -378 1425 -366
rect 1346 -379 1361 -378
rect 1346 -433 1357 -379
rect 1412 -430 1425 -378
rect 1411 -433 1425 -430
rect 1346 -445 1425 -433
rect 1669 -519 1715 -335
rect 1870 -336 1921 -190
rect 2077 -219 2123 -24
rect 2265 -123 2344 -110
rect 2265 -179 2276 -123
rect 2332 -179 2344 -123
rect 2265 -189 2344 -179
rect 2672 -123 2751 -111
rect 2672 -179 2684 -123
rect 2740 -179 2751 -123
rect 2278 -336 2329 -189
rect 2672 -190 2751 -179
rect 1958 -366 2036 -365
rect 2162 -366 2240 -365
rect 1958 -378 2037 -366
rect 1958 -379 1973 -378
rect 1958 -433 1969 -379
rect 2024 -430 2037 -378
rect 2023 -433 2037 -430
rect 1958 -445 2037 -433
rect 2162 -378 2241 -366
rect 2162 -379 2177 -378
rect 2162 -433 2173 -379
rect 2228 -430 2241 -378
rect 2227 -433 2241 -430
rect 2162 -445 2241 -433
rect 2485 -519 2531 -335
rect 2686 -336 2737 -190
rect 2893 -219 2939 -24
rect 3078 -123 3157 -111
rect 3078 -179 3089 -123
rect 3145 -179 3157 -123
rect 3078 -190 3157 -179
rect 3490 -123 3569 -111
rect 3490 -179 3501 -123
rect 3557 -179 3569 -123
rect 3490 -190 3569 -179
rect 3094 -336 3145 -190
rect 2774 -367 2852 -365
rect 2978 -367 3056 -365
rect 2774 -379 2853 -367
rect 2774 -435 2786 -379
rect 2842 -435 2853 -379
rect 2774 -446 2853 -435
rect 2978 -379 3057 -367
rect 2978 -435 2990 -379
rect 3046 -435 3057 -379
rect 2978 -446 3057 -435
rect 3301 -519 3347 -335
rect 3502 -336 3552 -190
rect 3709 -223 3755 -24
rect 3897 -123 3976 -111
rect 3897 -179 3908 -123
rect 3964 -179 3976 -123
rect 3897 -190 3976 -179
rect 4302 -123 4381 -110
rect 4302 -179 4314 -123
rect 4370 -179 4381 -123
rect 4302 -189 4381 -179
rect 3910 -336 3960 -190
rect 3590 -367 3668 -365
rect 3794 -366 3872 -364
rect 3590 -379 3669 -367
rect 3590 -435 3602 -379
rect 3658 -435 3669 -379
rect 3590 -446 3669 -435
rect 3794 -378 3873 -366
rect 3794 -434 3806 -378
rect 3862 -434 3873 -378
rect 3794 -445 3873 -434
rect 4117 -519 4163 -301
rect 4318 -336 4368 -189
rect 4525 -223 4571 -24
rect 4712 -123 4791 -111
rect 4712 -179 4723 -123
rect 4779 -179 4791 -123
rect 4712 -190 4791 -179
rect 5118 -123 5202 -109
rect 5118 -179 5133 -123
rect 5189 -179 5202 -123
rect 5118 -189 5202 -179
rect 4726 -336 4776 -190
rect 4406 -367 4484 -365
rect 4406 -379 4485 -367
rect 4610 -368 4688 -365
rect 4406 -435 4418 -379
rect 4474 -435 4485 -379
rect 4406 -446 4485 -435
rect 4609 -379 4688 -368
rect 4609 -380 4625 -379
rect 4676 -380 4688 -379
rect 4609 -436 4621 -380
rect 4677 -436 4688 -380
rect 4609 -447 4688 -436
rect 4933 -519 4979 -301
rect 5134 -336 5184 -189
rect 5341 -223 5387 -24
rect 5530 -113 5607 -112
rect 5525 -123 5607 -113
rect 5525 -179 5538 -123
rect 5594 -179 5607 -123
rect 5525 -186 5607 -179
rect 5933 -123 6014 -113
rect 5933 -179 5945 -123
rect 6001 -179 6014 -123
rect 5525 -187 5602 -186
rect 5933 -187 6014 -179
rect 5542 -336 5592 -187
rect 5222 -368 5300 -366
rect 5222 -380 5306 -368
rect 5426 -373 5504 -366
rect 5426 -374 5507 -373
rect 5222 -438 5237 -380
rect 5288 -382 5306 -380
rect 5293 -438 5306 -382
rect 5222 -448 5306 -438
rect 5425 -380 5507 -374
rect 5425 -384 5441 -380
rect 5492 -384 5507 -380
rect 5425 -440 5438 -384
rect 5494 -440 5507 -384
rect 5425 -447 5507 -440
rect 5425 -448 5502 -447
rect 5749 -519 5795 -308
rect 5950 -336 6000 -187
rect 6157 -225 6203 -24
rect 6349 -123 6426 -114
rect 6349 -179 6359 -123
rect 6415 -179 6426 -123
rect 6349 -188 6426 -179
rect 6358 -336 6408 -188
rect 6038 -374 6116 -366
rect 6242 -374 6320 -367
rect 6038 -380 6119 -374
rect 6038 -384 6053 -380
rect 6104 -384 6119 -380
rect 6038 -440 6050 -384
rect 6106 -440 6119 -384
rect 6038 -448 6119 -440
rect 6242 -381 6324 -374
rect 6242 -384 6257 -381
rect 6308 -384 6324 -381
rect 6242 -440 6255 -384
rect 6311 -440 6324 -384
rect 6242 -446 6324 -440
rect 6243 -448 6324 -446
rect 6565 -519 6611 -318
rect 0 -587 6685 -519
rect 0 -631 6682 -587
<< via1 >>
rect 125 306 179 335
rect 125 281 151 306
rect 151 281 179 306
rect 237 137 291 191
rect 741 343 797 345
rect 741 290 744 343
rect 744 290 792 343
rect 792 290 797 343
rect 947 285 1010 346
rect 645 140 699 194
rect 1053 141 1107 195
rect 1558 285 1617 348
rect 1764 287 1826 347
rect 1461 141 1515 195
rect 1869 139 1923 193
rect 2372 286 2440 349
rect 2577 285 2640 349
rect 2276 141 2330 195
rect 2683 139 2737 193
rect 3188 286 3256 350
rect 3389 283 3461 352
rect 3093 144 3147 198
rect 3500 139 3554 193
rect 4004 284 4069 350
rect 4207 284 4274 349
rect 3908 143 3962 197
rect 4316 148 4370 202
rect 4825 286 4883 341
rect 5030 285 5088 340
rect 4724 146 4778 200
rect 5643 294 5701 349
rect 5846 293 5904 347
rect 5131 129 5185 183
rect 5540 162 5594 216
rect 5948 160 6002 214
rect 6468 340 6524 344
rect 6468 291 6472 340
rect 6472 291 6518 340
rect 6518 291 6524 340
rect 6468 288 6524 291
rect 6356 165 6410 219
rect 237 -178 291 -124
rect 644 -179 700 -123
rect 1047 -179 1103 -123
rect 337 -430 341 -380
rect 341 -430 391 -380
rect 337 -434 391 -430
rect 541 -430 545 -379
rect 545 -430 595 -379
rect 541 -433 595 -430
rect 1463 -179 1519 -123
rect 1866 -179 1922 -123
rect 1153 -430 1157 -379
rect 1157 -430 1207 -379
rect 1153 -433 1207 -430
rect 1357 -430 1361 -379
rect 1361 -430 1411 -379
rect 1357 -433 1411 -430
rect 2276 -179 2332 -123
rect 2684 -179 2740 -123
rect 1969 -430 1973 -379
rect 1973 -430 2023 -379
rect 1969 -433 2023 -430
rect 2173 -430 2177 -379
rect 2177 -430 2227 -379
rect 2173 -433 2227 -430
rect 3089 -179 3145 -123
rect 3501 -179 3557 -123
rect 2786 -430 2789 -379
rect 2789 -430 2840 -379
rect 2840 -430 2842 -379
rect 2786 -435 2842 -430
rect 2990 -430 2993 -379
rect 2993 -430 3044 -379
rect 3044 -430 3046 -379
rect 2990 -435 3046 -430
rect 3908 -179 3964 -123
rect 4314 -179 4370 -123
rect 3602 -430 3605 -379
rect 3605 -430 3656 -379
rect 3656 -430 3658 -379
rect 3602 -435 3658 -430
rect 3806 -429 3809 -378
rect 3809 -429 3860 -378
rect 3860 -429 3862 -378
rect 3806 -434 3862 -429
rect 4723 -179 4779 -123
rect 5133 -179 5189 -123
rect 4418 -430 4421 -379
rect 4421 -430 4472 -379
rect 4472 -430 4474 -379
rect 4418 -435 4474 -430
rect 4621 -430 4625 -380
rect 4625 -430 4676 -380
rect 4676 -430 4677 -380
rect 4621 -436 4677 -430
rect 5538 -179 5594 -123
rect 5945 -179 6001 -123
rect 5237 -431 5288 -382
rect 5288 -431 5293 -382
rect 5237 -438 5293 -431
rect 5438 -431 5441 -384
rect 5441 -431 5492 -384
rect 5492 -431 5494 -384
rect 5438 -440 5494 -431
rect 6359 -179 6415 -123
rect 6050 -431 6053 -384
rect 6053 -431 6104 -384
rect 6104 -431 6106 -384
rect 6050 -440 6106 -431
rect 6255 -432 6257 -384
rect 6257 -432 6308 -384
rect 6308 -432 6311 -384
rect 6255 -440 6311 -432
<< metal2 >>
rect 114 344 195 348
rect 732 345 811 356
rect 732 344 741 345
rect 114 335 741 344
rect 114 281 125 335
rect 179 290 741 335
rect 797 344 811 345
rect 934 346 1025 360
rect 934 344 947 346
rect 797 290 947 344
rect 179 288 947 290
rect 179 281 195 288
rect 114 269 195 281
rect 732 277 811 288
rect 934 285 947 288
rect 1010 344 1025 346
rect 1546 348 1634 360
rect 1546 344 1558 348
rect 1010 288 1558 344
rect 1010 285 1025 288
rect 934 273 1025 285
rect 1546 285 1558 288
rect 1617 344 1634 348
rect 1752 347 1839 361
rect 1752 344 1764 347
rect 1617 288 1764 344
rect 1617 285 1634 288
rect 1546 272 1634 285
rect 1752 287 1764 288
rect 1826 344 1839 347
rect 2357 349 2455 364
rect 2357 344 2372 349
rect 1826 288 2372 344
rect 1826 287 1839 288
rect 1752 275 1839 287
rect 2357 286 2372 288
rect 2440 344 2455 349
rect 2565 349 2656 366
rect 2565 344 2577 349
rect 2440 288 2577 344
rect 2440 286 2455 288
rect 2357 273 2455 286
rect 2565 285 2577 288
rect 2640 344 2656 349
rect 3174 350 3270 364
rect 3174 344 3188 350
rect 2640 288 3188 344
rect 2640 285 2656 288
rect 2565 272 2656 285
rect 3174 286 3188 288
rect 3256 344 3270 350
rect 3377 352 3473 364
rect 3377 344 3389 352
rect 3256 288 3389 344
rect 3256 286 3270 288
rect 3174 273 3270 286
rect 3377 283 3389 288
rect 3461 344 3473 352
rect 3991 350 4085 364
rect 3991 344 4004 350
rect 3461 288 4004 344
rect 3461 283 3473 288
rect 3377 270 3473 283
rect 3991 284 4004 288
rect 4069 344 4085 350
rect 4192 349 4290 365
rect 4192 344 4207 349
rect 4069 288 4207 344
rect 4069 284 4085 288
rect 3991 270 4085 284
rect 4192 284 4207 288
rect 4274 344 4290 349
rect 4814 344 4897 353
rect 5017 344 5100 353
rect 5628 349 5715 360
rect 5628 344 5643 349
rect 4274 341 5643 344
rect 4274 288 4825 341
rect 4274 284 4290 288
rect 4192 270 4290 284
rect 4814 286 4825 288
rect 4883 340 5643 341
rect 4883 288 5030 340
rect 4883 286 4897 288
rect 4814 274 4897 286
rect 5017 285 5030 288
rect 5088 294 5643 340
rect 5701 344 5715 349
rect 5831 347 5918 361
rect 5831 344 5846 347
rect 5701 294 5846 344
rect 5088 293 5846 294
rect 5904 344 5918 347
rect 6456 344 6537 356
rect 5904 293 6468 344
rect 5088 288 6468 293
rect 6524 288 6537 344
rect 5088 285 5100 288
rect 5017 274 5100 285
rect 5628 282 5715 288
rect 5831 284 5918 288
rect 6456 280 6537 288
rect 5529 216 5606 227
rect 224 191 301 202
rect 224 137 237 191
rect 291 137 301 191
rect 224 128 301 137
rect 634 194 711 209
rect 634 140 645 194
rect 699 140 711 194
rect 634 128 711 140
rect 1041 195 1118 207
rect 1041 141 1053 195
rect 1107 141 1118 195
rect 1041 133 1118 141
rect 1450 195 1527 207
rect 1450 141 1461 195
rect 1515 141 1527 195
rect 1450 133 1527 141
rect 1858 193 1935 205
rect 1858 139 1869 193
rect 1923 139 1935 193
rect 236 -111 292 128
rect 644 -110 700 128
rect 1052 -110 1108 133
rect 226 -123 307 -111
rect 631 -123 710 -110
rect 1035 -123 1114 -110
rect 1460 -111 1516 133
rect 1858 131 1935 139
rect 2265 195 2342 206
rect 2265 141 2276 195
rect 2330 141 2342 195
rect 2265 132 2342 141
rect 2671 193 2748 204
rect 2671 139 2683 193
rect 2737 139 2748 193
rect 1868 -111 1924 131
rect 2276 -110 2332 132
rect 2671 130 2748 139
rect 3082 198 3159 208
rect 3082 144 3093 198
rect 3147 144 3159 198
rect 3082 134 3159 144
rect 3488 193 3565 202
rect 3488 139 3500 193
rect 3554 139 3565 193
rect 1451 -123 1530 -111
rect 1854 -123 1933 -111
rect 2265 -123 2344 -110
rect 2683 -111 2739 130
rect 3092 -111 3148 134
rect 3488 128 3565 139
rect 3896 197 3973 208
rect 3896 143 3908 197
rect 3962 143 3973 197
rect 3896 135 3973 143
rect 4305 202 4382 214
rect 4305 148 4316 202
rect 4370 148 4382 202
rect 4305 140 4382 148
rect 4712 200 4789 211
rect 4712 146 4724 200
rect 4778 146 4789 200
rect 3499 -111 3555 128
rect 3907 -111 3963 135
rect 4315 -110 4371 140
rect 4712 137 4789 146
rect 5122 183 5199 193
rect 2672 -123 2751 -111
rect 3078 -123 3157 -111
rect 3490 -123 3569 -111
rect 3897 -123 3976 -111
rect 4302 -123 4381 -110
rect 4723 -111 4779 137
rect 5122 129 5131 183
rect 5185 129 5199 183
rect 5529 162 5540 216
rect 5594 162 5606 216
rect 5529 153 5606 162
rect 5936 214 6013 227
rect 5936 160 5948 214
rect 6002 160 6013 214
rect 5122 119 5199 129
rect 5131 -109 5187 119
rect 4712 -123 4791 -111
rect 5118 -123 5202 -109
rect 5539 -112 5595 153
rect 5936 150 6013 160
rect 6346 219 6423 231
rect 6346 165 6356 219
rect 6410 165 6423 219
rect 6346 157 6423 165
rect 5530 -113 5607 -112
rect 5947 -113 6003 150
rect 5525 -123 5607 -113
rect 5933 -123 6014 -113
rect 6355 -114 6411 157
rect 6349 -123 6426 -114
rect 226 -124 644 -123
rect 226 -178 237 -124
rect 291 -178 644 -124
rect 226 -179 644 -178
rect 700 -179 1047 -123
rect 1103 -179 1463 -123
rect 1519 -179 1866 -123
rect 1922 -179 2276 -123
rect 2332 -179 2684 -123
rect 2740 -179 3089 -123
rect 3145 -179 3501 -123
rect 3557 -179 3908 -123
rect 3964 -179 4314 -123
rect 4370 -179 4723 -123
rect 4779 -179 5133 -123
rect 5189 -179 5538 -123
rect 5594 -179 5945 -123
rect 6001 -179 6359 -123
rect 6415 -179 6426 -123
rect 226 -190 307 -179
rect 631 -189 710 -179
rect 1035 -189 1114 -179
rect 1451 -190 1530 -179
rect 1854 -190 1933 -179
rect 2265 -189 2344 -179
rect 2672 -190 2751 -179
rect 3078 -190 3157 -179
rect 3490 -190 3569 -179
rect 3897 -190 3976 -179
rect 4302 -189 4381 -179
rect 4712 -190 4791 -179
rect 5118 -189 5202 -179
rect 5525 -186 5607 -179
rect 5525 -187 5602 -186
rect 5933 -187 6014 -179
rect 6349 -188 6426 -179
rect 326 -380 405 -367
rect 326 -434 337 -380
rect 391 -385 405 -380
rect 530 -379 609 -366
rect 530 -385 541 -379
rect 391 -433 541 -385
rect 595 -385 609 -379
rect 1142 -379 1221 -366
rect 1142 -385 1153 -379
rect 595 -433 1153 -385
rect 1207 -385 1221 -379
rect 1346 -379 1425 -366
rect 1346 -385 1357 -379
rect 1207 -433 1357 -385
rect 1411 -385 1425 -379
rect 1958 -379 2037 -366
rect 1958 -385 1969 -379
rect 1411 -433 1969 -385
rect 2023 -385 2037 -379
rect 2162 -379 2241 -366
rect 2162 -385 2173 -379
rect 2023 -433 2173 -385
rect 2227 -385 2241 -379
rect 2774 -379 2853 -367
rect 2774 -385 2786 -379
rect 2227 -433 2786 -385
rect 391 -434 2786 -433
rect 326 -435 2786 -434
rect 2842 -385 2853 -379
rect 2978 -379 3057 -367
rect 2978 -385 2990 -379
rect 2842 -435 2990 -385
rect 3046 -385 3057 -379
rect 3590 -379 3669 -367
rect 3590 -385 3602 -379
rect 3046 -435 3602 -385
rect 3658 -385 3669 -379
rect 3794 -378 3873 -366
rect 3794 -385 3806 -378
rect 3658 -434 3806 -385
rect 3862 -385 3873 -378
rect 4406 -379 4485 -367
rect 4406 -385 4418 -379
rect 3862 -434 4418 -385
rect 3658 -435 4418 -434
rect 4474 -385 4485 -379
rect 4609 -380 4688 -368
rect 4609 -385 4621 -380
rect 4474 -435 4621 -385
rect 326 -436 4621 -435
rect 4677 -385 4688 -380
rect 5222 -382 5306 -368
rect 5430 -374 5507 -373
rect 5222 -385 5237 -382
rect 4677 -436 5237 -385
rect 326 -438 5237 -436
rect 5293 -385 5306 -382
rect 5425 -384 5507 -374
rect 5425 -385 5438 -384
rect 5293 -438 5438 -385
rect 326 -440 5438 -438
rect 5494 -385 5507 -384
rect 6038 -384 6119 -374
rect 6038 -385 6050 -384
rect 5494 -440 6050 -385
rect 6106 -385 6119 -384
rect 6243 -384 6324 -374
rect 6243 -385 6255 -384
rect 6106 -440 6255 -385
rect 6311 -440 6324 -384
rect 326 -441 6324 -440
rect 326 -446 405 -441
rect 530 -445 609 -441
rect 1142 -445 1221 -441
rect 1346 -445 1425 -441
rect 1958 -445 2037 -441
rect 2162 -445 2241 -441
rect 2774 -446 2853 -441
rect 2978 -446 3057 -441
rect 3590 -446 3669 -441
rect 3794 -445 3873 -441
rect 4406 -446 4485 -441
rect 4609 -447 4688 -441
rect 5222 -448 5306 -441
rect 5425 -447 5507 -441
rect 5425 -448 5502 -447
rect 6038 -448 6119 -441
rect 6243 -448 6324 -441
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_0
timestamp 1691401996
transform 1 0 2406 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_1
timestamp 1691401996
transform 1 0 162 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_2
timestamp 1691401996
transform 1 0 366 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_3
timestamp 1691401996
transform 1 0 570 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_4
timestamp 1691401996
transform 1 0 774 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_5
timestamp 1691401996
transform 1 0 978 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_6
timestamp 1691401996
transform 1 0 1182 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_7
timestamp 1691401996
transform 1 0 1386 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_8
timestamp 1691401996
transform 1 0 1590 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_9
timestamp 1691401996
transform 1 0 1794 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_10
timestamp 1691401996
transform 1 0 1998 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_11
timestamp 1691401996
transform 1 0 2202 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_12
timestamp 1691401996
transform 1 0 2814 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_13
timestamp 1691401996
transform 1 0 2610 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_14
timestamp 1691401996
transform 1 0 3018 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_15
timestamp 1691401996
transform 1 0 3222 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_16
timestamp 1691401996
transform 1 0 3630 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_17
timestamp 1691401996
transform 1 0 3426 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_18
timestamp 1691401996
transform 1 0 3834 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_19
timestamp 1691401996
transform 1 0 4242 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_20
timestamp 1691401996
transform 1 0 4038 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_21
timestamp 1691401996
transform 1 0 4446 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_22
timestamp 1691401996
transform 1 0 4854 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_23
timestamp 1691401996
transform 1 0 4650 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_24
timestamp 1691401996
transform 1 0 5058 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_25
timestamp 1691401996
transform 1 0 5466 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_26
timestamp 1691401996
transform 1 0 5262 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_27
timestamp 1691401996
transform 1 0 6078 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_28
timestamp 1691401996
transform 1 0 5670 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_29
timestamp 1691401996
transform 1 0 5874 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_30
timestamp 1691401996
transform 1 0 6486 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_31
timestamp 1691401996
transform 1 0 6282 0 1 -277
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_0
timestamp 1691392065
transform 1 0 1998 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_1
timestamp 1691392065
transform 1 0 162 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_2
timestamp 1691392065
transform 1 0 366 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_3
timestamp 1691392065
transform 1 0 570 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_4
timestamp 1691392065
transform 1 0 774 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_5
timestamp 1691392065
transform 1 0 978 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_6
timestamp 1691392065
transform 1 0 1182 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_7
timestamp 1691392065
transform 1 0 1386 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_8
timestamp 1691392065
transform 1 0 1590 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_9
timestamp 1691392065
transform 1 0 1794 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_10
timestamp 1691392065
transform 1 0 3222 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_11
timestamp 1691392065
transform 1 0 2202 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_12
timestamp 1691392065
transform 1 0 2406 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_13
timestamp 1691392065
transform 1 0 2610 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_14
timestamp 1691392065
transform 1 0 2814 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_15
timestamp 1691392065
transform 1 0 3018 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_16
timestamp 1691392065
transform 1 0 5466 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_17
timestamp 1691392065
transform 1 0 3426 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_18
timestamp 1691392065
transform 1 0 3630 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_19
timestamp 1691392065
transform 1 0 3834 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_20
timestamp 1691392065
transform 1 0 4038 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_21
timestamp 1691392065
transform 1 0 4242 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_22
timestamp 1691392065
transform 1 0 4446 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_23
timestamp 1691392065
transform 1 0 4650 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_24
timestamp 1691392065
transform 1 0 4854 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_25
timestamp 1691392065
transform 1 0 5058 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_26
timestamp 1691392065
transform 1 0 5262 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_27
timestamp 1691392065
transform 1 0 6078 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_28
timestamp 1691392065
transform 1 0 5670 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_29
timestamp 1691392065
transform 1 0 5874 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_30
timestamp 1691392065
transform 1 0 6486 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_31
timestamp 1691392065
transform 1 0 6282 0 1 128
box -162 -128 162 128
<< end >>
