magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2230 -2614 2230 2614
<< nwell >>
rect -230 -614 230 614
<< pmos >>
rect -56 344 56 484
rect -56 68 56 208
rect -56 -208 56 -68
rect -56 -484 56 -344
<< pdiff >>
rect -144 437 -56 484
rect -144 391 -131 437
rect -85 391 -56 437
rect -144 344 -56 391
rect 56 437 144 484
rect 56 391 85 437
rect 131 391 144 437
rect 56 344 144 391
rect -144 161 -56 208
rect -144 115 -131 161
rect -85 115 -56 161
rect -144 68 -56 115
rect 56 161 144 208
rect 56 115 85 161
rect 131 115 144 161
rect 56 68 144 115
rect -144 -115 -56 -68
rect -144 -161 -131 -115
rect -85 -161 -56 -115
rect -144 -208 -56 -161
rect 56 -115 144 -68
rect 56 -161 85 -115
rect 131 -161 144 -115
rect 56 -208 144 -161
rect -144 -391 -56 -344
rect -144 -437 -131 -391
rect -85 -437 -56 -391
rect -144 -484 -56 -437
rect 56 -391 144 -344
rect 56 -437 85 -391
rect 131 -437 144 -391
rect 56 -484 144 -437
<< pdiffc >>
rect -131 391 -85 437
rect 85 391 131 437
rect -131 115 -85 161
rect 85 115 131 161
rect -131 -161 -85 -115
rect 85 -161 131 -115
rect -131 -437 -85 -391
rect 85 -437 131 -391
<< polysilicon >>
rect -56 484 56 528
rect -56 300 56 344
rect -56 208 56 252
rect -56 24 56 68
rect -56 -68 56 -24
rect -56 -252 56 -208
rect -56 -344 56 -300
rect -56 -528 56 -484
<< metal1 >>
rect -131 437 -85 482
rect -131 346 -85 391
rect 85 437 131 482
rect 85 346 131 391
rect -131 161 -85 206
rect -131 70 -85 115
rect 85 161 131 206
rect 85 70 131 115
rect -131 -115 -85 -70
rect -131 -206 -85 -161
rect 85 -115 131 -70
rect 85 -206 131 -161
rect -131 -391 -85 -346
rect -131 -482 -85 -437
rect 85 -391 131 -346
rect 85 -482 131 -437
<< end >>
