** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/7b_divider_tb.sch
**.subckt 7b_divider_tb
V1 VSS GND 0
V2 VDD VSS 3.3
V3 CLK VSS pulse(0 3.3 0 10p 10p 5n 10n)
V5 D2_1 VSS 0
V9 D2_4 VSS 3.3
V7 D2_7 VSS 0
V10 D2_6 VSS 0
V8 D2_5 VSS 0
V4 D2_3 VSS 0
V6 D2_2 VSS 0
x1 VDD LD D2_7 Q1 D2_6 Q2 D2_5 D2_4 Q3 Q4 D2_3 D2_2 Q5 D2_1 Q6 Q7 CLK VSS OUT1 P2 pex_7b_divider_magic
**** begin user architecture code


*.option savecurrents
.include pex_7b_divider_magic.spice
.control
save all

tran 100n 5u
set xbrushwidth=2
set xfontsize=3
plot v(CLK) v(Q3)+3.5 v(Q2)+7 v(Q1)+10.5 v(P2)+14 v(x1.P0)+17.5 v(OUT1)+21 v(LD)+24.5 v(Q4)+28 v(Q5)+31.5
plot v(Q1)
plot v(Q2)
plot v(Q3) v(Q2) v(Q1)
write 7b_divider_tb.raw
*write test_nfet_03v3.raw
.endc



.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical

**** end user architecture code
**.ends
.GLOBAL GND
.end
