magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1205 -1329 1205 1329
<< metal1 >>
rect -205 323 205 329
rect -205 297 -199 323
rect -173 297 -137 323
rect -111 297 -75 323
rect -49 297 -13 323
rect 13 297 49 323
rect 75 297 111 323
rect 137 297 173 323
rect 199 297 205 323
rect -205 261 205 297
rect -205 235 -199 261
rect -173 235 -137 261
rect -111 235 -75 261
rect -49 235 -13 261
rect 13 235 49 261
rect 75 235 111 261
rect 137 235 173 261
rect 199 235 205 261
rect -205 199 205 235
rect -205 173 -199 199
rect -173 173 -137 199
rect -111 173 -75 199
rect -49 173 -13 199
rect 13 173 49 199
rect 75 173 111 199
rect 137 173 173 199
rect 199 173 205 199
rect -205 137 205 173
rect -205 111 -199 137
rect -173 111 -137 137
rect -111 111 -75 137
rect -49 111 -13 137
rect 13 111 49 137
rect 75 111 111 137
rect 137 111 173 137
rect 199 111 205 137
rect -205 75 205 111
rect -205 49 -199 75
rect -173 49 -137 75
rect -111 49 -75 75
rect -49 49 -13 75
rect 13 49 49 75
rect 75 49 111 75
rect 137 49 173 75
rect 199 49 205 75
rect -205 13 205 49
rect -205 -13 -199 13
rect -173 -13 -137 13
rect -111 -13 -75 13
rect -49 -13 -13 13
rect 13 -13 49 13
rect 75 -13 111 13
rect 137 -13 173 13
rect 199 -13 205 13
rect -205 -49 205 -13
rect -205 -75 -199 -49
rect -173 -75 -137 -49
rect -111 -75 -75 -49
rect -49 -75 -13 -49
rect 13 -75 49 -49
rect 75 -75 111 -49
rect 137 -75 173 -49
rect 199 -75 205 -49
rect -205 -111 205 -75
rect -205 -137 -199 -111
rect -173 -137 -137 -111
rect -111 -137 -75 -111
rect -49 -137 -13 -111
rect 13 -137 49 -111
rect 75 -137 111 -111
rect 137 -137 173 -111
rect 199 -137 205 -111
rect -205 -173 205 -137
rect -205 -199 -199 -173
rect -173 -199 -137 -173
rect -111 -199 -75 -173
rect -49 -199 -13 -173
rect 13 -199 49 -173
rect 75 -199 111 -173
rect 137 -199 173 -173
rect 199 -199 205 -173
rect -205 -235 205 -199
rect -205 -261 -199 -235
rect -173 -261 -137 -235
rect -111 -261 -75 -235
rect -49 -261 -13 -235
rect 13 -261 49 -235
rect 75 -261 111 -235
rect 137 -261 173 -235
rect 199 -261 205 -235
rect -205 -297 205 -261
rect -205 -323 -199 -297
rect -173 -323 -137 -297
rect -111 -323 -75 -297
rect -49 -323 -13 -297
rect 13 -323 49 -297
rect 75 -323 111 -297
rect 137 -323 173 -297
rect 199 -323 205 -297
rect -205 -329 205 -323
<< via1 >>
rect -199 297 -173 323
rect -137 297 -111 323
rect -75 297 -49 323
rect -13 297 13 323
rect 49 297 75 323
rect 111 297 137 323
rect 173 297 199 323
rect -199 235 -173 261
rect -137 235 -111 261
rect -75 235 -49 261
rect -13 235 13 261
rect 49 235 75 261
rect 111 235 137 261
rect 173 235 199 261
rect -199 173 -173 199
rect -137 173 -111 199
rect -75 173 -49 199
rect -13 173 13 199
rect 49 173 75 199
rect 111 173 137 199
rect 173 173 199 199
rect -199 111 -173 137
rect -137 111 -111 137
rect -75 111 -49 137
rect -13 111 13 137
rect 49 111 75 137
rect 111 111 137 137
rect 173 111 199 137
rect -199 49 -173 75
rect -137 49 -111 75
rect -75 49 -49 75
rect -13 49 13 75
rect 49 49 75 75
rect 111 49 137 75
rect 173 49 199 75
rect -199 -13 -173 13
rect -137 -13 -111 13
rect -75 -13 -49 13
rect -13 -13 13 13
rect 49 -13 75 13
rect 111 -13 137 13
rect 173 -13 199 13
rect -199 -75 -173 -49
rect -137 -75 -111 -49
rect -75 -75 -49 -49
rect -13 -75 13 -49
rect 49 -75 75 -49
rect 111 -75 137 -49
rect 173 -75 199 -49
rect -199 -137 -173 -111
rect -137 -137 -111 -111
rect -75 -137 -49 -111
rect -13 -137 13 -111
rect 49 -137 75 -111
rect 111 -137 137 -111
rect 173 -137 199 -111
rect -199 -199 -173 -173
rect -137 -199 -111 -173
rect -75 -199 -49 -173
rect -13 -199 13 -173
rect 49 -199 75 -173
rect 111 -199 137 -173
rect 173 -199 199 -173
rect -199 -261 -173 -235
rect -137 -261 -111 -235
rect -75 -261 -49 -235
rect -13 -261 13 -235
rect 49 -261 75 -235
rect 111 -261 137 -235
rect 173 -261 199 -235
rect -199 -323 -173 -297
rect -137 -323 -111 -297
rect -75 -323 -49 -297
rect -13 -323 13 -297
rect 49 -323 75 -297
rect 111 -323 137 -297
rect 173 -323 199 -297
<< metal2 >>
rect -205 323 205 329
rect -205 297 -199 323
rect -173 297 -137 323
rect -111 297 -75 323
rect -49 297 -13 323
rect 13 297 49 323
rect 75 297 111 323
rect 137 297 173 323
rect 199 297 205 323
rect -205 261 205 297
rect -205 235 -199 261
rect -173 235 -137 261
rect -111 235 -75 261
rect -49 235 -13 261
rect 13 235 49 261
rect 75 235 111 261
rect 137 235 173 261
rect 199 235 205 261
rect -205 199 205 235
rect -205 173 -199 199
rect -173 173 -137 199
rect -111 173 -75 199
rect -49 173 -13 199
rect 13 173 49 199
rect 75 173 111 199
rect 137 173 173 199
rect 199 173 205 199
rect -205 137 205 173
rect -205 111 -199 137
rect -173 111 -137 137
rect -111 111 -75 137
rect -49 111 -13 137
rect 13 111 49 137
rect 75 111 111 137
rect 137 111 173 137
rect 199 111 205 137
rect -205 75 205 111
rect -205 49 -199 75
rect -173 49 -137 75
rect -111 49 -75 75
rect -49 49 -13 75
rect 13 49 49 75
rect 75 49 111 75
rect 137 49 173 75
rect 199 49 205 75
rect -205 13 205 49
rect -205 -13 -199 13
rect -173 -13 -137 13
rect -111 -13 -75 13
rect -49 -13 -13 13
rect 13 -13 49 13
rect 75 -13 111 13
rect 137 -13 173 13
rect 199 -13 205 13
rect -205 -49 205 -13
rect -205 -75 -199 -49
rect -173 -75 -137 -49
rect -111 -75 -75 -49
rect -49 -75 -13 -49
rect 13 -75 49 -49
rect 75 -75 111 -49
rect 137 -75 173 -49
rect 199 -75 205 -49
rect -205 -111 205 -75
rect -205 -137 -199 -111
rect -173 -137 -137 -111
rect -111 -137 -75 -111
rect -49 -137 -13 -111
rect 13 -137 49 -111
rect 75 -137 111 -111
rect 137 -137 173 -111
rect 199 -137 205 -111
rect -205 -173 205 -137
rect -205 -199 -199 -173
rect -173 -199 -137 -173
rect -111 -199 -75 -173
rect -49 -199 -13 -173
rect 13 -199 49 -173
rect 75 -199 111 -173
rect 137 -199 173 -173
rect 199 -199 205 -173
rect -205 -235 205 -199
rect -205 -261 -199 -235
rect -173 -261 -137 -235
rect -111 -261 -75 -235
rect -49 -261 -13 -235
rect 13 -261 49 -235
rect 75 -261 111 -235
rect 137 -261 173 -235
rect 199 -261 205 -235
rect -205 -297 205 -261
rect -205 -323 -199 -297
rect -173 -323 -137 -297
rect -111 -323 -75 -297
rect -49 -323 -13 -297
rect 13 -323 49 -297
rect 75 -323 111 -297
rect 137 -323 173 -297
rect 199 -323 205 -297
rect -205 -329 205 -323
<< end >>
