magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1357 1019 1357
<< metal1 >>
rect -19 351 19 357
rect -19 -351 -13 351
rect 13 -351 19 351
rect -19 -357 19 -351
<< via1 >>
rect -13 -351 13 351
<< metal2 >>
rect -19 351 19 357
rect -19 -351 -13 351
rect 13 -351 19 351
rect -19 -357 19 -351
<< end >>
