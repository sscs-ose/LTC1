magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1123 1019 1123
<< metal1 >>
rect -19 117 19 123
rect -19 -117 -13 117
rect 13 -117 19 117
rect -19 -123 19 -117
<< via1 >>
rect -13 -117 13 117
<< metal2 >>
rect -19 117 19 123
rect -19 -117 -13 117
rect 13 -117 19 117
rect -19 -123 19 -117
<< end >>
