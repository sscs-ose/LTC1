magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2145 -7045 2145 7045
<< psubdiff >>
rect -145 5005 145 5045
rect -145 -5005 -117 5005
rect 117 -5005 145 5005
rect -145 -5045 145 -5005
<< psubdiffcont >>
rect -117 -5005 117 5005
<< metal1 >>
rect -134 5005 134 5034
rect -134 -5005 -117 5005
rect 117 -5005 134 5005
rect -134 -5034 134 -5005
<< end >>
