magic
tech gf180mcuC
magscale 1 10
timestamp 1692950565
<< error_s >>
rect -3306 -4270 -3182 -4246
rect -1330 -4270 -1206 -4246
rect -3282 -4294 -3206 -4270
rect -1306 -4294 -1230 -4270
rect -1726 -4406 -1664 -4404
rect -1726 -4463 -1724 -4406
rect -1666 -4463 -1664 -4406
rect -1726 -4465 -1664 -4463
rect -2593 -4684 -2537 -4682
rect -2593 -4736 -2591 -4684
rect -2539 -4736 -2537 -4684
rect -2593 -4738 -2537 -4736
rect -1952 -4684 -1896 -4682
rect -1952 -4736 -1950 -4684
rect -1898 -4736 -1896 -4684
rect -1952 -4738 -1896 -4736
rect -2753 -4841 -2697 -4839
rect -2113 -4840 -2057 -4838
rect -2753 -4893 -2751 -4841
rect -2699 -4893 -2697 -4841
rect -2753 -4895 -2697 -4893
rect -2433 -4842 -2377 -4840
rect -2433 -4894 -2431 -4842
rect -2379 -4894 -2377 -4842
rect -2113 -4892 -2111 -4840
rect -2059 -4892 -2057 -4840
rect -2113 -4894 -2057 -4892
rect -1793 -4841 -1737 -4839
rect -1793 -4893 -1791 -4841
rect -1739 -4893 -1737 -4841
rect -2433 -4896 -2377 -4894
rect -1793 -4895 -1737 -4893
rect -3074 -4991 -3018 -4989
rect -3074 -5043 -3072 -4991
rect -3020 -5043 -3018 -4991
rect -3074 -5045 -3018 -5043
rect -2913 -4991 -2857 -4989
rect -2913 -5043 -2911 -4991
rect -2859 -5043 -2857 -4991
rect -2913 -5045 -2857 -5043
rect -2274 -4991 -2216 -4989
rect -2274 -5043 -2272 -4991
rect -2218 -5043 -2216 -4991
rect -2274 -5045 -2216 -5043
rect -1633 -4991 -1577 -4989
rect -1633 -5043 -1631 -4991
rect -1579 -5043 -1577 -4991
rect -1633 -5045 -1577 -5043
rect -1473 -4991 -1417 -4989
rect -1473 -5043 -1471 -4991
rect -1419 -5043 -1417 -4991
rect -1473 -5045 -1417 -5043
rect -2830 -5268 -2774 -5266
rect -2830 -5320 -2828 -5268
rect -2776 -5320 -2774 -5268
rect -2830 -5322 -2774 -5320
rect -2593 -5544 -2537 -5542
rect -2593 -5596 -2591 -5544
rect -2539 -5596 -2537 -5544
rect -2593 -5598 -2537 -5596
rect -1952 -5544 -1896 -5542
rect -1952 -5596 -1950 -5544
rect -1898 -5596 -1896 -5544
rect -1952 -5598 -1896 -5596
rect -2755 -5696 -2699 -5694
rect -2755 -5748 -2753 -5696
rect -2701 -5748 -2699 -5696
rect -2755 -5750 -2699 -5748
rect -2433 -5695 -2377 -5693
rect -2433 -5747 -2431 -5695
rect -2379 -5747 -2377 -5695
rect -2433 -5749 -2377 -5747
rect -2115 -5695 -2059 -5693
rect -2115 -5747 -2113 -5695
rect -2061 -5747 -2059 -5695
rect -2115 -5749 -2059 -5747
rect -1792 -5695 -1736 -5693
rect -1792 -5747 -1790 -5695
rect -1738 -5747 -1736 -5695
rect -1792 -5749 -1736 -5747
rect -3074 -5851 -3018 -5849
rect -3074 -5903 -3072 -5851
rect -3020 -5903 -3018 -5851
rect -3074 -5905 -3018 -5903
rect -2913 -5851 -2857 -5849
rect -2913 -5903 -2911 -5851
rect -2859 -5903 -2857 -5851
rect -2913 -5905 -2857 -5903
rect -2274 -5851 -2216 -5849
rect -2274 -5903 -2272 -5851
rect -2218 -5903 -2216 -5851
rect -2274 -5905 -2216 -5903
rect -1633 -5851 -1577 -5849
rect -1633 -5903 -1631 -5851
rect -1579 -5903 -1577 -5851
rect -1633 -5905 -1577 -5903
rect -1473 -5851 -1417 -5849
rect -1473 -5903 -1471 -5851
rect -1419 -5903 -1417 -5851
rect -1473 -5905 -1417 -5903
rect -1721 -6089 -1665 -6087
rect -1721 -6141 -1719 -6089
rect -1667 -6141 -1665 -6089
rect -1721 -6143 -1665 -6141
<< nwell >>
rect -3327 -6363 -1192 -4270
<< nsubdiff >>
rect -3282 -4286 -3206 -4270
rect -3282 -4332 -3267 -4286
rect -3221 -4332 -3206 -4286
rect -3282 -4380 -3206 -4332
rect -1306 -4286 -1230 -4270
rect -1306 -4332 -1291 -4286
rect -1245 -4332 -1230 -4286
rect -3282 -4426 -3267 -4380
rect -3221 -4426 -3206 -4380
rect -3282 -4474 -3206 -4426
rect -3282 -4520 -3267 -4474
rect -3221 -4520 -3206 -4474
rect -1306 -4380 -1230 -4332
rect -1306 -4426 -1291 -4380
rect -1245 -4426 -1230 -4380
rect -3282 -4568 -3206 -4520
rect -3282 -4614 -3267 -4568
rect -3221 -4614 -3206 -4568
rect -1306 -4474 -1230 -4426
rect -1306 -4520 -1291 -4474
rect -1245 -4520 -1230 -4474
rect -1306 -4568 -1230 -4520
rect -3282 -4662 -3206 -4614
rect -3282 -4708 -3267 -4662
rect -3221 -4708 -3206 -4662
rect -3282 -4756 -3206 -4708
rect -3282 -4802 -3267 -4756
rect -3221 -4802 -3206 -4756
rect -3282 -4850 -3206 -4802
rect -3282 -4896 -3267 -4850
rect -3221 -4896 -3206 -4850
rect -3282 -4944 -3206 -4896
rect -3282 -4990 -3267 -4944
rect -3221 -4990 -3206 -4944
rect -3282 -5038 -3206 -4990
rect -3282 -5084 -3267 -5038
rect -3221 -5084 -3206 -5038
rect -3282 -5132 -3206 -5084
rect -3282 -5178 -3267 -5132
rect -3221 -5178 -3206 -5132
rect -1306 -4614 -1291 -4568
rect -1245 -4614 -1230 -4568
rect -1306 -4662 -1230 -4614
rect -1306 -4708 -1291 -4662
rect -1245 -4708 -1230 -4662
rect -1306 -4756 -1230 -4708
rect -1306 -4802 -1291 -4756
rect -1245 -4802 -1230 -4756
rect -1306 -4850 -1230 -4802
rect -1306 -4896 -1291 -4850
rect -1245 -4896 -1230 -4850
rect -1306 -4944 -1230 -4896
rect -1306 -4990 -1291 -4944
rect -1245 -4990 -1230 -4944
rect -1306 -5038 -1230 -4990
rect -1306 -5084 -1291 -5038
rect -1245 -5084 -1230 -5038
rect -1306 -5132 -1230 -5084
rect -3282 -5226 -3206 -5178
rect -3282 -5272 -3267 -5226
rect -3221 -5272 -3206 -5226
rect -3282 -5320 -3206 -5272
rect -1306 -5178 -1291 -5132
rect -1245 -5178 -1230 -5132
rect -3282 -5366 -3267 -5320
rect -3221 -5366 -3206 -5320
rect -1306 -5226 -1230 -5178
rect -1306 -5272 -1291 -5226
rect -1245 -5272 -1230 -5226
rect -1306 -5320 -1230 -5272
rect -3282 -5414 -3206 -5366
rect -3282 -5460 -3267 -5414
rect -3221 -5460 -3206 -5414
rect -1306 -5366 -1291 -5320
rect -1245 -5366 -1230 -5320
rect -1306 -5414 -1230 -5366
rect -3282 -5508 -3206 -5460
rect -3282 -5554 -3267 -5508
rect -3221 -5554 -3206 -5508
rect -3282 -5602 -3206 -5554
rect -3282 -5648 -3267 -5602
rect -3221 -5648 -3206 -5602
rect -3282 -5696 -3206 -5648
rect -3282 -5742 -3267 -5696
rect -3221 -5742 -3206 -5696
rect -3282 -5790 -3206 -5742
rect -3282 -5836 -3267 -5790
rect -3221 -5836 -3206 -5790
rect -3282 -5884 -3206 -5836
rect -3282 -5930 -3267 -5884
rect -3221 -5930 -3206 -5884
rect -3282 -5978 -3206 -5930
rect -3282 -6024 -3267 -5978
rect -3221 -6024 -3206 -5978
rect -1306 -5460 -1291 -5414
rect -1245 -5460 -1230 -5414
rect -1306 -5508 -1230 -5460
rect -1306 -5554 -1291 -5508
rect -1245 -5554 -1230 -5508
rect -1306 -5602 -1230 -5554
rect -1306 -5648 -1291 -5602
rect -1245 -5648 -1230 -5602
rect -1306 -5696 -1230 -5648
rect -1306 -5742 -1291 -5696
rect -1245 -5742 -1230 -5696
rect -1306 -5790 -1230 -5742
rect -1306 -5836 -1291 -5790
rect -1245 -5836 -1230 -5790
rect -1306 -5884 -1230 -5836
rect -1306 -5930 -1291 -5884
rect -1245 -5930 -1230 -5884
rect -1306 -5978 -1230 -5930
rect -3282 -6072 -3206 -6024
rect -3282 -6118 -3267 -6072
rect -3221 -6118 -3206 -6072
rect -3282 -6166 -3206 -6118
rect -1306 -6024 -1291 -5978
rect -1245 -6024 -1230 -5978
rect -1306 -6072 -1230 -6024
rect -1306 -6118 -1291 -6072
rect -1245 -6118 -1230 -6072
rect -3282 -6212 -3267 -6166
rect -3221 -6212 -3206 -6166
rect -3282 -6245 -3206 -6212
rect -1306 -6166 -1230 -6118
rect -1306 -6212 -1291 -6166
rect -1245 -6212 -1230 -6166
rect -1306 -6245 -1230 -6212
rect -3282 -6260 -1230 -6245
rect -3282 -6306 -3266 -6260
rect -3220 -6306 -3172 -6260
rect -3126 -6306 -3078 -6260
rect -3032 -6306 -2984 -6260
rect -2938 -6306 -2890 -6260
rect -2844 -6306 -2796 -6260
rect -2750 -6306 -2702 -6260
rect -2656 -6306 -2608 -6260
rect -2562 -6306 -2514 -6260
rect -2468 -6306 -2420 -6260
rect -2374 -6306 -2326 -6260
rect -2280 -6306 -2232 -6260
rect -2186 -6306 -2138 -6260
rect -2092 -6306 -2044 -6260
rect -1998 -6306 -1950 -6260
rect -1904 -6306 -1856 -6260
rect -1810 -6306 -1762 -6260
rect -1716 -6306 -1668 -6260
rect -1622 -6306 -1574 -6260
rect -1528 -6306 -1480 -6260
rect -1434 -6306 -1386 -6260
rect -1340 -6306 -1292 -6260
rect -1246 -6306 -1230 -6260
rect -3282 -6321 -1230 -6306
<< nsubdiffcont >>
rect -3267 -4332 -3221 -4286
rect -1291 -4332 -1245 -4286
rect -3267 -4426 -3221 -4380
rect -3267 -4520 -3221 -4474
rect -1291 -4426 -1245 -4380
rect -3267 -4614 -3221 -4568
rect -1291 -4520 -1245 -4474
rect -3267 -4708 -3221 -4662
rect -3267 -4802 -3221 -4756
rect -3267 -4896 -3221 -4850
rect -3267 -4990 -3221 -4944
rect -3267 -5084 -3221 -5038
rect -3267 -5178 -3221 -5132
rect -1291 -4614 -1245 -4568
rect -1291 -4708 -1245 -4662
rect -1291 -4802 -1245 -4756
rect -1291 -4896 -1245 -4850
rect -1291 -4990 -1245 -4944
rect -1291 -5084 -1245 -5038
rect -3267 -5272 -3221 -5226
rect -1291 -5178 -1245 -5132
rect -3267 -5366 -3221 -5320
rect -1291 -5272 -1245 -5226
rect -3267 -5460 -3221 -5414
rect -1291 -5366 -1245 -5320
rect -3267 -5554 -3221 -5508
rect -3267 -5648 -3221 -5602
rect -3267 -5742 -3221 -5696
rect -3267 -5836 -3221 -5790
rect -3267 -5930 -3221 -5884
rect -3267 -6024 -3221 -5978
rect -1291 -5460 -1245 -5414
rect -1291 -5554 -1245 -5508
rect -1291 -5648 -1245 -5602
rect -1291 -5742 -1245 -5696
rect -1291 -5836 -1245 -5790
rect -1291 -5930 -1245 -5884
rect -3267 -6118 -3221 -6072
rect -1291 -6024 -1245 -5978
rect -1291 -6118 -1245 -6072
rect -3267 -6212 -3221 -6166
rect -1291 -6212 -1245 -6166
rect -3266 -6306 -3220 -6260
rect -3172 -6306 -3126 -6260
rect -3078 -6306 -3032 -6260
rect -2984 -6306 -2938 -6260
rect -2890 -6306 -2844 -6260
rect -2796 -6306 -2750 -6260
rect -2702 -6306 -2656 -6260
rect -2608 -6306 -2562 -6260
rect -2514 -6306 -2468 -6260
rect -2420 -6306 -2374 -6260
rect -2326 -6306 -2280 -6260
rect -2232 -6306 -2186 -6260
rect -2138 -6306 -2092 -6260
rect -2044 -6306 -1998 -6260
rect -1950 -6306 -1904 -6260
rect -1856 -6306 -1810 -6260
rect -1762 -6306 -1716 -6260
rect -1668 -6306 -1622 -6260
rect -1574 -6306 -1528 -6260
rect -1480 -6306 -1434 -6260
rect -1386 -6306 -1340 -6260
rect -1292 -6306 -1246 -6260
<< polysilicon >>
rect -3086 -4380 -2937 -4361
rect -3086 -4426 -3068 -4380
rect -3022 -4426 -2937 -4380
rect -2673 -4402 -2617 -4361
rect -3086 -4453 -2937 -4426
rect -2688 -4420 -2601 -4402
rect -2513 -4403 -2457 -4361
rect -2033 -4403 -1977 -4361
rect -1873 -4402 -1817 -4361
rect -1553 -4381 -1396 -4361
rect -2688 -4466 -2667 -4420
rect -2621 -4466 -2601 -4420
rect -2688 -4484 -2601 -4466
rect -2529 -4420 -2442 -4403
rect -2529 -4466 -2507 -4420
rect -2461 -4466 -2442 -4420
rect -2529 -4483 -2442 -4466
rect -2048 -4420 -1961 -4403
rect -2048 -4466 -2029 -4420
rect -1983 -4466 -1961 -4420
rect -2048 -4483 -1961 -4466
rect -1889 -4420 -1802 -4402
rect -1889 -4466 -1869 -4420
rect -1823 -4466 -1802 -4420
rect -1553 -4427 -1468 -4381
rect -1422 -4427 -1396 -4381
rect -1553 -4448 -1396 -4427
rect -2993 -4569 -2937 -4525
rect -2833 -4569 -2777 -4525
rect -2673 -4569 -2617 -4484
rect -2513 -4569 -2457 -4483
rect -2353 -4569 -2297 -4525
rect -2193 -4569 -2137 -4525
rect -2033 -4569 -1977 -4483
rect -1889 -4484 -1802 -4466
rect -1873 -4569 -1817 -4484
rect -1713 -4569 -1657 -4525
rect -1553 -4569 -1497 -4525
rect -2993 -5213 -2937 -5169
rect -3083 -5231 -2937 -5213
rect -3083 -5277 -3068 -5231
rect -3022 -5277 -2937 -5231
rect -2833 -5246 -2777 -5169
rect -2673 -5213 -2617 -5169
rect -2513 -5213 -2457 -5169
rect -2353 -5246 -2297 -5169
rect -2193 -5246 -2137 -5169
rect -2033 -5213 -1977 -5169
rect -1873 -5213 -1817 -5169
rect -1713 -5246 -1657 -5169
rect -1553 -5213 -1497 -5169
rect -1553 -5232 -1403 -5213
rect -3083 -5296 -2937 -5277
rect -2845 -5260 -2767 -5246
rect -2845 -5306 -2829 -5260
rect -2783 -5306 -2767 -5260
rect -2363 -5263 -2285 -5246
rect -2845 -5323 -2767 -5306
rect -2684 -5281 -2606 -5267
rect -2684 -5327 -2668 -5281
rect -2622 -5327 -2606 -5281
rect -2684 -5344 -2606 -5327
rect -2524 -5282 -2446 -5267
rect -2524 -5328 -2508 -5282
rect -2462 -5328 -2446 -5282
rect -2363 -5309 -2348 -5263
rect -2302 -5309 -2285 -5263
rect -2363 -5323 -2285 -5309
rect -2205 -5263 -2127 -5246
rect -2205 -5309 -2188 -5263
rect -2142 -5309 -2127 -5263
rect -1723 -5260 -1645 -5246
rect -2205 -5323 -2127 -5309
rect -2044 -5282 -1966 -5267
rect -2524 -5344 -2446 -5328
rect -2044 -5328 -2028 -5282
rect -1982 -5328 -1966 -5282
rect -2044 -5344 -1966 -5328
rect -1884 -5281 -1806 -5267
rect -1884 -5327 -1868 -5281
rect -1822 -5327 -1806 -5281
rect -1723 -5306 -1707 -5260
rect -1661 -5306 -1645 -5260
rect -1553 -5278 -1468 -5232
rect -1422 -5278 -1403 -5232
rect -1553 -5305 -1403 -5278
rect -1723 -5323 -1645 -5306
rect -1884 -5344 -1806 -5327
rect -2993 -5421 -2937 -5377
rect -2833 -5421 -2777 -5377
rect -2673 -5421 -2617 -5344
rect -2513 -5421 -2457 -5344
rect -2353 -5421 -2297 -5377
rect -2193 -5421 -2137 -5377
rect -2033 -5421 -1977 -5344
rect -1873 -5421 -1817 -5344
rect -1713 -5421 -1657 -5377
rect -1553 -5421 -1497 -5377
rect -2993 -6065 -2937 -6021
rect -3086 -6081 -2937 -6065
rect -2833 -6073 -2777 -6021
rect -2673 -6065 -2617 -6021
rect -2513 -6065 -2457 -6021
rect -3086 -6127 -3068 -6081
rect -3022 -6127 -2937 -6081
rect -3086 -6147 -2937 -6127
rect -2849 -6093 -2762 -6073
rect -2353 -6075 -2297 -6021
rect -2193 -6075 -2137 -6021
rect -2033 -6065 -1977 -6021
rect -1873 -6065 -1817 -6021
rect -1713 -6073 -1657 -6021
rect -1553 -6065 -1497 -6021
rect -2849 -6139 -2828 -6093
rect -2782 -6139 -2762 -6093
rect -2849 -6153 -2762 -6139
rect -2370 -6093 -2283 -6075
rect -2370 -6139 -2348 -6093
rect -2302 -6139 -2283 -6093
rect -2370 -6155 -2283 -6139
rect -2207 -6093 -2120 -6075
rect -2207 -6139 -2188 -6093
rect -2142 -6139 -2120 -6093
rect -2207 -6155 -2120 -6139
rect -1728 -6093 -1641 -6073
rect -1728 -6139 -1708 -6093
rect -1662 -6139 -1641 -6093
rect -1728 -6153 -1641 -6139
rect -1553 -6085 -1403 -6065
rect -1553 -6131 -1468 -6085
rect -1422 -6131 -1403 -6085
rect -1553 -6152 -1403 -6131
<< polycontact >>
rect -3068 -4426 -3022 -4380
rect -2667 -4466 -2621 -4420
rect -2507 -4466 -2461 -4420
rect -2029 -4466 -1983 -4420
rect -1869 -4466 -1823 -4420
rect -1468 -4427 -1422 -4381
rect -3068 -5277 -3022 -5231
rect -2829 -5306 -2783 -5260
rect -2668 -5327 -2622 -5281
rect -2508 -5328 -2462 -5282
rect -2348 -5309 -2302 -5263
rect -2188 -5309 -2142 -5263
rect -2028 -5328 -1982 -5282
rect -1868 -5327 -1822 -5281
rect -1707 -5306 -1661 -5260
rect -1468 -5278 -1422 -5232
rect -3068 -6127 -3022 -6081
rect -2828 -6139 -2782 -6093
rect -2348 -6139 -2302 -6093
rect -2188 -6139 -2142 -6093
rect -1708 -6139 -1662 -6093
rect -1468 -6131 -1422 -6085
<< metal1 >>
rect -3293 -4286 -3195 -4270
rect -3293 -4332 -3267 -4286
rect -3221 -4332 -3195 -4286
rect -1317 -4286 -1219 -4270
rect -3293 -4380 -3195 -4332
rect -3068 -4373 -3022 -4315
rect -1468 -4369 -1422 -4315
rect -1317 -4332 -1291 -4286
rect -1245 -4332 -1219 -4286
rect -3293 -4426 -3267 -4380
rect -3221 -4426 -3195 -4380
rect -3293 -4474 -3195 -4426
rect -3080 -4380 -3010 -4373
rect -3080 -4426 -3068 -4380
rect -3022 -4426 -3010 -4380
rect -1480 -4381 -1410 -4369
rect -1745 -4404 -1644 -4386
rect -1745 -4415 -1726 -4404
rect -3080 -4439 -3010 -4426
rect -2688 -4420 -1726 -4415
rect -2688 -4466 -2667 -4420
rect -2621 -4466 -2507 -4420
rect -2461 -4466 -2029 -4420
rect -1983 -4466 -1869 -4420
rect -1823 -4465 -1726 -4420
rect -1664 -4465 -1644 -4404
rect -1480 -4427 -1468 -4381
rect -1422 -4427 -1410 -4381
rect -1480 -4439 -1410 -4427
rect -1317 -4380 -1219 -4332
rect -1317 -4426 -1291 -4380
rect -1245 -4426 -1219 -4380
rect -1823 -4466 -1644 -4465
rect -2688 -4471 -1644 -4466
rect -3293 -4520 -3267 -4474
rect -3221 -4520 -3195 -4474
rect -1745 -4483 -1644 -4471
rect -1317 -4474 -1219 -4426
rect -3293 -4568 -3195 -4520
rect -3293 -4614 -3267 -4568
rect -3221 -4614 -3195 -4568
rect -1317 -4520 -1291 -4474
rect -1245 -4520 -1219 -4474
rect -1317 -4568 -1219 -4520
rect -3068 -4582 -3022 -4571
rect -2908 -4582 -2862 -4571
rect -2748 -4582 -2702 -4571
rect -2588 -4582 -2542 -4571
rect -2428 -4582 -2382 -4571
rect -2268 -4582 -2222 -4571
rect -2108 -4582 -2062 -4571
rect -1948 -4582 -1902 -4571
rect -1788 -4582 -1742 -4571
rect -1628 -4582 -1582 -4571
rect -1468 -4582 -1422 -4571
rect -3293 -4662 -3195 -4614
rect -3293 -4708 -3267 -4662
rect -3221 -4708 -3195 -4662
rect -1317 -4614 -1291 -4568
rect -1245 -4614 -1219 -4568
rect -1317 -4619 -1219 -4614
rect -1317 -4662 -1170 -4619
rect -3293 -4756 -3195 -4708
rect -2607 -4682 -2524 -4668
rect -2607 -4738 -2593 -4682
rect -2537 -4738 -2524 -4682
rect -2607 -4750 -2524 -4738
rect -1965 -4682 -1882 -4669
rect -1965 -4738 -1952 -4682
rect -1896 -4738 -1882 -4682
rect -1965 -4751 -1882 -4738
rect -1317 -4708 -1291 -4662
rect -1245 -4708 -1170 -4662
rect -3293 -4802 -3267 -4756
rect -3221 -4802 -3195 -4756
rect -3293 -4850 -3195 -4802
rect -1317 -4756 -1170 -4708
rect -1317 -4802 -1291 -4756
rect -1245 -4766 -1170 -4756
rect -1245 -4802 -1219 -4766
rect -3293 -4896 -3267 -4850
rect -3221 -4896 -3195 -4850
rect -3293 -4944 -3195 -4896
rect -2767 -4839 -2684 -4825
rect -2767 -4895 -2753 -4839
rect -2697 -4895 -2684 -4839
rect -2767 -4907 -2684 -4895
rect -2447 -4840 -2364 -4826
rect -2447 -4896 -2433 -4840
rect -2377 -4896 -2364 -4840
rect -2447 -4908 -2364 -4896
rect -2127 -4838 -2044 -4824
rect -2127 -4894 -2113 -4838
rect -2057 -4894 -2044 -4838
rect -2127 -4906 -2044 -4894
rect -1807 -4839 -1724 -4825
rect -1807 -4895 -1793 -4839
rect -1737 -4895 -1724 -4839
rect -1807 -4907 -1724 -4895
rect -1317 -4850 -1219 -4802
rect -1317 -4896 -1291 -4850
rect -1245 -4896 -1219 -4850
rect -3293 -4990 -3267 -4944
rect -3221 -4990 -3195 -4944
rect -1317 -4944 -1219 -4896
rect -3293 -5038 -3195 -4990
rect -3293 -5084 -3267 -5038
rect -3221 -5084 -3195 -5038
rect -3088 -4989 -3004 -4975
rect -3088 -5045 -3074 -4989
rect -3018 -5045 -3004 -4989
rect -3088 -5059 -3004 -5045
rect -2927 -4989 -2843 -4974
rect -2927 -5045 -2913 -4989
rect -2857 -5045 -2843 -4989
rect -2927 -5058 -2843 -5045
rect -2288 -4989 -2202 -4975
rect -2288 -5045 -2274 -4989
rect -2216 -5045 -2202 -4989
rect -2288 -5059 -2202 -5045
rect -1647 -4989 -1563 -4974
rect -1647 -5045 -1633 -4989
rect -1577 -5045 -1563 -4989
rect -1647 -5058 -1563 -5045
rect -1487 -4989 -1403 -4975
rect -1487 -5045 -1473 -4989
rect -1417 -5045 -1403 -4989
rect -1487 -5059 -1403 -5045
rect -1317 -4990 -1291 -4944
rect -1245 -4990 -1219 -4944
rect -1317 -5038 -1219 -4990
rect -3293 -5132 -3195 -5084
rect -3293 -5178 -3267 -5132
rect -3221 -5178 -3195 -5132
rect -1317 -5084 -1291 -5038
rect -1245 -5084 -1219 -5038
rect -1317 -5132 -1219 -5084
rect -3293 -5226 -3195 -5178
rect -3068 -5219 -3022 -5156
rect -2908 -5167 -2862 -5156
rect -2748 -5167 -2702 -5156
rect -2588 -5167 -2542 -5156
rect -2428 -5167 -2382 -5156
rect -2268 -5167 -2222 -5156
rect -2108 -5167 -2062 -5156
rect -1948 -5167 -1902 -5156
rect -1788 -5167 -1742 -5156
rect -1628 -5167 -1582 -5156
rect -3293 -5272 -3267 -5226
rect -3221 -5272 -3195 -5226
rect -3293 -5320 -3195 -5272
rect -3081 -5231 -3009 -5219
rect -1468 -5223 -1422 -5156
rect -1317 -5178 -1291 -5132
rect -1245 -5178 -1219 -5132
rect -3081 -5277 -3068 -5231
rect -3022 -5277 -3009 -5231
rect -1480 -5232 -1410 -5223
rect -3081 -5289 -3009 -5277
rect -2851 -5260 -2750 -5245
rect -2851 -5266 -2829 -5260
rect -2783 -5266 -2750 -5260
rect -3293 -5366 -3267 -5320
rect -3221 -5366 -3195 -5320
rect -2851 -5322 -2830 -5266
rect -2774 -5267 -2750 -5266
rect -2363 -5263 -2285 -5246
rect -2363 -5267 -2348 -5263
rect -2774 -5281 -2348 -5267
rect -2774 -5322 -2668 -5281
rect -2851 -5323 -2668 -5322
rect -2851 -5342 -2750 -5323
rect -2684 -5327 -2668 -5323
rect -2622 -5282 -2348 -5281
rect -2622 -5323 -2508 -5282
rect -2622 -5327 -2606 -5323
rect -2684 -5344 -2606 -5327
rect -2524 -5328 -2508 -5323
rect -2462 -5309 -2348 -5282
rect -2302 -5267 -2285 -5263
rect -2205 -5263 -2127 -5246
rect -2205 -5267 -2188 -5263
rect -2302 -5309 -2188 -5267
rect -2142 -5267 -2127 -5263
rect -1723 -5260 -1645 -5246
rect -1723 -5267 -1707 -5260
rect -2142 -5281 -1707 -5267
rect -2142 -5282 -1868 -5281
rect -2142 -5309 -2028 -5282
rect -2462 -5323 -2028 -5309
rect -2462 -5328 -2446 -5323
rect -2524 -5344 -2446 -5328
rect -2044 -5328 -2028 -5323
rect -1982 -5323 -1868 -5282
rect -1982 -5328 -1966 -5323
rect -2044 -5344 -1966 -5328
rect -1884 -5327 -1868 -5323
rect -1822 -5306 -1707 -5281
rect -1661 -5306 -1645 -5260
rect -1480 -5278 -1468 -5232
rect -1422 -5278 -1410 -5232
rect -1480 -5291 -1410 -5278
rect -1317 -5226 -1219 -5178
rect -1317 -5272 -1291 -5226
rect -1245 -5272 -1219 -5226
rect -1822 -5323 -1645 -5306
rect -1317 -5320 -1219 -5272
rect -1822 -5327 -1806 -5323
rect -1884 -5344 -1806 -5327
rect -3293 -5414 -3195 -5366
rect -3293 -5460 -3267 -5414
rect -3221 -5460 -3195 -5414
rect -1317 -5366 -1291 -5320
rect -1245 -5366 -1219 -5320
rect -1317 -5414 -1219 -5366
rect -3068 -5434 -3022 -5423
rect -2908 -5434 -2862 -5423
rect -2748 -5434 -2702 -5423
rect -2588 -5434 -2542 -5423
rect -2428 -5434 -2382 -5423
rect -2268 -5434 -2222 -5423
rect -2108 -5434 -2062 -5423
rect -1948 -5434 -1902 -5423
rect -1788 -5434 -1742 -5423
rect -1628 -5434 -1582 -5423
rect -1468 -5434 -1422 -5423
rect -3293 -5508 -3195 -5460
rect -3293 -5554 -3267 -5508
rect -3221 -5554 -3195 -5508
rect -1317 -5460 -1291 -5414
rect -1245 -5460 -1219 -5414
rect -1317 -5469 -1219 -5460
rect -1317 -5508 -1170 -5469
rect -3293 -5602 -3195 -5554
rect -3293 -5648 -3267 -5602
rect -3221 -5648 -3195 -5602
rect -2607 -5542 -2524 -5528
rect -2607 -5598 -2593 -5542
rect -2537 -5598 -2524 -5542
rect -2607 -5610 -2524 -5598
rect -1965 -5542 -1882 -5527
rect -1965 -5598 -1952 -5542
rect -1896 -5598 -1882 -5542
rect -1965 -5611 -1882 -5598
rect -1317 -5554 -1291 -5508
rect -1245 -5554 -1170 -5508
rect -1317 -5602 -1170 -5554
rect -3293 -5696 -3195 -5648
rect -1317 -5648 -1291 -5602
rect -1245 -5616 -1170 -5602
rect -1245 -5648 -1219 -5616
rect -3293 -5742 -3267 -5696
rect -3221 -5742 -3195 -5696
rect -3293 -5790 -3195 -5742
rect -2769 -5694 -2686 -5680
rect -2769 -5750 -2755 -5694
rect -2699 -5750 -2686 -5694
rect -2769 -5762 -2686 -5750
rect -2447 -5693 -2364 -5679
rect -2447 -5749 -2433 -5693
rect -2377 -5749 -2364 -5693
rect -2447 -5761 -2364 -5749
rect -2129 -5693 -2046 -5679
rect -2129 -5749 -2115 -5693
rect -2059 -5749 -2046 -5693
rect -2129 -5761 -2046 -5749
rect -1806 -5693 -1723 -5679
rect -1806 -5749 -1792 -5693
rect -1736 -5749 -1723 -5693
rect -1806 -5761 -1723 -5749
rect -1317 -5696 -1219 -5648
rect -1317 -5742 -1291 -5696
rect -1245 -5742 -1219 -5696
rect -3293 -5836 -3267 -5790
rect -3221 -5836 -3195 -5790
rect -1317 -5790 -1219 -5742
rect -3293 -5884 -3195 -5836
rect -3293 -5930 -3267 -5884
rect -3221 -5930 -3195 -5884
rect -3088 -5849 -3004 -5835
rect -3088 -5905 -3074 -5849
rect -3018 -5905 -3004 -5849
rect -3088 -5919 -3004 -5905
rect -2927 -5849 -2843 -5834
rect -2927 -5905 -2913 -5849
rect -2857 -5905 -2843 -5849
rect -2927 -5918 -2843 -5905
rect -2288 -5849 -2202 -5835
rect -2288 -5905 -2274 -5849
rect -2216 -5905 -2202 -5849
rect -2288 -5919 -2202 -5905
rect -1647 -5849 -1563 -5834
rect -1647 -5905 -1633 -5849
rect -1577 -5905 -1563 -5849
rect -1647 -5918 -1563 -5905
rect -1487 -5849 -1403 -5835
rect -1487 -5905 -1473 -5849
rect -1417 -5905 -1403 -5849
rect -1487 -5919 -1403 -5905
rect -1317 -5836 -1291 -5790
rect -1245 -5836 -1219 -5790
rect -1317 -5884 -1219 -5836
rect -3293 -5978 -3195 -5930
rect -3293 -6024 -3267 -5978
rect -3221 -6024 -3195 -5978
rect -1317 -5930 -1291 -5884
rect -1245 -5930 -1219 -5884
rect -1317 -5978 -1219 -5930
rect -3293 -6072 -3195 -6024
rect -3068 -6069 -3022 -6008
rect -2908 -6019 -2862 -6008
rect -2748 -6019 -2702 -6008
rect -2588 -6019 -2542 -6008
rect -2428 -6019 -2382 -6008
rect -2268 -6019 -2222 -6008
rect -2108 -6019 -2062 -6008
rect -1948 -6019 -1902 -6008
rect -1788 -6019 -1742 -6008
rect -1628 -6019 -1582 -6008
rect -3293 -6118 -3267 -6072
rect -3221 -6118 -3195 -6072
rect -3293 -6166 -3195 -6118
rect -3080 -6081 -3011 -6069
rect -3080 -6127 -3068 -6081
rect -3022 -6127 -3011 -6081
rect -1742 -6087 -1641 -6066
rect -1468 -6074 -1422 -6008
rect -1317 -6024 -1291 -5978
rect -1245 -6011 -1219 -5978
rect -1245 -6024 -1170 -6011
rect -1317 -6072 -1170 -6024
rect -3080 -6139 -3011 -6127
rect -2849 -6093 -1721 -6087
rect -1665 -6093 -1641 -6087
rect -2849 -6139 -2828 -6093
rect -2782 -6139 -2348 -6093
rect -2302 -6139 -2188 -6093
rect -2142 -6139 -1721 -6093
rect -1662 -6139 -1641 -6093
rect -2849 -6143 -1721 -6139
rect -1665 -6143 -1641 -6139
rect -1481 -6085 -1410 -6074
rect -1481 -6131 -1468 -6085
rect -1422 -6131 -1410 -6085
rect -1481 -6143 -1410 -6131
rect -1317 -6118 -1291 -6072
rect -1245 -6118 -1170 -6072
rect -1742 -6163 -1641 -6143
rect -1317 -6158 -1170 -6118
rect -3293 -6212 -3267 -6166
rect -3221 -6212 -3195 -6166
rect -3293 -6234 -3195 -6212
rect -1317 -6166 -1219 -6158
rect -1317 -6212 -1291 -6166
rect -1245 -6212 -1219 -6166
rect -1317 -6234 -1219 -6212
rect -3293 -6260 -1219 -6234
rect -3293 -6306 -3266 -6260
rect -3220 -6306 -3172 -6260
rect -3126 -6306 -3078 -6260
rect -3032 -6306 -2984 -6260
rect -2938 -6306 -2890 -6260
rect -2844 -6306 -2796 -6260
rect -2750 -6306 -2702 -6260
rect -2656 -6306 -2608 -6260
rect -2562 -6306 -2514 -6260
rect -2468 -6306 -2420 -6260
rect -2374 -6306 -2326 -6260
rect -2280 -6306 -2232 -6260
rect -2186 -6306 -2138 -6260
rect -2092 -6306 -2044 -6260
rect -1998 -6306 -1950 -6260
rect -1904 -6306 -1856 -6260
rect -1810 -6306 -1762 -6260
rect -1716 -6306 -1668 -6260
rect -1622 -6306 -1574 -6260
rect -1528 -6306 -1480 -6260
rect -1434 -6306 -1386 -6260
rect -1340 -6306 -1292 -6260
rect -1246 -6306 -1219 -6260
rect -3293 -6332 -1219 -6306
<< via1 >>
rect -1726 -4465 -1664 -4404
rect -2593 -4738 -2537 -4682
rect -1952 -4738 -1896 -4682
rect -2753 -4895 -2697 -4839
rect -2433 -4896 -2377 -4840
rect -2113 -4894 -2057 -4838
rect -1793 -4895 -1737 -4839
rect -3074 -5045 -3018 -4989
rect -2913 -5045 -2857 -4989
rect -2274 -5045 -2216 -4989
rect -1633 -5045 -1577 -4989
rect -1473 -5045 -1417 -4989
rect -2830 -5306 -2829 -5266
rect -2829 -5306 -2783 -5266
rect -2783 -5306 -2774 -5266
rect -2830 -5322 -2774 -5306
rect -2593 -5598 -2537 -5542
rect -1952 -5598 -1896 -5542
rect -2755 -5750 -2699 -5694
rect -2433 -5749 -2377 -5693
rect -2115 -5749 -2059 -5693
rect -1792 -5749 -1736 -5693
rect -3074 -5905 -3018 -5849
rect -2913 -5905 -2857 -5849
rect -2274 -5905 -2216 -5849
rect -1633 -5905 -1577 -5849
rect -1473 -5905 -1417 -5849
rect -1721 -6093 -1665 -6087
rect -1721 -6139 -1708 -6093
rect -1708 -6139 -1665 -6093
rect -1721 -6143 -1665 -6139
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_2
timestamp 1692683681
transform -1 0 -1925 0 -1 -4869
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_3
timestamp 1692683681
transform -1 0 -1925 0 -1 -5721
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_4
timestamp 1692683681
transform 1 0 -2565 0 -1 -4869
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_5
timestamp 1692683681
transform 1 0 -2565 0 -1 -5721
box -282 -430 282 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_8
timestamp 1692683681
transform -1 0 -1525 0 -1 -4869
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_9
timestamp 1692683681
transform -1 0 -1685 0 -1 -4869
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_10
timestamp 1692683681
transform -1 0 -2165 0 -1 -4869
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_11
timestamp 1692683681
transform -1 0 -1685 0 -1 -5721
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_12
timestamp 1692683681
transform -1 0 -1525 0 -1 -5721
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_13
timestamp 1692683681
transform -1 0 -2165 0 -1 -5721
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_16
timestamp 1692683681
transform 1 0 -2805 0 -1 -4869
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_17
timestamp 1692683681
transform 1 0 -2965 0 -1 -4869
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_18
timestamp 1692683681
transform 1 0 -2325 0 -1 -4869
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_20
timestamp 1692683681
transform 1 0 -2805 0 -1 -5721
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_21
timestamp 1692683681
transform 1 0 -2965 0 -1 -5721
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_22
timestamp 1692683681
transform 1 0 -2325 0 -1 -5721
box -202 -430 202 430
<< end >>
