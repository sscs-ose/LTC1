magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1305 1019 1305
<< metal1 >>
rect -19 299 19 305
rect -19 -299 -13 299
rect 13 -299 19 299
rect -19 -305 19 -299
<< via1 >>
rect -13 -299 13 299
<< metal2 >>
rect -19 299 19 305
rect -19 -299 -13 299
rect 13 -299 19 299
rect -19 -305 19 -299
<< end >>
