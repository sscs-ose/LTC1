magic
tech gf180mcuC
magscale 1 10
timestamp 1694760847
<< metal1 >>
rect 8531 9224 8884 9253
rect 8531 9048 8575 9224
rect 8830 9048 8884 9224
rect 8531 9005 8884 9048
rect 7909 -453 8620 -372
rect 7909 -774 7971 -453
rect 8552 -774 8620 -453
rect 7909 -826 8620 -774
<< via1 >>
rect 8575 9048 8830 9224
rect 7971 -774 8552 -453
<< metal2 >>
rect 8531 9224 8884 9253
rect 8531 9048 8575 9224
rect 8830 9048 8884 9224
rect 8531 9005 8884 9048
rect 7909 -453 8620 -372
rect 7909 -774 7971 -453
rect 8552 -774 8620 -453
rect 7909 -826 8620 -774
<< via2 >>
rect 8575 9048 8830 9224
rect 7971 -774 8552 -453
<< metal3 >>
rect 8531 9224 8884 9253
rect 8531 9048 8575 9224
rect 8830 9048 8884 9224
rect 8531 9005 8884 9048
rect 7909 -453 8620 -372
rect 7909 -774 7971 -453
rect 8552 -774 8620 -453
rect 7909 -826 8620 -774
<< via3 >>
rect 8575 9048 8830 9224
rect 7971 -774 8552 -453
<< metal4 >>
rect 8531 9224 8884 9253
rect 8531 9048 8575 9224
rect 8830 9048 8884 9224
rect 8531 9005 8884 9048
rect 7909 -453 8620 -372
rect 7909 -774 7971 -453
rect 8552 -774 8620 -453
rect 7909 -826 8620 -774
<< via4 >>
rect 8575 9048 8830 9224
rect 7971 -774 8552 -453
<< metal5 >>
rect 8531 9224 8884 9253
rect 8531 9048 8575 9224
rect 8830 9048 8884 9224
rect 8531 9005 8884 9048
rect 8710 8683 8798 9005
rect 8078 -372 8409 217
rect 7909 -453 8620 -372
rect 7909 -774 7971 -453
rect 8552 -774 8620 -453
rect 7909 -826 8620 -774
use mim_2p0fF_WS3THJ  mim_2p0fF_WS3THJ_0
timestamp 1694760847
transform 1 0 4370 0 1 4370
box -4490 -4370 4490 4370
<< labels >>
flabel via4 8135 -616 8135 -616 0 FreeSans 800 0 0 0 Pp
port 0 nsew
flabel via4 8665 9137 8665 9137 0 FreeSans 800 0 0 0 Nn
port 1 nsew
<< end >>
