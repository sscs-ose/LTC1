magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2395 -11745 2395 11745
<< psubdiff >>
rect -395 9723 395 9745
rect -395 -9723 -373 9723
rect 373 -9723 395 9723
rect -395 -9745 395 -9723
<< psubdiffcont >>
rect -373 -9723 373 9723
<< metal1 >>
rect -384 9723 384 9734
rect -384 -9723 -373 9723
rect 373 -9723 384 9723
rect -384 -9734 384 -9723
<< end >>
