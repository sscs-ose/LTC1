magic
tech gf180mcuC
magscale 1 10
timestamp 1692681704
<< nwell >>
rect 0 0 580 468
<< pwell >>
rect 0 -228 580 -30
<< nmos >>
rect 178 -154 234 -104
rect 346 -154 402 -104
<< pmos >>
rect 178 136 234 186
rect 346 136 402 186
<< ndiff >>
rect 86 -104 158 -93
rect 254 -104 326 -93
rect 422 -104 494 -93
rect 86 -106 178 -104
rect 86 -152 99 -106
rect 145 -152 178 -106
rect 86 -154 178 -152
rect 234 -106 346 -104
rect 234 -152 267 -106
rect 313 -152 346 -106
rect 234 -154 346 -152
rect 402 -106 494 -104
rect 402 -152 435 -106
rect 481 -152 494 -106
rect 402 -154 494 -152
rect 86 -165 158 -154
rect 254 -165 326 -154
rect 422 -165 494 -154
<< pdiff >>
rect 86 186 158 197
rect 254 186 326 197
rect 422 186 494 197
rect 86 184 178 186
rect 86 138 99 184
rect 145 138 178 184
rect 86 136 178 138
rect 234 184 346 186
rect 234 138 267 184
rect 313 138 346 184
rect 234 136 346 138
rect 402 184 494 186
rect 402 138 435 184
rect 481 138 494 184
rect 402 136 494 138
rect 86 125 158 136
rect 254 125 326 136
rect 422 125 494 136
<< ndiffc >>
rect 99 -152 145 -106
rect 267 -152 313 -106
rect 435 -152 481 -106
<< pdiffc >>
rect 99 138 145 184
rect 267 138 313 184
rect 435 138 481 184
<< psubdiff >>
rect 26 -324 554 -311
rect 26 -370 39 -324
rect 85 -370 150 -324
rect 196 -370 261 -324
rect 307 -370 372 -324
rect 418 -370 483 -324
rect 529 -370 554 -324
rect 26 -383 554 -370
<< nsubdiff >>
rect 26 431 554 444
rect 26 385 39 431
rect 85 385 150 431
rect 196 385 261 431
rect 307 385 372 431
rect 418 385 483 431
rect 529 385 554 431
rect 26 372 554 385
<< psubdiffcont >>
rect 39 -370 85 -324
rect 150 -370 196 -324
rect 261 -370 307 -324
rect 372 -370 418 -324
rect 483 -370 529 -324
<< nsubdiffcont >>
rect 39 385 85 431
rect 150 385 196 431
rect 261 385 307 431
rect 372 385 418 431
rect 483 385 529 431
<< polysilicon >>
rect 148 308 234 321
rect 148 262 161 308
rect 207 262 234 308
rect 148 249 234 262
rect 178 186 234 249
rect 346 186 402 230
rect 178 102 234 136
rect 346 102 402 136
rect 178 63 402 102
rect 178 -104 234 -60
rect 346 -104 402 63
rect 178 -198 234 -154
rect 346 -198 402 -154
rect 170 -211 242 -198
rect 170 -257 183 -211
rect 229 -257 242 -211
rect 170 -270 242 -257
<< polycontact >>
rect 161 262 207 308
rect 183 -257 229 -211
<< metal1 >>
rect 16 431 564 448
rect 16 385 39 431
rect 85 385 150 431
rect 196 385 261 431
rect 307 385 372 431
rect 418 385 483 431
rect 529 385 564 431
rect 16 368 564 385
rect 148 308 220 321
rect -34 262 161 308
rect 207 262 220 308
rect 148 249 220 262
rect 267 184 313 368
rect 88 138 99 184
rect 145 138 156 184
rect 256 138 267 184
rect 313 138 324 184
rect 424 138 435 184
rect 481 138 492 184
rect 99 90 145 138
rect 435 90 481 138
rect 99 44 481 90
rect 435 39 481 44
rect 435 -7 617 39
rect 435 -106 481 -7
rect 88 -152 99 -106
rect 145 -152 156 -106
rect 256 -152 267 -106
rect 313 -152 324 -106
rect 424 -152 435 -106
rect 481 -152 492 -106
rect 99 -198 145 -152
rect 267 -198 313 -152
rect 99 -211 313 -198
rect 99 -254 183 -211
rect 170 -257 183 -254
rect 229 -254 313 -211
rect 229 -257 242 -254
rect 170 -261 242 -257
rect 183 -307 229 -261
rect 16 -324 564 -307
rect 16 -370 39 -324
rect 85 -370 150 -324
rect 196 -370 261 -324
rect 307 -370 372 -324
rect 418 -370 483 -324
rect 529 -370 564 -324
rect 16 -387 564 -370
<< labels >>
flabel metal1 -12 285 -12 285 0 FreeSans 480 0 0 0 IN
port 0 nsew
flabel metal1 551 16 551 16 0 FreeSans 480 0 0 0 OUT
port 1 nsew
flabel nsubdiffcont 284 410 284 410 0 FreeSans 480 0 0 0 VDD
port 2 nsew
flabel psubdiffcont 284 -348 284 -348 0 FreeSans 480 0 0 0 VSS
port 3 nsew
<< end >>
