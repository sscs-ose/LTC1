magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1513 -3641 1513 3641
<< metal1 >>
rect -513 2635 513 2641
rect -513 2609 -507 2635
rect -481 2609 -431 2635
rect -405 2609 -355 2635
rect -329 2609 -279 2635
rect -253 2609 -203 2635
rect -177 2609 -127 2635
rect -101 2609 -51 2635
rect -25 2609 25 2635
rect 51 2609 101 2635
rect 127 2609 177 2635
rect 203 2609 253 2635
rect 279 2609 329 2635
rect 355 2609 405 2635
rect 431 2609 481 2635
rect 507 2609 513 2635
rect -513 2559 513 2609
rect -513 2533 -507 2559
rect -481 2533 -431 2559
rect -405 2533 -355 2559
rect -329 2533 -279 2559
rect -253 2533 -203 2559
rect -177 2533 -127 2559
rect -101 2533 -51 2559
rect -25 2533 25 2559
rect 51 2533 101 2559
rect 127 2533 177 2559
rect 203 2533 253 2559
rect 279 2533 329 2559
rect 355 2533 405 2559
rect 431 2533 481 2559
rect 507 2533 513 2559
rect -513 2483 513 2533
rect -513 2457 -507 2483
rect -481 2457 -431 2483
rect -405 2457 -355 2483
rect -329 2457 -279 2483
rect -253 2457 -203 2483
rect -177 2457 -127 2483
rect -101 2457 -51 2483
rect -25 2457 25 2483
rect 51 2457 101 2483
rect 127 2457 177 2483
rect 203 2457 253 2483
rect 279 2457 329 2483
rect 355 2457 405 2483
rect 431 2457 481 2483
rect 507 2457 513 2483
rect -513 2407 513 2457
rect -513 2381 -507 2407
rect -481 2381 -431 2407
rect -405 2381 -355 2407
rect -329 2381 -279 2407
rect -253 2381 -203 2407
rect -177 2381 -127 2407
rect -101 2381 -51 2407
rect -25 2381 25 2407
rect 51 2381 101 2407
rect 127 2381 177 2407
rect 203 2381 253 2407
rect 279 2381 329 2407
rect 355 2381 405 2407
rect 431 2381 481 2407
rect 507 2381 513 2407
rect -513 2331 513 2381
rect -513 2305 -507 2331
rect -481 2305 -431 2331
rect -405 2305 -355 2331
rect -329 2305 -279 2331
rect -253 2305 -203 2331
rect -177 2305 -127 2331
rect -101 2305 -51 2331
rect -25 2305 25 2331
rect 51 2305 101 2331
rect 127 2305 177 2331
rect 203 2305 253 2331
rect 279 2305 329 2331
rect 355 2305 405 2331
rect 431 2305 481 2331
rect 507 2305 513 2331
rect -513 2255 513 2305
rect -513 2229 -507 2255
rect -481 2229 -431 2255
rect -405 2229 -355 2255
rect -329 2229 -279 2255
rect -253 2229 -203 2255
rect -177 2229 -127 2255
rect -101 2229 -51 2255
rect -25 2229 25 2255
rect 51 2229 101 2255
rect 127 2229 177 2255
rect 203 2229 253 2255
rect 279 2229 329 2255
rect 355 2229 405 2255
rect 431 2229 481 2255
rect 507 2229 513 2255
rect -513 2179 513 2229
rect -513 2153 -507 2179
rect -481 2153 -431 2179
rect -405 2153 -355 2179
rect -329 2153 -279 2179
rect -253 2153 -203 2179
rect -177 2153 -127 2179
rect -101 2153 -51 2179
rect -25 2153 25 2179
rect 51 2153 101 2179
rect 127 2153 177 2179
rect 203 2153 253 2179
rect 279 2153 329 2179
rect 355 2153 405 2179
rect 431 2153 481 2179
rect 507 2153 513 2179
rect -513 2103 513 2153
rect -513 2077 -507 2103
rect -481 2077 -431 2103
rect -405 2077 -355 2103
rect -329 2077 -279 2103
rect -253 2077 -203 2103
rect -177 2077 -127 2103
rect -101 2077 -51 2103
rect -25 2077 25 2103
rect 51 2077 101 2103
rect 127 2077 177 2103
rect 203 2077 253 2103
rect 279 2077 329 2103
rect 355 2077 405 2103
rect 431 2077 481 2103
rect 507 2077 513 2103
rect -513 2027 513 2077
rect -513 2001 -507 2027
rect -481 2001 -431 2027
rect -405 2001 -355 2027
rect -329 2001 -279 2027
rect -253 2001 -203 2027
rect -177 2001 -127 2027
rect -101 2001 -51 2027
rect -25 2001 25 2027
rect 51 2001 101 2027
rect 127 2001 177 2027
rect 203 2001 253 2027
rect 279 2001 329 2027
rect 355 2001 405 2027
rect 431 2001 481 2027
rect 507 2001 513 2027
rect -513 1951 513 2001
rect -513 1925 -507 1951
rect -481 1925 -431 1951
rect -405 1925 -355 1951
rect -329 1925 -279 1951
rect -253 1925 -203 1951
rect -177 1925 -127 1951
rect -101 1925 -51 1951
rect -25 1925 25 1951
rect 51 1925 101 1951
rect 127 1925 177 1951
rect 203 1925 253 1951
rect 279 1925 329 1951
rect 355 1925 405 1951
rect 431 1925 481 1951
rect 507 1925 513 1951
rect -513 1875 513 1925
rect -513 1849 -507 1875
rect -481 1849 -431 1875
rect -405 1849 -355 1875
rect -329 1849 -279 1875
rect -253 1849 -203 1875
rect -177 1849 -127 1875
rect -101 1849 -51 1875
rect -25 1849 25 1875
rect 51 1849 101 1875
rect 127 1849 177 1875
rect 203 1849 253 1875
rect 279 1849 329 1875
rect 355 1849 405 1875
rect 431 1849 481 1875
rect 507 1849 513 1875
rect -513 1799 513 1849
rect -513 1773 -507 1799
rect -481 1773 -431 1799
rect -405 1773 -355 1799
rect -329 1773 -279 1799
rect -253 1773 -203 1799
rect -177 1773 -127 1799
rect -101 1773 -51 1799
rect -25 1773 25 1799
rect 51 1773 101 1799
rect 127 1773 177 1799
rect 203 1773 253 1799
rect 279 1773 329 1799
rect 355 1773 405 1799
rect 431 1773 481 1799
rect 507 1773 513 1799
rect -513 1723 513 1773
rect -513 1697 -507 1723
rect -481 1697 -431 1723
rect -405 1697 -355 1723
rect -329 1697 -279 1723
rect -253 1697 -203 1723
rect -177 1697 -127 1723
rect -101 1697 -51 1723
rect -25 1697 25 1723
rect 51 1697 101 1723
rect 127 1697 177 1723
rect 203 1697 253 1723
rect 279 1697 329 1723
rect 355 1697 405 1723
rect 431 1697 481 1723
rect 507 1697 513 1723
rect -513 1647 513 1697
rect -513 1621 -507 1647
rect -481 1621 -431 1647
rect -405 1621 -355 1647
rect -329 1621 -279 1647
rect -253 1621 -203 1647
rect -177 1621 -127 1647
rect -101 1621 -51 1647
rect -25 1621 25 1647
rect 51 1621 101 1647
rect 127 1621 177 1647
rect 203 1621 253 1647
rect 279 1621 329 1647
rect 355 1621 405 1647
rect 431 1621 481 1647
rect 507 1621 513 1647
rect -513 1571 513 1621
rect -513 1545 -507 1571
rect -481 1545 -431 1571
rect -405 1545 -355 1571
rect -329 1545 -279 1571
rect -253 1545 -203 1571
rect -177 1545 -127 1571
rect -101 1545 -51 1571
rect -25 1545 25 1571
rect 51 1545 101 1571
rect 127 1545 177 1571
rect 203 1545 253 1571
rect 279 1545 329 1571
rect 355 1545 405 1571
rect 431 1545 481 1571
rect 507 1545 513 1571
rect -513 1495 513 1545
rect -513 1469 -507 1495
rect -481 1469 -431 1495
rect -405 1469 -355 1495
rect -329 1469 -279 1495
rect -253 1469 -203 1495
rect -177 1469 -127 1495
rect -101 1469 -51 1495
rect -25 1469 25 1495
rect 51 1469 101 1495
rect 127 1469 177 1495
rect 203 1469 253 1495
rect 279 1469 329 1495
rect 355 1469 405 1495
rect 431 1469 481 1495
rect 507 1469 513 1495
rect -513 1419 513 1469
rect -513 1393 -507 1419
rect -481 1393 -431 1419
rect -405 1393 -355 1419
rect -329 1393 -279 1419
rect -253 1393 -203 1419
rect -177 1393 -127 1419
rect -101 1393 -51 1419
rect -25 1393 25 1419
rect 51 1393 101 1419
rect 127 1393 177 1419
rect 203 1393 253 1419
rect 279 1393 329 1419
rect 355 1393 405 1419
rect 431 1393 481 1419
rect 507 1393 513 1419
rect -513 1343 513 1393
rect -513 1317 -507 1343
rect -481 1317 -431 1343
rect -405 1317 -355 1343
rect -329 1317 -279 1343
rect -253 1317 -203 1343
rect -177 1317 -127 1343
rect -101 1317 -51 1343
rect -25 1317 25 1343
rect 51 1317 101 1343
rect 127 1317 177 1343
rect 203 1317 253 1343
rect 279 1317 329 1343
rect 355 1317 405 1343
rect 431 1317 481 1343
rect 507 1317 513 1343
rect -513 1267 513 1317
rect -513 1241 -507 1267
rect -481 1241 -431 1267
rect -405 1241 -355 1267
rect -329 1241 -279 1267
rect -253 1241 -203 1267
rect -177 1241 -127 1267
rect -101 1241 -51 1267
rect -25 1241 25 1267
rect 51 1241 101 1267
rect 127 1241 177 1267
rect 203 1241 253 1267
rect 279 1241 329 1267
rect 355 1241 405 1267
rect 431 1241 481 1267
rect 507 1241 513 1267
rect -513 1191 513 1241
rect -513 1165 -507 1191
rect -481 1165 -431 1191
rect -405 1165 -355 1191
rect -329 1165 -279 1191
rect -253 1165 -203 1191
rect -177 1165 -127 1191
rect -101 1165 -51 1191
rect -25 1165 25 1191
rect 51 1165 101 1191
rect 127 1165 177 1191
rect 203 1165 253 1191
rect 279 1165 329 1191
rect 355 1165 405 1191
rect 431 1165 481 1191
rect 507 1165 513 1191
rect -513 1115 513 1165
rect -513 1089 -507 1115
rect -481 1089 -431 1115
rect -405 1089 -355 1115
rect -329 1089 -279 1115
rect -253 1089 -203 1115
rect -177 1089 -127 1115
rect -101 1089 -51 1115
rect -25 1089 25 1115
rect 51 1089 101 1115
rect 127 1089 177 1115
rect 203 1089 253 1115
rect 279 1089 329 1115
rect 355 1089 405 1115
rect 431 1089 481 1115
rect 507 1089 513 1115
rect -513 1039 513 1089
rect -513 1013 -507 1039
rect -481 1013 -431 1039
rect -405 1013 -355 1039
rect -329 1013 -279 1039
rect -253 1013 -203 1039
rect -177 1013 -127 1039
rect -101 1013 -51 1039
rect -25 1013 25 1039
rect 51 1013 101 1039
rect 127 1013 177 1039
rect 203 1013 253 1039
rect 279 1013 329 1039
rect 355 1013 405 1039
rect 431 1013 481 1039
rect 507 1013 513 1039
rect -513 963 513 1013
rect -513 937 -507 963
rect -481 937 -431 963
rect -405 937 -355 963
rect -329 937 -279 963
rect -253 937 -203 963
rect -177 937 -127 963
rect -101 937 -51 963
rect -25 937 25 963
rect 51 937 101 963
rect 127 937 177 963
rect 203 937 253 963
rect 279 937 329 963
rect 355 937 405 963
rect 431 937 481 963
rect 507 937 513 963
rect -513 887 513 937
rect -513 861 -507 887
rect -481 861 -431 887
rect -405 861 -355 887
rect -329 861 -279 887
rect -253 861 -203 887
rect -177 861 -127 887
rect -101 861 -51 887
rect -25 861 25 887
rect 51 861 101 887
rect 127 861 177 887
rect 203 861 253 887
rect 279 861 329 887
rect 355 861 405 887
rect 431 861 481 887
rect 507 861 513 887
rect -513 811 513 861
rect -513 785 -507 811
rect -481 785 -431 811
rect -405 785 -355 811
rect -329 785 -279 811
rect -253 785 -203 811
rect -177 785 -127 811
rect -101 785 -51 811
rect -25 785 25 811
rect 51 785 101 811
rect 127 785 177 811
rect 203 785 253 811
rect 279 785 329 811
rect 355 785 405 811
rect 431 785 481 811
rect 507 785 513 811
rect -513 735 513 785
rect -513 709 -507 735
rect -481 709 -431 735
rect -405 709 -355 735
rect -329 709 -279 735
rect -253 709 -203 735
rect -177 709 -127 735
rect -101 709 -51 735
rect -25 709 25 735
rect 51 709 101 735
rect 127 709 177 735
rect 203 709 253 735
rect 279 709 329 735
rect 355 709 405 735
rect 431 709 481 735
rect 507 709 513 735
rect -513 659 513 709
rect -513 633 -507 659
rect -481 633 -431 659
rect -405 633 -355 659
rect -329 633 -279 659
rect -253 633 -203 659
rect -177 633 -127 659
rect -101 633 -51 659
rect -25 633 25 659
rect 51 633 101 659
rect 127 633 177 659
rect 203 633 253 659
rect 279 633 329 659
rect 355 633 405 659
rect 431 633 481 659
rect 507 633 513 659
rect -513 583 513 633
rect -513 557 -507 583
rect -481 557 -431 583
rect -405 557 -355 583
rect -329 557 -279 583
rect -253 557 -203 583
rect -177 557 -127 583
rect -101 557 -51 583
rect -25 557 25 583
rect 51 557 101 583
rect 127 557 177 583
rect 203 557 253 583
rect 279 557 329 583
rect 355 557 405 583
rect 431 557 481 583
rect 507 557 513 583
rect -513 507 513 557
rect -513 481 -507 507
rect -481 481 -431 507
rect -405 481 -355 507
rect -329 481 -279 507
rect -253 481 -203 507
rect -177 481 -127 507
rect -101 481 -51 507
rect -25 481 25 507
rect 51 481 101 507
rect 127 481 177 507
rect 203 481 253 507
rect 279 481 329 507
rect 355 481 405 507
rect 431 481 481 507
rect 507 481 513 507
rect -513 431 513 481
rect -513 405 -507 431
rect -481 405 -431 431
rect -405 405 -355 431
rect -329 405 -279 431
rect -253 405 -203 431
rect -177 405 -127 431
rect -101 405 -51 431
rect -25 405 25 431
rect 51 405 101 431
rect 127 405 177 431
rect 203 405 253 431
rect 279 405 329 431
rect 355 405 405 431
rect 431 405 481 431
rect 507 405 513 431
rect -513 355 513 405
rect -513 329 -507 355
rect -481 329 -431 355
rect -405 329 -355 355
rect -329 329 -279 355
rect -253 329 -203 355
rect -177 329 -127 355
rect -101 329 -51 355
rect -25 329 25 355
rect 51 329 101 355
rect 127 329 177 355
rect 203 329 253 355
rect 279 329 329 355
rect 355 329 405 355
rect 431 329 481 355
rect 507 329 513 355
rect -513 279 513 329
rect -513 253 -507 279
rect -481 253 -431 279
rect -405 253 -355 279
rect -329 253 -279 279
rect -253 253 -203 279
rect -177 253 -127 279
rect -101 253 -51 279
rect -25 253 25 279
rect 51 253 101 279
rect 127 253 177 279
rect 203 253 253 279
rect 279 253 329 279
rect 355 253 405 279
rect 431 253 481 279
rect 507 253 513 279
rect -513 203 513 253
rect -513 177 -507 203
rect -481 177 -431 203
rect -405 177 -355 203
rect -329 177 -279 203
rect -253 177 -203 203
rect -177 177 -127 203
rect -101 177 -51 203
rect -25 177 25 203
rect 51 177 101 203
rect 127 177 177 203
rect 203 177 253 203
rect 279 177 329 203
rect 355 177 405 203
rect 431 177 481 203
rect 507 177 513 203
rect -513 127 513 177
rect -513 101 -507 127
rect -481 101 -431 127
rect -405 101 -355 127
rect -329 101 -279 127
rect -253 101 -203 127
rect -177 101 -127 127
rect -101 101 -51 127
rect -25 101 25 127
rect 51 101 101 127
rect 127 101 177 127
rect 203 101 253 127
rect 279 101 329 127
rect 355 101 405 127
rect 431 101 481 127
rect 507 101 513 127
rect -513 51 513 101
rect -513 25 -507 51
rect -481 25 -431 51
rect -405 25 -355 51
rect -329 25 -279 51
rect -253 25 -203 51
rect -177 25 -127 51
rect -101 25 -51 51
rect -25 25 25 51
rect 51 25 101 51
rect 127 25 177 51
rect 203 25 253 51
rect 279 25 329 51
rect 355 25 405 51
rect 431 25 481 51
rect 507 25 513 51
rect -513 -25 513 25
rect -513 -51 -507 -25
rect -481 -51 -431 -25
rect -405 -51 -355 -25
rect -329 -51 -279 -25
rect -253 -51 -203 -25
rect -177 -51 -127 -25
rect -101 -51 -51 -25
rect -25 -51 25 -25
rect 51 -51 101 -25
rect 127 -51 177 -25
rect 203 -51 253 -25
rect 279 -51 329 -25
rect 355 -51 405 -25
rect 431 -51 481 -25
rect 507 -51 513 -25
rect -513 -101 513 -51
rect -513 -127 -507 -101
rect -481 -127 -431 -101
rect -405 -127 -355 -101
rect -329 -127 -279 -101
rect -253 -127 -203 -101
rect -177 -127 -127 -101
rect -101 -127 -51 -101
rect -25 -127 25 -101
rect 51 -127 101 -101
rect 127 -127 177 -101
rect 203 -127 253 -101
rect 279 -127 329 -101
rect 355 -127 405 -101
rect 431 -127 481 -101
rect 507 -127 513 -101
rect -513 -177 513 -127
rect -513 -203 -507 -177
rect -481 -203 -431 -177
rect -405 -203 -355 -177
rect -329 -203 -279 -177
rect -253 -203 -203 -177
rect -177 -203 -127 -177
rect -101 -203 -51 -177
rect -25 -203 25 -177
rect 51 -203 101 -177
rect 127 -203 177 -177
rect 203 -203 253 -177
rect 279 -203 329 -177
rect 355 -203 405 -177
rect 431 -203 481 -177
rect 507 -203 513 -177
rect -513 -253 513 -203
rect -513 -279 -507 -253
rect -481 -279 -431 -253
rect -405 -279 -355 -253
rect -329 -279 -279 -253
rect -253 -279 -203 -253
rect -177 -279 -127 -253
rect -101 -279 -51 -253
rect -25 -279 25 -253
rect 51 -279 101 -253
rect 127 -279 177 -253
rect 203 -279 253 -253
rect 279 -279 329 -253
rect 355 -279 405 -253
rect 431 -279 481 -253
rect 507 -279 513 -253
rect -513 -329 513 -279
rect -513 -355 -507 -329
rect -481 -355 -431 -329
rect -405 -355 -355 -329
rect -329 -355 -279 -329
rect -253 -355 -203 -329
rect -177 -355 -127 -329
rect -101 -355 -51 -329
rect -25 -355 25 -329
rect 51 -355 101 -329
rect 127 -355 177 -329
rect 203 -355 253 -329
rect 279 -355 329 -329
rect 355 -355 405 -329
rect 431 -355 481 -329
rect 507 -355 513 -329
rect -513 -405 513 -355
rect -513 -431 -507 -405
rect -481 -431 -431 -405
rect -405 -431 -355 -405
rect -329 -431 -279 -405
rect -253 -431 -203 -405
rect -177 -431 -127 -405
rect -101 -431 -51 -405
rect -25 -431 25 -405
rect 51 -431 101 -405
rect 127 -431 177 -405
rect 203 -431 253 -405
rect 279 -431 329 -405
rect 355 -431 405 -405
rect 431 -431 481 -405
rect 507 -431 513 -405
rect -513 -481 513 -431
rect -513 -507 -507 -481
rect -481 -507 -431 -481
rect -405 -507 -355 -481
rect -329 -507 -279 -481
rect -253 -507 -203 -481
rect -177 -507 -127 -481
rect -101 -507 -51 -481
rect -25 -507 25 -481
rect 51 -507 101 -481
rect 127 -507 177 -481
rect 203 -507 253 -481
rect 279 -507 329 -481
rect 355 -507 405 -481
rect 431 -507 481 -481
rect 507 -507 513 -481
rect -513 -557 513 -507
rect -513 -583 -507 -557
rect -481 -583 -431 -557
rect -405 -583 -355 -557
rect -329 -583 -279 -557
rect -253 -583 -203 -557
rect -177 -583 -127 -557
rect -101 -583 -51 -557
rect -25 -583 25 -557
rect 51 -583 101 -557
rect 127 -583 177 -557
rect 203 -583 253 -557
rect 279 -583 329 -557
rect 355 -583 405 -557
rect 431 -583 481 -557
rect 507 -583 513 -557
rect -513 -633 513 -583
rect -513 -659 -507 -633
rect -481 -659 -431 -633
rect -405 -659 -355 -633
rect -329 -659 -279 -633
rect -253 -659 -203 -633
rect -177 -659 -127 -633
rect -101 -659 -51 -633
rect -25 -659 25 -633
rect 51 -659 101 -633
rect 127 -659 177 -633
rect 203 -659 253 -633
rect 279 -659 329 -633
rect 355 -659 405 -633
rect 431 -659 481 -633
rect 507 -659 513 -633
rect -513 -709 513 -659
rect -513 -735 -507 -709
rect -481 -735 -431 -709
rect -405 -735 -355 -709
rect -329 -735 -279 -709
rect -253 -735 -203 -709
rect -177 -735 -127 -709
rect -101 -735 -51 -709
rect -25 -735 25 -709
rect 51 -735 101 -709
rect 127 -735 177 -709
rect 203 -735 253 -709
rect 279 -735 329 -709
rect 355 -735 405 -709
rect 431 -735 481 -709
rect 507 -735 513 -709
rect -513 -785 513 -735
rect -513 -811 -507 -785
rect -481 -811 -431 -785
rect -405 -811 -355 -785
rect -329 -811 -279 -785
rect -253 -811 -203 -785
rect -177 -811 -127 -785
rect -101 -811 -51 -785
rect -25 -811 25 -785
rect 51 -811 101 -785
rect 127 -811 177 -785
rect 203 -811 253 -785
rect 279 -811 329 -785
rect 355 -811 405 -785
rect 431 -811 481 -785
rect 507 -811 513 -785
rect -513 -861 513 -811
rect -513 -887 -507 -861
rect -481 -887 -431 -861
rect -405 -887 -355 -861
rect -329 -887 -279 -861
rect -253 -887 -203 -861
rect -177 -887 -127 -861
rect -101 -887 -51 -861
rect -25 -887 25 -861
rect 51 -887 101 -861
rect 127 -887 177 -861
rect 203 -887 253 -861
rect 279 -887 329 -861
rect 355 -887 405 -861
rect 431 -887 481 -861
rect 507 -887 513 -861
rect -513 -937 513 -887
rect -513 -963 -507 -937
rect -481 -963 -431 -937
rect -405 -963 -355 -937
rect -329 -963 -279 -937
rect -253 -963 -203 -937
rect -177 -963 -127 -937
rect -101 -963 -51 -937
rect -25 -963 25 -937
rect 51 -963 101 -937
rect 127 -963 177 -937
rect 203 -963 253 -937
rect 279 -963 329 -937
rect 355 -963 405 -937
rect 431 -963 481 -937
rect 507 -963 513 -937
rect -513 -1013 513 -963
rect -513 -1039 -507 -1013
rect -481 -1039 -431 -1013
rect -405 -1039 -355 -1013
rect -329 -1039 -279 -1013
rect -253 -1039 -203 -1013
rect -177 -1039 -127 -1013
rect -101 -1039 -51 -1013
rect -25 -1039 25 -1013
rect 51 -1039 101 -1013
rect 127 -1039 177 -1013
rect 203 -1039 253 -1013
rect 279 -1039 329 -1013
rect 355 -1039 405 -1013
rect 431 -1039 481 -1013
rect 507 -1039 513 -1013
rect -513 -1089 513 -1039
rect -513 -1115 -507 -1089
rect -481 -1115 -431 -1089
rect -405 -1115 -355 -1089
rect -329 -1115 -279 -1089
rect -253 -1115 -203 -1089
rect -177 -1115 -127 -1089
rect -101 -1115 -51 -1089
rect -25 -1115 25 -1089
rect 51 -1115 101 -1089
rect 127 -1115 177 -1089
rect 203 -1115 253 -1089
rect 279 -1115 329 -1089
rect 355 -1115 405 -1089
rect 431 -1115 481 -1089
rect 507 -1115 513 -1089
rect -513 -1165 513 -1115
rect -513 -1191 -507 -1165
rect -481 -1191 -431 -1165
rect -405 -1191 -355 -1165
rect -329 -1191 -279 -1165
rect -253 -1191 -203 -1165
rect -177 -1191 -127 -1165
rect -101 -1191 -51 -1165
rect -25 -1191 25 -1165
rect 51 -1191 101 -1165
rect 127 -1191 177 -1165
rect 203 -1191 253 -1165
rect 279 -1191 329 -1165
rect 355 -1191 405 -1165
rect 431 -1191 481 -1165
rect 507 -1191 513 -1165
rect -513 -1241 513 -1191
rect -513 -1267 -507 -1241
rect -481 -1267 -431 -1241
rect -405 -1267 -355 -1241
rect -329 -1267 -279 -1241
rect -253 -1267 -203 -1241
rect -177 -1267 -127 -1241
rect -101 -1267 -51 -1241
rect -25 -1267 25 -1241
rect 51 -1267 101 -1241
rect 127 -1267 177 -1241
rect 203 -1267 253 -1241
rect 279 -1267 329 -1241
rect 355 -1267 405 -1241
rect 431 -1267 481 -1241
rect 507 -1267 513 -1241
rect -513 -1317 513 -1267
rect -513 -1343 -507 -1317
rect -481 -1343 -431 -1317
rect -405 -1343 -355 -1317
rect -329 -1343 -279 -1317
rect -253 -1343 -203 -1317
rect -177 -1343 -127 -1317
rect -101 -1343 -51 -1317
rect -25 -1343 25 -1317
rect 51 -1343 101 -1317
rect 127 -1343 177 -1317
rect 203 -1343 253 -1317
rect 279 -1343 329 -1317
rect 355 -1343 405 -1317
rect 431 -1343 481 -1317
rect 507 -1343 513 -1317
rect -513 -1393 513 -1343
rect -513 -1419 -507 -1393
rect -481 -1419 -431 -1393
rect -405 -1419 -355 -1393
rect -329 -1419 -279 -1393
rect -253 -1419 -203 -1393
rect -177 -1419 -127 -1393
rect -101 -1419 -51 -1393
rect -25 -1419 25 -1393
rect 51 -1419 101 -1393
rect 127 -1419 177 -1393
rect 203 -1419 253 -1393
rect 279 -1419 329 -1393
rect 355 -1419 405 -1393
rect 431 -1419 481 -1393
rect 507 -1419 513 -1393
rect -513 -1469 513 -1419
rect -513 -1495 -507 -1469
rect -481 -1495 -431 -1469
rect -405 -1495 -355 -1469
rect -329 -1495 -279 -1469
rect -253 -1495 -203 -1469
rect -177 -1495 -127 -1469
rect -101 -1495 -51 -1469
rect -25 -1495 25 -1469
rect 51 -1495 101 -1469
rect 127 -1495 177 -1469
rect 203 -1495 253 -1469
rect 279 -1495 329 -1469
rect 355 -1495 405 -1469
rect 431 -1495 481 -1469
rect 507 -1495 513 -1469
rect -513 -1545 513 -1495
rect -513 -1571 -507 -1545
rect -481 -1571 -431 -1545
rect -405 -1571 -355 -1545
rect -329 -1571 -279 -1545
rect -253 -1571 -203 -1545
rect -177 -1571 -127 -1545
rect -101 -1571 -51 -1545
rect -25 -1571 25 -1545
rect 51 -1571 101 -1545
rect 127 -1571 177 -1545
rect 203 -1571 253 -1545
rect 279 -1571 329 -1545
rect 355 -1571 405 -1545
rect 431 -1571 481 -1545
rect 507 -1571 513 -1545
rect -513 -1621 513 -1571
rect -513 -1647 -507 -1621
rect -481 -1647 -431 -1621
rect -405 -1647 -355 -1621
rect -329 -1647 -279 -1621
rect -253 -1647 -203 -1621
rect -177 -1647 -127 -1621
rect -101 -1647 -51 -1621
rect -25 -1647 25 -1621
rect 51 -1647 101 -1621
rect 127 -1647 177 -1621
rect 203 -1647 253 -1621
rect 279 -1647 329 -1621
rect 355 -1647 405 -1621
rect 431 -1647 481 -1621
rect 507 -1647 513 -1621
rect -513 -1697 513 -1647
rect -513 -1723 -507 -1697
rect -481 -1723 -431 -1697
rect -405 -1723 -355 -1697
rect -329 -1723 -279 -1697
rect -253 -1723 -203 -1697
rect -177 -1723 -127 -1697
rect -101 -1723 -51 -1697
rect -25 -1723 25 -1697
rect 51 -1723 101 -1697
rect 127 -1723 177 -1697
rect 203 -1723 253 -1697
rect 279 -1723 329 -1697
rect 355 -1723 405 -1697
rect 431 -1723 481 -1697
rect 507 -1723 513 -1697
rect -513 -1773 513 -1723
rect -513 -1799 -507 -1773
rect -481 -1799 -431 -1773
rect -405 -1799 -355 -1773
rect -329 -1799 -279 -1773
rect -253 -1799 -203 -1773
rect -177 -1799 -127 -1773
rect -101 -1799 -51 -1773
rect -25 -1799 25 -1773
rect 51 -1799 101 -1773
rect 127 -1799 177 -1773
rect 203 -1799 253 -1773
rect 279 -1799 329 -1773
rect 355 -1799 405 -1773
rect 431 -1799 481 -1773
rect 507 -1799 513 -1773
rect -513 -1849 513 -1799
rect -513 -1875 -507 -1849
rect -481 -1875 -431 -1849
rect -405 -1875 -355 -1849
rect -329 -1875 -279 -1849
rect -253 -1875 -203 -1849
rect -177 -1875 -127 -1849
rect -101 -1875 -51 -1849
rect -25 -1875 25 -1849
rect 51 -1875 101 -1849
rect 127 -1875 177 -1849
rect 203 -1875 253 -1849
rect 279 -1875 329 -1849
rect 355 -1875 405 -1849
rect 431 -1875 481 -1849
rect 507 -1875 513 -1849
rect -513 -1925 513 -1875
rect -513 -1951 -507 -1925
rect -481 -1951 -431 -1925
rect -405 -1951 -355 -1925
rect -329 -1951 -279 -1925
rect -253 -1951 -203 -1925
rect -177 -1951 -127 -1925
rect -101 -1951 -51 -1925
rect -25 -1951 25 -1925
rect 51 -1951 101 -1925
rect 127 -1951 177 -1925
rect 203 -1951 253 -1925
rect 279 -1951 329 -1925
rect 355 -1951 405 -1925
rect 431 -1951 481 -1925
rect 507 -1951 513 -1925
rect -513 -2001 513 -1951
rect -513 -2027 -507 -2001
rect -481 -2027 -431 -2001
rect -405 -2027 -355 -2001
rect -329 -2027 -279 -2001
rect -253 -2027 -203 -2001
rect -177 -2027 -127 -2001
rect -101 -2027 -51 -2001
rect -25 -2027 25 -2001
rect 51 -2027 101 -2001
rect 127 -2027 177 -2001
rect 203 -2027 253 -2001
rect 279 -2027 329 -2001
rect 355 -2027 405 -2001
rect 431 -2027 481 -2001
rect 507 -2027 513 -2001
rect -513 -2077 513 -2027
rect -513 -2103 -507 -2077
rect -481 -2103 -431 -2077
rect -405 -2103 -355 -2077
rect -329 -2103 -279 -2077
rect -253 -2103 -203 -2077
rect -177 -2103 -127 -2077
rect -101 -2103 -51 -2077
rect -25 -2103 25 -2077
rect 51 -2103 101 -2077
rect 127 -2103 177 -2077
rect 203 -2103 253 -2077
rect 279 -2103 329 -2077
rect 355 -2103 405 -2077
rect 431 -2103 481 -2077
rect 507 -2103 513 -2077
rect -513 -2153 513 -2103
rect -513 -2179 -507 -2153
rect -481 -2179 -431 -2153
rect -405 -2179 -355 -2153
rect -329 -2179 -279 -2153
rect -253 -2179 -203 -2153
rect -177 -2179 -127 -2153
rect -101 -2179 -51 -2153
rect -25 -2179 25 -2153
rect 51 -2179 101 -2153
rect 127 -2179 177 -2153
rect 203 -2179 253 -2153
rect 279 -2179 329 -2153
rect 355 -2179 405 -2153
rect 431 -2179 481 -2153
rect 507 -2179 513 -2153
rect -513 -2229 513 -2179
rect -513 -2255 -507 -2229
rect -481 -2255 -431 -2229
rect -405 -2255 -355 -2229
rect -329 -2255 -279 -2229
rect -253 -2255 -203 -2229
rect -177 -2255 -127 -2229
rect -101 -2255 -51 -2229
rect -25 -2255 25 -2229
rect 51 -2255 101 -2229
rect 127 -2255 177 -2229
rect 203 -2255 253 -2229
rect 279 -2255 329 -2229
rect 355 -2255 405 -2229
rect 431 -2255 481 -2229
rect 507 -2255 513 -2229
rect -513 -2305 513 -2255
rect -513 -2331 -507 -2305
rect -481 -2331 -431 -2305
rect -405 -2331 -355 -2305
rect -329 -2331 -279 -2305
rect -253 -2331 -203 -2305
rect -177 -2331 -127 -2305
rect -101 -2331 -51 -2305
rect -25 -2331 25 -2305
rect 51 -2331 101 -2305
rect 127 -2331 177 -2305
rect 203 -2331 253 -2305
rect 279 -2331 329 -2305
rect 355 -2331 405 -2305
rect 431 -2331 481 -2305
rect 507 -2331 513 -2305
rect -513 -2381 513 -2331
rect -513 -2407 -507 -2381
rect -481 -2407 -431 -2381
rect -405 -2407 -355 -2381
rect -329 -2407 -279 -2381
rect -253 -2407 -203 -2381
rect -177 -2407 -127 -2381
rect -101 -2407 -51 -2381
rect -25 -2407 25 -2381
rect 51 -2407 101 -2381
rect 127 -2407 177 -2381
rect 203 -2407 253 -2381
rect 279 -2407 329 -2381
rect 355 -2407 405 -2381
rect 431 -2407 481 -2381
rect 507 -2407 513 -2381
rect -513 -2457 513 -2407
rect -513 -2483 -507 -2457
rect -481 -2483 -431 -2457
rect -405 -2483 -355 -2457
rect -329 -2483 -279 -2457
rect -253 -2483 -203 -2457
rect -177 -2483 -127 -2457
rect -101 -2483 -51 -2457
rect -25 -2483 25 -2457
rect 51 -2483 101 -2457
rect 127 -2483 177 -2457
rect 203 -2483 253 -2457
rect 279 -2483 329 -2457
rect 355 -2483 405 -2457
rect 431 -2483 481 -2457
rect 507 -2483 513 -2457
rect -513 -2533 513 -2483
rect -513 -2559 -507 -2533
rect -481 -2559 -431 -2533
rect -405 -2559 -355 -2533
rect -329 -2559 -279 -2533
rect -253 -2559 -203 -2533
rect -177 -2559 -127 -2533
rect -101 -2559 -51 -2533
rect -25 -2559 25 -2533
rect 51 -2559 101 -2533
rect 127 -2559 177 -2533
rect 203 -2559 253 -2533
rect 279 -2559 329 -2533
rect 355 -2559 405 -2533
rect 431 -2559 481 -2533
rect 507 -2559 513 -2533
rect -513 -2609 513 -2559
rect -513 -2635 -507 -2609
rect -481 -2635 -431 -2609
rect -405 -2635 -355 -2609
rect -329 -2635 -279 -2609
rect -253 -2635 -203 -2609
rect -177 -2635 -127 -2609
rect -101 -2635 -51 -2609
rect -25 -2635 25 -2609
rect 51 -2635 101 -2609
rect 127 -2635 177 -2609
rect 203 -2635 253 -2609
rect 279 -2635 329 -2609
rect 355 -2635 405 -2609
rect 431 -2635 481 -2609
rect 507 -2635 513 -2609
rect -513 -2641 513 -2635
<< via1 >>
rect -507 2609 -481 2635
rect -431 2609 -405 2635
rect -355 2609 -329 2635
rect -279 2609 -253 2635
rect -203 2609 -177 2635
rect -127 2609 -101 2635
rect -51 2609 -25 2635
rect 25 2609 51 2635
rect 101 2609 127 2635
rect 177 2609 203 2635
rect 253 2609 279 2635
rect 329 2609 355 2635
rect 405 2609 431 2635
rect 481 2609 507 2635
rect -507 2533 -481 2559
rect -431 2533 -405 2559
rect -355 2533 -329 2559
rect -279 2533 -253 2559
rect -203 2533 -177 2559
rect -127 2533 -101 2559
rect -51 2533 -25 2559
rect 25 2533 51 2559
rect 101 2533 127 2559
rect 177 2533 203 2559
rect 253 2533 279 2559
rect 329 2533 355 2559
rect 405 2533 431 2559
rect 481 2533 507 2559
rect -507 2457 -481 2483
rect -431 2457 -405 2483
rect -355 2457 -329 2483
rect -279 2457 -253 2483
rect -203 2457 -177 2483
rect -127 2457 -101 2483
rect -51 2457 -25 2483
rect 25 2457 51 2483
rect 101 2457 127 2483
rect 177 2457 203 2483
rect 253 2457 279 2483
rect 329 2457 355 2483
rect 405 2457 431 2483
rect 481 2457 507 2483
rect -507 2381 -481 2407
rect -431 2381 -405 2407
rect -355 2381 -329 2407
rect -279 2381 -253 2407
rect -203 2381 -177 2407
rect -127 2381 -101 2407
rect -51 2381 -25 2407
rect 25 2381 51 2407
rect 101 2381 127 2407
rect 177 2381 203 2407
rect 253 2381 279 2407
rect 329 2381 355 2407
rect 405 2381 431 2407
rect 481 2381 507 2407
rect -507 2305 -481 2331
rect -431 2305 -405 2331
rect -355 2305 -329 2331
rect -279 2305 -253 2331
rect -203 2305 -177 2331
rect -127 2305 -101 2331
rect -51 2305 -25 2331
rect 25 2305 51 2331
rect 101 2305 127 2331
rect 177 2305 203 2331
rect 253 2305 279 2331
rect 329 2305 355 2331
rect 405 2305 431 2331
rect 481 2305 507 2331
rect -507 2229 -481 2255
rect -431 2229 -405 2255
rect -355 2229 -329 2255
rect -279 2229 -253 2255
rect -203 2229 -177 2255
rect -127 2229 -101 2255
rect -51 2229 -25 2255
rect 25 2229 51 2255
rect 101 2229 127 2255
rect 177 2229 203 2255
rect 253 2229 279 2255
rect 329 2229 355 2255
rect 405 2229 431 2255
rect 481 2229 507 2255
rect -507 2153 -481 2179
rect -431 2153 -405 2179
rect -355 2153 -329 2179
rect -279 2153 -253 2179
rect -203 2153 -177 2179
rect -127 2153 -101 2179
rect -51 2153 -25 2179
rect 25 2153 51 2179
rect 101 2153 127 2179
rect 177 2153 203 2179
rect 253 2153 279 2179
rect 329 2153 355 2179
rect 405 2153 431 2179
rect 481 2153 507 2179
rect -507 2077 -481 2103
rect -431 2077 -405 2103
rect -355 2077 -329 2103
rect -279 2077 -253 2103
rect -203 2077 -177 2103
rect -127 2077 -101 2103
rect -51 2077 -25 2103
rect 25 2077 51 2103
rect 101 2077 127 2103
rect 177 2077 203 2103
rect 253 2077 279 2103
rect 329 2077 355 2103
rect 405 2077 431 2103
rect 481 2077 507 2103
rect -507 2001 -481 2027
rect -431 2001 -405 2027
rect -355 2001 -329 2027
rect -279 2001 -253 2027
rect -203 2001 -177 2027
rect -127 2001 -101 2027
rect -51 2001 -25 2027
rect 25 2001 51 2027
rect 101 2001 127 2027
rect 177 2001 203 2027
rect 253 2001 279 2027
rect 329 2001 355 2027
rect 405 2001 431 2027
rect 481 2001 507 2027
rect -507 1925 -481 1951
rect -431 1925 -405 1951
rect -355 1925 -329 1951
rect -279 1925 -253 1951
rect -203 1925 -177 1951
rect -127 1925 -101 1951
rect -51 1925 -25 1951
rect 25 1925 51 1951
rect 101 1925 127 1951
rect 177 1925 203 1951
rect 253 1925 279 1951
rect 329 1925 355 1951
rect 405 1925 431 1951
rect 481 1925 507 1951
rect -507 1849 -481 1875
rect -431 1849 -405 1875
rect -355 1849 -329 1875
rect -279 1849 -253 1875
rect -203 1849 -177 1875
rect -127 1849 -101 1875
rect -51 1849 -25 1875
rect 25 1849 51 1875
rect 101 1849 127 1875
rect 177 1849 203 1875
rect 253 1849 279 1875
rect 329 1849 355 1875
rect 405 1849 431 1875
rect 481 1849 507 1875
rect -507 1773 -481 1799
rect -431 1773 -405 1799
rect -355 1773 -329 1799
rect -279 1773 -253 1799
rect -203 1773 -177 1799
rect -127 1773 -101 1799
rect -51 1773 -25 1799
rect 25 1773 51 1799
rect 101 1773 127 1799
rect 177 1773 203 1799
rect 253 1773 279 1799
rect 329 1773 355 1799
rect 405 1773 431 1799
rect 481 1773 507 1799
rect -507 1697 -481 1723
rect -431 1697 -405 1723
rect -355 1697 -329 1723
rect -279 1697 -253 1723
rect -203 1697 -177 1723
rect -127 1697 -101 1723
rect -51 1697 -25 1723
rect 25 1697 51 1723
rect 101 1697 127 1723
rect 177 1697 203 1723
rect 253 1697 279 1723
rect 329 1697 355 1723
rect 405 1697 431 1723
rect 481 1697 507 1723
rect -507 1621 -481 1647
rect -431 1621 -405 1647
rect -355 1621 -329 1647
rect -279 1621 -253 1647
rect -203 1621 -177 1647
rect -127 1621 -101 1647
rect -51 1621 -25 1647
rect 25 1621 51 1647
rect 101 1621 127 1647
rect 177 1621 203 1647
rect 253 1621 279 1647
rect 329 1621 355 1647
rect 405 1621 431 1647
rect 481 1621 507 1647
rect -507 1545 -481 1571
rect -431 1545 -405 1571
rect -355 1545 -329 1571
rect -279 1545 -253 1571
rect -203 1545 -177 1571
rect -127 1545 -101 1571
rect -51 1545 -25 1571
rect 25 1545 51 1571
rect 101 1545 127 1571
rect 177 1545 203 1571
rect 253 1545 279 1571
rect 329 1545 355 1571
rect 405 1545 431 1571
rect 481 1545 507 1571
rect -507 1469 -481 1495
rect -431 1469 -405 1495
rect -355 1469 -329 1495
rect -279 1469 -253 1495
rect -203 1469 -177 1495
rect -127 1469 -101 1495
rect -51 1469 -25 1495
rect 25 1469 51 1495
rect 101 1469 127 1495
rect 177 1469 203 1495
rect 253 1469 279 1495
rect 329 1469 355 1495
rect 405 1469 431 1495
rect 481 1469 507 1495
rect -507 1393 -481 1419
rect -431 1393 -405 1419
rect -355 1393 -329 1419
rect -279 1393 -253 1419
rect -203 1393 -177 1419
rect -127 1393 -101 1419
rect -51 1393 -25 1419
rect 25 1393 51 1419
rect 101 1393 127 1419
rect 177 1393 203 1419
rect 253 1393 279 1419
rect 329 1393 355 1419
rect 405 1393 431 1419
rect 481 1393 507 1419
rect -507 1317 -481 1343
rect -431 1317 -405 1343
rect -355 1317 -329 1343
rect -279 1317 -253 1343
rect -203 1317 -177 1343
rect -127 1317 -101 1343
rect -51 1317 -25 1343
rect 25 1317 51 1343
rect 101 1317 127 1343
rect 177 1317 203 1343
rect 253 1317 279 1343
rect 329 1317 355 1343
rect 405 1317 431 1343
rect 481 1317 507 1343
rect -507 1241 -481 1267
rect -431 1241 -405 1267
rect -355 1241 -329 1267
rect -279 1241 -253 1267
rect -203 1241 -177 1267
rect -127 1241 -101 1267
rect -51 1241 -25 1267
rect 25 1241 51 1267
rect 101 1241 127 1267
rect 177 1241 203 1267
rect 253 1241 279 1267
rect 329 1241 355 1267
rect 405 1241 431 1267
rect 481 1241 507 1267
rect -507 1165 -481 1191
rect -431 1165 -405 1191
rect -355 1165 -329 1191
rect -279 1165 -253 1191
rect -203 1165 -177 1191
rect -127 1165 -101 1191
rect -51 1165 -25 1191
rect 25 1165 51 1191
rect 101 1165 127 1191
rect 177 1165 203 1191
rect 253 1165 279 1191
rect 329 1165 355 1191
rect 405 1165 431 1191
rect 481 1165 507 1191
rect -507 1089 -481 1115
rect -431 1089 -405 1115
rect -355 1089 -329 1115
rect -279 1089 -253 1115
rect -203 1089 -177 1115
rect -127 1089 -101 1115
rect -51 1089 -25 1115
rect 25 1089 51 1115
rect 101 1089 127 1115
rect 177 1089 203 1115
rect 253 1089 279 1115
rect 329 1089 355 1115
rect 405 1089 431 1115
rect 481 1089 507 1115
rect -507 1013 -481 1039
rect -431 1013 -405 1039
rect -355 1013 -329 1039
rect -279 1013 -253 1039
rect -203 1013 -177 1039
rect -127 1013 -101 1039
rect -51 1013 -25 1039
rect 25 1013 51 1039
rect 101 1013 127 1039
rect 177 1013 203 1039
rect 253 1013 279 1039
rect 329 1013 355 1039
rect 405 1013 431 1039
rect 481 1013 507 1039
rect -507 937 -481 963
rect -431 937 -405 963
rect -355 937 -329 963
rect -279 937 -253 963
rect -203 937 -177 963
rect -127 937 -101 963
rect -51 937 -25 963
rect 25 937 51 963
rect 101 937 127 963
rect 177 937 203 963
rect 253 937 279 963
rect 329 937 355 963
rect 405 937 431 963
rect 481 937 507 963
rect -507 861 -481 887
rect -431 861 -405 887
rect -355 861 -329 887
rect -279 861 -253 887
rect -203 861 -177 887
rect -127 861 -101 887
rect -51 861 -25 887
rect 25 861 51 887
rect 101 861 127 887
rect 177 861 203 887
rect 253 861 279 887
rect 329 861 355 887
rect 405 861 431 887
rect 481 861 507 887
rect -507 785 -481 811
rect -431 785 -405 811
rect -355 785 -329 811
rect -279 785 -253 811
rect -203 785 -177 811
rect -127 785 -101 811
rect -51 785 -25 811
rect 25 785 51 811
rect 101 785 127 811
rect 177 785 203 811
rect 253 785 279 811
rect 329 785 355 811
rect 405 785 431 811
rect 481 785 507 811
rect -507 709 -481 735
rect -431 709 -405 735
rect -355 709 -329 735
rect -279 709 -253 735
rect -203 709 -177 735
rect -127 709 -101 735
rect -51 709 -25 735
rect 25 709 51 735
rect 101 709 127 735
rect 177 709 203 735
rect 253 709 279 735
rect 329 709 355 735
rect 405 709 431 735
rect 481 709 507 735
rect -507 633 -481 659
rect -431 633 -405 659
rect -355 633 -329 659
rect -279 633 -253 659
rect -203 633 -177 659
rect -127 633 -101 659
rect -51 633 -25 659
rect 25 633 51 659
rect 101 633 127 659
rect 177 633 203 659
rect 253 633 279 659
rect 329 633 355 659
rect 405 633 431 659
rect 481 633 507 659
rect -507 557 -481 583
rect -431 557 -405 583
rect -355 557 -329 583
rect -279 557 -253 583
rect -203 557 -177 583
rect -127 557 -101 583
rect -51 557 -25 583
rect 25 557 51 583
rect 101 557 127 583
rect 177 557 203 583
rect 253 557 279 583
rect 329 557 355 583
rect 405 557 431 583
rect 481 557 507 583
rect -507 481 -481 507
rect -431 481 -405 507
rect -355 481 -329 507
rect -279 481 -253 507
rect -203 481 -177 507
rect -127 481 -101 507
rect -51 481 -25 507
rect 25 481 51 507
rect 101 481 127 507
rect 177 481 203 507
rect 253 481 279 507
rect 329 481 355 507
rect 405 481 431 507
rect 481 481 507 507
rect -507 405 -481 431
rect -431 405 -405 431
rect -355 405 -329 431
rect -279 405 -253 431
rect -203 405 -177 431
rect -127 405 -101 431
rect -51 405 -25 431
rect 25 405 51 431
rect 101 405 127 431
rect 177 405 203 431
rect 253 405 279 431
rect 329 405 355 431
rect 405 405 431 431
rect 481 405 507 431
rect -507 329 -481 355
rect -431 329 -405 355
rect -355 329 -329 355
rect -279 329 -253 355
rect -203 329 -177 355
rect -127 329 -101 355
rect -51 329 -25 355
rect 25 329 51 355
rect 101 329 127 355
rect 177 329 203 355
rect 253 329 279 355
rect 329 329 355 355
rect 405 329 431 355
rect 481 329 507 355
rect -507 253 -481 279
rect -431 253 -405 279
rect -355 253 -329 279
rect -279 253 -253 279
rect -203 253 -177 279
rect -127 253 -101 279
rect -51 253 -25 279
rect 25 253 51 279
rect 101 253 127 279
rect 177 253 203 279
rect 253 253 279 279
rect 329 253 355 279
rect 405 253 431 279
rect 481 253 507 279
rect -507 177 -481 203
rect -431 177 -405 203
rect -355 177 -329 203
rect -279 177 -253 203
rect -203 177 -177 203
rect -127 177 -101 203
rect -51 177 -25 203
rect 25 177 51 203
rect 101 177 127 203
rect 177 177 203 203
rect 253 177 279 203
rect 329 177 355 203
rect 405 177 431 203
rect 481 177 507 203
rect -507 101 -481 127
rect -431 101 -405 127
rect -355 101 -329 127
rect -279 101 -253 127
rect -203 101 -177 127
rect -127 101 -101 127
rect -51 101 -25 127
rect 25 101 51 127
rect 101 101 127 127
rect 177 101 203 127
rect 253 101 279 127
rect 329 101 355 127
rect 405 101 431 127
rect 481 101 507 127
rect -507 25 -481 51
rect -431 25 -405 51
rect -355 25 -329 51
rect -279 25 -253 51
rect -203 25 -177 51
rect -127 25 -101 51
rect -51 25 -25 51
rect 25 25 51 51
rect 101 25 127 51
rect 177 25 203 51
rect 253 25 279 51
rect 329 25 355 51
rect 405 25 431 51
rect 481 25 507 51
rect -507 -51 -481 -25
rect -431 -51 -405 -25
rect -355 -51 -329 -25
rect -279 -51 -253 -25
rect -203 -51 -177 -25
rect -127 -51 -101 -25
rect -51 -51 -25 -25
rect 25 -51 51 -25
rect 101 -51 127 -25
rect 177 -51 203 -25
rect 253 -51 279 -25
rect 329 -51 355 -25
rect 405 -51 431 -25
rect 481 -51 507 -25
rect -507 -127 -481 -101
rect -431 -127 -405 -101
rect -355 -127 -329 -101
rect -279 -127 -253 -101
rect -203 -127 -177 -101
rect -127 -127 -101 -101
rect -51 -127 -25 -101
rect 25 -127 51 -101
rect 101 -127 127 -101
rect 177 -127 203 -101
rect 253 -127 279 -101
rect 329 -127 355 -101
rect 405 -127 431 -101
rect 481 -127 507 -101
rect -507 -203 -481 -177
rect -431 -203 -405 -177
rect -355 -203 -329 -177
rect -279 -203 -253 -177
rect -203 -203 -177 -177
rect -127 -203 -101 -177
rect -51 -203 -25 -177
rect 25 -203 51 -177
rect 101 -203 127 -177
rect 177 -203 203 -177
rect 253 -203 279 -177
rect 329 -203 355 -177
rect 405 -203 431 -177
rect 481 -203 507 -177
rect -507 -279 -481 -253
rect -431 -279 -405 -253
rect -355 -279 -329 -253
rect -279 -279 -253 -253
rect -203 -279 -177 -253
rect -127 -279 -101 -253
rect -51 -279 -25 -253
rect 25 -279 51 -253
rect 101 -279 127 -253
rect 177 -279 203 -253
rect 253 -279 279 -253
rect 329 -279 355 -253
rect 405 -279 431 -253
rect 481 -279 507 -253
rect -507 -355 -481 -329
rect -431 -355 -405 -329
rect -355 -355 -329 -329
rect -279 -355 -253 -329
rect -203 -355 -177 -329
rect -127 -355 -101 -329
rect -51 -355 -25 -329
rect 25 -355 51 -329
rect 101 -355 127 -329
rect 177 -355 203 -329
rect 253 -355 279 -329
rect 329 -355 355 -329
rect 405 -355 431 -329
rect 481 -355 507 -329
rect -507 -431 -481 -405
rect -431 -431 -405 -405
rect -355 -431 -329 -405
rect -279 -431 -253 -405
rect -203 -431 -177 -405
rect -127 -431 -101 -405
rect -51 -431 -25 -405
rect 25 -431 51 -405
rect 101 -431 127 -405
rect 177 -431 203 -405
rect 253 -431 279 -405
rect 329 -431 355 -405
rect 405 -431 431 -405
rect 481 -431 507 -405
rect -507 -507 -481 -481
rect -431 -507 -405 -481
rect -355 -507 -329 -481
rect -279 -507 -253 -481
rect -203 -507 -177 -481
rect -127 -507 -101 -481
rect -51 -507 -25 -481
rect 25 -507 51 -481
rect 101 -507 127 -481
rect 177 -507 203 -481
rect 253 -507 279 -481
rect 329 -507 355 -481
rect 405 -507 431 -481
rect 481 -507 507 -481
rect -507 -583 -481 -557
rect -431 -583 -405 -557
rect -355 -583 -329 -557
rect -279 -583 -253 -557
rect -203 -583 -177 -557
rect -127 -583 -101 -557
rect -51 -583 -25 -557
rect 25 -583 51 -557
rect 101 -583 127 -557
rect 177 -583 203 -557
rect 253 -583 279 -557
rect 329 -583 355 -557
rect 405 -583 431 -557
rect 481 -583 507 -557
rect -507 -659 -481 -633
rect -431 -659 -405 -633
rect -355 -659 -329 -633
rect -279 -659 -253 -633
rect -203 -659 -177 -633
rect -127 -659 -101 -633
rect -51 -659 -25 -633
rect 25 -659 51 -633
rect 101 -659 127 -633
rect 177 -659 203 -633
rect 253 -659 279 -633
rect 329 -659 355 -633
rect 405 -659 431 -633
rect 481 -659 507 -633
rect -507 -735 -481 -709
rect -431 -735 -405 -709
rect -355 -735 -329 -709
rect -279 -735 -253 -709
rect -203 -735 -177 -709
rect -127 -735 -101 -709
rect -51 -735 -25 -709
rect 25 -735 51 -709
rect 101 -735 127 -709
rect 177 -735 203 -709
rect 253 -735 279 -709
rect 329 -735 355 -709
rect 405 -735 431 -709
rect 481 -735 507 -709
rect -507 -811 -481 -785
rect -431 -811 -405 -785
rect -355 -811 -329 -785
rect -279 -811 -253 -785
rect -203 -811 -177 -785
rect -127 -811 -101 -785
rect -51 -811 -25 -785
rect 25 -811 51 -785
rect 101 -811 127 -785
rect 177 -811 203 -785
rect 253 -811 279 -785
rect 329 -811 355 -785
rect 405 -811 431 -785
rect 481 -811 507 -785
rect -507 -887 -481 -861
rect -431 -887 -405 -861
rect -355 -887 -329 -861
rect -279 -887 -253 -861
rect -203 -887 -177 -861
rect -127 -887 -101 -861
rect -51 -887 -25 -861
rect 25 -887 51 -861
rect 101 -887 127 -861
rect 177 -887 203 -861
rect 253 -887 279 -861
rect 329 -887 355 -861
rect 405 -887 431 -861
rect 481 -887 507 -861
rect -507 -963 -481 -937
rect -431 -963 -405 -937
rect -355 -963 -329 -937
rect -279 -963 -253 -937
rect -203 -963 -177 -937
rect -127 -963 -101 -937
rect -51 -963 -25 -937
rect 25 -963 51 -937
rect 101 -963 127 -937
rect 177 -963 203 -937
rect 253 -963 279 -937
rect 329 -963 355 -937
rect 405 -963 431 -937
rect 481 -963 507 -937
rect -507 -1039 -481 -1013
rect -431 -1039 -405 -1013
rect -355 -1039 -329 -1013
rect -279 -1039 -253 -1013
rect -203 -1039 -177 -1013
rect -127 -1039 -101 -1013
rect -51 -1039 -25 -1013
rect 25 -1039 51 -1013
rect 101 -1039 127 -1013
rect 177 -1039 203 -1013
rect 253 -1039 279 -1013
rect 329 -1039 355 -1013
rect 405 -1039 431 -1013
rect 481 -1039 507 -1013
rect -507 -1115 -481 -1089
rect -431 -1115 -405 -1089
rect -355 -1115 -329 -1089
rect -279 -1115 -253 -1089
rect -203 -1115 -177 -1089
rect -127 -1115 -101 -1089
rect -51 -1115 -25 -1089
rect 25 -1115 51 -1089
rect 101 -1115 127 -1089
rect 177 -1115 203 -1089
rect 253 -1115 279 -1089
rect 329 -1115 355 -1089
rect 405 -1115 431 -1089
rect 481 -1115 507 -1089
rect -507 -1191 -481 -1165
rect -431 -1191 -405 -1165
rect -355 -1191 -329 -1165
rect -279 -1191 -253 -1165
rect -203 -1191 -177 -1165
rect -127 -1191 -101 -1165
rect -51 -1191 -25 -1165
rect 25 -1191 51 -1165
rect 101 -1191 127 -1165
rect 177 -1191 203 -1165
rect 253 -1191 279 -1165
rect 329 -1191 355 -1165
rect 405 -1191 431 -1165
rect 481 -1191 507 -1165
rect -507 -1267 -481 -1241
rect -431 -1267 -405 -1241
rect -355 -1267 -329 -1241
rect -279 -1267 -253 -1241
rect -203 -1267 -177 -1241
rect -127 -1267 -101 -1241
rect -51 -1267 -25 -1241
rect 25 -1267 51 -1241
rect 101 -1267 127 -1241
rect 177 -1267 203 -1241
rect 253 -1267 279 -1241
rect 329 -1267 355 -1241
rect 405 -1267 431 -1241
rect 481 -1267 507 -1241
rect -507 -1343 -481 -1317
rect -431 -1343 -405 -1317
rect -355 -1343 -329 -1317
rect -279 -1343 -253 -1317
rect -203 -1343 -177 -1317
rect -127 -1343 -101 -1317
rect -51 -1343 -25 -1317
rect 25 -1343 51 -1317
rect 101 -1343 127 -1317
rect 177 -1343 203 -1317
rect 253 -1343 279 -1317
rect 329 -1343 355 -1317
rect 405 -1343 431 -1317
rect 481 -1343 507 -1317
rect -507 -1419 -481 -1393
rect -431 -1419 -405 -1393
rect -355 -1419 -329 -1393
rect -279 -1419 -253 -1393
rect -203 -1419 -177 -1393
rect -127 -1419 -101 -1393
rect -51 -1419 -25 -1393
rect 25 -1419 51 -1393
rect 101 -1419 127 -1393
rect 177 -1419 203 -1393
rect 253 -1419 279 -1393
rect 329 -1419 355 -1393
rect 405 -1419 431 -1393
rect 481 -1419 507 -1393
rect -507 -1495 -481 -1469
rect -431 -1495 -405 -1469
rect -355 -1495 -329 -1469
rect -279 -1495 -253 -1469
rect -203 -1495 -177 -1469
rect -127 -1495 -101 -1469
rect -51 -1495 -25 -1469
rect 25 -1495 51 -1469
rect 101 -1495 127 -1469
rect 177 -1495 203 -1469
rect 253 -1495 279 -1469
rect 329 -1495 355 -1469
rect 405 -1495 431 -1469
rect 481 -1495 507 -1469
rect -507 -1571 -481 -1545
rect -431 -1571 -405 -1545
rect -355 -1571 -329 -1545
rect -279 -1571 -253 -1545
rect -203 -1571 -177 -1545
rect -127 -1571 -101 -1545
rect -51 -1571 -25 -1545
rect 25 -1571 51 -1545
rect 101 -1571 127 -1545
rect 177 -1571 203 -1545
rect 253 -1571 279 -1545
rect 329 -1571 355 -1545
rect 405 -1571 431 -1545
rect 481 -1571 507 -1545
rect -507 -1647 -481 -1621
rect -431 -1647 -405 -1621
rect -355 -1647 -329 -1621
rect -279 -1647 -253 -1621
rect -203 -1647 -177 -1621
rect -127 -1647 -101 -1621
rect -51 -1647 -25 -1621
rect 25 -1647 51 -1621
rect 101 -1647 127 -1621
rect 177 -1647 203 -1621
rect 253 -1647 279 -1621
rect 329 -1647 355 -1621
rect 405 -1647 431 -1621
rect 481 -1647 507 -1621
rect -507 -1723 -481 -1697
rect -431 -1723 -405 -1697
rect -355 -1723 -329 -1697
rect -279 -1723 -253 -1697
rect -203 -1723 -177 -1697
rect -127 -1723 -101 -1697
rect -51 -1723 -25 -1697
rect 25 -1723 51 -1697
rect 101 -1723 127 -1697
rect 177 -1723 203 -1697
rect 253 -1723 279 -1697
rect 329 -1723 355 -1697
rect 405 -1723 431 -1697
rect 481 -1723 507 -1697
rect -507 -1799 -481 -1773
rect -431 -1799 -405 -1773
rect -355 -1799 -329 -1773
rect -279 -1799 -253 -1773
rect -203 -1799 -177 -1773
rect -127 -1799 -101 -1773
rect -51 -1799 -25 -1773
rect 25 -1799 51 -1773
rect 101 -1799 127 -1773
rect 177 -1799 203 -1773
rect 253 -1799 279 -1773
rect 329 -1799 355 -1773
rect 405 -1799 431 -1773
rect 481 -1799 507 -1773
rect -507 -1875 -481 -1849
rect -431 -1875 -405 -1849
rect -355 -1875 -329 -1849
rect -279 -1875 -253 -1849
rect -203 -1875 -177 -1849
rect -127 -1875 -101 -1849
rect -51 -1875 -25 -1849
rect 25 -1875 51 -1849
rect 101 -1875 127 -1849
rect 177 -1875 203 -1849
rect 253 -1875 279 -1849
rect 329 -1875 355 -1849
rect 405 -1875 431 -1849
rect 481 -1875 507 -1849
rect -507 -1951 -481 -1925
rect -431 -1951 -405 -1925
rect -355 -1951 -329 -1925
rect -279 -1951 -253 -1925
rect -203 -1951 -177 -1925
rect -127 -1951 -101 -1925
rect -51 -1951 -25 -1925
rect 25 -1951 51 -1925
rect 101 -1951 127 -1925
rect 177 -1951 203 -1925
rect 253 -1951 279 -1925
rect 329 -1951 355 -1925
rect 405 -1951 431 -1925
rect 481 -1951 507 -1925
rect -507 -2027 -481 -2001
rect -431 -2027 -405 -2001
rect -355 -2027 -329 -2001
rect -279 -2027 -253 -2001
rect -203 -2027 -177 -2001
rect -127 -2027 -101 -2001
rect -51 -2027 -25 -2001
rect 25 -2027 51 -2001
rect 101 -2027 127 -2001
rect 177 -2027 203 -2001
rect 253 -2027 279 -2001
rect 329 -2027 355 -2001
rect 405 -2027 431 -2001
rect 481 -2027 507 -2001
rect -507 -2103 -481 -2077
rect -431 -2103 -405 -2077
rect -355 -2103 -329 -2077
rect -279 -2103 -253 -2077
rect -203 -2103 -177 -2077
rect -127 -2103 -101 -2077
rect -51 -2103 -25 -2077
rect 25 -2103 51 -2077
rect 101 -2103 127 -2077
rect 177 -2103 203 -2077
rect 253 -2103 279 -2077
rect 329 -2103 355 -2077
rect 405 -2103 431 -2077
rect 481 -2103 507 -2077
rect -507 -2179 -481 -2153
rect -431 -2179 -405 -2153
rect -355 -2179 -329 -2153
rect -279 -2179 -253 -2153
rect -203 -2179 -177 -2153
rect -127 -2179 -101 -2153
rect -51 -2179 -25 -2153
rect 25 -2179 51 -2153
rect 101 -2179 127 -2153
rect 177 -2179 203 -2153
rect 253 -2179 279 -2153
rect 329 -2179 355 -2153
rect 405 -2179 431 -2153
rect 481 -2179 507 -2153
rect -507 -2255 -481 -2229
rect -431 -2255 -405 -2229
rect -355 -2255 -329 -2229
rect -279 -2255 -253 -2229
rect -203 -2255 -177 -2229
rect -127 -2255 -101 -2229
rect -51 -2255 -25 -2229
rect 25 -2255 51 -2229
rect 101 -2255 127 -2229
rect 177 -2255 203 -2229
rect 253 -2255 279 -2229
rect 329 -2255 355 -2229
rect 405 -2255 431 -2229
rect 481 -2255 507 -2229
rect -507 -2331 -481 -2305
rect -431 -2331 -405 -2305
rect -355 -2331 -329 -2305
rect -279 -2331 -253 -2305
rect -203 -2331 -177 -2305
rect -127 -2331 -101 -2305
rect -51 -2331 -25 -2305
rect 25 -2331 51 -2305
rect 101 -2331 127 -2305
rect 177 -2331 203 -2305
rect 253 -2331 279 -2305
rect 329 -2331 355 -2305
rect 405 -2331 431 -2305
rect 481 -2331 507 -2305
rect -507 -2407 -481 -2381
rect -431 -2407 -405 -2381
rect -355 -2407 -329 -2381
rect -279 -2407 -253 -2381
rect -203 -2407 -177 -2381
rect -127 -2407 -101 -2381
rect -51 -2407 -25 -2381
rect 25 -2407 51 -2381
rect 101 -2407 127 -2381
rect 177 -2407 203 -2381
rect 253 -2407 279 -2381
rect 329 -2407 355 -2381
rect 405 -2407 431 -2381
rect 481 -2407 507 -2381
rect -507 -2483 -481 -2457
rect -431 -2483 -405 -2457
rect -355 -2483 -329 -2457
rect -279 -2483 -253 -2457
rect -203 -2483 -177 -2457
rect -127 -2483 -101 -2457
rect -51 -2483 -25 -2457
rect 25 -2483 51 -2457
rect 101 -2483 127 -2457
rect 177 -2483 203 -2457
rect 253 -2483 279 -2457
rect 329 -2483 355 -2457
rect 405 -2483 431 -2457
rect 481 -2483 507 -2457
rect -507 -2559 -481 -2533
rect -431 -2559 -405 -2533
rect -355 -2559 -329 -2533
rect -279 -2559 -253 -2533
rect -203 -2559 -177 -2533
rect -127 -2559 -101 -2533
rect -51 -2559 -25 -2533
rect 25 -2559 51 -2533
rect 101 -2559 127 -2533
rect 177 -2559 203 -2533
rect 253 -2559 279 -2533
rect 329 -2559 355 -2533
rect 405 -2559 431 -2533
rect 481 -2559 507 -2533
rect -507 -2635 -481 -2609
rect -431 -2635 -405 -2609
rect -355 -2635 -329 -2609
rect -279 -2635 -253 -2609
rect -203 -2635 -177 -2609
rect -127 -2635 -101 -2609
rect -51 -2635 -25 -2609
rect 25 -2635 51 -2609
rect 101 -2635 127 -2609
rect 177 -2635 203 -2609
rect 253 -2635 279 -2609
rect 329 -2635 355 -2609
rect 405 -2635 431 -2609
rect 481 -2635 507 -2609
<< metal2 >>
rect -513 2635 513 2641
rect -513 2609 -507 2635
rect -481 2609 -431 2635
rect -405 2609 -355 2635
rect -329 2609 -279 2635
rect -253 2609 -203 2635
rect -177 2609 -127 2635
rect -101 2609 -51 2635
rect -25 2609 25 2635
rect 51 2609 101 2635
rect 127 2609 177 2635
rect 203 2609 253 2635
rect 279 2609 329 2635
rect 355 2609 405 2635
rect 431 2609 481 2635
rect 507 2609 513 2635
rect -513 2559 513 2609
rect -513 2533 -507 2559
rect -481 2533 -431 2559
rect -405 2533 -355 2559
rect -329 2533 -279 2559
rect -253 2533 -203 2559
rect -177 2533 -127 2559
rect -101 2533 -51 2559
rect -25 2533 25 2559
rect 51 2533 101 2559
rect 127 2533 177 2559
rect 203 2533 253 2559
rect 279 2533 329 2559
rect 355 2533 405 2559
rect 431 2533 481 2559
rect 507 2533 513 2559
rect -513 2483 513 2533
rect -513 2457 -507 2483
rect -481 2457 -431 2483
rect -405 2457 -355 2483
rect -329 2457 -279 2483
rect -253 2457 -203 2483
rect -177 2457 -127 2483
rect -101 2457 -51 2483
rect -25 2457 25 2483
rect 51 2457 101 2483
rect 127 2457 177 2483
rect 203 2457 253 2483
rect 279 2457 329 2483
rect 355 2457 405 2483
rect 431 2457 481 2483
rect 507 2457 513 2483
rect -513 2407 513 2457
rect -513 2381 -507 2407
rect -481 2381 -431 2407
rect -405 2381 -355 2407
rect -329 2381 -279 2407
rect -253 2381 -203 2407
rect -177 2381 -127 2407
rect -101 2381 -51 2407
rect -25 2381 25 2407
rect 51 2381 101 2407
rect 127 2381 177 2407
rect 203 2381 253 2407
rect 279 2381 329 2407
rect 355 2381 405 2407
rect 431 2381 481 2407
rect 507 2381 513 2407
rect -513 2331 513 2381
rect -513 2305 -507 2331
rect -481 2305 -431 2331
rect -405 2305 -355 2331
rect -329 2305 -279 2331
rect -253 2305 -203 2331
rect -177 2305 -127 2331
rect -101 2305 -51 2331
rect -25 2305 25 2331
rect 51 2305 101 2331
rect 127 2305 177 2331
rect 203 2305 253 2331
rect 279 2305 329 2331
rect 355 2305 405 2331
rect 431 2305 481 2331
rect 507 2305 513 2331
rect -513 2255 513 2305
rect -513 2229 -507 2255
rect -481 2229 -431 2255
rect -405 2229 -355 2255
rect -329 2229 -279 2255
rect -253 2229 -203 2255
rect -177 2229 -127 2255
rect -101 2229 -51 2255
rect -25 2229 25 2255
rect 51 2229 101 2255
rect 127 2229 177 2255
rect 203 2229 253 2255
rect 279 2229 329 2255
rect 355 2229 405 2255
rect 431 2229 481 2255
rect 507 2229 513 2255
rect -513 2179 513 2229
rect -513 2153 -507 2179
rect -481 2153 -431 2179
rect -405 2153 -355 2179
rect -329 2153 -279 2179
rect -253 2153 -203 2179
rect -177 2153 -127 2179
rect -101 2153 -51 2179
rect -25 2153 25 2179
rect 51 2153 101 2179
rect 127 2153 177 2179
rect 203 2153 253 2179
rect 279 2153 329 2179
rect 355 2153 405 2179
rect 431 2153 481 2179
rect 507 2153 513 2179
rect -513 2103 513 2153
rect -513 2077 -507 2103
rect -481 2077 -431 2103
rect -405 2077 -355 2103
rect -329 2077 -279 2103
rect -253 2077 -203 2103
rect -177 2077 -127 2103
rect -101 2077 -51 2103
rect -25 2077 25 2103
rect 51 2077 101 2103
rect 127 2077 177 2103
rect 203 2077 253 2103
rect 279 2077 329 2103
rect 355 2077 405 2103
rect 431 2077 481 2103
rect 507 2077 513 2103
rect -513 2027 513 2077
rect -513 2001 -507 2027
rect -481 2001 -431 2027
rect -405 2001 -355 2027
rect -329 2001 -279 2027
rect -253 2001 -203 2027
rect -177 2001 -127 2027
rect -101 2001 -51 2027
rect -25 2001 25 2027
rect 51 2001 101 2027
rect 127 2001 177 2027
rect 203 2001 253 2027
rect 279 2001 329 2027
rect 355 2001 405 2027
rect 431 2001 481 2027
rect 507 2001 513 2027
rect -513 1951 513 2001
rect -513 1925 -507 1951
rect -481 1925 -431 1951
rect -405 1925 -355 1951
rect -329 1925 -279 1951
rect -253 1925 -203 1951
rect -177 1925 -127 1951
rect -101 1925 -51 1951
rect -25 1925 25 1951
rect 51 1925 101 1951
rect 127 1925 177 1951
rect 203 1925 253 1951
rect 279 1925 329 1951
rect 355 1925 405 1951
rect 431 1925 481 1951
rect 507 1925 513 1951
rect -513 1875 513 1925
rect -513 1849 -507 1875
rect -481 1849 -431 1875
rect -405 1849 -355 1875
rect -329 1849 -279 1875
rect -253 1849 -203 1875
rect -177 1849 -127 1875
rect -101 1849 -51 1875
rect -25 1849 25 1875
rect 51 1849 101 1875
rect 127 1849 177 1875
rect 203 1849 253 1875
rect 279 1849 329 1875
rect 355 1849 405 1875
rect 431 1849 481 1875
rect 507 1849 513 1875
rect -513 1799 513 1849
rect -513 1773 -507 1799
rect -481 1773 -431 1799
rect -405 1773 -355 1799
rect -329 1773 -279 1799
rect -253 1773 -203 1799
rect -177 1773 -127 1799
rect -101 1773 -51 1799
rect -25 1773 25 1799
rect 51 1773 101 1799
rect 127 1773 177 1799
rect 203 1773 253 1799
rect 279 1773 329 1799
rect 355 1773 405 1799
rect 431 1773 481 1799
rect 507 1773 513 1799
rect -513 1723 513 1773
rect -513 1697 -507 1723
rect -481 1697 -431 1723
rect -405 1697 -355 1723
rect -329 1697 -279 1723
rect -253 1697 -203 1723
rect -177 1697 -127 1723
rect -101 1697 -51 1723
rect -25 1697 25 1723
rect 51 1697 101 1723
rect 127 1697 177 1723
rect 203 1697 253 1723
rect 279 1697 329 1723
rect 355 1697 405 1723
rect 431 1697 481 1723
rect 507 1697 513 1723
rect -513 1647 513 1697
rect -513 1621 -507 1647
rect -481 1621 -431 1647
rect -405 1621 -355 1647
rect -329 1621 -279 1647
rect -253 1621 -203 1647
rect -177 1621 -127 1647
rect -101 1621 -51 1647
rect -25 1621 25 1647
rect 51 1621 101 1647
rect 127 1621 177 1647
rect 203 1621 253 1647
rect 279 1621 329 1647
rect 355 1621 405 1647
rect 431 1621 481 1647
rect 507 1621 513 1647
rect -513 1571 513 1621
rect -513 1545 -507 1571
rect -481 1545 -431 1571
rect -405 1545 -355 1571
rect -329 1545 -279 1571
rect -253 1545 -203 1571
rect -177 1545 -127 1571
rect -101 1545 -51 1571
rect -25 1545 25 1571
rect 51 1545 101 1571
rect 127 1545 177 1571
rect 203 1545 253 1571
rect 279 1545 329 1571
rect 355 1545 405 1571
rect 431 1545 481 1571
rect 507 1545 513 1571
rect -513 1495 513 1545
rect -513 1469 -507 1495
rect -481 1469 -431 1495
rect -405 1469 -355 1495
rect -329 1469 -279 1495
rect -253 1469 -203 1495
rect -177 1469 -127 1495
rect -101 1469 -51 1495
rect -25 1469 25 1495
rect 51 1469 101 1495
rect 127 1469 177 1495
rect 203 1469 253 1495
rect 279 1469 329 1495
rect 355 1469 405 1495
rect 431 1469 481 1495
rect 507 1469 513 1495
rect -513 1419 513 1469
rect -513 1393 -507 1419
rect -481 1393 -431 1419
rect -405 1393 -355 1419
rect -329 1393 -279 1419
rect -253 1393 -203 1419
rect -177 1393 -127 1419
rect -101 1393 -51 1419
rect -25 1393 25 1419
rect 51 1393 101 1419
rect 127 1393 177 1419
rect 203 1393 253 1419
rect 279 1393 329 1419
rect 355 1393 405 1419
rect 431 1393 481 1419
rect 507 1393 513 1419
rect -513 1343 513 1393
rect -513 1317 -507 1343
rect -481 1317 -431 1343
rect -405 1317 -355 1343
rect -329 1317 -279 1343
rect -253 1317 -203 1343
rect -177 1317 -127 1343
rect -101 1317 -51 1343
rect -25 1317 25 1343
rect 51 1317 101 1343
rect 127 1317 177 1343
rect 203 1317 253 1343
rect 279 1317 329 1343
rect 355 1317 405 1343
rect 431 1317 481 1343
rect 507 1317 513 1343
rect -513 1267 513 1317
rect -513 1241 -507 1267
rect -481 1241 -431 1267
rect -405 1241 -355 1267
rect -329 1241 -279 1267
rect -253 1241 -203 1267
rect -177 1241 -127 1267
rect -101 1241 -51 1267
rect -25 1241 25 1267
rect 51 1241 101 1267
rect 127 1241 177 1267
rect 203 1241 253 1267
rect 279 1241 329 1267
rect 355 1241 405 1267
rect 431 1241 481 1267
rect 507 1241 513 1267
rect -513 1191 513 1241
rect -513 1165 -507 1191
rect -481 1165 -431 1191
rect -405 1165 -355 1191
rect -329 1165 -279 1191
rect -253 1165 -203 1191
rect -177 1165 -127 1191
rect -101 1165 -51 1191
rect -25 1165 25 1191
rect 51 1165 101 1191
rect 127 1165 177 1191
rect 203 1165 253 1191
rect 279 1165 329 1191
rect 355 1165 405 1191
rect 431 1165 481 1191
rect 507 1165 513 1191
rect -513 1115 513 1165
rect -513 1089 -507 1115
rect -481 1089 -431 1115
rect -405 1089 -355 1115
rect -329 1089 -279 1115
rect -253 1089 -203 1115
rect -177 1089 -127 1115
rect -101 1089 -51 1115
rect -25 1089 25 1115
rect 51 1089 101 1115
rect 127 1089 177 1115
rect 203 1089 253 1115
rect 279 1089 329 1115
rect 355 1089 405 1115
rect 431 1089 481 1115
rect 507 1089 513 1115
rect -513 1039 513 1089
rect -513 1013 -507 1039
rect -481 1013 -431 1039
rect -405 1013 -355 1039
rect -329 1013 -279 1039
rect -253 1013 -203 1039
rect -177 1013 -127 1039
rect -101 1013 -51 1039
rect -25 1013 25 1039
rect 51 1013 101 1039
rect 127 1013 177 1039
rect 203 1013 253 1039
rect 279 1013 329 1039
rect 355 1013 405 1039
rect 431 1013 481 1039
rect 507 1013 513 1039
rect -513 963 513 1013
rect -513 937 -507 963
rect -481 937 -431 963
rect -405 937 -355 963
rect -329 937 -279 963
rect -253 937 -203 963
rect -177 937 -127 963
rect -101 937 -51 963
rect -25 937 25 963
rect 51 937 101 963
rect 127 937 177 963
rect 203 937 253 963
rect 279 937 329 963
rect 355 937 405 963
rect 431 937 481 963
rect 507 937 513 963
rect -513 887 513 937
rect -513 861 -507 887
rect -481 861 -431 887
rect -405 861 -355 887
rect -329 861 -279 887
rect -253 861 -203 887
rect -177 861 -127 887
rect -101 861 -51 887
rect -25 861 25 887
rect 51 861 101 887
rect 127 861 177 887
rect 203 861 253 887
rect 279 861 329 887
rect 355 861 405 887
rect 431 861 481 887
rect 507 861 513 887
rect -513 811 513 861
rect -513 785 -507 811
rect -481 785 -431 811
rect -405 785 -355 811
rect -329 785 -279 811
rect -253 785 -203 811
rect -177 785 -127 811
rect -101 785 -51 811
rect -25 785 25 811
rect 51 785 101 811
rect 127 785 177 811
rect 203 785 253 811
rect 279 785 329 811
rect 355 785 405 811
rect 431 785 481 811
rect 507 785 513 811
rect -513 735 513 785
rect -513 709 -507 735
rect -481 709 -431 735
rect -405 709 -355 735
rect -329 709 -279 735
rect -253 709 -203 735
rect -177 709 -127 735
rect -101 709 -51 735
rect -25 709 25 735
rect 51 709 101 735
rect 127 709 177 735
rect 203 709 253 735
rect 279 709 329 735
rect 355 709 405 735
rect 431 709 481 735
rect 507 709 513 735
rect -513 659 513 709
rect -513 633 -507 659
rect -481 633 -431 659
rect -405 633 -355 659
rect -329 633 -279 659
rect -253 633 -203 659
rect -177 633 -127 659
rect -101 633 -51 659
rect -25 633 25 659
rect 51 633 101 659
rect 127 633 177 659
rect 203 633 253 659
rect 279 633 329 659
rect 355 633 405 659
rect 431 633 481 659
rect 507 633 513 659
rect -513 583 513 633
rect -513 557 -507 583
rect -481 557 -431 583
rect -405 557 -355 583
rect -329 557 -279 583
rect -253 557 -203 583
rect -177 557 -127 583
rect -101 557 -51 583
rect -25 557 25 583
rect 51 557 101 583
rect 127 557 177 583
rect 203 557 253 583
rect 279 557 329 583
rect 355 557 405 583
rect 431 557 481 583
rect 507 557 513 583
rect -513 507 513 557
rect -513 481 -507 507
rect -481 481 -431 507
rect -405 481 -355 507
rect -329 481 -279 507
rect -253 481 -203 507
rect -177 481 -127 507
rect -101 481 -51 507
rect -25 481 25 507
rect 51 481 101 507
rect 127 481 177 507
rect 203 481 253 507
rect 279 481 329 507
rect 355 481 405 507
rect 431 481 481 507
rect 507 481 513 507
rect -513 431 513 481
rect -513 405 -507 431
rect -481 405 -431 431
rect -405 405 -355 431
rect -329 405 -279 431
rect -253 405 -203 431
rect -177 405 -127 431
rect -101 405 -51 431
rect -25 405 25 431
rect 51 405 101 431
rect 127 405 177 431
rect 203 405 253 431
rect 279 405 329 431
rect 355 405 405 431
rect 431 405 481 431
rect 507 405 513 431
rect -513 355 513 405
rect -513 329 -507 355
rect -481 329 -431 355
rect -405 329 -355 355
rect -329 329 -279 355
rect -253 329 -203 355
rect -177 329 -127 355
rect -101 329 -51 355
rect -25 329 25 355
rect 51 329 101 355
rect 127 329 177 355
rect 203 329 253 355
rect 279 329 329 355
rect 355 329 405 355
rect 431 329 481 355
rect 507 329 513 355
rect -513 279 513 329
rect -513 253 -507 279
rect -481 253 -431 279
rect -405 253 -355 279
rect -329 253 -279 279
rect -253 253 -203 279
rect -177 253 -127 279
rect -101 253 -51 279
rect -25 253 25 279
rect 51 253 101 279
rect 127 253 177 279
rect 203 253 253 279
rect 279 253 329 279
rect 355 253 405 279
rect 431 253 481 279
rect 507 253 513 279
rect -513 203 513 253
rect -513 177 -507 203
rect -481 177 -431 203
rect -405 177 -355 203
rect -329 177 -279 203
rect -253 177 -203 203
rect -177 177 -127 203
rect -101 177 -51 203
rect -25 177 25 203
rect 51 177 101 203
rect 127 177 177 203
rect 203 177 253 203
rect 279 177 329 203
rect 355 177 405 203
rect 431 177 481 203
rect 507 177 513 203
rect -513 127 513 177
rect -513 101 -507 127
rect -481 101 -431 127
rect -405 101 -355 127
rect -329 101 -279 127
rect -253 101 -203 127
rect -177 101 -127 127
rect -101 101 -51 127
rect -25 101 25 127
rect 51 101 101 127
rect 127 101 177 127
rect 203 101 253 127
rect 279 101 329 127
rect 355 101 405 127
rect 431 101 481 127
rect 507 101 513 127
rect -513 51 513 101
rect -513 25 -507 51
rect -481 25 -431 51
rect -405 25 -355 51
rect -329 25 -279 51
rect -253 25 -203 51
rect -177 25 -127 51
rect -101 25 -51 51
rect -25 25 25 51
rect 51 25 101 51
rect 127 25 177 51
rect 203 25 253 51
rect 279 25 329 51
rect 355 25 405 51
rect 431 25 481 51
rect 507 25 513 51
rect -513 -25 513 25
rect -513 -51 -507 -25
rect -481 -51 -431 -25
rect -405 -51 -355 -25
rect -329 -51 -279 -25
rect -253 -51 -203 -25
rect -177 -51 -127 -25
rect -101 -51 -51 -25
rect -25 -51 25 -25
rect 51 -51 101 -25
rect 127 -51 177 -25
rect 203 -51 253 -25
rect 279 -51 329 -25
rect 355 -51 405 -25
rect 431 -51 481 -25
rect 507 -51 513 -25
rect -513 -101 513 -51
rect -513 -127 -507 -101
rect -481 -127 -431 -101
rect -405 -127 -355 -101
rect -329 -127 -279 -101
rect -253 -127 -203 -101
rect -177 -127 -127 -101
rect -101 -127 -51 -101
rect -25 -127 25 -101
rect 51 -127 101 -101
rect 127 -127 177 -101
rect 203 -127 253 -101
rect 279 -127 329 -101
rect 355 -127 405 -101
rect 431 -127 481 -101
rect 507 -127 513 -101
rect -513 -177 513 -127
rect -513 -203 -507 -177
rect -481 -203 -431 -177
rect -405 -203 -355 -177
rect -329 -203 -279 -177
rect -253 -203 -203 -177
rect -177 -203 -127 -177
rect -101 -203 -51 -177
rect -25 -203 25 -177
rect 51 -203 101 -177
rect 127 -203 177 -177
rect 203 -203 253 -177
rect 279 -203 329 -177
rect 355 -203 405 -177
rect 431 -203 481 -177
rect 507 -203 513 -177
rect -513 -253 513 -203
rect -513 -279 -507 -253
rect -481 -279 -431 -253
rect -405 -279 -355 -253
rect -329 -279 -279 -253
rect -253 -279 -203 -253
rect -177 -279 -127 -253
rect -101 -279 -51 -253
rect -25 -279 25 -253
rect 51 -279 101 -253
rect 127 -279 177 -253
rect 203 -279 253 -253
rect 279 -279 329 -253
rect 355 -279 405 -253
rect 431 -279 481 -253
rect 507 -279 513 -253
rect -513 -329 513 -279
rect -513 -355 -507 -329
rect -481 -355 -431 -329
rect -405 -355 -355 -329
rect -329 -355 -279 -329
rect -253 -355 -203 -329
rect -177 -355 -127 -329
rect -101 -355 -51 -329
rect -25 -355 25 -329
rect 51 -355 101 -329
rect 127 -355 177 -329
rect 203 -355 253 -329
rect 279 -355 329 -329
rect 355 -355 405 -329
rect 431 -355 481 -329
rect 507 -355 513 -329
rect -513 -405 513 -355
rect -513 -431 -507 -405
rect -481 -431 -431 -405
rect -405 -431 -355 -405
rect -329 -431 -279 -405
rect -253 -431 -203 -405
rect -177 -431 -127 -405
rect -101 -431 -51 -405
rect -25 -431 25 -405
rect 51 -431 101 -405
rect 127 -431 177 -405
rect 203 -431 253 -405
rect 279 -431 329 -405
rect 355 -431 405 -405
rect 431 -431 481 -405
rect 507 -431 513 -405
rect -513 -481 513 -431
rect -513 -507 -507 -481
rect -481 -507 -431 -481
rect -405 -507 -355 -481
rect -329 -507 -279 -481
rect -253 -507 -203 -481
rect -177 -507 -127 -481
rect -101 -507 -51 -481
rect -25 -507 25 -481
rect 51 -507 101 -481
rect 127 -507 177 -481
rect 203 -507 253 -481
rect 279 -507 329 -481
rect 355 -507 405 -481
rect 431 -507 481 -481
rect 507 -507 513 -481
rect -513 -557 513 -507
rect -513 -583 -507 -557
rect -481 -583 -431 -557
rect -405 -583 -355 -557
rect -329 -583 -279 -557
rect -253 -583 -203 -557
rect -177 -583 -127 -557
rect -101 -583 -51 -557
rect -25 -583 25 -557
rect 51 -583 101 -557
rect 127 -583 177 -557
rect 203 -583 253 -557
rect 279 -583 329 -557
rect 355 -583 405 -557
rect 431 -583 481 -557
rect 507 -583 513 -557
rect -513 -633 513 -583
rect -513 -659 -507 -633
rect -481 -659 -431 -633
rect -405 -659 -355 -633
rect -329 -659 -279 -633
rect -253 -659 -203 -633
rect -177 -659 -127 -633
rect -101 -659 -51 -633
rect -25 -659 25 -633
rect 51 -659 101 -633
rect 127 -659 177 -633
rect 203 -659 253 -633
rect 279 -659 329 -633
rect 355 -659 405 -633
rect 431 -659 481 -633
rect 507 -659 513 -633
rect -513 -709 513 -659
rect -513 -735 -507 -709
rect -481 -735 -431 -709
rect -405 -735 -355 -709
rect -329 -735 -279 -709
rect -253 -735 -203 -709
rect -177 -735 -127 -709
rect -101 -735 -51 -709
rect -25 -735 25 -709
rect 51 -735 101 -709
rect 127 -735 177 -709
rect 203 -735 253 -709
rect 279 -735 329 -709
rect 355 -735 405 -709
rect 431 -735 481 -709
rect 507 -735 513 -709
rect -513 -785 513 -735
rect -513 -811 -507 -785
rect -481 -811 -431 -785
rect -405 -811 -355 -785
rect -329 -811 -279 -785
rect -253 -811 -203 -785
rect -177 -811 -127 -785
rect -101 -811 -51 -785
rect -25 -811 25 -785
rect 51 -811 101 -785
rect 127 -811 177 -785
rect 203 -811 253 -785
rect 279 -811 329 -785
rect 355 -811 405 -785
rect 431 -811 481 -785
rect 507 -811 513 -785
rect -513 -861 513 -811
rect -513 -887 -507 -861
rect -481 -887 -431 -861
rect -405 -887 -355 -861
rect -329 -887 -279 -861
rect -253 -887 -203 -861
rect -177 -887 -127 -861
rect -101 -887 -51 -861
rect -25 -887 25 -861
rect 51 -887 101 -861
rect 127 -887 177 -861
rect 203 -887 253 -861
rect 279 -887 329 -861
rect 355 -887 405 -861
rect 431 -887 481 -861
rect 507 -887 513 -861
rect -513 -937 513 -887
rect -513 -963 -507 -937
rect -481 -963 -431 -937
rect -405 -963 -355 -937
rect -329 -963 -279 -937
rect -253 -963 -203 -937
rect -177 -963 -127 -937
rect -101 -963 -51 -937
rect -25 -963 25 -937
rect 51 -963 101 -937
rect 127 -963 177 -937
rect 203 -963 253 -937
rect 279 -963 329 -937
rect 355 -963 405 -937
rect 431 -963 481 -937
rect 507 -963 513 -937
rect -513 -1013 513 -963
rect -513 -1039 -507 -1013
rect -481 -1039 -431 -1013
rect -405 -1039 -355 -1013
rect -329 -1039 -279 -1013
rect -253 -1039 -203 -1013
rect -177 -1039 -127 -1013
rect -101 -1039 -51 -1013
rect -25 -1039 25 -1013
rect 51 -1039 101 -1013
rect 127 -1039 177 -1013
rect 203 -1039 253 -1013
rect 279 -1039 329 -1013
rect 355 -1039 405 -1013
rect 431 -1039 481 -1013
rect 507 -1039 513 -1013
rect -513 -1089 513 -1039
rect -513 -1115 -507 -1089
rect -481 -1115 -431 -1089
rect -405 -1115 -355 -1089
rect -329 -1115 -279 -1089
rect -253 -1115 -203 -1089
rect -177 -1115 -127 -1089
rect -101 -1115 -51 -1089
rect -25 -1115 25 -1089
rect 51 -1115 101 -1089
rect 127 -1115 177 -1089
rect 203 -1115 253 -1089
rect 279 -1115 329 -1089
rect 355 -1115 405 -1089
rect 431 -1115 481 -1089
rect 507 -1115 513 -1089
rect -513 -1165 513 -1115
rect -513 -1191 -507 -1165
rect -481 -1191 -431 -1165
rect -405 -1191 -355 -1165
rect -329 -1191 -279 -1165
rect -253 -1191 -203 -1165
rect -177 -1191 -127 -1165
rect -101 -1191 -51 -1165
rect -25 -1191 25 -1165
rect 51 -1191 101 -1165
rect 127 -1191 177 -1165
rect 203 -1191 253 -1165
rect 279 -1191 329 -1165
rect 355 -1191 405 -1165
rect 431 -1191 481 -1165
rect 507 -1191 513 -1165
rect -513 -1241 513 -1191
rect -513 -1267 -507 -1241
rect -481 -1267 -431 -1241
rect -405 -1267 -355 -1241
rect -329 -1267 -279 -1241
rect -253 -1267 -203 -1241
rect -177 -1267 -127 -1241
rect -101 -1267 -51 -1241
rect -25 -1267 25 -1241
rect 51 -1267 101 -1241
rect 127 -1267 177 -1241
rect 203 -1267 253 -1241
rect 279 -1267 329 -1241
rect 355 -1267 405 -1241
rect 431 -1267 481 -1241
rect 507 -1267 513 -1241
rect -513 -1317 513 -1267
rect -513 -1343 -507 -1317
rect -481 -1343 -431 -1317
rect -405 -1343 -355 -1317
rect -329 -1343 -279 -1317
rect -253 -1343 -203 -1317
rect -177 -1343 -127 -1317
rect -101 -1343 -51 -1317
rect -25 -1343 25 -1317
rect 51 -1343 101 -1317
rect 127 -1343 177 -1317
rect 203 -1343 253 -1317
rect 279 -1343 329 -1317
rect 355 -1343 405 -1317
rect 431 -1343 481 -1317
rect 507 -1343 513 -1317
rect -513 -1393 513 -1343
rect -513 -1419 -507 -1393
rect -481 -1419 -431 -1393
rect -405 -1419 -355 -1393
rect -329 -1419 -279 -1393
rect -253 -1419 -203 -1393
rect -177 -1419 -127 -1393
rect -101 -1419 -51 -1393
rect -25 -1419 25 -1393
rect 51 -1419 101 -1393
rect 127 -1419 177 -1393
rect 203 -1419 253 -1393
rect 279 -1419 329 -1393
rect 355 -1419 405 -1393
rect 431 -1419 481 -1393
rect 507 -1419 513 -1393
rect -513 -1469 513 -1419
rect -513 -1495 -507 -1469
rect -481 -1495 -431 -1469
rect -405 -1495 -355 -1469
rect -329 -1495 -279 -1469
rect -253 -1495 -203 -1469
rect -177 -1495 -127 -1469
rect -101 -1495 -51 -1469
rect -25 -1495 25 -1469
rect 51 -1495 101 -1469
rect 127 -1495 177 -1469
rect 203 -1495 253 -1469
rect 279 -1495 329 -1469
rect 355 -1495 405 -1469
rect 431 -1495 481 -1469
rect 507 -1495 513 -1469
rect -513 -1545 513 -1495
rect -513 -1571 -507 -1545
rect -481 -1571 -431 -1545
rect -405 -1571 -355 -1545
rect -329 -1571 -279 -1545
rect -253 -1571 -203 -1545
rect -177 -1571 -127 -1545
rect -101 -1571 -51 -1545
rect -25 -1571 25 -1545
rect 51 -1571 101 -1545
rect 127 -1571 177 -1545
rect 203 -1571 253 -1545
rect 279 -1571 329 -1545
rect 355 -1571 405 -1545
rect 431 -1571 481 -1545
rect 507 -1571 513 -1545
rect -513 -1621 513 -1571
rect -513 -1647 -507 -1621
rect -481 -1647 -431 -1621
rect -405 -1647 -355 -1621
rect -329 -1647 -279 -1621
rect -253 -1647 -203 -1621
rect -177 -1647 -127 -1621
rect -101 -1647 -51 -1621
rect -25 -1647 25 -1621
rect 51 -1647 101 -1621
rect 127 -1647 177 -1621
rect 203 -1647 253 -1621
rect 279 -1647 329 -1621
rect 355 -1647 405 -1621
rect 431 -1647 481 -1621
rect 507 -1647 513 -1621
rect -513 -1697 513 -1647
rect -513 -1723 -507 -1697
rect -481 -1723 -431 -1697
rect -405 -1723 -355 -1697
rect -329 -1723 -279 -1697
rect -253 -1723 -203 -1697
rect -177 -1723 -127 -1697
rect -101 -1723 -51 -1697
rect -25 -1723 25 -1697
rect 51 -1723 101 -1697
rect 127 -1723 177 -1697
rect 203 -1723 253 -1697
rect 279 -1723 329 -1697
rect 355 -1723 405 -1697
rect 431 -1723 481 -1697
rect 507 -1723 513 -1697
rect -513 -1773 513 -1723
rect -513 -1799 -507 -1773
rect -481 -1799 -431 -1773
rect -405 -1799 -355 -1773
rect -329 -1799 -279 -1773
rect -253 -1799 -203 -1773
rect -177 -1799 -127 -1773
rect -101 -1799 -51 -1773
rect -25 -1799 25 -1773
rect 51 -1799 101 -1773
rect 127 -1799 177 -1773
rect 203 -1799 253 -1773
rect 279 -1799 329 -1773
rect 355 -1799 405 -1773
rect 431 -1799 481 -1773
rect 507 -1799 513 -1773
rect -513 -1849 513 -1799
rect -513 -1875 -507 -1849
rect -481 -1875 -431 -1849
rect -405 -1875 -355 -1849
rect -329 -1875 -279 -1849
rect -253 -1875 -203 -1849
rect -177 -1875 -127 -1849
rect -101 -1875 -51 -1849
rect -25 -1875 25 -1849
rect 51 -1875 101 -1849
rect 127 -1875 177 -1849
rect 203 -1875 253 -1849
rect 279 -1875 329 -1849
rect 355 -1875 405 -1849
rect 431 -1875 481 -1849
rect 507 -1875 513 -1849
rect -513 -1925 513 -1875
rect -513 -1951 -507 -1925
rect -481 -1951 -431 -1925
rect -405 -1951 -355 -1925
rect -329 -1951 -279 -1925
rect -253 -1951 -203 -1925
rect -177 -1951 -127 -1925
rect -101 -1951 -51 -1925
rect -25 -1951 25 -1925
rect 51 -1951 101 -1925
rect 127 -1951 177 -1925
rect 203 -1951 253 -1925
rect 279 -1951 329 -1925
rect 355 -1951 405 -1925
rect 431 -1951 481 -1925
rect 507 -1951 513 -1925
rect -513 -2001 513 -1951
rect -513 -2027 -507 -2001
rect -481 -2027 -431 -2001
rect -405 -2027 -355 -2001
rect -329 -2027 -279 -2001
rect -253 -2027 -203 -2001
rect -177 -2027 -127 -2001
rect -101 -2027 -51 -2001
rect -25 -2027 25 -2001
rect 51 -2027 101 -2001
rect 127 -2027 177 -2001
rect 203 -2027 253 -2001
rect 279 -2027 329 -2001
rect 355 -2027 405 -2001
rect 431 -2027 481 -2001
rect 507 -2027 513 -2001
rect -513 -2077 513 -2027
rect -513 -2103 -507 -2077
rect -481 -2103 -431 -2077
rect -405 -2103 -355 -2077
rect -329 -2103 -279 -2077
rect -253 -2103 -203 -2077
rect -177 -2103 -127 -2077
rect -101 -2103 -51 -2077
rect -25 -2103 25 -2077
rect 51 -2103 101 -2077
rect 127 -2103 177 -2077
rect 203 -2103 253 -2077
rect 279 -2103 329 -2077
rect 355 -2103 405 -2077
rect 431 -2103 481 -2077
rect 507 -2103 513 -2077
rect -513 -2153 513 -2103
rect -513 -2179 -507 -2153
rect -481 -2179 -431 -2153
rect -405 -2179 -355 -2153
rect -329 -2179 -279 -2153
rect -253 -2179 -203 -2153
rect -177 -2179 -127 -2153
rect -101 -2179 -51 -2153
rect -25 -2179 25 -2153
rect 51 -2179 101 -2153
rect 127 -2179 177 -2153
rect 203 -2179 253 -2153
rect 279 -2179 329 -2153
rect 355 -2179 405 -2153
rect 431 -2179 481 -2153
rect 507 -2179 513 -2153
rect -513 -2229 513 -2179
rect -513 -2255 -507 -2229
rect -481 -2255 -431 -2229
rect -405 -2255 -355 -2229
rect -329 -2255 -279 -2229
rect -253 -2255 -203 -2229
rect -177 -2255 -127 -2229
rect -101 -2255 -51 -2229
rect -25 -2255 25 -2229
rect 51 -2255 101 -2229
rect 127 -2255 177 -2229
rect 203 -2255 253 -2229
rect 279 -2255 329 -2229
rect 355 -2255 405 -2229
rect 431 -2255 481 -2229
rect 507 -2255 513 -2229
rect -513 -2305 513 -2255
rect -513 -2331 -507 -2305
rect -481 -2331 -431 -2305
rect -405 -2331 -355 -2305
rect -329 -2331 -279 -2305
rect -253 -2331 -203 -2305
rect -177 -2331 -127 -2305
rect -101 -2331 -51 -2305
rect -25 -2331 25 -2305
rect 51 -2331 101 -2305
rect 127 -2331 177 -2305
rect 203 -2331 253 -2305
rect 279 -2331 329 -2305
rect 355 -2331 405 -2305
rect 431 -2331 481 -2305
rect 507 -2331 513 -2305
rect -513 -2381 513 -2331
rect -513 -2407 -507 -2381
rect -481 -2407 -431 -2381
rect -405 -2407 -355 -2381
rect -329 -2407 -279 -2381
rect -253 -2407 -203 -2381
rect -177 -2407 -127 -2381
rect -101 -2407 -51 -2381
rect -25 -2407 25 -2381
rect 51 -2407 101 -2381
rect 127 -2407 177 -2381
rect 203 -2407 253 -2381
rect 279 -2407 329 -2381
rect 355 -2407 405 -2381
rect 431 -2407 481 -2381
rect 507 -2407 513 -2381
rect -513 -2457 513 -2407
rect -513 -2483 -507 -2457
rect -481 -2483 -431 -2457
rect -405 -2483 -355 -2457
rect -329 -2483 -279 -2457
rect -253 -2483 -203 -2457
rect -177 -2483 -127 -2457
rect -101 -2483 -51 -2457
rect -25 -2483 25 -2457
rect 51 -2483 101 -2457
rect 127 -2483 177 -2457
rect 203 -2483 253 -2457
rect 279 -2483 329 -2457
rect 355 -2483 405 -2457
rect 431 -2483 481 -2457
rect 507 -2483 513 -2457
rect -513 -2533 513 -2483
rect -513 -2559 -507 -2533
rect -481 -2559 -431 -2533
rect -405 -2559 -355 -2533
rect -329 -2559 -279 -2533
rect -253 -2559 -203 -2533
rect -177 -2559 -127 -2533
rect -101 -2559 -51 -2533
rect -25 -2559 25 -2533
rect 51 -2559 101 -2533
rect 127 -2559 177 -2533
rect 203 -2559 253 -2533
rect 279 -2559 329 -2533
rect 355 -2559 405 -2533
rect 431 -2559 481 -2533
rect 507 -2559 513 -2533
rect -513 -2609 513 -2559
rect -513 -2635 -507 -2609
rect -481 -2635 -431 -2609
rect -405 -2635 -355 -2609
rect -329 -2635 -279 -2609
rect -253 -2635 -203 -2609
rect -177 -2635 -127 -2609
rect -101 -2635 -51 -2609
rect -25 -2635 25 -2609
rect 51 -2635 101 -2609
rect 127 -2635 177 -2609
rect 203 -2635 253 -2609
rect 279 -2635 329 -2609
rect 355 -2635 405 -2609
rect 431 -2635 481 -2609
rect 507 -2635 513 -2609
rect -513 -2641 513 -2635
<< end >>
