* NGSPICE file created from /home/shahid/GF180Projects/Layout/Magic/VCO1/INV_2/DFF_3_mag.ext - technology: gf180mcuC

.subckt pmos_3p3_YMKZL5 a_n138_n84# a_50_n84# a_n50_n128# w_n224_n214#
X0 a_50_n84# a_n50_n128# a_n138_n84# w_n224_n214# pfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
.ends

.subckt nmos_3p3_UKFAHE a_n138_n84# a_50_n84# a_n50_n128# VSUBS
X0 a_50_n84# a_n50_n128# a_n138_n84# VSUBS nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
.ends

.subckt Tr_Gate VSS OUT CLK VDD IN
Xpmos_3p3_YMKZL5_0 OUT IN a_174_n81# VDD pmos_3p3_YMKZL5
Xpmos_3p3_YMKZL5_1 IN OUT a_174_n81# VDD pmos_3p3_YMKZL5
Xpmos_3p3_YMKZL5_2 OUT IN a_174_n81# VDD pmos_3p3_YMKZL5
Xpmos_3p3_YMKZL5_3 IN OUT a_174_n81# VDD pmos_3p3_YMKZL5
Xpmos_3p3_YMKZL5_4 a_174_n81# VDD CLK VDD pmos_3p3_YMKZL5
Xpmos_3p3_YMKZL5_5 VDD a_174_n81# CLK VDD pmos_3p3_YMKZL5
Xnmos_3p3_UKFAHE_0 OUT IN CLK VSS nmos_3p3_UKFAHE
Xpmos_3p3_YMKZL5_6 a_174_n81# VDD CLK VDD pmos_3p3_YMKZL5
Xnmos_3p3_UKFAHE_1 IN OUT CLK VSS nmos_3p3_UKFAHE
Xpmos_3p3_YMKZL5_7 VDD a_174_n81# CLK VDD pmos_3p3_YMKZL5
Xnmos_3p3_UKFAHE_2 OUT IN CLK VSS nmos_3p3_UKFAHE
Xnmos_3p3_UKFAHE_3 OUT IN CLK VSS nmos_3p3_UKFAHE
Xnmos_3p3_UKFAHE_5 a_174_n81# VSS CLK VSS nmos_3p3_UKFAHE
Xnmos_3p3_UKFAHE_4 VSS a_174_n81# CLK VSS nmos_3p3_UKFAHE
.ends

.subckt nmos_3p3_6FEA4B a_n52_n50# a_256_n94# a_52_n94# a_356_n50# a_n256_n50# a_n444_n50#
+ a_152_n50# a_n356_n94# a_n152_n94# VSUBS
X0 a_152_n50# a_52_n94# a_n52_n50# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1 a_n52_n50# a_n152_n94# a_n256_n50# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X2 a_n256_n50# a_n356_n94# a_n444_n50# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X3 a_356_n50# a_256_n94# a_152_n50# VSUBS nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
.ends

.subckt pmos_3p3_KYEELV a_152_68# a_n444_n168# a_n256_68# a_n52_68# a_52_24# a_152_n168#
+ a_n444_68# a_356_68# a_256_n212# a_n256_n168# a_n356_n212# a_n152_24# w_n530_n298#
+ a_52_n212# a_n52_n168# a_n152_n212# a_n356_24# a_356_n168# a_256_24#
X0 a_n256_n168# a_n356_n212# a_n444_n168# w_n530_n298# pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X1 a_356_n168# a_256_n212# a_152_n168# w_n530_n298# pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X2 a_152_68# a_52_24# a_n52_68# w_n530_n298# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X3 a_n52_68# a_n152_24# a_n256_68# w_n530_n298# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X4 a_152_n168# a_52_n212# a_n52_n168# w_n530_n298# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X5 a_356_68# a_256_24# a_152_68# w_n530_n298# pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X6 a_n52_n168# a_n152_n212# a_n256_n168# w_n530_n298# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X7 a_n256_68# a_n356_24# a_n444_68# w_n530_n298# pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
.ends

.subckt INV_2 VDD VSS IN OUT
Xnmos_3p3_6FEA4B_0 VSS IN IN VSS OUT VSS OUT IN IN VSS nmos_3p3_6FEA4B
Xpmos_3p3_KYEELV_0 OUT VDD OUT VDD IN OUT VDD VDD IN OUT IN IN VDD IN VDD IN IN VDD
+ IN pmos_3p3_KYEELV
.ends

.subckt x/home/shahid/GF180Projects/Layout/Magic/VCO1/INV_2/DFF_3_mag D CLK Q Q- VSS
+ VDD
XTr_Gate_3 VSS INV_2_1/IN CLK VDD INV_2_5/OUT Tr_Gate
XINV_2_0 VDD VSS CLK INV_2_0/OUT INV_2
XINV_2_1 VDD VSS INV_2_1/IN INV_2_5/IN INV_2
XINV_2_2 VDD VSS Q Q- INV_2
XINV_2_3 VDD VSS INV_2_3/IN Q INV_2
XINV_2_4 VDD VSS Q INV_2_4/OUT INV_2
XINV_2_5 VDD VSS INV_2_5/IN INV_2_5/OUT INV_2
XTr_Gate_0 VSS INV_2_3/IN INV_2_0/OUT VDD INV_2_4/OUT Tr_Gate
XTr_Gate_1 VSS INV_2_3/IN CLK VDD INV_2_5/IN Tr_Gate
XTr_Gate_2 VSS INV_2_1/IN INV_2_0/OUT VDD D Tr_Gate
.ends

