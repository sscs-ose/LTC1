magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2205 -2083 7981 10547
<< isosubstrate >>
rect -83 -83 5981 8547
<< nwell >>
rect -83 6391 5981 8547
rect 454 3720 5444 5844
rect -83 2617 5981 3173
rect -83 473 473 2617
rect 5425 473 5981 2617
rect -83 -83 5981 473
<< psubdiff >>
rect 537 2280 5361 2524
rect 537 1744 781 2280
rect 5117 1744 5361 2280
rect 537 1346 5361 1744
rect 537 810 781 1346
rect 5117 810 5361 1346
rect 537 566 5361 810
<< nsubdiff >>
rect 537 5517 5361 5761
rect 537 4981 781 5517
rect 5117 4981 5361 5517
rect 537 4583 5361 4981
rect 537 4047 781 4583
rect 5117 4047 5361 4583
rect 537 3803 5361 4047
<< metal1 >>
rect 379 8085 465 8453
rect 5433 8085 5519 8453
rect 1771 7781 4127 7961
rect 1771 6977 4127 7157
rect 379 6485 465 6853
rect 5433 6485 5519 6853
rect 379 5948 465 6316
rect 5433 5948 5519 6316
rect 548 5528 5350 5750
rect 548 4970 770 5528
rect 5128 4970 5350 5528
rect 548 4594 5350 4970
rect 548 4036 770 4594
rect 5128 4036 5350 4594
rect 548 3814 5350 4036
rect 379 3248 465 3616
rect 5433 3248 5519 3616
rect 379 2711 465 3079
rect 5433 2711 5519 3079
rect 548 2291 5350 2513
rect 548 1733 770 2291
rect 5128 1733 5350 2291
rect 548 1357 5350 1733
rect 548 799 770 1357
rect 5128 799 5350 1357
rect 548 577 5350 799
rect 379 11 465 379
rect 5433 11 5519 379
<< metal2 >>
rect 11 8085 2582 8453
rect 3316 8085 5887 8453
rect 11 6485 379 8085
rect 1766 7781 4130 7961
rect 949 6485 4949 7157
rect 5519 6485 5887 8085
rect 548 4859 770 5750
rect 11 3539 379 4659
rect 949 3439 1395 6485
rect 1455 3814 1901 5750
rect 1961 3439 2407 6485
rect 2467 3814 2913 5750
rect 2985 3814 3431 5750
rect 3491 3439 3937 6485
rect 3997 3814 4443 5750
rect 4503 3439 4949 6485
rect 5128 4859 5350 5750
rect -205 2939 4949 3439
rect 5519 3259 5887 4659
rect 11 1659 379 2839
rect 548 780 770 1428
rect 949 978 1395 2939
rect 1455 780 1901 2513
rect 1961 978 2407 2939
rect 2514 780 2754 2513
rect 3145 780 3385 2513
rect 3491 978 3937 2939
rect 3997 780 4443 2513
rect 4503 978 4949 2939
rect 5519 1659 5887 3059
rect 5130 780 5348 1428
rect 548 579 2774 780
rect 3124 579 5348 780
use M1_NACTIVE_CDNS_69033583165629  M1_NACTIVE_CDNS_69033583165629_0
timestamp 1713338890
transform 1 0 2949 0 1 3848
box -2395 -45 2395 45
use M1_NACTIVE_CDNS_69033583165629  M1_NACTIVE_CDNS_69033583165629_1
timestamp 1713338890
transform 1 0 2949 0 1 5716
box -2395 -45 2395 45
use M1_NACTIVE_CDNS_69033583165635  M1_NACTIVE_CDNS_69033583165635_0
timestamp 1713338890
transform 1 0 2949 0 1 195
box -2495 -195 2495 195
use M1_NACTIVE_CDNS_69033583165635  M1_NACTIVE_CDNS_69033583165635_1
timestamp 1713338890
transform 1 0 2949 0 1 2895
box -2495 -195 2495 195
use M1_NACTIVE_CDNS_69033583165635  M1_NACTIVE_CDNS_69033583165635_2
timestamp 1713338890
transform 1 0 2949 0 1 8269
box -2495 -195 2495 195
use M1_NACTIVE_CDNS_69033583165635  M1_NACTIVE_CDNS_69033583165635_3
timestamp 1713338890
transform 1 0 2949 0 1 6669
box -2495 -195 2495 195
use M1_NACTIVE_CDNS_69033583165641  M1_NACTIVE_CDNS_69033583165641_0
timestamp 1713338890
transform 1 0 582 0 1 4782
box -45 -797 45 797
use M1_NACTIVE_CDNS_69033583165641  M1_NACTIVE_CDNS_69033583165641_1
timestamp 1713338890
transform 1 0 5316 0 1 4782
box -45 -797 45 797
use M1_NACTIVE_CDNS_69033583165642  M1_NACTIVE_CDNS_69033583165642_0
timestamp 1713338890
transform 1 0 2949 0 1 4782
box -2254 -45 2254 45
use M1_NACTIVE_CDNS_69033583165643  M1_NACTIVE_CDNS_69033583165643_0
timestamp 1713338890
transform 1 0 5162 0 1 4318
box -45 -327 45 327
use M1_NACTIVE_CDNS_69033583165643  M1_NACTIVE_CDNS_69033583165643_1
timestamp 1713338890
transform 1 0 736 0 1 4318
box -45 -327 45 327
use M1_NACTIVE_CDNS_69033583165643  M1_NACTIVE_CDNS_69033583165643_2
timestamp 1713338890
transform 1 0 736 0 1 5252
box -45 -327 45 327
use M1_NACTIVE_CDNS_69033583165643  M1_NACTIVE_CDNS_69033583165643_3
timestamp 1713338890
transform 1 0 5162 0 1 5252
box -45 -327 45 327
use M1_NACTIVE_CDNS_69033583165644  M1_NACTIVE_CDNS_69033583165644_0
timestamp 1713338890
transform 1 0 2949 0 1 4628
box -2113 -45 2113 45
use M1_NACTIVE_CDNS_69033583165644  M1_NACTIVE_CDNS_69033583165644_1
timestamp 1713338890
transform 1 0 2949 0 1 4002
box -2113 -45 2113 45
use M1_NACTIVE_CDNS_69033583165644  M1_NACTIVE_CDNS_69033583165644_2
timestamp 1713338890
transform 1 0 2949 0 1 4936
box -2113 -45 2113 45
use M1_NACTIVE_CDNS_69033583165644  M1_NACTIVE_CDNS_69033583165644_3
timestamp 1713338890
transform 1 0 2949 0 1 5562
box -2113 -45 2113 45
use M1_NACTIVE_CDNS_69033583165647  M1_NACTIVE_CDNS_69033583165647_0
timestamp 1713338890
transform 1 0 195 0 1 7469
box -195 -995 195 995
use M1_NACTIVE_CDNS_69033583165647  M1_NACTIVE_CDNS_69033583165647_1
timestamp 1713338890
transform 1 0 5703 0 1 7469
box -195 -995 195 995
use M1_NACTIVE_CDNS_69033583165655  M1_NACTIVE_CDNS_69033583165655_0
timestamp 1713338890
transform 1 0 195 0 1 1545
box -195 -1545 195 1545
use M1_NACTIVE_CDNS_69033583165655  M1_NACTIVE_CDNS_69033583165655_1
timestamp 1713338890
transform 1 0 5703 0 1 1545
box -195 -1545 195 1545
use M1_PSUB_CDNS_6903358316545  M1_PSUB_CDNS_6903358316545_0
timestamp 1713338890
transform 1 0 736 0 1 1081
box -45 -327 45 327
use M1_PSUB_CDNS_6903358316545  M1_PSUB_CDNS_6903358316545_1
timestamp 1713338890
transform 1 0 5162 0 1 1081
box -45 -327 45 327
use M1_PSUB_CDNS_6903358316545  M1_PSUB_CDNS_6903358316545_2
timestamp 1713338890
transform 1 0 736 0 1 2015
box -45 -327 45 327
use M1_PSUB_CDNS_6903358316545  M1_PSUB_CDNS_6903358316545_3
timestamp 1713338890
transform 1 0 5162 0 1 2015
box -45 -327 45 327
use M1_PSUB_CDNS_69033583165599  M1_PSUB_CDNS_69033583165599_0
timestamp 1713338890
transform 1 0 582 0 1 1545
box -45 -797 45 797
use M1_PSUB_CDNS_69033583165599  M1_PSUB_CDNS_69033583165599_1
timestamp 1713338890
transform 1 0 5316 0 1 1545
box -45 -797 45 797
use M1_PSUB_CDNS_69033583165630  M1_PSUB_CDNS_69033583165630_0
timestamp 1713338890
transform 1 0 195 0 1 4782
box -195 -1545 195 1545
use M1_PSUB_CDNS_69033583165630  M1_PSUB_CDNS_69033583165630_1
timestamp 1713338890
transform 1 0 5703 0 1 4782
box -195 -1545 195 1545
use M1_PSUB_CDNS_69033583165636  M1_PSUB_CDNS_69033583165636_0
timestamp 1713338890
transform 1 0 2949 0 1 3432
box -2495 -195 2495 195
use M1_PSUB_CDNS_69033583165636  M1_PSUB_CDNS_69033583165636_1
timestamp 1713338890
transform 1 0 2949 0 1 6132
box -2495 -195 2495 195
use M1_PSUB_CDNS_69033583165637  M1_PSUB_CDNS_69033583165637_0
timestamp 1713338890
transform 1 0 2949 0 1 1545
box -2254 -45 2254 45
use M1_PSUB_CDNS_69033583165638  M1_PSUB_CDNS_69033583165638_0
timestamp 1713338890
transform 1 0 2949 0 1 765
box -2113 -45 2113 45
use M1_PSUB_CDNS_69033583165638  M1_PSUB_CDNS_69033583165638_1
timestamp 1713338890
transform 1 0 2949 0 1 1391
box -2113 -45 2113 45
use M1_PSUB_CDNS_69033583165638  M1_PSUB_CDNS_69033583165638_2
timestamp 1713338890
transform 1 0 2949 0 1 1699
box -2113 -45 2113 45
use M1_PSUB_CDNS_69033583165638  M1_PSUB_CDNS_69033583165638_3
timestamp 1713338890
transform 1 0 2949 0 1 2325
box -2113 -45 2113 45
use M1_PSUB_CDNS_69033583165639  M1_PSUB_CDNS_69033583165639_0
timestamp 1713338890
transform 1 0 2949 0 1 611
box -2395 -45 2395 45
use M1_PSUB_CDNS_69033583165639  M1_PSUB_CDNS_69033583165639_1
timestamp 1713338890
transform 1 0 2949 0 1 2479
box -2395 -45 2395 45
use M2_M1_CDNS_69033583165538  M2_M1_CDNS_69033583165538_0
timestamp 1713338890
transform 1 0 2634 0 1 2402
box -90 -90 90 90
use M2_M1_CDNS_69033583165538  M2_M1_CDNS_69033583165538_1
timestamp 1713338890
transform 1 0 3265 0 1 2402
box -90 -90 90 90
use M2_M1_CDNS_69033583165574  M2_M1_CDNS_69033583165574_0
timestamp 1713338890
transform 1 0 1678 0 1 1545
box -194 -142 194 142
use M2_M1_CDNS_69033583165574  M2_M1_CDNS_69033583165574_1
timestamp 1713338890
transform 1 0 4220 0 1 1545
box -194 -142 194 142
use M2_M1_CDNS_69033583165574  M2_M1_CDNS_69033583165574_2
timestamp 1713338890
transform 1 0 1678 0 1 4782
box -194 -142 194 142
use M2_M1_CDNS_69033583165574  M2_M1_CDNS_69033583165574_3
timestamp 1713338890
transform 1 0 2690 0 1 4782
box -194 -142 194 142
use M2_M1_CDNS_69033583165574  M2_M1_CDNS_69033583165574_4
timestamp 1713338890
transform 1 0 3208 0 1 4782
box -194 -142 194 142
use M2_M1_CDNS_69033583165574  M2_M1_CDNS_69033583165574_5
timestamp 1713338890
transform 1 0 4220 0 1 4782
box -194 -142 194 142
use M2_M1_CDNS_69033583165631  M2_M1_CDNS_69033583165631_0
timestamp 1713338890
transform 1 0 2948 0 1 7871
box -1182 -90 1182 90
use M2_M1_CDNS_69033583165631  M2_M1_CDNS_69033583165631_1
timestamp 1713338890
transform 1 0 2948 0 -1 7067
box -1182 -90 1182 90
use M2_M1_CDNS_69033583165633  M2_M1_CDNS_69033583165633_0
timestamp 1713338890
transform 1 0 5703 0 1 2359
box -146 -686 146 686
use M2_M1_CDNS_69033583165633  M2_M1_CDNS_69033583165633_1
timestamp 1713338890
transform 1 0 5703 0 1 3959
box -146 -686 146 686
use M2_M1_CDNS_69033583165634  M2_M1_CDNS_69033583165634_0
timestamp 1713338890
transform 1 0 195 0 1 4099
box -146 -524 146 524
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_0
timestamp 1713338890
transform 1 0 1172 0 1 1078
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_1
timestamp 1713338890
transform 1 0 2184 0 1 1078
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_2
timestamp 1713338890
transform 1 0 4726 0 1 1078
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_3
timestamp 1713338890
transform 1 0 3714 0 1 1078
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_4
timestamp 1713338890
transform 1 0 1172 0 1 2012
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_5
timestamp 1713338890
transform 1 0 2184 0 1 2012
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_6
timestamp 1713338890
transform 1 0 4726 0 1 2012
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_7
timestamp 1713338890
transform 1 0 3714 0 1 2012
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_8
timestamp 1713338890
transform 1 0 1678 0 1 2402
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_9
timestamp 1713338890
transform 1 0 4220 0 1 2402
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_10
timestamp 1713338890
transform 1 0 1678 0 1 3925
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_11
timestamp 1713338890
transform 1 0 2690 0 1 3925
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_12
timestamp 1713338890
transform 1 0 3208 0 1 3925
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_13
timestamp 1713338890
transform 1 0 4220 0 1 3925
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_14
timestamp 1713338890
transform 1 0 3714 0 1 4315
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_15
timestamp 1713338890
transform 1 0 1172 0 1 4315
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_16
timestamp 1713338890
transform 1 0 2184 0 1 4315
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_17
timestamp 1713338890
transform 1 0 4726 0 1 4315
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_18
timestamp 1713338890
transform 1 0 1172 0 1 5249
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_19
timestamp 1713338890
transform 1 0 1678 0 1 5639
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_20
timestamp 1713338890
transform 1 0 2184 0 1 5249
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_21
timestamp 1713338890
transform 1 0 2690 0 1 5639
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_22
timestamp 1713338890
transform 1 0 3208 0 1 5639
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_23
timestamp 1713338890
transform 1 0 3714 0 1 5249
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_24
timestamp 1713338890
transform 1 0 4220 0 1 5639
box -194 -90 194 90
use M2_M1_CDNS_69033583165640  M2_M1_CDNS_69033583165640_25
timestamp 1713338890
transform 1 0 4726 0 1 5249
box -194 -90 194 90
use M2_M1_CDNS_69033583165646  M2_M1_CDNS_69033583165646_0
timestamp 1713338890
transform 0 1 195 -1 0 7469
box -956 -146 956 146
use M2_M1_CDNS_69033583165646  M2_M1_CDNS_69033583165646_1
timestamp 1713338890
transform 0 1 5703 -1 0 7469
box -956 -146 956 146
use M2_M1_CDNS_69033583165648  M2_M1_CDNS_69033583165648_0
timestamp 1713338890
transform 1 0 1518 0 1 8269
box -1064 -146 1064 146
use M2_M1_CDNS_69033583165648  M2_M1_CDNS_69033583165648_1
timestamp 1713338890
transform 1 0 4380 0 1 8269
box -1064 -146 1064 146
use M2_M1_CDNS_69033583165651  M2_M1_CDNS_69033583165651_0
timestamp 1713338890
transform 1 0 659 0 1 1012
box -92 -416 92 416
use M2_M1_CDNS_69033583165651  M2_M1_CDNS_69033583165651_1
timestamp 1713338890
transform 1 0 5239 0 1 1012
box -92 -416 92 416
use M2_M1_CDNS_69033583165651  M2_M1_CDNS_69033583165651_2
timestamp 1713338890
transform 1 0 659 0 1 5304
box -92 -416 92 416
use M2_M1_CDNS_69033583165651  M2_M1_CDNS_69033583165651_3
timestamp 1713338890
transform 1 0 5239 0 1 5304
box -92 -416 92 416
use M2_M1_CDNS_69033583165652  M2_M1_CDNS_69033583165652_0
timestamp 1713338890
transform 1 0 1761 0 1 688
box -956 -92 956 92
use M2_M1_CDNS_69033583165652  M2_M1_CDNS_69033583165652_1
timestamp 1713338890
transform 1 0 4137 0 1 688
box -956 -92 956 92
use M2_M1_CDNS_69033583165653  M2_M1_CDNS_69033583165653_0
timestamp 1713338890
transform 1 0 2632 0 1 1545
box -90 -142 90 142
use M2_M1_CDNS_69033583165653  M2_M1_CDNS_69033583165653_1
timestamp 1713338890
transform 1 0 3263 0 1 1545
box -90 -142 90 142
use M2_M1_CDNS_69033583165656  M2_M1_CDNS_69033583165656_0
timestamp 1713338890
transform 1 0 195 0 1 2255
box -146 -578 146 578
use M3_M2_CDNS_69033583165560  M3_M2_CDNS_69033583165560_0
timestamp 1713338890
transform 1 0 5703 0 1 2366
box -180 -677 180 677
use M3_M2_CDNS_69033583165560  M3_M2_CDNS_69033583165560_1
timestamp 1713338890
transform 1 0 5703 0 1 3959
box -180 -677 180 677
use M3_M2_CDNS_69033583165560  M3_M2_CDNS_69033583165560_2
timestamp 1713338890
transform 1 0 195 0 1 7168
box -180 -677 180 677
use M3_M2_CDNS_69033583165560  M3_M2_CDNS_69033583165560_3
timestamp 1713338890
transform 1 0 5703 0 1 7168
box -180 -677 180 677
use M3_M2_CDNS_69033583165632  M3_M2_CDNS_69033583165632_0
timestamp 1713338890
transform 1 0 195 0 1 2254
box -180 -535 180 535
use M3_M2_CDNS_69033583165632  M3_M2_CDNS_69033583165632_1
timestamp 1713338890
transform 1 0 195 0 1 4099
box -180 -535 180 535
use M3_M2_CDNS_69033583165645  M3_M2_CDNS_69033583165645_0
timestamp 1713338890
transform 1 0 659 0 1 5305
box -109 -393 109 393
use M3_M2_CDNS_69033583165645  M3_M2_CDNS_69033583165645_1
timestamp 1713338890
transform 1 0 5239 0 1 5305
box -109 -393 109 393
use M3_M2_CDNS_69033583165649  M3_M2_CDNS_69033583165649_0
timestamp 1713338890
transform 1 0 1260 0 1 8269
box -1245 -180 1245 180
use M3_M2_CDNS_69033583165649  M3_M2_CDNS_69033583165649_1
timestamp 1713338890
transform 1 0 4638 0 1 8269
box -1245 -180 1245 180
use M3_M2_CDNS_69033583165650  M3_M2_CDNS_69033583165650_0
timestamp 1713338890
transform 1 0 1678 0 1 5305
box -180 -393 180 393
use M3_M2_CDNS_69033583165650  M3_M2_CDNS_69033583165650_1
timestamp 1713338890
transform 1 0 2690 0 1 5305
box -180 -393 180 393
use M3_M2_CDNS_69033583165650  M3_M2_CDNS_69033583165650_2
timestamp 1713338890
transform 1 0 3208 0 1 5305
box -180 -393 180 393
use M3_M2_CDNS_69033583165650  M3_M2_CDNS_69033583165650_3
timestamp 1713338890
transform 1 0 4220 0 1 5305
box -180 -393 180 393
use M3_M2_CDNS_69033583165654  M3_M2_CDNS_69033583165654_0
timestamp 1713338890
transform 1 0 1671 0 1 688
box -1103 -109 1103 109
use M3_M2_CDNS_69033583165654  M3_M2_CDNS_69033583165654_1
timestamp 1713338890
transform 1 0 4227 0 1 688
box -1103 -109 1103 109
use M3_M2_CDNS_69033583165657  M3_M2_CDNS_69033583165657_0
timestamp 1713338890
transform 1 0 659 0 1 1177
box -109 -251 109 251
use M3_M2_CDNS_69033583165657  M3_M2_CDNS_69033583165657_1
timestamp 1713338890
transform 1 0 2634 0 1 1177
box -109 -251 109 251
use M3_M2_CDNS_69033583165657  M3_M2_CDNS_69033583165657_2
timestamp 1713338890
transform 1 0 3265 0 1 1177
box -109 -251 109 251
use M3_M2_CDNS_69033583165657  M3_M2_CDNS_69033583165657_3
timestamp 1713338890
transform 1 0 5239 0 1 1177
box -109 -251 109 251
use M3_M2_CDNS_69033583165658  M3_M2_CDNS_69033583165658_0
timestamp 1713338890
transform 1 0 1678 0 1 1177
box -180 -251 180 251
use M3_M2_CDNS_69033583165658  M3_M2_CDNS_69033583165658_1
timestamp 1713338890
transform 1 0 4220 0 1 1177
box -180 -251 180 251
use np_6p0_CDNS_4066195314526  np_6p0_CDNS_4066195314526_0
timestamp 1713338890
transform 0 1 949 -1 0 1178
box 0 0 200 4000
use np_6p0_CDNS_4066195314526  np_6p0_CDNS_4066195314526_1
timestamp 1713338890
transform 0 1 949 -1 0 2112
box 0 0 200 4000
use pn_6p0_CDNS_4066195314527  pn_6p0_CDNS_4066195314527_0
timestamp 1713338890
transform 0 1 949 -1 0 4415
box -120 -120 320 4120
use pn_6p0_CDNS_4066195314527  pn_6p0_CDNS_4066195314527_1
timestamp 1713338890
transform 0 1 949 -1 0 5349
box -120 -120 320 4120
use ppolyf_u_CDNS_4066195314525  ppolyf_u_CDNS_4066195314525_0
timestamp 1713338890
transform 0 1 2389 -1 0 7851
box 0 0 764 500
use ppolyf_u_CDNS_4066195314525  ppolyf_u_CDNS_4066195314525_1
timestamp 1713338890
transform 0 1 1769 -1 0 7851
box 0 0 764 500
use ppolyf_u_CDNS_4066195314525  ppolyf_u_CDNS_4066195314525_2
timestamp 1713338890
transform 0 1 3629 -1 0 7851
box 0 0 764 500
use ppolyf_u_CDNS_4066195314525  ppolyf_u_CDNS_4066195314525_3
timestamp 1713338890
transform 0 1 3009 -1 0 7851
box 0 0 764 500
<< labels >>
rlabel metal1 s 494 6132 494 6132 4 DVSS
port 1 nsew
rlabel metal1 s 494 8257 494 8257 4 DVDD
port 2 nsew
rlabel metal2 s 2965 7877 2965 7877 4 PAD
port 3 nsew
rlabel metal2 s 2965 6784 2965 6784 4 IP_IN
port 4 nsew
<< end >>
