magic
tech gf180mcuC
magscale 1 10
timestamp 1695284343
<< pwell >>
rect -446 3978 4332 7401
rect -446 3967 3704 3978
rect -446 3898 3732 3967
rect 3783 3963 4332 3978
rect 3798 3898 4332 3963
rect -446 3633 4332 3898
<< psubdiff >>
rect -422 7360 4308 7377
rect -422 7270 -407 7360
rect -307 7270 -207 7360
rect -107 7270 -7 7360
rect 93 7270 193 7360
rect 293 7270 393 7360
rect 493 7270 593 7360
rect 693 7270 793 7360
rect 893 7270 993 7360
rect 1093 7270 1193 7360
rect 1293 7270 1393 7360
rect 1493 7270 1593 7360
rect 1693 7270 1793 7360
rect 1893 7270 1993 7360
rect 2093 7270 2193 7360
rect 2293 7270 2393 7360
rect 2493 7270 2593 7360
rect 2693 7270 2793 7360
rect 2893 7270 2993 7360
rect 3093 7270 3193 7360
rect 3293 7270 3393 7360
rect 3493 7270 3593 7360
rect 3693 7270 3793 7360
rect 3893 7270 3993 7360
rect 4093 7270 4193 7360
rect 4293 7270 4308 7360
rect -422 7257 4308 7270
rect -422 7160 -292 7257
rect -422 7070 -407 7160
rect -307 7070 -292 7160
rect -422 6960 -292 7070
rect -422 6870 -407 6960
rect -307 6870 -292 6960
rect -422 6760 -292 6870
rect -422 6670 -407 6760
rect -307 6670 -292 6760
rect -422 6560 -292 6670
rect -422 6470 -407 6560
rect -307 6470 -292 6560
rect -422 6360 -292 6470
rect -422 6270 -407 6360
rect -307 6270 -292 6360
rect -422 6160 -292 6270
rect -422 6070 -407 6160
rect -307 6070 -292 6160
rect -422 5960 -292 6070
rect -422 5870 -407 5960
rect -307 5870 -292 5960
rect -422 5760 -292 5870
rect -422 5670 -407 5760
rect -307 5670 -292 5760
rect -422 5560 -292 5670
rect -422 5470 -407 5560
rect -307 5470 -292 5560
rect -422 5360 -292 5470
rect -422 5270 -407 5360
rect -307 5270 -292 5360
rect -422 5160 -292 5270
rect -422 5070 -407 5160
rect -307 5070 -292 5160
rect -422 4960 -292 5070
rect -422 4870 -407 4960
rect -307 4870 -292 4960
rect -422 4760 -292 4870
rect -422 4670 -407 4760
rect -307 4670 -292 4760
rect -422 4560 -292 4670
rect -422 4470 -407 4560
rect -307 4470 -292 4560
rect -422 4360 -292 4470
rect -422 4270 -407 4360
rect -307 4270 -292 4360
rect -422 4160 -292 4270
rect -422 4070 -407 4160
rect -307 4070 -292 4160
rect -422 3960 -292 4070
rect 4178 7160 4308 7257
rect 4178 7070 4193 7160
rect 4293 7070 4308 7160
rect 4178 6960 4308 7070
rect 4178 6870 4193 6960
rect 4293 6870 4308 6960
rect 4178 6760 4308 6870
rect 4178 6670 4193 6760
rect 4293 6670 4308 6760
rect 4178 6560 4308 6670
rect 4178 6470 4193 6560
rect 4293 6470 4308 6560
rect 4178 6360 4308 6470
rect 4178 6270 4193 6360
rect 4293 6270 4308 6360
rect 4178 6160 4308 6270
rect 4178 6070 4193 6160
rect 4293 6070 4308 6160
rect 4178 5960 4308 6070
rect 4178 5870 4193 5960
rect 4293 5870 4308 5960
rect 4178 5760 4308 5870
rect 4178 5670 4193 5760
rect 4293 5670 4308 5760
rect 4178 5560 4308 5670
rect 4178 5470 4193 5560
rect 4293 5470 4308 5560
rect 4178 5360 4308 5470
rect 4178 5270 4193 5360
rect 4293 5270 4308 5360
rect 4178 5160 4308 5270
rect 4178 5070 4193 5160
rect 4293 5070 4308 5160
rect 4178 4960 4308 5070
rect 4178 4870 4193 4960
rect 4293 4870 4308 4960
rect 4178 4760 4308 4870
rect 4178 4670 4193 4760
rect 4293 4670 4308 4760
rect 4178 4560 4308 4670
rect 4178 4470 4193 4560
rect 4293 4470 4308 4560
rect 4178 4360 4308 4470
rect 4178 4270 4193 4360
rect 4293 4270 4308 4360
rect 4178 4160 4308 4270
rect 4178 4070 4193 4160
rect 4293 4070 4308 4160
rect -422 3870 -407 3960
rect -307 3870 -292 3960
rect 4178 3960 4308 4070
rect -422 3777 -292 3870
rect 4178 3870 4193 3960
rect 4293 3870 4308 3960
rect 4178 3777 4308 3870
rect -422 3760 4308 3777
rect -422 3670 -407 3760
rect -307 3670 -207 3760
rect -107 3670 -7 3760
rect 93 3670 193 3760
rect 293 3670 393 3760
rect 493 3670 593 3760
rect 693 3670 793 3760
rect 893 3670 993 3760
rect 1093 3670 1193 3760
rect 1293 3670 1393 3760
rect 1493 3670 1593 3760
rect 1693 3670 1793 3760
rect 1893 3670 1993 3760
rect 2093 3670 2193 3760
rect 2293 3670 2393 3760
rect 2493 3670 2593 3760
rect 2693 3670 2793 3760
rect 2893 3670 2993 3760
rect 3093 3670 3193 3760
rect 3293 3670 3393 3760
rect 3493 3670 3593 3760
rect 3693 3670 3793 3760
rect 3893 3670 3993 3760
rect 4093 3670 4193 3760
rect 4293 3670 4308 3760
rect -422 3657 4308 3670
<< psubdiffcont >>
rect -407 7270 -307 7360
rect -207 7270 -107 7360
rect -7 7270 93 7360
rect 193 7270 293 7360
rect 393 7270 493 7360
rect 593 7270 693 7360
rect 793 7270 893 7360
rect 993 7270 1093 7360
rect 1193 7270 1293 7360
rect 1393 7270 1493 7360
rect 1593 7270 1693 7360
rect 1793 7270 1893 7360
rect 1993 7270 2093 7360
rect 2193 7270 2293 7360
rect 2393 7270 2493 7360
rect 2593 7270 2693 7360
rect 2793 7270 2893 7360
rect 2993 7270 3093 7360
rect 3193 7270 3293 7360
rect 3393 7270 3493 7360
rect 3593 7270 3693 7360
rect 3793 7270 3893 7360
rect 3993 7270 4093 7360
rect 4193 7270 4293 7360
rect -407 7070 -307 7160
rect -407 6870 -307 6960
rect -407 6670 -307 6760
rect -407 6470 -307 6560
rect -407 6270 -307 6360
rect -407 6070 -307 6160
rect -407 5870 -307 5960
rect -407 5670 -307 5760
rect -407 5470 -307 5560
rect -407 5270 -307 5360
rect -407 5070 -307 5160
rect -407 4870 -307 4960
rect -407 4670 -307 4760
rect -407 4470 -307 4560
rect -407 4270 -307 4360
rect -407 4070 -307 4160
rect 4193 7070 4293 7160
rect 4193 6870 4293 6960
rect 4193 6670 4293 6760
rect 4193 6470 4293 6560
rect 4193 6270 4293 6360
rect 4193 6070 4293 6160
rect 4193 5870 4293 5960
rect 4193 5670 4293 5760
rect 4193 5470 4293 5560
rect 4193 5270 4293 5360
rect 4193 5070 4293 5160
rect 4193 4870 4293 4960
rect 4193 4670 4293 4760
rect 4193 4470 4293 4560
rect 4193 4270 4293 4360
rect 4193 4070 4293 4160
rect -407 3870 -307 3960
rect 4193 3870 4293 3960
rect -407 3670 -307 3760
rect -207 3670 -107 3760
rect -7 3670 93 3760
rect 193 3670 293 3760
rect 393 3670 493 3760
rect 593 3670 693 3760
rect 793 3670 893 3760
rect 993 3670 1093 3760
rect 1193 3670 1293 3760
rect 1393 3670 1493 3760
rect 1593 3670 1693 3760
rect 1793 3670 1893 3760
rect 1993 3670 2093 3760
rect 2193 3670 2293 3760
rect 2393 3670 2493 3760
rect 2593 3670 2693 3760
rect 2793 3670 2893 3760
rect 2993 3670 3093 3760
rect 3193 3670 3293 3760
rect 3393 3670 3493 3760
rect 3593 3670 3693 3760
rect 3793 3670 3893 3760
rect 3993 3670 4093 3760
rect 4193 3670 4293 3760
<< polysilicon >>
rect 75 3960 167 3981
rect 75 3909 95 3960
rect 146 3949 167 3960
rect 146 3909 697 3949
rect 75 3899 697 3909
rect 75 3889 167 3899
<< polycontact >>
rect 95 3909 146 3960
<< metal1 >>
rect 3645 7677 3729 7689
rect 3645 7621 3661 7677
rect 3716 7621 3729 7677
rect 3645 7608 3729 7621
rect 3846 7674 3930 7686
rect 3846 7618 3862 7674
rect 3917 7618 3930 7674
rect 3846 7605 3930 7618
rect 3643 7543 3727 7555
rect 3643 7487 3659 7543
rect 3714 7487 3727 7543
rect 3643 7474 3727 7487
rect 3851 7538 3935 7550
rect 3851 7482 3867 7538
rect 3922 7482 3935 7538
rect 3851 7469 3935 7482
rect -422 7360 -292 7377
rect -422 7270 -407 7360
rect -307 7343 -292 7360
rect -222 7360 -92 7377
rect -222 7343 -207 7360
rect -307 7297 -207 7343
rect -307 7270 -292 7297
rect -422 7257 -292 7270
rect -222 7270 -207 7297
rect -107 7343 -92 7360
rect -22 7360 108 7377
rect -22 7343 -7 7360
rect -107 7297 -7 7343
rect -107 7270 -92 7297
rect -222 7257 -92 7270
rect -22 7270 -7 7297
rect 93 7343 108 7360
rect 178 7360 308 7377
rect 178 7343 193 7360
rect 93 7297 193 7343
rect 93 7270 108 7297
rect -22 7257 108 7270
rect 178 7270 193 7297
rect 293 7343 308 7360
rect 378 7360 508 7377
rect 378 7343 393 7360
rect 293 7297 393 7343
rect 293 7270 308 7297
rect 178 7257 308 7270
rect 378 7270 393 7297
rect 493 7343 508 7360
rect 578 7360 708 7377
rect 578 7343 593 7360
rect 493 7297 593 7343
rect 493 7270 508 7297
rect 378 7257 508 7270
rect 578 7270 593 7297
rect 693 7343 708 7360
rect 778 7360 908 7377
rect 778 7343 793 7360
rect 693 7297 793 7343
rect 693 7270 708 7297
rect 578 7257 708 7270
rect 778 7270 793 7297
rect 893 7343 908 7360
rect 978 7360 1108 7377
rect 978 7343 993 7360
rect 893 7297 993 7343
rect 893 7270 908 7297
rect 778 7257 908 7270
rect 978 7270 993 7297
rect 1093 7343 1108 7360
rect 1178 7360 1308 7377
rect 1178 7343 1193 7360
rect 1093 7297 1193 7343
rect 1093 7270 1108 7297
rect 978 7257 1108 7270
rect 1178 7270 1193 7297
rect 1293 7343 1308 7360
rect 1378 7360 1508 7377
rect 1378 7343 1393 7360
rect 1293 7297 1393 7343
rect 1293 7270 1308 7297
rect 1178 7257 1308 7270
rect 1378 7270 1393 7297
rect 1493 7343 1508 7360
rect 1578 7360 1708 7377
rect 1578 7343 1593 7360
rect 1493 7297 1593 7343
rect 1493 7270 1508 7297
rect 1378 7257 1508 7270
rect 1578 7270 1593 7297
rect 1693 7343 1708 7360
rect 1778 7360 1908 7377
rect 1778 7343 1793 7360
rect 1693 7297 1793 7343
rect 1693 7270 1708 7297
rect 1578 7257 1708 7270
rect 1778 7270 1793 7297
rect 1893 7343 1908 7360
rect 1978 7360 2108 7377
rect 1978 7343 1993 7360
rect 1893 7297 1993 7343
rect 1893 7270 1908 7297
rect 1778 7257 1908 7270
rect 1978 7270 1993 7297
rect 2093 7343 2108 7360
rect 2178 7360 2308 7377
rect 2178 7343 2193 7360
rect 2093 7297 2193 7343
rect 2093 7270 2108 7297
rect 1978 7257 2108 7270
rect 2178 7270 2193 7297
rect 2293 7343 2308 7360
rect 2378 7360 2508 7377
rect 2378 7343 2393 7360
rect 2293 7297 2393 7343
rect 2293 7270 2308 7297
rect 2178 7257 2308 7270
rect 2378 7270 2393 7297
rect 2493 7343 2508 7360
rect 2578 7360 2708 7377
rect 2578 7343 2593 7360
rect 2493 7297 2593 7343
rect 2493 7270 2508 7297
rect 2378 7257 2508 7270
rect 2578 7270 2593 7297
rect 2693 7343 2708 7360
rect 2778 7360 2908 7377
rect 2778 7343 2793 7360
rect 2693 7297 2793 7343
rect 2693 7270 2708 7297
rect 2578 7257 2708 7270
rect 2778 7270 2793 7297
rect 2893 7343 2908 7360
rect 2978 7360 3108 7377
rect 2978 7343 2993 7360
rect 2893 7297 2993 7343
rect 2893 7270 2908 7297
rect 2778 7257 2908 7270
rect 2978 7270 2993 7297
rect 3093 7343 3108 7360
rect 3178 7360 3308 7377
rect 3178 7343 3193 7360
rect 3093 7297 3193 7343
rect 3093 7270 3108 7297
rect 2978 7257 3108 7270
rect 3178 7270 3193 7297
rect 3293 7343 3308 7360
rect 3378 7360 3508 7377
rect 3378 7343 3393 7360
rect 3293 7297 3393 7343
rect 3293 7270 3308 7297
rect 3178 7257 3308 7270
rect 3378 7270 3393 7297
rect 3493 7343 3508 7360
rect 3578 7360 3708 7377
rect 3578 7343 3593 7360
rect 3493 7297 3593 7343
rect 3493 7270 3508 7297
rect 3378 7257 3508 7270
rect 3578 7270 3593 7297
rect 3693 7343 3708 7360
rect 3778 7360 3908 7377
rect 3778 7343 3793 7360
rect 3693 7297 3793 7343
rect 3693 7270 3708 7297
rect 3578 7257 3708 7270
rect 3778 7270 3793 7297
rect 3893 7343 3908 7360
rect 3978 7360 4108 7377
rect 3978 7343 3993 7360
rect 3893 7297 3993 7343
rect 3893 7270 3908 7297
rect 3778 7257 3908 7270
rect 3978 7270 3993 7297
rect 4093 7343 4108 7360
rect 4178 7360 4308 7377
rect 4178 7343 4193 7360
rect 4093 7297 4193 7343
rect 4093 7270 4108 7297
rect 3978 7257 4108 7270
rect 4178 7270 4193 7297
rect 4293 7270 4308 7360
rect 4178 7257 4308 7270
rect -393 7177 -347 7257
rect 4220 7177 4266 7257
rect -422 7160 -292 7177
rect -422 7070 -407 7160
rect -307 7070 -292 7160
rect 454 7124 3348 7170
rect -422 7057 -292 7070
rect 81 7101 159 7113
rect -393 6977 -347 7057
rect 81 7047 93 7101
rect 147 7097 159 7101
rect 147 7051 281 7097
rect 147 7047 159 7051
rect 81 7039 159 7047
rect -422 6960 -292 6977
rect -422 6870 -407 6960
rect -307 6870 -292 6960
rect -422 6857 -292 6870
rect -393 6777 -347 6857
rect -422 6760 -292 6777
rect -422 6670 -407 6760
rect -307 6670 -292 6760
rect -422 6657 -292 6670
rect -90 6692 -12 6704
rect -393 6577 -347 6657
rect -90 6638 -78 6692
rect -24 6688 -12 6692
rect -24 6642 172 6688
rect -24 6638 -12 6642
rect -90 6632 -12 6638
rect -422 6560 -292 6577
rect -422 6470 -407 6560
rect -307 6470 -292 6560
rect -3641 6452 -2588 6462
rect -422 6457 -292 6470
rect -3641 6336 -2549 6452
rect -393 6377 -347 6457
rect -422 6360 -292 6377
rect -3641 6312 -2588 6336
rect -422 6270 -407 6360
rect -307 6270 -292 6360
rect -422 6257 -292 6270
rect 80 6302 158 6311
rect -393 6177 -347 6257
rect 80 6246 92 6302
rect 148 6246 284 6302
rect 80 6237 158 6246
rect -422 6160 -292 6177
rect -422 6070 -407 6160
rect -307 6070 -292 6160
rect -422 6057 -292 6070
rect -602 5992 -488 6038
rect -393 5977 -347 6057
rect -422 5960 -292 5977
rect -3625 5942 -2835 5960
rect -3625 5896 -2825 5942
rect -3625 5878 -2835 5896
rect -422 5870 -407 5960
rect -307 5870 -292 5960
rect -422 5857 -292 5870
rect -93 5887 -15 5894
rect -393 5777 -347 5857
rect -93 5831 -79 5887
rect -23 5831 163 5887
rect -93 5822 -15 5831
rect -422 5760 -292 5777
rect -422 5670 -407 5760
rect -307 5670 -292 5760
rect -422 5657 -292 5670
rect -393 5577 -347 5657
rect -422 5560 -292 5577
rect -422 5470 -407 5560
rect -307 5470 -292 5560
rect -422 5457 -292 5470
rect 80 5506 158 5517
rect -393 5377 -347 5457
rect 80 5450 92 5506
rect 148 5450 284 5506
rect 80 5443 158 5450
rect -422 5360 -292 5377
rect -422 5270 -407 5360
rect -307 5270 -292 5360
rect -422 5257 -292 5270
rect -393 5177 -347 5257
rect -422 5160 -292 5177
rect -422 5070 -407 5160
rect -307 5070 -292 5160
rect -422 5057 -292 5070
rect -94 5095 -11 5101
rect -2887 5007 -2815 5023
rect -716 5015 -551 5043
rect -2887 4991 -2804 5007
rect -716 4997 -617 5015
rect -3642 4917 -2790 4991
rect -673 4965 -617 4997
rect -630 4961 -617 4965
rect -563 4961 -551 5015
rect -393 4977 -347 5057
rect -94 5039 -79 5095
rect -23 5039 183 5095
rect -94 5029 -11 5039
rect -630 4954 -551 4961
rect -422 4960 -292 4977
rect -2887 4912 -2804 4917
rect -422 4870 -407 4960
rect -307 4870 -292 4960
rect -422 4857 -292 4870
rect -393 4777 -347 4857
rect -245 4838 -173 4852
rect -245 4782 -238 4838
rect -182 4782 128 4838
rect -422 4760 -292 4777
rect -245 4770 -173 4782
rect -422 4670 -407 4760
rect -307 4670 -292 4760
rect -422 4657 -292 4670
rect 72 4721 128 4782
rect 72 4711 156 4721
rect -393 4577 -347 4657
rect 72 4655 92 4711
rect 148 4655 280 4711
rect 72 4652 156 4655
rect 78 4647 156 4652
rect -422 4560 -292 4577
rect -422 4470 -407 4560
rect -307 4470 -292 4560
rect -422 4457 -292 4470
rect -393 4377 -347 4457
rect -422 4360 -292 4377
rect -422 4270 -407 4360
rect -307 4270 -292 4360
rect -422 4257 -292 4270
rect -92 4293 -10 4300
rect -393 4177 -347 4257
rect -92 4237 -79 4293
rect -23 4237 158 4293
rect -92 4228 -10 4237
rect -422 4160 -292 4177
rect -422 4070 -407 4160
rect -307 4070 -292 4160
rect -422 4057 -292 4070
rect -3573 4003 -2810 4019
rect -3573 3957 -2795 4003
rect -393 3977 -347 4057
rect 1234 3982 1325 7105
rect 1643 3982 1734 7105
rect 2058 3982 2149 7105
rect 2461 3982 2552 7111
rect 3302 7009 3348 7124
rect 4178 7160 4308 7177
rect 4178 7070 4193 7160
rect 4293 7070 4308 7160
rect 4178 7057 4308 7070
rect 4220 6977 4266 7057
rect 4178 6960 4308 6977
rect 4178 6870 4193 6960
rect 4293 6870 4308 6960
rect 4178 6857 4308 6870
rect 3824 6796 3906 6812
rect 3824 6792 3837 6796
rect 3494 6746 3837 6792
rect 3824 6742 3837 6746
rect 3891 6742 3906 6796
rect 4220 6777 4266 6857
rect 3824 6736 3906 6742
rect 4178 6760 4308 6777
rect 4178 6670 4193 6760
rect 4293 6670 4308 6760
rect 4178 6657 4308 6670
rect 4220 6577 4266 6657
rect 4178 6560 4308 6577
rect 4178 6470 4193 6560
rect 4293 6470 4308 6560
rect 4178 6457 4308 6470
rect 4220 6377 4266 6457
rect 4178 6360 4308 6377
rect 4178 6270 4193 6360
rect 4293 6270 4308 6360
rect 4178 6257 4308 6270
rect 4220 6177 4266 6257
rect 4178 6160 4308 6177
rect 4178 6070 4193 6160
rect 4293 6070 4308 6160
rect 4178 6057 4308 6070
rect 3824 5998 3906 6009
rect 3824 5995 3836 5998
rect 3526 5949 3836 5995
rect 3824 5942 3836 5949
rect 3892 5942 3906 5998
rect 4220 5977 4266 6057
rect 3824 5933 3906 5942
rect 4178 5960 4308 5977
rect 4178 5870 4193 5960
rect 4293 5870 4308 5960
rect 4178 5857 4308 5870
rect 4220 5777 4266 5857
rect 4178 5760 4308 5777
rect 4178 5670 4193 5760
rect 4293 5670 4308 5760
rect 4178 5657 4308 5670
rect 4220 5577 4266 5657
rect 4178 5560 4308 5577
rect 4178 5470 4193 5560
rect 4293 5470 4308 5560
rect 4178 5457 4308 5470
rect 4220 5377 4266 5457
rect 4178 5360 4308 5377
rect 4178 5270 4193 5360
rect 4293 5270 4308 5360
rect 4178 5257 4308 5270
rect 3822 5200 3904 5213
rect 3822 5198 3836 5200
rect 3495 5152 3836 5198
rect 3822 5144 3836 5152
rect 3892 5144 3904 5200
rect 4220 5177 4266 5257
rect 3822 5137 3904 5144
rect 4178 5160 4308 5177
rect 4178 5070 4193 5160
rect 4293 5070 4308 5160
rect 4178 5057 4308 5070
rect 4220 4977 4266 5057
rect 4178 4960 4308 4977
rect 4178 4870 4193 4960
rect 4293 4870 4308 4960
rect 4178 4857 4308 4870
rect 4220 4777 4266 4857
rect 4178 4760 4308 4777
rect 4178 4670 4193 4760
rect 4293 4670 4308 4760
rect 4178 4657 4308 4670
rect 4220 4577 4266 4657
rect 4178 4560 4308 4577
rect 4178 4470 4193 4560
rect 4293 4470 4308 4560
rect 4178 4457 4308 4470
rect 3826 4402 3908 4413
rect 3826 4401 3836 4402
rect 3507 4355 3836 4401
rect 3826 4346 3836 4355
rect 3892 4346 3908 4402
rect 4220 4377 4266 4457
rect 3826 4337 3908 4346
rect 4178 4360 4308 4377
rect 4178 4270 4193 4360
rect 4293 4270 4308 4360
rect 4178 4257 4308 4270
rect 4220 4177 4266 4257
rect 4178 4160 4308 4177
rect 4178 4070 4193 4160
rect 4293 4070 4308 4160
rect 4178 4057 4308 4070
rect 3618 4020 4015 4037
rect 3618 3982 3790 4020
rect -422 3960 -292 3977
rect -3573 3941 -2810 3957
rect -422 3870 -407 3960
rect -307 3870 -292 3960
rect 75 3963 167 3981
rect 75 3907 92 3963
rect 148 3907 167 3963
rect 75 3889 167 3907
rect 451 3966 3790 3982
rect 3844 3966 4015 4020
rect 4220 3977 4266 4057
rect 451 3952 4015 3966
rect 451 3898 3657 3952
rect 3711 3943 4015 3952
rect 3711 3898 3917 3943
rect 451 3891 3917 3898
rect 3618 3889 3917 3891
rect 3971 3889 4015 3943
rect 3618 3870 4015 3889
rect 4178 3960 4308 3977
rect 4178 3870 4193 3960
rect 4293 3870 4308 3960
rect -422 3857 -292 3870
rect 4178 3857 4308 3870
rect -393 3777 -347 3857
rect 4220 3777 4266 3857
rect -422 3760 -292 3777
rect -2784 3687 -2655 3699
rect -422 3698 -407 3760
rect -3538 3662 -2591 3687
rect -2361 3662 -2225 3673
rect -3538 3656 -2225 3662
rect -988 3670 -407 3698
rect -307 3743 -292 3760
rect -222 3760 -92 3777
rect -222 3743 -207 3760
rect -307 3670 -207 3743
rect -107 3743 -92 3760
rect -22 3760 108 3777
rect -22 3743 -7 3760
rect -107 3670 -7 3743
rect 93 3743 108 3760
rect 178 3760 308 3777
rect 178 3743 193 3760
rect 93 3670 193 3743
rect 293 3743 308 3760
rect 378 3760 508 3777
rect 378 3743 393 3760
rect 293 3670 393 3743
rect 493 3743 508 3760
rect 578 3760 708 3777
rect 578 3743 593 3760
rect 493 3670 593 3743
rect 693 3743 708 3760
rect 778 3760 908 3777
rect 778 3743 793 3760
rect 693 3670 793 3743
rect 893 3743 908 3760
rect 978 3760 1108 3777
rect 978 3743 993 3760
rect 893 3670 993 3743
rect 1093 3743 1108 3760
rect 1178 3760 1308 3777
rect 1178 3743 1193 3760
rect 1093 3670 1193 3743
rect 1293 3743 1308 3760
rect 1378 3760 1508 3777
rect 1378 3743 1393 3760
rect 1293 3670 1393 3743
rect 1493 3743 1508 3760
rect 1578 3760 1708 3777
rect 1578 3743 1593 3760
rect 1493 3670 1593 3743
rect 1693 3743 1708 3760
rect 1778 3760 1908 3777
rect 1778 3743 1793 3760
rect 1693 3670 1793 3743
rect 1893 3743 1908 3760
rect 1978 3760 2108 3777
rect 1978 3743 1993 3760
rect 1893 3670 1993 3743
rect 2093 3743 2108 3760
rect 2178 3760 2308 3777
rect 2178 3743 2193 3760
rect 2093 3670 2193 3743
rect 2293 3743 2308 3760
rect 2378 3760 2508 3777
rect 2378 3743 2393 3760
rect 2293 3670 2393 3743
rect 2493 3743 2508 3760
rect 2578 3760 2708 3777
rect 2578 3743 2593 3760
rect 2493 3670 2593 3743
rect 2693 3743 2708 3760
rect 2778 3760 2908 3777
rect 2778 3743 2793 3760
rect 2693 3670 2793 3743
rect 2893 3743 2908 3760
rect 2978 3760 3108 3777
rect 2978 3743 2993 3760
rect 2893 3670 2993 3743
rect 3093 3743 3108 3760
rect 3178 3760 3308 3777
rect 3178 3743 3193 3760
rect 3093 3670 3193 3743
rect 3293 3743 3308 3760
rect 3378 3760 3508 3777
rect 3378 3743 3393 3760
rect 3293 3670 3393 3743
rect 3493 3743 3508 3760
rect 3578 3760 3708 3777
rect 3578 3743 3593 3760
rect 3493 3670 3593 3743
rect 3693 3743 3708 3760
rect 3778 3760 3908 3777
rect 3778 3743 3793 3760
rect 3693 3670 3793 3743
rect 3893 3743 3908 3760
rect 3978 3760 4108 3777
rect 3978 3743 3993 3760
rect 3893 3697 3993 3743
rect 3893 3670 3908 3697
rect -988 3657 3908 3670
rect 3978 3670 3993 3697
rect 4093 3743 4108 3760
rect 4178 3760 4308 3777
rect 4178 3743 4193 3760
rect 4093 3697 4193 3743
rect 4093 3670 4108 3697
rect 3978 3657 4108 3670
rect 4178 3670 4193 3697
rect 4293 3670 4308 3760
rect 4178 3657 4308 3670
rect -988 3656 3879 3657
rect -3538 3570 3879 3656
rect -2784 3450 3879 3570
rect 4031 3524 4129 3540
rect 4031 3454 4046 3524
rect 4116 3454 4129 3524
rect -2784 3303 -2655 3450
rect 4031 3444 4129 3454
rect -3538 3196 -2939 3264
rect 4045 2769 4117 3444
rect -2997 2737 -2943 2738
rect -3513 2660 -2931 2737
rect 3984 2697 4117 2769
<< via1 >>
rect 3661 7621 3716 7677
rect 3862 7618 3917 7674
rect 3659 7487 3714 7543
rect 3867 7482 3922 7538
rect 93 7047 147 7101
rect -78 6638 -24 6692
rect 92 6246 148 6302
rect -79 5831 -23 5887
rect 92 5450 148 5506
rect -617 4961 -563 5015
rect -79 5039 -23 5095
rect -238 4782 -182 4838
rect 92 4655 148 4711
rect -79 4237 -23 4293
rect 3837 6742 3891 6796
rect 3836 5942 3892 5998
rect 3836 5144 3892 5200
rect 3836 4346 3892 4402
rect 92 3960 148 3963
rect 92 3909 95 3960
rect 95 3909 146 3960
rect 146 3909 148 3960
rect 92 3907 148 3909
rect 3790 3966 3844 4020
rect 3657 3898 3711 3952
rect 3917 3889 3971 3943
rect 4046 3454 4116 3524
<< metal2 >>
rect 3633 7677 3738 7695
rect 3633 7621 3661 7677
rect 3716 7621 3738 7677
rect 3633 7543 3738 7621
rect 3633 7487 3659 7543
rect 3714 7487 3738 7543
rect 81 7101 159 7113
rect 81 7047 93 7101
rect 147 7047 159 7101
rect 81 7039 159 7047
rect -90 6692 -12 6704
rect -90 6638 -78 6692
rect -24 6638 -12 6692
rect -90 6632 -12 6638
rect -79 6038 -23 6632
rect 92 6311 148 7039
rect 3633 6610 3738 7487
rect 3836 7674 3944 7693
rect 3836 7618 3862 7674
rect 3917 7618 3944 7674
rect 3836 7538 3944 7618
rect 3836 7482 3867 7538
rect 3922 7482 3944 7538
rect 3836 6812 3944 7482
rect 3824 6796 3944 6812
rect 3824 6742 3837 6796
rect 3891 6742 3944 6796
rect 3824 6736 3944 6742
rect 3531 6554 3738 6610
rect 80 6302 158 6311
rect 80 6246 92 6302
rect 148 6246 158 6302
rect 80 6237 158 6246
rect -618 5982 -23 6038
rect -79 5894 -23 5982
rect -93 5887 -15 5894
rect -93 5831 -79 5887
rect -23 5831 -15 5887
rect -93 5822 -15 5831
rect -79 5101 -23 5822
rect 92 5517 148 6237
rect 3633 5808 3738 6554
rect 3836 6009 3944 6736
rect 3824 5998 3944 6009
rect 3824 5942 3836 5998
rect 3892 5942 3944 5998
rect 3824 5933 3944 5942
rect 3530 5752 3738 5808
rect 80 5506 158 5517
rect 80 5450 92 5506
rect 148 5450 158 5506
rect 80 5443 158 5450
rect -94 5095 -11 5101
rect -94 5039 -79 5095
rect -23 5039 -11 5095
rect -94 5029 -11 5039
rect -630 5015 -551 5027
rect -630 4961 -617 5015
rect -563 4961 -551 5015
rect -630 4954 -551 4961
rect -618 4838 -562 4954
rect -245 4838 -173 4852
rect -618 4782 -238 4838
rect -182 4782 -173 4838
rect -245 4774 -173 4782
rect -245 4770 -175 4774
rect -79 4300 -23 5029
rect 92 4721 148 5443
rect 3633 5008 3738 5752
rect 3836 5213 3944 5933
rect 3822 5200 3944 5213
rect 3822 5144 3836 5200
rect 3892 5144 3944 5200
rect 3822 5137 3944 5144
rect 3544 4952 3738 5008
rect 78 4711 156 4721
rect 78 4655 92 4711
rect 148 4655 156 4711
rect 78 4647 156 4655
rect -92 4293 -10 4300
rect -92 4237 -79 4293
rect -23 4237 -10 4293
rect -92 4228 -10 4237
rect 92 3981 148 4647
rect 3633 4208 3738 4952
rect 3836 4413 3944 5137
rect 3826 4402 3944 4413
rect 3826 4346 3836 4402
rect 3892 4357 3944 4402
rect 3892 4346 3908 4357
rect 3826 4337 3908 4346
rect 3538 4152 3738 4208
rect 3605 4020 4117 4043
rect 75 3963 167 3981
rect 75 3907 92 3963
rect 148 3907 167 3963
rect 75 3889 167 3907
rect 3605 3966 3790 4020
rect 3844 3966 4117 4020
rect 3605 3952 4117 3966
rect 3605 3898 3657 3952
rect 3711 3943 4117 3952
rect 3711 3898 3917 3943
rect 3605 3889 3917 3898
rect 3971 3889 4117 3943
rect 3605 3870 4117 3889
rect 4045 3540 4117 3870
rect 4031 3524 4129 3540
rect 4031 3454 4046 3524
rect 4116 3454 4129 3524
rect 4031 3444 4129 3454
rect -2995 3104 -2937 3259
rect -569 2452 -512 2619
use CM_MSB_V2  CM_MSB_V2_0
timestamp 1693309239
transform 1 0 -2839 0 1 2178
box -171 -208 6915 1285
use Local_Enc  Local_Enc_0
timestamp 1694584912
transform 1 0 -2914 0 1 3601
box -304 -1 2426 2861
use MSB_Unit_Cell_p2  MSB_Unit_Cell_p2_0
timestamp 1691476851
transform 1 0 205 0 1 5176
box -74 -480 3384 367
use MSB_Unit_Cell_p2  MSB_Unit_Cell_p2_1
timestamp 1691476851
transform 1 0 205 0 1 4379
box -74 -480 3384 367
use MSB_Unit_Cell_p2  MSB_Unit_Cell_p2_2
timestamp 1691476851
transform 1 0 205 0 1 5973
box -74 -480 3384 367
use MSB_Unit_Cell_p2  MSB_Unit_Cell_p2_3
timestamp 1691476851
transform 1 0 205 0 1 6770
box -74 -480 3384 367
<< labels >>
flabel metal1 -3384 3241 -3384 3241 0 FreeSans 1600 0 0 0 IM_T
port 0 nsew
flabel metal1 -3340 2694 -3340 2694 0 FreeSans 1600 0 0 0 IM
port 1 nsew
flabel metal1 -3423 3612 -3423 3612 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
flabel metal1 -3204 3981 -3204 3981 0 FreeSans 1600 0 0 0 Ri
port 3 nsew
flabel metal1 -3431 4954 -3431 4954 0 FreeSans 1600 0 0 0 Ci
port 4 nsew
flabel metal1 -3540 5919 -3540 5919 0 FreeSans 1600 0 0 0 Ri-1
port 5 nsew
flabel metal1 -3483 6325 -3483 6325 0 FreeSans 1600 0 0 0 VDD
port 6 nsew
flabel metal2 -517 6019 -517 6019 0 FreeSans 1600 0 0 0 QB
port 7 nsew
flabel via1 -589 4973 -589 4973 0 FreeSans 1600 0 0 0 Q
port 8 nsew
flabel metal1 4074 2797 4074 2797 0 FreeSans 1600 0 0 0 OUT
port 9 nsew
flabel via1 3898 7510 3898 7510 0 FreeSans 1600 0 0 0 OUT+
port 10 nsew
flabel via1 3681 7653 3681 7653 0 FreeSans 1600 0 0 0 OUT-
port 11 nsew
flabel metal2 -540 2480 -540 2480 0 FreeSans 1600 0 0 0 SD
port 12 nsew
<< end >>
