magic
tech gf180mcuC
magscale 1 10
timestamp 1699871744
<< nwell >>
rect -1264 -986 1264 986
<< nsubdiff >>
rect -1240 890 1240 962
rect -1240 846 -1168 890
rect -1240 -846 -1227 846
rect -1181 -846 -1168 846
rect 1168 846 1240 890
rect -1240 -890 -1168 -846
rect 1168 -846 1181 846
rect 1227 -846 1240 846
rect 1168 -890 1240 -846
rect -1240 -962 1240 -890
<< nsubdiffcont >>
rect -1227 -846 -1181 846
rect 1181 -846 1227 846
<< polysilicon >>
rect -1080 789 -880 802
rect -1080 743 -1067 789
rect -893 743 -880 789
rect -1080 700 -880 743
rect -1080 -743 -880 -700
rect -1080 -789 -1067 -743
rect -893 -789 -880 -743
rect -1080 -802 -880 -789
rect -800 789 -600 802
rect -800 743 -787 789
rect -613 743 -600 789
rect -800 700 -600 743
rect -800 -743 -600 -700
rect -800 -789 -787 -743
rect -613 -789 -600 -743
rect -800 -802 -600 -789
rect -520 789 -320 802
rect -520 743 -507 789
rect -333 743 -320 789
rect -520 700 -320 743
rect -520 -743 -320 -700
rect -520 -789 -507 -743
rect -333 -789 -320 -743
rect -520 -802 -320 -789
rect -240 789 -40 802
rect -240 743 -227 789
rect -53 743 -40 789
rect -240 700 -40 743
rect -240 -743 -40 -700
rect -240 -789 -227 -743
rect -53 -789 -40 -743
rect -240 -802 -40 -789
rect 40 789 240 802
rect 40 743 53 789
rect 227 743 240 789
rect 40 700 240 743
rect 40 -743 240 -700
rect 40 -789 53 -743
rect 227 -789 240 -743
rect 40 -802 240 -789
rect 320 789 520 802
rect 320 743 333 789
rect 507 743 520 789
rect 320 700 520 743
rect 320 -743 520 -700
rect 320 -789 333 -743
rect 507 -789 520 -743
rect 320 -802 520 -789
rect 600 789 800 802
rect 600 743 613 789
rect 787 743 800 789
rect 600 700 800 743
rect 600 -743 800 -700
rect 600 -789 613 -743
rect 787 -789 800 -743
rect 600 -802 800 -789
rect 880 789 1080 802
rect 880 743 893 789
rect 1067 743 1080 789
rect 880 700 1080 743
rect 880 -743 1080 -700
rect 880 -789 893 -743
rect 1067 -789 1080 -743
rect 880 -802 1080 -789
<< polycontact >>
rect -1067 743 -893 789
rect -1067 -789 -893 -743
rect -787 743 -613 789
rect -787 -789 -613 -743
rect -507 743 -333 789
rect -507 -789 -333 -743
rect -227 743 -53 789
rect -227 -789 -53 -743
rect 53 743 227 789
rect 53 -789 227 -743
rect 333 743 507 789
rect 333 -789 507 -743
rect 613 743 787 789
rect 613 -789 787 -743
rect 893 743 1067 789
rect 893 -789 1067 -743
<< ppolyres >>
rect -1080 -700 -880 700
rect -800 -700 -600 700
rect -520 -700 -320 700
rect -240 -700 -40 700
rect 40 -700 240 700
rect 320 -700 520 700
rect 600 -700 800 700
rect 880 -700 1080 700
<< metal1 >>
rect -1227 903 1227 949
rect -1227 846 -1181 903
rect 1181 846 1227 903
rect -1078 743 -1067 789
rect -893 743 -882 789
rect -798 743 -787 789
rect -613 743 -602 789
rect -518 743 -507 789
rect -333 743 -322 789
rect -238 743 -227 789
rect -53 743 -42 789
rect 42 743 53 789
rect 227 743 238 789
rect 322 743 333 789
rect 507 743 518 789
rect 602 743 613 789
rect 787 743 798 789
rect 882 743 893 789
rect 1067 743 1078 789
rect -1078 -789 -1067 -743
rect -893 -789 -882 -743
rect -798 -789 -787 -743
rect -613 -789 -602 -743
rect -518 -789 -507 -743
rect -333 -789 -322 -743
rect -238 -789 -227 -743
rect -53 -789 -42 -743
rect 42 -789 53 -743
rect 227 -789 238 -743
rect 322 -789 333 -743
rect 507 -789 518 -743
rect 602 -789 613 -743
rect 787 -789 798 -743
rect 882 -789 893 -743
rect 1067 -789 1078 -743
rect -1227 -903 -1181 -846
rect 1181 -903 1227 -846
rect -1227 -949 1227 -903
<< properties >>
string FIXED_BBOX -1204 -926 1204 926
string gencell ppolyf_u
string library gf180mcu
string parameters w 1.0 l 7.0 m 1 nx 8 wmin 0.80 lmin 1.00 rho 315 val 2.37k dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 1 grc 1 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 1
<< end >>
