magic
tech gf180mcuC
magscale 1 10
timestamp 1692268103
<< mimcap >>
rect -5041 920 -3041 1000
rect -5041 -920 -4961 920
rect -3121 -920 -3041 920
rect -5041 -1000 -3041 -920
rect -2427 920 -427 1000
rect -2427 -920 -2347 920
rect -507 -920 -427 920
rect -2427 -1000 -427 -920
rect 187 920 2187 1000
rect 187 -920 267 920
rect 2107 -920 2187 920
rect 187 -1000 2187 -920
rect 2801 920 4801 1000
rect 2801 -920 2881 920
rect 4721 -920 4801 920
rect 2801 -1000 4801 -920
<< mimcapcontact >>
rect -4961 -920 -3121 920
rect -2347 -920 -507 920
rect 267 -920 2107 920
rect 2881 -920 4721 920
<< metal4 >>
rect -5161 1053 -2681 1120
rect -5161 1000 -2831 1053
rect -5161 -1000 -5041 1000
rect -3041 -1000 -2831 1000
rect -5161 -1053 -2831 -1000
rect -2743 -1053 -2681 1053
rect -5161 -1120 -2681 -1053
rect -2547 1053 -67 1120
rect -2547 1000 -217 1053
rect -2547 -1000 -2427 1000
rect -427 -1000 -217 1000
rect -2547 -1053 -217 -1000
rect -129 -1053 -67 1053
rect -2547 -1120 -67 -1053
rect 67 1053 2547 1120
rect 67 1000 2397 1053
rect 67 -1000 187 1000
rect 2187 -1000 2397 1000
rect 67 -1053 2397 -1000
rect 2485 -1053 2547 1053
rect 67 -1120 2547 -1053
rect 2681 1053 5161 1120
rect 2681 1000 5011 1053
rect 2681 -1000 2801 1000
rect 4801 -1000 5011 1000
rect 2681 -1053 5011 -1000
rect 5099 -1053 5161 1053
rect 2681 -1120 5161 -1053
<< via4 >>
rect -2831 -1053 -2743 1053
rect -217 -1053 -129 1053
rect 2397 -1053 2485 1053
rect 5011 -1053 5099 1053
<< metal5 >>
rect -2831 1053 -2743 1063
rect -217 1053 -129 1063
rect -2831 -1063 -2743 -1053
rect 2397 1053 2485 1063
rect -217 -1063 -129 -1053
rect 5011 1053 5099 1063
rect 2397 -1063 2485 -1053
rect 5011 -1063 5099 -1053
<< properties >>
string FIXED_BBOX 2681 -1120 4921 1120
string gencell mim_2p0fF
string library gf180mcu
string parameters w 10 l 10 val 3.3k carea 25.00 cperi 20.00 nx 4 ny 1 dummy 0 square 0 lmin 5.00 wmin 5.00 lmax 100.0 wmax 100.0 dc 0 bconnect 1 tconnect 1
<< end >>
