* NGSPICE file created from Inverter_Layout_flat.ext - technology: gf180mcuC

.subckt Inverter_Layout_flat IN OUT VSS VDD
X0 OUT IN.t0 VDD.t1 VDD.t0 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X1 OUT IN.t1 VSS.t1 VSS.t0 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
R0 IN.n0 IN.t0 34.6755
R1 IN IN.n0 17.6692
R2 IN.n0 IN.t1 13.0362
R3 VDD.n1 VDD.t0 611.386
R4 VDD.n3 VDD.t1 4.7942
R5 VDD.n5 VDD.n4 3.1505
R6 VDD VDD.n2 1.6259
R7 VDD.n2 VDD.n1 1.58417
R8 VDD.n1 VDD.n0 0.684132
R9 VDD VDD.n5 0.0382679
R10 VDD.n5 VDD.n3 0.0270179
R11 OUT.n2 OUT.n1 6.88041
R12 OUT.n2 OUT.n0 4.70224
R13 OUT OUT.n2 0.115935
R14 VSS.n3 VSS.t0 1496.29
R15 VSS.n2 VSS.n1 9.13939
R16 VSS.n0 VSS.t1 6.68085
R17 VSS.n1 VSS.n0 2.61175
R18 VSS VSS.n4 1.31259
R19 VSS.n4 VSS.n3 1.30969
R20 VSS.n4 VSS.n2 0.50294
R21 VSS VSS.n0 0.0647857
C0 IN OUT 0.0407f
C1 VDD IN 0.162f
C2 VDD OUT 0.145f
.ends

