** sch_path: /home/shahid/GF180Projects/PLL_pakistan2/top/xschem/pex_PLL_13_TB.sch
**.subckt pex_PLL_13_TB
C1 Output1 VSS 100f m=1
C2 Output2 VSS 100f m=1
C3 Output_test VSS 100f m=1
C5 LP_op_test VSS 100f m=1
C4 net1 VSS 80.14p m=1
C6 LP_ext VSS 3.77p m=1
R2 LP_ext net1 48.84k m=1
V1 P1 VSS 0
.save i(v1)
V14 P0 VSS 0
.save i(v14)
VCNTL Vref VSS pulse(3.3 0 0 100p 100p 250n 500n)
.save i(vcntl)
V23 VDD_VCO VSS PWL( 0 0 100n 0 100.001n 3.3)
.save i(v23)
V27 VDD VSS 3.3
.save i(v27)
V28 VSS GND 0
.save i(v28)
V29 RST_DIV VSS PWL( 0 0 10n 0 10.001n 3)
.save i(v29)
V30 F1 VSS 3.3
.save i(v30)
V31 F0 VSS 3.3
.save i(v31)
V32 F2 VSS 3.3
.save i(v32)
V33 OPA0 VSS 3.3
.save i(v33)
V34 OPA1 VSS 3.3
.save i(v34)
V35 OPB0 VSS 3.3
.save i(v35)
V36 OPB1 VSS 0
.save i(v36)
I3 VDD Iref 100u
V37 S1 VSS 3.3
.save i(v37)
V38 S0 VSS 3.3
.save i(v38)
V39 S2 VSS 0
.save i(v39)
V40 T1 VSS 0
.save i(v40)
V41 T0 VSS 0
.save i(v41)
V42 vcntl_test VSS 1.08
.save i(v42)
V43 Vo_test VSS PWL( 0 0 10n 0 10.001n 3)
.save i(v43)
V44 Vdiv_test VSS pulse(3.3 0 20n 100p 100p 50n 100n)
.save i(v44)
V45 PU_test VSS pulse(3.3 0 50n 100p 100p 75n 100n)
.save i(v45)
V46 PD_test VSS pulse(3.3 0 0 100p 100p 75n 100n)
.save i(v46)
V2 VDD_BUFF VSS 3.3
.save i(v2)
x1 Iref LP_ext VDD_BUFF VDD VDD_VCO VSS RST_DIV Vref S2 T0 S0 S1 F2 F0 T1 F1 OPA1 OPA0 OPB1 P1 OPB0
+ P0 Vo_test PD_test vcntl_test PU_test Vdiv_test Output1 Output2 Output_test LP_op_test pex_pll_13_mag
**** begin user architecture code


.include pex_pll_13_mag.spice
.control
save F2  F1  LP_op_test  Vref  Output1  Output2  RST_DIV  x1.pu_mux_op_int.t4  x1.pu_int.t9
+  x1.pu_test.n0  x1.pd_int.t11  x1.vco_op_bar.t6  x1.vco_op.t39  x1.vdiv_fb_mux_int.n33  x1.vdiv_fb_mux_int.n33
+  x1.pfd_vref_in_int.t3  x1.pfd_vdiv_in_int.t4

tran 20n 45u
plot v(Output_test) v(LP_op_test)+4
plot v(Output1) v(Output1B)+4 v(Output2)+8
plot v(Vref)
write pex_PLL_13_TB.raw
.endc




.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice cap_mim
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice moscap_typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice mimcap_typical
* .lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_statistical

**** end user architecture code
**.ends
.GLOBAL GND
.end
