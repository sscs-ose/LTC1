magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1955 1019 1955
<< metal1 >>
rect -19 949 19 955
rect -19 -949 -13 949
rect 13 -949 19 949
rect -19 -955 19 -949
<< via1 >>
rect -13 -949 13 949
<< metal2 >>
rect -19 949 19 955
rect -19 -949 -13 949
rect 13 -949 19 949
rect -19 -955 19 -949
<< end >>
