* NGSPICE file created from GF_INV_MAG_flat.ext - technology: gf180mcuC

.subckt GF_INV_MAG_flat VDD VSS IN OUT
X0 OUT IN.t0 VDD.t1 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1 OUT IN.t1 VSS.t1 VSS.t0 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
R0 IN.n0 IN.t0 25.2177
R1 IN.n0 IN.t1 14.6587
R2 IN IN.n0 4.20675
R3 VDD.n0 VDD.t0 483.349
R4 VDD VDD.n0 6.3005
R5 VDD VDD.n0 6.3005
R6 VDD VDD.t1 5.16454
R7 OUT.n2 OUT.n1 9.33985
R8 OUT.n2 OUT.n0 5.17836
R9 OUT OUT.n2 0.115328
R10 VSS.n1 VSS.t0 1249.51
R11 VSS.n2 VSS.t1 9.3736
R12 VSS.n2 VSS.n1 2.6005
R13 VSS.n1 VSS.n0 0.194944
R14 VSS VSS.n2 0.00219811
C0 IN OUT 0.101f
C1 VDD IN 0.195f
C2 VDD OUT 0.152f
.ends

