magic
tech gf180mcuC
magscale 1 10
timestamp 1690200015
<< nwell >>
rect 38 813 846 891
rect 1398 813 2206 891
rect 38 424 1250 813
rect 1398 424 3508 813
rect 846 391 1250 424
rect 2206 391 3508 424
rect 846 372 1050 391
rect 2206 372 2410 391
rect 2610 372 2904 391
rect 3104 372 3308 391
rect 38 -126 846 -48
rect 38 -515 1250 -126
rect 846 -548 1250 -515
rect 1371 -548 2179 -126
rect 2503 -548 3311 -126
rect 846 -567 1050 -548
rect 1371 -567 1575 -548
rect 1775 -567 1979 -548
rect 2503 -567 2707 -548
rect 2907 -567 3111 -548
rect 38 -1009 1734 -988
rect 38 -1087 2459 -1009
rect 38 -1456 3682 -1087
rect 1166 -1476 3682 -1456
rect 1166 -1509 1570 -1476
rect 2459 -1509 3682 -1476
rect 1166 -1528 1370 -1509
rect 2459 -1528 2663 -1509
rect 2863 -1528 3078 -1509
rect 3278 -1528 3482 -1509
rect 38 -2024 846 -1946
rect 1249 -2024 2859 -1946
rect 38 -2045 2859 -2024
rect 38 -2413 3678 -2045
rect 846 -2414 3678 -2413
rect 846 -2446 1250 -2414
rect 846 -2465 1050 -2446
rect 2455 -2467 3678 -2414
rect 2455 -2486 2659 -2467
rect 2859 -2486 3074 -2467
rect 3274 -2486 3478 -2467
rect 38 -3005 1590 -2906
rect 38 -3374 2389 -3005
rect 1166 -3427 2389 -3374
rect 1166 -3446 1370 -3427
rect 1581 -3446 1785 -3427
rect 1985 -3446 2189 -3427
rect 38 -4336 3142 -3868
rect 1166 -4389 1570 -4336
rect 2738 -4389 3142 -4336
rect 3303 -4389 4111 -3967
rect 1166 -4408 1370 -4389
rect 2738 -4408 2942 -4389
rect 3303 -4408 3507 -4389
rect 3707 -4408 3911 -4389
<< pwell >>
rect 100 147 784 383
rect 904 148 1192 346
rect 1460 147 2144 383
rect 2264 148 2552 346
rect 2758 148 3046 346
rect 3162 148 3450 346
rect 100 -792 784 -556
rect 904 -791 1192 -593
rect 1429 -791 1717 -593
rect 1833 -791 2121 -593
rect 2561 -791 2849 -593
rect 2965 -791 3253 -593
rect 256 -1750 948 -1552
rect 1224 -1752 1512 -1554
rect 1713 -1753 2397 -1517
rect 2517 -1752 2805 -1554
rect 2932 -1752 3220 -1554
rect 3336 -1752 3624 -1554
rect 100 -2690 784 -2454
rect 904 -2689 1192 -2491
rect 1545 -2708 2237 -2510
rect 2513 -2710 2801 -2512
rect 2928 -2710 3216 -2512
rect 3332 -2710 3620 -2512
rect 256 -3668 948 -3470
rect 1224 -3670 1512 -3472
rect 1639 -3670 1927 -3472
rect 2043 -3670 2331 -3472
rect 256 -4630 948 -4432
rect 1224 -4632 1512 -4434
rect 1828 -4630 2520 -4432
rect 2796 -4632 3084 -4434
rect 3361 -4632 3649 -4434
rect 3765 -4632 4053 -4434
<< nmos >>
rect 212 215 268 315
rect 616 215 672 315
rect 1020 222 1076 272
rect 1572 215 1628 315
rect 1976 215 2032 315
rect 2380 222 2436 272
rect 2874 222 2930 272
rect 3278 222 3334 272
rect 212 -724 268 -624
rect 616 -724 672 -624
rect 1020 -717 1076 -667
rect 1545 -717 1601 -667
rect 1949 -717 2005 -667
rect 2677 -717 2733 -667
rect 3081 -717 3137 -667
rect 372 -1676 428 -1626
rect 776 -1676 832 -1626
rect 1340 -1678 1396 -1628
rect 1825 -1685 1881 -1585
rect 2229 -1685 2285 -1585
rect 2633 -1678 2689 -1628
rect 3048 -1678 3104 -1628
rect 3452 -1678 3508 -1628
rect 212 -2622 268 -2522
rect 616 -2622 672 -2522
rect 1020 -2615 1076 -2565
rect 1661 -2634 1717 -2584
rect 2065 -2634 2121 -2584
rect 2629 -2636 2685 -2586
rect 3044 -2636 3100 -2586
rect 3448 -2636 3504 -2586
rect 372 -3594 428 -3544
rect 776 -3594 832 -3544
rect 1340 -3596 1396 -3546
rect 1755 -3596 1811 -3546
rect 2159 -3596 2215 -3546
rect 372 -4556 428 -4506
rect 776 -4556 832 -4506
rect 1340 -4558 1396 -4508
rect 1944 -4556 2000 -4506
rect 2348 -4556 2404 -4506
rect 2912 -4558 2968 -4508
rect 3477 -4558 3533 -4508
rect 3881 -4558 3937 -4508
<< pmos >>
rect 212 554 268 654
rect 616 554 672 654
rect 1020 521 1076 621
rect 1572 554 1628 654
rect 1976 554 2032 654
rect 2380 521 2436 621
rect 2874 521 2930 621
rect 3278 521 3334 621
rect 212 -385 268 -285
rect 616 -385 672 -285
rect 1020 -418 1076 -318
rect 1545 -418 1601 -318
rect 1949 -418 2005 -318
rect 2677 -418 2733 -318
rect 3081 -418 3137 -318
rect 212 -1326 268 -1226
rect 372 -1326 428 -1226
rect 776 -1326 832 -1226
rect 936 -1326 992 -1226
rect 1340 -1379 1396 -1279
rect 1825 -1346 1881 -1246
rect 2229 -1346 2285 -1246
rect 2633 -1379 2689 -1279
rect 3048 -1379 3104 -1279
rect 3452 -1379 3508 -1279
rect 212 -2283 268 -2183
rect 616 -2283 672 -2183
rect 1020 -2316 1076 -2216
rect 1501 -2284 1557 -2184
rect 1661 -2284 1717 -2184
rect 2065 -2284 2121 -2184
rect 2225 -2284 2281 -2184
rect 2629 -2337 2685 -2237
rect 3044 -2337 3100 -2237
rect 3448 -2337 3504 -2237
rect 212 -3244 268 -3144
rect 372 -3244 428 -3144
rect 776 -3244 832 -3144
rect 936 -3244 992 -3144
rect 1340 -3297 1396 -3197
rect 1755 -3297 1811 -3197
rect 2159 -3297 2215 -3197
rect 212 -4206 268 -4106
rect 372 -4206 428 -4106
rect 776 -4206 832 -4106
rect 936 -4206 992 -4106
rect 1340 -4259 1396 -4159
rect 1784 -4206 1840 -4106
rect 1944 -4206 2000 -4106
rect 2348 -4206 2404 -4106
rect 2508 -4206 2564 -4106
rect 2912 -4259 2968 -4159
rect 3477 -4259 3533 -4159
rect 3881 -4259 3937 -4159
<< ndiff >>
rect 124 302 212 315
rect 124 228 137 302
rect 183 228 212 302
rect 124 215 212 228
rect 268 302 356 315
rect 268 228 297 302
rect 343 228 356 302
rect 268 215 356 228
rect 528 302 616 315
rect 528 228 541 302
rect 587 228 616 302
rect 528 215 616 228
rect 672 302 760 315
rect 672 228 701 302
rect 747 228 760 302
rect 672 215 760 228
rect 928 272 1000 283
rect 1484 302 1572 315
rect 1096 272 1168 283
rect 928 270 1020 272
rect 928 224 941 270
rect 987 224 1020 270
rect 928 222 1020 224
rect 1076 270 1168 272
rect 1076 224 1109 270
rect 1155 224 1168 270
rect 1076 222 1168 224
rect 928 211 1000 222
rect 1096 211 1168 222
rect 1484 228 1497 302
rect 1543 228 1572 302
rect 1484 215 1572 228
rect 1628 302 1716 315
rect 1628 228 1657 302
rect 1703 228 1716 302
rect 1628 215 1716 228
rect 1888 302 1976 315
rect 1888 228 1901 302
rect 1947 228 1976 302
rect 1888 215 1976 228
rect 2032 302 2120 315
rect 2032 228 2061 302
rect 2107 228 2120 302
rect 2032 215 2120 228
rect 2288 272 2360 283
rect 2456 272 2528 283
rect 2288 270 2380 272
rect 2288 224 2301 270
rect 2347 224 2380 270
rect 2288 222 2380 224
rect 2436 270 2528 272
rect 2436 224 2469 270
rect 2515 224 2528 270
rect 2436 222 2528 224
rect 2288 211 2360 222
rect 2456 211 2528 222
rect 2782 272 2854 283
rect 2950 272 3022 283
rect 2782 270 2874 272
rect 2782 224 2795 270
rect 2841 224 2874 270
rect 2782 222 2874 224
rect 2930 270 3022 272
rect 2930 224 2963 270
rect 3009 224 3022 270
rect 2930 222 3022 224
rect 2782 211 2854 222
rect 2950 211 3022 222
rect 3186 272 3258 283
rect 3354 272 3426 283
rect 3186 270 3278 272
rect 3186 224 3199 270
rect 3245 224 3278 270
rect 3186 222 3278 224
rect 3334 270 3426 272
rect 3334 224 3367 270
rect 3413 224 3426 270
rect 3334 222 3426 224
rect 3186 211 3258 222
rect 3354 211 3426 222
rect 124 -637 212 -624
rect 124 -711 137 -637
rect 183 -711 212 -637
rect 124 -724 212 -711
rect 268 -637 356 -624
rect 268 -711 297 -637
rect 343 -711 356 -637
rect 268 -724 356 -711
rect 528 -637 616 -624
rect 528 -711 541 -637
rect 587 -711 616 -637
rect 528 -724 616 -711
rect 672 -637 760 -624
rect 672 -711 701 -637
rect 747 -711 760 -637
rect 672 -724 760 -711
rect 928 -667 1000 -656
rect 1096 -667 1168 -656
rect 928 -669 1020 -667
rect 928 -715 941 -669
rect 987 -715 1020 -669
rect 928 -717 1020 -715
rect 1076 -669 1168 -667
rect 1076 -715 1109 -669
rect 1155 -715 1168 -669
rect 1076 -717 1168 -715
rect 928 -728 1000 -717
rect 1096 -728 1168 -717
rect 1453 -667 1525 -656
rect 1621 -667 1693 -656
rect 1453 -669 1545 -667
rect 1453 -715 1466 -669
rect 1512 -715 1545 -669
rect 1453 -717 1545 -715
rect 1601 -669 1693 -667
rect 1601 -715 1634 -669
rect 1680 -715 1693 -669
rect 1601 -717 1693 -715
rect 1453 -728 1525 -717
rect 1621 -728 1693 -717
rect 1857 -667 1929 -656
rect 2025 -667 2097 -656
rect 1857 -669 1949 -667
rect 1857 -715 1870 -669
rect 1916 -715 1949 -669
rect 1857 -717 1949 -715
rect 2005 -669 2097 -667
rect 2005 -715 2038 -669
rect 2084 -715 2097 -669
rect 2005 -717 2097 -715
rect 1857 -728 1929 -717
rect 2025 -728 2097 -717
rect 2585 -667 2657 -656
rect 2753 -667 2825 -656
rect 2585 -669 2677 -667
rect 2585 -715 2598 -669
rect 2644 -715 2677 -669
rect 2585 -717 2677 -715
rect 2733 -669 2825 -667
rect 2733 -715 2766 -669
rect 2812 -715 2825 -669
rect 2733 -717 2825 -715
rect 2585 -728 2657 -717
rect 2753 -728 2825 -717
rect 2989 -667 3061 -656
rect 3157 -667 3229 -656
rect 2989 -669 3081 -667
rect 2989 -715 3002 -669
rect 3048 -715 3081 -669
rect 2989 -717 3081 -715
rect 3137 -669 3229 -667
rect 3137 -715 3170 -669
rect 3216 -715 3229 -669
rect 3137 -717 3229 -715
rect 2989 -728 3061 -717
rect 3157 -728 3229 -717
rect 280 -1626 352 -1615
rect 448 -1626 520 -1615
rect 280 -1628 372 -1626
rect 280 -1674 293 -1628
rect 339 -1674 372 -1628
rect 280 -1676 372 -1674
rect 428 -1628 520 -1626
rect 428 -1674 461 -1628
rect 507 -1674 520 -1628
rect 428 -1676 520 -1674
rect 280 -1687 352 -1676
rect 448 -1687 520 -1676
rect 684 -1626 756 -1615
rect 852 -1626 924 -1615
rect 684 -1628 776 -1626
rect 684 -1674 697 -1628
rect 743 -1674 776 -1628
rect 684 -1676 776 -1674
rect 832 -1628 924 -1626
rect 832 -1674 865 -1628
rect 911 -1674 924 -1628
rect 832 -1676 924 -1674
rect 684 -1687 756 -1676
rect 852 -1687 924 -1676
rect 1248 -1628 1320 -1617
rect 1737 -1598 1825 -1585
rect 1416 -1628 1488 -1617
rect 1248 -1630 1340 -1628
rect 1248 -1676 1261 -1630
rect 1307 -1676 1340 -1630
rect 1248 -1678 1340 -1676
rect 1396 -1630 1488 -1628
rect 1396 -1676 1429 -1630
rect 1475 -1676 1488 -1630
rect 1396 -1678 1488 -1676
rect 1248 -1689 1320 -1678
rect 1416 -1689 1488 -1678
rect 1737 -1672 1750 -1598
rect 1796 -1672 1825 -1598
rect 1737 -1685 1825 -1672
rect 1881 -1598 1969 -1585
rect 1881 -1672 1910 -1598
rect 1956 -1672 1969 -1598
rect 1881 -1685 1969 -1672
rect 2141 -1598 2229 -1585
rect 2141 -1672 2154 -1598
rect 2200 -1672 2229 -1598
rect 2141 -1685 2229 -1672
rect 2285 -1598 2373 -1585
rect 2285 -1672 2314 -1598
rect 2360 -1672 2373 -1598
rect 2285 -1685 2373 -1672
rect 2541 -1628 2613 -1617
rect 2709 -1628 2781 -1617
rect 2541 -1630 2633 -1628
rect 2541 -1676 2554 -1630
rect 2600 -1676 2633 -1630
rect 2541 -1678 2633 -1676
rect 2689 -1630 2781 -1628
rect 2689 -1676 2722 -1630
rect 2768 -1676 2781 -1630
rect 2689 -1678 2781 -1676
rect 2541 -1689 2613 -1678
rect 2709 -1689 2781 -1678
rect 2956 -1628 3028 -1617
rect 3124 -1628 3196 -1617
rect 2956 -1630 3048 -1628
rect 2956 -1676 2969 -1630
rect 3015 -1676 3048 -1630
rect 2956 -1678 3048 -1676
rect 3104 -1630 3196 -1628
rect 3104 -1676 3137 -1630
rect 3183 -1676 3196 -1630
rect 3104 -1678 3196 -1676
rect 2956 -1689 3028 -1678
rect 3124 -1689 3196 -1678
rect 3360 -1628 3432 -1617
rect 3528 -1628 3600 -1617
rect 3360 -1630 3452 -1628
rect 3360 -1676 3373 -1630
rect 3419 -1676 3452 -1630
rect 3360 -1678 3452 -1676
rect 3508 -1630 3600 -1628
rect 3508 -1676 3541 -1630
rect 3587 -1676 3600 -1630
rect 3508 -1678 3600 -1676
rect 3360 -1689 3432 -1678
rect 3528 -1689 3600 -1678
rect 124 -2535 212 -2522
rect 124 -2609 137 -2535
rect 183 -2609 212 -2535
rect 124 -2622 212 -2609
rect 268 -2535 356 -2522
rect 268 -2609 297 -2535
rect 343 -2609 356 -2535
rect 268 -2622 356 -2609
rect 528 -2535 616 -2522
rect 528 -2609 541 -2535
rect 587 -2609 616 -2535
rect 528 -2622 616 -2609
rect 672 -2535 760 -2522
rect 672 -2609 701 -2535
rect 747 -2609 760 -2535
rect 672 -2622 760 -2609
rect 928 -2565 1000 -2554
rect 1096 -2565 1168 -2554
rect 928 -2567 1020 -2565
rect 928 -2613 941 -2567
rect 987 -2613 1020 -2567
rect 928 -2615 1020 -2613
rect 1076 -2567 1168 -2565
rect 1076 -2613 1109 -2567
rect 1155 -2613 1168 -2567
rect 1076 -2615 1168 -2613
rect 928 -2626 1000 -2615
rect 1096 -2626 1168 -2615
rect 1569 -2584 1641 -2573
rect 1737 -2584 1809 -2573
rect 1569 -2586 1661 -2584
rect 1569 -2632 1582 -2586
rect 1628 -2632 1661 -2586
rect 1569 -2634 1661 -2632
rect 1717 -2586 1809 -2584
rect 1717 -2632 1750 -2586
rect 1796 -2632 1809 -2586
rect 1717 -2634 1809 -2632
rect 1569 -2645 1641 -2634
rect 1737 -2645 1809 -2634
rect 1973 -2584 2045 -2573
rect 2141 -2584 2213 -2573
rect 1973 -2586 2065 -2584
rect 1973 -2632 1986 -2586
rect 2032 -2632 2065 -2586
rect 1973 -2634 2065 -2632
rect 2121 -2586 2213 -2584
rect 2121 -2632 2154 -2586
rect 2200 -2632 2213 -2586
rect 2121 -2634 2213 -2632
rect 1973 -2645 2045 -2634
rect 2141 -2645 2213 -2634
rect 2537 -2586 2609 -2575
rect 2705 -2586 2777 -2575
rect 2537 -2588 2629 -2586
rect 2537 -2634 2550 -2588
rect 2596 -2634 2629 -2588
rect 2537 -2636 2629 -2634
rect 2685 -2588 2777 -2586
rect 2685 -2634 2718 -2588
rect 2764 -2634 2777 -2588
rect 2685 -2636 2777 -2634
rect 2537 -2647 2609 -2636
rect 2705 -2647 2777 -2636
rect 2952 -2586 3024 -2575
rect 3120 -2586 3192 -2575
rect 2952 -2588 3044 -2586
rect 2952 -2634 2965 -2588
rect 3011 -2634 3044 -2588
rect 2952 -2636 3044 -2634
rect 3100 -2588 3192 -2586
rect 3100 -2634 3133 -2588
rect 3179 -2634 3192 -2588
rect 3100 -2636 3192 -2634
rect 2952 -2647 3024 -2636
rect 3120 -2647 3192 -2636
rect 3356 -2586 3428 -2575
rect 3524 -2586 3596 -2575
rect 3356 -2588 3448 -2586
rect 3356 -2634 3369 -2588
rect 3415 -2634 3448 -2588
rect 3356 -2636 3448 -2634
rect 3504 -2588 3596 -2586
rect 3504 -2634 3537 -2588
rect 3583 -2634 3596 -2588
rect 3504 -2636 3596 -2634
rect 3356 -2647 3428 -2636
rect 3524 -2647 3596 -2636
rect 280 -3544 352 -3533
rect 448 -3544 520 -3533
rect 280 -3546 372 -3544
rect 280 -3592 293 -3546
rect 339 -3592 372 -3546
rect 280 -3594 372 -3592
rect 428 -3546 520 -3544
rect 428 -3592 461 -3546
rect 507 -3592 520 -3546
rect 428 -3594 520 -3592
rect 280 -3605 352 -3594
rect 448 -3605 520 -3594
rect 684 -3544 756 -3533
rect 852 -3544 924 -3533
rect 684 -3546 776 -3544
rect 684 -3592 697 -3546
rect 743 -3592 776 -3546
rect 684 -3594 776 -3592
rect 832 -3546 924 -3544
rect 832 -3592 865 -3546
rect 911 -3592 924 -3546
rect 832 -3594 924 -3592
rect 684 -3605 756 -3594
rect 852 -3605 924 -3594
rect 1248 -3546 1320 -3535
rect 1416 -3546 1488 -3535
rect 1248 -3548 1340 -3546
rect 1248 -3594 1261 -3548
rect 1307 -3594 1340 -3548
rect 1248 -3596 1340 -3594
rect 1396 -3548 1488 -3546
rect 1396 -3594 1429 -3548
rect 1475 -3594 1488 -3548
rect 1396 -3596 1488 -3594
rect 1248 -3607 1320 -3596
rect 1416 -3607 1488 -3596
rect 1663 -3546 1735 -3535
rect 1831 -3546 1903 -3535
rect 1663 -3548 1755 -3546
rect 1663 -3594 1676 -3548
rect 1722 -3594 1755 -3548
rect 1663 -3596 1755 -3594
rect 1811 -3548 1903 -3546
rect 1811 -3594 1844 -3548
rect 1890 -3594 1903 -3548
rect 1811 -3596 1903 -3594
rect 1663 -3607 1735 -3596
rect 1831 -3607 1903 -3596
rect 2067 -3546 2139 -3535
rect 2235 -3546 2307 -3535
rect 2067 -3548 2159 -3546
rect 2067 -3594 2080 -3548
rect 2126 -3594 2159 -3548
rect 2067 -3596 2159 -3594
rect 2215 -3548 2307 -3546
rect 2215 -3594 2248 -3548
rect 2294 -3594 2307 -3548
rect 2215 -3596 2307 -3594
rect 2067 -3607 2139 -3596
rect 2235 -3607 2307 -3596
rect 280 -4506 352 -4495
rect 448 -4506 520 -4495
rect 280 -4508 372 -4506
rect 280 -4554 293 -4508
rect 339 -4554 372 -4508
rect 280 -4556 372 -4554
rect 428 -4508 520 -4506
rect 428 -4554 461 -4508
rect 507 -4554 520 -4508
rect 428 -4556 520 -4554
rect 280 -4567 352 -4556
rect 448 -4567 520 -4556
rect 684 -4506 756 -4495
rect 852 -4506 924 -4495
rect 684 -4508 776 -4506
rect 684 -4554 697 -4508
rect 743 -4554 776 -4508
rect 684 -4556 776 -4554
rect 832 -4508 924 -4506
rect 832 -4554 865 -4508
rect 911 -4554 924 -4508
rect 832 -4556 924 -4554
rect 684 -4567 756 -4556
rect 852 -4567 924 -4556
rect 1248 -4508 1320 -4497
rect 1416 -4508 1488 -4497
rect 1248 -4510 1340 -4508
rect 1248 -4556 1261 -4510
rect 1307 -4556 1340 -4510
rect 1248 -4558 1340 -4556
rect 1396 -4510 1488 -4508
rect 1396 -4556 1429 -4510
rect 1475 -4556 1488 -4510
rect 1396 -4558 1488 -4556
rect 1248 -4569 1320 -4558
rect 1416 -4569 1488 -4558
rect 1852 -4506 1924 -4495
rect 2020 -4506 2092 -4495
rect 1852 -4508 1944 -4506
rect 1852 -4554 1865 -4508
rect 1911 -4554 1944 -4508
rect 1852 -4556 1944 -4554
rect 2000 -4508 2092 -4506
rect 2000 -4554 2033 -4508
rect 2079 -4554 2092 -4508
rect 2000 -4556 2092 -4554
rect 1852 -4567 1924 -4556
rect 2020 -4567 2092 -4556
rect 2256 -4506 2328 -4495
rect 2424 -4506 2496 -4495
rect 2256 -4508 2348 -4506
rect 2256 -4554 2269 -4508
rect 2315 -4554 2348 -4508
rect 2256 -4556 2348 -4554
rect 2404 -4508 2496 -4506
rect 2404 -4554 2437 -4508
rect 2483 -4554 2496 -4508
rect 2404 -4556 2496 -4554
rect 2256 -4567 2328 -4556
rect 2424 -4567 2496 -4556
rect 2820 -4508 2892 -4497
rect 2988 -4508 3060 -4497
rect 2820 -4510 2912 -4508
rect 2820 -4556 2833 -4510
rect 2879 -4556 2912 -4510
rect 2820 -4558 2912 -4556
rect 2968 -4510 3060 -4508
rect 2968 -4556 3001 -4510
rect 3047 -4556 3060 -4510
rect 2968 -4558 3060 -4556
rect 2820 -4569 2892 -4558
rect 2988 -4569 3060 -4558
rect 3385 -4508 3457 -4497
rect 3553 -4508 3625 -4497
rect 3385 -4510 3477 -4508
rect 3385 -4556 3398 -4510
rect 3444 -4556 3477 -4510
rect 3385 -4558 3477 -4556
rect 3533 -4510 3625 -4508
rect 3533 -4556 3566 -4510
rect 3612 -4556 3625 -4510
rect 3533 -4558 3625 -4556
rect 3385 -4569 3457 -4558
rect 3553 -4569 3625 -4558
rect 3789 -4508 3861 -4497
rect 3957 -4508 4029 -4497
rect 3789 -4510 3881 -4508
rect 3789 -4556 3802 -4510
rect 3848 -4556 3881 -4510
rect 3789 -4558 3881 -4556
rect 3937 -4510 4029 -4508
rect 3937 -4556 3970 -4510
rect 4016 -4556 4029 -4510
rect 3937 -4558 4029 -4556
rect 3789 -4569 3861 -4558
rect 3957 -4569 4029 -4558
<< pdiff >>
rect 124 641 212 654
rect 124 567 137 641
rect 183 567 212 641
rect 124 554 212 567
rect 268 641 356 654
rect 268 567 297 641
rect 343 567 356 641
rect 268 554 356 567
rect 528 641 616 654
rect 528 567 541 641
rect 587 567 616 641
rect 528 554 616 567
rect 672 641 760 654
rect 672 567 701 641
rect 747 567 760 641
rect 1484 641 1572 654
rect 672 554 760 567
rect 932 608 1020 621
rect 932 534 945 608
rect 991 534 1020 608
rect 932 521 1020 534
rect 1076 608 1164 621
rect 1076 534 1105 608
rect 1151 534 1164 608
rect 1076 521 1164 534
rect 1484 567 1497 641
rect 1543 567 1572 641
rect 1484 554 1572 567
rect 1628 641 1716 654
rect 1628 567 1657 641
rect 1703 567 1716 641
rect 1628 554 1716 567
rect 1888 641 1976 654
rect 1888 567 1901 641
rect 1947 567 1976 641
rect 1888 554 1976 567
rect 2032 641 2120 654
rect 2032 567 2061 641
rect 2107 567 2120 641
rect 2032 554 2120 567
rect 2292 608 2380 621
rect 2292 534 2305 608
rect 2351 534 2380 608
rect 2292 521 2380 534
rect 2436 608 2524 621
rect 2436 534 2465 608
rect 2511 534 2524 608
rect 2436 521 2524 534
rect 2786 608 2874 621
rect 2786 534 2799 608
rect 2845 534 2874 608
rect 2786 521 2874 534
rect 2930 608 3018 621
rect 2930 534 2959 608
rect 3005 534 3018 608
rect 2930 521 3018 534
rect 3190 608 3278 621
rect 3190 534 3203 608
rect 3249 534 3278 608
rect 3190 521 3278 534
rect 3334 608 3422 621
rect 3334 534 3363 608
rect 3409 534 3422 608
rect 3334 521 3422 534
rect 124 -298 212 -285
rect 124 -372 137 -298
rect 183 -372 212 -298
rect 124 -385 212 -372
rect 268 -298 356 -285
rect 268 -372 297 -298
rect 343 -372 356 -298
rect 268 -385 356 -372
rect 528 -298 616 -285
rect 528 -372 541 -298
rect 587 -372 616 -298
rect 528 -385 616 -372
rect 672 -298 760 -285
rect 672 -372 701 -298
rect 747 -372 760 -298
rect 672 -385 760 -372
rect 932 -331 1020 -318
rect 932 -405 945 -331
rect 991 -405 1020 -331
rect 932 -418 1020 -405
rect 1076 -331 1164 -318
rect 1076 -405 1105 -331
rect 1151 -405 1164 -331
rect 1076 -418 1164 -405
rect 1457 -331 1545 -318
rect 1457 -405 1470 -331
rect 1516 -405 1545 -331
rect 1457 -418 1545 -405
rect 1601 -331 1689 -318
rect 1601 -405 1630 -331
rect 1676 -405 1689 -331
rect 1601 -418 1689 -405
rect 1861 -331 1949 -318
rect 1861 -405 1874 -331
rect 1920 -405 1949 -331
rect 1861 -418 1949 -405
rect 2005 -331 2093 -318
rect 2005 -405 2034 -331
rect 2080 -405 2093 -331
rect 2005 -418 2093 -405
rect 2589 -331 2677 -318
rect 2589 -405 2602 -331
rect 2648 -405 2677 -331
rect 2589 -418 2677 -405
rect 2733 -331 2821 -318
rect 2733 -405 2762 -331
rect 2808 -405 2821 -331
rect 2733 -418 2821 -405
rect 2993 -331 3081 -318
rect 2993 -405 3006 -331
rect 3052 -405 3081 -331
rect 2993 -418 3081 -405
rect 3137 -331 3225 -318
rect 3137 -405 3166 -331
rect 3212 -405 3225 -331
rect 3137 -418 3225 -405
rect 124 -1239 212 -1226
rect 124 -1313 137 -1239
rect 183 -1313 212 -1239
rect 124 -1326 212 -1313
rect 268 -1239 372 -1226
rect 268 -1313 297 -1239
rect 343 -1313 372 -1239
rect 268 -1326 372 -1313
rect 428 -1239 516 -1226
rect 428 -1313 457 -1239
rect 503 -1313 516 -1239
rect 428 -1326 516 -1313
rect 688 -1239 776 -1226
rect 688 -1313 701 -1239
rect 747 -1313 776 -1239
rect 688 -1326 776 -1313
rect 832 -1239 936 -1226
rect 832 -1313 861 -1239
rect 907 -1313 936 -1239
rect 832 -1326 936 -1313
rect 992 -1239 1080 -1226
rect 992 -1313 1021 -1239
rect 1067 -1313 1080 -1239
rect 1737 -1259 1825 -1246
rect 992 -1326 1080 -1313
rect 1252 -1292 1340 -1279
rect 1252 -1366 1265 -1292
rect 1311 -1366 1340 -1292
rect 1252 -1379 1340 -1366
rect 1396 -1292 1484 -1279
rect 1396 -1366 1425 -1292
rect 1471 -1366 1484 -1292
rect 1396 -1379 1484 -1366
rect 1737 -1333 1750 -1259
rect 1796 -1333 1825 -1259
rect 1737 -1346 1825 -1333
rect 1881 -1259 1969 -1246
rect 1881 -1333 1910 -1259
rect 1956 -1333 1969 -1259
rect 1881 -1346 1969 -1333
rect 2141 -1259 2229 -1246
rect 2141 -1333 2154 -1259
rect 2200 -1333 2229 -1259
rect 2141 -1346 2229 -1333
rect 2285 -1259 2373 -1246
rect 2285 -1333 2314 -1259
rect 2360 -1333 2373 -1259
rect 2285 -1346 2373 -1333
rect 2545 -1292 2633 -1279
rect 2545 -1366 2558 -1292
rect 2604 -1366 2633 -1292
rect 2545 -1379 2633 -1366
rect 2689 -1292 2777 -1279
rect 2689 -1366 2718 -1292
rect 2764 -1366 2777 -1292
rect 2689 -1379 2777 -1366
rect 2960 -1292 3048 -1279
rect 2960 -1366 2973 -1292
rect 3019 -1366 3048 -1292
rect 2960 -1379 3048 -1366
rect 3104 -1292 3192 -1279
rect 3104 -1366 3133 -1292
rect 3179 -1366 3192 -1292
rect 3104 -1379 3192 -1366
rect 3364 -1292 3452 -1279
rect 3364 -1366 3377 -1292
rect 3423 -1366 3452 -1292
rect 3364 -1379 3452 -1366
rect 3508 -1292 3596 -1279
rect 3508 -1366 3537 -1292
rect 3583 -1366 3596 -1292
rect 3508 -1379 3596 -1366
rect 124 -2196 212 -2183
rect 124 -2270 137 -2196
rect 183 -2270 212 -2196
rect 124 -2283 212 -2270
rect 268 -2196 356 -2183
rect 268 -2270 297 -2196
rect 343 -2270 356 -2196
rect 268 -2283 356 -2270
rect 528 -2196 616 -2183
rect 528 -2270 541 -2196
rect 587 -2270 616 -2196
rect 528 -2283 616 -2270
rect 672 -2196 760 -2183
rect 672 -2270 701 -2196
rect 747 -2270 760 -2196
rect 1413 -2197 1501 -2184
rect 672 -2283 760 -2270
rect 932 -2229 1020 -2216
rect 932 -2303 945 -2229
rect 991 -2303 1020 -2229
rect 932 -2316 1020 -2303
rect 1076 -2229 1164 -2216
rect 1076 -2303 1105 -2229
rect 1151 -2303 1164 -2229
rect 1413 -2271 1426 -2197
rect 1472 -2271 1501 -2197
rect 1413 -2284 1501 -2271
rect 1557 -2197 1661 -2184
rect 1557 -2271 1586 -2197
rect 1632 -2271 1661 -2197
rect 1557 -2284 1661 -2271
rect 1717 -2197 1805 -2184
rect 1717 -2271 1746 -2197
rect 1792 -2271 1805 -2197
rect 1717 -2284 1805 -2271
rect 1977 -2197 2065 -2184
rect 1977 -2271 1990 -2197
rect 2036 -2271 2065 -2197
rect 1977 -2284 2065 -2271
rect 2121 -2197 2225 -2184
rect 2121 -2271 2150 -2197
rect 2196 -2271 2225 -2197
rect 2121 -2284 2225 -2271
rect 2281 -2197 2369 -2184
rect 2281 -2271 2310 -2197
rect 2356 -2271 2369 -2197
rect 2281 -2284 2369 -2271
rect 2541 -2250 2629 -2237
rect 1076 -2316 1164 -2303
rect 2541 -2324 2554 -2250
rect 2600 -2324 2629 -2250
rect 2541 -2337 2629 -2324
rect 2685 -2250 2773 -2237
rect 2685 -2324 2714 -2250
rect 2760 -2324 2773 -2250
rect 2685 -2337 2773 -2324
rect 2956 -2250 3044 -2237
rect 2956 -2324 2969 -2250
rect 3015 -2324 3044 -2250
rect 2956 -2337 3044 -2324
rect 3100 -2250 3188 -2237
rect 3100 -2324 3129 -2250
rect 3175 -2324 3188 -2250
rect 3100 -2337 3188 -2324
rect 3360 -2250 3448 -2237
rect 3360 -2324 3373 -2250
rect 3419 -2324 3448 -2250
rect 3360 -2337 3448 -2324
rect 3504 -2250 3592 -2237
rect 3504 -2324 3533 -2250
rect 3579 -2324 3592 -2250
rect 3504 -2337 3592 -2324
rect 124 -3157 212 -3144
rect 124 -3231 137 -3157
rect 183 -3231 212 -3157
rect 124 -3244 212 -3231
rect 268 -3157 372 -3144
rect 268 -3231 297 -3157
rect 343 -3231 372 -3157
rect 268 -3244 372 -3231
rect 428 -3157 516 -3144
rect 428 -3231 457 -3157
rect 503 -3231 516 -3157
rect 428 -3244 516 -3231
rect 688 -3157 776 -3144
rect 688 -3231 701 -3157
rect 747 -3231 776 -3157
rect 688 -3244 776 -3231
rect 832 -3157 936 -3144
rect 832 -3231 861 -3157
rect 907 -3231 936 -3157
rect 832 -3244 936 -3231
rect 992 -3157 1080 -3144
rect 992 -3231 1021 -3157
rect 1067 -3231 1080 -3157
rect 992 -3244 1080 -3231
rect 1252 -3210 1340 -3197
rect 1252 -3284 1265 -3210
rect 1311 -3284 1340 -3210
rect 1252 -3297 1340 -3284
rect 1396 -3210 1484 -3197
rect 1396 -3284 1425 -3210
rect 1471 -3284 1484 -3210
rect 1396 -3297 1484 -3284
rect 1667 -3210 1755 -3197
rect 1667 -3284 1680 -3210
rect 1726 -3284 1755 -3210
rect 1667 -3297 1755 -3284
rect 1811 -3210 1899 -3197
rect 1811 -3284 1840 -3210
rect 1886 -3284 1899 -3210
rect 1811 -3297 1899 -3284
rect 2071 -3210 2159 -3197
rect 2071 -3284 2084 -3210
rect 2130 -3284 2159 -3210
rect 2071 -3297 2159 -3284
rect 2215 -3210 2303 -3197
rect 2215 -3284 2244 -3210
rect 2290 -3284 2303 -3210
rect 2215 -3297 2303 -3284
rect 124 -4119 212 -4106
rect 124 -4193 137 -4119
rect 183 -4193 212 -4119
rect 124 -4206 212 -4193
rect 268 -4119 372 -4106
rect 268 -4193 297 -4119
rect 343 -4193 372 -4119
rect 268 -4206 372 -4193
rect 428 -4119 516 -4106
rect 428 -4193 457 -4119
rect 503 -4193 516 -4119
rect 428 -4206 516 -4193
rect 688 -4119 776 -4106
rect 688 -4193 701 -4119
rect 747 -4193 776 -4119
rect 688 -4206 776 -4193
rect 832 -4119 936 -4106
rect 832 -4193 861 -4119
rect 907 -4193 936 -4119
rect 832 -4206 936 -4193
rect 992 -4119 1080 -4106
rect 992 -4193 1021 -4119
rect 1067 -4193 1080 -4119
rect 1696 -4119 1784 -4106
rect 992 -4206 1080 -4193
rect 1252 -4172 1340 -4159
rect 1252 -4246 1265 -4172
rect 1311 -4246 1340 -4172
rect 1252 -4259 1340 -4246
rect 1396 -4172 1484 -4159
rect 1396 -4246 1425 -4172
rect 1471 -4246 1484 -4172
rect 1696 -4193 1709 -4119
rect 1755 -4193 1784 -4119
rect 1696 -4206 1784 -4193
rect 1840 -4119 1944 -4106
rect 1840 -4193 1869 -4119
rect 1915 -4193 1944 -4119
rect 1840 -4206 1944 -4193
rect 2000 -4119 2088 -4106
rect 2000 -4193 2029 -4119
rect 2075 -4193 2088 -4119
rect 2000 -4206 2088 -4193
rect 2260 -4119 2348 -4106
rect 2260 -4193 2273 -4119
rect 2319 -4193 2348 -4119
rect 2260 -4206 2348 -4193
rect 2404 -4119 2508 -4106
rect 2404 -4193 2433 -4119
rect 2479 -4193 2508 -4119
rect 2404 -4206 2508 -4193
rect 2564 -4119 2652 -4106
rect 2564 -4193 2593 -4119
rect 2639 -4193 2652 -4119
rect 2564 -4206 2652 -4193
rect 2824 -4172 2912 -4159
rect 1396 -4259 1484 -4246
rect 2824 -4246 2837 -4172
rect 2883 -4246 2912 -4172
rect 2824 -4259 2912 -4246
rect 2968 -4172 3056 -4159
rect 2968 -4246 2997 -4172
rect 3043 -4246 3056 -4172
rect 2968 -4259 3056 -4246
rect 3389 -4172 3477 -4159
rect 3389 -4246 3402 -4172
rect 3448 -4246 3477 -4172
rect 3389 -4259 3477 -4246
rect 3533 -4172 3621 -4159
rect 3533 -4246 3562 -4172
rect 3608 -4246 3621 -4172
rect 3533 -4259 3621 -4246
rect 3793 -4172 3881 -4159
rect 3793 -4246 3806 -4172
rect 3852 -4246 3881 -4172
rect 3793 -4259 3881 -4246
rect 3937 -4172 4025 -4159
rect 3937 -4246 3966 -4172
rect 4012 -4246 4025 -4172
rect 3937 -4259 4025 -4246
<< ndiffc >>
rect 137 228 183 302
rect 297 228 343 302
rect 541 228 587 302
rect 701 228 747 302
rect 941 224 987 270
rect 1109 224 1155 270
rect 1497 228 1543 302
rect 1657 228 1703 302
rect 1901 228 1947 302
rect 2061 228 2107 302
rect 2301 224 2347 270
rect 2469 224 2515 270
rect 2795 224 2841 270
rect 2963 224 3009 270
rect 3199 224 3245 270
rect 3367 224 3413 270
rect 137 -711 183 -637
rect 297 -711 343 -637
rect 541 -711 587 -637
rect 701 -711 747 -637
rect 941 -715 987 -669
rect 1109 -715 1155 -669
rect 1466 -715 1512 -669
rect 1634 -715 1680 -669
rect 1870 -715 1916 -669
rect 2038 -715 2084 -669
rect 2598 -715 2644 -669
rect 2766 -715 2812 -669
rect 3002 -715 3048 -669
rect 3170 -715 3216 -669
rect 293 -1674 339 -1628
rect 461 -1674 507 -1628
rect 697 -1674 743 -1628
rect 865 -1674 911 -1628
rect 1261 -1676 1307 -1630
rect 1429 -1676 1475 -1630
rect 1750 -1672 1796 -1598
rect 1910 -1672 1956 -1598
rect 2154 -1672 2200 -1598
rect 2314 -1672 2360 -1598
rect 2554 -1676 2600 -1630
rect 2722 -1676 2768 -1630
rect 2969 -1676 3015 -1630
rect 3137 -1676 3183 -1630
rect 3373 -1676 3419 -1630
rect 3541 -1676 3587 -1630
rect 137 -2609 183 -2535
rect 297 -2609 343 -2535
rect 541 -2609 587 -2535
rect 701 -2609 747 -2535
rect 941 -2613 987 -2567
rect 1109 -2613 1155 -2567
rect 1582 -2632 1628 -2586
rect 1750 -2632 1796 -2586
rect 1986 -2632 2032 -2586
rect 2154 -2632 2200 -2586
rect 2550 -2634 2596 -2588
rect 2718 -2634 2764 -2588
rect 2965 -2634 3011 -2588
rect 3133 -2634 3179 -2588
rect 3369 -2634 3415 -2588
rect 3537 -2634 3583 -2588
rect 293 -3592 339 -3546
rect 461 -3592 507 -3546
rect 697 -3592 743 -3546
rect 865 -3592 911 -3546
rect 1261 -3594 1307 -3548
rect 1429 -3594 1475 -3548
rect 1676 -3594 1722 -3548
rect 1844 -3594 1890 -3548
rect 2080 -3594 2126 -3548
rect 2248 -3594 2294 -3548
rect 293 -4554 339 -4508
rect 461 -4554 507 -4508
rect 697 -4554 743 -4508
rect 865 -4554 911 -4508
rect 1261 -4556 1307 -4510
rect 1429 -4556 1475 -4510
rect 1865 -4554 1911 -4508
rect 2033 -4554 2079 -4508
rect 2269 -4554 2315 -4508
rect 2437 -4554 2483 -4508
rect 2833 -4556 2879 -4510
rect 3001 -4556 3047 -4510
rect 3398 -4556 3444 -4510
rect 3566 -4556 3612 -4510
rect 3802 -4556 3848 -4510
rect 3970 -4556 4016 -4510
<< pdiffc >>
rect 137 567 183 641
rect 297 567 343 641
rect 541 567 587 641
rect 701 567 747 641
rect 945 534 991 608
rect 1105 534 1151 608
rect 1497 567 1543 641
rect 1657 567 1703 641
rect 1901 567 1947 641
rect 2061 567 2107 641
rect 2305 534 2351 608
rect 2465 534 2511 608
rect 2799 534 2845 608
rect 2959 534 3005 608
rect 3203 534 3249 608
rect 3363 534 3409 608
rect 137 -372 183 -298
rect 297 -372 343 -298
rect 541 -372 587 -298
rect 701 -372 747 -298
rect 945 -405 991 -331
rect 1105 -405 1151 -331
rect 1470 -405 1516 -331
rect 1630 -405 1676 -331
rect 1874 -405 1920 -331
rect 2034 -405 2080 -331
rect 2602 -405 2648 -331
rect 2762 -405 2808 -331
rect 3006 -405 3052 -331
rect 3166 -405 3212 -331
rect 137 -1313 183 -1239
rect 297 -1313 343 -1239
rect 457 -1313 503 -1239
rect 701 -1313 747 -1239
rect 861 -1313 907 -1239
rect 1021 -1313 1067 -1239
rect 1265 -1366 1311 -1292
rect 1425 -1366 1471 -1292
rect 1750 -1333 1796 -1259
rect 1910 -1333 1956 -1259
rect 2154 -1333 2200 -1259
rect 2314 -1333 2360 -1259
rect 2558 -1366 2604 -1292
rect 2718 -1366 2764 -1292
rect 2973 -1366 3019 -1292
rect 3133 -1366 3179 -1292
rect 3377 -1366 3423 -1292
rect 3537 -1366 3583 -1292
rect 137 -2270 183 -2196
rect 297 -2270 343 -2196
rect 541 -2270 587 -2196
rect 701 -2270 747 -2196
rect 945 -2303 991 -2229
rect 1105 -2303 1151 -2229
rect 1426 -2271 1472 -2197
rect 1586 -2271 1632 -2197
rect 1746 -2271 1792 -2197
rect 1990 -2271 2036 -2197
rect 2150 -2271 2196 -2197
rect 2310 -2271 2356 -2197
rect 2554 -2324 2600 -2250
rect 2714 -2324 2760 -2250
rect 2969 -2324 3015 -2250
rect 3129 -2324 3175 -2250
rect 3373 -2324 3419 -2250
rect 3533 -2324 3579 -2250
rect 137 -3231 183 -3157
rect 297 -3231 343 -3157
rect 457 -3231 503 -3157
rect 701 -3231 747 -3157
rect 861 -3231 907 -3157
rect 1021 -3231 1067 -3157
rect 1265 -3284 1311 -3210
rect 1425 -3284 1471 -3210
rect 1680 -3284 1726 -3210
rect 1840 -3284 1886 -3210
rect 2084 -3284 2130 -3210
rect 2244 -3284 2290 -3210
rect 137 -4193 183 -4119
rect 297 -4193 343 -4119
rect 457 -4193 503 -4119
rect 701 -4193 747 -4119
rect 861 -4193 907 -4119
rect 1021 -4193 1067 -4119
rect 1265 -4246 1311 -4172
rect 1425 -4246 1471 -4172
rect 1709 -4193 1755 -4119
rect 1869 -4193 1915 -4119
rect 2029 -4193 2075 -4119
rect 2273 -4193 2319 -4119
rect 2433 -4193 2479 -4119
rect 2593 -4193 2639 -4119
rect 2837 -4246 2883 -4172
rect 2997 -4246 3043 -4172
rect 3402 -4246 3448 -4172
rect 3562 -4246 3608 -4172
rect 3806 -4246 3852 -4172
rect 3966 -4246 4012 -4172
<< psubdiff >>
rect 64 91 891 97
rect 1424 91 2251 97
rect 64 83 1220 91
rect 64 37 87 83
rect 794 78 1220 83
rect 794 37 891 78
rect 64 29 891 37
rect 1200 29 1220 78
rect 64 24 1220 29
rect 1424 83 2580 91
rect 1424 37 1447 83
rect 2154 78 2580 83
rect 2154 37 2251 78
rect 1424 29 2251 37
rect 2560 29 2580 78
rect 1424 24 2580 29
rect 815 21 1220 24
rect 2175 21 2580 24
rect 872 14 1220 21
rect 2232 14 2580 21
rect 2726 78 3074 91
rect 2726 29 2745 78
rect 3054 29 3074 78
rect 2726 14 3074 29
rect 3130 78 3478 91
rect 3130 29 3149 78
rect 3458 29 3478 78
rect 3130 14 3478 29
rect 64 -848 891 -842
rect 64 -856 1220 -848
rect 64 -902 87 -856
rect 794 -861 1220 -856
rect 794 -902 891 -861
rect 64 -910 891 -902
rect 1200 -910 1220 -861
rect 64 -915 1220 -910
rect 815 -918 1220 -915
rect 872 -925 1220 -918
rect 1397 -861 1745 -848
rect 1397 -910 1416 -861
rect 1725 -910 1745 -861
rect 1397 -925 1745 -910
rect 1801 -861 2149 -848
rect 1801 -910 1820 -861
rect 2129 -910 2149 -861
rect 1801 -925 2149 -910
rect 2529 -861 2877 -848
rect 2529 -910 2548 -861
rect 2857 -910 2877 -861
rect 2529 -925 2877 -910
rect 2933 -861 3281 -848
rect 2933 -910 2952 -861
rect 3261 -910 3281 -861
rect 2933 -925 3281 -910
rect 72 -1822 1115 -1807
rect 1677 -1809 2504 -1803
rect 72 -1868 102 -1822
rect 1086 -1868 1115 -1822
rect 72 -1883 1115 -1868
rect 1192 -1822 1540 -1809
rect 1192 -1871 1211 -1822
rect 1520 -1871 1540 -1822
rect 1192 -1886 1540 -1871
rect 1677 -1817 2833 -1809
rect 1677 -1863 1700 -1817
rect 2407 -1822 2833 -1817
rect 2407 -1863 2504 -1822
rect 1677 -1871 2504 -1863
rect 2813 -1871 2833 -1822
rect 1677 -1876 2833 -1871
rect 2428 -1879 2833 -1876
rect 2485 -1886 2833 -1879
rect 2900 -1822 3248 -1809
rect 2900 -1871 2919 -1822
rect 3228 -1871 3248 -1822
rect 2900 -1886 3248 -1871
rect 3304 -1822 3652 -1809
rect 3304 -1871 3323 -1822
rect 3632 -1871 3652 -1822
rect 3304 -1886 3652 -1871
rect 64 -2746 891 -2740
rect 64 -2754 1220 -2746
rect 64 -2800 87 -2754
rect 794 -2759 1220 -2754
rect 794 -2800 891 -2759
rect 64 -2808 891 -2800
rect 1200 -2808 1220 -2759
rect 64 -2813 1220 -2808
rect 815 -2816 1220 -2813
rect 872 -2823 1220 -2816
rect 1361 -2780 2404 -2765
rect 1361 -2826 1391 -2780
rect 2375 -2826 2404 -2780
rect 1361 -2841 2404 -2826
rect 2481 -2780 2829 -2767
rect 2481 -2829 2500 -2780
rect 2809 -2829 2829 -2780
rect 2481 -2844 2829 -2829
rect 2896 -2780 3244 -2767
rect 2896 -2829 2915 -2780
rect 3224 -2829 3244 -2780
rect 2896 -2844 3244 -2829
rect 3300 -2780 3648 -2767
rect 3300 -2829 3319 -2780
rect 3628 -2829 3648 -2780
rect 3300 -2844 3648 -2829
rect 72 -3740 1115 -3725
rect 72 -3786 102 -3740
rect 1086 -3786 1115 -3740
rect 72 -3801 1115 -3786
rect 1192 -3740 1540 -3727
rect 1192 -3789 1211 -3740
rect 1520 -3789 1540 -3740
rect 1192 -3804 1540 -3789
rect 1607 -3740 1955 -3727
rect 1607 -3789 1626 -3740
rect 1935 -3789 1955 -3740
rect 1607 -3804 1955 -3789
rect 2011 -3740 2359 -3727
rect 2011 -3789 2030 -3740
rect 2339 -3789 2359 -3740
rect 2011 -3804 2359 -3789
rect 72 -4702 1115 -4687
rect 72 -4748 102 -4702
rect 1086 -4748 1115 -4702
rect 72 -4763 1115 -4748
rect 1192 -4702 1540 -4689
rect 1192 -4751 1211 -4702
rect 1520 -4751 1540 -4702
rect 1192 -4766 1540 -4751
rect 1644 -4702 2687 -4687
rect 1644 -4748 1674 -4702
rect 2658 -4748 2687 -4702
rect 1644 -4763 2687 -4748
rect 2764 -4702 3112 -4689
rect 2764 -4751 2783 -4702
rect 3092 -4751 3112 -4702
rect 2764 -4766 3112 -4751
rect 3329 -4702 3677 -4689
rect 3329 -4751 3348 -4702
rect 3657 -4751 3677 -4702
rect 3329 -4766 3677 -4751
rect 3733 -4702 4081 -4689
rect 3733 -4751 3752 -4702
rect 4061 -4751 4081 -4702
rect 3733 -4766 4081 -4751
<< nsubdiff >>
rect 67 851 808 866
rect 67 799 88 851
rect 787 799 808 851
rect 67 782 808 799
rect 1427 851 2168 866
rect 1427 799 1448 851
rect 2147 799 2168 851
rect 886 769 1178 786
rect 1427 782 2168 799
rect 886 718 906 769
rect 1156 718 1178 769
rect 886 701 1178 718
rect 2246 769 2538 786
rect 2246 718 2266 769
rect 2516 718 2538 769
rect 2246 701 2538 718
rect 2740 769 3032 786
rect 2740 718 2760 769
rect 3010 718 3032 769
rect 2740 701 3032 718
rect 3144 769 3436 786
rect 3144 718 3164 769
rect 3414 718 3436 769
rect 3144 701 3436 718
rect 67 -88 808 -73
rect 67 -140 88 -88
rect 787 -140 808 -88
rect 67 -157 808 -140
rect 886 -170 1178 -153
rect 886 -221 906 -170
rect 1156 -221 1178 -170
rect 886 -238 1178 -221
rect 1411 -170 1703 -153
rect 1411 -221 1431 -170
rect 1681 -221 1703 -170
rect 1411 -238 1703 -221
rect 1815 -170 2107 -153
rect 1815 -221 1835 -170
rect 2085 -221 2107 -170
rect 1815 -238 2107 -221
rect 2543 -170 2835 -153
rect 2543 -221 2563 -170
rect 2813 -221 2835 -170
rect 2543 -238 2835 -221
rect 2947 -170 3239 -153
rect 2947 -221 2967 -170
rect 3217 -221 3239 -170
rect 2947 -238 3239 -221
rect 62 -1025 1134 -1012
rect 62 -1072 83 -1025
rect 1105 -1072 1134 -1025
rect 62 -1087 1134 -1072
rect 1680 -1049 2421 -1034
rect 1680 -1101 1701 -1049
rect 2400 -1101 2421 -1049
rect 1206 -1131 1498 -1114
rect 1680 -1118 2421 -1101
rect 1206 -1182 1226 -1131
rect 1476 -1182 1498 -1131
rect 1206 -1199 1498 -1182
rect 2499 -1131 2791 -1114
rect 2499 -1182 2519 -1131
rect 2769 -1182 2791 -1131
rect 2499 -1199 2791 -1182
rect 2914 -1131 3206 -1114
rect 2914 -1182 2934 -1131
rect 3184 -1182 3206 -1131
rect 2914 -1199 3206 -1182
rect 3318 -1131 3610 -1114
rect 3318 -1182 3338 -1131
rect 3588 -1182 3610 -1131
rect 3318 -1199 3610 -1182
rect 67 -1986 808 -1971
rect 67 -2038 88 -1986
rect 787 -2038 808 -1986
rect 67 -2055 808 -2038
rect 1351 -1983 2423 -1970
rect 1351 -2030 1372 -1983
rect 2394 -2030 2423 -1983
rect 1351 -2045 2423 -2030
rect 886 -2068 1178 -2051
rect 886 -2119 906 -2068
rect 1156 -2119 1178 -2068
rect 2495 -2089 2787 -2072
rect 886 -2136 1178 -2119
rect 2495 -2140 2515 -2089
rect 2765 -2140 2787 -2089
rect 2495 -2157 2787 -2140
rect 2910 -2089 3202 -2072
rect 2910 -2140 2930 -2089
rect 3180 -2140 3202 -2089
rect 2910 -2157 3202 -2140
rect 3314 -2089 3606 -2072
rect 3314 -2140 3334 -2089
rect 3584 -2140 3606 -2089
rect 3314 -2157 3606 -2140
rect 62 -2943 1134 -2930
rect 62 -2990 83 -2943
rect 1105 -2990 1134 -2943
rect 62 -3005 1134 -2990
rect 1206 -3049 1498 -3032
rect 1206 -3100 1226 -3049
rect 1476 -3100 1498 -3049
rect 1206 -3117 1498 -3100
rect 1621 -3049 1913 -3032
rect 1621 -3100 1641 -3049
rect 1891 -3100 1913 -3049
rect 1621 -3117 1913 -3100
rect 2025 -3049 2317 -3032
rect 2025 -3100 2045 -3049
rect 2295 -3100 2317 -3049
rect 2025 -3117 2317 -3100
rect 62 -3905 1134 -3892
rect 62 -3952 83 -3905
rect 1105 -3952 1134 -3905
rect 62 -3967 1134 -3952
rect 1634 -3905 2706 -3892
rect 1634 -3952 1655 -3905
rect 2677 -3952 2706 -3905
rect 1634 -3967 2706 -3952
rect 1206 -4011 1498 -3994
rect 1206 -4062 1226 -4011
rect 1476 -4062 1498 -4011
rect 2778 -4011 3070 -3994
rect 1206 -4079 1498 -4062
rect 2778 -4062 2798 -4011
rect 3048 -4062 3070 -4011
rect 2778 -4079 3070 -4062
rect 3343 -4011 3635 -3994
rect 3343 -4062 3363 -4011
rect 3613 -4062 3635 -4011
rect 3343 -4079 3635 -4062
rect 3747 -4011 4039 -3994
rect 3747 -4062 3767 -4011
rect 4017 -4062 4039 -4011
rect 3747 -4079 4039 -4062
<< psubdiffcont >>
rect 87 37 794 83
rect 891 29 1200 78
rect 1447 37 2154 83
rect 2251 29 2560 78
rect 2745 29 3054 78
rect 3149 29 3458 78
rect 87 -902 794 -856
rect 891 -910 1200 -861
rect 1416 -910 1725 -861
rect 1820 -910 2129 -861
rect 2548 -910 2857 -861
rect 2952 -910 3261 -861
rect 102 -1868 1086 -1822
rect 1211 -1871 1520 -1822
rect 1700 -1863 2407 -1817
rect 2504 -1871 2813 -1822
rect 2919 -1871 3228 -1822
rect 3323 -1871 3632 -1822
rect 87 -2800 794 -2754
rect 891 -2808 1200 -2759
rect 1391 -2826 2375 -2780
rect 2500 -2829 2809 -2780
rect 2915 -2829 3224 -2780
rect 3319 -2829 3628 -2780
rect 102 -3786 1086 -3740
rect 1211 -3789 1520 -3740
rect 1626 -3789 1935 -3740
rect 2030 -3789 2339 -3740
rect 102 -4748 1086 -4702
rect 1211 -4751 1520 -4702
rect 1674 -4748 2658 -4702
rect 2783 -4751 3092 -4702
rect 3348 -4751 3657 -4702
rect 3752 -4751 4061 -4702
<< nsubdiffcont >>
rect 88 799 787 851
rect 1448 799 2147 851
rect 906 718 1156 769
rect 2266 718 2516 769
rect 2760 718 3010 769
rect 3164 718 3414 769
rect 88 -140 787 -88
rect 906 -221 1156 -170
rect 1431 -221 1681 -170
rect 1835 -221 2085 -170
rect 2563 -221 2813 -170
rect 2967 -221 3217 -170
rect 83 -1072 1105 -1025
rect 1701 -1101 2400 -1049
rect 1226 -1182 1476 -1131
rect 2519 -1182 2769 -1131
rect 2934 -1182 3184 -1131
rect 3338 -1182 3588 -1131
rect 88 -2038 787 -1986
rect 1372 -2030 2394 -1983
rect 906 -2119 1156 -2068
rect 2515 -2140 2765 -2089
rect 2930 -2140 3180 -2089
rect 3334 -2140 3584 -2089
rect 83 -2990 1105 -2943
rect 1226 -3100 1476 -3049
rect 1641 -3100 1891 -3049
rect 2045 -3100 2295 -3049
rect 83 -3952 1105 -3905
rect 1655 -3952 2677 -3905
rect 1226 -4062 1476 -4011
rect 2798 -4062 3048 -4011
rect 3363 -4062 3613 -4011
rect 3767 -4062 4017 -4011
<< polysilicon >>
rect 212 654 268 698
rect 616 654 672 698
rect 0 566 89 579
rect 0 507 13 566
rect 76 528 89 566
rect 1020 621 1076 665
rect 1572 654 1628 698
rect 1976 654 2032 698
rect 212 528 268 554
rect 76 507 268 528
rect 0 492 268 507
rect 212 315 268 492
rect 401 418 490 431
rect 401 359 414 418
rect 477 381 490 418
rect 616 381 672 554
rect 1360 566 1449 579
rect 1020 459 1076 521
rect 1360 507 1373 566
rect 1436 528 1449 566
rect 2380 621 2436 665
rect 2874 621 2930 665
rect 3278 621 3334 665
rect 1572 528 1628 554
rect 1436 507 1628 528
rect 1360 492 1628 507
rect 477 359 672 381
rect 961 445 1076 459
rect 961 386 975 445
rect 1038 386 1076 445
rect 961 372 1076 386
rect 401 344 672 359
rect 616 315 672 344
rect 1020 272 1076 372
rect 1572 315 1628 492
rect 1761 418 1850 431
rect 1761 359 1774 418
rect 1837 381 1850 418
rect 1976 381 2032 554
rect 2380 459 2436 521
rect 2874 459 2930 521
rect 3278 459 3334 521
rect 1837 359 2032 381
rect 2321 445 2436 459
rect 2321 386 2335 445
rect 2398 386 2436 445
rect 2321 372 2436 386
rect 2815 445 2930 459
rect 2815 386 2829 445
rect 2892 386 2930 445
rect 2815 372 2930 386
rect 3219 445 3334 459
rect 3219 386 3233 445
rect 3296 386 3334 445
rect 3219 372 3334 386
rect 1761 344 2032 359
rect 1976 315 2032 344
rect 212 171 268 215
rect 616 171 672 215
rect 1020 178 1076 222
rect 2380 272 2436 372
rect 1572 171 1628 215
rect 1976 171 2032 215
rect 2380 178 2436 222
rect 2874 272 2930 372
rect 2874 178 2930 222
rect 3278 272 3334 372
rect 3278 178 3334 222
rect 212 -285 268 -241
rect 616 -285 672 -241
rect 0 -373 89 -360
rect 0 -432 13 -373
rect 76 -411 89 -373
rect 1020 -318 1076 -274
rect 1545 -318 1601 -274
rect 1949 -318 2005 -274
rect 2677 -318 2733 -274
rect 3081 -318 3137 -274
rect 212 -411 268 -385
rect 76 -432 268 -411
rect 0 -447 268 -432
rect 212 -624 268 -447
rect 401 -521 490 -508
rect 401 -580 414 -521
rect 477 -558 490 -521
rect 616 -558 672 -385
rect 1020 -480 1076 -418
rect 1545 -480 1601 -418
rect 1949 -480 2005 -418
rect 2677 -480 2733 -418
rect 3081 -480 3137 -418
rect 477 -580 672 -558
rect 961 -494 1076 -480
rect 961 -553 975 -494
rect 1038 -553 1076 -494
rect 961 -567 1076 -553
rect 1486 -494 1601 -480
rect 1486 -553 1500 -494
rect 1563 -553 1601 -494
rect 1486 -567 1601 -553
rect 1890 -494 2005 -480
rect 1890 -553 1904 -494
rect 1967 -553 2005 -494
rect 1890 -567 2005 -553
rect 2618 -494 2733 -480
rect 2618 -553 2632 -494
rect 2695 -553 2733 -494
rect 2618 -567 2733 -553
rect 3022 -494 3137 -480
rect 3022 -553 3036 -494
rect 3099 -553 3137 -494
rect 3022 -567 3137 -553
rect 401 -595 672 -580
rect 616 -624 672 -595
rect 1020 -667 1076 -567
rect 212 -768 268 -724
rect 616 -768 672 -724
rect 1020 -761 1076 -717
rect 1545 -667 1601 -567
rect 1545 -761 1601 -717
rect 1949 -667 2005 -567
rect 1949 -761 2005 -717
rect 2677 -667 2733 -567
rect 2677 -761 2733 -717
rect 3081 -667 3137 -567
rect 3081 -761 3137 -717
rect 212 -1198 428 -1162
rect 212 -1226 268 -1198
rect 372 -1226 428 -1198
rect 776 -1199 992 -1160
rect 776 -1226 832 -1199
rect 936 -1226 992 -1199
rect 1340 -1279 1396 -1235
rect 1825 -1246 1881 -1202
rect 2229 -1246 2285 -1202
rect 212 -1370 268 -1326
rect 372 -1488 428 -1326
rect 776 -1373 832 -1326
rect 936 -1370 992 -1326
rect 697 -1387 832 -1373
rect 1613 -1334 1702 -1321
rect 697 -1446 710 -1387
rect 773 -1446 832 -1387
rect 1340 -1441 1396 -1379
rect 1613 -1393 1626 -1334
rect 1689 -1372 1702 -1334
rect 2633 -1279 2689 -1235
rect 3048 -1279 3104 -1235
rect 3452 -1279 3508 -1235
rect 1825 -1372 1881 -1346
rect 1689 -1393 1881 -1372
rect 1613 -1408 1881 -1393
rect 697 -1460 832 -1446
rect 296 -1501 428 -1488
rect 296 -1560 310 -1501
rect 373 -1560 428 -1501
rect 296 -1575 428 -1560
rect 372 -1626 428 -1575
rect 372 -1720 428 -1676
rect 776 -1626 832 -1460
rect 1281 -1455 1396 -1441
rect 1281 -1514 1295 -1455
rect 1358 -1514 1396 -1455
rect 1281 -1528 1396 -1514
rect 776 -1720 832 -1676
rect 1340 -1628 1396 -1528
rect 1825 -1585 1881 -1408
rect 2014 -1482 2103 -1469
rect 2014 -1541 2027 -1482
rect 2090 -1519 2103 -1482
rect 2229 -1519 2285 -1346
rect 2633 -1441 2689 -1379
rect 3048 -1441 3104 -1379
rect 3452 -1441 3508 -1379
rect 2090 -1541 2285 -1519
rect 2574 -1455 2689 -1441
rect 2574 -1514 2588 -1455
rect 2651 -1514 2689 -1455
rect 2574 -1528 2689 -1514
rect 2989 -1455 3104 -1441
rect 2989 -1514 3003 -1455
rect 3066 -1514 3104 -1455
rect 2989 -1528 3104 -1514
rect 3393 -1455 3508 -1441
rect 3393 -1514 3407 -1455
rect 3470 -1514 3508 -1455
rect 3393 -1528 3508 -1514
rect 2014 -1556 2285 -1541
rect 2229 -1585 2285 -1556
rect 1340 -1722 1396 -1678
rect 2633 -1628 2689 -1528
rect 1825 -1729 1881 -1685
rect 2229 -1729 2285 -1685
rect 2633 -1722 2689 -1678
rect 3048 -1628 3104 -1528
rect 3048 -1722 3104 -1678
rect 3452 -1628 3508 -1528
rect 3452 -1722 3508 -1678
rect 212 -2183 268 -2139
rect 616 -2183 672 -2139
rect 1501 -2156 1717 -2120
rect 0 -2271 89 -2258
rect 0 -2330 13 -2271
rect 76 -2309 89 -2271
rect 1020 -2216 1076 -2172
rect 1501 -2184 1557 -2156
rect 1661 -2184 1717 -2156
rect 2065 -2157 2281 -2118
rect 2065 -2184 2121 -2157
rect 2225 -2184 2281 -2157
rect 212 -2309 268 -2283
rect 76 -2330 268 -2309
rect 0 -2345 268 -2330
rect 212 -2522 268 -2345
rect 401 -2419 490 -2406
rect 401 -2478 414 -2419
rect 477 -2456 490 -2419
rect 616 -2456 672 -2283
rect 2629 -2237 2685 -2193
rect 3044 -2237 3100 -2193
rect 3448 -2237 3504 -2193
rect 1020 -2378 1076 -2316
rect 1501 -2328 1557 -2284
rect 477 -2478 672 -2456
rect 961 -2392 1076 -2378
rect 961 -2451 975 -2392
rect 1038 -2451 1076 -2392
rect 1661 -2446 1717 -2284
rect 2065 -2331 2121 -2284
rect 2225 -2328 2281 -2284
rect 1986 -2345 2121 -2331
rect 1986 -2404 1999 -2345
rect 2062 -2404 2121 -2345
rect 2629 -2399 2685 -2337
rect 3044 -2399 3100 -2337
rect 3448 -2399 3504 -2337
rect 1986 -2418 2121 -2404
rect 961 -2465 1076 -2451
rect 401 -2493 672 -2478
rect 616 -2522 672 -2493
rect 1020 -2565 1076 -2465
rect 1585 -2459 1717 -2446
rect 1585 -2518 1599 -2459
rect 1662 -2518 1717 -2459
rect 1585 -2533 1717 -2518
rect 212 -2666 268 -2622
rect 616 -2666 672 -2622
rect 1020 -2659 1076 -2615
rect 1661 -2584 1717 -2533
rect 1661 -2678 1717 -2634
rect 2065 -2584 2121 -2418
rect 2570 -2413 2685 -2399
rect 2570 -2472 2584 -2413
rect 2647 -2472 2685 -2413
rect 2570 -2486 2685 -2472
rect 2985 -2413 3100 -2399
rect 2985 -2472 2999 -2413
rect 3062 -2472 3100 -2413
rect 2985 -2486 3100 -2472
rect 3389 -2413 3504 -2399
rect 3389 -2472 3403 -2413
rect 3466 -2472 3504 -2413
rect 3389 -2486 3504 -2472
rect 2065 -2678 2121 -2634
rect 2629 -2586 2685 -2486
rect 2629 -2680 2685 -2636
rect 3044 -2586 3100 -2486
rect 3044 -2680 3100 -2636
rect 3448 -2586 3504 -2486
rect 3448 -2680 3504 -2636
rect 212 -3116 428 -3080
rect 212 -3144 268 -3116
rect 372 -3144 428 -3116
rect 776 -3117 992 -3078
rect 776 -3144 832 -3117
rect 936 -3144 992 -3117
rect 1340 -3197 1396 -3153
rect 1755 -3197 1811 -3153
rect 2159 -3197 2215 -3153
rect 212 -3288 268 -3244
rect 372 -3406 428 -3244
rect 776 -3291 832 -3244
rect 936 -3288 992 -3244
rect 697 -3305 832 -3291
rect 697 -3364 710 -3305
rect 773 -3364 832 -3305
rect 1340 -3359 1396 -3297
rect 1755 -3359 1811 -3297
rect 2159 -3359 2215 -3297
rect 697 -3378 832 -3364
rect 296 -3419 428 -3406
rect 296 -3478 310 -3419
rect 373 -3478 428 -3419
rect 296 -3493 428 -3478
rect 372 -3544 428 -3493
rect 372 -3638 428 -3594
rect 776 -3544 832 -3378
rect 1281 -3373 1396 -3359
rect 1281 -3432 1295 -3373
rect 1358 -3432 1396 -3373
rect 1281 -3446 1396 -3432
rect 1696 -3373 1811 -3359
rect 1696 -3432 1710 -3373
rect 1773 -3432 1811 -3373
rect 1696 -3446 1811 -3432
rect 2100 -3373 2215 -3359
rect 2100 -3432 2114 -3373
rect 2177 -3432 2215 -3373
rect 2100 -3446 2215 -3432
rect 776 -3638 832 -3594
rect 1340 -3546 1396 -3446
rect 1340 -3640 1396 -3596
rect 1755 -3546 1811 -3446
rect 1755 -3640 1811 -3596
rect 2159 -3546 2215 -3446
rect 2159 -3640 2215 -3596
rect 212 -4078 428 -4042
rect 212 -4106 268 -4078
rect 372 -4106 428 -4078
rect 776 -4079 992 -4040
rect 1784 -4078 2000 -4042
rect 776 -4106 832 -4079
rect 936 -4106 992 -4079
rect 1784 -4106 1840 -4078
rect 1944 -4106 2000 -4078
rect 2348 -4079 2564 -4040
rect 2348 -4106 2404 -4079
rect 2508 -4106 2564 -4079
rect 1340 -4159 1396 -4115
rect 212 -4250 268 -4206
rect 372 -4368 428 -4206
rect 776 -4253 832 -4206
rect 936 -4250 992 -4206
rect 697 -4267 832 -4253
rect 2912 -4159 2968 -4115
rect 3477 -4159 3533 -4115
rect 3881 -4159 3937 -4115
rect 1784 -4250 1840 -4206
rect 697 -4326 710 -4267
rect 773 -4326 832 -4267
rect 1340 -4321 1396 -4259
rect 697 -4340 832 -4326
rect 296 -4381 428 -4368
rect 296 -4440 310 -4381
rect 373 -4440 428 -4381
rect 296 -4455 428 -4440
rect 372 -4506 428 -4455
rect 372 -4600 428 -4556
rect 776 -4506 832 -4340
rect 1281 -4335 1396 -4321
rect 1281 -4394 1295 -4335
rect 1358 -4394 1396 -4335
rect 1944 -4368 2000 -4206
rect 2348 -4253 2404 -4206
rect 2508 -4250 2564 -4206
rect 2269 -4267 2404 -4253
rect 2269 -4326 2282 -4267
rect 2345 -4326 2404 -4267
rect 2912 -4321 2968 -4259
rect 3477 -4321 3533 -4259
rect 3881 -4321 3937 -4259
rect 2269 -4340 2404 -4326
rect 1281 -4408 1396 -4394
rect 776 -4600 832 -4556
rect 1340 -4508 1396 -4408
rect 1868 -4381 2000 -4368
rect 1868 -4440 1882 -4381
rect 1945 -4440 2000 -4381
rect 1868 -4455 2000 -4440
rect 1340 -4602 1396 -4558
rect 1944 -4506 2000 -4455
rect 1944 -4600 2000 -4556
rect 2348 -4506 2404 -4340
rect 2853 -4335 2968 -4321
rect 2853 -4394 2867 -4335
rect 2930 -4394 2968 -4335
rect 2853 -4408 2968 -4394
rect 3418 -4335 3533 -4321
rect 3418 -4394 3432 -4335
rect 3495 -4394 3533 -4335
rect 3418 -4408 3533 -4394
rect 3822 -4335 3937 -4321
rect 3822 -4394 3836 -4335
rect 3899 -4394 3937 -4335
rect 3822 -4408 3937 -4394
rect 2348 -4600 2404 -4556
rect 2912 -4508 2968 -4408
rect 2912 -4602 2968 -4558
rect 3477 -4508 3533 -4408
rect 3477 -4602 3533 -4558
rect 3881 -4508 3937 -4408
rect 3881 -4602 3937 -4558
<< polycontact >>
rect 13 507 76 566
rect 414 359 477 418
rect 1373 507 1436 566
rect 975 386 1038 445
rect 1774 359 1837 418
rect 2335 386 2398 445
rect 2829 386 2892 445
rect 3233 386 3296 445
rect 13 -432 76 -373
rect 414 -580 477 -521
rect 975 -553 1038 -494
rect 1500 -553 1563 -494
rect 1904 -553 1967 -494
rect 2632 -553 2695 -494
rect 3036 -553 3099 -494
rect 710 -1446 773 -1387
rect 1626 -1393 1689 -1334
rect 310 -1560 373 -1501
rect 1295 -1514 1358 -1455
rect 2027 -1541 2090 -1482
rect 2588 -1514 2651 -1455
rect 3003 -1514 3066 -1455
rect 3407 -1514 3470 -1455
rect 13 -2330 76 -2271
rect 414 -2478 477 -2419
rect 975 -2451 1038 -2392
rect 1999 -2404 2062 -2345
rect 1599 -2518 1662 -2459
rect 2584 -2472 2647 -2413
rect 2999 -2472 3062 -2413
rect 3403 -2472 3466 -2413
rect 710 -3364 773 -3305
rect 310 -3478 373 -3419
rect 1295 -3432 1358 -3373
rect 1710 -3432 1773 -3373
rect 2114 -3432 2177 -3373
rect 710 -4326 773 -4267
rect 310 -4440 373 -4381
rect 1295 -4394 1358 -4335
rect 2282 -4326 2345 -4267
rect 1882 -4440 1945 -4381
rect 2867 -4394 2930 -4335
rect 3432 -4394 3495 -4335
rect 3836 -4394 3899 -4335
<< metal1 >>
rect -821 847 -747 856
rect 38 851 3508 891
rect 38 847 88 851
rect -821 791 -812 847
rect -756 799 88 847
rect 787 799 1448 851
rect 2147 799 3508 851
rect -756 791 3508 799
rect -821 781 -747 791
rect 38 773 3508 791
rect 137 641 183 773
rect -655 576 -581 585
rect -10 576 89 579
rect -655 520 -646 576
rect -590 566 89 576
rect -590 520 13 566
rect -655 511 -581 520
rect -10 507 13 520
rect 76 507 89 566
rect 137 556 183 567
rect 297 641 343 652
rect 541 641 587 652
rect 343 586 541 632
rect 297 556 343 567
rect -10 492 89 507
rect 541 500 587 567
rect 701 641 747 773
rect 846 769 1250 773
rect 846 718 906 769
rect 1156 718 1250 769
rect 846 700 1250 718
rect 701 556 747 567
rect 922 608 992 700
rect 1497 641 1543 773
rect 922 534 945 608
rect 991 534 992 608
rect 922 519 992 534
rect 1104 608 1168 621
rect 1104 534 1105 608
rect 1151 534 1168 608
rect 541 454 747 500
rect -489 426 -417 435
rect -489 372 -480 426
rect -426 422 -417 426
rect 401 422 490 431
rect -426 418 490 422
rect -426 376 414 418
rect -426 372 -417 376
rect -489 363 -417 372
rect 401 359 414 376
rect 477 359 490 418
rect 401 344 490 359
rect 701 428 747 454
rect 846 445 1050 453
rect 846 428 975 445
rect 701 386 975 428
rect 1038 386 1050 445
rect 701 382 1050 386
rect -12 299 68 308
rect -12 243 0 299
rect 56 243 68 299
rect -12 234 68 243
rect 137 302 183 313
rect 137 118 183 228
rect 297 302 343 313
rect 541 302 587 313
rect 343 244 541 290
rect 297 217 343 228
rect 541 217 587 228
rect 701 302 747 382
rect 846 372 1050 382
rect 1104 418 1168 534
rect 1360 566 1449 579
rect 1360 507 1373 566
rect 1436 507 1449 566
rect 1497 556 1543 567
rect 1657 641 1703 652
rect 1901 641 1947 652
rect 1703 586 1901 632
rect 1657 556 1703 567
rect 1360 492 1449 507
rect 1901 500 1947 567
rect 2061 641 2107 773
rect 2206 769 3508 773
rect 2206 718 2266 769
rect 2516 718 2760 769
rect 3010 718 3164 769
rect 3414 718 3508 769
rect 2206 700 3508 718
rect 2061 556 2107 567
rect 2282 608 2352 700
rect 2282 534 2305 608
rect 2351 534 2352 608
rect 2282 519 2352 534
rect 2464 608 2528 621
rect 2464 534 2465 608
rect 2511 534 2528 608
rect 1901 454 2107 500
rect 1761 422 1850 431
rect 1314 418 1850 422
rect 1104 376 1774 418
rect 1104 371 1360 376
rect 701 217 747 228
rect 919 270 1000 275
rect 1104 270 1168 371
rect 1761 359 1774 376
rect 1837 359 1850 418
rect 1761 344 1850 359
rect 2061 428 2107 454
rect 2206 445 2410 453
rect 2206 428 2335 445
rect 2061 386 2335 428
rect 2398 386 2410 445
rect 2061 382 2410 386
rect 919 224 941 270
rect 987 224 1000 270
rect 1098 224 1109 270
rect 1155 224 1168 270
rect 38 113 846 118
rect 919 113 1000 224
rect 1104 223 1168 224
rect 1497 302 1543 313
rect 1497 118 1543 228
rect 1657 302 1703 313
rect 1901 302 1947 313
rect 1703 244 1901 290
rect 1657 217 1703 228
rect 1901 217 1947 228
rect 2061 302 2107 382
rect 2206 372 2410 382
rect 2464 418 2528 534
rect 2776 608 2846 700
rect 2776 534 2799 608
rect 2845 534 2846 608
rect 2776 519 2846 534
rect 2958 608 3022 621
rect 2958 534 2959 608
rect 3005 534 3022 608
rect 2610 445 2904 453
rect 2610 418 2829 445
rect 2464 386 2829 418
rect 2892 386 2904 445
rect 2464 372 2904 386
rect 2958 418 3022 534
rect 3180 608 3250 700
rect 3180 534 3203 608
rect 3249 534 3250 608
rect 3180 519 3250 534
rect 3362 608 3426 621
rect 3362 534 3363 608
rect 3409 534 3426 608
rect 3104 445 3308 453
rect 3104 418 3233 445
rect 2958 386 3233 418
rect 3296 386 3308 445
rect 2958 372 3308 386
rect 3362 418 3426 534
rect 2464 371 2641 372
rect 2958 371 3127 372
rect 3362 371 3568 418
rect 2061 217 2107 228
rect 2279 270 2360 275
rect 2464 270 2528 371
rect 2279 224 2301 270
rect 2347 224 2360 270
rect 2458 224 2469 270
rect 2515 224 2528 270
rect 1250 113 2206 118
rect 2279 113 2360 224
rect 2464 223 2528 224
rect 2773 270 2854 275
rect 2958 270 3022 371
rect 2773 224 2795 270
rect 2841 224 2854 270
rect 2952 224 2963 270
rect 3009 224 3022 270
rect 2773 113 2854 224
rect 2958 223 3022 224
rect 3177 270 3258 275
rect 3362 270 3426 371
rect 3177 224 3199 270
rect 3245 224 3258 270
rect 3356 224 3367 270
rect 3413 224 3426 270
rect 3177 113 3258 224
rect 3362 223 3426 224
rect -198 100 -126 109
rect -198 46 -189 100
rect -135 97 -126 100
rect 38 97 3508 113
rect -135 83 3508 97
rect -135 48 87 83
rect -135 46 -126 48
rect -198 37 -126 46
rect 38 37 87 48
rect 794 78 1447 83
rect 794 37 891 78
rect 38 29 891 37
rect 1200 37 1447 78
rect 2154 78 3508 83
rect 2154 37 2251 78
rect 1200 29 2251 37
rect 2560 29 2745 78
rect 3054 29 3149 78
rect 3458 29 3508 78
rect 38 0 3508 29
rect -822 -84 -748 -75
rect 38 -84 3311 -48
rect -822 -140 -812 -84
rect -756 -88 3311 -84
rect -756 -140 88 -88
rect 787 -126 3311 -88
rect 787 -140 2179 -126
rect -822 -149 -748 -140
rect 38 -166 2179 -140
rect 137 -298 183 -166
rect -658 -375 -587 -363
rect -4 -370 89 -360
rect -21 -373 89 -370
rect -21 -375 13 -373
rect -658 -431 -646 -375
rect -590 -376 13 -375
rect -590 -430 7 -376
rect -590 -431 13 -430
rect -658 -443 -587 -431
rect -21 -432 13 -431
rect 76 -432 89 -373
rect 137 -383 183 -372
rect 297 -298 343 -287
rect 541 -298 587 -287
rect 343 -353 541 -307
rect 297 -383 343 -372
rect -21 -446 89 -432
rect -4 -447 89 -446
rect 541 -439 587 -372
rect 701 -298 747 -166
rect 846 -170 2179 -166
rect 846 -221 906 -170
rect 1156 -221 1431 -170
rect 1681 -221 1835 -170
rect 2085 -221 2179 -170
rect 846 -239 2179 -221
rect 2492 -170 3311 -126
rect 2492 -221 2563 -170
rect 2813 -221 2967 -170
rect 3217 -221 3311 -170
rect 2492 -239 3311 -221
rect 701 -383 747 -372
rect 922 -331 992 -239
rect 922 -405 945 -331
rect 991 -405 992 -331
rect 922 -420 992 -405
rect 1104 -331 1168 -318
rect 1104 -405 1105 -331
rect 1151 -405 1168 -331
rect 541 -485 747 -439
rect -500 -513 -428 -504
rect -500 -567 -491 -513
rect -437 -517 -428 -513
rect 401 -517 490 -508
rect -437 -521 490 -517
rect -437 -563 414 -521
rect -437 -567 -428 -563
rect -500 -576 -428 -567
rect 401 -580 414 -563
rect 477 -580 490 -521
rect 401 -595 490 -580
rect 701 -511 747 -485
rect 846 -494 1050 -486
rect 846 -511 975 -494
rect 701 -553 975 -511
rect 1038 -553 1050 -494
rect 701 -557 1050 -553
rect 137 -637 183 -626
rect 137 -821 183 -711
rect 297 -637 343 -626
rect 541 -637 587 -626
rect 343 -695 541 -649
rect 297 -722 343 -711
rect 541 -722 587 -711
rect 701 -637 747 -557
rect 846 -567 1050 -557
rect 1104 -521 1168 -405
rect 1447 -331 1517 -239
rect 1447 -405 1470 -331
rect 1516 -405 1517 -331
rect 1447 -420 1517 -405
rect 1629 -331 1693 -318
rect 1629 -405 1630 -331
rect 1676 -405 1693 -331
rect 1281 -494 1575 -486
rect 1281 -521 1500 -494
rect 1104 -553 1500 -521
rect 1563 -553 1575 -494
rect 1104 -567 1575 -553
rect 1629 -521 1693 -405
rect 1851 -331 1921 -239
rect 1851 -405 1874 -331
rect 1920 -405 1921 -331
rect 1851 -420 1921 -405
rect 2033 -331 2097 -318
rect 2033 -405 2034 -331
rect 2080 -405 2097 -331
rect 1775 -494 1979 -486
rect 1775 -521 1904 -494
rect 1629 -553 1904 -521
rect 1967 -553 1979 -494
rect 1629 -567 1979 -553
rect 2033 -521 2097 -405
rect 2579 -331 2649 -239
rect 2579 -405 2602 -331
rect 2648 -405 2649 -331
rect 2579 -420 2649 -405
rect 2761 -331 2825 -318
rect 2761 -405 2762 -331
rect 2808 -405 2825 -331
rect 2413 -494 2707 -486
rect 2413 -501 2632 -494
rect 2380 -509 2632 -501
rect 2208 -521 2255 -520
rect 1104 -568 1281 -567
rect 1629 -568 1798 -567
rect 2033 -568 2264 -521
rect 2380 -565 2399 -509
rect 2455 -553 2632 -509
rect 2695 -553 2707 -494
rect 2455 -565 2707 -553
rect 2380 -567 2707 -565
rect 2761 -521 2825 -405
rect 2983 -331 3053 -239
rect 2983 -405 3006 -331
rect 3052 -405 3053 -331
rect 2983 -420 3053 -405
rect 3165 -331 3229 -318
rect 3165 -405 3166 -331
rect 3212 -405 3229 -331
rect 2907 -494 3111 -486
rect 2907 -521 3036 -494
rect 2761 -553 3036 -521
rect 3099 -553 3111 -494
rect 2761 -567 3111 -553
rect 3165 -521 3229 -405
rect 3333 -344 3410 -329
rect 3333 -400 3340 -344
rect 3396 -400 3410 -344
rect 3333 -414 3410 -400
rect 701 -722 747 -711
rect 919 -669 1000 -664
rect 1104 -669 1168 -568
rect 919 -715 941 -669
rect 987 -715 1000 -669
rect 1098 -715 1109 -669
rect 1155 -715 1168 -669
rect 38 -826 846 -821
rect 919 -826 1000 -715
rect 1104 -716 1168 -715
rect 1444 -669 1525 -664
rect 1629 -669 1693 -568
rect 1444 -715 1466 -669
rect 1512 -715 1525 -669
rect 1623 -715 1634 -669
rect 1680 -715 1693 -669
rect 1444 -826 1525 -715
rect 1629 -716 1693 -715
rect 1848 -669 1929 -664
rect 2033 -669 2097 -568
rect 1848 -715 1870 -669
rect 1916 -715 1929 -669
rect 2027 -715 2038 -669
rect 2084 -715 2097 -669
rect 2208 -657 2255 -568
rect 2380 -577 2466 -567
rect 2761 -568 2930 -567
rect 3165 -568 3407 -521
rect 2358 -653 2452 -635
rect 2358 -657 2382 -653
rect 2208 -704 2382 -657
rect 1848 -826 1929 -715
rect 2033 -716 2097 -715
rect 2358 -707 2382 -704
rect 2436 -707 2452 -653
rect 2358 -726 2452 -707
rect 2576 -669 2657 -664
rect 2761 -669 2825 -568
rect 2576 -715 2598 -669
rect 2644 -715 2657 -669
rect 2755 -715 2766 -669
rect 2812 -715 2825 -669
rect 2576 -826 2657 -715
rect 2761 -716 2825 -715
rect 2980 -669 3061 -664
rect 3165 -669 3229 -568
rect 2980 -715 3002 -669
rect 3048 -715 3061 -669
rect 3159 -715 3170 -669
rect 3216 -715 3229 -669
rect 2980 -826 3061 -715
rect 3165 -716 3229 -715
rect -201 -854 -127 -846
rect 38 -849 3311 -826
rect -19 -854 3311 -849
rect -201 -910 -190 -854
rect -134 -856 3311 -854
rect -134 -902 87 -856
rect 794 -861 3311 -856
rect 794 -902 891 -861
rect -134 -910 891 -902
rect 1200 -910 1416 -861
rect 1725 -910 1820 -861
rect 2129 -910 2548 -861
rect 2857 -910 2952 -861
rect 3261 -910 3311 -861
rect -201 -918 -127 -910
rect -19 -913 3311 -910
rect 38 -939 3311 -913
rect -825 -1013 -747 -1005
rect 38 -1013 3682 -988
rect -825 -1069 -812 -1013
rect -756 -1025 3682 -1013
rect -756 -1069 83 -1025
rect -825 -1081 -747 -1069
rect 38 -1072 83 -1069
rect 1105 -1049 3682 -1025
rect 1105 -1072 1701 -1049
rect 38 -1087 1701 -1072
rect -658 -1193 -583 -1187
rect -57 -1193 19 -1185
rect -658 -1194 19 -1193
rect -658 -1249 -646 -1194
rect -591 -1249 -48 -1194
rect -658 -1250 -48 -1249
rect -658 -1260 -583 -1250
rect -57 -1251 -48 -1250
rect 9 -1251 19 -1194
rect -57 -1260 19 -1251
rect 137 -1239 183 -1087
rect 280 -1138 359 -1136
rect 280 -1192 293 -1138
rect 347 -1192 359 -1138
rect 280 -1200 359 -1192
rect 137 -1324 183 -1313
rect 297 -1239 343 -1200
rect 297 -1324 343 -1313
rect 457 -1239 503 -1087
rect 1166 -1131 1570 -1087
rect 1651 -1101 1701 -1087
rect 2400 -1101 3682 -1049
rect 1651 -1127 3682 -1101
rect 687 -1136 761 -1134
rect 687 -1147 1067 -1136
rect 687 -1201 697 -1147
rect 751 -1182 1067 -1147
rect 751 -1201 761 -1182
rect 687 -1214 761 -1201
rect 457 -1324 503 -1313
rect 701 -1239 747 -1214
rect 701 -1324 747 -1313
rect 861 -1239 907 -1228
rect -502 -1370 -424 -1361
rect -502 -1424 -491 -1370
rect -437 -1374 -424 -1370
rect 697 -1374 786 -1373
rect -437 -1387 786 -1374
rect -437 -1420 710 -1387
rect -437 -1424 -424 -1420
rect -502 -1433 -424 -1424
rect 697 -1446 710 -1420
rect 773 -1446 786 -1387
rect 697 -1460 786 -1446
rect -354 -1505 -274 -1496
rect -354 -1559 -344 -1505
rect -290 -1509 -274 -1505
rect 296 -1501 385 -1488
rect 296 -1509 310 -1501
rect -290 -1555 310 -1509
rect -290 -1559 -274 -1555
rect -354 -1569 -274 -1559
rect 296 -1560 310 -1555
rect 373 -1560 385 -1501
rect 861 -1536 907 -1313
rect 1021 -1239 1067 -1182
rect 1166 -1182 1226 -1131
rect 1476 -1182 1570 -1131
rect 1166 -1200 1570 -1182
rect 1021 -1324 1067 -1313
rect 1242 -1292 1312 -1200
rect 1750 -1259 1796 -1127
rect 1242 -1366 1265 -1292
rect 1311 -1366 1312 -1292
rect 1242 -1381 1312 -1366
rect 1424 -1292 1488 -1279
rect 1424 -1366 1425 -1292
rect 1471 -1366 1488 -1292
rect 296 -1575 385 -1560
rect 457 -1582 907 -1536
rect 457 -1628 503 -1582
rect 861 -1588 907 -1582
rect 1126 -1455 1370 -1447
rect 1126 -1514 1295 -1455
rect 1358 -1514 1370 -1455
rect 1126 -1528 1370 -1514
rect 1424 -1482 1488 -1366
rect 1613 -1334 1702 -1321
rect 1613 -1393 1626 -1334
rect 1689 -1393 1702 -1334
rect 1750 -1344 1796 -1333
rect 1910 -1259 1956 -1248
rect 2154 -1259 2200 -1248
rect 1956 -1314 2154 -1268
rect 1910 -1344 1956 -1333
rect 1613 -1408 1702 -1393
rect 2154 -1400 2200 -1333
rect 2314 -1259 2360 -1127
rect 2459 -1131 3682 -1127
rect 2459 -1182 2519 -1131
rect 2769 -1182 2934 -1131
rect 3184 -1182 3338 -1131
rect 3588 -1182 3682 -1131
rect 2459 -1200 3682 -1182
rect 2314 -1344 2360 -1333
rect 2535 -1292 2605 -1200
rect 2535 -1366 2558 -1292
rect 2604 -1366 2605 -1292
rect 2535 -1381 2605 -1366
rect 2717 -1292 2781 -1279
rect 2717 -1366 2718 -1292
rect 2764 -1366 2781 -1292
rect 2154 -1446 2360 -1400
rect 2014 -1478 2103 -1469
rect 1613 -1482 2103 -1478
rect 1424 -1524 2027 -1482
rect 1126 -1588 1172 -1528
rect 861 -1628 1172 -1588
rect 1424 -1529 1676 -1524
rect 282 -1674 293 -1628
rect 339 -1674 350 -1628
rect 450 -1674 461 -1628
rect 507 -1674 518 -1628
rect 686 -1674 697 -1628
rect 743 -1674 754 -1628
rect 854 -1674 865 -1628
rect 911 -1634 1172 -1628
rect 1239 -1630 1320 -1625
rect 1424 -1630 1488 -1529
rect 2014 -1541 2027 -1524
rect 2090 -1541 2103 -1482
rect 2014 -1556 2103 -1541
rect 2314 -1472 2360 -1446
rect 2717 -1447 2781 -1366
rect 2950 -1292 3020 -1200
rect 2950 -1366 2973 -1292
rect 3019 -1366 3020 -1292
rect 2950 -1381 3020 -1366
rect 3132 -1292 3196 -1279
rect 3132 -1366 3133 -1292
rect 3179 -1366 3196 -1292
rect 2459 -1455 2663 -1447
rect 2459 -1472 2588 -1455
rect 2314 -1514 2588 -1472
rect 2651 -1514 2663 -1455
rect 2314 -1518 2663 -1514
rect 911 -1674 922 -1634
rect 282 -1782 350 -1674
rect 686 -1782 754 -1674
rect 1239 -1676 1261 -1630
rect 1307 -1676 1320 -1630
rect 1418 -1676 1429 -1630
rect 1475 -1676 1488 -1630
rect 1239 -1782 1320 -1676
rect 1424 -1677 1488 -1676
rect 1750 -1598 1796 -1587
rect 1750 -1782 1796 -1672
rect 1910 -1598 1956 -1587
rect 2154 -1598 2200 -1587
rect 1956 -1656 2154 -1610
rect 1910 -1683 1956 -1672
rect 2154 -1683 2200 -1672
rect 2314 -1598 2360 -1518
rect 2459 -1528 2663 -1518
rect 2717 -1455 3078 -1447
rect 2717 -1514 3003 -1455
rect 3066 -1514 3078 -1455
rect 2717 -1528 3078 -1514
rect 3132 -1482 3196 -1366
rect 3354 -1292 3424 -1200
rect 3354 -1366 3377 -1292
rect 3423 -1366 3424 -1292
rect 3354 -1381 3424 -1366
rect 3536 -1292 3600 -1279
rect 3536 -1366 3537 -1292
rect 3583 -1366 3600 -1292
rect 3278 -1455 3482 -1447
rect 3278 -1482 3407 -1455
rect 3132 -1514 3407 -1482
rect 3470 -1514 3482 -1455
rect 3132 -1528 3482 -1514
rect 3536 -1482 3600 -1366
rect 2717 -1529 2894 -1528
rect 3132 -1529 3301 -1528
rect 3536 -1529 3759 -1482
rect 2314 -1683 2360 -1672
rect 2532 -1630 2613 -1625
rect 2717 -1630 2781 -1529
rect 2532 -1676 2554 -1630
rect 2600 -1676 2613 -1630
rect 2711 -1676 2722 -1630
rect 2768 -1676 2781 -1630
rect 2532 -1782 2613 -1676
rect 2717 -1677 2781 -1676
rect 2947 -1630 3028 -1625
rect 3132 -1630 3196 -1529
rect 2947 -1676 2969 -1630
rect 3015 -1676 3028 -1630
rect 3126 -1676 3137 -1630
rect 3183 -1676 3196 -1630
rect 2947 -1782 3028 -1676
rect 3132 -1677 3196 -1676
rect 3351 -1630 3432 -1625
rect 3536 -1630 3600 -1529
rect 3351 -1676 3373 -1630
rect 3419 -1676 3432 -1630
rect 3530 -1676 3541 -1630
rect 3587 -1676 3600 -1630
rect 3351 -1782 3432 -1676
rect 3536 -1677 3600 -1676
rect 51 -1787 3669 -1782
rect -200 -1809 -127 -1800
rect -200 -1863 -191 -1809
rect -137 -1812 -127 -1809
rect 38 -1812 3682 -1787
rect -137 -1817 3682 -1812
rect -137 -1822 1700 -1817
rect -137 -1861 102 -1822
rect -137 -1863 -127 -1861
rect -200 -1873 -127 -1863
rect 38 -1868 102 -1861
rect 1086 -1868 1211 -1822
rect 38 -1871 1211 -1868
rect 1520 -1863 1700 -1822
rect 2407 -1822 3682 -1817
rect 2407 -1863 2504 -1822
rect 1520 -1871 2504 -1863
rect 2813 -1871 2919 -1822
rect 3228 -1871 3323 -1822
rect 3632 -1871 3682 -1822
rect 38 -1900 3682 -1871
rect -823 -1980 -749 -1969
rect 38 -1980 3678 -1946
rect -823 -2036 -812 -1980
rect -756 -1983 3678 -1980
rect -756 -1986 1372 -1983
rect -756 -2036 88 -1986
rect -823 -2046 -749 -2036
rect 38 -2038 88 -2036
rect 787 -2030 1372 -1986
rect 2394 -2030 3678 -1983
rect 787 -2038 3678 -2030
rect 38 -2045 3678 -2038
rect 38 -2064 1250 -2045
rect 137 -2196 183 -2064
rect -499 -2269 -421 -2258
rect 0 -2269 89 -2258
rect -499 -2325 -487 -2269
rect -431 -2271 89 -2269
rect -431 -2325 13 -2271
rect -499 -2334 -421 -2325
rect 0 -2330 13 -2325
rect 76 -2330 89 -2271
rect 137 -2281 183 -2270
rect 297 -2196 343 -2185
rect 541 -2196 587 -2185
rect 343 -2251 541 -2205
rect 297 -2281 343 -2270
rect 0 -2345 89 -2330
rect 541 -2337 587 -2270
rect 701 -2196 747 -2064
rect 846 -2068 1250 -2064
rect 846 -2119 906 -2068
rect 1156 -2119 1250 -2068
rect 846 -2137 1250 -2119
rect 701 -2281 747 -2270
rect 922 -2229 992 -2137
rect 1426 -2197 1472 -2045
rect 1569 -2096 1648 -2094
rect 1569 -2150 1582 -2096
rect 1636 -2150 1648 -2096
rect 1569 -2158 1648 -2150
rect 922 -2303 945 -2229
rect 991 -2303 992 -2229
rect 922 -2318 992 -2303
rect 1104 -2229 1168 -2216
rect 1104 -2303 1105 -2229
rect 1151 -2303 1168 -2229
rect 541 -2383 747 -2337
rect -356 -2411 -275 -2401
rect -356 -2465 -343 -2411
rect -289 -2415 -275 -2411
rect 401 -2415 490 -2406
rect -289 -2419 490 -2415
rect -289 -2461 414 -2419
rect -289 -2465 -275 -2461
rect -356 -2474 -275 -2465
rect 401 -2478 414 -2461
rect 477 -2478 490 -2419
rect 401 -2493 490 -2478
rect 701 -2409 747 -2383
rect 846 -2392 1050 -2384
rect 846 -2409 975 -2392
rect 701 -2451 975 -2409
rect 1038 -2451 1050 -2392
rect 701 -2455 1050 -2451
rect -662 -2551 -583 -2541
rect -15 -2547 67 -2532
rect -15 -2551 2 -2547
rect -662 -2607 -646 -2551
rect -590 -2603 2 -2551
rect 58 -2603 67 -2547
rect -590 -2607 67 -2603
rect -662 -2617 -583 -2607
rect -15 -2623 67 -2607
rect 137 -2535 183 -2524
rect 137 -2719 183 -2609
rect 297 -2535 343 -2524
rect 541 -2535 587 -2524
rect 343 -2593 541 -2547
rect 297 -2620 343 -2609
rect 541 -2620 587 -2609
rect 701 -2535 747 -2455
rect 846 -2465 1050 -2455
rect 1104 -2419 1168 -2303
rect 1253 -2250 1328 -2240
rect 1253 -2251 1329 -2250
rect 1253 -2305 1266 -2251
rect 1320 -2255 1329 -2251
rect 1320 -2305 1373 -2255
rect 1426 -2282 1472 -2271
rect 1586 -2197 1632 -2158
rect 1586 -2282 1632 -2271
rect 1746 -2197 1792 -2045
rect 2455 -2089 3678 -2045
rect 1976 -2094 2050 -2092
rect 1976 -2105 2356 -2094
rect 1976 -2159 1986 -2105
rect 2040 -2140 2356 -2105
rect 2040 -2159 2050 -2140
rect 1976 -2172 2050 -2159
rect 1746 -2282 1792 -2271
rect 1990 -2197 2036 -2172
rect 1990 -2282 2036 -2271
rect 2150 -2197 2196 -2186
rect 1253 -2315 1373 -2305
rect 1327 -2332 1373 -2315
rect 1986 -2332 2075 -2331
rect 1327 -2345 2075 -2332
rect 1327 -2378 1999 -2345
rect 1986 -2404 1999 -2378
rect 2062 -2404 2075 -2345
rect 1986 -2418 2075 -2404
rect 1104 -2464 1281 -2419
rect 1585 -2459 1674 -2446
rect 1104 -2466 1370 -2464
rect 701 -2620 747 -2609
rect 919 -2567 1000 -2562
rect 1104 -2567 1168 -2466
rect 1233 -2467 1370 -2466
rect 1585 -2467 1599 -2459
rect 1233 -2511 1599 -2467
rect 1327 -2513 1599 -2511
rect 1585 -2518 1599 -2513
rect 1662 -2518 1674 -2459
rect 2150 -2494 2196 -2271
rect 2310 -2197 2356 -2140
rect 2455 -2140 2515 -2089
rect 2765 -2140 2930 -2089
rect 3180 -2140 3334 -2089
rect 3584 -2140 3678 -2089
rect 2455 -2158 3678 -2140
rect 2310 -2282 2356 -2271
rect 2531 -2250 2601 -2158
rect 2531 -2324 2554 -2250
rect 2600 -2324 2601 -2250
rect 2531 -2339 2601 -2324
rect 2713 -2250 2777 -2237
rect 2713 -2324 2714 -2250
rect 2760 -2324 2777 -2250
rect 2713 -2405 2777 -2324
rect 2946 -2250 3016 -2158
rect 2946 -2324 2969 -2250
rect 3015 -2324 3016 -2250
rect 2946 -2339 3016 -2324
rect 3128 -2250 3192 -2237
rect 3128 -2324 3129 -2250
rect 3175 -2324 3192 -2250
rect 1585 -2533 1674 -2518
rect 919 -2613 941 -2567
rect 987 -2613 1000 -2567
rect 1098 -2613 1109 -2567
rect 1155 -2613 1168 -2567
rect 1746 -2540 2196 -2494
rect 1746 -2586 1792 -2540
rect 2150 -2546 2196 -2540
rect 2415 -2413 2659 -2405
rect 2415 -2472 2584 -2413
rect 2647 -2472 2659 -2413
rect 2415 -2486 2659 -2472
rect 2713 -2413 3074 -2405
rect 2713 -2472 2999 -2413
rect 3062 -2472 3074 -2413
rect 2713 -2486 3074 -2472
rect 3128 -2440 3192 -2324
rect 3350 -2250 3420 -2158
rect 3350 -2324 3373 -2250
rect 3419 -2324 3420 -2250
rect 3350 -2339 3420 -2324
rect 3532 -2250 3596 -2237
rect 3532 -2324 3533 -2250
rect 3579 -2324 3596 -2250
rect 3274 -2413 3478 -2405
rect 3274 -2440 3403 -2413
rect 3128 -2472 3403 -2440
rect 3466 -2472 3478 -2413
rect 3128 -2486 3478 -2472
rect 3532 -2440 3596 -2324
rect 2415 -2546 2461 -2486
rect 2150 -2586 2461 -2546
rect 2713 -2487 2893 -2486
rect 3128 -2487 3297 -2486
rect 3532 -2487 3761 -2440
rect 38 -2724 846 -2719
rect 919 -2724 1000 -2613
rect 1104 -2614 1168 -2613
rect 1571 -2632 1582 -2586
rect 1628 -2632 1639 -2586
rect 1739 -2632 1750 -2586
rect 1796 -2632 1807 -2586
rect 1975 -2632 1986 -2586
rect 2032 -2632 2043 -2586
rect 2143 -2632 2154 -2586
rect 2200 -2592 2461 -2586
rect 2528 -2588 2609 -2583
rect 2713 -2588 2777 -2487
rect 2200 -2632 2211 -2592
rect -202 -2750 -121 -2738
rect 38 -2745 1250 -2724
rect 1571 -2745 1639 -2632
rect 1975 -2745 2043 -2632
rect 2528 -2634 2550 -2588
rect 2596 -2634 2609 -2588
rect 2707 -2634 2718 -2588
rect 2764 -2634 2777 -2588
rect 2528 -2745 2609 -2634
rect 2713 -2635 2777 -2634
rect 2943 -2588 3024 -2583
rect 3128 -2588 3192 -2487
rect 2943 -2634 2965 -2588
rect 3011 -2634 3024 -2588
rect 3122 -2634 3133 -2588
rect 3179 -2634 3192 -2588
rect 2943 -2745 3024 -2634
rect 3128 -2635 3192 -2634
rect 3347 -2588 3428 -2583
rect 3532 -2588 3596 -2487
rect 3347 -2634 3369 -2588
rect 3415 -2634 3428 -2588
rect 3526 -2634 3537 -2588
rect 3583 -2634 3596 -2588
rect 3347 -2745 3428 -2634
rect 3532 -2635 3596 -2634
rect 38 -2750 3678 -2745
rect -202 -2806 -190 -2750
rect -134 -2754 3678 -2750
rect -134 -2800 87 -2754
rect 794 -2759 3678 -2754
rect 794 -2800 891 -2759
rect -134 -2806 891 -2800
rect -202 -2817 -121 -2806
rect 38 -2808 891 -2806
rect 1200 -2780 3678 -2759
rect 1200 -2808 1391 -2780
rect 38 -2826 1391 -2808
rect 2375 -2826 2500 -2780
rect 38 -2829 2500 -2826
rect 2809 -2829 2915 -2780
rect 3224 -2829 3319 -2780
rect 3628 -2829 3678 -2780
rect 38 -2858 3678 -2829
rect -842 -2925 -744 -2912
rect 38 -2925 2389 -2906
rect -842 -2981 -812 -2925
rect -756 -2943 2389 -2925
rect -756 -2981 83 -2943
rect -842 -2999 -744 -2981
rect 38 -2990 83 -2981
rect 1105 -2990 2389 -2943
rect 38 -3005 2389 -2990
rect 137 -3157 183 -3005
rect 280 -3056 359 -3054
rect 280 -3110 293 -3056
rect 347 -3110 359 -3056
rect 280 -3118 359 -3110
rect 137 -3242 183 -3231
rect 297 -3157 343 -3118
rect 297 -3242 343 -3231
rect 457 -3157 503 -3005
rect 1166 -3049 2389 -3005
rect 687 -3054 761 -3052
rect 687 -3065 1067 -3054
rect 687 -3119 697 -3065
rect 751 -3100 1067 -3065
rect 751 -3119 761 -3100
rect 687 -3132 761 -3119
rect 457 -3242 503 -3231
rect 701 -3157 747 -3132
rect 701 -3242 747 -3231
rect 861 -3157 907 -3146
rect -664 -3288 -582 -3278
rect -664 -3342 -649 -3288
rect -595 -3292 -582 -3288
rect 697 -3292 786 -3291
rect -595 -3305 786 -3292
rect -595 -3338 710 -3305
rect -595 -3342 -582 -3338
rect -664 -3351 -582 -3342
rect 697 -3364 710 -3338
rect 773 -3364 786 -3305
rect 697 -3378 786 -3364
rect -503 -3423 -422 -3413
rect -503 -3477 -490 -3423
rect -436 -3427 -422 -3423
rect 296 -3419 385 -3406
rect 296 -3427 310 -3419
rect -436 -3473 310 -3427
rect -436 -3477 -422 -3473
rect -503 -3488 -422 -3477
rect 296 -3478 310 -3473
rect 373 -3478 385 -3419
rect 861 -3454 907 -3231
rect 1021 -3157 1067 -3100
rect 1166 -3100 1226 -3049
rect 1476 -3100 1641 -3049
rect 1891 -3100 2045 -3049
rect 2295 -3100 2389 -3049
rect 1166 -3118 2389 -3100
rect 1021 -3242 1067 -3231
rect 1242 -3210 1312 -3118
rect 1242 -3284 1265 -3210
rect 1311 -3284 1312 -3210
rect 1242 -3299 1312 -3284
rect 1424 -3210 1488 -3197
rect 1424 -3284 1425 -3210
rect 1471 -3284 1488 -3210
rect 1424 -3365 1488 -3284
rect 1657 -3210 1727 -3118
rect 1657 -3284 1680 -3210
rect 1726 -3284 1727 -3210
rect 1657 -3299 1727 -3284
rect 1839 -3210 1903 -3197
rect 1839 -3284 1840 -3210
rect 1886 -3284 1903 -3210
rect 296 -3493 385 -3478
rect 457 -3500 907 -3454
rect 457 -3546 503 -3500
rect 861 -3506 907 -3500
rect 1126 -3373 1370 -3365
rect 1126 -3432 1295 -3373
rect 1358 -3432 1370 -3373
rect 1126 -3446 1370 -3432
rect 1424 -3373 1785 -3365
rect 1424 -3432 1710 -3373
rect 1773 -3432 1785 -3373
rect 1424 -3446 1785 -3432
rect 1839 -3400 1903 -3284
rect 2061 -3210 2131 -3118
rect 2061 -3284 2084 -3210
rect 2130 -3284 2131 -3210
rect 2061 -3299 2131 -3284
rect 2243 -3210 2307 -3197
rect 2243 -3284 2244 -3210
rect 2290 -3284 2307 -3210
rect 1985 -3373 2189 -3365
rect 1985 -3400 2114 -3373
rect 1839 -3432 2114 -3400
rect 2177 -3432 2189 -3373
rect 1839 -3446 2189 -3432
rect 2243 -3400 2307 -3284
rect 1126 -3506 1172 -3446
rect 861 -3546 1172 -3506
rect 1424 -3447 1604 -3446
rect 1839 -3447 2008 -3446
rect 2243 -3447 2485 -3400
rect 282 -3592 293 -3546
rect 339 -3592 350 -3546
rect 450 -3592 461 -3546
rect 507 -3592 518 -3546
rect 686 -3592 697 -3546
rect 743 -3592 754 -3546
rect 854 -3592 865 -3546
rect 911 -3552 1172 -3546
rect 1239 -3548 1320 -3543
rect 1424 -3548 1488 -3447
rect 911 -3592 922 -3552
rect 282 -3705 350 -3592
rect 686 -3705 754 -3592
rect 1239 -3594 1261 -3548
rect 1307 -3594 1320 -3548
rect 1418 -3594 1429 -3548
rect 1475 -3594 1488 -3548
rect 1239 -3705 1320 -3594
rect 1424 -3595 1488 -3594
rect 1654 -3548 1735 -3543
rect 1839 -3548 1903 -3447
rect 1654 -3594 1676 -3548
rect 1722 -3594 1735 -3548
rect 1833 -3594 1844 -3548
rect 1890 -3594 1903 -3548
rect 1654 -3705 1735 -3594
rect 1839 -3595 1903 -3594
rect 2058 -3548 2139 -3543
rect 2243 -3548 2307 -3447
rect 2058 -3594 2080 -3548
rect 2126 -3594 2139 -3548
rect 2237 -3594 2248 -3548
rect 2294 -3594 2307 -3548
rect 2058 -3705 2139 -3594
rect 2243 -3595 2307 -3594
rect -202 -3742 -127 -3733
rect 38 -3740 2389 -3705
rect 38 -3742 102 -3740
rect -202 -3798 -190 -3742
rect -134 -3786 102 -3742
rect 1086 -3786 1211 -3740
rect -134 -3789 1211 -3786
rect 1520 -3789 1626 -3740
rect 1935 -3789 2030 -3740
rect 2339 -3789 2389 -3740
rect -134 -3798 2389 -3789
rect -202 -3814 -127 -3798
rect 38 -3818 2389 -3798
rect -825 -3896 -750 -3884
rect 38 -3896 4110 -3868
rect -825 -3952 -812 -3896
rect -756 -3905 4110 -3896
rect -756 -3952 83 -3905
rect 1105 -3952 1655 -3905
rect 2677 -3952 4110 -3905
rect -825 -3967 -750 -3952
rect 38 -3967 4110 -3952
rect 137 -4119 183 -3967
rect 280 -4018 359 -4016
rect 280 -4072 293 -4018
rect 347 -4072 359 -4018
rect 280 -4080 359 -4072
rect 137 -4204 183 -4193
rect 297 -4119 343 -4080
rect 297 -4204 343 -4193
rect 457 -4119 503 -3967
rect 1166 -4011 1570 -3967
rect 687 -4016 761 -4014
rect 687 -4027 1067 -4016
rect 687 -4081 697 -4027
rect 751 -4062 1067 -4027
rect 751 -4081 761 -4062
rect 687 -4094 761 -4081
rect 457 -4204 503 -4193
rect 701 -4119 747 -4094
rect 701 -4204 747 -4193
rect 861 -4119 907 -4108
rect -664 -4250 -583 -4241
rect -664 -4304 -651 -4250
rect -597 -4254 -583 -4250
rect 697 -4254 786 -4253
rect -597 -4267 786 -4254
rect -597 -4300 710 -4267
rect -597 -4304 -583 -4300
rect -664 -4315 -583 -4304
rect 697 -4326 710 -4300
rect 773 -4326 786 -4267
rect 697 -4340 786 -4326
rect -508 -4385 -428 -4375
rect -508 -4439 -493 -4385
rect -439 -4389 -428 -4385
rect 296 -4381 385 -4368
rect 296 -4389 310 -4381
rect -439 -4435 310 -4389
rect -439 -4439 -428 -4435
rect -508 -4450 -428 -4439
rect 296 -4440 310 -4435
rect 373 -4440 385 -4381
rect 861 -4416 907 -4193
rect 1021 -4119 1067 -4062
rect 1166 -4062 1226 -4011
rect 1476 -4062 1570 -4011
rect 1166 -4080 1570 -4062
rect 1021 -4204 1067 -4193
rect 1242 -4172 1312 -4080
rect 1709 -4119 1755 -3967
rect 1852 -4018 1931 -4016
rect 1852 -4072 1865 -4018
rect 1919 -4072 1931 -4018
rect 1852 -4080 1931 -4072
rect 1242 -4246 1265 -4172
rect 1311 -4246 1312 -4172
rect 1242 -4261 1312 -4246
rect 1424 -4172 1488 -4159
rect 1424 -4246 1425 -4172
rect 1471 -4246 1488 -4172
rect 296 -4455 385 -4440
rect 457 -4462 907 -4416
rect -355 -4502 -274 -4490
rect 19 -4502 92 -4500
rect -355 -4558 -340 -4502
rect -284 -4512 92 -4502
rect 457 -4508 503 -4462
rect 861 -4468 907 -4462
rect 1126 -4335 1370 -4327
rect 1126 -4394 1295 -4335
rect 1358 -4394 1370 -4335
rect 1126 -4408 1370 -4394
rect 1424 -4362 1488 -4246
rect 1534 -4174 1607 -4163
rect 1534 -4228 1543 -4174
rect 1597 -4228 1607 -4174
rect 1709 -4204 1755 -4193
rect 1869 -4119 1915 -4080
rect 1869 -4204 1915 -4193
rect 2029 -4119 2075 -3967
rect 2738 -4011 4111 -3967
rect 2259 -4016 2333 -4014
rect 2259 -4027 2639 -4016
rect 2259 -4081 2269 -4027
rect 2323 -4062 2639 -4027
rect 2323 -4081 2333 -4062
rect 2259 -4094 2333 -4081
rect 2029 -4204 2075 -4193
rect 2273 -4119 2319 -4094
rect 2273 -4204 2319 -4193
rect 2433 -4119 2479 -4108
rect 1534 -4254 1607 -4228
rect 2269 -4254 2358 -4253
rect 1534 -4255 2358 -4254
rect 1543 -4267 2358 -4255
rect 1543 -4300 2282 -4267
rect 2269 -4326 2282 -4300
rect 2345 -4326 2358 -4267
rect 2269 -4340 2358 -4326
rect 1424 -4389 1604 -4362
rect 1868 -4381 1957 -4368
rect 1868 -4389 1882 -4381
rect 1126 -4468 1172 -4408
rect 861 -4508 1172 -4468
rect 1424 -4409 1882 -4389
rect -284 -4558 30 -4512
rect -355 -4572 -274 -4558
rect 19 -4568 30 -4558
rect 86 -4568 92 -4512
rect 19 -4580 92 -4568
rect 282 -4554 293 -4508
rect 339 -4554 350 -4508
rect 450 -4554 461 -4508
rect 507 -4554 518 -4508
rect 686 -4554 697 -4508
rect 743 -4554 754 -4508
rect 854 -4554 865 -4508
rect 911 -4514 1172 -4508
rect 1239 -4510 1320 -4505
rect 1424 -4510 1488 -4409
rect 1534 -4435 1882 -4409
rect 1868 -4440 1882 -4435
rect 1945 -4440 1957 -4381
rect 2433 -4416 2479 -4193
rect 2593 -4119 2639 -4062
rect 2738 -4062 2798 -4011
rect 3048 -4062 3142 -4011
rect 2738 -4080 3142 -4062
rect 3292 -4062 3363 -4011
rect 3613 -4062 3767 -4011
rect 4017 -4062 4111 -4011
rect 3292 -4080 4111 -4062
rect 2593 -4204 2639 -4193
rect 2814 -4172 2884 -4080
rect 2814 -4246 2837 -4172
rect 2883 -4246 2884 -4172
rect 2814 -4261 2884 -4246
rect 2996 -4172 3060 -4159
rect 2996 -4246 2997 -4172
rect 3043 -4246 3060 -4172
rect 1868 -4455 1957 -4440
rect 2029 -4462 2479 -4416
rect 2029 -4508 2075 -4462
rect 2433 -4468 2479 -4462
rect 2698 -4335 2942 -4327
rect 2698 -4394 2867 -4335
rect 2930 -4394 2942 -4335
rect 2698 -4408 2942 -4394
rect 2996 -4362 3060 -4246
rect 3379 -4172 3449 -4080
rect 3379 -4246 3402 -4172
rect 3448 -4246 3449 -4172
rect 3379 -4261 3449 -4246
rect 3561 -4172 3625 -4159
rect 3561 -4246 3562 -4172
rect 3608 -4246 3625 -4172
rect 3213 -4335 3507 -4327
rect 3213 -4362 3432 -4335
rect 2996 -4394 3432 -4362
rect 3495 -4394 3507 -4335
rect 2996 -4408 3507 -4394
rect 3561 -4362 3625 -4246
rect 3783 -4172 3853 -4080
rect 3783 -4246 3806 -4172
rect 3852 -4246 3853 -4172
rect 3783 -4261 3853 -4246
rect 3965 -4172 4029 -4159
rect 3965 -4246 3966 -4172
rect 4012 -4246 4029 -4172
rect 3707 -4335 3911 -4327
rect 3707 -4362 3836 -4335
rect 3561 -4394 3836 -4362
rect 3899 -4394 3911 -4335
rect 3561 -4408 3911 -4394
rect 3965 -4362 4029 -4246
rect 2698 -4468 2744 -4408
rect 2433 -4508 2744 -4468
rect 2996 -4409 3244 -4408
rect 3561 -4409 3730 -4408
rect 3965 -4409 4210 -4362
rect 911 -4554 922 -4514
rect -204 -4670 -124 -4658
rect 282 -4667 350 -4554
rect 686 -4667 754 -4554
rect 1239 -4556 1261 -4510
rect 1307 -4556 1320 -4510
rect 1418 -4556 1429 -4510
rect 1475 -4556 1488 -4510
rect 1239 -4667 1320 -4556
rect 1424 -4557 1488 -4556
rect 1854 -4554 1865 -4508
rect 1911 -4554 1922 -4508
rect 2022 -4554 2033 -4508
rect 2079 -4554 2090 -4508
rect 2258 -4554 2269 -4508
rect 2315 -4554 2326 -4508
rect 2426 -4554 2437 -4508
rect 2483 -4514 2744 -4508
rect 2811 -4510 2892 -4505
rect 2996 -4510 3060 -4409
rect 2483 -4554 2494 -4514
rect 1854 -4667 1922 -4554
rect 2258 -4667 2326 -4554
rect 2811 -4556 2833 -4510
rect 2879 -4556 2892 -4510
rect 2990 -4556 3001 -4510
rect 3047 -4556 3060 -4510
rect 2811 -4667 2892 -4556
rect 2996 -4557 3060 -4556
rect 3376 -4510 3457 -4505
rect 3561 -4510 3625 -4409
rect 3376 -4556 3398 -4510
rect 3444 -4556 3457 -4510
rect 3555 -4556 3566 -4510
rect 3612 -4556 3625 -4510
rect 3376 -4667 3457 -4556
rect 3561 -4557 3625 -4556
rect 3780 -4510 3861 -4505
rect 3965 -4510 4029 -4409
rect 3780 -4556 3802 -4510
rect 3848 -4556 3861 -4510
rect 3959 -4556 3970 -4510
rect 4016 -4556 4029 -4510
rect 3780 -4667 3861 -4556
rect 3965 -4557 4029 -4556
rect 38 -4670 4111 -4667
rect -204 -4726 -190 -4670
rect -134 -4702 4111 -4670
rect -134 -4726 102 -4702
rect -204 -4742 -124 -4726
rect 38 -4748 102 -4726
rect 1086 -4748 1211 -4702
rect 38 -4751 1211 -4748
rect 1520 -4748 1674 -4702
rect 2658 -4748 2783 -4702
rect 1520 -4751 2783 -4748
rect 3092 -4751 3348 -4702
rect 3657 -4751 3752 -4702
rect 4061 -4751 4111 -4702
rect 38 -4780 4111 -4751
<< via1 >>
rect -812 791 -756 847
rect -646 520 -590 576
rect -480 372 -426 426
rect 0 243 56 299
rect 1373 507 1436 566
rect -189 46 -135 100
rect -812 -140 -756 -84
rect -646 -431 -590 -375
rect 7 -430 13 -376
rect 13 -430 61 -376
rect -491 -567 -437 -513
rect 2399 -565 2455 -509
rect 3340 -400 3396 -344
rect 2382 -707 2436 -653
rect -190 -910 -134 -854
rect -812 -1069 -756 -1013
rect -646 -1249 -591 -1194
rect -48 -1251 9 -1194
rect 293 -1192 347 -1138
rect 697 -1201 751 -1147
rect -491 -1424 -437 -1370
rect -344 -1559 -290 -1505
rect 1626 -1393 1689 -1334
rect -191 -1863 -137 -1809
rect -812 -2036 -756 -1980
rect -487 -2325 -431 -2269
rect 1582 -2150 1636 -2096
rect -343 -2465 -289 -2411
rect -646 -2607 -590 -2551
rect 2 -2603 58 -2547
rect 1266 -2305 1320 -2251
rect 1986 -2159 2040 -2105
rect -190 -2806 -134 -2750
rect -812 -2981 -756 -2925
rect 293 -3110 347 -3056
rect 697 -3119 751 -3065
rect -649 -3342 -595 -3288
rect -490 -3477 -436 -3423
rect -190 -3798 -134 -3742
rect -812 -3952 -756 -3896
rect 293 -4072 347 -4018
rect 697 -4081 751 -4027
rect -651 -4304 -597 -4250
rect -493 -4439 -439 -4385
rect 1865 -4072 1919 -4018
rect -340 -4558 -284 -4502
rect 1543 -4228 1597 -4174
rect 2269 -4081 2323 -4027
rect 30 -4568 86 -4512
rect -190 -4726 -134 -4670
<< metal2 >>
rect -821 847 -747 856
rect -821 791 -812 847
rect -756 791 -747 847
rect -821 781 -747 791
rect -812 -75 -756 781
rect -655 576 -581 585
rect -655 520 -646 576
rect -590 520 -581 576
rect -655 511 -581 520
rect 200 566 1449 579
rect 200 523 1373 566
rect -822 -84 -748 -75
rect -822 -140 -812 -84
rect -756 -140 -748 -84
rect -822 -149 -748 -140
rect -812 -1005 -756 -149
rect -646 -363 -590 511
rect -489 426 -417 435
rect -489 372 -480 426
rect -426 372 -417 426
rect -489 363 -417 372
rect -658 -375 -587 -363
rect -658 -431 -646 -375
rect -590 -431 -587 -375
rect -658 -443 -587 -431
rect -825 -1013 -747 -1005
rect -825 -1069 -812 -1013
rect -756 -1069 -747 -1013
rect -825 -1081 -747 -1069
rect -812 -1969 -756 -1081
rect -646 -1187 -590 -443
rect -487 -504 -431 363
rect -12 299 68 308
rect 200 299 256 523
rect 1329 521 1373 523
rect 1360 507 1373 521
rect 1436 507 1449 566
rect 1360 492 1449 507
rect -340 243 0 299
rect 56 243 256 299
rect -500 -513 -428 -504
rect -500 -567 -491 -513
rect -437 -567 -428 -513
rect -500 -576 -428 -567
rect -658 -1194 -583 -1187
rect -658 -1249 -646 -1194
rect -591 -1249 -583 -1194
rect -658 -1260 -583 -1249
rect -823 -1980 -749 -1969
rect -823 -2036 -812 -1980
rect -756 -2036 -749 -1980
rect -823 -2046 -749 -2036
rect -812 -2912 -756 -2046
rect -646 -2541 -590 -1260
rect -487 -1361 -431 -576
rect -502 -1370 -424 -1361
rect -502 -1424 -491 -1370
rect -437 -1424 -424 -1370
rect -502 -1433 -424 -1424
rect -487 -2258 -431 -1433
rect -340 -1496 -284 243
rect -12 234 68 243
rect -198 100 -126 109
rect -198 46 -189 100
rect -135 46 -126 100
rect -198 37 -126 46
rect -190 -846 -134 37
rect 6 -312 2455 -256
rect 6 -370 62 -312
rect -21 -376 73 -370
rect -21 -430 7 -376
rect 61 -430 73 -376
rect -21 -446 73 -430
rect 2399 -501 2455 -312
rect 3333 -344 3410 -329
rect 2648 -400 3340 -344
rect 3396 -400 3410 -344
rect 2380 -509 2466 -501
rect 2380 -565 2399 -509
rect 2455 -565 2466 -509
rect 2380 -577 2466 -565
rect 2358 -652 2452 -635
rect 2648 -652 2704 -400
rect 3333 -414 3410 -400
rect 2358 -653 2704 -652
rect 2358 -707 2382 -653
rect 2436 -707 2704 -653
rect 2358 -708 2704 -707
rect 2358 -726 2452 -708
rect -201 -854 -127 -846
rect -201 -910 -190 -854
rect -134 -910 -127 -854
rect -201 -918 -127 -910
rect -354 -1505 -274 -1496
rect -354 -1559 -344 -1505
rect -290 -1559 -274 -1505
rect -354 -1569 -274 -1559
rect -499 -2269 -421 -2258
rect -499 -2325 -487 -2269
rect -431 -2325 -421 -2269
rect -499 -2334 -421 -2325
rect -662 -2551 -583 -2541
rect -662 -2607 -646 -2551
rect -590 -2607 -583 -2551
rect -662 -2617 -583 -2607
rect -842 -2925 -744 -2912
rect -842 -2981 -812 -2925
rect -756 -2981 -744 -2925
rect -842 -2999 -744 -2981
rect -812 -3884 -756 -2999
rect -646 -3278 -590 -2617
rect -664 -3288 -582 -3278
rect -664 -3342 -649 -3288
rect -595 -3342 -582 -3288
rect -664 -3351 -582 -3342
rect -825 -3896 -750 -3884
rect -825 -3952 -812 -3896
rect -756 -3952 -750 -3896
rect -825 -3967 -750 -3952
rect -646 -4241 -590 -3351
rect -487 -3413 -431 -2334
rect -340 -2401 -284 -1569
rect -190 -1800 -134 -918
rect 277 -1136 361 -1126
rect 687 -1136 761 -1134
rect 277 -1138 761 -1136
rect -57 -1194 19 -1185
rect 277 -1192 293 -1138
rect 347 -1147 761 -1138
rect 347 -1192 697 -1147
rect -57 -1251 -48 -1194
rect 9 -1251 130 -1194
rect 277 -1209 361 -1192
rect 687 -1201 697 -1192
rect 751 -1201 761 -1147
rect 687 -1214 761 -1201
rect -57 -1260 130 -1251
rect 73 -1332 130 -1260
rect 1613 -1332 1702 -1321
rect 73 -1334 1702 -1332
rect 73 -1389 1626 -1334
rect 1613 -1393 1626 -1389
rect 1689 -1393 1702 -1334
rect 1613 -1408 1702 -1393
rect -200 -1809 -127 -1800
rect -200 -1863 -191 -1809
rect -137 -1863 -127 -1809
rect -200 -1873 -127 -1863
rect -356 -2411 -275 -2401
rect -356 -2465 -343 -2411
rect -289 -2465 -275 -2411
rect -356 -2474 -275 -2465
rect -503 -3423 -422 -3413
rect -503 -3477 -490 -3423
rect -436 -3477 -422 -3423
rect -503 -3488 -422 -3477
rect -664 -4250 -583 -4241
rect -664 -4304 -651 -4250
rect -597 -4304 -583 -4250
rect -664 -4315 -583 -4304
rect -487 -4371 -431 -3488
rect -509 -4385 -426 -4371
rect -509 -4439 -493 -4385
rect -439 -4439 -426 -4385
rect -509 -4453 -426 -4439
rect -340 -4490 -284 -2474
rect -190 -2738 -134 -1873
rect 1566 -2094 1650 -2084
rect 1976 -2094 2050 -2092
rect 1566 -2096 2050 -2094
rect 1566 -2150 1582 -2096
rect 1636 -2105 2050 -2096
rect 1636 -2150 1986 -2105
rect 1566 -2167 1650 -2150
rect 1976 -2159 1986 -2150
rect 2040 -2159 2050 -2105
rect 1976 -2172 2050 -2159
rect 1253 -2250 1328 -2240
rect 258 -2251 1328 -2250
rect 258 -2305 1266 -2251
rect 1320 -2305 1328 -2251
rect 258 -2306 1328 -2305
rect -15 -2547 67 -2532
rect 258 -2547 314 -2306
rect 1253 -2315 1328 -2306
rect -15 -2603 2 -2547
rect 58 -2603 314 -2547
rect -15 -2623 67 -2603
rect -202 -2750 -121 -2738
rect -202 -2806 -190 -2750
rect -134 -2806 -121 -2750
rect -202 -2817 -121 -2806
rect -190 -3733 -134 -2817
rect 277 -3054 361 -3044
rect 687 -3054 761 -3052
rect 277 -3056 761 -3054
rect 277 -3110 293 -3056
rect 347 -3065 761 -3056
rect 347 -3110 697 -3065
rect 277 -3127 361 -3110
rect 687 -3119 697 -3110
rect 751 -3119 761 -3065
rect 687 -3132 761 -3119
rect -202 -3742 -127 -3733
rect -202 -3798 -190 -3742
rect -134 -3798 -127 -3742
rect -202 -3814 -127 -3798
rect -355 -4502 -274 -4490
rect -355 -4558 -340 -4502
rect -284 -4558 -274 -4502
rect -355 -4572 -274 -4558
rect -190 -4658 -134 -3814
rect 277 -4016 361 -4006
rect 687 -4016 761 -4014
rect 277 -4018 761 -4016
rect 277 -4072 293 -4018
rect 347 -4027 761 -4018
rect 347 -4072 697 -4027
rect 277 -4089 361 -4072
rect 687 -4081 697 -4072
rect 751 -4081 761 -4027
rect 687 -4094 761 -4081
rect 1849 -4016 1933 -4006
rect 2259 -4016 2333 -4014
rect 1849 -4018 2333 -4016
rect 1849 -4072 1865 -4018
rect 1919 -4027 2333 -4018
rect 1919 -4072 2269 -4027
rect 1849 -4089 1933 -4072
rect 2259 -4081 2269 -4072
rect 2323 -4081 2333 -4027
rect 2259 -4094 2333 -4081
rect 1533 -4174 1607 -4163
rect 1533 -4200 1543 -4174
rect 261 -4228 1543 -4200
rect 1597 -4228 1607 -4174
rect 261 -4255 1607 -4228
rect 261 -4256 1570 -4255
rect 19 -4512 92 -4500
rect 261 -4512 317 -4256
rect 19 -4568 30 -4512
rect 86 -4568 317 -4512
rect 19 -4580 92 -4568
rect -204 -4670 -124 -4658
rect -204 -4726 -190 -4670
rect -134 -4726 -124 -4670
rect -204 -4742 -124 -4726
<< labels >>
flabel metal1 34 536 34 536 0 FreeSans 640 0 0 0 B1
port 0 nsew
flabel metal1 4 398 4 398 0 FreeSans 640 0 0 0 B2
port 1 nsew
flabel via1 18 270 18 270 0 FreeSans 640 0 0 0 B3
port 2 nsew
flabel metal1 1320 841 1320 841 0 FreeSans 640 0 0 0 VDD
port 3 nsew
flabel metal1 1314 46 1314 46 0 FreeSans 640 0 0 0 VSS
port 4 nsew
flabel metal1 3562 396 3562 396 0 FreeSans 640 0 0 0 D1
port 5 nsew
flabel via1 3367 -373 3367 -373 0 FreeSans 640 0 0 0 D2
port 6 nsew
flabel metal1 3372 -543 3372 -543 0 FreeSans 640 0 0 0 D4
port 7 nsew
flabel metal1 3741 -1506 3741 -1506 0 FreeSans 640 0 0 0 D3
port 8 nsew
flabel metal1 3737 -2461 3737 -2461 0 FreeSans 640 0 0 0 D5
port 9 nsew
flabel metal1 2471 -3426 2471 -3426 0 FreeSans 640 0 0 0 D6
port 11 nsew
flabel metal1 4200 -4382 4200 -4382 0 FreeSans 640 0 0 0 D7
port 12 nsew
flabel metal1 1532 -3411 1532 -3411 0 FreeSans 640 0 0 0 INV_BUFF_5.IN
flabel metal1 2423 -3425 2423 -3425 0 FreeSans 640 0 0 0 INV_BUFF_5.OUT
flabel metal1 1961 -3058 1961 -3058 0 FreeSans 640 0 0 0 INV_BUFF_5.VDD
flabel metal1 1981 -3778 1981 -3778 0 FreeSans 640 0 0 0 INV_BUFF_5.VSS
flabel nsubdiffcont 2170 -3074 2170 -3074 0 FreeSans 640 0 0 0 INV_BUFF_5.Inverter_0.VDD
flabel psubdiffcont 2184 -3766 2184 -3766 0 FreeSans 640 0 0 0 INV_BUFF_5.Inverter_0.VSS
flabel metal1 2008 -3405 2008 -3405 0 FreeSans 640 0 0 0 INV_BUFF_5.Inverter_0.IN
flabel metal1 2375 -3432 2375 -3432 0 FreeSans 640 0 0 0 INV_BUFF_5.Inverter_0.OUT
flabel nsubdiffcont 1766 -3074 1766 -3074 0 FreeSans 640 0 0 0 INV_BUFF_5.Inverter_1.VDD
flabel psubdiffcont 1780 -3766 1780 -3766 0 FreeSans 640 0 0 0 INV_BUFF_5.Inverter_1.VSS
flabel metal1 1604 -3405 1604 -3405 0 FreeSans 640 0 0 0 INV_BUFF_5.Inverter_1.IN
flabel metal1 1971 -3432 1971 -3432 0 FreeSans 640 0 0 0 INV_BUFF_5.Inverter_1.OUT
flabel nsubdiffcont 381 -2021 451 -1998 0 FreeSans 640 0 0 0 AND_4.VDD
flabel psubdiffcont 422 -2788 492 -2765 0 FreeSans 640 0 0 0 AND_4.VSS
flabel metal1 39 -2445 109 -2422 0 FreeSans 640 0 0 0 AND_4.B
flabel polycontact 38 -2300 38 -2300 0 FreeSans 640 0 0 0 AND_4.A
flabel metal1 1258 -2440 1258 -2440 0 FreeSans 640 0 0 0 AND_4.OUT
flabel nsubdiffcont 1031 -2093 1031 -2093 0 FreeSans 640 0 0 0 AND_4.Inverter_0.VDD
flabel psubdiffcont 1045 -2785 1045 -2785 0 FreeSans 640 0 0 0 AND_4.Inverter_0.VSS
flabel metal1 869 -2424 869 -2424 0 FreeSans 640 0 0 0 AND_4.Inverter_0.IN
flabel metal1 1236 -2451 1236 -2451 0 FreeSans 640 0 0 0 AND_4.Inverter_0.OUT
flabel metal1 2821 -2451 2821 -2451 0 FreeSans 640 0 0 0 INV_BUFF_4.IN
flabel metal1 3712 -2465 3712 -2465 0 FreeSans 640 0 0 0 INV_BUFF_4.OUT
flabel metal1 3250 -2098 3250 -2098 0 FreeSans 640 0 0 0 INV_BUFF_4.VDD
flabel metal1 3270 -2818 3270 -2818 0 FreeSans 640 0 0 0 INV_BUFF_4.VSS
flabel nsubdiffcont 3459 -2114 3459 -2114 0 FreeSans 640 0 0 0 INV_BUFF_4.Inverter_0.VDD
flabel psubdiffcont 3473 -2806 3473 -2806 0 FreeSans 640 0 0 0 INV_BUFF_4.Inverter_0.VSS
flabel metal1 3297 -2445 3297 -2445 0 FreeSans 640 0 0 0 INV_BUFF_4.Inverter_0.IN
flabel metal1 3664 -2472 3664 -2472 0 FreeSans 640 0 0 0 INV_BUFF_4.Inverter_0.OUT
flabel nsubdiffcont 3055 -2114 3055 -2114 0 FreeSans 640 0 0 0 INV_BUFF_4.Inverter_1.VDD
flabel psubdiffcont 3069 -2806 3069 -2806 0 FreeSans 640 0 0 0 INV_BUFF_4.Inverter_1.VSS
flabel metal1 2893 -2445 2893 -2445 0 FreeSans 640 0 0 0 INV_BUFF_4.Inverter_1.IN
flabel metal1 3260 -2472 3260 -2472 0 FreeSans 640 0 0 0 INV_BUFF_4.Inverter_1.OUT
flabel nsubdiffcont 1994 -1084 2064 -1061 0 FreeSans 640 0 0 0 AND_3.VDD
flabel psubdiffcont 2035 -1851 2105 -1828 0 FreeSans 640 0 0 0 AND_3.VSS
flabel metal1 1652 -1508 1722 -1485 0 FreeSans 640 0 0 0 AND_3.B
flabel polycontact 1651 -1363 1651 -1363 0 FreeSans 640 0 0 0 AND_3.A
flabel metal1 2871 -1503 2871 -1503 0 FreeSans 640 0 0 0 AND_3.OUT
flabel nsubdiffcont 2644 -1156 2644 -1156 0 FreeSans 640 0 0 0 AND_3.Inverter_0.VDD
flabel psubdiffcont 2658 -1848 2658 -1848 0 FreeSans 640 0 0 0 AND_3.Inverter_0.VSS
flabel metal1 2482 -1487 2482 -1487 0 FreeSans 640 0 0 0 AND_3.Inverter_0.IN
flabel metal1 2849 -1514 2849 -1514 0 FreeSans 640 0 0 0 AND_3.Inverter_0.OUT
flabel metal1 2825 -1493 2825 -1493 0 FreeSans 640 0 0 0 INV_BUFF_2.IN
flabel metal1 3716 -1507 3716 -1507 0 FreeSans 640 0 0 0 INV_BUFF_2.OUT
flabel metal1 3254 -1140 3254 -1140 0 FreeSans 640 0 0 0 INV_BUFF_2.VDD
flabel metal1 3274 -1860 3274 -1860 0 FreeSans 640 0 0 0 INV_BUFF_2.VSS
flabel nsubdiffcont 3463 -1156 3463 -1156 0 FreeSans 640 0 0 0 INV_BUFF_2.Inverter_0.VDD
flabel psubdiffcont 3477 -1848 3477 -1848 0 FreeSans 640 0 0 0 INV_BUFF_2.Inverter_0.VSS
flabel metal1 3301 -1487 3301 -1487 0 FreeSans 640 0 0 0 INV_BUFF_2.Inverter_0.IN
flabel metal1 3668 -1514 3668 -1514 0 FreeSans 640 0 0 0 INV_BUFF_2.Inverter_0.OUT
flabel nsubdiffcont 3059 -1156 3059 -1156 0 FreeSans 640 0 0 0 INV_BUFF_2.Inverter_1.VDD
flabel psubdiffcont 3073 -1848 3073 -1848 0 FreeSans 640 0 0 0 INV_BUFF_2.Inverter_1.VSS
flabel metal1 2897 -1487 2897 -1487 0 FreeSans 640 0 0 0 INV_BUFF_2.Inverter_1.IN
flabel metal1 3264 -1514 3264 -1514 0 FreeSans 640 0 0 0 INV_BUFF_2.Inverter_1.OUT
flabel nsubdiffcont 381 -123 451 -100 0 FreeSans 640 0 0 0 AND_2.VDD
flabel psubdiffcont 422 -890 492 -867 0 FreeSans 640 0 0 0 AND_2.VSS
flabel metal1 39 -547 109 -524 0 FreeSans 640 0 0 0 AND_2.B
flabel polycontact 38 -402 38 -402 0 FreeSans 640 0 0 0 AND_2.A
flabel metal1 1258 -542 1258 -542 0 FreeSans 640 0 0 0 AND_2.OUT
flabel nsubdiffcont 1031 -195 1031 -195 0 FreeSans 640 0 0 0 AND_2.Inverter_0.VDD
flabel psubdiffcont 1045 -887 1045 -887 0 FreeSans 640 0 0 0 AND_2.Inverter_0.VSS
flabel metal1 869 -526 869 -526 0 FreeSans 640 0 0 0 AND_2.Inverter_0.IN
flabel metal1 1236 -553 1236 -553 0 FreeSans 640 0 0 0 AND_2.Inverter_0.OUT
flabel metal1 1322 -532 1322 -532 0 FreeSans 640 0 0 0 INV_BUFF_1.IN
flabel metal1 2213 -546 2213 -546 0 FreeSans 640 0 0 0 INV_BUFF_1.OUT
flabel metal1 1751 -179 1751 -179 0 FreeSans 640 0 0 0 INV_BUFF_1.VDD
flabel metal1 1771 -899 1771 -899 0 FreeSans 640 0 0 0 INV_BUFF_1.VSS
flabel nsubdiffcont 1960 -195 1960 -195 0 FreeSans 640 0 0 0 INV_BUFF_1.Inverter_0.VDD
flabel psubdiffcont 1974 -887 1974 -887 0 FreeSans 640 0 0 0 INV_BUFF_1.Inverter_0.VSS
flabel metal1 1798 -526 1798 -526 0 FreeSans 640 0 0 0 INV_BUFF_1.Inverter_0.IN
flabel metal1 2165 -553 2165 -553 0 FreeSans 640 0 0 0 INV_BUFF_1.Inverter_0.OUT
flabel nsubdiffcont 1556 -195 1556 -195 0 FreeSans 640 0 0 0 INV_BUFF_1.Inverter_1.VDD
flabel psubdiffcont 1570 -887 1570 -887 0 FreeSans 640 0 0 0 INV_BUFF_1.Inverter_1.VSS
flabel metal1 1394 -526 1394 -526 0 FreeSans 640 0 0 0 INV_BUFF_1.Inverter_1.IN
flabel metal1 1761 -553 1761 -553 0 FreeSans 640 0 0 0 INV_BUFF_1.Inverter_1.OUT
flabel metal1 2454 -532 2454 -532 0 FreeSans 640 0 0 0 INV_BUFF_3.IN
flabel metal1 3345 -546 3345 -546 0 FreeSans 640 0 0 0 INV_BUFF_3.OUT
flabel metal1 2883 -179 2883 -179 0 FreeSans 640 0 0 0 INV_BUFF_3.VDD
flabel metal1 2903 -899 2903 -899 0 FreeSans 640 0 0 0 INV_BUFF_3.VSS
flabel nsubdiffcont 3092 -195 3092 -195 0 FreeSans 640 0 0 0 INV_BUFF_3.Inverter_0.VDD
flabel psubdiffcont 3106 -887 3106 -887 0 FreeSans 640 0 0 0 INV_BUFF_3.Inverter_0.VSS
flabel metal1 2930 -526 2930 -526 0 FreeSans 640 0 0 0 INV_BUFF_3.Inverter_0.IN
flabel metal1 3297 -553 3297 -553 0 FreeSans 640 0 0 0 INV_BUFF_3.Inverter_0.OUT
flabel nsubdiffcont 2688 -195 2688 -195 0 FreeSans 640 0 0 0 INV_BUFF_3.Inverter_1.VDD
flabel psubdiffcont 2702 -887 2702 -887 0 FreeSans 640 0 0 0 INV_BUFF_3.Inverter_1.VSS
flabel metal1 2526 -526 2526 -526 0 FreeSans 640 0 0 0 INV_BUFF_3.Inverter_1.IN
flabel metal1 2893 -553 2893 -553 0 FreeSans 640 0 0 0 INV_BUFF_3.Inverter_1.OUT
flabel nsubdiffcont 1741 816 1811 839 0 FreeSans 640 0 0 0 AND_0.VDD
flabel psubdiffcont 1782 49 1852 72 0 FreeSans 640 0 0 0 AND_0.VSS
flabel metal1 1399 392 1469 415 0 FreeSans 640 0 0 0 AND_0.B
flabel polycontact 1398 537 1398 537 0 FreeSans 640 0 0 0 AND_0.A
flabel metal1 2618 397 2618 397 0 FreeSans 640 0 0 0 AND_0.OUT
flabel nsubdiffcont 2391 744 2391 744 0 FreeSans 640 0 0 0 AND_0.Inverter_0.VDD
flabel psubdiffcont 2405 52 2405 52 0 FreeSans 640 0 0 0 AND_0.Inverter_0.VSS
flabel metal1 2229 413 2229 413 0 FreeSans 640 0 0 0 AND_0.Inverter_0.IN
flabel metal1 2596 386 2596 386 0 FreeSans 640 0 0 0 AND_0.Inverter_0.OUT
flabel nsubdiffcont 381 816 451 839 0 FreeSans 640 0 0 0 AND_1.VDD
flabel psubdiffcont 422 49 492 72 0 FreeSans 640 0 0 0 AND_1.VSS
flabel metal1 39 392 109 415 0 FreeSans 640 0 0 0 AND_1.B
flabel polycontact 38 537 38 537 0 FreeSans 640 0 0 0 AND_1.A
flabel metal1 1258 397 1258 397 0 FreeSans 640 0 0 0 AND_1.OUT
flabel nsubdiffcont 1031 744 1031 744 0 FreeSans 640 0 0 0 AND_1.Inverter_0.VDD
flabel psubdiffcont 1045 52 1045 52 0 FreeSans 640 0 0 0 AND_1.Inverter_0.VSS
flabel metal1 869 413 869 413 0 FreeSans 640 0 0 0 AND_1.Inverter_0.IN
flabel metal1 1236 386 1236 386 0 FreeSans 640 0 0 0 AND_1.Inverter_0.OUT
flabel metal1 2651 407 2651 407 0 FreeSans 640 0 0 0 INV_BUFF_0.IN
flabel metal1 3542 393 3542 393 0 FreeSans 640 0 0 0 INV_BUFF_0.OUT
flabel metal1 3080 760 3080 760 0 FreeSans 640 0 0 0 INV_BUFF_0.VDD
flabel metal1 3100 40 3100 40 0 FreeSans 640 0 0 0 INV_BUFF_0.VSS
flabel nsubdiffcont 3289 744 3289 744 0 FreeSans 640 0 0 0 INV_BUFF_0.Inverter_0.VDD
flabel psubdiffcont 3303 52 3303 52 0 FreeSans 640 0 0 0 INV_BUFF_0.Inverter_0.VSS
flabel metal1 3127 413 3127 413 0 FreeSans 640 0 0 0 INV_BUFF_0.Inverter_0.IN
flabel metal1 3494 386 3494 386 0 FreeSans 640 0 0 0 INV_BUFF_0.Inverter_0.OUT
flabel nsubdiffcont 2885 744 2885 744 0 FreeSans 640 0 0 0 INV_BUFF_0.Inverter_1.VDD
flabel psubdiffcont 2899 52 2899 52 0 FreeSans 640 0 0 0 INV_BUFF_0.Inverter_1.VSS
flabel metal1 2723 413 2723 413 0 FreeSans 640 0 0 0 INV_BUFF_0.Inverter_1.IN
flabel metal1 3090 386 3090 386 0 FreeSans 640 0 0 0 INV_BUFF_0.Inverter_1.OUT
flabel metal1 51 -1397 51 -1397 0 FreeSans 640 0 0 0 OR_0.A
flabel metal1 59 -1533 59 -1533 0 FreeSans 640 0 0 0 OR_0.B
flabel psubdiffcont 594 -1844 594 -1844 0 FreeSans 640 0 0 0 OR_0.VSS
flabel nsubdiffcont 593 -1047 593 -1047 0 FreeSans 640 0 0 0 OR_0.VDD
flabel metal1 1580 -1511 1580 -1511 0 FreeSans 640 0 0 0 OR_0.OUT
flabel nsubdiffcont 1351 -1156 1351 -1156 0 FreeSans 640 0 0 0 OR_0.Inverter_0.VDD
flabel psubdiffcont 1365 -1848 1365 -1848 0 FreeSans 640 0 0 0 OR_0.Inverter_0.VSS
flabel metal1 1189 -1487 1189 -1487 0 FreeSans 640 0 0 0 OR_0.Inverter_0.IN
flabel metal1 1556 -1514 1556 -1514 0 FreeSans 640 0 0 0 OR_0.Inverter_0.OUT
flabel metal1 1340 -2355 1340 -2355 0 FreeSans 640 0 0 0 OR_1.A
flabel metal1 1348 -2491 1348 -2491 0 FreeSans 640 0 0 0 OR_1.B
flabel psubdiffcont 1883 -2802 1883 -2802 0 FreeSans 640 0 0 0 OR_1.VSS
flabel nsubdiffcont 1882 -2005 1882 -2005 0 FreeSans 640 0 0 0 OR_1.VDD
flabel metal1 2869 -2469 2869 -2469 0 FreeSans 640 0 0 0 OR_1.OUT
flabel nsubdiffcont 2640 -2114 2640 -2114 0 FreeSans 640 0 0 0 OR_1.Inverter_0.VDD
flabel psubdiffcont 2654 -2806 2654 -2806 0 FreeSans 640 0 0 0 OR_1.Inverter_0.VSS
flabel metal1 2478 -2445 2478 -2445 0 FreeSans 640 0 0 0 OR_1.Inverter_0.IN
flabel metal1 2845 -2472 2845 -2472 0 FreeSans 640 0 0 0 OR_1.Inverter_0.OUT
flabel metal1 51 -3315 51 -3315 0 FreeSans 640 0 0 0 OR_2.A
flabel metal1 59 -3451 59 -3451 0 FreeSans 640 0 0 0 OR_2.B
flabel psubdiffcont 594 -3762 594 -3762 0 FreeSans 640 0 0 0 OR_2.VSS
flabel nsubdiffcont 593 -2965 593 -2965 0 FreeSans 640 0 0 0 OR_2.VDD
flabel metal1 1580 -3429 1580 -3429 0 FreeSans 640 0 0 0 OR_2.OUT
flabel nsubdiffcont 1351 -3074 1351 -3074 0 FreeSans 640 0 0 0 OR_2.Inverter_0.VDD
flabel psubdiffcont 1365 -3766 1365 -3766 0 FreeSans 640 0 0 0 OR_2.Inverter_0.VSS
flabel metal1 1189 -3405 1189 -3405 0 FreeSans 640 0 0 0 OR_2.Inverter_0.IN
flabel metal1 1556 -3432 1556 -3432 0 FreeSans 640 0 0 0 OR_2.Inverter_0.OUT
flabel metal1 1623 -4277 1623 -4277 0 FreeSans 640 0 0 0 OR_3.A
flabel metal1 1631 -4413 1631 -4413 0 FreeSans 640 0 0 0 OR_3.B
flabel psubdiffcont 2166 -4724 2166 -4724 0 FreeSans 640 0 0 0 OR_3.VSS
flabel nsubdiffcont 2165 -3927 2165 -3927 0 FreeSans 640 0 0 0 OR_3.VDD
flabel metal1 3152 -4391 3152 -4391 0 FreeSans 640 0 0 0 OR_3.OUT
flabel nsubdiffcont 2923 -4036 2923 -4036 0 FreeSans 640 0 0 0 OR_3.Inverter_0.VDD
flabel psubdiffcont 2937 -4728 2937 -4728 0 FreeSans 640 0 0 0 OR_3.Inverter_0.VSS
flabel metal1 2761 -4367 2761 -4367 0 FreeSans 640 0 0 0 OR_3.Inverter_0.IN
flabel metal1 3128 -4394 3128 -4394 0 FreeSans 640 0 0 0 OR_3.Inverter_0.OUT
flabel metal1 51 -4277 51 -4277 0 FreeSans 640 0 0 0 OR_4.A
flabel metal1 59 -4413 59 -4413 0 FreeSans 640 0 0 0 OR_4.B
flabel psubdiffcont 594 -4724 594 -4724 0 FreeSans 640 0 0 0 OR_4.VSS
flabel nsubdiffcont 593 -3927 593 -3927 0 FreeSans 640 0 0 0 OR_4.VDD
flabel metal1 1580 -4391 1580 -4391 0 FreeSans 640 0 0 0 OR_4.OUT
flabel nsubdiffcont 1351 -4036 1351 -4036 0 FreeSans 640 0 0 0 OR_4.Inverter_0.VDD
flabel psubdiffcont 1365 -4728 1365 -4728 0 FreeSans 640 0 0 0 OR_4.Inverter_0.VSS
flabel metal1 1189 -4367 1189 -4367 0 FreeSans 640 0 0 0 OR_4.Inverter_0.IN
flabel metal1 1556 -4394 1556 -4394 0 FreeSans 640 0 0 0 OR_4.Inverter_0.OUT
flabel metal1 3254 -4373 3254 -4373 0 FreeSans 640 0 0 0 INV_BUFF_6.IN
flabel metal1 4145 -4387 4145 -4387 0 FreeSans 640 0 0 0 INV_BUFF_6.OUT
flabel metal1 3683 -4020 3683 -4020 0 FreeSans 640 0 0 0 INV_BUFF_6.VDD
flabel metal1 3703 -4740 3703 -4740 0 FreeSans 640 0 0 0 INV_BUFF_6.VSS
flabel nsubdiffcont 3892 -4036 3892 -4036 0 FreeSans 640 0 0 0 INV_BUFF_6.Inverter_0.VDD
flabel psubdiffcont 3906 -4728 3906 -4728 0 FreeSans 640 0 0 0 INV_BUFF_6.Inverter_0.VSS
flabel metal1 3730 -4367 3730 -4367 0 FreeSans 640 0 0 0 INV_BUFF_6.Inverter_0.IN
flabel metal1 4097 -4394 4097 -4394 0 FreeSans 640 0 0 0 INV_BUFF_6.Inverter_0.OUT
flabel nsubdiffcont 3488 -4036 3488 -4036 0 FreeSans 640 0 0 0 INV_BUFF_6.Inverter_1.VDD
flabel psubdiffcont 3502 -4728 3502 -4728 0 FreeSans 640 0 0 0 INV_BUFF_6.Inverter_1.VSS
flabel metal1 3326 -4367 3326 -4367 0 FreeSans 640 0 0 0 INV_BUFF_6.Inverter_1.IN
flabel metal1 3693 -4394 3693 -4394 0 FreeSans 640 0 0 0 INV_BUFF_6.Inverter_1.OUT
<< end >>
