magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2128 -2598 2128 2598
<< nwell >>
rect -128 -598 128 598
<< nsubdiff >>
rect -45 493 45 515
rect -45 -493 -23 493
rect 23 -493 45 493
rect -45 -515 45 -493
<< nsubdiffcont >>
rect -23 -493 23 493
<< metal1 >>
rect -34 493 34 504
rect -34 -493 -23 493
rect 23 -493 34 493
rect -34 -504 34 -493
<< end >>
