* NGSPICE file created from res_48k_flat.ext - technology: gf180mcuC

.subckt res_48k_flat A B VDD
X0 a_364_2227# a_124_124# VDD.t2 ppolyf_u r_width=0.8u r_length=10u
X1 a_844_2227# a_604_124# VDD.t7 ppolyf_u r_width=0.8u r_length=10u
X2 a_1324_2227# a_1084_124# VDD.t1 ppolyf_u r_width=0.8u r_length=10u
X3 a_1804_2227# a_1564_124# VDD.t0 ppolyf_u r_width=0.8u r_length=10u
X4 a_1804_2227# a_2044_124# VDD.t3 ppolyf_u r_width=0.8u r_length=10u
X5 a_2284_2227# a_2524_124# VDD.t10 ppolyf_u r_width=0.8u r_length=10u
X6 a_844_2227# a_1084_124# VDD.t4 ppolyf_u r_width=0.8u r_length=10u
X7 a_1324_2227# a_1564_124# VDD.t11 ppolyf_u r_width=0.8u r_length=10u
X8 A.t0 a_124_124# VDD.t6 ppolyf_u r_width=0.8u r_length=10u
X9 a_364_2227# a_604_124# VDD.t8 ppolyf_u r_width=0.8u r_length=10u
X10 a_2284_2227# a_2044_124# VDD.t9 ppolyf_u r_width=0.8u r_length=10u
X11 B.t0 a_2524_124# VDD.t5 ppolyf_u r_width=0.8u r_length=10u
R0 VDD.t10 VDD.t5 85.7761
R1 VDD.t9 VDD.t10 85.7761
R2 VDD.t3 VDD.t9 85.7761
R3 VDD.t0 VDD.t3 85.7761
R4 VDD.t11 VDD.t1 85.7761
R5 VDD.t1 VDD.t4 85.7761
R6 VDD.t4 VDD.t7 85.7761
R7 VDD.t7 VDD.t8 85.7761
R8 VDD.t8 VDD.t2 85.7761
R9 VDD.t2 VDD.t6 85.7761
R10 VDD.n0 VDD.t0 76.8411
R11 VDD.n0 VDD.t11 8.93545
R12 VDD VDD.n2 3.15339
R13 VDD.n2 VDD.n0 3.1505
R14 VDD.n2 VDD.n1 0.448216
R15 A A.t0 7.19856
R16 B B.t0 7.19406
C0 a_2524_124# VDD 0.261f
C1 a_1564_124# a_2044_124# 0.0416f
C2 a_2284_2227# a_1804_2227# 0.0416f
C3 VDD B 0.182f
C4 a_364_2227# VDD 0.235f
C5 A a_844_2227# 0.00112f
C6 a_2524_124# a_2044_124# 0.0416f
C7 A a_1804_2227# 5.24e-20
C8 a_1324_2227# a_844_2227# 0.0416f
C9 a_124_124# a_604_124# 0.0416f
C10 a_1324_2227# a_1804_2227# 0.0416f
C11 a_1084_124# a_604_124# 0.0416f
C12 a_1564_124# a_1084_124# 0.0416f
C13 VDD a_2044_124# 0.253f
C14 A a_1324_2227# 4.21e-19
C15 VDD a_844_2227# 0.235f
C16 a_124_124# VDD 0.261f
C17 a_844_2227# B 5.34e-20
C18 VDD a_1804_2227# 0.235f
C19 VDD a_1084_124# 0.253f
C20 a_364_2227# a_844_2227# 0.0416f
C21 VDD a_2284_2227# 0.235f
C22 B a_1804_2227# 0.00114f
C23 a_2284_2227# B 0.049f
C24 A VDD 0.182f
C25 a_364_2227# A 0.0489f
C26 VDD a_604_124# 0.253f
C27 a_1324_2227# VDD 0.235f
C28 a_1564_124# VDD 0.321f
C29 a_1324_2227# B 4.29e-19
C30 B VSUBS 0.192f
C31 A VSUBS 0.193f
C32 VDD VSUBS 26.7f
C33 a_2524_124# VSUBS 0.227f
C34 a_2044_124# VSUBS 0.213f
C35 a_2284_2227# VSUBS 0.231f
C36 a_1564_124# VSUBS 0.18f
C37 a_1804_2227# VSUBS 0.231f
C38 a_1084_124# VSUBS 0.213f
C39 a_1324_2227# VSUBS 0.231f
C40 a_604_124# VSUBS 0.213f
C41 a_844_2227# VSUBS 0.231f
C42 a_124_124# VSUBS 0.227f
C43 a_364_2227# VSUBS 0.231f
.ends

