magic
tech gf180mcuC
magscale 1 10
timestamp 1714126980
<< pwell >>
rect -168 -168 168 168
<< nmos >>
rect -56 -100 56 100
<< ndiff >>
rect -144 87 -56 100
rect -144 -87 -131 87
rect -85 -87 -56 87
rect -144 -100 -56 -87
rect 56 87 144 100
rect 56 -87 85 87
rect 131 -87 144 87
rect 56 -100 144 -87
<< ndiffc >>
rect -131 -87 -85 87
rect 85 -87 131 87
<< polysilicon >>
rect -56 100 56 144
rect -56 -144 56 -100
<< metal1 >>
rect -131 87 -85 98
rect -131 -98 -85 -87
rect 85 87 131 98
rect 85 -98 131 -87
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 1 l 0.56 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
