magic
tech gf180mcuC
magscale 1 10
timestamp 1698947120
<< nwell >>
rect 3407 10933 5689 14411
rect -7770 4277 -3759 10715
rect 493 7241 5689 10933
rect 11863 7241 17059 11779
rect 32592 7342 40984 12256
rect 42288 7342 50680 12256
rect 51984 7342 60376 12256
rect 61680 7342 65936 12256
rect 872 1399 5074 4849
rect 18076 939 31918 5811
<< pwell >>
rect 6425 13632 6705 14344
rect 6713 13632 8113 14344
rect 8121 13632 8401 14344
rect 6425 12770 6705 13482
rect 6713 12770 8113 13482
rect 8121 12770 8401 13482
rect 6425 11908 6705 12620
rect 6713 11908 8113 12620
rect 8121 11908 8401 12620
rect 18675 12521 18955 13257
rect 18963 12521 20363 13257
rect 20371 12521 20651 13257
rect 23827 12521 24107 13257
rect 24115 12521 25515 13257
rect 25523 12521 25803 13257
rect 27796 12521 28076 13257
rect 28084 12521 29484 13257
rect 29492 12521 29772 13257
rect 6425 11046 6705 11758
rect 6713 11046 8113 11758
rect 8121 11046 8401 11758
rect 6425 10184 6705 10896
rect 6713 10184 8113 10896
rect 8121 10184 8401 10896
rect 8660 10165 8940 10877
rect 8948 10165 9228 10877
rect 9236 10165 9676 10877
rect 9684 10165 10124 10877
rect 10132 10165 10572 10877
rect 10580 10165 10860 10877
rect 10868 10165 11148 10877
rect 6425 9322 6705 10034
rect 6713 9322 8113 10034
rect 8121 9322 8401 10034
rect 8660 9303 8940 10015
rect 8948 9303 9228 10015
rect 9236 9303 9676 10015
rect 9684 9303 10124 10015
rect 10132 9303 10572 10015
rect 10580 9303 10860 10015
rect 10868 9303 11148 10015
rect 6425 8460 6705 9172
rect 6713 8460 8113 9172
rect 8121 8460 8401 9172
rect 8660 8441 8940 9153
rect 8948 8441 9228 9153
rect 9236 8441 9676 9153
rect 9684 8441 10124 9153
rect 10132 8441 10572 9153
rect 10580 8441 10860 9153
rect 10868 8441 11148 9153
rect 6425 7598 6705 8310
rect 6713 7598 8113 8310
rect 8121 7598 8401 8310
rect 8660 7579 8940 8291
rect 8948 7579 9228 8291
rect 9236 7579 9676 8291
rect 9684 7579 10124 8291
rect 10132 7579 10572 8291
rect 10580 7579 10860 8291
rect 10868 7579 11148 8291
rect 18675 11585 18955 12321
rect 18963 11585 20363 12321
rect 20371 11585 20651 12321
rect 23827 11585 24107 12321
rect 24115 11585 25515 12321
rect 25523 11585 25803 12321
rect 27796 11585 28076 12321
rect 28084 11585 29484 12321
rect 29492 11585 29772 12321
rect 18675 10649 18955 11385
rect 18963 10649 20363 11385
rect 20371 10649 20651 11385
rect 23827 10649 24107 11385
rect 24115 10649 25515 11385
rect 25523 10649 25803 11385
rect 27796 10649 28076 11385
rect 28084 10649 29484 11385
rect 29492 10649 29772 11385
rect 18675 9713 18955 10449
rect 18963 9713 20363 10449
rect 20371 9713 20651 10449
rect 23827 9713 24107 10449
rect 24115 9713 25515 10449
rect 25523 9713 25803 10449
rect 27796 9713 28076 10449
rect 28084 9713 29484 10449
rect 29492 9713 29772 10449
rect 18675 8777 18955 9513
rect 18963 8777 20363 9513
rect 20371 8777 20651 9513
rect 23827 8777 24107 9513
rect 24115 8777 25515 9513
rect 25523 8777 25803 9513
rect 27796 8777 28076 9513
rect 28084 8777 29484 9513
rect 29492 8777 29772 9513
rect 18675 7841 18955 8577
rect 18963 7841 20363 8577
rect 20371 7841 20651 8577
rect 23827 7841 24107 8577
rect 24115 7841 25515 8577
rect 25523 7841 25803 8577
rect 27796 7841 28076 8577
rect 28084 7841 29484 8577
rect 29492 7841 29772 8577
rect 7359 5470 7639 5806
rect 7647 5470 9367 5806
rect 9375 5470 9655 5806
rect 7359 4934 7639 5270
rect 7647 4934 9367 5270
rect 9375 4934 9655 5270
rect 7359 4398 7639 4734
rect 7647 4398 9367 4734
rect 9375 4398 9655 4734
rect 7359 3862 7639 4198
rect 7647 3862 9367 4198
rect 9375 3862 9655 4198
rect 7359 3326 7639 3662
rect 7647 3326 9367 3662
rect 9375 3326 9655 3662
rect 7359 2790 7639 3126
rect 7647 2790 9367 3126
rect 9375 2790 9655 3126
rect 12646 2777 13070 3849
rect 13078 2777 15022 3849
rect 15030 2777 16974 3849
rect 6112 2161 6392 2497
rect 6400 2161 9400 2497
rect 9408 2161 10904 2497
rect 12646 1941 13070 2477
rect 13078 1941 15022 2477
rect 15030 1941 16974 2477
rect 6112 1524 6392 1860
rect 6400 1524 9800 1860
rect 9824 1524 10904 1860
<< nmos >>
rect 6537 13700 6593 14276
rect 6825 13700 6881 14276
rect 6985 13700 7041 14276
rect 7145 13700 7201 14276
rect 7305 13700 7361 14276
rect 7465 13700 7521 14276
rect 7625 13700 7681 14276
rect 7785 13700 7841 14276
rect 7945 13700 8001 14276
rect 8233 13700 8289 14276
rect 6537 12838 6593 13414
rect 6825 12838 6881 13414
rect 6985 12838 7041 13414
rect 7145 12838 7201 13414
rect 7305 12838 7361 13414
rect 7465 12838 7521 13414
rect 7625 12838 7681 13414
rect 7785 12838 7841 13414
rect 7945 12838 8001 13414
rect 8233 12838 8289 13414
rect 6537 11976 6593 12552
rect 6825 11976 6881 12552
rect 6985 11976 7041 12552
rect 7145 11976 7201 12552
rect 7305 11976 7361 12552
rect 7465 11976 7521 12552
rect 7625 11976 7681 12552
rect 7785 11976 7841 12552
rect 7945 11976 8001 12552
rect 8233 11976 8289 12552
rect 18787 12589 18843 13189
rect 19075 12589 19131 13189
rect 19235 12589 19291 13189
rect 19395 12589 19451 13189
rect 19555 12589 19611 13189
rect 19715 12589 19771 13189
rect 19875 12589 19931 13189
rect 20035 12589 20091 13189
rect 20195 12589 20251 13189
rect 20483 12589 20539 13189
rect 6537 11114 6593 11690
rect 6825 11114 6881 11690
rect 6985 11114 7041 11690
rect 7145 11114 7201 11690
rect 7305 11114 7361 11690
rect 7465 11114 7521 11690
rect 7625 11114 7681 11690
rect 7785 11114 7841 11690
rect 7945 11114 8001 11690
rect 8233 11114 8289 11690
rect 6537 10252 6593 10828
rect 6825 10252 6881 10828
rect 6985 10252 7041 10828
rect 7145 10252 7201 10828
rect 7305 10252 7361 10828
rect 7465 10252 7521 10828
rect 7625 10252 7681 10828
rect 7785 10252 7841 10828
rect 7945 10252 8001 10828
rect 8233 10252 8289 10828
rect 8772 10233 8828 10809
rect 9060 10233 9116 10809
rect 9348 10233 9404 10809
rect 9508 10233 9564 10809
rect 9796 10233 9852 10809
rect 9956 10233 10012 10809
rect 10244 10233 10300 10809
rect 10404 10233 10460 10809
rect 10692 10233 10748 10809
rect 10980 10233 11036 10809
rect 6537 9390 6593 9966
rect 6825 9390 6881 9966
rect 6985 9390 7041 9966
rect 7145 9390 7201 9966
rect 7305 9390 7361 9966
rect 7465 9390 7521 9966
rect 7625 9390 7681 9966
rect 7785 9390 7841 9966
rect 7945 9390 8001 9966
rect 8233 9390 8289 9966
rect 8772 9371 8828 9947
rect 9060 9371 9116 9947
rect 9348 9371 9404 9947
rect 9508 9371 9564 9947
rect 9796 9371 9852 9947
rect 9956 9371 10012 9947
rect 10244 9371 10300 9947
rect 10404 9371 10460 9947
rect 10692 9371 10748 9947
rect 10980 9371 11036 9947
rect 6537 8528 6593 9104
rect 6825 8528 6881 9104
rect 6985 8528 7041 9104
rect 7145 8528 7201 9104
rect 7305 8528 7361 9104
rect 7465 8528 7521 9104
rect 7625 8528 7681 9104
rect 7785 8528 7841 9104
rect 7945 8528 8001 9104
rect 8233 8528 8289 9104
rect 8772 8509 8828 9085
rect 9060 8509 9116 9085
rect 9348 8509 9404 9085
rect 9508 8509 9564 9085
rect 9796 8509 9852 9085
rect 9956 8509 10012 9085
rect 10244 8509 10300 9085
rect 10404 8509 10460 9085
rect 10692 8509 10748 9085
rect 10980 8509 11036 9085
rect 6537 7666 6593 8242
rect 6825 7666 6881 8242
rect 6985 7666 7041 8242
rect 7145 7666 7201 8242
rect 7305 7666 7361 8242
rect 7465 7666 7521 8242
rect 7625 7666 7681 8242
rect 7785 7666 7841 8242
rect 7945 7666 8001 8242
rect 8233 7666 8289 8242
rect 8772 7647 8828 8223
rect 9060 7647 9116 8223
rect 9348 7647 9404 8223
rect 9508 7647 9564 8223
rect 9796 7647 9852 8223
rect 9956 7647 10012 8223
rect 10244 7647 10300 8223
rect 10404 7647 10460 8223
rect 10692 7647 10748 8223
rect 10980 7647 11036 8223
rect 18787 11653 18843 12253
rect 19075 11653 19131 12253
rect 19235 11653 19291 12253
rect 19395 11653 19451 12253
rect 19555 11653 19611 12253
rect 19715 11653 19771 12253
rect 19875 11653 19931 12253
rect 20035 11653 20091 12253
rect 20195 11653 20251 12253
rect 20483 11653 20539 12253
rect 18787 10717 18843 11317
rect 19075 10717 19131 11317
rect 19235 10717 19291 11317
rect 19395 10717 19451 11317
rect 19555 10717 19611 11317
rect 19715 10717 19771 11317
rect 19875 10717 19931 11317
rect 20035 10717 20091 11317
rect 20195 10717 20251 11317
rect 20483 10717 20539 11317
rect 18787 9781 18843 10381
rect 19075 9781 19131 10381
rect 19235 9781 19291 10381
rect 19395 9781 19451 10381
rect 19555 9781 19611 10381
rect 19715 9781 19771 10381
rect 19875 9781 19931 10381
rect 20035 9781 20091 10381
rect 20195 9781 20251 10381
rect 20483 9781 20539 10381
rect 18787 8845 18843 9445
rect 19075 8845 19131 9445
rect 19235 8845 19291 9445
rect 19395 8845 19451 9445
rect 19555 8845 19611 9445
rect 19715 8845 19771 9445
rect 19875 8845 19931 9445
rect 20035 8845 20091 9445
rect 20195 8845 20251 9445
rect 20483 8845 20539 9445
rect 18787 7909 18843 8509
rect 19075 7909 19131 8509
rect 19235 7909 19291 8509
rect 19395 7909 19451 8509
rect 19555 7909 19611 8509
rect 19715 7909 19771 8509
rect 19875 7909 19931 8509
rect 20035 7909 20091 8509
rect 20195 7909 20251 8509
rect 20483 7909 20539 8509
rect 23939 12589 23995 13189
rect 24227 12589 24283 13189
rect 24387 12589 24443 13189
rect 24547 12589 24603 13189
rect 24707 12589 24763 13189
rect 24867 12589 24923 13189
rect 25027 12589 25083 13189
rect 25187 12589 25243 13189
rect 25347 12589 25403 13189
rect 25635 12589 25691 13189
rect 23939 11653 23995 12253
rect 24227 11653 24283 12253
rect 24387 11653 24443 12253
rect 24547 11653 24603 12253
rect 24707 11653 24763 12253
rect 24867 11653 24923 12253
rect 25027 11653 25083 12253
rect 25187 11653 25243 12253
rect 25347 11653 25403 12253
rect 25635 11653 25691 12253
rect 23939 10717 23995 11317
rect 24227 10717 24283 11317
rect 24387 10717 24443 11317
rect 24547 10717 24603 11317
rect 24707 10717 24763 11317
rect 24867 10717 24923 11317
rect 25027 10717 25083 11317
rect 25187 10717 25243 11317
rect 25347 10717 25403 11317
rect 25635 10717 25691 11317
rect 23939 9781 23995 10381
rect 24227 9781 24283 10381
rect 24387 9781 24443 10381
rect 24547 9781 24603 10381
rect 24707 9781 24763 10381
rect 24867 9781 24923 10381
rect 25027 9781 25083 10381
rect 25187 9781 25243 10381
rect 25347 9781 25403 10381
rect 25635 9781 25691 10381
rect 23939 8845 23995 9445
rect 24227 8845 24283 9445
rect 24387 8845 24443 9445
rect 24547 8845 24603 9445
rect 24707 8845 24763 9445
rect 24867 8845 24923 9445
rect 25027 8845 25083 9445
rect 25187 8845 25243 9445
rect 25347 8845 25403 9445
rect 25635 8845 25691 9445
rect 23939 7909 23995 8509
rect 24227 7909 24283 8509
rect 24387 7909 24443 8509
rect 24547 7909 24603 8509
rect 24707 7909 24763 8509
rect 24867 7909 24923 8509
rect 25027 7909 25083 8509
rect 25187 7909 25243 8509
rect 25347 7909 25403 8509
rect 25635 7909 25691 8509
rect 27908 12589 27964 13189
rect 28196 12589 28252 13189
rect 28356 12589 28412 13189
rect 28516 12589 28572 13189
rect 28676 12589 28732 13189
rect 28836 12589 28892 13189
rect 28996 12589 29052 13189
rect 29156 12589 29212 13189
rect 29316 12589 29372 13189
rect 29604 12589 29660 13189
rect 27908 11653 27964 12253
rect 28196 11653 28252 12253
rect 28356 11653 28412 12253
rect 28516 11653 28572 12253
rect 28676 11653 28732 12253
rect 28836 11653 28892 12253
rect 28996 11653 29052 12253
rect 29156 11653 29212 12253
rect 29316 11653 29372 12253
rect 29604 11653 29660 12253
rect 27908 10717 27964 11317
rect 28196 10717 28252 11317
rect 28356 10717 28412 11317
rect 28516 10717 28572 11317
rect 28676 10717 28732 11317
rect 28836 10717 28892 11317
rect 28996 10717 29052 11317
rect 29156 10717 29212 11317
rect 29316 10717 29372 11317
rect 29604 10717 29660 11317
rect 27908 9781 27964 10381
rect 28196 9781 28252 10381
rect 28356 9781 28412 10381
rect 28516 9781 28572 10381
rect 28676 9781 28732 10381
rect 28836 9781 28892 10381
rect 28996 9781 29052 10381
rect 29156 9781 29212 10381
rect 29316 9781 29372 10381
rect 29604 9781 29660 10381
rect 27908 8845 27964 9445
rect 28196 8845 28252 9445
rect 28356 8845 28412 9445
rect 28516 8845 28572 9445
rect 28676 8845 28732 9445
rect 28836 8845 28892 9445
rect 28996 8845 29052 9445
rect 29156 8845 29212 9445
rect 29316 8845 29372 9445
rect 29604 8845 29660 9445
rect 27908 7909 27964 8509
rect 28196 7909 28252 8509
rect 28356 7909 28412 8509
rect 28516 7909 28572 8509
rect 28676 7909 28732 8509
rect 28836 7909 28892 8509
rect 28996 7909 29052 8509
rect 29156 7909 29212 8509
rect 29316 7909 29372 8509
rect 29604 7909 29660 8509
rect 7471 5538 7527 5738
rect 7759 5538 7815 5738
rect 7919 5538 7975 5738
rect 8079 5538 8135 5738
rect 8239 5538 8295 5738
rect 8399 5538 8455 5738
rect 8559 5538 8615 5738
rect 8719 5538 8775 5738
rect 8879 5538 8935 5738
rect 9039 5538 9095 5738
rect 9199 5538 9255 5738
rect 9487 5538 9543 5738
rect 7471 5002 7527 5202
rect 7759 5002 7815 5202
rect 7919 5002 7975 5202
rect 8079 5002 8135 5202
rect 8239 5002 8295 5202
rect 8399 5002 8455 5202
rect 8559 5002 8615 5202
rect 8719 5002 8775 5202
rect 8879 5002 8935 5202
rect 9039 5002 9095 5202
rect 9199 5002 9255 5202
rect 9487 5002 9543 5202
rect 7471 4466 7527 4666
rect 7759 4466 7815 4666
rect 7919 4466 7975 4666
rect 8079 4466 8135 4666
rect 8239 4466 8295 4666
rect 8399 4466 8455 4666
rect 8559 4466 8615 4666
rect 8719 4466 8775 4666
rect 8879 4466 8935 4666
rect 9039 4466 9095 4666
rect 9199 4466 9255 4666
rect 9487 4466 9543 4666
rect 7471 3930 7527 4130
rect 7759 3930 7815 4130
rect 7919 3930 7975 4130
rect 8079 3930 8135 4130
rect 8239 3930 8295 4130
rect 8399 3930 8455 4130
rect 8559 3930 8615 4130
rect 8719 3930 8775 4130
rect 8879 3930 8935 4130
rect 9039 3930 9095 4130
rect 9199 3930 9255 4130
rect 9487 3930 9543 4130
rect 7471 3394 7527 3594
rect 7759 3394 7815 3594
rect 7919 3394 7975 3594
rect 8079 3394 8135 3594
rect 8239 3394 8295 3594
rect 8399 3394 8455 3594
rect 8559 3394 8615 3594
rect 8719 3394 8775 3594
rect 8879 3394 8935 3594
rect 9039 3394 9095 3594
rect 9199 3394 9255 3594
rect 9487 3394 9543 3594
rect 7471 2858 7527 3058
rect 7759 2858 7815 3058
rect 7919 2858 7975 3058
rect 8079 2858 8135 3058
rect 8239 2858 8295 3058
rect 8399 2858 8455 3058
rect 8559 2858 8615 3058
rect 8719 2858 8775 3058
rect 8879 2858 8935 3058
rect 9039 2858 9095 3058
rect 9199 2858 9255 3058
rect 9487 2858 9543 3058
rect 12758 3381 12958 3781
rect 13190 3381 13390 3781
rect 13494 3381 13694 3781
rect 13798 3381 13998 3781
rect 14102 3381 14302 3781
rect 14406 3381 14606 3781
rect 14710 3381 14910 3781
rect 15142 3381 15342 3781
rect 15446 3381 15646 3781
rect 15750 3381 15950 3781
rect 16054 3381 16254 3781
rect 16358 3381 16558 3781
rect 16662 3381 16862 3781
rect 6224 2229 6280 2429
rect 6512 2229 6568 2429
rect 6672 2229 6728 2429
rect 6832 2229 6888 2429
rect 6992 2229 7048 2429
rect 7152 2229 7208 2429
rect 7312 2229 7368 2429
rect 7472 2229 7528 2429
rect 7632 2229 7688 2429
rect 7792 2229 7848 2429
rect 7952 2229 8008 2429
rect 8112 2229 8168 2429
rect 8272 2229 8328 2429
rect 8432 2229 8488 2429
rect 8592 2229 8648 2429
rect 8752 2229 8808 2429
rect 8912 2229 8968 2429
rect 9072 2229 9128 2429
rect 9232 2229 9288 2429
rect 9520 2229 9720 2429
rect 9824 2229 10024 2429
rect 10128 2229 10328 2429
rect 10432 2229 10632 2429
rect 10736 2229 10792 2429
rect 6224 1592 6280 1792
rect 6512 1592 6624 1792
rect 6728 1592 6840 1792
rect 6944 1592 7056 1792
rect 7160 1592 7272 1792
rect 7376 1592 7488 1792
rect 7592 1592 7704 1792
rect 7808 1592 7920 1792
rect 8024 1592 8136 1792
rect 8240 1592 8352 1792
rect 8456 1592 8568 1792
rect 8672 1592 8728 1792
rect 8832 1592 8888 1792
rect 8992 1592 9048 1792
rect 9152 1592 9208 1792
rect 9312 1592 9368 1792
rect 9472 1592 9528 1792
rect 9632 1592 9688 1792
rect 9936 1592 9992 1792
rect 10096 1592 10152 1792
rect 10256 1592 10312 1792
rect 10416 1592 10472 1792
rect 10576 1592 10632 1792
rect 10736 1592 10792 1792
rect 12758 2845 12958 3245
rect 13190 2845 13390 3245
rect 13494 2845 13694 3245
rect 13798 2845 13998 3245
rect 14102 2845 14302 3245
rect 14406 2845 14606 3245
rect 14710 2845 14910 3245
rect 15142 2845 15342 3245
rect 15446 2845 15646 3245
rect 15750 2845 15950 3245
rect 16054 2845 16254 3245
rect 16358 2845 16558 3245
rect 16662 2845 16862 3245
rect 12758 2009 12958 2409
rect 13190 2009 13390 2409
rect 13494 2009 13694 2409
rect 13798 2009 13998 2409
rect 14102 2009 14302 2409
rect 14406 2009 14606 2409
rect 14710 2009 14910 2409
rect 15142 2009 15342 2409
rect 15446 2009 15646 2409
rect 15750 2009 15950 2409
rect 16054 2009 16254 2409
rect 16358 2009 16558 2409
rect 16662 2009 16862 2409
<< pmos >>
rect 3672 13276 3728 14026
rect 3960 13276 4016 14026
rect 4120 13276 4176 14026
rect 4280 13276 4336 14026
rect 4440 13276 4496 14026
rect 4600 13276 4656 14026
rect 4760 13276 4816 14026
rect 4920 13276 4976 14026
rect 5080 13276 5136 14026
rect 5368 13276 5424 14026
rect 3672 12146 3728 12896
rect 3960 12146 4016 12896
rect 4120 12146 4176 12896
rect 4280 12146 4336 12896
rect 4440 12146 4496 12896
rect 4600 12146 4656 12896
rect 4760 12146 4816 12896
rect 4920 12146 4976 12896
rect 5080 12146 5136 12896
rect 5368 12146 5424 12896
rect 3672 11016 3728 11766
rect 3960 11016 4016 11766
rect 4120 11016 4176 11766
rect 4280 11016 4336 11766
rect 4440 11016 4496 11766
rect 4600 11016 4656 11766
rect 4760 11016 4816 11766
rect 4920 11016 4976 11766
rect 5080 11016 5136 11766
rect 5368 11016 5424 11766
rect 986 9932 1098 10558
rect 1202 9932 1314 10558
rect 1418 9932 1530 10558
rect 1634 9932 1746 10558
rect 1850 9932 1962 10558
rect 2066 9932 2178 10558
rect 2282 9932 2394 10558
rect 2498 9932 2610 10558
rect 2714 9932 2826 10558
rect 2930 9932 3042 10558
rect 3672 9886 3728 10636
rect 3960 9886 4016 10636
rect 4120 9886 4176 10636
rect 4280 9886 4336 10636
rect 4440 9886 4496 10636
rect 4600 9886 4656 10636
rect 4760 9886 4816 10636
rect 4920 9886 4976 10636
rect 5080 9886 5136 10636
rect 5368 9886 5424 10636
rect 986 9170 1098 9796
rect 1202 9170 1314 9796
rect 1418 9170 1530 9796
rect 1634 9170 1746 9796
rect 1850 9170 1962 9796
rect 2066 9170 2178 9796
rect 2282 9170 2394 9796
rect 2498 9170 2610 9796
rect 2714 9170 2826 9796
rect 2930 9170 3042 9796
rect 986 8408 1098 9034
rect 1202 8408 1314 9034
rect 1418 8408 1530 9034
rect 1634 8408 1746 9034
rect 1850 8408 1962 9034
rect 2066 8408 2178 9034
rect 2282 8408 2394 9034
rect 2498 8408 2610 9034
rect 2714 8408 2826 9034
rect 2930 8408 3042 9034
rect 3672 8756 3728 9506
rect 3960 8756 4016 9506
rect 4120 8756 4176 9506
rect 4280 8756 4336 9506
rect 4440 8756 4496 9506
rect 4600 8756 4656 9506
rect 4760 8756 4816 9506
rect 4920 8756 4976 9506
rect 5080 8756 5136 9506
rect 5368 8756 5424 9506
rect 986 7646 1098 8272
rect 1202 7646 1314 8272
rect 1418 7646 1530 8272
rect 1634 7646 1746 8272
rect 1850 7646 1962 8272
rect 2066 7646 2178 8272
rect 2282 7646 2394 8272
rect 2498 7646 2610 8272
rect 2714 7646 2826 8272
rect 2930 7646 3042 8272
rect 3672 7626 3728 8376
rect 3960 7626 4016 8376
rect 4120 7626 4176 8376
rect 4280 7626 4336 8376
rect 4440 7626 4496 8376
rect 4600 7626 4656 8376
rect 4760 7626 4816 8376
rect 4920 7626 4976 8376
rect 5080 7626 5136 8376
rect 5368 7626 5424 8376
rect 12154 10751 12210 11377
rect 12442 10751 12498 11377
rect 12730 10751 12786 11377
rect 12890 10751 12946 11377
rect 13178 10751 13234 11377
rect 13338 10751 13394 11377
rect 13626 10751 13682 11377
rect 13786 10751 13842 11377
rect 14074 10751 14130 11377
rect 14362 10751 14418 11377
rect 14948 10751 15004 11377
rect 15236 10751 15292 11377
rect 15396 10751 15452 11377
rect 15556 10751 15612 11377
rect 15716 10751 15772 11377
rect 15876 10751 15932 11377
rect 16036 10751 16092 11377
rect 16196 10751 16252 11377
rect 16356 10751 16412 11377
rect 16644 10751 16700 11377
rect 12154 9715 12210 10341
rect 12442 9715 12498 10341
rect 12730 9715 12786 10341
rect 12890 9715 12946 10341
rect 13178 9715 13234 10341
rect 13338 9715 13394 10341
rect 13626 9715 13682 10341
rect 13786 9715 13842 10341
rect 14074 9715 14130 10341
rect 14362 9715 14418 10341
rect 14948 9715 15004 10341
rect 15236 9715 15292 10341
rect 15396 9715 15452 10341
rect 15556 9715 15612 10341
rect 15716 9715 15772 10341
rect 15876 9715 15932 10341
rect 16036 9715 16092 10341
rect 16196 9715 16252 10341
rect 16356 9715 16412 10341
rect 16644 9715 16700 10341
rect 12154 8679 12210 9305
rect 12442 8679 12498 9305
rect 12730 8679 12786 9305
rect 12890 8679 12946 9305
rect 13178 8679 13234 9305
rect 13338 8679 13394 9305
rect 13626 8679 13682 9305
rect 13786 8679 13842 9305
rect 14074 8679 14130 9305
rect 14362 8679 14418 9305
rect 14948 8679 15004 9305
rect 15236 8679 15292 9305
rect 15396 8679 15452 9305
rect 15556 8679 15612 9305
rect 15716 8679 15772 9305
rect 15876 8679 15932 9305
rect 16036 8679 16092 9305
rect 16196 8679 16252 9305
rect 16356 8679 16412 9305
rect 16644 8679 16700 9305
rect 12154 7643 12210 8269
rect 12442 7643 12498 8269
rect 12730 7643 12786 8269
rect 12890 7643 12946 8269
rect 13178 7643 13234 8269
rect 13338 7643 13394 8269
rect 13626 7643 13682 8269
rect 13786 7643 13842 8269
rect 14074 7643 14130 8269
rect 14362 7643 14418 8269
rect 14948 7643 15004 8269
rect 15236 7643 15292 8269
rect 15396 7643 15452 8269
rect 15556 7643 15612 8269
rect 15716 7643 15772 8269
rect 15876 7643 15932 8269
rect 16036 7643 16092 8269
rect 16196 7643 16252 8269
rect 16356 7643 16412 8269
rect 16644 7643 16700 8269
rect 33204 11089 33260 11689
rect 33492 11089 33548 11689
rect 33652 11089 33708 11689
rect 33812 11089 33868 11689
rect 33972 11089 34028 11689
rect 34132 11089 34188 11689
rect 34292 11089 34348 11689
rect 34452 11089 34508 11689
rect 34612 11089 34668 11689
rect 34772 11089 34828 11689
rect 34932 11089 34988 11689
rect 35092 11089 35148 11689
rect 35252 11089 35308 11689
rect 35412 11089 35468 11689
rect 35572 11089 35628 11689
rect 35732 11089 35788 11689
rect 35892 11089 35948 11689
rect 36180 11089 36236 11689
rect 37340 11089 37396 11689
rect 37628 11089 37684 11689
rect 37788 11089 37844 11689
rect 37948 11089 38004 11689
rect 38108 11089 38164 11689
rect 38268 11089 38324 11689
rect 38428 11089 38484 11689
rect 38588 11089 38644 11689
rect 38748 11089 38804 11689
rect 38908 11089 38964 11689
rect 39068 11089 39124 11689
rect 39228 11089 39284 11689
rect 39388 11089 39444 11689
rect 39548 11089 39604 11689
rect 39708 11089 39764 11689
rect 39868 11089 39924 11689
rect 40028 11089 40084 11689
rect 40316 11089 40372 11689
rect 33204 10029 33260 10629
rect 33492 10029 33548 10629
rect 33652 10029 33708 10629
rect 33812 10029 33868 10629
rect 33972 10029 34028 10629
rect 34132 10029 34188 10629
rect 34292 10029 34348 10629
rect 34452 10029 34508 10629
rect 34612 10029 34668 10629
rect 34772 10029 34828 10629
rect 34932 10029 34988 10629
rect 35092 10029 35148 10629
rect 35252 10029 35308 10629
rect 35412 10029 35468 10629
rect 35572 10029 35628 10629
rect 35732 10029 35788 10629
rect 35892 10029 35948 10629
rect 36180 10029 36236 10629
rect 37340 10029 37396 10629
rect 37628 10029 37684 10629
rect 37788 10029 37844 10629
rect 37948 10029 38004 10629
rect 38108 10029 38164 10629
rect 38268 10029 38324 10629
rect 38428 10029 38484 10629
rect 38588 10029 38644 10629
rect 38748 10029 38804 10629
rect 38908 10029 38964 10629
rect 39068 10029 39124 10629
rect 39228 10029 39284 10629
rect 39388 10029 39444 10629
rect 39548 10029 39604 10629
rect 39708 10029 39764 10629
rect 39868 10029 39924 10629
rect 40028 10029 40084 10629
rect 40316 10029 40372 10629
rect 33204 8969 33260 9569
rect 33492 8969 33548 9569
rect 33652 8969 33708 9569
rect 33812 8969 33868 9569
rect 33972 8969 34028 9569
rect 34132 8969 34188 9569
rect 34292 8969 34348 9569
rect 34452 8969 34508 9569
rect 34612 8969 34668 9569
rect 34772 8969 34828 9569
rect 34932 8969 34988 9569
rect 35092 8969 35148 9569
rect 35252 8969 35308 9569
rect 35412 8969 35468 9569
rect 35572 8969 35628 9569
rect 35732 8969 35788 9569
rect 35892 8969 35948 9569
rect 36180 8969 36236 9569
rect 37340 8969 37396 9569
rect 37628 8969 37684 9569
rect 37788 8969 37844 9569
rect 37948 8969 38004 9569
rect 38108 8969 38164 9569
rect 38268 8969 38324 9569
rect 38428 8969 38484 9569
rect 38588 8969 38644 9569
rect 38748 8969 38804 9569
rect 38908 8969 38964 9569
rect 39068 8969 39124 9569
rect 39228 8969 39284 9569
rect 39388 8969 39444 9569
rect 39548 8969 39604 9569
rect 39708 8969 39764 9569
rect 39868 8969 39924 9569
rect 40028 8969 40084 9569
rect 40316 8969 40372 9569
rect 33204 7909 33260 8509
rect 33492 7909 33548 8509
rect 33652 7909 33708 8509
rect 33812 7909 33868 8509
rect 33972 7909 34028 8509
rect 34132 7909 34188 8509
rect 34292 7909 34348 8509
rect 34452 7909 34508 8509
rect 34612 7909 34668 8509
rect 34772 7909 34828 8509
rect 34932 7909 34988 8509
rect 35092 7909 35148 8509
rect 35252 7909 35308 8509
rect 35412 7909 35468 8509
rect 35572 7909 35628 8509
rect 35732 7909 35788 8509
rect 35892 7909 35948 8509
rect 36180 7909 36236 8509
rect 37340 7909 37396 8509
rect 37628 7909 37684 8509
rect 37788 7909 37844 8509
rect 37948 7909 38004 8509
rect 38108 7909 38164 8509
rect 38268 7909 38324 8509
rect 38428 7909 38484 8509
rect 38588 7909 38644 8509
rect 38748 7909 38804 8509
rect 38908 7909 38964 8509
rect 39068 7909 39124 8509
rect 39228 7909 39284 8509
rect 39388 7909 39444 8509
rect 39548 7909 39604 8509
rect 39708 7909 39764 8509
rect 39868 7909 39924 8509
rect 40028 7909 40084 8509
rect 40316 7909 40372 8509
rect 42900 11089 42956 11689
rect 43188 11089 43244 11689
rect 43348 11089 43404 11689
rect 43508 11089 43564 11689
rect 43668 11089 43724 11689
rect 43828 11089 43884 11689
rect 43988 11089 44044 11689
rect 44148 11089 44204 11689
rect 44308 11089 44364 11689
rect 44468 11089 44524 11689
rect 44628 11089 44684 11689
rect 44788 11089 44844 11689
rect 44948 11089 45004 11689
rect 45108 11089 45164 11689
rect 45268 11089 45324 11689
rect 45428 11089 45484 11689
rect 45588 11089 45644 11689
rect 45876 11089 45932 11689
rect 47036 11089 47092 11689
rect 47324 11089 47380 11689
rect 47484 11089 47540 11689
rect 47644 11089 47700 11689
rect 47804 11089 47860 11689
rect 47964 11089 48020 11689
rect 48124 11089 48180 11689
rect 48284 11089 48340 11689
rect 48444 11089 48500 11689
rect 48604 11089 48660 11689
rect 48764 11089 48820 11689
rect 48924 11089 48980 11689
rect 49084 11089 49140 11689
rect 49244 11089 49300 11689
rect 49404 11089 49460 11689
rect 49564 11089 49620 11689
rect 49724 11089 49780 11689
rect 50012 11089 50068 11689
rect 42900 10029 42956 10629
rect 43188 10029 43244 10629
rect 43348 10029 43404 10629
rect 43508 10029 43564 10629
rect 43668 10029 43724 10629
rect 43828 10029 43884 10629
rect 43988 10029 44044 10629
rect 44148 10029 44204 10629
rect 44308 10029 44364 10629
rect 44468 10029 44524 10629
rect 44628 10029 44684 10629
rect 44788 10029 44844 10629
rect 44948 10029 45004 10629
rect 45108 10029 45164 10629
rect 45268 10029 45324 10629
rect 45428 10029 45484 10629
rect 45588 10029 45644 10629
rect 45876 10029 45932 10629
rect 47036 10029 47092 10629
rect 47324 10029 47380 10629
rect 47484 10029 47540 10629
rect 47644 10029 47700 10629
rect 47804 10029 47860 10629
rect 47964 10029 48020 10629
rect 48124 10029 48180 10629
rect 48284 10029 48340 10629
rect 48444 10029 48500 10629
rect 48604 10029 48660 10629
rect 48764 10029 48820 10629
rect 48924 10029 48980 10629
rect 49084 10029 49140 10629
rect 49244 10029 49300 10629
rect 49404 10029 49460 10629
rect 49564 10029 49620 10629
rect 49724 10029 49780 10629
rect 50012 10029 50068 10629
rect 42900 8969 42956 9569
rect 43188 8969 43244 9569
rect 43348 8969 43404 9569
rect 43508 8969 43564 9569
rect 43668 8969 43724 9569
rect 43828 8969 43884 9569
rect 43988 8969 44044 9569
rect 44148 8969 44204 9569
rect 44308 8969 44364 9569
rect 44468 8969 44524 9569
rect 44628 8969 44684 9569
rect 44788 8969 44844 9569
rect 44948 8969 45004 9569
rect 45108 8969 45164 9569
rect 45268 8969 45324 9569
rect 45428 8969 45484 9569
rect 45588 8969 45644 9569
rect 45876 8969 45932 9569
rect 47036 8969 47092 9569
rect 47324 8969 47380 9569
rect 47484 8969 47540 9569
rect 47644 8969 47700 9569
rect 47804 8969 47860 9569
rect 47964 8969 48020 9569
rect 48124 8969 48180 9569
rect 48284 8969 48340 9569
rect 48444 8969 48500 9569
rect 48604 8969 48660 9569
rect 48764 8969 48820 9569
rect 48924 8969 48980 9569
rect 49084 8969 49140 9569
rect 49244 8969 49300 9569
rect 49404 8969 49460 9569
rect 49564 8969 49620 9569
rect 49724 8969 49780 9569
rect 50012 8969 50068 9569
rect 42900 7909 42956 8509
rect 43188 7909 43244 8509
rect 43348 7909 43404 8509
rect 43508 7909 43564 8509
rect 43668 7909 43724 8509
rect 43828 7909 43884 8509
rect 43988 7909 44044 8509
rect 44148 7909 44204 8509
rect 44308 7909 44364 8509
rect 44468 7909 44524 8509
rect 44628 7909 44684 8509
rect 44788 7909 44844 8509
rect 44948 7909 45004 8509
rect 45108 7909 45164 8509
rect 45268 7909 45324 8509
rect 45428 7909 45484 8509
rect 45588 7909 45644 8509
rect 45876 7909 45932 8509
rect 47036 7909 47092 8509
rect 47324 7909 47380 8509
rect 47484 7909 47540 8509
rect 47644 7909 47700 8509
rect 47804 7909 47860 8509
rect 47964 7909 48020 8509
rect 48124 7909 48180 8509
rect 48284 7909 48340 8509
rect 48444 7909 48500 8509
rect 48604 7909 48660 8509
rect 48764 7909 48820 8509
rect 48924 7909 48980 8509
rect 49084 7909 49140 8509
rect 49244 7909 49300 8509
rect 49404 7909 49460 8509
rect 49564 7909 49620 8509
rect 49724 7909 49780 8509
rect 50012 7909 50068 8509
rect 52596 11089 52652 11689
rect 52884 11089 52940 11689
rect 53044 11089 53100 11689
rect 53204 11089 53260 11689
rect 53364 11089 53420 11689
rect 53524 11089 53580 11689
rect 53684 11089 53740 11689
rect 53844 11089 53900 11689
rect 54004 11089 54060 11689
rect 54164 11089 54220 11689
rect 54324 11089 54380 11689
rect 54484 11089 54540 11689
rect 54644 11089 54700 11689
rect 54804 11089 54860 11689
rect 54964 11089 55020 11689
rect 55124 11089 55180 11689
rect 55284 11089 55340 11689
rect 55572 11089 55628 11689
rect 56732 11089 56788 11689
rect 57020 11089 57076 11689
rect 57180 11089 57236 11689
rect 57340 11089 57396 11689
rect 57500 11089 57556 11689
rect 57660 11089 57716 11689
rect 57820 11089 57876 11689
rect 57980 11089 58036 11689
rect 58140 11089 58196 11689
rect 58300 11089 58356 11689
rect 58460 11089 58516 11689
rect 58620 11089 58676 11689
rect 58780 11089 58836 11689
rect 58940 11089 58996 11689
rect 59100 11089 59156 11689
rect 59260 11089 59316 11689
rect 59420 11089 59476 11689
rect 59708 11089 59764 11689
rect 52596 10029 52652 10629
rect 52884 10029 52940 10629
rect 53044 10029 53100 10629
rect 53204 10029 53260 10629
rect 53364 10029 53420 10629
rect 53524 10029 53580 10629
rect 53684 10029 53740 10629
rect 53844 10029 53900 10629
rect 54004 10029 54060 10629
rect 54164 10029 54220 10629
rect 54324 10029 54380 10629
rect 54484 10029 54540 10629
rect 54644 10029 54700 10629
rect 54804 10029 54860 10629
rect 54964 10029 55020 10629
rect 55124 10029 55180 10629
rect 55284 10029 55340 10629
rect 55572 10029 55628 10629
rect 56732 10029 56788 10629
rect 57020 10029 57076 10629
rect 57180 10029 57236 10629
rect 57340 10029 57396 10629
rect 57500 10029 57556 10629
rect 57660 10029 57716 10629
rect 57820 10029 57876 10629
rect 57980 10029 58036 10629
rect 58140 10029 58196 10629
rect 58300 10029 58356 10629
rect 58460 10029 58516 10629
rect 58620 10029 58676 10629
rect 58780 10029 58836 10629
rect 58940 10029 58996 10629
rect 59100 10029 59156 10629
rect 59260 10029 59316 10629
rect 59420 10029 59476 10629
rect 59708 10029 59764 10629
rect 52596 8969 52652 9569
rect 52884 8969 52940 9569
rect 53044 8969 53100 9569
rect 53204 8969 53260 9569
rect 53364 8969 53420 9569
rect 53524 8969 53580 9569
rect 53684 8969 53740 9569
rect 53844 8969 53900 9569
rect 54004 8969 54060 9569
rect 54164 8969 54220 9569
rect 54324 8969 54380 9569
rect 54484 8969 54540 9569
rect 54644 8969 54700 9569
rect 54804 8969 54860 9569
rect 54964 8969 55020 9569
rect 55124 8969 55180 9569
rect 55284 8969 55340 9569
rect 55572 8969 55628 9569
rect 56732 8969 56788 9569
rect 57020 8969 57076 9569
rect 57180 8969 57236 9569
rect 57340 8969 57396 9569
rect 57500 8969 57556 9569
rect 57660 8969 57716 9569
rect 57820 8969 57876 9569
rect 57980 8969 58036 9569
rect 58140 8969 58196 9569
rect 58300 8969 58356 9569
rect 58460 8969 58516 9569
rect 58620 8969 58676 9569
rect 58780 8969 58836 9569
rect 58940 8969 58996 9569
rect 59100 8969 59156 9569
rect 59260 8969 59316 9569
rect 59420 8969 59476 9569
rect 59708 8969 59764 9569
rect 52596 7909 52652 8509
rect 52884 7909 52940 8509
rect 53044 7909 53100 8509
rect 53204 7909 53260 8509
rect 53364 7909 53420 8509
rect 53524 7909 53580 8509
rect 53684 7909 53740 8509
rect 53844 7909 53900 8509
rect 54004 7909 54060 8509
rect 54164 7909 54220 8509
rect 54324 7909 54380 8509
rect 54484 7909 54540 8509
rect 54644 7909 54700 8509
rect 54804 7909 54860 8509
rect 54964 7909 55020 8509
rect 55124 7909 55180 8509
rect 55284 7909 55340 8509
rect 55572 7909 55628 8509
rect 56732 7909 56788 8509
rect 57020 7909 57076 8509
rect 57180 7909 57236 8509
rect 57340 7909 57396 8509
rect 57500 7909 57556 8509
rect 57660 7909 57716 8509
rect 57820 7909 57876 8509
rect 57980 7909 58036 8509
rect 58140 7909 58196 8509
rect 58300 7909 58356 8509
rect 58460 7909 58516 8509
rect 58620 7909 58676 8509
rect 58780 7909 58836 8509
rect 58940 7909 58996 8509
rect 59100 7909 59156 8509
rect 59260 7909 59316 8509
rect 59420 7909 59476 8509
rect 59708 7909 59764 8509
rect 62292 11089 62348 11689
rect 62580 11089 62636 11689
rect 62740 11089 62796 11689
rect 62900 11089 62956 11689
rect 63060 11089 63116 11689
rect 63220 11089 63276 11689
rect 63380 11089 63436 11689
rect 63540 11089 63596 11689
rect 63700 11089 63756 11689
rect 63860 11089 63916 11689
rect 64020 11089 64076 11689
rect 64180 11089 64236 11689
rect 64340 11089 64396 11689
rect 64500 11089 64556 11689
rect 64660 11089 64716 11689
rect 64820 11089 64876 11689
rect 64980 11089 65036 11689
rect 65268 11089 65324 11689
rect 62292 10029 62348 10629
rect 62580 10029 62636 10629
rect 62740 10029 62796 10629
rect 62900 10029 62956 10629
rect 63060 10029 63116 10629
rect 63220 10029 63276 10629
rect 63380 10029 63436 10629
rect 63540 10029 63596 10629
rect 63700 10029 63756 10629
rect 63860 10029 63916 10629
rect 64020 10029 64076 10629
rect 64180 10029 64236 10629
rect 64340 10029 64396 10629
rect 64500 10029 64556 10629
rect 64660 10029 64716 10629
rect 64820 10029 64876 10629
rect 64980 10029 65036 10629
rect 65268 10029 65324 10629
rect 62292 8969 62348 9569
rect 62580 8969 62636 9569
rect 62740 8969 62796 9569
rect 62900 8969 62956 9569
rect 63060 8969 63116 9569
rect 63220 8969 63276 9569
rect 63380 8969 63436 9569
rect 63540 8969 63596 9569
rect 63700 8969 63756 9569
rect 63860 8969 63916 9569
rect 64020 8969 64076 9569
rect 64180 8969 64236 9569
rect 64340 8969 64396 9569
rect 64500 8969 64556 9569
rect 64660 8969 64716 9569
rect 64820 8969 64876 9569
rect 64980 8969 65036 9569
rect 65268 8969 65324 9569
rect 62292 7909 62348 8509
rect 62580 7909 62636 8509
rect 62740 7909 62796 8509
rect 62900 7909 62956 8509
rect 63060 7909 63116 8509
rect 63220 7909 63276 8509
rect 63380 7909 63436 8509
rect 63540 7909 63596 8509
rect 63700 7909 63756 8509
rect 63860 7909 63916 8509
rect 64020 7909 64076 8509
rect 64180 7909 64236 8509
rect 64340 7909 64396 8509
rect 64500 7909 64556 8509
rect 64660 7909 64716 8509
rect 64820 7909 64876 8509
rect 64980 7909 65036 8509
rect 65268 7909 65324 8509
rect 1365 3634 1421 4434
rect 1653 3634 1709 4434
rect 1941 3634 2053 4434
rect 2157 3634 2269 4434
rect 2373 3634 2485 4434
rect 2589 3634 2701 4434
rect 2805 3634 2917 4434
rect 3021 3634 3133 4434
rect 3237 3634 3349 4434
rect 3453 3634 3565 4434
rect 3669 3634 3781 4434
rect 3885 3634 3997 4434
rect 4101 3634 4213 4434
rect 4317 3634 4373 4434
rect 4477 3634 4533 4434
rect 1365 2374 1421 3174
rect 1661 2374 1717 3174
rect 1949 2374 2061 3174
rect 2165 2374 2277 3174
rect 2381 2374 2493 3174
rect 2597 2374 2709 3174
rect 2813 2374 2925 3174
rect 3029 2374 3085 3174
rect 3189 2374 3245 3174
rect 3349 2374 3405 3174
rect 3509 2374 3565 3174
rect 3669 2374 3781 3174
rect 4013 2374 4125 3174
rect 4229 2374 4285 3174
rect 4525 2374 4581 3174
rect 1365 1814 1421 1914
rect 1661 1814 1717 1914
rect 1821 1814 1877 1914
rect 1981 1814 2037 1914
rect 2141 1814 2197 1914
rect 2301 1814 2357 1914
rect 2461 1814 2517 1914
rect 2621 1814 2677 1914
rect 2781 1814 2837 1914
rect 2941 1814 2997 1914
rect 3101 1814 3157 1914
rect 3261 1814 3317 1914
rect 3421 1814 3477 1914
rect 3581 1814 3637 1914
rect 3741 1814 3797 1914
rect 3901 1814 3957 1914
rect 4061 1814 4117 1914
rect 4221 1814 4421 1914
rect 4525 1814 4581 1914
rect 18870 4179 18926 4779
rect 19030 4179 19086 4779
rect 19190 4179 19246 4779
rect 19350 4179 19406 4779
rect 19510 4179 19566 4779
rect 19670 4179 19726 4779
rect 19830 4179 19886 4779
rect 19990 4179 20046 4779
rect 20150 4179 20206 4779
rect 20310 4179 20366 4779
rect 20470 4179 20526 4779
rect 20630 4179 20686 4779
rect 20790 4179 20846 4779
rect 20950 4179 21006 4779
rect 21110 4179 21166 4779
rect 21270 4179 21326 4779
rect 21430 4179 21486 4779
rect 21590 4179 21646 4779
rect 21750 4179 21806 4779
rect 22038 4179 22094 4779
rect 22326 4179 22382 4779
rect 18870 3443 18926 4043
rect 19030 3443 19086 4043
rect 19190 3443 19246 4043
rect 19350 3443 19406 4043
rect 19510 3443 19566 4043
rect 19670 3443 19726 4043
rect 19830 3443 19886 4043
rect 19990 3443 20046 4043
rect 20150 3443 20206 4043
rect 20310 3443 20366 4043
rect 20470 3443 20526 4043
rect 20630 3443 20686 4043
rect 20790 3443 20846 4043
rect 20950 3443 21006 4043
rect 21110 3443 21166 4043
rect 21270 3443 21326 4043
rect 21430 3443 21486 4043
rect 21590 3443 21646 4043
rect 21750 3443 21806 4043
rect 22038 3443 22094 4043
rect 22326 3443 22382 4043
rect 18870 2707 18926 3307
rect 19030 2707 19086 3307
rect 19190 2707 19246 3307
rect 19350 2707 19406 3307
rect 19510 2707 19566 3307
rect 19670 2707 19726 3307
rect 19830 2707 19886 3307
rect 19990 2707 20046 3307
rect 20150 2707 20206 3307
rect 20310 2707 20366 3307
rect 20470 2707 20526 3307
rect 20630 2707 20686 3307
rect 20790 2707 20846 3307
rect 20950 2707 21006 3307
rect 21110 2707 21166 3307
rect 21270 2707 21326 3307
rect 21430 2707 21486 3307
rect 21590 2707 21646 3307
rect 21750 2707 21806 3307
rect 22038 2707 22094 3207
rect 22326 2707 22382 3307
rect 18870 1971 18926 2571
rect 19030 1971 19086 2571
rect 19190 1971 19246 2571
rect 19350 1971 19406 2571
rect 19510 1971 19566 2571
rect 19670 1971 19726 2571
rect 19830 1971 19886 2571
rect 19990 1971 20046 2571
rect 20150 1971 20206 2571
rect 20310 1971 20366 2571
rect 20470 1971 20526 2571
rect 20630 1971 20686 2571
rect 20790 1971 20846 2571
rect 20950 1971 21006 2571
rect 21110 1971 21166 2571
rect 21270 1971 21326 2571
rect 21430 1971 21486 2571
rect 21590 1971 21646 2571
rect 21750 1971 21806 2571
rect 22038 1971 22094 2471
rect 22326 1971 22382 2571
<< ndiff >>
rect 6449 14263 6537 14276
rect 6449 13713 6462 14263
rect 6508 13713 6537 14263
rect 6449 13700 6537 13713
rect 6593 14263 6681 14276
rect 6593 13713 6622 14263
rect 6668 13713 6681 14263
rect 6593 13700 6681 13713
rect 6737 14263 6825 14276
rect 6737 13713 6750 14263
rect 6796 13713 6825 14263
rect 6737 13700 6825 13713
rect 6881 14263 6985 14276
rect 6881 13713 6910 14263
rect 6956 13713 6985 14263
rect 6881 13700 6985 13713
rect 7041 14263 7145 14276
rect 7041 13713 7070 14263
rect 7116 13713 7145 14263
rect 7041 13700 7145 13713
rect 7201 14263 7305 14276
rect 7201 13713 7230 14263
rect 7276 13713 7305 14263
rect 7201 13700 7305 13713
rect 7361 14263 7465 14276
rect 7361 13713 7390 14263
rect 7436 13713 7465 14263
rect 7361 13700 7465 13713
rect 7521 14263 7625 14276
rect 7521 13713 7550 14263
rect 7596 13713 7625 14263
rect 7521 13700 7625 13713
rect 7681 14263 7785 14276
rect 7681 13713 7710 14263
rect 7756 13713 7785 14263
rect 7681 13700 7785 13713
rect 7841 14263 7945 14276
rect 7841 13713 7870 14263
rect 7916 13713 7945 14263
rect 7841 13700 7945 13713
rect 8001 14263 8089 14276
rect 8001 13713 8030 14263
rect 8076 13713 8089 14263
rect 8001 13700 8089 13713
rect 8145 14263 8233 14276
rect 8145 13713 8158 14263
rect 8204 13713 8233 14263
rect 8145 13700 8233 13713
rect 8289 14263 8377 14276
rect 8289 13713 8318 14263
rect 8364 13713 8377 14263
rect 8289 13700 8377 13713
rect 6449 13401 6537 13414
rect 6449 12851 6462 13401
rect 6508 12851 6537 13401
rect 6449 12838 6537 12851
rect 6593 13401 6681 13414
rect 6593 12851 6622 13401
rect 6668 12851 6681 13401
rect 6593 12838 6681 12851
rect 6737 13401 6825 13414
rect 6737 12851 6750 13401
rect 6796 12851 6825 13401
rect 6737 12838 6825 12851
rect 6881 13401 6985 13414
rect 6881 12851 6910 13401
rect 6956 12851 6985 13401
rect 6881 12838 6985 12851
rect 7041 13401 7145 13414
rect 7041 12851 7070 13401
rect 7116 12851 7145 13401
rect 7041 12838 7145 12851
rect 7201 13401 7305 13414
rect 7201 12851 7230 13401
rect 7276 12851 7305 13401
rect 7201 12838 7305 12851
rect 7361 13401 7465 13414
rect 7361 12851 7390 13401
rect 7436 12851 7465 13401
rect 7361 12838 7465 12851
rect 7521 13401 7625 13414
rect 7521 12851 7550 13401
rect 7596 12851 7625 13401
rect 7521 12838 7625 12851
rect 7681 13401 7785 13414
rect 7681 12851 7710 13401
rect 7756 12851 7785 13401
rect 7681 12838 7785 12851
rect 7841 13401 7945 13414
rect 7841 12851 7870 13401
rect 7916 12851 7945 13401
rect 7841 12838 7945 12851
rect 8001 13401 8089 13414
rect 8001 12851 8030 13401
rect 8076 12851 8089 13401
rect 8001 12838 8089 12851
rect 8145 13401 8233 13414
rect 8145 12851 8158 13401
rect 8204 12851 8233 13401
rect 8145 12838 8233 12851
rect 8289 13401 8377 13414
rect 8289 12851 8318 13401
rect 8364 12851 8377 13401
rect 8289 12838 8377 12851
rect 6449 12539 6537 12552
rect 6449 11989 6462 12539
rect 6508 11989 6537 12539
rect 6449 11976 6537 11989
rect 6593 12539 6681 12552
rect 6593 11989 6622 12539
rect 6668 11989 6681 12539
rect 6593 11976 6681 11989
rect 6737 12539 6825 12552
rect 6737 11989 6750 12539
rect 6796 11989 6825 12539
rect 6737 11976 6825 11989
rect 6881 12539 6985 12552
rect 6881 11989 6910 12539
rect 6956 11989 6985 12539
rect 6881 11976 6985 11989
rect 7041 12539 7145 12552
rect 7041 11989 7070 12539
rect 7116 11989 7145 12539
rect 7041 11976 7145 11989
rect 7201 12539 7305 12552
rect 7201 11989 7230 12539
rect 7276 11989 7305 12539
rect 7201 11976 7305 11989
rect 7361 12539 7465 12552
rect 7361 11989 7390 12539
rect 7436 11989 7465 12539
rect 7361 11976 7465 11989
rect 7521 12539 7625 12552
rect 7521 11989 7550 12539
rect 7596 11989 7625 12539
rect 7521 11976 7625 11989
rect 7681 12539 7785 12552
rect 7681 11989 7710 12539
rect 7756 11989 7785 12539
rect 7681 11976 7785 11989
rect 7841 12539 7945 12552
rect 7841 11989 7870 12539
rect 7916 11989 7945 12539
rect 7841 11976 7945 11989
rect 8001 12539 8089 12552
rect 8001 11989 8030 12539
rect 8076 11989 8089 12539
rect 8001 11976 8089 11989
rect 8145 12539 8233 12552
rect 8145 11989 8158 12539
rect 8204 11989 8233 12539
rect 8145 11976 8233 11989
rect 8289 12539 8377 12552
rect 8289 11989 8318 12539
rect 8364 11989 8377 12539
rect 8289 11976 8377 11989
rect 18699 13176 18787 13189
rect 18699 12602 18712 13176
rect 18758 12602 18787 13176
rect 18699 12589 18787 12602
rect 18843 13176 18931 13189
rect 18843 12602 18872 13176
rect 18918 12602 18931 13176
rect 18843 12589 18931 12602
rect 18987 13176 19075 13189
rect 18987 12602 19000 13176
rect 19046 12602 19075 13176
rect 18987 12589 19075 12602
rect 19131 13176 19235 13189
rect 19131 12602 19160 13176
rect 19206 12602 19235 13176
rect 19131 12589 19235 12602
rect 19291 13176 19395 13189
rect 19291 12602 19320 13176
rect 19366 12602 19395 13176
rect 19291 12589 19395 12602
rect 19451 13176 19555 13189
rect 19451 12602 19480 13176
rect 19526 12602 19555 13176
rect 19451 12589 19555 12602
rect 19611 13176 19715 13189
rect 19611 12602 19640 13176
rect 19686 12602 19715 13176
rect 19611 12589 19715 12602
rect 19771 13176 19875 13189
rect 19771 12602 19800 13176
rect 19846 12602 19875 13176
rect 19771 12589 19875 12602
rect 19931 13176 20035 13189
rect 19931 12602 19960 13176
rect 20006 12602 20035 13176
rect 19931 12589 20035 12602
rect 20091 13176 20195 13189
rect 20091 12602 20120 13176
rect 20166 12602 20195 13176
rect 20091 12589 20195 12602
rect 20251 13176 20339 13189
rect 20251 12602 20280 13176
rect 20326 12602 20339 13176
rect 20251 12589 20339 12602
rect 20395 13176 20483 13189
rect 20395 12602 20408 13176
rect 20454 12602 20483 13176
rect 20395 12589 20483 12602
rect 20539 13176 20627 13189
rect 20539 12602 20568 13176
rect 20614 12602 20627 13176
rect 20539 12589 20627 12602
rect 6449 11677 6537 11690
rect 6449 11127 6462 11677
rect 6508 11127 6537 11677
rect 6449 11114 6537 11127
rect 6593 11677 6681 11690
rect 6593 11127 6622 11677
rect 6668 11127 6681 11677
rect 6593 11114 6681 11127
rect 6737 11677 6825 11690
rect 6737 11127 6750 11677
rect 6796 11127 6825 11677
rect 6737 11114 6825 11127
rect 6881 11677 6985 11690
rect 6881 11127 6910 11677
rect 6956 11127 6985 11677
rect 6881 11114 6985 11127
rect 7041 11677 7145 11690
rect 7041 11127 7070 11677
rect 7116 11127 7145 11677
rect 7041 11114 7145 11127
rect 7201 11677 7305 11690
rect 7201 11127 7230 11677
rect 7276 11127 7305 11677
rect 7201 11114 7305 11127
rect 7361 11677 7465 11690
rect 7361 11127 7390 11677
rect 7436 11127 7465 11677
rect 7361 11114 7465 11127
rect 7521 11677 7625 11690
rect 7521 11127 7550 11677
rect 7596 11127 7625 11677
rect 7521 11114 7625 11127
rect 7681 11677 7785 11690
rect 7681 11127 7710 11677
rect 7756 11127 7785 11677
rect 7681 11114 7785 11127
rect 7841 11677 7945 11690
rect 7841 11127 7870 11677
rect 7916 11127 7945 11677
rect 7841 11114 7945 11127
rect 8001 11677 8089 11690
rect 8001 11127 8030 11677
rect 8076 11127 8089 11677
rect 8001 11114 8089 11127
rect 8145 11677 8233 11690
rect 8145 11127 8158 11677
rect 8204 11127 8233 11677
rect 8145 11114 8233 11127
rect 8289 11677 8377 11690
rect 8289 11127 8318 11677
rect 8364 11127 8377 11677
rect 8289 11114 8377 11127
rect 6449 10815 6537 10828
rect 6449 10265 6462 10815
rect 6508 10265 6537 10815
rect 6449 10252 6537 10265
rect 6593 10815 6681 10828
rect 6593 10265 6622 10815
rect 6668 10265 6681 10815
rect 6593 10252 6681 10265
rect 6737 10815 6825 10828
rect 6737 10265 6750 10815
rect 6796 10265 6825 10815
rect 6737 10252 6825 10265
rect 6881 10815 6985 10828
rect 6881 10265 6910 10815
rect 6956 10265 6985 10815
rect 6881 10252 6985 10265
rect 7041 10815 7145 10828
rect 7041 10265 7070 10815
rect 7116 10265 7145 10815
rect 7041 10252 7145 10265
rect 7201 10815 7305 10828
rect 7201 10265 7230 10815
rect 7276 10265 7305 10815
rect 7201 10252 7305 10265
rect 7361 10815 7465 10828
rect 7361 10265 7390 10815
rect 7436 10265 7465 10815
rect 7361 10252 7465 10265
rect 7521 10815 7625 10828
rect 7521 10265 7550 10815
rect 7596 10265 7625 10815
rect 7521 10252 7625 10265
rect 7681 10815 7785 10828
rect 7681 10265 7710 10815
rect 7756 10265 7785 10815
rect 7681 10252 7785 10265
rect 7841 10815 7945 10828
rect 7841 10265 7870 10815
rect 7916 10265 7945 10815
rect 7841 10252 7945 10265
rect 8001 10815 8089 10828
rect 8001 10265 8030 10815
rect 8076 10265 8089 10815
rect 8001 10252 8089 10265
rect 8145 10815 8233 10828
rect 8145 10265 8158 10815
rect 8204 10265 8233 10815
rect 8145 10252 8233 10265
rect 8289 10815 8377 10828
rect 8289 10265 8318 10815
rect 8364 10265 8377 10815
rect 8289 10252 8377 10265
rect 8684 10796 8772 10809
rect 8684 10246 8697 10796
rect 8743 10246 8772 10796
rect 8684 10233 8772 10246
rect 8828 10796 8916 10809
rect 8828 10246 8857 10796
rect 8903 10246 8916 10796
rect 8828 10233 8916 10246
rect 8972 10796 9060 10809
rect 8972 10246 8985 10796
rect 9031 10246 9060 10796
rect 8972 10233 9060 10246
rect 9116 10796 9204 10809
rect 9116 10246 9145 10796
rect 9191 10246 9204 10796
rect 9116 10233 9204 10246
rect 9260 10796 9348 10809
rect 9260 10246 9273 10796
rect 9319 10246 9348 10796
rect 9260 10233 9348 10246
rect 9404 10796 9508 10809
rect 9404 10246 9433 10796
rect 9479 10246 9508 10796
rect 9404 10233 9508 10246
rect 9564 10796 9652 10809
rect 9564 10246 9593 10796
rect 9639 10246 9652 10796
rect 9564 10233 9652 10246
rect 9708 10796 9796 10809
rect 9708 10246 9721 10796
rect 9767 10246 9796 10796
rect 9708 10233 9796 10246
rect 9852 10796 9956 10809
rect 9852 10246 9881 10796
rect 9927 10246 9956 10796
rect 9852 10233 9956 10246
rect 10012 10796 10100 10809
rect 10012 10246 10041 10796
rect 10087 10246 10100 10796
rect 10012 10233 10100 10246
rect 10156 10796 10244 10809
rect 10156 10246 10169 10796
rect 10215 10246 10244 10796
rect 10156 10233 10244 10246
rect 10300 10796 10404 10809
rect 10300 10246 10329 10796
rect 10375 10246 10404 10796
rect 10300 10233 10404 10246
rect 10460 10796 10548 10809
rect 10460 10246 10489 10796
rect 10535 10246 10548 10796
rect 10460 10233 10548 10246
rect 10604 10796 10692 10809
rect 10604 10246 10617 10796
rect 10663 10246 10692 10796
rect 10604 10233 10692 10246
rect 10748 10796 10836 10809
rect 10748 10246 10777 10796
rect 10823 10246 10836 10796
rect 10748 10233 10836 10246
rect 10892 10796 10980 10809
rect 10892 10246 10905 10796
rect 10951 10246 10980 10796
rect 10892 10233 10980 10246
rect 11036 10796 11124 10809
rect 11036 10246 11065 10796
rect 11111 10246 11124 10796
rect 11036 10233 11124 10246
rect 6449 9953 6537 9966
rect 6449 9403 6462 9953
rect 6508 9403 6537 9953
rect 6449 9390 6537 9403
rect 6593 9953 6681 9966
rect 6593 9403 6622 9953
rect 6668 9403 6681 9953
rect 6593 9390 6681 9403
rect 6737 9953 6825 9966
rect 6737 9403 6750 9953
rect 6796 9403 6825 9953
rect 6737 9390 6825 9403
rect 6881 9953 6985 9966
rect 6881 9403 6910 9953
rect 6956 9403 6985 9953
rect 6881 9390 6985 9403
rect 7041 9953 7145 9966
rect 7041 9403 7070 9953
rect 7116 9403 7145 9953
rect 7041 9390 7145 9403
rect 7201 9953 7305 9966
rect 7201 9403 7230 9953
rect 7276 9403 7305 9953
rect 7201 9390 7305 9403
rect 7361 9953 7465 9966
rect 7361 9403 7390 9953
rect 7436 9403 7465 9953
rect 7361 9390 7465 9403
rect 7521 9953 7625 9966
rect 7521 9403 7550 9953
rect 7596 9403 7625 9953
rect 7521 9390 7625 9403
rect 7681 9953 7785 9966
rect 7681 9403 7710 9953
rect 7756 9403 7785 9953
rect 7681 9390 7785 9403
rect 7841 9953 7945 9966
rect 7841 9403 7870 9953
rect 7916 9403 7945 9953
rect 7841 9390 7945 9403
rect 8001 9953 8089 9966
rect 8001 9403 8030 9953
rect 8076 9403 8089 9953
rect 8001 9390 8089 9403
rect 8145 9953 8233 9966
rect 8145 9403 8158 9953
rect 8204 9403 8233 9953
rect 8145 9390 8233 9403
rect 8289 9953 8377 9966
rect 8289 9403 8318 9953
rect 8364 9403 8377 9953
rect 8289 9390 8377 9403
rect 8684 9934 8772 9947
rect 8684 9384 8697 9934
rect 8743 9384 8772 9934
rect 8684 9371 8772 9384
rect 8828 9934 8916 9947
rect 8828 9384 8857 9934
rect 8903 9384 8916 9934
rect 8828 9371 8916 9384
rect 8972 9934 9060 9947
rect 8972 9384 8985 9934
rect 9031 9384 9060 9934
rect 8972 9371 9060 9384
rect 9116 9934 9204 9947
rect 9116 9384 9145 9934
rect 9191 9384 9204 9934
rect 9116 9371 9204 9384
rect 9260 9934 9348 9947
rect 9260 9384 9273 9934
rect 9319 9384 9348 9934
rect 9260 9371 9348 9384
rect 9404 9934 9508 9947
rect 9404 9384 9433 9934
rect 9479 9384 9508 9934
rect 9404 9371 9508 9384
rect 9564 9934 9652 9947
rect 9564 9384 9593 9934
rect 9639 9384 9652 9934
rect 9564 9371 9652 9384
rect 9708 9934 9796 9947
rect 9708 9384 9721 9934
rect 9767 9384 9796 9934
rect 9708 9371 9796 9384
rect 9852 9934 9956 9947
rect 9852 9384 9881 9934
rect 9927 9384 9956 9934
rect 9852 9371 9956 9384
rect 10012 9934 10100 9947
rect 10012 9384 10041 9934
rect 10087 9384 10100 9934
rect 10012 9371 10100 9384
rect 10156 9934 10244 9947
rect 10156 9384 10169 9934
rect 10215 9384 10244 9934
rect 10156 9371 10244 9384
rect 10300 9934 10404 9947
rect 10300 9384 10329 9934
rect 10375 9384 10404 9934
rect 10300 9371 10404 9384
rect 10460 9934 10548 9947
rect 10460 9384 10489 9934
rect 10535 9384 10548 9934
rect 10460 9371 10548 9384
rect 10604 9934 10692 9947
rect 10604 9384 10617 9934
rect 10663 9384 10692 9934
rect 10604 9371 10692 9384
rect 10748 9934 10836 9947
rect 10748 9384 10777 9934
rect 10823 9384 10836 9934
rect 10748 9371 10836 9384
rect 10892 9934 10980 9947
rect 10892 9384 10905 9934
rect 10951 9384 10980 9934
rect 10892 9371 10980 9384
rect 11036 9934 11124 9947
rect 11036 9384 11065 9934
rect 11111 9384 11124 9934
rect 11036 9371 11124 9384
rect 6449 9091 6537 9104
rect 6449 8541 6462 9091
rect 6508 8541 6537 9091
rect 6449 8528 6537 8541
rect 6593 9091 6681 9104
rect 6593 8541 6622 9091
rect 6668 8541 6681 9091
rect 6593 8528 6681 8541
rect 6737 9091 6825 9104
rect 6737 8541 6750 9091
rect 6796 8541 6825 9091
rect 6737 8528 6825 8541
rect 6881 9091 6985 9104
rect 6881 8541 6910 9091
rect 6956 8541 6985 9091
rect 6881 8528 6985 8541
rect 7041 9091 7145 9104
rect 7041 8541 7070 9091
rect 7116 8541 7145 9091
rect 7041 8528 7145 8541
rect 7201 9091 7305 9104
rect 7201 8541 7230 9091
rect 7276 8541 7305 9091
rect 7201 8528 7305 8541
rect 7361 9091 7465 9104
rect 7361 8541 7390 9091
rect 7436 8541 7465 9091
rect 7361 8528 7465 8541
rect 7521 9091 7625 9104
rect 7521 8541 7550 9091
rect 7596 8541 7625 9091
rect 7521 8528 7625 8541
rect 7681 9091 7785 9104
rect 7681 8541 7710 9091
rect 7756 8541 7785 9091
rect 7681 8528 7785 8541
rect 7841 9091 7945 9104
rect 7841 8541 7870 9091
rect 7916 8541 7945 9091
rect 7841 8528 7945 8541
rect 8001 9091 8089 9104
rect 8001 8541 8030 9091
rect 8076 8541 8089 9091
rect 8001 8528 8089 8541
rect 8145 9091 8233 9104
rect 8145 8541 8158 9091
rect 8204 8541 8233 9091
rect 8145 8528 8233 8541
rect 8289 9091 8377 9104
rect 8289 8541 8318 9091
rect 8364 8541 8377 9091
rect 8289 8528 8377 8541
rect 8684 9072 8772 9085
rect 8684 8522 8697 9072
rect 8743 8522 8772 9072
rect 8684 8509 8772 8522
rect 8828 9072 8916 9085
rect 8828 8522 8857 9072
rect 8903 8522 8916 9072
rect 8828 8509 8916 8522
rect 8972 9072 9060 9085
rect 8972 8522 8985 9072
rect 9031 8522 9060 9072
rect 8972 8509 9060 8522
rect 9116 9072 9204 9085
rect 9116 8522 9145 9072
rect 9191 8522 9204 9072
rect 9116 8509 9204 8522
rect 9260 9072 9348 9085
rect 9260 8522 9273 9072
rect 9319 8522 9348 9072
rect 9260 8509 9348 8522
rect 9404 9072 9508 9085
rect 9404 8522 9433 9072
rect 9479 8522 9508 9072
rect 9404 8509 9508 8522
rect 9564 9072 9652 9085
rect 9564 8522 9593 9072
rect 9639 8522 9652 9072
rect 9564 8509 9652 8522
rect 9708 9072 9796 9085
rect 9708 8522 9721 9072
rect 9767 8522 9796 9072
rect 9708 8509 9796 8522
rect 9852 9072 9956 9085
rect 9852 8522 9881 9072
rect 9927 8522 9956 9072
rect 9852 8509 9956 8522
rect 10012 9072 10100 9085
rect 10012 8522 10041 9072
rect 10087 8522 10100 9072
rect 10012 8509 10100 8522
rect 10156 9072 10244 9085
rect 10156 8522 10169 9072
rect 10215 8522 10244 9072
rect 10156 8509 10244 8522
rect 10300 9072 10404 9085
rect 10300 8522 10329 9072
rect 10375 8522 10404 9072
rect 10300 8509 10404 8522
rect 10460 9072 10548 9085
rect 10460 8522 10489 9072
rect 10535 8522 10548 9072
rect 10460 8509 10548 8522
rect 10604 9072 10692 9085
rect 10604 8522 10617 9072
rect 10663 8522 10692 9072
rect 10604 8509 10692 8522
rect 10748 9072 10836 9085
rect 10748 8522 10777 9072
rect 10823 8522 10836 9072
rect 10748 8509 10836 8522
rect 10892 9072 10980 9085
rect 10892 8522 10905 9072
rect 10951 8522 10980 9072
rect 10892 8509 10980 8522
rect 11036 9072 11124 9085
rect 11036 8522 11065 9072
rect 11111 8522 11124 9072
rect 11036 8509 11124 8522
rect 6449 8229 6537 8242
rect 6449 7679 6462 8229
rect 6508 7679 6537 8229
rect 6449 7666 6537 7679
rect 6593 8229 6681 8242
rect 6593 7679 6622 8229
rect 6668 7679 6681 8229
rect 6593 7666 6681 7679
rect 6737 8229 6825 8242
rect 6737 7679 6750 8229
rect 6796 7679 6825 8229
rect 6737 7666 6825 7679
rect 6881 8229 6985 8242
rect 6881 7679 6910 8229
rect 6956 7679 6985 8229
rect 6881 7666 6985 7679
rect 7041 8229 7145 8242
rect 7041 7679 7070 8229
rect 7116 7679 7145 8229
rect 7041 7666 7145 7679
rect 7201 8229 7305 8242
rect 7201 7679 7230 8229
rect 7276 7679 7305 8229
rect 7201 7666 7305 7679
rect 7361 8229 7465 8242
rect 7361 7679 7390 8229
rect 7436 7679 7465 8229
rect 7361 7666 7465 7679
rect 7521 8229 7625 8242
rect 7521 7679 7550 8229
rect 7596 7679 7625 8229
rect 7521 7666 7625 7679
rect 7681 8229 7785 8242
rect 7681 7679 7710 8229
rect 7756 7679 7785 8229
rect 7681 7666 7785 7679
rect 7841 8229 7945 8242
rect 7841 7679 7870 8229
rect 7916 7679 7945 8229
rect 7841 7666 7945 7679
rect 8001 8229 8089 8242
rect 8001 7679 8030 8229
rect 8076 7679 8089 8229
rect 8001 7666 8089 7679
rect 8145 8229 8233 8242
rect 8145 7679 8158 8229
rect 8204 7679 8233 8229
rect 8145 7666 8233 7679
rect 8289 8229 8377 8242
rect 8289 7679 8318 8229
rect 8364 7679 8377 8229
rect 8289 7666 8377 7679
rect 8684 8210 8772 8223
rect 8684 7660 8697 8210
rect 8743 7660 8772 8210
rect 8684 7647 8772 7660
rect 8828 8210 8916 8223
rect 8828 7660 8857 8210
rect 8903 7660 8916 8210
rect 8828 7647 8916 7660
rect 8972 8210 9060 8223
rect 8972 7660 8985 8210
rect 9031 7660 9060 8210
rect 8972 7647 9060 7660
rect 9116 8210 9204 8223
rect 9116 7660 9145 8210
rect 9191 7660 9204 8210
rect 9116 7647 9204 7660
rect 9260 8210 9348 8223
rect 9260 7660 9273 8210
rect 9319 7660 9348 8210
rect 9260 7647 9348 7660
rect 9404 8210 9508 8223
rect 9404 7660 9433 8210
rect 9479 7660 9508 8210
rect 9404 7647 9508 7660
rect 9564 8210 9652 8223
rect 9564 7660 9593 8210
rect 9639 7660 9652 8210
rect 9564 7647 9652 7660
rect 9708 8210 9796 8223
rect 9708 7660 9721 8210
rect 9767 7660 9796 8210
rect 9708 7647 9796 7660
rect 9852 8210 9956 8223
rect 9852 7660 9881 8210
rect 9927 7660 9956 8210
rect 9852 7647 9956 7660
rect 10012 8210 10100 8223
rect 10012 7660 10041 8210
rect 10087 7660 10100 8210
rect 10012 7647 10100 7660
rect 10156 8210 10244 8223
rect 10156 7660 10169 8210
rect 10215 7660 10244 8210
rect 10156 7647 10244 7660
rect 10300 8210 10404 8223
rect 10300 7660 10329 8210
rect 10375 7660 10404 8210
rect 10300 7647 10404 7660
rect 10460 8210 10548 8223
rect 10460 7660 10489 8210
rect 10535 7660 10548 8210
rect 10460 7647 10548 7660
rect 10604 8210 10692 8223
rect 10604 7660 10617 8210
rect 10663 7660 10692 8210
rect 10604 7647 10692 7660
rect 10748 8210 10836 8223
rect 10748 7660 10777 8210
rect 10823 7660 10836 8210
rect 10748 7647 10836 7660
rect 10892 8210 10980 8223
rect 10892 7660 10905 8210
rect 10951 7660 10980 8210
rect 10892 7647 10980 7660
rect 11036 8210 11124 8223
rect 11036 7660 11065 8210
rect 11111 7660 11124 8210
rect 11036 7647 11124 7660
rect 18699 12240 18787 12253
rect 18699 11666 18712 12240
rect 18758 11666 18787 12240
rect 18699 11653 18787 11666
rect 18843 12240 18931 12253
rect 18843 11666 18872 12240
rect 18918 11666 18931 12240
rect 18843 11653 18931 11666
rect 18987 12240 19075 12253
rect 18987 11666 19000 12240
rect 19046 11666 19075 12240
rect 18987 11653 19075 11666
rect 19131 12240 19235 12253
rect 19131 11666 19160 12240
rect 19206 11666 19235 12240
rect 19131 11653 19235 11666
rect 19291 12240 19395 12253
rect 19291 11666 19320 12240
rect 19366 11666 19395 12240
rect 19291 11653 19395 11666
rect 19451 12240 19555 12253
rect 19451 11666 19480 12240
rect 19526 11666 19555 12240
rect 19451 11653 19555 11666
rect 19611 12240 19715 12253
rect 19611 11666 19640 12240
rect 19686 11666 19715 12240
rect 19611 11653 19715 11666
rect 19771 12240 19875 12253
rect 19771 11666 19800 12240
rect 19846 11666 19875 12240
rect 19771 11653 19875 11666
rect 19931 12240 20035 12253
rect 19931 11666 19960 12240
rect 20006 11666 20035 12240
rect 19931 11653 20035 11666
rect 20091 12240 20195 12253
rect 20091 11666 20120 12240
rect 20166 11666 20195 12240
rect 20091 11653 20195 11666
rect 20251 12240 20339 12253
rect 20251 11666 20280 12240
rect 20326 11666 20339 12240
rect 20251 11653 20339 11666
rect 20395 12240 20483 12253
rect 20395 11666 20408 12240
rect 20454 11666 20483 12240
rect 20395 11653 20483 11666
rect 20539 12240 20627 12253
rect 20539 11666 20568 12240
rect 20614 11666 20627 12240
rect 20539 11653 20627 11666
rect 18699 11304 18787 11317
rect 18699 10730 18712 11304
rect 18758 10730 18787 11304
rect 18699 10717 18787 10730
rect 18843 11304 18931 11317
rect 18843 10730 18872 11304
rect 18918 10730 18931 11304
rect 18843 10717 18931 10730
rect 18987 11304 19075 11317
rect 18987 10730 19000 11304
rect 19046 10730 19075 11304
rect 18987 10717 19075 10730
rect 19131 11304 19235 11317
rect 19131 10730 19160 11304
rect 19206 10730 19235 11304
rect 19131 10717 19235 10730
rect 19291 11304 19395 11317
rect 19291 10730 19320 11304
rect 19366 10730 19395 11304
rect 19291 10717 19395 10730
rect 19451 11304 19555 11317
rect 19451 10730 19480 11304
rect 19526 10730 19555 11304
rect 19451 10717 19555 10730
rect 19611 11304 19715 11317
rect 19611 10730 19640 11304
rect 19686 10730 19715 11304
rect 19611 10717 19715 10730
rect 19771 11304 19875 11317
rect 19771 10730 19800 11304
rect 19846 10730 19875 11304
rect 19771 10717 19875 10730
rect 19931 11304 20035 11317
rect 19931 10730 19960 11304
rect 20006 10730 20035 11304
rect 19931 10717 20035 10730
rect 20091 11304 20195 11317
rect 20091 10730 20120 11304
rect 20166 10730 20195 11304
rect 20091 10717 20195 10730
rect 20251 11304 20339 11317
rect 20251 10730 20280 11304
rect 20326 10730 20339 11304
rect 20251 10717 20339 10730
rect 20395 11304 20483 11317
rect 20395 10730 20408 11304
rect 20454 10730 20483 11304
rect 20395 10717 20483 10730
rect 20539 11304 20627 11317
rect 20539 10730 20568 11304
rect 20614 10730 20627 11304
rect 20539 10717 20627 10730
rect 18699 10368 18787 10381
rect 18699 9794 18712 10368
rect 18758 9794 18787 10368
rect 18699 9781 18787 9794
rect 18843 10368 18931 10381
rect 18843 9794 18872 10368
rect 18918 9794 18931 10368
rect 18843 9781 18931 9794
rect 18987 10368 19075 10381
rect 18987 9794 19000 10368
rect 19046 9794 19075 10368
rect 18987 9781 19075 9794
rect 19131 10368 19235 10381
rect 19131 9794 19160 10368
rect 19206 9794 19235 10368
rect 19131 9781 19235 9794
rect 19291 10368 19395 10381
rect 19291 9794 19320 10368
rect 19366 9794 19395 10368
rect 19291 9781 19395 9794
rect 19451 10368 19555 10381
rect 19451 9794 19480 10368
rect 19526 9794 19555 10368
rect 19451 9781 19555 9794
rect 19611 10368 19715 10381
rect 19611 9794 19640 10368
rect 19686 9794 19715 10368
rect 19611 9781 19715 9794
rect 19771 10368 19875 10381
rect 19771 9794 19800 10368
rect 19846 9794 19875 10368
rect 19771 9781 19875 9794
rect 19931 10368 20035 10381
rect 19931 9794 19960 10368
rect 20006 9794 20035 10368
rect 19931 9781 20035 9794
rect 20091 10368 20195 10381
rect 20091 9794 20120 10368
rect 20166 9794 20195 10368
rect 20091 9781 20195 9794
rect 20251 10368 20339 10381
rect 20251 9794 20280 10368
rect 20326 9794 20339 10368
rect 20251 9781 20339 9794
rect 20395 10368 20483 10381
rect 20395 9794 20408 10368
rect 20454 9794 20483 10368
rect 20395 9781 20483 9794
rect 20539 10368 20627 10381
rect 20539 9794 20568 10368
rect 20614 9794 20627 10368
rect 20539 9781 20627 9794
rect 18699 9432 18787 9445
rect 18699 8858 18712 9432
rect 18758 8858 18787 9432
rect 18699 8845 18787 8858
rect 18843 9432 18931 9445
rect 18843 8858 18872 9432
rect 18918 8858 18931 9432
rect 18843 8845 18931 8858
rect 18987 9432 19075 9445
rect 18987 8858 19000 9432
rect 19046 8858 19075 9432
rect 18987 8845 19075 8858
rect 19131 9432 19235 9445
rect 19131 8858 19160 9432
rect 19206 8858 19235 9432
rect 19131 8845 19235 8858
rect 19291 9432 19395 9445
rect 19291 8858 19320 9432
rect 19366 8858 19395 9432
rect 19291 8845 19395 8858
rect 19451 9432 19555 9445
rect 19451 8858 19480 9432
rect 19526 8858 19555 9432
rect 19451 8845 19555 8858
rect 19611 9432 19715 9445
rect 19611 8858 19640 9432
rect 19686 8858 19715 9432
rect 19611 8845 19715 8858
rect 19771 9432 19875 9445
rect 19771 8858 19800 9432
rect 19846 8858 19875 9432
rect 19771 8845 19875 8858
rect 19931 9432 20035 9445
rect 19931 8858 19960 9432
rect 20006 8858 20035 9432
rect 19931 8845 20035 8858
rect 20091 9432 20195 9445
rect 20091 8858 20120 9432
rect 20166 8858 20195 9432
rect 20091 8845 20195 8858
rect 20251 9432 20339 9445
rect 20251 8858 20280 9432
rect 20326 8858 20339 9432
rect 20251 8845 20339 8858
rect 20395 9432 20483 9445
rect 20395 8858 20408 9432
rect 20454 8858 20483 9432
rect 20395 8845 20483 8858
rect 20539 9432 20627 9445
rect 20539 8858 20568 9432
rect 20614 8858 20627 9432
rect 20539 8845 20627 8858
rect 18699 8496 18787 8509
rect 18699 7922 18712 8496
rect 18758 7922 18787 8496
rect 18699 7909 18787 7922
rect 18843 8496 18931 8509
rect 18843 7922 18872 8496
rect 18918 7922 18931 8496
rect 18843 7909 18931 7922
rect 18987 8496 19075 8509
rect 18987 7922 19000 8496
rect 19046 7922 19075 8496
rect 18987 7909 19075 7922
rect 19131 8496 19235 8509
rect 19131 7922 19160 8496
rect 19206 7922 19235 8496
rect 19131 7909 19235 7922
rect 19291 8496 19395 8509
rect 19291 7922 19320 8496
rect 19366 7922 19395 8496
rect 19291 7909 19395 7922
rect 19451 8496 19555 8509
rect 19451 7922 19480 8496
rect 19526 7922 19555 8496
rect 19451 7909 19555 7922
rect 19611 8496 19715 8509
rect 19611 7922 19640 8496
rect 19686 7922 19715 8496
rect 19611 7909 19715 7922
rect 19771 8496 19875 8509
rect 19771 7922 19800 8496
rect 19846 7922 19875 8496
rect 19771 7909 19875 7922
rect 19931 8496 20035 8509
rect 19931 7922 19960 8496
rect 20006 7922 20035 8496
rect 19931 7909 20035 7922
rect 20091 8496 20195 8509
rect 20091 7922 20120 8496
rect 20166 7922 20195 8496
rect 20091 7909 20195 7922
rect 20251 8496 20339 8509
rect 20251 7922 20280 8496
rect 20326 7922 20339 8496
rect 20251 7909 20339 7922
rect 20395 8496 20483 8509
rect 20395 7922 20408 8496
rect 20454 7922 20483 8496
rect 20395 7909 20483 7922
rect 20539 8496 20627 8509
rect 20539 7922 20568 8496
rect 20614 7922 20627 8496
rect 20539 7909 20627 7922
rect 23851 13176 23939 13189
rect 23851 12602 23864 13176
rect 23910 12602 23939 13176
rect 23851 12589 23939 12602
rect 23995 13176 24083 13189
rect 23995 12602 24024 13176
rect 24070 12602 24083 13176
rect 23995 12589 24083 12602
rect 24139 13176 24227 13189
rect 24139 12602 24152 13176
rect 24198 12602 24227 13176
rect 24139 12589 24227 12602
rect 24283 13176 24387 13189
rect 24283 12602 24312 13176
rect 24358 12602 24387 13176
rect 24283 12589 24387 12602
rect 24443 13176 24547 13189
rect 24443 12602 24472 13176
rect 24518 12602 24547 13176
rect 24443 12589 24547 12602
rect 24603 13176 24707 13189
rect 24603 12602 24632 13176
rect 24678 12602 24707 13176
rect 24603 12589 24707 12602
rect 24763 13176 24867 13189
rect 24763 12602 24792 13176
rect 24838 12602 24867 13176
rect 24763 12589 24867 12602
rect 24923 13176 25027 13189
rect 24923 12602 24952 13176
rect 24998 12602 25027 13176
rect 24923 12589 25027 12602
rect 25083 13176 25187 13189
rect 25083 12602 25112 13176
rect 25158 12602 25187 13176
rect 25083 12589 25187 12602
rect 25243 13176 25347 13189
rect 25243 12602 25272 13176
rect 25318 12602 25347 13176
rect 25243 12589 25347 12602
rect 25403 13176 25491 13189
rect 25403 12602 25432 13176
rect 25478 12602 25491 13176
rect 25403 12589 25491 12602
rect 25547 13176 25635 13189
rect 25547 12602 25560 13176
rect 25606 12602 25635 13176
rect 25547 12589 25635 12602
rect 25691 13176 25779 13189
rect 25691 12602 25720 13176
rect 25766 12602 25779 13176
rect 25691 12589 25779 12602
rect 23851 12240 23939 12253
rect 23851 11666 23864 12240
rect 23910 11666 23939 12240
rect 23851 11653 23939 11666
rect 23995 12240 24083 12253
rect 23995 11666 24024 12240
rect 24070 11666 24083 12240
rect 23995 11653 24083 11666
rect 24139 12240 24227 12253
rect 24139 11666 24152 12240
rect 24198 11666 24227 12240
rect 24139 11653 24227 11666
rect 24283 12240 24387 12253
rect 24283 11666 24312 12240
rect 24358 11666 24387 12240
rect 24283 11653 24387 11666
rect 24443 12240 24547 12253
rect 24443 11666 24472 12240
rect 24518 11666 24547 12240
rect 24443 11653 24547 11666
rect 24603 12240 24707 12253
rect 24603 11666 24632 12240
rect 24678 11666 24707 12240
rect 24603 11653 24707 11666
rect 24763 12240 24867 12253
rect 24763 11666 24792 12240
rect 24838 11666 24867 12240
rect 24763 11653 24867 11666
rect 24923 12240 25027 12253
rect 24923 11666 24952 12240
rect 24998 11666 25027 12240
rect 24923 11653 25027 11666
rect 25083 12240 25187 12253
rect 25083 11666 25112 12240
rect 25158 11666 25187 12240
rect 25083 11653 25187 11666
rect 25243 12240 25347 12253
rect 25243 11666 25272 12240
rect 25318 11666 25347 12240
rect 25243 11653 25347 11666
rect 25403 12240 25491 12253
rect 25403 11666 25432 12240
rect 25478 11666 25491 12240
rect 25403 11653 25491 11666
rect 25547 12240 25635 12253
rect 25547 11666 25560 12240
rect 25606 11666 25635 12240
rect 25547 11653 25635 11666
rect 25691 12240 25779 12253
rect 25691 11666 25720 12240
rect 25766 11666 25779 12240
rect 25691 11653 25779 11666
rect 23851 11304 23939 11317
rect 23851 10730 23864 11304
rect 23910 10730 23939 11304
rect 23851 10717 23939 10730
rect 23995 11304 24083 11317
rect 23995 10730 24024 11304
rect 24070 10730 24083 11304
rect 23995 10717 24083 10730
rect 24139 11304 24227 11317
rect 24139 10730 24152 11304
rect 24198 10730 24227 11304
rect 24139 10717 24227 10730
rect 24283 11304 24387 11317
rect 24283 10730 24312 11304
rect 24358 10730 24387 11304
rect 24283 10717 24387 10730
rect 24443 11304 24547 11317
rect 24443 10730 24472 11304
rect 24518 10730 24547 11304
rect 24443 10717 24547 10730
rect 24603 11304 24707 11317
rect 24603 10730 24632 11304
rect 24678 10730 24707 11304
rect 24603 10717 24707 10730
rect 24763 11304 24867 11317
rect 24763 10730 24792 11304
rect 24838 10730 24867 11304
rect 24763 10717 24867 10730
rect 24923 11304 25027 11317
rect 24923 10730 24952 11304
rect 24998 10730 25027 11304
rect 24923 10717 25027 10730
rect 25083 11304 25187 11317
rect 25083 10730 25112 11304
rect 25158 10730 25187 11304
rect 25083 10717 25187 10730
rect 25243 11304 25347 11317
rect 25243 10730 25272 11304
rect 25318 10730 25347 11304
rect 25243 10717 25347 10730
rect 25403 11304 25491 11317
rect 25403 10730 25432 11304
rect 25478 10730 25491 11304
rect 25403 10717 25491 10730
rect 25547 11304 25635 11317
rect 25547 10730 25560 11304
rect 25606 10730 25635 11304
rect 25547 10717 25635 10730
rect 25691 11304 25779 11317
rect 25691 10730 25720 11304
rect 25766 10730 25779 11304
rect 25691 10717 25779 10730
rect 23851 10368 23939 10381
rect 23851 9794 23864 10368
rect 23910 9794 23939 10368
rect 23851 9781 23939 9794
rect 23995 10368 24083 10381
rect 23995 9794 24024 10368
rect 24070 9794 24083 10368
rect 23995 9781 24083 9794
rect 24139 10368 24227 10381
rect 24139 9794 24152 10368
rect 24198 9794 24227 10368
rect 24139 9781 24227 9794
rect 24283 10368 24387 10381
rect 24283 9794 24312 10368
rect 24358 9794 24387 10368
rect 24283 9781 24387 9794
rect 24443 10368 24547 10381
rect 24443 9794 24472 10368
rect 24518 9794 24547 10368
rect 24443 9781 24547 9794
rect 24603 10368 24707 10381
rect 24603 9794 24632 10368
rect 24678 9794 24707 10368
rect 24603 9781 24707 9794
rect 24763 10368 24867 10381
rect 24763 9794 24792 10368
rect 24838 9794 24867 10368
rect 24763 9781 24867 9794
rect 24923 10368 25027 10381
rect 24923 9794 24952 10368
rect 24998 9794 25027 10368
rect 24923 9781 25027 9794
rect 25083 10368 25187 10381
rect 25083 9794 25112 10368
rect 25158 9794 25187 10368
rect 25083 9781 25187 9794
rect 25243 10368 25347 10381
rect 25243 9794 25272 10368
rect 25318 9794 25347 10368
rect 25243 9781 25347 9794
rect 25403 10368 25491 10381
rect 25403 9794 25432 10368
rect 25478 9794 25491 10368
rect 25403 9781 25491 9794
rect 25547 10368 25635 10381
rect 25547 9794 25560 10368
rect 25606 9794 25635 10368
rect 25547 9781 25635 9794
rect 25691 10368 25779 10381
rect 25691 9794 25720 10368
rect 25766 9794 25779 10368
rect 25691 9781 25779 9794
rect 23851 9432 23939 9445
rect 23851 8858 23864 9432
rect 23910 8858 23939 9432
rect 23851 8845 23939 8858
rect 23995 9432 24083 9445
rect 23995 8858 24024 9432
rect 24070 8858 24083 9432
rect 23995 8845 24083 8858
rect 24139 9432 24227 9445
rect 24139 8858 24152 9432
rect 24198 8858 24227 9432
rect 24139 8845 24227 8858
rect 24283 9432 24387 9445
rect 24283 8858 24312 9432
rect 24358 8858 24387 9432
rect 24283 8845 24387 8858
rect 24443 9432 24547 9445
rect 24443 8858 24472 9432
rect 24518 8858 24547 9432
rect 24443 8845 24547 8858
rect 24603 9432 24707 9445
rect 24603 8858 24632 9432
rect 24678 8858 24707 9432
rect 24603 8845 24707 8858
rect 24763 9432 24867 9445
rect 24763 8858 24792 9432
rect 24838 8858 24867 9432
rect 24763 8845 24867 8858
rect 24923 9432 25027 9445
rect 24923 8858 24952 9432
rect 24998 8858 25027 9432
rect 24923 8845 25027 8858
rect 25083 9432 25187 9445
rect 25083 8858 25112 9432
rect 25158 8858 25187 9432
rect 25083 8845 25187 8858
rect 25243 9432 25347 9445
rect 25243 8858 25272 9432
rect 25318 8858 25347 9432
rect 25243 8845 25347 8858
rect 25403 9432 25491 9445
rect 25403 8858 25432 9432
rect 25478 8858 25491 9432
rect 25403 8845 25491 8858
rect 25547 9432 25635 9445
rect 25547 8858 25560 9432
rect 25606 8858 25635 9432
rect 25547 8845 25635 8858
rect 25691 9432 25779 9445
rect 25691 8858 25720 9432
rect 25766 8858 25779 9432
rect 25691 8845 25779 8858
rect 23851 8496 23939 8509
rect 23851 7922 23864 8496
rect 23910 7922 23939 8496
rect 23851 7909 23939 7922
rect 23995 8496 24083 8509
rect 23995 7922 24024 8496
rect 24070 7922 24083 8496
rect 23995 7909 24083 7922
rect 24139 8496 24227 8509
rect 24139 7922 24152 8496
rect 24198 7922 24227 8496
rect 24139 7909 24227 7922
rect 24283 8496 24387 8509
rect 24283 7922 24312 8496
rect 24358 7922 24387 8496
rect 24283 7909 24387 7922
rect 24443 8496 24547 8509
rect 24443 7922 24472 8496
rect 24518 7922 24547 8496
rect 24443 7909 24547 7922
rect 24603 8496 24707 8509
rect 24603 7922 24632 8496
rect 24678 7922 24707 8496
rect 24603 7909 24707 7922
rect 24763 8496 24867 8509
rect 24763 7922 24792 8496
rect 24838 7922 24867 8496
rect 24763 7909 24867 7922
rect 24923 8496 25027 8509
rect 24923 7922 24952 8496
rect 24998 7922 25027 8496
rect 24923 7909 25027 7922
rect 25083 8496 25187 8509
rect 25083 7922 25112 8496
rect 25158 7922 25187 8496
rect 25083 7909 25187 7922
rect 25243 8496 25347 8509
rect 25243 7922 25272 8496
rect 25318 7922 25347 8496
rect 25243 7909 25347 7922
rect 25403 8496 25491 8509
rect 25403 7922 25432 8496
rect 25478 7922 25491 8496
rect 25403 7909 25491 7922
rect 25547 8496 25635 8509
rect 25547 7922 25560 8496
rect 25606 7922 25635 8496
rect 25547 7909 25635 7922
rect 25691 8496 25779 8509
rect 25691 7922 25720 8496
rect 25766 7922 25779 8496
rect 25691 7909 25779 7922
rect 27820 13176 27908 13189
rect 27820 12602 27833 13176
rect 27879 12602 27908 13176
rect 27820 12589 27908 12602
rect 27964 13176 28052 13189
rect 27964 12602 27993 13176
rect 28039 12602 28052 13176
rect 27964 12589 28052 12602
rect 28108 13176 28196 13189
rect 28108 12602 28121 13176
rect 28167 12602 28196 13176
rect 28108 12589 28196 12602
rect 28252 13176 28356 13189
rect 28252 12602 28281 13176
rect 28327 12602 28356 13176
rect 28252 12589 28356 12602
rect 28412 13176 28516 13189
rect 28412 12602 28441 13176
rect 28487 12602 28516 13176
rect 28412 12589 28516 12602
rect 28572 13176 28676 13189
rect 28572 12602 28601 13176
rect 28647 12602 28676 13176
rect 28572 12589 28676 12602
rect 28732 13176 28836 13189
rect 28732 12602 28761 13176
rect 28807 12602 28836 13176
rect 28732 12589 28836 12602
rect 28892 13176 28996 13189
rect 28892 12602 28921 13176
rect 28967 12602 28996 13176
rect 28892 12589 28996 12602
rect 29052 13176 29156 13189
rect 29052 12602 29081 13176
rect 29127 12602 29156 13176
rect 29052 12589 29156 12602
rect 29212 13176 29316 13189
rect 29212 12602 29241 13176
rect 29287 12602 29316 13176
rect 29212 12589 29316 12602
rect 29372 13176 29460 13189
rect 29372 12602 29401 13176
rect 29447 12602 29460 13176
rect 29372 12589 29460 12602
rect 29516 13176 29604 13189
rect 29516 12602 29529 13176
rect 29575 12602 29604 13176
rect 29516 12589 29604 12602
rect 29660 13176 29748 13189
rect 29660 12602 29689 13176
rect 29735 12602 29748 13176
rect 29660 12589 29748 12602
rect 27820 12240 27908 12253
rect 27820 11666 27833 12240
rect 27879 11666 27908 12240
rect 27820 11653 27908 11666
rect 27964 12240 28052 12253
rect 27964 11666 27993 12240
rect 28039 11666 28052 12240
rect 27964 11653 28052 11666
rect 28108 12240 28196 12253
rect 28108 11666 28121 12240
rect 28167 11666 28196 12240
rect 28108 11653 28196 11666
rect 28252 12240 28356 12253
rect 28252 11666 28281 12240
rect 28327 11666 28356 12240
rect 28252 11653 28356 11666
rect 28412 12240 28516 12253
rect 28412 11666 28441 12240
rect 28487 11666 28516 12240
rect 28412 11653 28516 11666
rect 28572 12240 28676 12253
rect 28572 11666 28601 12240
rect 28647 11666 28676 12240
rect 28572 11653 28676 11666
rect 28732 12240 28836 12253
rect 28732 11666 28761 12240
rect 28807 11666 28836 12240
rect 28732 11653 28836 11666
rect 28892 12240 28996 12253
rect 28892 11666 28921 12240
rect 28967 11666 28996 12240
rect 28892 11653 28996 11666
rect 29052 12240 29156 12253
rect 29052 11666 29081 12240
rect 29127 11666 29156 12240
rect 29052 11653 29156 11666
rect 29212 12240 29316 12253
rect 29212 11666 29241 12240
rect 29287 11666 29316 12240
rect 29212 11653 29316 11666
rect 29372 12240 29460 12253
rect 29372 11666 29401 12240
rect 29447 11666 29460 12240
rect 29372 11653 29460 11666
rect 29516 12240 29604 12253
rect 29516 11666 29529 12240
rect 29575 11666 29604 12240
rect 29516 11653 29604 11666
rect 29660 12240 29748 12253
rect 29660 11666 29689 12240
rect 29735 11666 29748 12240
rect 29660 11653 29748 11666
rect 27820 11304 27908 11317
rect 27820 10730 27833 11304
rect 27879 10730 27908 11304
rect 27820 10717 27908 10730
rect 27964 11304 28052 11317
rect 27964 10730 27993 11304
rect 28039 10730 28052 11304
rect 27964 10717 28052 10730
rect 28108 11304 28196 11317
rect 28108 10730 28121 11304
rect 28167 10730 28196 11304
rect 28108 10717 28196 10730
rect 28252 11304 28356 11317
rect 28252 10730 28281 11304
rect 28327 10730 28356 11304
rect 28252 10717 28356 10730
rect 28412 11304 28516 11317
rect 28412 10730 28441 11304
rect 28487 10730 28516 11304
rect 28412 10717 28516 10730
rect 28572 11304 28676 11317
rect 28572 10730 28601 11304
rect 28647 10730 28676 11304
rect 28572 10717 28676 10730
rect 28732 11304 28836 11317
rect 28732 10730 28761 11304
rect 28807 10730 28836 11304
rect 28732 10717 28836 10730
rect 28892 11304 28996 11317
rect 28892 10730 28921 11304
rect 28967 10730 28996 11304
rect 28892 10717 28996 10730
rect 29052 11304 29156 11317
rect 29052 10730 29081 11304
rect 29127 10730 29156 11304
rect 29052 10717 29156 10730
rect 29212 11304 29316 11317
rect 29212 10730 29241 11304
rect 29287 10730 29316 11304
rect 29212 10717 29316 10730
rect 29372 11304 29460 11317
rect 29372 10730 29401 11304
rect 29447 10730 29460 11304
rect 29372 10717 29460 10730
rect 29516 11304 29604 11317
rect 29516 10730 29529 11304
rect 29575 10730 29604 11304
rect 29516 10717 29604 10730
rect 29660 11304 29748 11317
rect 29660 10730 29689 11304
rect 29735 10730 29748 11304
rect 29660 10717 29748 10730
rect 27820 10368 27908 10381
rect 27820 9794 27833 10368
rect 27879 9794 27908 10368
rect 27820 9781 27908 9794
rect 27964 10368 28052 10381
rect 27964 9794 27993 10368
rect 28039 9794 28052 10368
rect 27964 9781 28052 9794
rect 28108 10368 28196 10381
rect 28108 9794 28121 10368
rect 28167 9794 28196 10368
rect 28108 9781 28196 9794
rect 28252 10368 28356 10381
rect 28252 9794 28281 10368
rect 28327 9794 28356 10368
rect 28252 9781 28356 9794
rect 28412 10368 28516 10381
rect 28412 9794 28441 10368
rect 28487 9794 28516 10368
rect 28412 9781 28516 9794
rect 28572 10368 28676 10381
rect 28572 9794 28601 10368
rect 28647 9794 28676 10368
rect 28572 9781 28676 9794
rect 28732 10368 28836 10381
rect 28732 9794 28761 10368
rect 28807 9794 28836 10368
rect 28732 9781 28836 9794
rect 28892 10368 28996 10381
rect 28892 9794 28921 10368
rect 28967 9794 28996 10368
rect 28892 9781 28996 9794
rect 29052 10368 29156 10381
rect 29052 9794 29081 10368
rect 29127 9794 29156 10368
rect 29052 9781 29156 9794
rect 29212 10368 29316 10381
rect 29212 9794 29241 10368
rect 29287 9794 29316 10368
rect 29212 9781 29316 9794
rect 29372 10368 29460 10381
rect 29372 9794 29401 10368
rect 29447 9794 29460 10368
rect 29372 9781 29460 9794
rect 29516 10368 29604 10381
rect 29516 9794 29529 10368
rect 29575 9794 29604 10368
rect 29516 9781 29604 9794
rect 29660 10368 29748 10381
rect 29660 9794 29689 10368
rect 29735 9794 29748 10368
rect 29660 9781 29748 9794
rect 27820 9432 27908 9445
rect 27820 8858 27833 9432
rect 27879 8858 27908 9432
rect 27820 8845 27908 8858
rect 27964 9432 28052 9445
rect 27964 8858 27993 9432
rect 28039 8858 28052 9432
rect 27964 8845 28052 8858
rect 28108 9432 28196 9445
rect 28108 8858 28121 9432
rect 28167 8858 28196 9432
rect 28108 8845 28196 8858
rect 28252 9432 28356 9445
rect 28252 8858 28281 9432
rect 28327 8858 28356 9432
rect 28252 8845 28356 8858
rect 28412 9432 28516 9445
rect 28412 8858 28441 9432
rect 28487 8858 28516 9432
rect 28412 8845 28516 8858
rect 28572 9432 28676 9445
rect 28572 8858 28601 9432
rect 28647 8858 28676 9432
rect 28572 8845 28676 8858
rect 28732 9432 28836 9445
rect 28732 8858 28761 9432
rect 28807 8858 28836 9432
rect 28732 8845 28836 8858
rect 28892 9432 28996 9445
rect 28892 8858 28921 9432
rect 28967 8858 28996 9432
rect 28892 8845 28996 8858
rect 29052 9432 29156 9445
rect 29052 8858 29081 9432
rect 29127 8858 29156 9432
rect 29052 8845 29156 8858
rect 29212 9432 29316 9445
rect 29212 8858 29241 9432
rect 29287 8858 29316 9432
rect 29212 8845 29316 8858
rect 29372 9432 29460 9445
rect 29372 8858 29401 9432
rect 29447 8858 29460 9432
rect 29372 8845 29460 8858
rect 29516 9432 29604 9445
rect 29516 8858 29529 9432
rect 29575 8858 29604 9432
rect 29516 8845 29604 8858
rect 29660 9432 29748 9445
rect 29660 8858 29689 9432
rect 29735 8858 29748 9432
rect 29660 8845 29748 8858
rect 27820 8496 27908 8509
rect 27820 7922 27833 8496
rect 27879 7922 27908 8496
rect 27820 7909 27908 7922
rect 27964 8496 28052 8509
rect 27964 7922 27993 8496
rect 28039 7922 28052 8496
rect 27964 7909 28052 7922
rect 28108 8496 28196 8509
rect 28108 7922 28121 8496
rect 28167 7922 28196 8496
rect 28108 7909 28196 7922
rect 28252 8496 28356 8509
rect 28252 7922 28281 8496
rect 28327 7922 28356 8496
rect 28252 7909 28356 7922
rect 28412 8496 28516 8509
rect 28412 7922 28441 8496
rect 28487 7922 28516 8496
rect 28412 7909 28516 7922
rect 28572 8496 28676 8509
rect 28572 7922 28601 8496
rect 28647 7922 28676 8496
rect 28572 7909 28676 7922
rect 28732 8496 28836 8509
rect 28732 7922 28761 8496
rect 28807 7922 28836 8496
rect 28732 7909 28836 7922
rect 28892 8496 28996 8509
rect 28892 7922 28921 8496
rect 28967 7922 28996 8496
rect 28892 7909 28996 7922
rect 29052 8496 29156 8509
rect 29052 7922 29081 8496
rect 29127 7922 29156 8496
rect 29052 7909 29156 7922
rect 29212 8496 29316 8509
rect 29212 7922 29241 8496
rect 29287 7922 29316 8496
rect 29212 7909 29316 7922
rect 29372 8496 29460 8509
rect 29372 7922 29401 8496
rect 29447 7922 29460 8496
rect 29372 7909 29460 7922
rect 29516 8496 29604 8509
rect 29516 7922 29529 8496
rect 29575 7922 29604 8496
rect 29516 7909 29604 7922
rect 29660 8496 29748 8509
rect 29660 7922 29689 8496
rect 29735 7922 29748 8496
rect 29660 7909 29748 7922
rect 7383 5725 7471 5738
rect 7383 5551 7396 5725
rect 7442 5551 7471 5725
rect 7383 5538 7471 5551
rect 7527 5725 7615 5738
rect 7527 5551 7556 5725
rect 7602 5551 7615 5725
rect 7527 5538 7615 5551
rect 7671 5725 7759 5738
rect 7671 5551 7684 5725
rect 7730 5551 7759 5725
rect 7671 5538 7759 5551
rect 7815 5725 7919 5738
rect 7815 5551 7844 5725
rect 7890 5551 7919 5725
rect 7815 5538 7919 5551
rect 7975 5725 8079 5738
rect 7975 5551 8004 5725
rect 8050 5551 8079 5725
rect 7975 5538 8079 5551
rect 8135 5725 8239 5738
rect 8135 5551 8164 5725
rect 8210 5551 8239 5725
rect 8135 5538 8239 5551
rect 8295 5725 8399 5738
rect 8295 5551 8324 5725
rect 8370 5551 8399 5725
rect 8295 5538 8399 5551
rect 8455 5725 8559 5738
rect 8455 5551 8484 5725
rect 8530 5551 8559 5725
rect 8455 5538 8559 5551
rect 8615 5725 8719 5738
rect 8615 5551 8644 5725
rect 8690 5551 8719 5725
rect 8615 5538 8719 5551
rect 8775 5725 8879 5738
rect 8775 5551 8804 5725
rect 8850 5551 8879 5725
rect 8775 5538 8879 5551
rect 8935 5725 9039 5738
rect 8935 5551 8964 5725
rect 9010 5551 9039 5725
rect 8935 5538 9039 5551
rect 9095 5725 9199 5738
rect 9095 5551 9124 5725
rect 9170 5551 9199 5725
rect 9095 5538 9199 5551
rect 9255 5725 9343 5738
rect 9255 5551 9284 5725
rect 9330 5551 9343 5725
rect 9255 5538 9343 5551
rect 9399 5725 9487 5738
rect 9399 5551 9412 5725
rect 9458 5551 9487 5725
rect 9399 5538 9487 5551
rect 9543 5725 9631 5738
rect 9543 5551 9572 5725
rect 9618 5551 9631 5725
rect 9543 5538 9631 5551
rect 7383 5189 7471 5202
rect 7383 5015 7396 5189
rect 7442 5015 7471 5189
rect 7383 5002 7471 5015
rect 7527 5189 7615 5202
rect 7527 5015 7556 5189
rect 7602 5015 7615 5189
rect 7527 5002 7615 5015
rect 7671 5189 7759 5202
rect 7671 5015 7684 5189
rect 7730 5015 7759 5189
rect 7671 5002 7759 5015
rect 7815 5189 7919 5202
rect 7815 5015 7844 5189
rect 7890 5015 7919 5189
rect 7815 5002 7919 5015
rect 7975 5189 8079 5202
rect 7975 5015 8004 5189
rect 8050 5015 8079 5189
rect 7975 5002 8079 5015
rect 8135 5189 8239 5202
rect 8135 5015 8164 5189
rect 8210 5015 8239 5189
rect 8135 5002 8239 5015
rect 8295 5189 8399 5202
rect 8295 5015 8324 5189
rect 8370 5015 8399 5189
rect 8295 5002 8399 5015
rect 8455 5189 8559 5202
rect 8455 5015 8484 5189
rect 8530 5015 8559 5189
rect 8455 5002 8559 5015
rect 8615 5189 8719 5202
rect 8615 5015 8644 5189
rect 8690 5015 8719 5189
rect 8615 5002 8719 5015
rect 8775 5189 8879 5202
rect 8775 5015 8804 5189
rect 8850 5015 8879 5189
rect 8775 5002 8879 5015
rect 8935 5189 9039 5202
rect 8935 5015 8964 5189
rect 9010 5015 9039 5189
rect 8935 5002 9039 5015
rect 9095 5189 9199 5202
rect 9095 5015 9124 5189
rect 9170 5015 9199 5189
rect 9095 5002 9199 5015
rect 9255 5189 9343 5202
rect 9255 5015 9284 5189
rect 9330 5015 9343 5189
rect 9255 5002 9343 5015
rect 9399 5189 9487 5202
rect 9399 5015 9412 5189
rect 9458 5015 9487 5189
rect 9399 5002 9487 5015
rect 9543 5189 9631 5202
rect 9543 5015 9572 5189
rect 9618 5015 9631 5189
rect 9543 5002 9631 5015
rect 7383 4653 7471 4666
rect 7383 4479 7396 4653
rect 7442 4479 7471 4653
rect 7383 4466 7471 4479
rect 7527 4653 7615 4666
rect 7527 4479 7556 4653
rect 7602 4479 7615 4653
rect 7527 4466 7615 4479
rect 7671 4653 7759 4666
rect 7671 4479 7684 4653
rect 7730 4479 7759 4653
rect 7671 4466 7759 4479
rect 7815 4653 7919 4666
rect 7815 4479 7844 4653
rect 7890 4479 7919 4653
rect 7815 4466 7919 4479
rect 7975 4653 8079 4666
rect 7975 4479 8004 4653
rect 8050 4479 8079 4653
rect 7975 4466 8079 4479
rect 8135 4653 8239 4666
rect 8135 4479 8164 4653
rect 8210 4479 8239 4653
rect 8135 4466 8239 4479
rect 8295 4653 8399 4666
rect 8295 4479 8324 4653
rect 8370 4479 8399 4653
rect 8295 4466 8399 4479
rect 8455 4653 8559 4666
rect 8455 4479 8484 4653
rect 8530 4479 8559 4653
rect 8455 4466 8559 4479
rect 8615 4653 8719 4666
rect 8615 4479 8644 4653
rect 8690 4479 8719 4653
rect 8615 4466 8719 4479
rect 8775 4653 8879 4666
rect 8775 4479 8804 4653
rect 8850 4479 8879 4653
rect 8775 4466 8879 4479
rect 8935 4653 9039 4666
rect 8935 4479 8964 4653
rect 9010 4479 9039 4653
rect 8935 4466 9039 4479
rect 9095 4653 9199 4666
rect 9095 4479 9124 4653
rect 9170 4479 9199 4653
rect 9095 4466 9199 4479
rect 9255 4653 9343 4666
rect 9255 4479 9284 4653
rect 9330 4479 9343 4653
rect 9255 4466 9343 4479
rect 9399 4653 9487 4666
rect 9399 4479 9412 4653
rect 9458 4479 9487 4653
rect 9399 4466 9487 4479
rect 9543 4653 9631 4666
rect 9543 4479 9572 4653
rect 9618 4479 9631 4653
rect 9543 4466 9631 4479
rect 7383 4117 7471 4130
rect 7383 3943 7396 4117
rect 7442 3943 7471 4117
rect 7383 3930 7471 3943
rect 7527 4117 7615 4130
rect 7527 3943 7556 4117
rect 7602 3943 7615 4117
rect 7527 3930 7615 3943
rect 7671 4117 7759 4130
rect 7671 3943 7684 4117
rect 7730 3943 7759 4117
rect 7671 3930 7759 3943
rect 7815 4117 7919 4130
rect 7815 3943 7844 4117
rect 7890 3943 7919 4117
rect 7815 3930 7919 3943
rect 7975 4117 8079 4130
rect 7975 3943 8004 4117
rect 8050 3943 8079 4117
rect 7975 3930 8079 3943
rect 8135 4117 8239 4130
rect 8135 3943 8164 4117
rect 8210 3943 8239 4117
rect 8135 3930 8239 3943
rect 8295 4117 8399 4130
rect 8295 3943 8324 4117
rect 8370 3943 8399 4117
rect 8295 3930 8399 3943
rect 8455 4117 8559 4130
rect 8455 3943 8484 4117
rect 8530 3943 8559 4117
rect 8455 3930 8559 3943
rect 8615 4117 8719 4130
rect 8615 3943 8644 4117
rect 8690 3943 8719 4117
rect 8615 3930 8719 3943
rect 8775 4117 8879 4130
rect 8775 3943 8804 4117
rect 8850 3943 8879 4117
rect 8775 3930 8879 3943
rect 8935 4117 9039 4130
rect 8935 3943 8964 4117
rect 9010 3943 9039 4117
rect 8935 3930 9039 3943
rect 9095 4117 9199 4130
rect 9095 3943 9124 4117
rect 9170 3943 9199 4117
rect 9095 3930 9199 3943
rect 9255 4117 9343 4130
rect 9255 3943 9284 4117
rect 9330 3943 9343 4117
rect 9255 3930 9343 3943
rect 9399 4117 9487 4130
rect 9399 3943 9412 4117
rect 9458 3943 9487 4117
rect 9399 3930 9487 3943
rect 9543 4117 9631 4130
rect 9543 3943 9572 4117
rect 9618 3943 9631 4117
rect 9543 3930 9631 3943
rect 7383 3581 7471 3594
rect 7383 3407 7396 3581
rect 7442 3407 7471 3581
rect 7383 3394 7471 3407
rect 7527 3581 7615 3594
rect 7527 3407 7556 3581
rect 7602 3407 7615 3581
rect 7527 3394 7615 3407
rect 7671 3581 7759 3594
rect 7671 3407 7684 3581
rect 7730 3407 7759 3581
rect 7671 3394 7759 3407
rect 7815 3581 7919 3594
rect 7815 3407 7844 3581
rect 7890 3407 7919 3581
rect 7815 3394 7919 3407
rect 7975 3581 8079 3594
rect 7975 3407 8004 3581
rect 8050 3407 8079 3581
rect 7975 3394 8079 3407
rect 8135 3581 8239 3594
rect 8135 3407 8164 3581
rect 8210 3407 8239 3581
rect 8135 3394 8239 3407
rect 8295 3581 8399 3594
rect 8295 3407 8324 3581
rect 8370 3407 8399 3581
rect 8295 3394 8399 3407
rect 8455 3581 8559 3594
rect 8455 3407 8484 3581
rect 8530 3407 8559 3581
rect 8455 3394 8559 3407
rect 8615 3581 8719 3594
rect 8615 3407 8644 3581
rect 8690 3407 8719 3581
rect 8615 3394 8719 3407
rect 8775 3581 8879 3594
rect 8775 3407 8804 3581
rect 8850 3407 8879 3581
rect 8775 3394 8879 3407
rect 8935 3581 9039 3594
rect 8935 3407 8964 3581
rect 9010 3407 9039 3581
rect 8935 3394 9039 3407
rect 9095 3581 9199 3594
rect 9095 3407 9124 3581
rect 9170 3407 9199 3581
rect 9095 3394 9199 3407
rect 9255 3581 9343 3594
rect 9255 3407 9284 3581
rect 9330 3407 9343 3581
rect 9255 3394 9343 3407
rect 9399 3581 9487 3594
rect 9399 3407 9412 3581
rect 9458 3407 9487 3581
rect 9399 3394 9487 3407
rect 9543 3581 9631 3594
rect 9543 3407 9572 3581
rect 9618 3407 9631 3581
rect 9543 3394 9631 3407
rect 7383 3045 7471 3058
rect 7383 2871 7396 3045
rect 7442 2871 7471 3045
rect 7383 2858 7471 2871
rect 7527 3045 7615 3058
rect 7527 2871 7556 3045
rect 7602 2871 7615 3045
rect 7527 2858 7615 2871
rect 7671 3045 7759 3058
rect 7671 2871 7684 3045
rect 7730 2871 7759 3045
rect 7671 2858 7759 2871
rect 7815 3045 7919 3058
rect 7815 2871 7844 3045
rect 7890 2871 7919 3045
rect 7815 2858 7919 2871
rect 7975 3045 8079 3058
rect 7975 2871 8004 3045
rect 8050 2871 8079 3045
rect 7975 2858 8079 2871
rect 8135 3045 8239 3058
rect 8135 2871 8164 3045
rect 8210 2871 8239 3045
rect 8135 2858 8239 2871
rect 8295 3045 8399 3058
rect 8295 2871 8324 3045
rect 8370 2871 8399 3045
rect 8295 2858 8399 2871
rect 8455 3045 8559 3058
rect 8455 2871 8484 3045
rect 8530 2871 8559 3045
rect 8455 2858 8559 2871
rect 8615 3045 8719 3058
rect 8615 2871 8644 3045
rect 8690 2871 8719 3045
rect 8615 2858 8719 2871
rect 8775 3045 8879 3058
rect 8775 2871 8804 3045
rect 8850 2871 8879 3045
rect 8775 2858 8879 2871
rect 8935 3045 9039 3058
rect 8935 2871 8964 3045
rect 9010 2871 9039 3045
rect 8935 2858 9039 2871
rect 9095 3045 9199 3058
rect 9095 2871 9124 3045
rect 9170 2871 9199 3045
rect 9095 2858 9199 2871
rect 9255 3045 9343 3058
rect 9255 2871 9284 3045
rect 9330 2871 9343 3045
rect 9255 2858 9343 2871
rect 9399 3045 9487 3058
rect 9399 2871 9412 3045
rect 9458 2871 9487 3045
rect 9399 2858 9487 2871
rect 9543 3045 9631 3058
rect 9543 2871 9572 3045
rect 9618 2871 9631 3045
rect 9543 2858 9631 2871
rect 12670 3768 12758 3781
rect 12670 3394 12683 3768
rect 12729 3394 12758 3768
rect 12670 3381 12758 3394
rect 12958 3768 13046 3781
rect 12958 3394 12987 3768
rect 13033 3394 13046 3768
rect 12958 3381 13046 3394
rect 13102 3768 13190 3781
rect 13102 3394 13115 3768
rect 13161 3394 13190 3768
rect 13102 3381 13190 3394
rect 13390 3768 13494 3781
rect 13390 3394 13419 3768
rect 13465 3394 13494 3768
rect 13390 3381 13494 3394
rect 13694 3768 13798 3781
rect 13694 3394 13723 3768
rect 13769 3394 13798 3768
rect 13694 3381 13798 3394
rect 13998 3768 14102 3781
rect 13998 3394 14027 3768
rect 14073 3394 14102 3768
rect 13998 3381 14102 3394
rect 14302 3768 14406 3781
rect 14302 3394 14331 3768
rect 14377 3394 14406 3768
rect 14302 3381 14406 3394
rect 14606 3768 14710 3781
rect 14606 3394 14635 3768
rect 14681 3394 14710 3768
rect 14606 3381 14710 3394
rect 14910 3768 14998 3781
rect 14910 3394 14939 3768
rect 14985 3394 14998 3768
rect 14910 3381 14998 3394
rect 15054 3768 15142 3781
rect 15054 3394 15067 3768
rect 15113 3394 15142 3768
rect 15054 3381 15142 3394
rect 15342 3768 15446 3781
rect 15342 3394 15371 3768
rect 15417 3394 15446 3768
rect 15342 3381 15446 3394
rect 15646 3768 15750 3781
rect 15646 3394 15675 3768
rect 15721 3394 15750 3768
rect 15646 3381 15750 3394
rect 15950 3768 16054 3781
rect 15950 3394 15979 3768
rect 16025 3394 16054 3768
rect 15950 3381 16054 3394
rect 16254 3768 16358 3781
rect 16254 3394 16283 3768
rect 16329 3394 16358 3768
rect 16254 3381 16358 3394
rect 16558 3768 16662 3781
rect 16558 3394 16587 3768
rect 16633 3394 16662 3768
rect 16558 3381 16662 3394
rect 16862 3768 16950 3781
rect 16862 3394 16891 3768
rect 16937 3394 16950 3768
rect 16862 3381 16950 3394
rect 6136 2416 6224 2429
rect 6136 2242 6149 2416
rect 6195 2242 6224 2416
rect 6136 2229 6224 2242
rect 6280 2416 6368 2429
rect 6280 2242 6309 2416
rect 6355 2242 6368 2416
rect 6280 2229 6368 2242
rect 6424 2416 6512 2429
rect 6424 2242 6437 2416
rect 6483 2242 6512 2416
rect 6424 2229 6512 2242
rect 6568 2416 6672 2429
rect 6568 2242 6597 2416
rect 6643 2242 6672 2416
rect 6568 2229 6672 2242
rect 6728 2416 6832 2429
rect 6728 2242 6757 2416
rect 6803 2242 6832 2416
rect 6728 2229 6832 2242
rect 6888 2416 6992 2429
rect 6888 2242 6917 2416
rect 6963 2242 6992 2416
rect 6888 2229 6992 2242
rect 7048 2416 7152 2429
rect 7048 2242 7077 2416
rect 7123 2242 7152 2416
rect 7048 2229 7152 2242
rect 7208 2416 7312 2429
rect 7208 2242 7237 2416
rect 7283 2242 7312 2416
rect 7208 2229 7312 2242
rect 7368 2416 7472 2429
rect 7368 2242 7397 2416
rect 7443 2242 7472 2416
rect 7368 2229 7472 2242
rect 7528 2416 7632 2429
rect 7528 2242 7557 2416
rect 7603 2242 7632 2416
rect 7528 2229 7632 2242
rect 7688 2416 7792 2429
rect 7688 2242 7717 2416
rect 7763 2242 7792 2416
rect 7688 2229 7792 2242
rect 7848 2416 7952 2429
rect 7848 2242 7877 2416
rect 7923 2242 7952 2416
rect 7848 2229 7952 2242
rect 8008 2416 8112 2429
rect 8008 2242 8037 2416
rect 8083 2242 8112 2416
rect 8008 2229 8112 2242
rect 8168 2416 8272 2429
rect 8168 2242 8197 2416
rect 8243 2242 8272 2416
rect 8168 2229 8272 2242
rect 8328 2416 8432 2429
rect 8328 2242 8357 2416
rect 8403 2242 8432 2416
rect 8328 2229 8432 2242
rect 8488 2416 8592 2429
rect 8488 2242 8517 2416
rect 8563 2242 8592 2416
rect 8488 2229 8592 2242
rect 8648 2416 8752 2429
rect 8648 2242 8677 2416
rect 8723 2242 8752 2416
rect 8648 2229 8752 2242
rect 8808 2416 8912 2429
rect 8808 2242 8837 2416
rect 8883 2242 8912 2416
rect 8808 2229 8912 2242
rect 8968 2416 9072 2429
rect 8968 2242 8997 2416
rect 9043 2242 9072 2416
rect 8968 2229 9072 2242
rect 9128 2416 9232 2429
rect 9128 2242 9157 2416
rect 9203 2242 9232 2416
rect 9128 2229 9232 2242
rect 9288 2416 9376 2429
rect 9288 2242 9317 2416
rect 9363 2242 9376 2416
rect 9288 2229 9376 2242
rect 9432 2416 9520 2429
rect 9432 2242 9445 2416
rect 9491 2242 9520 2416
rect 9432 2229 9520 2242
rect 9720 2416 9824 2429
rect 9720 2242 9749 2416
rect 9795 2242 9824 2416
rect 9720 2229 9824 2242
rect 10024 2416 10128 2429
rect 10024 2242 10053 2416
rect 10099 2242 10128 2416
rect 10024 2229 10128 2242
rect 10328 2416 10432 2429
rect 10328 2242 10357 2416
rect 10403 2242 10432 2416
rect 10328 2229 10432 2242
rect 10632 2416 10736 2429
rect 10632 2242 10661 2416
rect 10707 2242 10736 2416
rect 10632 2229 10736 2242
rect 10792 2416 10880 2429
rect 10792 2242 10821 2416
rect 10867 2242 10880 2416
rect 10792 2229 10880 2242
rect 6136 1779 6224 1792
rect 6136 1605 6149 1779
rect 6195 1605 6224 1779
rect 6136 1592 6224 1605
rect 6280 1779 6368 1792
rect 6280 1605 6309 1779
rect 6355 1605 6368 1779
rect 6280 1592 6368 1605
rect 6424 1779 6512 1792
rect 6424 1605 6437 1779
rect 6483 1605 6512 1779
rect 6424 1592 6512 1605
rect 6624 1779 6728 1792
rect 6624 1605 6653 1779
rect 6699 1605 6728 1779
rect 6624 1592 6728 1605
rect 6840 1779 6944 1792
rect 6840 1605 6869 1779
rect 6915 1605 6944 1779
rect 6840 1592 6944 1605
rect 7056 1779 7160 1792
rect 7056 1605 7085 1779
rect 7131 1605 7160 1779
rect 7056 1592 7160 1605
rect 7272 1779 7376 1792
rect 7272 1605 7301 1779
rect 7347 1605 7376 1779
rect 7272 1592 7376 1605
rect 7488 1779 7592 1792
rect 7488 1605 7517 1779
rect 7563 1605 7592 1779
rect 7488 1592 7592 1605
rect 7704 1779 7808 1792
rect 7704 1605 7733 1779
rect 7779 1605 7808 1779
rect 7704 1592 7808 1605
rect 7920 1779 8024 1792
rect 7920 1605 7949 1779
rect 7995 1605 8024 1779
rect 7920 1592 8024 1605
rect 8136 1779 8240 1792
rect 8136 1605 8165 1779
rect 8211 1605 8240 1779
rect 8136 1592 8240 1605
rect 8352 1779 8456 1792
rect 8352 1605 8381 1779
rect 8427 1605 8456 1779
rect 8352 1592 8456 1605
rect 8568 1779 8672 1792
rect 8568 1605 8597 1779
rect 8643 1605 8672 1779
rect 8568 1592 8672 1605
rect 8728 1779 8832 1792
rect 8728 1605 8757 1779
rect 8803 1605 8832 1779
rect 8728 1592 8832 1605
rect 8888 1779 8992 1792
rect 8888 1605 8917 1779
rect 8963 1605 8992 1779
rect 8888 1592 8992 1605
rect 9048 1779 9152 1792
rect 9048 1605 9077 1779
rect 9123 1605 9152 1779
rect 9048 1592 9152 1605
rect 9208 1779 9312 1792
rect 9208 1605 9237 1779
rect 9283 1605 9312 1779
rect 9208 1592 9312 1605
rect 9368 1779 9472 1792
rect 9368 1605 9397 1779
rect 9443 1605 9472 1779
rect 9368 1592 9472 1605
rect 9528 1779 9632 1792
rect 9528 1605 9557 1779
rect 9603 1605 9632 1779
rect 9528 1592 9632 1605
rect 9688 1779 9776 1792
rect 9688 1605 9717 1779
rect 9763 1605 9776 1779
rect 9688 1592 9776 1605
rect 9848 1779 9936 1792
rect 9848 1605 9861 1779
rect 9907 1605 9936 1779
rect 9848 1592 9936 1605
rect 9992 1779 10096 1792
rect 9992 1605 10021 1779
rect 10067 1605 10096 1779
rect 9992 1592 10096 1605
rect 10152 1779 10256 1792
rect 10152 1605 10181 1779
rect 10227 1605 10256 1779
rect 10152 1592 10256 1605
rect 10312 1779 10416 1792
rect 10312 1605 10341 1779
rect 10387 1605 10416 1779
rect 10312 1592 10416 1605
rect 10472 1779 10576 1792
rect 10472 1605 10501 1779
rect 10547 1605 10576 1779
rect 10472 1592 10576 1605
rect 10632 1779 10736 1792
rect 10632 1605 10661 1779
rect 10707 1605 10736 1779
rect 10632 1592 10736 1605
rect 10792 1779 10880 1792
rect 10792 1605 10821 1779
rect 10867 1605 10880 1779
rect 10792 1592 10880 1605
rect 12670 3232 12758 3245
rect 12670 2858 12683 3232
rect 12729 2858 12758 3232
rect 12670 2845 12758 2858
rect 12958 3232 13046 3245
rect 12958 2858 12987 3232
rect 13033 2858 13046 3232
rect 12958 2845 13046 2858
rect 13102 3232 13190 3245
rect 13102 2858 13115 3232
rect 13161 2858 13190 3232
rect 13102 2845 13190 2858
rect 13390 3232 13494 3245
rect 13390 2858 13419 3232
rect 13465 2858 13494 3232
rect 13390 2845 13494 2858
rect 13694 3232 13798 3245
rect 13694 2858 13723 3232
rect 13769 2858 13798 3232
rect 13694 2845 13798 2858
rect 13998 3232 14102 3245
rect 13998 2858 14027 3232
rect 14073 2858 14102 3232
rect 13998 2845 14102 2858
rect 14302 3232 14406 3245
rect 14302 2858 14331 3232
rect 14377 2858 14406 3232
rect 14302 2845 14406 2858
rect 14606 3232 14710 3245
rect 14606 2858 14635 3232
rect 14681 2858 14710 3232
rect 14606 2845 14710 2858
rect 14910 3232 14998 3245
rect 14910 2858 14939 3232
rect 14985 2858 14998 3232
rect 14910 2845 14998 2858
rect 15054 3232 15142 3245
rect 15054 2858 15067 3232
rect 15113 2858 15142 3232
rect 15054 2845 15142 2858
rect 15342 3232 15446 3245
rect 15342 2858 15371 3232
rect 15417 2858 15446 3232
rect 15342 2845 15446 2858
rect 15646 3232 15750 3245
rect 15646 2858 15675 3232
rect 15721 2858 15750 3232
rect 15646 2845 15750 2858
rect 15950 3232 16054 3245
rect 15950 2858 15979 3232
rect 16025 2858 16054 3232
rect 15950 2845 16054 2858
rect 16254 3232 16358 3245
rect 16254 2858 16283 3232
rect 16329 2858 16358 3232
rect 16254 2845 16358 2858
rect 16558 3232 16662 3245
rect 16558 2858 16587 3232
rect 16633 2858 16662 3232
rect 16558 2845 16662 2858
rect 16862 3232 16950 3245
rect 16862 2858 16891 3232
rect 16937 2858 16950 3232
rect 16862 2845 16950 2858
rect 12670 2396 12758 2409
rect 12670 2022 12683 2396
rect 12729 2022 12758 2396
rect 12670 2009 12758 2022
rect 12958 2396 13046 2409
rect 12958 2022 12987 2396
rect 13033 2022 13046 2396
rect 12958 2009 13046 2022
rect 13102 2396 13190 2409
rect 13102 2022 13115 2396
rect 13161 2022 13190 2396
rect 13102 2009 13190 2022
rect 13390 2396 13494 2409
rect 13390 2022 13419 2396
rect 13465 2022 13494 2396
rect 13390 2009 13494 2022
rect 13694 2396 13798 2409
rect 13694 2022 13723 2396
rect 13769 2022 13798 2396
rect 13694 2009 13798 2022
rect 13998 2396 14102 2409
rect 13998 2022 14027 2396
rect 14073 2022 14102 2396
rect 13998 2009 14102 2022
rect 14302 2396 14406 2409
rect 14302 2022 14331 2396
rect 14377 2022 14406 2396
rect 14302 2009 14406 2022
rect 14606 2396 14710 2409
rect 14606 2022 14635 2396
rect 14681 2022 14710 2396
rect 14606 2009 14710 2022
rect 14910 2396 14998 2409
rect 14910 2022 14939 2396
rect 14985 2022 14998 2396
rect 14910 2009 14998 2022
rect 15054 2396 15142 2409
rect 15054 2022 15067 2396
rect 15113 2022 15142 2396
rect 15054 2009 15142 2022
rect 15342 2396 15446 2409
rect 15342 2022 15371 2396
rect 15417 2022 15446 2396
rect 15342 2009 15446 2022
rect 15646 2396 15750 2409
rect 15646 2022 15675 2396
rect 15721 2022 15750 2396
rect 15646 2009 15750 2022
rect 15950 2396 16054 2409
rect 15950 2022 15979 2396
rect 16025 2022 16054 2396
rect 15950 2009 16054 2022
rect 16254 2396 16358 2409
rect 16254 2022 16283 2396
rect 16329 2022 16358 2396
rect 16254 2009 16358 2022
rect 16558 2396 16662 2409
rect 16558 2022 16587 2396
rect 16633 2022 16662 2396
rect 16558 2009 16662 2022
rect 16862 2396 16950 2409
rect 16862 2022 16891 2396
rect 16937 2022 16950 2396
rect 16862 2009 16950 2022
<< pdiff >>
rect 3584 14013 3672 14026
rect 3584 13289 3597 14013
rect 3643 13289 3672 14013
rect 3584 13276 3672 13289
rect 3728 14013 3816 14026
rect 3728 13289 3757 14013
rect 3803 13289 3816 14013
rect 3728 13276 3816 13289
rect 3872 14013 3960 14026
rect 3872 13289 3885 14013
rect 3931 13289 3960 14013
rect 3872 13276 3960 13289
rect 4016 14013 4120 14026
rect 4016 13289 4045 14013
rect 4091 13289 4120 14013
rect 4016 13276 4120 13289
rect 4176 14013 4280 14026
rect 4176 13289 4205 14013
rect 4251 13289 4280 14013
rect 4176 13276 4280 13289
rect 4336 14013 4440 14026
rect 4336 13289 4365 14013
rect 4411 13289 4440 14013
rect 4336 13276 4440 13289
rect 4496 14013 4600 14026
rect 4496 13289 4525 14013
rect 4571 13289 4600 14013
rect 4496 13276 4600 13289
rect 4656 14013 4760 14026
rect 4656 13289 4685 14013
rect 4731 13289 4760 14013
rect 4656 13276 4760 13289
rect 4816 14013 4920 14026
rect 4816 13289 4845 14013
rect 4891 13289 4920 14013
rect 4816 13276 4920 13289
rect 4976 14013 5080 14026
rect 4976 13289 5005 14013
rect 5051 13289 5080 14013
rect 4976 13276 5080 13289
rect 5136 14013 5224 14026
rect 5136 13289 5165 14013
rect 5211 13289 5224 14013
rect 5136 13276 5224 13289
rect 5280 14013 5368 14026
rect 5280 13289 5293 14013
rect 5339 13289 5368 14013
rect 5280 13276 5368 13289
rect 5424 14013 5512 14026
rect 5424 13289 5453 14013
rect 5499 13289 5512 14013
rect 5424 13276 5512 13289
rect 3584 12883 3672 12896
rect 3584 12159 3597 12883
rect 3643 12159 3672 12883
rect 3584 12146 3672 12159
rect 3728 12883 3816 12896
rect 3728 12159 3757 12883
rect 3803 12159 3816 12883
rect 3728 12146 3816 12159
rect 3872 12883 3960 12896
rect 3872 12159 3885 12883
rect 3931 12159 3960 12883
rect 3872 12146 3960 12159
rect 4016 12883 4120 12896
rect 4016 12159 4045 12883
rect 4091 12159 4120 12883
rect 4016 12146 4120 12159
rect 4176 12883 4280 12896
rect 4176 12159 4205 12883
rect 4251 12159 4280 12883
rect 4176 12146 4280 12159
rect 4336 12883 4440 12896
rect 4336 12159 4365 12883
rect 4411 12159 4440 12883
rect 4336 12146 4440 12159
rect 4496 12883 4600 12896
rect 4496 12159 4525 12883
rect 4571 12159 4600 12883
rect 4496 12146 4600 12159
rect 4656 12883 4760 12896
rect 4656 12159 4685 12883
rect 4731 12159 4760 12883
rect 4656 12146 4760 12159
rect 4816 12883 4920 12896
rect 4816 12159 4845 12883
rect 4891 12159 4920 12883
rect 4816 12146 4920 12159
rect 4976 12883 5080 12896
rect 4976 12159 5005 12883
rect 5051 12159 5080 12883
rect 4976 12146 5080 12159
rect 5136 12883 5224 12896
rect 5136 12159 5165 12883
rect 5211 12159 5224 12883
rect 5136 12146 5224 12159
rect 5280 12883 5368 12896
rect 5280 12159 5293 12883
rect 5339 12159 5368 12883
rect 5280 12146 5368 12159
rect 5424 12883 5512 12896
rect 5424 12159 5453 12883
rect 5499 12159 5512 12883
rect 5424 12146 5512 12159
rect 3584 11753 3672 11766
rect 3584 11029 3597 11753
rect 3643 11029 3672 11753
rect 3584 11016 3672 11029
rect 3728 11753 3816 11766
rect 3728 11029 3757 11753
rect 3803 11029 3816 11753
rect 3728 11016 3816 11029
rect 3872 11753 3960 11766
rect 3872 11029 3885 11753
rect 3931 11029 3960 11753
rect 3872 11016 3960 11029
rect 4016 11753 4120 11766
rect 4016 11029 4045 11753
rect 4091 11029 4120 11753
rect 4016 11016 4120 11029
rect 4176 11753 4280 11766
rect 4176 11029 4205 11753
rect 4251 11029 4280 11753
rect 4176 11016 4280 11029
rect 4336 11753 4440 11766
rect 4336 11029 4365 11753
rect 4411 11029 4440 11753
rect 4336 11016 4440 11029
rect 4496 11753 4600 11766
rect 4496 11029 4525 11753
rect 4571 11029 4600 11753
rect 4496 11016 4600 11029
rect 4656 11753 4760 11766
rect 4656 11029 4685 11753
rect 4731 11029 4760 11753
rect 4656 11016 4760 11029
rect 4816 11753 4920 11766
rect 4816 11029 4845 11753
rect 4891 11029 4920 11753
rect 4816 11016 4920 11029
rect 4976 11753 5080 11766
rect 4976 11029 5005 11753
rect 5051 11029 5080 11753
rect 4976 11016 5080 11029
rect 5136 11753 5224 11766
rect 5136 11029 5165 11753
rect 5211 11029 5224 11753
rect 5136 11016 5224 11029
rect 5280 11753 5368 11766
rect 5280 11029 5293 11753
rect 5339 11029 5368 11753
rect 5280 11016 5368 11029
rect 5424 11753 5512 11766
rect 5424 11029 5453 11753
rect 5499 11029 5512 11753
rect 5424 11016 5512 11029
rect 898 10545 986 10558
rect 898 9945 911 10545
rect 957 9945 986 10545
rect 898 9932 986 9945
rect 1098 10545 1202 10558
rect 1098 9945 1127 10545
rect 1173 9945 1202 10545
rect 1098 9932 1202 9945
rect 1314 10545 1418 10558
rect 1314 9945 1343 10545
rect 1389 9945 1418 10545
rect 1314 9932 1418 9945
rect 1530 10545 1634 10558
rect 1530 9945 1559 10545
rect 1605 9945 1634 10545
rect 1530 9932 1634 9945
rect 1746 10545 1850 10558
rect 1746 9945 1775 10545
rect 1821 9945 1850 10545
rect 1746 9932 1850 9945
rect 1962 10545 2066 10558
rect 1962 9945 1991 10545
rect 2037 9945 2066 10545
rect 1962 9932 2066 9945
rect 2178 10545 2282 10558
rect 2178 9945 2207 10545
rect 2253 9945 2282 10545
rect 2178 9932 2282 9945
rect 2394 10545 2498 10558
rect 2394 9945 2423 10545
rect 2469 9945 2498 10545
rect 2394 9932 2498 9945
rect 2610 10545 2714 10558
rect 2610 9945 2639 10545
rect 2685 9945 2714 10545
rect 2610 9932 2714 9945
rect 2826 10545 2930 10558
rect 2826 9945 2855 10545
rect 2901 9945 2930 10545
rect 2826 9932 2930 9945
rect 3042 10545 3130 10558
rect 3042 9945 3071 10545
rect 3117 9945 3130 10545
rect 3042 9932 3130 9945
rect 3584 10623 3672 10636
rect 3584 9899 3597 10623
rect 3643 9899 3672 10623
rect 3584 9886 3672 9899
rect 3728 10623 3816 10636
rect 3728 9899 3757 10623
rect 3803 9899 3816 10623
rect 3728 9886 3816 9899
rect 3872 10623 3960 10636
rect 3872 9899 3885 10623
rect 3931 9899 3960 10623
rect 3872 9886 3960 9899
rect 4016 10623 4120 10636
rect 4016 9899 4045 10623
rect 4091 9899 4120 10623
rect 4016 9886 4120 9899
rect 4176 10623 4280 10636
rect 4176 9899 4205 10623
rect 4251 9899 4280 10623
rect 4176 9886 4280 9899
rect 4336 10623 4440 10636
rect 4336 9899 4365 10623
rect 4411 9899 4440 10623
rect 4336 9886 4440 9899
rect 4496 10623 4600 10636
rect 4496 9899 4525 10623
rect 4571 9899 4600 10623
rect 4496 9886 4600 9899
rect 4656 10623 4760 10636
rect 4656 9899 4685 10623
rect 4731 9899 4760 10623
rect 4656 9886 4760 9899
rect 4816 10623 4920 10636
rect 4816 9899 4845 10623
rect 4891 9899 4920 10623
rect 4816 9886 4920 9899
rect 4976 10623 5080 10636
rect 4976 9899 5005 10623
rect 5051 9899 5080 10623
rect 4976 9886 5080 9899
rect 5136 10623 5224 10636
rect 5136 9899 5165 10623
rect 5211 9899 5224 10623
rect 5136 9886 5224 9899
rect 5280 10623 5368 10636
rect 5280 9899 5293 10623
rect 5339 9899 5368 10623
rect 5280 9886 5368 9899
rect 5424 10623 5512 10636
rect 5424 9899 5453 10623
rect 5499 9899 5512 10623
rect 5424 9886 5512 9899
rect 898 9783 986 9796
rect 898 9183 911 9783
rect 957 9183 986 9783
rect 898 9170 986 9183
rect 1098 9783 1202 9796
rect 1098 9183 1127 9783
rect 1173 9183 1202 9783
rect 1098 9170 1202 9183
rect 1314 9783 1418 9796
rect 1314 9183 1343 9783
rect 1389 9183 1418 9783
rect 1314 9170 1418 9183
rect 1530 9783 1634 9796
rect 1530 9183 1559 9783
rect 1605 9183 1634 9783
rect 1530 9170 1634 9183
rect 1746 9783 1850 9796
rect 1746 9183 1775 9783
rect 1821 9183 1850 9783
rect 1746 9170 1850 9183
rect 1962 9783 2066 9796
rect 1962 9183 1991 9783
rect 2037 9183 2066 9783
rect 1962 9170 2066 9183
rect 2178 9783 2282 9796
rect 2178 9183 2207 9783
rect 2253 9183 2282 9783
rect 2178 9170 2282 9183
rect 2394 9783 2498 9796
rect 2394 9183 2423 9783
rect 2469 9183 2498 9783
rect 2394 9170 2498 9183
rect 2610 9783 2714 9796
rect 2610 9183 2639 9783
rect 2685 9183 2714 9783
rect 2610 9170 2714 9183
rect 2826 9783 2930 9796
rect 2826 9183 2855 9783
rect 2901 9183 2930 9783
rect 2826 9170 2930 9183
rect 3042 9783 3130 9796
rect 3042 9183 3071 9783
rect 3117 9183 3130 9783
rect 3042 9170 3130 9183
rect 898 9021 986 9034
rect 898 8421 911 9021
rect 957 8421 986 9021
rect 898 8408 986 8421
rect 1098 9021 1202 9034
rect 1098 8421 1127 9021
rect 1173 8421 1202 9021
rect 1098 8408 1202 8421
rect 1314 9021 1418 9034
rect 1314 8421 1343 9021
rect 1389 8421 1418 9021
rect 1314 8408 1418 8421
rect 1530 9021 1634 9034
rect 1530 8421 1559 9021
rect 1605 8421 1634 9021
rect 1530 8408 1634 8421
rect 1746 9021 1850 9034
rect 1746 8421 1775 9021
rect 1821 8421 1850 9021
rect 1746 8408 1850 8421
rect 1962 9021 2066 9034
rect 1962 8421 1991 9021
rect 2037 8421 2066 9021
rect 1962 8408 2066 8421
rect 2178 9021 2282 9034
rect 2178 8421 2207 9021
rect 2253 8421 2282 9021
rect 2178 8408 2282 8421
rect 2394 9021 2498 9034
rect 2394 8421 2423 9021
rect 2469 8421 2498 9021
rect 2394 8408 2498 8421
rect 2610 9021 2714 9034
rect 2610 8421 2639 9021
rect 2685 8421 2714 9021
rect 2610 8408 2714 8421
rect 2826 9021 2930 9034
rect 2826 8421 2855 9021
rect 2901 8421 2930 9021
rect 2826 8408 2930 8421
rect 3042 9021 3130 9034
rect 3042 8421 3071 9021
rect 3117 8421 3130 9021
rect 3042 8408 3130 8421
rect 3584 9493 3672 9506
rect 3584 8769 3597 9493
rect 3643 8769 3672 9493
rect 3584 8756 3672 8769
rect 3728 9493 3816 9506
rect 3728 8769 3757 9493
rect 3803 8769 3816 9493
rect 3728 8756 3816 8769
rect 3872 9493 3960 9506
rect 3872 8769 3885 9493
rect 3931 8769 3960 9493
rect 3872 8756 3960 8769
rect 4016 9493 4120 9506
rect 4016 8769 4045 9493
rect 4091 8769 4120 9493
rect 4016 8756 4120 8769
rect 4176 9493 4280 9506
rect 4176 8769 4205 9493
rect 4251 8769 4280 9493
rect 4176 8756 4280 8769
rect 4336 9493 4440 9506
rect 4336 8769 4365 9493
rect 4411 8769 4440 9493
rect 4336 8756 4440 8769
rect 4496 9493 4600 9506
rect 4496 8769 4525 9493
rect 4571 8769 4600 9493
rect 4496 8756 4600 8769
rect 4656 9493 4760 9506
rect 4656 8769 4685 9493
rect 4731 8769 4760 9493
rect 4656 8756 4760 8769
rect 4816 9493 4920 9506
rect 4816 8769 4845 9493
rect 4891 8769 4920 9493
rect 4816 8756 4920 8769
rect 4976 9493 5080 9506
rect 4976 8769 5005 9493
rect 5051 8769 5080 9493
rect 4976 8756 5080 8769
rect 5136 9493 5224 9506
rect 5136 8769 5165 9493
rect 5211 8769 5224 9493
rect 5136 8756 5224 8769
rect 5280 9493 5368 9506
rect 5280 8769 5293 9493
rect 5339 8769 5368 9493
rect 5280 8756 5368 8769
rect 5424 9493 5512 9506
rect 5424 8769 5453 9493
rect 5499 8769 5512 9493
rect 5424 8756 5512 8769
rect 898 8259 986 8272
rect 898 7659 911 8259
rect 957 7659 986 8259
rect 898 7646 986 7659
rect 1098 8259 1202 8272
rect 1098 7659 1127 8259
rect 1173 7659 1202 8259
rect 1098 7646 1202 7659
rect 1314 8259 1418 8272
rect 1314 7659 1343 8259
rect 1389 7659 1418 8259
rect 1314 7646 1418 7659
rect 1530 8259 1634 8272
rect 1530 7659 1559 8259
rect 1605 7659 1634 8259
rect 1530 7646 1634 7659
rect 1746 8259 1850 8272
rect 1746 7659 1775 8259
rect 1821 7659 1850 8259
rect 1746 7646 1850 7659
rect 1962 8259 2066 8272
rect 1962 7659 1991 8259
rect 2037 7659 2066 8259
rect 1962 7646 2066 7659
rect 2178 8259 2282 8272
rect 2178 7659 2207 8259
rect 2253 7659 2282 8259
rect 2178 7646 2282 7659
rect 2394 8259 2498 8272
rect 2394 7659 2423 8259
rect 2469 7659 2498 8259
rect 2394 7646 2498 7659
rect 2610 8259 2714 8272
rect 2610 7659 2639 8259
rect 2685 7659 2714 8259
rect 2610 7646 2714 7659
rect 2826 8259 2930 8272
rect 2826 7659 2855 8259
rect 2901 7659 2930 8259
rect 2826 7646 2930 7659
rect 3042 8259 3130 8272
rect 3042 7659 3071 8259
rect 3117 7659 3130 8259
rect 3042 7646 3130 7659
rect 3584 8363 3672 8376
rect 3584 7639 3597 8363
rect 3643 7639 3672 8363
rect 3584 7626 3672 7639
rect 3728 8363 3816 8376
rect 3728 7639 3757 8363
rect 3803 7639 3816 8363
rect 3728 7626 3816 7639
rect 3872 8363 3960 8376
rect 3872 7639 3885 8363
rect 3931 7639 3960 8363
rect 3872 7626 3960 7639
rect 4016 8363 4120 8376
rect 4016 7639 4045 8363
rect 4091 7639 4120 8363
rect 4016 7626 4120 7639
rect 4176 8363 4280 8376
rect 4176 7639 4205 8363
rect 4251 7639 4280 8363
rect 4176 7626 4280 7639
rect 4336 8363 4440 8376
rect 4336 7639 4365 8363
rect 4411 7639 4440 8363
rect 4336 7626 4440 7639
rect 4496 8363 4600 8376
rect 4496 7639 4525 8363
rect 4571 7639 4600 8363
rect 4496 7626 4600 7639
rect 4656 8363 4760 8376
rect 4656 7639 4685 8363
rect 4731 7639 4760 8363
rect 4656 7626 4760 7639
rect 4816 8363 4920 8376
rect 4816 7639 4845 8363
rect 4891 7639 4920 8363
rect 4816 7626 4920 7639
rect 4976 8363 5080 8376
rect 4976 7639 5005 8363
rect 5051 7639 5080 8363
rect 4976 7626 5080 7639
rect 5136 8363 5224 8376
rect 5136 7639 5165 8363
rect 5211 7639 5224 8363
rect 5136 7626 5224 7639
rect 5280 8363 5368 8376
rect 5280 7639 5293 8363
rect 5339 7639 5368 8363
rect 5280 7626 5368 7639
rect 5424 8363 5512 8376
rect 5424 7639 5453 8363
rect 5499 7639 5512 8363
rect 5424 7626 5512 7639
rect 12066 11364 12154 11377
rect 12066 10764 12079 11364
rect 12125 10764 12154 11364
rect 12066 10751 12154 10764
rect 12210 11364 12298 11377
rect 12210 10764 12239 11364
rect 12285 10764 12298 11364
rect 12210 10751 12298 10764
rect 12354 11364 12442 11377
rect 12354 10764 12367 11364
rect 12413 10764 12442 11364
rect 12354 10751 12442 10764
rect 12498 11364 12586 11377
rect 12498 10764 12527 11364
rect 12573 10764 12586 11364
rect 12498 10751 12586 10764
rect 12642 11364 12730 11377
rect 12642 10764 12655 11364
rect 12701 10764 12730 11364
rect 12642 10751 12730 10764
rect 12786 11364 12890 11377
rect 12786 10764 12815 11364
rect 12861 10764 12890 11364
rect 12786 10751 12890 10764
rect 12946 11364 13034 11377
rect 12946 10764 12975 11364
rect 13021 10764 13034 11364
rect 12946 10751 13034 10764
rect 13090 11364 13178 11377
rect 13090 10764 13103 11364
rect 13149 10764 13178 11364
rect 13090 10751 13178 10764
rect 13234 11364 13338 11377
rect 13234 10764 13263 11364
rect 13309 10764 13338 11364
rect 13234 10751 13338 10764
rect 13394 11364 13482 11377
rect 13394 10764 13423 11364
rect 13469 10764 13482 11364
rect 13394 10751 13482 10764
rect 13538 11364 13626 11377
rect 13538 10764 13551 11364
rect 13597 10764 13626 11364
rect 13538 10751 13626 10764
rect 13682 11364 13786 11377
rect 13682 10764 13711 11364
rect 13757 10764 13786 11364
rect 13682 10751 13786 10764
rect 13842 11364 13930 11377
rect 13842 10764 13871 11364
rect 13917 10764 13930 11364
rect 13842 10751 13930 10764
rect 13986 11364 14074 11377
rect 13986 10764 13999 11364
rect 14045 10764 14074 11364
rect 13986 10751 14074 10764
rect 14130 11364 14218 11377
rect 14130 10764 14159 11364
rect 14205 10764 14218 11364
rect 14130 10751 14218 10764
rect 14274 11364 14362 11377
rect 14274 10764 14287 11364
rect 14333 10764 14362 11364
rect 14274 10751 14362 10764
rect 14418 11364 14506 11377
rect 14418 10764 14447 11364
rect 14493 10764 14506 11364
rect 14418 10751 14506 10764
rect 14860 11364 14948 11377
rect 14860 10764 14873 11364
rect 14919 10764 14948 11364
rect 14860 10751 14948 10764
rect 15004 11364 15092 11377
rect 15004 10764 15033 11364
rect 15079 10764 15092 11364
rect 15004 10751 15092 10764
rect 15148 11364 15236 11377
rect 15148 10764 15161 11364
rect 15207 10764 15236 11364
rect 15148 10751 15236 10764
rect 15292 11364 15396 11377
rect 15292 10764 15321 11364
rect 15367 10764 15396 11364
rect 15292 10751 15396 10764
rect 15452 11364 15556 11377
rect 15452 10764 15481 11364
rect 15527 10764 15556 11364
rect 15452 10751 15556 10764
rect 15612 11364 15716 11377
rect 15612 10764 15641 11364
rect 15687 10764 15716 11364
rect 15612 10751 15716 10764
rect 15772 11364 15876 11377
rect 15772 10764 15801 11364
rect 15847 10764 15876 11364
rect 15772 10751 15876 10764
rect 15932 11364 16036 11377
rect 15932 10764 15961 11364
rect 16007 10764 16036 11364
rect 15932 10751 16036 10764
rect 16092 11364 16196 11377
rect 16092 10764 16121 11364
rect 16167 10764 16196 11364
rect 16092 10751 16196 10764
rect 16252 11364 16356 11377
rect 16252 10764 16281 11364
rect 16327 10764 16356 11364
rect 16252 10751 16356 10764
rect 16412 11364 16500 11377
rect 16412 10764 16441 11364
rect 16487 10764 16500 11364
rect 16412 10751 16500 10764
rect 16556 11364 16644 11377
rect 16556 10764 16569 11364
rect 16615 10764 16644 11364
rect 16556 10751 16644 10764
rect 16700 11364 16788 11377
rect 16700 10764 16729 11364
rect 16775 10764 16788 11364
rect 16700 10751 16788 10764
rect 12066 10328 12154 10341
rect 12066 9728 12079 10328
rect 12125 9728 12154 10328
rect 12066 9715 12154 9728
rect 12210 10328 12298 10341
rect 12210 9728 12239 10328
rect 12285 9728 12298 10328
rect 12210 9715 12298 9728
rect 12354 10328 12442 10341
rect 12354 9728 12367 10328
rect 12413 9728 12442 10328
rect 12354 9715 12442 9728
rect 12498 10328 12586 10341
rect 12498 9728 12527 10328
rect 12573 9728 12586 10328
rect 12498 9715 12586 9728
rect 12642 10328 12730 10341
rect 12642 9728 12655 10328
rect 12701 9728 12730 10328
rect 12642 9715 12730 9728
rect 12786 10328 12890 10341
rect 12786 9728 12815 10328
rect 12861 9728 12890 10328
rect 12786 9715 12890 9728
rect 12946 10328 13034 10341
rect 12946 9728 12975 10328
rect 13021 9728 13034 10328
rect 12946 9715 13034 9728
rect 13090 10328 13178 10341
rect 13090 9728 13103 10328
rect 13149 9728 13178 10328
rect 13090 9715 13178 9728
rect 13234 10328 13338 10341
rect 13234 9728 13263 10328
rect 13309 9728 13338 10328
rect 13234 9715 13338 9728
rect 13394 10328 13482 10341
rect 13394 9728 13423 10328
rect 13469 9728 13482 10328
rect 13394 9715 13482 9728
rect 13538 10328 13626 10341
rect 13538 9728 13551 10328
rect 13597 9728 13626 10328
rect 13538 9715 13626 9728
rect 13682 10328 13786 10341
rect 13682 9728 13711 10328
rect 13757 9728 13786 10328
rect 13682 9715 13786 9728
rect 13842 10328 13930 10341
rect 13842 9728 13871 10328
rect 13917 9728 13930 10328
rect 13842 9715 13930 9728
rect 13986 10328 14074 10341
rect 13986 9728 13999 10328
rect 14045 9728 14074 10328
rect 13986 9715 14074 9728
rect 14130 10328 14218 10341
rect 14130 9728 14159 10328
rect 14205 9728 14218 10328
rect 14130 9715 14218 9728
rect 14274 10328 14362 10341
rect 14274 9728 14287 10328
rect 14333 9728 14362 10328
rect 14274 9715 14362 9728
rect 14418 10328 14506 10341
rect 14418 9728 14447 10328
rect 14493 9728 14506 10328
rect 14418 9715 14506 9728
rect 14860 10328 14948 10341
rect 14860 9728 14873 10328
rect 14919 9728 14948 10328
rect 14860 9715 14948 9728
rect 15004 10328 15092 10341
rect 15004 9728 15033 10328
rect 15079 9728 15092 10328
rect 15004 9715 15092 9728
rect 15148 10328 15236 10341
rect 15148 9728 15161 10328
rect 15207 9728 15236 10328
rect 15148 9715 15236 9728
rect 15292 10328 15396 10341
rect 15292 9728 15321 10328
rect 15367 9728 15396 10328
rect 15292 9715 15396 9728
rect 15452 10328 15556 10341
rect 15452 9728 15481 10328
rect 15527 9728 15556 10328
rect 15452 9715 15556 9728
rect 15612 10328 15716 10341
rect 15612 9728 15641 10328
rect 15687 9728 15716 10328
rect 15612 9715 15716 9728
rect 15772 10328 15876 10341
rect 15772 9728 15801 10328
rect 15847 9728 15876 10328
rect 15772 9715 15876 9728
rect 15932 10328 16036 10341
rect 15932 9728 15961 10328
rect 16007 9728 16036 10328
rect 15932 9715 16036 9728
rect 16092 10328 16196 10341
rect 16092 9728 16121 10328
rect 16167 9728 16196 10328
rect 16092 9715 16196 9728
rect 16252 10328 16356 10341
rect 16252 9728 16281 10328
rect 16327 9728 16356 10328
rect 16252 9715 16356 9728
rect 16412 10328 16500 10341
rect 16412 9728 16441 10328
rect 16487 9728 16500 10328
rect 16412 9715 16500 9728
rect 16556 10328 16644 10341
rect 16556 9728 16569 10328
rect 16615 9728 16644 10328
rect 16556 9715 16644 9728
rect 16700 10328 16788 10341
rect 16700 9728 16729 10328
rect 16775 9728 16788 10328
rect 16700 9715 16788 9728
rect 12066 9292 12154 9305
rect 12066 8692 12079 9292
rect 12125 8692 12154 9292
rect 12066 8679 12154 8692
rect 12210 9292 12298 9305
rect 12210 8692 12239 9292
rect 12285 8692 12298 9292
rect 12210 8679 12298 8692
rect 12354 9292 12442 9305
rect 12354 8692 12367 9292
rect 12413 8692 12442 9292
rect 12354 8679 12442 8692
rect 12498 9292 12586 9305
rect 12498 8692 12527 9292
rect 12573 8692 12586 9292
rect 12498 8679 12586 8692
rect 12642 9292 12730 9305
rect 12642 8692 12655 9292
rect 12701 8692 12730 9292
rect 12642 8679 12730 8692
rect 12786 9292 12890 9305
rect 12786 8692 12815 9292
rect 12861 8692 12890 9292
rect 12786 8679 12890 8692
rect 12946 9292 13034 9305
rect 12946 8692 12975 9292
rect 13021 8692 13034 9292
rect 12946 8679 13034 8692
rect 13090 9292 13178 9305
rect 13090 8692 13103 9292
rect 13149 8692 13178 9292
rect 13090 8679 13178 8692
rect 13234 9292 13338 9305
rect 13234 8692 13263 9292
rect 13309 8692 13338 9292
rect 13234 8679 13338 8692
rect 13394 9292 13482 9305
rect 13394 8692 13423 9292
rect 13469 8692 13482 9292
rect 13394 8679 13482 8692
rect 13538 9292 13626 9305
rect 13538 8692 13551 9292
rect 13597 8692 13626 9292
rect 13538 8679 13626 8692
rect 13682 9292 13786 9305
rect 13682 8692 13711 9292
rect 13757 8692 13786 9292
rect 13682 8679 13786 8692
rect 13842 9292 13930 9305
rect 13842 8692 13871 9292
rect 13917 8692 13930 9292
rect 13842 8679 13930 8692
rect 13986 9292 14074 9305
rect 13986 8692 13999 9292
rect 14045 8692 14074 9292
rect 13986 8679 14074 8692
rect 14130 9292 14218 9305
rect 14130 8692 14159 9292
rect 14205 8692 14218 9292
rect 14130 8679 14218 8692
rect 14274 9292 14362 9305
rect 14274 8692 14287 9292
rect 14333 8692 14362 9292
rect 14274 8679 14362 8692
rect 14418 9292 14506 9305
rect 14418 8692 14447 9292
rect 14493 8692 14506 9292
rect 14418 8679 14506 8692
rect 14860 9292 14948 9305
rect 14860 8692 14873 9292
rect 14919 8692 14948 9292
rect 14860 8679 14948 8692
rect 15004 9292 15092 9305
rect 15004 8692 15033 9292
rect 15079 8692 15092 9292
rect 15004 8679 15092 8692
rect 15148 9292 15236 9305
rect 15148 8692 15161 9292
rect 15207 8692 15236 9292
rect 15148 8679 15236 8692
rect 15292 9292 15396 9305
rect 15292 8692 15321 9292
rect 15367 8692 15396 9292
rect 15292 8679 15396 8692
rect 15452 9292 15556 9305
rect 15452 8692 15481 9292
rect 15527 8692 15556 9292
rect 15452 8679 15556 8692
rect 15612 9292 15716 9305
rect 15612 8692 15641 9292
rect 15687 8692 15716 9292
rect 15612 8679 15716 8692
rect 15772 9292 15876 9305
rect 15772 8692 15801 9292
rect 15847 8692 15876 9292
rect 15772 8679 15876 8692
rect 15932 9292 16036 9305
rect 15932 8692 15961 9292
rect 16007 8692 16036 9292
rect 15932 8679 16036 8692
rect 16092 9292 16196 9305
rect 16092 8692 16121 9292
rect 16167 8692 16196 9292
rect 16092 8679 16196 8692
rect 16252 9292 16356 9305
rect 16252 8692 16281 9292
rect 16327 8692 16356 9292
rect 16252 8679 16356 8692
rect 16412 9292 16500 9305
rect 16412 8692 16441 9292
rect 16487 8692 16500 9292
rect 16412 8679 16500 8692
rect 16556 9292 16644 9305
rect 16556 8692 16569 9292
rect 16615 8692 16644 9292
rect 16556 8679 16644 8692
rect 16700 9292 16788 9305
rect 16700 8692 16729 9292
rect 16775 8692 16788 9292
rect 16700 8679 16788 8692
rect 12066 8256 12154 8269
rect 12066 7656 12079 8256
rect 12125 7656 12154 8256
rect 12066 7643 12154 7656
rect 12210 8256 12298 8269
rect 12210 7656 12239 8256
rect 12285 7656 12298 8256
rect 12210 7643 12298 7656
rect 12354 8256 12442 8269
rect 12354 7656 12367 8256
rect 12413 7656 12442 8256
rect 12354 7643 12442 7656
rect 12498 8256 12586 8269
rect 12498 7656 12527 8256
rect 12573 7656 12586 8256
rect 12498 7643 12586 7656
rect 12642 8256 12730 8269
rect 12642 7656 12655 8256
rect 12701 7656 12730 8256
rect 12642 7643 12730 7656
rect 12786 8256 12890 8269
rect 12786 7656 12815 8256
rect 12861 7656 12890 8256
rect 12786 7643 12890 7656
rect 12946 8256 13034 8269
rect 12946 7656 12975 8256
rect 13021 7656 13034 8256
rect 12946 7643 13034 7656
rect 13090 8256 13178 8269
rect 13090 7656 13103 8256
rect 13149 7656 13178 8256
rect 13090 7643 13178 7656
rect 13234 8256 13338 8269
rect 13234 7656 13263 8256
rect 13309 7656 13338 8256
rect 13234 7643 13338 7656
rect 13394 8256 13482 8269
rect 13394 7656 13423 8256
rect 13469 7656 13482 8256
rect 13394 7643 13482 7656
rect 13538 8256 13626 8269
rect 13538 7656 13551 8256
rect 13597 7656 13626 8256
rect 13538 7643 13626 7656
rect 13682 8256 13786 8269
rect 13682 7656 13711 8256
rect 13757 7656 13786 8256
rect 13682 7643 13786 7656
rect 13842 8256 13930 8269
rect 13842 7656 13871 8256
rect 13917 7656 13930 8256
rect 13842 7643 13930 7656
rect 13986 8256 14074 8269
rect 13986 7656 13999 8256
rect 14045 7656 14074 8256
rect 13986 7643 14074 7656
rect 14130 8256 14218 8269
rect 14130 7656 14159 8256
rect 14205 7656 14218 8256
rect 14130 7643 14218 7656
rect 14274 8256 14362 8269
rect 14274 7656 14287 8256
rect 14333 7656 14362 8256
rect 14274 7643 14362 7656
rect 14418 8256 14506 8269
rect 14418 7656 14447 8256
rect 14493 7656 14506 8256
rect 14418 7643 14506 7656
rect 14860 8256 14948 8269
rect 14860 7656 14873 8256
rect 14919 7656 14948 8256
rect 14860 7643 14948 7656
rect 15004 8256 15092 8269
rect 15004 7656 15033 8256
rect 15079 7656 15092 8256
rect 15004 7643 15092 7656
rect 15148 8256 15236 8269
rect 15148 7656 15161 8256
rect 15207 7656 15236 8256
rect 15148 7643 15236 7656
rect 15292 8256 15396 8269
rect 15292 7656 15321 8256
rect 15367 7656 15396 8256
rect 15292 7643 15396 7656
rect 15452 8256 15556 8269
rect 15452 7656 15481 8256
rect 15527 7656 15556 8256
rect 15452 7643 15556 7656
rect 15612 8256 15716 8269
rect 15612 7656 15641 8256
rect 15687 7656 15716 8256
rect 15612 7643 15716 7656
rect 15772 8256 15876 8269
rect 15772 7656 15801 8256
rect 15847 7656 15876 8256
rect 15772 7643 15876 7656
rect 15932 8256 16036 8269
rect 15932 7656 15961 8256
rect 16007 7656 16036 8256
rect 15932 7643 16036 7656
rect 16092 8256 16196 8269
rect 16092 7656 16121 8256
rect 16167 7656 16196 8256
rect 16092 7643 16196 7656
rect 16252 8256 16356 8269
rect 16252 7656 16281 8256
rect 16327 7656 16356 8256
rect 16252 7643 16356 7656
rect 16412 8256 16500 8269
rect 16412 7656 16441 8256
rect 16487 7656 16500 8256
rect 16412 7643 16500 7656
rect 16556 8256 16644 8269
rect 16556 7656 16569 8256
rect 16615 7656 16644 8256
rect 16556 7643 16644 7656
rect 16700 8256 16788 8269
rect 16700 7656 16729 8256
rect 16775 7656 16788 8256
rect 16700 7643 16788 7656
rect 33116 11676 33204 11689
rect 33116 11102 33129 11676
rect 33175 11102 33204 11676
rect 33116 11089 33204 11102
rect 33260 11676 33348 11689
rect 33260 11102 33289 11676
rect 33335 11102 33348 11676
rect 33260 11089 33348 11102
rect 33404 11676 33492 11689
rect 33404 11102 33417 11676
rect 33463 11102 33492 11676
rect 33404 11089 33492 11102
rect 33548 11676 33652 11689
rect 33548 11102 33577 11676
rect 33623 11102 33652 11676
rect 33548 11089 33652 11102
rect 33708 11676 33812 11689
rect 33708 11102 33737 11676
rect 33783 11102 33812 11676
rect 33708 11089 33812 11102
rect 33868 11676 33972 11689
rect 33868 11102 33897 11676
rect 33943 11102 33972 11676
rect 33868 11089 33972 11102
rect 34028 11676 34132 11689
rect 34028 11102 34057 11676
rect 34103 11102 34132 11676
rect 34028 11089 34132 11102
rect 34188 11676 34292 11689
rect 34188 11102 34217 11676
rect 34263 11102 34292 11676
rect 34188 11089 34292 11102
rect 34348 11676 34452 11689
rect 34348 11102 34377 11676
rect 34423 11102 34452 11676
rect 34348 11089 34452 11102
rect 34508 11676 34612 11689
rect 34508 11102 34537 11676
rect 34583 11102 34612 11676
rect 34508 11089 34612 11102
rect 34668 11676 34772 11689
rect 34668 11102 34697 11676
rect 34743 11102 34772 11676
rect 34668 11089 34772 11102
rect 34828 11676 34932 11689
rect 34828 11102 34857 11676
rect 34903 11102 34932 11676
rect 34828 11089 34932 11102
rect 34988 11676 35092 11689
rect 34988 11102 35017 11676
rect 35063 11102 35092 11676
rect 34988 11089 35092 11102
rect 35148 11676 35252 11689
rect 35148 11102 35177 11676
rect 35223 11102 35252 11676
rect 35148 11089 35252 11102
rect 35308 11676 35412 11689
rect 35308 11102 35337 11676
rect 35383 11102 35412 11676
rect 35308 11089 35412 11102
rect 35468 11676 35572 11689
rect 35468 11102 35497 11676
rect 35543 11102 35572 11676
rect 35468 11089 35572 11102
rect 35628 11676 35732 11689
rect 35628 11102 35657 11676
rect 35703 11102 35732 11676
rect 35628 11089 35732 11102
rect 35788 11676 35892 11689
rect 35788 11102 35817 11676
rect 35863 11102 35892 11676
rect 35788 11089 35892 11102
rect 35948 11676 36036 11689
rect 35948 11102 35977 11676
rect 36023 11102 36036 11676
rect 35948 11089 36036 11102
rect 36092 11676 36180 11689
rect 36092 11102 36105 11676
rect 36151 11102 36180 11676
rect 36092 11089 36180 11102
rect 36236 11676 36324 11689
rect 36236 11102 36265 11676
rect 36311 11102 36324 11676
rect 36236 11089 36324 11102
rect 37252 11676 37340 11689
rect 37252 11102 37265 11676
rect 37311 11102 37340 11676
rect 37252 11089 37340 11102
rect 37396 11676 37484 11689
rect 37396 11102 37425 11676
rect 37471 11102 37484 11676
rect 37396 11089 37484 11102
rect 37540 11676 37628 11689
rect 37540 11102 37553 11676
rect 37599 11102 37628 11676
rect 37540 11089 37628 11102
rect 37684 11676 37788 11689
rect 37684 11102 37713 11676
rect 37759 11102 37788 11676
rect 37684 11089 37788 11102
rect 37844 11676 37948 11689
rect 37844 11102 37873 11676
rect 37919 11102 37948 11676
rect 37844 11089 37948 11102
rect 38004 11676 38108 11689
rect 38004 11102 38033 11676
rect 38079 11102 38108 11676
rect 38004 11089 38108 11102
rect 38164 11676 38268 11689
rect 38164 11102 38193 11676
rect 38239 11102 38268 11676
rect 38164 11089 38268 11102
rect 38324 11676 38428 11689
rect 38324 11102 38353 11676
rect 38399 11102 38428 11676
rect 38324 11089 38428 11102
rect 38484 11676 38588 11689
rect 38484 11102 38513 11676
rect 38559 11102 38588 11676
rect 38484 11089 38588 11102
rect 38644 11676 38748 11689
rect 38644 11102 38673 11676
rect 38719 11102 38748 11676
rect 38644 11089 38748 11102
rect 38804 11676 38908 11689
rect 38804 11102 38833 11676
rect 38879 11102 38908 11676
rect 38804 11089 38908 11102
rect 38964 11676 39068 11689
rect 38964 11102 38993 11676
rect 39039 11102 39068 11676
rect 38964 11089 39068 11102
rect 39124 11676 39228 11689
rect 39124 11102 39153 11676
rect 39199 11102 39228 11676
rect 39124 11089 39228 11102
rect 39284 11676 39388 11689
rect 39284 11102 39313 11676
rect 39359 11102 39388 11676
rect 39284 11089 39388 11102
rect 39444 11676 39548 11689
rect 39444 11102 39473 11676
rect 39519 11102 39548 11676
rect 39444 11089 39548 11102
rect 39604 11676 39708 11689
rect 39604 11102 39633 11676
rect 39679 11102 39708 11676
rect 39604 11089 39708 11102
rect 39764 11676 39868 11689
rect 39764 11102 39793 11676
rect 39839 11102 39868 11676
rect 39764 11089 39868 11102
rect 39924 11676 40028 11689
rect 39924 11102 39953 11676
rect 39999 11102 40028 11676
rect 39924 11089 40028 11102
rect 40084 11676 40172 11689
rect 40084 11102 40113 11676
rect 40159 11102 40172 11676
rect 40084 11089 40172 11102
rect 40228 11676 40316 11689
rect 40228 11102 40241 11676
rect 40287 11102 40316 11676
rect 40228 11089 40316 11102
rect 40372 11676 40460 11689
rect 40372 11102 40401 11676
rect 40447 11102 40460 11676
rect 40372 11089 40460 11102
rect 33116 10616 33204 10629
rect 33116 10042 33129 10616
rect 33175 10042 33204 10616
rect 33116 10029 33204 10042
rect 33260 10616 33348 10629
rect 33260 10042 33289 10616
rect 33335 10042 33348 10616
rect 33260 10029 33348 10042
rect 33404 10616 33492 10629
rect 33404 10042 33417 10616
rect 33463 10042 33492 10616
rect 33404 10029 33492 10042
rect 33548 10616 33652 10629
rect 33548 10042 33577 10616
rect 33623 10042 33652 10616
rect 33548 10029 33652 10042
rect 33708 10616 33812 10629
rect 33708 10042 33737 10616
rect 33783 10042 33812 10616
rect 33708 10029 33812 10042
rect 33868 10616 33972 10629
rect 33868 10042 33897 10616
rect 33943 10042 33972 10616
rect 33868 10029 33972 10042
rect 34028 10616 34132 10629
rect 34028 10042 34057 10616
rect 34103 10042 34132 10616
rect 34028 10029 34132 10042
rect 34188 10616 34292 10629
rect 34188 10042 34217 10616
rect 34263 10042 34292 10616
rect 34188 10029 34292 10042
rect 34348 10616 34452 10629
rect 34348 10042 34377 10616
rect 34423 10042 34452 10616
rect 34348 10029 34452 10042
rect 34508 10616 34612 10629
rect 34508 10042 34537 10616
rect 34583 10042 34612 10616
rect 34508 10029 34612 10042
rect 34668 10616 34772 10629
rect 34668 10042 34697 10616
rect 34743 10042 34772 10616
rect 34668 10029 34772 10042
rect 34828 10616 34932 10629
rect 34828 10042 34857 10616
rect 34903 10042 34932 10616
rect 34828 10029 34932 10042
rect 34988 10616 35092 10629
rect 34988 10042 35017 10616
rect 35063 10042 35092 10616
rect 34988 10029 35092 10042
rect 35148 10616 35252 10629
rect 35148 10042 35177 10616
rect 35223 10042 35252 10616
rect 35148 10029 35252 10042
rect 35308 10616 35412 10629
rect 35308 10042 35337 10616
rect 35383 10042 35412 10616
rect 35308 10029 35412 10042
rect 35468 10616 35572 10629
rect 35468 10042 35497 10616
rect 35543 10042 35572 10616
rect 35468 10029 35572 10042
rect 35628 10616 35732 10629
rect 35628 10042 35657 10616
rect 35703 10042 35732 10616
rect 35628 10029 35732 10042
rect 35788 10616 35892 10629
rect 35788 10042 35817 10616
rect 35863 10042 35892 10616
rect 35788 10029 35892 10042
rect 35948 10616 36036 10629
rect 35948 10042 35977 10616
rect 36023 10042 36036 10616
rect 35948 10029 36036 10042
rect 36092 10616 36180 10629
rect 36092 10042 36105 10616
rect 36151 10042 36180 10616
rect 36092 10029 36180 10042
rect 36236 10616 36324 10629
rect 36236 10042 36265 10616
rect 36311 10042 36324 10616
rect 36236 10029 36324 10042
rect 37252 10616 37340 10629
rect 37252 10042 37265 10616
rect 37311 10042 37340 10616
rect 37252 10029 37340 10042
rect 37396 10616 37484 10629
rect 37396 10042 37425 10616
rect 37471 10042 37484 10616
rect 37396 10029 37484 10042
rect 37540 10616 37628 10629
rect 37540 10042 37553 10616
rect 37599 10042 37628 10616
rect 37540 10029 37628 10042
rect 37684 10616 37788 10629
rect 37684 10042 37713 10616
rect 37759 10042 37788 10616
rect 37684 10029 37788 10042
rect 37844 10616 37948 10629
rect 37844 10042 37873 10616
rect 37919 10042 37948 10616
rect 37844 10029 37948 10042
rect 38004 10616 38108 10629
rect 38004 10042 38033 10616
rect 38079 10042 38108 10616
rect 38004 10029 38108 10042
rect 38164 10616 38268 10629
rect 38164 10042 38193 10616
rect 38239 10042 38268 10616
rect 38164 10029 38268 10042
rect 38324 10616 38428 10629
rect 38324 10042 38353 10616
rect 38399 10042 38428 10616
rect 38324 10029 38428 10042
rect 38484 10616 38588 10629
rect 38484 10042 38513 10616
rect 38559 10042 38588 10616
rect 38484 10029 38588 10042
rect 38644 10616 38748 10629
rect 38644 10042 38673 10616
rect 38719 10042 38748 10616
rect 38644 10029 38748 10042
rect 38804 10616 38908 10629
rect 38804 10042 38833 10616
rect 38879 10042 38908 10616
rect 38804 10029 38908 10042
rect 38964 10616 39068 10629
rect 38964 10042 38993 10616
rect 39039 10042 39068 10616
rect 38964 10029 39068 10042
rect 39124 10616 39228 10629
rect 39124 10042 39153 10616
rect 39199 10042 39228 10616
rect 39124 10029 39228 10042
rect 39284 10616 39388 10629
rect 39284 10042 39313 10616
rect 39359 10042 39388 10616
rect 39284 10029 39388 10042
rect 39444 10616 39548 10629
rect 39444 10042 39473 10616
rect 39519 10042 39548 10616
rect 39444 10029 39548 10042
rect 39604 10616 39708 10629
rect 39604 10042 39633 10616
rect 39679 10042 39708 10616
rect 39604 10029 39708 10042
rect 39764 10616 39868 10629
rect 39764 10042 39793 10616
rect 39839 10042 39868 10616
rect 39764 10029 39868 10042
rect 39924 10616 40028 10629
rect 39924 10042 39953 10616
rect 39999 10042 40028 10616
rect 39924 10029 40028 10042
rect 40084 10616 40172 10629
rect 40084 10042 40113 10616
rect 40159 10042 40172 10616
rect 40084 10029 40172 10042
rect 40228 10616 40316 10629
rect 40228 10042 40241 10616
rect 40287 10042 40316 10616
rect 40228 10029 40316 10042
rect 40372 10616 40460 10629
rect 40372 10042 40401 10616
rect 40447 10042 40460 10616
rect 40372 10029 40460 10042
rect 33116 9556 33204 9569
rect 33116 8982 33129 9556
rect 33175 8982 33204 9556
rect 33116 8969 33204 8982
rect 33260 9556 33348 9569
rect 33260 8982 33289 9556
rect 33335 8982 33348 9556
rect 33260 8969 33348 8982
rect 33404 9556 33492 9569
rect 33404 8982 33417 9556
rect 33463 8982 33492 9556
rect 33404 8969 33492 8982
rect 33548 9556 33652 9569
rect 33548 8982 33577 9556
rect 33623 8982 33652 9556
rect 33548 8969 33652 8982
rect 33708 9556 33812 9569
rect 33708 8982 33737 9556
rect 33783 8982 33812 9556
rect 33708 8969 33812 8982
rect 33868 9556 33972 9569
rect 33868 8982 33897 9556
rect 33943 8982 33972 9556
rect 33868 8969 33972 8982
rect 34028 9556 34132 9569
rect 34028 8982 34057 9556
rect 34103 8982 34132 9556
rect 34028 8969 34132 8982
rect 34188 9556 34292 9569
rect 34188 8982 34217 9556
rect 34263 8982 34292 9556
rect 34188 8969 34292 8982
rect 34348 9556 34452 9569
rect 34348 8982 34377 9556
rect 34423 8982 34452 9556
rect 34348 8969 34452 8982
rect 34508 9556 34612 9569
rect 34508 8982 34537 9556
rect 34583 8982 34612 9556
rect 34508 8969 34612 8982
rect 34668 9556 34772 9569
rect 34668 8982 34697 9556
rect 34743 8982 34772 9556
rect 34668 8969 34772 8982
rect 34828 9556 34932 9569
rect 34828 8982 34857 9556
rect 34903 8982 34932 9556
rect 34828 8969 34932 8982
rect 34988 9556 35092 9569
rect 34988 8982 35017 9556
rect 35063 8982 35092 9556
rect 34988 8969 35092 8982
rect 35148 9556 35252 9569
rect 35148 8982 35177 9556
rect 35223 8982 35252 9556
rect 35148 8969 35252 8982
rect 35308 9556 35412 9569
rect 35308 8982 35337 9556
rect 35383 8982 35412 9556
rect 35308 8969 35412 8982
rect 35468 9556 35572 9569
rect 35468 8982 35497 9556
rect 35543 8982 35572 9556
rect 35468 8969 35572 8982
rect 35628 9556 35732 9569
rect 35628 8982 35657 9556
rect 35703 8982 35732 9556
rect 35628 8969 35732 8982
rect 35788 9556 35892 9569
rect 35788 8982 35817 9556
rect 35863 8982 35892 9556
rect 35788 8969 35892 8982
rect 35948 9556 36036 9569
rect 35948 8982 35977 9556
rect 36023 8982 36036 9556
rect 35948 8969 36036 8982
rect 36092 9556 36180 9569
rect 36092 8982 36105 9556
rect 36151 8982 36180 9556
rect 36092 8969 36180 8982
rect 36236 9556 36324 9569
rect 36236 8982 36265 9556
rect 36311 8982 36324 9556
rect 36236 8969 36324 8982
rect 37252 9556 37340 9569
rect 37252 8982 37265 9556
rect 37311 8982 37340 9556
rect 37252 8969 37340 8982
rect 37396 9556 37484 9569
rect 37396 8982 37425 9556
rect 37471 8982 37484 9556
rect 37396 8969 37484 8982
rect 37540 9556 37628 9569
rect 37540 8982 37553 9556
rect 37599 8982 37628 9556
rect 37540 8969 37628 8982
rect 37684 9556 37788 9569
rect 37684 8982 37713 9556
rect 37759 8982 37788 9556
rect 37684 8969 37788 8982
rect 37844 9556 37948 9569
rect 37844 8982 37873 9556
rect 37919 8982 37948 9556
rect 37844 8969 37948 8982
rect 38004 9556 38108 9569
rect 38004 8982 38033 9556
rect 38079 8982 38108 9556
rect 38004 8969 38108 8982
rect 38164 9556 38268 9569
rect 38164 8982 38193 9556
rect 38239 8982 38268 9556
rect 38164 8969 38268 8982
rect 38324 9556 38428 9569
rect 38324 8982 38353 9556
rect 38399 8982 38428 9556
rect 38324 8969 38428 8982
rect 38484 9556 38588 9569
rect 38484 8982 38513 9556
rect 38559 8982 38588 9556
rect 38484 8969 38588 8982
rect 38644 9556 38748 9569
rect 38644 8982 38673 9556
rect 38719 8982 38748 9556
rect 38644 8969 38748 8982
rect 38804 9556 38908 9569
rect 38804 8982 38833 9556
rect 38879 8982 38908 9556
rect 38804 8969 38908 8982
rect 38964 9556 39068 9569
rect 38964 8982 38993 9556
rect 39039 8982 39068 9556
rect 38964 8969 39068 8982
rect 39124 9556 39228 9569
rect 39124 8982 39153 9556
rect 39199 8982 39228 9556
rect 39124 8969 39228 8982
rect 39284 9556 39388 9569
rect 39284 8982 39313 9556
rect 39359 8982 39388 9556
rect 39284 8969 39388 8982
rect 39444 9556 39548 9569
rect 39444 8982 39473 9556
rect 39519 8982 39548 9556
rect 39444 8969 39548 8982
rect 39604 9556 39708 9569
rect 39604 8982 39633 9556
rect 39679 8982 39708 9556
rect 39604 8969 39708 8982
rect 39764 9556 39868 9569
rect 39764 8982 39793 9556
rect 39839 8982 39868 9556
rect 39764 8969 39868 8982
rect 39924 9556 40028 9569
rect 39924 8982 39953 9556
rect 39999 8982 40028 9556
rect 39924 8969 40028 8982
rect 40084 9556 40172 9569
rect 40084 8982 40113 9556
rect 40159 8982 40172 9556
rect 40084 8969 40172 8982
rect 40228 9556 40316 9569
rect 40228 8982 40241 9556
rect 40287 8982 40316 9556
rect 40228 8969 40316 8982
rect 40372 9556 40460 9569
rect 40372 8982 40401 9556
rect 40447 8982 40460 9556
rect 40372 8969 40460 8982
rect 33116 8496 33204 8509
rect 33116 7922 33129 8496
rect 33175 7922 33204 8496
rect 33116 7909 33204 7922
rect 33260 8496 33348 8509
rect 33260 7922 33289 8496
rect 33335 7922 33348 8496
rect 33260 7909 33348 7922
rect 33404 8496 33492 8509
rect 33404 7922 33417 8496
rect 33463 7922 33492 8496
rect 33404 7909 33492 7922
rect 33548 8496 33652 8509
rect 33548 7922 33577 8496
rect 33623 7922 33652 8496
rect 33548 7909 33652 7922
rect 33708 8496 33812 8509
rect 33708 7922 33737 8496
rect 33783 7922 33812 8496
rect 33708 7909 33812 7922
rect 33868 8496 33972 8509
rect 33868 7922 33897 8496
rect 33943 7922 33972 8496
rect 33868 7909 33972 7922
rect 34028 8496 34132 8509
rect 34028 7922 34057 8496
rect 34103 7922 34132 8496
rect 34028 7909 34132 7922
rect 34188 8496 34292 8509
rect 34188 7922 34217 8496
rect 34263 7922 34292 8496
rect 34188 7909 34292 7922
rect 34348 8496 34452 8509
rect 34348 7922 34377 8496
rect 34423 7922 34452 8496
rect 34348 7909 34452 7922
rect 34508 8496 34612 8509
rect 34508 7922 34537 8496
rect 34583 7922 34612 8496
rect 34508 7909 34612 7922
rect 34668 8496 34772 8509
rect 34668 7922 34697 8496
rect 34743 7922 34772 8496
rect 34668 7909 34772 7922
rect 34828 8496 34932 8509
rect 34828 7922 34857 8496
rect 34903 7922 34932 8496
rect 34828 7909 34932 7922
rect 34988 8496 35092 8509
rect 34988 7922 35017 8496
rect 35063 7922 35092 8496
rect 34988 7909 35092 7922
rect 35148 8496 35252 8509
rect 35148 7922 35177 8496
rect 35223 7922 35252 8496
rect 35148 7909 35252 7922
rect 35308 8496 35412 8509
rect 35308 7922 35337 8496
rect 35383 7922 35412 8496
rect 35308 7909 35412 7922
rect 35468 8496 35572 8509
rect 35468 7922 35497 8496
rect 35543 7922 35572 8496
rect 35468 7909 35572 7922
rect 35628 8496 35732 8509
rect 35628 7922 35657 8496
rect 35703 7922 35732 8496
rect 35628 7909 35732 7922
rect 35788 8496 35892 8509
rect 35788 7922 35817 8496
rect 35863 7922 35892 8496
rect 35788 7909 35892 7922
rect 35948 8496 36036 8509
rect 35948 7922 35977 8496
rect 36023 7922 36036 8496
rect 35948 7909 36036 7922
rect 36092 8496 36180 8509
rect 36092 7922 36105 8496
rect 36151 7922 36180 8496
rect 36092 7909 36180 7922
rect 36236 8496 36324 8509
rect 36236 7922 36265 8496
rect 36311 7922 36324 8496
rect 36236 7909 36324 7922
rect 37252 8496 37340 8509
rect 37252 7922 37265 8496
rect 37311 7922 37340 8496
rect 37252 7909 37340 7922
rect 37396 8496 37484 8509
rect 37396 7922 37425 8496
rect 37471 7922 37484 8496
rect 37396 7909 37484 7922
rect 37540 8496 37628 8509
rect 37540 7922 37553 8496
rect 37599 7922 37628 8496
rect 37540 7909 37628 7922
rect 37684 8496 37788 8509
rect 37684 7922 37713 8496
rect 37759 7922 37788 8496
rect 37684 7909 37788 7922
rect 37844 8496 37948 8509
rect 37844 7922 37873 8496
rect 37919 7922 37948 8496
rect 37844 7909 37948 7922
rect 38004 8496 38108 8509
rect 38004 7922 38033 8496
rect 38079 7922 38108 8496
rect 38004 7909 38108 7922
rect 38164 8496 38268 8509
rect 38164 7922 38193 8496
rect 38239 7922 38268 8496
rect 38164 7909 38268 7922
rect 38324 8496 38428 8509
rect 38324 7922 38353 8496
rect 38399 7922 38428 8496
rect 38324 7909 38428 7922
rect 38484 8496 38588 8509
rect 38484 7922 38513 8496
rect 38559 7922 38588 8496
rect 38484 7909 38588 7922
rect 38644 8496 38748 8509
rect 38644 7922 38673 8496
rect 38719 7922 38748 8496
rect 38644 7909 38748 7922
rect 38804 8496 38908 8509
rect 38804 7922 38833 8496
rect 38879 7922 38908 8496
rect 38804 7909 38908 7922
rect 38964 8496 39068 8509
rect 38964 7922 38993 8496
rect 39039 7922 39068 8496
rect 38964 7909 39068 7922
rect 39124 8496 39228 8509
rect 39124 7922 39153 8496
rect 39199 7922 39228 8496
rect 39124 7909 39228 7922
rect 39284 8496 39388 8509
rect 39284 7922 39313 8496
rect 39359 7922 39388 8496
rect 39284 7909 39388 7922
rect 39444 8496 39548 8509
rect 39444 7922 39473 8496
rect 39519 7922 39548 8496
rect 39444 7909 39548 7922
rect 39604 8496 39708 8509
rect 39604 7922 39633 8496
rect 39679 7922 39708 8496
rect 39604 7909 39708 7922
rect 39764 8496 39868 8509
rect 39764 7922 39793 8496
rect 39839 7922 39868 8496
rect 39764 7909 39868 7922
rect 39924 8496 40028 8509
rect 39924 7922 39953 8496
rect 39999 7922 40028 8496
rect 39924 7909 40028 7922
rect 40084 8496 40172 8509
rect 40084 7922 40113 8496
rect 40159 7922 40172 8496
rect 40084 7909 40172 7922
rect 40228 8496 40316 8509
rect 40228 7922 40241 8496
rect 40287 7922 40316 8496
rect 40228 7909 40316 7922
rect 40372 8496 40460 8509
rect 40372 7922 40401 8496
rect 40447 7922 40460 8496
rect 40372 7909 40460 7922
rect 42812 11676 42900 11689
rect 42812 11102 42825 11676
rect 42871 11102 42900 11676
rect 42812 11089 42900 11102
rect 42956 11676 43044 11689
rect 42956 11102 42985 11676
rect 43031 11102 43044 11676
rect 42956 11089 43044 11102
rect 43100 11676 43188 11689
rect 43100 11102 43113 11676
rect 43159 11102 43188 11676
rect 43100 11089 43188 11102
rect 43244 11676 43348 11689
rect 43244 11102 43273 11676
rect 43319 11102 43348 11676
rect 43244 11089 43348 11102
rect 43404 11676 43508 11689
rect 43404 11102 43433 11676
rect 43479 11102 43508 11676
rect 43404 11089 43508 11102
rect 43564 11676 43668 11689
rect 43564 11102 43593 11676
rect 43639 11102 43668 11676
rect 43564 11089 43668 11102
rect 43724 11676 43828 11689
rect 43724 11102 43753 11676
rect 43799 11102 43828 11676
rect 43724 11089 43828 11102
rect 43884 11676 43988 11689
rect 43884 11102 43913 11676
rect 43959 11102 43988 11676
rect 43884 11089 43988 11102
rect 44044 11676 44148 11689
rect 44044 11102 44073 11676
rect 44119 11102 44148 11676
rect 44044 11089 44148 11102
rect 44204 11676 44308 11689
rect 44204 11102 44233 11676
rect 44279 11102 44308 11676
rect 44204 11089 44308 11102
rect 44364 11676 44468 11689
rect 44364 11102 44393 11676
rect 44439 11102 44468 11676
rect 44364 11089 44468 11102
rect 44524 11676 44628 11689
rect 44524 11102 44553 11676
rect 44599 11102 44628 11676
rect 44524 11089 44628 11102
rect 44684 11676 44788 11689
rect 44684 11102 44713 11676
rect 44759 11102 44788 11676
rect 44684 11089 44788 11102
rect 44844 11676 44948 11689
rect 44844 11102 44873 11676
rect 44919 11102 44948 11676
rect 44844 11089 44948 11102
rect 45004 11676 45108 11689
rect 45004 11102 45033 11676
rect 45079 11102 45108 11676
rect 45004 11089 45108 11102
rect 45164 11676 45268 11689
rect 45164 11102 45193 11676
rect 45239 11102 45268 11676
rect 45164 11089 45268 11102
rect 45324 11676 45428 11689
rect 45324 11102 45353 11676
rect 45399 11102 45428 11676
rect 45324 11089 45428 11102
rect 45484 11676 45588 11689
rect 45484 11102 45513 11676
rect 45559 11102 45588 11676
rect 45484 11089 45588 11102
rect 45644 11676 45732 11689
rect 45644 11102 45673 11676
rect 45719 11102 45732 11676
rect 45644 11089 45732 11102
rect 45788 11676 45876 11689
rect 45788 11102 45801 11676
rect 45847 11102 45876 11676
rect 45788 11089 45876 11102
rect 45932 11676 46020 11689
rect 45932 11102 45961 11676
rect 46007 11102 46020 11676
rect 45932 11089 46020 11102
rect 46948 11676 47036 11689
rect 46948 11102 46961 11676
rect 47007 11102 47036 11676
rect 46948 11089 47036 11102
rect 47092 11676 47180 11689
rect 47092 11102 47121 11676
rect 47167 11102 47180 11676
rect 47092 11089 47180 11102
rect 47236 11676 47324 11689
rect 47236 11102 47249 11676
rect 47295 11102 47324 11676
rect 47236 11089 47324 11102
rect 47380 11676 47484 11689
rect 47380 11102 47409 11676
rect 47455 11102 47484 11676
rect 47380 11089 47484 11102
rect 47540 11676 47644 11689
rect 47540 11102 47569 11676
rect 47615 11102 47644 11676
rect 47540 11089 47644 11102
rect 47700 11676 47804 11689
rect 47700 11102 47729 11676
rect 47775 11102 47804 11676
rect 47700 11089 47804 11102
rect 47860 11676 47964 11689
rect 47860 11102 47889 11676
rect 47935 11102 47964 11676
rect 47860 11089 47964 11102
rect 48020 11676 48124 11689
rect 48020 11102 48049 11676
rect 48095 11102 48124 11676
rect 48020 11089 48124 11102
rect 48180 11676 48284 11689
rect 48180 11102 48209 11676
rect 48255 11102 48284 11676
rect 48180 11089 48284 11102
rect 48340 11676 48444 11689
rect 48340 11102 48369 11676
rect 48415 11102 48444 11676
rect 48340 11089 48444 11102
rect 48500 11676 48604 11689
rect 48500 11102 48529 11676
rect 48575 11102 48604 11676
rect 48500 11089 48604 11102
rect 48660 11676 48764 11689
rect 48660 11102 48689 11676
rect 48735 11102 48764 11676
rect 48660 11089 48764 11102
rect 48820 11676 48924 11689
rect 48820 11102 48849 11676
rect 48895 11102 48924 11676
rect 48820 11089 48924 11102
rect 48980 11676 49084 11689
rect 48980 11102 49009 11676
rect 49055 11102 49084 11676
rect 48980 11089 49084 11102
rect 49140 11676 49244 11689
rect 49140 11102 49169 11676
rect 49215 11102 49244 11676
rect 49140 11089 49244 11102
rect 49300 11676 49404 11689
rect 49300 11102 49329 11676
rect 49375 11102 49404 11676
rect 49300 11089 49404 11102
rect 49460 11676 49564 11689
rect 49460 11102 49489 11676
rect 49535 11102 49564 11676
rect 49460 11089 49564 11102
rect 49620 11676 49724 11689
rect 49620 11102 49649 11676
rect 49695 11102 49724 11676
rect 49620 11089 49724 11102
rect 49780 11676 49868 11689
rect 49780 11102 49809 11676
rect 49855 11102 49868 11676
rect 49780 11089 49868 11102
rect 49924 11676 50012 11689
rect 49924 11102 49937 11676
rect 49983 11102 50012 11676
rect 49924 11089 50012 11102
rect 50068 11676 50156 11689
rect 50068 11102 50097 11676
rect 50143 11102 50156 11676
rect 50068 11089 50156 11102
rect 42812 10616 42900 10629
rect 42812 10042 42825 10616
rect 42871 10042 42900 10616
rect 42812 10029 42900 10042
rect 42956 10616 43044 10629
rect 42956 10042 42985 10616
rect 43031 10042 43044 10616
rect 42956 10029 43044 10042
rect 43100 10616 43188 10629
rect 43100 10042 43113 10616
rect 43159 10042 43188 10616
rect 43100 10029 43188 10042
rect 43244 10616 43348 10629
rect 43244 10042 43273 10616
rect 43319 10042 43348 10616
rect 43244 10029 43348 10042
rect 43404 10616 43508 10629
rect 43404 10042 43433 10616
rect 43479 10042 43508 10616
rect 43404 10029 43508 10042
rect 43564 10616 43668 10629
rect 43564 10042 43593 10616
rect 43639 10042 43668 10616
rect 43564 10029 43668 10042
rect 43724 10616 43828 10629
rect 43724 10042 43753 10616
rect 43799 10042 43828 10616
rect 43724 10029 43828 10042
rect 43884 10616 43988 10629
rect 43884 10042 43913 10616
rect 43959 10042 43988 10616
rect 43884 10029 43988 10042
rect 44044 10616 44148 10629
rect 44044 10042 44073 10616
rect 44119 10042 44148 10616
rect 44044 10029 44148 10042
rect 44204 10616 44308 10629
rect 44204 10042 44233 10616
rect 44279 10042 44308 10616
rect 44204 10029 44308 10042
rect 44364 10616 44468 10629
rect 44364 10042 44393 10616
rect 44439 10042 44468 10616
rect 44364 10029 44468 10042
rect 44524 10616 44628 10629
rect 44524 10042 44553 10616
rect 44599 10042 44628 10616
rect 44524 10029 44628 10042
rect 44684 10616 44788 10629
rect 44684 10042 44713 10616
rect 44759 10042 44788 10616
rect 44684 10029 44788 10042
rect 44844 10616 44948 10629
rect 44844 10042 44873 10616
rect 44919 10042 44948 10616
rect 44844 10029 44948 10042
rect 45004 10616 45108 10629
rect 45004 10042 45033 10616
rect 45079 10042 45108 10616
rect 45004 10029 45108 10042
rect 45164 10616 45268 10629
rect 45164 10042 45193 10616
rect 45239 10042 45268 10616
rect 45164 10029 45268 10042
rect 45324 10616 45428 10629
rect 45324 10042 45353 10616
rect 45399 10042 45428 10616
rect 45324 10029 45428 10042
rect 45484 10616 45588 10629
rect 45484 10042 45513 10616
rect 45559 10042 45588 10616
rect 45484 10029 45588 10042
rect 45644 10616 45732 10629
rect 45644 10042 45673 10616
rect 45719 10042 45732 10616
rect 45644 10029 45732 10042
rect 45788 10616 45876 10629
rect 45788 10042 45801 10616
rect 45847 10042 45876 10616
rect 45788 10029 45876 10042
rect 45932 10616 46020 10629
rect 45932 10042 45961 10616
rect 46007 10042 46020 10616
rect 45932 10029 46020 10042
rect 46948 10616 47036 10629
rect 46948 10042 46961 10616
rect 47007 10042 47036 10616
rect 46948 10029 47036 10042
rect 47092 10616 47180 10629
rect 47092 10042 47121 10616
rect 47167 10042 47180 10616
rect 47092 10029 47180 10042
rect 47236 10616 47324 10629
rect 47236 10042 47249 10616
rect 47295 10042 47324 10616
rect 47236 10029 47324 10042
rect 47380 10616 47484 10629
rect 47380 10042 47409 10616
rect 47455 10042 47484 10616
rect 47380 10029 47484 10042
rect 47540 10616 47644 10629
rect 47540 10042 47569 10616
rect 47615 10042 47644 10616
rect 47540 10029 47644 10042
rect 47700 10616 47804 10629
rect 47700 10042 47729 10616
rect 47775 10042 47804 10616
rect 47700 10029 47804 10042
rect 47860 10616 47964 10629
rect 47860 10042 47889 10616
rect 47935 10042 47964 10616
rect 47860 10029 47964 10042
rect 48020 10616 48124 10629
rect 48020 10042 48049 10616
rect 48095 10042 48124 10616
rect 48020 10029 48124 10042
rect 48180 10616 48284 10629
rect 48180 10042 48209 10616
rect 48255 10042 48284 10616
rect 48180 10029 48284 10042
rect 48340 10616 48444 10629
rect 48340 10042 48369 10616
rect 48415 10042 48444 10616
rect 48340 10029 48444 10042
rect 48500 10616 48604 10629
rect 48500 10042 48529 10616
rect 48575 10042 48604 10616
rect 48500 10029 48604 10042
rect 48660 10616 48764 10629
rect 48660 10042 48689 10616
rect 48735 10042 48764 10616
rect 48660 10029 48764 10042
rect 48820 10616 48924 10629
rect 48820 10042 48849 10616
rect 48895 10042 48924 10616
rect 48820 10029 48924 10042
rect 48980 10616 49084 10629
rect 48980 10042 49009 10616
rect 49055 10042 49084 10616
rect 48980 10029 49084 10042
rect 49140 10616 49244 10629
rect 49140 10042 49169 10616
rect 49215 10042 49244 10616
rect 49140 10029 49244 10042
rect 49300 10616 49404 10629
rect 49300 10042 49329 10616
rect 49375 10042 49404 10616
rect 49300 10029 49404 10042
rect 49460 10616 49564 10629
rect 49460 10042 49489 10616
rect 49535 10042 49564 10616
rect 49460 10029 49564 10042
rect 49620 10616 49724 10629
rect 49620 10042 49649 10616
rect 49695 10042 49724 10616
rect 49620 10029 49724 10042
rect 49780 10616 49868 10629
rect 49780 10042 49809 10616
rect 49855 10042 49868 10616
rect 49780 10029 49868 10042
rect 49924 10616 50012 10629
rect 49924 10042 49937 10616
rect 49983 10042 50012 10616
rect 49924 10029 50012 10042
rect 50068 10616 50156 10629
rect 50068 10042 50097 10616
rect 50143 10042 50156 10616
rect 50068 10029 50156 10042
rect 42812 9556 42900 9569
rect 42812 8982 42825 9556
rect 42871 8982 42900 9556
rect 42812 8969 42900 8982
rect 42956 9556 43044 9569
rect 42956 8982 42985 9556
rect 43031 8982 43044 9556
rect 42956 8969 43044 8982
rect 43100 9556 43188 9569
rect 43100 8982 43113 9556
rect 43159 8982 43188 9556
rect 43100 8969 43188 8982
rect 43244 9556 43348 9569
rect 43244 8982 43273 9556
rect 43319 8982 43348 9556
rect 43244 8969 43348 8982
rect 43404 9556 43508 9569
rect 43404 8982 43433 9556
rect 43479 8982 43508 9556
rect 43404 8969 43508 8982
rect 43564 9556 43668 9569
rect 43564 8982 43593 9556
rect 43639 8982 43668 9556
rect 43564 8969 43668 8982
rect 43724 9556 43828 9569
rect 43724 8982 43753 9556
rect 43799 8982 43828 9556
rect 43724 8969 43828 8982
rect 43884 9556 43988 9569
rect 43884 8982 43913 9556
rect 43959 8982 43988 9556
rect 43884 8969 43988 8982
rect 44044 9556 44148 9569
rect 44044 8982 44073 9556
rect 44119 8982 44148 9556
rect 44044 8969 44148 8982
rect 44204 9556 44308 9569
rect 44204 8982 44233 9556
rect 44279 8982 44308 9556
rect 44204 8969 44308 8982
rect 44364 9556 44468 9569
rect 44364 8982 44393 9556
rect 44439 8982 44468 9556
rect 44364 8969 44468 8982
rect 44524 9556 44628 9569
rect 44524 8982 44553 9556
rect 44599 8982 44628 9556
rect 44524 8969 44628 8982
rect 44684 9556 44788 9569
rect 44684 8982 44713 9556
rect 44759 8982 44788 9556
rect 44684 8969 44788 8982
rect 44844 9556 44948 9569
rect 44844 8982 44873 9556
rect 44919 8982 44948 9556
rect 44844 8969 44948 8982
rect 45004 9556 45108 9569
rect 45004 8982 45033 9556
rect 45079 8982 45108 9556
rect 45004 8969 45108 8982
rect 45164 9556 45268 9569
rect 45164 8982 45193 9556
rect 45239 8982 45268 9556
rect 45164 8969 45268 8982
rect 45324 9556 45428 9569
rect 45324 8982 45353 9556
rect 45399 8982 45428 9556
rect 45324 8969 45428 8982
rect 45484 9556 45588 9569
rect 45484 8982 45513 9556
rect 45559 8982 45588 9556
rect 45484 8969 45588 8982
rect 45644 9556 45732 9569
rect 45644 8982 45673 9556
rect 45719 8982 45732 9556
rect 45644 8969 45732 8982
rect 45788 9556 45876 9569
rect 45788 8982 45801 9556
rect 45847 8982 45876 9556
rect 45788 8969 45876 8982
rect 45932 9556 46020 9569
rect 45932 8982 45961 9556
rect 46007 8982 46020 9556
rect 45932 8969 46020 8982
rect 46948 9556 47036 9569
rect 46948 8982 46961 9556
rect 47007 8982 47036 9556
rect 46948 8969 47036 8982
rect 47092 9556 47180 9569
rect 47092 8982 47121 9556
rect 47167 8982 47180 9556
rect 47092 8969 47180 8982
rect 47236 9556 47324 9569
rect 47236 8982 47249 9556
rect 47295 8982 47324 9556
rect 47236 8969 47324 8982
rect 47380 9556 47484 9569
rect 47380 8982 47409 9556
rect 47455 8982 47484 9556
rect 47380 8969 47484 8982
rect 47540 9556 47644 9569
rect 47540 8982 47569 9556
rect 47615 8982 47644 9556
rect 47540 8969 47644 8982
rect 47700 9556 47804 9569
rect 47700 8982 47729 9556
rect 47775 8982 47804 9556
rect 47700 8969 47804 8982
rect 47860 9556 47964 9569
rect 47860 8982 47889 9556
rect 47935 8982 47964 9556
rect 47860 8969 47964 8982
rect 48020 9556 48124 9569
rect 48020 8982 48049 9556
rect 48095 8982 48124 9556
rect 48020 8969 48124 8982
rect 48180 9556 48284 9569
rect 48180 8982 48209 9556
rect 48255 8982 48284 9556
rect 48180 8969 48284 8982
rect 48340 9556 48444 9569
rect 48340 8982 48369 9556
rect 48415 8982 48444 9556
rect 48340 8969 48444 8982
rect 48500 9556 48604 9569
rect 48500 8982 48529 9556
rect 48575 8982 48604 9556
rect 48500 8969 48604 8982
rect 48660 9556 48764 9569
rect 48660 8982 48689 9556
rect 48735 8982 48764 9556
rect 48660 8969 48764 8982
rect 48820 9556 48924 9569
rect 48820 8982 48849 9556
rect 48895 8982 48924 9556
rect 48820 8969 48924 8982
rect 48980 9556 49084 9569
rect 48980 8982 49009 9556
rect 49055 8982 49084 9556
rect 48980 8969 49084 8982
rect 49140 9556 49244 9569
rect 49140 8982 49169 9556
rect 49215 8982 49244 9556
rect 49140 8969 49244 8982
rect 49300 9556 49404 9569
rect 49300 8982 49329 9556
rect 49375 8982 49404 9556
rect 49300 8969 49404 8982
rect 49460 9556 49564 9569
rect 49460 8982 49489 9556
rect 49535 8982 49564 9556
rect 49460 8969 49564 8982
rect 49620 9556 49724 9569
rect 49620 8982 49649 9556
rect 49695 8982 49724 9556
rect 49620 8969 49724 8982
rect 49780 9556 49868 9569
rect 49780 8982 49809 9556
rect 49855 8982 49868 9556
rect 49780 8969 49868 8982
rect 49924 9556 50012 9569
rect 49924 8982 49937 9556
rect 49983 8982 50012 9556
rect 49924 8969 50012 8982
rect 50068 9556 50156 9569
rect 50068 8982 50097 9556
rect 50143 8982 50156 9556
rect 50068 8969 50156 8982
rect 42812 8496 42900 8509
rect 42812 7922 42825 8496
rect 42871 7922 42900 8496
rect 42812 7909 42900 7922
rect 42956 8496 43044 8509
rect 42956 7922 42985 8496
rect 43031 7922 43044 8496
rect 42956 7909 43044 7922
rect 43100 8496 43188 8509
rect 43100 7922 43113 8496
rect 43159 7922 43188 8496
rect 43100 7909 43188 7922
rect 43244 8496 43348 8509
rect 43244 7922 43273 8496
rect 43319 7922 43348 8496
rect 43244 7909 43348 7922
rect 43404 8496 43508 8509
rect 43404 7922 43433 8496
rect 43479 7922 43508 8496
rect 43404 7909 43508 7922
rect 43564 8496 43668 8509
rect 43564 7922 43593 8496
rect 43639 7922 43668 8496
rect 43564 7909 43668 7922
rect 43724 8496 43828 8509
rect 43724 7922 43753 8496
rect 43799 7922 43828 8496
rect 43724 7909 43828 7922
rect 43884 8496 43988 8509
rect 43884 7922 43913 8496
rect 43959 7922 43988 8496
rect 43884 7909 43988 7922
rect 44044 8496 44148 8509
rect 44044 7922 44073 8496
rect 44119 7922 44148 8496
rect 44044 7909 44148 7922
rect 44204 8496 44308 8509
rect 44204 7922 44233 8496
rect 44279 7922 44308 8496
rect 44204 7909 44308 7922
rect 44364 8496 44468 8509
rect 44364 7922 44393 8496
rect 44439 7922 44468 8496
rect 44364 7909 44468 7922
rect 44524 8496 44628 8509
rect 44524 7922 44553 8496
rect 44599 7922 44628 8496
rect 44524 7909 44628 7922
rect 44684 8496 44788 8509
rect 44684 7922 44713 8496
rect 44759 7922 44788 8496
rect 44684 7909 44788 7922
rect 44844 8496 44948 8509
rect 44844 7922 44873 8496
rect 44919 7922 44948 8496
rect 44844 7909 44948 7922
rect 45004 8496 45108 8509
rect 45004 7922 45033 8496
rect 45079 7922 45108 8496
rect 45004 7909 45108 7922
rect 45164 8496 45268 8509
rect 45164 7922 45193 8496
rect 45239 7922 45268 8496
rect 45164 7909 45268 7922
rect 45324 8496 45428 8509
rect 45324 7922 45353 8496
rect 45399 7922 45428 8496
rect 45324 7909 45428 7922
rect 45484 8496 45588 8509
rect 45484 7922 45513 8496
rect 45559 7922 45588 8496
rect 45484 7909 45588 7922
rect 45644 8496 45732 8509
rect 45644 7922 45673 8496
rect 45719 7922 45732 8496
rect 45644 7909 45732 7922
rect 45788 8496 45876 8509
rect 45788 7922 45801 8496
rect 45847 7922 45876 8496
rect 45788 7909 45876 7922
rect 45932 8496 46020 8509
rect 45932 7922 45961 8496
rect 46007 7922 46020 8496
rect 45932 7909 46020 7922
rect 46948 8496 47036 8509
rect 46948 7922 46961 8496
rect 47007 7922 47036 8496
rect 46948 7909 47036 7922
rect 47092 8496 47180 8509
rect 47092 7922 47121 8496
rect 47167 7922 47180 8496
rect 47092 7909 47180 7922
rect 47236 8496 47324 8509
rect 47236 7922 47249 8496
rect 47295 7922 47324 8496
rect 47236 7909 47324 7922
rect 47380 8496 47484 8509
rect 47380 7922 47409 8496
rect 47455 7922 47484 8496
rect 47380 7909 47484 7922
rect 47540 8496 47644 8509
rect 47540 7922 47569 8496
rect 47615 7922 47644 8496
rect 47540 7909 47644 7922
rect 47700 8496 47804 8509
rect 47700 7922 47729 8496
rect 47775 7922 47804 8496
rect 47700 7909 47804 7922
rect 47860 8496 47964 8509
rect 47860 7922 47889 8496
rect 47935 7922 47964 8496
rect 47860 7909 47964 7922
rect 48020 8496 48124 8509
rect 48020 7922 48049 8496
rect 48095 7922 48124 8496
rect 48020 7909 48124 7922
rect 48180 8496 48284 8509
rect 48180 7922 48209 8496
rect 48255 7922 48284 8496
rect 48180 7909 48284 7922
rect 48340 8496 48444 8509
rect 48340 7922 48369 8496
rect 48415 7922 48444 8496
rect 48340 7909 48444 7922
rect 48500 8496 48604 8509
rect 48500 7922 48529 8496
rect 48575 7922 48604 8496
rect 48500 7909 48604 7922
rect 48660 8496 48764 8509
rect 48660 7922 48689 8496
rect 48735 7922 48764 8496
rect 48660 7909 48764 7922
rect 48820 8496 48924 8509
rect 48820 7922 48849 8496
rect 48895 7922 48924 8496
rect 48820 7909 48924 7922
rect 48980 8496 49084 8509
rect 48980 7922 49009 8496
rect 49055 7922 49084 8496
rect 48980 7909 49084 7922
rect 49140 8496 49244 8509
rect 49140 7922 49169 8496
rect 49215 7922 49244 8496
rect 49140 7909 49244 7922
rect 49300 8496 49404 8509
rect 49300 7922 49329 8496
rect 49375 7922 49404 8496
rect 49300 7909 49404 7922
rect 49460 8496 49564 8509
rect 49460 7922 49489 8496
rect 49535 7922 49564 8496
rect 49460 7909 49564 7922
rect 49620 8496 49724 8509
rect 49620 7922 49649 8496
rect 49695 7922 49724 8496
rect 49620 7909 49724 7922
rect 49780 8496 49868 8509
rect 49780 7922 49809 8496
rect 49855 7922 49868 8496
rect 49780 7909 49868 7922
rect 49924 8496 50012 8509
rect 49924 7922 49937 8496
rect 49983 7922 50012 8496
rect 49924 7909 50012 7922
rect 50068 8496 50156 8509
rect 50068 7922 50097 8496
rect 50143 7922 50156 8496
rect 50068 7909 50156 7922
rect 52508 11676 52596 11689
rect 52508 11102 52521 11676
rect 52567 11102 52596 11676
rect 52508 11089 52596 11102
rect 52652 11676 52740 11689
rect 52652 11102 52681 11676
rect 52727 11102 52740 11676
rect 52652 11089 52740 11102
rect 52796 11676 52884 11689
rect 52796 11102 52809 11676
rect 52855 11102 52884 11676
rect 52796 11089 52884 11102
rect 52940 11676 53044 11689
rect 52940 11102 52969 11676
rect 53015 11102 53044 11676
rect 52940 11089 53044 11102
rect 53100 11676 53204 11689
rect 53100 11102 53129 11676
rect 53175 11102 53204 11676
rect 53100 11089 53204 11102
rect 53260 11676 53364 11689
rect 53260 11102 53289 11676
rect 53335 11102 53364 11676
rect 53260 11089 53364 11102
rect 53420 11676 53524 11689
rect 53420 11102 53449 11676
rect 53495 11102 53524 11676
rect 53420 11089 53524 11102
rect 53580 11676 53684 11689
rect 53580 11102 53609 11676
rect 53655 11102 53684 11676
rect 53580 11089 53684 11102
rect 53740 11676 53844 11689
rect 53740 11102 53769 11676
rect 53815 11102 53844 11676
rect 53740 11089 53844 11102
rect 53900 11676 54004 11689
rect 53900 11102 53929 11676
rect 53975 11102 54004 11676
rect 53900 11089 54004 11102
rect 54060 11676 54164 11689
rect 54060 11102 54089 11676
rect 54135 11102 54164 11676
rect 54060 11089 54164 11102
rect 54220 11676 54324 11689
rect 54220 11102 54249 11676
rect 54295 11102 54324 11676
rect 54220 11089 54324 11102
rect 54380 11676 54484 11689
rect 54380 11102 54409 11676
rect 54455 11102 54484 11676
rect 54380 11089 54484 11102
rect 54540 11676 54644 11689
rect 54540 11102 54569 11676
rect 54615 11102 54644 11676
rect 54540 11089 54644 11102
rect 54700 11676 54804 11689
rect 54700 11102 54729 11676
rect 54775 11102 54804 11676
rect 54700 11089 54804 11102
rect 54860 11676 54964 11689
rect 54860 11102 54889 11676
rect 54935 11102 54964 11676
rect 54860 11089 54964 11102
rect 55020 11676 55124 11689
rect 55020 11102 55049 11676
rect 55095 11102 55124 11676
rect 55020 11089 55124 11102
rect 55180 11676 55284 11689
rect 55180 11102 55209 11676
rect 55255 11102 55284 11676
rect 55180 11089 55284 11102
rect 55340 11676 55428 11689
rect 55340 11102 55369 11676
rect 55415 11102 55428 11676
rect 55340 11089 55428 11102
rect 55484 11676 55572 11689
rect 55484 11102 55497 11676
rect 55543 11102 55572 11676
rect 55484 11089 55572 11102
rect 55628 11676 55716 11689
rect 55628 11102 55657 11676
rect 55703 11102 55716 11676
rect 55628 11089 55716 11102
rect 56644 11676 56732 11689
rect 56644 11102 56657 11676
rect 56703 11102 56732 11676
rect 56644 11089 56732 11102
rect 56788 11676 56876 11689
rect 56788 11102 56817 11676
rect 56863 11102 56876 11676
rect 56788 11089 56876 11102
rect 56932 11676 57020 11689
rect 56932 11102 56945 11676
rect 56991 11102 57020 11676
rect 56932 11089 57020 11102
rect 57076 11676 57180 11689
rect 57076 11102 57105 11676
rect 57151 11102 57180 11676
rect 57076 11089 57180 11102
rect 57236 11676 57340 11689
rect 57236 11102 57265 11676
rect 57311 11102 57340 11676
rect 57236 11089 57340 11102
rect 57396 11676 57500 11689
rect 57396 11102 57425 11676
rect 57471 11102 57500 11676
rect 57396 11089 57500 11102
rect 57556 11676 57660 11689
rect 57556 11102 57585 11676
rect 57631 11102 57660 11676
rect 57556 11089 57660 11102
rect 57716 11676 57820 11689
rect 57716 11102 57745 11676
rect 57791 11102 57820 11676
rect 57716 11089 57820 11102
rect 57876 11676 57980 11689
rect 57876 11102 57905 11676
rect 57951 11102 57980 11676
rect 57876 11089 57980 11102
rect 58036 11676 58140 11689
rect 58036 11102 58065 11676
rect 58111 11102 58140 11676
rect 58036 11089 58140 11102
rect 58196 11676 58300 11689
rect 58196 11102 58225 11676
rect 58271 11102 58300 11676
rect 58196 11089 58300 11102
rect 58356 11676 58460 11689
rect 58356 11102 58385 11676
rect 58431 11102 58460 11676
rect 58356 11089 58460 11102
rect 58516 11676 58620 11689
rect 58516 11102 58545 11676
rect 58591 11102 58620 11676
rect 58516 11089 58620 11102
rect 58676 11676 58780 11689
rect 58676 11102 58705 11676
rect 58751 11102 58780 11676
rect 58676 11089 58780 11102
rect 58836 11676 58940 11689
rect 58836 11102 58865 11676
rect 58911 11102 58940 11676
rect 58836 11089 58940 11102
rect 58996 11676 59100 11689
rect 58996 11102 59025 11676
rect 59071 11102 59100 11676
rect 58996 11089 59100 11102
rect 59156 11676 59260 11689
rect 59156 11102 59185 11676
rect 59231 11102 59260 11676
rect 59156 11089 59260 11102
rect 59316 11676 59420 11689
rect 59316 11102 59345 11676
rect 59391 11102 59420 11676
rect 59316 11089 59420 11102
rect 59476 11676 59564 11689
rect 59476 11102 59505 11676
rect 59551 11102 59564 11676
rect 59476 11089 59564 11102
rect 59620 11676 59708 11689
rect 59620 11102 59633 11676
rect 59679 11102 59708 11676
rect 59620 11089 59708 11102
rect 59764 11676 59852 11689
rect 59764 11102 59793 11676
rect 59839 11102 59852 11676
rect 59764 11089 59852 11102
rect 52508 10616 52596 10629
rect 52508 10042 52521 10616
rect 52567 10042 52596 10616
rect 52508 10029 52596 10042
rect 52652 10616 52740 10629
rect 52652 10042 52681 10616
rect 52727 10042 52740 10616
rect 52652 10029 52740 10042
rect 52796 10616 52884 10629
rect 52796 10042 52809 10616
rect 52855 10042 52884 10616
rect 52796 10029 52884 10042
rect 52940 10616 53044 10629
rect 52940 10042 52969 10616
rect 53015 10042 53044 10616
rect 52940 10029 53044 10042
rect 53100 10616 53204 10629
rect 53100 10042 53129 10616
rect 53175 10042 53204 10616
rect 53100 10029 53204 10042
rect 53260 10616 53364 10629
rect 53260 10042 53289 10616
rect 53335 10042 53364 10616
rect 53260 10029 53364 10042
rect 53420 10616 53524 10629
rect 53420 10042 53449 10616
rect 53495 10042 53524 10616
rect 53420 10029 53524 10042
rect 53580 10616 53684 10629
rect 53580 10042 53609 10616
rect 53655 10042 53684 10616
rect 53580 10029 53684 10042
rect 53740 10616 53844 10629
rect 53740 10042 53769 10616
rect 53815 10042 53844 10616
rect 53740 10029 53844 10042
rect 53900 10616 54004 10629
rect 53900 10042 53929 10616
rect 53975 10042 54004 10616
rect 53900 10029 54004 10042
rect 54060 10616 54164 10629
rect 54060 10042 54089 10616
rect 54135 10042 54164 10616
rect 54060 10029 54164 10042
rect 54220 10616 54324 10629
rect 54220 10042 54249 10616
rect 54295 10042 54324 10616
rect 54220 10029 54324 10042
rect 54380 10616 54484 10629
rect 54380 10042 54409 10616
rect 54455 10042 54484 10616
rect 54380 10029 54484 10042
rect 54540 10616 54644 10629
rect 54540 10042 54569 10616
rect 54615 10042 54644 10616
rect 54540 10029 54644 10042
rect 54700 10616 54804 10629
rect 54700 10042 54729 10616
rect 54775 10042 54804 10616
rect 54700 10029 54804 10042
rect 54860 10616 54964 10629
rect 54860 10042 54889 10616
rect 54935 10042 54964 10616
rect 54860 10029 54964 10042
rect 55020 10616 55124 10629
rect 55020 10042 55049 10616
rect 55095 10042 55124 10616
rect 55020 10029 55124 10042
rect 55180 10616 55284 10629
rect 55180 10042 55209 10616
rect 55255 10042 55284 10616
rect 55180 10029 55284 10042
rect 55340 10616 55428 10629
rect 55340 10042 55369 10616
rect 55415 10042 55428 10616
rect 55340 10029 55428 10042
rect 55484 10616 55572 10629
rect 55484 10042 55497 10616
rect 55543 10042 55572 10616
rect 55484 10029 55572 10042
rect 55628 10616 55716 10629
rect 55628 10042 55657 10616
rect 55703 10042 55716 10616
rect 55628 10029 55716 10042
rect 56644 10616 56732 10629
rect 56644 10042 56657 10616
rect 56703 10042 56732 10616
rect 56644 10029 56732 10042
rect 56788 10616 56876 10629
rect 56788 10042 56817 10616
rect 56863 10042 56876 10616
rect 56788 10029 56876 10042
rect 56932 10616 57020 10629
rect 56932 10042 56945 10616
rect 56991 10042 57020 10616
rect 56932 10029 57020 10042
rect 57076 10616 57180 10629
rect 57076 10042 57105 10616
rect 57151 10042 57180 10616
rect 57076 10029 57180 10042
rect 57236 10616 57340 10629
rect 57236 10042 57265 10616
rect 57311 10042 57340 10616
rect 57236 10029 57340 10042
rect 57396 10616 57500 10629
rect 57396 10042 57425 10616
rect 57471 10042 57500 10616
rect 57396 10029 57500 10042
rect 57556 10616 57660 10629
rect 57556 10042 57585 10616
rect 57631 10042 57660 10616
rect 57556 10029 57660 10042
rect 57716 10616 57820 10629
rect 57716 10042 57745 10616
rect 57791 10042 57820 10616
rect 57716 10029 57820 10042
rect 57876 10616 57980 10629
rect 57876 10042 57905 10616
rect 57951 10042 57980 10616
rect 57876 10029 57980 10042
rect 58036 10616 58140 10629
rect 58036 10042 58065 10616
rect 58111 10042 58140 10616
rect 58036 10029 58140 10042
rect 58196 10616 58300 10629
rect 58196 10042 58225 10616
rect 58271 10042 58300 10616
rect 58196 10029 58300 10042
rect 58356 10616 58460 10629
rect 58356 10042 58385 10616
rect 58431 10042 58460 10616
rect 58356 10029 58460 10042
rect 58516 10616 58620 10629
rect 58516 10042 58545 10616
rect 58591 10042 58620 10616
rect 58516 10029 58620 10042
rect 58676 10616 58780 10629
rect 58676 10042 58705 10616
rect 58751 10042 58780 10616
rect 58676 10029 58780 10042
rect 58836 10616 58940 10629
rect 58836 10042 58865 10616
rect 58911 10042 58940 10616
rect 58836 10029 58940 10042
rect 58996 10616 59100 10629
rect 58996 10042 59025 10616
rect 59071 10042 59100 10616
rect 58996 10029 59100 10042
rect 59156 10616 59260 10629
rect 59156 10042 59185 10616
rect 59231 10042 59260 10616
rect 59156 10029 59260 10042
rect 59316 10616 59420 10629
rect 59316 10042 59345 10616
rect 59391 10042 59420 10616
rect 59316 10029 59420 10042
rect 59476 10616 59564 10629
rect 59476 10042 59505 10616
rect 59551 10042 59564 10616
rect 59476 10029 59564 10042
rect 59620 10616 59708 10629
rect 59620 10042 59633 10616
rect 59679 10042 59708 10616
rect 59620 10029 59708 10042
rect 59764 10616 59852 10629
rect 59764 10042 59793 10616
rect 59839 10042 59852 10616
rect 59764 10029 59852 10042
rect 52508 9556 52596 9569
rect 52508 8982 52521 9556
rect 52567 8982 52596 9556
rect 52508 8969 52596 8982
rect 52652 9556 52740 9569
rect 52652 8982 52681 9556
rect 52727 8982 52740 9556
rect 52652 8969 52740 8982
rect 52796 9556 52884 9569
rect 52796 8982 52809 9556
rect 52855 8982 52884 9556
rect 52796 8969 52884 8982
rect 52940 9556 53044 9569
rect 52940 8982 52969 9556
rect 53015 8982 53044 9556
rect 52940 8969 53044 8982
rect 53100 9556 53204 9569
rect 53100 8982 53129 9556
rect 53175 8982 53204 9556
rect 53100 8969 53204 8982
rect 53260 9556 53364 9569
rect 53260 8982 53289 9556
rect 53335 8982 53364 9556
rect 53260 8969 53364 8982
rect 53420 9556 53524 9569
rect 53420 8982 53449 9556
rect 53495 8982 53524 9556
rect 53420 8969 53524 8982
rect 53580 9556 53684 9569
rect 53580 8982 53609 9556
rect 53655 8982 53684 9556
rect 53580 8969 53684 8982
rect 53740 9556 53844 9569
rect 53740 8982 53769 9556
rect 53815 8982 53844 9556
rect 53740 8969 53844 8982
rect 53900 9556 54004 9569
rect 53900 8982 53929 9556
rect 53975 8982 54004 9556
rect 53900 8969 54004 8982
rect 54060 9556 54164 9569
rect 54060 8982 54089 9556
rect 54135 8982 54164 9556
rect 54060 8969 54164 8982
rect 54220 9556 54324 9569
rect 54220 8982 54249 9556
rect 54295 8982 54324 9556
rect 54220 8969 54324 8982
rect 54380 9556 54484 9569
rect 54380 8982 54409 9556
rect 54455 8982 54484 9556
rect 54380 8969 54484 8982
rect 54540 9556 54644 9569
rect 54540 8982 54569 9556
rect 54615 8982 54644 9556
rect 54540 8969 54644 8982
rect 54700 9556 54804 9569
rect 54700 8982 54729 9556
rect 54775 8982 54804 9556
rect 54700 8969 54804 8982
rect 54860 9556 54964 9569
rect 54860 8982 54889 9556
rect 54935 8982 54964 9556
rect 54860 8969 54964 8982
rect 55020 9556 55124 9569
rect 55020 8982 55049 9556
rect 55095 8982 55124 9556
rect 55020 8969 55124 8982
rect 55180 9556 55284 9569
rect 55180 8982 55209 9556
rect 55255 8982 55284 9556
rect 55180 8969 55284 8982
rect 55340 9556 55428 9569
rect 55340 8982 55369 9556
rect 55415 8982 55428 9556
rect 55340 8969 55428 8982
rect 55484 9556 55572 9569
rect 55484 8982 55497 9556
rect 55543 8982 55572 9556
rect 55484 8969 55572 8982
rect 55628 9556 55716 9569
rect 55628 8982 55657 9556
rect 55703 8982 55716 9556
rect 55628 8969 55716 8982
rect 56644 9556 56732 9569
rect 56644 8982 56657 9556
rect 56703 8982 56732 9556
rect 56644 8969 56732 8982
rect 56788 9556 56876 9569
rect 56788 8982 56817 9556
rect 56863 8982 56876 9556
rect 56788 8969 56876 8982
rect 56932 9556 57020 9569
rect 56932 8982 56945 9556
rect 56991 8982 57020 9556
rect 56932 8969 57020 8982
rect 57076 9556 57180 9569
rect 57076 8982 57105 9556
rect 57151 8982 57180 9556
rect 57076 8969 57180 8982
rect 57236 9556 57340 9569
rect 57236 8982 57265 9556
rect 57311 8982 57340 9556
rect 57236 8969 57340 8982
rect 57396 9556 57500 9569
rect 57396 8982 57425 9556
rect 57471 8982 57500 9556
rect 57396 8969 57500 8982
rect 57556 9556 57660 9569
rect 57556 8982 57585 9556
rect 57631 8982 57660 9556
rect 57556 8969 57660 8982
rect 57716 9556 57820 9569
rect 57716 8982 57745 9556
rect 57791 8982 57820 9556
rect 57716 8969 57820 8982
rect 57876 9556 57980 9569
rect 57876 8982 57905 9556
rect 57951 8982 57980 9556
rect 57876 8969 57980 8982
rect 58036 9556 58140 9569
rect 58036 8982 58065 9556
rect 58111 8982 58140 9556
rect 58036 8969 58140 8982
rect 58196 9556 58300 9569
rect 58196 8982 58225 9556
rect 58271 8982 58300 9556
rect 58196 8969 58300 8982
rect 58356 9556 58460 9569
rect 58356 8982 58385 9556
rect 58431 8982 58460 9556
rect 58356 8969 58460 8982
rect 58516 9556 58620 9569
rect 58516 8982 58545 9556
rect 58591 8982 58620 9556
rect 58516 8969 58620 8982
rect 58676 9556 58780 9569
rect 58676 8982 58705 9556
rect 58751 8982 58780 9556
rect 58676 8969 58780 8982
rect 58836 9556 58940 9569
rect 58836 8982 58865 9556
rect 58911 8982 58940 9556
rect 58836 8969 58940 8982
rect 58996 9556 59100 9569
rect 58996 8982 59025 9556
rect 59071 8982 59100 9556
rect 58996 8969 59100 8982
rect 59156 9556 59260 9569
rect 59156 8982 59185 9556
rect 59231 8982 59260 9556
rect 59156 8969 59260 8982
rect 59316 9556 59420 9569
rect 59316 8982 59345 9556
rect 59391 8982 59420 9556
rect 59316 8969 59420 8982
rect 59476 9556 59564 9569
rect 59476 8982 59505 9556
rect 59551 8982 59564 9556
rect 59476 8969 59564 8982
rect 59620 9556 59708 9569
rect 59620 8982 59633 9556
rect 59679 8982 59708 9556
rect 59620 8969 59708 8982
rect 59764 9556 59852 9569
rect 59764 8982 59793 9556
rect 59839 8982 59852 9556
rect 59764 8969 59852 8982
rect 52508 8496 52596 8509
rect 52508 7922 52521 8496
rect 52567 7922 52596 8496
rect 52508 7909 52596 7922
rect 52652 8496 52740 8509
rect 52652 7922 52681 8496
rect 52727 7922 52740 8496
rect 52652 7909 52740 7922
rect 52796 8496 52884 8509
rect 52796 7922 52809 8496
rect 52855 7922 52884 8496
rect 52796 7909 52884 7922
rect 52940 8496 53044 8509
rect 52940 7922 52969 8496
rect 53015 7922 53044 8496
rect 52940 7909 53044 7922
rect 53100 8496 53204 8509
rect 53100 7922 53129 8496
rect 53175 7922 53204 8496
rect 53100 7909 53204 7922
rect 53260 8496 53364 8509
rect 53260 7922 53289 8496
rect 53335 7922 53364 8496
rect 53260 7909 53364 7922
rect 53420 8496 53524 8509
rect 53420 7922 53449 8496
rect 53495 7922 53524 8496
rect 53420 7909 53524 7922
rect 53580 8496 53684 8509
rect 53580 7922 53609 8496
rect 53655 7922 53684 8496
rect 53580 7909 53684 7922
rect 53740 8496 53844 8509
rect 53740 7922 53769 8496
rect 53815 7922 53844 8496
rect 53740 7909 53844 7922
rect 53900 8496 54004 8509
rect 53900 7922 53929 8496
rect 53975 7922 54004 8496
rect 53900 7909 54004 7922
rect 54060 8496 54164 8509
rect 54060 7922 54089 8496
rect 54135 7922 54164 8496
rect 54060 7909 54164 7922
rect 54220 8496 54324 8509
rect 54220 7922 54249 8496
rect 54295 7922 54324 8496
rect 54220 7909 54324 7922
rect 54380 8496 54484 8509
rect 54380 7922 54409 8496
rect 54455 7922 54484 8496
rect 54380 7909 54484 7922
rect 54540 8496 54644 8509
rect 54540 7922 54569 8496
rect 54615 7922 54644 8496
rect 54540 7909 54644 7922
rect 54700 8496 54804 8509
rect 54700 7922 54729 8496
rect 54775 7922 54804 8496
rect 54700 7909 54804 7922
rect 54860 8496 54964 8509
rect 54860 7922 54889 8496
rect 54935 7922 54964 8496
rect 54860 7909 54964 7922
rect 55020 8496 55124 8509
rect 55020 7922 55049 8496
rect 55095 7922 55124 8496
rect 55020 7909 55124 7922
rect 55180 8496 55284 8509
rect 55180 7922 55209 8496
rect 55255 7922 55284 8496
rect 55180 7909 55284 7922
rect 55340 8496 55428 8509
rect 55340 7922 55369 8496
rect 55415 7922 55428 8496
rect 55340 7909 55428 7922
rect 55484 8496 55572 8509
rect 55484 7922 55497 8496
rect 55543 7922 55572 8496
rect 55484 7909 55572 7922
rect 55628 8496 55716 8509
rect 55628 7922 55657 8496
rect 55703 7922 55716 8496
rect 55628 7909 55716 7922
rect 56644 8496 56732 8509
rect 56644 7922 56657 8496
rect 56703 7922 56732 8496
rect 56644 7909 56732 7922
rect 56788 8496 56876 8509
rect 56788 7922 56817 8496
rect 56863 7922 56876 8496
rect 56788 7909 56876 7922
rect 56932 8496 57020 8509
rect 56932 7922 56945 8496
rect 56991 7922 57020 8496
rect 56932 7909 57020 7922
rect 57076 8496 57180 8509
rect 57076 7922 57105 8496
rect 57151 7922 57180 8496
rect 57076 7909 57180 7922
rect 57236 8496 57340 8509
rect 57236 7922 57265 8496
rect 57311 7922 57340 8496
rect 57236 7909 57340 7922
rect 57396 8496 57500 8509
rect 57396 7922 57425 8496
rect 57471 7922 57500 8496
rect 57396 7909 57500 7922
rect 57556 8496 57660 8509
rect 57556 7922 57585 8496
rect 57631 7922 57660 8496
rect 57556 7909 57660 7922
rect 57716 8496 57820 8509
rect 57716 7922 57745 8496
rect 57791 7922 57820 8496
rect 57716 7909 57820 7922
rect 57876 8496 57980 8509
rect 57876 7922 57905 8496
rect 57951 7922 57980 8496
rect 57876 7909 57980 7922
rect 58036 8496 58140 8509
rect 58036 7922 58065 8496
rect 58111 7922 58140 8496
rect 58036 7909 58140 7922
rect 58196 8496 58300 8509
rect 58196 7922 58225 8496
rect 58271 7922 58300 8496
rect 58196 7909 58300 7922
rect 58356 8496 58460 8509
rect 58356 7922 58385 8496
rect 58431 7922 58460 8496
rect 58356 7909 58460 7922
rect 58516 8496 58620 8509
rect 58516 7922 58545 8496
rect 58591 7922 58620 8496
rect 58516 7909 58620 7922
rect 58676 8496 58780 8509
rect 58676 7922 58705 8496
rect 58751 7922 58780 8496
rect 58676 7909 58780 7922
rect 58836 8496 58940 8509
rect 58836 7922 58865 8496
rect 58911 7922 58940 8496
rect 58836 7909 58940 7922
rect 58996 8496 59100 8509
rect 58996 7922 59025 8496
rect 59071 7922 59100 8496
rect 58996 7909 59100 7922
rect 59156 8496 59260 8509
rect 59156 7922 59185 8496
rect 59231 7922 59260 8496
rect 59156 7909 59260 7922
rect 59316 8496 59420 8509
rect 59316 7922 59345 8496
rect 59391 7922 59420 8496
rect 59316 7909 59420 7922
rect 59476 8496 59564 8509
rect 59476 7922 59505 8496
rect 59551 7922 59564 8496
rect 59476 7909 59564 7922
rect 59620 8496 59708 8509
rect 59620 7922 59633 8496
rect 59679 7922 59708 8496
rect 59620 7909 59708 7922
rect 59764 8496 59852 8509
rect 59764 7922 59793 8496
rect 59839 7922 59852 8496
rect 59764 7909 59852 7922
rect 62204 11676 62292 11689
rect 62204 11102 62217 11676
rect 62263 11102 62292 11676
rect 62204 11089 62292 11102
rect 62348 11676 62436 11689
rect 62348 11102 62377 11676
rect 62423 11102 62436 11676
rect 62348 11089 62436 11102
rect 62492 11676 62580 11689
rect 62492 11102 62505 11676
rect 62551 11102 62580 11676
rect 62492 11089 62580 11102
rect 62636 11676 62740 11689
rect 62636 11102 62665 11676
rect 62711 11102 62740 11676
rect 62636 11089 62740 11102
rect 62796 11676 62900 11689
rect 62796 11102 62825 11676
rect 62871 11102 62900 11676
rect 62796 11089 62900 11102
rect 62956 11676 63060 11689
rect 62956 11102 62985 11676
rect 63031 11102 63060 11676
rect 62956 11089 63060 11102
rect 63116 11676 63220 11689
rect 63116 11102 63145 11676
rect 63191 11102 63220 11676
rect 63116 11089 63220 11102
rect 63276 11676 63380 11689
rect 63276 11102 63305 11676
rect 63351 11102 63380 11676
rect 63276 11089 63380 11102
rect 63436 11676 63540 11689
rect 63436 11102 63465 11676
rect 63511 11102 63540 11676
rect 63436 11089 63540 11102
rect 63596 11676 63700 11689
rect 63596 11102 63625 11676
rect 63671 11102 63700 11676
rect 63596 11089 63700 11102
rect 63756 11676 63860 11689
rect 63756 11102 63785 11676
rect 63831 11102 63860 11676
rect 63756 11089 63860 11102
rect 63916 11676 64020 11689
rect 63916 11102 63945 11676
rect 63991 11102 64020 11676
rect 63916 11089 64020 11102
rect 64076 11676 64180 11689
rect 64076 11102 64105 11676
rect 64151 11102 64180 11676
rect 64076 11089 64180 11102
rect 64236 11676 64340 11689
rect 64236 11102 64265 11676
rect 64311 11102 64340 11676
rect 64236 11089 64340 11102
rect 64396 11676 64500 11689
rect 64396 11102 64425 11676
rect 64471 11102 64500 11676
rect 64396 11089 64500 11102
rect 64556 11676 64660 11689
rect 64556 11102 64585 11676
rect 64631 11102 64660 11676
rect 64556 11089 64660 11102
rect 64716 11676 64820 11689
rect 64716 11102 64745 11676
rect 64791 11102 64820 11676
rect 64716 11089 64820 11102
rect 64876 11676 64980 11689
rect 64876 11102 64905 11676
rect 64951 11102 64980 11676
rect 64876 11089 64980 11102
rect 65036 11676 65124 11689
rect 65036 11102 65065 11676
rect 65111 11102 65124 11676
rect 65036 11089 65124 11102
rect 65180 11676 65268 11689
rect 65180 11102 65193 11676
rect 65239 11102 65268 11676
rect 65180 11089 65268 11102
rect 65324 11676 65412 11689
rect 65324 11102 65353 11676
rect 65399 11102 65412 11676
rect 65324 11089 65412 11102
rect 62204 10616 62292 10629
rect 62204 10042 62217 10616
rect 62263 10042 62292 10616
rect 62204 10029 62292 10042
rect 62348 10616 62436 10629
rect 62348 10042 62377 10616
rect 62423 10042 62436 10616
rect 62348 10029 62436 10042
rect 62492 10616 62580 10629
rect 62492 10042 62505 10616
rect 62551 10042 62580 10616
rect 62492 10029 62580 10042
rect 62636 10616 62740 10629
rect 62636 10042 62665 10616
rect 62711 10042 62740 10616
rect 62636 10029 62740 10042
rect 62796 10616 62900 10629
rect 62796 10042 62825 10616
rect 62871 10042 62900 10616
rect 62796 10029 62900 10042
rect 62956 10616 63060 10629
rect 62956 10042 62985 10616
rect 63031 10042 63060 10616
rect 62956 10029 63060 10042
rect 63116 10616 63220 10629
rect 63116 10042 63145 10616
rect 63191 10042 63220 10616
rect 63116 10029 63220 10042
rect 63276 10616 63380 10629
rect 63276 10042 63305 10616
rect 63351 10042 63380 10616
rect 63276 10029 63380 10042
rect 63436 10616 63540 10629
rect 63436 10042 63465 10616
rect 63511 10042 63540 10616
rect 63436 10029 63540 10042
rect 63596 10616 63700 10629
rect 63596 10042 63625 10616
rect 63671 10042 63700 10616
rect 63596 10029 63700 10042
rect 63756 10616 63860 10629
rect 63756 10042 63785 10616
rect 63831 10042 63860 10616
rect 63756 10029 63860 10042
rect 63916 10616 64020 10629
rect 63916 10042 63945 10616
rect 63991 10042 64020 10616
rect 63916 10029 64020 10042
rect 64076 10616 64180 10629
rect 64076 10042 64105 10616
rect 64151 10042 64180 10616
rect 64076 10029 64180 10042
rect 64236 10616 64340 10629
rect 64236 10042 64265 10616
rect 64311 10042 64340 10616
rect 64236 10029 64340 10042
rect 64396 10616 64500 10629
rect 64396 10042 64425 10616
rect 64471 10042 64500 10616
rect 64396 10029 64500 10042
rect 64556 10616 64660 10629
rect 64556 10042 64585 10616
rect 64631 10042 64660 10616
rect 64556 10029 64660 10042
rect 64716 10616 64820 10629
rect 64716 10042 64745 10616
rect 64791 10042 64820 10616
rect 64716 10029 64820 10042
rect 64876 10616 64980 10629
rect 64876 10042 64905 10616
rect 64951 10042 64980 10616
rect 64876 10029 64980 10042
rect 65036 10616 65124 10629
rect 65036 10042 65065 10616
rect 65111 10042 65124 10616
rect 65036 10029 65124 10042
rect 65180 10616 65268 10629
rect 65180 10042 65193 10616
rect 65239 10042 65268 10616
rect 65180 10029 65268 10042
rect 65324 10616 65412 10629
rect 65324 10042 65353 10616
rect 65399 10042 65412 10616
rect 65324 10029 65412 10042
rect 62204 9556 62292 9569
rect 62204 8982 62217 9556
rect 62263 8982 62292 9556
rect 62204 8969 62292 8982
rect 62348 9556 62436 9569
rect 62348 8982 62377 9556
rect 62423 8982 62436 9556
rect 62348 8969 62436 8982
rect 62492 9556 62580 9569
rect 62492 8982 62505 9556
rect 62551 8982 62580 9556
rect 62492 8969 62580 8982
rect 62636 9556 62740 9569
rect 62636 8982 62665 9556
rect 62711 8982 62740 9556
rect 62636 8969 62740 8982
rect 62796 9556 62900 9569
rect 62796 8982 62825 9556
rect 62871 8982 62900 9556
rect 62796 8969 62900 8982
rect 62956 9556 63060 9569
rect 62956 8982 62985 9556
rect 63031 8982 63060 9556
rect 62956 8969 63060 8982
rect 63116 9556 63220 9569
rect 63116 8982 63145 9556
rect 63191 8982 63220 9556
rect 63116 8969 63220 8982
rect 63276 9556 63380 9569
rect 63276 8982 63305 9556
rect 63351 8982 63380 9556
rect 63276 8969 63380 8982
rect 63436 9556 63540 9569
rect 63436 8982 63465 9556
rect 63511 8982 63540 9556
rect 63436 8969 63540 8982
rect 63596 9556 63700 9569
rect 63596 8982 63625 9556
rect 63671 8982 63700 9556
rect 63596 8969 63700 8982
rect 63756 9556 63860 9569
rect 63756 8982 63785 9556
rect 63831 8982 63860 9556
rect 63756 8969 63860 8982
rect 63916 9556 64020 9569
rect 63916 8982 63945 9556
rect 63991 8982 64020 9556
rect 63916 8969 64020 8982
rect 64076 9556 64180 9569
rect 64076 8982 64105 9556
rect 64151 8982 64180 9556
rect 64076 8969 64180 8982
rect 64236 9556 64340 9569
rect 64236 8982 64265 9556
rect 64311 8982 64340 9556
rect 64236 8969 64340 8982
rect 64396 9556 64500 9569
rect 64396 8982 64425 9556
rect 64471 8982 64500 9556
rect 64396 8969 64500 8982
rect 64556 9556 64660 9569
rect 64556 8982 64585 9556
rect 64631 8982 64660 9556
rect 64556 8969 64660 8982
rect 64716 9556 64820 9569
rect 64716 8982 64745 9556
rect 64791 8982 64820 9556
rect 64716 8969 64820 8982
rect 64876 9556 64980 9569
rect 64876 8982 64905 9556
rect 64951 8982 64980 9556
rect 64876 8969 64980 8982
rect 65036 9556 65124 9569
rect 65036 8982 65065 9556
rect 65111 8982 65124 9556
rect 65036 8969 65124 8982
rect 65180 9556 65268 9569
rect 65180 8982 65193 9556
rect 65239 8982 65268 9556
rect 65180 8969 65268 8982
rect 65324 9556 65412 9569
rect 65324 8982 65353 9556
rect 65399 8982 65412 9556
rect 65324 8969 65412 8982
rect 62204 8496 62292 8509
rect 62204 7922 62217 8496
rect 62263 7922 62292 8496
rect 62204 7909 62292 7922
rect 62348 8496 62436 8509
rect 62348 7922 62377 8496
rect 62423 7922 62436 8496
rect 62348 7909 62436 7922
rect 62492 8496 62580 8509
rect 62492 7922 62505 8496
rect 62551 7922 62580 8496
rect 62492 7909 62580 7922
rect 62636 8496 62740 8509
rect 62636 7922 62665 8496
rect 62711 7922 62740 8496
rect 62636 7909 62740 7922
rect 62796 8496 62900 8509
rect 62796 7922 62825 8496
rect 62871 7922 62900 8496
rect 62796 7909 62900 7922
rect 62956 8496 63060 8509
rect 62956 7922 62985 8496
rect 63031 7922 63060 8496
rect 62956 7909 63060 7922
rect 63116 8496 63220 8509
rect 63116 7922 63145 8496
rect 63191 7922 63220 8496
rect 63116 7909 63220 7922
rect 63276 8496 63380 8509
rect 63276 7922 63305 8496
rect 63351 7922 63380 8496
rect 63276 7909 63380 7922
rect 63436 8496 63540 8509
rect 63436 7922 63465 8496
rect 63511 7922 63540 8496
rect 63436 7909 63540 7922
rect 63596 8496 63700 8509
rect 63596 7922 63625 8496
rect 63671 7922 63700 8496
rect 63596 7909 63700 7922
rect 63756 8496 63860 8509
rect 63756 7922 63785 8496
rect 63831 7922 63860 8496
rect 63756 7909 63860 7922
rect 63916 8496 64020 8509
rect 63916 7922 63945 8496
rect 63991 7922 64020 8496
rect 63916 7909 64020 7922
rect 64076 8496 64180 8509
rect 64076 7922 64105 8496
rect 64151 7922 64180 8496
rect 64076 7909 64180 7922
rect 64236 8496 64340 8509
rect 64236 7922 64265 8496
rect 64311 7922 64340 8496
rect 64236 7909 64340 7922
rect 64396 8496 64500 8509
rect 64396 7922 64425 8496
rect 64471 7922 64500 8496
rect 64396 7909 64500 7922
rect 64556 8496 64660 8509
rect 64556 7922 64585 8496
rect 64631 7922 64660 8496
rect 64556 7909 64660 7922
rect 64716 8496 64820 8509
rect 64716 7922 64745 8496
rect 64791 7922 64820 8496
rect 64716 7909 64820 7922
rect 64876 8496 64980 8509
rect 64876 7922 64905 8496
rect 64951 7922 64980 8496
rect 64876 7909 64980 7922
rect 65036 8496 65124 8509
rect 65036 7922 65065 8496
rect 65111 7922 65124 8496
rect 65036 7909 65124 7922
rect 65180 8496 65268 8509
rect 65180 7922 65193 8496
rect 65239 7922 65268 8496
rect 65180 7909 65268 7922
rect 65324 8496 65412 8509
rect 65324 7922 65353 8496
rect 65399 7922 65412 8496
rect 65324 7909 65412 7922
rect 1277 4421 1365 4434
rect 1277 3647 1290 4421
rect 1336 3647 1365 4421
rect 1277 3634 1365 3647
rect 1421 4421 1509 4434
rect 1421 3647 1450 4421
rect 1496 3647 1509 4421
rect 1421 3634 1509 3647
rect 1565 4421 1653 4434
rect 1565 3647 1578 4421
rect 1624 3647 1653 4421
rect 1565 3634 1653 3647
rect 1709 4421 1797 4434
rect 1709 3647 1738 4421
rect 1784 3647 1797 4421
rect 1709 3634 1797 3647
rect 1853 4421 1941 4434
rect 1853 3647 1866 4421
rect 1912 3647 1941 4421
rect 1853 3634 1941 3647
rect 2053 4421 2157 4434
rect 2053 3647 2082 4421
rect 2128 3647 2157 4421
rect 2053 3634 2157 3647
rect 2269 4421 2373 4434
rect 2269 3647 2298 4421
rect 2344 3647 2373 4421
rect 2269 3634 2373 3647
rect 2485 4421 2589 4434
rect 2485 3647 2514 4421
rect 2560 3647 2589 4421
rect 2485 3634 2589 3647
rect 2701 4421 2805 4434
rect 2701 3647 2730 4421
rect 2776 3647 2805 4421
rect 2701 3634 2805 3647
rect 2917 4421 3021 4434
rect 2917 3647 2946 4421
rect 2992 3647 3021 4421
rect 2917 3634 3021 3647
rect 3133 4421 3237 4434
rect 3133 3647 3162 4421
rect 3208 3647 3237 4421
rect 3133 3634 3237 3647
rect 3349 4421 3453 4434
rect 3349 3647 3378 4421
rect 3424 3647 3453 4421
rect 3349 3634 3453 3647
rect 3565 4421 3669 4434
rect 3565 3647 3594 4421
rect 3640 3647 3669 4421
rect 3565 3634 3669 3647
rect 3781 4421 3885 4434
rect 3781 3647 3810 4421
rect 3856 3647 3885 4421
rect 3781 3634 3885 3647
rect 3997 4421 4101 4434
rect 3997 3647 4026 4421
rect 4072 3647 4101 4421
rect 3997 3634 4101 3647
rect 4213 4421 4317 4434
rect 4213 3647 4242 4421
rect 4288 3647 4317 4421
rect 4213 3634 4317 3647
rect 4373 4421 4477 4434
rect 4373 3647 4402 4421
rect 4448 3647 4477 4421
rect 4373 3634 4477 3647
rect 4533 4421 4621 4434
rect 4533 3647 4562 4421
rect 4608 3647 4621 4421
rect 4533 3634 4621 3647
rect 1277 3161 1365 3174
rect 1277 2387 1290 3161
rect 1336 2387 1365 3161
rect 1277 2374 1365 2387
rect 1421 3161 1509 3174
rect 1421 2387 1450 3161
rect 1496 2387 1509 3161
rect 1421 2374 1509 2387
rect 1573 3161 1661 3174
rect 1573 2387 1586 3161
rect 1632 2387 1661 3161
rect 1573 2374 1661 2387
rect 1717 3161 1805 3174
rect 1717 2387 1746 3161
rect 1792 2387 1805 3161
rect 1717 2374 1805 2387
rect 1861 3161 1949 3174
rect 1861 2387 1874 3161
rect 1920 2387 1949 3161
rect 1861 2374 1949 2387
rect 2061 3161 2165 3174
rect 2061 2387 2090 3161
rect 2136 2387 2165 3161
rect 2061 2374 2165 2387
rect 2277 3161 2381 3174
rect 2277 2387 2306 3161
rect 2352 2387 2381 3161
rect 2277 2374 2381 2387
rect 2493 3161 2597 3174
rect 2493 2387 2522 3161
rect 2568 2387 2597 3161
rect 2493 2374 2597 2387
rect 2709 3161 2813 3174
rect 2709 2387 2738 3161
rect 2784 2387 2813 3161
rect 2709 2374 2813 2387
rect 2925 3161 3029 3174
rect 2925 2387 2954 3161
rect 3000 2387 3029 3161
rect 2925 2374 3029 2387
rect 3085 3161 3189 3174
rect 3085 2387 3114 3161
rect 3160 2387 3189 3161
rect 3085 2374 3189 2387
rect 3245 3161 3349 3174
rect 3245 2387 3274 3161
rect 3320 2387 3349 3161
rect 3245 2374 3349 2387
rect 3405 3161 3509 3174
rect 3405 2387 3434 3161
rect 3480 2387 3509 3161
rect 3405 2374 3509 2387
rect 3565 3161 3669 3174
rect 3565 2387 3594 3161
rect 3640 2387 3669 3161
rect 3565 2374 3669 2387
rect 3781 3161 3869 3174
rect 3781 2387 3810 3161
rect 3856 2387 3869 3161
rect 3781 2374 3869 2387
rect 3925 3161 4013 3174
rect 3925 2387 3938 3161
rect 3984 2387 4013 3161
rect 3925 2374 4013 2387
rect 4125 3161 4229 3174
rect 4125 2387 4154 3161
rect 4200 2387 4229 3161
rect 4125 2374 4229 2387
rect 4285 3161 4373 3174
rect 4285 2387 4314 3161
rect 4360 2387 4373 3161
rect 4285 2374 4373 2387
rect 4437 3161 4525 3174
rect 4437 2387 4450 3161
rect 4496 2387 4525 3161
rect 4437 2374 4525 2387
rect 4581 3161 4669 3174
rect 4581 2387 4610 3161
rect 4656 2387 4669 3161
rect 4581 2374 4669 2387
rect 1277 1901 1365 1914
rect 1277 1827 1290 1901
rect 1336 1827 1365 1901
rect 1277 1814 1365 1827
rect 1421 1901 1509 1914
rect 1421 1827 1450 1901
rect 1496 1827 1509 1901
rect 1421 1814 1509 1827
rect 1573 1901 1661 1914
rect 1573 1827 1586 1901
rect 1632 1827 1661 1901
rect 1573 1814 1661 1827
rect 1717 1901 1821 1914
rect 1717 1827 1746 1901
rect 1792 1827 1821 1901
rect 1717 1814 1821 1827
rect 1877 1901 1981 1914
rect 1877 1827 1906 1901
rect 1952 1827 1981 1901
rect 1877 1814 1981 1827
rect 2037 1901 2141 1914
rect 2037 1827 2066 1901
rect 2112 1827 2141 1901
rect 2037 1814 2141 1827
rect 2197 1901 2301 1914
rect 2197 1827 2226 1901
rect 2272 1827 2301 1901
rect 2197 1814 2301 1827
rect 2357 1901 2461 1914
rect 2357 1827 2386 1901
rect 2432 1827 2461 1901
rect 2357 1814 2461 1827
rect 2517 1901 2621 1914
rect 2517 1827 2546 1901
rect 2592 1827 2621 1901
rect 2517 1814 2621 1827
rect 2677 1901 2781 1914
rect 2677 1827 2706 1901
rect 2752 1827 2781 1901
rect 2677 1814 2781 1827
rect 2837 1901 2941 1914
rect 2837 1827 2866 1901
rect 2912 1827 2941 1901
rect 2837 1814 2941 1827
rect 2997 1901 3101 1914
rect 2997 1827 3026 1901
rect 3072 1827 3101 1901
rect 2997 1814 3101 1827
rect 3157 1901 3261 1914
rect 3157 1827 3186 1901
rect 3232 1827 3261 1901
rect 3157 1814 3261 1827
rect 3317 1901 3421 1914
rect 3317 1827 3346 1901
rect 3392 1827 3421 1901
rect 3317 1814 3421 1827
rect 3477 1901 3581 1914
rect 3477 1827 3506 1901
rect 3552 1827 3581 1901
rect 3477 1814 3581 1827
rect 3637 1901 3741 1914
rect 3637 1827 3666 1901
rect 3712 1827 3741 1901
rect 3637 1814 3741 1827
rect 3797 1901 3901 1914
rect 3797 1827 3826 1901
rect 3872 1827 3901 1901
rect 3797 1814 3901 1827
rect 3957 1901 4061 1914
rect 3957 1827 3986 1901
rect 4032 1827 4061 1901
rect 3957 1814 4061 1827
rect 4117 1901 4221 1914
rect 4117 1827 4146 1901
rect 4192 1827 4221 1901
rect 4117 1814 4221 1827
rect 4421 1901 4525 1914
rect 4421 1827 4450 1901
rect 4496 1827 4525 1901
rect 4421 1814 4525 1827
rect 4581 1901 4669 1914
rect 4581 1827 4610 1901
rect 4656 1827 4669 1901
rect 4581 1814 4669 1827
rect 18782 4766 18870 4779
rect 18782 4192 18795 4766
rect 18841 4192 18870 4766
rect 18782 4179 18870 4192
rect 18926 4766 19030 4779
rect 18926 4192 18955 4766
rect 19001 4192 19030 4766
rect 18926 4179 19030 4192
rect 19086 4766 19190 4779
rect 19086 4192 19115 4766
rect 19161 4192 19190 4766
rect 19086 4179 19190 4192
rect 19246 4766 19350 4779
rect 19246 4192 19275 4766
rect 19321 4192 19350 4766
rect 19246 4179 19350 4192
rect 19406 4766 19510 4779
rect 19406 4192 19435 4766
rect 19481 4192 19510 4766
rect 19406 4179 19510 4192
rect 19566 4766 19670 4779
rect 19566 4192 19595 4766
rect 19641 4192 19670 4766
rect 19566 4179 19670 4192
rect 19726 4766 19830 4779
rect 19726 4192 19755 4766
rect 19801 4192 19830 4766
rect 19726 4179 19830 4192
rect 19886 4766 19990 4779
rect 19886 4192 19915 4766
rect 19961 4192 19990 4766
rect 19886 4179 19990 4192
rect 20046 4766 20150 4779
rect 20046 4192 20075 4766
rect 20121 4192 20150 4766
rect 20046 4179 20150 4192
rect 20206 4766 20310 4779
rect 20206 4192 20235 4766
rect 20281 4192 20310 4766
rect 20206 4179 20310 4192
rect 20366 4766 20470 4779
rect 20366 4192 20395 4766
rect 20441 4192 20470 4766
rect 20366 4179 20470 4192
rect 20526 4766 20630 4779
rect 20526 4192 20555 4766
rect 20601 4192 20630 4766
rect 20526 4179 20630 4192
rect 20686 4766 20790 4779
rect 20686 4192 20715 4766
rect 20761 4192 20790 4766
rect 20686 4179 20790 4192
rect 20846 4766 20950 4779
rect 20846 4192 20875 4766
rect 20921 4192 20950 4766
rect 20846 4179 20950 4192
rect 21006 4766 21110 4779
rect 21006 4192 21035 4766
rect 21081 4192 21110 4766
rect 21006 4179 21110 4192
rect 21166 4766 21270 4779
rect 21166 4192 21195 4766
rect 21241 4192 21270 4766
rect 21166 4179 21270 4192
rect 21326 4766 21430 4779
rect 21326 4192 21355 4766
rect 21401 4192 21430 4766
rect 21326 4179 21430 4192
rect 21486 4766 21590 4779
rect 21486 4192 21515 4766
rect 21561 4192 21590 4766
rect 21486 4179 21590 4192
rect 21646 4766 21750 4779
rect 21646 4192 21675 4766
rect 21721 4192 21750 4766
rect 21646 4179 21750 4192
rect 21806 4766 21894 4779
rect 21806 4192 21835 4766
rect 21881 4192 21894 4766
rect 21806 4179 21894 4192
rect 21950 4766 22038 4779
rect 21950 4192 21963 4766
rect 22009 4192 22038 4766
rect 21950 4179 22038 4192
rect 22094 4766 22182 4779
rect 22094 4192 22123 4766
rect 22169 4192 22182 4766
rect 22094 4179 22182 4192
rect 22238 4766 22326 4779
rect 22238 4192 22251 4766
rect 22297 4192 22326 4766
rect 22238 4179 22326 4192
rect 22382 4766 22470 4779
rect 22382 4192 22411 4766
rect 22457 4192 22470 4766
rect 22382 4179 22470 4192
rect 18782 4030 18870 4043
rect 18782 3456 18795 4030
rect 18841 3456 18870 4030
rect 18782 3443 18870 3456
rect 18926 4030 19030 4043
rect 18926 3456 18955 4030
rect 19001 3456 19030 4030
rect 18926 3443 19030 3456
rect 19086 4030 19190 4043
rect 19086 3456 19115 4030
rect 19161 3456 19190 4030
rect 19086 3443 19190 3456
rect 19246 4030 19350 4043
rect 19246 3456 19275 4030
rect 19321 3456 19350 4030
rect 19246 3443 19350 3456
rect 19406 4030 19510 4043
rect 19406 3456 19435 4030
rect 19481 3456 19510 4030
rect 19406 3443 19510 3456
rect 19566 4030 19670 4043
rect 19566 3456 19595 4030
rect 19641 3456 19670 4030
rect 19566 3443 19670 3456
rect 19726 4030 19830 4043
rect 19726 3456 19755 4030
rect 19801 3456 19830 4030
rect 19726 3443 19830 3456
rect 19886 4030 19990 4043
rect 19886 3456 19915 4030
rect 19961 3456 19990 4030
rect 19886 3443 19990 3456
rect 20046 4030 20150 4043
rect 20046 3456 20075 4030
rect 20121 3456 20150 4030
rect 20046 3443 20150 3456
rect 20206 4030 20310 4043
rect 20206 3456 20235 4030
rect 20281 3456 20310 4030
rect 20206 3443 20310 3456
rect 20366 4030 20470 4043
rect 20366 3456 20395 4030
rect 20441 3456 20470 4030
rect 20366 3443 20470 3456
rect 20526 4030 20630 4043
rect 20526 3456 20555 4030
rect 20601 3456 20630 4030
rect 20526 3443 20630 3456
rect 20686 4030 20790 4043
rect 20686 3456 20715 4030
rect 20761 3456 20790 4030
rect 20686 3443 20790 3456
rect 20846 4030 20950 4043
rect 20846 3456 20875 4030
rect 20921 3456 20950 4030
rect 20846 3443 20950 3456
rect 21006 4030 21110 4043
rect 21006 3456 21035 4030
rect 21081 3456 21110 4030
rect 21006 3443 21110 3456
rect 21166 4030 21270 4043
rect 21166 3456 21195 4030
rect 21241 3456 21270 4030
rect 21166 3443 21270 3456
rect 21326 4030 21430 4043
rect 21326 3456 21355 4030
rect 21401 3456 21430 4030
rect 21326 3443 21430 3456
rect 21486 4030 21590 4043
rect 21486 3456 21515 4030
rect 21561 3456 21590 4030
rect 21486 3443 21590 3456
rect 21646 4030 21750 4043
rect 21646 3456 21675 4030
rect 21721 3456 21750 4030
rect 21646 3443 21750 3456
rect 21806 4030 21894 4043
rect 21806 3456 21835 4030
rect 21881 3456 21894 4030
rect 21806 3443 21894 3456
rect 21950 4030 22038 4043
rect 21950 3456 21963 4030
rect 22009 3456 22038 4030
rect 21950 3443 22038 3456
rect 22094 4030 22182 4043
rect 22094 3456 22123 4030
rect 22169 3456 22182 4030
rect 22094 3443 22182 3456
rect 22238 4030 22326 4043
rect 22238 3456 22251 4030
rect 22297 3456 22326 4030
rect 22238 3443 22326 3456
rect 22382 4030 22470 4043
rect 22382 3456 22411 4030
rect 22457 3456 22470 4030
rect 22382 3443 22470 3456
rect 18782 3294 18870 3307
rect 18782 2720 18795 3294
rect 18841 2720 18870 3294
rect 18782 2707 18870 2720
rect 18926 3294 19030 3307
rect 18926 2720 18955 3294
rect 19001 2720 19030 3294
rect 18926 2707 19030 2720
rect 19086 3294 19190 3307
rect 19086 2720 19115 3294
rect 19161 2720 19190 3294
rect 19086 2707 19190 2720
rect 19246 3294 19350 3307
rect 19246 2720 19275 3294
rect 19321 2720 19350 3294
rect 19246 2707 19350 2720
rect 19406 3294 19510 3307
rect 19406 2720 19435 3294
rect 19481 2720 19510 3294
rect 19406 2707 19510 2720
rect 19566 3294 19670 3307
rect 19566 2720 19595 3294
rect 19641 2720 19670 3294
rect 19566 2707 19670 2720
rect 19726 3294 19830 3307
rect 19726 2720 19755 3294
rect 19801 2720 19830 3294
rect 19726 2707 19830 2720
rect 19886 3294 19990 3307
rect 19886 2720 19915 3294
rect 19961 2720 19990 3294
rect 19886 2707 19990 2720
rect 20046 3294 20150 3307
rect 20046 2720 20075 3294
rect 20121 2720 20150 3294
rect 20046 2707 20150 2720
rect 20206 3294 20310 3307
rect 20206 2720 20235 3294
rect 20281 2720 20310 3294
rect 20206 2707 20310 2720
rect 20366 3294 20470 3307
rect 20366 2720 20395 3294
rect 20441 2720 20470 3294
rect 20366 2707 20470 2720
rect 20526 3294 20630 3307
rect 20526 2720 20555 3294
rect 20601 2720 20630 3294
rect 20526 2707 20630 2720
rect 20686 3294 20790 3307
rect 20686 2720 20715 3294
rect 20761 2720 20790 3294
rect 20686 2707 20790 2720
rect 20846 3294 20950 3307
rect 20846 2720 20875 3294
rect 20921 2720 20950 3294
rect 20846 2707 20950 2720
rect 21006 3294 21110 3307
rect 21006 2720 21035 3294
rect 21081 2720 21110 3294
rect 21006 2707 21110 2720
rect 21166 3294 21270 3307
rect 21166 2720 21195 3294
rect 21241 2720 21270 3294
rect 21166 2707 21270 2720
rect 21326 3294 21430 3307
rect 21326 2720 21355 3294
rect 21401 2720 21430 3294
rect 21326 2707 21430 2720
rect 21486 3294 21590 3307
rect 21486 2720 21515 3294
rect 21561 2720 21590 3294
rect 21486 2707 21590 2720
rect 21646 3294 21750 3307
rect 21646 2720 21675 3294
rect 21721 2720 21750 3294
rect 21646 2707 21750 2720
rect 21806 3294 21894 3307
rect 21806 2720 21835 3294
rect 21881 2720 21894 3294
rect 22238 3294 22326 3307
rect 21806 2707 21894 2720
rect 21950 3194 22038 3207
rect 21950 2720 21963 3194
rect 22009 2720 22038 3194
rect 21950 2707 22038 2720
rect 22094 3194 22182 3207
rect 22094 2720 22123 3194
rect 22169 2720 22182 3194
rect 22094 2707 22182 2720
rect 22238 2720 22251 3294
rect 22297 2720 22326 3294
rect 22238 2707 22326 2720
rect 22382 3294 22470 3307
rect 22382 2720 22411 3294
rect 22457 2720 22470 3294
rect 22382 2707 22470 2720
rect 18782 2558 18870 2571
rect 18782 1984 18795 2558
rect 18841 1984 18870 2558
rect 18782 1971 18870 1984
rect 18926 2558 19030 2571
rect 18926 1984 18955 2558
rect 19001 1984 19030 2558
rect 18926 1971 19030 1984
rect 19086 2558 19190 2571
rect 19086 1984 19115 2558
rect 19161 1984 19190 2558
rect 19086 1971 19190 1984
rect 19246 2558 19350 2571
rect 19246 1984 19275 2558
rect 19321 1984 19350 2558
rect 19246 1971 19350 1984
rect 19406 2558 19510 2571
rect 19406 1984 19435 2558
rect 19481 1984 19510 2558
rect 19406 1971 19510 1984
rect 19566 2558 19670 2571
rect 19566 1984 19595 2558
rect 19641 1984 19670 2558
rect 19566 1971 19670 1984
rect 19726 2558 19830 2571
rect 19726 1984 19755 2558
rect 19801 1984 19830 2558
rect 19726 1971 19830 1984
rect 19886 2558 19990 2571
rect 19886 1984 19915 2558
rect 19961 1984 19990 2558
rect 19886 1971 19990 1984
rect 20046 2558 20150 2571
rect 20046 1984 20075 2558
rect 20121 1984 20150 2558
rect 20046 1971 20150 1984
rect 20206 2558 20310 2571
rect 20206 1984 20235 2558
rect 20281 1984 20310 2558
rect 20206 1971 20310 1984
rect 20366 2558 20470 2571
rect 20366 1984 20395 2558
rect 20441 1984 20470 2558
rect 20366 1971 20470 1984
rect 20526 2558 20630 2571
rect 20526 1984 20555 2558
rect 20601 1984 20630 2558
rect 20526 1971 20630 1984
rect 20686 2558 20790 2571
rect 20686 1984 20715 2558
rect 20761 1984 20790 2558
rect 20686 1971 20790 1984
rect 20846 2558 20950 2571
rect 20846 1984 20875 2558
rect 20921 1984 20950 2558
rect 20846 1971 20950 1984
rect 21006 2558 21110 2571
rect 21006 1984 21035 2558
rect 21081 1984 21110 2558
rect 21006 1971 21110 1984
rect 21166 2558 21270 2571
rect 21166 1984 21195 2558
rect 21241 1984 21270 2558
rect 21166 1971 21270 1984
rect 21326 2558 21430 2571
rect 21326 1984 21355 2558
rect 21401 1984 21430 2558
rect 21326 1971 21430 1984
rect 21486 2558 21590 2571
rect 21486 1984 21515 2558
rect 21561 1984 21590 2558
rect 21486 1971 21590 1984
rect 21646 2558 21750 2571
rect 21646 1984 21675 2558
rect 21721 1984 21750 2558
rect 21646 1971 21750 1984
rect 21806 2558 21894 2571
rect 21806 1984 21835 2558
rect 21881 1984 21894 2558
rect 22238 2558 22326 2571
rect 21806 1971 21894 1984
rect 21950 2458 22038 2471
rect 21950 1984 21963 2458
rect 22009 1984 22038 2458
rect 21950 1971 22038 1984
rect 22094 2458 22182 2471
rect 22094 1984 22123 2458
rect 22169 1984 22182 2458
rect 22094 1971 22182 1984
rect 22238 1984 22251 2558
rect 22297 1984 22326 2558
rect 22238 1971 22326 1984
rect 22382 2558 22470 2571
rect 22382 1984 22411 2558
rect 22457 1984 22470 2558
rect 22382 1971 22470 1984
<< ndiffc >>
rect 6462 13713 6508 14263
rect 6622 13713 6668 14263
rect 6750 13713 6796 14263
rect 6910 13713 6956 14263
rect 7070 13713 7116 14263
rect 7230 13713 7276 14263
rect 7390 13713 7436 14263
rect 7550 13713 7596 14263
rect 7710 13713 7756 14263
rect 7870 13713 7916 14263
rect 8030 13713 8076 14263
rect 8158 13713 8204 14263
rect 8318 13713 8364 14263
rect 6462 12851 6508 13401
rect 6622 12851 6668 13401
rect 6750 12851 6796 13401
rect 6910 12851 6956 13401
rect 7070 12851 7116 13401
rect 7230 12851 7276 13401
rect 7390 12851 7436 13401
rect 7550 12851 7596 13401
rect 7710 12851 7756 13401
rect 7870 12851 7916 13401
rect 8030 12851 8076 13401
rect 8158 12851 8204 13401
rect 8318 12851 8364 13401
rect 6462 11989 6508 12539
rect 6622 11989 6668 12539
rect 6750 11989 6796 12539
rect 6910 11989 6956 12539
rect 7070 11989 7116 12539
rect 7230 11989 7276 12539
rect 7390 11989 7436 12539
rect 7550 11989 7596 12539
rect 7710 11989 7756 12539
rect 7870 11989 7916 12539
rect 8030 11989 8076 12539
rect 8158 11989 8204 12539
rect 8318 11989 8364 12539
rect 18712 12602 18758 13176
rect 18872 12602 18918 13176
rect 19000 12602 19046 13176
rect 19160 12602 19206 13176
rect 19320 12602 19366 13176
rect 19480 12602 19526 13176
rect 19640 12602 19686 13176
rect 19800 12602 19846 13176
rect 19960 12602 20006 13176
rect 20120 12602 20166 13176
rect 20280 12602 20326 13176
rect 20408 12602 20454 13176
rect 20568 12602 20614 13176
rect 6462 11127 6508 11677
rect 6622 11127 6668 11677
rect 6750 11127 6796 11677
rect 6910 11127 6956 11677
rect 7070 11127 7116 11677
rect 7230 11127 7276 11677
rect 7390 11127 7436 11677
rect 7550 11127 7596 11677
rect 7710 11127 7756 11677
rect 7870 11127 7916 11677
rect 8030 11127 8076 11677
rect 8158 11127 8204 11677
rect 8318 11127 8364 11677
rect 6462 10265 6508 10815
rect 6622 10265 6668 10815
rect 6750 10265 6796 10815
rect 6910 10265 6956 10815
rect 7070 10265 7116 10815
rect 7230 10265 7276 10815
rect 7390 10265 7436 10815
rect 7550 10265 7596 10815
rect 7710 10265 7756 10815
rect 7870 10265 7916 10815
rect 8030 10265 8076 10815
rect 8158 10265 8204 10815
rect 8318 10265 8364 10815
rect 8697 10246 8743 10796
rect 8857 10246 8903 10796
rect 8985 10246 9031 10796
rect 9145 10246 9191 10796
rect 9273 10246 9319 10796
rect 9433 10246 9479 10796
rect 9593 10246 9639 10796
rect 9721 10246 9767 10796
rect 9881 10246 9927 10796
rect 10041 10246 10087 10796
rect 10169 10246 10215 10796
rect 10329 10246 10375 10796
rect 10489 10246 10535 10796
rect 10617 10246 10663 10796
rect 10777 10246 10823 10796
rect 10905 10246 10951 10796
rect 11065 10246 11111 10796
rect 6462 9403 6508 9953
rect 6622 9403 6668 9953
rect 6750 9403 6796 9953
rect 6910 9403 6956 9953
rect 7070 9403 7116 9953
rect 7230 9403 7276 9953
rect 7390 9403 7436 9953
rect 7550 9403 7596 9953
rect 7710 9403 7756 9953
rect 7870 9403 7916 9953
rect 8030 9403 8076 9953
rect 8158 9403 8204 9953
rect 8318 9403 8364 9953
rect 8697 9384 8743 9934
rect 8857 9384 8903 9934
rect 8985 9384 9031 9934
rect 9145 9384 9191 9934
rect 9273 9384 9319 9934
rect 9433 9384 9479 9934
rect 9593 9384 9639 9934
rect 9721 9384 9767 9934
rect 9881 9384 9927 9934
rect 10041 9384 10087 9934
rect 10169 9384 10215 9934
rect 10329 9384 10375 9934
rect 10489 9384 10535 9934
rect 10617 9384 10663 9934
rect 10777 9384 10823 9934
rect 10905 9384 10951 9934
rect 11065 9384 11111 9934
rect 6462 8541 6508 9091
rect 6622 8541 6668 9091
rect 6750 8541 6796 9091
rect 6910 8541 6956 9091
rect 7070 8541 7116 9091
rect 7230 8541 7276 9091
rect 7390 8541 7436 9091
rect 7550 8541 7596 9091
rect 7710 8541 7756 9091
rect 7870 8541 7916 9091
rect 8030 8541 8076 9091
rect 8158 8541 8204 9091
rect 8318 8541 8364 9091
rect 8697 8522 8743 9072
rect 8857 8522 8903 9072
rect 8985 8522 9031 9072
rect 9145 8522 9191 9072
rect 9273 8522 9319 9072
rect 9433 8522 9479 9072
rect 9593 8522 9639 9072
rect 9721 8522 9767 9072
rect 9881 8522 9927 9072
rect 10041 8522 10087 9072
rect 10169 8522 10215 9072
rect 10329 8522 10375 9072
rect 10489 8522 10535 9072
rect 10617 8522 10663 9072
rect 10777 8522 10823 9072
rect 10905 8522 10951 9072
rect 11065 8522 11111 9072
rect 6462 7679 6508 8229
rect 6622 7679 6668 8229
rect 6750 7679 6796 8229
rect 6910 7679 6956 8229
rect 7070 7679 7116 8229
rect 7230 7679 7276 8229
rect 7390 7679 7436 8229
rect 7550 7679 7596 8229
rect 7710 7679 7756 8229
rect 7870 7679 7916 8229
rect 8030 7679 8076 8229
rect 8158 7679 8204 8229
rect 8318 7679 8364 8229
rect 8697 7660 8743 8210
rect 8857 7660 8903 8210
rect 8985 7660 9031 8210
rect 9145 7660 9191 8210
rect 9273 7660 9319 8210
rect 9433 7660 9479 8210
rect 9593 7660 9639 8210
rect 9721 7660 9767 8210
rect 9881 7660 9927 8210
rect 10041 7660 10087 8210
rect 10169 7660 10215 8210
rect 10329 7660 10375 8210
rect 10489 7660 10535 8210
rect 10617 7660 10663 8210
rect 10777 7660 10823 8210
rect 10905 7660 10951 8210
rect 11065 7660 11111 8210
rect 18712 11666 18758 12240
rect 18872 11666 18918 12240
rect 19000 11666 19046 12240
rect 19160 11666 19206 12240
rect 19320 11666 19366 12240
rect 19480 11666 19526 12240
rect 19640 11666 19686 12240
rect 19800 11666 19846 12240
rect 19960 11666 20006 12240
rect 20120 11666 20166 12240
rect 20280 11666 20326 12240
rect 20408 11666 20454 12240
rect 20568 11666 20614 12240
rect 18712 10730 18758 11304
rect 18872 10730 18918 11304
rect 19000 10730 19046 11304
rect 19160 10730 19206 11304
rect 19320 10730 19366 11304
rect 19480 10730 19526 11304
rect 19640 10730 19686 11304
rect 19800 10730 19846 11304
rect 19960 10730 20006 11304
rect 20120 10730 20166 11304
rect 20280 10730 20326 11304
rect 20408 10730 20454 11304
rect 20568 10730 20614 11304
rect 18712 9794 18758 10368
rect 18872 9794 18918 10368
rect 19000 9794 19046 10368
rect 19160 9794 19206 10368
rect 19320 9794 19366 10368
rect 19480 9794 19526 10368
rect 19640 9794 19686 10368
rect 19800 9794 19846 10368
rect 19960 9794 20006 10368
rect 20120 9794 20166 10368
rect 20280 9794 20326 10368
rect 20408 9794 20454 10368
rect 20568 9794 20614 10368
rect 18712 8858 18758 9432
rect 18872 8858 18918 9432
rect 19000 8858 19046 9432
rect 19160 8858 19206 9432
rect 19320 8858 19366 9432
rect 19480 8858 19526 9432
rect 19640 8858 19686 9432
rect 19800 8858 19846 9432
rect 19960 8858 20006 9432
rect 20120 8858 20166 9432
rect 20280 8858 20326 9432
rect 20408 8858 20454 9432
rect 20568 8858 20614 9432
rect 18712 7922 18758 8496
rect 18872 7922 18918 8496
rect 19000 7922 19046 8496
rect 19160 7922 19206 8496
rect 19320 7922 19366 8496
rect 19480 7922 19526 8496
rect 19640 7922 19686 8496
rect 19800 7922 19846 8496
rect 19960 7922 20006 8496
rect 20120 7922 20166 8496
rect 20280 7922 20326 8496
rect 20408 7922 20454 8496
rect 20568 7922 20614 8496
rect 23864 12602 23910 13176
rect 24024 12602 24070 13176
rect 24152 12602 24198 13176
rect 24312 12602 24358 13176
rect 24472 12602 24518 13176
rect 24632 12602 24678 13176
rect 24792 12602 24838 13176
rect 24952 12602 24998 13176
rect 25112 12602 25158 13176
rect 25272 12602 25318 13176
rect 25432 12602 25478 13176
rect 25560 12602 25606 13176
rect 25720 12602 25766 13176
rect 23864 11666 23910 12240
rect 24024 11666 24070 12240
rect 24152 11666 24198 12240
rect 24312 11666 24358 12240
rect 24472 11666 24518 12240
rect 24632 11666 24678 12240
rect 24792 11666 24838 12240
rect 24952 11666 24998 12240
rect 25112 11666 25158 12240
rect 25272 11666 25318 12240
rect 25432 11666 25478 12240
rect 25560 11666 25606 12240
rect 25720 11666 25766 12240
rect 23864 10730 23910 11304
rect 24024 10730 24070 11304
rect 24152 10730 24198 11304
rect 24312 10730 24358 11304
rect 24472 10730 24518 11304
rect 24632 10730 24678 11304
rect 24792 10730 24838 11304
rect 24952 10730 24998 11304
rect 25112 10730 25158 11304
rect 25272 10730 25318 11304
rect 25432 10730 25478 11304
rect 25560 10730 25606 11304
rect 25720 10730 25766 11304
rect 23864 9794 23910 10368
rect 24024 9794 24070 10368
rect 24152 9794 24198 10368
rect 24312 9794 24358 10368
rect 24472 9794 24518 10368
rect 24632 9794 24678 10368
rect 24792 9794 24838 10368
rect 24952 9794 24998 10368
rect 25112 9794 25158 10368
rect 25272 9794 25318 10368
rect 25432 9794 25478 10368
rect 25560 9794 25606 10368
rect 25720 9794 25766 10368
rect 23864 8858 23910 9432
rect 24024 8858 24070 9432
rect 24152 8858 24198 9432
rect 24312 8858 24358 9432
rect 24472 8858 24518 9432
rect 24632 8858 24678 9432
rect 24792 8858 24838 9432
rect 24952 8858 24998 9432
rect 25112 8858 25158 9432
rect 25272 8858 25318 9432
rect 25432 8858 25478 9432
rect 25560 8858 25606 9432
rect 25720 8858 25766 9432
rect 23864 7922 23910 8496
rect 24024 7922 24070 8496
rect 24152 7922 24198 8496
rect 24312 7922 24358 8496
rect 24472 7922 24518 8496
rect 24632 7922 24678 8496
rect 24792 7922 24838 8496
rect 24952 7922 24998 8496
rect 25112 7922 25158 8496
rect 25272 7922 25318 8496
rect 25432 7922 25478 8496
rect 25560 7922 25606 8496
rect 25720 7922 25766 8496
rect 27833 12602 27879 13176
rect 27993 12602 28039 13176
rect 28121 12602 28167 13176
rect 28281 12602 28327 13176
rect 28441 12602 28487 13176
rect 28601 12602 28647 13176
rect 28761 12602 28807 13176
rect 28921 12602 28967 13176
rect 29081 12602 29127 13176
rect 29241 12602 29287 13176
rect 29401 12602 29447 13176
rect 29529 12602 29575 13176
rect 29689 12602 29735 13176
rect 27833 11666 27879 12240
rect 27993 11666 28039 12240
rect 28121 11666 28167 12240
rect 28281 11666 28327 12240
rect 28441 11666 28487 12240
rect 28601 11666 28647 12240
rect 28761 11666 28807 12240
rect 28921 11666 28967 12240
rect 29081 11666 29127 12240
rect 29241 11666 29287 12240
rect 29401 11666 29447 12240
rect 29529 11666 29575 12240
rect 29689 11666 29735 12240
rect 27833 10730 27879 11304
rect 27993 10730 28039 11304
rect 28121 10730 28167 11304
rect 28281 10730 28327 11304
rect 28441 10730 28487 11304
rect 28601 10730 28647 11304
rect 28761 10730 28807 11304
rect 28921 10730 28967 11304
rect 29081 10730 29127 11304
rect 29241 10730 29287 11304
rect 29401 10730 29447 11304
rect 29529 10730 29575 11304
rect 29689 10730 29735 11304
rect 27833 9794 27879 10368
rect 27993 9794 28039 10368
rect 28121 9794 28167 10368
rect 28281 9794 28327 10368
rect 28441 9794 28487 10368
rect 28601 9794 28647 10368
rect 28761 9794 28807 10368
rect 28921 9794 28967 10368
rect 29081 9794 29127 10368
rect 29241 9794 29287 10368
rect 29401 9794 29447 10368
rect 29529 9794 29575 10368
rect 29689 9794 29735 10368
rect 27833 8858 27879 9432
rect 27993 8858 28039 9432
rect 28121 8858 28167 9432
rect 28281 8858 28327 9432
rect 28441 8858 28487 9432
rect 28601 8858 28647 9432
rect 28761 8858 28807 9432
rect 28921 8858 28967 9432
rect 29081 8858 29127 9432
rect 29241 8858 29287 9432
rect 29401 8858 29447 9432
rect 29529 8858 29575 9432
rect 29689 8858 29735 9432
rect 27833 7922 27879 8496
rect 27993 7922 28039 8496
rect 28121 7922 28167 8496
rect 28281 7922 28327 8496
rect 28441 7922 28487 8496
rect 28601 7922 28647 8496
rect 28761 7922 28807 8496
rect 28921 7922 28967 8496
rect 29081 7922 29127 8496
rect 29241 7922 29287 8496
rect 29401 7922 29447 8496
rect 29529 7922 29575 8496
rect 29689 7922 29735 8496
rect 7396 5551 7442 5725
rect 7556 5551 7602 5725
rect 7684 5551 7730 5725
rect 7844 5551 7890 5725
rect 8004 5551 8050 5725
rect 8164 5551 8210 5725
rect 8324 5551 8370 5725
rect 8484 5551 8530 5725
rect 8644 5551 8690 5725
rect 8804 5551 8850 5725
rect 8964 5551 9010 5725
rect 9124 5551 9170 5725
rect 9284 5551 9330 5725
rect 9412 5551 9458 5725
rect 9572 5551 9618 5725
rect 7396 5015 7442 5189
rect 7556 5015 7602 5189
rect 7684 5015 7730 5189
rect 7844 5015 7890 5189
rect 8004 5015 8050 5189
rect 8164 5015 8210 5189
rect 8324 5015 8370 5189
rect 8484 5015 8530 5189
rect 8644 5015 8690 5189
rect 8804 5015 8850 5189
rect 8964 5015 9010 5189
rect 9124 5015 9170 5189
rect 9284 5015 9330 5189
rect 9412 5015 9458 5189
rect 9572 5015 9618 5189
rect 7396 4479 7442 4653
rect 7556 4479 7602 4653
rect 7684 4479 7730 4653
rect 7844 4479 7890 4653
rect 8004 4479 8050 4653
rect 8164 4479 8210 4653
rect 8324 4479 8370 4653
rect 8484 4479 8530 4653
rect 8644 4479 8690 4653
rect 8804 4479 8850 4653
rect 8964 4479 9010 4653
rect 9124 4479 9170 4653
rect 9284 4479 9330 4653
rect 9412 4479 9458 4653
rect 9572 4479 9618 4653
rect 7396 3943 7442 4117
rect 7556 3943 7602 4117
rect 7684 3943 7730 4117
rect 7844 3943 7890 4117
rect 8004 3943 8050 4117
rect 8164 3943 8210 4117
rect 8324 3943 8370 4117
rect 8484 3943 8530 4117
rect 8644 3943 8690 4117
rect 8804 3943 8850 4117
rect 8964 3943 9010 4117
rect 9124 3943 9170 4117
rect 9284 3943 9330 4117
rect 9412 3943 9458 4117
rect 9572 3943 9618 4117
rect 7396 3407 7442 3581
rect 7556 3407 7602 3581
rect 7684 3407 7730 3581
rect 7844 3407 7890 3581
rect 8004 3407 8050 3581
rect 8164 3407 8210 3581
rect 8324 3407 8370 3581
rect 8484 3407 8530 3581
rect 8644 3407 8690 3581
rect 8804 3407 8850 3581
rect 8964 3407 9010 3581
rect 9124 3407 9170 3581
rect 9284 3407 9330 3581
rect 9412 3407 9458 3581
rect 9572 3407 9618 3581
rect 7396 2871 7442 3045
rect 7556 2871 7602 3045
rect 7684 2871 7730 3045
rect 7844 2871 7890 3045
rect 8004 2871 8050 3045
rect 8164 2871 8210 3045
rect 8324 2871 8370 3045
rect 8484 2871 8530 3045
rect 8644 2871 8690 3045
rect 8804 2871 8850 3045
rect 8964 2871 9010 3045
rect 9124 2871 9170 3045
rect 9284 2871 9330 3045
rect 9412 2871 9458 3045
rect 9572 2871 9618 3045
rect 12683 3394 12729 3768
rect 12987 3394 13033 3768
rect 13115 3394 13161 3768
rect 13419 3394 13465 3768
rect 13723 3394 13769 3768
rect 14027 3394 14073 3768
rect 14331 3394 14377 3768
rect 14635 3394 14681 3768
rect 14939 3394 14985 3768
rect 15067 3394 15113 3768
rect 15371 3394 15417 3768
rect 15675 3394 15721 3768
rect 15979 3394 16025 3768
rect 16283 3394 16329 3768
rect 16587 3394 16633 3768
rect 16891 3394 16937 3768
rect 6149 2242 6195 2416
rect 6309 2242 6355 2416
rect 6437 2242 6483 2416
rect 6597 2242 6643 2416
rect 6757 2242 6803 2416
rect 6917 2242 6963 2416
rect 7077 2242 7123 2416
rect 7237 2242 7283 2416
rect 7397 2242 7443 2416
rect 7557 2242 7603 2416
rect 7717 2242 7763 2416
rect 7877 2242 7923 2416
rect 8037 2242 8083 2416
rect 8197 2242 8243 2416
rect 8357 2242 8403 2416
rect 8517 2242 8563 2416
rect 8677 2242 8723 2416
rect 8837 2242 8883 2416
rect 8997 2242 9043 2416
rect 9157 2242 9203 2416
rect 9317 2242 9363 2416
rect 9445 2242 9491 2416
rect 9749 2242 9795 2416
rect 10053 2242 10099 2416
rect 10357 2242 10403 2416
rect 10661 2242 10707 2416
rect 10821 2242 10867 2416
rect 6149 1605 6195 1779
rect 6309 1605 6355 1779
rect 6437 1605 6483 1779
rect 6653 1605 6699 1779
rect 6869 1605 6915 1779
rect 7085 1605 7131 1779
rect 7301 1605 7347 1779
rect 7517 1605 7563 1779
rect 7733 1605 7779 1779
rect 7949 1605 7995 1779
rect 8165 1605 8211 1779
rect 8381 1605 8427 1779
rect 8597 1605 8643 1779
rect 8757 1605 8803 1779
rect 8917 1605 8963 1779
rect 9077 1605 9123 1779
rect 9237 1605 9283 1779
rect 9397 1605 9443 1779
rect 9557 1605 9603 1779
rect 9717 1605 9763 1779
rect 9861 1605 9907 1779
rect 10021 1605 10067 1779
rect 10181 1605 10227 1779
rect 10341 1605 10387 1779
rect 10501 1605 10547 1779
rect 10661 1605 10707 1779
rect 10821 1605 10867 1779
rect 12683 2858 12729 3232
rect 12987 2858 13033 3232
rect 13115 2858 13161 3232
rect 13419 2858 13465 3232
rect 13723 2858 13769 3232
rect 14027 2858 14073 3232
rect 14331 2858 14377 3232
rect 14635 2858 14681 3232
rect 14939 2858 14985 3232
rect 15067 2858 15113 3232
rect 15371 2858 15417 3232
rect 15675 2858 15721 3232
rect 15979 2858 16025 3232
rect 16283 2858 16329 3232
rect 16587 2858 16633 3232
rect 16891 2858 16937 3232
rect 12683 2022 12729 2396
rect 12987 2022 13033 2396
rect 13115 2022 13161 2396
rect 13419 2022 13465 2396
rect 13723 2022 13769 2396
rect 14027 2022 14073 2396
rect 14331 2022 14377 2396
rect 14635 2022 14681 2396
rect 14939 2022 14985 2396
rect 15067 2022 15113 2396
rect 15371 2022 15417 2396
rect 15675 2022 15721 2396
rect 15979 2022 16025 2396
rect 16283 2022 16329 2396
rect 16587 2022 16633 2396
rect 16891 2022 16937 2396
<< pdiffc >>
rect 3597 13289 3643 14013
rect 3757 13289 3803 14013
rect 3885 13289 3931 14013
rect 4045 13289 4091 14013
rect 4205 13289 4251 14013
rect 4365 13289 4411 14013
rect 4525 13289 4571 14013
rect 4685 13289 4731 14013
rect 4845 13289 4891 14013
rect 5005 13289 5051 14013
rect 5165 13289 5211 14013
rect 5293 13289 5339 14013
rect 5453 13289 5499 14013
rect 3597 12159 3643 12883
rect 3757 12159 3803 12883
rect 3885 12159 3931 12883
rect 4045 12159 4091 12883
rect 4205 12159 4251 12883
rect 4365 12159 4411 12883
rect 4525 12159 4571 12883
rect 4685 12159 4731 12883
rect 4845 12159 4891 12883
rect 5005 12159 5051 12883
rect 5165 12159 5211 12883
rect 5293 12159 5339 12883
rect 5453 12159 5499 12883
rect 3597 11029 3643 11753
rect 3757 11029 3803 11753
rect 3885 11029 3931 11753
rect 4045 11029 4091 11753
rect 4205 11029 4251 11753
rect 4365 11029 4411 11753
rect 4525 11029 4571 11753
rect 4685 11029 4731 11753
rect 4845 11029 4891 11753
rect 5005 11029 5051 11753
rect 5165 11029 5211 11753
rect 5293 11029 5339 11753
rect 5453 11029 5499 11753
rect 911 9945 957 10545
rect 1127 9945 1173 10545
rect 1343 9945 1389 10545
rect 1559 9945 1605 10545
rect 1775 9945 1821 10545
rect 1991 9945 2037 10545
rect 2207 9945 2253 10545
rect 2423 9945 2469 10545
rect 2639 9945 2685 10545
rect 2855 9945 2901 10545
rect 3071 9945 3117 10545
rect 3597 9899 3643 10623
rect 3757 9899 3803 10623
rect 3885 9899 3931 10623
rect 4045 9899 4091 10623
rect 4205 9899 4251 10623
rect 4365 9899 4411 10623
rect 4525 9899 4571 10623
rect 4685 9899 4731 10623
rect 4845 9899 4891 10623
rect 5005 9899 5051 10623
rect 5165 9899 5211 10623
rect 5293 9899 5339 10623
rect 5453 9899 5499 10623
rect 911 9183 957 9783
rect 1127 9183 1173 9783
rect 1343 9183 1389 9783
rect 1559 9183 1605 9783
rect 1775 9183 1821 9783
rect 1991 9183 2037 9783
rect 2207 9183 2253 9783
rect 2423 9183 2469 9783
rect 2639 9183 2685 9783
rect 2855 9183 2901 9783
rect 3071 9183 3117 9783
rect 911 8421 957 9021
rect 1127 8421 1173 9021
rect 1343 8421 1389 9021
rect 1559 8421 1605 9021
rect 1775 8421 1821 9021
rect 1991 8421 2037 9021
rect 2207 8421 2253 9021
rect 2423 8421 2469 9021
rect 2639 8421 2685 9021
rect 2855 8421 2901 9021
rect 3071 8421 3117 9021
rect 3597 8769 3643 9493
rect 3757 8769 3803 9493
rect 3885 8769 3931 9493
rect 4045 8769 4091 9493
rect 4205 8769 4251 9493
rect 4365 8769 4411 9493
rect 4525 8769 4571 9493
rect 4685 8769 4731 9493
rect 4845 8769 4891 9493
rect 5005 8769 5051 9493
rect 5165 8769 5211 9493
rect 5293 8769 5339 9493
rect 5453 8769 5499 9493
rect 911 7659 957 8259
rect 1127 7659 1173 8259
rect 1343 7659 1389 8259
rect 1559 7659 1605 8259
rect 1775 7659 1821 8259
rect 1991 7659 2037 8259
rect 2207 7659 2253 8259
rect 2423 7659 2469 8259
rect 2639 7659 2685 8259
rect 2855 7659 2901 8259
rect 3071 7659 3117 8259
rect 3597 7639 3643 8363
rect 3757 7639 3803 8363
rect 3885 7639 3931 8363
rect 4045 7639 4091 8363
rect 4205 7639 4251 8363
rect 4365 7639 4411 8363
rect 4525 7639 4571 8363
rect 4685 7639 4731 8363
rect 4845 7639 4891 8363
rect 5005 7639 5051 8363
rect 5165 7639 5211 8363
rect 5293 7639 5339 8363
rect 5453 7639 5499 8363
rect 12079 10764 12125 11364
rect 12239 10764 12285 11364
rect 12367 10764 12413 11364
rect 12527 10764 12573 11364
rect 12655 10764 12701 11364
rect 12815 10764 12861 11364
rect 12975 10764 13021 11364
rect 13103 10764 13149 11364
rect 13263 10764 13309 11364
rect 13423 10764 13469 11364
rect 13551 10764 13597 11364
rect 13711 10764 13757 11364
rect 13871 10764 13917 11364
rect 13999 10764 14045 11364
rect 14159 10764 14205 11364
rect 14287 10764 14333 11364
rect 14447 10764 14493 11364
rect 14873 10764 14919 11364
rect 15033 10764 15079 11364
rect 15161 10764 15207 11364
rect 15321 10764 15367 11364
rect 15481 10764 15527 11364
rect 15641 10764 15687 11364
rect 15801 10764 15847 11364
rect 15961 10764 16007 11364
rect 16121 10764 16167 11364
rect 16281 10764 16327 11364
rect 16441 10764 16487 11364
rect 16569 10764 16615 11364
rect 16729 10764 16775 11364
rect 12079 9728 12125 10328
rect 12239 9728 12285 10328
rect 12367 9728 12413 10328
rect 12527 9728 12573 10328
rect 12655 9728 12701 10328
rect 12815 9728 12861 10328
rect 12975 9728 13021 10328
rect 13103 9728 13149 10328
rect 13263 9728 13309 10328
rect 13423 9728 13469 10328
rect 13551 9728 13597 10328
rect 13711 9728 13757 10328
rect 13871 9728 13917 10328
rect 13999 9728 14045 10328
rect 14159 9728 14205 10328
rect 14287 9728 14333 10328
rect 14447 9728 14493 10328
rect 14873 9728 14919 10328
rect 15033 9728 15079 10328
rect 15161 9728 15207 10328
rect 15321 9728 15367 10328
rect 15481 9728 15527 10328
rect 15641 9728 15687 10328
rect 15801 9728 15847 10328
rect 15961 9728 16007 10328
rect 16121 9728 16167 10328
rect 16281 9728 16327 10328
rect 16441 9728 16487 10328
rect 16569 9728 16615 10328
rect 16729 9728 16775 10328
rect 12079 8692 12125 9292
rect 12239 8692 12285 9292
rect 12367 8692 12413 9292
rect 12527 8692 12573 9292
rect 12655 8692 12701 9292
rect 12815 8692 12861 9292
rect 12975 8692 13021 9292
rect 13103 8692 13149 9292
rect 13263 8692 13309 9292
rect 13423 8692 13469 9292
rect 13551 8692 13597 9292
rect 13711 8692 13757 9292
rect 13871 8692 13917 9292
rect 13999 8692 14045 9292
rect 14159 8692 14205 9292
rect 14287 8692 14333 9292
rect 14447 8692 14493 9292
rect 14873 8692 14919 9292
rect 15033 8692 15079 9292
rect 15161 8692 15207 9292
rect 15321 8692 15367 9292
rect 15481 8692 15527 9292
rect 15641 8692 15687 9292
rect 15801 8692 15847 9292
rect 15961 8692 16007 9292
rect 16121 8692 16167 9292
rect 16281 8692 16327 9292
rect 16441 8692 16487 9292
rect 16569 8692 16615 9292
rect 16729 8692 16775 9292
rect 12079 7656 12125 8256
rect 12239 7656 12285 8256
rect 12367 7656 12413 8256
rect 12527 7656 12573 8256
rect 12655 7656 12701 8256
rect 12815 7656 12861 8256
rect 12975 7656 13021 8256
rect 13103 7656 13149 8256
rect 13263 7656 13309 8256
rect 13423 7656 13469 8256
rect 13551 7656 13597 8256
rect 13711 7656 13757 8256
rect 13871 7656 13917 8256
rect 13999 7656 14045 8256
rect 14159 7656 14205 8256
rect 14287 7656 14333 8256
rect 14447 7656 14493 8256
rect 14873 7656 14919 8256
rect 15033 7656 15079 8256
rect 15161 7656 15207 8256
rect 15321 7656 15367 8256
rect 15481 7656 15527 8256
rect 15641 7656 15687 8256
rect 15801 7656 15847 8256
rect 15961 7656 16007 8256
rect 16121 7656 16167 8256
rect 16281 7656 16327 8256
rect 16441 7656 16487 8256
rect 16569 7656 16615 8256
rect 16729 7656 16775 8256
rect 33129 11102 33175 11676
rect 33289 11102 33335 11676
rect 33417 11102 33463 11676
rect 33577 11102 33623 11676
rect 33737 11102 33783 11676
rect 33897 11102 33943 11676
rect 34057 11102 34103 11676
rect 34217 11102 34263 11676
rect 34377 11102 34423 11676
rect 34537 11102 34583 11676
rect 34697 11102 34743 11676
rect 34857 11102 34903 11676
rect 35017 11102 35063 11676
rect 35177 11102 35223 11676
rect 35337 11102 35383 11676
rect 35497 11102 35543 11676
rect 35657 11102 35703 11676
rect 35817 11102 35863 11676
rect 35977 11102 36023 11676
rect 36105 11102 36151 11676
rect 36265 11102 36311 11676
rect 37265 11102 37311 11676
rect 37425 11102 37471 11676
rect 37553 11102 37599 11676
rect 37713 11102 37759 11676
rect 37873 11102 37919 11676
rect 38033 11102 38079 11676
rect 38193 11102 38239 11676
rect 38353 11102 38399 11676
rect 38513 11102 38559 11676
rect 38673 11102 38719 11676
rect 38833 11102 38879 11676
rect 38993 11102 39039 11676
rect 39153 11102 39199 11676
rect 39313 11102 39359 11676
rect 39473 11102 39519 11676
rect 39633 11102 39679 11676
rect 39793 11102 39839 11676
rect 39953 11102 39999 11676
rect 40113 11102 40159 11676
rect 40241 11102 40287 11676
rect 40401 11102 40447 11676
rect 33129 10042 33175 10616
rect 33289 10042 33335 10616
rect 33417 10042 33463 10616
rect 33577 10042 33623 10616
rect 33737 10042 33783 10616
rect 33897 10042 33943 10616
rect 34057 10042 34103 10616
rect 34217 10042 34263 10616
rect 34377 10042 34423 10616
rect 34537 10042 34583 10616
rect 34697 10042 34743 10616
rect 34857 10042 34903 10616
rect 35017 10042 35063 10616
rect 35177 10042 35223 10616
rect 35337 10042 35383 10616
rect 35497 10042 35543 10616
rect 35657 10042 35703 10616
rect 35817 10042 35863 10616
rect 35977 10042 36023 10616
rect 36105 10042 36151 10616
rect 36265 10042 36311 10616
rect 37265 10042 37311 10616
rect 37425 10042 37471 10616
rect 37553 10042 37599 10616
rect 37713 10042 37759 10616
rect 37873 10042 37919 10616
rect 38033 10042 38079 10616
rect 38193 10042 38239 10616
rect 38353 10042 38399 10616
rect 38513 10042 38559 10616
rect 38673 10042 38719 10616
rect 38833 10042 38879 10616
rect 38993 10042 39039 10616
rect 39153 10042 39199 10616
rect 39313 10042 39359 10616
rect 39473 10042 39519 10616
rect 39633 10042 39679 10616
rect 39793 10042 39839 10616
rect 39953 10042 39999 10616
rect 40113 10042 40159 10616
rect 40241 10042 40287 10616
rect 40401 10042 40447 10616
rect 33129 8982 33175 9556
rect 33289 8982 33335 9556
rect 33417 8982 33463 9556
rect 33577 8982 33623 9556
rect 33737 8982 33783 9556
rect 33897 8982 33943 9556
rect 34057 8982 34103 9556
rect 34217 8982 34263 9556
rect 34377 8982 34423 9556
rect 34537 8982 34583 9556
rect 34697 8982 34743 9556
rect 34857 8982 34903 9556
rect 35017 8982 35063 9556
rect 35177 8982 35223 9556
rect 35337 8982 35383 9556
rect 35497 8982 35543 9556
rect 35657 8982 35703 9556
rect 35817 8982 35863 9556
rect 35977 8982 36023 9556
rect 36105 8982 36151 9556
rect 36265 8982 36311 9556
rect 37265 8982 37311 9556
rect 37425 8982 37471 9556
rect 37553 8982 37599 9556
rect 37713 8982 37759 9556
rect 37873 8982 37919 9556
rect 38033 8982 38079 9556
rect 38193 8982 38239 9556
rect 38353 8982 38399 9556
rect 38513 8982 38559 9556
rect 38673 8982 38719 9556
rect 38833 8982 38879 9556
rect 38993 8982 39039 9556
rect 39153 8982 39199 9556
rect 39313 8982 39359 9556
rect 39473 8982 39519 9556
rect 39633 8982 39679 9556
rect 39793 8982 39839 9556
rect 39953 8982 39999 9556
rect 40113 8982 40159 9556
rect 40241 8982 40287 9556
rect 40401 8982 40447 9556
rect 33129 7922 33175 8496
rect 33289 7922 33335 8496
rect 33417 7922 33463 8496
rect 33577 7922 33623 8496
rect 33737 7922 33783 8496
rect 33897 7922 33943 8496
rect 34057 7922 34103 8496
rect 34217 7922 34263 8496
rect 34377 7922 34423 8496
rect 34537 7922 34583 8496
rect 34697 7922 34743 8496
rect 34857 7922 34903 8496
rect 35017 7922 35063 8496
rect 35177 7922 35223 8496
rect 35337 7922 35383 8496
rect 35497 7922 35543 8496
rect 35657 7922 35703 8496
rect 35817 7922 35863 8496
rect 35977 7922 36023 8496
rect 36105 7922 36151 8496
rect 36265 7922 36311 8496
rect 37265 7922 37311 8496
rect 37425 7922 37471 8496
rect 37553 7922 37599 8496
rect 37713 7922 37759 8496
rect 37873 7922 37919 8496
rect 38033 7922 38079 8496
rect 38193 7922 38239 8496
rect 38353 7922 38399 8496
rect 38513 7922 38559 8496
rect 38673 7922 38719 8496
rect 38833 7922 38879 8496
rect 38993 7922 39039 8496
rect 39153 7922 39199 8496
rect 39313 7922 39359 8496
rect 39473 7922 39519 8496
rect 39633 7922 39679 8496
rect 39793 7922 39839 8496
rect 39953 7922 39999 8496
rect 40113 7922 40159 8496
rect 40241 7922 40287 8496
rect 40401 7922 40447 8496
rect 42825 11102 42871 11676
rect 42985 11102 43031 11676
rect 43113 11102 43159 11676
rect 43273 11102 43319 11676
rect 43433 11102 43479 11676
rect 43593 11102 43639 11676
rect 43753 11102 43799 11676
rect 43913 11102 43959 11676
rect 44073 11102 44119 11676
rect 44233 11102 44279 11676
rect 44393 11102 44439 11676
rect 44553 11102 44599 11676
rect 44713 11102 44759 11676
rect 44873 11102 44919 11676
rect 45033 11102 45079 11676
rect 45193 11102 45239 11676
rect 45353 11102 45399 11676
rect 45513 11102 45559 11676
rect 45673 11102 45719 11676
rect 45801 11102 45847 11676
rect 45961 11102 46007 11676
rect 46961 11102 47007 11676
rect 47121 11102 47167 11676
rect 47249 11102 47295 11676
rect 47409 11102 47455 11676
rect 47569 11102 47615 11676
rect 47729 11102 47775 11676
rect 47889 11102 47935 11676
rect 48049 11102 48095 11676
rect 48209 11102 48255 11676
rect 48369 11102 48415 11676
rect 48529 11102 48575 11676
rect 48689 11102 48735 11676
rect 48849 11102 48895 11676
rect 49009 11102 49055 11676
rect 49169 11102 49215 11676
rect 49329 11102 49375 11676
rect 49489 11102 49535 11676
rect 49649 11102 49695 11676
rect 49809 11102 49855 11676
rect 49937 11102 49983 11676
rect 50097 11102 50143 11676
rect 42825 10042 42871 10616
rect 42985 10042 43031 10616
rect 43113 10042 43159 10616
rect 43273 10042 43319 10616
rect 43433 10042 43479 10616
rect 43593 10042 43639 10616
rect 43753 10042 43799 10616
rect 43913 10042 43959 10616
rect 44073 10042 44119 10616
rect 44233 10042 44279 10616
rect 44393 10042 44439 10616
rect 44553 10042 44599 10616
rect 44713 10042 44759 10616
rect 44873 10042 44919 10616
rect 45033 10042 45079 10616
rect 45193 10042 45239 10616
rect 45353 10042 45399 10616
rect 45513 10042 45559 10616
rect 45673 10042 45719 10616
rect 45801 10042 45847 10616
rect 45961 10042 46007 10616
rect 46961 10042 47007 10616
rect 47121 10042 47167 10616
rect 47249 10042 47295 10616
rect 47409 10042 47455 10616
rect 47569 10042 47615 10616
rect 47729 10042 47775 10616
rect 47889 10042 47935 10616
rect 48049 10042 48095 10616
rect 48209 10042 48255 10616
rect 48369 10042 48415 10616
rect 48529 10042 48575 10616
rect 48689 10042 48735 10616
rect 48849 10042 48895 10616
rect 49009 10042 49055 10616
rect 49169 10042 49215 10616
rect 49329 10042 49375 10616
rect 49489 10042 49535 10616
rect 49649 10042 49695 10616
rect 49809 10042 49855 10616
rect 49937 10042 49983 10616
rect 50097 10042 50143 10616
rect 42825 8982 42871 9556
rect 42985 8982 43031 9556
rect 43113 8982 43159 9556
rect 43273 8982 43319 9556
rect 43433 8982 43479 9556
rect 43593 8982 43639 9556
rect 43753 8982 43799 9556
rect 43913 8982 43959 9556
rect 44073 8982 44119 9556
rect 44233 8982 44279 9556
rect 44393 8982 44439 9556
rect 44553 8982 44599 9556
rect 44713 8982 44759 9556
rect 44873 8982 44919 9556
rect 45033 8982 45079 9556
rect 45193 8982 45239 9556
rect 45353 8982 45399 9556
rect 45513 8982 45559 9556
rect 45673 8982 45719 9556
rect 45801 8982 45847 9556
rect 45961 8982 46007 9556
rect 46961 8982 47007 9556
rect 47121 8982 47167 9556
rect 47249 8982 47295 9556
rect 47409 8982 47455 9556
rect 47569 8982 47615 9556
rect 47729 8982 47775 9556
rect 47889 8982 47935 9556
rect 48049 8982 48095 9556
rect 48209 8982 48255 9556
rect 48369 8982 48415 9556
rect 48529 8982 48575 9556
rect 48689 8982 48735 9556
rect 48849 8982 48895 9556
rect 49009 8982 49055 9556
rect 49169 8982 49215 9556
rect 49329 8982 49375 9556
rect 49489 8982 49535 9556
rect 49649 8982 49695 9556
rect 49809 8982 49855 9556
rect 49937 8982 49983 9556
rect 50097 8982 50143 9556
rect 42825 7922 42871 8496
rect 42985 7922 43031 8496
rect 43113 7922 43159 8496
rect 43273 7922 43319 8496
rect 43433 7922 43479 8496
rect 43593 7922 43639 8496
rect 43753 7922 43799 8496
rect 43913 7922 43959 8496
rect 44073 7922 44119 8496
rect 44233 7922 44279 8496
rect 44393 7922 44439 8496
rect 44553 7922 44599 8496
rect 44713 7922 44759 8496
rect 44873 7922 44919 8496
rect 45033 7922 45079 8496
rect 45193 7922 45239 8496
rect 45353 7922 45399 8496
rect 45513 7922 45559 8496
rect 45673 7922 45719 8496
rect 45801 7922 45847 8496
rect 45961 7922 46007 8496
rect 46961 7922 47007 8496
rect 47121 7922 47167 8496
rect 47249 7922 47295 8496
rect 47409 7922 47455 8496
rect 47569 7922 47615 8496
rect 47729 7922 47775 8496
rect 47889 7922 47935 8496
rect 48049 7922 48095 8496
rect 48209 7922 48255 8496
rect 48369 7922 48415 8496
rect 48529 7922 48575 8496
rect 48689 7922 48735 8496
rect 48849 7922 48895 8496
rect 49009 7922 49055 8496
rect 49169 7922 49215 8496
rect 49329 7922 49375 8496
rect 49489 7922 49535 8496
rect 49649 7922 49695 8496
rect 49809 7922 49855 8496
rect 49937 7922 49983 8496
rect 50097 7922 50143 8496
rect 52521 11102 52567 11676
rect 52681 11102 52727 11676
rect 52809 11102 52855 11676
rect 52969 11102 53015 11676
rect 53129 11102 53175 11676
rect 53289 11102 53335 11676
rect 53449 11102 53495 11676
rect 53609 11102 53655 11676
rect 53769 11102 53815 11676
rect 53929 11102 53975 11676
rect 54089 11102 54135 11676
rect 54249 11102 54295 11676
rect 54409 11102 54455 11676
rect 54569 11102 54615 11676
rect 54729 11102 54775 11676
rect 54889 11102 54935 11676
rect 55049 11102 55095 11676
rect 55209 11102 55255 11676
rect 55369 11102 55415 11676
rect 55497 11102 55543 11676
rect 55657 11102 55703 11676
rect 56657 11102 56703 11676
rect 56817 11102 56863 11676
rect 56945 11102 56991 11676
rect 57105 11102 57151 11676
rect 57265 11102 57311 11676
rect 57425 11102 57471 11676
rect 57585 11102 57631 11676
rect 57745 11102 57791 11676
rect 57905 11102 57951 11676
rect 58065 11102 58111 11676
rect 58225 11102 58271 11676
rect 58385 11102 58431 11676
rect 58545 11102 58591 11676
rect 58705 11102 58751 11676
rect 58865 11102 58911 11676
rect 59025 11102 59071 11676
rect 59185 11102 59231 11676
rect 59345 11102 59391 11676
rect 59505 11102 59551 11676
rect 59633 11102 59679 11676
rect 59793 11102 59839 11676
rect 52521 10042 52567 10616
rect 52681 10042 52727 10616
rect 52809 10042 52855 10616
rect 52969 10042 53015 10616
rect 53129 10042 53175 10616
rect 53289 10042 53335 10616
rect 53449 10042 53495 10616
rect 53609 10042 53655 10616
rect 53769 10042 53815 10616
rect 53929 10042 53975 10616
rect 54089 10042 54135 10616
rect 54249 10042 54295 10616
rect 54409 10042 54455 10616
rect 54569 10042 54615 10616
rect 54729 10042 54775 10616
rect 54889 10042 54935 10616
rect 55049 10042 55095 10616
rect 55209 10042 55255 10616
rect 55369 10042 55415 10616
rect 55497 10042 55543 10616
rect 55657 10042 55703 10616
rect 56657 10042 56703 10616
rect 56817 10042 56863 10616
rect 56945 10042 56991 10616
rect 57105 10042 57151 10616
rect 57265 10042 57311 10616
rect 57425 10042 57471 10616
rect 57585 10042 57631 10616
rect 57745 10042 57791 10616
rect 57905 10042 57951 10616
rect 58065 10042 58111 10616
rect 58225 10042 58271 10616
rect 58385 10042 58431 10616
rect 58545 10042 58591 10616
rect 58705 10042 58751 10616
rect 58865 10042 58911 10616
rect 59025 10042 59071 10616
rect 59185 10042 59231 10616
rect 59345 10042 59391 10616
rect 59505 10042 59551 10616
rect 59633 10042 59679 10616
rect 59793 10042 59839 10616
rect 52521 8982 52567 9556
rect 52681 8982 52727 9556
rect 52809 8982 52855 9556
rect 52969 8982 53015 9556
rect 53129 8982 53175 9556
rect 53289 8982 53335 9556
rect 53449 8982 53495 9556
rect 53609 8982 53655 9556
rect 53769 8982 53815 9556
rect 53929 8982 53975 9556
rect 54089 8982 54135 9556
rect 54249 8982 54295 9556
rect 54409 8982 54455 9556
rect 54569 8982 54615 9556
rect 54729 8982 54775 9556
rect 54889 8982 54935 9556
rect 55049 8982 55095 9556
rect 55209 8982 55255 9556
rect 55369 8982 55415 9556
rect 55497 8982 55543 9556
rect 55657 8982 55703 9556
rect 56657 8982 56703 9556
rect 56817 8982 56863 9556
rect 56945 8982 56991 9556
rect 57105 8982 57151 9556
rect 57265 8982 57311 9556
rect 57425 8982 57471 9556
rect 57585 8982 57631 9556
rect 57745 8982 57791 9556
rect 57905 8982 57951 9556
rect 58065 8982 58111 9556
rect 58225 8982 58271 9556
rect 58385 8982 58431 9556
rect 58545 8982 58591 9556
rect 58705 8982 58751 9556
rect 58865 8982 58911 9556
rect 59025 8982 59071 9556
rect 59185 8982 59231 9556
rect 59345 8982 59391 9556
rect 59505 8982 59551 9556
rect 59633 8982 59679 9556
rect 59793 8982 59839 9556
rect 52521 7922 52567 8496
rect 52681 7922 52727 8496
rect 52809 7922 52855 8496
rect 52969 7922 53015 8496
rect 53129 7922 53175 8496
rect 53289 7922 53335 8496
rect 53449 7922 53495 8496
rect 53609 7922 53655 8496
rect 53769 7922 53815 8496
rect 53929 7922 53975 8496
rect 54089 7922 54135 8496
rect 54249 7922 54295 8496
rect 54409 7922 54455 8496
rect 54569 7922 54615 8496
rect 54729 7922 54775 8496
rect 54889 7922 54935 8496
rect 55049 7922 55095 8496
rect 55209 7922 55255 8496
rect 55369 7922 55415 8496
rect 55497 7922 55543 8496
rect 55657 7922 55703 8496
rect 56657 7922 56703 8496
rect 56817 7922 56863 8496
rect 56945 7922 56991 8496
rect 57105 7922 57151 8496
rect 57265 7922 57311 8496
rect 57425 7922 57471 8496
rect 57585 7922 57631 8496
rect 57745 7922 57791 8496
rect 57905 7922 57951 8496
rect 58065 7922 58111 8496
rect 58225 7922 58271 8496
rect 58385 7922 58431 8496
rect 58545 7922 58591 8496
rect 58705 7922 58751 8496
rect 58865 7922 58911 8496
rect 59025 7922 59071 8496
rect 59185 7922 59231 8496
rect 59345 7922 59391 8496
rect 59505 7922 59551 8496
rect 59633 7922 59679 8496
rect 59793 7922 59839 8496
rect 62217 11102 62263 11676
rect 62377 11102 62423 11676
rect 62505 11102 62551 11676
rect 62665 11102 62711 11676
rect 62825 11102 62871 11676
rect 62985 11102 63031 11676
rect 63145 11102 63191 11676
rect 63305 11102 63351 11676
rect 63465 11102 63511 11676
rect 63625 11102 63671 11676
rect 63785 11102 63831 11676
rect 63945 11102 63991 11676
rect 64105 11102 64151 11676
rect 64265 11102 64311 11676
rect 64425 11102 64471 11676
rect 64585 11102 64631 11676
rect 64745 11102 64791 11676
rect 64905 11102 64951 11676
rect 65065 11102 65111 11676
rect 65193 11102 65239 11676
rect 65353 11102 65399 11676
rect 62217 10042 62263 10616
rect 62377 10042 62423 10616
rect 62505 10042 62551 10616
rect 62665 10042 62711 10616
rect 62825 10042 62871 10616
rect 62985 10042 63031 10616
rect 63145 10042 63191 10616
rect 63305 10042 63351 10616
rect 63465 10042 63511 10616
rect 63625 10042 63671 10616
rect 63785 10042 63831 10616
rect 63945 10042 63991 10616
rect 64105 10042 64151 10616
rect 64265 10042 64311 10616
rect 64425 10042 64471 10616
rect 64585 10042 64631 10616
rect 64745 10042 64791 10616
rect 64905 10042 64951 10616
rect 65065 10042 65111 10616
rect 65193 10042 65239 10616
rect 65353 10042 65399 10616
rect 62217 8982 62263 9556
rect 62377 8982 62423 9556
rect 62505 8982 62551 9556
rect 62665 8982 62711 9556
rect 62825 8982 62871 9556
rect 62985 8982 63031 9556
rect 63145 8982 63191 9556
rect 63305 8982 63351 9556
rect 63465 8982 63511 9556
rect 63625 8982 63671 9556
rect 63785 8982 63831 9556
rect 63945 8982 63991 9556
rect 64105 8982 64151 9556
rect 64265 8982 64311 9556
rect 64425 8982 64471 9556
rect 64585 8982 64631 9556
rect 64745 8982 64791 9556
rect 64905 8982 64951 9556
rect 65065 8982 65111 9556
rect 65193 8982 65239 9556
rect 65353 8982 65399 9556
rect 62217 7922 62263 8496
rect 62377 7922 62423 8496
rect 62505 7922 62551 8496
rect 62665 7922 62711 8496
rect 62825 7922 62871 8496
rect 62985 7922 63031 8496
rect 63145 7922 63191 8496
rect 63305 7922 63351 8496
rect 63465 7922 63511 8496
rect 63625 7922 63671 8496
rect 63785 7922 63831 8496
rect 63945 7922 63991 8496
rect 64105 7922 64151 8496
rect 64265 7922 64311 8496
rect 64425 7922 64471 8496
rect 64585 7922 64631 8496
rect 64745 7922 64791 8496
rect 64905 7922 64951 8496
rect 65065 7922 65111 8496
rect 65193 7922 65239 8496
rect 65353 7922 65399 8496
rect 1290 3647 1336 4421
rect 1450 3647 1496 4421
rect 1578 3647 1624 4421
rect 1738 3647 1784 4421
rect 1866 3647 1912 4421
rect 2082 3647 2128 4421
rect 2298 3647 2344 4421
rect 2514 3647 2560 4421
rect 2730 3647 2776 4421
rect 2946 3647 2992 4421
rect 3162 3647 3208 4421
rect 3378 3647 3424 4421
rect 3594 3647 3640 4421
rect 3810 3647 3856 4421
rect 4026 3647 4072 4421
rect 4242 3647 4288 4421
rect 4402 3647 4448 4421
rect 4562 3647 4608 4421
rect 1290 2387 1336 3161
rect 1450 2387 1496 3161
rect 1586 2387 1632 3161
rect 1746 2387 1792 3161
rect 1874 2387 1920 3161
rect 2090 2387 2136 3161
rect 2306 2387 2352 3161
rect 2522 2387 2568 3161
rect 2738 2387 2784 3161
rect 2954 2387 3000 3161
rect 3114 2387 3160 3161
rect 3274 2387 3320 3161
rect 3434 2387 3480 3161
rect 3594 2387 3640 3161
rect 3810 2387 3856 3161
rect 3938 2387 3984 3161
rect 4154 2387 4200 3161
rect 4314 2387 4360 3161
rect 4450 2387 4496 3161
rect 4610 2387 4656 3161
rect 1290 1827 1336 1901
rect 1450 1827 1496 1901
rect 1586 1827 1632 1901
rect 1746 1827 1792 1901
rect 1906 1827 1952 1901
rect 2066 1827 2112 1901
rect 2226 1827 2272 1901
rect 2386 1827 2432 1901
rect 2546 1827 2592 1901
rect 2706 1827 2752 1901
rect 2866 1827 2912 1901
rect 3026 1827 3072 1901
rect 3186 1827 3232 1901
rect 3346 1827 3392 1901
rect 3506 1827 3552 1901
rect 3666 1827 3712 1901
rect 3826 1827 3872 1901
rect 3986 1827 4032 1901
rect 4146 1827 4192 1901
rect 4450 1827 4496 1901
rect 4610 1827 4656 1901
rect 18795 4192 18841 4766
rect 18955 4192 19001 4766
rect 19115 4192 19161 4766
rect 19275 4192 19321 4766
rect 19435 4192 19481 4766
rect 19595 4192 19641 4766
rect 19755 4192 19801 4766
rect 19915 4192 19961 4766
rect 20075 4192 20121 4766
rect 20235 4192 20281 4766
rect 20395 4192 20441 4766
rect 20555 4192 20601 4766
rect 20715 4192 20761 4766
rect 20875 4192 20921 4766
rect 21035 4192 21081 4766
rect 21195 4192 21241 4766
rect 21355 4192 21401 4766
rect 21515 4192 21561 4766
rect 21675 4192 21721 4766
rect 21835 4192 21881 4766
rect 21963 4192 22009 4766
rect 22123 4192 22169 4766
rect 22251 4192 22297 4766
rect 22411 4192 22457 4766
rect 18795 3456 18841 4030
rect 18955 3456 19001 4030
rect 19115 3456 19161 4030
rect 19275 3456 19321 4030
rect 19435 3456 19481 4030
rect 19595 3456 19641 4030
rect 19755 3456 19801 4030
rect 19915 3456 19961 4030
rect 20075 3456 20121 4030
rect 20235 3456 20281 4030
rect 20395 3456 20441 4030
rect 20555 3456 20601 4030
rect 20715 3456 20761 4030
rect 20875 3456 20921 4030
rect 21035 3456 21081 4030
rect 21195 3456 21241 4030
rect 21355 3456 21401 4030
rect 21515 3456 21561 4030
rect 21675 3456 21721 4030
rect 21835 3456 21881 4030
rect 21963 3456 22009 4030
rect 22123 3456 22169 4030
rect 22251 3456 22297 4030
rect 22411 3456 22457 4030
rect 18795 2720 18841 3294
rect 18955 2720 19001 3294
rect 19115 2720 19161 3294
rect 19275 2720 19321 3294
rect 19435 2720 19481 3294
rect 19595 2720 19641 3294
rect 19755 2720 19801 3294
rect 19915 2720 19961 3294
rect 20075 2720 20121 3294
rect 20235 2720 20281 3294
rect 20395 2720 20441 3294
rect 20555 2720 20601 3294
rect 20715 2720 20761 3294
rect 20875 2720 20921 3294
rect 21035 2720 21081 3294
rect 21195 2720 21241 3294
rect 21355 2720 21401 3294
rect 21515 2720 21561 3294
rect 21675 2720 21721 3294
rect 21835 2720 21881 3294
rect 21963 2720 22009 3194
rect 22123 2720 22169 3194
rect 22251 2720 22297 3294
rect 22411 2720 22457 3294
rect 18795 1984 18841 2558
rect 18955 1984 19001 2558
rect 19115 1984 19161 2558
rect 19275 1984 19321 2558
rect 19435 1984 19481 2558
rect 19595 1984 19641 2558
rect 19755 1984 19801 2558
rect 19915 1984 19961 2558
rect 20075 1984 20121 2558
rect 20235 1984 20281 2558
rect 20395 1984 20441 2558
rect 20555 1984 20601 2558
rect 20715 1984 20761 2558
rect 20875 1984 20921 2558
rect 21035 1984 21081 2558
rect 21195 1984 21241 2558
rect 21355 1984 21401 2558
rect 21515 1984 21561 2558
rect 21675 1984 21721 2558
rect 21835 1984 21881 2558
rect 21963 1984 22009 2458
rect 22123 1984 22169 2458
rect 22251 1984 22297 2558
rect 22411 1984 22457 2558
<< psubdiff >>
rect 6249 14665 8577 14678
rect 6249 14619 6262 14665
rect 6308 14619 6356 14665
rect 6402 14619 6450 14665
rect 6496 14619 6544 14665
rect 6590 14619 6638 14665
rect 6684 14619 6732 14665
rect 6778 14619 6826 14665
rect 6872 14619 6920 14665
rect 6966 14619 7014 14665
rect 7060 14619 7108 14665
rect 7154 14619 7202 14665
rect 7248 14619 7296 14665
rect 7342 14619 7390 14665
rect 7436 14619 7484 14665
rect 7530 14619 7578 14665
rect 7624 14619 7672 14665
rect 7718 14619 7766 14665
rect 7812 14619 7860 14665
rect 7906 14619 7954 14665
rect 8000 14619 8048 14665
rect 8094 14619 8142 14665
rect 8188 14619 8236 14665
rect 8282 14619 8330 14665
rect 8376 14619 8424 14665
rect 8470 14619 8518 14665
rect 8564 14619 8577 14665
rect 6249 14606 8577 14619
rect 6249 14571 6321 14606
rect 6249 14525 6262 14571
rect 6308 14525 6321 14571
rect 6249 14477 6321 14525
rect 6249 14431 6262 14477
rect 6308 14431 6321 14477
rect 6249 14383 6321 14431
rect 6249 14337 6262 14383
rect 6308 14337 6321 14383
rect 6249 14289 6321 14337
rect 8505 14571 8577 14606
rect 8505 14525 8518 14571
rect 8564 14525 8577 14571
rect 8505 14477 8577 14525
rect 8505 14431 8518 14477
rect 8564 14431 8577 14477
rect 8505 14383 8577 14431
rect 8505 14337 8518 14383
rect 8564 14337 8577 14383
rect 6249 14243 6262 14289
rect 6308 14243 6321 14289
rect 8505 14289 8577 14337
rect 6249 14195 6321 14243
rect 6249 14149 6262 14195
rect 6308 14149 6321 14195
rect 6249 14101 6321 14149
rect 6249 14055 6262 14101
rect 6308 14055 6321 14101
rect 6249 14007 6321 14055
rect 6249 13961 6262 14007
rect 6308 13961 6321 14007
rect 6249 13913 6321 13961
rect 6249 13867 6262 13913
rect 6308 13867 6321 13913
rect 6249 13819 6321 13867
rect 6249 13773 6262 13819
rect 6308 13773 6321 13819
rect 6249 13725 6321 13773
rect 6249 13679 6262 13725
rect 6308 13679 6321 13725
rect 8505 14243 8518 14289
rect 8564 14243 8577 14289
rect 8505 14195 8577 14243
rect 8505 14149 8518 14195
rect 8564 14149 8577 14195
rect 8505 14101 8577 14149
rect 8505 14055 8518 14101
rect 8564 14055 8577 14101
rect 8505 14007 8577 14055
rect 8505 13961 8518 14007
rect 8564 13961 8577 14007
rect 8505 13913 8577 13961
rect 8505 13867 8518 13913
rect 8564 13867 8577 13913
rect 8505 13819 8577 13867
rect 8505 13773 8518 13819
rect 8564 13773 8577 13819
rect 8505 13725 8577 13773
rect 6249 13631 6321 13679
rect 6249 13585 6262 13631
rect 6308 13585 6321 13631
rect 6249 13537 6321 13585
rect 6249 13491 6262 13537
rect 6308 13491 6321 13537
rect 6249 13443 6321 13491
rect 6249 13397 6262 13443
rect 6308 13397 6321 13443
rect 8505 13679 8518 13725
rect 8564 13679 8577 13725
rect 8505 13631 8577 13679
rect 8505 13585 8518 13631
rect 8564 13585 8577 13631
rect 8505 13537 8577 13585
rect 8505 13491 8518 13537
rect 8564 13491 8577 13537
rect 8505 13443 8577 13491
rect 6249 13349 6321 13397
rect 6249 13303 6262 13349
rect 6308 13303 6321 13349
rect 6249 13255 6321 13303
rect 6249 13209 6262 13255
rect 6308 13209 6321 13255
rect 6249 13161 6321 13209
rect 6249 13115 6262 13161
rect 6308 13115 6321 13161
rect 6249 13067 6321 13115
rect 6249 13021 6262 13067
rect 6308 13021 6321 13067
rect 6249 12973 6321 13021
rect 6249 12927 6262 12973
rect 6308 12927 6321 12973
rect 6249 12879 6321 12927
rect 6249 12833 6262 12879
rect 6308 12833 6321 12879
rect 8505 13397 8518 13443
rect 8564 13397 8577 13443
rect 8505 13349 8577 13397
rect 8505 13303 8518 13349
rect 8564 13303 8577 13349
rect 8505 13255 8577 13303
rect 8505 13209 8518 13255
rect 8564 13209 8577 13255
rect 8505 13161 8577 13209
rect 8505 13115 8518 13161
rect 8564 13115 8577 13161
rect 8505 13067 8577 13115
rect 8505 13021 8518 13067
rect 8564 13021 8577 13067
rect 8505 12973 8577 13021
rect 8505 12927 8518 12973
rect 8564 12927 8577 12973
rect 8505 12879 8577 12927
rect 6249 12785 6321 12833
rect 6249 12739 6262 12785
rect 6308 12739 6321 12785
rect 6249 12691 6321 12739
rect 6249 12645 6262 12691
rect 6308 12645 6321 12691
rect 6249 12597 6321 12645
rect 6249 12551 6262 12597
rect 6308 12551 6321 12597
rect 8505 12833 8518 12879
rect 8564 12833 8577 12879
rect 8505 12785 8577 12833
rect 8505 12739 8518 12785
rect 8564 12739 8577 12785
rect 8505 12691 8577 12739
rect 8505 12645 8518 12691
rect 8564 12645 8577 12691
rect 8505 12597 8577 12645
rect 6249 12503 6321 12551
rect 6249 12448 6262 12503
rect 6308 12448 6321 12503
rect 6249 12400 6321 12448
rect 6249 12354 6262 12400
rect 6308 12354 6321 12400
rect 6249 12306 6321 12354
rect 6249 12260 6262 12306
rect 6308 12260 6321 12306
rect 6249 12212 6321 12260
rect 6249 12166 6262 12212
rect 6308 12166 6321 12212
rect 6249 12118 6321 12166
rect 6249 12072 6262 12118
rect 6308 12072 6321 12118
rect 6249 12024 6321 12072
rect 6249 11978 6262 12024
rect 6308 11978 6321 12024
rect 6249 11930 6321 11978
rect 8505 12551 8518 12597
rect 8564 12551 8577 12597
rect 8505 12503 8577 12551
rect 8505 12448 8518 12503
rect 8564 12448 8577 12503
rect 8505 12400 8577 12448
rect 8505 12354 8518 12400
rect 8564 12354 8577 12400
rect 8505 12306 8577 12354
rect 8505 12260 8518 12306
rect 8564 12260 8577 12306
rect 8505 12212 8577 12260
rect 8505 12166 8518 12212
rect 8564 12166 8577 12212
rect 8505 12118 8577 12166
rect 8505 12072 8518 12118
rect 8564 12072 8577 12118
rect 8505 12024 8577 12072
rect 8505 11978 8518 12024
rect 8564 11978 8577 12024
rect 6249 11884 6262 11930
rect 6308 11884 6321 11930
rect 6249 11836 6321 11884
rect 6249 11790 6262 11836
rect 6308 11790 6321 11836
rect 6249 11742 6321 11790
rect 6249 11696 6262 11742
rect 6308 11696 6321 11742
rect 6249 11648 6321 11696
rect 8505 11930 8577 11978
rect 8505 11884 8518 11930
rect 8564 11884 8577 11930
rect 8505 11836 8577 11884
rect 8505 11790 8518 11836
rect 8564 11790 8577 11836
rect 8505 11742 8577 11790
rect 18123 13768 21203 13781
rect 18123 13722 18136 13768
rect 18182 13722 18230 13768
rect 18276 13722 18324 13768
rect 18370 13722 18418 13768
rect 18464 13722 18512 13768
rect 18558 13722 18606 13768
rect 18652 13722 18700 13768
rect 18746 13722 18794 13768
rect 18840 13722 18888 13768
rect 18934 13722 18982 13768
rect 19028 13722 19076 13768
rect 19122 13722 19170 13768
rect 19216 13722 19264 13768
rect 19310 13722 19358 13768
rect 19404 13722 19452 13768
rect 19498 13722 19546 13768
rect 19592 13722 19640 13768
rect 19686 13722 19734 13768
rect 19780 13722 19828 13768
rect 19874 13722 19922 13768
rect 19968 13722 20016 13768
rect 20062 13722 20110 13768
rect 20156 13722 20204 13768
rect 20250 13722 20298 13768
rect 20344 13722 20392 13768
rect 20438 13722 20486 13768
rect 20532 13722 20580 13768
rect 20626 13722 20674 13768
rect 20720 13722 20768 13768
rect 20814 13722 20862 13768
rect 20908 13722 20956 13768
rect 21002 13722 21050 13768
rect 21096 13722 21144 13768
rect 21190 13722 21203 13768
rect 18123 13709 21203 13722
rect 18123 13674 18195 13709
rect 18123 13628 18136 13674
rect 18182 13628 18195 13674
rect 18123 13580 18195 13628
rect 18123 13534 18136 13580
rect 18182 13534 18195 13580
rect 18123 13486 18195 13534
rect 18123 13440 18136 13486
rect 18182 13440 18195 13486
rect 18123 13392 18195 13440
rect 21131 13674 21203 13709
rect 21131 13628 21144 13674
rect 21190 13628 21203 13674
rect 21131 13580 21203 13628
rect 21131 13534 21144 13580
rect 21190 13534 21203 13580
rect 21131 13486 21203 13534
rect 21131 13440 21144 13486
rect 21190 13440 21203 13486
rect 18123 13346 18136 13392
rect 18182 13346 18195 13392
rect 18123 13298 18195 13346
rect 21131 13392 21203 13440
rect 21131 13346 21144 13392
rect 21190 13346 21203 13392
rect 18123 13252 18136 13298
rect 18182 13252 18195 13298
rect 18123 13204 18195 13252
rect 18123 13158 18136 13204
rect 18182 13158 18195 13204
rect 21131 13298 21203 13346
rect 21131 13252 21144 13298
rect 21190 13252 21203 13298
rect 21131 13204 21203 13252
rect 18123 13110 18195 13158
rect 18123 13064 18136 13110
rect 18182 13064 18195 13110
rect 18123 13016 18195 13064
rect 18123 12970 18136 13016
rect 18182 12970 18195 13016
rect 18123 12922 18195 12970
rect 18123 12876 18136 12922
rect 18182 12876 18195 12922
rect 18123 12828 18195 12876
rect 18123 12782 18136 12828
rect 18182 12782 18195 12828
rect 18123 12734 18195 12782
rect 18123 12688 18136 12734
rect 18182 12688 18195 12734
rect 18123 12640 18195 12688
rect 18123 12594 18136 12640
rect 18182 12594 18195 12640
rect 18123 12546 18195 12594
rect 21131 13158 21144 13204
rect 21190 13158 21203 13204
rect 21131 13110 21203 13158
rect 21131 13064 21144 13110
rect 21190 13064 21203 13110
rect 21131 13016 21203 13064
rect 21131 12970 21144 13016
rect 21190 12970 21203 13016
rect 21131 12922 21203 12970
rect 21131 12876 21144 12922
rect 21190 12876 21203 12922
rect 21131 12828 21203 12876
rect 21131 12782 21144 12828
rect 21190 12782 21203 12828
rect 21131 12734 21203 12782
rect 21131 12688 21144 12734
rect 21190 12688 21203 12734
rect 21131 12640 21203 12688
rect 21131 12594 21144 12640
rect 21190 12594 21203 12640
rect 18123 12500 18136 12546
rect 18182 12500 18195 12546
rect 18123 12452 18195 12500
rect 18123 12406 18136 12452
rect 18182 12406 18195 12452
rect 18123 12358 18195 12406
rect 21131 12546 21203 12594
rect 21131 12500 21144 12546
rect 21190 12500 21203 12546
rect 18123 12312 18136 12358
rect 18182 12312 18195 12358
rect 18123 12264 18195 12312
rect 18123 12218 18136 12264
rect 18182 12218 18195 12264
rect 21131 12452 21203 12500
rect 21131 12406 21144 12452
rect 21190 12406 21203 12452
rect 21131 12358 21203 12406
rect 21131 12312 21144 12358
rect 21190 12312 21203 12358
rect 21131 12264 21203 12312
rect 18123 12170 18195 12218
rect 18123 12124 18136 12170
rect 18182 12124 18195 12170
rect 18123 12076 18195 12124
rect 18123 12030 18136 12076
rect 18182 12030 18195 12076
rect 18123 11982 18195 12030
rect 18123 11936 18136 11982
rect 18182 11936 18195 11982
rect 18123 11888 18195 11936
rect 18123 11842 18136 11888
rect 18182 11842 18195 11888
rect 18123 11794 18195 11842
rect 8505 11696 8518 11742
rect 8564 11696 8577 11742
rect 6249 11602 6262 11648
rect 6308 11602 6321 11648
rect 6249 11554 6321 11602
rect 6249 11508 6262 11554
rect 6308 11508 6321 11554
rect 6249 11460 6321 11508
rect 6249 11414 6262 11460
rect 6308 11414 6321 11460
rect 6249 11366 6321 11414
rect 6249 11320 6262 11366
rect 6308 11320 6321 11366
rect 6249 11272 6321 11320
rect 6249 11226 6262 11272
rect 6308 11226 6321 11272
rect 6249 11178 6321 11226
rect 6249 11132 6262 11178
rect 6308 11132 6321 11178
rect 6249 11084 6321 11132
rect 8505 11648 8577 11696
rect 8505 11602 8518 11648
rect 8564 11602 8577 11648
rect 8505 11554 8577 11602
rect 8505 11508 8518 11554
rect 8564 11508 8577 11554
rect 8505 11460 8577 11508
rect 8505 11414 8518 11460
rect 8564 11414 8577 11460
rect 8505 11366 8577 11414
rect 8505 11320 8518 11366
rect 8564 11320 8577 11366
rect 8505 11272 8577 11320
rect 8505 11226 8518 11272
rect 8564 11226 8577 11272
rect 8505 11191 8577 11226
rect 8505 11178 11303 11191
rect 8505 11132 8518 11178
rect 8564 11132 8612 11178
rect 8658 11132 8706 11178
rect 8752 11132 8800 11178
rect 8846 11132 8894 11178
rect 8940 11132 8988 11178
rect 9034 11132 9082 11178
rect 9128 11132 9176 11178
rect 9222 11132 9270 11178
rect 9316 11132 9364 11178
rect 9410 11132 9458 11178
rect 9504 11132 9552 11178
rect 9598 11132 9646 11178
rect 9692 11132 9740 11178
rect 9786 11132 9834 11178
rect 9880 11132 9928 11178
rect 9974 11132 10022 11178
rect 10068 11132 10116 11178
rect 10162 11132 10210 11178
rect 10256 11132 10304 11178
rect 10350 11132 10398 11178
rect 10444 11132 10492 11178
rect 10538 11132 10586 11178
rect 10632 11132 10680 11178
rect 10726 11132 10774 11178
rect 10820 11132 10868 11178
rect 10914 11132 10962 11178
rect 11008 11132 11056 11178
rect 11102 11132 11150 11178
rect 11196 11132 11244 11178
rect 11290 11132 11303 11178
rect 8505 11119 11303 11132
rect 6249 11038 6262 11084
rect 6308 11038 6321 11084
rect 6249 10990 6321 11038
rect 6249 10944 6262 10990
rect 6308 10944 6321 10990
rect 6249 10896 6321 10944
rect 6249 10850 6262 10896
rect 6308 10850 6321 10896
rect 6249 10802 6321 10850
rect 8505 11084 8577 11119
rect 8505 11038 8518 11084
rect 8564 11038 8577 11084
rect 8505 10990 8577 11038
rect 8505 10944 8518 10990
rect 8564 10944 8577 10990
rect 8505 10896 8577 10944
rect 8505 10850 8518 10896
rect 8564 10850 8577 10896
rect 11231 11084 11303 11119
rect 11231 11038 11244 11084
rect 11290 11038 11303 11084
rect 11231 10990 11303 11038
rect 11231 10944 11244 10990
rect 11290 10944 11303 10990
rect 11231 10896 11303 10944
rect 6249 10756 6262 10802
rect 6308 10756 6321 10802
rect 6249 10708 6321 10756
rect 6249 10662 6262 10708
rect 6308 10662 6321 10708
rect 6249 10614 6321 10662
rect 6249 10568 6262 10614
rect 6308 10568 6321 10614
rect 6249 10520 6321 10568
rect 6249 10474 6262 10520
rect 6308 10474 6321 10520
rect 6249 10426 6321 10474
rect 6249 10380 6262 10426
rect 6308 10380 6321 10426
rect 6249 10332 6321 10380
rect 6249 10286 6262 10332
rect 6308 10286 6321 10332
rect 6249 10238 6321 10286
rect 8505 10802 8577 10850
rect 11231 10850 11244 10896
rect 11290 10850 11303 10896
rect 8505 10756 8518 10802
rect 8564 10756 8577 10802
rect 8505 10708 8577 10756
rect 8505 10662 8518 10708
rect 8564 10662 8577 10708
rect 8505 10614 8577 10662
rect 8505 10568 8518 10614
rect 8564 10568 8577 10614
rect 8505 10520 8577 10568
rect 8505 10474 8518 10520
rect 8564 10474 8577 10520
rect 8505 10426 8577 10474
rect 8505 10380 8518 10426
rect 8564 10380 8577 10426
rect 8505 10332 8577 10380
rect 8505 10286 8518 10332
rect 8564 10286 8577 10332
rect 6249 10192 6262 10238
rect 6308 10192 6321 10238
rect 6249 10144 6321 10192
rect 6249 10098 6262 10144
rect 6308 10098 6321 10144
rect 6249 10050 6321 10098
rect 6249 10004 6262 10050
rect 6308 10004 6321 10050
rect 6249 9956 6321 10004
rect 8505 10238 8577 10286
rect 8505 10192 8518 10238
rect 8564 10192 8577 10238
rect 11231 10802 11303 10850
rect 11231 10756 11244 10802
rect 11290 10756 11303 10802
rect 11231 10708 11303 10756
rect 11231 10662 11244 10708
rect 11290 10662 11303 10708
rect 11231 10614 11303 10662
rect 11231 10568 11244 10614
rect 11290 10568 11303 10614
rect 11231 10520 11303 10568
rect 11231 10474 11244 10520
rect 11290 10474 11303 10520
rect 11231 10426 11303 10474
rect 11231 10380 11244 10426
rect 11290 10380 11303 10426
rect 11231 10332 11303 10380
rect 11231 10286 11244 10332
rect 11290 10286 11303 10332
rect 11231 10238 11303 10286
rect 8505 10144 8577 10192
rect 8505 10098 8518 10144
rect 8564 10098 8577 10144
rect 8505 10050 8577 10098
rect 8505 10004 8518 10050
rect 8564 10004 8577 10050
rect 6249 9910 6262 9956
rect 6308 9910 6321 9956
rect 6249 9862 6321 9910
rect 6249 9816 6262 9862
rect 6308 9816 6321 9862
rect 6249 9768 6321 9816
rect 6249 9722 6262 9768
rect 6308 9722 6321 9768
rect 6249 9674 6321 9722
rect 6249 9628 6262 9674
rect 6308 9628 6321 9674
rect 6249 9580 6321 9628
rect 6249 9534 6262 9580
rect 6308 9534 6321 9580
rect 6249 9486 6321 9534
rect 6249 9440 6262 9486
rect 6308 9440 6321 9486
rect 6249 9392 6321 9440
rect 6249 9346 6262 9392
rect 6308 9346 6321 9392
rect 8505 9956 8577 10004
rect 8505 9910 8518 9956
rect 8564 9910 8577 9956
rect 11231 10192 11244 10238
rect 11290 10192 11303 10238
rect 11231 10144 11303 10192
rect 11231 10098 11244 10144
rect 11290 10098 11303 10144
rect 11231 10050 11303 10098
rect 11231 10004 11244 10050
rect 11290 10004 11303 10050
rect 11231 9956 11303 10004
rect 8505 9862 8577 9910
rect 8505 9816 8518 9862
rect 8564 9816 8577 9862
rect 8505 9768 8577 9816
rect 8505 9722 8518 9768
rect 8564 9722 8577 9768
rect 8505 9674 8577 9722
rect 8505 9628 8518 9674
rect 8564 9628 8577 9674
rect 8505 9580 8577 9628
rect 8505 9534 8518 9580
rect 8564 9534 8577 9580
rect 8505 9486 8577 9534
rect 8505 9440 8518 9486
rect 8564 9440 8577 9486
rect 8505 9392 8577 9440
rect 6249 9298 6321 9346
rect 6249 9252 6262 9298
rect 6308 9252 6321 9298
rect 6249 9204 6321 9252
rect 6249 9158 6262 9204
rect 6308 9158 6321 9204
rect 6249 9110 6321 9158
rect 6249 9064 6262 9110
rect 6308 9064 6321 9110
rect 8505 9346 8518 9392
rect 8564 9346 8577 9392
rect 11231 9910 11244 9956
rect 11290 9910 11303 9956
rect 11231 9862 11303 9910
rect 11231 9816 11244 9862
rect 11290 9816 11303 9862
rect 11231 9768 11303 9816
rect 11231 9722 11244 9768
rect 11290 9722 11303 9768
rect 11231 9674 11303 9722
rect 11231 9628 11244 9674
rect 11290 9628 11303 9674
rect 11231 9580 11303 9628
rect 11231 9534 11244 9580
rect 11290 9534 11303 9580
rect 11231 9486 11303 9534
rect 11231 9440 11244 9486
rect 11290 9440 11303 9486
rect 11231 9392 11303 9440
rect 8505 9298 8577 9346
rect 8505 9252 8518 9298
rect 8564 9252 8577 9298
rect 8505 9204 8577 9252
rect 8505 9158 8518 9204
rect 8564 9158 8577 9204
rect 8505 9110 8577 9158
rect 6249 9016 6321 9064
rect 6249 8970 6262 9016
rect 6308 8970 6321 9016
rect 6249 8922 6321 8970
rect 6249 8876 6262 8922
rect 6308 8876 6321 8922
rect 6249 8828 6321 8876
rect 6249 8782 6262 8828
rect 6308 8782 6321 8828
rect 6249 8734 6321 8782
rect 6249 8688 6262 8734
rect 6308 8688 6321 8734
rect 6249 8640 6321 8688
rect 6249 8594 6262 8640
rect 6308 8594 6321 8640
rect 6249 8546 6321 8594
rect 6249 8500 6262 8546
rect 6308 8500 6321 8546
rect 8505 9064 8518 9110
rect 8564 9064 8577 9110
rect 11231 9346 11244 9392
rect 11290 9346 11303 9392
rect 11231 9298 11303 9346
rect 11231 9252 11244 9298
rect 11290 9252 11303 9298
rect 11231 9204 11303 9252
rect 11231 9158 11244 9204
rect 11290 9158 11303 9204
rect 11231 9110 11303 9158
rect 8505 9016 8577 9064
rect 8505 8970 8518 9016
rect 8564 8970 8577 9016
rect 8505 8922 8577 8970
rect 8505 8876 8518 8922
rect 8564 8876 8577 8922
rect 8505 8828 8577 8876
rect 8505 8782 8518 8828
rect 8564 8782 8577 8828
rect 8505 8734 8577 8782
rect 8505 8688 8518 8734
rect 8564 8688 8577 8734
rect 8505 8640 8577 8688
rect 8505 8594 8518 8640
rect 8564 8594 8577 8640
rect 8505 8546 8577 8594
rect 6249 8452 6321 8500
rect 6249 8406 6262 8452
rect 6308 8406 6321 8452
rect 6249 8358 6321 8406
rect 6249 8312 6262 8358
rect 6308 8312 6321 8358
rect 8505 8500 8518 8546
rect 8564 8500 8577 8546
rect 11231 9064 11244 9110
rect 11290 9064 11303 9110
rect 11231 9016 11303 9064
rect 11231 8970 11244 9016
rect 11290 8970 11303 9016
rect 11231 8922 11303 8970
rect 11231 8876 11244 8922
rect 11290 8876 11303 8922
rect 11231 8828 11303 8876
rect 11231 8782 11244 8828
rect 11290 8782 11303 8828
rect 11231 8734 11303 8782
rect 11231 8688 11244 8734
rect 11290 8688 11303 8734
rect 11231 8640 11303 8688
rect 11231 8594 11244 8640
rect 11290 8594 11303 8640
rect 11231 8546 11303 8594
rect 8505 8452 8577 8500
rect 6249 8264 6321 8312
rect 6249 8218 6262 8264
rect 6308 8218 6321 8264
rect 8505 8406 8518 8452
rect 8564 8406 8577 8452
rect 8505 8358 8577 8406
rect 8505 8312 8518 8358
rect 8564 8312 8577 8358
rect 11231 8500 11244 8546
rect 11290 8500 11303 8546
rect 11231 8452 11303 8500
rect 11231 8406 11244 8452
rect 11290 8406 11303 8452
rect 8505 8264 8577 8312
rect 6249 8170 6321 8218
rect 6249 8124 6262 8170
rect 6308 8124 6321 8170
rect 6249 8076 6321 8124
rect 6249 8030 6262 8076
rect 6308 8030 6321 8076
rect 6249 7982 6321 8030
rect 6249 7936 6262 7982
rect 6308 7936 6321 7982
rect 6249 7888 6321 7936
rect 6249 7842 6262 7888
rect 6308 7842 6321 7888
rect 6249 7794 6321 7842
rect 6249 7748 6262 7794
rect 6308 7748 6321 7794
rect 6249 7700 6321 7748
rect 6249 7654 6262 7700
rect 6308 7654 6321 7700
rect 8505 8218 8518 8264
rect 8564 8218 8577 8264
rect 11231 8358 11303 8406
rect 11231 8312 11244 8358
rect 11290 8312 11303 8358
rect 11231 8264 11303 8312
rect 8505 8170 8577 8218
rect 8505 8124 8518 8170
rect 8564 8124 8577 8170
rect 8505 8076 8577 8124
rect 8505 8030 8518 8076
rect 8564 8030 8577 8076
rect 8505 7982 8577 8030
rect 8505 7936 8518 7982
rect 8564 7936 8577 7982
rect 8505 7888 8577 7936
rect 8505 7842 8518 7888
rect 8564 7842 8577 7888
rect 8505 7794 8577 7842
rect 8505 7748 8518 7794
rect 8564 7748 8577 7794
rect 8505 7700 8577 7748
rect 6249 7606 6321 7654
rect 8505 7654 8518 7700
rect 8564 7654 8577 7700
rect 6249 7560 6262 7606
rect 6308 7560 6321 7606
rect 6249 7512 6321 7560
rect 6249 7466 6262 7512
rect 6308 7466 6321 7512
rect 6249 7418 6321 7466
rect 6249 7372 6262 7418
rect 6308 7372 6321 7418
rect 6249 7337 6321 7372
rect 8505 7606 8577 7654
rect 11231 8218 11244 8264
rect 11290 8218 11303 8264
rect 11231 8170 11303 8218
rect 11231 8124 11244 8170
rect 11290 8124 11303 8170
rect 11231 8076 11303 8124
rect 11231 8030 11244 8076
rect 11290 8030 11303 8076
rect 11231 7982 11303 8030
rect 11231 7936 11244 7982
rect 11290 7936 11303 7982
rect 11231 7888 11303 7936
rect 11231 7842 11244 7888
rect 11290 7842 11303 7888
rect 11231 7794 11303 7842
rect 11231 7748 11244 7794
rect 11290 7748 11303 7794
rect 11231 7700 11303 7748
rect 11231 7654 11244 7700
rect 11290 7654 11303 7700
rect 8505 7560 8518 7606
rect 8564 7560 8577 7606
rect 11231 7606 11303 7654
rect 8505 7512 8577 7560
rect 8505 7466 8518 7512
rect 8564 7466 8577 7512
rect 8505 7418 8577 7466
rect 8505 7372 8518 7418
rect 8564 7372 8577 7418
rect 8505 7337 8577 7372
rect 11231 7560 11244 7606
rect 11290 7560 11303 7606
rect 11231 7512 11303 7560
rect 11231 7466 11244 7512
rect 11290 7466 11303 7512
rect 11231 7418 11303 7466
rect 11231 7372 11244 7418
rect 11290 7372 11303 7418
rect 11231 7337 11303 7372
rect 6249 7324 11303 7337
rect 6249 7278 6262 7324
rect 6308 7278 6356 7324
rect 6402 7278 6450 7324
rect 6496 7278 6544 7324
rect 6590 7278 6638 7324
rect 6684 7278 6732 7324
rect 6778 7278 6826 7324
rect 6872 7278 6920 7324
rect 6966 7278 7014 7324
rect 7060 7278 7108 7324
rect 7154 7278 7202 7324
rect 7248 7278 7296 7324
rect 7342 7278 7390 7324
rect 7436 7278 7484 7324
rect 7530 7278 7578 7324
rect 7624 7278 7672 7324
rect 7718 7278 7766 7324
rect 7812 7278 7860 7324
rect 7906 7278 7954 7324
rect 8000 7278 8048 7324
rect 8094 7278 8142 7324
rect 8188 7278 8236 7324
rect 8282 7278 8330 7324
rect 8376 7278 8424 7324
rect 8470 7278 8518 7324
rect 8564 7278 8612 7324
rect 8658 7278 8706 7324
rect 8752 7278 8800 7324
rect 8846 7278 8894 7324
rect 8940 7278 8988 7324
rect 9034 7278 9082 7324
rect 9128 7278 9176 7324
rect 9222 7278 9270 7324
rect 9316 7278 9364 7324
rect 9410 7278 9458 7324
rect 9504 7278 9552 7324
rect 9598 7278 9646 7324
rect 9692 7278 9740 7324
rect 9786 7278 9834 7324
rect 9880 7278 9928 7324
rect 9974 7278 10022 7324
rect 10068 7278 10116 7324
rect 10162 7278 10210 7324
rect 10256 7278 10304 7324
rect 10350 7278 10398 7324
rect 10444 7278 10492 7324
rect 10538 7278 10586 7324
rect 10632 7278 10680 7324
rect 10726 7278 10774 7324
rect 10820 7278 10868 7324
rect 10914 7278 10962 7324
rect 11008 7278 11056 7324
rect 11102 7278 11150 7324
rect 11196 7278 11244 7324
rect 11290 7278 11303 7324
rect 6249 7265 11303 7278
rect 18123 11748 18136 11794
rect 18182 11748 18195 11794
rect 18123 11700 18195 11748
rect 18123 11654 18136 11700
rect 18182 11654 18195 11700
rect 18123 11606 18195 11654
rect 21131 12218 21144 12264
rect 21190 12218 21203 12264
rect 21131 12170 21203 12218
rect 21131 12124 21144 12170
rect 21190 12124 21203 12170
rect 21131 12076 21203 12124
rect 21131 12030 21144 12076
rect 21190 12030 21203 12076
rect 21131 11982 21203 12030
rect 21131 11936 21144 11982
rect 21190 11936 21203 11982
rect 21131 11888 21203 11936
rect 21131 11842 21144 11888
rect 21190 11842 21203 11888
rect 21131 11794 21203 11842
rect 21131 11748 21144 11794
rect 21190 11748 21203 11794
rect 21131 11700 21203 11748
rect 21131 11654 21144 11700
rect 21190 11654 21203 11700
rect 18123 11560 18136 11606
rect 18182 11560 18195 11606
rect 18123 11512 18195 11560
rect 18123 11466 18136 11512
rect 18182 11466 18195 11512
rect 18123 11418 18195 11466
rect 18123 11372 18136 11418
rect 18182 11372 18195 11418
rect 18123 11324 18195 11372
rect 18123 11278 18136 11324
rect 18182 11278 18195 11324
rect 21131 11606 21203 11654
rect 21131 11560 21144 11606
rect 21190 11560 21203 11606
rect 21131 11512 21203 11560
rect 21131 11466 21144 11512
rect 21190 11466 21203 11512
rect 21131 11418 21203 11466
rect 21131 11372 21144 11418
rect 21190 11372 21203 11418
rect 21131 11324 21203 11372
rect 18123 11230 18195 11278
rect 18123 11184 18136 11230
rect 18182 11184 18195 11230
rect 18123 11136 18195 11184
rect 18123 11090 18136 11136
rect 18182 11090 18195 11136
rect 18123 11042 18195 11090
rect 18123 10996 18136 11042
rect 18182 10996 18195 11042
rect 18123 10948 18195 10996
rect 18123 10902 18136 10948
rect 18182 10902 18195 10948
rect 18123 10854 18195 10902
rect 18123 10808 18136 10854
rect 18182 10808 18195 10854
rect 18123 10760 18195 10808
rect 18123 10714 18136 10760
rect 18182 10714 18195 10760
rect 21131 11278 21144 11324
rect 21190 11278 21203 11324
rect 21131 11230 21203 11278
rect 21131 11184 21144 11230
rect 21190 11184 21203 11230
rect 21131 11136 21203 11184
rect 21131 11090 21144 11136
rect 21190 11090 21203 11136
rect 21131 11042 21203 11090
rect 21131 10996 21144 11042
rect 21190 10996 21203 11042
rect 21131 10948 21203 10996
rect 21131 10902 21144 10948
rect 21190 10902 21203 10948
rect 21131 10854 21203 10902
rect 21131 10808 21144 10854
rect 21190 10808 21203 10854
rect 21131 10760 21203 10808
rect 18123 10666 18195 10714
rect 18123 10620 18136 10666
rect 18182 10620 18195 10666
rect 18123 10572 18195 10620
rect 18123 10526 18136 10572
rect 18182 10526 18195 10572
rect 18123 10478 18195 10526
rect 18123 10432 18136 10478
rect 18182 10432 18195 10478
rect 18123 10384 18195 10432
rect 18123 10338 18136 10384
rect 18182 10338 18195 10384
rect 21131 10714 21144 10760
rect 21190 10714 21203 10760
rect 21131 10666 21203 10714
rect 21131 10620 21144 10666
rect 21190 10620 21203 10666
rect 21131 10572 21203 10620
rect 21131 10526 21144 10572
rect 21190 10526 21203 10572
rect 21131 10478 21203 10526
rect 21131 10432 21144 10478
rect 21190 10432 21203 10478
rect 21131 10384 21203 10432
rect 18123 10290 18195 10338
rect 18123 10244 18136 10290
rect 18182 10244 18195 10290
rect 18123 10196 18195 10244
rect 18123 10150 18136 10196
rect 18182 10150 18195 10196
rect 18123 10102 18195 10150
rect 18123 10056 18136 10102
rect 18182 10056 18195 10102
rect 18123 10008 18195 10056
rect 18123 9962 18136 10008
rect 18182 9962 18195 10008
rect 18123 9914 18195 9962
rect 18123 9868 18136 9914
rect 18182 9868 18195 9914
rect 18123 9820 18195 9868
rect 18123 9774 18136 9820
rect 18182 9774 18195 9820
rect 21131 10338 21144 10384
rect 21190 10338 21203 10384
rect 21131 10290 21203 10338
rect 21131 10244 21144 10290
rect 21190 10244 21203 10290
rect 21131 10196 21203 10244
rect 21131 10150 21144 10196
rect 21190 10150 21203 10196
rect 21131 10102 21203 10150
rect 21131 10056 21144 10102
rect 21190 10056 21203 10102
rect 21131 10008 21203 10056
rect 21131 9962 21144 10008
rect 21190 9962 21203 10008
rect 21131 9914 21203 9962
rect 21131 9868 21144 9914
rect 21190 9868 21203 9914
rect 21131 9820 21203 9868
rect 18123 9726 18195 9774
rect 18123 9680 18136 9726
rect 18182 9680 18195 9726
rect 18123 9632 18195 9680
rect 18123 9586 18136 9632
rect 18182 9586 18195 9632
rect 18123 9538 18195 9586
rect 18123 9492 18136 9538
rect 18182 9492 18195 9538
rect 18123 9444 18195 9492
rect 21131 9774 21144 9820
rect 21190 9774 21203 9820
rect 21131 9726 21203 9774
rect 21131 9680 21144 9726
rect 21190 9680 21203 9726
rect 21131 9632 21203 9680
rect 21131 9586 21144 9632
rect 21190 9586 21203 9632
rect 21131 9538 21203 9586
rect 21131 9492 21144 9538
rect 21190 9492 21203 9538
rect 18123 9398 18136 9444
rect 18182 9398 18195 9444
rect 18123 9350 18195 9398
rect 18123 9304 18136 9350
rect 18182 9304 18195 9350
rect 18123 9256 18195 9304
rect 18123 9210 18136 9256
rect 18182 9210 18195 9256
rect 18123 9162 18195 9210
rect 18123 9116 18136 9162
rect 18182 9116 18195 9162
rect 18123 9068 18195 9116
rect 18123 9022 18136 9068
rect 18182 9022 18195 9068
rect 18123 8974 18195 9022
rect 18123 8928 18136 8974
rect 18182 8928 18195 8974
rect 18123 8880 18195 8928
rect 18123 8834 18136 8880
rect 18182 8834 18195 8880
rect 21131 9444 21203 9492
rect 21131 9398 21144 9444
rect 21190 9398 21203 9444
rect 21131 9350 21203 9398
rect 21131 9304 21144 9350
rect 21190 9304 21203 9350
rect 21131 9256 21203 9304
rect 21131 9210 21144 9256
rect 21190 9210 21203 9256
rect 21131 9162 21203 9210
rect 21131 9116 21144 9162
rect 21190 9116 21203 9162
rect 21131 9068 21203 9116
rect 21131 9022 21144 9068
rect 21190 9022 21203 9068
rect 21131 8974 21203 9022
rect 21131 8928 21144 8974
rect 21190 8928 21203 8974
rect 21131 8880 21203 8928
rect 18123 8786 18195 8834
rect 18123 8740 18136 8786
rect 18182 8740 18195 8786
rect 18123 8692 18195 8740
rect 18123 8646 18136 8692
rect 18182 8646 18195 8692
rect 18123 8598 18195 8646
rect 21131 8834 21144 8880
rect 21190 8834 21203 8880
rect 21131 8786 21203 8834
rect 21131 8740 21144 8786
rect 21190 8740 21203 8786
rect 18123 8552 18136 8598
rect 18182 8552 18195 8598
rect 18123 8504 18195 8552
rect 21131 8692 21203 8740
rect 21131 8646 21144 8692
rect 21190 8646 21203 8692
rect 21131 8598 21203 8646
rect 21131 8552 21144 8598
rect 21190 8552 21203 8598
rect 18123 8458 18136 8504
rect 18182 8458 18195 8504
rect 18123 8410 18195 8458
rect 18123 8364 18136 8410
rect 18182 8364 18195 8410
rect 18123 8316 18195 8364
rect 18123 8270 18136 8316
rect 18182 8270 18195 8316
rect 18123 8222 18195 8270
rect 18123 8176 18136 8222
rect 18182 8176 18195 8222
rect 18123 8128 18195 8176
rect 18123 8082 18136 8128
rect 18182 8082 18195 8128
rect 18123 8034 18195 8082
rect 18123 7988 18136 8034
rect 18182 7988 18195 8034
rect 18123 7940 18195 7988
rect 18123 7894 18136 7940
rect 18182 7894 18195 7940
rect 21131 8504 21203 8552
rect 21131 8458 21144 8504
rect 21190 8458 21203 8504
rect 21131 8410 21203 8458
rect 21131 8364 21144 8410
rect 21190 8364 21203 8410
rect 21131 8316 21203 8364
rect 21131 8270 21144 8316
rect 21190 8270 21203 8316
rect 21131 8222 21203 8270
rect 21131 8176 21144 8222
rect 21190 8176 21203 8222
rect 21131 8128 21203 8176
rect 21131 8082 21144 8128
rect 21190 8082 21203 8128
rect 21131 8034 21203 8082
rect 21131 7988 21144 8034
rect 21190 7988 21203 8034
rect 21131 7940 21203 7988
rect 18123 7846 18195 7894
rect 18123 7800 18136 7846
rect 18182 7800 18195 7846
rect 18123 7752 18195 7800
rect 21131 7894 21144 7940
rect 21190 7894 21203 7940
rect 21131 7846 21203 7894
rect 21131 7800 21144 7846
rect 21190 7800 21203 7846
rect 18123 7706 18136 7752
rect 18182 7706 18195 7752
rect 18123 7658 18195 7706
rect 21131 7752 21203 7800
rect 21131 7706 21144 7752
rect 21190 7706 21203 7752
rect 18123 7612 18136 7658
rect 18182 7612 18195 7658
rect 18123 7564 18195 7612
rect 18123 7518 18136 7564
rect 18182 7518 18195 7564
rect 18123 7470 18195 7518
rect 18123 7424 18136 7470
rect 18182 7424 18195 7470
rect 18123 7389 18195 7424
rect 21131 7658 21203 7706
rect 21131 7612 21144 7658
rect 21190 7612 21203 7658
rect 21131 7564 21203 7612
rect 21131 7518 21144 7564
rect 21190 7518 21203 7564
rect 21131 7470 21203 7518
rect 21131 7424 21144 7470
rect 21190 7424 21203 7470
rect 21131 7389 21203 7424
rect 18123 7376 21203 7389
rect 18123 7330 18136 7376
rect 18182 7330 18230 7376
rect 18276 7330 18324 7376
rect 18370 7330 18418 7376
rect 18464 7330 18512 7376
rect 18558 7330 18606 7376
rect 18652 7330 18700 7376
rect 18746 7330 18794 7376
rect 18840 7330 18888 7376
rect 18934 7330 18982 7376
rect 19028 7330 19076 7376
rect 19122 7330 19170 7376
rect 19216 7330 19264 7376
rect 19310 7330 19358 7376
rect 19404 7330 19452 7376
rect 19498 7330 19546 7376
rect 19592 7330 19640 7376
rect 19686 7330 19734 7376
rect 19780 7330 19828 7376
rect 19874 7330 19922 7376
rect 19968 7330 20016 7376
rect 20062 7330 20110 7376
rect 20156 7330 20204 7376
rect 20250 7330 20298 7376
rect 20344 7330 20392 7376
rect 20438 7330 20486 7376
rect 20532 7330 20580 7376
rect 20626 7330 20674 7376
rect 20720 7330 20768 7376
rect 20814 7330 20862 7376
rect 20908 7330 20956 7376
rect 21002 7330 21050 7376
rect 21096 7330 21144 7376
rect 21190 7330 21203 7376
rect 18123 7317 21203 7330
rect 23275 13768 26355 13781
rect 23275 13722 23288 13768
rect 23334 13722 23382 13768
rect 23428 13722 23476 13768
rect 23522 13722 23570 13768
rect 23616 13722 23664 13768
rect 23710 13722 23758 13768
rect 23804 13722 23852 13768
rect 23898 13722 23946 13768
rect 23992 13722 24040 13768
rect 24086 13722 24134 13768
rect 24180 13722 24228 13768
rect 24274 13722 24322 13768
rect 24368 13722 24416 13768
rect 24462 13722 24510 13768
rect 24556 13722 24604 13768
rect 24650 13722 24698 13768
rect 24744 13722 24792 13768
rect 24838 13722 24886 13768
rect 24932 13722 24980 13768
rect 25026 13722 25074 13768
rect 25120 13722 25168 13768
rect 25214 13722 25262 13768
rect 25308 13722 25356 13768
rect 25402 13722 25450 13768
rect 25496 13722 25544 13768
rect 25590 13722 25638 13768
rect 25684 13722 25732 13768
rect 25778 13722 25826 13768
rect 25872 13722 25920 13768
rect 25966 13722 26014 13768
rect 26060 13722 26108 13768
rect 26154 13722 26202 13768
rect 26248 13722 26296 13768
rect 26342 13722 26355 13768
rect 23275 13709 26355 13722
rect 23275 13674 23347 13709
rect 23275 13628 23288 13674
rect 23334 13628 23347 13674
rect 23275 13580 23347 13628
rect 23275 13534 23288 13580
rect 23334 13534 23347 13580
rect 23275 13486 23347 13534
rect 23275 13440 23288 13486
rect 23334 13440 23347 13486
rect 23275 13392 23347 13440
rect 26283 13674 26355 13709
rect 26283 13628 26296 13674
rect 26342 13628 26355 13674
rect 26283 13580 26355 13628
rect 26283 13534 26296 13580
rect 26342 13534 26355 13580
rect 26283 13486 26355 13534
rect 26283 13440 26296 13486
rect 26342 13440 26355 13486
rect 23275 13346 23288 13392
rect 23334 13346 23347 13392
rect 23275 13298 23347 13346
rect 26283 13392 26355 13440
rect 26283 13346 26296 13392
rect 26342 13346 26355 13392
rect 23275 13252 23288 13298
rect 23334 13252 23347 13298
rect 23275 13204 23347 13252
rect 23275 13158 23288 13204
rect 23334 13158 23347 13204
rect 26283 13298 26355 13346
rect 26283 13252 26296 13298
rect 26342 13252 26355 13298
rect 26283 13204 26355 13252
rect 23275 13110 23347 13158
rect 23275 13064 23288 13110
rect 23334 13064 23347 13110
rect 23275 13016 23347 13064
rect 23275 12970 23288 13016
rect 23334 12970 23347 13016
rect 23275 12922 23347 12970
rect 23275 12876 23288 12922
rect 23334 12876 23347 12922
rect 23275 12828 23347 12876
rect 23275 12782 23288 12828
rect 23334 12782 23347 12828
rect 23275 12734 23347 12782
rect 23275 12688 23288 12734
rect 23334 12688 23347 12734
rect 23275 12640 23347 12688
rect 23275 12594 23288 12640
rect 23334 12594 23347 12640
rect 23275 12546 23347 12594
rect 26283 13158 26296 13204
rect 26342 13158 26355 13204
rect 26283 13110 26355 13158
rect 26283 13064 26296 13110
rect 26342 13064 26355 13110
rect 26283 13016 26355 13064
rect 26283 12970 26296 13016
rect 26342 12970 26355 13016
rect 26283 12922 26355 12970
rect 26283 12876 26296 12922
rect 26342 12876 26355 12922
rect 26283 12828 26355 12876
rect 26283 12782 26296 12828
rect 26342 12782 26355 12828
rect 26283 12734 26355 12782
rect 26283 12688 26296 12734
rect 26342 12688 26355 12734
rect 26283 12640 26355 12688
rect 26283 12594 26296 12640
rect 26342 12594 26355 12640
rect 23275 12500 23288 12546
rect 23334 12500 23347 12546
rect 23275 12452 23347 12500
rect 23275 12406 23288 12452
rect 23334 12406 23347 12452
rect 23275 12358 23347 12406
rect 26283 12546 26355 12594
rect 26283 12500 26296 12546
rect 26342 12500 26355 12546
rect 23275 12312 23288 12358
rect 23334 12312 23347 12358
rect 23275 12264 23347 12312
rect 23275 12218 23288 12264
rect 23334 12218 23347 12264
rect 26283 12452 26355 12500
rect 26283 12406 26296 12452
rect 26342 12406 26355 12452
rect 26283 12358 26355 12406
rect 26283 12312 26296 12358
rect 26342 12312 26355 12358
rect 26283 12264 26355 12312
rect 23275 12170 23347 12218
rect 23275 12124 23288 12170
rect 23334 12124 23347 12170
rect 23275 12076 23347 12124
rect 23275 12030 23288 12076
rect 23334 12030 23347 12076
rect 23275 11982 23347 12030
rect 23275 11936 23288 11982
rect 23334 11936 23347 11982
rect 23275 11888 23347 11936
rect 23275 11842 23288 11888
rect 23334 11842 23347 11888
rect 23275 11794 23347 11842
rect 23275 11748 23288 11794
rect 23334 11748 23347 11794
rect 23275 11700 23347 11748
rect 23275 11654 23288 11700
rect 23334 11654 23347 11700
rect 23275 11606 23347 11654
rect 26283 12218 26296 12264
rect 26342 12218 26355 12264
rect 26283 12170 26355 12218
rect 26283 12124 26296 12170
rect 26342 12124 26355 12170
rect 26283 12076 26355 12124
rect 26283 12030 26296 12076
rect 26342 12030 26355 12076
rect 26283 11982 26355 12030
rect 26283 11936 26296 11982
rect 26342 11936 26355 11982
rect 26283 11888 26355 11936
rect 26283 11842 26296 11888
rect 26342 11842 26355 11888
rect 26283 11794 26355 11842
rect 26283 11748 26296 11794
rect 26342 11748 26355 11794
rect 26283 11700 26355 11748
rect 26283 11654 26296 11700
rect 26342 11654 26355 11700
rect 23275 11560 23288 11606
rect 23334 11560 23347 11606
rect 23275 11512 23347 11560
rect 23275 11466 23288 11512
rect 23334 11466 23347 11512
rect 23275 11418 23347 11466
rect 23275 11372 23288 11418
rect 23334 11372 23347 11418
rect 23275 11324 23347 11372
rect 23275 11278 23288 11324
rect 23334 11278 23347 11324
rect 26283 11606 26355 11654
rect 26283 11560 26296 11606
rect 26342 11560 26355 11606
rect 26283 11512 26355 11560
rect 26283 11466 26296 11512
rect 26342 11466 26355 11512
rect 26283 11418 26355 11466
rect 26283 11372 26296 11418
rect 26342 11372 26355 11418
rect 26283 11324 26355 11372
rect 23275 11230 23347 11278
rect 23275 11184 23288 11230
rect 23334 11184 23347 11230
rect 23275 11136 23347 11184
rect 23275 11090 23288 11136
rect 23334 11090 23347 11136
rect 23275 11042 23347 11090
rect 23275 10996 23288 11042
rect 23334 10996 23347 11042
rect 23275 10948 23347 10996
rect 23275 10902 23288 10948
rect 23334 10902 23347 10948
rect 23275 10854 23347 10902
rect 23275 10808 23288 10854
rect 23334 10808 23347 10854
rect 23275 10760 23347 10808
rect 23275 10714 23288 10760
rect 23334 10714 23347 10760
rect 26283 11278 26296 11324
rect 26342 11278 26355 11324
rect 26283 11230 26355 11278
rect 26283 11184 26296 11230
rect 26342 11184 26355 11230
rect 26283 11136 26355 11184
rect 26283 11090 26296 11136
rect 26342 11090 26355 11136
rect 26283 11042 26355 11090
rect 26283 10996 26296 11042
rect 26342 10996 26355 11042
rect 26283 10948 26355 10996
rect 26283 10902 26296 10948
rect 26342 10902 26355 10948
rect 26283 10854 26355 10902
rect 26283 10808 26296 10854
rect 26342 10808 26355 10854
rect 26283 10760 26355 10808
rect 23275 10666 23347 10714
rect 23275 10620 23288 10666
rect 23334 10620 23347 10666
rect 23275 10572 23347 10620
rect 23275 10526 23288 10572
rect 23334 10526 23347 10572
rect 23275 10478 23347 10526
rect 23275 10432 23288 10478
rect 23334 10432 23347 10478
rect 23275 10384 23347 10432
rect 23275 10338 23288 10384
rect 23334 10338 23347 10384
rect 26283 10714 26296 10760
rect 26342 10714 26355 10760
rect 26283 10666 26355 10714
rect 26283 10620 26296 10666
rect 26342 10620 26355 10666
rect 26283 10572 26355 10620
rect 26283 10526 26296 10572
rect 26342 10526 26355 10572
rect 26283 10478 26355 10526
rect 26283 10432 26296 10478
rect 26342 10432 26355 10478
rect 26283 10384 26355 10432
rect 23275 10290 23347 10338
rect 23275 10244 23288 10290
rect 23334 10244 23347 10290
rect 23275 10196 23347 10244
rect 23275 10150 23288 10196
rect 23334 10150 23347 10196
rect 23275 10102 23347 10150
rect 23275 10056 23288 10102
rect 23334 10056 23347 10102
rect 23275 10008 23347 10056
rect 23275 9962 23288 10008
rect 23334 9962 23347 10008
rect 23275 9914 23347 9962
rect 23275 9868 23288 9914
rect 23334 9868 23347 9914
rect 23275 9820 23347 9868
rect 23275 9774 23288 9820
rect 23334 9774 23347 9820
rect 26283 10338 26296 10384
rect 26342 10338 26355 10384
rect 26283 10290 26355 10338
rect 26283 10244 26296 10290
rect 26342 10244 26355 10290
rect 26283 10196 26355 10244
rect 26283 10150 26296 10196
rect 26342 10150 26355 10196
rect 26283 10102 26355 10150
rect 26283 10056 26296 10102
rect 26342 10056 26355 10102
rect 26283 10008 26355 10056
rect 26283 9962 26296 10008
rect 26342 9962 26355 10008
rect 26283 9914 26355 9962
rect 26283 9868 26296 9914
rect 26342 9868 26355 9914
rect 26283 9820 26355 9868
rect 23275 9726 23347 9774
rect 23275 9680 23288 9726
rect 23334 9680 23347 9726
rect 23275 9632 23347 9680
rect 23275 9586 23288 9632
rect 23334 9586 23347 9632
rect 23275 9538 23347 9586
rect 23275 9492 23288 9538
rect 23334 9492 23347 9538
rect 23275 9444 23347 9492
rect 26283 9774 26296 9820
rect 26342 9774 26355 9820
rect 26283 9726 26355 9774
rect 26283 9680 26296 9726
rect 26342 9680 26355 9726
rect 26283 9632 26355 9680
rect 26283 9586 26296 9632
rect 26342 9586 26355 9632
rect 26283 9538 26355 9586
rect 26283 9492 26296 9538
rect 26342 9492 26355 9538
rect 23275 9398 23288 9444
rect 23334 9398 23347 9444
rect 23275 9350 23347 9398
rect 23275 9304 23288 9350
rect 23334 9304 23347 9350
rect 23275 9256 23347 9304
rect 23275 9210 23288 9256
rect 23334 9210 23347 9256
rect 23275 9162 23347 9210
rect 23275 9116 23288 9162
rect 23334 9116 23347 9162
rect 23275 9068 23347 9116
rect 23275 9022 23288 9068
rect 23334 9022 23347 9068
rect 23275 8974 23347 9022
rect 23275 8928 23288 8974
rect 23334 8928 23347 8974
rect 23275 8880 23347 8928
rect 23275 8834 23288 8880
rect 23334 8834 23347 8880
rect 26283 9444 26355 9492
rect 26283 9398 26296 9444
rect 26342 9398 26355 9444
rect 26283 9350 26355 9398
rect 26283 9304 26296 9350
rect 26342 9304 26355 9350
rect 26283 9256 26355 9304
rect 26283 9210 26296 9256
rect 26342 9210 26355 9256
rect 26283 9162 26355 9210
rect 26283 9116 26296 9162
rect 26342 9116 26355 9162
rect 26283 9068 26355 9116
rect 26283 9022 26296 9068
rect 26342 9022 26355 9068
rect 26283 8974 26355 9022
rect 26283 8928 26296 8974
rect 26342 8928 26355 8974
rect 26283 8880 26355 8928
rect 23275 8786 23347 8834
rect 23275 8740 23288 8786
rect 23334 8740 23347 8786
rect 23275 8692 23347 8740
rect 23275 8646 23288 8692
rect 23334 8646 23347 8692
rect 23275 8598 23347 8646
rect 26283 8834 26296 8880
rect 26342 8834 26355 8880
rect 26283 8786 26355 8834
rect 26283 8740 26296 8786
rect 26342 8740 26355 8786
rect 23275 8552 23288 8598
rect 23334 8552 23347 8598
rect 23275 8504 23347 8552
rect 26283 8692 26355 8740
rect 26283 8646 26296 8692
rect 26342 8646 26355 8692
rect 26283 8598 26355 8646
rect 26283 8552 26296 8598
rect 26342 8552 26355 8598
rect 23275 8458 23288 8504
rect 23334 8458 23347 8504
rect 23275 8410 23347 8458
rect 23275 8364 23288 8410
rect 23334 8364 23347 8410
rect 23275 8316 23347 8364
rect 23275 8270 23288 8316
rect 23334 8270 23347 8316
rect 23275 8222 23347 8270
rect 23275 8176 23288 8222
rect 23334 8176 23347 8222
rect 23275 8128 23347 8176
rect 23275 8082 23288 8128
rect 23334 8082 23347 8128
rect 23275 8034 23347 8082
rect 23275 7988 23288 8034
rect 23334 7988 23347 8034
rect 23275 7940 23347 7988
rect 23275 7894 23288 7940
rect 23334 7894 23347 7940
rect 26283 8504 26355 8552
rect 26283 8458 26296 8504
rect 26342 8458 26355 8504
rect 26283 8410 26355 8458
rect 26283 8364 26296 8410
rect 26342 8364 26355 8410
rect 26283 8316 26355 8364
rect 26283 8270 26296 8316
rect 26342 8270 26355 8316
rect 26283 8222 26355 8270
rect 26283 8176 26296 8222
rect 26342 8176 26355 8222
rect 26283 8128 26355 8176
rect 26283 8082 26296 8128
rect 26342 8082 26355 8128
rect 26283 8034 26355 8082
rect 26283 7988 26296 8034
rect 26342 7988 26355 8034
rect 26283 7940 26355 7988
rect 23275 7846 23347 7894
rect 23275 7800 23288 7846
rect 23334 7800 23347 7846
rect 26283 7894 26296 7940
rect 26342 7894 26355 7940
rect 23275 7752 23347 7800
rect 26283 7846 26355 7894
rect 26283 7800 26296 7846
rect 26342 7800 26355 7846
rect 23275 7706 23288 7752
rect 23334 7706 23347 7752
rect 23275 7658 23347 7706
rect 26283 7752 26355 7800
rect 26283 7706 26296 7752
rect 26342 7706 26355 7752
rect 23275 7612 23288 7658
rect 23334 7612 23347 7658
rect 23275 7564 23347 7612
rect 23275 7518 23288 7564
rect 23334 7518 23347 7564
rect 23275 7470 23347 7518
rect 23275 7424 23288 7470
rect 23334 7424 23347 7470
rect 23275 7389 23347 7424
rect 26283 7658 26355 7706
rect 26283 7612 26296 7658
rect 26342 7612 26355 7658
rect 26283 7564 26355 7612
rect 26283 7518 26296 7564
rect 26342 7518 26355 7564
rect 26283 7470 26355 7518
rect 26283 7424 26296 7470
rect 26342 7424 26355 7470
rect 26283 7389 26355 7424
rect 23275 7376 26355 7389
rect 23275 7330 23288 7376
rect 23334 7330 23382 7376
rect 23428 7330 23476 7376
rect 23522 7330 23570 7376
rect 23616 7330 23664 7376
rect 23710 7330 23758 7376
rect 23804 7330 23852 7376
rect 23898 7330 23946 7376
rect 23992 7330 24040 7376
rect 24086 7330 24134 7376
rect 24180 7330 24228 7376
rect 24274 7330 24322 7376
rect 24368 7330 24416 7376
rect 24462 7330 24510 7376
rect 24556 7330 24604 7376
rect 24650 7330 24698 7376
rect 24744 7330 24792 7376
rect 24838 7330 24886 7376
rect 24932 7330 24980 7376
rect 25026 7330 25074 7376
rect 25120 7330 25168 7376
rect 25214 7330 25262 7376
rect 25308 7330 25356 7376
rect 25402 7330 25450 7376
rect 25496 7330 25544 7376
rect 25590 7330 25638 7376
rect 25684 7330 25732 7376
rect 25778 7330 25826 7376
rect 25872 7330 25920 7376
rect 25966 7330 26014 7376
rect 26060 7330 26108 7376
rect 26154 7330 26202 7376
rect 26248 7330 26296 7376
rect 26342 7330 26355 7376
rect 23275 7317 26355 7330
rect 27244 13768 30324 13781
rect 27244 13722 27257 13768
rect 27303 13722 27351 13768
rect 27397 13722 27445 13768
rect 27491 13722 27539 13768
rect 27585 13722 27633 13768
rect 27679 13722 27727 13768
rect 27773 13722 27821 13768
rect 27867 13722 27915 13768
rect 27961 13722 28009 13768
rect 28055 13722 28103 13768
rect 28149 13722 28197 13768
rect 28243 13722 28291 13768
rect 28337 13722 28385 13768
rect 28431 13722 28479 13768
rect 28525 13722 28573 13768
rect 28619 13722 28667 13768
rect 28713 13722 28761 13768
rect 28807 13722 28855 13768
rect 28901 13722 28949 13768
rect 28995 13722 29043 13768
rect 29089 13722 29137 13768
rect 29183 13722 29231 13768
rect 29277 13722 29325 13768
rect 29371 13722 29419 13768
rect 29465 13722 29513 13768
rect 29559 13722 29607 13768
rect 29653 13722 29701 13768
rect 29747 13722 29795 13768
rect 29841 13722 29889 13768
rect 29935 13722 29983 13768
rect 30029 13722 30077 13768
rect 30123 13722 30171 13768
rect 30217 13722 30265 13768
rect 30311 13722 30324 13768
rect 27244 13709 30324 13722
rect 27244 13674 27316 13709
rect 27244 13628 27257 13674
rect 27303 13628 27316 13674
rect 27244 13580 27316 13628
rect 27244 13534 27257 13580
rect 27303 13534 27316 13580
rect 27244 13486 27316 13534
rect 27244 13440 27257 13486
rect 27303 13440 27316 13486
rect 27244 13392 27316 13440
rect 30252 13674 30324 13709
rect 30252 13628 30265 13674
rect 30311 13628 30324 13674
rect 30252 13580 30324 13628
rect 30252 13534 30265 13580
rect 30311 13534 30324 13580
rect 30252 13486 30324 13534
rect 30252 13440 30265 13486
rect 30311 13440 30324 13486
rect 27244 13346 27257 13392
rect 27303 13346 27316 13392
rect 27244 13298 27316 13346
rect 30252 13392 30324 13440
rect 30252 13346 30265 13392
rect 30311 13346 30324 13392
rect 27244 13252 27257 13298
rect 27303 13252 27316 13298
rect 27244 13204 27316 13252
rect 27244 13158 27257 13204
rect 27303 13158 27316 13204
rect 30252 13298 30324 13346
rect 30252 13252 30265 13298
rect 30311 13252 30324 13298
rect 30252 13204 30324 13252
rect 27244 13110 27316 13158
rect 27244 13064 27257 13110
rect 27303 13064 27316 13110
rect 27244 13016 27316 13064
rect 27244 12970 27257 13016
rect 27303 12970 27316 13016
rect 27244 12922 27316 12970
rect 27244 12876 27257 12922
rect 27303 12876 27316 12922
rect 27244 12828 27316 12876
rect 27244 12782 27257 12828
rect 27303 12782 27316 12828
rect 27244 12734 27316 12782
rect 27244 12688 27257 12734
rect 27303 12688 27316 12734
rect 27244 12640 27316 12688
rect 27244 12594 27257 12640
rect 27303 12594 27316 12640
rect 27244 12546 27316 12594
rect 30252 13158 30265 13204
rect 30311 13158 30324 13204
rect 30252 13110 30324 13158
rect 30252 13064 30265 13110
rect 30311 13064 30324 13110
rect 30252 13016 30324 13064
rect 30252 12970 30265 13016
rect 30311 12970 30324 13016
rect 30252 12922 30324 12970
rect 30252 12876 30265 12922
rect 30311 12876 30324 12922
rect 30252 12828 30324 12876
rect 30252 12782 30265 12828
rect 30311 12782 30324 12828
rect 30252 12734 30324 12782
rect 30252 12688 30265 12734
rect 30311 12688 30324 12734
rect 30252 12640 30324 12688
rect 30252 12594 30265 12640
rect 30311 12594 30324 12640
rect 27244 12500 27257 12546
rect 27303 12500 27316 12546
rect 27244 12452 27316 12500
rect 27244 12406 27257 12452
rect 27303 12406 27316 12452
rect 27244 12358 27316 12406
rect 30252 12546 30324 12594
rect 30252 12500 30265 12546
rect 30311 12500 30324 12546
rect 27244 12312 27257 12358
rect 27303 12312 27316 12358
rect 27244 12264 27316 12312
rect 27244 12218 27257 12264
rect 27303 12218 27316 12264
rect 30252 12452 30324 12500
rect 30252 12406 30265 12452
rect 30311 12406 30324 12452
rect 30252 12358 30324 12406
rect 30252 12312 30265 12358
rect 30311 12312 30324 12358
rect 30252 12264 30324 12312
rect 27244 12170 27316 12218
rect 27244 12124 27257 12170
rect 27303 12124 27316 12170
rect 27244 12076 27316 12124
rect 27244 12030 27257 12076
rect 27303 12030 27316 12076
rect 27244 11982 27316 12030
rect 27244 11936 27257 11982
rect 27303 11936 27316 11982
rect 27244 11888 27316 11936
rect 27244 11842 27257 11888
rect 27303 11842 27316 11888
rect 27244 11794 27316 11842
rect 27244 11748 27257 11794
rect 27303 11748 27316 11794
rect 27244 11700 27316 11748
rect 27244 11654 27257 11700
rect 27303 11654 27316 11700
rect 27244 11606 27316 11654
rect 30252 12218 30265 12264
rect 30311 12218 30324 12264
rect 30252 12170 30324 12218
rect 30252 12124 30265 12170
rect 30311 12124 30324 12170
rect 30252 12076 30324 12124
rect 30252 12030 30265 12076
rect 30311 12030 30324 12076
rect 30252 11982 30324 12030
rect 30252 11936 30265 11982
rect 30311 11936 30324 11982
rect 30252 11888 30324 11936
rect 30252 11842 30265 11888
rect 30311 11842 30324 11888
rect 30252 11794 30324 11842
rect 30252 11748 30265 11794
rect 30311 11748 30324 11794
rect 30252 11700 30324 11748
rect 30252 11654 30265 11700
rect 30311 11654 30324 11700
rect 27244 11560 27257 11606
rect 27303 11560 27316 11606
rect 27244 11512 27316 11560
rect 27244 11466 27257 11512
rect 27303 11466 27316 11512
rect 27244 11418 27316 11466
rect 27244 11372 27257 11418
rect 27303 11372 27316 11418
rect 27244 11324 27316 11372
rect 27244 11278 27257 11324
rect 27303 11278 27316 11324
rect 30252 11606 30324 11654
rect 30252 11560 30265 11606
rect 30311 11560 30324 11606
rect 30252 11512 30324 11560
rect 30252 11466 30265 11512
rect 30311 11466 30324 11512
rect 30252 11418 30324 11466
rect 30252 11372 30265 11418
rect 30311 11372 30324 11418
rect 30252 11324 30324 11372
rect 27244 11230 27316 11278
rect 27244 11184 27257 11230
rect 27303 11184 27316 11230
rect 27244 11136 27316 11184
rect 27244 11090 27257 11136
rect 27303 11090 27316 11136
rect 27244 11042 27316 11090
rect 27244 10996 27257 11042
rect 27303 10996 27316 11042
rect 27244 10948 27316 10996
rect 27244 10902 27257 10948
rect 27303 10902 27316 10948
rect 27244 10854 27316 10902
rect 27244 10808 27257 10854
rect 27303 10808 27316 10854
rect 27244 10760 27316 10808
rect 27244 10714 27257 10760
rect 27303 10714 27316 10760
rect 30252 11278 30265 11324
rect 30311 11278 30324 11324
rect 30252 11230 30324 11278
rect 30252 11184 30265 11230
rect 30311 11184 30324 11230
rect 30252 11136 30324 11184
rect 30252 11090 30265 11136
rect 30311 11090 30324 11136
rect 30252 11042 30324 11090
rect 30252 10996 30265 11042
rect 30311 10996 30324 11042
rect 30252 10948 30324 10996
rect 30252 10902 30265 10948
rect 30311 10902 30324 10948
rect 30252 10854 30324 10902
rect 30252 10808 30265 10854
rect 30311 10808 30324 10854
rect 30252 10760 30324 10808
rect 27244 10666 27316 10714
rect 27244 10620 27257 10666
rect 27303 10620 27316 10666
rect 27244 10572 27316 10620
rect 27244 10526 27257 10572
rect 27303 10526 27316 10572
rect 27244 10478 27316 10526
rect 27244 10432 27257 10478
rect 27303 10432 27316 10478
rect 27244 10384 27316 10432
rect 27244 10338 27257 10384
rect 27303 10338 27316 10384
rect 30252 10714 30265 10760
rect 30311 10714 30324 10760
rect 30252 10666 30324 10714
rect 30252 10620 30265 10666
rect 30311 10620 30324 10666
rect 30252 10572 30324 10620
rect 30252 10526 30265 10572
rect 30311 10526 30324 10572
rect 30252 10478 30324 10526
rect 30252 10432 30265 10478
rect 30311 10432 30324 10478
rect 30252 10384 30324 10432
rect 27244 10290 27316 10338
rect 27244 10244 27257 10290
rect 27303 10244 27316 10290
rect 27244 10196 27316 10244
rect 27244 10150 27257 10196
rect 27303 10150 27316 10196
rect 27244 10102 27316 10150
rect 27244 10056 27257 10102
rect 27303 10056 27316 10102
rect 27244 10008 27316 10056
rect 27244 9962 27257 10008
rect 27303 9962 27316 10008
rect 27244 9914 27316 9962
rect 27244 9868 27257 9914
rect 27303 9868 27316 9914
rect 27244 9820 27316 9868
rect 27244 9774 27257 9820
rect 27303 9774 27316 9820
rect 30252 10338 30265 10384
rect 30311 10338 30324 10384
rect 30252 10290 30324 10338
rect 30252 10244 30265 10290
rect 30311 10244 30324 10290
rect 30252 10196 30324 10244
rect 30252 10150 30265 10196
rect 30311 10150 30324 10196
rect 30252 10102 30324 10150
rect 30252 10056 30265 10102
rect 30311 10056 30324 10102
rect 30252 10008 30324 10056
rect 30252 9962 30265 10008
rect 30311 9962 30324 10008
rect 30252 9914 30324 9962
rect 30252 9868 30265 9914
rect 30311 9868 30324 9914
rect 30252 9820 30324 9868
rect 27244 9726 27316 9774
rect 27244 9680 27257 9726
rect 27303 9680 27316 9726
rect 27244 9632 27316 9680
rect 27244 9586 27257 9632
rect 27303 9586 27316 9632
rect 27244 9538 27316 9586
rect 27244 9492 27257 9538
rect 27303 9492 27316 9538
rect 27244 9444 27316 9492
rect 30252 9774 30265 9820
rect 30311 9774 30324 9820
rect 30252 9726 30324 9774
rect 30252 9680 30265 9726
rect 30311 9680 30324 9726
rect 30252 9632 30324 9680
rect 30252 9586 30265 9632
rect 30311 9586 30324 9632
rect 30252 9538 30324 9586
rect 30252 9492 30265 9538
rect 30311 9492 30324 9538
rect 27244 9398 27257 9444
rect 27303 9398 27316 9444
rect 27244 9350 27316 9398
rect 27244 9304 27257 9350
rect 27303 9304 27316 9350
rect 27244 9256 27316 9304
rect 27244 9210 27257 9256
rect 27303 9210 27316 9256
rect 27244 9162 27316 9210
rect 27244 9116 27257 9162
rect 27303 9116 27316 9162
rect 27244 9068 27316 9116
rect 27244 9022 27257 9068
rect 27303 9022 27316 9068
rect 27244 8974 27316 9022
rect 27244 8928 27257 8974
rect 27303 8928 27316 8974
rect 27244 8880 27316 8928
rect 27244 8834 27257 8880
rect 27303 8834 27316 8880
rect 30252 9444 30324 9492
rect 30252 9398 30265 9444
rect 30311 9398 30324 9444
rect 30252 9350 30324 9398
rect 30252 9304 30265 9350
rect 30311 9304 30324 9350
rect 30252 9256 30324 9304
rect 30252 9210 30265 9256
rect 30311 9210 30324 9256
rect 30252 9162 30324 9210
rect 30252 9116 30265 9162
rect 30311 9116 30324 9162
rect 30252 9068 30324 9116
rect 30252 9022 30265 9068
rect 30311 9022 30324 9068
rect 30252 8974 30324 9022
rect 30252 8928 30265 8974
rect 30311 8928 30324 8974
rect 30252 8880 30324 8928
rect 27244 8786 27316 8834
rect 27244 8740 27257 8786
rect 27303 8740 27316 8786
rect 27244 8692 27316 8740
rect 27244 8646 27257 8692
rect 27303 8646 27316 8692
rect 27244 8598 27316 8646
rect 30252 8834 30265 8880
rect 30311 8834 30324 8880
rect 30252 8786 30324 8834
rect 30252 8740 30265 8786
rect 30311 8740 30324 8786
rect 27244 8552 27257 8598
rect 27303 8552 27316 8598
rect 27244 8504 27316 8552
rect 30252 8692 30324 8740
rect 30252 8646 30265 8692
rect 30311 8646 30324 8692
rect 30252 8598 30324 8646
rect 30252 8552 30265 8598
rect 30311 8552 30324 8598
rect 27244 8458 27257 8504
rect 27303 8458 27316 8504
rect 27244 8410 27316 8458
rect 27244 8364 27257 8410
rect 27303 8364 27316 8410
rect 27244 8316 27316 8364
rect 27244 8270 27257 8316
rect 27303 8270 27316 8316
rect 27244 8222 27316 8270
rect 27244 8176 27257 8222
rect 27303 8176 27316 8222
rect 27244 8128 27316 8176
rect 27244 8082 27257 8128
rect 27303 8082 27316 8128
rect 27244 8034 27316 8082
rect 27244 7988 27257 8034
rect 27303 7988 27316 8034
rect 27244 7940 27316 7988
rect 27244 7894 27257 7940
rect 27303 7894 27316 7940
rect 30252 8504 30324 8552
rect 30252 8458 30265 8504
rect 30311 8458 30324 8504
rect 30252 8410 30324 8458
rect 30252 8364 30265 8410
rect 30311 8364 30324 8410
rect 30252 8316 30324 8364
rect 30252 8270 30265 8316
rect 30311 8270 30324 8316
rect 30252 8222 30324 8270
rect 30252 8176 30265 8222
rect 30311 8176 30324 8222
rect 30252 8128 30324 8176
rect 30252 8082 30265 8128
rect 30311 8082 30324 8128
rect 30252 8034 30324 8082
rect 30252 7988 30265 8034
rect 30311 7988 30324 8034
rect 30252 7940 30324 7988
rect 27244 7846 27316 7894
rect 27244 7800 27257 7846
rect 27303 7800 27316 7846
rect 27244 7752 27316 7800
rect 30252 7894 30265 7940
rect 30311 7894 30324 7940
rect 30252 7846 30324 7894
rect 30252 7800 30265 7846
rect 30311 7800 30324 7846
rect 27244 7706 27257 7752
rect 27303 7706 27316 7752
rect 27244 7658 27316 7706
rect 30252 7752 30324 7800
rect 30252 7706 30265 7752
rect 30311 7706 30324 7752
rect 27244 7612 27257 7658
rect 27303 7612 27316 7658
rect 27244 7564 27316 7612
rect 27244 7518 27257 7564
rect 27303 7518 27316 7564
rect 27244 7470 27316 7518
rect 27244 7424 27257 7470
rect 27303 7424 27316 7470
rect 27244 7389 27316 7424
rect 30252 7658 30324 7706
rect 30252 7612 30265 7658
rect 30311 7612 30324 7658
rect 30252 7564 30324 7612
rect 30252 7518 30265 7564
rect 30311 7518 30324 7564
rect 30252 7470 30324 7518
rect 30252 7424 30265 7470
rect 30311 7424 30324 7470
rect 30252 7389 30324 7424
rect 27244 7376 30324 7389
rect 27244 7330 27257 7376
rect 27303 7330 27351 7376
rect 27397 7330 27445 7376
rect 27491 7330 27539 7376
rect 27585 7330 27633 7376
rect 27679 7330 27727 7376
rect 27773 7330 27821 7376
rect 27867 7330 27915 7376
rect 27961 7330 28009 7376
rect 28055 7330 28103 7376
rect 28149 7330 28197 7376
rect 28243 7330 28291 7376
rect 28337 7330 28385 7376
rect 28431 7330 28479 7376
rect 28525 7330 28573 7376
rect 28619 7330 28667 7376
rect 28713 7330 28761 7376
rect 28807 7330 28855 7376
rect 28901 7330 28949 7376
rect 28995 7330 29043 7376
rect 29089 7330 29137 7376
rect 29183 7330 29231 7376
rect 29277 7330 29325 7376
rect 29371 7330 29419 7376
rect 29465 7330 29513 7376
rect 29559 7330 29607 7376
rect 29653 7330 29701 7376
rect 29747 7330 29795 7376
rect 29841 7330 29889 7376
rect 29935 7330 29983 7376
rect 30029 7330 30077 7376
rect 30123 7330 30171 7376
rect 30217 7330 30265 7376
rect 30311 7330 30324 7376
rect 27244 7317 30324 7330
rect 6921 6118 10095 6131
rect 6921 6072 6934 6118
rect 6980 6072 7028 6118
rect 7074 6072 7122 6118
rect 7168 6072 7216 6118
rect 7262 6072 7310 6118
rect 7356 6072 7404 6118
rect 7450 6072 7498 6118
rect 7544 6072 7592 6118
rect 7638 6072 7686 6118
rect 7732 6072 7780 6118
rect 7826 6072 7874 6118
rect 7920 6072 7968 6118
rect 8014 6072 8062 6118
rect 8108 6072 8156 6118
rect 8202 6072 8250 6118
rect 8296 6072 8344 6118
rect 8390 6072 8438 6118
rect 8484 6072 8532 6118
rect 8578 6072 8626 6118
rect 8672 6072 8720 6118
rect 8766 6072 8814 6118
rect 8860 6072 8908 6118
rect 8954 6072 9002 6118
rect 9048 6072 9096 6118
rect 9142 6072 9190 6118
rect 9236 6072 9284 6118
rect 9330 6072 9378 6118
rect 9424 6072 9472 6118
rect 9518 6072 9566 6118
rect 9612 6072 9660 6118
rect 9706 6072 9754 6118
rect 9800 6072 9848 6118
rect 9894 6072 9942 6118
rect 9988 6072 10036 6118
rect 10082 6072 10095 6118
rect 6921 6059 10095 6072
rect 6921 6024 6993 6059
rect 6921 5978 6934 6024
rect 6980 5978 6993 6024
rect 6921 5930 6993 5978
rect 10023 6024 10095 6059
rect 10023 5978 10036 6024
rect 10082 5978 10095 6024
rect 6921 5884 6934 5930
rect 6980 5884 6993 5930
rect 6921 5836 6993 5884
rect 6921 5790 6934 5836
rect 6980 5790 6993 5836
rect 6921 5742 6993 5790
rect 6921 5696 6934 5742
rect 6980 5696 6993 5742
rect 10023 5930 10095 5978
rect 10023 5884 10036 5930
rect 10082 5884 10095 5930
rect 10023 5836 10095 5884
rect 10023 5790 10036 5836
rect 10082 5790 10095 5836
rect 10023 5742 10095 5790
rect 6921 5648 6993 5696
rect 6921 5602 6934 5648
rect 6980 5602 6993 5648
rect 6921 5554 6993 5602
rect 6921 5508 6934 5554
rect 6980 5508 6993 5554
rect 10023 5696 10036 5742
rect 10082 5696 10095 5742
rect 10023 5648 10095 5696
rect 10023 5602 10036 5648
rect 10082 5602 10095 5648
rect 10023 5554 10095 5602
rect 6921 5460 6993 5508
rect 6921 5414 6934 5460
rect 6980 5414 6993 5460
rect 6921 5366 6993 5414
rect 6921 5320 6934 5366
rect 6980 5320 6993 5366
rect 6921 5272 6993 5320
rect 6921 5226 6934 5272
rect 6980 5226 6993 5272
rect 6921 5178 6993 5226
rect 10023 5508 10036 5554
rect 10082 5508 10095 5554
rect 10023 5460 10095 5508
rect 10023 5414 10036 5460
rect 10082 5414 10095 5460
rect 10023 5366 10095 5414
rect 10023 5320 10036 5366
rect 10082 5320 10095 5366
rect 10023 5272 10095 5320
rect 10023 5226 10036 5272
rect 10082 5226 10095 5272
rect 6921 5132 6934 5178
rect 6980 5132 6993 5178
rect 6921 5084 6993 5132
rect 6921 5038 6934 5084
rect 6980 5038 6993 5084
rect 6921 4990 6993 5038
rect 10023 5178 10095 5226
rect 10023 5132 10036 5178
rect 10082 5132 10095 5178
rect 10023 5084 10095 5132
rect 10023 5038 10036 5084
rect 10082 5038 10095 5084
rect 6921 4944 6934 4990
rect 6980 4944 6993 4990
rect 6921 4896 6993 4944
rect 6921 4850 6934 4896
rect 6980 4850 6993 4896
rect 6921 4802 6993 4850
rect 6921 4756 6934 4802
rect 6980 4756 6993 4802
rect 6921 4708 6993 4756
rect 6921 4662 6934 4708
rect 6980 4662 6993 4708
rect 10023 4990 10095 5038
rect 10023 4944 10036 4990
rect 10082 4944 10095 4990
rect 10023 4896 10095 4944
rect 10023 4850 10036 4896
rect 10082 4850 10095 4896
rect 10023 4802 10095 4850
rect 10023 4756 10036 4802
rect 10082 4756 10095 4802
rect 10023 4708 10095 4756
rect 6921 4614 6993 4662
rect 6921 4568 6934 4614
rect 6980 4568 6993 4614
rect 6921 4520 6993 4568
rect 6921 4474 6934 4520
rect 6980 4474 6993 4520
rect 6921 4426 6993 4474
rect 10023 4662 10036 4708
rect 10082 4662 10095 4708
rect 10023 4614 10095 4662
rect 10023 4568 10036 4614
rect 10082 4568 10095 4614
rect 10023 4520 10095 4568
rect 10023 4474 10036 4520
rect 10082 4474 10095 4520
rect 6921 4380 6934 4426
rect 6980 4380 6993 4426
rect 6921 4332 6993 4380
rect 6921 4286 6934 4332
rect 6980 4286 6993 4332
rect 6921 4238 6993 4286
rect 6921 4192 6934 4238
rect 6980 4192 6993 4238
rect 6921 4144 6993 4192
rect 6921 4098 6934 4144
rect 6980 4098 6993 4144
rect 10023 4426 10095 4474
rect 10023 4380 10036 4426
rect 10082 4380 10095 4426
rect 10023 4332 10095 4380
rect 10023 4286 10036 4332
rect 10082 4286 10095 4332
rect 10023 4238 10095 4286
rect 10023 4192 10036 4238
rect 10082 4192 10095 4238
rect 10023 4144 10095 4192
rect 6921 4050 6993 4098
rect 6921 4004 6934 4050
rect 6980 4004 6993 4050
rect 6921 3956 6993 4004
rect 6921 3910 6934 3956
rect 6980 3910 6993 3956
rect 10023 4098 10036 4144
rect 10082 4098 10095 4144
rect 10023 4050 10095 4098
rect 10023 4004 10036 4050
rect 10082 4004 10095 4050
rect 10023 3956 10095 4004
rect 6921 3862 6993 3910
rect 6921 3816 6934 3862
rect 6980 3816 6993 3862
rect 6921 3768 6993 3816
rect 6921 3722 6934 3768
rect 6980 3722 6993 3768
rect 6921 3674 6993 3722
rect 6921 3628 6934 3674
rect 6980 3628 6993 3674
rect 6921 3580 6993 3628
rect 10023 3910 10036 3956
rect 10082 3910 10095 3956
rect 10023 3862 10095 3910
rect 10023 3816 10036 3862
rect 10082 3816 10095 3862
rect 10023 3768 10095 3816
rect 10023 3722 10036 3768
rect 10082 3722 10095 3768
rect 10023 3674 10095 3722
rect 10023 3628 10036 3674
rect 10082 3628 10095 3674
rect 6921 3534 6934 3580
rect 6980 3534 6993 3580
rect 6921 3486 6993 3534
rect 6921 3440 6934 3486
rect 6980 3440 6993 3486
rect 6921 3392 6993 3440
rect 10023 3580 10095 3628
rect 10023 3534 10036 3580
rect 10082 3534 10095 3580
rect 10023 3486 10095 3534
rect 10023 3440 10036 3486
rect 10082 3440 10095 3486
rect 6921 3346 6934 3392
rect 6980 3346 6993 3392
rect 6921 3298 6993 3346
rect 6921 3252 6934 3298
rect 6980 3252 6993 3298
rect 6921 3204 6993 3252
rect 6921 3158 6934 3204
rect 6980 3158 6993 3204
rect 6921 3110 6993 3158
rect 6921 3064 6934 3110
rect 6980 3064 6993 3110
rect 6921 3016 6993 3064
rect 10023 3392 10095 3440
rect 10023 3346 10036 3392
rect 10082 3346 10095 3392
rect 10023 3298 10095 3346
rect 10023 3252 10036 3298
rect 10082 3252 10095 3298
rect 10023 3204 10095 3252
rect 10023 3158 10036 3204
rect 10082 3158 10095 3204
rect 10023 3110 10095 3158
rect 10023 3064 10036 3110
rect 10082 3064 10095 3110
rect 6921 2970 6934 3016
rect 6980 2970 6993 3016
rect 6921 2922 6993 2970
rect 6921 2876 6934 2922
rect 6980 2876 6993 2922
rect 6921 2841 6993 2876
rect 10023 3016 10095 3064
rect 10023 2970 10036 3016
rect 10082 2970 10095 3016
rect 10023 2922 10095 2970
rect 10023 2876 10036 2922
rect 10082 2876 10095 2922
rect 5887 2828 6993 2841
rect 5887 2782 5900 2828
rect 5946 2782 5994 2828
rect 6040 2782 6088 2828
rect 6134 2782 6182 2828
rect 6228 2782 6276 2828
rect 6322 2782 6370 2828
rect 6416 2782 6464 2828
rect 6510 2782 6558 2828
rect 6604 2782 6652 2828
rect 6698 2782 6746 2828
rect 6792 2782 6840 2828
rect 6886 2782 6934 2828
rect 6980 2782 6993 2828
rect 5887 2769 6993 2782
rect 10023 2841 10095 2876
rect 12001 4469 17619 4482
rect 12001 4423 12014 4469
rect 12060 4423 12108 4469
rect 12154 4423 12202 4469
rect 12248 4423 12296 4469
rect 12342 4423 12390 4469
rect 12436 4423 12484 4469
rect 12530 4423 12578 4469
rect 12624 4423 12672 4469
rect 12718 4423 12766 4469
rect 12812 4423 12860 4469
rect 12906 4423 12954 4469
rect 13000 4423 13048 4469
rect 13094 4423 13142 4469
rect 13188 4423 13236 4469
rect 13282 4423 13330 4469
rect 13376 4423 13424 4469
rect 13470 4423 13518 4469
rect 13564 4423 13612 4469
rect 13658 4423 13706 4469
rect 13752 4423 13800 4469
rect 13846 4423 13894 4469
rect 13940 4423 13988 4469
rect 14034 4423 14082 4469
rect 14128 4423 14176 4469
rect 14222 4423 14270 4469
rect 14316 4423 14364 4469
rect 14410 4423 14458 4469
rect 14504 4423 14552 4469
rect 14598 4423 14646 4469
rect 14692 4423 14740 4469
rect 14786 4423 14834 4469
rect 14880 4423 14928 4469
rect 14974 4423 15022 4469
rect 15068 4423 15116 4469
rect 15162 4423 15210 4469
rect 15256 4423 15304 4469
rect 15350 4423 15398 4469
rect 15444 4423 15492 4469
rect 15538 4423 15586 4469
rect 15632 4423 15680 4469
rect 15726 4423 15774 4469
rect 15820 4423 15868 4469
rect 15914 4423 15962 4469
rect 16008 4423 16056 4469
rect 16102 4423 16150 4469
rect 16196 4423 16244 4469
rect 16290 4423 16338 4469
rect 16384 4423 16432 4469
rect 16478 4423 16526 4469
rect 16572 4423 16620 4469
rect 16666 4423 16714 4469
rect 16760 4423 16808 4469
rect 16854 4423 16902 4469
rect 16948 4423 16996 4469
rect 17042 4423 17090 4469
rect 17136 4423 17184 4469
rect 17230 4423 17278 4469
rect 17324 4423 17372 4469
rect 17418 4423 17466 4469
rect 17512 4423 17560 4469
rect 17606 4423 17619 4469
rect 12001 4410 17619 4423
rect 12001 4375 12073 4410
rect 12001 4329 12014 4375
rect 12060 4329 12073 4375
rect 12001 4281 12073 4329
rect 12001 4235 12014 4281
rect 12060 4235 12073 4281
rect 12001 4187 12073 4235
rect 12001 4141 12014 4187
rect 12060 4141 12073 4187
rect 12001 4093 12073 4141
rect 12001 4047 12014 4093
rect 12060 4047 12073 4093
rect 17547 4375 17619 4410
rect 17547 4329 17560 4375
rect 17606 4329 17619 4375
rect 17547 4281 17619 4329
rect 17547 4235 17560 4281
rect 17606 4235 17619 4281
rect 17547 4187 17619 4235
rect 17547 4141 17560 4187
rect 17606 4141 17619 4187
rect 17547 4093 17619 4141
rect 12001 3999 12073 4047
rect 12001 3953 12014 3999
rect 12060 3953 12073 3999
rect 12001 3905 12073 3953
rect 12001 3859 12014 3905
rect 12060 3859 12073 3905
rect 12001 3811 12073 3859
rect 12001 3765 12014 3811
rect 12060 3765 12073 3811
rect 17547 4047 17560 4093
rect 17606 4047 17619 4093
rect 17547 3999 17619 4047
rect 17547 3953 17560 3999
rect 17606 3953 17619 3999
rect 17547 3905 17619 3953
rect 17547 3859 17560 3905
rect 17606 3859 17619 3905
rect 17547 3811 17619 3859
rect 12001 3717 12073 3765
rect 12001 3671 12014 3717
rect 12060 3671 12073 3717
rect 12001 3623 12073 3671
rect 12001 3577 12014 3623
rect 12060 3577 12073 3623
rect 12001 3529 12073 3577
rect 12001 3483 12014 3529
rect 12060 3483 12073 3529
rect 12001 3435 12073 3483
rect 12001 3389 12014 3435
rect 12060 3389 12073 3435
rect 12001 3341 12073 3389
rect 17547 3765 17560 3811
rect 17606 3765 17619 3811
rect 17547 3717 17619 3765
rect 17547 3671 17560 3717
rect 17606 3671 17619 3717
rect 17547 3623 17619 3671
rect 17547 3577 17560 3623
rect 17606 3577 17619 3623
rect 17547 3529 17619 3577
rect 17547 3483 17560 3529
rect 17606 3483 17619 3529
rect 17547 3435 17619 3483
rect 17547 3389 17560 3435
rect 17606 3389 17619 3435
rect 12001 3295 12014 3341
rect 12060 3295 12073 3341
rect 12001 3247 12073 3295
rect 12001 3201 12014 3247
rect 12060 3201 12073 3247
rect 17547 3341 17619 3389
rect 17547 3295 17560 3341
rect 17606 3295 17619 3341
rect 17547 3247 17619 3295
rect 12001 3153 12073 3201
rect 12001 3107 12014 3153
rect 12060 3107 12073 3153
rect 12001 3059 12073 3107
rect 12001 3013 12014 3059
rect 12060 3013 12073 3059
rect 12001 2965 12073 3013
rect 12001 2919 12014 2965
rect 12060 2919 12073 2965
rect 12001 2871 12073 2919
rect 10023 2828 11129 2841
rect 10023 2782 10036 2828
rect 10082 2782 10130 2828
rect 10176 2782 10224 2828
rect 10270 2782 10318 2828
rect 10364 2782 10412 2828
rect 10458 2782 10506 2828
rect 10552 2782 10600 2828
rect 10646 2782 10694 2828
rect 10740 2782 10788 2828
rect 10834 2782 10882 2828
rect 10928 2782 10976 2828
rect 11022 2782 11070 2828
rect 11116 2782 11129 2828
rect 5887 2734 5959 2769
rect 10023 2769 11129 2782
rect 11057 2734 11129 2769
rect 5887 2688 5900 2734
rect 5946 2688 5959 2734
rect 5887 2640 5959 2688
rect 11057 2688 11070 2734
rect 11116 2688 11129 2734
rect 5887 2594 5900 2640
rect 5946 2594 5959 2640
rect 5887 2546 5959 2594
rect 5887 2500 5900 2546
rect 5946 2500 5959 2546
rect 5887 2452 5959 2500
rect 5887 2406 5900 2452
rect 5946 2406 5959 2452
rect 11057 2640 11129 2688
rect 11057 2594 11070 2640
rect 11116 2594 11129 2640
rect 11057 2546 11129 2594
rect 11057 2500 11070 2546
rect 11116 2500 11129 2546
rect 11057 2452 11129 2500
rect 5887 2358 5959 2406
rect 5887 2312 5900 2358
rect 5946 2312 5959 2358
rect 5887 2264 5959 2312
rect 5887 2218 5900 2264
rect 5946 2218 5959 2264
rect 11057 2406 11070 2452
rect 11116 2406 11129 2452
rect 11057 2358 11129 2406
rect 11057 2312 11070 2358
rect 11116 2312 11129 2358
rect 11057 2264 11129 2312
rect 5887 2170 5959 2218
rect 5887 2124 5900 2170
rect 5946 2124 5959 2170
rect 5887 2076 5959 2124
rect 5887 2030 5900 2076
rect 5946 2030 5959 2076
rect 11057 2218 11070 2264
rect 11116 2218 11129 2264
rect 11057 2170 11129 2218
rect 11057 2124 11070 2170
rect 11116 2124 11129 2170
rect 11057 2076 11129 2124
rect 5887 1982 5959 2030
rect 5887 1936 5900 1982
rect 5946 1936 5959 1982
rect 11057 2030 11070 2076
rect 11116 2030 11129 2076
rect 11057 1982 11129 2030
rect 5887 1888 5959 1936
rect 5887 1842 5900 1888
rect 5946 1842 5959 1888
rect 5887 1794 5959 1842
rect 5887 1748 5900 1794
rect 5946 1748 5959 1794
rect 11057 1936 11070 1982
rect 11116 1936 11129 1982
rect 11057 1888 11129 1936
rect 11057 1842 11070 1888
rect 11116 1842 11129 1888
rect 11057 1794 11129 1842
rect 5887 1700 5959 1748
rect 5887 1654 5900 1700
rect 5946 1654 5959 1700
rect 5887 1606 5959 1654
rect 5887 1560 5900 1606
rect 5946 1560 5959 1606
rect 11057 1748 11070 1794
rect 11116 1748 11129 1794
rect 11057 1700 11129 1748
rect 11057 1654 11070 1700
rect 11116 1654 11129 1700
rect 11057 1606 11129 1654
rect 5887 1512 5959 1560
rect 11057 1560 11070 1606
rect 11116 1560 11129 1606
rect 5887 1466 5900 1512
rect 5946 1466 5959 1512
rect 5887 1418 5959 1466
rect 5887 1372 5900 1418
rect 5946 1372 5959 1418
rect 5887 1337 5959 1372
rect 11057 1512 11129 1560
rect 11057 1466 11070 1512
rect 11116 1466 11129 1512
rect 11057 1418 11129 1466
rect 11057 1372 11070 1418
rect 11116 1372 11129 1418
rect 11057 1337 11129 1372
rect 5887 1324 11129 1337
rect 5887 1278 5900 1324
rect 5946 1278 5994 1324
rect 6040 1278 6088 1324
rect 6134 1278 6182 1324
rect 6228 1278 6276 1324
rect 6322 1278 6370 1324
rect 6416 1278 6464 1324
rect 6510 1278 6558 1324
rect 6604 1278 6652 1324
rect 6698 1278 6746 1324
rect 6792 1278 6840 1324
rect 6886 1278 6934 1324
rect 6980 1278 7028 1324
rect 7074 1278 7122 1324
rect 7168 1278 7216 1324
rect 7262 1278 7310 1324
rect 7356 1278 7404 1324
rect 7450 1278 7498 1324
rect 7544 1278 7592 1324
rect 7638 1278 7686 1324
rect 7732 1278 7780 1324
rect 7826 1278 7874 1324
rect 7920 1278 7968 1324
rect 8014 1278 8062 1324
rect 8108 1278 8156 1324
rect 8202 1278 8250 1324
rect 8296 1278 8344 1324
rect 8390 1278 8438 1324
rect 8484 1278 8532 1324
rect 8578 1278 8626 1324
rect 8672 1278 8720 1324
rect 8766 1278 8814 1324
rect 8860 1278 8908 1324
rect 8954 1278 9002 1324
rect 9048 1278 9096 1324
rect 9142 1278 9190 1324
rect 9236 1278 9284 1324
rect 9330 1278 9378 1324
rect 9424 1278 9472 1324
rect 9518 1278 9566 1324
rect 9612 1278 9660 1324
rect 9706 1278 9754 1324
rect 9800 1278 9848 1324
rect 9894 1278 9942 1324
rect 9988 1278 10036 1324
rect 10082 1278 10130 1324
rect 10176 1278 10224 1324
rect 10270 1278 10318 1324
rect 10364 1278 10412 1324
rect 10458 1278 10506 1324
rect 10552 1278 10600 1324
rect 10646 1278 10694 1324
rect 10740 1278 10788 1324
rect 10834 1278 10882 1324
rect 10928 1278 10976 1324
rect 11022 1278 11070 1324
rect 11116 1278 11129 1324
rect 12001 2825 12014 2871
rect 12060 2825 12073 2871
rect 17547 3201 17560 3247
rect 17606 3201 17619 3247
rect 17547 3153 17619 3201
rect 17547 3107 17560 3153
rect 17606 3107 17619 3153
rect 17547 3059 17619 3107
rect 17547 3013 17560 3059
rect 17606 3013 17619 3059
rect 17547 2965 17619 3013
rect 17547 2919 17560 2965
rect 17606 2919 17619 2965
rect 17547 2871 17619 2919
rect 12001 2777 12073 2825
rect 12001 2731 12014 2777
rect 12060 2731 12073 2777
rect 12001 2683 12073 2731
rect 12001 2637 12014 2683
rect 12060 2637 12073 2683
rect 12001 2589 12073 2637
rect 12001 2543 12014 2589
rect 12060 2543 12073 2589
rect 12001 2495 12073 2543
rect 12001 2449 12014 2495
rect 12060 2449 12073 2495
rect 12001 2401 12073 2449
rect 17547 2825 17560 2871
rect 17606 2825 17619 2871
rect 17547 2777 17619 2825
rect 17547 2731 17560 2777
rect 17606 2731 17619 2777
rect 17547 2683 17619 2731
rect 17547 2637 17560 2683
rect 17606 2637 17619 2683
rect 17547 2589 17619 2637
rect 17547 2543 17560 2589
rect 17606 2543 17619 2589
rect 17547 2495 17619 2543
rect 17547 2449 17560 2495
rect 17606 2449 17619 2495
rect 12001 2355 12014 2401
rect 12060 2355 12073 2401
rect 12001 2307 12073 2355
rect 12001 2261 12014 2307
rect 12060 2261 12073 2307
rect 12001 2213 12073 2261
rect 12001 2167 12014 2213
rect 12060 2167 12073 2213
rect 12001 2119 12073 2167
rect 12001 2073 12014 2119
rect 12060 2073 12073 2119
rect 12001 2025 12073 2073
rect 12001 1979 12014 2025
rect 12060 1979 12073 2025
rect 17547 2401 17619 2449
rect 17547 2355 17560 2401
rect 17606 2355 17619 2401
rect 17547 2307 17619 2355
rect 17547 2261 17560 2307
rect 17606 2261 17619 2307
rect 17547 2213 17619 2261
rect 17547 2167 17560 2213
rect 17606 2167 17619 2213
rect 17547 2119 17619 2167
rect 17547 2073 17560 2119
rect 17606 2073 17619 2119
rect 17547 2025 17619 2073
rect 12001 1931 12073 1979
rect 12001 1885 12014 1931
rect 12060 1885 12073 1931
rect 12001 1837 12073 1885
rect 12001 1791 12014 1837
rect 12060 1791 12073 1837
rect 12001 1743 12073 1791
rect 12001 1697 12014 1743
rect 12060 1697 12073 1743
rect 12001 1649 12073 1697
rect 12001 1603 12014 1649
rect 12060 1603 12073 1649
rect 17547 1979 17560 2025
rect 17606 1979 17619 2025
rect 17547 1931 17619 1979
rect 17547 1885 17560 1931
rect 17606 1885 17619 1931
rect 17547 1837 17619 1885
rect 17547 1791 17560 1837
rect 17606 1791 17619 1837
rect 17547 1743 17619 1791
rect 17547 1697 17560 1743
rect 17606 1697 17619 1743
rect 17547 1649 17619 1697
rect 12001 1555 12073 1603
rect 12001 1509 12014 1555
rect 12060 1509 12073 1555
rect 12001 1461 12073 1509
rect 12001 1415 12014 1461
rect 12060 1415 12073 1461
rect 12001 1380 12073 1415
rect 17547 1603 17560 1649
rect 17606 1603 17619 1649
rect 17547 1555 17619 1603
rect 17547 1509 17560 1555
rect 17606 1509 17619 1555
rect 17547 1461 17619 1509
rect 17547 1415 17560 1461
rect 17606 1415 17619 1461
rect 17547 1380 17619 1415
rect 12001 1367 17619 1380
rect 12001 1321 12014 1367
rect 12060 1321 12108 1367
rect 12154 1321 12202 1367
rect 12248 1321 12296 1367
rect 12342 1321 12390 1367
rect 12436 1321 12484 1367
rect 12530 1321 12578 1367
rect 12624 1321 12672 1367
rect 12718 1321 12766 1367
rect 12812 1321 12860 1367
rect 12906 1321 12954 1367
rect 13000 1321 13048 1367
rect 13094 1321 13142 1367
rect 13188 1321 13236 1367
rect 13282 1321 13330 1367
rect 13376 1321 13424 1367
rect 13470 1321 13518 1367
rect 13564 1321 13612 1367
rect 13658 1321 13706 1367
rect 13752 1321 13800 1367
rect 13846 1321 13894 1367
rect 13940 1321 13988 1367
rect 14034 1321 14082 1367
rect 14128 1321 14176 1367
rect 14222 1321 14270 1367
rect 14316 1321 14364 1367
rect 14410 1321 14458 1367
rect 14504 1321 14552 1367
rect 14598 1321 14646 1367
rect 14692 1321 14740 1367
rect 14786 1321 14834 1367
rect 14880 1321 14928 1367
rect 14974 1321 15022 1367
rect 15068 1321 15116 1367
rect 15162 1321 15210 1367
rect 15256 1321 15304 1367
rect 15350 1321 15398 1367
rect 15444 1321 15492 1367
rect 15538 1321 15586 1367
rect 15632 1321 15680 1367
rect 15726 1321 15774 1367
rect 15820 1321 15868 1367
rect 15914 1321 15962 1367
rect 16008 1321 16056 1367
rect 16102 1321 16150 1367
rect 16196 1321 16244 1367
rect 16290 1321 16338 1367
rect 16384 1321 16432 1367
rect 16478 1321 16526 1367
rect 16572 1321 16620 1367
rect 16666 1321 16714 1367
rect 16760 1321 16808 1367
rect 16854 1321 16902 1367
rect 16948 1321 16996 1367
rect 17042 1321 17090 1367
rect 17136 1321 17184 1367
rect 17230 1321 17278 1367
rect 17324 1321 17372 1367
rect 17418 1321 17466 1367
rect 17512 1321 17560 1367
rect 17606 1321 17619 1367
rect 12001 1308 17619 1321
rect 5887 1265 11129 1278
<< nsubdiff >>
rect 3431 14374 5665 14387
rect 3431 14328 3444 14374
rect 3490 14328 3538 14374
rect 3584 14328 3632 14374
rect 3678 14328 3726 14374
rect 3772 14328 3820 14374
rect 3866 14328 3914 14374
rect 3960 14328 4008 14374
rect 4054 14328 4102 14374
rect 4148 14328 4196 14374
rect 4242 14328 4290 14374
rect 4336 14328 4384 14374
rect 4430 14328 4478 14374
rect 4524 14328 4572 14374
rect 4618 14328 4666 14374
rect 4712 14328 4760 14374
rect 4806 14328 4854 14374
rect 4900 14328 4948 14374
rect 4994 14328 5042 14374
rect 5088 14328 5136 14374
rect 5182 14328 5230 14374
rect 5276 14328 5324 14374
rect 5370 14328 5418 14374
rect 5464 14328 5512 14374
rect 5558 14328 5606 14374
rect 5652 14328 5665 14374
rect 3431 14315 5665 14328
rect 3431 14280 3503 14315
rect 3431 14234 3444 14280
rect 3490 14234 3503 14280
rect 3431 14186 3503 14234
rect 5593 14280 5665 14315
rect 5593 14234 5606 14280
rect 5652 14234 5665 14280
rect 3431 14140 3444 14186
rect 3490 14140 3503 14186
rect 5593 14186 5665 14234
rect 3431 14092 3503 14140
rect 3431 14046 3444 14092
rect 3490 14046 3503 14092
rect 3431 13998 3503 14046
rect 5593 14140 5606 14186
rect 5652 14140 5665 14186
rect 5593 14092 5665 14140
rect 5593 14046 5606 14092
rect 5652 14046 5665 14092
rect 3431 13952 3444 13998
rect 3490 13952 3503 13998
rect 3431 13904 3503 13952
rect 3431 13858 3444 13904
rect 3490 13858 3503 13904
rect 3431 13810 3503 13858
rect 3431 13764 3444 13810
rect 3490 13764 3503 13810
rect 3431 13716 3503 13764
rect 3431 13670 3444 13716
rect 3490 13670 3503 13716
rect 3431 13622 3503 13670
rect 3431 13576 3444 13622
rect 3490 13576 3503 13622
rect 3431 13528 3503 13576
rect 3431 13482 3444 13528
rect 3490 13482 3503 13528
rect 3431 13434 3503 13482
rect 3431 13388 3444 13434
rect 3490 13388 3503 13434
rect 3431 13340 3503 13388
rect 3431 13294 3444 13340
rect 3490 13294 3503 13340
rect 3431 13246 3503 13294
rect 5593 13998 5665 14046
rect 5593 13952 5606 13998
rect 5652 13952 5665 13998
rect 5593 13904 5665 13952
rect 5593 13858 5606 13904
rect 5652 13858 5665 13904
rect 5593 13810 5665 13858
rect 5593 13764 5606 13810
rect 5652 13764 5665 13810
rect 5593 13716 5665 13764
rect 5593 13670 5606 13716
rect 5652 13670 5665 13716
rect 5593 13622 5665 13670
rect 5593 13576 5606 13622
rect 5652 13576 5665 13622
rect 5593 13528 5665 13576
rect 5593 13482 5606 13528
rect 5652 13482 5665 13528
rect 5593 13434 5665 13482
rect 5593 13388 5606 13434
rect 5652 13388 5665 13434
rect 5593 13340 5665 13388
rect 5593 13294 5606 13340
rect 5652 13294 5665 13340
rect 3431 13200 3444 13246
rect 3490 13200 3503 13246
rect 3431 13152 3503 13200
rect 3431 13106 3444 13152
rect 3490 13106 3503 13152
rect 3431 13058 3503 13106
rect 3431 13012 3444 13058
rect 3490 13012 3503 13058
rect 3431 12964 3503 13012
rect 3431 12918 3444 12964
rect 3490 12918 3503 12964
rect 3431 12870 3503 12918
rect 5593 13246 5665 13294
rect 5593 13200 5606 13246
rect 5652 13200 5665 13246
rect 5593 13152 5665 13200
rect 5593 13106 5606 13152
rect 5652 13106 5665 13152
rect 5593 13058 5665 13106
rect 5593 13012 5606 13058
rect 5652 13012 5665 13058
rect 5593 12964 5665 13012
rect 5593 12918 5606 12964
rect 5652 12918 5665 12964
rect 3431 12824 3444 12870
rect 3490 12824 3503 12870
rect 3431 12776 3503 12824
rect 3431 12730 3444 12776
rect 3490 12730 3503 12776
rect 3431 12682 3503 12730
rect 3431 12636 3444 12682
rect 3490 12636 3503 12682
rect 3431 12588 3503 12636
rect 3431 12542 3444 12588
rect 3490 12542 3503 12588
rect 3431 12494 3503 12542
rect 3431 12448 3444 12494
rect 3490 12448 3503 12494
rect 3431 12400 3503 12448
rect 3431 12354 3444 12400
rect 3490 12354 3503 12400
rect 3431 12306 3503 12354
rect 3431 12260 3444 12306
rect 3490 12260 3503 12306
rect 3431 12212 3503 12260
rect 3431 12166 3444 12212
rect 3490 12166 3503 12212
rect 3431 12118 3503 12166
rect 5593 12870 5665 12918
rect 5593 12824 5606 12870
rect 5652 12824 5665 12870
rect 5593 12776 5665 12824
rect 5593 12730 5606 12776
rect 5652 12730 5665 12776
rect 5593 12682 5665 12730
rect 5593 12636 5606 12682
rect 5652 12636 5665 12682
rect 5593 12588 5665 12636
rect 5593 12542 5606 12588
rect 5652 12542 5665 12588
rect 5593 12494 5665 12542
rect 5593 12448 5606 12494
rect 5652 12448 5665 12494
rect 5593 12400 5665 12448
rect 5593 12354 5606 12400
rect 5652 12354 5665 12400
rect 5593 12306 5665 12354
rect 5593 12260 5606 12306
rect 5652 12260 5665 12306
rect 5593 12212 5665 12260
rect 5593 12166 5606 12212
rect 5652 12166 5665 12212
rect 3431 12072 3444 12118
rect 3490 12072 3503 12118
rect 3431 12024 3503 12072
rect 3431 11978 3444 12024
rect 3490 11978 3503 12024
rect 3431 11930 3503 11978
rect 3431 11884 3444 11930
rect 3490 11884 3503 11930
rect 3431 11836 3503 11884
rect 3431 11790 3444 11836
rect 3490 11790 3503 11836
rect 3431 11742 3503 11790
rect 5593 12118 5665 12166
rect 5593 12072 5606 12118
rect 5652 12072 5665 12118
rect 5593 12024 5665 12072
rect 5593 11978 5606 12024
rect 5652 11978 5665 12024
rect 5593 11930 5665 11978
rect 5593 11884 5606 11930
rect 5652 11884 5665 11930
rect 5593 11836 5665 11884
rect 5593 11790 5606 11836
rect 5652 11790 5665 11836
rect 3431 11696 3444 11742
rect 3490 11696 3503 11742
rect 3431 11648 3503 11696
rect 3431 11602 3444 11648
rect 3490 11602 3503 11648
rect 3431 11554 3503 11602
rect 3431 11508 3444 11554
rect 3490 11508 3503 11554
rect 3431 11460 3503 11508
rect 3431 11414 3444 11460
rect 3490 11414 3503 11460
rect 3431 11366 3503 11414
rect 3431 11320 3444 11366
rect 3490 11320 3503 11366
rect 3431 11272 3503 11320
rect 3431 11226 3444 11272
rect 3490 11226 3503 11272
rect 3431 11178 3503 11226
rect 3431 11132 3444 11178
rect 3490 11132 3503 11178
rect 3431 11084 3503 11132
rect 3431 11038 3444 11084
rect 3490 11038 3503 11084
rect 3431 10990 3503 11038
rect 5593 11742 5665 11790
rect 5593 11696 5606 11742
rect 5652 11696 5665 11742
rect 5593 11648 5665 11696
rect 5593 11602 5606 11648
rect 5652 11602 5665 11648
rect 5593 11554 5665 11602
rect 5593 11508 5606 11554
rect 5652 11508 5665 11554
rect 5593 11460 5665 11508
rect 5593 11414 5606 11460
rect 5652 11414 5665 11460
rect 5593 11366 5665 11414
rect 5593 11320 5606 11366
rect 5652 11320 5665 11366
rect 5593 11272 5665 11320
rect 5593 11226 5606 11272
rect 5652 11226 5665 11272
rect 5593 11178 5665 11226
rect 5593 11132 5606 11178
rect 5652 11132 5665 11178
rect 5593 11084 5665 11132
rect 5593 11038 5606 11084
rect 5652 11038 5665 11084
rect 3431 10944 3444 10990
rect 3490 10944 3503 10990
rect 3431 10909 3503 10944
rect 517 10896 3503 10909
rect 517 10850 530 10896
rect 576 10850 624 10896
rect 670 10850 718 10896
rect 764 10850 812 10896
rect 858 10850 906 10896
rect 952 10850 1000 10896
rect 1046 10850 1094 10896
rect 1140 10850 1188 10896
rect 1234 10850 1282 10896
rect 1328 10850 1376 10896
rect 1422 10850 1470 10896
rect 1516 10850 1564 10896
rect 1610 10850 1658 10896
rect 1704 10850 1752 10896
rect 1798 10850 1846 10896
rect 1892 10850 1940 10896
rect 1986 10850 2034 10896
rect 2080 10850 2128 10896
rect 2174 10850 2222 10896
rect 2268 10850 2316 10896
rect 2362 10850 2410 10896
rect 2456 10850 2504 10896
rect 2550 10850 2598 10896
rect 2644 10850 2692 10896
rect 2738 10850 2786 10896
rect 2832 10850 2880 10896
rect 2926 10850 2974 10896
rect 3020 10850 3068 10896
rect 3114 10850 3162 10896
rect 3208 10850 3256 10896
rect 3302 10850 3350 10896
rect 3396 10850 3444 10896
rect 3490 10850 3503 10896
rect 517 10837 3503 10850
rect 517 10802 589 10837
rect 517 10756 530 10802
rect 576 10756 589 10802
rect 517 10708 589 10756
rect -7720 10648 -3809 10665
rect -7720 10602 -7703 10648
rect -7657 10602 -7605 10648
rect -7559 10602 -7507 10648
rect -7461 10602 -7409 10648
rect -7363 10602 -7311 10648
rect -7265 10602 -7213 10648
rect -7167 10602 -7115 10648
rect -7069 10602 -7017 10648
rect -6971 10602 -6919 10648
rect -6873 10602 -6821 10648
rect -6775 10602 -6723 10648
rect -6677 10602 -6625 10648
rect -6579 10602 -6527 10648
rect -6481 10602 -6429 10648
rect -6383 10602 -6331 10648
rect -6285 10602 -6233 10648
rect -6187 10602 -6135 10648
rect -6089 10602 -6037 10648
rect -5991 10602 -5939 10648
rect -5893 10602 -5841 10648
rect -5795 10602 -5743 10648
rect -5697 10602 -5645 10648
rect -5599 10602 -5547 10648
rect -5501 10602 -5449 10648
rect -5403 10602 -5351 10648
rect -5305 10602 -5253 10648
rect -5207 10602 -5155 10648
rect -5109 10602 -5057 10648
rect -5011 10602 -4959 10648
rect -4913 10602 -4861 10648
rect -4815 10602 -4763 10648
rect -4717 10602 -4665 10648
rect -4619 10602 -4567 10648
rect -4521 10602 -4469 10648
rect -4423 10602 -4371 10648
rect -4325 10602 -4273 10648
rect -4227 10602 -4175 10648
rect -4129 10602 -4077 10648
rect -4031 10602 -3979 10648
rect -3933 10602 -3872 10648
rect -3826 10602 -3809 10648
rect -7720 10585 -3809 10602
rect -7720 10540 -7640 10585
rect -7720 10494 -7703 10540
rect -7657 10494 -7640 10540
rect -3889 10540 -3809 10585
rect -7720 10442 -7640 10494
rect -7720 10396 -7703 10442
rect -7657 10396 -7640 10442
rect -7720 10344 -7640 10396
rect -7720 10298 -7703 10344
rect -7657 10298 -7640 10344
rect -7720 10246 -7640 10298
rect -7720 10200 -7703 10246
rect -7657 10200 -7640 10246
rect -7720 10148 -7640 10200
rect -7720 10102 -7703 10148
rect -7657 10102 -7640 10148
rect -7720 10050 -7640 10102
rect -7720 10004 -7703 10050
rect -7657 10004 -7640 10050
rect -7720 9952 -7640 10004
rect -7720 9906 -7703 9952
rect -7657 9906 -7640 9952
rect -7720 9854 -7640 9906
rect -7720 9808 -7703 9854
rect -7657 9808 -7640 9854
rect -7720 9756 -7640 9808
rect -7720 9710 -7703 9756
rect -7657 9710 -7640 9756
rect -7720 9658 -7640 9710
rect -7720 9612 -7703 9658
rect -7657 9612 -7640 9658
rect -7720 9560 -7640 9612
rect -7720 9514 -7703 9560
rect -7657 9514 -7640 9560
rect -7720 9462 -7640 9514
rect -7720 9416 -7703 9462
rect -7657 9416 -7640 9462
rect -7720 9364 -7640 9416
rect -7720 9318 -7703 9364
rect -7657 9318 -7640 9364
rect -7720 9266 -7640 9318
rect -7720 9220 -7703 9266
rect -7657 9220 -7640 9266
rect -7720 9168 -7640 9220
rect -7720 9122 -7703 9168
rect -7657 9122 -7640 9168
rect -7720 9070 -7640 9122
rect -7720 9024 -7703 9070
rect -7657 9024 -7640 9070
rect -7720 8972 -7640 9024
rect -7720 8926 -7703 8972
rect -7657 8926 -7640 8972
rect -7720 8874 -7640 8926
rect -7720 8828 -7703 8874
rect -7657 8828 -7640 8874
rect -7720 8776 -7640 8828
rect -7720 8730 -7703 8776
rect -7657 8730 -7640 8776
rect -7720 8678 -7640 8730
rect -7720 8632 -7703 8678
rect -7657 8632 -7640 8678
rect -7720 8580 -7640 8632
rect -7720 8534 -7703 8580
rect -7657 8534 -7640 8580
rect -7720 8482 -7640 8534
rect -7720 8436 -7703 8482
rect -7657 8436 -7640 8482
rect -7720 8384 -7640 8436
rect -7720 8338 -7703 8384
rect -7657 8338 -7640 8384
rect -7720 8286 -7640 8338
rect -7720 8240 -7703 8286
rect -7657 8240 -7640 8286
rect -7720 8188 -7640 8240
rect -7720 8142 -7703 8188
rect -7657 8142 -7640 8188
rect -7720 8090 -7640 8142
rect -7720 8044 -7703 8090
rect -7657 8044 -7640 8090
rect -7720 7992 -7640 8044
rect -7720 7946 -7703 7992
rect -7657 7946 -7640 7992
rect -7720 7894 -7640 7946
rect -7720 7848 -7703 7894
rect -7657 7848 -7640 7894
rect -7720 7796 -7640 7848
rect -7720 7750 -7703 7796
rect -7657 7750 -7640 7796
rect -7720 7698 -7640 7750
rect -7546 10457 -3946 10529
rect -7546 9617 -7474 10457
rect -4018 9617 -3946 10457
rect -7546 9540 -3946 9617
rect -7546 8700 -7474 9540
rect -4018 8700 -3946 9540
rect -7546 8623 -3946 8700
rect -7546 7783 -7474 8623
rect -4018 7783 -3946 8623
rect -7546 7711 -3946 7783
rect -3889 10494 -3872 10540
rect -3826 10494 -3809 10540
rect -3889 10442 -3809 10494
rect -3889 10396 -3872 10442
rect -3826 10396 -3809 10442
rect -3889 10344 -3809 10396
rect -3889 10298 -3872 10344
rect -3826 10298 -3809 10344
rect -3889 10246 -3809 10298
rect -3889 10200 -3872 10246
rect -3826 10200 -3809 10246
rect -3889 10148 -3809 10200
rect -3889 10102 -3872 10148
rect -3826 10102 -3809 10148
rect -3889 10050 -3809 10102
rect -3889 10004 -3872 10050
rect -3826 10004 -3809 10050
rect -3889 9952 -3809 10004
rect -3889 9906 -3872 9952
rect -3826 9906 -3809 9952
rect -3889 9854 -3809 9906
rect -3889 9808 -3872 9854
rect -3826 9808 -3809 9854
rect -3889 9756 -3809 9808
rect -3889 9710 -3872 9756
rect -3826 9710 -3809 9756
rect -3889 9658 -3809 9710
rect -3889 9612 -3872 9658
rect -3826 9612 -3809 9658
rect -3889 9560 -3809 9612
rect -3889 9514 -3872 9560
rect -3826 9514 -3809 9560
rect -3889 9462 -3809 9514
rect -3889 9416 -3872 9462
rect -3826 9416 -3809 9462
rect -3889 9364 -3809 9416
rect -3889 9318 -3872 9364
rect -3826 9318 -3809 9364
rect -3889 9266 -3809 9318
rect -3889 9220 -3872 9266
rect -3826 9220 -3809 9266
rect -3889 9168 -3809 9220
rect -3889 9122 -3872 9168
rect -3826 9122 -3809 9168
rect -3889 9070 -3809 9122
rect -3889 9024 -3872 9070
rect -3826 9024 -3809 9070
rect -3889 8972 -3809 9024
rect -3889 8926 -3872 8972
rect -3826 8926 -3809 8972
rect -3889 8874 -3809 8926
rect -3889 8828 -3872 8874
rect -3826 8828 -3809 8874
rect -3889 8776 -3809 8828
rect -3889 8730 -3872 8776
rect -3826 8730 -3809 8776
rect -3889 8678 -3809 8730
rect -3889 8632 -3872 8678
rect -3826 8632 -3809 8678
rect -3889 8580 -3809 8632
rect -3889 8534 -3872 8580
rect -3826 8534 -3809 8580
rect -3889 8482 -3809 8534
rect -3889 8436 -3872 8482
rect -3826 8436 -3809 8482
rect -3889 8384 -3809 8436
rect -3889 8338 -3872 8384
rect -3826 8338 -3809 8384
rect -3889 8286 -3809 8338
rect -3889 8240 -3872 8286
rect -3826 8240 -3809 8286
rect -3889 8188 -3809 8240
rect -3889 8142 -3872 8188
rect -3826 8142 -3809 8188
rect -3889 8090 -3809 8142
rect -3889 8044 -3872 8090
rect -3826 8044 -3809 8090
rect -3889 7992 -3809 8044
rect -3889 7946 -3872 7992
rect -3826 7946 -3809 7992
rect -3889 7894 -3809 7946
rect -3889 7848 -3872 7894
rect -3826 7848 -3809 7894
rect -3889 7796 -3809 7848
rect -3889 7750 -3872 7796
rect -3826 7750 -3809 7796
rect -7720 7652 -7703 7698
rect -7657 7652 -7640 7698
rect -7720 7617 -7640 7652
rect -3889 7698 -3809 7750
rect -3889 7652 -3872 7698
rect -3826 7652 -3809 7698
rect -3889 7617 -3809 7652
rect -7720 7600 -3809 7617
rect -7720 7554 -7703 7600
rect -7657 7554 -7605 7600
rect -7559 7554 -7507 7600
rect -7461 7554 -7409 7600
rect -7363 7554 -7311 7600
rect -7265 7554 -7213 7600
rect -7167 7554 -7115 7600
rect -7069 7554 -7017 7600
rect -6971 7554 -6919 7600
rect -6873 7554 -6821 7600
rect -6775 7554 -6723 7600
rect -6677 7554 -6625 7600
rect -6579 7554 -6527 7600
rect -6481 7554 -6429 7600
rect -6383 7554 -6331 7600
rect -6285 7554 -6233 7600
rect -6187 7554 -6135 7600
rect -6089 7554 -6037 7600
rect -5991 7554 -5939 7600
rect -5893 7554 -5841 7600
rect -5795 7554 -5743 7600
rect -5697 7554 -5645 7600
rect -5599 7554 -5547 7600
rect -5501 7554 -5449 7600
rect -5403 7554 -5351 7600
rect -5305 7554 -5253 7600
rect -5207 7554 -5155 7600
rect -5109 7554 -5057 7600
rect -5011 7554 -4959 7600
rect -4913 7554 -4861 7600
rect -4815 7554 -4763 7600
rect -4717 7554 -4665 7600
rect -4619 7554 -4567 7600
rect -4521 7554 -4469 7600
rect -4423 7554 -4371 7600
rect -4325 7554 -4273 7600
rect -4227 7554 -4175 7600
rect -4129 7554 -4077 7600
rect -4031 7554 -3979 7600
rect -3933 7554 -3872 7600
rect -3826 7554 -3809 7600
rect -7720 7537 -3809 7554
rect 517 10662 530 10708
rect 576 10662 589 10708
rect 517 10614 589 10662
rect 517 10568 530 10614
rect 576 10568 589 10614
rect 3431 10802 3503 10837
rect 3431 10756 3444 10802
rect 3490 10756 3503 10802
rect 3431 10708 3503 10756
rect 3431 10662 3444 10708
rect 3490 10662 3503 10708
rect 3431 10614 3503 10662
rect 5593 10990 5665 11038
rect 5593 10944 5606 10990
rect 5652 10944 5665 10990
rect 5593 10896 5665 10944
rect 5593 10850 5606 10896
rect 5652 10850 5665 10896
rect 5593 10802 5665 10850
rect 5593 10756 5606 10802
rect 5652 10756 5665 10802
rect 5593 10708 5665 10756
rect 5593 10662 5606 10708
rect 5652 10662 5665 10708
rect 517 10520 589 10568
rect 3431 10568 3444 10614
rect 3490 10568 3503 10614
rect 517 10474 530 10520
rect 576 10474 589 10520
rect 517 10426 589 10474
rect 517 10380 530 10426
rect 576 10380 589 10426
rect 517 10332 589 10380
rect 517 10286 530 10332
rect 576 10286 589 10332
rect 517 10238 589 10286
rect 517 10192 530 10238
rect 576 10192 589 10238
rect 517 10144 589 10192
rect 517 10098 530 10144
rect 576 10098 589 10144
rect 517 10050 589 10098
rect 517 10004 530 10050
rect 576 10004 589 10050
rect 517 9956 589 10004
rect 517 9910 530 9956
rect 576 9910 589 9956
rect 3431 10520 3503 10568
rect 3431 10474 3444 10520
rect 3490 10474 3503 10520
rect 3431 10426 3503 10474
rect 3431 10380 3444 10426
rect 3490 10380 3503 10426
rect 3431 10332 3503 10380
rect 3431 10286 3444 10332
rect 3490 10286 3503 10332
rect 3431 10238 3503 10286
rect 3431 10192 3444 10238
rect 3490 10192 3503 10238
rect 3431 10144 3503 10192
rect 3431 10098 3444 10144
rect 3490 10098 3503 10144
rect 3431 10050 3503 10098
rect 3431 10004 3444 10050
rect 3490 10004 3503 10050
rect 3431 9956 3503 10004
rect 517 9862 589 9910
rect 517 9816 530 9862
rect 576 9816 589 9862
rect 517 9768 589 9816
rect 3431 9910 3444 9956
rect 3490 9910 3503 9956
rect 3431 9862 3503 9910
rect 5593 10614 5665 10662
rect 5593 10568 5606 10614
rect 5652 10568 5665 10614
rect 5593 10520 5665 10568
rect 5593 10474 5606 10520
rect 5652 10474 5665 10520
rect 5593 10426 5665 10474
rect 5593 10380 5606 10426
rect 5652 10380 5665 10426
rect 5593 10332 5665 10380
rect 5593 10286 5606 10332
rect 5652 10286 5665 10332
rect 5593 10238 5665 10286
rect 5593 10192 5606 10238
rect 5652 10192 5665 10238
rect 5593 10144 5665 10192
rect 5593 10098 5606 10144
rect 5652 10098 5665 10144
rect 5593 10050 5665 10098
rect 5593 10004 5606 10050
rect 5652 10004 5665 10050
rect 5593 9956 5665 10004
rect 5593 9910 5606 9956
rect 5652 9910 5665 9956
rect 3431 9816 3444 9862
rect 3490 9816 3503 9862
rect 517 9722 530 9768
rect 576 9722 589 9768
rect 517 9674 589 9722
rect 517 9628 530 9674
rect 576 9628 589 9674
rect 517 9580 589 9628
rect 517 9534 530 9580
rect 576 9534 589 9580
rect 517 9486 589 9534
rect 517 9440 530 9486
rect 576 9440 589 9486
rect 517 9392 589 9440
rect 517 9346 530 9392
rect 576 9346 589 9392
rect 517 9298 589 9346
rect 517 9252 530 9298
rect 576 9252 589 9298
rect 517 9204 589 9252
rect 517 9158 530 9204
rect 576 9158 589 9204
rect 3431 9768 3503 9816
rect 3431 9722 3444 9768
rect 3490 9722 3503 9768
rect 3431 9674 3503 9722
rect 3431 9628 3444 9674
rect 3490 9628 3503 9674
rect 3431 9580 3503 9628
rect 3431 9534 3444 9580
rect 3490 9534 3503 9580
rect 3431 9486 3503 9534
rect 5593 9862 5665 9910
rect 5593 9816 5606 9862
rect 5652 9816 5665 9862
rect 5593 9768 5665 9816
rect 5593 9722 5606 9768
rect 5652 9722 5665 9768
rect 5593 9674 5665 9722
rect 5593 9628 5606 9674
rect 5652 9628 5665 9674
rect 5593 9580 5665 9628
rect 5593 9534 5606 9580
rect 5652 9534 5665 9580
rect 3431 9440 3444 9486
rect 3490 9440 3503 9486
rect 3431 9392 3503 9440
rect 3431 9346 3444 9392
rect 3490 9346 3503 9392
rect 3431 9298 3503 9346
rect 3431 9252 3444 9298
rect 3490 9252 3503 9298
rect 3431 9204 3503 9252
rect 517 9110 589 9158
rect 517 9064 530 9110
rect 576 9064 589 9110
rect 517 9016 589 9064
rect 3431 9158 3444 9204
rect 3490 9158 3503 9204
rect 3431 9110 3503 9158
rect 3431 9064 3444 9110
rect 3490 9064 3503 9110
rect 517 8970 530 9016
rect 576 8970 589 9016
rect 517 8922 589 8970
rect 517 8876 530 8922
rect 576 8876 589 8922
rect 517 8828 589 8876
rect 517 8782 530 8828
rect 576 8782 589 8828
rect 517 8734 589 8782
rect 517 8688 530 8734
rect 576 8688 589 8734
rect 517 8640 589 8688
rect 517 8594 530 8640
rect 576 8594 589 8640
rect 517 8546 589 8594
rect 517 8500 530 8546
rect 576 8500 589 8546
rect 517 8452 589 8500
rect 517 8406 530 8452
rect 576 8406 589 8452
rect 3431 9016 3503 9064
rect 3431 8970 3444 9016
rect 3490 8970 3503 9016
rect 3431 8922 3503 8970
rect 3431 8876 3444 8922
rect 3490 8876 3503 8922
rect 3431 8828 3503 8876
rect 3431 8782 3444 8828
rect 3490 8782 3503 8828
rect 3431 8734 3503 8782
rect 5593 9486 5665 9534
rect 5593 9440 5606 9486
rect 5652 9440 5665 9486
rect 5593 9392 5665 9440
rect 5593 9346 5606 9392
rect 5652 9346 5665 9392
rect 5593 9298 5665 9346
rect 5593 9252 5606 9298
rect 5652 9252 5665 9298
rect 5593 9204 5665 9252
rect 5593 9158 5606 9204
rect 5652 9158 5665 9204
rect 5593 9110 5665 9158
rect 5593 9064 5606 9110
rect 5652 9064 5665 9110
rect 5593 9016 5665 9064
rect 5593 8970 5606 9016
rect 5652 8970 5665 9016
rect 5593 8922 5665 8970
rect 5593 8876 5606 8922
rect 5652 8876 5665 8922
rect 5593 8828 5665 8876
rect 5593 8782 5606 8828
rect 5652 8782 5665 8828
rect 3431 8688 3444 8734
rect 3490 8688 3503 8734
rect 3431 8640 3503 8688
rect 3431 8594 3444 8640
rect 3490 8594 3503 8640
rect 3431 8546 3503 8594
rect 3431 8500 3444 8546
rect 3490 8500 3503 8546
rect 5593 8734 5665 8782
rect 5593 8688 5606 8734
rect 5652 8688 5665 8734
rect 5593 8640 5665 8688
rect 3431 8452 3503 8500
rect 517 8358 589 8406
rect 517 8312 530 8358
rect 576 8312 589 8358
rect 517 8264 589 8312
rect 3431 8406 3444 8452
rect 3490 8406 3503 8452
rect 3431 8358 3503 8406
rect 5593 8594 5606 8640
rect 5652 8594 5665 8640
rect 5593 8546 5665 8594
rect 5593 8500 5606 8546
rect 5652 8500 5665 8546
rect 5593 8452 5665 8500
rect 5593 8406 5606 8452
rect 5652 8406 5665 8452
rect 3431 8312 3444 8358
rect 3490 8312 3503 8358
rect 517 8218 530 8264
rect 576 8218 589 8264
rect 517 8170 589 8218
rect 517 8124 530 8170
rect 576 8124 589 8170
rect 517 8076 589 8124
rect 517 8030 530 8076
rect 576 8030 589 8076
rect 517 7982 589 8030
rect 517 7936 530 7982
rect 576 7936 589 7982
rect 517 7888 589 7936
rect 517 7842 530 7888
rect 576 7842 589 7888
rect 517 7794 589 7842
rect 517 7748 530 7794
rect 576 7748 589 7794
rect 517 7700 589 7748
rect 517 7654 530 7700
rect 576 7654 589 7700
rect 517 7606 589 7654
rect 3431 8264 3503 8312
rect 3431 8218 3444 8264
rect 3490 8218 3503 8264
rect 3431 8170 3503 8218
rect 3431 8124 3444 8170
rect 3490 8124 3503 8170
rect 3431 8076 3503 8124
rect 3431 8030 3444 8076
rect 3490 8030 3503 8076
rect 3431 7982 3503 8030
rect 3431 7936 3444 7982
rect 3490 7936 3503 7982
rect 3431 7888 3503 7936
rect 3431 7842 3444 7888
rect 3490 7842 3503 7888
rect 3431 7794 3503 7842
rect 3431 7748 3444 7794
rect 3490 7748 3503 7794
rect 3431 7700 3503 7748
rect 3431 7654 3444 7700
rect 3490 7654 3503 7700
rect 517 7560 530 7606
rect 576 7560 589 7606
rect 517 7512 589 7560
rect 3431 7606 3503 7654
rect 5593 8358 5665 8406
rect 5593 8312 5606 8358
rect 5652 8312 5665 8358
rect 5593 8264 5665 8312
rect 5593 8218 5606 8264
rect 5652 8218 5665 8264
rect 5593 8170 5665 8218
rect 5593 8124 5606 8170
rect 5652 8124 5665 8170
rect 5593 8076 5665 8124
rect 5593 8030 5606 8076
rect 5652 8030 5665 8076
rect 5593 7982 5665 8030
rect 5593 7936 5606 7982
rect 5652 7936 5665 7982
rect 5593 7888 5665 7936
rect 5593 7842 5606 7888
rect 5652 7842 5665 7888
rect 5593 7794 5665 7842
rect 5593 7748 5606 7794
rect 5652 7748 5665 7794
rect 5593 7700 5665 7748
rect 5593 7654 5606 7700
rect 5652 7654 5665 7700
rect 3431 7560 3444 7606
rect 3490 7560 3503 7606
rect 517 7466 530 7512
rect 576 7466 589 7512
rect -7720 7438 -3809 7455
rect -7720 7392 -7703 7438
rect -7657 7392 -7605 7438
rect -7559 7392 -7507 7438
rect -7461 7392 -7409 7438
rect -7363 7392 -7311 7438
rect -7265 7392 -7213 7438
rect -7167 7392 -7115 7438
rect -7069 7392 -7017 7438
rect -6971 7392 -6919 7438
rect -6873 7392 -6821 7438
rect -6775 7392 -6723 7438
rect -6677 7392 -6625 7438
rect -6579 7392 -6527 7438
rect -6481 7392 -6429 7438
rect -6383 7392 -6331 7438
rect -6285 7392 -6233 7438
rect -6187 7392 -6135 7438
rect -6089 7392 -6037 7438
rect -5991 7392 -5939 7438
rect -5893 7392 -5841 7438
rect -5795 7392 -5743 7438
rect -5697 7392 -5645 7438
rect -5599 7392 -5547 7438
rect -5501 7392 -5449 7438
rect -5403 7392 -5351 7438
rect -5305 7392 -5253 7438
rect -5207 7392 -5155 7438
rect -5109 7392 -5057 7438
rect -5011 7392 -4959 7438
rect -4913 7392 -4861 7438
rect -4815 7392 -4763 7438
rect -4717 7392 -4665 7438
rect -4619 7392 -4567 7438
rect -4521 7392 -4469 7438
rect -4423 7392 -4371 7438
rect -4325 7392 -4273 7438
rect -4227 7392 -4175 7438
rect -4129 7392 -4077 7438
rect -4031 7392 -3979 7438
rect -3933 7392 -3872 7438
rect -3826 7392 -3809 7438
rect -7720 7375 -3809 7392
rect -7720 7340 -7640 7375
rect -7720 7294 -7703 7340
rect -7657 7294 -7640 7340
rect -7720 7242 -7640 7294
rect -3889 7340 -3809 7375
rect -3889 7294 -3872 7340
rect -3826 7294 -3809 7340
rect -7720 7196 -7703 7242
rect -7657 7196 -7640 7242
rect -7720 7144 -7640 7196
rect -7720 7098 -7703 7144
rect -7657 7098 -7640 7144
rect -7720 7046 -7640 7098
rect -7720 7000 -7703 7046
rect -7657 7000 -7640 7046
rect -7720 6948 -7640 7000
rect -7720 6902 -7703 6948
rect -7657 6902 -7640 6948
rect -7720 6850 -7640 6902
rect -7720 6804 -7703 6850
rect -7657 6804 -7640 6850
rect -7720 6752 -7640 6804
rect -7720 6706 -7703 6752
rect -7657 6706 -7640 6752
rect -7720 6654 -7640 6706
rect -7720 6608 -7703 6654
rect -7657 6608 -7640 6654
rect -7720 6556 -7640 6608
rect -7720 6510 -7703 6556
rect -7657 6510 -7640 6556
rect -7720 6458 -7640 6510
rect -7720 6412 -7703 6458
rect -7657 6412 -7640 6458
rect -7720 6360 -7640 6412
rect -7720 6314 -7703 6360
rect -7657 6314 -7640 6360
rect -7720 6262 -7640 6314
rect -7720 6216 -7703 6262
rect -7657 6216 -7640 6262
rect -7720 6164 -7640 6216
rect -7720 6118 -7703 6164
rect -7657 6118 -7640 6164
rect -7720 6066 -7640 6118
rect -7720 6020 -7703 6066
rect -7657 6020 -7640 6066
rect -7720 5968 -7640 6020
rect -7720 5922 -7703 5968
rect -7657 5922 -7640 5968
rect -7720 5870 -7640 5922
rect -7720 5824 -7703 5870
rect -7657 5824 -7640 5870
rect -7720 5772 -7640 5824
rect -7720 5726 -7703 5772
rect -7657 5726 -7640 5772
rect -7720 5674 -7640 5726
rect -7720 5628 -7703 5674
rect -7657 5628 -7640 5674
rect -7720 5576 -7640 5628
rect -7720 5530 -7703 5576
rect -7657 5530 -7640 5576
rect -7720 5478 -7640 5530
rect -7720 5432 -7703 5478
rect -7657 5432 -7640 5478
rect -7720 5380 -7640 5432
rect -7720 5334 -7703 5380
rect -7657 5334 -7640 5380
rect -7720 5282 -7640 5334
rect -7720 5236 -7703 5282
rect -7657 5236 -7640 5282
rect -7720 5184 -7640 5236
rect -7720 5138 -7703 5184
rect -7657 5138 -7640 5184
rect -7720 5086 -7640 5138
rect -7720 5040 -7703 5086
rect -7657 5040 -7640 5086
rect -7720 4988 -7640 5040
rect -7720 4942 -7703 4988
rect -7657 4942 -7640 4988
rect -7720 4890 -7640 4942
rect -7720 4844 -7703 4890
rect -7657 4844 -7640 4890
rect -7720 4792 -7640 4844
rect -7720 4746 -7703 4792
rect -7657 4746 -7640 4792
rect -7720 4694 -7640 4746
rect -7720 4648 -7703 4694
rect -7657 4648 -7640 4694
rect -7720 4596 -7640 4648
rect -7720 4550 -7703 4596
rect -7657 4550 -7640 4596
rect -7720 4498 -7640 4550
rect -7720 4452 -7703 4498
rect -7657 4452 -7640 4498
rect -7546 7209 -3946 7281
rect -7546 6369 -7474 7209
rect -4018 6369 -3946 7209
rect -7546 6292 -3946 6369
rect -7546 5452 -7474 6292
rect -4018 5452 -3946 6292
rect -7546 5375 -3946 5452
rect -7546 4535 -7474 5375
rect -4018 4535 -3946 5375
rect -7546 4463 -3946 4535
rect -3889 7242 -3809 7294
rect 517 7418 589 7466
rect 517 7372 530 7418
rect 576 7372 589 7418
rect 517 7337 589 7372
rect 3431 7512 3503 7560
rect 3431 7466 3444 7512
rect 3490 7466 3503 7512
rect 5593 7606 5665 7654
rect 5593 7560 5606 7606
rect 5652 7560 5665 7606
rect 5593 7512 5665 7560
rect 3431 7418 3503 7466
rect 5593 7466 5606 7512
rect 5652 7466 5665 7512
rect 3431 7372 3444 7418
rect 3490 7372 3503 7418
rect 3431 7337 3503 7372
rect 5593 7418 5665 7466
rect 5593 7372 5606 7418
rect 5652 7372 5665 7418
rect 5593 7337 5665 7372
rect 517 7324 5665 7337
rect 517 7278 530 7324
rect 576 7278 624 7324
rect 670 7278 718 7324
rect 764 7278 812 7324
rect 858 7278 906 7324
rect 952 7278 1000 7324
rect 1046 7278 1094 7324
rect 1140 7278 1188 7324
rect 1234 7278 1282 7324
rect 1328 7278 1376 7324
rect 1422 7278 1470 7324
rect 1516 7278 1564 7324
rect 1610 7278 1658 7324
rect 1704 7278 1752 7324
rect 1798 7278 1846 7324
rect 1892 7278 1940 7324
rect 1986 7278 2034 7324
rect 2080 7278 2128 7324
rect 2174 7278 2222 7324
rect 2268 7278 2316 7324
rect 2362 7278 2410 7324
rect 2456 7278 2504 7324
rect 2550 7278 2598 7324
rect 2644 7278 2692 7324
rect 2738 7278 2786 7324
rect 2832 7278 2880 7324
rect 2926 7278 2974 7324
rect 3020 7278 3068 7324
rect 3114 7278 3162 7324
rect 3208 7278 3256 7324
rect 3302 7278 3350 7324
rect 3396 7278 3444 7324
rect 3490 7278 3538 7324
rect 3584 7278 3632 7324
rect 3678 7278 3726 7324
rect 3772 7278 3820 7324
rect 3866 7278 3914 7324
rect 3960 7278 4008 7324
rect 4054 7278 4102 7324
rect 4148 7278 4196 7324
rect 4242 7278 4290 7324
rect 4336 7278 4384 7324
rect 4430 7278 4478 7324
rect 4524 7278 4572 7324
rect 4618 7278 4666 7324
rect 4712 7278 4760 7324
rect 4806 7278 4854 7324
rect 4900 7278 4948 7324
rect 4994 7278 5042 7324
rect 5088 7278 5136 7324
rect 5182 7278 5230 7324
rect 5276 7278 5324 7324
rect 5370 7278 5418 7324
rect 5464 7278 5512 7324
rect 5558 7278 5606 7324
rect 5652 7278 5665 7324
rect 517 7265 5665 7278
rect 11887 11742 17035 11755
rect 11887 11696 11900 11742
rect 11946 11696 11994 11742
rect 12040 11696 12088 11742
rect 12134 11696 12182 11742
rect 12228 11696 12276 11742
rect 12322 11696 12370 11742
rect 12416 11696 12464 11742
rect 12510 11696 12558 11742
rect 12604 11696 12652 11742
rect 12698 11696 12746 11742
rect 12792 11696 12840 11742
rect 12886 11696 12934 11742
rect 12980 11696 13028 11742
rect 13074 11696 13122 11742
rect 13168 11696 13216 11742
rect 13262 11696 13310 11742
rect 13356 11696 13404 11742
rect 13450 11696 13498 11742
rect 13544 11696 13592 11742
rect 13638 11696 13686 11742
rect 13732 11696 13780 11742
rect 13826 11696 13874 11742
rect 13920 11696 13968 11742
rect 14014 11696 14062 11742
rect 14108 11696 14156 11742
rect 14202 11696 14250 11742
rect 14296 11696 14344 11742
rect 14390 11696 14438 11742
rect 14484 11696 14532 11742
rect 14578 11696 14626 11742
rect 14672 11696 14720 11742
rect 14766 11696 14814 11742
rect 14860 11696 14908 11742
rect 14954 11696 15002 11742
rect 15048 11696 15096 11742
rect 15142 11696 15190 11742
rect 15236 11696 15284 11742
rect 15330 11696 15378 11742
rect 15424 11696 15472 11742
rect 15518 11696 15566 11742
rect 15612 11696 15660 11742
rect 15706 11696 15754 11742
rect 15800 11696 15848 11742
rect 15894 11696 15942 11742
rect 15988 11696 16036 11742
rect 16082 11696 16130 11742
rect 16176 11696 16224 11742
rect 16270 11696 16318 11742
rect 16364 11696 16412 11742
rect 16458 11696 16506 11742
rect 16552 11696 16600 11742
rect 16646 11696 16694 11742
rect 16740 11696 16788 11742
rect 16834 11696 16882 11742
rect 16928 11696 16976 11742
rect 17022 11696 17035 11742
rect 11887 11683 17035 11696
rect 11887 11648 11959 11683
rect 11887 11602 11900 11648
rect 11946 11602 11959 11648
rect 11887 11554 11959 11602
rect 11887 11508 11900 11554
rect 11946 11508 11959 11554
rect 11887 11460 11959 11508
rect 11887 11414 11900 11460
rect 11946 11414 11959 11460
rect 14613 11648 14685 11683
rect 14613 11602 14626 11648
rect 14672 11602 14685 11648
rect 14613 11554 14685 11602
rect 14613 11508 14626 11554
rect 14672 11508 14685 11554
rect 14613 11460 14685 11508
rect 11887 11366 11959 11414
rect 14613 11414 14626 11460
rect 14672 11414 14685 11460
rect 16963 11648 17035 11683
rect 16963 11602 16976 11648
rect 17022 11602 17035 11648
rect 16963 11554 17035 11602
rect 16963 11508 16976 11554
rect 17022 11508 17035 11554
rect 16963 11460 17035 11508
rect 11887 11320 11900 11366
rect 11946 11320 11959 11366
rect 11887 11272 11959 11320
rect 11887 11226 11900 11272
rect 11946 11226 11959 11272
rect 11887 11178 11959 11226
rect 11887 11132 11900 11178
rect 11946 11132 11959 11178
rect 11887 11084 11959 11132
rect 11887 11038 11900 11084
rect 11946 11038 11959 11084
rect 11887 10990 11959 11038
rect 11887 10944 11900 10990
rect 11946 10944 11959 10990
rect 11887 10896 11959 10944
rect 11887 10850 11900 10896
rect 11946 10850 11959 10896
rect 11887 10802 11959 10850
rect 11887 10756 11900 10802
rect 11946 10756 11959 10802
rect 11887 10708 11959 10756
rect 14613 11366 14685 11414
rect 16963 11414 16976 11460
rect 17022 11414 17035 11460
rect 14613 11320 14626 11366
rect 14672 11320 14685 11366
rect 14613 11272 14685 11320
rect 14613 11226 14626 11272
rect 14672 11226 14685 11272
rect 14613 11178 14685 11226
rect 14613 11132 14626 11178
rect 14672 11132 14685 11178
rect 14613 11084 14685 11132
rect 14613 11038 14626 11084
rect 14672 11038 14685 11084
rect 14613 10990 14685 11038
rect 14613 10944 14626 10990
rect 14672 10944 14685 10990
rect 14613 10896 14685 10944
rect 14613 10850 14626 10896
rect 14672 10850 14685 10896
rect 14613 10802 14685 10850
rect 14613 10756 14626 10802
rect 14672 10756 14685 10802
rect 11887 10662 11900 10708
rect 11946 10662 11959 10708
rect 11887 10614 11959 10662
rect 11887 10568 11900 10614
rect 11946 10568 11959 10614
rect 11887 10520 11959 10568
rect 11887 10474 11900 10520
rect 11946 10474 11959 10520
rect 11887 10426 11959 10474
rect 11887 10380 11900 10426
rect 11946 10380 11959 10426
rect 11887 10332 11959 10380
rect 14613 10708 14685 10756
rect 16963 11366 17035 11414
rect 16963 11320 16976 11366
rect 17022 11320 17035 11366
rect 16963 11272 17035 11320
rect 16963 11226 16976 11272
rect 17022 11226 17035 11272
rect 16963 11178 17035 11226
rect 16963 11132 16976 11178
rect 17022 11132 17035 11178
rect 16963 11084 17035 11132
rect 16963 11038 16976 11084
rect 17022 11038 17035 11084
rect 16963 10990 17035 11038
rect 16963 10944 16976 10990
rect 17022 10944 17035 10990
rect 16963 10896 17035 10944
rect 16963 10850 16976 10896
rect 17022 10850 17035 10896
rect 16963 10802 17035 10850
rect 16963 10756 16976 10802
rect 17022 10756 17035 10802
rect 14613 10662 14626 10708
rect 14672 10662 14685 10708
rect 14613 10614 14685 10662
rect 14613 10568 14626 10614
rect 14672 10568 14685 10614
rect 14613 10520 14685 10568
rect 14613 10474 14626 10520
rect 14672 10474 14685 10520
rect 14613 10426 14685 10474
rect 14613 10380 14626 10426
rect 14672 10380 14685 10426
rect 11887 10286 11900 10332
rect 11946 10286 11959 10332
rect 11887 10238 11959 10286
rect 11887 10192 11900 10238
rect 11946 10192 11959 10238
rect 11887 10144 11959 10192
rect 11887 10098 11900 10144
rect 11946 10098 11959 10144
rect 11887 10050 11959 10098
rect 11887 10004 11900 10050
rect 11946 10004 11959 10050
rect 11887 9956 11959 10004
rect 11887 9910 11900 9956
rect 11946 9910 11959 9956
rect 11887 9862 11959 9910
rect 11887 9816 11900 9862
rect 11946 9816 11959 9862
rect 11887 9768 11959 9816
rect 11887 9722 11900 9768
rect 11946 9722 11959 9768
rect 11887 9674 11959 9722
rect 14613 10332 14685 10380
rect 16963 10708 17035 10756
rect 16963 10662 16976 10708
rect 17022 10662 17035 10708
rect 16963 10614 17035 10662
rect 16963 10568 16976 10614
rect 17022 10568 17035 10614
rect 16963 10520 17035 10568
rect 16963 10474 16976 10520
rect 17022 10474 17035 10520
rect 16963 10426 17035 10474
rect 16963 10380 16976 10426
rect 17022 10380 17035 10426
rect 14613 10286 14626 10332
rect 14672 10286 14685 10332
rect 14613 10238 14685 10286
rect 14613 10192 14626 10238
rect 14672 10192 14685 10238
rect 14613 10144 14685 10192
rect 14613 10098 14626 10144
rect 14672 10098 14685 10144
rect 14613 10050 14685 10098
rect 14613 10004 14626 10050
rect 14672 10004 14685 10050
rect 14613 9956 14685 10004
rect 14613 9910 14626 9956
rect 14672 9910 14685 9956
rect 14613 9862 14685 9910
rect 14613 9816 14626 9862
rect 14672 9816 14685 9862
rect 14613 9768 14685 9816
rect 14613 9722 14626 9768
rect 14672 9722 14685 9768
rect 11887 9628 11900 9674
rect 11946 9628 11959 9674
rect 11887 9580 11959 9628
rect 11887 9534 11900 9580
rect 11946 9534 11959 9580
rect 11887 9486 11959 9534
rect 11887 9440 11900 9486
rect 11946 9440 11959 9486
rect 11887 9392 11959 9440
rect 11887 9346 11900 9392
rect 11946 9346 11959 9392
rect 11887 9298 11959 9346
rect 14613 9674 14685 9722
rect 16963 10332 17035 10380
rect 16963 10286 16976 10332
rect 17022 10286 17035 10332
rect 16963 10238 17035 10286
rect 16963 10192 16976 10238
rect 17022 10192 17035 10238
rect 16963 10144 17035 10192
rect 16963 10098 16976 10144
rect 17022 10098 17035 10144
rect 16963 10050 17035 10098
rect 16963 10004 16976 10050
rect 17022 10004 17035 10050
rect 16963 9956 17035 10004
rect 16963 9910 16976 9956
rect 17022 9910 17035 9956
rect 16963 9862 17035 9910
rect 16963 9816 16976 9862
rect 17022 9816 17035 9862
rect 16963 9768 17035 9816
rect 16963 9722 16976 9768
rect 17022 9722 17035 9768
rect 14613 9628 14626 9674
rect 14672 9628 14685 9674
rect 14613 9580 14685 9628
rect 14613 9534 14626 9580
rect 14672 9534 14685 9580
rect 14613 9486 14685 9534
rect 14613 9440 14626 9486
rect 14672 9440 14685 9486
rect 14613 9392 14685 9440
rect 14613 9346 14626 9392
rect 14672 9346 14685 9392
rect 11887 9252 11900 9298
rect 11946 9252 11959 9298
rect 11887 9204 11959 9252
rect 11887 9158 11900 9204
rect 11946 9158 11959 9204
rect 11887 9110 11959 9158
rect 11887 9064 11900 9110
rect 11946 9064 11959 9110
rect 11887 9016 11959 9064
rect 11887 8970 11900 9016
rect 11946 8970 11959 9016
rect 11887 8922 11959 8970
rect 11887 8876 11900 8922
rect 11946 8876 11959 8922
rect 11887 8828 11959 8876
rect 11887 8782 11900 8828
rect 11946 8782 11959 8828
rect 11887 8734 11959 8782
rect 11887 8688 11900 8734
rect 11946 8688 11959 8734
rect 11887 8640 11959 8688
rect 14613 9298 14685 9346
rect 16963 9674 17035 9722
rect 16963 9628 16976 9674
rect 17022 9628 17035 9674
rect 16963 9580 17035 9628
rect 16963 9534 16976 9580
rect 17022 9534 17035 9580
rect 16963 9486 17035 9534
rect 16963 9440 16976 9486
rect 17022 9440 17035 9486
rect 16963 9392 17035 9440
rect 16963 9346 16976 9392
rect 17022 9346 17035 9392
rect 14613 9252 14626 9298
rect 14672 9252 14685 9298
rect 14613 9204 14685 9252
rect 14613 9158 14626 9204
rect 14672 9158 14685 9204
rect 14613 9110 14685 9158
rect 14613 9064 14626 9110
rect 14672 9064 14685 9110
rect 14613 9016 14685 9064
rect 14613 8970 14626 9016
rect 14672 8970 14685 9016
rect 14613 8922 14685 8970
rect 14613 8876 14626 8922
rect 14672 8876 14685 8922
rect 14613 8828 14685 8876
rect 14613 8782 14626 8828
rect 14672 8782 14685 8828
rect 14613 8734 14685 8782
rect 14613 8688 14626 8734
rect 14672 8688 14685 8734
rect 11887 8594 11900 8640
rect 11946 8594 11959 8640
rect 11887 8546 11959 8594
rect 11887 8500 11900 8546
rect 11946 8500 11959 8546
rect 11887 8452 11959 8500
rect 11887 8406 11900 8452
rect 11946 8406 11959 8452
rect 11887 8358 11959 8406
rect 14613 8640 14685 8688
rect 16963 9298 17035 9346
rect 16963 9252 16976 9298
rect 17022 9252 17035 9298
rect 16963 9204 17035 9252
rect 16963 9158 16976 9204
rect 17022 9158 17035 9204
rect 16963 9110 17035 9158
rect 16963 9064 16976 9110
rect 17022 9064 17035 9110
rect 16963 9016 17035 9064
rect 16963 8970 16976 9016
rect 17022 8970 17035 9016
rect 16963 8922 17035 8970
rect 16963 8876 16976 8922
rect 17022 8876 17035 8922
rect 16963 8828 17035 8876
rect 16963 8782 16976 8828
rect 17022 8782 17035 8828
rect 16963 8734 17035 8782
rect 16963 8688 16976 8734
rect 17022 8688 17035 8734
rect 14613 8594 14626 8640
rect 14672 8594 14685 8640
rect 14613 8546 14685 8594
rect 14613 8500 14626 8546
rect 14672 8500 14685 8546
rect 14613 8452 14685 8500
rect 11887 8312 11900 8358
rect 11946 8312 11959 8358
rect 11887 8264 11959 8312
rect 14613 8406 14626 8452
rect 14672 8406 14685 8452
rect 14613 8358 14685 8406
rect 16963 8640 17035 8688
rect 16963 8594 16976 8640
rect 17022 8594 17035 8640
rect 16963 8546 17035 8594
rect 16963 8500 16976 8546
rect 17022 8500 17035 8546
rect 16963 8452 17035 8500
rect 14613 8312 14626 8358
rect 14672 8312 14685 8358
rect 11887 8218 11900 8264
rect 11946 8218 11959 8264
rect 11887 8170 11959 8218
rect 11887 8124 11900 8170
rect 11946 8124 11959 8170
rect 11887 8076 11959 8124
rect 11887 8030 11900 8076
rect 11946 8030 11959 8076
rect 11887 7982 11959 8030
rect 11887 7936 11900 7982
rect 11946 7936 11959 7982
rect 11887 7888 11959 7936
rect 11887 7842 11900 7888
rect 11946 7842 11959 7888
rect 11887 7794 11959 7842
rect 11887 7748 11900 7794
rect 11946 7748 11959 7794
rect 11887 7700 11959 7748
rect 11887 7654 11900 7700
rect 11946 7654 11959 7700
rect 11887 7606 11959 7654
rect 14613 8264 14685 8312
rect 16963 8406 16976 8452
rect 17022 8406 17035 8452
rect 16963 8358 17035 8406
rect 16963 8312 16976 8358
rect 17022 8312 17035 8358
rect 14613 8218 14626 8264
rect 14672 8218 14685 8264
rect 14613 8170 14685 8218
rect 14613 8124 14626 8170
rect 14672 8124 14685 8170
rect 14613 8076 14685 8124
rect 14613 8030 14626 8076
rect 14672 8030 14685 8076
rect 14613 7982 14685 8030
rect 14613 7936 14626 7982
rect 14672 7936 14685 7982
rect 14613 7888 14685 7936
rect 14613 7842 14626 7888
rect 14672 7842 14685 7888
rect 14613 7794 14685 7842
rect 14613 7748 14626 7794
rect 14672 7748 14685 7794
rect 14613 7700 14685 7748
rect 14613 7654 14626 7700
rect 14672 7654 14685 7700
rect 11887 7560 11900 7606
rect 11946 7560 11959 7606
rect 14613 7606 14685 7654
rect 16963 8264 17035 8312
rect 16963 8218 16976 8264
rect 17022 8218 17035 8264
rect 16963 8170 17035 8218
rect 16963 8124 16976 8170
rect 17022 8124 17035 8170
rect 16963 8076 17035 8124
rect 16963 8030 16976 8076
rect 17022 8030 17035 8076
rect 16963 7982 17035 8030
rect 16963 7936 16976 7982
rect 17022 7936 17035 7982
rect 16963 7888 17035 7936
rect 16963 7842 16976 7888
rect 17022 7842 17035 7888
rect 16963 7794 17035 7842
rect 16963 7748 16976 7794
rect 17022 7748 17035 7794
rect 16963 7700 17035 7748
rect 16963 7654 16976 7700
rect 17022 7654 17035 7700
rect 11887 7512 11959 7560
rect 11887 7466 11900 7512
rect 11946 7466 11959 7512
rect 11887 7418 11959 7466
rect 11887 7372 11900 7418
rect 11946 7372 11959 7418
rect 11887 7337 11959 7372
rect 14613 7560 14626 7606
rect 14672 7560 14685 7606
rect 16963 7606 17035 7654
rect 14613 7512 14685 7560
rect 14613 7466 14626 7512
rect 14672 7466 14685 7512
rect 14613 7418 14685 7466
rect 14613 7372 14626 7418
rect 14672 7372 14685 7418
rect 14613 7337 14685 7372
rect 16963 7560 16976 7606
rect 17022 7560 17035 7606
rect 16963 7512 17035 7560
rect 16963 7466 16976 7512
rect 17022 7466 17035 7512
rect 16963 7418 17035 7466
rect 16963 7372 16976 7418
rect 17022 7372 17035 7418
rect 16963 7337 17035 7372
rect 11887 7324 17035 7337
rect 11887 7278 11900 7324
rect 11946 7278 11994 7324
rect 12040 7278 12088 7324
rect 12134 7278 12182 7324
rect 12228 7278 12276 7324
rect 12322 7278 12370 7324
rect 12416 7278 12464 7324
rect 12510 7278 12558 7324
rect 12604 7278 12652 7324
rect 12698 7278 12746 7324
rect 12792 7278 12840 7324
rect 12886 7278 12934 7324
rect 12980 7278 13028 7324
rect 13074 7278 13122 7324
rect 13168 7278 13216 7324
rect 13262 7278 13310 7324
rect 13356 7278 13404 7324
rect 13450 7278 13498 7324
rect 13544 7278 13592 7324
rect 13638 7278 13686 7324
rect 13732 7278 13780 7324
rect 13826 7278 13874 7324
rect 13920 7278 13968 7324
rect 14014 7278 14062 7324
rect 14108 7278 14156 7324
rect 14202 7278 14250 7324
rect 14296 7278 14344 7324
rect 14390 7278 14438 7324
rect 14484 7278 14532 7324
rect 14578 7278 14626 7324
rect 14672 7278 14720 7324
rect 14766 7278 14814 7324
rect 14860 7278 14908 7324
rect 14954 7278 15002 7324
rect 15048 7278 15096 7324
rect 15142 7278 15190 7324
rect 15236 7278 15284 7324
rect 15330 7278 15378 7324
rect 15424 7278 15472 7324
rect 15518 7278 15566 7324
rect 15612 7278 15660 7324
rect 15706 7278 15754 7324
rect 15800 7278 15848 7324
rect 15894 7278 15942 7324
rect 15988 7278 16036 7324
rect 16082 7278 16130 7324
rect 16176 7278 16224 7324
rect 16270 7278 16318 7324
rect 16364 7278 16412 7324
rect 16458 7278 16506 7324
rect 16552 7278 16600 7324
rect 16646 7278 16694 7324
rect 16740 7278 16788 7324
rect 16834 7278 16882 7324
rect 16928 7278 16976 7324
rect 17022 7278 17035 7324
rect 32616 12219 40960 12232
rect 32616 12173 32629 12219
rect 32675 12173 32723 12219
rect 32769 12173 32817 12219
rect 32863 12173 32911 12219
rect 32957 12173 33005 12219
rect 33051 12173 33099 12219
rect 33145 12173 33193 12219
rect 33239 12173 33287 12219
rect 33333 12173 33381 12219
rect 33427 12173 33475 12219
rect 33521 12173 33569 12219
rect 33615 12173 33663 12219
rect 33709 12173 33757 12219
rect 33803 12173 33851 12219
rect 33897 12173 33945 12219
rect 33991 12173 34039 12219
rect 34085 12173 34133 12219
rect 34179 12173 34227 12219
rect 34273 12173 34321 12219
rect 34367 12173 34415 12219
rect 34461 12173 34509 12219
rect 34555 12173 34603 12219
rect 34649 12173 34697 12219
rect 34743 12173 34791 12219
rect 34837 12173 34885 12219
rect 34931 12173 34979 12219
rect 35025 12173 35073 12219
rect 35119 12173 35167 12219
rect 35213 12173 35261 12219
rect 35307 12173 35355 12219
rect 35401 12173 35449 12219
rect 35495 12173 35543 12219
rect 35589 12173 35637 12219
rect 35683 12173 35731 12219
rect 35777 12173 35825 12219
rect 35871 12173 35919 12219
rect 35965 12173 36013 12219
rect 36059 12173 36107 12219
rect 36153 12173 36201 12219
rect 36247 12173 36295 12219
rect 36341 12173 36389 12219
rect 36435 12173 36483 12219
rect 36529 12173 36577 12219
rect 36623 12173 36671 12219
rect 36717 12173 36765 12219
rect 36811 12173 36859 12219
rect 36905 12173 36953 12219
rect 36999 12173 37047 12219
rect 37093 12173 37141 12219
rect 37187 12173 37235 12219
rect 37281 12173 37329 12219
rect 37375 12173 37423 12219
rect 37469 12173 37517 12219
rect 37563 12173 37611 12219
rect 37657 12173 37705 12219
rect 37751 12173 37799 12219
rect 37845 12173 37893 12219
rect 37939 12173 37987 12219
rect 38033 12173 38081 12219
rect 38127 12173 38175 12219
rect 38221 12173 38269 12219
rect 38315 12173 38363 12219
rect 38409 12173 38457 12219
rect 38503 12173 38551 12219
rect 38597 12173 38645 12219
rect 38691 12173 38739 12219
rect 38785 12173 38833 12219
rect 38879 12173 38927 12219
rect 38973 12173 39021 12219
rect 39067 12173 39115 12219
rect 39161 12173 39209 12219
rect 39255 12173 39303 12219
rect 39349 12173 39397 12219
rect 39443 12173 39491 12219
rect 39537 12173 39585 12219
rect 39631 12173 39679 12219
rect 39725 12173 39773 12219
rect 39819 12173 39867 12219
rect 39913 12173 39961 12219
rect 40007 12173 40055 12219
rect 40101 12173 40149 12219
rect 40195 12173 40243 12219
rect 40289 12173 40337 12219
rect 40383 12173 40431 12219
rect 40477 12173 40525 12219
rect 40571 12173 40619 12219
rect 40665 12173 40713 12219
rect 40759 12173 40807 12219
rect 40853 12173 40901 12219
rect 40947 12173 40960 12219
rect 32616 12160 40960 12173
rect 32616 12125 32688 12160
rect 32616 12079 32629 12125
rect 32675 12079 32688 12125
rect 32616 12031 32688 12079
rect 32616 11985 32629 12031
rect 32675 11985 32688 12031
rect 32616 11937 32688 11985
rect 32616 11891 32629 11937
rect 32675 11891 32688 11937
rect 32616 11843 32688 11891
rect 32616 11797 32629 11843
rect 32675 11797 32688 11843
rect 36752 12125 36824 12160
rect 36752 12079 36765 12125
rect 36811 12079 36824 12125
rect 36752 12031 36824 12079
rect 36752 11985 36765 12031
rect 36811 11985 36824 12031
rect 36752 11937 36824 11985
rect 36752 11891 36765 11937
rect 36811 11891 36824 11937
rect 36752 11843 36824 11891
rect 32616 11749 32688 11797
rect 36752 11797 36765 11843
rect 36811 11797 36824 11843
rect 40888 12125 40960 12160
rect 40888 12079 40901 12125
rect 40947 12079 40960 12125
rect 40888 12031 40960 12079
rect 40888 11985 40901 12031
rect 40947 11985 40960 12031
rect 40888 11937 40960 11985
rect 40888 11891 40901 11937
rect 40947 11891 40960 11937
rect 40888 11843 40960 11891
rect 32616 11703 32629 11749
rect 32675 11703 32688 11749
rect 32616 11655 32688 11703
rect 36752 11749 36824 11797
rect 40888 11797 40901 11843
rect 40947 11797 40960 11843
rect 36752 11703 36765 11749
rect 36811 11703 36824 11749
rect 32616 11609 32629 11655
rect 32675 11609 32688 11655
rect 32616 11561 32688 11609
rect 32616 11515 32629 11561
rect 32675 11515 32688 11561
rect 32616 11467 32688 11515
rect 32616 11421 32629 11467
rect 32675 11421 32688 11467
rect 32616 11373 32688 11421
rect 32616 11327 32629 11373
rect 32675 11327 32688 11373
rect 32616 11279 32688 11327
rect 32616 11233 32629 11279
rect 32675 11233 32688 11279
rect 32616 11185 32688 11233
rect 32616 11139 32629 11185
rect 32675 11139 32688 11185
rect 32616 11091 32688 11139
rect 32616 11045 32629 11091
rect 32675 11045 32688 11091
rect 36752 11655 36824 11703
rect 40888 11749 40960 11797
rect 40888 11703 40901 11749
rect 40947 11703 40960 11749
rect 36752 11609 36765 11655
rect 36811 11609 36824 11655
rect 36752 11561 36824 11609
rect 36752 11515 36765 11561
rect 36811 11515 36824 11561
rect 36752 11467 36824 11515
rect 36752 11421 36765 11467
rect 36811 11421 36824 11467
rect 36752 11373 36824 11421
rect 36752 11327 36765 11373
rect 36811 11327 36824 11373
rect 36752 11279 36824 11327
rect 36752 11233 36765 11279
rect 36811 11233 36824 11279
rect 36752 11185 36824 11233
rect 36752 11139 36765 11185
rect 36811 11139 36824 11185
rect 36752 11091 36824 11139
rect 32616 10997 32688 11045
rect 32616 10951 32629 10997
rect 32675 10951 32688 10997
rect 32616 10903 32688 10951
rect 32616 10857 32629 10903
rect 32675 10857 32688 10903
rect 32616 10809 32688 10857
rect 32616 10763 32629 10809
rect 32675 10763 32688 10809
rect 32616 10715 32688 10763
rect 32616 10669 32629 10715
rect 32675 10669 32688 10715
rect 32616 10621 32688 10669
rect 36752 11045 36765 11091
rect 36811 11045 36824 11091
rect 40888 11655 40960 11703
rect 40888 11609 40901 11655
rect 40947 11609 40960 11655
rect 40888 11561 40960 11609
rect 40888 11515 40901 11561
rect 40947 11515 40960 11561
rect 40888 11467 40960 11515
rect 40888 11421 40901 11467
rect 40947 11421 40960 11467
rect 40888 11373 40960 11421
rect 40888 11327 40901 11373
rect 40947 11327 40960 11373
rect 40888 11279 40960 11327
rect 40888 11233 40901 11279
rect 40947 11233 40960 11279
rect 40888 11185 40960 11233
rect 40888 11139 40901 11185
rect 40947 11139 40960 11185
rect 40888 11091 40960 11139
rect 36752 10997 36824 11045
rect 36752 10951 36765 10997
rect 36811 10951 36824 10997
rect 36752 10903 36824 10951
rect 36752 10857 36765 10903
rect 36811 10857 36824 10903
rect 36752 10809 36824 10857
rect 36752 10763 36765 10809
rect 36811 10763 36824 10809
rect 36752 10715 36824 10763
rect 36752 10669 36765 10715
rect 36811 10669 36824 10715
rect 32616 10575 32629 10621
rect 32675 10575 32688 10621
rect 32616 10527 32688 10575
rect 32616 10481 32629 10527
rect 32675 10481 32688 10527
rect 32616 10433 32688 10481
rect 32616 10387 32629 10433
rect 32675 10387 32688 10433
rect 32616 10339 32688 10387
rect 32616 10293 32629 10339
rect 32675 10293 32688 10339
rect 32616 10245 32688 10293
rect 32616 10199 32629 10245
rect 32675 10199 32688 10245
rect 32616 10151 32688 10199
rect 32616 10105 32629 10151
rect 32675 10105 32688 10151
rect 32616 10057 32688 10105
rect 32616 10011 32629 10057
rect 32675 10011 32688 10057
rect 36752 10621 36824 10669
rect 40888 11045 40901 11091
rect 40947 11045 40960 11091
rect 40888 10997 40960 11045
rect 40888 10951 40901 10997
rect 40947 10951 40960 10997
rect 40888 10903 40960 10951
rect 40888 10857 40901 10903
rect 40947 10857 40960 10903
rect 40888 10809 40960 10857
rect 40888 10763 40901 10809
rect 40947 10763 40960 10809
rect 40888 10715 40960 10763
rect 40888 10669 40901 10715
rect 40947 10669 40960 10715
rect 36752 10575 36765 10621
rect 36811 10575 36824 10621
rect 36752 10527 36824 10575
rect 36752 10481 36765 10527
rect 36811 10481 36824 10527
rect 36752 10433 36824 10481
rect 36752 10387 36765 10433
rect 36811 10387 36824 10433
rect 36752 10339 36824 10387
rect 36752 10293 36765 10339
rect 36811 10293 36824 10339
rect 36752 10245 36824 10293
rect 36752 10199 36765 10245
rect 36811 10199 36824 10245
rect 36752 10151 36824 10199
rect 36752 10105 36765 10151
rect 36811 10105 36824 10151
rect 36752 10057 36824 10105
rect 32616 9963 32688 10011
rect 32616 9917 32629 9963
rect 32675 9917 32688 9963
rect 32616 9869 32688 9917
rect 32616 9823 32629 9869
rect 32675 9823 32688 9869
rect 32616 9775 32688 9823
rect 32616 9729 32629 9775
rect 32675 9729 32688 9775
rect 32616 9681 32688 9729
rect 32616 9635 32629 9681
rect 32675 9635 32688 9681
rect 32616 9587 32688 9635
rect 32616 9541 32629 9587
rect 32675 9541 32688 9587
rect 36752 10011 36765 10057
rect 36811 10011 36824 10057
rect 40888 10621 40960 10669
rect 40888 10575 40901 10621
rect 40947 10575 40960 10621
rect 40888 10527 40960 10575
rect 40888 10481 40901 10527
rect 40947 10481 40960 10527
rect 40888 10433 40960 10481
rect 40888 10387 40901 10433
rect 40947 10387 40960 10433
rect 40888 10339 40960 10387
rect 40888 10293 40901 10339
rect 40947 10293 40960 10339
rect 40888 10245 40960 10293
rect 40888 10199 40901 10245
rect 40947 10199 40960 10245
rect 40888 10151 40960 10199
rect 40888 10105 40901 10151
rect 40947 10105 40960 10151
rect 40888 10057 40960 10105
rect 36752 9963 36824 10011
rect 36752 9917 36765 9963
rect 36811 9917 36824 9963
rect 36752 9869 36824 9917
rect 36752 9823 36765 9869
rect 36811 9823 36824 9869
rect 36752 9775 36824 9823
rect 36752 9729 36765 9775
rect 36811 9729 36824 9775
rect 36752 9681 36824 9729
rect 36752 9635 36765 9681
rect 36811 9635 36824 9681
rect 36752 9587 36824 9635
rect 32616 9493 32688 9541
rect 32616 9447 32629 9493
rect 32675 9447 32688 9493
rect 32616 9399 32688 9447
rect 32616 9353 32629 9399
rect 32675 9353 32688 9399
rect 32616 9305 32688 9353
rect 32616 9259 32629 9305
rect 32675 9259 32688 9305
rect 32616 9211 32688 9259
rect 32616 9165 32629 9211
rect 32675 9165 32688 9211
rect 32616 9117 32688 9165
rect 32616 9071 32629 9117
rect 32675 9071 32688 9117
rect 32616 9023 32688 9071
rect 32616 8977 32629 9023
rect 32675 8977 32688 9023
rect 32616 8929 32688 8977
rect 36752 9541 36765 9587
rect 36811 9541 36824 9587
rect 40888 10011 40901 10057
rect 40947 10011 40960 10057
rect 40888 9963 40960 10011
rect 40888 9917 40901 9963
rect 40947 9917 40960 9963
rect 40888 9869 40960 9917
rect 40888 9823 40901 9869
rect 40947 9823 40960 9869
rect 40888 9775 40960 9823
rect 40888 9729 40901 9775
rect 40947 9729 40960 9775
rect 40888 9681 40960 9729
rect 40888 9635 40901 9681
rect 40947 9635 40960 9681
rect 40888 9587 40960 9635
rect 36752 9493 36824 9541
rect 36752 9447 36765 9493
rect 36811 9447 36824 9493
rect 36752 9399 36824 9447
rect 36752 9353 36765 9399
rect 36811 9353 36824 9399
rect 36752 9305 36824 9353
rect 36752 9259 36765 9305
rect 36811 9259 36824 9305
rect 36752 9211 36824 9259
rect 36752 9165 36765 9211
rect 36811 9165 36824 9211
rect 36752 9117 36824 9165
rect 36752 9071 36765 9117
rect 36811 9071 36824 9117
rect 36752 9023 36824 9071
rect 36752 8977 36765 9023
rect 36811 8977 36824 9023
rect 32616 8883 32629 8929
rect 32675 8883 32688 8929
rect 32616 8835 32688 8883
rect 32616 8789 32629 8835
rect 32675 8789 32688 8835
rect 32616 8741 32688 8789
rect 32616 8695 32629 8741
rect 32675 8695 32688 8741
rect 32616 8647 32688 8695
rect 32616 8601 32629 8647
rect 32675 8601 32688 8647
rect 32616 8553 32688 8601
rect 32616 8507 32629 8553
rect 32675 8507 32688 8553
rect 36752 8929 36824 8977
rect 40888 9541 40901 9587
rect 40947 9541 40960 9587
rect 40888 9493 40960 9541
rect 40888 9447 40901 9493
rect 40947 9447 40960 9493
rect 40888 9399 40960 9447
rect 40888 9353 40901 9399
rect 40947 9353 40960 9399
rect 40888 9305 40960 9353
rect 40888 9259 40901 9305
rect 40947 9259 40960 9305
rect 40888 9211 40960 9259
rect 40888 9165 40901 9211
rect 40947 9165 40960 9211
rect 40888 9117 40960 9165
rect 40888 9071 40901 9117
rect 40947 9071 40960 9117
rect 40888 9023 40960 9071
rect 40888 8977 40901 9023
rect 40947 8977 40960 9023
rect 36752 8883 36765 8929
rect 36811 8883 36824 8929
rect 36752 8835 36824 8883
rect 36752 8789 36765 8835
rect 36811 8789 36824 8835
rect 36752 8741 36824 8789
rect 36752 8695 36765 8741
rect 36811 8695 36824 8741
rect 36752 8647 36824 8695
rect 36752 8601 36765 8647
rect 36811 8601 36824 8647
rect 36752 8553 36824 8601
rect 32616 8459 32688 8507
rect 32616 8413 32629 8459
rect 32675 8413 32688 8459
rect 32616 8365 32688 8413
rect 32616 8319 32629 8365
rect 32675 8319 32688 8365
rect 32616 8271 32688 8319
rect 32616 8225 32629 8271
rect 32675 8225 32688 8271
rect 32616 8177 32688 8225
rect 32616 8131 32629 8177
rect 32675 8131 32688 8177
rect 32616 8083 32688 8131
rect 32616 8037 32629 8083
rect 32675 8037 32688 8083
rect 32616 7989 32688 8037
rect 32616 7943 32629 7989
rect 32675 7943 32688 7989
rect 32616 7895 32688 7943
rect 36752 8507 36765 8553
rect 36811 8507 36824 8553
rect 40888 8929 40960 8977
rect 40888 8883 40901 8929
rect 40947 8883 40960 8929
rect 40888 8835 40960 8883
rect 40888 8789 40901 8835
rect 40947 8789 40960 8835
rect 40888 8741 40960 8789
rect 40888 8695 40901 8741
rect 40947 8695 40960 8741
rect 40888 8647 40960 8695
rect 40888 8601 40901 8647
rect 40947 8601 40960 8647
rect 40888 8553 40960 8601
rect 36752 8459 36824 8507
rect 36752 8413 36765 8459
rect 36811 8413 36824 8459
rect 36752 8365 36824 8413
rect 36752 8319 36765 8365
rect 36811 8319 36824 8365
rect 36752 8271 36824 8319
rect 36752 8225 36765 8271
rect 36811 8225 36824 8271
rect 36752 8177 36824 8225
rect 36752 8131 36765 8177
rect 36811 8131 36824 8177
rect 36752 8083 36824 8131
rect 36752 8037 36765 8083
rect 36811 8037 36824 8083
rect 36752 7989 36824 8037
rect 36752 7943 36765 7989
rect 36811 7943 36824 7989
rect 32616 7849 32629 7895
rect 32675 7849 32688 7895
rect 36752 7895 36824 7943
rect 40888 8507 40901 8553
rect 40947 8507 40960 8553
rect 40888 8459 40960 8507
rect 40888 8413 40901 8459
rect 40947 8413 40960 8459
rect 40888 8365 40960 8413
rect 40888 8319 40901 8365
rect 40947 8319 40960 8365
rect 40888 8271 40960 8319
rect 40888 8225 40901 8271
rect 40947 8225 40960 8271
rect 40888 8177 40960 8225
rect 40888 8131 40901 8177
rect 40947 8131 40960 8177
rect 40888 8083 40960 8131
rect 40888 8037 40901 8083
rect 40947 8037 40960 8083
rect 40888 7989 40960 8037
rect 40888 7943 40901 7989
rect 40947 7943 40960 7989
rect 32616 7801 32688 7849
rect 32616 7755 32629 7801
rect 32675 7755 32688 7801
rect 32616 7707 32688 7755
rect 32616 7661 32629 7707
rect 32675 7661 32688 7707
rect 32616 7613 32688 7661
rect 32616 7567 32629 7613
rect 32675 7567 32688 7613
rect 32616 7519 32688 7567
rect 32616 7473 32629 7519
rect 32675 7473 32688 7519
rect 32616 7438 32688 7473
rect 36752 7849 36765 7895
rect 36811 7849 36824 7895
rect 40888 7895 40960 7943
rect 36752 7801 36824 7849
rect 36752 7755 36765 7801
rect 36811 7755 36824 7801
rect 36752 7707 36824 7755
rect 36752 7661 36765 7707
rect 36811 7661 36824 7707
rect 36752 7613 36824 7661
rect 36752 7567 36765 7613
rect 36811 7567 36824 7613
rect 36752 7519 36824 7567
rect 36752 7473 36765 7519
rect 36811 7473 36824 7519
rect 36752 7438 36824 7473
rect 40888 7849 40901 7895
rect 40947 7849 40960 7895
rect 40888 7801 40960 7849
rect 40888 7755 40901 7801
rect 40947 7755 40960 7801
rect 40888 7707 40960 7755
rect 40888 7661 40901 7707
rect 40947 7661 40960 7707
rect 40888 7613 40960 7661
rect 40888 7567 40901 7613
rect 40947 7567 40960 7613
rect 40888 7519 40960 7567
rect 40888 7473 40901 7519
rect 40947 7473 40960 7519
rect 40888 7438 40960 7473
rect 32616 7425 40960 7438
rect 32616 7379 32629 7425
rect 32675 7379 32723 7425
rect 32769 7379 32817 7425
rect 32863 7379 32911 7425
rect 32957 7379 33005 7425
rect 33051 7379 33099 7425
rect 33145 7379 33193 7425
rect 33239 7379 33287 7425
rect 33333 7379 33381 7425
rect 33427 7379 33475 7425
rect 33521 7379 33569 7425
rect 33615 7379 33663 7425
rect 33709 7379 33757 7425
rect 33803 7379 33851 7425
rect 33897 7379 33945 7425
rect 33991 7379 34039 7425
rect 34085 7379 34133 7425
rect 34179 7379 34227 7425
rect 34273 7379 34321 7425
rect 34367 7379 34415 7425
rect 34461 7379 34509 7425
rect 34555 7379 34603 7425
rect 34649 7379 34697 7425
rect 34743 7379 34791 7425
rect 34837 7379 34885 7425
rect 34931 7379 34979 7425
rect 35025 7379 35073 7425
rect 35119 7379 35167 7425
rect 35213 7379 35261 7425
rect 35307 7379 35355 7425
rect 35401 7379 35449 7425
rect 35495 7379 35543 7425
rect 35589 7379 35637 7425
rect 35683 7379 35731 7425
rect 35777 7379 35825 7425
rect 35871 7379 35919 7425
rect 35965 7379 36013 7425
rect 36059 7379 36107 7425
rect 36153 7379 36201 7425
rect 36247 7379 36295 7425
rect 36341 7379 36389 7425
rect 36435 7379 36483 7425
rect 36529 7379 36577 7425
rect 36623 7379 36671 7425
rect 36717 7379 36765 7425
rect 36811 7379 36859 7425
rect 36905 7379 36953 7425
rect 36999 7379 37047 7425
rect 37093 7379 37141 7425
rect 37187 7379 37235 7425
rect 37281 7379 37329 7425
rect 37375 7379 37423 7425
rect 37469 7379 37517 7425
rect 37563 7379 37611 7425
rect 37657 7379 37705 7425
rect 37751 7379 37799 7425
rect 37845 7379 37893 7425
rect 37939 7379 37987 7425
rect 38033 7379 38081 7425
rect 38127 7379 38175 7425
rect 38221 7379 38269 7425
rect 38315 7379 38363 7425
rect 38409 7379 38457 7425
rect 38503 7379 38551 7425
rect 38597 7379 38645 7425
rect 38691 7379 38739 7425
rect 38785 7379 38833 7425
rect 38879 7379 38927 7425
rect 38973 7379 39021 7425
rect 39067 7379 39115 7425
rect 39161 7379 39209 7425
rect 39255 7379 39303 7425
rect 39349 7379 39397 7425
rect 39443 7379 39491 7425
rect 39537 7379 39585 7425
rect 39631 7379 39679 7425
rect 39725 7379 39773 7425
rect 39819 7379 39867 7425
rect 39913 7379 39961 7425
rect 40007 7379 40055 7425
rect 40101 7379 40149 7425
rect 40195 7379 40243 7425
rect 40289 7379 40337 7425
rect 40383 7379 40431 7425
rect 40477 7379 40525 7425
rect 40571 7379 40619 7425
rect 40665 7379 40713 7425
rect 40759 7379 40807 7425
rect 40853 7379 40901 7425
rect 40947 7379 40960 7425
rect 32616 7366 40960 7379
rect 42312 12219 50656 12232
rect 42312 12173 42325 12219
rect 42371 12173 42419 12219
rect 42465 12173 42513 12219
rect 42559 12173 42607 12219
rect 42653 12173 42701 12219
rect 42747 12173 42795 12219
rect 42841 12173 42889 12219
rect 42935 12173 42983 12219
rect 43029 12173 43077 12219
rect 43123 12173 43171 12219
rect 43217 12173 43265 12219
rect 43311 12173 43359 12219
rect 43405 12173 43453 12219
rect 43499 12173 43547 12219
rect 43593 12173 43641 12219
rect 43687 12173 43735 12219
rect 43781 12173 43829 12219
rect 43875 12173 43923 12219
rect 43969 12173 44017 12219
rect 44063 12173 44111 12219
rect 44157 12173 44205 12219
rect 44251 12173 44299 12219
rect 44345 12173 44393 12219
rect 44439 12173 44487 12219
rect 44533 12173 44581 12219
rect 44627 12173 44675 12219
rect 44721 12173 44769 12219
rect 44815 12173 44863 12219
rect 44909 12173 44957 12219
rect 45003 12173 45051 12219
rect 45097 12173 45145 12219
rect 45191 12173 45239 12219
rect 45285 12173 45333 12219
rect 45379 12173 45427 12219
rect 45473 12173 45521 12219
rect 45567 12173 45615 12219
rect 45661 12173 45709 12219
rect 45755 12173 45803 12219
rect 45849 12173 45897 12219
rect 45943 12173 45991 12219
rect 46037 12173 46085 12219
rect 46131 12173 46179 12219
rect 46225 12173 46273 12219
rect 46319 12173 46367 12219
rect 46413 12173 46461 12219
rect 46507 12173 46555 12219
rect 46601 12173 46649 12219
rect 46695 12173 46743 12219
rect 46789 12173 46837 12219
rect 46883 12173 46931 12219
rect 46977 12173 47025 12219
rect 47071 12173 47119 12219
rect 47165 12173 47213 12219
rect 47259 12173 47307 12219
rect 47353 12173 47401 12219
rect 47447 12173 47495 12219
rect 47541 12173 47589 12219
rect 47635 12173 47683 12219
rect 47729 12173 47777 12219
rect 47823 12173 47871 12219
rect 47917 12173 47965 12219
rect 48011 12173 48059 12219
rect 48105 12173 48153 12219
rect 48199 12173 48247 12219
rect 48293 12173 48341 12219
rect 48387 12173 48435 12219
rect 48481 12173 48529 12219
rect 48575 12173 48623 12219
rect 48669 12173 48717 12219
rect 48763 12173 48811 12219
rect 48857 12173 48905 12219
rect 48951 12173 48999 12219
rect 49045 12173 49093 12219
rect 49139 12173 49187 12219
rect 49233 12173 49281 12219
rect 49327 12173 49375 12219
rect 49421 12173 49469 12219
rect 49515 12173 49563 12219
rect 49609 12173 49657 12219
rect 49703 12173 49751 12219
rect 49797 12173 49845 12219
rect 49891 12173 49939 12219
rect 49985 12173 50033 12219
rect 50079 12173 50127 12219
rect 50173 12173 50221 12219
rect 50267 12173 50315 12219
rect 50361 12173 50409 12219
rect 50455 12173 50503 12219
rect 50549 12173 50597 12219
rect 50643 12173 50656 12219
rect 42312 12160 50656 12173
rect 42312 12125 42384 12160
rect 42312 12079 42325 12125
rect 42371 12079 42384 12125
rect 42312 12031 42384 12079
rect 42312 11985 42325 12031
rect 42371 11985 42384 12031
rect 42312 11937 42384 11985
rect 42312 11891 42325 11937
rect 42371 11891 42384 11937
rect 42312 11843 42384 11891
rect 42312 11797 42325 11843
rect 42371 11797 42384 11843
rect 46448 12125 46520 12160
rect 46448 12079 46461 12125
rect 46507 12079 46520 12125
rect 46448 12031 46520 12079
rect 46448 11985 46461 12031
rect 46507 11985 46520 12031
rect 46448 11937 46520 11985
rect 46448 11891 46461 11937
rect 46507 11891 46520 11937
rect 46448 11843 46520 11891
rect 42312 11749 42384 11797
rect 46448 11797 46461 11843
rect 46507 11797 46520 11843
rect 50584 12125 50656 12160
rect 50584 12079 50597 12125
rect 50643 12079 50656 12125
rect 50584 12031 50656 12079
rect 50584 11985 50597 12031
rect 50643 11985 50656 12031
rect 50584 11937 50656 11985
rect 50584 11891 50597 11937
rect 50643 11891 50656 11937
rect 50584 11843 50656 11891
rect 42312 11703 42325 11749
rect 42371 11703 42384 11749
rect 42312 11655 42384 11703
rect 46448 11749 46520 11797
rect 50584 11797 50597 11843
rect 50643 11797 50656 11843
rect 46448 11703 46461 11749
rect 46507 11703 46520 11749
rect 42312 11609 42325 11655
rect 42371 11609 42384 11655
rect 42312 11561 42384 11609
rect 42312 11515 42325 11561
rect 42371 11515 42384 11561
rect 42312 11467 42384 11515
rect 42312 11421 42325 11467
rect 42371 11421 42384 11467
rect 42312 11373 42384 11421
rect 42312 11327 42325 11373
rect 42371 11327 42384 11373
rect 42312 11279 42384 11327
rect 42312 11233 42325 11279
rect 42371 11233 42384 11279
rect 42312 11185 42384 11233
rect 42312 11139 42325 11185
rect 42371 11139 42384 11185
rect 42312 11091 42384 11139
rect 42312 11045 42325 11091
rect 42371 11045 42384 11091
rect 46448 11655 46520 11703
rect 50584 11749 50656 11797
rect 50584 11703 50597 11749
rect 50643 11703 50656 11749
rect 46448 11609 46461 11655
rect 46507 11609 46520 11655
rect 46448 11561 46520 11609
rect 46448 11515 46461 11561
rect 46507 11515 46520 11561
rect 46448 11467 46520 11515
rect 46448 11421 46461 11467
rect 46507 11421 46520 11467
rect 46448 11373 46520 11421
rect 46448 11327 46461 11373
rect 46507 11327 46520 11373
rect 46448 11279 46520 11327
rect 46448 11233 46461 11279
rect 46507 11233 46520 11279
rect 46448 11185 46520 11233
rect 46448 11139 46461 11185
rect 46507 11139 46520 11185
rect 46448 11091 46520 11139
rect 42312 10997 42384 11045
rect 42312 10951 42325 10997
rect 42371 10951 42384 10997
rect 42312 10903 42384 10951
rect 42312 10857 42325 10903
rect 42371 10857 42384 10903
rect 42312 10809 42384 10857
rect 42312 10763 42325 10809
rect 42371 10763 42384 10809
rect 42312 10715 42384 10763
rect 42312 10669 42325 10715
rect 42371 10669 42384 10715
rect 42312 10621 42384 10669
rect 46448 11045 46461 11091
rect 46507 11045 46520 11091
rect 50584 11655 50656 11703
rect 50584 11609 50597 11655
rect 50643 11609 50656 11655
rect 50584 11561 50656 11609
rect 50584 11515 50597 11561
rect 50643 11515 50656 11561
rect 50584 11467 50656 11515
rect 50584 11421 50597 11467
rect 50643 11421 50656 11467
rect 50584 11373 50656 11421
rect 50584 11327 50597 11373
rect 50643 11327 50656 11373
rect 50584 11279 50656 11327
rect 50584 11233 50597 11279
rect 50643 11233 50656 11279
rect 50584 11185 50656 11233
rect 50584 11139 50597 11185
rect 50643 11139 50656 11185
rect 50584 11091 50656 11139
rect 46448 10997 46520 11045
rect 46448 10951 46461 10997
rect 46507 10951 46520 10997
rect 46448 10903 46520 10951
rect 46448 10857 46461 10903
rect 46507 10857 46520 10903
rect 46448 10809 46520 10857
rect 46448 10763 46461 10809
rect 46507 10763 46520 10809
rect 46448 10715 46520 10763
rect 46448 10669 46461 10715
rect 46507 10669 46520 10715
rect 42312 10575 42325 10621
rect 42371 10575 42384 10621
rect 42312 10527 42384 10575
rect 42312 10481 42325 10527
rect 42371 10481 42384 10527
rect 42312 10433 42384 10481
rect 42312 10387 42325 10433
rect 42371 10387 42384 10433
rect 42312 10339 42384 10387
rect 42312 10293 42325 10339
rect 42371 10293 42384 10339
rect 42312 10245 42384 10293
rect 42312 10199 42325 10245
rect 42371 10199 42384 10245
rect 42312 10151 42384 10199
rect 42312 10105 42325 10151
rect 42371 10105 42384 10151
rect 42312 10057 42384 10105
rect 42312 10011 42325 10057
rect 42371 10011 42384 10057
rect 46448 10621 46520 10669
rect 50584 11045 50597 11091
rect 50643 11045 50656 11091
rect 50584 10997 50656 11045
rect 50584 10951 50597 10997
rect 50643 10951 50656 10997
rect 50584 10903 50656 10951
rect 50584 10857 50597 10903
rect 50643 10857 50656 10903
rect 50584 10809 50656 10857
rect 50584 10763 50597 10809
rect 50643 10763 50656 10809
rect 50584 10715 50656 10763
rect 50584 10669 50597 10715
rect 50643 10669 50656 10715
rect 46448 10575 46461 10621
rect 46507 10575 46520 10621
rect 46448 10527 46520 10575
rect 46448 10481 46461 10527
rect 46507 10481 46520 10527
rect 46448 10433 46520 10481
rect 46448 10387 46461 10433
rect 46507 10387 46520 10433
rect 46448 10339 46520 10387
rect 46448 10293 46461 10339
rect 46507 10293 46520 10339
rect 46448 10245 46520 10293
rect 46448 10199 46461 10245
rect 46507 10199 46520 10245
rect 46448 10151 46520 10199
rect 46448 10105 46461 10151
rect 46507 10105 46520 10151
rect 46448 10057 46520 10105
rect 42312 9963 42384 10011
rect 42312 9917 42325 9963
rect 42371 9917 42384 9963
rect 42312 9869 42384 9917
rect 42312 9823 42325 9869
rect 42371 9823 42384 9869
rect 42312 9775 42384 9823
rect 42312 9729 42325 9775
rect 42371 9729 42384 9775
rect 42312 9681 42384 9729
rect 42312 9635 42325 9681
rect 42371 9635 42384 9681
rect 42312 9587 42384 9635
rect 42312 9541 42325 9587
rect 42371 9541 42384 9587
rect 46448 10011 46461 10057
rect 46507 10011 46520 10057
rect 50584 10621 50656 10669
rect 50584 10575 50597 10621
rect 50643 10575 50656 10621
rect 50584 10527 50656 10575
rect 50584 10481 50597 10527
rect 50643 10481 50656 10527
rect 50584 10433 50656 10481
rect 50584 10387 50597 10433
rect 50643 10387 50656 10433
rect 50584 10339 50656 10387
rect 50584 10293 50597 10339
rect 50643 10293 50656 10339
rect 50584 10245 50656 10293
rect 50584 10199 50597 10245
rect 50643 10199 50656 10245
rect 50584 10151 50656 10199
rect 50584 10105 50597 10151
rect 50643 10105 50656 10151
rect 50584 10057 50656 10105
rect 46448 9963 46520 10011
rect 46448 9917 46461 9963
rect 46507 9917 46520 9963
rect 46448 9869 46520 9917
rect 46448 9823 46461 9869
rect 46507 9823 46520 9869
rect 46448 9775 46520 9823
rect 46448 9729 46461 9775
rect 46507 9729 46520 9775
rect 46448 9681 46520 9729
rect 46448 9635 46461 9681
rect 46507 9635 46520 9681
rect 46448 9587 46520 9635
rect 42312 9493 42384 9541
rect 42312 9447 42325 9493
rect 42371 9447 42384 9493
rect 42312 9399 42384 9447
rect 42312 9353 42325 9399
rect 42371 9353 42384 9399
rect 42312 9305 42384 9353
rect 42312 9259 42325 9305
rect 42371 9259 42384 9305
rect 42312 9211 42384 9259
rect 42312 9165 42325 9211
rect 42371 9165 42384 9211
rect 42312 9117 42384 9165
rect 42312 9071 42325 9117
rect 42371 9071 42384 9117
rect 42312 9023 42384 9071
rect 42312 8977 42325 9023
rect 42371 8977 42384 9023
rect 42312 8929 42384 8977
rect 46448 9541 46461 9587
rect 46507 9541 46520 9587
rect 50584 10011 50597 10057
rect 50643 10011 50656 10057
rect 50584 9963 50656 10011
rect 50584 9917 50597 9963
rect 50643 9917 50656 9963
rect 50584 9869 50656 9917
rect 50584 9823 50597 9869
rect 50643 9823 50656 9869
rect 50584 9775 50656 9823
rect 50584 9729 50597 9775
rect 50643 9729 50656 9775
rect 50584 9681 50656 9729
rect 50584 9635 50597 9681
rect 50643 9635 50656 9681
rect 50584 9587 50656 9635
rect 46448 9493 46520 9541
rect 46448 9447 46461 9493
rect 46507 9447 46520 9493
rect 46448 9399 46520 9447
rect 46448 9353 46461 9399
rect 46507 9353 46520 9399
rect 46448 9305 46520 9353
rect 46448 9259 46461 9305
rect 46507 9259 46520 9305
rect 46448 9211 46520 9259
rect 46448 9165 46461 9211
rect 46507 9165 46520 9211
rect 46448 9117 46520 9165
rect 46448 9071 46461 9117
rect 46507 9071 46520 9117
rect 46448 9023 46520 9071
rect 46448 8977 46461 9023
rect 46507 8977 46520 9023
rect 42312 8883 42325 8929
rect 42371 8883 42384 8929
rect 42312 8835 42384 8883
rect 42312 8789 42325 8835
rect 42371 8789 42384 8835
rect 42312 8741 42384 8789
rect 42312 8695 42325 8741
rect 42371 8695 42384 8741
rect 42312 8647 42384 8695
rect 42312 8601 42325 8647
rect 42371 8601 42384 8647
rect 42312 8553 42384 8601
rect 42312 8507 42325 8553
rect 42371 8507 42384 8553
rect 46448 8929 46520 8977
rect 50584 9541 50597 9587
rect 50643 9541 50656 9587
rect 50584 9493 50656 9541
rect 50584 9447 50597 9493
rect 50643 9447 50656 9493
rect 50584 9399 50656 9447
rect 50584 9353 50597 9399
rect 50643 9353 50656 9399
rect 50584 9305 50656 9353
rect 50584 9259 50597 9305
rect 50643 9259 50656 9305
rect 50584 9211 50656 9259
rect 50584 9165 50597 9211
rect 50643 9165 50656 9211
rect 50584 9117 50656 9165
rect 50584 9071 50597 9117
rect 50643 9071 50656 9117
rect 50584 9023 50656 9071
rect 50584 8977 50597 9023
rect 50643 8977 50656 9023
rect 46448 8883 46461 8929
rect 46507 8883 46520 8929
rect 46448 8835 46520 8883
rect 46448 8789 46461 8835
rect 46507 8789 46520 8835
rect 46448 8741 46520 8789
rect 46448 8695 46461 8741
rect 46507 8695 46520 8741
rect 46448 8647 46520 8695
rect 46448 8601 46461 8647
rect 46507 8601 46520 8647
rect 46448 8553 46520 8601
rect 42312 8459 42384 8507
rect 42312 8413 42325 8459
rect 42371 8413 42384 8459
rect 42312 8365 42384 8413
rect 42312 8319 42325 8365
rect 42371 8319 42384 8365
rect 42312 8271 42384 8319
rect 42312 8225 42325 8271
rect 42371 8225 42384 8271
rect 42312 8177 42384 8225
rect 42312 8131 42325 8177
rect 42371 8131 42384 8177
rect 42312 8083 42384 8131
rect 42312 8037 42325 8083
rect 42371 8037 42384 8083
rect 42312 7989 42384 8037
rect 42312 7943 42325 7989
rect 42371 7943 42384 7989
rect 42312 7895 42384 7943
rect 46448 8507 46461 8553
rect 46507 8507 46520 8553
rect 50584 8929 50656 8977
rect 50584 8883 50597 8929
rect 50643 8883 50656 8929
rect 50584 8835 50656 8883
rect 50584 8789 50597 8835
rect 50643 8789 50656 8835
rect 50584 8741 50656 8789
rect 50584 8695 50597 8741
rect 50643 8695 50656 8741
rect 50584 8647 50656 8695
rect 50584 8601 50597 8647
rect 50643 8601 50656 8647
rect 50584 8553 50656 8601
rect 46448 8459 46520 8507
rect 46448 8413 46461 8459
rect 46507 8413 46520 8459
rect 46448 8365 46520 8413
rect 46448 8319 46461 8365
rect 46507 8319 46520 8365
rect 46448 8271 46520 8319
rect 46448 8225 46461 8271
rect 46507 8225 46520 8271
rect 46448 8177 46520 8225
rect 46448 8131 46461 8177
rect 46507 8131 46520 8177
rect 46448 8083 46520 8131
rect 46448 8037 46461 8083
rect 46507 8037 46520 8083
rect 46448 7989 46520 8037
rect 46448 7943 46461 7989
rect 46507 7943 46520 7989
rect 42312 7849 42325 7895
rect 42371 7849 42384 7895
rect 46448 7895 46520 7943
rect 50584 8507 50597 8553
rect 50643 8507 50656 8553
rect 50584 8459 50656 8507
rect 50584 8413 50597 8459
rect 50643 8413 50656 8459
rect 50584 8365 50656 8413
rect 50584 8319 50597 8365
rect 50643 8319 50656 8365
rect 50584 8271 50656 8319
rect 50584 8225 50597 8271
rect 50643 8225 50656 8271
rect 50584 8177 50656 8225
rect 50584 8131 50597 8177
rect 50643 8131 50656 8177
rect 50584 8083 50656 8131
rect 50584 8037 50597 8083
rect 50643 8037 50656 8083
rect 50584 7989 50656 8037
rect 50584 7943 50597 7989
rect 50643 7943 50656 7989
rect 42312 7801 42384 7849
rect 42312 7755 42325 7801
rect 42371 7755 42384 7801
rect 42312 7707 42384 7755
rect 42312 7661 42325 7707
rect 42371 7661 42384 7707
rect 42312 7613 42384 7661
rect 42312 7567 42325 7613
rect 42371 7567 42384 7613
rect 42312 7519 42384 7567
rect 42312 7473 42325 7519
rect 42371 7473 42384 7519
rect 42312 7438 42384 7473
rect 46448 7849 46461 7895
rect 46507 7849 46520 7895
rect 50584 7895 50656 7943
rect 46448 7801 46520 7849
rect 46448 7755 46461 7801
rect 46507 7755 46520 7801
rect 46448 7707 46520 7755
rect 46448 7661 46461 7707
rect 46507 7661 46520 7707
rect 46448 7613 46520 7661
rect 46448 7567 46461 7613
rect 46507 7567 46520 7613
rect 46448 7519 46520 7567
rect 46448 7473 46461 7519
rect 46507 7473 46520 7519
rect 46448 7438 46520 7473
rect 50584 7849 50597 7895
rect 50643 7849 50656 7895
rect 50584 7801 50656 7849
rect 50584 7755 50597 7801
rect 50643 7755 50656 7801
rect 50584 7707 50656 7755
rect 50584 7661 50597 7707
rect 50643 7661 50656 7707
rect 50584 7613 50656 7661
rect 50584 7567 50597 7613
rect 50643 7567 50656 7613
rect 50584 7519 50656 7567
rect 50584 7473 50597 7519
rect 50643 7473 50656 7519
rect 50584 7438 50656 7473
rect 42312 7425 50656 7438
rect 42312 7379 42325 7425
rect 42371 7379 42419 7425
rect 42465 7379 42513 7425
rect 42559 7379 42607 7425
rect 42653 7379 42701 7425
rect 42747 7379 42795 7425
rect 42841 7379 42889 7425
rect 42935 7379 42983 7425
rect 43029 7379 43077 7425
rect 43123 7379 43171 7425
rect 43217 7379 43265 7425
rect 43311 7379 43359 7425
rect 43405 7379 43453 7425
rect 43499 7379 43547 7425
rect 43593 7379 43641 7425
rect 43687 7379 43735 7425
rect 43781 7379 43829 7425
rect 43875 7379 43923 7425
rect 43969 7379 44017 7425
rect 44063 7379 44111 7425
rect 44157 7379 44205 7425
rect 44251 7379 44299 7425
rect 44345 7379 44393 7425
rect 44439 7379 44487 7425
rect 44533 7379 44581 7425
rect 44627 7379 44675 7425
rect 44721 7379 44769 7425
rect 44815 7379 44863 7425
rect 44909 7379 44957 7425
rect 45003 7379 45051 7425
rect 45097 7379 45145 7425
rect 45191 7379 45239 7425
rect 45285 7379 45333 7425
rect 45379 7379 45427 7425
rect 45473 7379 45521 7425
rect 45567 7379 45615 7425
rect 45661 7379 45709 7425
rect 45755 7379 45803 7425
rect 45849 7379 45897 7425
rect 45943 7379 45991 7425
rect 46037 7379 46085 7425
rect 46131 7379 46179 7425
rect 46225 7379 46273 7425
rect 46319 7379 46367 7425
rect 46413 7379 46461 7425
rect 46507 7379 46555 7425
rect 46601 7379 46649 7425
rect 46695 7379 46743 7425
rect 46789 7379 46837 7425
rect 46883 7379 46931 7425
rect 46977 7379 47025 7425
rect 47071 7379 47119 7425
rect 47165 7379 47213 7425
rect 47259 7379 47307 7425
rect 47353 7379 47401 7425
rect 47447 7379 47495 7425
rect 47541 7379 47589 7425
rect 47635 7379 47683 7425
rect 47729 7379 47777 7425
rect 47823 7379 47871 7425
rect 47917 7379 47965 7425
rect 48011 7379 48059 7425
rect 48105 7379 48153 7425
rect 48199 7379 48247 7425
rect 48293 7379 48341 7425
rect 48387 7379 48435 7425
rect 48481 7379 48529 7425
rect 48575 7379 48623 7425
rect 48669 7379 48717 7425
rect 48763 7379 48811 7425
rect 48857 7379 48905 7425
rect 48951 7379 48999 7425
rect 49045 7379 49093 7425
rect 49139 7379 49187 7425
rect 49233 7379 49281 7425
rect 49327 7379 49375 7425
rect 49421 7379 49469 7425
rect 49515 7379 49563 7425
rect 49609 7379 49657 7425
rect 49703 7379 49751 7425
rect 49797 7379 49845 7425
rect 49891 7379 49939 7425
rect 49985 7379 50033 7425
rect 50079 7379 50127 7425
rect 50173 7379 50221 7425
rect 50267 7379 50315 7425
rect 50361 7379 50409 7425
rect 50455 7379 50503 7425
rect 50549 7379 50597 7425
rect 50643 7379 50656 7425
rect 42312 7366 50656 7379
rect 52008 12219 60352 12232
rect 52008 12173 52021 12219
rect 52067 12173 52115 12219
rect 52161 12173 52209 12219
rect 52255 12173 52303 12219
rect 52349 12173 52397 12219
rect 52443 12173 52491 12219
rect 52537 12173 52585 12219
rect 52631 12173 52679 12219
rect 52725 12173 52773 12219
rect 52819 12173 52867 12219
rect 52913 12173 52961 12219
rect 53007 12173 53055 12219
rect 53101 12173 53149 12219
rect 53195 12173 53243 12219
rect 53289 12173 53337 12219
rect 53383 12173 53431 12219
rect 53477 12173 53525 12219
rect 53571 12173 53619 12219
rect 53665 12173 53713 12219
rect 53759 12173 53807 12219
rect 53853 12173 53901 12219
rect 53947 12173 53995 12219
rect 54041 12173 54089 12219
rect 54135 12173 54183 12219
rect 54229 12173 54277 12219
rect 54323 12173 54371 12219
rect 54417 12173 54465 12219
rect 54511 12173 54559 12219
rect 54605 12173 54653 12219
rect 54699 12173 54747 12219
rect 54793 12173 54841 12219
rect 54887 12173 54935 12219
rect 54981 12173 55029 12219
rect 55075 12173 55123 12219
rect 55169 12173 55217 12219
rect 55263 12173 55311 12219
rect 55357 12173 55405 12219
rect 55451 12173 55499 12219
rect 55545 12173 55593 12219
rect 55639 12173 55687 12219
rect 55733 12173 55781 12219
rect 55827 12173 55875 12219
rect 55921 12173 55969 12219
rect 56015 12173 56063 12219
rect 56109 12173 56157 12219
rect 56203 12173 56251 12219
rect 56297 12173 56345 12219
rect 56391 12173 56439 12219
rect 56485 12173 56533 12219
rect 56579 12173 56627 12219
rect 56673 12173 56721 12219
rect 56767 12173 56815 12219
rect 56861 12173 56909 12219
rect 56955 12173 57003 12219
rect 57049 12173 57097 12219
rect 57143 12173 57191 12219
rect 57237 12173 57285 12219
rect 57331 12173 57379 12219
rect 57425 12173 57473 12219
rect 57519 12173 57567 12219
rect 57613 12173 57661 12219
rect 57707 12173 57755 12219
rect 57801 12173 57849 12219
rect 57895 12173 57943 12219
rect 57989 12173 58037 12219
rect 58083 12173 58131 12219
rect 58177 12173 58225 12219
rect 58271 12173 58319 12219
rect 58365 12173 58413 12219
rect 58459 12173 58507 12219
rect 58553 12173 58601 12219
rect 58647 12173 58695 12219
rect 58741 12173 58789 12219
rect 58835 12173 58883 12219
rect 58929 12173 58977 12219
rect 59023 12173 59071 12219
rect 59117 12173 59165 12219
rect 59211 12173 59259 12219
rect 59305 12173 59353 12219
rect 59399 12173 59447 12219
rect 59493 12173 59541 12219
rect 59587 12173 59635 12219
rect 59681 12173 59729 12219
rect 59775 12173 59823 12219
rect 59869 12173 59917 12219
rect 59963 12173 60011 12219
rect 60057 12173 60105 12219
rect 60151 12173 60199 12219
rect 60245 12173 60293 12219
rect 60339 12173 60352 12219
rect 52008 12160 60352 12173
rect 52008 12125 52080 12160
rect 52008 12079 52021 12125
rect 52067 12079 52080 12125
rect 52008 12031 52080 12079
rect 52008 11985 52021 12031
rect 52067 11985 52080 12031
rect 52008 11937 52080 11985
rect 52008 11891 52021 11937
rect 52067 11891 52080 11937
rect 52008 11843 52080 11891
rect 52008 11797 52021 11843
rect 52067 11797 52080 11843
rect 56144 12125 56216 12160
rect 56144 12079 56157 12125
rect 56203 12079 56216 12125
rect 56144 12031 56216 12079
rect 56144 11985 56157 12031
rect 56203 11985 56216 12031
rect 56144 11937 56216 11985
rect 56144 11891 56157 11937
rect 56203 11891 56216 11937
rect 56144 11843 56216 11891
rect 52008 11749 52080 11797
rect 56144 11797 56157 11843
rect 56203 11797 56216 11843
rect 60280 12125 60352 12160
rect 60280 12079 60293 12125
rect 60339 12079 60352 12125
rect 60280 12031 60352 12079
rect 60280 11985 60293 12031
rect 60339 11985 60352 12031
rect 60280 11937 60352 11985
rect 60280 11891 60293 11937
rect 60339 11891 60352 11937
rect 60280 11843 60352 11891
rect 52008 11703 52021 11749
rect 52067 11703 52080 11749
rect 52008 11655 52080 11703
rect 56144 11749 56216 11797
rect 60280 11797 60293 11843
rect 60339 11797 60352 11843
rect 56144 11703 56157 11749
rect 56203 11703 56216 11749
rect 52008 11609 52021 11655
rect 52067 11609 52080 11655
rect 52008 11561 52080 11609
rect 52008 11515 52021 11561
rect 52067 11515 52080 11561
rect 52008 11467 52080 11515
rect 52008 11421 52021 11467
rect 52067 11421 52080 11467
rect 52008 11373 52080 11421
rect 52008 11327 52021 11373
rect 52067 11327 52080 11373
rect 52008 11279 52080 11327
rect 52008 11233 52021 11279
rect 52067 11233 52080 11279
rect 52008 11185 52080 11233
rect 52008 11139 52021 11185
rect 52067 11139 52080 11185
rect 52008 11091 52080 11139
rect 52008 11045 52021 11091
rect 52067 11045 52080 11091
rect 56144 11655 56216 11703
rect 60280 11749 60352 11797
rect 60280 11703 60293 11749
rect 60339 11703 60352 11749
rect 56144 11609 56157 11655
rect 56203 11609 56216 11655
rect 56144 11561 56216 11609
rect 56144 11515 56157 11561
rect 56203 11515 56216 11561
rect 56144 11467 56216 11515
rect 56144 11421 56157 11467
rect 56203 11421 56216 11467
rect 56144 11373 56216 11421
rect 56144 11327 56157 11373
rect 56203 11327 56216 11373
rect 56144 11279 56216 11327
rect 56144 11233 56157 11279
rect 56203 11233 56216 11279
rect 56144 11185 56216 11233
rect 56144 11139 56157 11185
rect 56203 11139 56216 11185
rect 56144 11091 56216 11139
rect 52008 10997 52080 11045
rect 52008 10951 52021 10997
rect 52067 10951 52080 10997
rect 52008 10903 52080 10951
rect 52008 10857 52021 10903
rect 52067 10857 52080 10903
rect 52008 10809 52080 10857
rect 52008 10763 52021 10809
rect 52067 10763 52080 10809
rect 52008 10715 52080 10763
rect 52008 10669 52021 10715
rect 52067 10669 52080 10715
rect 52008 10621 52080 10669
rect 56144 11045 56157 11091
rect 56203 11045 56216 11091
rect 60280 11655 60352 11703
rect 60280 11609 60293 11655
rect 60339 11609 60352 11655
rect 60280 11561 60352 11609
rect 60280 11515 60293 11561
rect 60339 11515 60352 11561
rect 60280 11467 60352 11515
rect 60280 11421 60293 11467
rect 60339 11421 60352 11467
rect 60280 11373 60352 11421
rect 60280 11327 60293 11373
rect 60339 11327 60352 11373
rect 60280 11279 60352 11327
rect 60280 11233 60293 11279
rect 60339 11233 60352 11279
rect 60280 11185 60352 11233
rect 60280 11139 60293 11185
rect 60339 11139 60352 11185
rect 60280 11091 60352 11139
rect 56144 10997 56216 11045
rect 56144 10951 56157 10997
rect 56203 10951 56216 10997
rect 56144 10903 56216 10951
rect 56144 10857 56157 10903
rect 56203 10857 56216 10903
rect 56144 10809 56216 10857
rect 56144 10763 56157 10809
rect 56203 10763 56216 10809
rect 56144 10715 56216 10763
rect 56144 10669 56157 10715
rect 56203 10669 56216 10715
rect 52008 10575 52021 10621
rect 52067 10575 52080 10621
rect 52008 10527 52080 10575
rect 52008 10481 52021 10527
rect 52067 10481 52080 10527
rect 52008 10433 52080 10481
rect 52008 10387 52021 10433
rect 52067 10387 52080 10433
rect 52008 10339 52080 10387
rect 52008 10293 52021 10339
rect 52067 10293 52080 10339
rect 52008 10245 52080 10293
rect 52008 10199 52021 10245
rect 52067 10199 52080 10245
rect 52008 10151 52080 10199
rect 52008 10105 52021 10151
rect 52067 10105 52080 10151
rect 52008 10057 52080 10105
rect 52008 10011 52021 10057
rect 52067 10011 52080 10057
rect 56144 10621 56216 10669
rect 60280 11045 60293 11091
rect 60339 11045 60352 11091
rect 60280 10997 60352 11045
rect 60280 10951 60293 10997
rect 60339 10951 60352 10997
rect 60280 10903 60352 10951
rect 60280 10857 60293 10903
rect 60339 10857 60352 10903
rect 60280 10809 60352 10857
rect 60280 10763 60293 10809
rect 60339 10763 60352 10809
rect 60280 10715 60352 10763
rect 60280 10669 60293 10715
rect 60339 10669 60352 10715
rect 56144 10575 56157 10621
rect 56203 10575 56216 10621
rect 56144 10527 56216 10575
rect 56144 10481 56157 10527
rect 56203 10481 56216 10527
rect 56144 10433 56216 10481
rect 56144 10387 56157 10433
rect 56203 10387 56216 10433
rect 56144 10339 56216 10387
rect 56144 10293 56157 10339
rect 56203 10293 56216 10339
rect 56144 10245 56216 10293
rect 56144 10199 56157 10245
rect 56203 10199 56216 10245
rect 56144 10151 56216 10199
rect 56144 10105 56157 10151
rect 56203 10105 56216 10151
rect 56144 10057 56216 10105
rect 52008 9963 52080 10011
rect 52008 9917 52021 9963
rect 52067 9917 52080 9963
rect 52008 9869 52080 9917
rect 52008 9823 52021 9869
rect 52067 9823 52080 9869
rect 52008 9775 52080 9823
rect 52008 9729 52021 9775
rect 52067 9729 52080 9775
rect 52008 9681 52080 9729
rect 52008 9635 52021 9681
rect 52067 9635 52080 9681
rect 52008 9587 52080 9635
rect 52008 9541 52021 9587
rect 52067 9541 52080 9587
rect 56144 10011 56157 10057
rect 56203 10011 56216 10057
rect 60280 10621 60352 10669
rect 60280 10575 60293 10621
rect 60339 10575 60352 10621
rect 60280 10527 60352 10575
rect 60280 10481 60293 10527
rect 60339 10481 60352 10527
rect 60280 10433 60352 10481
rect 60280 10387 60293 10433
rect 60339 10387 60352 10433
rect 60280 10339 60352 10387
rect 60280 10293 60293 10339
rect 60339 10293 60352 10339
rect 60280 10245 60352 10293
rect 60280 10199 60293 10245
rect 60339 10199 60352 10245
rect 60280 10151 60352 10199
rect 60280 10105 60293 10151
rect 60339 10105 60352 10151
rect 60280 10057 60352 10105
rect 56144 9963 56216 10011
rect 56144 9917 56157 9963
rect 56203 9917 56216 9963
rect 56144 9869 56216 9917
rect 56144 9823 56157 9869
rect 56203 9823 56216 9869
rect 56144 9775 56216 9823
rect 56144 9729 56157 9775
rect 56203 9729 56216 9775
rect 56144 9681 56216 9729
rect 56144 9635 56157 9681
rect 56203 9635 56216 9681
rect 56144 9587 56216 9635
rect 52008 9493 52080 9541
rect 52008 9447 52021 9493
rect 52067 9447 52080 9493
rect 52008 9399 52080 9447
rect 52008 9353 52021 9399
rect 52067 9353 52080 9399
rect 52008 9305 52080 9353
rect 52008 9259 52021 9305
rect 52067 9259 52080 9305
rect 52008 9211 52080 9259
rect 52008 9165 52021 9211
rect 52067 9165 52080 9211
rect 52008 9117 52080 9165
rect 52008 9071 52021 9117
rect 52067 9071 52080 9117
rect 52008 9023 52080 9071
rect 52008 8977 52021 9023
rect 52067 8977 52080 9023
rect 52008 8929 52080 8977
rect 56144 9541 56157 9587
rect 56203 9541 56216 9587
rect 60280 10011 60293 10057
rect 60339 10011 60352 10057
rect 60280 9963 60352 10011
rect 60280 9917 60293 9963
rect 60339 9917 60352 9963
rect 60280 9869 60352 9917
rect 60280 9823 60293 9869
rect 60339 9823 60352 9869
rect 60280 9775 60352 9823
rect 60280 9729 60293 9775
rect 60339 9729 60352 9775
rect 60280 9681 60352 9729
rect 60280 9635 60293 9681
rect 60339 9635 60352 9681
rect 60280 9587 60352 9635
rect 56144 9493 56216 9541
rect 56144 9447 56157 9493
rect 56203 9447 56216 9493
rect 56144 9399 56216 9447
rect 56144 9353 56157 9399
rect 56203 9353 56216 9399
rect 56144 9305 56216 9353
rect 56144 9259 56157 9305
rect 56203 9259 56216 9305
rect 56144 9211 56216 9259
rect 56144 9165 56157 9211
rect 56203 9165 56216 9211
rect 56144 9117 56216 9165
rect 56144 9071 56157 9117
rect 56203 9071 56216 9117
rect 56144 9023 56216 9071
rect 56144 8977 56157 9023
rect 56203 8977 56216 9023
rect 52008 8883 52021 8929
rect 52067 8883 52080 8929
rect 52008 8835 52080 8883
rect 52008 8789 52021 8835
rect 52067 8789 52080 8835
rect 52008 8741 52080 8789
rect 52008 8695 52021 8741
rect 52067 8695 52080 8741
rect 52008 8647 52080 8695
rect 52008 8601 52021 8647
rect 52067 8601 52080 8647
rect 52008 8553 52080 8601
rect 52008 8507 52021 8553
rect 52067 8507 52080 8553
rect 56144 8929 56216 8977
rect 60280 9541 60293 9587
rect 60339 9541 60352 9587
rect 60280 9493 60352 9541
rect 60280 9447 60293 9493
rect 60339 9447 60352 9493
rect 60280 9399 60352 9447
rect 60280 9353 60293 9399
rect 60339 9353 60352 9399
rect 60280 9305 60352 9353
rect 60280 9259 60293 9305
rect 60339 9259 60352 9305
rect 60280 9211 60352 9259
rect 60280 9165 60293 9211
rect 60339 9165 60352 9211
rect 60280 9117 60352 9165
rect 60280 9071 60293 9117
rect 60339 9071 60352 9117
rect 60280 9023 60352 9071
rect 60280 8977 60293 9023
rect 60339 8977 60352 9023
rect 56144 8883 56157 8929
rect 56203 8883 56216 8929
rect 56144 8835 56216 8883
rect 56144 8789 56157 8835
rect 56203 8789 56216 8835
rect 56144 8741 56216 8789
rect 56144 8695 56157 8741
rect 56203 8695 56216 8741
rect 56144 8647 56216 8695
rect 56144 8601 56157 8647
rect 56203 8601 56216 8647
rect 56144 8553 56216 8601
rect 52008 8459 52080 8507
rect 52008 8413 52021 8459
rect 52067 8413 52080 8459
rect 52008 8365 52080 8413
rect 52008 8319 52021 8365
rect 52067 8319 52080 8365
rect 52008 8271 52080 8319
rect 52008 8225 52021 8271
rect 52067 8225 52080 8271
rect 52008 8177 52080 8225
rect 52008 8131 52021 8177
rect 52067 8131 52080 8177
rect 52008 8083 52080 8131
rect 52008 8037 52021 8083
rect 52067 8037 52080 8083
rect 52008 7989 52080 8037
rect 52008 7943 52021 7989
rect 52067 7943 52080 7989
rect 52008 7895 52080 7943
rect 56144 8507 56157 8553
rect 56203 8507 56216 8553
rect 60280 8929 60352 8977
rect 60280 8883 60293 8929
rect 60339 8883 60352 8929
rect 60280 8835 60352 8883
rect 60280 8789 60293 8835
rect 60339 8789 60352 8835
rect 60280 8741 60352 8789
rect 60280 8695 60293 8741
rect 60339 8695 60352 8741
rect 60280 8647 60352 8695
rect 60280 8601 60293 8647
rect 60339 8601 60352 8647
rect 60280 8553 60352 8601
rect 56144 8459 56216 8507
rect 56144 8413 56157 8459
rect 56203 8413 56216 8459
rect 56144 8365 56216 8413
rect 56144 8319 56157 8365
rect 56203 8319 56216 8365
rect 56144 8271 56216 8319
rect 56144 8225 56157 8271
rect 56203 8225 56216 8271
rect 56144 8177 56216 8225
rect 56144 8131 56157 8177
rect 56203 8131 56216 8177
rect 56144 8083 56216 8131
rect 56144 8037 56157 8083
rect 56203 8037 56216 8083
rect 56144 7989 56216 8037
rect 56144 7943 56157 7989
rect 56203 7943 56216 7989
rect 52008 7849 52021 7895
rect 52067 7849 52080 7895
rect 56144 7895 56216 7943
rect 60280 8507 60293 8553
rect 60339 8507 60352 8553
rect 60280 8459 60352 8507
rect 60280 8413 60293 8459
rect 60339 8413 60352 8459
rect 60280 8365 60352 8413
rect 60280 8319 60293 8365
rect 60339 8319 60352 8365
rect 60280 8271 60352 8319
rect 60280 8225 60293 8271
rect 60339 8225 60352 8271
rect 60280 8177 60352 8225
rect 60280 8131 60293 8177
rect 60339 8131 60352 8177
rect 60280 8083 60352 8131
rect 60280 8037 60293 8083
rect 60339 8037 60352 8083
rect 60280 7989 60352 8037
rect 60280 7943 60293 7989
rect 60339 7943 60352 7989
rect 52008 7801 52080 7849
rect 52008 7755 52021 7801
rect 52067 7755 52080 7801
rect 52008 7707 52080 7755
rect 52008 7661 52021 7707
rect 52067 7661 52080 7707
rect 52008 7613 52080 7661
rect 52008 7567 52021 7613
rect 52067 7567 52080 7613
rect 52008 7519 52080 7567
rect 52008 7473 52021 7519
rect 52067 7473 52080 7519
rect 52008 7438 52080 7473
rect 56144 7849 56157 7895
rect 56203 7849 56216 7895
rect 60280 7895 60352 7943
rect 56144 7801 56216 7849
rect 56144 7755 56157 7801
rect 56203 7755 56216 7801
rect 56144 7707 56216 7755
rect 56144 7661 56157 7707
rect 56203 7661 56216 7707
rect 56144 7613 56216 7661
rect 56144 7567 56157 7613
rect 56203 7567 56216 7613
rect 56144 7519 56216 7567
rect 56144 7473 56157 7519
rect 56203 7473 56216 7519
rect 56144 7438 56216 7473
rect 60280 7849 60293 7895
rect 60339 7849 60352 7895
rect 60280 7801 60352 7849
rect 60280 7755 60293 7801
rect 60339 7755 60352 7801
rect 60280 7707 60352 7755
rect 60280 7661 60293 7707
rect 60339 7661 60352 7707
rect 60280 7613 60352 7661
rect 60280 7567 60293 7613
rect 60339 7567 60352 7613
rect 60280 7519 60352 7567
rect 60280 7473 60293 7519
rect 60339 7473 60352 7519
rect 60280 7438 60352 7473
rect 52008 7425 60352 7438
rect 52008 7379 52021 7425
rect 52067 7379 52115 7425
rect 52161 7379 52209 7425
rect 52255 7379 52303 7425
rect 52349 7379 52397 7425
rect 52443 7379 52491 7425
rect 52537 7379 52585 7425
rect 52631 7379 52679 7425
rect 52725 7379 52773 7425
rect 52819 7379 52867 7425
rect 52913 7379 52961 7425
rect 53007 7379 53055 7425
rect 53101 7379 53149 7425
rect 53195 7379 53243 7425
rect 53289 7379 53337 7425
rect 53383 7379 53431 7425
rect 53477 7379 53525 7425
rect 53571 7379 53619 7425
rect 53665 7379 53713 7425
rect 53759 7379 53807 7425
rect 53853 7379 53901 7425
rect 53947 7379 53995 7425
rect 54041 7379 54089 7425
rect 54135 7379 54183 7425
rect 54229 7379 54277 7425
rect 54323 7379 54371 7425
rect 54417 7379 54465 7425
rect 54511 7379 54559 7425
rect 54605 7379 54653 7425
rect 54699 7379 54747 7425
rect 54793 7379 54841 7425
rect 54887 7379 54935 7425
rect 54981 7379 55029 7425
rect 55075 7379 55123 7425
rect 55169 7379 55217 7425
rect 55263 7379 55311 7425
rect 55357 7379 55405 7425
rect 55451 7379 55499 7425
rect 55545 7379 55593 7425
rect 55639 7379 55687 7425
rect 55733 7379 55781 7425
rect 55827 7379 55875 7425
rect 55921 7379 55969 7425
rect 56015 7379 56063 7425
rect 56109 7379 56157 7425
rect 56203 7379 56251 7425
rect 56297 7379 56345 7425
rect 56391 7379 56439 7425
rect 56485 7379 56533 7425
rect 56579 7379 56627 7425
rect 56673 7379 56721 7425
rect 56767 7379 56815 7425
rect 56861 7379 56909 7425
rect 56955 7379 57003 7425
rect 57049 7379 57097 7425
rect 57143 7379 57191 7425
rect 57237 7379 57285 7425
rect 57331 7379 57379 7425
rect 57425 7379 57473 7425
rect 57519 7379 57567 7425
rect 57613 7379 57661 7425
rect 57707 7379 57755 7425
rect 57801 7379 57849 7425
rect 57895 7379 57943 7425
rect 57989 7379 58037 7425
rect 58083 7379 58131 7425
rect 58177 7379 58225 7425
rect 58271 7379 58319 7425
rect 58365 7379 58413 7425
rect 58459 7379 58507 7425
rect 58553 7379 58601 7425
rect 58647 7379 58695 7425
rect 58741 7379 58789 7425
rect 58835 7379 58883 7425
rect 58929 7379 58977 7425
rect 59023 7379 59071 7425
rect 59117 7379 59165 7425
rect 59211 7379 59259 7425
rect 59305 7379 59353 7425
rect 59399 7379 59447 7425
rect 59493 7379 59541 7425
rect 59587 7379 59635 7425
rect 59681 7379 59729 7425
rect 59775 7379 59823 7425
rect 59869 7379 59917 7425
rect 59963 7379 60011 7425
rect 60057 7379 60105 7425
rect 60151 7379 60199 7425
rect 60245 7379 60293 7425
rect 60339 7379 60352 7425
rect 52008 7366 60352 7379
rect 61704 12219 65912 12232
rect 61704 12173 61717 12219
rect 61763 12173 61811 12219
rect 61857 12173 61905 12219
rect 61951 12173 61999 12219
rect 62045 12173 62093 12219
rect 62139 12173 62187 12219
rect 62233 12173 62281 12219
rect 62327 12173 62375 12219
rect 62421 12173 62469 12219
rect 62515 12173 62563 12219
rect 62609 12173 62657 12219
rect 62703 12173 62751 12219
rect 62797 12173 62845 12219
rect 62891 12173 62939 12219
rect 62985 12173 63033 12219
rect 63079 12173 63127 12219
rect 63173 12173 63221 12219
rect 63267 12173 63315 12219
rect 63361 12173 63409 12219
rect 63455 12173 63503 12219
rect 63549 12173 63597 12219
rect 63643 12173 63691 12219
rect 63737 12173 63785 12219
rect 63831 12173 63879 12219
rect 63925 12173 63973 12219
rect 64019 12173 64067 12219
rect 64113 12173 64161 12219
rect 64207 12173 64255 12219
rect 64301 12173 64349 12219
rect 64395 12173 64443 12219
rect 64489 12173 64537 12219
rect 64583 12173 64631 12219
rect 64677 12173 64725 12219
rect 64771 12173 64819 12219
rect 64865 12173 64913 12219
rect 64959 12173 65007 12219
rect 65053 12173 65101 12219
rect 65147 12173 65195 12219
rect 65241 12173 65289 12219
rect 65335 12173 65383 12219
rect 65429 12173 65477 12219
rect 65523 12173 65571 12219
rect 65617 12173 65665 12219
rect 65711 12173 65759 12219
rect 65805 12173 65853 12219
rect 65899 12173 65912 12219
rect 61704 12160 65912 12173
rect 61704 12125 61776 12160
rect 61704 12079 61717 12125
rect 61763 12079 61776 12125
rect 61704 12031 61776 12079
rect 61704 11985 61717 12031
rect 61763 11985 61776 12031
rect 61704 11937 61776 11985
rect 61704 11891 61717 11937
rect 61763 11891 61776 11937
rect 61704 11843 61776 11891
rect 61704 11797 61717 11843
rect 61763 11797 61776 11843
rect 65840 12125 65912 12160
rect 65840 12079 65853 12125
rect 65899 12079 65912 12125
rect 65840 12031 65912 12079
rect 65840 11985 65853 12031
rect 65899 11985 65912 12031
rect 65840 11937 65912 11985
rect 65840 11891 65853 11937
rect 65899 11891 65912 11937
rect 65840 11843 65912 11891
rect 61704 11749 61776 11797
rect 65840 11797 65853 11843
rect 65899 11797 65912 11843
rect 61704 11703 61717 11749
rect 61763 11703 61776 11749
rect 61704 11655 61776 11703
rect 65840 11749 65912 11797
rect 65840 11703 65853 11749
rect 65899 11703 65912 11749
rect 61704 11609 61717 11655
rect 61763 11609 61776 11655
rect 61704 11561 61776 11609
rect 61704 11515 61717 11561
rect 61763 11515 61776 11561
rect 61704 11467 61776 11515
rect 61704 11421 61717 11467
rect 61763 11421 61776 11467
rect 61704 11373 61776 11421
rect 61704 11327 61717 11373
rect 61763 11327 61776 11373
rect 61704 11279 61776 11327
rect 61704 11233 61717 11279
rect 61763 11233 61776 11279
rect 61704 11185 61776 11233
rect 61704 11139 61717 11185
rect 61763 11139 61776 11185
rect 61704 11091 61776 11139
rect 61704 11045 61717 11091
rect 61763 11045 61776 11091
rect 65840 11655 65912 11703
rect 65840 11609 65853 11655
rect 65899 11609 65912 11655
rect 65840 11561 65912 11609
rect 65840 11515 65853 11561
rect 65899 11515 65912 11561
rect 65840 11467 65912 11515
rect 65840 11421 65853 11467
rect 65899 11421 65912 11467
rect 65840 11373 65912 11421
rect 65840 11327 65853 11373
rect 65899 11327 65912 11373
rect 65840 11279 65912 11327
rect 65840 11233 65853 11279
rect 65899 11233 65912 11279
rect 65840 11185 65912 11233
rect 65840 11139 65853 11185
rect 65899 11139 65912 11185
rect 65840 11091 65912 11139
rect 61704 10997 61776 11045
rect 61704 10951 61717 10997
rect 61763 10951 61776 10997
rect 61704 10903 61776 10951
rect 61704 10857 61717 10903
rect 61763 10857 61776 10903
rect 61704 10809 61776 10857
rect 61704 10763 61717 10809
rect 61763 10763 61776 10809
rect 61704 10715 61776 10763
rect 61704 10669 61717 10715
rect 61763 10669 61776 10715
rect 61704 10621 61776 10669
rect 65840 11045 65853 11091
rect 65899 11045 65912 11091
rect 65840 10997 65912 11045
rect 65840 10951 65853 10997
rect 65899 10951 65912 10997
rect 65840 10903 65912 10951
rect 65840 10857 65853 10903
rect 65899 10857 65912 10903
rect 65840 10809 65912 10857
rect 65840 10763 65853 10809
rect 65899 10763 65912 10809
rect 65840 10715 65912 10763
rect 65840 10669 65853 10715
rect 65899 10669 65912 10715
rect 61704 10575 61717 10621
rect 61763 10575 61776 10621
rect 61704 10527 61776 10575
rect 61704 10481 61717 10527
rect 61763 10481 61776 10527
rect 61704 10433 61776 10481
rect 61704 10387 61717 10433
rect 61763 10387 61776 10433
rect 61704 10339 61776 10387
rect 61704 10293 61717 10339
rect 61763 10293 61776 10339
rect 61704 10245 61776 10293
rect 61704 10199 61717 10245
rect 61763 10199 61776 10245
rect 61704 10151 61776 10199
rect 61704 10105 61717 10151
rect 61763 10105 61776 10151
rect 61704 10057 61776 10105
rect 61704 10011 61717 10057
rect 61763 10011 61776 10057
rect 65840 10621 65912 10669
rect 65840 10575 65853 10621
rect 65899 10575 65912 10621
rect 65840 10527 65912 10575
rect 65840 10481 65853 10527
rect 65899 10481 65912 10527
rect 65840 10433 65912 10481
rect 65840 10387 65853 10433
rect 65899 10387 65912 10433
rect 65840 10339 65912 10387
rect 65840 10293 65853 10339
rect 65899 10293 65912 10339
rect 65840 10245 65912 10293
rect 65840 10199 65853 10245
rect 65899 10199 65912 10245
rect 65840 10151 65912 10199
rect 65840 10105 65853 10151
rect 65899 10105 65912 10151
rect 65840 10057 65912 10105
rect 61704 9963 61776 10011
rect 61704 9917 61717 9963
rect 61763 9917 61776 9963
rect 61704 9869 61776 9917
rect 61704 9823 61717 9869
rect 61763 9823 61776 9869
rect 61704 9775 61776 9823
rect 61704 9729 61717 9775
rect 61763 9729 61776 9775
rect 61704 9681 61776 9729
rect 61704 9635 61717 9681
rect 61763 9635 61776 9681
rect 61704 9587 61776 9635
rect 61704 9541 61717 9587
rect 61763 9541 61776 9587
rect 65840 10011 65853 10057
rect 65899 10011 65912 10057
rect 65840 9963 65912 10011
rect 65840 9917 65853 9963
rect 65899 9917 65912 9963
rect 65840 9869 65912 9917
rect 65840 9823 65853 9869
rect 65899 9823 65912 9869
rect 65840 9775 65912 9823
rect 65840 9729 65853 9775
rect 65899 9729 65912 9775
rect 65840 9681 65912 9729
rect 65840 9635 65853 9681
rect 65899 9635 65912 9681
rect 65840 9587 65912 9635
rect 61704 9493 61776 9541
rect 61704 9447 61717 9493
rect 61763 9447 61776 9493
rect 61704 9399 61776 9447
rect 61704 9353 61717 9399
rect 61763 9353 61776 9399
rect 61704 9305 61776 9353
rect 61704 9259 61717 9305
rect 61763 9259 61776 9305
rect 61704 9211 61776 9259
rect 61704 9165 61717 9211
rect 61763 9165 61776 9211
rect 61704 9117 61776 9165
rect 61704 9071 61717 9117
rect 61763 9071 61776 9117
rect 61704 9023 61776 9071
rect 61704 8977 61717 9023
rect 61763 8977 61776 9023
rect 61704 8929 61776 8977
rect 65840 9541 65853 9587
rect 65899 9541 65912 9587
rect 65840 9493 65912 9541
rect 65840 9447 65853 9493
rect 65899 9447 65912 9493
rect 65840 9399 65912 9447
rect 65840 9353 65853 9399
rect 65899 9353 65912 9399
rect 65840 9305 65912 9353
rect 65840 9259 65853 9305
rect 65899 9259 65912 9305
rect 65840 9211 65912 9259
rect 65840 9165 65853 9211
rect 65899 9165 65912 9211
rect 65840 9117 65912 9165
rect 65840 9071 65853 9117
rect 65899 9071 65912 9117
rect 65840 9023 65912 9071
rect 65840 8977 65853 9023
rect 65899 8977 65912 9023
rect 61704 8883 61717 8929
rect 61763 8883 61776 8929
rect 61704 8835 61776 8883
rect 61704 8789 61717 8835
rect 61763 8789 61776 8835
rect 61704 8741 61776 8789
rect 61704 8695 61717 8741
rect 61763 8695 61776 8741
rect 61704 8647 61776 8695
rect 61704 8601 61717 8647
rect 61763 8601 61776 8647
rect 61704 8553 61776 8601
rect 61704 8507 61717 8553
rect 61763 8507 61776 8553
rect 65840 8929 65912 8977
rect 65840 8883 65853 8929
rect 65899 8883 65912 8929
rect 65840 8835 65912 8883
rect 65840 8789 65853 8835
rect 65899 8789 65912 8835
rect 65840 8741 65912 8789
rect 65840 8695 65853 8741
rect 65899 8695 65912 8741
rect 65840 8647 65912 8695
rect 65840 8601 65853 8647
rect 65899 8601 65912 8647
rect 65840 8553 65912 8601
rect 61704 8459 61776 8507
rect 61704 8413 61717 8459
rect 61763 8413 61776 8459
rect 61704 8365 61776 8413
rect 61704 8319 61717 8365
rect 61763 8319 61776 8365
rect 61704 8271 61776 8319
rect 61704 8225 61717 8271
rect 61763 8225 61776 8271
rect 61704 8177 61776 8225
rect 61704 8131 61717 8177
rect 61763 8131 61776 8177
rect 61704 8083 61776 8131
rect 61704 8037 61717 8083
rect 61763 8037 61776 8083
rect 61704 7989 61776 8037
rect 61704 7943 61717 7989
rect 61763 7943 61776 7989
rect 61704 7895 61776 7943
rect 65840 8507 65853 8553
rect 65899 8507 65912 8553
rect 65840 8459 65912 8507
rect 65840 8413 65853 8459
rect 65899 8413 65912 8459
rect 65840 8365 65912 8413
rect 65840 8319 65853 8365
rect 65899 8319 65912 8365
rect 65840 8271 65912 8319
rect 65840 8225 65853 8271
rect 65899 8225 65912 8271
rect 65840 8177 65912 8225
rect 65840 8131 65853 8177
rect 65899 8131 65912 8177
rect 65840 8083 65912 8131
rect 65840 8037 65853 8083
rect 65899 8037 65912 8083
rect 65840 7989 65912 8037
rect 65840 7943 65853 7989
rect 65899 7943 65912 7989
rect 61704 7849 61717 7895
rect 61763 7849 61776 7895
rect 65840 7895 65912 7943
rect 61704 7801 61776 7849
rect 61704 7755 61717 7801
rect 61763 7755 61776 7801
rect 61704 7707 61776 7755
rect 61704 7661 61717 7707
rect 61763 7661 61776 7707
rect 61704 7613 61776 7661
rect 61704 7567 61717 7613
rect 61763 7567 61776 7613
rect 61704 7519 61776 7567
rect 61704 7473 61717 7519
rect 61763 7473 61776 7519
rect 61704 7438 61776 7473
rect 65840 7849 65853 7895
rect 65899 7849 65912 7895
rect 65840 7801 65912 7849
rect 65840 7755 65853 7801
rect 65899 7755 65912 7801
rect 65840 7707 65912 7755
rect 65840 7661 65853 7707
rect 65899 7661 65912 7707
rect 65840 7613 65912 7661
rect 65840 7567 65853 7613
rect 65899 7567 65912 7613
rect 65840 7519 65912 7567
rect 65840 7473 65853 7519
rect 65899 7473 65912 7519
rect 65840 7438 65912 7473
rect 61704 7425 65912 7438
rect 61704 7379 61717 7425
rect 61763 7379 61811 7425
rect 61857 7379 61905 7425
rect 61951 7379 61999 7425
rect 62045 7379 62093 7425
rect 62139 7379 62187 7425
rect 62233 7379 62281 7425
rect 62327 7379 62375 7425
rect 62421 7379 62469 7425
rect 62515 7379 62563 7425
rect 62609 7379 62657 7425
rect 62703 7379 62751 7425
rect 62797 7379 62845 7425
rect 62891 7379 62939 7425
rect 62985 7379 63033 7425
rect 63079 7379 63127 7425
rect 63173 7379 63221 7425
rect 63267 7379 63315 7425
rect 63361 7379 63409 7425
rect 63455 7379 63503 7425
rect 63549 7379 63597 7425
rect 63643 7379 63691 7425
rect 63737 7379 63785 7425
rect 63831 7379 63879 7425
rect 63925 7379 63973 7425
rect 64019 7379 64067 7425
rect 64113 7379 64161 7425
rect 64207 7379 64255 7425
rect 64301 7379 64349 7425
rect 64395 7379 64443 7425
rect 64489 7379 64537 7425
rect 64583 7379 64631 7425
rect 64677 7379 64725 7425
rect 64771 7379 64819 7425
rect 64865 7379 64913 7425
rect 64959 7379 65007 7425
rect 65053 7379 65101 7425
rect 65147 7379 65195 7425
rect 65241 7379 65289 7425
rect 65335 7379 65383 7425
rect 65429 7379 65477 7425
rect 65523 7379 65571 7425
rect 65617 7379 65665 7425
rect 65711 7379 65759 7425
rect 65805 7379 65853 7425
rect 65899 7379 65912 7425
rect 61704 7366 65912 7379
rect 11887 7265 17035 7278
rect -3889 7196 -3872 7242
rect -3826 7196 -3809 7242
rect -3889 7144 -3809 7196
rect -3889 7098 -3872 7144
rect -3826 7098 -3809 7144
rect -3889 7046 -3809 7098
rect -3889 7000 -3872 7046
rect -3826 7000 -3809 7046
rect -3889 6948 -3809 7000
rect -3889 6902 -3872 6948
rect -3826 6902 -3809 6948
rect -3889 6850 -3809 6902
rect -3889 6804 -3872 6850
rect -3826 6804 -3809 6850
rect -3889 6752 -3809 6804
rect -3889 6706 -3872 6752
rect -3826 6706 -3809 6752
rect -3889 6654 -3809 6706
rect -3889 6608 -3872 6654
rect -3826 6608 -3809 6654
rect -3889 6556 -3809 6608
rect -3889 6510 -3872 6556
rect -3826 6510 -3809 6556
rect -3889 6458 -3809 6510
rect -3889 6412 -3872 6458
rect -3826 6412 -3809 6458
rect -3889 6360 -3809 6412
rect -3889 6314 -3872 6360
rect -3826 6314 -3809 6360
rect -3889 6262 -3809 6314
rect -3889 6216 -3872 6262
rect -3826 6216 -3809 6262
rect -3889 6164 -3809 6216
rect -3889 6118 -3872 6164
rect -3826 6118 -3809 6164
rect -3889 6066 -3809 6118
rect -3889 6020 -3872 6066
rect -3826 6020 -3809 6066
rect -3889 5968 -3809 6020
rect -3889 5922 -3872 5968
rect -3826 5922 -3809 5968
rect -3889 5870 -3809 5922
rect -3889 5824 -3872 5870
rect -3826 5824 -3809 5870
rect -3889 5772 -3809 5824
rect -3889 5726 -3872 5772
rect -3826 5726 -3809 5772
rect -3889 5674 -3809 5726
rect -3889 5628 -3872 5674
rect -3826 5628 -3809 5674
rect -3889 5576 -3809 5628
rect -3889 5530 -3872 5576
rect -3826 5530 -3809 5576
rect -3889 5478 -3809 5530
rect -3889 5432 -3872 5478
rect -3826 5432 -3809 5478
rect -3889 5380 -3809 5432
rect -3889 5334 -3872 5380
rect -3826 5334 -3809 5380
rect -3889 5282 -3809 5334
rect -3889 5236 -3872 5282
rect -3826 5236 -3809 5282
rect -3889 5184 -3809 5236
rect -3889 5138 -3872 5184
rect -3826 5138 -3809 5184
rect -3889 5086 -3809 5138
rect -3889 5040 -3872 5086
rect -3826 5040 -3809 5086
rect -3889 4988 -3809 5040
rect -3889 4942 -3872 4988
rect -3826 4942 -3809 4988
rect -3889 4890 -3809 4942
rect -3889 4844 -3872 4890
rect -3826 4844 -3809 4890
rect -3889 4792 -3809 4844
rect -3889 4746 -3872 4792
rect -3826 4746 -3809 4792
rect -3889 4694 -3809 4746
rect -3889 4648 -3872 4694
rect -3826 4648 -3809 4694
rect -3889 4596 -3809 4648
rect -3889 4550 -3872 4596
rect -3826 4550 -3809 4596
rect -3889 4498 -3809 4550
rect -7720 4407 -7640 4452
rect -3889 4452 -3872 4498
rect -3826 4452 -3809 4498
rect -3889 4407 -3809 4452
rect -7720 4390 -3809 4407
rect -7720 4344 -7703 4390
rect -7657 4344 -7605 4390
rect -7559 4344 -7507 4390
rect -7461 4344 -7409 4390
rect -7363 4344 -7311 4390
rect -7265 4344 -7213 4390
rect -7167 4344 -7115 4390
rect -7069 4344 -7017 4390
rect -6971 4344 -6919 4390
rect -6873 4344 -6821 4390
rect -6775 4344 -6723 4390
rect -6677 4344 -6625 4390
rect -6579 4344 -6527 4390
rect -6481 4344 -6429 4390
rect -6383 4344 -6331 4390
rect -6285 4344 -6233 4390
rect -6187 4344 -6135 4390
rect -6089 4344 -6037 4390
rect -5991 4344 -5939 4390
rect -5893 4344 -5841 4390
rect -5795 4344 -5743 4390
rect -5697 4344 -5645 4390
rect -5599 4344 -5547 4390
rect -5501 4344 -5449 4390
rect -5403 4344 -5351 4390
rect -5305 4344 -5253 4390
rect -5207 4344 -5155 4390
rect -5109 4344 -5057 4390
rect -5011 4344 -4959 4390
rect -4913 4344 -4861 4390
rect -4815 4344 -4763 4390
rect -4717 4344 -4665 4390
rect -4619 4344 -4567 4390
rect -4521 4344 -4469 4390
rect -4423 4344 -4371 4390
rect -4325 4344 -4273 4390
rect -4227 4344 -4175 4390
rect -4129 4344 -4077 4390
rect -4031 4344 -3979 4390
rect -3933 4344 -3872 4390
rect -3826 4344 -3809 4390
rect -7720 4327 -3809 4344
rect 916 4792 5030 4805
rect 916 4746 929 4792
rect 975 4746 1023 4792
rect 1069 4746 1117 4792
rect 1163 4746 1211 4792
rect 1257 4746 1305 4792
rect 1351 4746 1399 4792
rect 1445 4746 1493 4792
rect 1539 4746 1587 4792
rect 1633 4746 1681 4792
rect 1727 4746 1775 4792
rect 1821 4746 1869 4792
rect 1915 4746 1963 4792
rect 2009 4746 2057 4792
rect 2103 4746 2151 4792
rect 2197 4746 2245 4792
rect 2291 4746 2339 4792
rect 2385 4746 2433 4792
rect 2479 4746 2527 4792
rect 2573 4746 2621 4792
rect 2667 4746 2715 4792
rect 2761 4746 2809 4792
rect 2855 4746 2903 4792
rect 2949 4746 2997 4792
rect 3043 4746 3091 4792
rect 3137 4746 3185 4792
rect 3231 4746 3279 4792
rect 3325 4746 3373 4792
rect 3419 4746 3467 4792
rect 3513 4746 3561 4792
rect 3607 4746 3655 4792
rect 3701 4746 3749 4792
rect 3795 4746 3843 4792
rect 3889 4746 3937 4792
rect 3983 4746 4031 4792
rect 4077 4746 4125 4792
rect 4171 4746 4219 4792
rect 4265 4746 4313 4792
rect 4359 4746 4407 4792
rect 4453 4746 4501 4792
rect 4547 4746 4595 4792
rect 4641 4746 4689 4792
rect 4735 4746 4783 4792
rect 4829 4746 4877 4792
rect 4923 4746 4971 4792
rect 5017 4746 5030 4792
rect 916 4733 5030 4746
rect 916 4698 988 4733
rect 916 4652 929 4698
rect 975 4652 988 4698
rect 916 4604 988 4652
rect 916 4558 929 4604
rect 975 4558 988 4604
rect 4958 4698 5030 4733
rect 4958 4652 4971 4698
rect 5017 4652 5030 4698
rect 4958 4604 5030 4652
rect 916 4510 988 4558
rect 916 4464 929 4510
rect 975 4464 988 4510
rect 916 4416 988 4464
rect 4958 4558 4971 4604
rect 5017 4558 5030 4604
rect 4958 4510 5030 4558
rect 4958 4464 4971 4510
rect 5017 4464 5030 4510
rect 916 4370 929 4416
rect 975 4370 988 4416
rect 916 4322 988 4370
rect 916 4276 929 4322
rect 975 4276 988 4322
rect 916 4228 988 4276
rect 916 4182 929 4228
rect 975 4182 988 4228
rect 916 4134 988 4182
rect 916 4088 929 4134
rect 975 4088 988 4134
rect 916 4040 988 4088
rect 916 3994 929 4040
rect 975 3994 988 4040
rect 916 3946 988 3994
rect 916 3900 929 3946
rect 975 3900 988 3946
rect 916 3852 988 3900
rect 916 3806 929 3852
rect 975 3806 988 3852
rect 916 3758 988 3806
rect 916 3712 929 3758
rect 975 3712 988 3758
rect 916 3664 988 3712
rect 916 3618 929 3664
rect 975 3618 988 3664
rect 4958 4416 5030 4464
rect 4958 4370 4971 4416
rect 5017 4370 5030 4416
rect 4958 4322 5030 4370
rect 4958 4276 4971 4322
rect 5017 4276 5030 4322
rect 4958 4228 5030 4276
rect 4958 4182 4971 4228
rect 5017 4182 5030 4228
rect 4958 4134 5030 4182
rect 4958 4088 4971 4134
rect 5017 4088 5030 4134
rect 4958 4040 5030 4088
rect 4958 3994 4971 4040
rect 5017 3994 5030 4040
rect 4958 3946 5030 3994
rect 4958 3900 4971 3946
rect 5017 3900 5030 3946
rect 4958 3852 5030 3900
rect 4958 3806 4971 3852
rect 5017 3806 5030 3852
rect 4958 3758 5030 3806
rect 4958 3712 4971 3758
rect 5017 3712 5030 3758
rect 4958 3664 5030 3712
rect 916 3570 988 3618
rect 916 3524 929 3570
rect 975 3524 988 3570
rect 916 3476 988 3524
rect 916 3430 929 3476
rect 975 3430 988 3476
rect 916 3382 988 3430
rect 916 3336 929 3382
rect 975 3336 988 3382
rect 916 3288 988 3336
rect 916 3242 929 3288
rect 975 3242 988 3288
rect 916 3194 988 3242
rect 916 3148 929 3194
rect 975 3148 988 3194
rect 4958 3618 4971 3664
rect 5017 3618 5030 3664
rect 4958 3570 5030 3618
rect 4958 3524 4971 3570
rect 5017 3524 5030 3570
rect 4958 3476 5030 3524
rect 4958 3430 4971 3476
rect 5017 3430 5030 3476
rect 4958 3382 5030 3430
rect 4958 3336 4971 3382
rect 5017 3336 5030 3382
rect 4958 3288 5030 3336
rect 4958 3242 4971 3288
rect 5017 3242 5030 3288
rect 4958 3194 5030 3242
rect 916 3100 988 3148
rect 916 3054 929 3100
rect 975 3054 988 3100
rect 916 3006 988 3054
rect 916 2960 929 3006
rect 975 2960 988 3006
rect 916 2912 988 2960
rect 916 2866 929 2912
rect 975 2866 988 2912
rect 916 2818 988 2866
rect 916 2772 929 2818
rect 975 2772 988 2818
rect 916 2724 988 2772
rect 916 2678 929 2724
rect 975 2678 988 2724
rect 916 2630 988 2678
rect 916 2584 929 2630
rect 975 2584 988 2630
rect 916 2536 988 2584
rect 916 2490 929 2536
rect 975 2490 988 2536
rect 916 2442 988 2490
rect 916 2396 929 2442
rect 975 2396 988 2442
rect 916 2348 988 2396
rect 4958 3148 4971 3194
rect 5017 3148 5030 3194
rect 4958 3100 5030 3148
rect 4958 3054 4971 3100
rect 5017 3054 5030 3100
rect 4958 3006 5030 3054
rect 4958 2960 4971 3006
rect 5017 2960 5030 3006
rect 4958 2912 5030 2960
rect 4958 2866 4971 2912
rect 5017 2866 5030 2912
rect 4958 2818 5030 2866
rect 18193 5701 31801 5714
rect 18193 5655 18206 5701
rect 18252 5655 18300 5701
rect 18346 5655 18394 5701
rect 18440 5655 18488 5701
rect 18534 5655 18582 5701
rect 18628 5655 18676 5701
rect 18722 5655 18770 5701
rect 18816 5655 18864 5701
rect 18910 5655 18958 5701
rect 19004 5655 19052 5701
rect 19098 5655 19146 5701
rect 19192 5655 19240 5701
rect 19286 5655 19334 5701
rect 19380 5655 19428 5701
rect 19474 5655 19522 5701
rect 19568 5655 19616 5701
rect 19662 5655 19710 5701
rect 19756 5655 19804 5701
rect 19850 5655 19898 5701
rect 19944 5655 19992 5701
rect 20038 5655 20086 5701
rect 20132 5655 20180 5701
rect 20226 5655 20274 5701
rect 20320 5655 20368 5701
rect 20414 5655 20462 5701
rect 20508 5655 20556 5701
rect 20602 5655 20650 5701
rect 20696 5655 20744 5701
rect 20790 5655 20838 5701
rect 20884 5655 20932 5701
rect 20978 5655 21026 5701
rect 21072 5655 21120 5701
rect 21166 5655 21214 5701
rect 21260 5655 21308 5701
rect 21354 5655 21402 5701
rect 21448 5655 21496 5701
rect 21542 5655 21590 5701
rect 21636 5655 21684 5701
rect 21730 5655 21778 5701
rect 21824 5655 21872 5701
rect 21918 5655 21966 5701
rect 22012 5655 22060 5701
rect 22106 5655 22154 5701
rect 22200 5655 22248 5701
rect 22294 5655 22342 5701
rect 22388 5655 22436 5701
rect 22482 5655 22530 5701
rect 22576 5655 22624 5701
rect 22670 5655 22718 5701
rect 22764 5655 22812 5701
rect 22858 5655 22906 5701
rect 22952 5655 23000 5701
rect 23046 5655 23094 5701
rect 23140 5655 23188 5701
rect 23234 5655 23282 5701
rect 23328 5655 23376 5701
rect 23422 5655 23470 5701
rect 23516 5655 23564 5701
rect 23610 5655 23658 5701
rect 23704 5655 23752 5701
rect 23798 5655 23846 5701
rect 23892 5655 23940 5701
rect 23986 5655 24034 5701
rect 24080 5655 24128 5701
rect 24174 5655 24222 5701
rect 24268 5655 24316 5701
rect 24362 5655 24410 5701
rect 24456 5655 24504 5701
rect 24550 5655 24598 5701
rect 24644 5655 24692 5701
rect 24738 5655 24786 5701
rect 24832 5655 24880 5701
rect 24926 5655 24974 5701
rect 25020 5655 25068 5701
rect 25114 5655 25162 5701
rect 25208 5655 25256 5701
rect 25302 5655 25350 5701
rect 25396 5655 25444 5701
rect 25490 5655 25538 5701
rect 25584 5655 25632 5701
rect 25678 5655 25726 5701
rect 25772 5655 25820 5701
rect 25866 5655 25914 5701
rect 25960 5655 26008 5701
rect 26054 5655 26102 5701
rect 26148 5655 26196 5701
rect 26242 5655 26290 5701
rect 26336 5655 26384 5701
rect 26430 5655 26478 5701
rect 26524 5655 26572 5701
rect 26618 5655 26666 5701
rect 26712 5655 26760 5701
rect 26806 5655 26854 5701
rect 26900 5655 26948 5701
rect 26994 5655 27042 5701
rect 27088 5655 27136 5701
rect 27182 5655 27230 5701
rect 27276 5655 27324 5701
rect 27370 5655 27418 5701
rect 27464 5655 27512 5701
rect 27558 5655 27606 5701
rect 27652 5655 27700 5701
rect 27746 5655 27794 5701
rect 27840 5655 27888 5701
rect 27934 5655 27982 5701
rect 28028 5655 28076 5701
rect 28122 5655 28170 5701
rect 28216 5655 28264 5701
rect 28310 5655 28358 5701
rect 28404 5655 28452 5701
rect 28498 5655 28546 5701
rect 28592 5655 28640 5701
rect 28686 5655 28734 5701
rect 28780 5655 28828 5701
rect 28874 5655 28922 5701
rect 28968 5655 29016 5701
rect 29062 5655 29110 5701
rect 29156 5655 29204 5701
rect 29250 5655 29298 5701
rect 29344 5655 29392 5701
rect 29438 5655 29486 5701
rect 29532 5655 29580 5701
rect 29626 5655 29674 5701
rect 29720 5655 29768 5701
rect 29814 5655 29862 5701
rect 29908 5655 29956 5701
rect 30002 5655 30050 5701
rect 30096 5655 30144 5701
rect 30190 5655 30238 5701
rect 30284 5655 30332 5701
rect 30378 5655 30426 5701
rect 30472 5655 30520 5701
rect 30566 5655 30614 5701
rect 30660 5655 30708 5701
rect 30754 5655 30802 5701
rect 30848 5655 30896 5701
rect 30942 5655 30990 5701
rect 31036 5655 31084 5701
rect 31130 5655 31178 5701
rect 31224 5655 31272 5701
rect 31318 5655 31366 5701
rect 31412 5655 31460 5701
rect 31506 5655 31554 5701
rect 31600 5655 31648 5701
rect 31694 5655 31742 5701
rect 31788 5655 31801 5701
rect 18193 5642 31801 5655
rect 18193 5607 18265 5642
rect 18193 5561 18206 5607
rect 18252 5561 18265 5607
rect 18193 5513 18265 5561
rect 18193 5467 18206 5513
rect 18252 5467 18265 5513
rect 18193 5419 18265 5467
rect 18193 5373 18206 5419
rect 18252 5373 18265 5419
rect 18193 5325 18265 5373
rect 18193 5279 18206 5325
rect 18252 5279 18265 5325
rect 18193 5231 18265 5279
rect 18193 5185 18206 5231
rect 18252 5185 18265 5231
rect 18193 5137 18265 5185
rect 18193 5091 18206 5137
rect 18252 5091 18265 5137
rect 18193 5043 18265 5091
rect 18193 4997 18206 5043
rect 18252 4997 18265 5043
rect 18193 4949 18265 4997
rect 18193 4903 18206 4949
rect 18252 4903 18265 4949
rect 22987 5607 23059 5642
rect 22987 5561 23000 5607
rect 23046 5561 23059 5607
rect 22987 5513 23059 5561
rect 22987 5467 23000 5513
rect 23046 5467 23059 5513
rect 22987 5419 23059 5467
rect 22987 5373 23000 5419
rect 23046 5373 23059 5419
rect 22987 5325 23059 5373
rect 22987 5279 23000 5325
rect 23046 5279 23059 5325
rect 22987 5231 23059 5279
rect 22987 5185 23000 5231
rect 23046 5185 23059 5231
rect 22987 5137 23059 5185
rect 22987 5091 23000 5137
rect 23046 5091 23059 5137
rect 22987 5043 23059 5091
rect 28721 5607 28793 5642
rect 28721 5561 28734 5607
rect 28780 5561 28793 5607
rect 28721 5513 28793 5561
rect 28721 5467 28734 5513
rect 28780 5467 28793 5513
rect 28721 5419 28793 5467
rect 28721 5373 28734 5419
rect 28780 5373 28793 5419
rect 28721 5325 28793 5373
rect 28721 5279 28734 5325
rect 28780 5279 28793 5325
rect 28721 5231 28793 5279
rect 31729 5607 31801 5642
rect 31729 5561 31742 5607
rect 31788 5561 31801 5607
rect 31729 5513 31801 5561
rect 31729 5467 31742 5513
rect 31788 5467 31801 5513
rect 31729 5419 31801 5467
rect 31729 5373 31742 5419
rect 31788 5373 31801 5419
rect 31729 5325 31801 5373
rect 31729 5279 31742 5325
rect 31788 5279 31801 5325
rect 28721 5185 28734 5231
rect 28780 5185 28793 5231
rect 28721 5137 28793 5185
rect 28721 5091 28734 5137
rect 28780 5091 28793 5137
rect 22987 4997 23000 5043
rect 23046 4997 23059 5043
rect 22987 4949 23059 4997
rect 18193 4855 18265 4903
rect 18193 4809 18206 4855
rect 18252 4809 18265 4855
rect 18193 4761 18265 4809
rect 22987 4903 23000 4949
rect 23046 4903 23059 4949
rect 22987 4855 23059 4903
rect 22987 4809 23000 4855
rect 23046 4809 23059 4855
rect 18193 4715 18206 4761
rect 18252 4715 18265 4761
rect 18193 4667 18265 4715
rect 18193 4621 18206 4667
rect 18252 4621 18265 4667
rect 18193 4573 18265 4621
rect 18193 4527 18206 4573
rect 18252 4527 18265 4573
rect 4958 2772 4971 2818
rect 5017 2772 5030 2818
rect 4958 2724 5030 2772
rect 4958 2678 4971 2724
rect 5017 2678 5030 2724
rect 4958 2630 5030 2678
rect 4958 2584 4971 2630
rect 5017 2584 5030 2630
rect 4958 2536 5030 2584
rect 4958 2490 4971 2536
rect 5017 2490 5030 2536
rect 4958 2442 5030 2490
rect 4958 2396 4971 2442
rect 5017 2396 5030 2442
rect 916 2302 929 2348
rect 975 2302 988 2348
rect 916 2254 988 2302
rect 916 2208 929 2254
rect 975 2208 988 2254
rect 916 2160 988 2208
rect 916 2114 929 2160
rect 975 2114 988 2160
rect 916 2066 988 2114
rect 916 2020 929 2066
rect 975 2020 988 2066
rect 916 1972 988 2020
rect 916 1926 929 1972
rect 975 1926 988 1972
rect 916 1878 988 1926
rect 4958 2348 5030 2396
rect 4958 2302 4971 2348
rect 5017 2302 5030 2348
rect 4958 2254 5030 2302
rect 4958 2208 4971 2254
rect 5017 2208 5030 2254
rect 4958 2160 5030 2208
rect 4958 2114 4971 2160
rect 5017 2114 5030 2160
rect 4958 2066 5030 2114
rect 4958 2020 4971 2066
rect 5017 2020 5030 2066
rect 4958 1972 5030 2020
rect 4958 1926 4971 1972
rect 5017 1926 5030 1972
rect 916 1832 929 1878
rect 975 1832 988 1878
rect 916 1784 988 1832
rect 4958 1878 5030 1926
rect 4958 1832 4971 1878
rect 5017 1832 5030 1878
rect 916 1738 929 1784
rect 975 1738 988 1784
rect 4958 1784 5030 1832
rect 916 1690 988 1738
rect 4958 1738 4971 1784
rect 5017 1738 5030 1784
rect 916 1644 929 1690
rect 975 1644 988 1690
rect 916 1596 988 1644
rect 916 1550 929 1596
rect 975 1550 988 1596
rect 916 1515 988 1550
rect 4958 1690 5030 1738
rect 4958 1644 4971 1690
rect 5017 1644 5030 1690
rect 4958 1596 5030 1644
rect 4958 1550 4971 1596
rect 5017 1550 5030 1596
rect 4958 1515 5030 1550
rect 916 1502 5030 1515
rect 916 1456 929 1502
rect 975 1456 1023 1502
rect 1069 1456 1117 1502
rect 1163 1456 1211 1502
rect 1257 1456 1305 1502
rect 1351 1456 1399 1502
rect 1445 1456 1493 1502
rect 1539 1456 1587 1502
rect 1633 1456 1681 1502
rect 1727 1456 1775 1502
rect 1821 1456 1869 1502
rect 1915 1456 1963 1502
rect 2009 1456 2057 1502
rect 2103 1456 2151 1502
rect 2197 1456 2245 1502
rect 2291 1456 2339 1502
rect 2385 1456 2433 1502
rect 2479 1456 2527 1502
rect 2573 1456 2621 1502
rect 2667 1456 2715 1502
rect 2761 1456 2809 1502
rect 2855 1456 2903 1502
rect 2949 1456 2997 1502
rect 3043 1456 3091 1502
rect 3137 1456 3185 1502
rect 3231 1456 3279 1502
rect 3325 1456 3373 1502
rect 3419 1456 3467 1502
rect 3513 1456 3561 1502
rect 3607 1456 3655 1502
rect 3701 1456 3749 1502
rect 3795 1456 3843 1502
rect 3889 1456 3937 1502
rect 3983 1456 4031 1502
rect 4077 1456 4125 1502
rect 4171 1456 4219 1502
rect 4265 1456 4313 1502
rect 4359 1456 4407 1502
rect 4453 1456 4501 1502
rect 4547 1456 4595 1502
rect 4641 1456 4689 1502
rect 4735 1456 4783 1502
rect 4829 1456 4877 1502
rect 4923 1456 4971 1502
rect 5017 1456 5030 1502
rect 916 1443 5030 1456
rect 18193 4479 18265 4527
rect 18193 4433 18206 4479
rect 18252 4433 18265 4479
rect 18193 4385 18265 4433
rect 18193 4339 18206 4385
rect 18252 4339 18265 4385
rect 18193 4291 18265 4339
rect 18193 4245 18206 4291
rect 18252 4245 18265 4291
rect 18193 4197 18265 4245
rect 18193 4151 18206 4197
rect 18252 4151 18265 4197
rect 22987 4761 23059 4809
rect 22987 4715 23000 4761
rect 23046 4715 23059 4761
rect 22987 4667 23059 4715
rect 22987 4621 23000 4667
rect 23046 4621 23059 4667
rect 22987 4573 23059 4621
rect 22987 4527 23000 4573
rect 23046 4527 23059 4573
rect 22987 4479 23059 4527
rect 22987 4433 23000 4479
rect 23046 4433 23059 4479
rect 22987 4385 23059 4433
rect 22987 4339 23000 4385
rect 23046 4339 23059 4385
rect 22987 4291 23059 4339
rect 22987 4245 23000 4291
rect 23046 4245 23059 4291
rect 22987 4197 23059 4245
rect 18193 4103 18265 4151
rect 18193 4057 18206 4103
rect 18252 4057 18265 4103
rect 18193 4009 18265 4057
rect 22987 4151 23000 4197
rect 23046 4151 23059 4197
rect 22987 4103 23059 4151
rect 22987 4057 23000 4103
rect 23046 4057 23059 4103
rect 18193 3963 18206 4009
rect 18252 3963 18265 4009
rect 18193 3915 18265 3963
rect 18193 3869 18206 3915
rect 18252 3869 18265 3915
rect 18193 3821 18265 3869
rect 18193 3775 18206 3821
rect 18252 3775 18265 3821
rect 18193 3727 18265 3775
rect 18193 3681 18206 3727
rect 18252 3681 18265 3727
rect 18193 3633 18265 3681
rect 18193 3587 18206 3633
rect 18252 3587 18265 3633
rect 18193 3539 18265 3587
rect 18193 3493 18206 3539
rect 18252 3493 18265 3539
rect 18193 3445 18265 3493
rect 18193 3399 18206 3445
rect 18252 3399 18265 3445
rect 22987 4009 23059 4057
rect 22987 3963 23000 4009
rect 23046 3963 23059 4009
rect 22987 3915 23059 3963
rect 22987 3869 23000 3915
rect 23046 3869 23059 3915
rect 22987 3821 23059 3869
rect 22987 3775 23000 3821
rect 23046 3775 23059 3821
rect 22987 3727 23059 3775
rect 22987 3681 23000 3727
rect 23046 3681 23059 3727
rect 22987 3633 23059 3681
rect 22987 3587 23000 3633
rect 23046 3587 23059 3633
rect 22987 3539 23059 3587
rect 23500 5007 28300 5079
rect 23500 3627 23572 5007
rect 23948 3627 24020 5007
rect 24396 3627 24468 5007
rect 25124 3627 25196 5007
rect 25852 3627 25924 5007
rect 26580 3627 26652 5007
rect 27308 3627 27380 5007
rect 27756 3627 27852 5007
rect 28228 3627 28300 5007
rect 23500 3555 28300 3627
rect 28721 5043 28793 5091
rect 28721 4997 28734 5043
rect 28780 4997 28793 5043
rect 28721 4949 28793 4997
rect 28721 4903 28734 4949
rect 28780 4903 28793 4949
rect 28721 4855 28793 4903
rect 28721 4809 28734 4855
rect 28780 4809 28793 4855
rect 28721 4761 28793 4809
rect 28721 4715 28734 4761
rect 28780 4715 28793 4761
rect 28721 4667 28793 4715
rect 28721 4621 28734 4667
rect 28780 4621 28793 4667
rect 28721 4573 28793 4621
rect 28721 4527 28734 4573
rect 28780 4527 28793 4573
rect 28721 4479 28793 4527
rect 28721 4433 28734 4479
rect 28780 4433 28793 4479
rect 28721 4385 28793 4433
rect 28721 4339 28734 4385
rect 28780 4339 28793 4385
rect 28721 4291 28793 4339
rect 28721 4245 28734 4291
rect 28780 4245 28793 4291
rect 28721 4197 28793 4245
rect 28721 4151 28734 4197
rect 28780 4151 28793 4197
rect 28721 4103 28793 4151
rect 28721 4057 28734 4103
rect 28780 4057 28793 4103
rect 28721 4009 28793 4057
rect 28721 3963 28734 4009
rect 28780 3963 28793 4009
rect 28721 3915 28793 3963
rect 28721 3869 28734 3915
rect 28780 3869 28793 3915
rect 28721 3821 28793 3869
rect 28721 3775 28734 3821
rect 28780 3775 28793 3821
rect 28721 3727 28793 3775
rect 28721 3681 28734 3727
rect 28780 3681 28793 3727
rect 28721 3633 28793 3681
rect 28721 3587 28734 3633
rect 28780 3587 28793 3633
rect 22987 3493 23000 3539
rect 23046 3493 23059 3539
rect 22987 3445 23059 3493
rect 18193 3351 18265 3399
rect 18193 3305 18206 3351
rect 18252 3305 18265 3351
rect 22987 3399 23000 3445
rect 23046 3399 23059 3445
rect 22987 3351 23059 3399
rect 18193 3257 18265 3305
rect 18193 3211 18206 3257
rect 18252 3211 18265 3257
rect 18193 3163 18265 3211
rect 18193 3117 18206 3163
rect 18252 3117 18265 3163
rect 18193 3069 18265 3117
rect 18193 3023 18206 3069
rect 18252 3023 18265 3069
rect 18193 2975 18265 3023
rect 18193 2929 18206 2975
rect 18252 2929 18265 2975
rect 18193 2881 18265 2929
rect 18193 2835 18206 2881
rect 18252 2835 18265 2881
rect 18193 2787 18265 2835
rect 18193 2741 18206 2787
rect 18252 2741 18265 2787
rect 18193 2693 18265 2741
rect 22987 3305 23000 3351
rect 23046 3305 23059 3351
rect 22987 3257 23059 3305
rect 22987 3211 23000 3257
rect 23046 3211 23059 3257
rect 22987 3163 23059 3211
rect 22987 3117 23000 3163
rect 23046 3117 23059 3163
rect 22987 3069 23059 3117
rect 28721 3539 28793 3587
rect 28721 3493 28734 3539
rect 28780 3493 28793 3539
rect 29126 5191 31382 5263
rect 29126 3571 29198 5191
rect 29574 3571 29646 5191
rect 30862 3571 30934 5191
rect 31310 3571 31382 5191
rect 29126 3499 31382 3571
rect 31729 5231 31801 5279
rect 31729 5185 31742 5231
rect 31788 5185 31801 5231
rect 31729 5137 31801 5185
rect 31729 5091 31742 5137
rect 31788 5091 31801 5137
rect 31729 5043 31801 5091
rect 31729 4997 31742 5043
rect 31788 4997 31801 5043
rect 31729 4949 31801 4997
rect 31729 4903 31742 4949
rect 31788 4903 31801 4949
rect 31729 4855 31801 4903
rect 31729 4809 31742 4855
rect 31788 4809 31801 4855
rect 31729 4761 31801 4809
rect 31729 4715 31742 4761
rect 31788 4715 31801 4761
rect 31729 4667 31801 4715
rect 31729 4621 31742 4667
rect 31788 4621 31801 4667
rect 31729 4573 31801 4621
rect 31729 4527 31742 4573
rect 31788 4527 31801 4573
rect 31729 4479 31801 4527
rect 31729 4433 31742 4479
rect 31788 4433 31801 4479
rect 31729 4385 31801 4433
rect 31729 4339 31742 4385
rect 31788 4339 31801 4385
rect 31729 4291 31801 4339
rect 31729 4245 31742 4291
rect 31788 4245 31801 4291
rect 31729 4197 31801 4245
rect 31729 4151 31742 4197
rect 31788 4151 31801 4197
rect 31729 4103 31801 4151
rect 31729 4057 31742 4103
rect 31788 4057 31801 4103
rect 31729 4009 31801 4057
rect 31729 3963 31742 4009
rect 31788 3963 31801 4009
rect 31729 3915 31801 3963
rect 31729 3869 31742 3915
rect 31788 3869 31801 3915
rect 31729 3821 31801 3869
rect 31729 3775 31742 3821
rect 31788 3775 31801 3821
rect 31729 3727 31801 3775
rect 31729 3681 31742 3727
rect 31788 3681 31801 3727
rect 31729 3633 31801 3681
rect 31729 3587 31742 3633
rect 31788 3587 31801 3633
rect 31729 3539 31801 3587
rect 28721 3445 28793 3493
rect 28721 3399 28734 3445
rect 28780 3399 28793 3445
rect 28721 3351 28793 3399
rect 28721 3305 28734 3351
rect 28780 3305 28793 3351
rect 28721 3257 28793 3305
rect 28721 3211 28734 3257
rect 28780 3211 28793 3257
rect 31729 3493 31742 3539
rect 31788 3493 31801 3539
rect 31729 3445 31801 3493
rect 31729 3399 31742 3445
rect 31788 3399 31801 3445
rect 31729 3351 31801 3399
rect 31729 3305 31742 3351
rect 31788 3305 31801 3351
rect 31729 3257 31801 3305
rect 28721 3163 28793 3211
rect 28721 3117 28734 3163
rect 28780 3117 28793 3163
rect 22987 3023 23000 3069
rect 23046 3023 23059 3069
rect 22987 2975 23059 3023
rect 22987 2929 23000 2975
rect 23046 2929 23059 2975
rect 22987 2881 23059 2929
rect 22987 2835 23000 2881
rect 23046 2835 23059 2881
rect 22987 2787 23059 2835
rect 22987 2741 23000 2787
rect 23046 2741 23059 2787
rect 18193 2647 18206 2693
rect 18252 2647 18265 2693
rect 18193 2599 18265 2647
rect 18193 2553 18206 2599
rect 18252 2553 18265 2599
rect 18193 2505 18265 2553
rect 18193 2459 18206 2505
rect 18252 2459 18265 2505
rect 18193 2411 18265 2459
rect 18193 2365 18206 2411
rect 18252 2365 18265 2411
rect 18193 2317 18265 2365
rect 18193 2271 18206 2317
rect 18252 2271 18265 2317
rect 18193 2223 18265 2271
rect 18193 2177 18206 2223
rect 18252 2177 18265 2223
rect 18193 2129 18265 2177
rect 18193 2083 18206 2129
rect 18252 2083 18265 2129
rect 18193 2035 18265 2083
rect 18193 1989 18206 2035
rect 18252 1989 18265 2035
rect 18193 1941 18265 1989
rect 22987 2693 23059 2741
rect 22987 2647 23000 2693
rect 23046 2647 23059 2693
rect 22987 2599 23059 2647
rect 22987 2553 23000 2599
rect 23046 2553 23059 2599
rect 22987 2505 23059 2553
rect 22987 2459 23000 2505
rect 23046 2459 23059 2505
rect 22987 2411 23059 2459
rect 22987 2365 23000 2411
rect 23046 2365 23059 2411
rect 22987 2317 23059 2365
rect 22987 2271 23000 2317
rect 23046 2271 23059 2317
rect 22987 2223 23059 2271
rect 22987 2177 23000 2223
rect 23046 2177 23059 2223
rect 22987 2129 23059 2177
rect 22987 2083 23000 2129
rect 23046 2083 23059 2129
rect 22987 2035 23059 2083
rect 22987 1989 23000 2035
rect 23046 1989 23059 2035
rect 18193 1895 18206 1941
rect 18252 1895 18265 1941
rect 18193 1847 18265 1895
rect 18193 1801 18206 1847
rect 18252 1801 18265 1847
rect 22987 1941 23059 1989
rect 22987 1895 23000 1941
rect 23046 1895 23059 1941
rect 22987 1847 23059 1895
rect 18193 1753 18265 1801
rect 18193 1707 18206 1753
rect 18252 1707 18265 1753
rect 18193 1659 18265 1707
rect 18193 1613 18206 1659
rect 18252 1613 18265 1659
rect 18193 1565 18265 1613
rect 18193 1519 18206 1565
rect 18252 1519 18265 1565
rect 18193 1471 18265 1519
rect 18193 1425 18206 1471
rect 18252 1425 18265 1471
rect 18193 1377 18265 1425
rect 18193 1331 18206 1377
rect 18252 1331 18265 1377
rect 18193 1283 18265 1331
rect 18193 1237 18206 1283
rect 18252 1237 18265 1283
rect 18193 1189 18265 1237
rect 18193 1143 18206 1189
rect 18252 1143 18265 1189
rect 18193 1108 18265 1143
rect 22987 1801 23000 1847
rect 23046 1801 23059 1847
rect 22987 1753 23059 1801
rect 22987 1707 23000 1753
rect 23046 1707 23059 1753
rect 22987 1659 23059 1707
rect 22987 1613 23000 1659
rect 23046 1613 23059 1659
rect 22987 1565 23059 1613
rect 23500 3035 28300 3107
rect 23500 1655 23572 3035
rect 23948 1655 24020 3035
rect 24396 1655 24468 3035
rect 25124 1655 25196 3035
rect 25852 1655 25924 3035
rect 26580 1655 26652 3035
rect 27308 1655 27380 3035
rect 27756 1655 27852 3035
rect 28228 1655 28300 3035
rect 23500 1583 28300 1655
rect 28721 3069 28793 3117
rect 28721 3023 28734 3069
rect 28780 3023 28793 3069
rect 28721 2975 28793 3023
rect 28721 2929 28734 2975
rect 28780 2929 28793 2975
rect 28721 2881 28793 2929
rect 28721 2835 28734 2881
rect 28780 2835 28793 2881
rect 28721 2787 28793 2835
rect 28721 2741 28734 2787
rect 28780 2741 28793 2787
rect 28721 2693 28793 2741
rect 28721 2647 28734 2693
rect 28780 2647 28793 2693
rect 28721 2599 28793 2647
rect 28721 2553 28734 2599
rect 28780 2553 28793 2599
rect 28721 2505 28793 2553
rect 28721 2459 28734 2505
rect 28780 2459 28793 2505
rect 28721 2411 28793 2459
rect 28721 2365 28734 2411
rect 28780 2365 28793 2411
rect 28721 2317 28793 2365
rect 28721 2271 28734 2317
rect 28780 2271 28793 2317
rect 28721 2223 28793 2271
rect 28721 2177 28734 2223
rect 28780 2177 28793 2223
rect 28721 2129 28793 2177
rect 28721 2083 28734 2129
rect 28780 2083 28793 2129
rect 28721 2035 28793 2083
rect 28721 1989 28734 2035
rect 28780 1989 28793 2035
rect 28721 1941 28793 1989
rect 28721 1895 28734 1941
rect 28780 1895 28793 1941
rect 28721 1847 28793 1895
rect 28721 1801 28734 1847
rect 28780 1801 28793 1847
rect 28721 1753 28793 1801
rect 28721 1707 28734 1753
rect 28780 1707 28793 1753
rect 28721 1659 28793 1707
rect 28721 1613 28734 1659
rect 28780 1613 28793 1659
rect 22987 1519 23000 1565
rect 23046 1519 23059 1565
rect 22987 1471 23059 1519
rect 22987 1425 23000 1471
rect 23046 1425 23059 1471
rect 22987 1377 23059 1425
rect 22987 1331 23000 1377
rect 23046 1331 23059 1377
rect 22987 1283 23059 1331
rect 22987 1237 23000 1283
rect 23046 1237 23059 1283
rect 22987 1189 23059 1237
rect 22987 1143 23000 1189
rect 23046 1143 23059 1189
rect 22987 1108 23059 1143
rect 28721 1565 28793 1613
rect 28721 1519 28734 1565
rect 28780 1519 28793 1565
rect 28721 1471 28793 1519
rect 29126 3179 31382 3251
rect 29126 1559 29198 3179
rect 29574 1559 29646 3179
rect 30862 1559 30934 3179
rect 31310 1559 31382 3179
rect 29126 1487 31382 1559
rect 31729 3211 31742 3257
rect 31788 3211 31801 3257
rect 31729 3163 31801 3211
rect 31729 3117 31742 3163
rect 31788 3117 31801 3163
rect 31729 3069 31801 3117
rect 31729 3023 31742 3069
rect 31788 3023 31801 3069
rect 31729 2975 31801 3023
rect 31729 2929 31742 2975
rect 31788 2929 31801 2975
rect 31729 2881 31801 2929
rect 31729 2835 31742 2881
rect 31788 2835 31801 2881
rect 31729 2787 31801 2835
rect 31729 2741 31742 2787
rect 31788 2741 31801 2787
rect 31729 2693 31801 2741
rect 31729 2647 31742 2693
rect 31788 2647 31801 2693
rect 31729 2599 31801 2647
rect 31729 2553 31742 2599
rect 31788 2553 31801 2599
rect 31729 2505 31801 2553
rect 31729 2459 31742 2505
rect 31788 2459 31801 2505
rect 31729 2411 31801 2459
rect 31729 2365 31742 2411
rect 31788 2365 31801 2411
rect 31729 2317 31801 2365
rect 31729 2271 31742 2317
rect 31788 2271 31801 2317
rect 31729 2223 31801 2271
rect 31729 2177 31742 2223
rect 31788 2177 31801 2223
rect 31729 2129 31801 2177
rect 31729 2083 31742 2129
rect 31788 2083 31801 2129
rect 31729 2035 31801 2083
rect 31729 1989 31742 2035
rect 31788 1989 31801 2035
rect 31729 1941 31801 1989
rect 31729 1895 31742 1941
rect 31788 1895 31801 1941
rect 31729 1847 31801 1895
rect 31729 1801 31742 1847
rect 31788 1801 31801 1847
rect 31729 1753 31801 1801
rect 31729 1707 31742 1753
rect 31788 1707 31801 1753
rect 31729 1659 31801 1707
rect 31729 1613 31742 1659
rect 31788 1613 31801 1659
rect 31729 1565 31801 1613
rect 31729 1519 31742 1565
rect 31788 1519 31801 1565
rect 28721 1425 28734 1471
rect 28780 1425 28793 1471
rect 28721 1377 28793 1425
rect 28721 1331 28734 1377
rect 28780 1331 28793 1377
rect 28721 1283 28793 1331
rect 28721 1237 28734 1283
rect 28780 1237 28793 1283
rect 28721 1189 28793 1237
rect 28721 1143 28734 1189
rect 28780 1143 28793 1189
rect 28721 1108 28793 1143
rect 31729 1471 31801 1519
rect 31729 1425 31742 1471
rect 31788 1425 31801 1471
rect 31729 1377 31801 1425
rect 31729 1331 31742 1377
rect 31788 1331 31801 1377
rect 31729 1283 31801 1331
rect 31729 1237 31742 1283
rect 31788 1237 31801 1283
rect 31729 1189 31801 1237
rect 31729 1143 31742 1189
rect 31788 1143 31801 1189
rect 31729 1108 31801 1143
rect 18193 1095 31801 1108
rect 18193 1049 18206 1095
rect 18252 1049 18300 1095
rect 18346 1049 18394 1095
rect 18440 1049 18488 1095
rect 18534 1049 18582 1095
rect 18628 1049 18676 1095
rect 18722 1049 18770 1095
rect 18816 1049 18864 1095
rect 18910 1049 18958 1095
rect 19004 1049 19052 1095
rect 19098 1049 19146 1095
rect 19192 1049 19240 1095
rect 19286 1049 19334 1095
rect 19380 1049 19428 1095
rect 19474 1049 19522 1095
rect 19568 1049 19616 1095
rect 19662 1049 19710 1095
rect 19756 1049 19804 1095
rect 19850 1049 19898 1095
rect 19944 1049 19992 1095
rect 20038 1049 20086 1095
rect 20132 1049 20180 1095
rect 20226 1049 20274 1095
rect 20320 1049 20368 1095
rect 20414 1049 20462 1095
rect 20508 1049 20556 1095
rect 20602 1049 20650 1095
rect 20696 1049 20744 1095
rect 20790 1049 20838 1095
rect 20884 1049 20932 1095
rect 20978 1049 21026 1095
rect 21072 1049 21120 1095
rect 21166 1049 21214 1095
rect 21260 1049 21308 1095
rect 21354 1049 21402 1095
rect 21448 1049 21496 1095
rect 21542 1049 21590 1095
rect 21636 1049 21684 1095
rect 21730 1049 21778 1095
rect 21824 1049 21872 1095
rect 21918 1049 21966 1095
rect 22012 1049 22060 1095
rect 22106 1049 22154 1095
rect 22200 1049 22248 1095
rect 22294 1049 22342 1095
rect 22388 1049 22436 1095
rect 22482 1049 22530 1095
rect 22576 1049 22624 1095
rect 22670 1049 22718 1095
rect 22764 1049 22812 1095
rect 22858 1049 22906 1095
rect 22952 1049 23000 1095
rect 23046 1049 23094 1095
rect 23140 1049 23188 1095
rect 23234 1049 23282 1095
rect 23328 1049 23376 1095
rect 23422 1049 23470 1095
rect 23516 1049 23564 1095
rect 23610 1049 23658 1095
rect 23704 1049 23752 1095
rect 23798 1049 23846 1095
rect 23892 1049 23940 1095
rect 23986 1049 24034 1095
rect 24080 1049 24128 1095
rect 24174 1049 24222 1095
rect 24268 1049 24316 1095
rect 24362 1049 24410 1095
rect 24456 1049 24504 1095
rect 24550 1049 24598 1095
rect 24644 1049 24692 1095
rect 24738 1049 24786 1095
rect 24832 1049 24880 1095
rect 24926 1049 24974 1095
rect 25020 1049 25068 1095
rect 25114 1049 25162 1095
rect 25208 1049 25256 1095
rect 25302 1049 25350 1095
rect 25396 1049 25444 1095
rect 25490 1049 25538 1095
rect 25584 1049 25632 1095
rect 25678 1049 25726 1095
rect 25772 1049 25820 1095
rect 25866 1049 25914 1095
rect 25960 1049 26008 1095
rect 26054 1049 26102 1095
rect 26148 1049 26196 1095
rect 26242 1049 26290 1095
rect 26336 1049 26384 1095
rect 26430 1049 26478 1095
rect 26524 1049 26572 1095
rect 26618 1049 26666 1095
rect 26712 1049 26760 1095
rect 26806 1049 26854 1095
rect 26900 1049 26948 1095
rect 26994 1049 27042 1095
rect 27088 1049 27136 1095
rect 27182 1049 27230 1095
rect 27276 1049 27324 1095
rect 27370 1049 27418 1095
rect 27464 1049 27512 1095
rect 27558 1049 27606 1095
rect 27652 1049 27700 1095
rect 27746 1049 27794 1095
rect 27840 1049 27888 1095
rect 27934 1049 27982 1095
rect 28028 1049 28076 1095
rect 28122 1049 28170 1095
rect 28216 1049 28264 1095
rect 28310 1049 28358 1095
rect 28404 1049 28452 1095
rect 28498 1049 28546 1095
rect 28592 1049 28640 1095
rect 28686 1049 28734 1095
rect 28780 1049 28828 1095
rect 28874 1049 28922 1095
rect 28968 1049 29016 1095
rect 29062 1049 29110 1095
rect 29156 1049 29204 1095
rect 29250 1049 29298 1095
rect 29344 1049 29392 1095
rect 29438 1049 29486 1095
rect 29532 1049 29580 1095
rect 29626 1049 29674 1095
rect 29720 1049 29768 1095
rect 29814 1049 29862 1095
rect 29908 1049 29956 1095
rect 30002 1049 30050 1095
rect 30096 1049 30144 1095
rect 30190 1049 30238 1095
rect 30284 1049 30332 1095
rect 30378 1049 30426 1095
rect 30472 1049 30520 1095
rect 30566 1049 30614 1095
rect 30660 1049 30708 1095
rect 30754 1049 30802 1095
rect 30848 1049 30896 1095
rect 30942 1049 30990 1095
rect 31036 1049 31084 1095
rect 31130 1049 31178 1095
rect 31224 1049 31272 1095
rect 31318 1049 31366 1095
rect 31412 1049 31460 1095
rect 31506 1049 31554 1095
rect 31600 1049 31648 1095
rect 31694 1049 31742 1095
rect 31788 1049 31801 1095
rect 18193 1036 31801 1049
<< psubdiffcont >>
rect 6262 14619 6308 14665
rect 6356 14619 6402 14665
rect 6450 14619 6496 14665
rect 6544 14619 6590 14665
rect 6638 14619 6684 14665
rect 6732 14619 6778 14665
rect 6826 14619 6872 14665
rect 6920 14619 6966 14665
rect 7014 14619 7060 14665
rect 7108 14619 7154 14665
rect 7202 14619 7248 14665
rect 7296 14619 7342 14665
rect 7390 14619 7436 14665
rect 7484 14619 7530 14665
rect 7578 14619 7624 14665
rect 7672 14619 7718 14665
rect 7766 14619 7812 14665
rect 7860 14619 7906 14665
rect 7954 14619 8000 14665
rect 8048 14619 8094 14665
rect 8142 14619 8188 14665
rect 8236 14619 8282 14665
rect 8330 14619 8376 14665
rect 8424 14619 8470 14665
rect 8518 14619 8564 14665
rect 6262 14525 6308 14571
rect 6262 14431 6308 14477
rect 6262 14337 6308 14383
rect 8518 14525 8564 14571
rect 8518 14431 8564 14477
rect 8518 14337 8564 14383
rect 6262 14243 6308 14289
rect 6262 14149 6308 14195
rect 6262 14055 6308 14101
rect 6262 13961 6308 14007
rect 6262 13867 6308 13913
rect 6262 13773 6308 13819
rect 6262 13679 6308 13725
rect 8518 14243 8564 14289
rect 8518 14149 8564 14195
rect 8518 14055 8564 14101
rect 8518 13961 8564 14007
rect 8518 13867 8564 13913
rect 8518 13773 8564 13819
rect 6262 13585 6308 13631
rect 6262 13491 6308 13537
rect 6262 13397 6308 13443
rect 8518 13679 8564 13725
rect 8518 13585 8564 13631
rect 8518 13491 8564 13537
rect 6262 13303 6308 13349
rect 6262 13209 6308 13255
rect 6262 13115 6308 13161
rect 6262 13021 6308 13067
rect 6262 12927 6308 12973
rect 6262 12833 6308 12879
rect 8518 13397 8564 13443
rect 8518 13303 8564 13349
rect 8518 13209 8564 13255
rect 8518 13115 8564 13161
rect 8518 13021 8564 13067
rect 8518 12927 8564 12973
rect 6262 12739 6308 12785
rect 6262 12645 6308 12691
rect 6262 12551 6308 12597
rect 8518 12833 8564 12879
rect 8518 12739 8564 12785
rect 8518 12645 8564 12691
rect 6262 12448 6308 12503
rect 6262 12354 6308 12400
rect 6262 12260 6308 12306
rect 6262 12166 6308 12212
rect 6262 12072 6308 12118
rect 6262 11978 6308 12024
rect 8518 12551 8564 12597
rect 8518 12448 8564 12503
rect 8518 12354 8564 12400
rect 8518 12260 8564 12306
rect 8518 12166 8564 12212
rect 8518 12072 8564 12118
rect 8518 11978 8564 12024
rect 6262 11884 6308 11930
rect 6262 11790 6308 11836
rect 6262 11696 6308 11742
rect 8518 11884 8564 11930
rect 8518 11790 8564 11836
rect 18136 13722 18182 13768
rect 18230 13722 18276 13768
rect 18324 13722 18370 13768
rect 18418 13722 18464 13768
rect 18512 13722 18558 13768
rect 18606 13722 18652 13768
rect 18700 13722 18746 13768
rect 18794 13722 18840 13768
rect 18888 13722 18934 13768
rect 18982 13722 19028 13768
rect 19076 13722 19122 13768
rect 19170 13722 19216 13768
rect 19264 13722 19310 13768
rect 19358 13722 19404 13768
rect 19452 13722 19498 13768
rect 19546 13722 19592 13768
rect 19640 13722 19686 13768
rect 19734 13722 19780 13768
rect 19828 13722 19874 13768
rect 19922 13722 19968 13768
rect 20016 13722 20062 13768
rect 20110 13722 20156 13768
rect 20204 13722 20250 13768
rect 20298 13722 20344 13768
rect 20392 13722 20438 13768
rect 20486 13722 20532 13768
rect 20580 13722 20626 13768
rect 20674 13722 20720 13768
rect 20768 13722 20814 13768
rect 20862 13722 20908 13768
rect 20956 13722 21002 13768
rect 21050 13722 21096 13768
rect 21144 13722 21190 13768
rect 18136 13628 18182 13674
rect 18136 13534 18182 13580
rect 18136 13440 18182 13486
rect 21144 13628 21190 13674
rect 21144 13534 21190 13580
rect 21144 13440 21190 13486
rect 18136 13346 18182 13392
rect 21144 13346 21190 13392
rect 18136 13252 18182 13298
rect 18136 13158 18182 13204
rect 21144 13252 21190 13298
rect 18136 13064 18182 13110
rect 18136 12970 18182 13016
rect 18136 12876 18182 12922
rect 18136 12782 18182 12828
rect 18136 12688 18182 12734
rect 18136 12594 18182 12640
rect 21144 13158 21190 13204
rect 21144 13064 21190 13110
rect 21144 12970 21190 13016
rect 21144 12876 21190 12922
rect 21144 12782 21190 12828
rect 21144 12688 21190 12734
rect 21144 12594 21190 12640
rect 18136 12500 18182 12546
rect 18136 12406 18182 12452
rect 21144 12500 21190 12546
rect 18136 12312 18182 12358
rect 18136 12218 18182 12264
rect 21144 12406 21190 12452
rect 21144 12312 21190 12358
rect 18136 12124 18182 12170
rect 18136 12030 18182 12076
rect 18136 11936 18182 11982
rect 18136 11842 18182 11888
rect 8518 11696 8564 11742
rect 6262 11602 6308 11648
rect 6262 11508 6308 11554
rect 6262 11414 6308 11460
rect 6262 11320 6308 11366
rect 6262 11226 6308 11272
rect 6262 11132 6308 11178
rect 8518 11602 8564 11648
rect 8518 11508 8564 11554
rect 8518 11414 8564 11460
rect 8518 11320 8564 11366
rect 8518 11226 8564 11272
rect 8518 11132 8564 11178
rect 8612 11132 8658 11178
rect 8706 11132 8752 11178
rect 8800 11132 8846 11178
rect 8894 11132 8940 11178
rect 8988 11132 9034 11178
rect 9082 11132 9128 11178
rect 9176 11132 9222 11178
rect 9270 11132 9316 11178
rect 9364 11132 9410 11178
rect 9458 11132 9504 11178
rect 9552 11132 9598 11178
rect 9646 11132 9692 11178
rect 9740 11132 9786 11178
rect 9834 11132 9880 11178
rect 9928 11132 9974 11178
rect 10022 11132 10068 11178
rect 10116 11132 10162 11178
rect 10210 11132 10256 11178
rect 10304 11132 10350 11178
rect 10398 11132 10444 11178
rect 10492 11132 10538 11178
rect 10586 11132 10632 11178
rect 10680 11132 10726 11178
rect 10774 11132 10820 11178
rect 10868 11132 10914 11178
rect 10962 11132 11008 11178
rect 11056 11132 11102 11178
rect 11150 11132 11196 11178
rect 11244 11132 11290 11178
rect 6262 11038 6308 11084
rect 6262 10944 6308 10990
rect 6262 10850 6308 10896
rect 8518 11038 8564 11084
rect 8518 10944 8564 10990
rect 8518 10850 8564 10896
rect 11244 11038 11290 11084
rect 11244 10944 11290 10990
rect 6262 10756 6308 10802
rect 6262 10662 6308 10708
rect 6262 10568 6308 10614
rect 6262 10474 6308 10520
rect 6262 10380 6308 10426
rect 6262 10286 6308 10332
rect 11244 10850 11290 10896
rect 8518 10756 8564 10802
rect 8518 10662 8564 10708
rect 8518 10568 8564 10614
rect 8518 10474 8564 10520
rect 8518 10380 8564 10426
rect 8518 10286 8564 10332
rect 6262 10192 6308 10238
rect 6262 10098 6308 10144
rect 6262 10004 6308 10050
rect 8518 10192 8564 10238
rect 11244 10756 11290 10802
rect 11244 10662 11290 10708
rect 11244 10568 11290 10614
rect 11244 10474 11290 10520
rect 11244 10380 11290 10426
rect 11244 10286 11290 10332
rect 8518 10098 8564 10144
rect 8518 10004 8564 10050
rect 6262 9910 6308 9956
rect 6262 9816 6308 9862
rect 6262 9722 6308 9768
rect 6262 9628 6308 9674
rect 6262 9534 6308 9580
rect 6262 9440 6308 9486
rect 6262 9346 6308 9392
rect 8518 9910 8564 9956
rect 11244 10192 11290 10238
rect 11244 10098 11290 10144
rect 11244 10004 11290 10050
rect 8518 9816 8564 9862
rect 8518 9722 8564 9768
rect 8518 9628 8564 9674
rect 8518 9534 8564 9580
rect 8518 9440 8564 9486
rect 6262 9252 6308 9298
rect 6262 9158 6308 9204
rect 6262 9064 6308 9110
rect 8518 9346 8564 9392
rect 11244 9910 11290 9956
rect 11244 9816 11290 9862
rect 11244 9722 11290 9768
rect 11244 9628 11290 9674
rect 11244 9534 11290 9580
rect 11244 9440 11290 9486
rect 8518 9252 8564 9298
rect 8518 9158 8564 9204
rect 6262 8970 6308 9016
rect 6262 8876 6308 8922
rect 6262 8782 6308 8828
rect 6262 8688 6308 8734
rect 6262 8594 6308 8640
rect 6262 8500 6308 8546
rect 8518 9064 8564 9110
rect 11244 9346 11290 9392
rect 11244 9252 11290 9298
rect 11244 9158 11290 9204
rect 8518 8970 8564 9016
rect 8518 8876 8564 8922
rect 8518 8782 8564 8828
rect 8518 8688 8564 8734
rect 8518 8594 8564 8640
rect 6262 8406 6308 8452
rect 6262 8312 6308 8358
rect 8518 8500 8564 8546
rect 11244 9064 11290 9110
rect 11244 8970 11290 9016
rect 11244 8876 11290 8922
rect 11244 8782 11290 8828
rect 11244 8688 11290 8734
rect 11244 8594 11290 8640
rect 6262 8218 6308 8264
rect 8518 8406 8564 8452
rect 8518 8312 8564 8358
rect 11244 8500 11290 8546
rect 11244 8406 11290 8452
rect 6262 8124 6308 8170
rect 6262 8030 6308 8076
rect 6262 7936 6308 7982
rect 6262 7842 6308 7888
rect 6262 7748 6308 7794
rect 6262 7654 6308 7700
rect 8518 8218 8564 8264
rect 11244 8312 11290 8358
rect 8518 8124 8564 8170
rect 8518 8030 8564 8076
rect 8518 7936 8564 7982
rect 8518 7842 8564 7888
rect 8518 7748 8564 7794
rect 8518 7654 8564 7700
rect 6262 7560 6308 7606
rect 6262 7466 6308 7512
rect 6262 7372 6308 7418
rect 11244 8218 11290 8264
rect 11244 8124 11290 8170
rect 11244 8030 11290 8076
rect 11244 7936 11290 7982
rect 11244 7842 11290 7888
rect 11244 7748 11290 7794
rect 11244 7654 11290 7700
rect 8518 7560 8564 7606
rect 8518 7466 8564 7512
rect 8518 7372 8564 7418
rect 11244 7560 11290 7606
rect 11244 7466 11290 7512
rect 11244 7372 11290 7418
rect 6262 7278 6308 7324
rect 6356 7278 6402 7324
rect 6450 7278 6496 7324
rect 6544 7278 6590 7324
rect 6638 7278 6684 7324
rect 6732 7278 6778 7324
rect 6826 7278 6872 7324
rect 6920 7278 6966 7324
rect 7014 7278 7060 7324
rect 7108 7278 7154 7324
rect 7202 7278 7248 7324
rect 7296 7278 7342 7324
rect 7390 7278 7436 7324
rect 7484 7278 7530 7324
rect 7578 7278 7624 7324
rect 7672 7278 7718 7324
rect 7766 7278 7812 7324
rect 7860 7278 7906 7324
rect 7954 7278 8000 7324
rect 8048 7278 8094 7324
rect 8142 7278 8188 7324
rect 8236 7278 8282 7324
rect 8330 7278 8376 7324
rect 8424 7278 8470 7324
rect 8518 7278 8564 7324
rect 8612 7278 8658 7324
rect 8706 7278 8752 7324
rect 8800 7278 8846 7324
rect 8894 7278 8940 7324
rect 8988 7278 9034 7324
rect 9082 7278 9128 7324
rect 9176 7278 9222 7324
rect 9270 7278 9316 7324
rect 9364 7278 9410 7324
rect 9458 7278 9504 7324
rect 9552 7278 9598 7324
rect 9646 7278 9692 7324
rect 9740 7278 9786 7324
rect 9834 7278 9880 7324
rect 9928 7278 9974 7324
rect 10022 7278 10068 7324
rect 10116 7278 10162 7324
rect 10210 7278 10256 7324
rect 10304 7278 10350 7324
rect 10398 7278 10444 7324
rect 10492 7278 10538 7324
rect 10586 7278 10632 7324
rect 10680 7278 10726 7324
rect 10774 7278 10820 7324
rect 10868 7278 10914 7324
rect 10962 7278 11008 7324
rect 11056 7278 11102 7324
rect 11150 7278 11196 7324
rect 11244 7278 11290 7324
rect 18136 11748 18182 11794
rect 18136 11654 18182 11700
rect 21144 12218 21190 12264
rect 21144 12124 21190 12170
rect 21144 12030 21190 12076
rect 21144 11936 21190 11982
rect 21144 11842 21190 11888
rect 21144 11748 21190 11794
rect 21144 11654 21190 11700
rect 18136 11560 18182 11606
rect 18136 11466 18182 11512
rect 18136 11372 18182 11418
rect 18136 11278 18182 11324
rect 21144 11560 21190 11606
rect 21144 11466 21190 11512
rect 21144 11372 21190 11418
rect 18136 11184 18182 11230
rect 18136 11090 18182 11136
rect 18136 10996 18182 11042
rect 18136 10902 18182 10948
rect 18136 10808 18182 10854
rect 18136 10714 18182 10760
rect 21144 11278 21190 11324
rect 21144 11184 21190 11230
rect 21144 11090 21190 11136
rect 21144 10996 21190 11042
rect 21144 10902 21190 10948
rect 21144 10808 21190 10854
rect 18136 10620 18182 10666
rect 18136 10526 18182 10572
rect 18136 10432 18182 10478
rect 18136 10338 18182 10384
rect 21144 10714 21190 10760
rect 21144 10620 21190 10666
rect 21144 10526 21190 10572
rect 21144 10432 21190 10478
rect 18136 10244 18182 10290
rect 18136 10150 18182 10196
rect 18136 10056 18182 10102
rect 18136 9962 18182 10008
rect 18136 9868 18182 9914
rect 18136 9774 18182 9820
rect 21144 10338 21190 10384
rect 21144 10244 21190 10290
rect 21144 10150 21190 10196
rect 21144 10056 21190 10102
rect 21144 9962 21190 10008
rect 21144 9868 21190 9914
rect 18136 9680 18182 9726
rect 18136 9586 18182 9632
rect 18136 9492 18182 9538
rect 21144 9774 21190 9820
rect 21144 9680 21190 9726
rect 21144 9586 21190 9632
rect 21144 9492 21190 9538
rect 18136 9398 18182 9444
rect 18136 9304 18182 9350
rect 18136 9210 18182 9256
rect 18136 9116 18182 9162
rect 18136 9022 18182 9068
rect 18136 8928 18182 8974
rect 18136 8834 18182 8880
rect 21144 9398 21190 9444
rect 21144 9304 21190 9350
rect 21144 9210 21190 9256
rect 21144 9116 21190 9162
rect 21144 9022 21190 9068
rect 21144 8928 21190 8974
rect 18136 8740 18182 8786
rect 18136 8646 18182 8692
rect 21144 8834 21190 8880
rect 21144 8740 21190 8786
rect 18136 8552 18182 8598
rect 21144 8646 21190 8692
rect 21144 8552 21190 8598
rect 18136 8458 18182 8504
rect 18136 8364 18182 8410
rect 18136 8270 18182 8316
rect 18136 8176 18182 8222
rect 18136 8082 18182 8128
rect 18136 7988 18182 8034
rect 18136 7894 18182 7940
rect 21144 8458 21190 8504
rect 21144 8364 21190 8410
rect 21144 8270 21190 8316
rect 21144 8176 21190 8222
rect 21144 8082 21190 8128
rect 21144 7988 21190 8034
rect 18136 7800 18182 7846
rect 21144 7894 21190 7940
rect 21144 7800 21190 7846
rect 18136 7706 18182 7752
rect 21144 7706 21190 7752
rect 18136 7612 18182 7658
rect 18136 7518 18182 7564
rect 18136 7424 18182 7470
rect 21144 7612 21190 7658
rect 21144 7518 21190 7564
rect 21144 7424 21190 7470
rect 18136 7330 18182 7376
rect 18230 7330 18276 7376
rect 18324 7330 18370 7376
rect 18418 7330 18464 7376
rect 18512 7330 18558 7376
rect 18606 7330 18652 7376
rect 18700 7330 18746 7376
rect 18794 7330 18840 7376
rect 18888 7330 18934 7376
rect 18982 7330 19028 7376
rect 19076 7330 19122 7376
rect 19170 7330 19216 7376
rect 19264 7330 19310 7376
rect 19358 7330 19404 7376
rect 19452 7330 19498 7376
rect 19546 7330 19592 7376
rect 19640 7330 19686 7376
rect 19734 7330 19780 7376
rect 19828 7330 19874 7376
rect 19922 7330 19968 7376
rect 20016 7330 20062 7376
rect 20110 7330 20156 7376
rect 20204 7330 20250 7376
rect 20298 7330 20344 7376
rect 20392 7330 20438 7376
rect 20486 7330 20532 7376
rect 20580 7330 20626 7376
rect 20674 7330 20720 7376
rect 20768 7330 20814 7376
rect 20862 7330 20908 7376
rect 20956 7330 21002 7376
rect 21050 7330 21096 7376
rect 21144 7330 21190 7376
rect 23288 13722 23334 13768
rect 23382 13722 23428 13768
rect 23476 13722 23522 13768
rect 23570 13722 23616 13768
rect 23664 13722 23710 13768
rect 23758 13722 23804 13768
rect 23852 13722 23898 13768
rect 23946 13722 23992 13768
rect 24040 13722 24086 13768
rect 24134 13722 24180 13768
rect 24228 13722 24274 13768
rect 24322 13722 24368 13768
rect 24416 13722 24462 13768
rect 24510 13722 24556 13768
rect 24604 13722 24650 13768
rect 24698 13722 24744 13768
rect 24792 13722 24838 13768
rect 24886 13722 24932 13768
rect 24980 13722 25026 13768
rect 25074 13722 25120 13768
rect 25168 13722 25214 13768
rect 25262 13722 25308 13768
rect 25356 13722 25402 13768
rect 25450 13722 25496 13768
rect 25544 13722 25590 13768
rect 25638 13722 25684 13768
rect 25732 13722 25778 13768
rect 25826 13722 25872 13768
rect 25920 13722 25966 13768
rect 26014 13722 26060 13768
rect 26108 13722 26154 13768
rect 26202 13722 26248 13768
rect 26296 13722 26342 13768
rect 23288 13628 23334 13674
rect 23288 13534 23334 13580
rect 23288 13440 23334 13486
rect 26296 13628 26342 13674
rect 26296 13534 26342 13580
rect 26296 13440 26342 13486
rect 23288 13346 23334 13392
rect 26296 13346 26342 13392
rect 23288 13252 23334 13298
rect 23288 13158 23334 13204
rect 26296 13252 26342 13298
rect 23288 13064 23334 13110
rect 23288 12970 23334 13016
rect 23288 12876 23334 12922
rect 23288 12782 23334 12828
rect 23288 12688 23334 12734
rect 23288 12594 23334 12640
rect 26296 13158 26342 13204
rect 26296 13064 26342 13110
rect 26296 12970 26342 13016
rect 26296 12876 26342 12922
rect 26296 12782 26342 12828
rect 26296 12688 26342 12734
rect 26296 12594 26342 12640
rect 23288 12500 23334 12546
rect 23288 12406 23334 12452
rect 26296 12500 26342 12546
rect 23288 12312 23334 12358
rect 23288 12218 23334 12264
rect 26296 12406 26342 12452
rect 26296 12312 26342 12358
rect 23288 12124 23334 12170
rect 23288 12030 23334 12076
rect 23288 11936 23334 11982
rect 23288 11842 23334 11888
rect 23288 11748 23334 11794
rect 23288 11654 23334 11700
rect 26296 12218 26342 12264
rect 26296 12124 26342 12170
rect 26296 12030 26342 12076
rect 26296 11936 26342 11982
rect 26296 11842 26342 11888
rect 26296 11748 26342 11794
rect 26296 11654 26342 11700
rect 23288 11560 23334 11606
rect 23288 11466 23334 11512
rect 23288 11372 23334 11418
rect 23288 11278 23334 11324
rect 26296 11560 26342 11606
rect 26296 11466 26342 11512
rect 26296 11372 26342 11418
rect 23288 11184 23334 11230
rect 23288 11090 23334 11136
rect 23288 10996 23334 11042
rect 23288 10902 23334 10948
rect 23288 10808 23334 10854
rect 23288 10714 23334 10760
rect 26296 11278 26342 11324
rect 26296 11184 26342 11230
rect 26296 11090 26342 11136
rect 26296 10996 26342 11042
rect 26296 10902 26342 10948
rect 26296 10808 26342 10854
rect 23288 10620 23334 10666
rect 23288 10526 23334 10572
rect 23288 10432 23334 10478
rect 23288 10338 23334 10384
rect 26296 10714 26342 10760
rect 26296 10620 26342 10666
rect 26296 10526 26342 10572
rect 26296 10432 26342 10478
rect 23288 10244 23334 10290
rect 23288 10150 23334 10196
rect 23288 10056 23334 10102
rect 23288 9962 23334 10008
rect 23288 9868 23334 9914
rect 23288 9774 23334 9820
rect 26296 10338 26342 10384
rect 26296 10244 26342 10290
rect 26296 10150 26342 10196
rect 26296 10056 26342 10102
rect 26296 9962 26342 10008
rect 26296 9868 26342 9914
rect 23288 9680 23334 9726
rect 23288 9586 23334 9632
rect 23288 9492 23334 9538
rect 26296 9774 26342 9820
rect 26296 9680 26342 9726
rect 26296 9586 26342 9632
rect 26296 9492 26342 9538
rect 23288 9398 23334 9444
rect 23288 9304 23334 9350
rect 23288 9210 23334 9256
rect 23288 9116 23334 9162
rect 23288 9022 23334 9068
rect 23288 8928 23334 8974
rect 23288 8834 23334 8880
rect 26296 9398 26342 9444
rect 26296 9304 26342 9350
rect 26296 9210 26342 9256
rect 26296 9116 26342 9162
rect 26296 9022 26342 9068
rect 26296 8928 26342 8974
rect 23288 8740 23334 8786
rect 23288 8646 23334 8692
rect 26296 8834 26342 8880
rect 26296 8740 26342 8786
rect 23288 8552 23334 8598
rect 26296 8646 26342 8692
rect 26296 8552 26342 8598
rect 23288 8458 23334 8504
rect 23288 8364 23334 8410
rect 23288 8270 23334 8316
rect 23288 8176 23334 8222
rect 23288 8082 23334 8128
rect 23288 7988 23334 8034
rect 23288 7894 23334 7940
rect 26296 8458 26342 8504
rect 26296 8364 26342 8410
rect 26296 8270 26342 8316
rect 26296 8176 26342 8222
rect 26296 8082 26342 8128
rect 26296 7988 26342 8034
rect 23288 7800 23334 7846
rect 26296 7894 26342 7940
rect 26296 7800 26342 7846
rect 23288 7706 23334 7752
rect 26296 7706 26342 7752
rect 23288 7612 23334 7658
rect 23288 7518 23334 7564
rect 23288 7424 23334 7470
rect 26296 7612 26342 7658
rect 26296 7518 26342 7564
rect 26296 7424 26342 7470
rect 23288 7330 23334 7376
rect 23382 7330 23428 7376
rect 23476 7330 23522 7376
rect 23570 7330 23616 7376
rect 23664 7330 23710 7376
rect 23758 7330 23804 7376
rect 23852 7330 23898 7376
rect 23946 7330 23992 7376
rect 24040 7330 24086 7376
rect 24134 7330 24180 7376
rect 24228 7330 24274 7376
rect 24322 7330 24368 7376
rect 24416 7330 24462 7376
rect 24510 7330 24556 7376
rect 24604 7330 24650 7376
rect 24698 7330 24744 7376
rect 24792 7330 24838 7376
rect 24886 7330 24932 7376
rect 24980 7330 25026 7376
rect 25074 7330 25120 7376
rect 25168 7330 25214 7376
rect 25262 7330 25308 7376
rect 25356 7330 25402 7376
rect 25450 7330 25496 7376
rect 25544 7330 25590 7376
rect 25638 7330 25684 7376
rect 25732 7330 25778 7376
rect 25826 7330 25872 7376
rect 25920 7330 25966 7376
rect 26014 7330 26060 7376
rect 26108 7330 26154 7376
rect 26202 7330 26248 7376
rect 26296 7330 26342 7376
rect 27257 13722 27303 13768
rect 27351 13722 27397 13768
rect 27445 13722 27491 13768
rect 27539 13722 27585 13768
rect 27633 13722 27679 13768
rect 27727 13722 27773 13768
rect 27821 13722 27867 13768
rect 27915 13722 27961 13768
rect 28009 13722 28055 13768
rect 28103 13722 28149 13768
rect 28197 13722 28243 13768
rect 28291 13722 28337 13768
rect 28385 13722 28431 13768
rect 28479 13722 28525 13768
rect 28573 13722 28619 13768
rect 28667 13722 28713 13768
rect 28761 13722 28807 13768
rect 28855 13722 28901 13768
rect 28949 13722 28995 13768
rect 29043 13722 29089 13768
rect 29137 13722 29183 13768
rect 29231 13722 29277 13768
rect 29325 13722 29371 13768
rect 29419 13722 29465 13768
rect 29513 13722 29559 13768
rect 29607 13722 29653 13768
rect 29701 13722 29747 13768
rect 29795 13722 29841 13768
rect 29889 13722 29935 13768
rect 29983 13722 30029 13768
rect 30077 13722 30123 13768
rect 30171 13722 30217 13768
rect 30265 13722 30311 13768
rect 27257 13628 27303 13674
rect 27257 13534 27303 13580
rect 27257 13440 27303 13486
rect 30265 13628 30311 13674
rect 30265 13534 30311 13580
rect 30265 13440 30311 13486
rect 27257 13346 27303 13392
rect 30265 13346 30311 13392
rect 27257 13252 27303 13298
rect 27257 13158 27303 13204
rect 30265 13252 30311 13298
rect 27257 13064 27303 13110
rect 27257 12970 27303 13016
rect 27257 12876 27303 12922
rect 27257 12782 27303 12828
rect 27257 12688 27303 12734
rect 27257 12594 27303 12640
rect 30265 13158 30311 13204
rect 30265 13064 30311 13110
rect 30265 12970 30311 13016
rect 30265 12876 30311 12922
rect 30265 12782 30311 12828
rect 30265 12688 30311 12734
rect 30265 12594 30311 12640
rect 27257 12500 27303 12546
rect 27257 12406 27303 12452
rect 30265 12500 30311 12546
rect 27257 12312 27303 12358
rect 27257 12218 27303 12264
rect 30265 12406 30311 12452
rect 30265 12312 30311 12358
rect 27257 12124 27303 12170
rect 27257 12030 27303 12076
rect 27257 11936 27303 11982
rect 27257 11842 27303 11888
rect 27257 11748 27303 11794
rect 27257 11654 27303 11700
rect 30265 12218 30311 12264
rect 30265 12124 30311 12170
rect 30265 12030 30311 12076
rect 30265 11936 30311 11982
rect 30265 11842 30311 11888
rect 30265 11748 30311 11794
rect 30265 11654 30311 11700
rect 27257 11560 27303 11606
rect 27257 11466 27303 11512
rect 27257 11372 27303 11418
rect 27257 11278 27303 11324
rect 30265 11560 30311 11606
rect 30265 11466 30311 11512
rect 30265 11372 30311 11418
rect 27257 11184 27303 11230
rect 27257 11090 27303 11136
rect 27257 10996 27303 11042
rect 27257 10902 27303 10948
rect 27257 10808 27303 10854
rect 27257 10714 27303 10760
rect 30265 11278 30311 11324
rect 30265 11184 30311 11230
rect 30265 11090 30311 11136
rect 30265 10996 30311 11042
rect 30265 10902 30311 10948
rect 30265 10808 30311 10854
rect 27257 10620 27303 10666
rect 27257 10526 27303 10572
rect 27257 10432 27303 10478
rect 27257 10338 27303 10384
rect 30265 10714 30311 10760
rect 30265 10620 30311 10666
rect 30265 10526 30311 10572
rect 30265 10432 30311 10478
rect 27257 10244 27303 10290
rect 27257 10150 27303 10196
rect 27257 10056 27303 10102
rect 27257 9962 27303 10008
rect 27257 9868 27303 9914
rect 27257 9774 27303 9820
rect 30265 10338 30311 10384
rect 30265 10244 30311 10290
rect 30265 10150 30311 10196
rect 30265 10056 30311 10102
rect 30265 9962 30311 10008
rect 30265 9868 30311 9914
rect 27257 9680 27303 9726
rect 27257 9586 27303 9632
rect 27257 9492 27303 9538
rect 30265 9774 30311 9820
rect 30265 9680 30311 9726
rect 30265 9586 30311 9632
rect 30265 9492 30311 9538
rect 27257 9398 27303 9444
rect 27257 9304 27303 9350
rect 27257 9210 27303 9256
rect 27257 9116 27303 9162
rect 27257 9022 27303 9068
rect 27257 8928 27303 8974
rect 27257 8834 27303 8880
rect 30265 9398 30311 9444
rect 30265 9304 30311 9350
rect 30265 9210 30311 9256
rect 30265 9116 30311 9162
rect 30265 9022 30311 9068
rect 30265 8928 30311 8974
rect 27257 8740 27303 8786
rect 27257 8646 27303 8692
rect 30265 8834 30311 8880
rect 30265 8740 30311 8786
rect 27257 8552 27303 8598
rect 30265 8646 30311 8692
rect 30265 8552 30311 8598
rect 27257 8458 27303 8504
rect 27257 8364 27303 8410
rect 27257 8270 27303 8316
rect 27257 8176 27303 8222
rect 27257 8082 27303 8128
rect 27257 7988 27303 8034
rect 27257 7894 27303 7940
rect 30265 8458 30311 8504
rect 30265 8364 30311 8410
rect 30265 8270 30311 8316
rect 30265 8176 30311 8222
rect 30265 8082 30311 8128
rect 30265 7988 30311 8034
rect 27257 7800 27303 7846
rect 30265 7894 30311 7940
rect 30265 7800 30311 7846
rect 27257 7706 27303 7752
rect 30265 7706 30311 7752
rect 27257 7612 27303 7658
rect 27257 7518 27303 7564
rect 27257 7424 27303 7470
rect 30265 7612 30311 7658
rect 30265 7518 30311 7564
rect 30265 7424 30311 7470
rect 27257 7330 27303 7376
rect 27351 7330 27397 7376
rect 27445 7330 27491 7376
rect 27539 7330 27585 7376
rect 27633 7330 27679 7376
rect 27727 7330 27773 7376
rect 27821 7330 27867 7376
rect 27915 7330 27961 7376
rect 28009 7330 28055 7376
rect 28103 7330 28149 7376
rect 28197 7330 28243 7376
rect 28291 7330 28337 7376
rect 28385 7330 28431 7376
rect 28479 7330 28525 7376
rect 28573 7330 28619 7376
rect 28667 7330 28713 7376
rect 28761 7330 28807 7376
rect 28855 7330 28901 7376
rect 28949 7330 28995 7376
rect 29043 7330 29089 7376
rect 29137 7330 29183 7376
rect 29231 7330 29277 7376
rect 29325 7330 29371 7376
rect 29419 7330 29465 7376
rect 29513 7330 29559 7376
rect 29607 7330 29653 7376
rect 29701 7330 29747 7376
rect 29795 7330 29841 7376
rect 29889 7330 29935 7376
rect 29983 7330 30029 7376
rect 30077 7330 30123 7376
rect 30171 7330 30217 7376
rect 30265 7330 30311 7376
rect 6934 6072 6980 6118
rect 7028 6072 7074 6118
rect 7122 6072 7168 6118
rect 7216 6072 7262 6118
rect 7310 6072 7356 6118
rect 7404 6072 7450 6118
rect 7498 6072 7544 6118
rect 7592 6072 7638 6118
rect 7686 6072 7732 6118
rect 7780 6072 7826 6118
rect 7874 6072 7920 6118
rect 7968 6072 8014 6118
rect 8062 6072 8108 6118
rect 8156 6072 8202 6118
rect 8250 6072 8296 6118
rect 8344 6072 8390 6118
rect 8438 6072 8484 6118
rect 8532 6072 8578 6118
rect 8626 6072 8672 6118
rect 8720 6072 8766 6118
rect 8814 6072 8860 6118
rect 8908 6072 8954 6118
rect 9002 6072 9048 6118
rect 9096 6072 9142 6118
rect 9190 6072 9236 6118
rect 9284 6072 9330 6118
rect 9378 6072 9424 6118
rect 9472 6072 9518 6118
rect 9566 6072 9612 6118
rect 9660 6072 9706 6118
rect 9754 6072 9800 6118
rect 9848 6072 9894 6118
rect 9942 6072 9988 6118
rect 10036 6072 10082 6118
rect 6934 5978 6980 6024
rect 10036 5978 10082 6024
rect 6934 5884 6980 5930
rect 6934 5790 6980 5836
rect 6934 5696 6980 5742
rect 10036 5884 10082 5930
rect 10036 5790 10082 5836
rect 6934 5602 6980 5648
rect 6934 5508 6980 5554
rect 10036 5696 10082 5742
rect 10036 5602 10082 5648
rect 6934 5414 6980 5460
rect 6934 5320 6980 5366
rect 6934 5226 6980 5272
rect 10036 5508 10082 5554
rect 10036 5414 10082 5460
rect 10036 5320 10082 5366
rect 10036 5226 10082 5272
rect 6934 5132 6980 5178
rect 6934 5038 6980 5084
rect 10036 5132 10082 5178
rect 10036 5038 10082 5084
rect 6934 4944 6980 4990
rect 6934 4850 6980 4896
rect 6934 4756 6980 4802
rect 6934 4662 6980 4708
rect 10036 4944 10082 4990
rect 10036 4850 10082 4896
rect 10036 4756 10082 4802
rect 6934 4568 6980 4614
rect 6934 4474 6980 4520
rect 10036 4662 10082 4708
rect 10036 4568 10082 4614
rect 10036 4474 10082 4520
rect 6934 4380 6980 4426
rect 6934 4286 6980 4332
rect 6934 4192 6980 4238
rect 6934 4098 6980 4144
rect 10036 4380 10082 4426
rect 10036 4286 10082 4332
rect 10036 4192 10082 4238
rect 6934 4004 6980 4050
rect 6934 3910 6980 3956
rect 10036 4098 10082 4144
rect 10036 4004 10082 4050
rect 6934 3816 6980 3862
rect 6934 3722 6980 3768
rect 6934 3628 6980 3674
rect 10036 3910 10082 3956
rect 10036 3816 10082 3862
rect 10036 3722 10082 3768
rect 10036 3628 10082 3674
rect 6934 3534 6980 3580
rect 6934 3440 6980 3486
rect 10036 3534 10082 3580
rect 10036 3440 10082 3486
rect 6934 3346 6980 3392
rect 6934 3252 6980 3298
rect 6934 3158 6980 3204
rect 6934 3064 6980 3110
rect 10036 3346 10082 3392
rect 10036 3252 10082 3298
rect 10036 3158 10082 3204
rect 10036 3064 10082 3110
rect 6934 2970 6980 3016
rect 6934 2876 6980 2922
rect 10036 2970 10082 3016
rect 10036 2876 10082 2922
rect 5900 2782 5946 2828
rect 5994 2782 6040 2828
rect 6088 2782 6134 2828
rect 6182 2782 6228 2828
rect 6276 2782 6322 2828
rect 6370 2782 6416 2828
rect 6464 2782 6510 2828
rect 6558 2782 6604 2828
rect 6652 2782 6698 2828
rect 6746 2782 6792 2828
rect 6840 2782 6886 2828
rect 6934 2782 6980 2828
rect 12014 4423 12060 4469
rect 12108 4423 12154 4469
rect 12202 4423 12248 4469
rect 12296 4423 12342 4469
rect 12390 4423 12436 4469
rect 12484 4423 12530 4469
rect 12578 4423 12624 4469
rect 12672 4423 12718 4469
rect 12766 4423 12812 4469
rect 12860 4423 12906 4469
rect 12954 4423 13000 4469
rect 13048 4423 13094 4469
rect 13142 4423 13188 4469
rect 13236 4423 13282 4469
rect 13330 4423 13376 4469
rect 13424 4423 13470 4469
rect 13518 4423 13564 4469
rect 13612 4423 13658 4469
rect 13706 4423 13752 4469
rect 13800 4423 13846 4469
rect 13894 4423 13940 4469
rect 13988 4423 14034 4469
rect 14082 4423 14128 4469
rect 14176 4423 14222 4469
rect 14270 4423 14316 4469
rect 14364 4423 14410 4469
rect 14458 4423 14504 4469
rect 14552 4423 14598 4469
rect 14646 4423 14692 4469
rect 14740 4423 14786 4469
rect 14834 4423 14880 4469
rect 14928 4423 14974 4469
rect 15022 4423 15068 4469
rect 15116 4423 15162 4469
rect 15210 4423 15256 4469
rect 15304 4423 15350 4469
rect 15398 4423 15444 4469
rect 15492 4423 15538 4469
rect 15586 4423 15632 4469
rect 15680 4423 15726 4469
rect 15774 4423 15820 4469
rect 15868 4423 15914 4469
rect 15962 4423 16008 4469
rect 16056 4423 16102 4469
rect 16150 4423 16196 4469
rect 16244 4423 16290 4469
rect 16338 4423 16384 4469
rect 16432 4423 16478 4469
rect 16526 4423 16572 4469
rect 16620 4423 16666 4469
rect 16714 4423 16760 4469
rect 16808 4423 16854 4469
rect 16902 4423 16948 4469
rect 16996 4423 17042 4469
rect 17090 4423 17136 4469
rect 17184 4423 17230 4469
rect 17278 4423 17324 4469
rect 17372 4423 17418 4469
rect 17466 4423 17512 4469
rect 17560 4423 17606 4469
rect 12014 4329 12060 4375
rect 12014 4235 12060 4281
rect 12014 4141 12060 4187
rect 12014 4047 12060 4093
rect 17560 4329 17606 4375
rect 17560 4235 17606 4281
rect 17560 4141 17606 4187
rect 12014 3953 12060 3999
rect 12014 3859 12060 3905
rect 12014 3765 12060 3811
rect 17560 4047 17606 4093
rect 17560 3953 17606 3999
rect 17560 3859 17606 3905
rect 12014 3671 12060 3717
rect 12014 3577 12060 3623
rect 12014 3483 12060 3529
rect 12014 3389 12060 3435
rect 17560 3765 17606 3811
rect 17560 3671 17606 3717
rect 17560 3577 17606 3623
rect 17560 3483 17606 3529
rect 17560 3389 17606 3435
rect 12014 3295 12060 3341
rect 12014 3201 12060 3247
rect 17560 3295 17606 3341
rect 12014 3107 12060 3153
rect 12014 3013 12060 3059
rect 12014 2919 12060 2965
rect 10036 2782 10082 2828
rect 10130 2782 10176 2828
rect 10224 2782 10270 2828
rect 10318 2782 10364 2828
rect 10412 2782 10458 2828
rect 10506 2782 10552 2828
rect 10600 2782 10646 2828
rect 10694 2782 10740 2828
rect 10788 2782 10834 2828
rect 10882 2782 10928 2828
rect 10976 2782 11022 2828
rect 11070 2782 11116 2828
rect 5900 2688 5946 2734
rect 11070 2688 11116 2734
rect 5900 2594 5946 2640
rect 5900 2500 5946 2546
rect 5900 2406 5946 2452
rect 11070 2594 11116 2640
rect 11070 2500 11116 2546
rect 5900 2312 5946 2358
rect 5900 2218 5946 2264
rect 11070 2406 11116 2452
rect 11070 2312 11116 2358
rect 5900 2124 5946 2170
rect 5900 2030 5946 2076
rect 11070 2218 11116 2264
rect 11070 2124 11116 2170
rect 5900 1936 5946 1982
rect 11070 2030 11116 2076
rect 5900 1842 5946 1888
rect 5900 1748 5946 1794
rect 11070 1936 11116 1982
rect 11070 1842 11116 1888
rect 5900 1654 5946 1700
rect 5900 1560 5946 1606
rect 11070 1748 11116 1794
rect 11070 1654 11116 1700
rect 11070 1560 11116 1606
rect 5900 1466 5946 1512
rect 5900 1372 5946 1418
rect 11070 1466 11116 1512
rect 11070 1372 11116 1418
rect 5900 1278 5946 1324
rect 5994 1278 6040 1324
rect 6088 1278 6134 1324
rect 6182 1278 6228 1324
rect 6276 1278 6322 1324
rect 6370 1278 6416 1324
rect 6464 1278 6510 1324
rect 6558 1278 6604 1324
rect 6652 1278 6698 1324
rect 6746 1278 6792 1324
rect 6840 1278 6886 1324
rect 6934 1278 6980 1324
rect 7028 1278 7074 1324
rect 7122 1278 7168 1324
rect 7216 1278 7262 1324
rect 7310 1278 7356 1324
rect 7404 1278 7450 1324
rect 7498 1278 7544 1324
rect 7592 1278 7638 1324
rect 7686 1278 7732 1324
rect 7780 1278 7826 1324
rect 7874 1278 7920 1324
rect 7968 1278 8014 1324
rect 8062 1278 8108 1324
rect 8156 1278 8202 1324
rect 8250 1278 8296 1324
rect 8344 1278 8390 1324
rect 8438 1278 8484 1324
rect 8532 1278 8578 1324
rect 8626 1278 8672 1324
rect 8720 1278 8766 1324
rect 8814 1278 8860 1324
rect 8908 1278 8954 1324
rect 9002 1278 9048 1324
rect 9096 1278 9142 1324
rect 9190 1278 9236 1324
rect 9284 1278 9330 1324
rect 9378 1278 9424 1324
rect 9472 1278 9518 1324
rect 9566 1278 9612 1324
rect 9660 1278 9706 1324
rect 9754 1278 9800 1324
rect 9848 1278 9894 1324
rect 9942 1278 9988 1324
rect 10036 1278 10082 1324
rect 10130 1278 10176 1324
rect 10224 1278 10270 1324
rect 10318 1278 10364 1324
rect 10412 1278 10458 1324
rect 10506 1278 10552 1324
rect 10600 1278 10646 1324
rect 10694 1278 10740 1324
rect 10788 1278 10834 1324
rect 10882 1278 10928 1324
rect 10976 1278 11022 1324
rect 11070 1278 11116 1324
rect 12014 2825 12060 2871
rect 17560 3201 17606 3247
rect 17560 3107 17606 3153
rect 17560 3013 17606 3059
rect 17560 2919 17606 2965
rect 12014 2731 12060 2777
rect 12014 2637 12060 2683
rect 12014 2543 12060 2589
rect 12014 2449 12060 2495
rect 17560 2825 17606 2871
rect 17560 2731 17606 2777
rect 17560 2637 17606 2683
rect 17560 2543 17606 2589
rect 17560 2449 17606 2495
rect 12014 2355 12060 2401
rect 12014 2261 12060 2307
rect 12014 2167 12060 2213
rect 12014 2073 12060 2119
rect 12014 1979 12060 2025
rect 17560 2355 17606 2401
rect 17560 2261 17606 2307
rect 17560 2167 17606 2213
rect 17560 2073 17606 2119
rect 12014 1885 12060 1931
rect 12014 1791 12060 1837
rect 12014 1697 12060 1743
rect 12014 1603 12060 1649
rect 17560 1979 17606 2025
rect 17560 1885 17606 1931
rect 17560 1791 17606 1837
rect 17560 1697 17606 1743
rect 12014 1509 12060 1555
rect 12014 1415 12060 1461
rect 17560 1603 17606 1649
rect 17560 1509 17606 1555
rect 17560 1415 17606 1461
rect 12014 1321 12060 1367
rect 12108 1321 12154 1367
rect 12202 1321 12248 1367
rect 12296 1321 12342 1367
rect 12390 1321 12436 1367
rect 12484 1321 12530 1367
rect 12578 1321 12624 1367
rect 12672 1321 12718 1367
rect 12766 1321 12812 1367
rect 12860 1321 12906 1367
rect 12954 1321 13000 1367
rect 13048 1321 13094 1367
rect 13142 1321 13188 1367
rect 13236 1321 13282 1367
rect 13330 1321 13376 1367
rect 13424 1321 13470 1367
rect 13518 1321 13564 1367
rect 13612 1321 13658 1367
rect 13706 1321 13752 1367
rect 13800 1321 13846 1367
rect 13894 1321 13940 1367
rect 13988 1321 14034 1367
rect 14082 1321 14128 1367
rect 14176 1321 14222 1367
rect 14270 1321 14316 1367
rect 14364 1321 14410 1367
rect 14458 1321 14504 1367
rect 14552 1321 14598 1367
rect 14646 1321 14692 1367
rect 14740 1321 14786 1367
rect 14834 1321 14880 1367
rect 14928 1321 14974 1367
rect 15022 1321 15068 1367
rect 15116 1321 15162 1367
rect 15210 1321 15256 1367
rect 15304 1321 15350 1367
rect 15398 1321 15444 1367
rect 15492 1321 15538 1367
rect 15586 1321 15632 1367
rect 15680 1321 15726 1367
rect 15774 1321 15820 1367
rect 15868 1321 15914 1367
rect 15962 1321 16008 1367
rect 16056 1321 16102 1367
rect 16150 1321 16196 1367
rect 16244 1321 16290 1367
rect 16338 1321 16384 1367
rect 16432 1321 16478 1367
rect 16526 1321 16572 1367
rect 16620 1321 16666 1367
rect 16714 1321 16760 1367
rect 16808 1321 16854 1367
rect 16902 1321 16948 1367
rect 16996 1321 17042 1367
rect 17090 1321 17136 1367
rect 17184 1321 17230 1367
rect 17278 1321 17324 1367
rect 17372 1321 17418 1367
rect 17466 1321 17512 1367
rect 17560 1321 17606 1367
<< nsubdiffcont >>
rect 3444 14328 3490 14374
rect 3538 14328 3584 14374
rect 3632 14328 3678 14374
rect 3726 14328 3772 14374
rect 3820 14328 3866 14374
rect 3914 14328 3960 14374
rect 4008 14328 4054 14374
rect 4102 14328 4148 14374
rect 4196 14328 4242 14374
rect 4290 14328 4336 14374
rect 4384 14328 4430 14374
rect 4478 14328 4524 14374
rect 4572 14328 4618 14374
rect 4666 14328 4712 14374
rect 4760 14328 4806 14374
rect 4854 14328 4900 14374
rect 4948 14328 4994 14374
rect 5042 14328 5088 14374
rect 5136 14328 5182 14374
rect 5230 14328 5276 14374
rect 5324 14328 5370 14374
rect 5418 14328 5464 14374
rect 5512 14328 5558 14374
rect 5606 14328 5652 14374
rect 3444 14234 3490 14280
rect 5606 14234 5652 14280
rect 3444 14140 3490 14186
rect 3444 14046 3490 14092
rect 5606 14140 5652 14186
rect 5606 14046 5652 14092
rect 3444 13952 3490 13998
rect 3444 13858 3490 13904
rect 3444 13764 3490 13810
rect 3444 13670 3490 13716
rect 3444 13576 3490 13622
rect 3444 13482 3490 13528
rect 3444 13388 3490 13434
rect 3444 13294 3490 13340
rect 5606 13952 5652 13998
rect 5606 13858 5652 13904
rect 5606 13764 5652 13810
rect 5606 13670 5652 13716
rect 5606 13576 5652 13622
rect 5606 13482 5652 13528
rect 5606 13388 5652 13434
rect 5606 13294 5652 13340
rect 3444 13200 3490 13246
rect 3444 13106 3490 13152
rect 3444 13012 3490 13058
rect 3444 12918 3490 12964
rect 5606 13200 5652 13246
rect 5606 13106 5652 13152
rect 5606 13012 5652 13058
rect 5606 12918 5652 12964
rect 3444 12824 3490 12870
rect 3444 12730 3490 12776
rect 3444 12636 3490 12682
rect 3444 12542 3490 12588
rect 3444 12448 3490 12494
rect 3444 12354 3490 12400
rect 3444 12260 3490 12306
rect 3444 12166 3490 12212
rect 5606 12824 5652 12870
rect 5606 12730 5652 12776
rect 5606 12636 5652 12682
rect 5606 12542 5652 12588
rect 5606 12448 5652 12494
rect 5606 12354 5652 12400
rect 5606 12260 5652 12306
rect 5606 12166 5652 12212
rect 3444 12072 3490 12118
rect 3444 11978 3490 12024
rect 3444 11884 3490 11930
rect 3444 11790 3490 11836
rect 5606 12072 5652 12118
rect 5606 11978 5652 12024
rect 5606 11884 5652 11930
rect 5606 11790 5652 11836
rect 3444 11696 3490 11742
rect 3444 11602 3490 11648
rect 3444 11508 3490 11554
rect 3444 11414 3490 11460
rect 3444 11320 3490 11366
rect 3444 11226 3490 11272
rect 3444 11132 3490 11178
rect 3444 11038 3490 11084
rect 5606 11696 5652 11742
rect 5606 11602 5652 11648
rect 5606 11508 5652 11554
rect 5606 11414 5652 11460
rect 5606 11320 5652 11366
rect 5606 11226 5652 11272
rect 5606 11132 5652 11178
rect 5606 11038 5652 11084
rect 3444 10944 3490 10990
rect 530 10850 576 10896
rect 624 10850 670 10896
rect 718 10850 764 10896
rect 812 10850 858 10896
rect 906 10850 952 10896
rect 1000 10850 1046 10896
rect 1094 10850 1140 10896
rect 1188 10850 1234 10896
rect 1282 10850 1328 10896
rect 1376 10850 1422 10896
rect 1470 10850 1516 10896
rect 1564 10850 1610 10896
rect 1658 10850 1704 10896
rect 1752 10850 1798 10896
rect 1846 10850 1892 10896
rect 1940 10850 1986 10896
rect 2034 10850 2080 10896
rect 2128 10850 2174 10896
rect 2222 10850 2268 10896
rect 2316 10850 2362 10896
rect 2410 10850 2456 10896
rect 2504 10850 2550 10896
rect 2598 10850 2644 10896
rect 2692 10850 2738 10896
rect 2786 10850 2832 10896
rect 2880 10850 2926 10896
rect 2974 10850 3020 10896
rect 3068 10850 3114 10896
rect 3162 10850 3208 10896
rect 3256 10850 3302 10896
rect 3350 10850 3396 10896
rect 3444 10850 3490 10896
rect 530 10756 576 10802
rect -7703 10602 -7657 10648
rect -7605 10602 -7559 10648
rect -7507 10602 -7461 10648
rect -7409 10602 -7363 10648
rect -7311 10602 -7265 10648
rect -7213 10602 -7167 10648
rect -7115 10602 -7069 10648
rect -7017 10602 -6971 10648
rect -6919 10602 -6873 10648
rect -6821 10602 -6775 10648
rect -6723 10602 -6677 10648
rect -6625 10602 -6579 10648
rect -6527 10602 -6481 10648
rect -6429 10602 -6383 10648
rect -6331 10602 -6285 10648
rect -6233 10602 -6187 10648
rect -6135 10602 -6089 10648
rect -6037 10602 -5991 10648
rect -5939 10602 -5893 10648
rect -5841 10602 -5795 10648
rect -5743 10602 -5697 10648
rect -5645 10602 -5599 10648
rect -5547 10602 -5501 10648
rect -5449 10602 -5403 10648
rect -5351 10602 -5305 10648
rect -5253 10602 -5207 10648
rect -5155 10602 -5109 10648
rect -5057 10602 -5011 10648
rect -4959 10602 -4913 10648
rect -4861 10602 -4815 10648
rect -4763 10602 -4717 10648
rect -4665 10602 -4619 10648
rect -4567 10602 -4521 10648
rect -4469 10602 -4423 10648
rect -4371 10602 -4325 10648
rect -4273 10602 -4227 10648
rect -4175 10602 -4129 10648
rect -4077 10602 -4031 10648
rect -3979 10602 -3933 10648
rect -3872 10602 -3826 10648
rect -7703 10494 -7657 10540
rect -7703 10396 -7657 10442
rect -7703 10298 -7657 10344
rect -7703 10200 -7657 10246
rect -7703 10102 -7657 10148
rect -7703 10004 -7657 10050
rect -7703 9906 -7657 9952
rect -7703 9808 -7657 9854
rect -7703 9710 -7657 9756
rect -7703 9612 -7657 9658
rect -7703 9514 -7657 9560
rect -7703 9416 -7657 9462
rect -7703 9318 -7657 9364
rect -7703 9220 -7657 9266
rect -7703 9122 -7657 9168
rect -7703 9024 -7657 9070
rect -7703 8926 -7657 8972
rect -7703 8828 -7657 8874
rect -7703 8730 -7657 8776
rect -7703 8632 -7657 8678
rect -7703 8534 -7657 8580
rect -7703 8436 -7657 8482
rect -7703 8338 -7657 8384
rect -7703 8240 -7657 8286
rect -7703 8142 -7657 8188
rect -7703 8044 -7657 8090
rect -7703 7946 -7657 7992
rect -7703 7848 -7657 7894
rect -7703 7750 -7657 7796
rect -3872 10494 -3826 10540
rect -3872 10396 -3826 10442
rect -3872 10298 -3826 10344
rect -3872 10200 -3826 10246
rect -3872 10102 -3826 10148
rect -3872 10004 -3826 10050
rect -3872 9906 -3826 9952
rect -3872 9808 -3826 9854
rect -3872 9710 -3826 9756
rect -3872 9612 -3826 9658
rect -3872 9514 -3826 9560
rect -3872 9416 -3826 9462
rect -3872 9318 -3826 9364
rect -3872 9220 -3826 9266
rect -3872 9122 -3826 9168
rect -3872 9024 -3826 9070
rect -3872 8926 -3826 8972
rect -3872 8828 -3826 8874
rect -3872 8730 -3826 8776
rect -3872 8632 -3826 8678
rect -3872 8534 -3826 8580
rect -3872 8436 -3826 8482
rect -3872 8338 -3826 8384
rect -3872 8240 -3826 8286
rect -3872 8142 -3826 8188
rect -3872 8044 -3826 8090
rect -3872 7946 -3826 7992
rect -3872 7848 -3826 7894
rect -3872 7750 -3826 7796
rect -7703 7652 -7657 7698
rect -3872 7652 -3826 7698
rect -7703 7554 -7657 7600
rect -7605 7554 -7559 7600
rect -7507 7554 -7461 7600
rect -7409 7554 -7363 7600
rect -7311 7554 -7265 7600
rect -7213 7554 -7167 7600
rect -7115 7554 -7069 7600
rect -7017 7554 -6971 7600
rect -6919 7554 -6873 7600
rect -6821 7554 -6775 7600
rect -6723 7554 -6677 7600
rect -6625 7554 -6579 7600
rect -6527 7554 -6481 7600
rect -6429 7554 -6383 7600
rect -6331 7554 -6285 7600
rect -6233 7554 -6187 7600
rect -6135 7554 -6089 7600
rect -6037 7554 -5991 7600
rect -5939 7554 -5893 7600
rect -5841 7554 -5795 7600
rect -5743 7554 -5697 7600
rect -5645 7554 -5599 7600
rect -5547 7554 -5501 7600
rect -5449 7554 -5403 7600
rect -5351 7554 -5305 7600
rect -5253 7554 -5207 7600
rect -5155 7554 -5109 7600
rect -5057 7554 -5011 7600
rect -4959 7554 -4913 7600
rect -4861 7554 -4815 7600
rect -4763 7554 -4717 7600
rect -4665 7554 -4619 7600
rect -4567 7554 -4521 7600
rect -4469 7554 -4423 7600
rect -4371 7554 -4325 7600
rect -4273 7554 -4227 7600
rect -4175 7554 -4129 7600
rect -4077 7554 -4031 7600
rect -3979 7554 -3933 7600
rect -3872 7554 -3826 7600
rect 530 10662 576 10708
rect 530 10568 576 10614
rect 3444 10756 3490 10802
rect 3444 10662 3490 10708
rect 5606 10944 5652 10990
rect 5606 10850 5652 10896
rect 5606 10756 5652 10802
rect 5606 10662 5652 10708
rect 3444 10568 3490 10614
rect 530 10474 576 10520
rect 530 10380 576 10426
rect 530 10286 576 10332
rect 530 10192 576 10238
rect 530 10098 576 10144
rect 530 10004 576 10050
rect 530 9910 576 9956
rect 3444 10474 3490 10520
rect 3444 10380 3490 10426
rect 3444 10286 3490 10332
rect 3444 10192 3490 10238
rect 3444 10098 3490 10144
rect 3444 10004 3490 10050
rect 530 9816 576 9862
rect 3444 9910 3490 9956
rect 5606 10568 5652 10614
rect 5606 10474 5652 10520
rect 5606 10380 5652 10426
rect 5606 10286 5652 10332
rect 5606 10192 5652 10238
rect 5606 10098 5652 10144
rect 5606 10004 5652 10050
rect 5606 9910 5652 9956
rect 3444 9816 3490 9862
rect 530 9722 576 9768
rect 530 9628 576 9674
rect 530 9534 576 9580
rect 530 9440 576 9486
rect 530 9346 576 9392
rect 530 9252 576 9298
rect 530 9158 576 9204
rect 3444 9722 3490 9768
rect 3444 9628 3490 9674
rect 3444 9534 3490 9580
rect 5606 9816 5652 9862
rect 5606 9722 5652 9768
rect 5606 9628 5652 9674
rect 5606 9534 5652 9580
rect 3444 9440 3490 9486
rect 3444 9346 3490 9392
rect 3444 9252 3490 9298
rect 530 9064 576 9110
rect 3444 9158 3490 9204
rect 3444 9064 3490 9110
rect 530 8970 576 9016
rect 530 8876 576 8922
rect 530 8782 576 8828
rect 530 8688 576 8734
rect 530 8594 576 8640
rect 530 8500 576 8546
rect 530 8406 576 8452
rect 3444 8970 3490 9016
rect 3444 8876 3490 8922
rect 3444 8782 3490 8828
rect 5606 9440 5652 9486
rect 5606 9346 5652 9392
rect 5606 9252 5652 9298
rect 5606 9158 5652 9204
rect 5606 9064 5652 9110
rect 5606 8970 5652 9016
rect 5606 8876 5652 8922
rect 5606 8782 5652 8828
rect 3444 8688 3490 8734
rect 3444 8594 3490 8640
rect 3444 8500 3490 8546
rect 5606 8688 5652 8734
rect 530 8312 576 8358
rect 3444 8406 3490 8452
rect 5606 8594 5652 8640
rect 5606 8500 5652 8546
rect 5606 8406 5652 8452
rect 3444 8312 3490 8358
rect 530 8218 576 8264
rect 530 8124 576 8170
rect 530 8030 576 8076
rect 530 7936 576 7982
rect 530 7842 576 7888
rect 530 7748 576 7794
rect 530 7654 576 7700
rect 3444 8218 3490 8264
rect 3444 8124 3490 8170
rect 3444 8030 3490 8076
rect 3444 7936 3490 7982
rect 3444 7842 3490 7888
rect 3444 7748 3490 7794
rect 3444 7654 3490 7700
rect 530 7560 576 7606
rect 5606 8312 5652 8358
rect 5606 8218 5652 8264
rect 5606 8124 5652 8170
rect 5606 8030 5652 8076
rect 5606 7936 5652 7982
rect 5606 7842 5652 7888
rect 5606 7748 5652 7794
rect 5606 7654 5652 7700
rect 3444 7560 3490 7606
rect 530 7466 576 7512
rect -7703 7392 -7657 7438
rect -7605 7392 -7559 7438
rect -7507 7392 -7461 7438
rect -7409 7392 -7363 7438
rect -7311 7392 -7265 7438
rect -7213 7392 -7167 7438
rect -7115 7392 -7069 7438
rect -7017 7392 -6971 7438
rect -6919 7392 -6873 7438
rect -6821 7392 -6775 7438
rect -6723 7392 -6677 7438
rect -6625 7392 -6579 7438
rect -6527 7392 -6481 7438
rect -6429 7392 -6383 7438
rect -6331 7392 -6285 7438
rect -6233 7392 -6187 7438
rect -6135 7392 -6089 7438
rect -6037 7392 -5991 7438
rect -5939 7392 -5893 7438
rect -5841 7392 -5795 7438
rect -5743 7392 -5697 7438
rect -5645 7392 -5599 7438
rect -5547 7392 -5501 7438
rect -5449 7392 -5403 7438
rect -5351 7392 -5305 7438
rect -5253 7392 -5207 7438
rect -5155 7392 -5109 7438
rect -5057 7392 -5011 7438
rect -4959 7392 -4913 7438
rect -4861 7392 -4815 7438
rect -4763 7392 -4717 7438
rect -4665 7392 -4619 7438
rect -4567 7392 -4521 7438
rect -4469 7392 -4423 7438
rect -4371 7392 -4325 7438
rect -4273 7392 -4227 7438
rect -4175 7392 -4129 7438
rect -4077 7392 -4031 7438
rect -3979 7392 -3933 7438
rect -3872 7392 -3826 7438
rect -7703 7294 -7657 7340
rect -3872 7294 -3826 7340
rect -7703 7196 -7657 7242
rect -7703 7098 -7657 7144
rect -7703 7000 -7657 7046
rect -7703 6902 -7657 6948
rect -7703 6804 -7657 6850
rect -7703 6706 -7657 6752
rect -7703 6608 -7657 6654
rect -7703 6510 -7657 6556
rect -7703 6412 -7657 6458
rect -7703 6314 -7657 6360
rect -7703 6216 -7657 6262
rect -7703 6118 -7657 6164
rect -7703 6020 -7657 6066
rect -7703 5922 -7657 5968
rect -7703 5824 -7657 5870
rect -7703 5726 -7657 5772
rect -7703 5628 -7657 5674
rect -7703 5530 -7657 5576
rect -7703 5432 -7657 5478
rect -7703 5334 -7657 5380
rect -7703 5236 -7657 5282
rect -7703 5138 -7657 5184
rect -7703 5040 -7657 5086
rect -7703 4942 -7657 4988
rect -7703 4844 -7657 4890
rect -7703 4746 -7657 4792
rect -7703 4648 -7657 4694
rect -7703 4550 -7657 4596
rect -7703 4452 -7657 4498
rect 530 7372 576 7418
rect 3444 7466 3490 7512
rect 5606 7560 5652 7606
rect 5606 7466 5652 7512
rect 3444 7372 3490 7418
rect 5606 7372 5652 7418
rect 530 7278 576 7324
rect 624 7278 670 7324
rect 718 7278 764 7324
rect 812 7278 858 7324
rect 906 7278 952 7324
rect 1000 7278 1046 7324
rect 1094 7278 1140 7324
rect 1188 7278 1234 7324
rect 1282 7278 1328 7324
rect 1376 7278 1422 7324
rect 1470 7278 1516 7324
rect 1564 7278 1610 7324
rect 1658 7278 1704 7324
rect 1752 7278 1798 7324
rect 1846 7278 1892 7324
rect 1940 7278 1986 7324
rect 2034 7278 2080 7324
rect 2128 7278 2174 7324
rect 2222 7278 2268 7324
rect 2316 7278 2362 7324
rect 2410 7278 2456 7324
rect 2504 7278 2550 7324
rect 2598 7278 2644 7324
rect 2692 7278 2738 7324
rect 2786 7278 2832 7324
rect 2880 7278 2926 7324
rect 2974 7278 3020 7324
rect 3068 7278 3114 7324
rect 3162 7278 3208 7324
rect 3256 7278 3302 7324
rect 3350 7278 3396 7324
rect 3444 7278 3490 7324
rect 3538 7278 3584 7324
rect 3632 7278 3678 7324
rect 3726 7278 3772 7324
rect 3820 7278 3866 7324
rect 3914 7278 3960 7324
rect 4008 7278 4054 7324
rect 4102 7278 4148 7324
rect 4196 7278 4242 7324
rect 4290 7278 4336 7324
rect 4384 7278 4430 7324
rect 4478 7278 4524 7324
rect 4572 7278 4618 7324
rect 4666 7278 4712 7324
rect 4760 7278 4806 7324
rect 4854 7278 4900 7324
rect 4948 7278 4994 7324
rect 5042 7278 5088 7324
rect 5136 7278 5182 7324
rect 5230 7278 5276 7324
rect 5324 7278 5370 7324
rect 5418 7278 5464 7324
rect 5512 7278 5558 7324
rect 5606 7278 5652 7324
rect 11900 11696 11946 11742
rect 11994 11696 12040 11742
rect 12088 11696 12134 11742
rect 12182 11696 12228 11742
rect 12276 11696 12322 11742
rect 12370 11696 12416 11742
rect 12464 11696 12510 11742
rect 12558 11696 12604 11742
rect 12652 11696 12698 11742
rect 12746 11696 12792 11742
rect 12840 11696 12886 11742
rect 12934 11696 12980 11742
rect 13028 11696 13074 11742
rect 13122 11696 13168 11742
rect 13216 11696 13262 11742
rect 13310 11696 13356 11742
rect 13404 11696 13450 11742
rect 13498 11696 13544 11742
rect 13592 11696 13638 11742
rect 13686 11696 13732 11742
rect 13780 11696 13826 11742
rect 13874 11696 13920 11742
rect 13968 11696 14014 11742
rect 14062 11696 14108 11742
rect 14156 11696 14202 11742
rect 14250 11696 14296 11742
rect 14344 11696 14390 11742
rect 14438 11696 14484 11742
rect 14532 11696 14578 11742
rect 14626 11696 14672 11742
rect 14720 11696 14766 11742
rect 14814 11696 14860 11742
rect 14908 11696 14954 11742
rect 15002 11696 15048 11742
rect 15096 11696 15142 11742
rect 15190 11696 15236 11742
rect 15284 11696 15330 11742
rect 15378 11696 15424 11742
rect 15472 11696 15518 11742
rect 15566 11696 15612 11742
rect 15660 11696 15706 11742
rect 15754 11696 15800 11742
rect 15848 11696 15894 11742
rect 15942 11696 15988 11742
rect 16036 11696 16082 11742
rect 16130 11696 16176 11742
rect 16224 11696 16270 11742
rect 16318 11696 16364 11742
rect 16412 11696 16458 11742
rect 16506 11696 16552 11742
rect 16600 11696 16646 11742
rect 16694 11696 16740 11742
rect 16788 11696 16834 11742
rect 16882 11696 16928 11742
rect 16976 11696 17022 11742
rect 11900 11602 11946 11648
rect 11900 11508 11946 11554
rect 11900 11414 11946 11460
rect 14626 11602 14672 11648
rect 14626 11508 14672 11554
rect 14626 11414 14672 11460
rect 16976 11602 17022 11648
rect 16976 11508 17022 11554
rect 11900 11320 11946 11366
rect 11900 11226 11946 11272
rect 11900 11132 11946 11178
rect 11900 11038 11946 11084
rect 11900 10944 11946 10990
rect 11900 10850 11946 10896
rect 11900 10756 11946 10802
rect 16976 11414 17022 11460
rect 14626 11320 14672 11366
rect 14626 11226 14672 11272
rect 14626 11132 14672 11178
rect 14626 11038 14672 11084
rect 14626 10944 14672 10990
rect 14626 10850 14672 10896
rect 14626 10756 14672 10802
rect 11900 10662 11946 10708
rect 11900 10568 11946 10614
rect 11900 10474 11946 10520
rect 11900 10380 11946 10426
rect 16976 11320 17022 11366
rect 16976 11226 17022 11272
rect 16976 11132 17022 11178
rect 16976 11038 17022 11084
rect 16976 10944 17022 10990
rect 16976 10850 17022 10896
rect 16976 10756 17022 10802
rect 14626 10662 14672 10708
rect 14626 10568 14672 10614
rect 14626 10474 14672 10520
rect 14626 10380 14672 10426
rect 11900 10286 11946 10332
rect 11900 10192 11946 10238
rect 11900 10098 11946 10144
rect 11900 10004 11946 10050
rect 11900 9910 11946 9956
rect 11900 9816 11946 9862
rect 11900 9722 11946 9768
rect 16976 10662 17022 10708
rect 16976 10568 17022 10614
rect 16976 10474 17022 10520
rect 16976 10380 17022 10426
rect 14626 10286 14672 10332
rect 14626 10192 14672 10238
rect 14626 10098 14672 10144
rect 14626 10004 14672 10050
rect 14626 9910 14672 9956
rect 14626 9816 14672 9862
rect 14626 9722 14672 9768
rect 11900 9628 11946 9674
rect 11900 9534 11946 9580
rect 11900 9440 11946 9486
rect 11900 9346 11946 9392
rect 16976 10286 17022 10332
rect 16976 10192 17022 10238
rect 16976 10098 17022 10144
rect 16976 10004 17022 10050
rect 16976 9910 17022 9956
rect 16976 9816 17022 9862
rect 16976 9722 17022 9768
rect 14626 9628 14672 9674
rect 14626 9534 14672 9580
rect 14626 9440 14672 9486
rect 14626 9346 14672 9392
rect 11900 9252 11946 9298
rect 11900 9158 11946 9204
rect 11900 9064 11946 9110
rect 11900 8970 11946 9016
rect 11900 8876 11946 8922
rect 11900 8782 11946 8828
rect 11900 8688 11946 8734
rect 16976 9628 17022 9674
rect 16976 9534 17022 9580
rect 16976 9440 17022 9486
rect 16976 9346 17022 9392
rect 14626 9252 14672 9298
rect 14626 9158 14672 9204
rect 14626 9064 14672 9110
rect 14626 8970 14672 9016
rect 14626 8876 14672 8922
rect 14626 8782 14672 8828
rect 14626 8688 14672 8734
rect 11900 8594 11946 8640
rect 11900 8500 11946 8546
rect 11900 8406 11946 8452
rect 16976 9252 17022 9298
rect 16976 9158 17022 9204
rect 16976 9064 17022 9110
rect 16976 8970 17022 9016
rect 16976 8876 17022 8922
rect 16976 8782 17022 8828
rect 16976 8688 17022 8734
rect 14626 8594 14672 8640
rect 14626 8500 14672 8546
rect 11900 8312 11946 8358
rect 14626 8406 14672 8452
rect 16976 8594 17022 8640
rect 16976 8500 17022 8546
rect 14626 8312 14672 8358
rect 11900 8218 11946 8264
rect 11900 8124 11946 8170
rect 11900 8030 11946 8076
rect 11900 7936 11946 7982
rect 11900 7842 11946 7888
rect 11900 7748 11946 7794
rect 11900 7654 11946 7700
rect 16976 8406 17022 8452
rect 16976 8312 17022 8358
rect 14626 8218 14672 8264
rect 14626 8124 14672 8170
rect 14626 8030 14672 8076
rect 14626 7936 14672 7982
rect 14626 7842 14672 7888
rect 14626 7748 14672 7794
rect 14626 7654 14672 7700
rect 11900 7560 11946 7606
rect 16976 8218 17022 8264
rect 16976 8124 17022 8170
rect 16976 8030 17022 8076
rect 16976 7936 17022 7982
rect 16976 7842 17022 7888
rect 16976 7748 17022 7794
rect 16976 7654 17022 7700
rect 11900 7466 11946 7512
rect 11900 7372 11946 7418
rect 14626 7560 14672 7606
rect 14626 7466 14672 7512
rect 14626 7372 14672 7418
rect 16976 7560 17022 7606
rect 16976 7466 17022 7512
rect 16976 7372 17022 7418
rect 11900 7278 11946 7324
rect 11994 7278 12040 7324
rect 12088 7278 12134 7324
rect 12182 7278 12228 7324
rect 12276 7278 12322 7324
rect 12370 7278 12416 7324
rect 12464 7278 12510 7324
rect 12558 7278 12604 7324
rect 12652 7278 12698 7324
rect 12746 7278 12792 7324
rect 12840 7278 12886 7324
rect 12934 7278 12980 7324
rect 13028 7278 13074 7324
rect 13122 7278 13168 7324
rect 13216 7278 13262 7324
rect 13310 7278 13356 7324
rect 13404 7278 13450 7324
rect 13498 7278 13544 7324
rect 13592 7278 13638 7324
rect 13686 7278 13732 7324
rect 13780 7278 13826 7324
rect 13874 7278 13920 7324
rect 13968 7278 14014 7324
rect 14062 7278 14108 7324
rect 14156 7278 14202 7324
rect 14250 7278 14296 7324
rect 14344 7278 14390 7324
rect 14438 7278 14484 7324
rect 14532 7278 14578 7324
rect 14626 7278 14672 7324
rect 14720 7278 14766 7324
rect 14814 7278 14860 7324
rect 14908 7278 14954 7324
rect 15002 7278 15048 7324
rect 15096 7278 15142 7324
rect 15190 7278 15236 7324
rect 15284 7278 15330 7324
rect 15378 7278 15424 7324
rect 15472 7278 15518 7324
rect 15566 7278 15612 7324
rect 15660 7278 15706 7324
rect 15754 7278 15800 7324
rect 15848 7278 15894 7324
rect 15942 7278 15988 7324
rect 16036 7278 16082 7324
rect 16130 7278 16176 7324
rect 16224 7278 16270 7324
rect 16318 7278 16364 7324
rect 16412 7278 16458 7324
rect 16506 7278 16552 7324
rect 16600 7278 16646 7324
rect 16694 7278 16740 7324
rect 16788 7278 16834 7324
rect 16882 7278 16928 7324
rect 16976 7278 17022 7324
rect 32629 12173 32675 12219
rect 32723 12173 32769 12219
rect 32817 12173 32863 12219
rect 32911 12173 32957 12219
rect 33005 12173 33051 12219
rect 33099 12173 33145 12219
rect 33193 12173 33239 12219
rect 33287 12173 33333 12219
rect 33381 12173 33427 12219
rect 33475 12173 33521 12219
rect 33569 12173 33615 12219
rect 33663 12173 33709 12219
rect 33757 12173 33803 12219
rect 33851 12173 33897 12219
rect 33945 12173 33991 12219
rect 34039 12173 34085 12219
rect 34133 12173 34179 12219
rect 34227 12173 34273 12219
rect 34321 12173 34367 12219
rect 34415 12173 34461 12219
rect 34509 12173 34555 12219
rect 34603 12173 34649 12219
rect 34697 12173 34743 12219
rect 34791 12173 34837 12219
rect 34885 12173 34931 12219
rect 34979 12173 35025 12219
rect 35073 12173 35119 12219
rect 35167 12173 35213 12219
rect 35261 12173 35307 12219
rect 35355 12173 35401 12219
rect 35449 12173 35495 12219
rect 35543 12173 35589 12219
rect 35637 12173 35683 12219
rect 35731 12173 35777 12219
rect 35825 12173 35871 12219
rect 35919 12173 35965 12219
rect 36013 12173 36059 12219
rect 36107 12173 36153 12219
rect 36201 12173 36247 12219
rect 36295 12173 36341 12219
rect 36389 12173 36435 12219
rect 36483 12173 36529 12219
rect 36577 12173 36623 12219
rect 36671 12173 36717 12219
rect 36765 12173 36811 12219
rect 36859 12173 36905 12219
rect 36953 12173 36999 12219
rect 37047 12173 37093 12219
rect 37141 12173 37187 12219
rect 37235 12173 37281 12219
rect 37329 12173 37375 12219
rect 37423 12173 37469 12219
rect 37517 12173 37563 12219
rect 37611 12173 37657 12219
rect 37705 12173 37751 12219
rect 37799 12173 37845 12219
rect 37893 12173 37939 12219
rect 37987 12173 38033 12219
rect 38081 12173 38127 12219
rect 38175 12173 38221 12219
rect 38269 12173 38315 12219
rect 38363 12173 38409 12219
rect 38457 12173 38503 12219
rect 38551 12173 38597 12219
rect 38645 12173 38691 12219
rect 38739 12173 38785 12219
rect 38833 12173 38879 12219
rect 38927 12173 38973 12219
rect 39021 12173 39067 12219
rect 39115 12173 39161 12219
rect 39209 12173 39255 12219
rect 39303 12173 39349 12219
rect 39397 12173 39443 12219
rect 39491 12173 39537 12219
rect 39585 12173 39631 12219
rect 39679 12173 39725 12219
rect 39773 12173 39819 12219
rect 39867 12173 39913 12219
rect 39961 12173 40007 12219
rect 40055 12173 40101 12219
rect 40149 12173 40195 12219
rect 40243 12173 40289 12219
rect 40337 12173 40383 12219
rect 40431 12173 40477 12219
rect 40525 12173 40571 12219
rect 40619 12173 40665 12219
rect 40713 12173 40759 12219
rect 40807 12173 40853 12219
rect 40901 12173 40947 12219
rect 32629 12079 32675 12125
rect 32629 11985 32675 12031
rect 32629 11891 32675 11937
rect 32629 11797 32675 11843
rect 36765 12079 36811 12125
rect 36765 11985 36811 12031
rect 36765 11891 36811 11937
rect 36765 11797 36811 11843
rect 40901 12079 40947 12125
rect 40901 11985 40947 12031
rect 40901 11891 40947 11937
rect 32629 11703 32675 11749
rect 40901 11797 40947 11843
rect 36765 11703 36811 11749
rect 32629 11609 32675 11655
rect 32629 11515 32675 11561
rect 32629 11421 32675 11467
rect 32629 11327 32675 11373
rect 32629 11233 32675 11279
rect 32629 11139 32675 11185
rect 32629 11045 32675 11091
rect 40901 11703 40947 11749
rect 36765 11609 36811 11655
rect 36765 11515 36811 11561
rect 36765 11421 36811 11467
rect 36765 11327 36811 11373
rect 36765 11233 36811 11279
rect 36765 11139 36811 11185
rect 32629 10951 32675 10997
rect 32629 10857 32675 10903
rect 32629 10763 32675 10809
rect 32629 10669 32675 10715
rect 36765 11045 36811 11091
rect 40901 11609 40947 11655
rect 40901 11515 40947 11561
rect 40901 11421 40947 11467
rect 40901 11327 40947 11373
rect 40901 11233 40947 11279
rect 40901 11139 40947 11185
rect 36765 10951 36811 10997
rect 36765 10857 36811 10903
rect 36765 10763 36811 10809
rect 36765 10669 36811 10715
rect 32629 10575 32675 10621
rect 32629 10481 32675 10527
rect 32629 10387 32675 10433
rect 32629 10293 32675 10339
rect 32629 10199 32675 10245
rect 32629 10105 32675 10151
rect 32629 10011 32675 10057
rect 40901 11045 40947 11091
rect 40901 10951 40947 10997
rect 40901 10857 40947 10903
rect 40901 10763 40947 10809
rect 40901 10669 40947 10715
rect 36765 10575 36811 10621
rect 36765 10481 36811 10527
rect 36765 10387 36811 10433
rect 36765 10293 36811 10339
rect 36765 10199 36811 10245
rect 36765 10105 36811 10151
rect 32629 9917 32675 9963
rect 32629 9823 32675 9869
rect 32629 9729 32675 9775
rect 32629 9635 32675 9681
rect 32629 9541 32675 9587
rect 36765 10011 36811 10057
rect 40901 10575 40947 10621
rect 40901 10481 40947 10527
rect 40901 10387 40947 10433
rect 40901 10293 40947 10339
rect 40901 10199 40947 10245
rect 40901 10105 40947 10151
rect 36765 9917 36811 9963
rect 36765 9823 36811 9869
rect 36765 9729 36811 9775
rect 36765 9635 36811 9681
rect 32629 9447 32675 9493
rect 32629 9353 32675 9399
rect 32629 9259 32675 9305
rect 32629 9165 32675 9211
rect 32629 9071 32675 9117
rect 32629 8977 32675 9023
rect 36765 9541 36811 9587
rect 40901 10011 40947 10057
rect 40901 9917 40947 9963
rect 40901 9823 40947 9869
rect 40901 9729 40947 9775
rect 40901 9635 40947 9681
rect 36765 9447 36811 9493
rect 36765 9353 36811 9399
rect 36765 9259 36811 9305
rect 36765 9165 36811 9211
rect 36765 9071 36811 9117
rect 36765 8977 36811 9023
rect 32629 8883 32675 8929
rect 32629 8789 32675 8835
rect 32629 8695 32675 8741
rect 32629 8601 32675 8647
rect 32629 8507 32675 8553
rect 40901 9541 40947 9587
rect 40901 9447 40947 9493
rect 40901 9353 40947 9399
rect 40901 9259 40947 9305
rect 40901 9165 40947 9211
rect 40901 9071 40947 9117
rect 40901 8977 40947 9023
rect 36765 8883 36811 8929
rect 36765 8789 36811 8835
rect 36765 8695 36811 8741
rect 36765 8601 36811 8647
rect 32629 8413 32675 8459
rect 32629 8319 32675 8365
rect 32629 8225 32675 8271
rect 32629 8131 32675 8177
rect 32629 8037 32675 8083
rect 32629 7943 32675 7989
rect 36765 8507 36811 8553
rect 40901 8883 40947 8929
rect 40901 8789 40947 8835
rect 40901 8695 40947 8741
rect 40901 8601 40947 8647
rect 36765 8413 36811 8459
rect 36765 8319 36811 8365
rect 36765 8225 36811 8271
rect 36765 8131 36811 8177
rect 36765 8037 36811 8083
rect 36765 7943 36811 7989
rect 32629 7849 32675 7895
rect 40901 8507 40947 8553
rect 40901 8413 40947 8459
rect 40901 8319 40947 8365
rect 40901 8225 40947 8271
rect 40901 8131 40947 8177
rect 40901 8037 40947 8083
rect 40901 7943 40947 7989
rect 32629 7755 32675 7801
rect 32629 7661 32675 7707
rect 32629 7567 32675 7613
rect 32629 7473 32675 7519
rect 36765 7849 36811 7895
rect 36765 7755 36811 7801
rect 36765 7661 36811 7707
rect 36765 7567 36811 7613
rect 36765 7473 36811 7519
rect 40901 7849 40947 7895
rect 40901 7755 40947 7801
rect 40901 7661 40947 7707
rect 40901 7567 40947 7613
rect 40901 7473 40947 7519
rect 32629 7379 32675 7425
rect 32723 7379 32769 7425
rect 32817 7379 32863 7425
rect 32911 7379 32957 7425
rect 33005 7379 33051 7425
rect 33099 7379 33145 7425
rect 33193 7379 33239 7425
rect 33287 7379 33333 7425
rect 33381 7379 33427 7425
rect 33475 7379 33521 7425
rect 33569 7379 33615 7425
rect 33663 7379 33709 7425
rect 33757 7379 33803 7425
rect 33851 7379 33897 7425
rect 33945 7379 33991 7425
rect 34039 7379 34085 7425
rect 34133 7379 34179 7425
rect 34227 7379 34273 7425
rect 34321 7379 34367 7425
rect 34415 7379 34461 7425
rect 34509 7379 34555 7425
rect 34603 7379 34649 7425
rect 34697 7379 34743 7425
rect 34791 7379 34837 7425
rect 34885 7379 34931 7425
rect 34979 7379 35025 7425
rect 35073 7379 35119 7425
rect 35167 7379 35213 7425
rect 35261 7379 35307 7425
rect 35355 7379 35401 7425
rect 35449 7379 35495 7425
rect 35543 7379 35589 7425
rect 35637 7379 35683 7425
rect 35731 7379 35777 7425
rect 35825 7379 35871 7425
rect 35919 7379 35965 7425
rect 36013 7379 36059 7425
rect 36107 7379 36153 7425
rect 36201 7379 36247 7425
rect 36295 7379 36341 7425
rect 36389 7379 36435 7425
rect 36483 7379 36529 7425
rect 36577 7379 36623 7425
rect 36671 7379 36717 7425
rect 36765 7379 36811 7425
rect 36859 7379 36905 7425
rect 36953 7379 36999 7425
rect 37047 7379 37093 7425
rect 37141 7379 37187 7425
rect 37235 7379 37281 7425
rect 37329 7379 37375 7425
rect 37423 7379 37469 7425
rect 37517 7379 37563 7425
rect 37611 7379 37657 7425
rect 37705 7379 37751 7425
rect 37799 7379 37845 7425
rect 37893 7379 37939 7425
rect 37987 7379 38033 7425
rect 38081 7379 38127 7425
rect 38175 7379 38221 7425
rect 38269 7379 38315 7425
rect 38363 7379 38409 7425
rect 38457 7379 38503 7425
rect 38551 7379 38597 7425
rect 38645 7379 38691 7425
rect 38739 7379 38785 7425
rect 38833 7379 38879 7425
rect 38927 7379 38973 7425
rect 39021 7379 39067 7425
rect 39115 7379 39161 7425
rect 39209 7379 39255 7425
rect 39303 7379 39349 7425
rect 39397 7379 39443 7425
rect 39491 7379 39537 7425
rect 39585 7379 39631 7425
rect 39679 7379 39725 7425
rect 39773 7379 39819 7425
rect 39867 7379 39913 7425
rect 39961 7379 40007 7425
rect 40055 7379 40101 7425
rect 40149 7379 40195 7425
rect 40243 7379 40289 7425
rect 40337 7379 40383 7425
rect 40431 7379 40477 7425
rect 40525 7379 40571 7425
rect 40619 7379 40665 7425
rect 40713 7379 40759 7425
rect 40807 7379 40853 7425
rect 40901 7379 40947 7425
rect 42325 12173 42371 12219
rect 42419 12173 42465 12219
rect 42513 12173 42559 12219
rect 42607 12173 42653 12219
rect 42701 12173 42747 12219
rect 42795 12173 42841 12219
rect 42889 12173 42935 12219
rect 42983 12173 43029 12219
rect 43077 12173 43123 12219
rect 43171 12173 43217 12219
rect 43265 12173 43311 12219
rect 43359 12173 43405 12219
rect 43453 12173 43499 12219
rect 43547 12173 43593 12219
rect 43641 12173 43687 12219
rect 43735 12173 43781 12219
rect 43829 12173 43875 12219
rect 43923 12173 43969 12219
rect 44017 12173 44063 12219
rect 44111 12173 44157 12219
rect 44205 12173 44251 12219
rect 44299 12173 44345 12219
rect 44393 12173 44439 12219
rect 44487 12173 44533 12219
rect 44581 12173 44627 12219
rect 44675 12173 44721 12219
rect 44769 12173 44815 12219
rect 44863 12173 44909 12219
rect 44957 12173 45003 12219
rect 45051 12173 45097 12219
rect 45145 12173 45191 12219
rect 45239 12173 45285 12219
rect 45333 12173 45379 12219
rect 45427 12173 45473 12219
rect 45521 12173 45567 12219
rect 45615 12173 45661 12219
rect 45709 12173 45755 12219
rect 45803 12173 45849 12219
rect 45897 12173 45943 12219
rect 45991 12173 46037 12219
rect 46085 12173 46131 12219
rect 46179 12173 46225 12219
rect 46273 12173 46319 12219
rect 46367 12173 46413 12219
rect 46461 12173 46507 12219
rect 46555 12173 46601 12219
rect 46649 12173 46695 12219
rect 46743 12173 46789 12219
rect 46837 12173 46883 12219
rect 46931 12173 46977 12219
rect 47025 12173 47071 12219
rect 47119 12173 47165 12219
rect 47213 12173 47259 12219
rect 47307 12173 47353 12219
rect 47401 12173 47447 12219
rect 47495 12173 47541 12219
rect 47589 12173 47635 12219
rect 47683 12173 47729 12219
rect 47777 12173 47823 12219
rect 47871 12173 47917 12219
rect 47965 12173 48011 12219
rect 48059 12173 48105 12219
rect 48153 12173 48199 12219
rect 48247 12173 48293 12219
rect 48341 12173 48387 12219
rect 48435 12173 48481 12219
rect 48529 12173 48575 12219
rect 48623 12173 48669 12219
rect 48717 12173 48763 12219
rect 48811 12173 48857 12219
rect 48905 12173 48951 12219
rect 48999 12173 49045 12219
rect 49093 12173 49139 12219
rect 49187 12173 49233 12219
rect 49281 12173 49327 12219
rect 49375 12173 49421 12219
rect 49469 12173 49515 12219
rect 49563 12173 49609 12219
rect 49657 12173 49703 12219
rect 49751 12173 49797 12219
rect 49845 12173 49891 12219
rect 49939 12173 49985 12219
rect 50033 12173 50079 12219
rect 50127 12173 50173 12219
rect 50221 12173 50267 12219
rect 50315 12173 50361 12219
rect 50409 12173 50455 12219
rect 50503 12173 50549 12219
rect 50597 12173 50643 12219
rect 42325 12079 42371 12125
rect 42325 11985 42371 12031
rect 42325 11891 42371 11937
rect 42325 11797 42371 11843
rect 46461 12079 46507 12125
rect 46461 11985 46507 12031
rect 46461 11891 46507 11937
rect 46461 11797 46507 11843
rect 50597 12079 50643 12125
rect 50597 11985 50643 12031
rect 50597 11891 50643 11937
rect 42325 11703 42371 11749
rect 50597 11797 50643 11843
rect 46461 11703 46507 11749
rect 42325 11609 42371 11655
rect 42325 11515 42371 11561
rect 42325 11421 42371 11467
rect 42325 11327 42371 11373
rect 42325 11233 42371 11279
rect 42325 11139 42371 11185
rect 42325 11045 42371 11091
rect 50597 11703 50643 11749
rect 46461 11609 46507 11655
rect 46461 11515 46507 11561
rect 46461 11421 46507 11467
rect 46461 11327 46507 11373
rect 46461 11233 46507 11279
rect 46461 11139 46507 11185
rect 42325 10951 42371 10997
rect 42325 10857 42371 10903
rect 42325 10763 42371 10809
rect 42325 10669 42371 10715
rect 46461 11045 46507 11091
rect 50597 11609 50643 11655
rect 50597 11515 50643 11561
rect 50597 11421 50643 11467
rect 50597 11327 50643 11373
rect 50597 11233 50643 11279
rect 50597 11139 50643 11185
rect 46461 10951 46507 10997
rect 46461 10857 46507 10903
rect 46461 10763 46507 10809
rect 46461 10669 46507 10715
rect 42325 10575 42371 10621
rect 42325 10481 42371 10527
rect 42325 10387 42371 10433
rect 42325 10293 42371 10339
rect 42325 10199 42371 10245
rect 42325 10105 42371 10151
rect 42325 10011 42371 10057
rect 50597 11045 50643 11091
rect 50597 10951 50643 10997
rect 50597 10857 50643 10903
rect 50597 10763 50643 10809
rect 50597 10669 50643 10715
rect 46461 10575 46507 10621
rect 46461 10481 46507 10527
rect 46461 10387 46507 10433
rect 46461 10293 46507 10339
rect 46461 10199 46507 10245
rect 46461 10105 46507 10151
rect 42325 9917 42371 9963
rect 42325 9823 42371 9869
rect 42325 9729 42371 9775
rect 42325 9635 42371 9681
rect 42325 9541 42371 9587
rect 46461 10011 46507 10057
rect 50597 10575 50643 10621
rect 50597 10481 50643 10527
rect 50597 10387 50643 10433
rect 50597 10293 50643 10339
rect 50597 10199 50643 10245
rect 50597 10105 50643 10151
rect 46461 9917 46507 9963
rect 46461 9823 46507 9869
rect 46461 9729 46507 9775
rect 46461 9635 46507 9681
rect 42325 9447 42371 9493
rect 42325 9353 42371 9399
rect 42325 9259 42371 9305
rect 42325 9165 42371 9211
rect 42325 9071 42371 9117
rect 42325 8977 42371 9023
rect 46461 9541 46507 9587
rect 50597 10011 50643 10057
rect 50597 9917 50643 9963
rect 50597 9823 50643 9869
rect 50597 9729 50643 9775
rect 50597 9635 50643 9681
rect 46461 9447 46507 9493
rect 46461 9353 46507 9399
rect 46461 9259 46507 9305
rect 46461 9165 46507 9211
rect 46461 9071 46507 9117
rect 46461 8977 46507 9023
rect 42325 8883 42371 8929
rect 42325 8789 42371 8835
rect 42325 8695 42371 8741
rect 42325 8601 42371 8647
rect 42325 8507 42371 8553
rect 50597 9541 50643 9587
rect 50597 9447 50643 9493
rect 50597 9353 50643 9399
rect 50597 9259 50643 9305
rect 50597 9165 50643 9211
rect 50597 9071 50643 9117
rect 50597 8977 50643 9023
rect 46461 8883 46507 8929
rect 46461 8789 46507 8835
rect 46461 8695 46507 8741
rect 46461 8601 46507 8647
rect 42325 8413 42371 8459
rect 42325 8319 42371 8365
rect 42325 8225 42371 8271
rect 42325 8131 42371 8177
rect 42325 8037 42371 8083
rect 42325 7943 42371 7989
rect 46461 8507 46507 8553
rect 50597 8883 50643 8929
rect 50597 8789 50643 8835
rect 50597 8695 50643 8741
rect 50597 8601 50643 8647
rect 46461 8413 46507 8459
rect 46461 8319 46507 8365
rect 46461 8225 46507 8271
rect 46461 8131 46507 8177
rect 46461 8037 46507 8083
rect 46461 7943 46507 7989
rect 42325 7849 42371 7895
rect 50597 8507 50643 8553
rect 50597 8413 50643 8459
rect 50597 8319 50643 8365
rect 50597 8225 50643 8271
rect 50597 8131 50643 8177
rect 50597 8037 50643 8083
rect 50597 7943 50643 7989
rect 42325 7755 42371 7801
rect 42325 7661 42371 7707
rect 42325 7567 42371 7613
rect 42325 7473 42371 7519
rect 46461 7849 46507 7895
rect 46461 7755 46507 7801
rect 46461 7661 46507 7707
rect 46461 7567 46507 7613
rect 46461 7473 46507 7519
rect 50597 7849 50643 7895
rect 50597 7755 50643 7801
rect 50597 7661 50643 7707
rect 50597 7567 50643 7613
rect 50597 7473 50643 7519
rect 42325 7379 42371 7425
rect 42419 7379 42465 7425
rect 42513 7379 42559 7425
rect 42607 7379 42653 7425
rect 42701 7379 42747 7425
rect 42795 7379 42841 7425
rect 42889 7379 42935 7425
rect 42983 7379 43029 7425
rect 43077 7379 43123 7425
rect 43171 7379 43217 7425
rect 43265 7379 43311 7425
rect 43359 7379 43405 7425
rect 43453 7379 43499 7425
rect 43547 7379 43593 7425
rect 43641 7379 43687 7425
rect 43735 7379 43781 7425
rect 43829 7379 43875 7425
rect 43923 7379 43969 7425
rect 44017 7379 44063 7425
rect 44111 7379 44157 7425
rect 44205 7379 44251 7425
rect 44299 7379 44345 7425
rect 44393 7379 44439 7425
rect 44487 7379 44533 7425
rect 44581 7379 44627 7425
rect 44675 7379 44721 7425
rect 44769 7379 44815 7425
rect 44863 7379 44909 7425
rect 44957 7379 45003 7425
rect 45051 7379 45097 7425
rect 45145 7379 45191 7425
rect 45239 7379 45285 7425
rect 45333 7379 45379 7425
rect 45427 7379 45473 7425
rect 45521 7379 45567 7425
rect 45615 7379 45661 7425
rect 45709 7379 45755 7425
rect 45803 7379 45849 7425
rect 45897 7379 45943 7425
rect 45991 7379 46037 7425
rect 46085 7379 46131 7425
rect 46179 7379 46225 7425
rect 46273 7379 46319 7425
rect 46367 7379 46413 7425
rect 46461 7379 46507 7425
rect 46555 7379 46601 7425
rect 46649 7379 46695 7425
rect 46743 7379 46789 7425
rect 46837 7379 46883 7425
rect 46931 7379 46977 7425
rect 47025 7379 47071 7425
rect 47119 7379 47165 7425
rect 47213 7379 47259 7425
rect 47307 7379 47353 7425
rect 47401 7379 47447 7425
rect 47495 7379 47541 7425
rect 47589 7379 47635 7425
rect 47683 7379 47729 7425
rect 47777 7379 47823 7425
rect 47871 7379 47917 7425
rect 47965 7379 48011 7425
rect 48059 7379 48105 7425
rect 48153 7379 48199 7425
rect 48247 7379 48293 7425
rect 48341 7379 48387 7425
rect 48435 7379 48481 7425
rect 48529 7379 48575 7425
rect 48623 7379 48669 7425
rect 48717 7379 48763 7425
rect 48811 7379 48857 7425
rect 48905 7379 48951 7425
rect 48999 7379 49045 7425
rect 49093 7379 49139 7425
rect 49187 7379 49233 7425
rect 49281 7379 49327 7425
rect 49375 7379 49421 7425
rect 49469 7379 49515 7425
rect 49563 7379 49609 7425
rect 49657 7379 49703 7425
rect 49751 7379 49797 7425
rect 49845 7379 49891 7425
rect 49939 7379 49985 7425
rect 50033 7379 50079 7425
rect 50127 7379 50173 7425
rect 50221 7379 50267 7425
rect 50315 7379 50361 7425
rect 50409 7379 50455 7425
rect 50503 7379 50549 7425
rect 50597 7379 50643 7425
rect 52021 12173 52067 12219
rect 52115 12173 52161 12219
rect 52209 12173 52255 12219
rect 52303 12173 52349 12219
rect 52397 12173 52443 12219
rect 52491 12173 52537 12219
rect 52585 12173 52631 12219
rect 52679 12173 52725 12219
rect 52773 12173 52819 12219
rect 52867 12173 52913 12219
rect 52961 12173 53007 12219
rect 53055 12173 53101 12219
rect 53149 12173 53195 12219
rect 53243 12173 53289 12219
rect 53337 12173 53383 12219
rect 53431 12173 53477 12219
rect 53525 12173 53571 12219
rect 53619 12173 53665 12219
rect 53713 12173 53759 12219
rect 53807 12173 53853 12219
rect 53901 12173 53947 12219
rect 53995 12173 54041 12219
rect 54089 12173 54135 12219
rect 54183 12173 54229 12219
rect 54277 12173 54323 12219
rect 54371 12173 54417 12219
rect 54465 12173 54511 12219
rect 54559 12173 54605 12219
rect 54653 12173 54699 12219
rect 54747 12173 54793 12219
rect 54841 12173 54887 12219
rect 54935 12173 54981 12219
rect 55029 12173 55075 12219
rect 55123 12173 55169 12219
rect 55217 12173 55263 12219
rect 55311 12173 55357 12219
rect 55405 12173 55451 12219
rect 55499 12173 55545 12219
rect 55593 12173 55639 12219
rect 55687 12173 55733 12219
rect 55781 12173 55827 12219
rect 55875 12173 55921 12219
rect 55969 12173 56015 12219
rect 56063 12173 56109 12219
rect 56157 12173 56203 12219
rect 56251 12173 56297 12219
rect 56345 12173 56391 12219
rect 56439 12173 56485 12219
rect 56533 12173 56579 12219
rect 56627 12173 56673 12219
rect 56721 12173 56767 12219
rect 56815 12173 56861 12219
rect 56909 12173 56955 12219
rect 57003 12173 57049 12219
rect 57097 12173 57143 12219
rect 57191 12173 57237 12219
rect 57285 12173 57331 12219
rect 57379 12173 57425 12219
rect 57473 12173 57519 12219
rect 57567 12173 57613 12219
rect 57661 12173 57707 12219
rect 57755 12173 57801 12219
rect 57849 12173 57895 12219
rect 57943 12173 57989 12219
rect 58037 12173 58083 12219
rect 58131 12173 58177 12219
rect 58225 12173 58271 12219
rect 58319 12173 58365 12219
rect 58413 12173 58459 12219
rect 58507 12173 58553 12219
rect 58601 12173 58647 12219
rect 58695 12173 58741 12219
rect 58789 12173 58835 12219
rect 58883 12173 58929 12219
rect 58977 12173 59023 12219
rect 59071 12173 59117 12219
rect 59165 12173 59211 12219
rect 59259 12173 59305 12219
rect 59353 12173 59399 12219
rect 59447 12173 59493 12219
rect 59541 12173 59587 12219
rect 59635 12173 59681 12219
rect 59729 12173 59775 12219
rect 59823 12173 59869 12219
rect 59917 12173 59963 12219
rect 60011 12173 60057 12219
rect 60105 12173 60151 12219
rect 60199 12173 60245 12219
rect 60293 12173 60339 12219
rect 52021 12079 52067 12125
rect 52021 11985 52067 12031
rect 52021 11891 52067 11937
rect 52021 11797 52067 11843
rect 56157 12079 56203 12125
rect 56157 11985 56203 12031
rect 56157 11891 56203 11937
rect 56157 11797 56203 11843
rect 60293 12079 60339 12125
rect 60293 11985 60339 12031
rect 60293 11891 60339 11937
rect 52021 11703 52067 11749
rect 60293 11797 60339 11843
rect 56157 11703 56203 11749
rect 52021 11609 52067 11655
rect 52021 11515 52067 11561
rect 52021 11421 52067 11467
rect 52021 11327 52067 11373
rect 52021 11233 52067 11279
rect 52021 11139 52067 11185
rect 52021 11045 52067 11091
rect 60293 11703 60339 11749
rect 56157 11609 56203 11655
rect 56157 11515 56203 11561
rect 56157 11421 56203 11467
rect 56157 11327 56203 11373
rect 56157 11233 56203 11279
rect 56157 11139 56203 11185
rect 52021 10951 52067 10997
rect 52021 10857 52067 10903
rect 52021 10763 52067 10809
rect 52021 10669 52067 10715
rect 56157 11045 56203 11091
rect 60293 11609 60339 11655
rect 60293 11515 60339 11561
rect 60293 11421 60339 11467
rect 60293 11327 60339 11373
rect 60293 11233 60339 11279
rect 60293 11139 60339 11185
rect 56157 10951 56203 10997
rect 56157 10857 56203 10903
rect 56157 10763 56203 10809
rect 56157 10669 56203 10715
rect 52021 10575 52067 10621
rect 52021 10481 52067 10527
rect 52021 10387 52067 10433
rect 52021 10293 52067 10339
rect 52021 10199 52067 10245
rect 52021 10105 52067 10151
rect 52021 10011 52067 10057
rect 60293 11045 60339 11091
rect 60293 10951 60339 10997
rect 60293 10857 60339 10903
rect 60293 10763 60339 10809
rect 60293 10669 60339 10715
rect 56157 10575 56203 10621
rect 56157 10481 56203 10527
rect 56157 10387 56203 10433
rect 56157 10293 56203 10339
rect 56157 10199 56203 10245
rect 56157 10105 56203 10151
rect 52021 9917 52067 9963
rect 52021 9823 52067 9869
rect 52021 9729 52067 9775
rect 52021 9635 52067 9681
rect 52021 9541 52067 9587
rect 56157 10011 56203 10057
rect 60293 10575 60339 10621
rect 60293 10481 60339 10527
rect 60293 10387 60339 10433
rect 60293 10293 60339 10339
rect 60293 10199 60339 10245
rect 60293 10105 60339 10151
rect 56157 9917 56203 9963
rect 56157 9823 56203 9869
rect 56157 9729 56203 9775
rect 56157 9635 56203 9681
rect 52021 9447 52067 9493
rect 52021 9353 52067 9399
rect 52021 9259 52067 9305
rect 52021 9165 52067 9211
rect 52021 9071 52067 9117
rect 52021 8977 52067 9023
rect 56157 9541 56203 9587
rect 60293 10011 60339 10057
rect 60293 9917 60339 9963
rect 60293 9823 60339 9869
rect 60293 9729 60339 9775
rect 60293 9635 60339 9681
rect 56157 9447 56203 9493
rect 56157 9353 56203 9399
rect 56157 9259 56203 9305
rect 56157 9165 56203 9211
rect 56157 9071 56203 9117
rect 56157 8977 56203 9023
rect 52021 8883 52067 8929
rect 52021 8789 52067 8835
rect 52021 8695 52067 8741
rect 52021 8601 52067 8647
rect 52021 8507 52067 8553
rect 60293 9541 60339 9587
rect 60293 9447 60339 9493
rect 60293 9353 60339 9399
rect 60293 9259 60339 9305
rect 60293 9165 60339 9211
rect 60293 9071 60339 9117
rect 60293 8977 60339 9023
rect 56157 8883 56203 8929
rect 56157 8789 56203 8835
rect 56157 8695 56203 8741
rect 56157 8601 56203 8647
rect 52021 8413 52067 8459
rect 52021 8319 52067 8365
rect 52021 8225 52067 8271
rect 52021 8131 52067 8177
rect 52021 8037 52067 8083
rect 52021 7943 52067 7989
rect 56157 8507 56203 8553
rect 60293 8883 60339 8929
rect 60293 8789 60339 8835
rect 60293 8695 60339 8741
rect 60293 8601 60339 8647
rect 56157 8413 56203 8459
rect 56157 8319 56203 8365
rect 56157 8225 56203 8271
rect 56157 8131 56203 8177
rect 56157 8037 56203 8083
rect 56157 7943 56203 7989
rect 52021 7849 52067 7895
rect 60293 8507 60339 8553
rect 60293 8413 60339 8459
rect 60293 8319 60339 8365
rect 60293 8225 60339 8271
rect 60293 8131 60339 8177
rect 60293 8037 60339 8083
rect 60293 7943 60339 7989
rect 52021 7755 52067 7801
rect 52021 7661 52067 7707
rect 52021 7567 52067 7613
rect 52021 7473 52067 7519
rect 56157 7849 56203 7895
rect 56157 7755 56203 7801
rect 56157 7661 56203 7707
rect 56157 7567 56203 7613
rect 56157 7473 56203 7519
rect 60293 7849 60339 7895
rect 60293 7755 60339 7801
rect 60293 7661 60339 7707
rect 60293 7567 60339 7613
rect 60293 7473 60339 7519
rect 52021 7379 52067 7425
rect 52115 7379 52161 7425
rect 52209 7379 52255 7425
rect 52303 7379 52349 7425
rect 52397 7379 52443 7425
rect 52491 7379 52537 7425
rect 52585 7379 52631 7425
rect 52679 7379 52725 7425
rect 52773 7379 52819 7425
rect 52867 7379 52913 7425
rect 52961 7379 53007 7425
rect 53055 7379 53101 7425
rect 53149 7379 53195 7425
rect 53243 7379 53289 7425
rect 53337 7379 53383 7425
rect 53431 7379 53477 7425
rect 53525 7379 53571 7425
rect 53619 7379 53665 7425
rect 53713 7379 53759 7425
rect 53807 7379 53853 7425
rect 53901 7379 53947 7425
rect 53995 7379 54041 7425
rect 54089 7379 54135 7425
rect 54183 7379 54229 7425
rect 54277 7379 54323 7425
rect 54371 7379 54417 7425
rect 54465 7379 54511 7425
rect 54559 7379 54605 7425
rect 54653 7379 54699 7425
rect 54747 7379 54793 7425
rect 54841 7379 54887 7425
rect 54935 7379 54981 7425
rect 55029 7379 55075 7425
rect 55123 7379 55169 7425
rect 55217 7379 55263 7425
rect 55311 7379 55357 7425
rect 55405 7379 55451 7425
rect 55499 7379 55545 7425
rect 55593 7379 55639 7425
rect 55687 7379 55733 7425
rect 55781 7379 55827 7425
rect 55875 7379 55921 7425
rect 55969 7379 56015 7425
rect 56063 7379 56109 7425
rect 56157 7379 56203 7425
rect 56251 7379 56297 7425
rect 56345 7379 56391 7425
rect 56439 7379 56485 7425
rect 56533 7379 56579 7425
rect 56627 7379 56673 7425
rect 56721 7379 56767 7425
rect 56815 7379 56861 7425
rect 56909 7379 56955 7425
rect 57003 7379 57049 7425
rect 57097 7379 57143 7425
rect 57191 7379 57237 7425
rect 57285 7379 57331 7425
rect 57379 7379 57425 7425
rect 57473 7379 57519 7425
rect 57567 7379 57613 7425
rect 57661 7379 57707 7425
rect 57755 7379 57801 7425
rect 57849 7379 57895 7425
rect 57943 7379 57989 7425
rect 58037 7379 58083 7425
rect 58131 7379 58177 7425
rect 58225 7379 58271 7425
rect 58319 7379 58365 7425
rect 58413 7379 58459 7425
rect 58507 7379 58553 7425
rect 58601 7379 58647 7425
rect 58695 7379 58741 7425
rect 58789 7379 58835 7425
rect 58883 7379 58929 7425
rect 58977 7379 59023 7425
rect 59071 7379 59117 7425
rect 59165 7379 59211 7425
rect 59259 7379 59305 7425
rect 59353 7379 59399 7425
rect 59447 7379 59493 7425
rect 59541 7379 59587 7425
rect 59635 7379 59681 7425
rect 59729 7379 59775 7425
rect 59823 7379 59869 7425
rect 59917 7379 59963 7425
rect 60011 7379 60057 7425
rect 60105 7379 60151 7425
rect 60199 7379 60245 7425
rect 60293 7379 60339 7425
rect 61717 12173 61763 12219
rect 61811 12173 61857 12219
rect 61905 12173 61951 12219
rect 61999 12173 62045 12219
rect 62093 12173 62139 12219
rect 62187 12173 62233 12219
rect 62281 12173 62327 12219
rect 62375 12173 62421 12219
rect 62469 12173 62515 12219
rect 62563 12173 62609 12219
rect 62657 12173 62703 12219
rect 62751 12173 62797 12219
rect 62845 12173 62891 12219
rect 62939 12173 62985 12219
rect 63033 12173 63079 12219
rect 63127 12173 63173 12219
rect 63221 12173 63267 12219
rect 63315 12173 63361 12219
rect 63409 12173 63455 12219
rect 63503 12173 63549 12219
rect 63597 12173 63643 12219
rect 63691 12173 63737 12219
rect 63785 12173 63831 12219
rect 63879 12173 63925 12219
rect 63973 12173 64019 12219
rect 64067 12173 64113 12219
rect 64161 12173 64207 12219
rect 64255 12173 64301 12219
rect 64349 12173 64395 12219
rect 64443 12173 64489 12219
rect 64537 12173 64583 12219
rect 64631 12173 64677 12219
rect 64725 12173 64771 12219
rect 64819 12173 64865 12219
rect 64913 12173 64959 12219
rect 65007 12173 65053 12219
rect 65101 12173 65147 12219
rect 65195 12173 65241 12219
rect 65289 12173 65335 12219
rect 65383 12173 65429 12219
rect 65477 12173 65523 12219
rect 65571 12173 65617 12219
rect 65665 12173 65711 12219
rect 65759 12173 65805 12219
rect 65853 12173 65899 12219
rect 61717 12079 61763 12125
rect 61717 11985 61763 12031
rect 61717 11891 61763 11937
rect 61717 11797 61763 11843
rect 65853 12079 65899 12125
rect 65853 11985 65899 12031
rect 65853 11891 65899 11937
rect 65853 11797 65899 11843
rect 61717 11703 61763 11749
rect 65853 11703 65899 11749
rect 61717 11609 61763 11655
rect 61717 11515 61763 11561
rect 61717 11421 61763 11467
rect 61717 11327 61763 11373
rect 61717 11233 61763 11279
rect 61717 11139 61763 11185
rect 61717 11045 61763 11091
rect 65853 11609 65899 11655
rect 65853 11515 65899 11561
rect 65853 11421 65899 11467
rect 65853 11327 65899 11373
rect 65853 11233 65899 11279
rect 65853 11139 65899 11185
rect 61717 10951 61763 10997
rect 61717 10857 61763 10903
rect 61717 10763 61763 10809
rect 61717 10669 61763 10715
rect 65853 11045 65899 11091
rect 65853 10951 65899 10997
rect 65853 10857 65899 10903
rect 65853 10763 65899 10809
rect 65853 10669 65899 10715
rect 61717 10575 61763 10621
rect 61717 10481 61763 10527
rect 61717 10387 61763 10433
rect 61717 10293 61763 10339
rect 61717 10199 61763 10245
rect 61717 10105 61763 10151
rect 61717 10011 61763 10057
rect 65853 10575 65899 10621
rect 65853 10481 65899 10527
rect 65853 10387 65899 10433
rect 65853 10293 65899 10339
rect 65853 10199 65899 10245
rect 65853 10105 65899 10151
rect 61717 9917 61763 9963
rect 61717 9823 61763 9869
rect 61717 9729 61763 9775
rect 61717 9635 61763 9681
rect 61717 9541 61763 9587
rect 65853 10011 65899 10057
rect 65853 9917 65899 9963
rect 65853 9823 65899 9869
rect 65853 9729 65899 9775
rect 65853 9635 65899 9681
rect 61717 9447 61763 9493
rect 61717 9353 61763 9399
rect 61717 9259 61763 9305
rect 61717 9165 61763 9211
rect 61717 9071 61763 9117
rect 61717 8977 61763 9023
rect 65853 9541 65899 9587
rect 65853 9447 65899 9493
rect 65853 9353 65899 9399
rect 65853 9259 65899 9305
rect 65853 9165 65899 9211
rect 65853 9071 65899 9117
rect 65853 8977 65899 9023
rect 61717 8883 61763 8929
rect 61717 8789 61763 8835
rect 61717 8695 61763 8741
rect 61717 8601 61763 8647
rect 61717 8507 61763 8553
rect 65853 8883 65899 8929
rect 65853 8789 65899 8835
rect 65853 8695 65899 8741
rect 65853 8601 65899 8647
rect 61717 8413 61763 8459
rect 61717 8319 61763 8365
rect 61717 8225 61763 8271
rect 61717 8131 61763 8177
rect 61717 8037 61763 8083
rect 61717 7943 61763 7989
rect 65853 8507 65899 8553
rect 65853 8413 65899 8459
rect 65853 8319 65899 8365
rect 65853 8225 65899 8271
rect 65853 8131 65899 8177
rect 65853 8037 65899 8083
rect 65853 7943 65899 7989
rect 61717 7849 61763 7895
rect 61717 7755 61763 7801
rect 61717 7661 61763 7707
rect 61717 7567 61763 7613
rect 61717 7473 61763 7519
rect 65853 7849 65899 7895
rect 65853 7755 65899 7801
rect 65853 7661 65899 7707
rect 65853 7567 65899 7613
rect 65853 7473 65899 7519
rect 61717 7379 61763 7425
rect 61811 7379 61857 7425
rect 61905 7379 61951 7425
rect 61999 7379 62045 7425
rect 62093 7379 62139 7425
rect 62187 7379 62233 7425
rect 62281 7379 62327 7425
rect 62375 7379 62421 7425
rect 62469 7379 62515 7425
rect 62563 7379 62609 7425
rect 62657 7379 62703 7425
rect 62751 7379 62797 7425
rect 62845 7379 62891 7425
rect 62939 7379 62985 7425
rect 63033 7379 63079 7425
rect 63127 7379 63173 7425
rect 63221 7379 63267 7425
rect 63315 7379 63361 7425
rect 63409 7379 63455 7425
rect 63503 7379 63549 7425
rect 63597 7379 63643 7425
rect 63691 7379 63737 7425
rect 63785 7379 63831 7425
rect 63879 7379 63925 7425
rect 63973 7379 64019 7425
rect 64067 7379 64113 7425
rect 64161 7379 64207 7425
rect 64255 7379 64301 7425
rect 64349 7379 64395 7425
rect 64443 7379 64489 7425
rect 64537 7379 64583 7425
rect 64631 7379 64677 7425
rect 64725 7379 64771 7425
rect 64819 7379 64865 7425
rect 64913 7379 64959 7425
rect 65007 7379 65053 7425
rect 65101 7379 65147 7425
rect 65195 7379 65241 7425
rect 65289 7379 65335 7425
rect 65383 7379 65429 7425
rect 65477 7379 65523 7425
rect 65571 7379 65617 7425
rect 65665 7379 65711 7425
rect 65759 7379 65805 7425
rect 65853 7379 65899 7425
rect -3872 7196 -3826 7242
rect -3872 7098 -3826 7144
rect -3872 7000 -3826 7046
rect -3872 6902 -3826 6948
rect -3872 6804 -3826 6850
rect -3872 6706 -3826 6752
rect -3872 6608 -3826 6654
rect -3872 6510 -3826 6556
rect -3872 6412 -3826 6458
rect -3872 6314 -3826 6360
rect -3872 6216 -3826 6262
rect -3872 6118 -3826 6164
rect -3872 6020 -3826 6066
rect -3872 5922 -3826 5968
rect -3872 5824 -3826 5870
rect -3872 5726 -3826 5772
rect -3872 5628 -3826 5674
rect -3872 5530 -3826 5576
rect -3872 5432 -3826 5478
rect -3872 5334 -3826 5380
rect -3872 5236 -3826 5282
rect -3872 5138 -3826 5184
rect -3872 5040 -3826 5086
rect -3872 4942 -3826 4988
rect -3872 4844 -3826 4890
rect -3872 4746 -3826 4792
rect -3872 4648 -3826 4694
rect -3872 4550 -3826 4596
rect -3872 4452 -3826 4498
rect -7703 4344 -7657 4390
rect -7605 4344 -7559 4390
rect -7507 4344 -7461 4390
rect -7409 4344 -7363 4390
rect -7311 4344 -7265 4390
rect -7213 4344 -7167 4390
rect -7115 4344 -7069 4390
rect -7017 4344 -6971 4390
rect -6919 4344 -6873 4390
rect -6821 4344 -6775 4390
rect -6723 4344 -6677 4390
rect -6625 4344 -6579 4390
rect -6527 4344 -6481 4390
rect -6429 4344 -6383 4390
rect -6331 4344 -6285 4390
rect -6233 4344 -6187 4390
rect -6135 4344 -6089 4390
rect -6037 4344 -5991 4390
rect -5939 4344 -5893 4390
rect -5841 4344 -5795 4390
rect -5743 4344 -5697 4390
rect -5645 4344 -5599 4390
rect -5547 4344 -5501 4390
rect -5449 4344 -5403 4390
rect -5351 4344 -5305 4390
rect -5253 4344 -5207 4390
rect -5155 4344 -5109 4390
rect -5057 4344 -5011 4390
rect -4959 4344 -4913 4390
rect -4861 4344 -4815 4390
rect -4763 4344 -4717 4390
rect -4665 4344 -4619 4390
rect -4567 4344 -4521 4390
rect -4469 4344 -4423 4390
rect -4371 4344 -4325 4390
rect -4273 4344 -4227 4390
rect -4175 4344 -4129 4390
rect -4077 4344 -4031 4390
rect -3979 4344 -3933 4390
rect -3872 4344 -3826 4390
rect 929 4746 975 4792
rect 1023 4746 1069 4792
rect 1117 4746 1163 4792
rect 1211 4746 1257 4792
rect 1305 4746 1351 4792
rect 1399 4746 1445 4792
rect 1493 4746 1539 4792
rect 1587 4746 1633 4792
rect 1681 4746 1727 4792
rect 1775 4746 1821 4792
rect 1869 4746 1915 4792
rect 1963 4746 2009 4792
rect 2057 4746 2103 4792
rect 2151 4746 2197 4792
rect 2245 4746 2291 4792
rect 2339 4746 2385 4792
rect 2433 4746 2479 4792
rect 2527 4746 2573 4792
rect 2621 4746 2667 4792
rect 2715 4746 2761 4792
rect 2809 4746 2855 4792
rect 2903 4746 2949 4792
rect 2997 4746 3043 4792
rect 3091 4746 3137 4792
rect 3185 4746 3231 4792
rect 3279 4746 3325 4792
rect 3373 4746 3419 4792
rect 3467 4746 3513 4792
rect 3561 4746 3607 4792
rect 3655 4746 3701 4792
rect 3749 4746 3795 4792
rect 3843 4746 3889 4792
rect 3937 4746 3983 4792
rect 4031 4746 4077 4792
rect 4125 4746 4171 4792
rect 4219 4746 4265 4792
rect 4313 4746 4359 4792
rect 4407 4746 4453 4792
rect 4501 4746 4547 4792
rect 4595 4746 4641 4792
rect 4689 4746 4735 4792
rect 4783 4746 4829 4792
rect 4877 4746 4923 4792
rect 4971 4746 5017 4792
rect 929 4652 975 4698
rect 929 4558 975 4604
rect 4971 4652 5017 4698
rect 929 4464 975 4510
rect 4971 4558 5017 4604
rect 4971 4464 5017 4510
rect 929 4370 975 4416
rect 929 4276 975 4322
rect 929 4182 975 4228
rect 929 4088 975 4134
rect 929 3994 975 4040
rect 929 3900 975 3946
rect 929 3806 975 3852
rect 929 3712 975 3758
rect 929 3618 975 3664
rect 4971 4370 5017 4416
rect 4971 4276 5017 4322
rect 4971 4182 5017 4228
rect 4971 4088 5017 4134
rect 4971 3994 5017 4040
rect 4971 3900 5017 3946
rect 4971 3806 5017 3852
rect 4971 3712 5017 3758
rect 929 3524 975 3570
rect 929 3430 975 3476
rect 929 3336 975 3382
rect 929 3242 975 3288
rect 929 3148 975 3194
rect 4971 3618 5017 3664
rect 4971 3524 5017 3570
rect 4971 3430 5017 3476
rect 4971 3336 5017 3382
rect 4971 3242 5017 3288
rect 929 3054 975 3100
rect 929 2960 975 3006
rect 929 2866 975 2912
rect 929 2772 975 2818
rect 929 2678 975 2724
rect 929 2584 975 2630
rect 929 2490 975 2536
rect 929 2396 975 2442
rect 4971 3148 5017 3194
rect 4971 3054 5017 3100
rect 4971 2960 5017 3006
rect 4971 2866 5017 2912
rect 18206 5655 18252 5701
rect 18300 5655 18346 5701
rect 18394 5655 18440 5701
rect 18488 5655 18534 5701
rect 18582 5655 18628 5701
rect 18676 5655 18722 5701
rect 18770 5655 18816 5701
rect 18864 5655 18910 5701
rect 18958 5655 19004 5701
rect 19052 5655 19098 5701
rect 19146 5655 19192 5701
rect 19240 5655 19286 5701
rect 19334 5655 19380 5701
rect 19428 5655 19474 5701
rect 19522 5655 19568 5701
rect 19616 5655 19662 5701
rect 19710 5655 19756 5701
rect 19804 5655 19850 5701
rect 19898 5655 19944 5701
rect 19992 5655 20038 5701
rect 20086 5655 20132 5701
rect 20180 5655 20226 5701
rect 20274 5655 20320 5701
rect 20368 5655 20414 5701
rect 20462 5655 20508 5701
rect 20556 5655 20602 5701
rect 20650 5655 20696 5701
rect 20744 5655 20790 5701
rect 20838 5655 20884 5701
rect 20932 5655 20978 5701
rect 21026 5655 21072 5701
rect 21120 5655 21166 5701
rect 21214 5655 21260 5701
rect 21308 5655 21354 5701
rect 21402 5655 21448 5701
rect 21496 5655 21542 5701
rect 21590 5655 21636 5701
rect 21684 5655 21730 5701
rect 21778 5655 21824 5701
rect 21872 5655 21918 5701
rect 21966 5655 22012 5701
rect 22060 5655 22106 5701
rect 22154 5655 22200 5701
rect 22248 5655 22294 5701
rect 22342 5655 22388 5701
rect 22436 5655 22482 5701
rect 22530 5655 22576 5701
rect 22624 5655 22670 5701
rect 22718 5655 22764 5701
rect 22812 5655 22858 5701
rect 22906 5655 22952 5701
rect 23000 5655 23046 5701
rect 23094 5655 23140 5701
rect 23188 5655 23234 5701
rect 23282 5655 23328 5701
rect 23376 5655 23422 5701
rect 23470 5655 23516 5701
rect 23564 5655 23610 5701
rect 23658 5655 23704 5701
rect 23752 5655 23798 5701
rect 23846 5655 23892 5701
rect 23940 5655 23986 5701
rect 24034 5655 24080 5701
rect 24128 5655 24174 5701
rect 24222 5655 24268 5701
rect 24316 5655 24362 5701
rect 24410 5655 24456 5701
rect 24504 5655 24550 5701
rect 24598 5655 24644 5701
rect 24692 5655 24738 5701
rect 24786 5655 24832 5701
rect 24880 5655 24926 5701
rect 24974 5655 25020 5701
rect 25068 5655 25114 5701
rect 25162 5655 25208 5701
rect 25256 5655 25302 5701
rect 25350 5655 25396 5701
rect 25444 5655 25490 5701
rect 25538 5655 25584 5701
rect 25632 5655 25678 5701
rect 25726 5655 25772 5701
rect 25820 5655 25866 5701
rect 25914 5655 25960 5701
rect 26008 5655 26054 5701
rect 26102 5655 26148 5701
rect 26196 5655 26242 5701
rect 26290 5655 26336 5701
rect 26384 5655 26430 5701
rect 26478 5655 26524 5701
rect 26572 5655 26618 5701
rect 26666 5655 26712 5701
rect 26760 5655 26806 5701
rect 26854 5655 26900 5701
rect 26948 5655 26994 5701
rect 27042 5655 27088 5701
rect 27136 5655 27182 5701
rect 27230 5655 27276 5701
rect 27324 5655 27370 5701
rect 27418 5655 27464 5701
rect 27512 5655 27558 5701
rect 27606 5655 27652 5701
rect 27700 5655 27746 5701
rect 27794 5655 27840 5701
rect 27888 5655 27934 5701
rect 27982 5655 28028 5701
rect 28076 5655 28122 5701
rect 28170 5655 28216 5701
rect 28264 5655 28310 5701
rect 28358 5655 28404 5701
rect 28452 5655 28498 5701
rect 28546 5655 28592 5701
rect 28640 5655 28686 5701
rect 28734 5655 28780 5701
rect 28828 5655 28874 5701
rect 28922 5655 28968 5701
rect 29016 5655 29062 5701
rect 29110 5655 29156 5701
rect 29204 5655 29250 5701
rect 29298 5655 29344 5701
rect 29392 5655 29438 5701
rect 29486 5655 29532 5701
rect 29580 5655 29626 5701
rect 29674 5655 29720 5701
rect 29768 5655 29814 5701
rect 29862 5655 29908 5701
rect 29956 5655 30002 5701
rect 30050 5655 30096 5701
rect 30144 5655 30190 5701
rect 30238 5655 30284 5701
rect 30332 5655 30378 5701
rect 30426 5655 30472 5701
rect 30520 5655 30566 5701
rect 30614 5655 30660 5701
rect 30708 5655 30754 5701
rect 30802 5655 30848 5701
rect 30896 5655 30942 5701
rect 30990 5655 31036 5701
rect 31084 5655 31130 5701
rect 31178 5655 31224 5701
rect 31272 5655 31318 5701
rect 31366 5655 31412 5701
rect 31460 5655 31506 5701
rect 31554 5655 31600 5701
rect 31648 5655 31694 5701
rect 31742 5655 31788 5701
rect 18206 5561 18252 5607
rect 18206 5467 18252 5513
rect 18206 5373 18252 5419
rect 18206 5279 18252 5325
rect 18206 5185 18252 5231
rect 18206 5091 18252 5137
rect 18206 4997 18252 5043
rect 18206 4903 18252 4949
rect 23000 5561 23046 5607
rect 23000 5467 23046 5513
rect 23000 5373 23046 5419
rect 23000 5279 23046 5325
rect 23000 5185 23046 5231
rect 23000 5091 23046 5137
rect 28734 5561 28780 5607
rect 28734 5467 28780 5513
rect 28734 5373 28780 5419
rect 28734 5279 28780 5325
rect 31742 5561 31788 5607
rect 31742 5467 31788 5513
rect 31742 5373 31788 5419
rect 31742 5279 31788 5325
rect 28734 5185 28780 5231
rect 28734 5091 28780 5137
rect 23000 4997 23046 5043
rect 18206 4809 18252 4855
rect 23000 4903 23046 4949
rect 23000 4809 23046 4855
rect 18206 4715 18252 4761
rect 18206 4621 18252 4667
rect 18206 4527 18252 4573
rect 4971 2772 5017 2818
rect 4971 2678 5017 2724
rect 4971 2584 5017 2630
rect 4971 2490 5017 2536
rect 4971 2396 5017 2442
rect 929 2302 975 2348
rect 929 2208 975 2254
rect 929 2114 975 2160
rect 929 2020 975 2066
rect 929 1926 975 1972
rect 4971 2302 5017 2348
rect 4971 2208 5017 2254
rect 4971 2114 5017 2160
rect 4971 2020 5017 2066
rect 4971 1926 5017 1972
rect 929 1832 975 1878
rect 4971 1832 5017 1878
rect 929 1738 975 1784
rect 4971 1738 5017 1784
rect 929 1644 975 1690
rect 929 1550 975 1596
rect 4971 1644 5017 1690
rect 4971 1550 5017 1596
rect 929 1456 975 1502
rect 1023 1456 1069 1502
rect 1117 1456 1163 1502
rect 1211 1456 1257 1502
rect 1305 1456 1351 1502
rect 1399 1456 1445 1502
rect 1493 1456 1539 1502
rect 1587 1456 1633 1502
rect 1681 1456 1727 1502
rect 1775 1456 1821 1502
rect 1869 1456 1915 1502
rect 1963 1456 2009 1502
rect 2057 1456 2103 1502
rect 2151 1456 2197 1502
rect 2245 1456 2291 1502
rect 2339 1456 2385 1502
rect 2433 1456 2479 1502
rect 2527 1456 2573 1502
rect 2621 1456 2667 1502
rect 2715 1456 2761 1502
rect 2809 1456 2855 1502
rect 2903 1456 2949 1502
rect 2997 1456 3043 1502
rect 3091 1456 3137 1502
rect 3185 1456 3231 1502
rect 3279 1456 3325 1502
rect 3373 1456 3419 1502
rect 3467 1456 3513 1502
rect 3561 1456 3607 1502
rect 3655 1456 3701 1502
rect 3749 1456 3795 1502
rect 3843 1456 3889 1502
rect 3937 1456 3983 1502
rect 4031 1456 4077 1502
rect 4125 1456 4171 1502
rect 4219 1456 4265 1502
rect 4313 1456 4359 1502
rect 4407 1456 4453 1502
rect 4501 1456 4547 1502
rect 4595 1456 4641 1502
rect 4689 1456 4735 1502
rect 4783 1456 4829 1502
rect 4877 1456 4923 1502
rect 4971 1456 5017 1502
rect 18206 4433 18252 4479
rect 18206 4339 18252 4385
rect 18206 4245 18252 4291
rect 18206 4151 18252 4197
rect 23000 4715 23046 4761
rect 23000 4621 23046 4667
rect 23000 4527 23046 4573
rect 23000 4433 23046 4479
rect 23000 4339 23046 4385
rect 23000 4245 23046 4291
rect 18206 4057 18252 4103
rect 23000 4151 23046 4197
rect 23000 4057 23046 4103
rect 18206 3963 18252 4009
rect 18206 3869 18252 3915
rect 18206 3775 18252 3821
rect 18206 3681 18252 3727
rect 18206 3587 18252 3633
rect 18206 3493 18252 3539
rect 18206 3399 18252 3445
rect 23000 3963 23046 4009
rect 23000 3869 23046 3915
rect 23000 3775 23046 3821
rect 23000 3681 23046 3727
rect 23000 3587 23046 3633
rect 28734 4997 28780 5043
rect 28734 4903 28780 4949
rect 28734 4809 28780 4855
rect 28734 4715 28780 4761
rect 28734 4621 28780 4667
rect 28734 4527 28780 4573
rect 28734 4433 28780 4479
rect 28734 4339 28780 4385
rect 28734 4245 28780 4291
rect 28734 4151 28780 4197
rect 28734 4057 28780 4103
rect 28734 3963 28780 4009
rect 28734 3869 28780 3915
rect 28734 3775 28780 3821
rect 28734 3681 28780 3727
rect 28734 3587 28780 3633
rect 23000 3493 23046 3539
rect 18206 3305 18252 3351
rect 23000 3399 23046 3445
rect 18206 3211 18252 3257
rect 18206 3117 18252 3163
rect 18206 3023 18252 3069
rect 18206 2929 18252 2975
rect 18206 2835 18252 2881
rect 18206 2741 18252 2787
rect 23000 3305 23046 3351
rect 23000 3211 23046 3257
rect 23000 3117 23046 3163
rect 28734 3493 28780 3539
rect 31742 5185 31788 5231
rect 31742 5091 31788 5137
rect 31742 4997 31788 5043
rect 31742 4903 31788 4949
rect 31742 4809 31788 4855
rect 31742 4715 31788 4761
rect 31742 4621 31788 4667
rect 31742 4527 31788 4573
rect 31742 4433 31788 4479
rect 31742 4339 31788 4385
rect 31742 4245 31788 4291
rect 31742 4151 31788 4197
rect 31742 4057 31788 4103
rect 31742 3963 31788 4009
rect 31742 3869 31788 3915
rect 31742 3775 31788 3821
rect 31742 3681 31788 3727
rect 31742 3587 31788 3633
rect 28734 3399 28780 3445
rect 28734 3305 28780 3351
rect 28734 3211 28780 3257
rect 31742 3493 31788 3539
rect 31742 3399 31788 3445
rect 31742 3305 31788 3351
rect 28734 3117 28780 3163
rect 23000 3023 23046 3069
rect 23000 2929 23046 2975
rect 23000 2835 23046 2881
rect 23000 2741 23046 2787
rect 18206 2647 18252 2693
rect 18206 2553 18252 2599
rect 18206 2459 18252 2505
rect 18206 2365 18252 2411
rect 18206 2271 18252 2317
rect 18206 2177 18252 2223
rect 18206 2083 18252 2129
rect 18206 1989 18252 2035
rect 23000 2647 23046 2693
rect 23000 2553 23046 2599
rect 23000 2459 23046 2505
rect 23000 2365 23046 2411
rect 23000 2271 23046 2317
rect 23000 2177 23046 2223
rect 23000 2083 23046 2129
rect 23000 1989 23046 2035
rect 18206 1895 18252 1941
rect 18206 1801 18252 1847
rect 23000 1895 23046 1941
rect 18206 1707 18252 1753
rect 18206 1613 18252 1659
rect 18206 1519 18252 1565
rect 18206 1425 18252 1471
rect 18206 1331 18252 1377
rect 18206 1237 18252 1283
rect 18206 1143 18252 1189
rect 23000 1801 23046 1847
rect 23000 1707 23046 1753
rect 23000 1613 23046 1659
rect 28734 3023 28780 3069
rect 28734 2929 28780 2975
rect 28734 2835 28780 2881
rect 28734 2741 28780 2787
rect 28734 2647 28780 2693
rect 28734 2553 28780 2599
rect 28734 2459 28780 2505
rect 28734 2365 28780 2411
rect 28734 2271 28780 2317
rect 28734 2177 28780 2223
rect 28734 2083 28780 2129
rect 28734 1989 28780 2035
rect 28734 1895 28780 1941
rect 28734 1801 28780 1847
rect 28734 1707 28780 1753
rect 28734 1613 28780 1659
rect 23000 1519 23046 1565
rect 23000 1425 23046 1471
rect 23000 1331 23046 1377
rect 23000 1237 23046 1283
rect 23000 1143 23046 1189
rect 28734 1519 28780 1565
rect 31742 3211 31788 3257
rect 31742 3117 31788 3163
rect 31742 3023 31788 3069
rect 31742 2929 31788 2975
rect 31742 2835 31788 2881
rect 31742 2741 31788 2787
rect 31742 2647 31788 2693
rect 31742 2553 31788 2599
rect 31742 2459 31788 2505
rect 31742 2365 31788 2411
rect 31742 2271 31788 2317
rect 31742 2177 31788 2223
rect 31742 2083 31788 2129
rect 31742 1989 31788 2035
rect 31742 1895 31788 1941
rect 31742 1801 31788 1847
rect 31742 1707 31788 1753
rect 31742 1613 31788 1659
rect 31742 1519 31788 1565
rect 28734 1425 28780 1471
rect 28734 1331 28780 1377
rect 28734 1237 28780 1283
rect 28734 1143 28780 1189
rect 31742 1425 31788 1471
rect 31742 1331 31788 1377
rect 31742 1237 31788 1283
rect 31742 1143 31788 1189
rect 18206 1049 18252 1095
rect 18300 1049 18346 1095
rect 18394 1049 18440 1095
rect 18488 1049 18534 1095
rect 18582 1049 18628 1095
rect 18676 1049 18722 1095
rect 18770 1049 18816 1095
rect 18864 1049 18910 1095
rect 18958 1049 19004 1095
rect 19052 1049 19098 1095
rect 19146 1049 19192 1095
rect 19240 1049 19286 1095
rect 19334 1049 19380 1095
rect 19428 1049 19474 1095
rect 19522 1049 19568 1095
rect 19616 1049 19662 1095
rect 19710 1049 19756 1095
rect 19804 1049 19850 1095
rect 19898 1049 19944 1095
rect 19992 1049 20038 1095
rect 20086 1049 20132 1095
rect 20180 1049 20226 1095
rect 20274 1049 20320 1095
rect 20368 1049 20414 1095
rect 20462 1049 20508 1095
rect 20556 1049 20602 1095
rect 20650 1049 20696 1095
rect 20744 1049 20790 1095
rect 20838 1049 20884 1095
rect 20932 1049 20978 1095
rect 21026 1049 21072 1095
rect 21120 1049 21166 1095
rect 21214 1049 21260 1095
rect 21308 1049 21354 1095
rect 21402 1049 21448 1095
rect 21496 1049 21542 1095
rect 21590 1049 21636 1095
rect 21684 1049 21730 1095
rect 21778 1049 21824 1095
rect 21872 1049 21918 1095
rect 21966 1049 22012 1095
rect 22060 1049 22106 1095
rect 22154 1049 22200 1095
rect 22248 1049 22294 1095
rect 22342 1049 22388 1095
rect 22436 1049 22482 1095
rect 22530 1049 22576 1095
rect 22624 1049 22670 1095
rect 22718 1049 22764 1095
rect 22812 1049 22858 1095
rect 22906 1049 22952 1095
rect 23000 1049 23046 1095
rect 23094 1049 23140 1095
rect 23188 1049 23234 1095
rect 23282 1049 23328 1095
rect 23376 1049 23422 1095
rect 23470 1049 23516 1095
rect 23564 1049 23610 1095
rect 23658 1049 23704 1095
rect 23752 1049 23798 1095
rect 23846 1049 23892 1095
rect 23940 1049 23986 1095
rect 24034 1049 24080 1095
rect 24128 1049 24174 1095
rect 24222 1049 24268 1095
rect 24316 1049 24362 1095
rect 24410 1049 24456 1095
rect 24504 1049 24550 1095
rect 24598 1049 24644 1095
rect 24692 1049 24738 1095
rect 24786 1049 24832 1095
rect 24880 1049 24926 1095
rect 24974 1049 25020 1095
rect 25068 1049 25114 1095
rect 25162 1049 25208 1095
rect 25256 1049 25302 1095
rect 25350 1049 25396 1095
rect 25444 1049 25490 1095
rect 25538 1049 25584 1095
rect 25632 1049 25678 1095
rect 25726 1049 25772 1095
rect 25820 1049 25866 1095
rect 25914 1049 25960 1095
rect 26008 1049 26054 1095
rect 26102 1049 26148 1095
rect 26196 1049 26242 1095
rect 26290 1049 26336 1095
rect 26384 1049 26430 1095
rect 26478 1049 26524 1095
rect 26572 1049 26618 1095
rect 26666 1049 26712 1095
rect 26760 1049 26806 1095
rect 26854 1049 26900 1095
rect 26948 1049 26994 1095
rect 27042 1049 27088 1095
rect 27136 1049 27182 1095
rect 27230 1049 27276 1095
rect 27324 1049 27370 1095
rect 27418 1049 27464 1095
rect 27512 1049 27558 1095
rect 27606 1049 27652 1095
rect 27700 1049 27746 1095
rect 27794 1049 27840 1095
rect 27888 1049 27934 1095
rect 27982 1049 28028 1095
rect 28076 1049 28122 1095
rect 28170 1049 28216 1095
rect 28264 1049 28310 1095
rect 28358 1049 28404 1095
rect 28452 1049 28498 1095
rect 28546 1049 28592 1095
rect 28640 1049 28686 1095
rect 28734 1049 28780 1095
rect 28828 1049 28874 1095
rect 28922 1049 28968 1095
rect 29016 1049 29062 1095
rect 29110 1049 29156 1095
rect 29204 1049 29250 1095
rect 29298 1049 29344 1095
rect 29392 1049 29438 1095
rect 29486 1049 29532 1095
rect 29580 1049 29626 1095
rect 29674 1049 29720 1095
rect 29768 1049 29814 1095
rect 29862 1049 29908 1095
rect 29956 1049 30002 1095
rect 30050 1049 30096 1095
rect 30144 1049 30190 1095
rect 30238 1049 30284 1095
rect 30332 1049 30378 1095
rect 30426 1049 30472 1095
rect 30520 1049 30566 1095
rect 30614 1049 30660 1095
rect 30708 1049 30754 1095
rect 30802 1049 30848 1095
rect 30896 1049 30942 1095
rect 30990 1049 31036 1095
rect 31084 1049 31130 1095
rect 31178 1049 31224 1095
rect 31272 1049 31318 1095
rect 31366 1049 31412 1095
rect 31460 1049 31506 1095
rect 31554 1049 31600 1095
rect 31648 1049 31694 1095
rect 31742 1049 31788 1095
<< polysilicon >>
rect 3952 14219 4024 14232
rect 3952 14173 3965 14219
rect 4011 14173 4024 14219
rect 3952 14160 4024 14173
rect 4432 14219 4504 14232
rect 4432 14173 4445 14219
rect 4491 14173 4504 14219
rect 4432 14160 4504 14173
rect 5072 14219 5144 14232
rect 5072 14173 5085 14219
rect 5131 14173 5144 14219
rect 5072 14160 5144 14173
rect 3672 14026 3728 14070
rect 3960 14026 4016 14160
rect 4440 14102 4496 14160
rect 4120 14026 4176 14070
rect 4280 14026 4336 14070
rect 4440 14046 4656 14102
rect 4440 14026 4496 14046
rect 4600 14026 4656 14046
rect 4760 14026 4816 14070
rect 4920 14026 4976 14070
rect 5080 14026 5136 14160
rect 5368 14026 5424 14070
rect 3672 12896 3728 13276
rect 3960 13232 4016 13276
rect 4120 13256 4176 13276
rect 4280 13256 4336 13276
rect 4120 13200 4336 13256
rect 4440 13232 4496 13276
rect 4600 13232 4656 13276
rect 4760 13256 4816 13276
rect 4920 13256 4976 13276
rect 4760 13200 4976 13256
rect 5080 13232 5136 13276
rect 4120 13104 4176 13200
rect 4760 13104 4816 13200
rect 3952 13091 4024 13104
rect 3952 13045 3965 13091
rect 4011 13045 4024 13091
rect 3952 13032 4024 13045
rect 4112 13091 4184 13104
rect 4112 13045 4125 13091
rect 4171 13045 4184 13091
rect 4112 13032 4184 13045
rect 4432 13091 4504 13104
rect 4432 13045 4445 13091
rect 4491 13045 4504 13091
rect 4432 13032 4504 13045
rect 4752 13091 4824 13104
rect 4752 13045 4765 13091
rect 4811 13045 4824 13091
rect 4752 13032 4824 13045
rect 5072 13091 5144 13104
rect 5072 13045 5085 13091
rect 5131 13045 5144 13091
rect 5072 13032 5144 13045
rect 3960 12896 4016 13032
rect 4440 12972 4496 13032
rect 4120 12896 4176 12940
rect 4280 12896 4336 12940
rect 4440 12916 4656 12972
rect 4440 12896 4496 12916
rect 4600 12896 4656 12916
rect 4760 12896 4816 12940
rect 4920 12896 4976 12940
rect 5080 12896 5136 13032
rect 5368 12896 5424 13276
rect 3672 11766 3728 12146
rect 3960 12102 4016 12146
rect 4120 12126 4176 12146
rect 4280 12126 4336 12146
rect 4120 12070 4336 12126
rect 4440 12102 4496 12146
rect 4600 12102 4656 12146
rect 4760 12126 4816 12146
rect 4920 12126 4976 12146
rect 4760 12070 4976 12126
rect 5080 12102 5136 12146
rect 4120 11976 4176 12070
rect 4760 11976 4816 12070
rect 3952 11963 4024 11976
rect 3952 11917 3965 11963
rect 4011 11917 4024 11963
rect 3952 11902 4024 11917
rect 4112 11963 4184 11976
rect 4112 11917 4125 11963
rect 4171 11917 4184 11963
rect 4112 11904 4184 11917
rect 4432 11963 4504 11976
rect 4432 11917 4445 11963
rect 4491 11917 4504 11963
rect 4432 11902 4504 11917
rect 4752 11963 4824 11976
rect 4752 11917 4765 11963
rect 4811 11917 4824 11963
rect 4752 11904 4824 11917
rect 5072 11963 5144 11976
rect 5072 11917 5085 11963
rect 5131 11917 5144 11963
rect 5072 11902 5144 11917
rect 3960 11766 4016 11902
rect 4440 11842 4496 11902
rect 4120 11766 4176 11810
rect 4280 11766 4336 11810
rect 4440 11786 4656 11842
rect 4440 11766 4496 11786
rect 4600 11766 4656 11786
rect 4760 11766 4816 11810
rect 4920 11766 4976 11810
rect 5080 11766 5136 11902
rect 5368 11766 5424 12146
rect -7386 10356 -7186 10369
rect -7386 10310 -7373 10356
rect -7199 10310 -7186 10356
rect -7386 10267 -7186 10310
rect -7386 9764 -7186 9807
rect -7386 9718 -7373 9764
rect -7199 9718 -7186 9764
rect -7386 9705 -7186 9718
rect -7106 10356 -6906 10369
rect -7106 10310 -7093 10356
rect -6919 10310 -6906 10356
rect -7106 10267 -6906 10310
rect -7106 9764 -6906 9807
rect -7106 9718 -7093 9764
rect -6919 9718 -6906 9764
rect -7106 9705 -6906 9718
rect -6826 10356 -6626 10369
rect -6826 10310 -6813 10356
rect -6639 10310 -6626 10356
rect -6826 10267 -6626 10310
rect -6826 9764 -6626 9807
rect -6826 9718 -6813 9764
rect -6639 9718 -6626 9764
rect -6826 9705 -6626 9718
rect -6546 10356 -6346 10369
rect -6546 10310 -6533 10356
rect -6359 10310 -6346 10356
rect -6546 10267 -6346 10310
rect -6546 9764 -6346 9807
rect -6546 9718 -6533 9764
rect -6359 9718 -6346 9764
rect -6546 9705 -6346 9718
rect -6266 10356 -6066 10369
rect -6266 10310 -6253 10356
rect -6079 10310 -6066 10356
rect -6266 10267 -6066 10310
rect -6266 9764 -6066 9807
rect -6266 9718 -6253 9764
rect -6079 9718 -6066 9764
rect -6266 9705 -6066 9718
rect -5986 10356 -5786 10369
rect -5986 10310 -5973 10356
rect -5799 10310 -5786 10356
rect -5986 10267 -5786 10310
rect -5986 9764 -5786 9807
rect -5986 9718 -5973 9764
rect -5799 9718 -5786 9764
rect -5986 9705 -5786 9718
rect -5706 10356 -5506 10369
rect -5706 10310 -5693 10356
rect -5519 10310 -5506 10356
rect -5706 10267 -5506 10310
rect -5706 9764 -5506 9807
rect -5706 9718 -5693 9764
rect -5519 9718 -5506 9764
rect -5706 9705 -5506 9718
rect -5426 10356 -5226 10369
rect -5426 10310 -5413 10356
rect -5239 10310 -5226 10356
rect -5426 10267 -5226 10310
rect -5426 9764 -5226 9807
rect -5426 9718 -5413 9764
rect -5239 9718 -5226 9764
rect -5426 9705 -5226 9718
rect -5146 10356 -4946 10369
rect -5146 10310 -5133 10356
rect -4959 10310 -4946 10356
rect -5146 10267 -4946 10310
rect -5146 9764 -4946 9807
rect -5146 9718 -5133 9764
rect -4959 9718 -4946 9764
rect -5146 9705 -4946 9718
rect -4866 10356 -4666 10369
rect -4866 10310 -4853 10356
rect -4679 10310 -4666 10356
rect -4866 10267 -4666 10310
rect -4866 9764 -4666 9807
rect -4866 9718 -4853 9764
rect -4679 9718 -4666 9764
rect -4866 9705 -4666 9718
rect -4586 10356 -4386 10369
rect -4586 10310 -4573 10356
rect -4399 10310 -4386 10356
rect -4586 10267 -4386 10310
rect -4586 9764 -4386 9807
rect -4586 9718 -4573 9764
rect -4399 9718 -4386 9764
rect -4586 9705 -4386 9718
rect -4306 10356 -4106 10369
rect -4306 10310 -4293 10356
rect -4119 10310 -4106 10356
rect -4306 10267 -4106 10310
rect -4306 9764 -4106 9807
rect -4306 9718 -4293 9764
rect -4119 9718 -4106 9764
rect -4306 9705 -4106 9718
rect -7386 9439 -7186 9452
rect -7386 9393 -7373 9439
rect -7199 9393 -7186 9439
rect -7386 9350 -7186 9393
rect -7386 8847 -7186 8890
rect -7386 8801 -7373 8847
rect -7199 8801 -7186 8847
rect -7386 8788 -7186 8801
rect -7106 9439 -6906 9452
rect -7106 9393 -7093 9439
rect -6919 9393 -6906 9439
rect -7106 9350 -6906 9393
rect -7106 8847 -6906 8890
rect -7106 8801 -7093 8847
rect -6919 8801 -6906 8847
rect -7106 8788 -6906 8801
rect -6826 9439 -6626 9452
rect -6826 9393 -6813 9439
rect -6639 9393 -6626 9439
rect -6826 9350 -6626 9393
rect -6826 8847 -6626 8890
rect -6826 8801 -6813 8847
rect -6639 8801 -6626 8847
rect -6826 8788 -6626 8801
rect -6546 9439 -6346 9452
rect -6546 9393 -6533 9439
rect -6359 9393 -6346 9439
rect -6546 9350 -6346 9393
rect -6546 8847 -6346 8890
rect -6546 8801 -6533 8847
rect -6359 8801 -6346 8847
rect -6546 8788 -6346 8801
rect -6266 9439 -6066 9452
rect -6266 9393 -6253 9439
rect -6079 9393 -6066 9439
rect -6266 9350 -6066 9393
rect -6266 8847 -6066 8890
rect -6266 8801 -6253 8847
rect -6079 8801 -6066 8847
rect -6266 8788 -6066 8801
rect -5986 9439 -5786 9452
rect -5986 9393 -5973 9439
rect -5799 9393 -5786 9439
rect -5986 9350 -5786 9393
rect -5986 8847 -5786 8890
rect -5986 8801 -5973 8847
rect -5799 8801 -5786 8847
rect -5986 8788 -5786 8801
rect -5706 9439 -5506 9452
rect -5706 9393 -5693 9439
rect -5519 9393 -5506 9439
rect -5706 9350 -5506 9393
rect -5706 8847 -5506 8890
rect -5706 8801 -5693 8847
rect -5519 8801 -5506 8847
rect -5706 8788 -5506 8801
rect -5426 9439 -5226 9452
rect -5426 9393 -5413 9439
rect -5239 9393 -5226 9439
rect -5426 9350 -5226 9393
rect -5426 8847 -5226 8890
rect -5426 8801 -5413 8847
rect -5239 8801 -5226 8847
rect -5426 8788 -5226 8801
rect -5146 9439 -4946 9452
rect -5146 9393 -5133 9439
rect -4959 9393 -4946 9439
rect -5146 9350 -4946 9393
rect -5146 8847 -4946 8890
rect -5146 8801 -5133 8847
rect -4959 8801 -4946 8847
rect -5146 8788 -4946 8801
rect -4866 9439 -4666 9452
rect -4866 9393 -4853 9439
rect -4679 9393 -4666 9439
rect -4866 9350 -4666 9393
rect -4866 8847 -4666 8890
rect -4866 8801 -4853 8847
rect -4679 8801 -4666 8847
rect -4866 8788 -4666 8801
rect -4586 9439 -4386 9452
rect -4586 9393 -4573 9439
rect -4399 9393 -4386 9439
rect -4586 9350 -4386 9393
rect -4586 8847 -4386 8890
rect -4586 8801 -4573 8847
rect -4399 8801 -4386 8847
rect -4586 8788 -4386 8801
rect -4306 9439 -4106 9452
rect -4306 9393 -4293 9439
rect -4119 9393 -4106 9439
rect -4306 9350 -4106 9393
rect -4306 8847 -4106 8890
rect -4306 8801 -4293 8847
rect -4119 8801 -4106 8847
rect -4306 8788 -4106 8801
rect -7386 8522 -7186 8535
rect -7386 8476 -7373 8522
rect -7199 8476 -7186 8522
rect -7386 8433 -7186 8476
rect -7386 7930 -7186 7973
rect -7386 7884 -7373 7930
rect -7199 7884 -7186 7930
rect -7386 7871 -7186 7884
rect -7106 8522 -6906 8535
rect -7106 8476 -7093 8522
rect -6919 8476 -6906 8522
rect -7106 8433 -6906 8476
rect -7106 7930 -6906 7973
rect -7106 7884 -7093 7930
rect -6919 7884 -6906 7930
rect -7106 7871 -6906 7884
rect -6826 8522 -6626 8535
rect -6826 8476 -6813 8522
rect -6639 8476 -6626 8522
rect -6826 8433 -6626 8476
rect -6826 7930 -6626 7973
rect -6826 7884 -6813 7930
rect -6639 7884 -6626 7930
rect -6826 7871 -6626 7884
rect -6546 8522 -6346 8535
rect -6546 8476 -6533 8522
rect -6359 8476 -6346 8522
rect -6546 8433 -6346 8476
rect -6546 7930 -6346 7973
rect -6546 7884 -6533 7930
rect -6359 7884 -6346 7930
rect -6546 7871 -6346 7884
rect -6266 8522 -6066 8535
rect -6266 8476 -6253 8522
rect -6079 8476 -6066 8522
rect -6266 8433 -6066 8476
rect -6266 7930 -6066 7973
rect -6266 7884 -6253 7930
rect -6079 7884 -6066 7930
rect -6266 7871 -6066 7884
rect -5986 8522 -5786 8535
rect -5986 8476 -5973 8522
rect -5799 8476 -5786 8522
rect -5986 8433 -5786 8476
rect -5986 7930 -5786 7973
rect -5986 7884 -5973 7930
rect -5799 7884 -5786 7930
rect -5986 7871 -5786 7884
rect -5706 8522 -5506 8535
rect -5706 8476 -5693 8522
rect -5519 8476 -5506 8522
rect -5706 8433 -5506 8476
rect -5706 7930 -5506 7973
rect -5706 7884 -5693 7930
rect -5519 7884 -5506 7930
rect -5706 7871 -5506 7884
rect -5426 8522 -5226 8535
rect -5426 8476 -5413 8522
rect -5239 8476 -5226 8522
rect -5426 8433 -5226 8476
rect -5426 7930 -5226 7973
rect -5426 7884 -5413 7930
rect -5239 7884 -5226 7930
rect -5426 7871 -5226 7884
rect -5146 8522 -4946 8535
rect -5146 8476 -5133 8522
rect -4959 8476 -4946 8522
rect -5146 8433 -4946 8476
rect -5146 7930 -4946 7973
rect -5146 7884 -5133 7930
rect -4959 7884 -4946 7930
rect -5146 7871 -4946 7884
rect -4866 8522 -4666 8535
rect -4866 8476 -4853 8522
rect -4679 8476 -4666 8522
rect -4866 8433 -4666 8476
rect -4866 7930 -4666 7973
rect -4866 7884 -4853 7930
rect -4679 7884 -4666 7930
rect -4866 7871 -4666 7884
rect -4586 8522 -4386 8535
rect -4586 8476 -4573 8522
rect -4399 8476 -4386 8522
rect -4586 8433 -4386 8476
rect -4586 7930 -4386 7973
rect -4586 7884 -4573 7930
rect -4399 7884 -4386 7930
rect -4586 7871 -4386 7884
rect -4306 8522 -4106 8535
rect -4306 8476 -4293 8522
rect -4119 8476 -4106 8522
rect -4306 8433 -4106 8476
rect -4306 7930 -4106 7973
rect -4306 7884 -4293 7930
rect -4119 7884 -4106 7930
rect -4306 7871 -4106 7884
rect 3672 10636 3728 11016
rect 3960 10636 4016 11016
rect 4120 10636 4176 11016
rect 4280 10636 4336 11016
rect 4440 10636 4496 11016
rect 4600 10636 4656 11016
rect 4760 10636 4816 11016
rect 4920 10636 4976 11016
rect 5080 10636 5136 11016
rect 5368 10636 5424 11016
rect 986 10558 1098 10602
rect 1202 10558 1314 10602
rect 1418 10558 1530 10602
rect 1634 10558 1746 10602
rect 1850 10558 1962 10602
rect 2066 10558 2178 10602
rect 2282 10558 2394 10602
rect 2498 10558 2610 10602
rect 2714 10558 2826 10602
rect 2930 10558 3042 10602
rect 986 9796 1098 9932
rect 1202 9796 1314 9932
rect 1418 9796 1530 9932
rect 1634 9796 1746 9932
rect 1850 9796 1962 9932
rect 2066 9796 2178 9932
rect 2282 9796 2394 9932
rect 2498 9796 2610 9932
rect 2714 9796 2826 9932
rect 2930 9796 3042 9932
rect 3672 9506 3728 9886
rect 3960 9842 4016 9886
rect 4120 9866 4176 9886
rect 4280 9866 4336 9886
rect 4120 9810 4336 9866
rect 4440 9842 4496 9886
rect 4600 9842 4656 9886
rect 4760 9866 4816 9886
rect 4920 9866 4976 9886
rect 4760 9810 4976 9866
rect 5080 9842 5136 9886
rect 4120 9716 4176 9810
rect 4760 9716 4816 9810
rect 3952 9703 4024 9716
rect 3952 9657 3965 9703
rect 4011 9657 4024 9703
rect 3952 9642 4024 9657
rect 4112 9703 4184 9716
rect 4112 9657 4125 9703
rect 4171 9657 4184 9703
rect 4112 9644 4184 9657
rect 4432 9703 4504 9716
rect 4432 9657 4445 9703
rect 4491 9657 4504 9703
rect 4432 9642 4504 9657
rect 4752 9703 4824 9716
rect 4752 9657 4765 9703
rect 4811 9657 4824 9703
rect 4752 9644 4824 9657
rect 5072 9703 5144 9716
rect 5072 9657 5085 9703
rect 5131 9657 5144 9703
rect 5072 9642 5144 9657
rect 3960 9506 4016 9642
rect 4440 9582 4496 9642
rect 4120 9506 4176 9550
rect 4280 9506 4336 9550
rect 4440 9526 4656 9582
rect 4440 9506 4496 9526
rect 4600 9506 4656 9526
rect 4760 9506 4816 9550
rect 4920 9506 4976 9550
rect 5080 9506 5136 9642
rect 5368 9506 5424 9886
rect 986 9034 1098 9170
rect 1202 9034 1314 9170
rect 1418 9034 1530 9170
rect 1634 9034 1746 9170
rect 1850 9034 1962 9170
rect 2066 9034 2178 9170
rect 2282 9034 2394 9170
rect 2498 9034 2610 9170
rect 2714 9034 2826 9170
rect 2930 9034 3042 9170
rect 3672 8602 3728 8756
rect 3960 8712 4016 8756
rect 4120 8736 4176 8756
rect 4280 8736 4336 8756
rect 4120 8680 4336 8736
rect 4440 8712 4496 8756
rect 4600 8712 4656 8756
rect 4760 8736 4816 8756
rect 4920 8736 4976 8756
rect 4760 8680 4976 8736
rect 5080 8712 5136 8756
rect 3664 8589 3736 8602
rect 3664 8543 3677 8589
rect 3723 8543 3736 8589
rect 4120 8586 4176 8680
rect 4760 8586 4816 8680
rect 5368 8602 5424 8756
rect 5360 8589 5432 8602
rect 3664 8530 3736 8543
rect 3952 8573 4024 8586
rect 986 8363 1098 8408
rect 986 8317 1019 8363
rect 1065 8317 1098 8363
rect 986 8272 1098 8317
rect 1202 8272 1314 8408
rect 1418 8272 1530 8408
rect 1634 8272 1746 8408
rect 1850 8272 1962 8408
rect 2066 8272 2178 8408
rect 2282 8272 2394 8408
rect 2498 8272 2610 8408
rect 2714 8272 2826 8408
rect 2930 8363 3042 8408
rect 2930 8317 2963 8363
rect 3009 8317 3042 8363
rect 2930 8272 3042 8317
rect 3672 8376 3728 8530
rect 3952 8527 3965 8573
rect 4011 8527 4024 8573
rect 3952 8514 4024 8527
rect 4112 8573 4184 8586
rect 4112 8527 4125 8573
rect 4171 8527 4184 8573
rect 4112 8514 4184 8527
rect 4432 8573 4504 8586
rect 4432 8527 4445 8573
rect 4491 8527 4504 8573
rect 3960 8376 4016 8514
rect 4432 8512 4504 8527
rect 4752 8573 4824 8586
rect 4752 8527 4765 8573
rect 4811 8527 4824 8573
rect 4752 8514 4824 8527
rect 5072 8573 5144 8586
rect 5072 8527 5085 8573
rect 5131 8527 5144 8573
rect 5360 8543 5373 8589
rect 5419 8543 5432 8589
rect 5360 8530 5432 8543
rect 5072 8514 5144 8527
rect 4440 8452 4496 8512
rect 4120 8376 4176 8420
rect 4280 8376 4336 8420
rect 4440 8396 4656 8452
rect 4440 8376 4496 8396
rect 4600 8376 4656 8396
rect 4760 8376 4816 8420
rect 4920 8376 4976 8420
rect 5080 8376 5136 8514
rect 5368 8376 5424 8530
rect 986 7602 1098 7646
rect 1202 7626 1314 7646
rect 1418 7626 1530 7646
rect 1634 7626 1746 7646
rect 1850 7626 1962 7646
rect 2066 7626 2178 7646
rect 2282 7626 2394 7646
rect 2498 7626 2610 7646
rect 2714 7626 2826 7646
rect 1202 7580 2826 7626
rect 2930 7602 3042 7646
rect 1202 7534 1242 7580
rect 1288 7534 1346 7580
rect 1392 7534 2826 7580
rect 1202 7514 2826 7534
rect 3672 7582 3728 7626
rect 3960 7582 4016 7626
rect 4120 7606 4176 7626
rect 4280 7606 4336 7626
rect -7386 7108 -7186 7121
rect -7386 7062 -7373 7108
rect -7199 7062 -7186 7108
rect -7386 7019 -7186 7062
rect -7386 6516 -7186 6559
rect -7386 6470 -7373 6516
rect -7199 6470 -7186 6516
rect -7386 6457 -7186 6470
rect -7106 7108 -6906 7121
rect -7106 7062 -7093 7108
rect -6919 7062 -6906 7108
rect -7106 7019 -6906 7062
rect -7106 6516 -6906 6559
rect -7106 6470 -7093 6516
rect -6919 6470 -6906 6516
rect -7106 6457 -6906 6470
rect -6826 7108 -6626 7121
rect -6826 7062 -6813 7108
rect -6639 7062 -6626 7108
rect -6826 7019 -6626 7062
rect -6826 6516 -6626 6559
rect -6826 6470 -6813 6516
rect -6639 6470 -6626 6516
rect -6826 6457 -6626 6470
rect -6546 7108 -6346 7121
rect -6546 7062 -6533 7108
rect -6359 7062 -6346 7108
rect -6546 7019 -6346 7062
rect -6546 6516 -6346 6559
rect -6546 6470 -6533 6516
rect -6359 6470 -6346 6516
rect -6546 6457 -6346 6470
rect -6266 7108 -6066 7121
rect -6266 7062 -6253 7108
rect -6079 7062 -6066 7108
rect -6266 7019 -6066 7062
rect -6266 6516 -6066 6559
rect -6266 6470 -6253 6516
rect -6079 6470 -6066 6516
rect -6266 6457 -6066 6470
rect -5986 7108 -5786 7121
rect -5986 7062 -5973 7108
rect -5799 7062 -5786 7108
rect -5986 7019 -5786 7062
rect -5986 6516 -5786 6559
rect -5986 6470 -5973 6516
rect -5799 6470 -5786 6516
rect -5986 6457 -5786 6470
rect -5706 7108 -5506 7121
rect -5706 7062 -5693 7108
rect -5519 7062 -5506 7108
rect -5706 7019 -5506 7062
rect -5706 6516 -5506 6559
rect -5706 6470 -5693 6516
rect -5519 6470 -5506 6516
rect -5706 6457 -5506 6470
rect -5426 7108 -5226 7121
rect -5426 7062 -5413 7108
rect -5239 7062 -5226 7108
rect -5426 7019 -5226 7062
rect -5426 6516 -5226 6559
rect -5426 6470 -5413 6516
rect -5239 6470 -5226 6516
rect -5426 6457 -5226 6470
rect -5146 7108 -4946 7121
rect -5146 7062 -5133 7108
rect -4959 7062 -4946 7108
rect -5146 7019 -4946 7062
rect -5146 6516 -4946 6559
rect -5146 6470 -5133 6516
rect -4959 6470 -4946 6516
rect -5146 6457 -4946 6470
rect -4866 7108 -4666 7121
rect -4866 7062 -4853 7108
rect -4679 7062 -4666 7108
rect -4866 7019 -4666 7062
rect -4866 6516 -4666 6559
rect -4866 6470 -4853 6516
rect -4679 6470 -4666 6516
rect -4866 6457 -4666 6470
rect -4586 7108 -4386 7121
rect -4586 7062 -4573 7108
rect -4399 7062 -4386 7108
rect -4586 7019 -4386 7062
rect -4586 6516 -4386 6559
rect -4586 6470 -4573 6516
rect -4399 6470 -4386 6516
rect -4586 6457 -4386 6470
rect -4306 7108 -4106 7121
rect -4306 7062 -4293 7108
rect -4119 7062 -4106 7108
rect -4306 7019 -4106 7062
rect -4306 6516 -4106 6559
rect -4306 6470 -4293 6516
rect -4119 6470 -4106 6516
rect -4306 6457 -4106 6470
rect -7386 6191 -7186 6204
rect -7386 6145 -7373 6191
rect -7199 6145 -7186 6191
rect -7386 6102 -7186 6145
rect -7386 5599 -7186 5642
rect -7386 5553 -7373 5599
rect -7199 5553 -7186 5599
rect -7386 5540 -7186 5553
rect -7106 6191 -6906 6204
rect -7106 6145 -7093 6191
rect -6919 6145 -6906 6191
rect -7106 6102 -6906 6145
rect -7106 5599 -6906 5642
rect -7106 5553 -7093 5599
rect -6919 5553 -6906 5599
rect -7106 5540 -6906 5553
rect -6826 6191 -6626 6204
rect -6826 6145 -6813 6191
rect -6639 6145 -6626 6191
rect -6826 6102 -6626 6145
rect -6826 5599 -6626 5642
rect -6826 5553 -6813 5599
rect -6639 5553 -6626 5599
rect -6826 5540 -6626 5553
rect -6546 6191 -6346 6204
rect -6546 6145 -6533 6191
rect -6359 6145 -6346 6191
rect -6546 6102 -6346 6145
rect -6546 5599 -6346 5642
rect -6546 5553 -6533 5599
rect -6359 5553 -6346 5599
rect -6546 5540 -6346 5553
rect -6266 6191 -6066 6204
rect -6266 6145 -6253 6191
rect -6079 6145 -6066 6191
rect -6266 6102 -6066 6145
rect -6266 5599 -6066 5642
rect -6266 5553 -6253 5599
rect -6079 5553 -6066 5599
rect -6266 5540 -6066 5553
rect -5986 6191 -5786 6204
rect -5986 6145 -5973 6191
rect -5799 6145 -5786 6191
rect -5986 6102 -5786 6145
rect -5986 5599 -5786 5642
rect -5986 5553 -5973 5599
rect -5799 5553 -5786 5599
rect -5986 5540 -5786 5553
rect -5706 6191 -5506 6204
rect -5706 6145 -5693 6191
rect -5519 6145 -5506 6191
rect -5706 6102 -5506 6145
rect -5706 5599 -5506 5642
rect -5706 5553 -5693 5599
rect -5519 5553 -5506 5599
rect -5706 5540 -5506 5553
rect -5426 6191 -5226 6204
rect -5426 6145 -5413 6191
rect -5239 6145 -5226 6191
rect -5426 6102 -5226 6145
rect -5426 5599 -5226 5642
rect -5426 5553 -5413 5599
rect -5239 5553 -5226 5599
rect -5426 5540 -5226 5553
rect -5146 6191 -4946 6204
rect -5146 6145 -5133 6191
rect -4959 6145 -4946 6191
rect -5146 6102 -4946 6145
rect -5146 5599 -4946 5642
rect -5146 5553 -5133 5599
rect -4959 5553 -4946 5599
rect -5146 5540 -4946 5553
rect -4866 6191 -4666 6204
rect -4866 6145 -4853 6191
rect -4679 6145 -4666 6191
rect -4866 6102 -4666 6145
rect -4866 5599 -4666 5642
rect -4866 5553 -4853 5599
rect -4679 5553 -4666 5599
rect -4866 5540 -4666 5553
rect -4586 6191 -4386 6204
rect -4586 6145 -4573 6191
rect -4399 6145 -4386 6191
rect -4586 6102 -4386 6145
rect -4586 5599 -4386 5642
rect -4586 5553 -4573 5599
rect -4399 5553 -4386 5599
rect -4586 5540 -4386 5553
rect -4306 6191 -4106 6204
rect -4306 6145 -4293 6191
rect -4119 6145 -4106 6191
rect -4306 6102 -4106 6145
rect -4306 5599 -4106 5642
rect -4306 5553 -4293 5599
rect -4119 5553 -4106 5599
rect -4306 5540 -4106 5553
rect -7386 5274 -7186 5287
rect -7386 5228 -7373 5274
rect -7199 5228 -7186 5274
rect -7386 5185 -7186 5228
rect -7386 4682 -7186 4725
rect -7386 4636 -7373 4682
rect -7199 4636 -7186 4682
rect -7386 4623 -7186 4636
rect -7106 5274 -6906 5287
rect -7106 5228 -7093 5274
rect -6919 5228 -6906 5274
rect -7106 5185 -6906 5228
rect -7106 4682 -6906 4725
rect -7106 4636 -7093 4682
rect -6919 4636 -6906 4682
rect -7106 4623 -6906 4636
rect -6826 5274 -6626 5287
rect -6826 5228 -6813 5274
rect -6639 5228 -6626 5274
rect -6826 5185 -6626 5228
rect -6826 4682 -6626 4725
rect -6826 4636 -6813 4682
rect -6639 4636 -6626 4682
rect -6826 4623 -6626 4636
rect -6546 5274 -6346 5287
rect -6546 5228 -6533 5274
rect -6359 5228 -6346 5274
rect -6546 5185 -6346 5228
rect -6546 4682 -6346 4725
rect -6546 4636 -6533 4682
rect -6359 4636 -6346 4682
rect -6546 4623 -6346 4636
rect -6266 5274 -6066 5287
rect -6266 5228 -6253 5274
rect -6079 5228 -6066 5274
rect -6266 5185 -6066 5228
rect -6266 4682 -6066 4725
rect -6266 4636 -6253 4682
rect -6079 4636 -6066 4682
rect -6266 4623 -6066 4636
rect -5986 5274 -5786 5287
rect -5986 5228 -5973 5274
rect -5799 5228 -5786 5274
rect -5986 5185 -5786 5228
rect -5986 4682 -5786 4725
rect -5986 4636 -5973 4682
rect -5799 4636 -5786 4682
rect -5986 4623 -5786 4636
rect -5706 5274 -5506 5287
rect -5706 5228 -5693 5274
rect -5519 5228 -5506 5274
rect -5706 5185 -5506 5228
rect -5706 4682 -5506 4725
rect -5706 4636 -5693 4682
rect -5519 4636 -5506 4682
rect -5706 4623 -5506 4636
rect -5426 5274 -5226 5287
rect -5426 5228 -5413 5274
rect -5239 5228 -5226 5274
rect -5426 5185 -5226 5228
rect -5426 4682 -5226 4725
rect -5426 4636 -5413 4682
rect -5239 4636 -5226 4682
rect -5426 4623 -5226 4636
rect -5146 5274 -4946 5287
rect -5146 5228 -5133 5274
rect -4959 5228 -4946 5274
rect -5146 5185 -4946 5228
rect -5146 4682 -4946 4725
rect -5146 4636 -5133 4682
rect -4959 4636 -4946 4682
rect -5146 4623 -4946 4636
rect -4866 5274 -4666 5287
rect -4866 5228 -4853 5274
rect -4679 5228 -4666 5274
rect -4866 5185 -4666 5228
rect -4866 4682 -4666 4725
rect -4866 4636 -4853 4682
rect -4679 4636 -4666 4682
rect -4866 4623 -4666 4636
rect -4586 5274 -4386 5287
rect -4586 5228 -4573 5274
rect -4399 5228 -4386 5274
rect -4586 5185 -4386 5228
rect -4586 4682 -4386 4725
rect -4586 4636 -4573 4682
rect -4399 4636 -4386 4682
rect -4586 4623 -4386 4636
rect -4306 5274 -4106 5287
rect -4306 5228 -4293 5274
rect -4119 5228 -4106 5274
rect -4306 5185 -4106 5228
rect -4306 4682 -4106 4725
rect -4306 4636 -4293 4682
rect -4119 4636 -4106 4682
rect -4306 4623 -4106 4636
rect 4120 7550 4336 7606
rect 4440 7582 4496 7626
rect 4600 7582 4656 7626
rect 4760 7606 4816 7626
rect 4920 7606 4976 7626
rect 4760 7550 4976 7606
rect 5080 7582 5136 7626
rect 5368 7582 5424 7626
rect 4120 7502 4176 7550
rect 4760 7502 4816 7550
rect 4112 7489 4184 7502
rect 4112 7443 4125 7489
rect 4171 7443 4184 7489
rect 4112 7430 4184 7443
rect 4752 7489 4824 7502
rect 4752 7443 4765 7489
rect 4811 7443 4824 7489
rect 4752 7430 4824 7443
rect 6537 14276 6593 14320
rect 6825 14276 6881 14320
rect 6985 14276 7041 14320
rect 7145 14276 7201 14320
rect 7305 14276 7361 14320
rect 7465 14276 7521 14320
rect 7625 14276 7681 14320
rect 7785 14276 7841 14320
rect 7945 14276 8001 14320
rect 8233 14276 8289 14320
rect 6537 13414 6593 13700
rect 6825 13641 6881 13700
rect 6985 13641 7041 13700
rect 7145 13641 7201 13700
rect 7305 13641 7361 13700
rect 7465 13641 7521 13700
rect 7625 13641 7681 13700
rect 7785 13641 7841 13700
rect 7945 13641 8001 13700
rect 6825 13521 8001 13641
rect 6825 13414 6881 13521
rect 6985 13414 7041 13521
rect 7145 13414 7201 13521
rect 7305 13478 8001 13521
rect 7305 13414 7361 13478
rect 7465 13414 7521 13478
rect 7625 13414 7681 13478
rect 7785 13414 7841 13478
rect 7945 13414 8001 13478
rect 8233 13414 8289 13700
rect 6537 12552 6593 12838
rect 6825 12777 6881 12838
rect 6985 12777 7041 12838
rect 7145 12777 7201 12838
rect 7305 12777 7361 12838
rect 7465 12777 7521 12838
rect 7625 12777 7681 12838
rect 7785 12777 7841 12838
rect 7945 12777 8001 12838
rect 6825 12657 8001 12777
rect 6825 12552 6881 12657
rect 6985 12552 7041 12657
rect 7145 12552 7201 12657
rect 7305 12552 7361 12657
rect 7465 12552 7521 12657
rect 7625 12552 7681 12657
rect 7785 12552 7841 12657
rect 7945 12552 8001 12657
rect 8233 12552 8289 12838
rect 6537 11690 6593 11976
rect 6825 11907 6881 11976
rect 6985 11907 7041 11976
rect 7145 11907 7201 11976
rect 7305 11907 7361 11976
rect 7465 11907 7521 11976
rect 7625 11907 7681 11976
rect 7785 11907 7841 11976
rect 7945 11907 8001 11976
rect 6825 11787 8001 11907
rect 6825 11690 6881 11787
rect 6985 11690 7041 11787
rect 7145 11690 7201 11787
rect 7305 11690 7361 11787
rect 7465 11690 7521 11787
rect 7625 11690 7681 11787
rect 7785 11690 7841 11787
rect 7945 11690 8001 11787
rect 8233 11690 8289 11976
rect 19067 13402 19139 13415
rect 19067 13356 19080 13402
rect 19126 13356 19139 13402
rect 19067 13343 19139 13356
rect 19547 13402 19619 13415
rect 19547 13356 19560 13402
rect 19606 13356 19619 13402
rect 19547 13343 19619 13356
rect 20187 13402 20259 13415
rect 20187 13356 20200 13402
rect 20246 13356 20259 13402
rect 20187 13343 20259 13356
rect 18787 13189 18843 13233
rect 19075 13189 19131 13343
rect 19555 13265 19611 13343
rect 19235 13189 19291 13233
rect 19395 13189 19451 13233
rect 19555 13209 19771 13265
rect 19555 13189 19611 13209
rect 19715 13189 19771 13209
rect 19875 13189 19931 13233
rect 20035 13189 20091 13233
rect 20195 13189 20251 13343
rect 20483 13189 20539 13233
rect 18787 12457 18843 12589
rect 19075 12545 19131 12589
rect 19235 12569 19291 12589
rect 19395 12569 19451 12589
rect 19235 12513 19451 12569
rect 19555 12545 19611 12589
rect 19715 12545 19771 12589
rect 19875 12569 19931 12589
rect 20035 12569 20091 12589
rect 19875 12513 20091 12569
rect 20195 12545 20251 12589
rect 18779 12444 18851 12457
rect 19235 12449 19291 12513
rect 19875 12449 19931 12513
rect 20483 12457 20539 12589
rect 18779 12398 18792 12444
rect 18838 12398 18851 12444
rect 18779 12385 18851 12398
rect 19067 12436 19139 12449
rect 19067 12390 19080 12436
rect 19126 12390 19139 12436
rect 18787 12253 18843 12385
rect 19067 12377 19139 12390
rect 19227 12436 19299 12449
rect 19227 12390 19240 12436
rect 19286 12390 19299 12436
rect 19227 12377 19299 12390
rect 19547 12436 19619 12449
rect 19547 12390 19560 12436
rect 19606 12390 19619 12436
rect 19547 12377 19619 12390
rect 19867 12436 19939 12449
rect 19867 12390 19880 12436
rect 19926 12390 19939 12436
rect 19867 12377 19939 12390
rect 20187 12436 20259 12449
rect 20187 12390 20200 12436
rect 20246 12390 20259 12436
rect 20187 12377 20259 12390
rect 20475 12444 20547 12457
rect 20475 12398 20488 12444
rect 20534 12398 20547 12444
rect 20475 12385 20547 12398
rect 19075 12253 19131 12377
rect 19555 12329 19611 12377
rect 19235 12253 19291 12297
rect 19395 12253 19451 12297
rect 19555 12273 19771 12329
rect 19555 12253 19611 12273
rect 19715 12253 19771 12273
rect 19875 12253 19931 12297
rect 20035 12253 20091 12297
rect 20195 12253 20251 12377
rect 20483 12253 20539 12385
rect 12154 11377 12210 11421
rect 12442 11377 12498 11421
rect 12730 11377 12786 11421
rect 12890 11377 12946 11421
rect 13178 11377 13234 11421
rect 13338 11377 13394 11421
rect 13626 11377 13682 11421
rect 13786 11377 13842 11421
rect 14074 11377 14130 11421
rect 14362 11377 14418 11421
rect 6537 10828 6593 11114
rect 6825 11033 6881 11114
rect 6985 11033 7041 11114
rect 7145 11033 7201 11114
rect 7305 11033 7361 11114
rect 7465 11033 7521 11114
rect 7625 11033 7681 11114
rect 7785 11033 7841 11114
rect 7945 11033 8001 11114
rect 6825 10913 8001 11033
rect 6825 10828 6881 10913
rect 6985 10828 7041 10913
rect 7145 10828 7201 10913
rect 7305 10828 7361 10913
rect 7465 10828 7521 10913
rect 7625 10828 7681 10913
rect 7785 10828 7841 10913
rect 7945 10828 8001 10913
rect 8233 10828 8289 11114
rect 8772 10809 8828 10853
rect 9060 10809 9116 10853
rect 9348 10809 9404 10853
rect 9508 10809 9564 10853
rect 9796 10809 9852 10853
rect 9956 10809 10012 10853
rect 10244 10809 10300 10853
rect 10404 10809 10460 10853
rect 10692 10809 10748 10853
rect 10980 10809 11036 10853
rect 6537 9966 6593 10252
rect 6825 10173 6881 10252
rect 6985 10173 7041 10252
rect 7145 10173 7201 10252
rect 7305 10173 7361 10252
rect 7465 10173 7521 10252
rect 7625 10173 7681 10252
rect 7785 10173 7841 10252
rect 7945 10173 8001 10252
rect 6825 10053 8001 10173
rect 6825 9966 6881 10053
rect 6985 9966 7041 10053
rect 7145 9966 7201 10053
rect 7305 9966 7361 10053
rect 7465 9966 7521 10053
rect 7625 9966 7681 10053
rect 7785 9966 7841 10053
rect 7945 9966 8001 10053
rect 8233 9966 8289 10252
rect 8772 9947 8828 10233
rect 9060 10135 9116 10233
rect 9348 10135 9404 10233
rect 9508 10135 9564 10233
rect 9796 10135 9852 10233
rect 9956 10135 10012 10233
rect 10244 10135 10300 10233
rect 10404 10135 10460 10233
rect 10692 10135 10748 10233
rect 9060 10015 10748 10135
rect 9060 9947 9116 10015
rect 9348 9947 9404 10015
rect 9508 9947 9564 10015
rect 9796 9947 9852 10015
rect 9956 9947 10012 10015
rect 10244 9947 10300 10015
rect 10404 9947 10460 10015
rect 10692 9947 10748 10015
rect 10980 9947 11036 10233
rect 6537 9104 6593 9390
rect 6825 9317 6881 9390
rect 6985 9317 7041 9390
rect 7145 9317 7201 9390
rect 7305 9317 7361 9390
rect 7465 9317 7521 9390
rect 7625 9317 7681 9390
rect 7785 9317 7841 9390
rect 7945 9317 8001 9390
rect 6825 9197 8001 9317
rect 6825 9104 6881 9197
rect 6985 9104 7041 9197
rect 7145 9104 7201 9197
rect 7305 9104 7361 9197
rect 7465 9104 7521 9197
rect 7625 9104 7681 9197
rect 7785 9104 7841 9197
rect 7945 9104 8001 9197
rect 8233 9104 8289 9390
rect 8772 9085 8828 9371
rect 9060 9273 9116 9371
rect 9348 9273 9404 9371
rect 9508 9273 9564 9371
rect 9796 9273 9852 9371
rect 9956 9273 10012 9371
rect 10244 9273 10300 9371
rect 10404 9273 10460 9371
rect 10692 9273 10748 9371
rect 9060 9153 10748 9273
rect 9060 9085 9116 9153
rect 9348 9085 9404 9153
rect 9508 9085 9564 9153
rect 9796 9085 9852 9153
rect 9956 9085 10012 9153
rect 10244 9085 10300 9153
rect 10404 9085 10460 9153
rect 10692 9085 10748 9153
rect 10980 9085 11036 9371
rect 6537 8421 6593 8528
rect 6529 8408 6601 8421
rect 6529 8362 6542 8408
rect 6588 8362 6601 8408
rect 6529 8349 6601 8362
rect 6825 8416 6881 8528
rect 6985 8416 7041 8528
rect 7145 8416 7201 8528
rect 7305 8416 7361 8528
rect 7465 8416 7521 8528
rect 7625 8416 7681 8528
rect 7785 8416 7841 8528
rect 7945 8476 8001 8528
rect 7945 8474 8020 8476
rect 7945 8461 8063 8474
rect 7945 8416 8004 8461
rect 6825 8415 8004 8416
rect 8050 8415 8063 8461
rect 8233 8421 8289 8528
rect 6825 8357 8063 8415
rect 6537 8242 6593 8349
rect 6825 8311 8004 8357
rect 8050 8311 8063 8357
rect 8225 8408 8297 8421
rect 8225 8362 8238 8408
rect 8284 8362 8297 8408
rect 8225 8349 8297 8362
rect 8772 8402 8828 8509
rect 9060 8441 9116 8509
rect 9348 8441 9404 8509
rect 9508 8441 9564 8509
rect 9796 8441 9852 8509
rect 9956 8441 10012 8509
rect 10244 8441 10300 8509
rect 10404 8441 10460 8509
rect 10692 8463 10748 8509
rect 10692 8450 10796 8463
rect 10692 8441 10737 8450
rect 9060 8404 10737 8441
rect 10783 8404 10796 8450
rect 6825 8298 8063 8311
rect 6825 8296 8020 8298
rect 6825 8242 6881 8296
rect 6985 8242 7041 8296
rect 7145 8242 7201 8296
rect 7305 8242 7361 8296
rect 7465 8242 7521 8296
rect 7625 8242 7681 8296
rect 7785 8242 7841 8296
rect 7945 8242 8001 8296
rect 8233 8242 8289 8349
rect 8764 8389 8836 8402
rect 8764 8343 8777 8389
rect 8823 8343 8836 8389
rect 8764 8330 8836 8343
rect 9060 8346 10796 8404
rect 10980 8402 11036 8509
rect 8772 8223 8828 8330
rect 9060 8321 10737 8346
rect 9060 8223 9116 8321
rect 9348 8223 9404 8321
rect 9508 8223 9564 8321
rect 9796 8223 9852 8321
rect 9956 8223 10012 8321
rect 10244 8223 10300 8321
rect 10404 8223 10460 8321
rect 10692 8300 10737 8321
rect 10783 8300 10796 8346
rect 10972 8389 11044 8402
rect 10972 8343 10985 8389
rect 11031 8343 11044 8389
rect 10972 8330 11044 8343
rect 10692 8287 10796 8300
rect 10692 8223 10748 8287
rect 10980 8223 11036 8330
rect 6537 7622 6593 7666
rect 6825 7622 6881 7666
rect 6985 7622 7041 7666
rect 7145 7622 7201 7666
rect 7305 7622 7361 7666
rect 7465 7622 7521 7666
rect 7625 7622 7681 7666
rect 7785 7622 7841 7666
rect 7945 7622 8001 7666
rect 8233 7622 8289 7666
rect 8772 7603 8828 7647
rect 9060 7603 9116 7647
rect 9348 7603 9404 7647
rect 9508 7603 9564 7647
rect 9796 7603 9852 7647
rect 9956 7603 10012 7647
rect 10244 7603 10300 7647
rect 10404 7603 10460 7647
rect 10692 7603 10748 7647
rect 10980 7603 11036 7647
rect 14948 11377 15004 11421
rect 15236 11377 15292 11421
rect 15396 11377 15452 11421
rect 15556 11377 15612 11421
rect 15716 11377 15772 11421
rect 15876 11377 15932 11421
rect 16036 11377 16092 11421
rect 16196 11377 16252 11421
rect 16356 11377 16412 11421
rect 16644 11377 16700 11421
rect 12154 10341 12210 10751
rect 12442 10605 12498 10751
rect 12730 10605 12786 10751
rect 12890 10605 12946 10751
rect 13178 10605 13234 10751
rect 13338 10605 13394 10751
rect 13626 10605 13682 10751
rect 13786 10605 13842 10751
rect 14074 10605 14130 10751
rect 12442 10485 14130 10605
rect 12442 10341 12498 10485
rect 12730 10341 12786 10485
rect 12890 10341 12946 10485
rect 13178 10341 13234 10485
rect 13338 10341 13394 10485
rect 13626 10341 13682 10485
rect 13786 10341 13842 10485
rect 14074 10341 14130 10485
rect 14362 10341 14418 10751
rect 14948 10341 15004 10751
rect 15236 10590 15292 10751
rect 15396 10590 15452 10751
rect 15556 10590 15612 10751
rect 15716 10590 15772 10751
rect 15876 10590 15932 10751
rect 16036 10590 16092 10751
rect 16196 10590 16252 10751
rect 16356 10590 16412 10751
rect 15236 10470 16412 10590
rect 15236 10341 15292 10470
rect 15396 10341 15452 10470
rect 15556 10341 15612 10470
rect 15716 10341 15772 10470
rect 15876 10341 15932 10470
rect 16036 10341 16092 10470
rect 16196 10341 16252 10470
rect 16356 10341 16412 10470
rect 16644 10341 16700 10751
rect 12154 9305 12210 9715
rect 12442 9555 12498 9715
rect 12730 9555 12786 9715
rect 12890 9555 12946 9715
rect 13178 9555 13234 9715
rect 13338 9555 13394 9715
rect 13626 9555 13682 9715
rect 13786 9555 13842 9715
rect 14074 9555 14130 9715
rect 12442 9435 14130 9555
rect 12442 9305 12498 9435
rect 12730 9305 12786 9435
rect 12890 9305 12946 9435
rect 13178 9305 13234 9435
rect 13338 9305 13394 9435
rect 13626 9305 13682 9435
rect 13786 9305 13842 9435
rect 14074 9305 14130 9435
rect 14362 9305 14418 9715
rect 14948 9305 15004 9715
rect 15236 9563 15292 9715
rect 15396 9563 15452 9715
rect 15556 9563 15612 9715
rect 15716 9563 15772 9715
rect 15876 9563 15932 9715
rect 16036 9563 16092 9715
rect 16196 9563 16252 9715
rect 16356 9563 16412 9715
rect 15236 9443 16412 9563
rect 15236 9305 15292 9443
rect 15396 9305 15452 9443
rect 15556 9305 15612 9443
rect 15716 9305 15772 9443
rect 15876 9305 15932 9443
rect 16036 9305 16092 9443
rect 16196 9305 16252 9443
rect 16356 9305 16412 9443
rect 16644 9305 16700 9715
rect 12154 8448 12210 8679
rect 12442 8575 12498 8679
rect 12388 8560 12498 8575
rect 12388 8514 12403 8560
rect 12449 8515 12498 8560
rect 12730 8515 12786 8679
rect 12890 8515 12946 8679
rect 13178 8515 13234 8679
rect 13338 8515 13394 8679
rect 13626 8515 13682 8679
rect 13786 8515 13842 8679
rect 14074 8515 14130 8679
rect 12449 8514 14130 8515
rect 12388 8456 14130 8514
rect 12146 8435 12218 8448
rect 12146 8389 12159 8435
rect 12205 8389 12218 8435
rect 12388 8410 12403 8456
rect 12449 8410 14130 8456
rect 14362 8448 14418 8679
rect 12388 8395 14130 8410
rect 12146 8376 12218 8389
rect 12154 8269 12210 8376
rect 12442 8269 12498 8395
rect 12730 8269 12786 8395
rect 12890 8269 12946 8395
rect 13178 8269 13234 8395
rect 13338 8269 13394 8395
rect 13626 8269 13682 8395
rect 13786 8269 13842 8395
rect 14074 8269 14130 8395
rect 14354 8435 14426 8448
rect 14354 8389 14367 8435
rect 14413 8389 14426 8435
rect 14354 8376 14426 8389
rect 14948 8448 15004 8679
rect 15236 8580 15292 8679
rect 15174 8565 15292 8580
rect 15174 8519 15189 8565
rect 15235 8520 15292 8565
rect 15396 8520 15452 8679
rect 15556 8520 15612 8679
rect 15716 8520 15772 8679
rect 15876 8520 15932 8679
rect 16036 8520 16092 8679
rect 16196 8520 16252 8679
rect 16356 8520 16412 8679
rect 15235 8519 16412 8520
rect 15174 8461 16412 8519
rect 14362 8269 14418 8376
rect 14940 8435 15012 8448
rect 14940 8389 14953 8435
rect 14999 8389 15012 8435
rect 15174 8415 15189 8461
rect 15235 8415 16412 8461
rect 16644 8448 16700 8679
rect 15174 8400 16412 8415
rect 14940 8376 15012 8389
rect 14948 8269 15004 8376
rect 15236 8269 15292 8400
rect 15396 8269 15452 8400
rect 15556 8269 15612 8400
rect 15716 8269 15772 8400
rect 15876 8269 15932 8400
rect 16036 8269 16092 8400
rect 16196 8269 16252 8400
rect 16356 8269 16412 8400
rect 16636 8435 16708 8448
rect 16636 8389 16649 8435
rect 16695 8389 16708 8435
rect 16636 8376 16708 8389
rect 16644 8269 16700 8376
rect 12154 7599 12210 7643
rect 12442 7599 12498 7643
rect 12730 7599 12786 7643
rect 12890 7599 12946 7643
rect 13178 7599 13234 7643
rect 13338 7599 13394 7643
rect 13626 7599 13682 7643
rect 13786 7599 13842 7643
rect 14074 7599 14130 7643
rect 14362 7599 14418 7643
rect 14948 7599 15004 7643
rect 15236 7599 15292 7643
rect 15396 7599 15452 7643
rect 15556 7599 15612 7643
rect 15716 7599 15772 7643
rect 15876 7599 15932 7643
rect 16036 7599 16092 7643
rect 16196 7599 16252 7643
rect 16356 7599 16412 7643
rect 16644 7599 16700 7643
rect 18787 11317 18843 11653
rect 19075 11609 19131 11653
rect 19235 11633 19291 11653
rect 19395 11633 19451 11653
rect 19235 11577 19451 11633
rect 19555 11609 19611 11653
rect 19715 11609 19771 11653
rect 19875 11633 19931 11653
rect 20035 11633 20091 11653
rect 19875 11577 20091 11633
rect 20195 11609 20251 11653
rect 19235 11513 19291 11577
rect 19875 11513 19931 11577
rect 19067 11500 19139 11513
rect 19067 11454 19080 11500
rect 19126 11454 19139 11500
rect 19067 11441 19139 11454
rect 19227 11500 19299 11513
rect 19227 11454 19240 11500
rect 19286 11454 19299 11500
rect 19227 11441 19299 11454
rect 19547 11500 19619 11513
rect 19547 11454 19560 11500
rect 19606 11454 19619 11500
rect 19547 11441 19619 11454
rect 19867 11500 19939 11513
rect 19867 11454 19880 11500
rect 19926 11454 19939 11500
rect 19867 11441 19939 11454
rect 20187 11500 20259 11513
rect 20187 11454 20200 11500
rect 20246 11454 20259 11500
rect 20187 11441 20259 11454
rect 19075 11317 19131 11441
rect 19555 11393 19611 11441
rect 19235 11317 19291 11361
rect 19395 11317 19451 11361
rect 19555 11337 19771 11393
rect 19555 11317 19611 11337
rect 19715 11317 19771 11337
rect 19875 11317 19931 11361
rect 20035 11317 20091 11361
rect 20195 11317 20251 11441
rect 20483 11317 20539 11653
rect 18787 10381 18843 10717
rect 19075 10381 19131 10717
rect 19235 10381 19291 10717
rect 19395 10381 19451 10717
rect 19555 10381 19611 10717
rect 19715 10381 19771 10717
rect 19875 10381 19931 10717
rect 20035 10381 20091 10717
rect 20195 10381 20251 10717
rect 20483 10381 20539 10717
rect 18787 9445 18843 9781
rect 19075 9737 19131 9781
rect 19235 9761 19291 9781
rect 19395 9761 19451 9781
rect 19235 9705 19451 9761
rect 19555 9737 19611 9781
rect 19715 9737 19771 9781
rect 19875 9761 19931 9781
rect 20035 9761 20091 9781
rect 19875 9705 20091 9761
rect 20195 9737 20251 9781
rect 19235 9641 19291 9705
rect 19875 9641 19931 9705
rect 19067 9628 19139 9641
rect 19067 9582 19080 9628
rect 19126 9582 19139 9628
rect 19067 9569 19139 9582
rect 19227 9628 19299 9641
rect 19227 9582 19240 9628
rect 19286 9582 19299 9628
rect 19227 9569 19299 9582
rect 19547 9628 19619 9641
rect 19547 9582 19560 9628
rect 19606 9582 19619 9628
rect 19547 9569 19619 9582
rect 19867 9628 19939 9641
rect 19867 9582 19880 9628
rect 19926 9582 19939 9628
rect 19867 9569 19939 9582
rect 20187 9628 20259 9641
rect 20187 9582 20200 9628
rect 20246 9582 20259 9628
rect 20187 9569 20259 9582
rect 19075 9445 19131 9569
rect 19555 9521 19611 9569
rect 19235 9445 19291 9489
rect 19395 9445 19451 9489
rect 19555 9465 19771 9521
rect 19555 9445 19611 9465
rect 19715 9445 19771 9465
rect 19875 9445 19931 9489
rect 20035 9445 20091 9489
rect 20195 9445 20251 9569
rect 20483 9445 20539 9781
rect 18787 8713 18843 8845
rect 19075 8801 19131 8845
rect 19235 8825 19291 8845
rect 19395 8825 19451 8845
rect 19235 8769 19451 8825
rect 19555 8801 19611 8845
rect 19715 8801 19771 8845
rect 19875 8825 19931 8845
rect 20035 8825 20091 8845
rect 19875 8769 20091 8825
rect 20195 8801 20251 8845
rect 18779 8700 18851 8713
rect 19235 8705 19291 8769
rect 19875 8705 19931 8769
rect 20483 8713 20539 8845
rect 18779 8654 18792 8700
rect 18838 8654 18851 8700
rect 18779 8641 18851 8654
rect 19067 8692 19139 8705
rect 19067 8646 19080 8692
rect 19126 8646 19139 8692
rect 18787 8509 18843 8641
rect 19067 8633 19139 8646
rect 19227 8692 19299 8705
rect 19227 8646 19240 8692
rect 19286 8646 19299 8692
rect 19227 8633 19299 8646
rect 19547 8692 19619 8705
rect 19547 8646 19560 8692
rect 19606 8646 19619 8692
rect 19547 8633 19619 8646
rect 19867 8692 19939 8705
rect 19867 8646 19880 8692
rect 19926 8646 19939 8692
rect 19867 8633 19939 8646
rect 20187 8692 20259 8705
rect 20187 8646 20200 8692
rect 20246 8646 20259 8692
rect 20187 8633 20259 8646
rect 20475 8700 20547 8713
rect 20475 8654 20488 8700
rect 20534 8654 20547 8700
rect 20475 8641 20547 8654
rect 19075 8509 19131 8633
rect 19555 8585 19611 8633
rect 19235 8509 19291 8553
rect 19395 8509 19451 8553
rect 19555 8529 19771 8585
rect 19555 8509 19611 8529
rect 19715 8509 19771 8529
rect 19875 8509 19931 8553
rect 20035 8509 20091 8553
rect 20195 8509 20251 8633
rect 20483 8509 20539 8641
rect 18787 7865 18843 7909
rect 19075 7865 19131 7909
rect 19235 7889 19291 7909
rect 19395 7889 19451 7909
rect 19235 7833 19451 7889
rect 19555 7865 19611 7909
rect 19715 7865 19771 7909
rect 19875 7889 19931 7909
rect 20035 7889 20091 7909
rect 19875 7833 20091 7889
rect 20195 7865 20251 7909
rect 20483 7865 20539 7909
rect 19235 7769 19291 7833
rect 19875 7769 19931 7833
rect 19227 7756 19299 7769
rect 19227 7710 19240 7756
rect 19286 7710 19299 7756
rect 19227 7697 19299 7710
rect 19867 7756 19939 7769
rect 19867 7710 19880 7756
rect 19926 7710 19939 7756
rect 19867 7697 19939 7710
rect 24219 13402 24291 13415
rect 24219 13356 24232 13402
rect 24278 13356 24291 13402
rect 24219 13343 24291 13356
rect 24859 13402 24931 13415
rect 24859 13356 24872 13402
rect 24918 13356 24931 13402
rect 24859 13343 24931 13356
rect 25339 13402 25411 13415
rect 25339 13356 25352 13402
rect 25398 13356 25411 13402
rect 25339 13343 25411 13356
rect 23939 13189 23995 13233
rect 24227 13189 24283 13343
rect 24867 13265 24923 13343
rect 24387 13189 24443 13233
rect 24547 13189 24603 13233
rect 24707 13209 24923 13265
rect 24707 13189 24763 13209
rect 24867 13189 24923 13209
rect 25027 13189 25083 13233
rect 25187 13189 25243 13233
rect 25347 13189 25403 13343
rect 25635 13189 25691 13233
rect 23939 12457 23995 12589
rect 24227 12545 24283 12589
rect 24387 12569 24443 12589
rect 24547 12569 24603 12589
rect 24387 12513 24603 12569
rect 24707 12545 24763 12589
rect 24867 12545 24923 12589
rect 25027 12569 25083 12589
rect 25187 12569 25243 12589
rect 25027 12513 25243 12569
rect 25347 12545 25403 12589
rect 23931 12444 24003 12457
rect 24547 12449 24603 12513
rect 25187 12449 25243 12513
rect 25635 12457 25691 12589
rect 23931 12398 23944 12444
rect 23990 12398 24003 12444
rect 23931 12385 24003 12398
rect 24219 12436 24291 12449
rect 24219 12390 24232 12436
rect 24278 12390 24291 12436
rect 23939 12253 23995 12385
rect 24219 12377 24291 12390
rect 24539 12436 24611 12449
rect 24539 12390 24552 12436
rect 24598 12390 24611 12436
rect 24539 12377 24611 12390
rect 24859 12436 24931 12449
rect 24859 12390 24872 12436
rect 24918 12390 24931 12436
rect 24859 12377 24931 12390
rect 25179 12436 25251 12449
rect 25179 12390 25192 12436
rect 25238 12390 25251 12436
rect 25179 12377 25251 12390
rect 25339 12436 25411 12449
rect 25339 12390 25352 12436
rect 25398 12390 25411 12436
rect 25339 12377 25411 12390
rect 25627 12444 25699 12457
rect 25627 12398 25640 12444
rect 25686 12398 25699 12444
rect 25627 12385 25699 12398
rect 24227 12253 24283 12377
rect 24867 12329 24923 12377
rect 24387 12253 24443 12297
rect 24547 12253 24603 12297
rect 24707 12273 24923 12329
rect 24707 12253 24763 12273
rect 24867 12253 24923 12273
rect 25027 12253 25083 12297
rect 25187 12253 25243 12297
rect 25347 12253 25403 12377
rect 25635 12253 25691 12385
rect 23939 11317 23995 11653
rect 24227 11609 24283 11653
rect 24387 11633 24443 11653
rect 24547 11633 24603 11653
rect 24387 11577 24603 11633
rect 24707 11609 24763 11653
rect 24867 11609 24923 11653
rect 25027 11633 25083 11653
rect 25187 11633 25243 11653
rect 25027 11577 25243 11633
rect 25347 11609 25403 11653
rect 24547 11513 24603 11577
rect 25187 11513 25243 11577
rect 24219 11500 24291 11513
rect 24219 11454 24232 11500
rect 24278 11454 24291 11500
rect 24219 11441 24291 11454
rect 24539 11500 24611 11513
rect 24539 11454 24552 11500
rect 24598 11454 24611 11500
rect 24539 11441 24611 11454
rect 24859 11500 24931 11513
rect 24859 11454 24872 11500
rect 24918 11454 24931 11500
rect 24859 11441 24931 11454
rect 25179 11500 25251 11513
rect 25179 11454 25192 11500
rect 25238 11454 25251 11500
rect 25179 11441 25251 11454
rect 25339 11500 25411 11513
rect 25339 11454 25352 11500
rect 25398 11454 25411 11500
rect 25339 11441 25411 11454
rect 24227 11317 24283 11441
rect 24867 11393 24923 11441
rect 24387 11317 24443 11361
rect 24547 11317 24603 11361
rect 24707 11337 24923 11393
rect 24707 11317 24763 11337
rect 24867 11317 24923 11337
rect 25027 11317 25083 11361
rect 25187 11317 25243 11361
rect 25347 11317 25403 11441
rect 25635 11317 25691 11653
rect 23939 10381 23995 10717
rect 24227 10381 24283 10717
rect 24387 10381 24443 10717
rect 24547 10381 24603 10717
rect 24707 10381 24763 10717
rect 24867 10381 24923 10717
rect 25027 10381 25083 10717
rect 25187 10381 25243 10717
rect 25347 10381 25403 10717
rect 25635 10381 25691 10717
rect 23939 9445 23995 9781
rect 24227 9737 24283 9781
rect 24387 9761 24443 9781
rect 24547 9761 24603 9781
rect 24387 9705 24603 9761
rect 24707 9737 24763 9781
rect 24867 9737 24923 9781
rect 25027 9761 25083 9781
rect 25187 9761 25243 9781
rect 25027 9705 25243 9761
rect 25347 9737 25403 9781
rect 24547 9641 24603 9705
rect 25187 9641 25243 9705
rect 24219 9628 24291 9641
rect 24219 9582 24232 9628
rect 24278 9582 24291 9628
rect 24219 9569 24291 9582
rect 24539 9628 24611 9641
rect 24539 9582 24552 9628
rect 24598 9582 24611 9628
rect 24539 9569 24611 9582
rect 24859 9628 24931 9641
rect 24859 9582 24872 9628
rect 24918 9582 24931 9628
rect 24859 9569 24931 9582
rect 25179 9628 25251 9641
rect 25179 9582 25192 9628
rect 25238 9582 25251 9628
rect 25179 9569 25251 9582
rect 25339 9628 25411 9641
rect 25339 9582 25352 9628
rect 25398 9582 25411 9628
rect 25339 9569 25411 9582
rect 24227 9445 24283 9569
rect 24867 9521 24923 9569
rect 24387 9445 24443 9489
rect 24547 9445 24603 9489
rect 24707 9465 24923 9521
rect 24707 9445 24763 9465
rect 24867 9445 24923 9465
rect 25027 9445 25083 9489
rect 25187 9445 25243 9489
rect 25347 9445 25403 9569
rect 25635 9445 25691 9781
rect 23939 8713 23995 8845
rect 24227 8801 24283 8845
rect 24387 8825 24443 8845
rect 24547 8825 24603 8845
rect 24387 8769 24603 8825
rect 24707 8801 24763 8845
rect 24867 8801 24923 8845
rect 25027 8825 25083 8845
rect 25187 8825 25243 8845
rect 25027 8769 25243 8825
rect 25347 8801 25403 8845
rect 23931 8700 24003 8713
rect 24547 8705 24603 8769
rect 25187 8705 25243 8769
rect 25635 8713 25691 8845
rect 23931 8654 23944 8700
rect 23990 8654 24003 8700
rect 23931 8641 24003 8654
rect 24219 8692 24291 8705
rect 24219 8646 24232 8692
rect 24278 8646 24291 8692
rect 23939 8509 23995 8641
rect 24219 8633 24291 8646
rect 24539 8692 24611 8705
rect 24539 8646 24552 8692
rect 24598 8646 24611 8692
rect 24539 8633 24611 8646
rect 24859 8692 24931 8705
rect 24859 8646 24872 8692
rect 24918 8646 24931 8692
rect 24859 8633 24931 8646
rect 25179 8692 25251 8705
rect 25179 8646 25192 8692
rect 25238 8646 25251 8692
rect 25179 8633 25251 8646
rect 25339 8692 25411 8705
rect 25339 8646 25352 8692
rect 25398 8646 25411 8692
rect 25339 8633 25411 8646
rect 25627 8700 25699 8713
rect 25627 8654 25640 8700
rect 25686 8654 25699 8700
rect 25627 8641 25699 8654
rect 24227 8509 24283 8633
rect 24867 8585 24923 8633
rect 24387 8509 24443 8553
rect 24547 8509 24603 8553
rect 24707 8529 24923 8585
rect 24707 8509 24763 8529
rect 24867 8509 24923 8529
rect 25027 8509 25083 8553
rect 25187 8509 25243 8553
rect 25347 8509 25403 8633
rect 25635 8509 25691 8641
rect 23939 7865 23995 7909
rect 24227 7865 24283 7909
rect 24387 7889 24443 7909
rect 24547 7889 24603 7909
rect 24387 7833 24603 7889
rect 24707 7865 24763 7909
rect 24867 7865 24923 7909
rect 25027 7889 25083 7909
rect 25187 7889 25243 7909
rect 25027 7833 25243 7889
rect 25347 7865 25403 7909
rect 25635 7865 25691 7909
rect 24547 7769 24603 7833
rect 25187 7769 25243 7833
rect 24539 7756 24611 7769
rect 24539 7710 24552 7756
rect 24598 7710 24611 7756
rect 24539 7697 24611 7710
rect 25179 7756 25251 7769
rect 25179 7710 25192 7756
rect 25238 7710 25251 7756
rect 25179 7697 25251 7710
rect 28188 13402 28260 13415
rect 28188 13356 28201 13402
rect 28247 13356 28260 13402
rect 28188 13343 28260 13356
rect 28668 13402 28740 13415
rect 28668 13356 28681 13402
rect 28727 13356 28740 13402
rect 28668 13343 28740 13356
rect 29308 13402 29380 13415
rect 29308 13356 29321 13402
rect 29367 13356 29380 13402
rect 29308 13343 29380 13356
rect 27908 13189 27964 13233
rect 28196 13189 28252 13343
rect 28676 13265 28732 13343
rect 28356 13189 28412 13233
rect 28516 13189 28572 13233
rect 28676 13209 28892 13265
rect 28676 13189 28732 13209
rect 28836 13189 28892 13209
rect 28996 13189 29052 13233
rect 29156 13189 29212 13233
rect 29316 13189 29372 13343
rect 29604 13189 29660 13233
rect 27908 12457 27964 12589
rect 28196 12545 28252 12589
rect 28356 12569 28412 12589
rect 28516 12569 28572 12589
rect 28356 12513 28572 12569
rect 28676 12545 28732 12589
rect 28836 12545 28892 12589
rect 28996 12569 29052 12589
rect 29156 12569 29212 12589
rect 28996 12513 29212 12569
rect 29316 12545 29372 12589
rect 27900 12444 27972 12457
rect 28356 12449 28412 12513
rect 28996 12449 29052 12513
rect 29604 12457 29660 12589
rect 27900 12398 27913 12444
rect 27959 12398 27972 12444
rect 27900 12385 27972 12398
rect 28188 12436 28260 12449
rect 28188 12390 28201 12436
rect 28247 12390 28260 12436
rect 27908 12253 27964 12385
rect 28188 12377 28260 12390
rect 28348 12436 28420 12449
rect 28348 12390 28361 12436
rect 28407 12390 28420 12436
rect 28348 12377 28420 12390
rect 28668 12436 28740 12449
rect 28668 12390 28681 12436
rect 28727 12390 28740 12436
rect 28668 12377 28740 12390
rect 28988 12436 29060 12449
rect 28988 12390 29001 12436
rect 29047 12390 29060 12436
rect 28988 12377 29060 12390
rect 29308 12436 29380 12449
rect 29308 12390 29321 12436
rect 29367 12390 29380 12436
rect 29308 12377 29380 12390
rect 29596 12444 29668 12457
rect 29596 12398 29609 12444
rect 29655 12398 29668 12444
rect 29596 12385 29668 12398
rect 28196 12253 28252 12377
rect 28676 12329 28732 12377
rect 28356 12253 28412 12297
rect 28516 12253 28572 12297
rect 28676 12273 28892 12329
rect 28676 12253 28732 12273
rect 28836 12253 28892 12273
rect 28996 12253 29052 12297
rect 29156 12253 29212 12297
rect 29316 12253 29372 12377
rect 29604 12253 29660 12385
rect 27908 11317 27964 11653
rect 28196 11609 28252 11653
rect 28356 11633 28412 11653
rect 28516 11633 28572 11653
rect 28356 11577 28572 11633
rect 28676 11609 28732 11653
rect 28836 11609 28892 11653
rect 28996 11633 29052 11653
rect 29156 11633 29212 11653
rect 28996 11577 29212 11633
rect 29316 11609 29372 11653
rect 28356 11513 28412 11577
rect 28996 11513 29052 11577
rect 28188 11500 28260 11513
rect 28188 11454 28201 11500
rect 28247 11454 28260 11500
rect 28188 11441 28260 11454
rect 28348 11500 28420 11513
rect 28348 11454 28361 11500
rect 28407 11454 28420 11500
rect 28348 11441 28420 11454
rect 28668 11500 28740 11513
rect 28668 11454 28681 11500
rect 28727 11454 28740 11500
rect 28668 11441 28740 11454
rect 28988 11500 29060 11513
rect 28988 11454 29001 11500
rect 29047 11454 29060 11500
rect 28988 11441 29060 11454
rect 29308 11500 29380 11513
rect 29308 11454 29321 11500
rect 29367 11454 29380 11500
rect 29308 11441 29380 11454
rect 28196 11317 28252 11441
rect 28676 11393 28732 11441
rect 28356 11317 28412 11361
rect 28516 11317 28572 11361
rect 28676 11337 28892 11393
rect 28676 11317 28732 11337
rect 28836 11317 28892 11337
rect 28996 11317 29052 11361
rect 29156 11317 29212 11361
rect 29316 11317 29372 11441
rect 29604 11317 29660 11653
rect 27908 10381 27964 10717
rect 28196 10381 28252 10717
rect 28356 10381 28412 10717
rect 28516 10381 28572 10717
rect 28676 10381 28732 10717
rect 28836 10381 28892 10717
rect 28996 10381 29052 10717
rect 29156 10381 29212 10717
rect 29316 10381 29372 10717
rect 29604 10381 29660 10717
rect 27908 9445 27964 9781
rect 28196 9737 28252 9781
rect 28356 9761 28412 9781
rect 28516 9761 28572 9781
rect 28356 9705 28572 9761
rect 28676 9737 28732 9781
rect 28836 9737 28892 9781
rect 28996 9761 29052 9781
rect 29156 9761 29212 9781
rect 28996 9705 29212 9761
rect 29316 9737 29372 9781
rect 28356 9641 28412 9705
rect 28996 9641 29052 9705
rect 28188 9628 28260 9641
rect 28188 9582 28201 9628
rect 28247 9582 28260 9628
rect 28188 9569 28260 9582
rect 28348 9628 28420 9641
rect 28348 9582 28361 9628
rect 28407 9582 28420 9628
rect 28348 9569 28420 9582
rect 28668 9628 28740 9641
rect 28668 9582 28681 9628
rect 28727 9582 28740 9628
rect 28668 9569 28740 9582
rect 28988 9628 29060 9641
rect 28988 9582 29001 9628
rect 29047 9582 29060 9628
rect 28988 9569 29060 9582
rect 29308 9628 29380 9641
rect 29308 9582 29321 9628
rect 29367 9582 29380 9628
rect 29308 9569 29380 9582
rect 28196 9445 28252 9569
rect 28676 9521 28732 9569
rect 28356 9445 28412 9489
rect 28516 9445 28572 9489
rect 28676 9465 28892 9521
rect 28676 9445 28732 9465
rect 28836 9445 28892 9465
rect 28996 9445 29052 9489
rect 29156 9445 29212 9489
rect 29316 9445 29372 9569
rect 29604 9445 29660 9781
rect 27908 8713 27964 8845
rect 28196 8801 28252 8845
rect 28356 8825 28412 8845
rect 28516 8825 28572 8845
rect 28356 8769 28572 8825
rect 28676 8801 28732 8845
rect 28836 8801 28892 8845
rect 28996 8825 29052 8845
rect 29156 8825 29212 8845
rect 28996 8769 29212 8825
rect 29316 8801 29372 8845
rect 27900 8700 27972 8713
rect 28356 8705 28412 8769
rect 28996 8705 29052 8769
rect 29604 8713 29660 8845
rect 27900 8654 27913 8700
rect 27959 8654 27972 8700
rect 27900 8641 27972 8654
rect 28188 8692 28260 8705
rect 28188 8646 28201 8692
rect 28247 8646 28260 8692
rect 27908 8509 27964 8641
rect 28188 8633 28260 8646
rect 28348 8692 28420 8705
rect 28348 8646 28361 8692
rect 28407 8646 28420 8692
rect 28348 8633 28420 8646
rect 28668 8692 28740 8705
rect 28668 8646 28681 8692
rect 28727 8646 28740 8692
rect 28668 8633 28740 8646
rect 28988 8692 29060 8705
rect 28988 8646 29001 8692
rect 29047 8646 29060 8692
rect 28988 8633 29060 8646
rect 29308 8692 29380 8705
rect 29308 8646 29321 8692
rect 29367 8646 29380 8692
rect 29308 8633 29380 8646
rect 29596 8700 29668 8713
rect 29596 8654 29609 8700
rect 29655 8654 29668 8700
rect 29596 8641 29668 8654
rect 28196 8509 28252 8633
rect 28676 8585 28732 8633
rect 28356 8509 28412 8553
rect 28516 8509 28572 8553
rect 28676 8529 28892 8585
rect 28676 8509 28732 8529
rect 28836 8509 28892 8529
rect 28996 8509 29052 8553
rect 29156 8509 29212 8553
rect 29316 8509 29372 8633
rect 29604 8509 29660 8641
rect 27908 7865 27964 7909
rect 28196 7865 28252 7909
rect 28356 7889 28412 7909
rect 28516 7889 28572 7909
rect 28356 7833 28572 7889
rect 28676 7865 28732 7909
rect 28836 7865 28892 7909
rect 28996 7889 29052 7909
rect 29156 7889 29212 7909
rect 28996 7833 29212 7889
rect 29316 7865 29372 7909
rect 29604 7865 29660 7909
rect 28356 7769 28412 7833
rect 28996 7769 29052 7833
rect 28348 7756 28420 7769
rect 28348 7710 28361 7756
rect 28407 7710 28420 7756
rect 28348 7697 28420 7710
rect 28988 7756 29060 7769
rect 28988 7710 29001 7756
rect 29047 7710 29060 7756
rect 28988 7697 29060 7710
rect 34604 11809 34676 11822
rect 34604 11763 34617 11809
rect 34663 11763 34676 11809
rect 34604 11750 34676 11763
rect 34764 11809 34836 11822
rect 34764 11763 34777 11809
rect 34823 11763 34836 11809
rect 34764 11750 34836 11763
rect 33204 11689 33260 11733
rect 33492 11689 33548 11733
rect 33652 11689 33708 11733
rect 33812 11689 33868 11733
rect 33972 11689 34028 11733
rect 34132 11689 34188 11733
rect 34292 11689 34348 11733
rect 34452 11689 34508 11733
rect 34612 11689 34668 11750
rect 34772 11689 34828 11750
rect 38740 11809 38812 11822
rect 38740 11763 38753 11809
rect 38799 11763 38812 11809
rect 38740 11750 38812 11763
rect 38900 11809 38972 11822
rect 38900 11763 38913 11809
rect 38959 11763 38972 11809
rect 38900 11750 38972 11763
rect 34932 11689 34988 11733
rect 35092 11689 35148 11733
rect 35252 11689 35308 11733
rect 35412 11689 35468 11733
rect 35572 11689 35628 11733
rect 35732 11689 35788 11733
rect 35892 11689 35948 11733
rect 36180 11689 36236 11733
rect 37340 11689 37396 11733
rect 37628 11689 37684 11733
rect 37788 11689 37844 11733
rect 37948 11689 38004 11733
rect 38108 11689 38164 11733
rect 38268 11689 38324 11733
rect 38428 11689 38484 11733
rect 38588 11689 38644 11733
rect 38748 11689 38804 11750
rect 38908 11689 38964 11750
rect 39068 11689 39124 11733
rect 39228 11689 39284 11733
rect 39388 11689 39444 11733
rect 39548 11689 39604 11733
rect 39708 11689 39764 11733
rect 39868 11689 39924 11733
rect 40028 11689 40084 11733
rect 40316 11689 40372 11733
rect 33204 10895 33260 11089
rect 33196 10882 33268 10895
rect 33196 10836 33209 10882
rect 33255 10836 33268 10882
rect 33196 10823 33268 10836
rect 33204 10629 33260 10823
rect 33492 10762 33548 11089
rect 33652 10762 33708 11089
rect 33812 10762 33868 11089
rect 33972 10762 34028 11089
rect 34132 10762 34188 11089
rect 34292 10762 34348 11089
rect 34452 10762 34508 11089
rect 34612 10762 34668 11089
rect 34772 10762 34828 11089
rect 34932 10762 34988 11089
rect 35092 10762 35148 11089
rect 35252 10762 35308 11089
rect 35412 10762 35468 11089
rect 35572 10762 35628 11089
rect 35732 10762 35788 11089
rect 35892 10762 35948 11089
rect 36180 10895 36236 11089
rect 36172 10882 36244 10895
rect 36172 10836 36185 10882
rect 36231 10836 36244 10882
rect 36172 10823 36244 10836
rect 37340 10895 37396 11089
rect 33492 10749 35948 10762
rect 33492 10703 34617 10749
rect 34663 10703 34777 10749
rect 34823 10703 35948 10749
rect 33492 10690 35948 10703
rect 33492 10629 33548 10690
rect 33652 10629 33708 10690
rect 33812 10629 33868 10690
rect 33972 10629 34028 10690
rect 34132 10629 34188 10690
rect 34292 10629 34348 10690
rect 34452 10629 34508 10690
rect 34612 10629 34668 10690
rect 34772 10629 34828 10690
rect 34932 10629 34988 10690
rect 35092 10629 35148 10690
rect 35252 10629 35308 10690
rect 35412 10629 35468 10690
rect 35572 10629 35628 10690
rect 35732 10629 35788 10690
rect 35892 10629 35948 10690
rect 36180 10629 36236 10823
rect 37332 10882 37404 10895
rect 37332 10836 37345 10882
rect 37391 10836 37404 10882
rect 37332 10823 37404 10836
rect 37340 10629 37396 10823
rect 37628 10762 37684 11089
rect 37788 10762 37844 11089
rect 37948 10762 38004 11089
rect 38108 10762 38164 11089
rect 38268 10762 38324 11089
rect 38428 10762 38484 11089
rect 38588 10762 38644 11089
rect 38748 10762 38804 11089
rect 38908 10762 38964 11089
rect 39068 10762 39124 11089
rect 39228 10762 39284 11089
rect 39388 10762 39444 11089
rect 39548 10762 39604 11089
rect 39708 10762 39764 11089
rect 39868 10762 39924 11089
rect 40028 10762 40084 11089
rect 40316 10895 40372 11089
rect 40308 10882 40380 10895
rect 40308 10836 40321 10882
rect 40367 10836 40380 10882
rect 40308 10823 40380 10836
rect 37628 10749 40084 10762
rect 37628 10703 38753 10749
rect 38799 10703 38913 10749
rect 38959 10703 40084 10749
rect 37628 10690 40084 10703
rect 37628 10629 37684 10690
rect 37788 10629 37844 10690
rect 37948 10629 38004 10690
rect 38108 10629 38164 10690
rect 38268 10629 38324 10690
rect 38428 10629 38484 10690
rect 38588 10629 38644 10690
rect 38748 10629 38804 10690
rect 38908 10629 38964 10690
rect 39068 10629 39124 10690
rect 39228 10629 39284 10690
rect 39388 10629 39444 10690
rect 39548 10629 39604 10690
rect 39708 10629 39764 10690
rect 39868 10629 39924 10690
rect 40028 10629 40084 10690
rect 40316 10629 40372 10823
rect 33204 9569 33260 10029
rect 33492 9702 33548 10029
rect 33652 9702 33708 10029
rect 33812 9702 33868 10029
rect 33972 9702 34028 10029
rect 34132 9702 34188 10029
rect 34292 9702 34348 10029
rect 34452 9702 34508 10029
rect 34612 9702 34668 10029
rect 34772 9702 34828 10029
rect 34932 9702 34988 10029
rect 35092 9702 35148 10029
rect 35252 9702 35308 10029
rect 35412 9702 35468 10029
rect 35572 9702 35628 10029
rect 35732 9702 35788 10029
rect 35892 9702 35948 10029
rect 33492 9689 35948 9702
rect 33492 9643 34617 9689
rect 34663 9643 34777 9689
rect 34823 9643 35948 9689
rect 33492 9630 35948 9643
rect 33492 9569 33548 9630
rect 33652 9569 33708 9630
rect 33812 9569 33868 9630
rect 33972 9569 34028 9630
rect 34132 9569 34188 9630
rect 34292 9569 34348 9630
rect 34452 9569 34508 9630
rect 34612 9569 34668 9630
rect 34772 9569 34828 9630
rect 34932 9569 34988 9630
rect 35092 9569 35148 9630
rect 35252 9569 35308 9630
rect 35412 9569 35468 9630
rect 35572 9569 35628 9630
rect 35732 9569 35788 9630
rect 35892 9569 35948 9630
rect 36180 9569 36236 10029
rect 37340 9569 37396 10029
rect 37628 9702 37684 10029
rect 37788 9702 37844 10029
rect 37948 9702 38004 10029
rect 38108 9702 38164 10029
rect 38268 9702 38324 10029
rect 38428 9702 38484 10029
rect 38588 9702 38644 10029
rect 38748 9702 38804 10029
rect 38908 9702 38964 10029
rect 39068 9702 39124 10029
rect 39228 9702 39284 10029
rect 39388 9702 39444 10029
rect 39548 9702 39604 10029
rect 39708 9702 39764 10029
rect 39868 9702 39924 10029
rect 40028 9702 40084 10029
rect 37628 9689 40084 9702
rect 37628 9643 38753 9689
rect 38799 9643 38913 9689
rect 38959 9643 40084 9689
rect 37628 9630 40084 9643
rect 37628 9569 37684 9630
rect 37788 9569 37844 9630
rect 37948 9569 38004 9630
rect 38108 9569 38164 9630
rect 38268 9569 38324 9630
rect 38428 9569 38484 9630
rect 38588 9569 38644 9630
rect 38748 9569 38804 9630
rect 38908 9569 38964 9630
rect 39068 9569 39124 9630
rect 39228 9569 39284 9630
rect 39388 9569 39444 9630
rect 39548 9569 39604 9630
rect 39708 9569 39764 9630
rect 39868 9569 39924 9630
rect 40028 9569 40084 9630
rect 40316 9569 40372 10029
rect 33204 8775 33260 8969
rect 33196 8762 33268 8775
rect 33196 8716 33209 8762
rect 33255 8716 33268 8762
rect 33196 8703 33268 8716
rect 33204 8509 33260 8703
rect 33492 8642 33548 8969
rect 33652 8642 33708 8969
rect 33812 8642 33868 8969
rect 33972 8642 34028 8969
rect 34132 8642 34188 8969
rect 34292 8642 34348 8969
rect 34452 8642 34508 8969
rect 34612 8642 34668 8969
rect 34772 8642 34828 8969
rect 34932 8642 34988 8969
rect 35092 8642 35148 8969
rect 35252 8642 35308 8969
rect 35412 8642 35468 8969
rect 35572 8642 35628 8969
rect 35732 8642 35788 8969
rect 35892 8642 35948 8969
rect 36180 8775 36236 8969
rect 36172 8762 36244 8775
rect 36172 8716 36185 8762
rect 36231 8716 36244 8762
rect 36172 8703 36244 8716
rect 37340 8775 37396 8969
rect 33492 8629 35948 8642
rect 33492 8583 34617 8629
rect 34663 8583 34777 8629
rect 34823 8583 35948 8629
rect 33492 8570 35948 8583
rect 33492 8509 33548 8570
rect 33652 8509 33708 8570
rect 33812 8509 33868 8570
rect 33972 8509 34028 8570
rect 34132 8509 34188 8570
rect 34292 8509 34348 8570
rect 34452 8509 34508 8570
rect 34612 8509 34668 8570
rect 34772 8509 34828 8570
rect 34932 8509 34988 8570
rect 35092 8509 35148 8570
rect 35252 8509 35308 8570
rect 35412 8509 35468 8570
rect 35572 8509 35628 8570
rect 35732 8509 35788 8570
rect 35892 8509 35948 8570
rect 36180 8509 36236 8703
rect 37332 8762 37404 8775
rect 37332 8716 37345 8762
rect 37391 8716 37404 8762
rect 37332 8703 37404 8716
rect 37340 8509 37396 8703
rect 37628 8642 37684 8969
rect 37788 8642 37844 8969
rect 37948 8642 38004 8969
rect 38108 8642 38164 8969
rect 38268 8642 38324 8969
rect 38428 8642 38484 8969
rect 38588 8642 38644 8969
rect 38748 8642 38804 8969
rect 38908 8642 38964 8969
rect 39068 8642 39124 8969
rect 39228 8642 39284 8969
rect 39388 8642 39444 8969
rect 39548 8642 39604 8969
rect 39708 8642 39764 8969
rect 39868 8642 39924 8969
rect 40028 8642 40084 8969
rect 40316 8775 40372 8969
rect 40308 8762 40380 8775
rect 40308 8716 40321 8762
rect 40367 8716 40380 8762
rect 40308 8703 40380 8716
rect 37628 8629 40084 8642
rect 37628 8583 38753 8629
rect 38799 8583 38913 8629
rect 38959 8583 40084 8629
rect 37628 8570 40084 8583
rect 37628 8509 37684 8570
rect 37788 8509 37844 8570
rect 37948 8509 38004 8570
rect 38108 8509 38164 8570
rect 38268 8509 38324 8570
rect 38428 8509 38484 8570
rect 38588 8509 38644 8570
rect 38748 8509 38804 8570
rect 38908 8509 38964 8570
rect 39068 8509 39124 8570
rect 39228 8509 39284 8570
rect 39388 8509 39444 8570
rect 39548 8509 39604 8570
rect 39708 8509 39764 8570
rect 39868 8509 39924 8570
rect 40028 8509 40084 8570
rect 40316 8509 40372 8703
rect 33204 7865 33260 7909
rect 33492 7865 33548 7909
rect 33652 7865 33708 7909
rect 33812 7865 33868 7909
rect 33972 7865 34028 7909
rect 34132 7865 34188 7909
rect 34292 7865 34348 7909
rect 34452 7865 34508 7909
rect 34612 7865 34668 7909
rect 34772 7865 34828 7909
rect 34932 7865 34988 7909
rect 35092 7865 35148 7909
rect 35252 7865 35308 7909
rect 35412 7865 35468 7909
rect 35572 7865 35628 7909
rect 35732 7865 35788 7909
rect 35892 7865 35948 7909
rect 36180 7865 36236 7909
rect 37340 7865 37396 7909
rect 37628 7865 37684 7909
rect 37788 7865 37844 7909
rect 37948 7865 38004 7909
rect 38108 7865 38164 7909
rect 38268 7865 38324 7909
rect 38428 7865 38484 7909
rect 38588 7865 38644 7909
rect 38748 7865 38804 7909
rect 38908 7865 38964 7909
rect 39068 7865 39124 7909
rect 39228 7865 39284 7909
rect 39388 7865 39444 7909
rect 39548 7865 39604 7909
rect 39708 7865 39764 7909
rect 39868 7865 39924 7909
rect 40028 7865 40084 7909
rect 40316 7865 40372 7909
rect 44300 11809 44372 11822
rect 44300 11763 44313 11809
rect 44359 11763 44372 11809
rect 44300 11750 44372 11763
rect 44460 11809 44532 11822
rect 44460 11763 44473 11809
rect 44519 11763 44532 11809
rect 44460 11750 44532 11763
rect 42900 11689 42956 11733
rect 43188 11689 43244 11733
rect 43348 11689 43404 11733
rect 43508 11689 43564 11733
rect 43668 11689 43724 11733
rect 43828 11689 43884 11733
rect 43988 11689 44044 11733
rect 44148 11689 44204 11733
rect 44308 11689 44364 11750
rect 44468 11689 44524 11750
rect 48436 11809 48508 11822
rect 48436 11763 48449 11809
rect 48495 11763 48508 11809
rect 48436 11750 48508 11763
rect 48596 11809 48668 11822
rect 48596 11763 48609 11809
rect 48655 11763 48668 11809
rect 48596 11750 48668 11763
rect 44628 11689 44684 11733
rect 44788 11689 44844 11733
rect 44948 11689 45004 11733
rect 45108 11689 45164 11733
rect 45268 11689 45324 11733
rect 45428 11689 45484 11733
rect 45588 11689 45644 11733
rect 45876 11689 45932 11733
rect 47036 11689 47092 11733
rect 47324 11689 47380 11733
rect 47484 11689 47540 11733
rect 47644 11689 47700 11733
rect 47804 11689 47860 11733
rect 47964 11689 48020 11733
rect 48124 11689 48180 11733
rect 48284 11689 48340 11733
rect 48444 11689 48500 11750
rect 48604 11689 48660 11750
rect 48764 11689 48820 11733
rect 48924 11689 48980 11733
rect 49084 11689 49140 11733
rect 49244 11689 49300 11733
rect 49404 11689 49460 11733
rect 49564 11689 49620 11733
rect 49724 11689 49780 11733
rect 50012 11689 50068 11733
rect 42900 10895 42956 11089
rect 42892 10882 42964 10895
rect 42892 10836 42905 10882
rect 42951 10836 42964 10882
rect 42892 10823 42964 10836
rect 42900 10629 42956 10823
rect 43188 10762 43244 11089
rect 43348 10762 43404 11089
rect 43508 10762 43564 11089
rect 43668 10762 43724 11089
rect 43828 10762 43884 11089
rect 43988 10762 44044 11089
rect 44148 10762 44204 11089
rect 44308 10762 44364 11089
rect 44468 10762 44524 11089
rect 44628 10762 44684 11089
rect 44788 10762 44844 11089
rect 44948 10762 45004 11089
rect 45108 10762 45164 11089
rect 45268 10762 45324 11089
rect 45428 10762 45484 11089
rect 45588 10762 45644 11089
rect 45876 10895 45932 11089
rect 45868 10882 45940 10895
rect 45868 10836 45881 10882
rect 45927 10836 45940 10882
rect 45868 10823 45940 10836
rect 47036 10895 47092 11089
rect 43188 10749 45644 10762
rect 43188 10703 44313 10749
rect 44359 10703 44473 10749
rect 44519 10703 45644 10749
rect 43188 10690 45644 10703
rect 43188 10629 43244 10690
rect 43348 10629 43404 10690
rect 43508 10629 43564 10690
rect 43668 10629 43724 10690
rect 43828 10629 43884 10690
rect 43988 10629 44044 10690
rect 44148 10629 44204 10690
rect 44308 10629 44364 10690
rect 44468 10629 44524 10690
rect 44628 10629 44684 10690
rect 44788 10629 44844 10690
rect 44948 10629 45004 10690
rect 45108 10629 45164 10690
rect 45268 10629 45324 10690
rect 45428 10629 45484 10690
rect 45588 10629 45644 10690
rect 45876 10629 45932 10823
rect 47028 10882 47100 10895
rect 47028 10836 47041 10882
rect 47087 10836 47100 10882
rect 47028 10823 47100 10836
rect 47036 10629 47092 10823
rect 47324 10762 47380 11089
rect 47484 10762 47540 11089
rect 47644 10762 47700 11089
rect 47804 10762 47860 11089
rect 47964 10762 48020 11089
rect 48124 10762 48180 11089
rect 48284 10762 48340 11089
rect 48444 10762 48500 11089
rect 48604 10762 48660 11089
rect 48764 10762 48820 11089
rect 48924 10762 48980 11089
rect 49084 10762 49140 11089
rect 49244 10762 49300 11089
rect 49404 10762 49460 11089
rect 49564 10762 49620 11089
rect 49724 10762 49780 11089
rect 50012 10895 50068 11089
rect 50004 10882 50076 10895
rect 50004 10836 50017 10882
rect 50063 10836 50076 10882
rect 50004 10823 50076 10836
rect 47324 10749 49780 10762
rect 47324 10703 48449 10749
rect 48495 10703 48609 10749
rect 48655 10703 49780 10749
rect 47324 10690 49780 10703
rect 47324 10629 47380 10690
rect 47484 10629 47540 10690
rect 47644 10629 47700 10690
rect 47804 10629 47860 10690
rect 47964 10629 48020 10690
rect 48124 10629 48180 10690
rect 48284 10629 48340 10690
rect 48444 10629 48500 10690
rect 48604 10629 48660 10690
rect 48764 10629 48820 10690
rect 48924 10629 48980 10690
rect 49084 10629 49140 10690
rect 49244 10629 49300 10690
rect 49404 10629 49460 10690
rect 49564 10629 49620 10690
rect 49724 10629 49780 10690
rect 50012 10629 50068 10823
rect 42900 9569 42956 10029
rect 43188 9702 43244 10029
rect 43348 9702 43404 10029
rect 43508 9702 43564 10029
rect 43668 9702 43724 10029
rect 43828 9702 43884 10029
rect 43988 9702 44044 10029
rect 44148 9702 44204 10029
rect 44308 9702 44364 10029
rect 44468 9702 44524 10029
rect 44628 9702 44684 10029
rect 44788 9702 44844 10029
rect 44948 9702 45004 10029
rect 45108 9702 45164 10029
rect 45268 9702 45324 10029
rect 45428 9702 45484 10029
rect 45588 9702 45644 10029
rect 43188 9689 45644 9702
rect 43188 9643 44313 9689
rect 44359 9643 44473 9689
rect 44519 9643 45644 9689
rect 43188 9630 45644 9643
rect 43188 9569 43244 9630
rect 43348 9569 43404 9630
rect 43508 9569 43564 9630
rect 43668 9569 43724 9630
rect 43828 9569 43884 9630
rect 43988 9569 44044 9630
rect 44148 9569 44204 9630
rect 44308 9569 44364 9630
rect 44468 9569 44524 9630
rect 44628 9569 44684 9630
rect 44788 9569 44844 9630
rect 44948 9569 45004 9630
rect 45108 9569 45164 9630
rect 45268 9569 45324 9630
rect 45428 9569 45484 9630
rect 45588 9569 45644 9630
rect 45876 9569 45932 10029
rect 47036 9569 47092 10029
rect 47324 9702 47380 10029
rect 47484 9702 47540 10029
rect 47644 9702 47700 10029
rect 47804 9702 47860 10029
rect 47964 9702 48020 10029
rect 48124 9702 48180 10029
rect 48284 9702 48340 10029
rect 48444 9702 48500 10029
rect 48604 9702 48660 10029
rect 48764 9702 48820 10029
rect 48924 9702 48980 10029
rect 49084 9702 49140 10029
rect 49244 9702 49300 10029
rect 49404 9702 49460 10029
rect 49564 9702 49620 10029
rect 49724 9702 49780 10029
rect 47324 9689 49780 9702
rect 47324 9643 48449 9689
rect 48495 9643 48609 9689
rect 48655 9643 49780 9689
rect 47324 9630 49780 9643
rect 47324 9569 47380 9630
rect 47484 9569 47540 9630
rect 47644 9569 47700 9630
rect 47804 9569 47860 9630
rect 47964 9569 48020 9630
rect 48124 9569 48180 9630
rect 48284 9569 48340 9630
rect 48444 9569 48500 9630
rect 48604 9569 48660 9630
rect 48764 9569 48820 9630
rect 48924 9569 48980 9630
rect 49084 9569 49140 9630
rect 49244 9569 49300 9630
rect 49404 9569 49460 9630
rect 49564 9569 49620 9630
rect 49724 9569 49780 9630
rect 50012 9569 50068 10029
rect 42900 8775 42956 8969
rect 42892 8762 42964 8775
rect 42892 8716 42905 8762
rect 42951 8716 42964 8762
rect 42892 8703 42964 8716
rect 42900 8509 42956 8703
rect 43188 8642 43244 8969
rect 43348 8642 43404 8969
rect 43508 8642 43564 8969
rect 43668 8642 43724 8969
rect 43828 8642 43884 8969
rect 43988 8642 44044 8969
rect 44148 8642 44204 8969
rect 44308 8642 44364 8969
rect 44468 8642 44524 8969
rect 44628 8642 44684 8969
rect 44788 8642 44844 8969
rect 44948 8642 45004 8969
rect 45108 8642 45164 8969
rect 45268 8642 45324 8969
rect 45428 8642 45484 8969
rect 45588 8642 45644 8969
rect 45876 8775 45932 8969
rect 45868 8762 45940 8775
rect 45868 8716 45881 8762
rect 45927 8716 45940 8762
rect 45868 8703 45940 8716
rect 47036 8775 47092 8969
rect 43188 8629 45644 8642
rect 43188 8583 44313 8629
rect 44359 8583 44473 8629
rect 44519 8583 45644 8629
rect 43188 8570 45644 8583
rect 43188 8509 43244 8570
rect 43348 8509 43404 8570
rect 43508 8509 43564 8570
rect 43668 8509 43724 8570
rect 43828 8509 43884 8570
rect 43988 8509 44044 8570
rect 44148 8509 44204 8570
rect 44308 8509 44364 8570
rect 44468 8509 44524 8570
rect 44628 8509 44684 8570
rect 44788 8509 44844 8570
rect 44948 8509 45004 8570
rect 45108 8509 45164 8570
rect 45268 8509 45324 8570
rect 45428 8509 45484 8570
rect 45588 8509 45644 8570
rect 45876 8509 45932 8703
rect 47028 8762 47100 8775
rect 47028 8716 47041 8762
rect 47087 8716 47100 8762
rect 47028 8703 47100 8716
rect 47036 8509 47092 8703
rect 47324 8642 47380 8969
rect 47484 8642 47540 8969
rect 47644 8642 47700 8969
rect 47804 8642 47860 8969
rect 47964 8642 48020 8969
rect 48124 8642 48180 8969
rect 48284 8642 48340 8969
rect 48444 8642 48500 8969
rect 48604 8642 48660 8969
rect 48764 8642 48820 8969
rect 48924 8642 48980 8969
rect 49084 8642 49140 8969
rect 49244 8642 49300 8969
rect 49404 8642 49460 8969
rect 49564 8642 49620 8969
rect 49724 8642 49780 8969
rect 50012 8775 50068 8969
rect 50004 8762 50076 8775
rect 50004 8716 50017 8762
rect 50063 8716 50076 8762
rect 50004 8703 50076 8716
rect 47324 8629 49780 8642
rect 47324 8583 48449 8629
rect 48495 8583 48609 8629
rect 48655 8583 49780 8629
rect 47324 8570 49780 8583
rect 47324 8509 47380 8570
rect 47484 8509 47540 8570
rect 47644 8509 47700 8570
rect 47804 8509 47860 8570
rect 47964 8509 48020 8570
rect 48124 8509 48180 8570
rect 48284 8509 48340 8570
rect 48444 8509 48500 8570
rect 48604 8509 48660 8570
rect 48764 8509 48820 8570
rect 48924 8509 48980 8570
rect 49084 8509 49140 8570
rect 49244 8509 49300 8570
rect 49404 8509 49460 8570
rect 49564 8509 49620 8570
rect 49724 8509 49780 8570
rect 50012 8509 50068 8703
rect 42900 7865 42956 7909
rect 43188 7865 43244 7909
rect 43348 7865 43404 7909
rect 43508 7865 43564 7909
rect 43668 7865 43724 7909
rect 43828 7865 43884 7909
rect 43988 7865 44044 7909
rect 44148 7865 44204 7909
rect 44308 7865 44364 7909
rect 44468 7865 44524 7909
rect 44628 7865 44684 7909
rect 44788 7865 44844 7909
rect 44948 7865 45004 7909
rect 45108 7865 45164 7909
rect 45268 7865 45324 7909
rect 45428 7865 45484 7909
rect 45588 7865 45644 7909
rect 45876 7865 45932 7909
rect 47036 7865 47092 7909
rect 47324 7865 47380 7909
rect 47484 7865 47540 7909
rect 47644 7865 47700 7909
rect 47804 7865 47860 7909
rect 47964 7865 48020 7909
rect 48124 7865 48180 7909
rect 48284 7865 48340 7909
rect 48444 7865 48500 7909
rect 48604 7865 48660 7909
rect 48764 7865 48820 7909
rect 48924 7865 48980 7909
rect 49084 7865 49140 7909
rect 49244 7865 49300 7909
rect 49404 7865 49460 7909
rect 49564 7865 49620 7909
rect 49724 7865 49780 7909
rect 50012 7865 50068 7909
rect 53996 11809 54068 11822
rect 53996 11763 54009 11809
rect 54055 11763 54068 11809
rect 53996 11750 54068 11763
rect 54156 11809 54228 11822
rect 54156 11763 54169 11809
rect 54215 11763 54228 11809
rect 54156 11750 54228 11763
rect 52596 11689 52652 11733
rect 52884 11689 52940 11733
rect 53044 11689 53100 11733
rect 53204 11689 53260 11733
rect 53364 11689 53420 11733
rect 53524 11689 53580 11733
rect 53684 11689 53740 11733
rect 53844 11689 53900 11733
rect 54004 11689 54060 11750
rect 54164 11689 54220 11750
rect 58132 11809 58204 11822
rect 58132 11763 58145 11809
rect 58191 11763 58204 11809
rect 58132 11750 58204 11763
rect 58292 11809 58364 11822
rect 58292 11763 58305 11809
rect 58351 11763 58364 11809
rect 58292 11750 58364 11763
rect 54324 11689 54380 11733
rect 54484 11689 54540 11733
rect 54644 11689 54700 11733
rect 54804 11689 54860 11733
rect 54964 11689 55020 11733
rect 55124 11689 55180 11733
rect 55284 11689 55340 11733
rect 55572 11689 55628 11733
rect 56732 11689 56788 11733
rect 57020 11689 57076 11733
rect 57180 11689 57236 11733
rect 57340 11689 57396 11733
rect 57500 11689 57556 11733
rect 57660 11689 57716 11733
rect 57820 11689 57876 11733
rect 57980 11689 58036 11733
rect 58140 11689 58196 11750
rect 58300 11689 58356 11750
rect 58460 11689 58516 11733
rect 58620 11689 58676 11733
rect 58780 11689 58836 11733
rect 58940 11689 58996 11733
rect 59100 11689 59156 11733
rect 59260 11689 59316 11733
rect 59420 11689 59476 11733
rect 59708 11689 59764 11733
rect 52596 10895 52652 11089
rect 52588 10882 52660 10895
rect 52588 10836 52601 10882
rect 52647 10836 52660 10882
rect 52588 10823 52660 10836
rect 52596 10629 52652 10823
rect 52884 10762 52940 11089
rect 53044 10762 53100 11089
rect 53204 10762 53260 11089
rect 53364 10762 53420 11089
rect 53524 10762 53580 11089
rect 53684 10762 53740 11089
rect 53844 10762 53900 11089
rect 54004 10762 54060 11089
rect 54164 10762 54220 11089
rect 54324 10762 54380 11089
rect 54484 10762 54540 11089
rect 54644 10762 54700 11089
rect 54804 10762 54860 11089
rect 54964 10762 55020 11089
rect 55124 10762 55180 11089
rect 55284 10762 55340 11089
rect 55572 10895 55628 11089
rect 55564 10882 55636 10895
rect 55564 10836 55577 10882
rect 55623 10836 55636 10882
rect 55564 10823 55636 10836
rect 56732 10895 56788 11089
rect 52884 10749 55340 10762
rect 52884 10703 54009 10749
rect 54055 10703 54169 10749
rect 54215 10703 55340 10749
rect 52884 10690 55340 10703
rect 52884 10629 52940 10690
rect 53044 10629 53100 10690
rect 53204 10629 53260 10690
rect 53364 10629 53420 10690
rect 53524 10629 53580 10690
rect 53684 10629 53740 10690
rect 53844 10629 53900 10690
rect 54004 10629 54060 10690
rect 54164 10629 54220 10690
rect 54324 10629 54380 10690
rect 54484 10629 54540 10690
rect 54644 10629 54700 10690
rect 54804 10629 54860 10690
rect 54964 10629 55020 10690
rect 55124 10629 55180 10690
rect 55284 10629 55340 10690
rect 55572 10629 55628 10823
rect 56724 10882 56796 10895
rect 56724 10836 56737 10882
rect 56783 10836 56796 10882
rect 56724 10823 56796 10836
rect 56732 10629 56788 10823
rect 57020 10762 57076 11089
rect 57180 10762 57236 11089
rect 57340 10762 57396 11089
rect 57500 10762 57556 11089
rect 57660 10762 57716 11089
rect 57820 10762 57876 11089
rect 57980 10762 58036 11089
rect 58140 10762 58196 11089
rect 58300 10762 58356 11089
rect 58460 10762 58516 11089
rect 58620 10762 58676 11089
rect 58780 10762 58836 11089
rect 58940 10762 58996 11089
rect 59100 10762 59156 11089
rect 59260 10762 59316 11089
rect 59420 10762 59476 11089
rect 59708 10895 59764 11089
rect 59700 10882 59772 10895
rect 59700 10836 59713 10882
rect 59759 10836 59772 10882
rect 59700 10823 59772 10836
rect 57020 10749 59476 10762
rect 57020 10703 58145 10749
rect 58191 10703 58305 10749
rect 58351 10703 59476 10749
rect 57020 10690 59476 10703
rect 57020 10629 57076 10690
rect 57180 10629 57236 10690
rect 57340 10629 57396 10690
rect 57500 10629 57556 10690
rect 57660 10629 57716 10690
rect 57820 10629 57876 10690
rect 57980 10629 58036 10690
rect 58140 10629 58196 10690
rect 58300 10629 58356 10690
rect 58460 10629 58516 10690
rect 58620 10629 58676 10690
rect 58780 10629 58836 10690
rect 58940 10629 58996 10690
rect 59100 10629 59156 10690
rect 59260 10629 59316 10690
rect 59420 10629 59476 10690
rect 59708 10629 59764 10823
rect 52596 9569 52652 10029
rect 52884 9702 52940 10029
rect 53044 9702 53100 10029
rect 53204 9702 53260 10029
rect 53364 9702 53420 10029
rect 53524 9702 53580 10029
rect 53684 9702 53740 10029
rect 53844 9702 53900 10029
rect 54004 9702 54060 10029
rect 54164 9702 54220 10029
rect 54324 9702 54380 10029
rect 54484 9702 54540 10029
rect 54644 9702 54700 10029
rect 54804 9702 54860 10029
rect 54964 9702 55020 10029
rect 55124 9702 55180 10029
rect 55284 9702 55340 10029
rect 52884 9689 55340 9702
rect 52884 9643 54009 9689
rect 54055 9643 54169 9689
rect 54215 9643 55340 9689
rect 52884 9630 55340 9643
rect 52884 9569 52940 9630
rect 53044 9569 53100 9630
rect 53204 9569 53260 9630
rect 53364 9569 53420 9630
rect 53524 9569 53580 9630
rect 53684 9569 53740 9630
rect 53844 9569 53900 9630
rect 54004 9569 54060 9630
rect 54164 9569 54220 9630
rect 54324 9569 54380 9630
rect 54484 9569 54540 9630
rect 54644 9569 54700 9630
rect 54804 9569 54860 9630
rect 54964 9569 55020 9630
rect 55124 9569 55180 9630
rect 55284 9569 55340 9630
rect 55572 9569 55628 10029
rect 56732 9569 56788 10029
rect 57020 9702 57076 10029
rect 57180 9702 57236 10029
rect 57340 9702 57396 10029
rect 57500 9702 57556 10029
rect 57660 9702 57716 10029
rect 57820 9702 57876 10029
rect 57980 9702 58036 10029
rect 58140 9702 58196 10029
rect 58300 9702 58356 10029
rect 58460 9702 58516 10029
rect 58620 9702 58676 10029
rect 58780 9702 58836 10029
rect 58940 9702 58996 10029
rect 59100 9702 59156 10029
rect 59260 9702 59316 10029
rect 59420 9702 59476 10029
rect 57020 9689 59476 9702
rect 57020 9643 58145 9689
rect 58191 9643 58305 9689
rect 58351 9643 59476 9689
rect 57020 9630 59476 9643
rect 57020 9569 57076 9630
rect 57180 9569 57236 9630
rect 57340 9569 57396 9630
rect 57500 9569 57556 9630
rect 57660 9569 57716 9630
rect 57820 9569 57876 9630
rect 57980 9569 58036 9630
rect 58140 9569 58196 9630
rect 58300 9569 58356 9630
rect 58460 9569 58516 9630
rect 58620 9569 58676 9630
rect 58780 9569 58836 9630
rect 58940 9569 58996 9630
rect 59100 9569 59156 9630
rect 59260 9569 59316 9630
rect 59420 9569 59476 9630
rect 59708 9569 59764 10029
rect 52596 8775 52652 8969
rect 52588 8762 52660 8775
rect 52588 8716 52601 8762
rect 52647 8716 52660 8762
rect 52588 8703 52660 8716
rect 52596 8509 52652 8703
rect 52884 8642 52940 8969
rect 53044 8642 53100 8969
rect 53204 8642 53260 8969
rect 53364 8642 53420 8969
rect 53524 8642 53580 8969
rect 53684 8642 53740 8969
rect 53844 8642 53900 8969
rect 54004 8642 54060 8969
rect 54164 8642 54220 8969
rect 54324 8642 54380 8969
rect 54484 8642 54540 8969
rect 54644 8642 54700 8969
rect 54804 8642 54860 8969
rect 54964 8642 55020 8969
rect 55124 8642 55180 8969
rect 55284 8642 55340 8969
rect 55572 8775 55628 8969
rect 55564 8762 55636 8775
rect 55564 8716 55577 8762
rect 55623 8716 55636 8762
rect 55564 8703 55636 8716
rect 56732 8775 56788 8969
rect 52884 8629 55340 8642
rect 52884 8583 54009 8629
rect 54055 8583 54169 8629
rect 54215 8583 55340 8629
rect 52884 8570 55340 8583
rect 52884 8509 52940 8570
rect 53044 8509 53100 8570
rect 53204 8509 53260 8570
rect 53364 8509 53420 8570
rect 53524 8509 53580 8570
rect 53684 8509 53740 8570
rect 53844 8509 53900 8570
rect 54004 8509 54060 8570
rect 54164 8509 54220 8570
rect 54324 8509 54380 8570
rect 54484 8509 54540 8570
rect 54644 8509 54700 8570
rect 54804 8509 54860 8570
rect 54964 8509 55020 8570
rect 55124 8509 55180 8570
rect 55284 8509 55340 8570
rect 55572 8509 55628 8703
rect 56724 8762 56796 8775
rect 56724 8716 56737 8762
rect 56783 8716 56796 8762
rect 56724 8703 56796 8716
rect 56732 8509 56788 8703
rect 57020 8642 57076 8969
rect 57180 8642 57236 8969
rect 57340 8642 57396 8969
rect 57500 8642 57556 8969
rect 57660 8642 57716 8969
rect 57820 8642 57876 8969
rect 57980 8642 58036 8969
rect 58140 8642 58196 8969
rect 58300 8642 58356 8969
rect 58460 8642 58516 8969
rect 58620 8642 58676 8969
rect 58780 8642 58836 8969
rect 58940 8642 58996 8969
rect 59100 8642 59156 8969
rect 59260 8642 59316 8969
rect 59420 8642 59476 8969
rect 59708 8775 59764 8969
rect 59700 8762 59772 8775
rect 59700 8716 59713 8762
rect 59759 8716 59772 8762
rect 59700 8703 59772 8716
rect 57020 8629 59476 8642
rect 57020 8583 58145 8629
rect 58191 8583 58305 8629
rect 58351 8583 59476 8629
rect 57020 8570 59476 8583
rect 57020 8509 57076 8570
rect 57180 8509 57236 8570
rect 57340 8509 57396 8570
rect 57500 8509 57556 8570
rect 57660 8509 57716 8570
rect 57820 8509 57876 8570
rect 57980 8509 58036 8570
rect 58140 8509 58196 8570
rect 58300 8509 58356 8570
rect 58460 8509 58516 8570
rect 58620 8509 58676 8570
rect 58780 8509 58836 8570
rect 58940 8509 58996 8570
rect 59100 8509 59156 8570
rect 59260 8509 59316 8570
rect 59420 8509 59476 8570
rect 59708 8509 59764 8703
rect 52596 7865 52652 7909
rect 52884 7865 52940 7909
rect 53044 7865 53100 7909
rect 53204 7865 53260 7909
rect 53364 7865 53420 7909
rect 53524 7865 53580 7909
rect 53684 7865 53740 7909
rect 53844 7865 53900 7909
rect 54004 7865 54060 7909
rect 54164 7865 54220 7909
rect 54324 7865 54380 7909
rect 54484 7865 54540 7909
rect 54644 7865 54700 7909
rect 54804 7865 54860 7909
rect 54964 7865 55020 7909
rect 55124 7865 55180 7909
rect 55284 7865 55340 7909
rect 55572 7865 55628 7909
rect 56732 7865 56788 7909
rect 57020 7865 57076 7909
rect 57180 7865 57236 7909
rect 57340 7865 57396 7909
rect 57500 7865 57556 7909
rect 57660 7865 57716 7909
rect 57820 7865 57876 7909
rect 57980 7865 58036 7909
rect 58140 7865 58196 7909
rect 58300 7865 58356 7909
rect 58460 7865 58516 7909
rect 58620 7865 58676 7909
rect 58780 7865 58836 7909
rect 58940 7865 58996 7909
rect 59100 7865 59156 7909
rect 59260 7865 59316 7909
rect 59420 7865 59476 7909
rect 59708 7865 59764 7909
rect 63692 11809 63764 11822
rect 63692 11763 63705 11809
rect 63751 11763 63764 11809
rect 63692 11750 63764 11763
rect 63852 11809 63924 11822
rect 63852 11763 63865 11809
rect 63911 11763 63924 11809
rect 63852 11750 63924 11763
rect 62292 11689 62348 11733
rect 62580 11689 62636 11733
rect 62740 11689 62796 11733
rect 62900 11689 62956 11733
rect 63060 11689 63116 11733
rect 63220 11689 63276 11733
rect 63380 11689 63436 11733
rect 63540 11689 63596 11733
rect 63700 11689 63756 11750
rect 63860 11689 63916 11750
rect 64020 11689 64076 11733
rect 64180 11689 64236 11733
rect 64340 11689 64396 11733
rect 64500 11689 64556 11733
rect 64660 11689 64716 11733
rect 64820 11689 64876 11733
rect 64980 11689 65036 11733
rect 65268 11689 65324 11733
rect 62292 10895 62348 11089
rect 62284 10882 62356 10895
rect 62284 10836 62297 10882
rect 62343 10836 62356 10882
rect 62284 10823 62356 10836
rect 62292 10629 62348 10823
rect 62580 10762 62636 11089
rect 62740 10762 62796 11089
rect 62900 10762 62956 11089
rect 63060 10762 63116 11089
rect 63220 10762 63276 11089
rect 63380 10762 63436 11089
rect 63540 10762 63596 11089
rect 63700 10762 63756 11089
rect 63860 10762 63916 11089
rect 64020 10762 64076 11089
rect 64180 10762 64236 11089
rect 64340 10762 64396 11089
rect 64500 10762 64556 11089
rect 64660 10762 64716 11089
rect 64820 10762 64876 11089
rect 64980 10762 65036 11089
rect 65268 10895 65324 11089
rect 65260 10882 65332 10895
rect 65260 10836 65273 10882
rect 65319 10836 65332 10882
rect 65260 10823 65332 10836
rect 62580 10749 65036 10762
rect 62580 10703 63705 10749
rect 63751 10703 63865 10749
rect 63911 10703 65036 10749
rect 62580 10690 65036 10703
rect 62580 10629 62636 10690
rect 62740 10629 62796 10690
rect 62900 10629 62956 10690
rect 63060 10629 63116 10690
rect 63220 10629 63276 10690
rect 63380 10629 63436 10690
rect 63540 10629 63596 10690
rect 63700 10629 63756 10690
rect 63860 10629 63916 10690
rect 64020 10629 64076 10690
rect 64180 10629 64236 10690
rect 64340 10629 64396 10690
rect 64500 10629 64556 10690
rect 64660 10629 64716 10690
rect 64820 10629 64876 10690
rect 64980 10629 65036 10690
rect 65268 10629 65324 10823
rect 62292 9569 62348 10029
rect 62580 9702 62636 10029
rect 62740 9702 62796 10029
rect 62900 9702 62956 10029
rect 63060 9702 63116 10029
rect 63220 9702 63276 10029
rect 63380 9702 63436 10029
rect 63540 9702 63596 10029
rect 63700 9702 63756 10029
rect 63860 9702 63916 10029
rect 64020 9702 64076 10029
rect 64180 9702 64236 10029
rect 64340 9702 64396 10029
rect 64500 9702 64556 10029
rect 64660 9702 64716 10029
rect 64820 9702 64876 10029
rect 64980 9702 65036 10029
rect 62580 9689 65036 9702
rect 62580 9643 63705 9689
rect 63751 9643 63865 9689
rect 63911 9643 65036 9689
rect 62580 9630 65036 9643
rect 62580 9569 62636 9630
rect 62740 9569 62796 9630
rect 62900 9569 62956 9630
rect 63060 9569 63116 9630
rect 63220 9569 63276 9630
rect 63380 9569 63436 9630
rect 63540 9569 63596 9630
rect 63700 9569 63756 9630
rect 63860 9569 63916 9630
rect 64020 9569 64076 9630
rect 64180 9569 64236 9630
rect 64340 9569 64396 9630
rect 64500 9569 64556 9630
rect 64660 9569 64716 9630
rect 64820 9569 64876 9630
rect 64980 9569 65036 9630
rect 65268 9569 65324 10029
rect 62292 8775 62348 8969
rect 62284 8762 62356 8775
rect 62284 8716 62297 8762
rect 62343 8716 62356 8762
rect 62284 8703 62356 8716
rect 62292 8509 62348 8703
rect 62580 8642 62636 8969
rect 62740 8642 62796 8969
rect 62900 8642 62956 8969
rect 63060 8642 63116 8969
rect 63220 8642 63276 8969
rect 63380 8642 63436 8969
rect 63540 8642 63596 8969
rect 63700 8642 63756 8969
rect 63860 8642 63916 8969
rect 64020 8642 64076 8969
rect 64180 8642 64236 8969
rect 64340 8642 64396 8969
rect 64500 8642 64556 8969
rect 64660 8642 64716 8969
rect 64820 8642 64876 8969
rect 64980 8642 65036 8969
rect 65268 8775 65324 8969
rect 65260 8762 65332 8775
rect 65260 8716 65273 8762
rect 65319 8716 65332 8762
rect 65260 8703 65332 8716
rect 62580 8629 65036 8642
rect 62580 8583 63705 8629
rect 63751 8583 63865 8629
rect 63911 8583 65036 8629
rect 62580 8570 65036 8583
rect 62580 8509 62636 8570
rect 62740 8509 62796 8570
rect 62900 8509 62956 8570
rect 63060 8509 63116 8570
rect 63220 8509 63276 8570
rect 63380 8509 63436 8570
rect 63540 8509 63596 8570
rect 63700 8509 63756 8570
rect 63860 8509 63916 8570
rect 64020 8509 64076 8570
rect 64180 8509 64236 8570
rect 64340 8509 64396 8570
rect 64500 8509 64556 8570
rect 64660 8509 64716 8570
rect 64820 8509 64876 8570
rect 64980 8509 65036 8570
rect 65268 8509 65324 8703
rect 62292 7865 62348 7909
rect 62580 7865 62636 7909
rect 62740 7865 62796 7909
rect 62900 7865 62956 7909
rect 63060 7865 63116 7909
rect 63220 7865 63276 7909
rect 63380 7865 63436 7909
rect 63540 7865 63596 7909
rect 63700 7865 63756 7909
rect 63860 7865 63916 7909
rect 64020 7865 64076 7909
rect 64180 7865 64236 7909
rect 64340 7865 64396 7909
rect 64500 7865 64556 7909
rect 64660 7865 64716 7909
rect 64820 7865 64876 7909
rect 64980 7865 65036 7909
rect 65268 7865 65324 7909
rect 7751 5934 7823 5948
rect 7751 5888 7764 5934
rect 7810 5888 7823 5934
rect 7751 5876 7823 5888
rect 8231 5939 8303 5948
rect 8711 5939 8783 5948
rect 8231 5934 8783 5939
rect 8231 5888 8244 5934
rect 8290 5888 8724 5934
rect 8770 5888 8783 5934
rect 8231 5883 8783 5888
rect 8231 5876 8303 5883
rect 7471 5738 7527 5782
rect 7759 5738 7815 5876
rect 7919 5738 7975 5782
rect 8079 5738 8135 5782
rect 8239 5738 8295 5876
rect 8399 5738 8455 5883
rect 8559 5738 8615 5883
rect 8711 5876 8783 5883
rect 9191 5935 9263 5948
rect 9191 5889 9204 5935
rect 9250 5889 9263 5935
rect 9191 5876 9263 5889
rect 8719 5738 8775 5876
rect 8879 5738 8935 5782
rect 9039 5738 9095 5782
rect 9199 5738 9255 5876
rect 9487 5738 9543 5782
rect 7471 5202 7527 5538
rect 7759 5494 7815 5538
rect 7919 5504 7975 5538
rect 8079 5504 8135 5538
rect 7919 5448 8135 5504
rect 8239 5494 8295 5538
rect 8399 5494 8455 5538
rect 8559 5494 8615 5538
rect 8719 5494 8775 5538
rect 8879 5504 8935 5538
rect 9039 5504 9095 5538
rect 8879 5448 9095 5504
rect 9199 5494 9255 5538
rect 7919 5397 7975 5448
rect 8879 5397 8935 5448
rect 7751 5384 7823 5397
rect 7751 5338 7764 5384
rect 7810 5338 7823 5384
rect 7751 5325 7823 5338
rect 7911 5384 7983 5397
rect 7911 5338 7924 5384
rect 7970 5338 7983 5384
rect 7911 5325 7983 5338
rect 8231 5389 8303 5397
rect 8711 5389 8783 5397
rect 8231 5384 8783 5389
rect 8231 5338 8244 5384
rect 8290 5338 8724 5384
rect 8770 5338 8783 5384
rect 8231 5333 8783 5338
rect 8231 5325 8303 5333
rect 7759 5202 7815 5325
rect 7919 5202 7975 5246
rect 8079 5202 8135 5246
rect 8239 5202 8295 5325
rect 8399 5202 8455 5333
rect 8559 5202 8615 5333
rect 8711 5325 8783 5333
rect 8871 5384 8943 5397
rect 8871 5338 8884 5384
rect 8930 5338 8943 5384
rect 8871 5325 8943 5338
rect 9191 5384 9263 5397
rect 9191 5338 9204 5384
rect 9250 5338 9263 5384
rect 9191 5325 9263 5338
rect 8719 5202 8775 5325
rect 8879 5202 8935 5246
rect 9039 5202 9095 5246
rect 9199 5202 9255 5325
rect 9487 5202 9543 5538
rect 1941 4553 4213 4586
rect 1645 4515 1717 4528
rect 1365 4434 1421 4478
rect 1645 4469 1658 4515
rect 1704 4469 1717 4515
rect 1645 4456 1717 4469
rect 1941 4507 2190 4553
rect 2236 4507 2294 4553
rect 2340 4507 4213 4553
rect 1941 4474 4213 4507
rect 1653 4434 1709 4456
rect 1941 4434 2053 4474
rect 2157 4434 2269 4474
rect 2373 4434 2485 4474
rect 2589 4434 2701 4474
rect 2805 4434 2917 4474
rect 3021 4434 3133 4474
rect 3237 4434 3349 4474
rect 3453 4434 3565 4474
rect 3669 4434 3781 4474
rect 3885 4434 3997 4474
rect 4101 4434 4213 4474
rect 4309 4513 4381 4526
rect 4309 4467 4322 4513
rect 4368 4467 4381 4513
rect 4309 4454 4381 4467
rect 4469 4513 4541 4526
rect 4469 4467 4482 4513
rect 4528 4467 4541 4513
rect 4469 4454 4541 4467
rect 4317 4434 4373 4454
rect 4477 4434 4533 4454
rect 1365 3268 1421 3634
rect 1653 3590 1709 3634
rect 1941 3590 2053 3634
rect 2157 3590 2269 3634
rect 2373 3590 2485 3634
rect 2589 3590 2701 3634
rect 2805 3590 2917 3634
rect 3021 3590 3133 3634
rect 3237 3590 3349 3634
rect 3453 3590 3565 3634
rect 1949 3341 2925 3374
rect 1949 3295 2102 3341
rect 2148 3295 2206 3341
rect 2252 3295 2310 3341
rect 2356 3295 2414 3341
rect 2460 3295 2518 3341
rect 2564 3295 2622 3341
rect 2668 3295 2925 3341
rect 1357 3255 1429 3268
rect 1357 3209 1370 3255
rect 1416 3209 1429 3255
rect 1357 3196 1429 3209
rect 1653 3255 1725 3268
rect 1653 3209 1666 3255
rect 1712 3209 1725 3255
rect 1653 3196 1725 3209
rect 1949 3262 2925 3295
rect 1365 3174 1421 3196
rect 1661 3174 1717 3196
rect 1949 3174 2061 3262
rect 2165 3174 2277 3262
rect 2381 3174 2493 3262
rect 2597 3174 2709 3262
rect 2813 3174 2925 3262
rect 3029 3174 3085 3218
rect 3189 3174 3245 3218
rect 3349 3174 3405 3218
rect 3509 3174 3565 3218
rect 3669 3174 3781 3634
rect 3885 3590 3997 3634
rect 4101 3590 4213 3634
rect 4317 3590 4373 3634
rect 4477 3590 4533 3634
rect 4221 3264 4293 3277
rect 4221 3218 4234 3264
rect 4280 3218 4293 3264
rect 4013 3174 4125 3218
rect 4221 3205 4293 3218
rect 4517 3264 4589 3277
rect 4517 3218 4530 3264
rect 4576 3218 4589 3264
rect 4517 3205 4589 3218
rect 4229 3174 4285 3205
rect 4525 3174 4581 3205
rect 7471 4666 7527 5002
rect 7759 4958 7815 5002
rect 7919 4980 7975 5002
rect 8079 4980 8135 5002
rect 7919 4924 8135 4980
rect 8239 4958 8295 5002
rect 8399 4958 8455 5002
rect 8559 4958 8615 5002
rect 8719 4958 8775 5002
rect 8879 4980 8935 5002
rect 9039 4980 9095 5002
rect 8879 4924 9095 4980
rect 9199 4958 9255 5002
rect 7919 4876 7975 4924
rect 8879 4876 8935 4924
rect 7751 4863 7823 4876
rect 7751 4817 7764 4863
rect 7810 4817 7823 4863
rect 7751 4804 7823 4817
rect 7911 4863 7983 4876
rect 7911 4817 7924 4863
rect 7970 4817 7983 4863
rect 7911 4804 7983 4817
rect 8231 4868 8303 4876
rect 8711 4868 8783 4876
rect 8231 4863 8783 4868
rect 8231 4817 8244 4863
rect 8290 4817 8724 4863
rect 8770 4817 8783 4863
rect 8231 4812 8455 4817
rect 8231 4804 8303 4812
rect 7759 4666 7815 4804
rect 7919 4666 7975 4710
rect 8079 4666 8135 4710
rect 8239 4666 8295 4804
rect 8399 4666 8455 4812
rect 8559 4666 8615 4817
rect 8711 4804 8783 4817
rect 8871 4863 8943 4876
rect 8871 4817 8884 4863
rect 8930 4817 8943 4863
rect 8871 4804 8943 4817
rect 9191 4863 9263 4876
rect 9191 4817 9204 4863
rect 9250 4817 9263 4863
rect 9191 4804 9263 4817
rect 8719 4666 8775 4804
rect 8879 4666 8935 4710
rect 9039 4666 9095 4710
rect 9199 4666 9255 4804
rect 9487 4666 9543 5002
rect 19030 4915 21486 4928
rect 19030 4869 20662 4915
rect 20708 4869 20766 4915
rect 20812 4869 21355 4915
rect 21401 4869 21486 4915
rect 19030 4856 21486 4869
rect 18870 4779 18926 4823
rect 19030 4779 19086 4856
rect 19190 4779 19246 4856
rect 19350 4779 19406 4856
rect 19510 4779 19566 4856
rect 19670 4779 19726 4856
rect 19830 4779 19886 4856
rect 19990 4779 20046 4856
rect 20150 4779 20206 4856
rect 20310 4779 20366 4856
rect 20470 4779 20526 4856
rect 20630 4779 20686 4856
rect 20790 4779 20846 4856
rect 20950 4779 21006 4856
rect 21110 4779 21166 4856
rect 21270 4779 21326 4856
rect 21430 4779 21486 4856
rect 21590 4779 21646 4823
rect 21750 4779 21806 4823
rect 22038 4779 22094 4823
rect 22326 4779 22382 4823
rect 7471 4130 7527 4466
rect 7759 4422 7815 4466
rect 7919 4446 7975 4466
rect 8079 4446 8135 4466
rect 7919 4390 8135 4446
rect 8239 4422 8295 4466
rect 8399 4422 8455 4466
rect 8559 4422 8615 4466
rect 8719 4422 8775 4466
rect 8879 4446 8935 4466
rect 9039 4446 9095 4466
rect 8879 4390 9095 4446
rect 9199 4422 9255 4466
rect 7919 4342 7975 4390
rect 8879 4342 8935 4390
rect 7751 4329 7823 4342
rect 7751 4283 7764 4329
rect 7810 4283 7823 4329
rect 7751 4270 7823 4283
rect 7911 4329 7983 4342
rect 7911 4283 7924 4329
rect 7970 4283 7983 4329
rect 7911 4270 7983 4283
rect 8231 4334 8303 4342
rect 8711 4334 8783 4342
rect 8231 4329 8783 4334
rect 8231 4283 8244 4329
rect 8290 4283 8724 4329
rect 8770 4283 8783 4329
rect 8231 4270 8303 4283
rect 7759 4130 7815 4270
rect 7919 4130 7975 4174
rect 8079 4130 8135 4174
rect 8239 4130 8295 4270
rect 8399 4130 8455 4283
rect 8559 4130 8615 4283
rect 8711 4270 8783 4283
rect 8871 4329 8943 4342
rect 8871 4283 8884 4329
rect 8930 4283 8943 4329
rect 8871 4270 8943 4283
rect 9191 4329 9263 4342
rect 9191 4283 9204 4329
rect 9250 4283 9263 4329
rect 9191 4270 9263 4283
rect 8719 4130 8775 4270
rect 8879 4130 8935 4174
rect 9039 4130 9095 4174
rect 9199 4130 9255 4270
rect 9487 4130 9543 4466
rect 7471 3798 7527 3930
rect 7759 3886 7815 3930
rect 7919 3910 7975 3930
rect 8079 3910 8135 3930
rect 7919 3854 8135 3910
rect 8239 3886 8295 3930
rect 8399 3886 8455 3930
rect 8559 3886 8615 3930
rect 8719 3886 8775 3930
rect 8879 3910 8935 3930
rect 9039 3910 9095 3930
rect 8879 3854 9095 3910
rect 9199 3886 9255 3930
rect 7919 3806 7975 3854
rect 8879 3806 8935 3854
rect 7463 3785 7535 3798
rect 7463 3739 7476 3785
rect 7522 3739 7535 3785
rect 7463 3726 7535 3739
rect 7751 3793 7823 3806
rect 7751 3747 7764 3793
rect 7810 3747 7823 3793
rect 7751 3734 7823 3747
rect 7911 3793 7983 3806
rect 7911 3747 7924 3793
rect 7970 3747 7983 3793
rect 7911 3734 7983 3747
rect 8231 3798 8303 3806
rect 8711 3798 8783 3806
rect 8231 3793 8783 3798
rect 8231 3747 8244 3793
rect 8290 3747 8724 3793
rect 8770 3747 8783 3793
rect 8231 3734 8303 3747
rect 7471 3594 7527 3726
rect 7759 3594 7815 3734
rect 7919 3594 7975 3638
rect 8079 3594 8135 3638
rect 8239 3594 8295 3734
rect 8399 3594 8455 3747
rect 8559 3594 8615 3747
rect 8711 3734 8783 3747
rect 8871 3793 8943 3806
rect 8871 3747 8884 3793
rect 8930 3747 8943 3793
rect 8871 3734 8943 3747
rect 9191 3791 9263 3804
rect 9487 3798 9543 3930
rect 9191 3745 9204 3791
rect 9250 3745 9263 3791
rect 8719 3594 8775 3734
rect 9191 3732 9263 3745
rect 9478 3785 9551 3798
rect 9478 3739 9492 3785
rect 9538 3739 9551 3785
rect 8879 3594 8935 3638
rect 9039 3594 9095 3638
rect 9199 3594 9255 3732
rect 9478 3726 9551 3739
rect 9487 3594 9543 3726
rect 7471 3058 7527 3394
rect 7759 3350 7815 3394
rect 7919 3374 7975 3394
rect 8079 3374 8135 3394
rect 7919 3318 8135 3374
rect 8239 3350 8295 3394
rect 8399 3350 8455 3394
rect 8559 3350 8615 3394
rect 8719 3350 8775 3394
rect 8879 3374 8935 3394
rect 9039 3374 9095 3394
rect 8879 3318 9095 3374
rect 9199 3350 9255 3394
rect 7919 3270 7975 3318
rect 8879 3270 8935 3318
rect 7751 3257 7823 3270
rect 7751 3211 7764 3257
rect 7810 3211 7823 3257
rect 7751 3198 7823 3211
rect 7911 3257 7983 3270
rect 7911 3211 7924 3257
rect 7970 3211 7983 3257
rect 7911 3198 7983 3211
rect 8231 3262 8303 3270
rect 8711 3262 8783 3270
rect 8231 3257 8783 3262
rect 8231 3211 8244 3257
rect 8290 3211 8724 3257
rect 8770 3211 8783 3257
rect 8231 3198 8303 3211
rect 7759 3058 7815 3198
rect 7919 3058 7975 3102
rect 8079 3058 8135 3102
rect 8239 3058 8295 3198
rect 8399 3058 8455 3211
rect 8559 3058 8615 3211
rect 8711 3198 8783 3211
rect 8871 3257 8943 3270
rect 8871 3211 8884 3257
rect 8930 3211 8943 3257
rect 8871 3198 8943 3211
rect 9191 3255 9263 3268
rect 9191 3209 9204 3255
rect 9250 3209 9263 3255
rect 8719 3058 8775 3198
rect 9191 3196 9263 3209
rect 8879 3058 8935 3102
rect 9039 3058 9095 3102
rect 9199 3058 9255 3196
rect 9487 3058 9543 3394
rect 1365 1914 1421 2374
rect 1661 2330 1717 2374
rect 1949 2330 2061 2374
rect 2165 2330 2277 2374
rect 2381 2330 2493 2374
rect 2597 2330 2709 2374
rect 2813 2330 2925 2374
rect 3029 2352 3085 2374
rect 3189 2352 3245 2374
rect 3029 2339 3245 2352
rect 3029 2293 3114 2339
rect 3160 2293 3245 2339
rect 3029 2288 3245 2293
rect 3349 2352 3405 2374
rect 3509 2352 3565 2374
rect 3349 2339 3565 2352
rect 3349 2293 3434 2339
rect 3480 2293 3565 2339
rect 3349 2288 3565 2293
rect 3669 2354 3781 2374
rect 4013 2354 4125 2374
rect 3669 2341 4125 2354
rect 3669 2295 3702 2341
rect 3748 2295 4125 2341
rect 4229 2330 4285 2374
rect 3101 2280 3173 2288
rect 3421 2280 3493 2288
rect 3669 2262 4125 2295
rect 1661 1914 1717 1958
rect 1821 1914 1877 1958
rect 1981 1914 2037 1958
rect 2141 1914 2197 1958
rect 2301 1914 2357 1958
rect 2461 1914 2517 1958
rect 2621 1914 2677 1958
rect 2781 1914 2837 1958
rect 2941 1914 2997 1958
rect 3101 1914 3157 1958
rect 3261 1914 3317 1958
rect 3421 1914 3477 1958
rect 3581 1914 3637 1958
rect 3741 1914 3797 1958
rect 3901 1914 3957 1958
rect 4061 1914 4117 1958
rect 4221 1914 4421 1958
rect 4525 1914 4581 2374
rect 1365 1770 1421 1814
rect 1661 1775 1717 1814
rect 1821 1783 1877 1814
rect 1981 1783 2037 1814
rect 1813 1775 1885 1783
rect 1973 1775 2045 1783
rect 2141 1775 2197 1814
rect 2301 1775 2357 1814
rect 2461 1783 2517 1814
rect 2453 1775 2525 1783
rect 2621 1775 2677 1814
rect 2781 1775 2837 1814
rect 2941 1775 2997 1814
rect 3101 1783 3157 1814
rect 3093 1775 3165 1783
rect 3261 1775 3317 1814
rect 3421 1775 3477 1814
rect 3581 1775 3637 1814
rect 3741 1775 3797 1814
rect 3901 1775 3957 1814
rect 4061 1775 4117 1814
rect 4221 1775 4421 1814
rect 1661 1770 4421 1775
rect 4525 1770 4581 1814
rect 1661 1724 1826 1770
rect 1872 1724 1986 1770
rect 2032 1724 2466 1770
rect 2512 1724 3106 1770
rect 3152 1724 4421 1770
rect 1661 1719 4421 1724
rect 1813 1711 1885 1719
rect 1973 1711 2045 1719
rect 2453 1711 2525 1719
rect 3093 1711 3165 1719
rect 7471 2814 7527 2858
rect 7759 2814 7815 2858
rect 7919 2838 7975 2858
rect 8079 2838 8135 2858
rect 7919 2782 8135 2838
rect 8239 2814 8295 2858
rect 8399 2814 8455 2858
rect 8559 2814 8615 2858
rect 8719 2814 8775 2858
rect 8879 2838 8935 2858
rect 9039 2838 9095 2858
rect 8879 2782 9095 2838
rect 9199 2814 9255 2858
rect 9487 2814 9543 2858
rect 13190 4001 13390 4081
rect 13190 3955 13220 4001
rect 13266 3955 13314 4001
rect 13360 3955 13390 4001
rect 13190 3907 13390 3955
rect 13190 3861 13220 3907
rect 13266 3861 13314 3907
rect 13360 3861 13390 3907
rect 12758 3781 12958 3825
rect 13190 3781 13390 3861
rect 13494 3781 13694 3825
rect 13798 3781 13998 3825
rect 14102 3781 14302 3825
rect 14406 3781 14606 3825
rect 14710 3781 14910 3825
rect 15142 3781 15342 3825
rect 15446 3781 15646 3825
rect 15750 3781 15950 3825
rect 16054 3781 16254 3825
rect 16358 3781 16558 3825
rect 16662 3781 16862 3825
rect 12758 3245 12958 3381
rect 13190 3245 13390 3381
rect 13494 3245 13694 3381
rect 13798 3245 13998 3381
rect 14102 3245 14302 3381
rect 14406 3245 14606 3381
rect 14710 3245 14910 3381
rect 15142 3245 15342 3381
rect 15446 3245 15646 3381
rect 15750 3245 15950 3381
rect 16054 3245 16254 3381
rect 16358 3245 16558 3381
rect 16662 3245 16862 3381
rect 7919 2734 7975 2782
rect 8879 2734 8935 2782
rect 7911 2721 7983 2734
rect 7911 2675 7924 2721
rect 7970 2675 7983 2721
rect 7911 2662 7983 2675
rect 8871 2721 8943 2734
rect 8871 2675 8884 2721
rect 8930 2675 8943 2721
rect 8871 2662 8943 2675
rect 9520 2633 10632 2649
rect 9520 2587 10328 2633
rect 10374 2587 10432 2633
rect 10478 2587 10632 2633
rect 6664 2524 6736 2532
rect 6824 2524 6896 2532
rect 7144 2524 7216 2532
rect 7304 2524 7376 2532
rect 7464 2524 7536 2532
rect 7624 2524 7696 2532
rect 7784 2524 7856 2532
rect 7944 2524 8016 2532
rect 8104 2524 8176 2532
rect 8264 2524 8336 2532
rect 8424 2524 8496 2532
rect 8584 2524 8656 2532
rect 8744 2524 8816 2532
rect 8904 2524 8976 2532
rect 9064 2524 9136 2532
rect 9224 2524 9296 2532
rect 6512 2519 7048 2524
rect 6512 2473 6677 2519
rect 6723 2473 6837 2519
rect 6883 2473 7048 2519
rect 6224 2429 6280 2473
rect 6512 2468 7048 2473
rect 6512 2429 6568 2468
rect 6664 2460 6736 2468
rect 6824 2460 6896 2468
rect 6672 2429 6728 2460
rect 6832 2429 6888 2460
rect 6992 2429 7048 2468
rect 7144 2519 9296 2524
rect 7144 2473 7157 2519
rect 7203 2473 7317 2519
rect 7363 2473 7477 2519
rect 7523 2473 7637 2519
rect 7683 2473 7797 2519
rect 7843 2473 7957 2519
rect 8003 2473 8117 2519
rect 8163 2473 8277 2519
rect 8323 2473 8437 2519
rect 8483 2473 8597 2519
rect 8643 2473 8757 2519
rect 8803 2473 8917 2519
rect 8963 2473 9077 2519
rect 9123 2473 9237 2519
rect 9283 2473 9296 2519
rect 7144 2468 9296 2473
rect 7144 2460 7216 2468
rect 7304 2460 7376 2468
rect 7464 2460 7536 2468
rect 7624 2460 7696 2468
rect 7784 2460 7856 2468
rect 7944 2460 8016 2468
rect 8104 2460 8176 2468
rect 8264 2460 8336 2468
rect 8424 2460 8496 2468
rect 8584 2460 8656 2468
rect 8744 2460 8816 2468
rect 8904 2460 8976 2468
rect 9064 2460 9136 2468
rect 9224 2460 9296 2468
rect 9520 2529 10632 2587
rect 9520 2483 10328 2529
rect 10374 2483 10432 2529
rect 10478 2483 10632 2529
rect 7152 2429 7208 2460
rect 7312 2429 7368 2460
rect 7472 2429 7528 2460
rect 7632 2429 7688 2460
rect 7792 2429 7848 2460
rect 7952 2429 8008 2460
rect 8112 2429 8168 2460
rect 8272 2429 8328 2460
rect 8432 2429 8488 2460
rect 8592 2429 8648 2460
rect 8752 2429 8808 2460
rect 8912 2429 8968 2460
rect 9072 2429 9128 2460
rect 9232 2429 9288 2460
rect 9520 2449 10632 2483
rect 9520 2429 9720 2449
rect 9824 2429 10024 2449
rect 10128 2429 10328 2449
rect 10432 2429 10632 2449
rect 10736 2429 10792 2473
rect 6224 2046 6280 2229
rect 6512 2185 6568 2229
rect 6672 2185 6728 2229
rect 6832 2185 6888 2229
rect 6992 2185 7048 2229
rect 7152 2185 7208 2229
rect 7312 2185 7368 2229
rect 7472 2185 7528 2229
rect 7632 2185 7688 2229
rect 7792 2185 7848 2229
rect 7952 2185 8008 2229
rect 8112 2185 8168 2229
rect 8272 2185 8328 2229
rect 8432 2185 8488 2229
rect 8592 2185 8648 2229
rect 8752 2185 8808 2229
rect 8912 2185 8968 2229
rect 9072 2185 9128 2229
rect 9232 2185 9288 2229
rect 9520 2185 9720 2229
rect 9824 2185 10024 2229
rect 10128 2185 10328 2229
rect 10432 2185 10632 2229
rect 10736 2046 10792 2229
rect 6216 2033 6288 2046
rect 6216 1987 6229 2033
rect 6275 1987 6288 2033
rect 6216 1974 6288 1987
rect 10728 2033 10800 2046
rect 10728 1987 10741 2033
rect 10787 1987 10800 2033
rect 10728 1974 10800 1987
rect 6224 1792 6280 1974
rect 6512 1907 8352 1924
rect 6512 1861 6527 1907
rect 6573 1861 6631 1907
rect 6677 1891 8352 1907
rect 6677 1861 8071 1891
rect 6512 1845 8071 1861
rect 8117 1845 8165 1891
rect 8211 1845 8259 1891
rect 8305 1845 8352 1891
rect 6512 1812 8352 1845
rect 6512 1792 6624 1812
rect 6728 1792 6840 1812
rect 6944 1792 7056 1812
rect 7160 1792 7272 1812
rect 7376 1792 7488 1812
rect 7592 1792 7704 1812
rect 7808 1792 7920 1812
rect 8024 1792 8136 1812
rect 8240 1792 8352 1812
rect 8456 1882 9688 1924
rect 8456 1836 8757 1882
rect 8803 1836 8917 1882
rect 8963 1836 9077 1882
rect 9123 1836 9237 1882
rect 9283 1836 9397 1882
rect 9443 1836 9557 1882
rect 9603 1836 9688 1882
rect 10736 1868 10792 1974
rect 8456 1812 9688 1836
rect 8456 1792 8568 1812
rect 8672 1792 8728 1812
rect 8832 1792 8888 1812
rect 8992 1792 9048 1812
rect 9152 1792 9208 1812
rect 9312 1792 9368 1812
rect 9472 1792 9528 1812
rect 9632 1792 9688 1812
rect 9936 1812 10792 1868
rect 9936 1792 9992 1812
rect 10096 1792 10152 1812
rect 10256 1792 10312 1812
rect 10416 1792 10472 1812
rect 10576 1792 10632 1812
rect 10736 1792 10792 1812
rect 6224 1548 6280 1592
rect 6512 1548 6624 1592
rect 6728 1548 6840 1592
rect 6944 1548 7056 1592
rect 7160 1548 7272 1592
rect 7376 1548 7488 1592
rect 7592 1548 7704 1592
rect 7808 1548 7920 1592
rect 8024 1548 8136 1592
rect 8240 1548 8352 1592
rect 8456 1548 8568 1592
rect 8672 1548 8728 1592
rect 8832 1548 8888 1592
rect 8992 1548 9048 1592
rect 9152 1548 9208 1592
rect 9312 1548 9368 1592
rect 9472 1548 9528 1592
rect 9632 1548 9688 1592
rect 9936 1548 9992 1592
rect 10096 1548 10152 1592
rect 10256 1548 10312 1592
rect 10416 1548 10472 1592
rect 10576 1548 10632 1592
rect 10736 1548 10792 1592
rect 12758 2697 12958 2845
rect 13190 2801 13390 2845
rect 12758 2651 12788 2697
rect 12834 2651 12882 2697
rect 12928 2651 12958 2697
rect 12758 2603 12958 2651
rect 12758 2557 12788 2603
rect 12834 2557 12882 2603
rect 12928 2557 12958 2603
rect 13494 2785 13694 2845
rect 13798 2785 13998 2845
rect 14102 2785 14302 2845
rect 14406 2785 14606 2845
rect 14710 2785 14910 2845
rect 15142 2785 15342 2845
rect 15446 2785 15646 2845
rect 15750 2785 15950 2845
rect 16054 2785 16254 2845
rect 16358 2785 16558 2845
rect 13494 2760 16558 2785
rect 13494 2714 16186 2760
rect 16232 2714 16290 2760
rect 16336 2714 16394 2760
rect 16440 2714 16558 2760
rect 13494 2708 16558 2714
rect 13494 2662 13629 2708
rect 13675 2662 13723 2708
rect 13769 2662 13817 2708
rect 13863 2662 14237 2708
rect 14283 2662 14331 2708
rect 14377 2662 14425 2708
rect 14471 2662 14845 2708
rect 14891 2662 14939 2708
rect 14985 2662 15033 2708
rect 15079 2662 16558 2708
rect 13494 2656 16558 2662
rect 13494 2610 16186 2656
rect 16232 2610 16290 2656
rect 16336 2610 16394 2656
rect 16440 2610 16558 2656
rect 13494 2585 16558 2610
rect 16662 2697 16862 2845
rect 16662 2651 16692 2697
rect 16738 2651 16786 2697
rect 16832 2651 16862 2697
rect 16662 2603 16862 2651
rect 12758 2409 12958 2557
rect 16662 2557 16692 2603
rect 16738 2557 16786 2603
rect 16832 2557 16862 2603
rect 13190 2409 13390 2453
rect 13494 2409 13694 2453
rect 13798 2409 13998 2453
rect 14102 2409 14302 2453
rect 14406 2409 14606 2453
rect 14710 2409 14910 2453
rect 15142 2409 15342 2453
rect 15446 2409 15646 2453
rect 15750 2409 15950 2453
rect 16054 2409 16254 2453
rect 16358 2409 16558 2453
rect 16662 2409 16862 2557
rect 12758 1965 12958 2009
rect 13190 1812 13390 2009
rect 13190 1766 13215 1812
rect 13261 1766 13319 1812
rect 13365 1766 13390 1812
rect 13190 1708 13390 1766
rect 13494 1909 13694 2009
rect 13798 1909 13998 2009
rect 14102 1909 14302 2009
rect 14406 1909 14606 2009
rect 14710 1909 14910 2009
rect 15142 1909 15342 2009
rect 15446 1909 15646 2009
rect 15750 1909 15950 2009
rect 16054 1909 16254 2009
rect 16358 1909 16558 2009
rect 16662 1965 16862 2009
rect 13494 1832 16558 1909
rect 13494 1786 13629 1832
rect 13675 1786 13723 1832
rect 13769 1786 13817 1832
rect 13863 1786 14227 1832
rect 14273 1786 14331 1832
rect 14377 1786 14435 1832
rect 14481 1786 14845 1832
rect 14891 1786 14939 1832
rect 14985 1786 15033 1832
rect 15079 1786 16558 1832
rect 13494 1709 16558 1786
rect 13190 1662 13215 1708
rect 13261 1662 13319 1708
rect 13365 1662 13390 1708
rect 13190 1637 13390 1662
rect 18870 4147 18926 4179
rect 18862 4134 18934 4147
rect 18862 4088 18875 4134
rect 18921 4088 18934 4134
rect 18862 4075 18934 4088
rect 18870 4043 18926 4075
rect 19030 4043 19086 4179
rect 19190 4043 19246 4179
rect 19350 4043 19406 4179
rect 19510 4043 19566 4179
rect 19670 4043 19726 4179
rect 19830 4043 19886 4179
rect 19990 4043 20046 4179
rect 20150 4043 20206 4179
rect 20310 4043 20366 4179
rect 20470 4043 20526 4179
rect 20630 4043 20686 4179
rect 20790 4043 20846 4179
rect 20950 4043 21006 4179
rect 21110 4043 21166 4179
rect 21270 4043 21326 4179
rect 21430 4043 21486 4179
rect 21590 4043 21646 4179
rect 21750 4043 21806 4179
rect 22038 4147 22094 4179
rect 22326 4147 22382 4179
rect 22030 4134 22102 4147
rect 22030 4088 22043 4134
rect 22089 4088 22102 4134
rect 22030 4075 22102 4088
rect 22318 4134 22390 4147
rect 22318 4088 22331 4134
rect 22377 4088 22390 4134
rect 22318 4075 22390 4088
rect 22038 4043 22094 4075
rect 22326 4043 22382 4075
rect 23660 4906 23860 4919
rect 23660 4860 23673 4906
rect 23847 4860 23860 4906
rect 23660 4817 23860 4860
rect 23660 3774 23860 3817
rect 23660 3728 23673 3774
rect 23847 3728 23860 3774
rect 23660 3715 23860 3728
rect 24108 4906 24308 4919
rect 24108 4860 24121 4906
rect 24295 4860 24308 4906
rect 24108 4817 24308 4860
rect 24108 3774 24308 3817
rect 24108 3728 24121 3774
rect 24295 3728 24308 3774
rect 24108 3715 24308 3728
rect 24556 4906 24756 4919
rect 24556 4860 24569 4906
rect 24743 4860 24756 4906
rect 24556 4817 24756 4860
rect 24556 3774 24756 3817
rect 24556 3728 24569 3774
rect 24743 3728 24756 3774
rect 24556 3715 24756 3728
rect 24836 4906 25036 4919
rect 24836 4860 24849 4906
rect 25023 4860 25036 4906
rect 24836 4817 25036 4860
rect 24836 3774 25036 3817
rect 24836 3728 24849 3774
rect 25023 3728 25036 3774
rect 24836 3715 25036 3728
rect 25284 4906 25484 4919
rect 25284 4860 25297 4906
rect 25471 4860 25484 4906
rect 25284 4817 25484 4860
rect 25284 3774 25484 3817
rect 25284 3728 25297 3774
rect 25471 3728 25484 3774
rect 25284 3715 25484 3728
rect 25564 4906 25764 4919
rect 25564 4860 25577 4906
rect 25751 4860 25764 4906
rect 25564 4817 25764 4860
rect 25564 3774 25764 3817
rect 25564 3728 25577 3774
rect 25751 3728 25764 3774
rect 25564 3715 25764 3728
rect 26012 4906 26212 4919
rect 26012 4860 26025 4906
rect 26199 4860 26212 4906
rect 26012 4817 26212 4860
rect 26012 3774 26212 3817
rect 26012 3728 26025 3774
rect 26199 3728 26212 3774
rect 26012 3715 26212 3728
rect 26292 4906 26492 4919
rect 26292 4860 26305 4906
rect 26479 4860 26492 4906
rect 26292 4817 26492 4860
rect 26292 3774 26492 3817
rect 26292 3728 26305 3774
rect 26479 3728 26492 3774
rect 26292 3715 26492 3728
rect 26740 4906 26940 4919
rect 26740 4860 26753 4906
rect 26927 4860 26940 4906
rect 26740 4817 26940 4860
rect 26740 3774 26940 3817
rect 26740 3728 26753 3774
rect 26927 3728 26940 3774
rect 26740 3715 26940 3728
rect 27020 4906 27220 4919
rect 27020 4860 27033 4906
rect 27207 4860 27220 4906
rect 27020 4817 27220 4860
rect 27020 3774 27220 3817
rect 27020 3728 27033 3774
rect 27207 3728 27220 3774
rect 27020 3715 27220 3728
rect 27468 4906 27668 4919
rect 27468 4860 27481 4906
rect 27655 4860 27668 4906
rect 27468 4817 27668 4860
rect 27468 3774 27668 3817
rect 27468 3728 27481 3774
rect 27655 3728 27668 3774
rect 27468 3715 27668 3728
rect 27940 4906 28140 4919
rect 27940 4860 27953 4906
rect 28127 4860 28140 4906
rect 27940 4817 28140 4860
rect 27940 3774 28140 3817
rect 27940 3728 27953 3774
rect 28127 3728 28140 3774
rect 27940 3715 28140 3728
rect 18870 3307 18926 3443
rect 19030 3307 19086 3443
rect 19190 3307 19246 3443
rect 19350 3307 19406 3443
rect 19510 3307 19566 3443
rect 19670 3307 19726 3443
rect 19830 3307 19886 3443
rect 19990 3307 20046 3443
rect 20150 3307 20206 3443
rect 20310 3307 20366 3443
rect 20470 3307 20526 3443
rect 20630 3307 20686 3443
rect 20790 3307 20846 3443
rect 20950 3307 21006 3443
rect 21110 3307 21166 3443
rect 21270 3307 21326 3443
rect 21430 3307 21486 3443
rect 21590 3307 21646 3443
rect 21750 3307 21806 3443
rect 22038 3399 22094 3443
rect 22326 3307 22382 3443
rect 22038 3207 22094 3251
rect 29286 5090 29486 5103
rect 29286 5044 29299 5090
rect 29473 5044 29486 5090
rect 29286 5001 29486 5044
rect 29286 3718 29486 3761
rect 29286 3672 29299 3718
rect 29473 3672 29486 3718
rect 29286 3659 29486 3672
rect 29734 5090 29934 5103
rect 29734 5044 29747 5090
rect 29921 5044 29934 5090
rect 29734 5001 29934 5044
rect 29734 3718 29934 3761
rect 29734 3672 29747 3718
rect 29921 3672 29934 3718
rect 29734 3659 29934 3672
rect 30014 5090 30214 5103
rect 30014 5044 30027 5090
rect 30201 5044 30214 5090
rect 30014 5001 30214 5044
rect 30014 3718 30214 3761
rect 30014 3672 30027 3718
rect 30201 3672 30214 3718
rect 30014 3659 30214 3672
rect 30294 5090 30494 5103
rect 30294 5044 30307 5090
rect 30481 5044 30494 5090
rect 30294 5001 30494 5044
rect 30294 3718 30494 3761
rect 30294 3672 30307 3718
rect 30481 3672 30494 3718
rect 30294 3659 30494 3672
rect 30574 5090 30774 5103
rect 30574 5044 30587 5090
rect 30761 5044 30774 5090
rect 30574 5001 30774 5044
rect 30574 3718 30774 3761
rect 30574 3672 30587 3718
rect 30761 3672 30774 3718
rect 30574 3659 30774 3672
rect 31022 5090 31222 5103
rect 31022 5044 31035 5090
rect 31209 5044 31222 5090
rect 31022 5001 31222 5044
rect 31022 3718 31222 3761
rect 31022 3672 31035 3718
rect 31209 3672 31222 3718
rect 31022 3659 31222 3672
rect 18870 2675 18926 2707
rect 18862 2662 18934 2675
rect 18862 2616 18875 2662
rect 18921 2616 18934 2662
rect 18862 2603 18934 2616
rect 18870 2571 18926 2603
rect 19030 2571 19086 2707
rect 19190 2571 19246 2707
rect 19350 2571 19406 2707
rect 19510 2571 19566 2707
rect 19670 2571 19726 2707
rect 19830 2571 19886 2707
rect 19990 2571 20046 2707
rect 20150 2571 20206 2707
rect 20310 2571 20366 2707
rect 20470 2571 20526 2707
rect 20630 2571 20686 2707
rect 20790 2571 20846 2707
rect 20950 2571 21006 2707
rect 21110 2571 21166 2707
rect 21270 2571 21326 2707
rect 21430 2571 21486 2707
rect 21590 2571 21646 2707
rect 21750 2571 21806 2707
rect 22038 2471 22094 2707
rect 22326 2675 22382 2707
rect 22318 2662 22390 2675
rect 22318 2616 22331 2662
rect 22377 2616 22390 2662
rect 22318 2603 22390 2616
rect 22326 2571 22382 2603
rect 18870 1927 18926 1971
rect 19030 1927 19086 1971
rect 19190 1927 19246 1971
rect 19350 1927 19406 1971
rect 19510 1927 19566 1971
rect 19670 1927 19726 1971
rect 19830 1927 19886 1971
rect 19990 1927 20046 1971
rect 20150 1927 20206 1971
rect 20310 1927 20366 1971
rect 20470 1927 20526 1971
rect 20630 1927 20686 1971
rect 20790 1927 20846 1971
rect 20950 1927 21006 1971
rect 21110 1927 21166 1971
rect 21270 1927 21326 1971
rect 21430 1927 21486 1971
rect 21590 1914 21646 1971
rect 21750 1914 21806 1971
rect 22038 1914 22094 1971
rect 22326 1927 22382 1971
rect 21590 1901 22094 1914
rect 21590 1855 21646 1901
rect 21692 1855 21750 1901
rect 21796 1855 21854 1901
rect 21900 1855 21963 1901
rect 22009 1855 22094 1901
rect 21590 1842 22094 1855
rect 23660 2934 23860 2947
rect 23660 2888 23673 2934
rect 23847 2888 23860 2934
rect 23660 2845 23860 2888
rect 23660 1802 23860 1845
rect 23660 1756 23673 1802
rect 23847 1756 23860 1802
rect 23660 1743 23860 1756
rect 24108 2934 24308 2947
rect 24108 2888 24121 2934
rect 24295 2888 24308 2934
rect 24108 2845 24308 2888
rect 24108 1802 24308 1845
rect 24108 1756 24121 1802
rect 24295 1756 24308 1802
rect 24108 1743 24308 1756
rect 24556 2934 24756 2947
rect 24556 2888 24569 2934
rect 24743 2888 24756 2934
rect 24556 2845 24756 2888
rect 24556 1802 24756 1845
rect 24556 1756 24569 1802
rect 24743 1756 24756 1802
rect 24556 1743 24756 1756
rect 24836 2934 25036 2947
rect 24836 2888 24849 2934
rect 25023 2888 25036 2934
rect 24836 2845 25036 2888
rect 24836 1802 25036 1845
rect 24836 1756 24849 1802
rect 25023 1756 25036 1802
rect 24836 1743 25036 1756
rect 25284 2934 25484 2947
rect 25284 2888 25297 2934
rect 25471 2888 25484 2934
rect 25284 2845 25484 2888
rect 25284 1802 25484 1845
rect 25284 1756 25297 1802
rect 25471 1756 25484 1802
rect 25284 1743 25484 1756
rect 25564 2934 25764 2947
rect 25564 2888 25577 2934
rect 25751 2888 25764 2934
rect 25564 2845 25764 2888
rect 25564 1802 25764 1845
rect 25564 1756 25577 1802
rect 25751 1756 25764 1802
rect 25564 1743 25764 1756
rect 26012 2934 26212 2947
rect 26012 2888 26025 2934
rect 26199 2888 26212 2934
rect 26012 2845 26212 2888
rect 26012 1802 26212 1845
rect 26012 1756 26025 1802
rect 26199 1756 26212 1802
rect 26012 1743 26212 1756
rect 26292 2934 26492 2947
rect 26292 2888 26305 2934
rect 26479 2888 26492 2934
rect 26292 2845 26492 2888
rect 26292 1802 26492 1845
rect 26292 1756 26305 1802
rect 26479 1756 26492 1802
rect 26292 1743 26492 1756
rect 26740 2934 26940 2947
rect 26740 2888 26753 2934
rect 26927 2888 26940 2934
rect 26740 2845 26940 2888
rect 26740 1802 26940 1845
rect 26740 1756 26753 1802
rect 26927 1756 26940 1802
rect 26740 1743 26940 1756
rect 27020 2934 27220 2947
rect 27020 2888 27033 2934
rect 27207 2888 27220 2934
rect 27020 2845 27220 2888
rect 27020 1802 27220 1845
rect 27020 1756 27033 1802
rect 27207 1756 27220 1802
rect 27020 1743 27220 1756
rect 27468 2934 27668 2947
rect 27468 2888 27481 2934
rect 27655 2888 27668 2934
rect 27468 2845 27668 2888
rect 27468 1802 27668 1845
rect 27468 1756 27481 1802
rect 27655 1756 27668 1802
rect 27468 1743 27668 1756
rect 27940 2934 28140 2947
rect 27940 2888 27953 2934
rect 28127 2888 28140 2934
rect 27940 2845 28140 2888
rect 27940 1802 28140 1845
rect 27940 1756 27953 1802
rect 28127 1756 28140 1802
rect 27940 1743 28140 1756
rect 29286 3078 29486 3091
rect 29286 3032 29299 3078
rect 29473 3032 29486 3078
rect 29286 2989 29486 3032
rect 29286 1706 29486 1749
rect 29286 1660 29299 1706
rect 29473 1660 29486 1706
rect 29286 1647 29486 1660
rect 29734 3078 29934 3091
rect 29734 3032 29747 3078
rect 29921 3032 29934 3078
rect 29734 2989 29934 3032
rect 29734 1706 29934 1749
rect 29734 1660 29747 1706
rect 29921 1660 29934 1706
rect 29734 1647 29934 1660
rect 30014 3078 30214 3091
rect 30014 3032 30027 3078
rect 30201 3032 30214 3078
rect 30014 2989 30214 3032
rect 30014 1706 30214 1749
rect 30014 1660 30027 1706
rect 30201 1660 30214 1706
rect 30014 1647 30214 1660
rect 30294 3078 30494 3091
rect 30294 3032 30307 3078
rect 30481 3032 30494 3078
rect 30294 2989 30494 3032
rect 30294 1706 30494 1749
rect 30294 1660 30307 1706
rect 30481 1660 30494 1706
rect 30294 1647 30494 1660
rect 30574 3078 30774 3091
rect 30574 3032 30587 3078
rect 30761 3032 30774 3078
rect 30574 2989 30774 3032
rect 30574 1706 30774 1749
rect 30574 1660 30587 1706
rect 30761 1660 30774 1706
rect 30574 1647 30774 1660
rect 31022 3078 31222 3091
rect 31022 3032 31035 3078
rect 31209 3032 31222 3078
rect 31022 2989 31222 3032
rect 31022 1706 31222 1749
rect 31022 1660 31035 1706
rect 31209 1660 31222 1706
rect 31022 1647 31222 1660
<< polycontact >>
rect 3965 14173 4011 14219
rect 4445 14173 4491 14219
rect 5085 14173 5131 14219
rect 3965 13045 4011 13091
rect 4125 13045 4171 13091
rect 4445 13045 4491 13091
rect 4765 13045 4811 13091
rect 5085 13045 5131 13091
rect 3965 11917 4011 11963
rect 4125 11917 4171 11963
rect 4445 11917 4491 11963
rect 4765 11917 4811 11963
rect 5085 11917 5131 11963
rect -7373 10310 -7199 10356
rect -7373 9718 -7199 9764
rect -7093 10310 -6919 10356
rect -7093 9718 -6919 9764
rect -6813 10310 -6639 10356
rect -6813 9718 -6639 9764
rect -6533 10310 -6359 10356
rect -6533 9718 -6359 9764
rect -6253 10310 -6079 10356
rect -6253 9718 -6079 9764
rect -5973 10310 -5799 10356
rect -5973 9718 -5799 9764
rect -5693 10310 -5519 10356
rect -5693 9718 -5519 9764
rect -5413 10310 -5239 10356
rect -5413 9718 -5239 9764
rect -5133 10310 -4959 10356
rect -5133 9718 -4959 9764
rect -4853 10310 -4679 10356
rect -4853 9718 -4679 9764
rect -4573 10310 -4399 10356
rect -4573 9718 -4399 9764
rect -4293 10310 -4119 10356
rect -4293 9718 -4119 9764
rect -7373 9393 -7199 9439
rect -7373 8801 -7199 8847
rect -7093 9393 -6919 9439
rect -7093 8801 -6919 8847
rect -6813 9393 -6639 9439
rect -6813 8801 -6639 8847
rect -6533 9393 -6359 9439
rect -6533 8801 -6359 8847
rect -6253 9393 -6079 9439
rect -6253 8801 -6079 8847
rect -5973 9393 -5799 9439
rect -5973 8801 -5799 8847
rect -5693 9393 -5519 9439
rect -5693 8801 -5519 8847
rect -5413 9393 -5239 9439
rect -5413 8801 -5239 8847
rect -5133 9393 -4959 9439
rect -5133 8801 -4959 8847
rect -4853 9393 -4679 9439
rect -4853 8801 -4679 8847
rect -4573 9393 -4399 9439
rect -4573 8801 -4399 8847
rect -4293 9393 -4119 9439
rect -4293 8801 -4119 8847
rect -7373 8476 -7199 8522
rect -7373 7884 -7199 7930
rect -7093 8476 -6919 8522
rect -7093 7884 -6919 7930
rect -6813 8476 -6639 8522
rect -6813 7884 -6639 7930
rect -6533 8476 -6359 8522
rect -6533 7884 -6359 7930
rect -6253 8476 -6079 8522
rect -6253 7884 -6079 7930
rect -5973 8476 -5799 8522
rect -5973 7884 -5799 7930
rect -5693 8476 -5519 8522
rect -5693 7884 -5519 7930
rect -5413 8476 -5239 8522
rect -5413 7884 -5239 7930
rect -5133 8476 -4959 8522
rect -5133 7884 -4959 7930
rect -4853 8476 -4679 8522
rect -4853 7884 -4679 7930
rect -4573 8476 -4399 8522
rect -4573 7884 -4399 7930
rect -4293 8476 -4119 8522
rect -4293 7884 -4119 7930
rect 3965 9657 4011 9703
rect 4125 9657 4171 9703
rect 4445 9657 4491 9703
rect 4765 9657 4811 9703
rect 5085 9657 5131 9703
rect 3677 8543 3723 8589
rect 1019 8317 1065 8363
rect 2963 8317 3009 8363
rect 3965 8527 4011 8573
rect 4125 8527 4171 8573
rect 4445 8527 4491 8573
rect 4765 8527 4811 8573
rect 5085 8527 5131 8573
rect 5373 8543 5419 8589
rect 1242 7534 1288 7580
rect 1346 7534 1392 7580
rect -7373 7062 -7199 7108
rect -7373 6470 -7199 6516
rect -7093 7062 -6919 7108
rect -7093 6470 -6919 6516
rect -6813 7062 -6639 7108
rect -6813 6470 -6639 6516
rect -6533 7062 -6359 7108
rect -6533 6470 -6359 6516
rect -6253 7062 -6079 7108
rect -6253 6470 -6079 6516
rect -5973 7062 -5799 7108
rect -5973 6470 -5799 6516
rect -5693 7062 -5519 7108
rect -5693 6470 -5519 6516
rect -5413 7062 -5239 7108
rect -5413 6470 -5239 6516
rect -5133 7062 -4959 7108
rect -5133 6470 -4959 6516
rect -4853 7062 -4679 7108
rect -4853 6470 -4679 6516
rect -4573 7062 -4399 7108
rect -4573 6470 -4399 6516
rect -4293 7062 -4119 7108
rect -4293 6470 -4119 6516
rect -7373 6145 -7199 6191
rect -7373 5553 -7199 5599
rect -7093 6145 -6919 6191
rect -7093 5553 -6919 5599
rect -6813 6145 -6639 6191
rect -6813 5553 -6639 5599
rect -6533 6145 -6359 6191
rect -6533 5553 -6359 5599
rect -6253 6145 -6079 6191
rect -6253 5553 -6079 5599
rect -5973 6145 -5799 6191
rect -5973 5553 -5799 5599
rect -5693 6145 -5519 6191
rect -5693 5553 -5519 5599
rect -5413 6145 -5239 6191
rect -5413 5553 -5239 5599
rect -5133 6145 -4959 6191
rect -5133 5553 -4959 5599
rect -4853 6145 -4679 6191
rect -4853 5553 -4679 5599
rect -4573 6145 -4399 6191
rect -4573 5553 -4399 5599
rect -4293 6145 -4119 6191
rect -4293 5553 -4119 5599
rect -7373 5228 -7199 5274
rect -7373 4636 -7199 4682
rect -7093 5228 -6919 5274
rect -7093 4636 -6919 4682
rect -6813 5228 -6639 5274
rect -6813 4636 -6639 4682
rect -6533 5228 -6359 5274
rect -6533 4636 -6359 4682
rect -6253 5228 -6079 5274
rect -6253 4636 -6079 4682
rect -5973 5228 -5799 5274
rect -5973 4636 -5799 4682
rect -5693 5228 -5519 5274
rect -5693 4636 -5519 4682
rect -5413 5228 -5239 5274
rect -5413 4636 -5239 4682
rect -5133 5228 -4959 5274
rect -5133 4636 -4959 4682
rect -4853 5228 -4679 5274
rect -4853 4636 -4679 4682
rect -4573 5228 -4399 5274
rect -4573 4636 -4399 4682
rect -4293 5228 -4119 5274
rect -4293 4636 -4119 4682
rect 4125 7443 4171 7489
rect 4765 7443 4811 7489
rect 19080 13356 19126 13402
rect 19560 13356 19606 13402
rect 20200 13356 20246 13402
rect 18792 12398 18838 12444
rect 19080 12390 19126 12436
rect 19240 12390 19286 12436
rect 19560 12390 19606 12436
rect 19880 12390 19926 12436
rect 20200 12390 20246 12436
rect 20488 12398 20534 12444
rect 6542 8362 6588 8408
rect 8004 8415 8050 8461
rect 8004 8311 8050 8357
rect 8238 8362 8284 8408
rect 10737 8404 10783 8450
rect 8777 8343 8823 8389
rect 10737 8300 10783 8346
rect 10985 8343 11031 8389
rect 12403 8514 12449 8560
rect 12159 8389 12205 8435
rect 12403 8410 12449 8456
rect 14367 8389 14413 8435
rect 15189 8519 15235 8565
rect 14953 8389 14999 8435
rect 15189 8415 15235 8461
rect 16649 8389 16695 8435
rect 19080 11454 19126 11500
rect 19240 11454 19286 11500
rect 19560 11454 19606 11500
rect 19880 11454 19926 11500
rect 20200 11454 20246 11500
rect 19080 9582 19126 9628
rect 19240 9582 19286 9628
rect 19560 9582 19606 9628
rect 19880 9582 19926 9628
rect 20200 9582 20246 9628
rect 18792 8654 18838 8700
rect 19080 8646 19126 8692
rect 19240 8646 19286 8692
rect 19560 8646 19606 8692
rect 19880 8646 19926 8692
rect 20200 8646 20246 8692
rect 20488 8654 20534 8700
rect 19240 7710 19286 7756
rect 19880 7710 19926 7756
rect 24232 13356 24278 13402
rect 24872 13356 24918 13402
rect 25352 13356 25398 13402
rect 23944 12398 23990 12444
rect 24232 12390 24278 12436
rect 24552 12390 24598 12436
rect 24872 12390 24918 12436
rect 25192 12390 25238 12436
rect 25352 12390 25398 12436
rect 25640 12398 25686 12444
rect 24232 11454 24278 11500
rect 24552 11454 24598 11500
rect 24872 11454 24918 11500
rect 25192 11454 25238 11500
rect 25352 11454 25398 11500
rect 24232 9582 24278 9628
rect 24552 9582 24598 9628
rect 24872 9582 24918 9628
rect 25192 9582 25238 9628
rect 25352 9582 25398 9628
rect 23944 8654 23990 8700
rect 24232 8646 24278 8692
rect 24552 8646 24598 8692
rect 24872 8646 24918 8692
rect 25192 8646 25238 8692
rect 25352 8646 25398 8692
rect 25640 8654 25686 8700
rect 24552 7710 24598 7756
rect 25192 7710 25238 7756
rect 28201 13356 28247 13402
rect 28681 13356 28727 13402
rect 29321 13356 29367 13402
rect 27913 12398 27959 12444
rect 28201 12390 28247 12436
rect 28361 12390 28407 12436
rect 28681 12390 28727 12436
rect 29001 12390 29047 12436
rect 29321 12390 29367 12436
rect 29609 12398 29655 12444
rect 28201 11454 28247 11500
rect 28361 11454 28407 11500
rect 28681 11454 28727 11500
rect 29001 11454 29047 11500
rect 29321 11454 29367 11500
rect 28201 9582 28247 9628
rect 28361 9582 28407 9628
rect 28681 9582 28727 9628
rect 29001 9582 29047 9628
rect 29321 9582 29367 9628
rect 27913 8654 27959 8700
rect 28201 8646 28247 8692
rect 28361 8646 28407 8692
rect 28681 8646 28727 8692
rect 29001 8646 29047 8692
rect 29321 8646 29367 8692
rect 29609 8654 29655 8700
rect 28361 7710 28407 7756
rect 29001 7710 29047 7756
rect 34617 11763 34663 11809
rect 34777 11763 34823 11809
rect 38753 11763 38799 11809
rect 38913 11763 38959 11809
rect 33209 10836 33255 10882
rect 36185 10836 36231 10882
rect 34617 10703 34663 10749
rect 34777 10703 34823 10749
rect 37345 10836 37391 10882
rect 40321 10836 40367 10882
rect 38753 10703 38799 10749
rect 38913 10703 38959 10749
rect 34617 9643 34663 9689
rect 34777 9643 34823 9689
rect 38753 9643 38799 9689
rect 38913 9643 38959 9689
rect 33209 8716 33255 8762
rect 36185 8716 36231 8762
rect 34617 8583 34663 8629
rect 34777 8583 34823 8629
rect 37345 8716 37391 8762
rect 40321 8716 40367 8762
rect 38753 8583 38799 8629
rect 38913 8583 38959 8629
rect 44313 11763 44359 11809
rect 44473 11763 44519 11809
rect 48449 11763 48495 11809
rect 48609 11763 48655 11809
rect 42905 10836 42951 10882
rect 45881 10836 45927 10882
rect 44313 10703 44359 10749
rect 44473 10703 44519 10749
rect 47041 10836 47087 10882
rect 50017 10836 50063 10882
rect 48449 10703 48495 10749
rect 48609 10703 48655 10749
rect 44313 9643 44359 9689
rect 44473 9643 44519 9689
rect 48449 9643 48495 9689
rect 48609 9643 48655 9689
rect 42905 8716 42951 8762
rect 45881 8716 45927 8762
rect 44313 8583 44359 8629
rect 44473 8583 44519 8629
rect 47041 8716 47087 8762
rect 50017 8716 50063 8762
rect 48449 8583 48495 8629
rect 48609 8583 48655 8629
rect 54009 11763 54055 11809
rect 54169 11763 54215 11809
rect 58145 11763 58191 11809
rect 58305 11763 58351 11809
rect 52601 10836 52647 10882
rect 55577 10836 55623 10882
rect 54009 10703 54055 10749
rect 54169 10703 54215 10749
rect 56737 10836 56783 10882
rect 59713 10836 59759 10882
rect 58145 10703 58191 10749
rect 58305 10703 58351 10749
rect 54009 9643 54055 9689
rect 54169 9643 54215 9689
rect 58145 9643 58191 9689
rect 58305 9643 58351 9689
rect 52601 8716 52647 8762
rect 55577 8716 55623 8762
rect 54009 8583 54055 8629
rect 54169 8583 54215 8629
rect 56737 8716 56783 8762
rect 59713 8716 59759 8762
rect 58145 8583 58191 8629
rect 58305 8583 58351 8629
rect 63705 11763 63751 11809
rect 63865 11763 63911 11809
rect 62297 10836 62343 10882
rect 65273 10836 65319 10882
rect 63705 10703 63751 10749
rect 63865 10703 63911 10749
rect 63705 9643 63751 9689
rect 63865 9643 63911 9689
rect 62297 8716 62343 8762
rect 65273 8716 65319 8762
rect 63705 8583 63751 8629
rect 63865 8583 63911 8629
rect 7764 5888 7810 5934
rect 8244 5888 8290 5934
rect 8724 5888 8770 5934
rect 9204 5889 9250 5935
rect 7764 5338 7810 5384
rect 7924 5338 7970 5384
rect 8244 5338 8290 5384
rect 8724 5338 8770 5384
rect 8884 5338 8930 5384
rect 9204 5338 9250 5384
rect 1658 4469 1704 4515
rect 2190 4507 2236 4553
rect 2294 4507 2340 4553
rect 4322 4467 4368 4513
rect 4482 4467 4528 4513
rect 2102 3295 2148 3341
rect 2206 3295 2252 3341
rect 2310 3295 2356 3341
rect 2414 3295 2460 3341
rect 2518 3295 2564 3341
rect 2622 3295 2668 3341
rect 1370 3209 1416 3255
rect 1666 3209 1712 3255
rect 4234 3218 4280 3264
rect 4530 3218 4576 3264
rect 7764 4817 7810 4863
rect 7924 4817 7970 4863
rect 8244 4817 8290 4863
rect 8724 4817 8770 4863
rect 8884 4817 8930 4863
rect 9204 4817 9250 4863
rect 20662 4869 20708 4915
rect 20766 4869 20812 4915
rect 21355 4869 21401 4915
rect 7764 4283 7810 4329
rect 7924 4283 7970 4329
rect 8244 4283 8290 4329
rect 8724 4283 8770 4329
rect 8884 4283 8930 4329
rect 9204 4283 9250 4329
rect 7476 3739 7522 3785
rect 7764 3747 7810 3793
rect 7924 3747 7970 3793
rect 8244 3747 8290 3793
rect 8724 3747 8770 3793
rect 8884 3747 8930 3793
rect 9204 3745 9250 3791
rect 9492 3739 9538 3785
rect 7764 3211 7810 3257
rect 7924 3211 7970 3257
rect 8244 3211 8290 3257
rect 8724 3211 8770 3257
rect 8884 3211 8930 3257
rect 9204 3209 9250 3255
rect 3114 2293 3160 2339
rect 3434 2293 3480 2339
rect 3702 2295 3748 2341
rect 1826 1724 1872 1770
rect 1986 1724 2032 1770
rect 2466 1724 2512 1770
rect 3106 1724 3152 1770
rect 13220 3955 13266 4001
rect 13314 3955 13360 4001
rect 13220 3861 13266 3907
rect 13314 3861 13360 3907
rect 7924 2675 7970 2721
rect 8884 2675 8930 2721
rect 10328 2587 10374 2633
rect 10432 2587 10478 2633
rect 6677 2473 6723 2519
rect 6837 2473 6883 2519
rect 7157 2473 7203 2519
rect 7317 2473 7363 2519
rect 7477 2473 7523 2519
rect 7637 2473 7683 2519
rect 7797 2473 7843 2519
rect 7957 2473 8003 2519
rect 8117 2473 8163 2519
rect 8277 2473 8323 2519
rect 8437 2473 8483 2519
rect 8597 2473 8643 2519
rect 8757 2473 8803 2519
rect 8917 2473 8963 2519
rect 9077 2473 9123 2519
rect 9237 2473 9283 2519
rect 10328 2483 10374 2529
rect 10432 2483 10478 2529
rect 6229 1987 6275 2033
rect 10741 1987 10787 2033
rect 6527 1861 6573 1907
rect 6631 1861 6677 1907
rect 8071 1845 8117 1891
rect 8165 1845 8211 1891
rect 8259 1845 8305 1891
rect 8757 1836 8803 1882
rect 8917 1836 8963 1882
rect 9077 1836 9123 1882
rect 9237 1836 9283 1882
rect 9397 1836 9443 1882
rect 9557 1836 9603 1882
rect 12788 2651 12834 2697
rect 12882 2651 12928 2697
rect 12788 2557 12834 2603
rect 12882 2557 12928 2603
rect 16186 2714 16232 2760
rect 16290 2714 16336 2760
rect 16394 2714 16440 2760
rect 13629 2662 13675 2708
rect 13723 2662 13769 2708
rect 13817 2662 13863 2708
rect 14237 2662 14283 2708
rect 14331 2662 14377 2708
rect 14425 2662 14471 2708
rect 14845 2662 14891 2708
rect 14939 2662 14985 2708
rect 15033 2662 15079 2708
rect 16186 2610 16232 2656
rect 16290 2610 16336 2656
rect 16394 2610 16440 2656
rect 16692 2651 16738 2697
rect 16786 2651 16832 2697
rect 16692 2557 16738 2603
rect 16786 2557 16832 2603
rect 13215 1766 13261 1812
rect 13319 1766 13365 1812
rect 13629 1786 13675 1832
rect 13723 1786 13769 1832
rect 13817 1786 13863 1832
rect 14227 1786 14273 1832
rect 14331 1786 14377 1832
rect 14435 1786 14481 1832
rect 14845 1786 14891 1832
rect 14939 1786 14985 1832
rect 15033 1786 15079 1832
rect 13215 1662 13261 1708
rect 13319 1662 13365 1708
rect 18875 4088 18921 4134
rect 22043 4088 22089 4134
rect 22331 4088 22377 4134
rect 23673 4860 23847 4906
rect 23673 3728 23847 3774
rect 24121 4860 24295 4906
rect 24121 3728 24295 3774
rect 24569 4860 24743 4906
rect 24569 3728 24743 3774
rect 24849 4860 25023 4906
rect 24849 3728 25023 3774
rect 25297 4860 25471 4906
rect 25297 3728 25471 3774
rect 25577 4860 25751 4906
rect 25577 3728 25751 3774
rect 26025 4860 26199 4906
rect 26025 3728 26199 3774
rect 26305 4860 26479 4906
rect 26305 3728 26479 3774
rect 26753 4860 26927 4906
rect 26753 3728 26927 3774
rect 27033 4860 27207 4906
rect 27033 3728 27207 3774
rect 27481 4860 27655 4906
rect 27481 3728 27655 3774
rect 27953 4860 28127 4906
rect 27953 3728 28127 3774
rect 29299 5044 29473 5090
rect 29299 3672 29473 3718
rect 29747 5044 29921 5090
rect 29747 3672 29921 3718
rect 30027 5044 30201 5090
rect 30027 3672 30201 3718
rect 30307 5044 30481 5090
rect 30307 3672 30481 3718
rect 30587 5044 30761 5090
rect 30587 3672 30761 3718
rect 31035 5044 31209 5090
rect 31035 3672 31209 3718
rect 18875 2616 18921 2662
rect 22331 2616 22377 2662
rect 21646 1855 21692 1901
rect 21750 1855 21796 1901
rect 21854 1855 21900 1901
rect 21963 1855 22009 1901
rect 23673 2888 23847 2934
rect 23673 1756 23847 1802
rect 24121 2888 24295 2934
rect 24121 1756 24295 1802
rect 24569 2888 24743 2934
rect 24569 1756 24743 1802
rect 24849 2888 25023 2934
rect 24849 1756 25023 1802
rect 25297 2888 25471 2934
rect 25297 1756 25471 1802
rect 25577 2888 25751 2934
rect 25577 1756 25751 1802
rect 26025 2888 26199 2934
rect 26025 1756 26199 1802
rect 26305 2888 26479 2934
rect 26305 1756 26479 1802
rect 26753 2888 26927 2934
rect 26753 1756 26927 1802
rect 27033 2888 27207 2934
rect 27033 1756 27207 1802
rect 27481 2888 27655 2934
rect 27481 1756 27655 1802
rect 27953 2888 28127 2934
rect 27953 1756 28127 1802
rect 29299 3032 29473 3078
rect 29299 1660 29473 1706
rect 29747 3032 29921 3078
rect 29747 1660 29921 1706
rect 30027 3032 30201 3078
rect 30027 1660 30201 1706
rect 30307 3032 30481 3078
rect 30307 1660 30481 1706
rect 30587 3032 30761 3078
rect 30587 1660 30761 1706
rect 31035 3032 31209 3078
rect 31035 1660 31209 1706
<< ppolyres >>
rect -7386 9807 -7186 10267
rect -7106 9807 -6906 10267
rect -6826 9807 -6626 10267
rect -6546 9807 -6346 10267
rect -6266 9807 -6066 10267
rect -5986 9807 -5786 10267
rect -5706 9807 -5506 10267
rect -5426 9807 -5226 10267
rect -5146 9807 -4946 10267
rect -4866 9807 -4666 10267
rect -4586 9807 -4386 10267
rect -4306 9807 -4106 10267
rect -7386 8890 -7186 9350
rect -7106 8890 -6906 9350
rect -6826 8890 -6626 9350
rect -6546 8890 -6346 9350
rect -6266 8890 -6066 9350
rect -5986 8890 -5786 9350
rect -5706 8890 -5506 9350
rect -5426 8890 -5226 9350
rect -5146 8890 -4946 9350
rect -4866 8890 -4666 9350
rect -4586 8890 -4386 9350
rect -4306 8890 -4106 9350
rect -7386 7973 -7186 8433
rect -7106 7973 -6906 8433
rect -6826 7973 -6626 8433
rect -6546 7973 -6346 8433
rect -6266 7973 -6066 8433
rect -5986 7973 -5786 8433
rect -5706 7973 -5506 8433
rect -5426 7973 -5226 8433
rect -5146 7973 -4946 8433
rect -4866 7973 -4666 8433
rect -4586 7973 -4386 8433
rect -4306 7973 -4106 8433
rect -7386 6559 -7186 7019
rect -7106 6559 -6906 7019
rect -6826 6559 -6626 7019
rect -6546 6559 -6346 7019
rect -6266 6559 -6066 7019
rect -5986 6559 -5786 7019
rect -5706 6559 -5506 7019
rect -5426 6559 -5226 7019
rect -5146 6559 -4946 7019
rect -4866 6559 -4666 7019
rect -4586 6559 -4386 7019
rect -4306 6559 -4106 7019
rect -7386 5642 -7186 6102
rect -7106 5642 -6906 6102
rect -6826 5642 -6626 6102
rect -6546 5642 -6346 6102
rect -6266 5642 -6066 6102
rect -5986 5642 -5786 6102
rect -5706 5642 -5506 6102
rect -5426 5642 -5226 6102
rect -5146 5642 -4946 6102
rect -4866 5642 -4666 6102
rect -4586 5642 -4386 6102
rect -4306 5642 -4106 6102
rect -7386 4725 -7186 5185
rect -7106 4725 -6906 5185
rect -6826 4725 -6626 5185
rect -6546 4725 -6346 5185
rect -6266 4725 -6066 5185
rect -5986 4725 -5786 5185
rect -5706 4725 -5506 5185
rect -5426 4725 -5226 5185
rect -5146 4725 -4946 5185
rect -4866 4725 -4666 5185
rect -4586 4725 -4386 5185
rect -4306 4725 -4106 5185
rect 23660 3817 23860 4817
rect 24108 3817 24308 4817
rect 24556 3817 24756 4817
rect 24836 3817 25036 4817
rect 25284 3817 25484 4817
rect 25564 3817 25764 4817
rect 26012 3817 26212 4817
rect 26292 3817 26492 4817
rect 26740 3817 26940 4817
rect 27020 3817 27220 4817
rect 27468 3817 27668 4817
rect 27940 3817 28140 4817
rect 29286 3761 29486 5001
rect 29734 3761 29934 5001
rect 30014 3761 30214 5001
rect 30294 3761 30494 5001
rect 30574 3761 30774 5001
rect 31022 3761 31222 5001
rect 23660 1845 23860 2845
rect 24108 1845 24308 2845
rect 24556 1845 24756 2845
rect 24836 1845 25036 2845
rect 25284 1845 25484 2845
rect 25564 1845 25764 2845
rect 26012 1845 26212 2845
rect 26292 1845 26492 2845
rect 26740 1845 26940 2845
rect 27020 1845 27220 2845
rect 27468 1845 27668 2845
rect 27940 1845 28140 2845
rect 29286 1749 29486 2989
rect 29734 1749 29934 2989
rect 30014 1749 30214 2989
rect 30294 1749 30494 2989
rect 30574 1749 30774 2989
rect 31022 1749 31222 2989
<< metal1 >>
rect 31218 15717 31505 15718
rect 31218 15705 33394 15717
rect 31218 15653 31230 15705
rect 31282 15653 31334 15705
rect 31386 15653 31438 15705
rect 31490 15653 33394 15705
rect 31218 15601 33394 15653
rect 31218 15549 31230 15601
rect 31282 15549 31334 15601
rect 31386 15549 31438 15601
rect 31490 15549 33394 15601
rect 31218 15497 33394 15549
rect 31218 15445 31230 15497
rect 31282 15445 31334 15497
rect 31386 15445 31438 15497
rect 31490 15445 33394 15497
rect 31218 15433 33394 15445
rect 31218 15420 31505 15433
rect 32132 15119 34298 15131
rect 32132 15067 32144 15119
rect 32196 15067 32248 15119
rect 32300 15067 32352 15119
rect 32404 15067 34298 15119
rect 32132 15015 34298 15067
rect 32132 14963 32144 15015
rect 32196 14963 32248 15015
rect 32300 14963 32352 15015
rect 32404 14963 34298 15015
rect 32132 14911 34298 14963
rect 32132 14859 32144 14911
rect 32196 14859 32248 14911
rect 32300 14859 32352 14911
rect 32404 14859 34298 14911
rect 32132 14847 34298 14859
rect 15658 14722 17304 14728
rect 6229 14665 30392 14722
rect 6229 14619 6262 14665
rect 6308 14619 6356 14665
rect 6402 14619 6450 14665
rect 6496 14619 6544 14665
rect 6590 14619 6638 14665
rect 6684 14619 6732 14665
rect 6778 14619 6826 14665
rect 6872 14619 6920 14665
rect 6966 14619 7014 14665
rect 7060 14619 7108 14665
rect 7154 14619 7202 14665
rect 7248 14619 7296 14665
rect 7342 14619 7390 14665
rect 7436 14619 7484 14665
rect 7530 14619 7578 14665
rect 7624 14619 7672 14665
rect 7718 14619 7766 14665
rect 7812 14619 7860 14665
rect 7906 14619 7954 14665
rect 8000 14619 8048 14665
rect 8094 14619 8142 14665
rect 8188 14619 8236 14665
rect 8282 14619 8330 14665
rect 8376 14619 8424 14665
rect 8470 14619 8518 14665
rect 8564 14619 30392 14665
rect 6229 14571 30392 14619
rect 6229 14525 6262 14571
rect 6308 14562 8518 14571
rect 6308 14525 6341 14562
rect 3411 14374 5685 14441
rect 1805 14328 2238 14334
rect 3161 14328 3341 14338
rect 1805 14326 3341 14328
rect 1805 14321 3173 14326
rect 1802 14265 1812 14321
rect 1868 14265 1922 14321
rect 1978 14265 2032 14321
rect 2088 14265 2142 14321
rect 2198 14274 3173 14321
rect 3225 14274 3277 14326
rect 3329 14274 3341 14326
rect 2198 14265 3341 14274
rect 1805 14222 3341 14265
rect 1805 14211 3173 14222
rect 1805 14155 1812 14211
rect 1868 14155 1922 14211
rect 1978 14155 2032 14211
rect 2088 14155 2142 14211
rect 2198 14170 3173 14211
rect 3225 14170 3277 14222
rect 3329 14170 3341 14222
rect 2198 14168 3341 14170
rect 2198 14155 2238 14168
rect 3161 14158 3341 14168
rect 3411 14328 3444 14374
rect 3490 14328 3538 14374
rect 3584 14328 3632 14374
rect 3678 14328 3726 14374
rect 3772 14328 3820 14374
rect 3866 14328 3914 14374
rect 3960 14328 4008 14374
rect 4054 14328 4102 14374
rect 4148 14328 4196 14374
rect 4242 14328 4290 14374
rect 4336 14328 4384 14374
rect 4430 14328 4478 14374
rect 4524 14328 4572 14374
rect 4618 14328 4666 14374
rect 4712 14328 4760 14374
rect 4806 14328 4854 14374
rect 4900 14328 4948 14374
rect 4994 14328 5042 14374
rect 5088 14328 5136 14374
rect 5182 14328 5230 14374
rect 5276 14328 5324 14374
rect 5370 14328 5418 14374
rect 5464 14328 5512 14374
rect 5558 14328 5606 14374
rect 5652 14328 5685 14374
rect 3411 14281 5685 14328
rect 5741 14284 5901 14474
rect 3411 14280 3523 14281
rect 3411 14234 3444 14280
rect 3490 14234 3523 14280
rect 3411 14186 3523 14234
rect 1805 14101 2238 14155
rect 1805 14045 1812 14101
rect 1868 14045 1922 14101
rect 1978 14045 2032 14101
rect 2088 14045 2142 14101
rect 2198 14045 2238 14101
rect 1805 14031 2238 14045
rect 3411 14140 3444 14186
rect 3490 14140 3523 14186
rect 3411 14092 3523 14140
rect 3411 14046 3444 14092
rect 3490 14046 3523 14092
rect 3411 13998 3523 14046
rect 2520 13979 2700 13989
rect 2338 13977 2700 13979
rect 2338 13925 2532 13977
rect 2584 13925 2636 13977
rect 2688 13925 2700 13977
rect 2338 13873 2700 13925
rect 2338 13821 2532 13873
rect 2584 13821 2636 13873
rect 2688 13821 2700 13873
rect 2338 13819 2700 13821
rect 2520 13809 2700 13819
rect 3411 13952 3444 13998
rect 3490 13952 3523 13998
rect 3411 13904 3523 13952
rect 3411 13858 3444 13904
rect 3490 13858 3523 13904
rect 3411 13810 3523 13858
rect 3411 13764 3444 13810
rect 3490 13764 3523 13810
rect 3411 13716 3523 13764
rect 3411 13670 3444 13716
rect 3490 13670 3523 13716
rect 3411 13622 3523 13670
rect 3411 13576 3444 13622
rect 3490 13576 3523 13622
rect 3411 13528 3523 13576
rect 3411 13482 3444 13528
rect 3490 13482 3523 13528
rect 3411 13434 3523 13482
rect 3411 13388 3444 13434
rect 3490 13388 3523 13434
rect 3411 13340 3523 13388
rect 3411 13294 3444 13340
rect 3490 13294 3523 13340
rect 3411 13246 3523 13294
rect 2881 13200 3061 13210
rect -720 13198 3061 13200
rect -720 13146 2893 13198
rect 2945 13146 2997 13198
rect 3049 13146 3061 13198
rect -720 13122 3061 13146
rect -721 13094 3061 13122
rect -721 13042 2893 13094
rect 2945 13042 2997 13094
rect 3049 13042 3061 13094
rect -721 13030 3061 13042
rect 3411 13200 3444 13246
rect 3490 13200 3523 13246
rect 3411 13152 3523 13200
rect 3411 13106 3444 13152
rect 3490 13106 3523 13152
rect 3411 13058 3523 13106
rect -721 12962 2902 13030
rect -720 12801 2902 12962
rect 3411 13012 3444 13058
rect 3490 13012 3523 13058
rect 3411 12964 3523 13012
rect 3411 12918 3444 12964
rect 3490 12918 3523 12964
rect 3411 12870 3523 12918
rect 3411 12824 3444 12870
rect 3490 12824 3523 12870
rect -7720 10648 -3809 10665
rect -7720 10602 -7703 10648
rect -7657 10602 -7605 10648
rect -7559 10602 -7507 10648
rect -7461 10602 -7409 10648
rect -7363 10602 -7311 10648
rect -7265 10602 -7213 10648
rect -7167 10602 -7115 10648
rect -7069 10602 -7017 10648
rect -6971 10602 -6919 10648
rect -6873 10602 -6821 10648
rect -6775 10602 -6723 10648
rect -6677 10602 -6625 10648
rect -6579 10602 -6527 10648
rect -6481 10602 -6429 10648
rect -6383 10602 -6331 10648
rect -6285 10602 -6233 10648
rect -6187 10602 -6135 10648
rect -6089 10602 -6037 10648
rect -5991 10602 -5939 10648
rect -5893 10602 -5841 10648
rect -5795 10602 -5743 10648
rect -5697 10602 -5645 10648
rect -5599 10602 -5547 10648
rect -5501 10602 -5449 10648
rect -5403 10602 -5351 10648
rect -5305 10602 -5253 10648
rect -5207 10602 -5155 10648
rect -5109 10602 -5057 10648
rect -5011 10602 -4959 10648
rect -4913 10602 -4861 10648
rect -4815 10602 -4763 10648
rect -4717 10602 -4665 10648
rect -4619 10602 -4567 10648
rect -4521 10602 -4469 10648
rect -4423 10602 -4371 10648
rect -4325 10602 -4273 10648
rect -4227 10602 -4175 10648
rect -4129 10602 -4077 10648
rect -4031 10602 -3979 10648
rect -3933 10602 -3872 10648
rect -3826 10602 -3809 10648
rect -7720 10585 -3809 10602
rect -7720 10540 -7640 10585
rect -7720 10494 -7703 10540
rect -7657 10494 -7640 10540
rect -7720 10442 -7640 10494
rect -3889 10540 -3809 10585
rect -3889 10494 -3872 10540
rect -3826 10494 -3809 10540
rect -7720 10396 -7703 10442
rect -7657 10396 -7640 10442
rect -7720 10363 -7640 10396
rect -6446 10402 -5886 10470
rect -7720 10356 -7188 10363
rect -6446 10356 -6359 10402
rect -5973 10356 -5886 10402
rect -5326 10402 -4766 10470
rect -5326 10356 -5239 10402
rect -4853 10356 -4766 10402
rect -3889 10442 -3809 10494
rect -3889 10396 -3872 10442
rect -3826 10396 -3809 10442
rect -3602 10427 -3416 10435
rect -3889 10363 -3809 10396
rect -3604 10371 -3594 10427
rect -3538 10371 -3484 10427
rect -3428 10371 -3416 10427
rect -4303 10356 -3809 10363
rect -7720 10344 -7373 10356
rect -7720 10298 -7703 10344
rect -7657 10310 -7373 10344
rect -7199 10310 -7188 10356
rect -7657 10298 -7188 10310
rect -7720 10295 -7188 10298
rect -7106 10310 -7093 10356
rect -6919 10310 -6906 10356
rect -7720 10246 -7640 10295
rect -7106 10289 -7089 10310
rect -7033 10289 -6979 10310
rect -6923 10289 -6906 10310
rect -7106 10283 -6906 10289
rect -6826 10310 -6813 10356
rect -6639 10310 -6626 10356
rect -6544 10310 -6533 10356
rect -6359 10310 -6348 10356
rect -6264 10310 -6253 10356
rect -6079 10310 -6068 10356
rect -5984 10310 -5973 10356
rect -5799 10310 -5788 10356
rect -5704 10310 -5693 10356
rect -5519 10310 -5508 10356
rect -5424 10310 -5413 10356
rect -5239 10310 -5228 10356
rect -5144 10310 -5133 10356
rect -4959 10310 -4948 10356
rect -4864 10310 -4853 10356
rect -4679 10310 -4668 10356
rect -4584 10310 -4573 10356
rect -4399 10310 -4388 10356
rect -4304 10310 -4293 10356
rect -4119 10344 -3809 10356
rect -4119 10310 -3872 10344
rect -6826 10289 -6809 10310
rect -6753 10289 -6699 10310
rect -6643 10289 -6626 10310
rect -6826 10283 -6626 10289
rect -7720 10200 -7703 10246
rect -7657 10200 -7640 10246
rect -7720 10148 -7640 10200
rect -6167 10264 -6080 10310
rect -5694 10264 -5607 10310
rect -6167 10196 -5607 10264
rect -5047 10264 -4960 10310
rect -4574 10264 -4487 10310
rect -4303 10298 -3872 10310
rect -3826 10298 -3809 10344
rect -4303 10295 -3809 10298
rect -5047 10196 -4487 10264
rect -3889 10246 -3809 10295
rect -3889 10200 -3872 10246
rect -3826 10200 -3809 10246
rect -7720 10102 -7703 10148
rect -7657 10102 -7640 10148
rect -7720 10050 -7640 10102
rect -7720 10004 -7703 10050
rect -7657 10004 -7640 10050
rect -7720 9952 -7640 10004
rect -7720 9906 -7703 9952
rect -7657 9906 -7640 9952
rect -7720 9854 -7640 9906
rect -3889 10148 -3809 10200
rect -3889 10102 -3872 10148
rect -3826 10102 -3809 10148
rect -3889 10050 -3809 10102
rect -3889 10004 -3872 10050
rect -3826 10004 -3809 10050
rect -3889 9952 -3809 10004
rect -3889 9906 -3872 9952
rect -3826 9906 -3809 9952
rect -3602 10369 -3416 10371
rect -720 10369 -288 12801
rect 3411 12776 3523 12824
rect 3411 12730 3444 12776
rect 3490 12730 3523 12776
rect 3411 12682 3523 12730
rect 3411 12636 3444 12682
rect 3490 12636 3523 12682
rect 3411 12588 3523 12636
rect 3411 12542 3444 12588
rect 3490 12542 3523 12588
rect 3411 12494 3523 12542
rect 3411 12448 3444 12494
rect 3490 12448 3523 12494
rect 3411 12400 3523 12448
rect 3411 12354 3444 12400
rect 3490 12354 3523 12400
rect 3411 12306 3523 12354
rect 3411 12260 3444 12306
rect 3490 12260 3523 12306
rect 3411 12212 3523 12260
rect 3411 12166 3444 12212
rect 3490 12166 3523 12212
rect 3411 12118 3523 12166
rect 3411 12072 3444 12118
rect 3490 12072 3523 12118
rect 3411 12024 3523 12072
rect 3411 11978 3444 12024
rect 3490 11978 3523 12024
rect 3411 11930 3523 11978
rect 3411 11884 3444 11930
rect 3490 11884 3523 11930
rect 3411 11836 3523 11884
rect 3411 11790 3444 11836
rect 3490 11790 3523 11836
rect 3411 11742 3523 11790
rect 3411 11696 3444 11742
rect 3490 11696 3523 11742
rect 3411 11648 3523 11696
rect 3411 11602 3444 11648
rect 3490 11602 3523 11648
rect 3411 11554 3523 11602
rect 3411 11508 3444 11554
rect 3490 11508 3523 11554
rect 3411 11460 3523 11508
rect 3411 11414 3444 11460
rect 3490 11414 3523 11460
rect 3411 11366 3523 11414
rect 3411 11320 3444 11366
rect 3490 11320 3523 11366
rect 3411 11272 3523 11320
rect 3411 11226 3444 11272
rect 3490 11226 3523 11272
rect 3411 11178 3523 11226
rect 3411 11132 3444 11178
rect 3490 11132 3523 11178
rect 3411 11084 3523 11132
rect 3411 11038 3444 11084
rect 3490 11038 3523 11084
rect 3411 10990 3523 11038
rect 3411 10953 3444 10990
rect -3602 10317 -288 10369
rect -3602 10261 -3594 10317
rect -3538 10261 -3484 10317
rect -3428 10261 -288 10317
rect -3602 10207 -288 10261
rect -3602 10151 -3594 10207
rect -3538 10151 -3484 10207
rect -3428 10151 -288 10207
rect -3602 10097 -288 10151
rect -3602 10041 -3594 10097
rect -3538 10041 -3484 10097
rect -3428 10041 -288 10097
rect -3602 9987 -288 10041
rect -3602 9931 -3594 9987
rect -3538 9931 -3484 9987
rect -3428 9931 -288 9987
rect 497 10944 3444 10953
rect 3490 10944 3523 10990
rect 497 10896 3523 10944
rect 497 10850 530 10896
rect 576 10850 624 10896
rect 670 10850 718 10896
rect 764 10850 812 10896
rect 858 10850 906 10896
rect 952 10850 1000 10896
rect 1046 10850 1094 10896
rect 1140 10850 1188 10896
rect 1234 10850 1282 10896
rect 1328 10850 1376 10896
rect 1422 10850 1470 10896
rect 1516 10850 1564 10896
rect 1610 10850 1658 10896
rect 1704 10850 1752 10896
rect 1798 10850 1846 10896
rect 1892 10850 1940 10896
rect 1986 10850 2034 10896
rect 2080 10850 2128 10896
rect 2174 10850 2222 10896
rect 2268 10850 2316 10896
rect 2362 10850 2410 10896
rect 2456 10850 2504 10896
rect 2550 10850 2598 10896
rect 2644 10850 2692 10896
rect 2738 10850 2786 10896
rect 2832 10850 2880 10896
rect 2926 10850 2974 10896
rect 3020 10850 3068 10896
rect 3114 10850 3162 10896
rect 3208 10850 3256 10896
rect 3302 10850 3350 10896
rect 3396 10850 3444 10896
rect 3490 10850 3523 10896
rect 497 10802 3523 10850
rect 497 10756 530 10802
rect 576 10793 3444 10802
rect 576 10756 609 10793
rect 497 10708 609 10756
rect 497 10662 530 10708
rect 576 10662 609 10708
rect 497 10614 609 10662
rect 497 10568 530 10614
rect 576 10568 609 10614
rect 497 10520 609 10568
rect 497 10474 530 10520
rect 576 10474 609 10520
rect 497 10426 609 10474
rect 497 10380 530 10426
rect 576 10380 609 10426
rect 497 10332 609 10380
rect 497 10286 530 10332
rect 576 10286 609 10332
rect 497 10238 609 10286
rect 497 10192 530 10238
rect 576 10192 609 10238
rect 497 10144 609 10192
rect 497 10098 530 10144
rect 576 10098 609 10144
rect 497 10050 609 10098
rect 497 10004 530 10050
rect 576 10004 609 10050
rect 497 9956 609 10004
rect -3602 9916 -3416 9931
rect -7720 9808 -7703 9854
rect -7657 9808 -7640 9854
rect -7720 9787 -7640 9808
rect -6726 9810 -6166 9878
rect -7720 9764 -7187 9787
rect -6726 9764 -6639 9810
rect -6253 9764 -6166 9810
rect -5606 9810 -5046 9878
rect -5606 9764 -5519 9810
rect -5133 9764 -5046 9810
rect -3889 9854 -3809 9906
rect -3889 9808 -3872 9854
rect -3826 9808 -3809 9854
rect -4586 9780 -4386 9791
rect -4586 9764 -4569 9780
rect -4513 9764 -4459 9780
rect -4403 9764 -4386 9780
rect -3889 9776 -3809 9808
rect -7720 9756 -7373 9764
rect -7720 9710 -7703 9756
rect -7657 9719 -7373 9756
rect -7657 9710 -7640 9719
rect -7384 9718 -7373 9719
rect -7199 9719 -7187 9764
rect -7199 9718 -7188 9719
rect -7104 9718 -7093 9764
rect -6919 9718 -6908 9764
rect -6824 9718 -6813 9764
rect -6639 9718 -6628 9764
rect -6544 9718 -6533 9764
rect -6359 9718 -6348 9764
rect -6264 9718 -6253 9764
rect -6079 9718 -6068 9764
rect -5984 9718 -5973 9764
rect -5799 9718 -5788 9764
rect -5704 9718 -5693 9764
rect -5519 9718 -5508 9764
rect -5424 9718 -5413 9764
rect -5239 9718 -5228 9764
rect -5144 9718 -5133 9764
rect -4959 9718 -4948 9764
rect -4864 9718 -4853 9764
rect -4679 9718 -4668 9764
rect -4586 9718 -4573 9764
rect -4399 9718 -4386 9764
rect -4306 9764 -3809 9776
rect -4306 9718 -4293 9764
rect -4119 9756 -3809 9764
rect -4119 9718 -3872 9756
rect -7720 9658 -7640 9710
rect -7720 9612 -7703 9658
rect -7657 9612 -7640 9658
rect -7720 9560 -7640 9612
rect -7007 9672 -6920 9718
rect -6534 9672 -6447 9718
rect -7007 9604 -6447 9672
rect -5886 9672 -5799 9718
rect -5413 9672 -5326 9718
rect -5886 9604 -5326 9672
rect -4789 9671 -4702 9718
rect -4306 9710 -3872 9718
rect -3826 9710 -3809 9756
rect -4306 9708 -3809 9710
rect -4789 9603 -4505 9671
rect -7720 9514 -7703 9560
rect -7657 9514 -7640 9560
rect -7720 9462 -7640 9514
rect -7720 9416 -7703 9462
rect -7657 9439 -7640 9462
rect -6726 9485 -6166 9553
rect -6726 9439 -6639 9485
rect -6253 9439 -6166 9485
rect -5606 9485 -5046 9553
rect -5606 9439 -5519 9485
rect -5133 9439 -5046 9485
rect -4573 9439 -4505 9603
rect -3889 9658 -3809 9708
rect -3889 9612 -3872 9658
rect -3826 9612 -3809 9658
rect -3889 9560 -3809 9612
rect -3889 9514 -3872 9560
rect -3826 9529 -3809 9560
rect 497 9910 530 9956
rect 576 9910 609 9956
rect 497 9862 609 9910
rect 497 9816 530 9862
rect 576 9816 609 9862
rect 497 9768 609 9816
rect 497 9722 530 9768
rect 576 9722 609 9768
rect 497 9674 609 9722
rect 497 9628 530 9674
rect 576 9628 609 9674
rect 497 9580 609 9628
rect 497 9534 530 9580
rect 576 9534 609 9580
rect 497 9529 609 9534
rect -3826 9514 609 9529
rect -3889 9486 609 9514
rect -3889 9462 530 9486
rect -3889 9445 -3872 9462
rect -4305 9439 -3872 9445
rect -7657 9416 -7373 9439
rect -7720 9393 -7373 9416
rect -7199 9393 -7188 9439
rect -7720 9371 -7188 9393
rect -7106 9393 -7093 9439
rect -6919 9393 -6906 9439
rect -6824 9393 -6813 9439
rect -6639 9393 -6628 9439
rect -6544 9393 -6533 9439
rect -6359 9393 -6348 9439
rect -6264 9393 -6253 9439
rect -6079 9393 -6068 9439
rect -5984 9393 -5973 9439
rect -5799 9393 -5788 9439
rect -5704 9393 -5693 9439
rect -5519 9393 -5508 9439
rect -5426 9393 -5413 9439
rect -5239 9393 -5226 9439
rect -5144 9393 -5133 9439
rect -4959 9393 -4948 9439
rect -4864 9393 -4853 9439
rect -4679 9393 -4668 9439
rect -4586 9393 -4573 9439
rect -4399 9393 -4386 9439
rect -7106 9372 -7089 9393
rect -7033 9372 -6979 9393
rect -6923 9372 -6906 9393
rect -7720 9364 -7640 9371
rect -7106 9366 -6906 9372
rect -7720 9318 -7703 9364
rect -7657 9318 -7640 9364
rect -7720 9266 -7640 9318
rect -6517 9295 -6438 9393
rect -7720 9220 -7703 9266
rect -7657 9220 -7640 9266
rect -7720 9168 -7640 9220
rect -7720 9122 -7703 9168
rect -7657 9122 -7640 9168
rect -7720 9070 -7640 9122
rect -7720 9024 -7703 9070
rect -7657 9024 -7640 9070
rect -7720 8972 -7640 9024
rect -7720 8926 -7703 8972
rect -7657 8926 -7640 8972
rect -7720 8874 -7640 8926
rect -6786 9216 -6438 9295
rect -5886 9320 -5799 9393
rect -5426 9372 -5409 9393
rect -5353 9372 -5299 9393
rect -5243 9372 -5226 9393
rect -5426 9366 -5226 9372
rect -4808 9320 -4740 9393
rect -4586 9372 -4569 9393
rect -4513 9372 -4459 9393
rect -4403 9372 -4386 9393
rect -4305 9393 -4293 9439
rect -4119 9416 -3872 9439
rect -3826 9440 530 9462
rect 576 9440 609 9486
rect -3826 9416 609 9440
rect -4119 9393 609 9416
rect -4305 9392 609 9393
rect -4305 9377 530 9392
rect -4586 9366 -4386 9372
rect -5886 9252 -4740 9320
rect -3889 9364 530 9377
rect -3889 9318 -3872 9364
rect -3826 9346 530 9364
rect 576 9346 609 9392
rect -3826 9318 609 9346
rect -3889 9298 609 9318
rect -3889 9266 530 9298
rect -3889 9220 -3872 9266
rect -3826 9252 530 9266
rect 576 9252 609 9298
rect -3826 9220 609 9252
rect -6786 8874 -6707 9216
rect -3889 9204 609 9220
rect -3889 9168 530 9204
rect -3889 9122 -3872 9168
rect -3826 9158 530 9168
rect 576 9158 609 9204
rect -3826 9122 609 9158
rect -3889 9110 609 9122
rect -3889 9079 530 9110
rect -6446 9008 -5300 9076
rect -7720 8828 -7703 8874
rect -7657 8869 -7640 8874
rect -7657 8847 -7188 8869
rect -6826 8863 -6626 8874
rect -6826 8847 -6809 8863
rect -6753 8847 -6699 8863
rect -6643 8847 -6626 8863
rect -6446 8847 -6359 9008
rect -6166 8893 -5606 8961
rect -6166 8847 -6079 8893
rect -5693 8847 -5606 8893
rect -5368 8847 -5300 9008
rect -3889 9070 -3809 9079
rect -3889 9024 -3872 9070
rect -3826 9024 -3809 9070
rect -3889 8972 -3809 9024
rect -3889 8926 -3872 8972
rect -3826 8926 -3809 8972
rect -3889 8874 -3809 8926
rect -4866 8863 -4666 8874
rect -4866 8847 -4849 8863
rect -4793 8847 -4739 8863
rect -4683 8847 -4666 8863
rect -3889 8860 -3872 8874
rect -4306 8847 -3872 8860
rect -7657 8828 -7373 8847
rect -7720 8801 -7373 8828
rect -7199 8801 -7188 8847
rect -7104 8801 -7093 8847
rect -6919 8801 -6908 8847
rect -6826 8801 -6813 8847
rect -6639 8801 -6626 8847
rect -6544 8801 -6533 8847
rect -6359 8801 -6348 8847
rect -6264 8801 -6253 8847
rect -6079 8801 -6068 8847
rect -5984 8801 -5973 8847
rect -5799 8801 -5788 8847
rect -5704 8801 -5693 8847
rect -5519 8801 -5508 8847
rect -5424 8801 -5413 8847
rect -5239 8801 -5228 8847
rect -5144 8801 -5133 8847
rect -4959 8801 -4948 8847
rect -4866 8801 -4853 8847
rect -4679 8801 -4666 8847
rect -4584 8801 -4573 8847
rect -4399 8801 -4388 8847
rect -4306 8801 -4293 8847
rect -4119 8828 -3872 8847
rect -3826 8828 -3809 8874
rect -4119 8801 -3809 8828
rect -7720 8776 -7640 8801
rect -7720 8730 -7703 8776
rect -7657 8730 -7640 8776
rect -7720 8678 -7640 8730
rect -7005 8755 -6918 8801
rect -5946 8755 -5859 8801
rect -7005 8687 -5859 8755
rect -5046 8755 -4959 8801
rect -4573 8755 -4486 8801
rect -4306 8792 -3809 8801
rect -5046 8687 -4486 8755
rect -3889 8776 -3809 8792
rect -3889 8730 -3872 8776
rect -3826 8730 -3809 8776
rect -7720 8632 -7703 8678
rect -7657 8632 -7640 8678
rect -7720 8580 -7640 8632
rect -7720 8534 -7703 8580
rect -7657 8534 -7640 8580
rect -3889 8678 -3809 8730
rect -3889 8632 -3872 8678
rect -3826 8632 -3809 8678
rect -3889 8580 -3809 8632
rect -7720 8524 -7640 8534
rect -7720 8522 -7188 8524
rect -6828 8523 -6345 8536
rect -6828 8522 -6344 8523
rect -7720 8482 -7373 8522
rect -7720 8436 -7703 8482
rect -7657 8476 -7373 8482
rect -7199 8476 -7188 8522
rect -7657 8456 -7188 8476
rect -7106 8476 -7093 8522
rect -6919 8476 -6906 8522
rect -7657 8436 -7640 8456
rect -7106 8455 -7089 8476
rect -7033 8455 -6979 8476
rect -6923 8455 -6906 8476
rect -7106 8449 -6906 8455
rect -6828 8476 -6813 8522
rect -6639 8476 -6533 8522
rect -6359 8476 -6344 8522
rect -6828 8465 -6344 8476
rect -6268 8522 -5788 8524
rect -5710 8522 -5229 8536
rect -3889 8534 -3872 8580
rect -3826 8534 -3809 8580
rect -5150 8522 -4669 8532
rect -3889 8529 -3809 8534
rect -4306 8522 -3809 8529
rect -6268 8476 -6253 8522
rect -6079 8476 -5973 8522
rect -5799 8476 -5784 8522
rect -7720 8384 -7640 8436
rect -7720 8338 -7703 8384
rect -7657 8338 -7640 8384
rect -6828 8382 -6345 8465
rect -6268 8393 -5784 8476
rect -6267 8368 -5784 8393
rect -5710 8476 -5693 8522
rect -5519 8476 -5413 8522
rect -5239 8476 -5224 8522
rect -5710 8464 -5224 8476
rect -5150 8476 -5133 8522
rect -4959 8476 -4853 8522
rect -4679 8476 -4664 8522
rect -4586 8487 -4573 8522
rect -5150 8464 -4664 8476
rect -4590 8476 -4573 8487
rect -4399 8476 -4386 8522
rect -5710 8366 -5229 8464
rect -5150 8362 -4669 8464
rect -4590 8455 -4569 8476
rect -4513 8455 -4459 8476
rect -4403 8455 -4386 8476
rect -4306 8476 -4293 8522
rect -4119 8482 -3809 8522
rect -4119 8476 -3872 8482
rect -4306 8461 -3872 8476
rect -4590 8449 -4386 8455
rect -7720 8286 -7640 8338
rect -7720 8240 -7703 8286
rect -7657 8240 -7640 8286
rect -7720 8188 -7640 8240
rect -7720 8142 -7703 8188
rect -7657 8142 -7640 8188
rect -7720 8090 -7640 8142
rect -7720 8044 -7703 8090
rect -7657 8044 -7640 8090
rect -7720 7992 -7640 8044
rect -7720 7946 -7703 7992
rect -7657 7946 -7640 7992
rect -7720 7940 -7640 7946
rect -7720 7930 -7186 7940
rect -7720 7894 -7373 7930
rect -7720 7848 -7703 7894
rect -7657 7884 -7373 7894
rect -7199 7884 -7186 7930
rect -7657 7872 -7186 7884
rect -7106 7930 -6623 8024
rect -7106 7884 -7093 7930
rect -6919 7884 -6813 7930
rect -6639 7884 -6623 7930
rect -7657 7848 -7640 7872
rect -7106 7870 -6623 7884
rect -6548 7942 -6065 8025
rect -5987 7942 -5507 8006
rect -5429 7942 -4948 8043
rect -4819 8036 -4673 8362
rect -4590 8036 -4401 8449
rect -3889 8436 -3872 8461
rect -3826 8436 -3809 8482
rect -3889 8384 -3809 8436
rect -3889 8338 -3872 8384
rect -3826 8338 -3809 8384
rect -3889 8286 -3809 8338
rect -3889 8240 -3872 8286
rect -3826 8240 -3809 8286
rect -3889 8188 -3809 8240
rect -3889 8142 -3872 8188
rect -3826 8142 -3809 8188
rect -3889 8090 -3809 8142
rect -3889 8044 -3872 8090
rect -3826 8044 -3809 8090
rect -6548 7930 -6064 7942
rect -6548 7884 -6533 7930
rect -6359 7884 -6253 7930
rect -6079 7884 -6064 7930
rect -5987 7930 -5504 7942
rect -5987 7884 -5973 7930
rect -5799 7884 -5693 7930
rect -5519 7884 -5504 7930
rect -5429 7930 -4944 7942
rect -5429 7884 -5413 7930
rect -5239 7884 -5133 7930
rect -4959 7884 -4944 7930
rect -4865 7930 -4384 8036
rect -3889 7992 -3809 8044
rect -3889 7946 -3872 7992
rect -3826 7946 -3809 7992
rect -3889 7940 -3809 7946
rect -4865 7884 -4853 7930
rect -4679 7884 -4573 7930
rect -4399 7884 -4384 7930
rect -6548 7871 -6065 7884
rect -5987 7875 -5507 7884
rect -5429 7873 -4948 7884
rect -4865 7866 -4384 7884
rect -4306 7930 -3809 7940
rect -4306 7884 -4293 7930
rect -4119 7894 -3809 7930
rect -4119 7884 -3872 7894
rect -4306 7872 -3872 7884
rect -7720 7796 -7640 7848
rect -7720 7750 -7703 7796
rect -7657 7750 -7640 7796
rect -7720 7698 -7640 7750
rect -7720 7652 -7703 7698
rect -7657 7652 -7640 7698
rect -7720 7617 -7640 7652
rect -3889 7848 -3872 7872
rect -3826 7848 -3809 7894
rect -3889 7796 -3809 7848
rect -3889 7750 -3872 7796
rect -3826 7750 -3809 7796
rect -3889 7698 -3809 7750
rect -3889 7652 -3872 7698
rect -3826 7652 -3809 7698
rect -3889 7617 -3809 7652
rect -7720 7600 -3809 7617
rect -7720 7554 -7703 7600
rect -7657 7554 -7605 7600
rect -7559 7554 -7507 7600
rect -7461 7554 -7409 7600
rect -7363 7554 -7311 7600
rect -7265 7554 -7213 7600
rect -7167 7554 -7115 7600
rect -7069 7554 -7017 7600
rect -6971 7554 -6919 7600
rect -6873 7554 -6821 7600
rect -6775 7554 -6723 7600
rect -6677 7554 -6625 7600
rect -6579 7554 -6527 7600
rect -6481 7554 -6429 7600
rect -6383 7554 -6331 7600
rect -6285 7554 -6233 7600
rect -6187 7554 -6135 7600
rect -6089 7554 -6037 7600
rect -5991 7554 -5939 7600
rect -5893 7554 -5841 7600
rect -5795 7554 -5743 7600
rect -5697 7554 -5645 7600
rect -5599 7554 -5547 7600
rect -5501 7554 -5449 7600
rect -5403 7554 -5351 7600
rect -5305 7554 -5253 7600
rect -5207 7554 -5155 7600
rect -5109 7554 -5057 7600
rect -5011 7554 -4959 7600
rect -4913 7554 -4861 7600
rect -4815 7554 -4763 7600
rect -4717 7554 -4665 7600
rect -4619 7554 -4567 7600
rect -4521 7554 -4469 7600
rect -4423 7554 -4371 7600
rect -4325 7554 -4273 7600
rect -4227 7554 -4175 7600
rect -4129 7554 -4077 7600
rect -4031 7554 -3979 7600
rect -3933 7554 -3872 7600
rect -3826 7554 -3809 7600
rect 497 9064 530 9079
rect 576 9064 609 9110
rect 497 9016 609 9064
rect 497 8970 530 9016
rect 576 8970 609 9016
rect 497 8922 609 8970
rect 497 8876 530 8922
rect 576 8876 609 8922
rect 497 8828 609 8876
rect 497 8782 530 8828
rect 576 8782 609 8828
rect 497 8734 609 8782
rect 497 8688 530 8734
rect 576 8688 609 8734
rect 497 8640 609 8688
rect 497 8594 530 8640
rect 576 8594 609 8640
rect 497 8546 609 8594
rect 497 8500 530 8546
rect 576 8500 609 8546
rect 497 8452 609 8500
rect 497 8406 530 8452
rect 576 8406 609 8452
rect 497 8358 609 8406
rect 497 8312 530 8358
rect 576 8312 609 8358
rect 497 8264 609 8312
rect 497 8218 530 8264
rect 576 8218 609 8264
rect 497 8170 609 8218
rect 497 8124 530 8170
rect 576 8124 609 8170
rect 497 8076 609 8124
rect 497 8030 530 8076
rect 576 8030 609 8076
rect 497 7982 609 8030
rect 497 7936 530 7982
rect 576 7936 609 7982
rect 497 7888 609 7936
rect 497 7842 530 7888
rect 576 7842 609 7888
rect 497 7794 609 7842
rect 497 7748 530 7794
rect 576 7748 609 7794
rect 497 7700 609 7748
rect 497 7654 530 7700
rect 576 7654 609 7700
rect 497 7606 609 7654
rect 226 7585 406 7595
rect -7720 7537 -3809 7554
rect 0 7583 406 7585
rect 0 7545 238 7583
rect -7612 7455 -3909 7537
rect -12 7531 238 7545
rect 290 7531 342 7583
rect 394 7531 406 7583
rect -12 7479 406 7531
rect -7720 7438 -3809 7455
rect -7720 7392 -7703 7438
rect -7657 7392 -7605 7438
rect -7559 7392 -7507 7438
rect -7461 7392 -7409 7438
rect -7363 7392 -7311 7438
rect -7265 7392 -7213 7438
rect -7167 7392 -7115 7438
rect -7069 7392 -7017 7438
rect -6971 7392 -6919 7438
rect -6873 7392 -6821 7438
rect -6775 7392 -6723 7438
rect -6677 7392 -6625 7438
rect -6579 7392 -6527 7438
rect -6481 7392 -6429 7438
rect -6383 7392 -6331 7438
rect -6285 7392 -6233 7438
rect -6187 7392 -6135 7438
rect -6089 7392 -6037 7438
rect -5991 7392 -5939 7438
rect -5893 7392 -5841 7438
rect -5795 7392 -5743 7438
rect -5697 7392 -5645 7438
rect -5599 7392 -5547 7438
rect -5501 7392 -5449 7438
rect -5403 7392 -5351 7438
rect -5305 7392 -5253 7438
rect -5207 7392 -5155 7438
rect -5109 7392 -5057 7438
rect -5011 7392 -4959 7438
rect -4913 7392 -4861 7438
rect -4815 7392 -4763 7438
rect -4717 7392 -4665 7438
rect -4619 7392 -4567 7438
rect -4521 7392 -4469 7438
rect -4423 7392 -4371 7438
rect -4325 7392 -4273 7438
rect -4227 7392 -4175 7438
rect -4129 7392 -4077 7438
rect -4031 7392 -3979 7438
rect -3933 7392 -3872 7438
rect -3826 7392 -3809 7438
rect -7720 7375 -3809 7392
rect -7720 7340 -7640 7375
rect -7720 7294 -7703 7340
rect -7657 7294 -7640 7340
rect -7720 7242 -7640 7294
rect -7720 7196 -7703 7242
rect -7657 7196 -7640 7242
rect -7720 7144 -7640 7196
rect -7720 7098 -7703 7144
rect -7657 7120 -7640 7144
rect -3889 7340 -3809 7375
rect -3889 7294 -3872 7340
rect -3826 7294 -3809 7340
rect -3889 7242 -3809 7294
rect -3889 7196 -3872 7242
rect -3826 7196 -3809 7242
rect -3889 7144 -3809 7196
rect -7657 7108 -7186 7120
rect -7657 7098 -7373 7108
rect -7720 7062 -7373 7098
rect -7199 7062 -7186 7108
rect -7720 7052 -7186 7062
rect -7109 7108 -6626 7118
rect -7109 7062 -7093 7108
rect -6919 7062 -6813 7108
rect -6639 7062 -6626 7108
rect -7720 7046 -7640 7052
rect -7720 7000 -7703 7046
rect -7657 7000 -7640 7046
rect -7720 6948 -7640 7000
rect -7109 6964 -6626 7062
rect -6547 7108 -6064 7124
rect -6547 7062 -6533 7108
rect -6359 7062 -6253 7108
rect -6079 7062 -6064 7108
rect -6547 6970 -6064 7062
rect -5987 7108 -5504 7124
rect -5987 7062 -5973 7108
rect -5799 7062 -5693 7108
rect -5519 7062 -5504 7108
rect -5987 6970 -5504 7062
rect -5427 7108 -4944 7121
rect -5427 7062 -5413 7108
rect -5239 7062 -5133 7108
rect -4959 7062 -4944 7108
rect -5427 6967 -4944 7062
rect -4866 7108 -4383 7123
rect -3889 7120 -3872 7144
rect -4866 7062 -4853 7108
rect -4679 7062 -4573 7108
rect -4399 7062 -4383 7108
rect -4866 6969 -4383 7062
rect -4306 7108 -3872 7120
rect -4306 7062 -4293 7108
rect -4119 7098 -3872 7108
rect -3826 7098 -3809 7144
rect -4119 7062 -3809 7098
rect -4306 7052 -3809 7062
rect -3889 7046 -3809 7052
rect -3889 7000 -3872 7046
rect -3826 7000 -3809 7046
rect -7720 6902 -7703 6948
rect -7657 6902 -7640 6948
rect -7720 6850 -7640 6902
rect -7720 6804 -7703 6850
rect -7657 6804 -7640 6850
rect -7720 6752 -7640 6804
rect -7720 6706 -7703 6752
rect -7657 6706 -7640 6752
rect -7720 6654 -7640 6706
rect -7720 6608 -7703 6654
rect -7657 6608 -7640 6654
rect -7720 6556 -7640 6608
rect -7720 6510 -7703 6556
rect -7657 6536 -7640 6556
rect -7106 6537 -6906 6543
rect -7657 6516 -7188 6536
rect -7657 6510 -7373 6516
rect -7720 6470 -7373 6510
rect -7199 6470 -7188 6516
rect -7106 6516 -7089 6537
rect -7033 6516 -6979 6537
rect -6923 6516 -6906 6537
rect -7106 6470 -7093 6516
rect -6919 6470 -6906 6516
rect -6826 6516 -6343 6612
rect -6826 6470 -6813 6516
rect -6639 6470 -6533 6516
rect -6359 6470 -6343 6516
rect -7720 6468 -7188 6470
rect -7720 6458 -7640 6468
rect -6826 6458 -6343 6470
rect -6266 6516 -5783 6612
rect -4846 6609 -4686 6969
rect -6266 6470 -6253 6516
rect -6079 6470 -5973 6516
rect -5799 6470 -5783 6516
rect -6266 6458 -5783 6470
rect -5704 6516 -5221 6609
rect -5704 6470 -5693 6516
rect -5519 6470 -5413 6516
rect -5239 6470 -5221 6516
rect -7720 6412 -7703 6458
rect -7657 6412 -7640 6458
rect -5704 6455 -5221 6470
rect -5147 6516 -4664 6609
rect -4568 6543 -4408 6969
rect -3889 6948 -3809 7000
rect -3889 6902 -3872 6948
rect -3826 6902 -3809 6948
rect -3889 6850 -3809 6902
rect -3889 6804 -3872 6850
rect -3826 6804 -3809 6850
rect -3889 6752 -3809 6804
rect -3889 6706 -3872 6752
rect -3826 6706 -3809 6752
rect -3889 6654 -3809 6706
rect -3889 6608 -3872 6654
rect -3826 6608 -3809 6654
rect -3889 6556 -3809 6608
rect -5147 6470 -5133 6516
rect -4959 6470 -4853 6516
rect -4679 6470 -4664 6516
rect -4586 6537 -4386 6543
rect -4586 6516 -4569 6537
rect -4513 6516 -4459 6537
rect -4403 6516 -4386 6537
rect -3889 6531 -3872 6556
rect -4586 6470 -4573 6516
rect -4399 6470 -4386 6516
rect -4306 6516 -3872 6531
rect -4306 6470 -4293 6516
rect -4119 6510 -3872 6516
rect -3826 6510 -3809 6556
rect -4119 6470 -3809 6510
rect -5147 6455 -4664 6470
rect -4306 6463 -3809 6470
rect -3889 6458 -3809 6463
rect -7720 6360 -7640 6412
rect -7720 6314 -7703 6360
rect -7657 6314 -7640 6360
rect -7720 6262 -7640 6314
rect -3889 6412 -3872 6458
rect -3826 6412 -3809 6458
rect -3889 6360 -3809 6412
rect -3889 6314 -3872 6360
rect -3826 6314 -3809 6360
rect -7720 6216 -7703 6262
rect -7657 6216 -7640 6262
rect -7720 6191 -7640 6216
rect -7005 6237 -5859 6305
rect -7005 6191 -6918 6237
rect -5946 6191 -5859 6237
rect -5046 6237 -4486 6305
rect -5046 6191 -4959 6237
rect -4573 6191 -4486 6237
rect -3889 6262 -3809 6314
rect -3889 6216 -3872 6262
rect -3826 6216 -3809 6262
rect -3889 6200 -3809 6216
rect -4306 6191 -3809 6200
rect -7720 6164 -7373 6191
rect -7720 6118 -7703 6164
rect -7657 6145 -7373 6164
rect -7199 6145 -7188 6191
rect -7104 6145 -7093 6191
rect -6919 6145 -6908 6191
rect -6826 6145 -6813 6191
rect -6639 6145 -6626 6191
rect -6544 6145 -6533 6191
rect -6359 6145 -6348 6191
rect -6264 6145 -6253 6191
rect -6079 6145 -6068 6191
rect -5984 6145 -5973 6191
rect -5799 6145 -5788 6191
rect -5704 6145 -5693 6191
rect -5519 6145 -5508 6191
rect -5424 6145 -5413 6191
rect -5239 6145 -5228 6191
rect -5144 6145 -5133 6191
rect -4959 6145 -4948 6191
rect -4866 6145 -4853 6191
rect -4679 6145 -4666 6191
rect -4584 6145 -4573 6191
rect -4399 6145 -4388 6191
rect -4306 6145 -4293 6191
rect -4119 6164 -3809 6191
rect -4119 6145 -3872 6164
rect -7657 6123 -7188 6145
rect -6826 6129 -6809 6145
rect -6753 6129 -6699 6145
rect -6643 6129 -6626 6145
rect -7657 6118 -7640 6123
rect -6826 6118 -6626 6129
rect -7720 6066 -7640 6118
rect -7720 6020 -7703 6066
rect -7657 6020 -7640 6066
rect -7720 5968 -7640 6020
rect -7720 5922 -7703 5968
rect -7657 5922 -7640 5968
rect -7720 5870 -7640 5922
rect -7720 5824 -7703 5870
rect -7657 5824 -7640 5870
rect -7720 5772 -7640 5824
rect -7720 5726 -7703 5772
rect -7657 5726 -7640 5772
rect -7720 5674 -7640 5726
rect -6786 5776 -6707 6118
rect -6446 5984 -6359 6145
rect -6166 6099 -6079 6145
rect -5693 6099 -5606 6145
rect -6166 6031 -5606 6099
rect -5368 5984 -5300 6145
rect -4866 6129 -4849 6145
rect -4793 6129 -4739 6145
rect -4683 6129 -4666 6145
rect -4306 6132 -3872 6145
rect -4866 6118 -4666 6129
rect -3889 6118 -3872 6132
rect -3826 6118 -3809 6164
rect -6446 5916 -5300 5984
rect -3889 6066 -3809 6118
rect -3889 6020 -3872 6066
rect -3826 6020 -3809 6066
rect -3889 5968 -3809 6020
rect -3889 5922 -3872 5968
rect -3826 5922 -3809 5968
rect -3889 5870 -3809 5922
rect -3889 5824 -3872 5870
rect -3826 5824 -3809 5870
rect -6786 5697 -6438 5776
rect -3889 5772 -3809 5824
rect -7720 5628 -7703 5674
rect -7657 5628 -7640 5674
rect -7720 5621 -7640 5628
rect -7720 5599 -7188 5621
rect -7720 5576 -7373 5599
rect -7720 5530 -7703 5576
rect -7657 5553 -7373 5576
rect -7199 5553 -7188 5599
rect -7106 5620 -6906 5626
rect -7106 5599 -7089 5620
rect -7033 5599 -6979 5620
rect -6923 5599 -6906 5620
rect -6517 5599 -6438 5697
rect -5886 5672 -4740 5740
rect -5886 5599 -5799 5672
rect -5426 5620 -5226 5626
rect -5426 5599 -5409 5620
rect -5353 5599 -5299 5620
rect -5243 5599 -5226 5620
rect -4808 5599 -4740 5672
rect -3889 5726 -3872 5772
rect -3826 5726 -3809 5772
rect -3889 5674 -3809 5726
rect -3889 5628 -3872 5674
rect -3826 5628 -3809 5674
rect -4586 5620 -4386 5626
rect -4586 5599 -4569 5620
rect -4513 5599 -4459 5620
rect -4403 5599 -4386 5620
rect -3889 5615 -3809 5628
rect -7106 5553 -7093 5599
rect -6919 5553 -6906 5599
rect -6824 5553 -6813 5599
rect -6639 5553 -6628 5599
rect -6544 5553 -6533 5599
rect -6359 5553 -6348 5599
rect -6264 5553 -6253 5599
rect -6079 5553 -6068 5599
rect -5984 5553 -5973 5599
rect -5799 5553 -5788 5599
rect -5704 5553 -5693 5599
rect -5519 5553 -5508 5599
rect -5426 5553 -5413 5599
rect -5239 5553 -5226 5599
rect -5144 5553 -5133 5599
rect -4959 5553 -4948 5599
rect -4864 5553 -4853 5599
rect -4679 5553 -4668 5599
rect -4586 5553 -4573 5599
rect -4399 5553 -4386 5599
rect -4305 5599 -3809 5615
rect -4305 5553 -4293 5599
rect -4119 5576 -3809 5599
rect -4119 5553 -3872 5576
rect -7657 5530 -7640 5553
rect -7720 5478 -7640 5530
rect -7720 5432 -7703 5478
rect -7657 5432 -7640 5478
rect -6726 5507 -6639 5553
rect -6253 5507 -6166 5553
rect -6726 5439 -6166 5507
rect -5606 5507 -5519 5553
rect -5133 5507 -5046 5553
rect -5606 5439 -5046 5507
rect -7720 5380 -7640 5432
rect -4573 5389 -4505 5553
rect -4305 5547 -3872 5553
rect -7720 5334 -7703 5380
rect -7657 5334 -7640 5380
rect -7720 5282 -7640 5334
rect -7720 5236 -7703 5282
rect -7657 5273 -7640 5282
rect -7007 5320 -6447 5388
rect -7007 5274 -6920 5320
rect -6534 5274 -6447 5320
rect -5886 5320 -5326 5388
rect -5886 5274 -5799 5320
rect -5413 5274 -5326 5320
rect -4789 5321 -4505 5389
rect -3889 5530 -3872 5547
rect -3826 5530 -3809 5576
rect -3889 5478 -3809 5530
rect -3889 5432 -3872 5478
rect -3826 5432 -3809 5478
rect -3889 5380 -3809 5432
rect -3889 5334 -3872 5380
rect -3826 5334 -3809 5380
rect -4789 5274 -4702 5321
rect -3889 5284 -3809 5334
rect -4306 5282 -3809 5284
rect -4306 5274 -3872 5282
rect -7384 5273 -7373 5274
rect -7657 5236 -7373 5273
rect -7720 5228 -7373 5236
rect -7199 5273 -7188 5274
rect -7199 5228 -7187 5273
rect -7104 5228 -7093 5274
rect -6919 5228 -6908 5274
rect -6824 5228 -6813 5274
rect -6639 5228 -6628 5274
rect -6544 5228 -6533 5274
rect -6359 5228 -6348 5274
rect -6264 5228 -6253 5274
rect -6079 5228 -6068 5274
rect -5984 5228 -5973 5274
rect -5799 5228 -5788 5274
rect -5704 5228 -5693 5274
rect -5519 5228 -5508 5274
rect -5424 5228 -5413 5274
rect -5239 5228 -5228 5274
rect -5144 5228 -5133 5274
rect -4959 5228 -4948 5274
rect -4864 5228 -4853 5274
rect -4679 5228 -4668 5274
rect -4586 5228 -4573 5274
rect -4399 5228 -4386 5274
rect -7720 5205 -7187 5228
rect -7720 5184 -7640 5205
rect -7720 5138 -7703 5184
rect -7657 5138 -7640 5184
rect -7720 5086 -7640 5138
rect -6726 5182 -6639 5228
rect -6253 5182 -6166 5228
rect -6726 5114 -6166 5182
rect -5606 5182 -5519 5228
rect -5133 5182 -5046 5228
rect -4586 5212 -4569 5228
rect -4513 5212 -4459 5228
rect -4403 5212 -4386 5228
rect -4306 5228 -4293 5274
rect -4119 5236 -3872 5274
rect -3826 5236 -3809 5282
rect -4119 5228 -3809 5236
rect -4306 5216 -3809 5228
rect -4586 5201 -4386 5212
rect -5606 5114 -5046 5182
rect -3889 5184 -3809 5216
rect -3889 5138 -3872 5184
rect -3826 5138 -3809 5184
rect -7720 5040 -7703 5086
rect -7657 5040 -7640 5086
rect -7720 4988 -7640 5040
rect -7720 4942 -7703 4988
rect -7657 4942 -7640 4988
rect -7720 4890 -7640 4942
rect -7720 4844 -7703 4890
rect -7657 4844 -7640 4890
rect -7720 4792 -7640 4844
rect -3889 5086 -3809 5138
rect -3889 5040 -3872 5086
rect -3826 5040 -3809 5086
rect -3889 4988 -3809 5040
rect -3889 4942 -3872 4988
rect -3826 4942 -3809 4988
rect -3889 4890 -3809 4942
rect -3889 4844 -3872 4890
rect -3826 4844 -3809 4890
rect -7720 4746 -7703 4792
rect -7657 4746 -7640 4792
rect -7720 4697 -7640 4746
rect -6167 4728 -5607 4796
rect -7106 4703 -6906 4709
rect -7720 4694 -7188 4697
rect -7720 4648 -7703 4694
rect -7657 4682 -7188 4694
rect -7657 4648 -7373 4682
rect -7720 4636 -7373 4648
rect -7199 4636 -7188 4682
rect -7106 4682 -7089 4703
rect -7033 4682 -6979 4703
rect -6923 4682 -6906 4703
rect -7106 4636 -7093 4682
rect -6919 4636 -6906 4682
rect -6826 4703 -6626 4709
rect -6826 4682 -6809 4703
rect -6753 4682 -6699 4703
rect -6643 4682 -6626 4703
rect -6167 4682 -6080 4728
rect -5694 4682 -5607 4728
rect -5047 4728 -4487 4796
rect -5047 4682 -4960 4728
rect -4574 4682 -4487 4728
rect -3889 4792 -3809 4844
rect -3889 4746 -3872 4792
rect -3826 4746 -3809 4792
rect -3889 4697 -3809 4746
rect -4303 4694 -3809 4697
rect -4303 4682 -3872 4694
rect -6826 4636 -6813 4682
rect -6639 4636 -6626 4682
rect -6544 4636 -6533 4682
rect -6359 4636 -6348 4682
rect -6264 4636 -6253 4682
rect -6079 4636 -6068 4682
rect -5984 4636 -5973 4682
rect -5799 4636 -5788 4682
rect -5704 4636 -5693 4682
rect -5519 4636 -5508 4682
rect -5424 4636 -5413 4682
rect -5239 4636 -5228 4682
rect -5144 4636 -5133 4682
rect -4959 4636 -4948 4682
rect -4864 4636 -4853 4682
rect -4679 4636 -4668 4682
rect -4584 4636 -4573 4682
rect -4399 4636 -4388 4682
rect -4304 4636 -4293 4682
rect -4119 4648 -3872 4682
rect -3826 4648 -3809 4694
rect -4119 4636 -3809 4648
rect -7720 4629 -7188 4636
rect -7720 4596 -7640 4629
rect -7720 4550 -7703 4596
rect -7657 4550 -7640 4596
rect -7720 4498 -7640 4550
rect -6446 4590 -6359 4636
rect -5973 4590 -5886 4636
rect -6446 4522 -5886 4590
rect -5326 4590 -5239 4636
rect -4853 4590 -4766 4636
rect -4303 4629 -3809 4636
rect -5326 4522 -4766 4590
rect -3889 4596 -3809 4629
rect -3889 4550 -3872 4596
rect -3826 4550 -3809 4596
rect -7720 4452 -7703 4498
rect -7657 4452 -7640 4498
rect -7720 4407 -7640 4452
rect -3889 4498 -3809 4550
rect -3889 4452 -3872 4498
rect -3826 4452 -3809 4498
rect -3889 4407 -3809 4452
rect -7720 4390 -3809 4407
rect -7720 4344 -7703 4390
rect -7657 4344 -7605 4390
rect -7559 4344 -7507 4390
rect -7461 4344 -7409 4390
rect -7363 4344 -7311 4390
rect -7265 4344 -7213 4390
rect -7167 4344 -7115 4390
rect -7069 4344 -7017 4390
rect -6971 4344 -6919 4390
rect -6873 4344 -6821 4390
rect -6775 4344 -6723 4390
rect -6677 4344 -6625 4390
rect -6579 4344 -6527 4390
rect -6481 4344 -6429 4390
rect -6383 4344 -6331 4390
rect -6285 4344 -6233 4390
rect -6187 4344 -6135 4390
rect -6089 4344 -6037 4390
rect -5991 4344 -5939 4390
rect -5893 4344 -5841 4390
rect -5795 4344 -5743 4390
rect -5697 4344 -5645 4390
rect -5599 4344 -5547 4390
rect -5501 4344 -5449 4390
rect -5403 4344 -5351 4390
rect -5305 4344 -5253 4390
rect -5207 4344 -5155 4390
rect -5109 4344 -5057 4390
rect -5011 4344 -4959 4390
rect -4913 4344 -4861 4390
rect -4815 4344 -4763 4390
rect -4717 4344 -4665 4390
rect -4619 4344 -4567 4390
rect -4521 4344 -4469 4390
rect -4423 4344 -4371 4390
rect -4325 4344 -4273 4390
rect -4227 4344 -4175 4390
rect -4129 4344 -4077 4390
rect -4031 4344 -3979 4390
rect -3933 4344 -3872 4390
rect -3826 4344 -3809 4390
rect -7720 4327 -3809 4344
rect -12 7427 238 7479
rect 290 7427 342 7479
rect 394 7427 406 7479
rect -12 7415 406 7427
rect 497 7560 530 7606
rect 576 7560 609 7606
rect 497 7512 609 7560
rect 497 7466 530 7512
rect 576 7466 609 7512
rect 497 7418 609 7466
rect -12 -83 292 7415
rect 497 7372 530 7418
rect 576 7381 609 7418
rect 911 10545 957 10793
rect 911 9783 957 9945
rect 911 9021 957 9183
rect 911 8363 957 8421
rect 1127 10545 1173 10793
rect 1127 9783 1173 9945
rect 1127 9021 1173 9183
rect 1008 8363 1076 8374
rect 1127 8363 1173 8421
rect 911 8317 1019 8363
rect 1065 8317 1173 8363
rect 911 8259 957 8317
rect 1008 8306 1076 8317
rect 911 7381 957 7659
rect 1127 8259 1173 8317
rect 1127 7381 1173 7659
rect 1343 10602 2685 10648
rect 1343 10545 1389 10602
rect 1343 9783 1389 9945
rect 1343 9021 1389 9183
rect 1343 8259 1389 8421
rect 1343 7648 1389 7659
rect 1559 10545 1605 10556
rect 1559 9783 1605 9945
rect 1559 9021 1605 9183
rect 1559 8259 1605 8421
rect 1227 7583 1407 7595
rect 1227 7531 1239 7583
rect 1291 7531 1343 7583
rect 1395 7531 1407 7583
rect 1227 7519 1407 7531
rect 1559 7381 1605 7659
rect 1775 10545 1821 10602
rect 1775 9783 1821 9945
rect 1775 9021 1821 9183
rect 1775 8259 1821 8421
rect 1775 7648 1821 7659
rect 1991 10545 2037 10556
rect 1991 9783 2037 9945
rect 1991 9021 2037 9183
rect 1991 8259 2037 8421
rect 1991 7381 2037 7659
rect 2207 10545 2253 10602
rect 2207 9783 2253 9945
rect 2207 9021 2253 9183
rect 2207 8259 2253 8421
rect 2207 7648 2253 7659
rect 2423 10545 2469 10556
rect 2639 10545 2685 10602
rect 2520 10323 2639 10335
rect 2855 10545 2901 10793
rect 2685 10323 2700 10335
rect 2520 10271 2532 10323
rect 2584 10271 2636 10323
rect 2688 10271 2700 10323
rect 2520 10219 2639 10271
rect 2685 10219 2700 10271
rect 2520 10167 2532 10219
rect 2584 10167 2636 10219
rect 2688 10167 2700 10219
rect 2520 10155 2639 10167
rect 2423 9783 2469 9945
rect 2685 10155 2700 10167
rect 2639 9783 2685 9945
rect 2624 9457 2639 9469
rect 2855 9783 2901 9945
rect 2685 9457 2700 9469
rect 2624 9405 2636 9457
rect 2688 9405 2700 9457
rect 2624 9353 2639 9405
rect 2685 9353 2700 9405
rect 2624 9301 2636 9353
rect 2688 9301 2700 9353
rect 2624 9289 2639 9301
rect 2423 9021 2469 9183
rect 2423 8259 2469 8421
rect 2685 9289 2700 9301
rect 2639 9021 2685 9183
rect 2639 8259 2685 8421
rect 2624 8127 2639 8139
rect 2855 9021 2901 9183
rect 2855 8363 2901 8421
rect 3071 10545 3117 10793
rect 3071 9783 3117 9945
rect 3071 9021 3117 9183
rect 2952 8363 3020 8374
rect 3071 8363 3117 8421
rect 2855 8317 2963 8363
rect 3009 8317 3117 8363
rect 2855 8259 2901 8317
rect 2952 8306 3020 8317
rect 2685 8127 2700 8139
rect 2624 8075 2636 8127
rect 2688 8075 2700 8127
rect 2624 8023 2639 8075
rect 2685 8023 2700 8075
rect 2624 7971 2636 8023
rect 2688 7971 2700 8023
rect 2624 7959 2639 7971
rect 2423 7381 2469 7659
rect 2685 7959 2700 7971
rect 2639 7648 2685 7659
rect 2855 7381 2901 7659
rect 3071 8259 3117 8317
rect 3071 7381 3117 7659
rect 3411 10756 3444 10793
rect 3490 10756 3523 10802
rect 3411 10708 3523 10756
rect 3411 10662 3444 10708
rect 3490 10662 3523 10708
rect 3411 10614 3523 10662
rect 3411 10568 3444 10614
rect 3490 10568 3523 10614
rect 3411 10520 3523 10568
rect 3411 10474 3444 10520
rect 3490 10474 3523 10520
rect 3411 10426 3523 10474
rect 3411 10380 3444 10426
rect 3490 10380 3523 10426
rect 3411 10332 3523 10380
rect 3411 10286 3444 10332
rect 3490 10286 3523 10332
rect 3411 10238 3523 10286
rect 3411 10192 3444 10238
rect 3490 10192 3523 10238
rect 3411 10144 3523 10192
rect 3411 10098 3444 10144
rect 3490 10098 3523 10144
rect 3411 10050 3523 10098
rect 3411 10004 3444 10050
rect 3490 10004 3523 10050
rect 3411 9956 3523 10004
rect 3411 9910 3444 9956
rect 3490 9910 3523 9956
rect 3411 9862 3523 9910
rect 3411 9816 3444 9862
rect 3490 9816 3523 9862
rect 3411 9768 3523 9816
rect 3411 9722 3444 9768
rect 3490 9722 3523 9768
rect 3411 9674 3523 9722
rect 3411 9628 3444 9674
rect 3490 9628 3523 9674
rect 3411 9580 3523 9628
rect 3411 9534 3444 9580
rect 3490 9534 3523 9580
rect 3411 9486 3523 9534
rect 3411 9440 3444 9486
rect 3490 9440 3523 9486
rect 3411 9392 3523 9440
rect 3411 9346 3444 9392
rect 3490 9346 3523 9392
rect 3411 9298 3523 9346
rect 3411 9252 3444 9298
rect 3490 9252 3523 9298
rect 3411 9204 3523 9252
rect 3411 9158 3444 9204
rect 3490 9158 3523 9204
rect 3411 9110 3523 9158
rect 3411 9064 3444 9110
rect 3490 9064 3523 9110
rect 3411 9016 3523 9064
rect 3411 8970 3444 9016
rect 3490 8970 3523 9016
rect 3411 8922 3523 8970
rect 3411 8876 3444 8922
rect 3490 8876 3523 8922
rect 3411 8828 3523 8876
rect 3411 8782 3444 8828
rect 3490 8782 3523 8828
rect 3411 8734 3523 8782
rect 3411 8688 3444 8734
rect 3490 8688 3523 8734
rect 3411 8640 3523 8688
rect 3411 8594 3444 8640
rect 3490 8594 3523 8640
rect 3411 8546 3523 8594
rect 3411 8500 3444 8546
rect 3490 8500 3523 8546
rect 3411 8452 3523 8500
rect 3411 8406 3444 8452
rect 3490 8406 3523 8452
rect 3411 8358 3523 8406
rect 3411 8312 3444 8358
rect 3490 8312 3523 8358
rect 3411 8264 3523 8312
rect 3411 8218 3444 8264
rect 3490 8218 3523 8264
rect 3411 8170 3523 8218
rect 3411 8124 3444 8170
rect 3490 8124 3523 8170
rect 3411 8076 3523 8124
rect 3411 8030 3444 8076
rect 3490 8030 3523 8076
rect 3411 7982 3523 8030
rect 3411 7936 3444 7982
rect 3490 7936 3523 7982
rect 3411 7888 3523 7936
rect 3411 7842 3444 7888
rect 3490 7842 3523 7888
rect 3411 7794 3523 7842
rect 3411 7748 3444 7794
rect 3490 7748 3523 7794
rect 3411 7700 3523 7748
rect 3411 7654 3444 7700
rect 3490 7654 3523 7700
rect 3411 7606 3523 7654
rect 3411 7560 3444 7606
rect 3490 7560 3523 7606
rect 3411 7512 3523 7560
rect 3411 7466 3444 7512
rect 3490 7466 3523 7512
rect 3411 7418 3523 7466
rect 3411 7381 3444 7418
rect 576 7372 3444 7381
rect 3490 7381 3523 7418
rect 3597 14013 3643 14281
rect 3597 12883 3643 13289
rect 3597 11753 3643 12159
rect 3597 10623 3643 11029
rect 3597 9493 3643 9899
rect 3597 8589 3643 8769
rect 3757 14013 3803 14281
rect 3950 14222 4026 14234
rect 3950 14170 3962 14222
rect 4014 14219 4026 14222
rect 4014 14173 4445 14219
rect 4491 14173 5085 14219
rect 5131 14173 5142 14219
rect 4014 14170 4026 14173
rect 3950 14158 4026 14170
rect 4045 14070 5051 14116
rect 3885 14013 3931 14024
rect 3870 13481 3885 13493
rect 4045 14013 4091 14070
rect 4030 13977 4045 13989
rect 4205 14013 4251 14024
rect 4091 13977 4106 13989
rect 4030 13925 4042 13977
rect 4094 13925 4106 13977
rect 4030 13873 4045 13925
rect 4091 13873 4106 13925
rect 4030 13821 4042 13873
rect 4094 13821 4106 13873
rect 4030 13809 4045 13821
rect 3931 13481 3946 13493
rect 3870 13429 3882 13481
rect 3934 13429 3946 13481
rect 3870 13377 3885 13429
rect 3931 13377 3946 13429
rect 3870 13325 3882 13377
rect 3934 13325 3946 13377
rect 3870 13313 3885 13325
rect 3757 12883 3803 13289
rect 3931 13313 3946 13325
rect 3885 13278 3931 13289
rect 4091 13809 4106 13821
rect 4190 13977 4205 13989
rect 4365 14013 4411 14070
rect 4251 13977 4266 13989
rect 4190 13925 4202 13977
rect 4254 13925 4266 13977
rect 4190 13873 4205 13925
rect 4251 13873 4266 13925
rect 4190 13821 4202 13873
rect 4254 13821 4266 13873
rect 4190 13809 4205 13821
rect 4045 13278 4091 13289
rect 4251 13809 4266 13821
rect 4205 13278 4251 13289
rect 4525 14013 4571 14024
rect 4510 13481 4525 13493
rect 4685 14013 4731 14070
rect 4571 13481 4586 13493
rect 4510 13429 4522 13481
rect 4574 13429 4586 13481
rect 4510 13377 4525 13429
rect 4571 13377 4586 13429
rect 4510 13325 4522 13377
rect 4574 13325 4586 13377
rect 4510 13313 4525 13325
rect 4365 13278 4411 13289
rect 4571 13313 4586 13325
rect 4525 13278 4571 13289
rect 4845 14013 4891 14024
rect 4831 13977 4845 13989
rect 5005 14013 5051 14070
rect 4891 13977 4907 13989
rect 4831 13925 4843 13977
rect 4895 13925 4907 13977
rect 4831 13873 4845 13925
rect 4891 13873 4907 13925
rect 4831 13821 4843 13873
rect 4895 13821 4907 13873
rect 4831 13809 4845 13821
rect 4685 13278 4731 13289
rect 4891 13809 4907 13821
rect 4845 13278 4891 13289
rect 5165 14013 5211 14024
rect 5150 13481 5165 13493
rect 5293 14013 5339 14281
rect 5211 13481 5226 13493
rect 5150 13429 5162 13481
rect 5214 13429 5226 13481
rect 5150 13377 5165 13429
rect 5211 13377 5226 13429
rect 5150 13325 5162 13377
rect 5214 13325 5226 13377
rect 5150 13313 5165 13325
rect 5005 13278 5051 13289
rect 5211 13313 5226 13325
rect 5165 13278 5211 13289
rect 3950 13198 4026 13210
rect 3950 13146 3962 13198
rect 4014 13146 4026 13198
rect 3950 13094 4026 13146
rect 3950 13042 3962 13094
rect 4014 13091 4026 13094
rect 4014 13045 4125 13091
rect 4171 13045 4445 13091
rect 4491 13045 4765 13091
rect 4811 13045 5085 13091
rect 5131 13045 5142 13091
rect 4014 13042 4026 13045
rect 3950 13030 4026 13042
rect 4045 12940 5051 12986
rect 3885 12883 3931 12894
rect 3870 12455 3885 12467
rect 4045 12883 4091 12940
rect 4030 12847 4045 12859
rect 4205 12883 4251 12894
rect 4091 12847 4106 12859
rect 4030 12795 4042 12847
rect 4094 12795 4106 12847
rect 4030 12743 4045 12795
rect 4091 12743 4106 12795
rect 4030 12691 4042 12743
rect 4094 12691 4106 12743
rect 4030 12679 4045 12691
rect 3931 12455 3946 12467
rect 3870 12403 3882 12455
rect 3934 12403 3946 12455
rect 3870 12351 3885 12403
rect 3931 12351 3946 12403
rect 3870 12299 3882 12351
rect 3934 12299 3946 12351
rect 3870 12287 3885 12299
rect 3757 11753 3803 12159
rect 3931 12287 3946 12299
rect 3885 12148 3931 12159
rect 4091 12679 4106 12691
rect 4190 12847 4205 12859
rect 4365 12883 4411 12940
rect 4251 12847 4266 12859
rect 4190 12795 4202 12847
rect 4254 12795 4266 12847
rect 4190 12743 4205 12795
rect 4251 12743 4266 12795
rect 4190 12691 4202 12743
rect 4254 12691 4266 12743
rect 4190 12679 4205 12691
rect 4045 12148 4091 12159
rect 4251 12679 4266 12691
rect 4205 12148 4251 12159
rect 4525 12883 4571 12894
rect 4510 12455 4525 12467
rect 4685 12883 4731 12940
rect 4571 12455 4586 12467
rect 4510 12403 4522 12455
rect 4574 12403 4586 12455
rect 4510 12351 4525 12403
rect 4571 12351 4586 12403
rect 4510 12299 4522 12351
rect 4574 12299 4586 12351
rect 4510 12287 4525 12299
rect 4365 12148 4411 12159
rect 4571 12287 4586 12299
rect 4525 12148 4571 12159
rect 4845 12883 4891 12894
rect 4831 12847 4845 12859
rect 5005 12883 5051 12940
rect 4891 12847 4907 12859
rect 4831 12795 4843 12847
rect 4895 12795 4907 12847
rect 4831 12743 4845 12795
rect 4891 12743 4907 12795
rect 4831 12691 4843 12743
rect 4895 12691 4907 12743
rect 4831 12679 4845 12691
rect 4685 12148 4731 12159
rect 4891 12679 4907 12691
rect 4845 12148 4891 12159
rect 5165 12883 5211 12894
rect 5150 12455 5165 12467
rect 5293 12883 5339 13289
rect 5211 12455 5226 12467
rect 5150 12403 5162 12455
rect 5214 12403 5226 12455
rect 5150 12351 5165 12403
rect 5211 12351 5226 12403
rect 5150 12299 5162 12351
rect 5214 12299 5226 12351
rect 5150 12287 5165 12299
rect 5005 12148 5051 12159
rect 5211 12287 5226 12299
rect 5165 12148 5211 12159
rect 3950 12068 4026 12080
rect 3950 12016 3962 12068
rect 4014 12016 4026 12068
rect 3950 11964 4026 12016
rect 3950 11912 3962 11964
rect 4014 11963 4026 11964
rect 4014 11917 4125 11963
rect 4171 11917 4445 11963
rect 4491 11917 4765 11963
rect 4811 11917 5085 11963
rect 5131 11917 5142 11963
rect 4014 11912 4026 11917
rect 3950 11900 4026 11912
rect 4045 11810 5051 11856
rect 3885 11753 3931 11764
rect 3870 11221 3885 11233
rect 4045 11753 4091 11810
rect 3931 11221 3946 11233
rect 3870 11169 3882 11221
rect 3934 11169 3946 11221
rect 3870 11117 3885 11169
rect 3931 11117 3946 11169
rect 3870 11065 3882 11117
rect 3934 11065 3946 11117
rect 3870 11053 3885 11065
rect 3757 10623 3803 11029
rect 3757 9493 3803 9899
rect 3931 11053 3946 11065
rect 3885 10623 3931 11029
rect 4205 11753 4251 11764
rect 4190 11717 4205 11729
rect 4365 11753 4411 11810
rect 4251 11717 4266 11729
rect 4190 11665 4202 11717
rect 4254 11665 4266 11717
rect 4190 11613 4205 11665
rect 4251 11613 4266 11665
rect 4190 11561 4202 11613
rect 4254 11561 4266 11613
rect 4190 11549 4205 11561
rect 4045 10623 4091 11029
rect 4030 10323 4045 10335
rect 4251 11549 4266 11561
rect 4205 10623 4251 11029
rect 4091 10323 4106 10335
rect 4030 10271 4042 10323
rect 4094 10271 4106 10323
rect 4030 10219 4045 10271
rect 4091 10219 4106 10271
rect 4030 10167 4042 10219
rect 4094 10167 4106 10219
rect 4030 10155 4045 10167
rect 3885 9888 3931 9899
rect 4091 10155 4106 10167
rect 4045 9888 4091 9899
rect 4205 9888 4251 9899
rect 4525 11753 4571 11764
rect 4510 11221 4525 11233
rect 4685 11753 4731 11810
rect 4571 11221 4586 11233
rect 4510 11169 4522 11221
rect 4574 11169 4586 11221
rect 4510 11117 4525 11169
rect 4571 11117 4586 11169
rect 4510 11065 4522 11117
rect 4574 11065 4586 11117
rect 4510 11053 4525 11065
rect 4365 10623 4411 11029
rect 4365 9888 4411 9899
rect 4571 11053 4586 11065
rect 4525 10623 4571 11029
rect 4525 9888 4571 9899
rect 4845 11753 4891 11764
rect 4831 11717 4845 11729
rect 5005 11753 5051 11810
rect 4891 11717 4907 11729
rect 4831 11665 4843 11717
rect 4895 11665 4907 11717
rect 4831 11613 4845 11665
rect 4891 11613 4907 11665
rect 4831 11561 4843 11613
rect 4895 11561 4907 11613
rect 4831 11549 4845 11561
rect 4685 10623 4731 11029
rect 4685 9888 4731 9899
rect 4891 11549 4907 11561
rect 4845 10623 4891 11029
rect 4845 9888 4891 9899
rect 5165 11753 5211 11764
rect 5150 11221 5165 11233
rect 5293 11753 5339 12159
rect 5211 11221 5226 11233
rect 5150 11169 5162 11221
rect 5214 11169 5226 11221
rect 5150 11117 5165 11169
rect 5211 11117 5226 11169
rect 5150 11065 5162 11117
rect 5214 11065 5226 11117
rect 5150 11053 5165 11065
rect 5005 10623 5051 11029
rect 5005 9888 5051 9899
rect 5211 11053 5226 11065
rect 5165 10623 5211 11029
rect 5165 9888 5211 9899
rect 5293 10623 5339 11029
rect 3950 9810 4026 9822
rect 3950 9758 3962 9810
rect 4014 9758 4026 9810
rect 3950 9706 4026 9758
rect 3950 9654 3962 9706
rect 4014 9703 4026 9706
rect 4014 9657 4125 9703
rect 4171 9657 4445 9703
rect 4491 9657 4765 9703
rect 4811 9657 5085 9703
rect 5131 9657 5142 9703
rect 4014 9654 4026 9657
rect 3950 9640 4026 9654
rect 4045 9550 5051 9596
rect 3885 9493 3931 9504
rect 3870 8961 3885 8973
rect 4045 9493 4091 9550
rect 4030 9457 4045 9469
rect 4205 9493 4251 9504
rect 4091 9457 4106 9469
rect 4030 9405 4042 9457
rect 4094 9405 4106 9457
rect 4030 9353 4045 9405
rect 4091 9353 4106 9405
rect 4030 9301 4042 9353
rect 4094 9301 4106 9353
rect 4030 9289 4045 9301
rect 3931 8961 3946 8973
rect 3870 8909 3882 8961
rect 3934 8909 3946 8961
rect 3870 8857 3885 8909
rect 3931 8857 3946 8909
rect 3870 8805 3882 8857
rect 3934 8805 3946 8857
rect 3870 8793 3885 8805
rect 3757 8589 3803 8769
rect 3931 8793 3946 8805
rect 3885 8758 3931 8769
rect 4091 9289 4106 9301
rect 4190 9457 4205 9469
rect 4365 9493 4411 9550
rect 4251 9457 4266 9469
rect 4190 9405 4202 9457
rect 4254 9405 4266 9457
rect 4190 9353 4205 9405
rect 4251 9353 4266 9405
rect 4190 9301 4202 9353
rect 4254 9301 4266 9353
rect 4190 9289 4205 9301
rect 4045 8758 4091 8769
rect 4251 9289 4266 9301
rect 4205 8758 4251 8769
rect 4525 9493 4571 9504
rect 4510 8961 4525 8973
rect 4685 9493 4731 9550
rect 4571 8961 4586 8973
rect 4510 8909 4522 8961
rect 4574 8909 4586 8961
rect 4510 8857 4525 8909
rect 4571 8857 4586 8909
rect 4510 8805 4522 8857
rect 4574 8805 4586 8857
rect 4510 8793 4525 8805
rect 4365 8758 4411 8769
rect 4571 8793 4586 8805
rect 4525 8758 4571 8769
rect 4845 9493 4891 9504
rect 4831 9457 4845 9469
rect 5005 9493 5051 9550
rect 4891 9457 4907 9469
rect 4831 9405 4843 9457
rect 4895 9405 4907 9457
rect 4831 9353 4845 9405
rect 4891 9353 4907 9405
rect 4831 9301 4843 9353
rect 4895 9301 4907 9353
rect 4831 9289 4845 9301
rect 4685 8758 4731 8769
rect 4891 9289 4907 9301
rect 4845 8758 4891 8769
rect 5165 9493 5211 9504
rect 5150 8961 5165 8973
rect 5293 9493 5339 9899
rect 5211 8961 5226 8973
rect 5150 8909 5162 8961
rect 5214 8909 5226 8961
rect 5150 8857 5165 8909
rect 5211 8857 5226 8909
rect 5150 8805 5162 8857
rect 5214 8805 5226 8857
rect 5150 8793 5165 8805
rect 5005 8758 5051 8769
rect 5211 8793 5226 8805
rect 5165 8758 5211 8769
rect 3597 8543 3677 8589
rect 3723 8543 3803 8589
rect 3597 8363 3643 8543
rect 3597 7381 3643 7639
rect 3757 8363 3803 8543
rect 3950 8680 4026 8692
rect 3950 8628 3962 8680
rect 4014 8628 4026 8680
rect 3950 8576 4026 8628
rect 3950 8524 3962 8576
rect 4014 8573 4026 8576
rect 5293 8589 5339 8769
rect 5453 14013 5499 14281
rect 5453 12883 5499 13289
rect 5453 11753 5499 12159
rect 5453 10623 5499 11029
rect 5453 9493 5499 9899
rect 5453 8589 5499 8769
rect 4014 8527 4125 8573
rect 4171 8527 4445 8573
rect 4491 8527 4765 8573
rect 4811 8527 5085 8573
rect 5131 8527 5142 8573
rect 5293 8543 5373 8589
rect 5419 8543 5499 8589
rect 4014 8524 4026 8527
rect 3950 8512 4026 8524
rect 4045 8420 5051 8466
rect 3885 8363 3931 8374
rect 3870 7831 3885 7843
rect 4045 8363 4091 8420
rect 4030 8127 4045 8139
rect 4205 8363 4251 8374
rect 4190 8327 4205 8339
rect 4365 8363 4411 8420
rect 4251 8327 4266 8339
rect 4190 8275 4202 8327
rect 4254 8275 4266 8327
rect 4190 8223 4205 8275
rect 4251 8223 4266 8275
rect 4190 8171 4202 8223
rect 4254 8171 4266 8223
rect 4190 8159 4205 8171
rect 4091 8127 4106 8139
rect 4030 8075 4042 8127
rect 4094 8075 4106 8127
rect 4030 8023 4045 8075
rect 4091 8023 4106 8075
rect 4030 7971 4042 8023
rect 4094 7971 4106 8023
rect 4030 7959 4045 7971
rect 3931 7831 3946 7843
rect 3870 7779 3882 7831
rect 3934 7779 3946 7831
rect 3870 7727 3885 7779
rect 3931 7727 3946 7779
rect 3870 7675 3882 7727
rect 3934 7675 3946 7727
rect 3870 7663 3885 7675
rect 3757 7381 3803 7639
rect 3931 7663 3946 7675
rect 3885 7628 3931 7639
rect 4091 7959 4106 7971
rect 4045 7628 4091 7639
rect 4251 8159 4266 8171
rect 4205 7628 4251 7639
rect 4525 8363 4571 8374
rect 4510 7831 4525 7843
rect 4685 8363 4731 8420
rect 4571 7831 4586 7843
rect 4510 7779 4522 7831
rect 4574 7779 4586 7831
rect 4510 7727 4525 7779
rect 4571 7727 4586 7779
rect 4510 7675 4522 7727
rect 4574 7675 4586 7727
rect 4510 7663 4525 7675
rect 4365 7628 4411 7639
rect 4571 7663 4586 7675
rect 4525 7628 4571 7639
rect 4845 8363 4891 8374
rect 4831 8327 4845 8339
rect 5005 8363 5051 8420
rect 4891 8327 4907 8339
rect 4831 8275 4843 8327
rect 4895 8275 4907 8327
rect 4831 8223 4845 8275
rect 4891 8223 4907 8275
rect 4831 8171 4843 8223
rect 4895 8171 4907 8223
rect 4831 8159 4845 8171
rect 4685 7628 4731 7639
rect 4891 8159 4907 8171
rect 4845 7628 4891 7639
rect 5165 8363 5211 8374
rect 5150 7831 5165 7843
rect 5293 8363 5339 8543
rect 5211 7831 5226 7843
rect 5150 7779 5162 7831
rect 5214 7779 5226 7831
rect 5150 7727 5165 7779
rect 5211 7727 5226 7779
rect 5150 7675 5162 7727
rect 5214 7675 5226 7727
rect 5150 7663 5165 7675
rect 5005 7628 5051 7639
rect 5211 7663 5226 7675
rect 5165 7628 5211 7639
rect 4110 7492 4186 7504
rect 4110 7440 4122 7492
rect 4174 7489 4186 7492
rect 4174 7443 4765 7489
rect 4811 7443 4822 7489
rect 4174 7440 4186 7443
rect 4110 7428 4186 7440
rect 5293 7381 5339 7639
rect 5453 8363 5499 8543
rect 5453 7381 5499 7639
rect 5573 14280 5685 14281
rect 5573 14234 5606 14280
rect 5652 14234 5685 14280
rect 5573 14186 5685 14234
rect 5573 14140 5606 14186
rect 5652 14140 5685 14186
rect 5573 14092 5685 14140
rect 5731 14272 5911 14284
rect 5731 14220 5743 14272
rect 5795 14220 5847 14272
rect 5899 14220 5911 14272
rect 5731 14168 5911 14220
rect 5731 14116 5743 14168
rect 5795 14116 5847 14168
rect 5899 14116 5911 14168
rect 5731 14104 5911 14116
rect 5573 14046 5606 14092
rect 5652 14046 5685 14092
rect 5573 13998 5685 14046
rect 5573 13952 5606 13998
rect 5652 13952 5685 13998
rect 6013 13989 6173 14490
rect 6229 14477 6341 14525
rect 6229 14431 6262 14477
rect 6308 14431 6341 14477
rect 6229 14383 6341 14431
rect 6229 14337 6262 14383
rect 6308 14337 6341 14383
rect 6229 14289 6341 14337
rect 6229 14243 6262 14289
rect 6308 14243 6341 14289
rect 6229 14195 6341 14243
rect 6229 14149 6262 14195
rect 6308 14149 6341 14195
rect 6229 14101 6341 14149
rect 6229 14055 6262 14101
rect 6308 14055 6341 14101
rect 6229 14007 6341 14055
rect 5573 13904 5685 13952
rect 5573 13858 5606 13904
rect 5652 13858 5685 13904
rect 5573 13810 5685 13858
rect 5573 13764 5606 13810
rect 5652 13764 5685 13810
rect 6003 13977 6183 13989
rect 6003 13925 6015 13977
rect 6067 13925 6119 13977
rect 6171 13925 6183 13977
rect 6003 13873 6183 13925
rect 6003 13821 6015 13873
rect 6067 13821 6119 13873
rect 6171 13821 6183 13873
rect 6003 13809 6183 13821
rect 6229 13961 6262 14007
rect 6308 13961 6341 14007
rect 6229 13913 6341 13961
rect 6229 13867 6262 13913
rect 6308 13867 6341 13913
rect 6229 13819 6341 13867
rect 5573 13716 5685 13764
rect 5573 13670 5606 13716
rect 5652 13670 5685 13716
rect 5573 13622 5685 13670
rect 5573 13576 5606 13622
rect 5652 13576 5685 13622
rect 5573 13528 5685 13576
rect 5573 13482 5606 13528
rect 5652 13482 5685 13528
rect 5573 13434 5685 13482
rect 5573 13388 5606 13434
rect 5652 13388 5685 13434
rect 5573 13340 5685 13388
rect 5573 13294 5606 13340
rect 5652 13294 5685 13340
rect 5573 13246 5685 13294
rect 5573 13200 5606 13246
rect 5652 13200 5685 13246
rect 5573 13152 5685 13200
rect 5573 13106 5606 13152
rect 5652 13106 5685 13152
rect 5573 13058 5685 13106
rect 5573 13012 5606 13058
rect 5652 13012 5685 13058
rect 5573 12964 5685 13012
rect 5573 12918 5606 12964
rect 5652 12918 5685 12964
rect 5573 12870 5685 12918
rect 5573 12824 5606 12870
rect 5652 12824 5685 12870
rect 5573 12776 5685 12824
rect 5573 12730 5606 12776
rect 5652 12730 5685 12776
rect 5573 12682 5685 12730
rect 5573 12636 5606 12682
rect 5652 12636 5685 12682
rect 5573 12588 5685 12636
rect 5573 12542 5606 12588
rect 5652 12542 5685 12588
rect 5573 12494 5685 12542
rect 5573 12448 5606 12494
rect 5652 12448 5685 12494
rect 5573 12400 5685 12448
rect 5573 12354 5606 12400
rect 5652 12354 5685 12400
rect 5573 12306 5685 12354
rect 5573 12260 5606 12306
rect 5652 12260 5685 12306
rect 5573 12212 5685 12260
rect 5573 12166 5606 12212
rect 5652 12166 5685 12212
rect 5573 12118 5685 12166
rect 5573 12072 5606 12118
rect 5652 12072 5685 12118
rect 5573 12024 5685 12072
rect 5573 11978 5606 12024
rect 5652 11978 5685 12024
rect 5573 11930 5685 11978
rect 5573 11884 5606 11930
rect 5652 11884 5685 11930
rect 5573 11836 5685 11884
rect 5573 11790 5606 11836
rect 5652 11790 5685 11836
rect 5573 11742 5685 11790
rect 5573 11696 5606 11742
rect 5652 11696 5685 11742
rect 5573 11648 5685 11696
rect 5573 11602 5606 11648
rect 5652 11602 5685 11648
rect 5573 11554 5685 11602
rect 5573 11508 5606 11554
rect 5652 11508 5685 11554
rect 5573 11460 5685 11508
rect 5573 11414 5606 11460
rect 5652 11414 5685 11460
rect 5573 11366 5685 11414
rect 5573 11320 5606 11366
rect 5652 11320 5685 11366
rect 5573 11272 5685 11320
rect 5573 11226 5606 11272
rect 5652 11226 5685 11272
rect 5573 11178 5685 11226
rect 5573 11132 5606 11178
rect 5652 11132 5685 11178
rect 5573 11084 5685 11132
rect 5573 11038 5606 11084
rect 5652 11038 5685 11084
rect 5573 10990 5685 11038
rect 5573 10944 5606 10990
rect 5652 10944 5685 10990
rect 5573 10896 5685 10944
rect 5573 10850 5606 10896
rect 5652 10850 5685 10896
rect 5573 10802 5685 10850
rect 5573 10756 5606 10802
rect 5652 10756 5685 10802
rect 5573 10708 5685 10756
rect 5573 10662 5606 10708
rect 5652 10662 5685 10708
rect 5573 10614 5685 10662
rect 5573 10568 5606 10614
rect 5652 10568 5685 10614
rect 5573 10520 5685 10568
rect 5573 10474 5606 10520
rect 5652 10474 5685 10520
rect 5573 10426 5685 10474
rect 5573 10380 5606 10426
rect 5652 10380 5685 10426
rect 5573 10332 5685 10380
rect 5573 10286 5606 10332
rect 5652 10286 5685 10332
rect 5573 10238 5685 10286
rect 5573 10192 5606 10238
rect 5652 10192 5685 10238
rect 5573 10144 5685 10192
rect 5573 10098 5606 10144
rect 5652 10098 5685 10144
rect 5573 10050 5685 10098
rect 5573 10004 5606 10050
rect 5652 10004 5685 10050
rect 5573 9956 5685 10004
rect 5573 9910 5606 9956
rect 5652 9910 5685 9956
rect 5573 9862 5685 9910
rect 5573 9816 5606 9862
rect 5652 9816 5685 9862
rect 5573 9768 5685 9816
rect 5573 9722 5606 9768
rect 5652 9722 5685 9768
rect 5573 9674 5685 9722
rect 5573 9628 5606 9674
rect 5652 9628 5685 9674
rect 5573 9580 5685 9628
rect 5573 9534 5606 9580
rect 5652 9534 5685 9580
rect 5573 9486 5685 9534
rect 5573 9440 5606 9486
rect 5652 9440 5685 9486
rect 5573 9392 5685 9440
rect 5573 9346 5606 9392
rect 5652 9346 5685 9392
rect 5573 9298 5685 9346
rect 5573 9252 5606 9298
rect 5652 9252 5685 9298
rect 5573 9204 5685 9252
rect 5573 9158 5606 9204
rect 5652 9158 5685 9204
rect 5573 9110 5685 9158
rect 5573 9064 5606 9110
rect 5652 9064 5685 9110
rect 5573 9016 5685 9064
rect 5573 8970 5606 9016
rect 5652 8970 5685 9016
rect 5573 8922 5685 8970
rect 5573 8876 5606 8922
rect 5652 8876 5685 8922
rect 5573 8828 5685 8876
rect 5573 8782 5606 8828
rect 5652 8782 5685 8828
rect 5573 8734 5685 8782
rect 5573 8688 5606 8734
rect 5652 8688 5685 8734
rect 5573 8640 5685 8688
rect 5573 8594 5606 8640
rect 5652 8594 5685 8640
rect 5573 8546 5685 8594
rect 5573 8500 5606 8546
rect 5652 8500 5685 8546
rect 5573 8452 5685 8500
rect 5573 8406 5606 8452
rect 5652 8406 5685 8452
rect 5573 8358 5685 8406
rect 5573 8312 5606 8358
rect 5652 8312 5685 8358
rect 5573 8264 5685 8312
rect 5573 8218 5606 8264
rect 5652 8218 5685 8264
rect 5573 8170 5685 8218
rect 5573 8124 5606 8170
rect 5652 8124 5685 8170
rect 5573 8076 5685 8124
rect 5573 8030 5606 8076
rect 5652 8030 5685 8076
rect 5573 7982 5685 8030
rect 5573 7936 5606 7982
rect 5652 7936 5685 7982
rect 5573 7888 5685 7936
rect 5573 7842 5606 7888
rect 5652 7842 5685 7888
rect 5573 7794 5685 7842
rect 5573 7748 5606 7794
rect 5652 7748 5685 7794
rect 5573 7700 5685 7748
rect 5573 7654 5606 7700
rect 5652 7654 5685 7700
rect 5573 7606 5685 7654
rect 5573 7560 5606 7606
rect 5652 7560 5685 7606
rect 5573 7512 5685 7560
rect 5573 7466 5606 7512
rect 5652 7466 5685 7512
rect 5573 7418 5685 7466
rect 5573 7381 5606 7418
rect 3490 7372 5606 7381
rect 5652 7372 5685 7418
rect 497 7324 5685 7372
rect 497 7278 530 7324
rect 576 7278 624 7324
rect 670 7278 718 7324
rect 764 7278 812 7324
rect 858 7278 906 7324
rect 952 7278 1000 7324
rect 1046 7278 1094 7324
rect 1140 7278 1188 7324
rect 1234 7278 1282 7324
rect 1328 7278 1376 7324
rect 1422 7278 1470 7324
rect 1516 7278 1564 7324
rect 1610 7278 1658 7324
rect 1704 7278 1752 7324
rect 1798 7278 1846 7324
rect 1892 7278 1940 7324
rect 1986 7278 2034 7324
rect 2080 7278 2128 7324
rect 2174 7278 2222 7324
rect 2268 7278 2316 7324
rect 2362 7278 2410 7324
rect 2456 7278 2504 7324
rect 2550 7278 2598 7324
rect 2644 7278 2692 7324
rect 2738 7278 2786 7324
rect 2832 7278 2880 7324
rect 2926 7278 2974 7324
rect 3020 7278 3068 7324
rect 3114 7278 3162 7324
rect 3208 7278 3256 7324
rect 3302 7278 3350 7324
rect 3396 7278 3444 7324
rect 3490 7278 3538 7324
rect 3584 7278 3632 7324
rect 3678 7278 3726 7324
rect 3772 7278 3820 7324
rect 3866 7278 3914 7324
rect 3960 7278 4008 7324
rect 4054 7278 4102 7324
rect 4148 7278 4196 7324
rect 4242 7278 4290 7324
rect 4336 7278 4384 7324
rect 4430 7278 4478 7324
rect 4524 7278 4572 7324
rect 4618 7278 4666 7324
rect 4712 7278 4760 7324
rect 4806 7278 4854 7324
rect 4900 7278 4948 7324
rect 4994 7278 5042 7324
rect 5088 7278 5136 7324
rect 5182 7278 5230 7324
rect 5276 7278 5324 7324
rect 5370 7278 5418 7324
rect 5464 7278 5512 7324
rect 5558 7278 5606 7324
rect 5652 7278 5685 7324
rect 497 7221 5685 7278
rect 6229 13773 6262 13819
rect 6308 13773 6341 13819
rect 6229 13725 6341 13773
rect 6229 13679 6262 13725
rect 6308 13679 6341 13725
rect 6229 13631 6341 13679
rect 6229 13585 6262 13631
rect 6308 13585 6341 13631
rect 6229 13537 6341 13585
rect 6229 13491 6262 13537
rect 6308 13491 6341 13537
rect 6229 13443 6341 13491
rect 6229 13397 6262 13443
rect 6308 13397 6341 13443
rect 6229 13349 6341 13397
rect 6229 13303 6262 13349
rect 6308 13303 6341 13349
rect 6229 13255 6341 13303
rect 6229 13209 6262 13255
rect 6308 13209 6341 13255
rect 6229 13161 6341 13209
rect 6229 13115 6262 13161
rect 6308 13115 6341 13161
rect 6229 13067 6341 13115
rect 6229 13021 6262 13067
rect 6308 13021 6341 13067
rect 6229 12973 6341 13021
rect 6229 12927 6262 12973
rect 6308 12927 6341 12973
rect 6229 12879 6341 12927
rect 6229 12833 6262 12879
rect 6308 12833 6341 12879
rect 6229 12785 6341 12833
rect 6229 12739 6262 12785
rect 6308 12739 6341 12785
rect 6229 12691 6341 12739
rect 6229 12645 6262 12691
rect 6308 12645 6341 12691
rect 6229 12597 6341 12645
rect 6229 12551 6262 12597
rect 6308 12551 6341 12597
rect 6229 12503 6341 12551
rect 6229 12448 6262 12503
rect 6308 12448 6341 12503
rect 6229 12400 6341 12448
rect 6229 12354 6262 12400
rect 6308 12354 6341 12400
rect 6229 12306 6341 12354
rect 6229 12260 6262 12306
rect 6308 12260 6341 12306
rect 6229 12212 6341 12260
rect 6229 12166 6262 12212
rect 6308 12166 6341 12212
rect 6229 12118 6341 12166
rect 6229 12072 6262 12118
rect 6308 12072 6341 12118
rect 6229 12024 6341 12072
rect 6229 11978 6262 12024
rect 6308 11978 6341 12024
rect 6229 11930 6341 11978
rect 6229 11884 6262 11930
rect 6308 11884 6341 11930
rect 6229 11836 6341 11884
rect 6229 11790 6262 11836
rect 6308 11790 6341 11836
rect 6229 11742 6341 11790
rect 6229 11696 6262 11742
rect 6308 11696 6341 11742
rect 6229 11648 6341 11696
rect 6229 11602 6262 11648
rect 6308 11602 6341 11648
rect 6229 11554 6341 11602
rect 6229 11508 6262 11554
rect 6308 11508 6341 11554
rect 6229 11460 6341 11508
rect 6229 11414 6262 11460
rect 6308 11414 6341 11460
rect 6229 11366 6341 11414
rect 6229 11320 6262 11366
rect 6308 11320 6341 11366
rect 6229 11272 6341 11320
rect 6229 11226 6262 11272
rect 6308 11226 6341 11272
rect 6229 11178 6341 11226
rect 6229 11132 6262 11178
rect 6308 11132 6341 11178
rect 6229 11084 6341 11132
rect 6229 11038 6262 11084
rect 6308 11038 6341 11084
rect 6229 10990 6341 11038
rect 6229 10944 6262 10990
rect 6308 10944 6341 10990
rect 6229 10896 6341 10944
rect 6229 10850 6262 10896
rect 6308 10850 6341 10896
rect 6229 10802 6341 10850
rect 6229 10756 6262 10802
rect 6308 10756 6341 10802
rect 6229 10708 6341 10756
rect 6229 10662 6262 10708
rect 6308 10662 6341 10708
rect 6229 10614 6341 10662
rect 6229 10568 6262 10614
rect 6308 10568 6341 10614
rect 6229 10520 6341 10568
rect 6229 10474 6262 10520
rect 6308 10474 6341 10520
rect 6229 10426 6341 10474
rect 6229 10380 6262 10426
rect 6308 10380 6341 10426
rect 6229 10332 6341 10380
rect 6229 10286 6262 10332
rect 6308 10286 6341 10332
rect 6229 10238 6341 10286
rect 6229 10192 6262 10238
rect 6308 10192 6341 10238
rect 6229 10144 6341 10192
rect 6229 10098 6262 10144
rect 6308 10098 6341 10144
rect 6229 10050 6341 10098
rect 6229 10004 6262 10050
rect 6308 10004 6341 10050
rect 6229 9956 6341 10004
rect 6229 9910 6262 9956
rect 6308 9910 6341 9956
rect 6229 9862 6341 9910
rect 6229 9816 6262 9862
rect 6308 9816 6341 9862
rect 6229 9768 6341 9816
rect 6229 9722 6262 9768
rect 6308 9722 6341 9768
rect 6229 9674 6341 9722
rect 6229 9628 6262 9674
rect 6308 9628 6341 9674
rect 6229 9580 6341 9628
rect 6229 9534 6262 9580
rect 6308 9534 6341 9580
rect 6229 9486 6341 9534
rect 6229 9440 6262 9486
rect 6308 9440 6341 9486
rect 6229 9392 6341 9440
rect 6229 9346 6262 9392
rect 6308 9346 6341 9392
rect 6229 9298 6341 9346
rect 6229 9252 6262 9298
rect 6308 9252 6341 9298
rect 6229 9204 6341 9252
rect 6229 9158 6262 9204
rect 6308 9158 6341 9204
rect 6229 9110 6341 9158
rect 6229 9064 6262 9110
rect 6308 9064 6341 9110
rect 6229 9016 6341 9064
rect 6229 8970 6262 9016
rect 6308 8970 6341 9016
rect 6229 8922 6341 8970
rect 6229 8876 6262 8922
rect 6308 8876 6341 8922
rect 6229 8828 6341 8876
rect 6229 8782 6262 8828
rect 6308 8782 6341 8828
rect 6229 8734 6341 8782
rect 6229 8688 6262 8734
rect 6308 8688 6341 8734
rect 6229 8640 6341 8688
rect 6229 8594 6262 8640
rect 6308 8594 6341 8640
rect 6229 8546 6341 8594
rect 6229 8500 6262 8546
rect 6308 8500 6341 8546
rect 6229 8452 6341 8500
rect 6229 8406 6262 8452
rect 6308 8406 6341 8452
rect 6229 8358 6341 8406
rect 6229 8312 6262 8358
rect 6308 8312 6341 8358
rect 6229 8264 6341 8312
rect 6229 8218 6262 8264
rect 6308 8218 6341 8264
rect 6229 8170 6341 8218
rect 6229 8124 6262 8170
rect 6308 8124 6341 8170
rect 6229 8076 6341 8124
rect 6229 8030 6262 8076
rect 6308 8030 6341 8076
rect 6229 7982 6341 8030
rect 6229 7936 6262 7982
rect 6308 7936 6341 7982
rect 6229 7888 6341 7936
rect 6229 7842 6262 7888
rect 6308 7842 6341 7888
rect 6229 7794 6341 7842
rect 6229 7748 6262 7794
rect 6308 7748 6341 7794
rect 6229 7700 6341 7748
rect 6229 7654 6262 7700
rect 6308 7654 6341 7700
rect 6229 7606 6341 7654
rect 6229 7560 6262 7606
rect 6308 7560 6341 7606
rect 6229 7512 6341 7560
rect 6229 7466 6262 7512
rect 6308 7466 6341 7512
rect 6229 7418 6341 7466
rect 6229 7372 6262 7418
rect 6308 7381 6341 7418
rect 6462 14263 6508 14562
rect 6462 13401 6508 13713
rect 6462 12539 6508 12851
rect 6462 11677 6508 11989
rect 6462 10815 6508 11127
rect 6462 9953 6508 10265
rect 6462 9091 6508 9403
rect 6462 8408 6508 8541
rect 6622 14263 6668 14562
rect 6735 14272 6811 14284
rect 6735 14220 6747 14272
rect 6799 14220 6811 14272
rect 6735 14168 6750 14220
rect 6796 14168 6811 14220
rect 6735 14116 6747 14168
rect 6799 14116 6811 14168
rect 6735 14104 6750 14116
rect 6622 13401 6668 13713
rect 6796 14104 6811 14116
rect 6910 14263 6956 14562
rect 6750 13702 6796 13713
rect 7070 14263 7116 14274
rect 7055 13977 7070 13989
rect 7230 14263 7276 14562
rect 7116 13977 7131 13989
rect 7055 13925 7067 13977
rect 7119 13925 7131 13977
rect 7055 13873 7070 13925
rect 7116 13873 7131 13925
rect 7055 13821 7067 13873
rect 7119 13821 7131 13873
rect 7055 13809 7070 13821
rect 6750 13401 6796 13412
rect 6622 12539 6668 12851
rect 6735 12998 6750 13010
rect 6910 13401 6956 13713
rect 7116 13809 7131 13821
rect 7070 13702 7116 13713
rect 7375 14272 7451 14284
rect 7375 14220 7387 14272
rect 7439 14220 7451 14272
rect 7375 14168 7390 14220
rect 7436 14168 7451 14220
rect 7375 14116 7387 14168
rect 7439 14116 7451 14168
rect 7375 14104 7390 14116
rect 6796 12998 6811 13010
rect 6735 12946 6747 12998
rect 6799 12946 6811 12998
rect 6735 12894 6750 12946
rect 6796 12894 6811 12946
rect 6735 12842 6747 12894
rect 6799 12842 6811 12894
rect 6735 12830 6811 12842
rect 7070 13401 7116 13412
rect 7055 13377 7070 13389
rect 7230 13401 7276 13713
rect 7436 14104 7451 14116
rect 7550 14263 7596 14562
rect 7390 13702 7436 13713
rect 7710 14263 7756 14274
rect 7695 13977 7710 13989
rect 7870 14263 7916 14562
rect 7756 13977 7771 13989
rect 7695 13925 7707 13977
rect 7759 13925 7771 13977
rect 7695 13873 7710 13925
rect 7756 13873 7771 13925
rect 7695 13821 7707 13873
rect 7759 13821 7771 13873
rect 7695 13809 7710 13821
rect 7116 13377 7131 13389
rect 7055 13325 7067 13377
rect 7119 13325 7131 13377
rect 7055 13273 7070 13325
rect 7116 13273 7131 13325
rect 7055 13221 7067 13273
rect 7119 13221 7131 13273
rect 7055 13209 7070 13221
rect 6750 12539 6796 12550
rect 6622 11677 6668 11989
rect 6735 12136 6750 12148
rect 6910 12539 6956 12851
rect 7116 13209 7131 13221
rect 7070 12840 7116 12851
rect 7390 13401 7436 13412
rect 6796 12136 6811 12148
rect 6735 12084 6747 12136
rect 6799 12084 6811 12136
rect 6735 12032 6750 12084
rect 6796 12032 6811 12084
rect 6735 11980 6747 12032
rect 6799 11980 6811 12032
rect 6735 11968 6811 11980
rect 7070 12539 7116 12550
rect 7055 12455 7070 12467
rect 7230 12539 7276 12851
rect 7375 12998 7390 13010
rect 7550 13401 7596 13713
rect 7756 13809 7771 13821
rect 7710 13702 7756 13713
rect 8015 14272 8091 14284
rect 8015 14220 8027 14272
rect 8079 14220 8091 14272
rect 8015 14168 8030 14220
rect 8076 14168 8091 14220
rect 8015 14116 8027 14168
rect 8079 14116 8091 14168
rect 8015 14104 8030 14116
rect 7436 12998 7451 13010
rect 7375 12946 7387 12998
rect 7439 12946 7451 12998
rect 7375 12894 7390 12946
rect 7436 12894 7451 12946
rect 7375 12842 7387 12894
rect 7439 12842 7451 12894
rect 7375 12830 7451 12842
rect 7710 13401 7756 13412
rect 7695 13377 7710 13389
rect 7870 13401 7916 13713
rect 8076 14104 8091 14116
rect 8158 14263 8204 14562
rect 8030 13702 8076 13713
rect 7756 13377 7771 13389
rect 7695 13325 7707 13377
rect 7759 13325 7771 13377
rect 7695 13273 7710 13325
rect 7756 13273 7771 13325
rect 7695 13221 7707 13273
rect 7759 13221 7771 13273
rect 7695 13209 7710 13221
rect 7116 12455 7131 12467
rect 7055 12403 7067 12455
rect 7119 12403 7131 12455
rect 7055 12351 7070 12403
rect 7116 12351 7131 12403
rect 7055 12299 7067 12351
rect 7119 12299 7131 12351
rect 7055 12287 7070 12299
rect 6750 11677 6796 11688
rect 6735 11613 6750 11625
rect 6910 11677 6956 11989
rect 7116 12287 7131 12299
rect 7070 11978 7116 11989
rect 7390 12539 7436 12550
rect 6796 11613 6811 11625
rect 6735 11561 6747 11613
rect 6799 11561 6811 11613
rect 6735 11509 6750 11561
rect 6796 11509 6811 11561
rect 6735 11457 6747 11509
rect 6799 11457 6811 11509
rect 6735 11445 6750 11457
rect 6622 10815 6668 11127
rect 6622 9953 6668 10265
rect 6796 11445 6811 11457
rect 6750 10815 6796 11127
rect 6750 10254 6796 10265
rect 7070 11677 7116 11688
rect 7055 11325 7070 11337
rect 7230 11677 7276 11989
rect 7375 12136 7390 12148
rect 7550 12539 7596 12851
rect 7756 13209 7771 13221
rect 7710 12840 7756 12851
rect 8030 13401 8076 13412
rect 7436 12136 7451 12148
rect 7375 12084 7387 12136
rect 7439 12084 7451 12136
rect 7375 12032 7390 12084
rect 7436 12032 7451 12084
rect 7375 11980 7387 12032
rect 7439 11980 7451 12032
rect 7375 11968 7451 11980
rect 7710 12539 7756 12550
rect 7695 12455 7710 12467
rect 7870 12539 7916 12851
rect 8015 12998 8030 13010
rect 8158 13401 8204 13713
rect 8076 12998 8091 13010
rect 8015 12946 8027 12998
rect 8079 12946 8091 12998
rect 8015 12894 8030 12946
rect 8076 12894 8091 12946
rect 8015 12842 8027 12894
rect 8079 12842 8091 12894
rect 8015 12830 8091 12842
rect 7756 12455 7771 12467
rect 7695 12403 7707 12455
rect 7759 12403 7771 12455
rect 7695 12351 7710 12403
rect 7756 12351 7771 12403
rect 7695 12299 7707 12351
rect 7759 12299 7771 12351
rect 7695 12287 7710 12299
rect 7116 11325 7131 11337
rect 7055 11273 7067 11325
rect 7119 11273 7131 11325
rect 7055 11221 7070 11273
rect 7116 11221 7131 11273
rect 7055 11169 7067 11221
rect 7119 11169 7131 11221
rect 7055 11157 7070 11169
rect 6910 10815 6956 11127
rect 6750 9953 6796 9964
rect 6622 9091 6668 9403
rect 6735 9561 6750 9573
rect 6910 9953 6956 10265
rect 7116 11157 7131 11169
rect 7070 10815 7116 11127
rect 7070 10254 7116 10265
rect 7390 11677 7436 11688
rect 7375 11613 7390 11625
rect 7550 11677 7596 11989
rect 7756 12287 7771 12299
rect 7710 11978 7756 11989
rect 8030 12539 8076 12550
rect 7436 11613 7451 11625
rect 7375 11561 7387 11613
rect 7439 11561 7451 11613
rect 7375 11509 7390 11561
rect 7436 11509 7451 11561
rect 7375 11457 7387 11509
rect 7439 11457 7451 11509
rect 7375 11445 7390 11457
rect 7230 10815 7276 11127
rect 6796 9561 6811 9573
rect 6735 9509 6747 9561
rect 6799 9509 6811 9561
rect 6735 9457 6750 9509
rect 6796 9457 6811 9509
rect 6735 9405 6747 9457
rect 6799 9405 6811 9457
rect 6735 9403 6750 9405
rect 6796 9403 6811 9405
rect 6735 9393 6811 9403
rect 7055 9962 7131 9974
rect 7055 9910 7067 9962
rect 7119 9910 7131 9962
rect 7055 9858 7070 9910
rect 7116 9858 7131 9910
rect 7055 9806 7067 9858
rect 7119 9806 7131 9858
rect 7055 9794 7070 9806
rect 6750 9392 6796 9393
rect 6750 9091 6796 9102
rect 6735 8961 6750 8973
rect 6910 9091 6956 9403
rect 7116 9794 7131 9806
rect 7230 9953 7276 10265
rect 7436 11445 7451 11457
rect 7390 10815 7436 11127
rect 7390 10254 7436 10265
rect 7710 11677 7756 11688
rect 7695 11325 7710 11337
rect 7870 11677 7916 11989
rect 8015 12136 8030 12148
rect 8158 12539 8204 12851
rect 8076 12136 8091 12148
rect 8015 12084 8027 12136
rect 8079 12084 8091 12136
rect 8015 12032 8030 12084
rect 8076 12032 8091 12084
rect 8015 11980 8027 12032
rect 8079 11980 8091 12032
rect 8015 11968 8091 11980
rect 7756 11325 7771 11337
rect 7695 11273 7707 11325
rect 7759 11273 7771 11325
rect 7695 11221 7710 11273
rect 7756 11221 7771 11273
rect 7695 11169 7707 11221
rect 7759 11169 7771 11221
rect 7695 11157 7710 11169
rect 7550 10815 7596 11127
rect 7070 9392 7116 9403
rect 7390 9953 7436 9964
rect 6796 8961 6811 8973
rect 6735 8909 6747 8961
rect 6799 8909 6811 8961
rect 6735 8857 6750 8909
rect 6796 8857 6811 8909
rect 6735 8805 6747 8857
rect 6799 8805 6811 8857
rect 6735 8793 6750 8805
rect 6622 8408 6668 8541
rect 6796 8793 6811 8805
rect 6750 8530 6796 8541
rect 7070 9091 7116 9102
rect 6462 8362 6542 8408
rect 6588 8362 6668 8408
rect 6462 8229 6508 8362
rect 6462 7381 6508 7679
rect 6622 8229 6668 8362
rect 6750 8229 6796 8240
rect 6622 7381 6668 7679
rect 6735 7831 6750 7843
rect 6910 8229 6956 8541
rect 7055 8688 7070 8700
rect 7230 9091 7276 9403
rect 7375 9561 7390 9573
rect 7550 9953 7596 10265
rect 7756 11157 7771 11169
rect 7710 10815 7756 11127
rect 7710 10254 7756 10265
rect 8030 11677 8076 11688
rect 8015 11613 8030 11625
rect 8158 11677 8204 11989
rect 8076 11613 8091 11625
rect 8015 11561 8027 11613
rect 8079 11561 8091 11613
rect 8015 11509 8030 11561
rect 8076 11509 8091 11561
rect 8015 11457 8027 11509
rect 8079 11457 8091 11509
rect 8015 11445 8030 11457
rect 7870 10815 7916 11127
rect 7436 9561 7451 9573
rect 7375 9509 7387 9561
rect 7439 9509 7451 9561
rect 7375 9457 7390 9509
rect 7436 9457 7451 9509
rect 7375 9405 7387 9457
rect 7439 9405 7451 9457
rect 7375 9403 7390 9405
rect 7436 9403 7451 9405
rect 7375 9393 7451 9403
rect 7695 9962 7771 9974
rect 7695 9910 7707 9962
rect 7759 9910 7771 9962
rect 7695 9858 7710 9910
rect 7756 9858 7771 9910
rect 7695 9806 7707 9858
rect 7759 9806 7771 9858
rect 7695 9794 7710 9806
rect 7390 9392 7436 9393
rect 7116 8688 7131 8700
rect 7055 8636 7067 8688
rect 7119 8636 7131 8688
rect 7055 8584 7070 8636
rect 7116 8584 7131 8636
rect 7055 8532 7067 8584
rect 7119 8532 7131 8584
rect 7055 8520 7131 8532
rect 7390 9091 7436 9102
rect 7375 8961 7390 8973
rect 7550 9091 7596 9403
rect 7756 9794 7771 9806
rect 7870 9953 7916 10265
rect 8076 11445 8091 11457
rect 8030 10815 8076 11127
rect 8030 10254 8076 10265
rect 8158 10815 8204 11127
rect 7710 9392 7756 9403
rect 8030 9953 8076 9964
rect 7436 8961 7451 8973
rect 7375 8909 7387 8961
rect 7439 8909 7451 8961
rect 7375 8857 7390 8909
rect 7436 8857 7451 8909
rect 7375 8805 7387 8857
rect 7439 8805 7451 8857
rect 7375 8793 7390 8805
rect 7070 8235 7116 8240
rect 6796 7831 6811 7843
rect 6735 7779 6747 7831
rect 6799 7779 6811 7831
rect 6735 7727 6750 7779
rect 6796 7727 6811 7779
rect 6735 7675 6747 7727
rect 6799 7675 6811 7727
rect 6735 7663 6811 7675
rect 7055 8229 7131 8235
rect 7055 8223 7070 8229
rect 7116 8223 7131 8229
rect 7055 8171 7067 8223
rect 7119 8171 7131 8223
rect 7055 8119 7070 8171
rect 7116 8119 7131 8171
rect 7055 8067 7067 8119
rect 7119 8067 7131 8119
rect 7055 8055 7070 8067
rect 6910 7391 6956 7679
rect 7116 8055 7131 8067
rect 7230 8229 7276 8541
rect 7436 8793 7451 8805
rect 7390 8530 7436 8541
rect 7710 9091 7756 9102
rect 7070 7668 7116 7679
rect 7390 8229 7436 8240
rect 6867 7381 7047 7391
rect 7230 7381 7276 7679
rect 7375 7831 7390 7843
rect 7550 8229 7596 8541
rect 7695 8688 7710 8700
rect 7870 9091 7916 9403
rect 8015 9561 8030 9573
rect 8158 9953 8204 10265
rect 8076 9561 8091 9573
rect 8015 9509 8027 9561
rect 8079 9509 8091 9561
rect 8015 9457 8030 9509
rect 8076 9457 8091 9509
rect 8015 9405 8027 9457
rect 8079 9405 8091 9457
rect 8015 9403 8030 9405
rect 8076 9403 8091 9405
rect 8015 9393 8091 9403
rect 8030 9392 8076 9393
rect 7756 8688 7771 8700
rect 7695 8636 7707 8688
rect 7759 8636 7771 8688
rect 7695 8584 7710 8636
rect 7756 8584 7771 8636
rect 7695 8532 7707 8584
rect 7759 8532 7771 8584
rect 7695 8520 7771 8532
rect 8030 9091 8076 9102
rect 8015 8961 8030 8973
rect 8158 9091 8204 9403
rect 8076 8961 8091 8973
rect 8015 8909 8027 8961
rect 8079 8909 8091 8961
rect 8015 8857 8030 8909
rect 8076 8857 8091 8909
rect 8015 8805 8027 8857
rect 8079 8805 8091 8857
rect 8015 8793 8030 8805
rect 7710 8235 7756 8240
rect 7436 7831 7451 7843
rect 7375 7779 7387 7831
rect 7439 7779 7451 7831
rect 7375 7727 7390 7779
rect 7436 7727 7451 7779
rect 7375 7675 7387 7727
rect 7439 7675 7451 7727
rect 7375 7663 7451 7675
rect 7695 8229 7771 8235
rect 7695 8223 7710 8229
rect 7756 8223 7771 8229
rect 7695 8171 7707 8223
rect 7759 8171 7771 8223
rect 7695 8119 7710 8171
rect 7756 8119 7771 8171
rect 7695 8067 7707 8119
rect 7759 8067 7771 8119
rect 7695 8055 7710 8067
rect 7550 7381 7596 7679
rect 7756 8055 7771 8067
rect 7870 8229 7916 8541
rect 8076 8793 8091 8805
rect 8030 8530 8076 8541
rect 7989 8464 8065 8476
rect 7989 8412 8001 8464
rect 8053 8412 8065 8464
rect 7989 8360 8065 8412
rect 7989 8308 8001 8360
rect 8053 8308 8065 8360
rect 7989 8296 8065 8308
rect 8158 8408 8204 8541
rect 8318 14263 8364 14562
rect 8318 13401 8364 13713
rect 8318 12539 8364 12851
rect 8318 11677 8364 11989
rect 8318 10815 8364 11127
rect 8318 9953 8364 10265
rect 8318 9091 8364 9403
rect 8318 8408 8364 8541
rect 8158 8362 8238 8408
rect 8284 8362 8364 8408
rect 7710 7668 7756 7679
rect 8030 8229 8076 8240
rect 7870 7381 7916 7679
rect 8015 7831 8030 7843
rect 8158 8229 8204 8362
rect 8076 7831 8091 7843
rect 8015 7779 8027 7831
rect 8079 7779 8091 7831
rect 8015 7727 8030 7779
rect 8076 7727 8091 7779
rect 8015 7675 8027 7727
rect 8079 7675 8091 7727
rect 8015 7663 8091 7675
rect 8158 7381 8204 7679
rect 8318 8229 8364 8362
rect 8318 7381 8364 7679
rect 8485 14525 8518 14562
rect 8564 14525 30392 14571
rect 8485 14477 30392 14525
rect 8485 14431 8518 14477
rect 8564 14431 30392 14477
rect 8485 14402 30392 14431
rect 8485 14383 8645 14402
rect 8485 14337 8518 14383
rect 8564 14337 8645 14383
rect 8485 14289 8645 14337
rect 8485 14243 8518 14289
rect 8564 14243 8645 14289
rect 8485 14195 8645 14243
rect 8485 14149 8518 14195
rect 8564 14149 8645 14195
rect 8485 14101 8645 14149
rect 8485 14055 8518 14101
rect 8564 14055 8645 14101
rect 8485 14007 8645 14055
rect 8485 13961 8518 14007
rect 8564 13961 8645 14007
rect 8485 13913 8645 13961
rect 8485 13867 8518 13913
rect 8564 13877 8645 13913
rect 9153 13877 9313 14402
rect 9858 13877 10018 14402
rect 10672 13877 10832 14402
rect 15658 14393 17304 14402
rect 22013 13877 22333 14402
rect 26650 13877 26970 14402
rect 30072 13877 30392 14402
rect 37919 14237 39343 14244
rect 8564 13867 30392 13877
rect 8485 13819 30392 13867
rect 8485 13773 8518 13819
rect 8564 13773 30392 13819
rect 8485 13768 30392 13773
rect 8485 13725 18136 13768
rect 8485 13679 8518 13725
rect 8564 13722 18136 13725
rect 18182 13722 18230 13768
rect 18276 13722 18324 13768
rect 18370 13722 18418 13768
rect 18464 13722 18512 13768
rect 18558 13722 18606 13768
rect 18652 13722 18700 13768
rect 18746 13722 18794 13768
rect 18840 13722 18888 13768
rect 18934 13722 18982 13768
rect 19028 13722 19076 13768
rect 19122 13722 19170 13768
rect 19216 13722 19264 13768
rect 19310 13722 19358 13768
rect 19404 13722 19452 13768
rect 19498 13722 19546 13768
rect 19592 13722 19640 13768
rect 19686 13722 19734 13768
rect 19780 13722 19828 13768
rect 19874 13722 19922 13768
rect 19968 13722 20016 13768
rect 20062 13722 20110 13768
rect 20156 13722 20204 13768
rect 20250 13722 20298 13768
rect 20344 13722 20392 13768
rect 20438 13722 20486 13768
rect 20532 13722 20580 13768
rect 20626 13722 20674 13768
rect 20720 13722 20768 13768
rect 20814 13722 20862 13768
rect 20908 13722 20956 13768
rect 21002 13722 21050 13768
rect 21096 13722 21144 13768
rect 21190 13722 23288 13768
rect 23334 13722 23382 13768
rect 23428 13722 23476 13768
rect 23522 13722 23570 13768
rect 23616 13722 23664 13768
rect 23710 13722 23758 13768
rect 23804 13722 23852 13768
rect 23898 13722 23946 13768
rect 23992 13722 24040 13768
rect 24086 13722 24134 13768
rect 24180 13722 24228 13768
rect 24274 13722 24322 13768
rect 24368 13722 24416 13768
rect 24462 13722 24510 13768
rect 24556 13722 24604 13768
rect 24650 13722 24698 13768
rect 24744 13722 24792 13768
rect 24838 13722 24886 13768
rect 24932 13722 24980 13768
rect 25026 13722 25074 13768
rect 25120 13722 25168 13768
rect 25214 13722 25262 13768
rect 25308 13722 25356 13768
rect 25402 13722 25450 13768
rect 25496 13722 25544 13768
rect 25590 13722 25638 13768
rect 25684 13722 25732 13768
rect 25778 13722 25826 13768
rect 25872 13722 25920 13768
rect 25966 13722 26014 13768
rect 26060 13722 26108 13768
rect 26154 13722 26202 13768
rect 26248 13722 26296 13768
rect 26342 13722 27257 13768
rect 27303 13722 27351 13768
rect 27397 13722 27445 13768
rect 27491 13722 27539 13768
rect 27585 13722 27633 13768
rect 27679 13722 27727 13768
rect 27773 13722 27821 13768
rect 27867 13722 27915 13768
rect 27961 13722 28009 13768
rect 28055 13722 28103 13768
rect 28149 13722 28197 13768
rect 28243 13722 28291 13768
rect 28337 13722 28385 13768
rect 28431 13722 28479 13768
rect 28525 13722 28573 13768
rect 28619 13722 28667 13768
rect 28713 13722 28761 13768
rect 28807 13722 28855 13768
rect 28901 13722 28949 13768
rect 28995 13722 29043 13768
rect 29089 13722 29137 13768
rect 29183 13722 29231 13768
rect 29277 13722 29325 13768
rect 29371 13722 29419 13768
rect 29465 13722 29513 13768
rect 29559 13722 29607 13768
rect 29653 13722 29701 13768
rect 29747 13722 29795 13768
rect 29841 13722 29889 13768
rect 29935 13722 29983 13768
rect 30029 13722 30077 13768
rect 30123 13722 30171 13768
rect 30217 13722 30265 13768
rect 30311 13722 30392 13768
rect 8564 13679 30392 13722
rect 8485 13674 30392 13679
rect 8485 13631 18136 13674
rect 8485 13585 8518 13631
rect 8564 13628 18136 13631
rect 18182 13628 21144 13674
rect 21190 13628 23288 13674
rect 23334 13628 26296 13674
rect 26342 13628 27257 13674
rect 27303 13628 30265 13674
rect 30311 13628 30392 13674
rect 8564 13585 30392 13628
rect 8485 13580 30392 13585
rect 8485 13557 18136 13580
rect 8485 13537 8645 13557
rect 8485 13491 8518 13537
rect 8564 13491 8645 13537
rect 8485 13443 8645 13491
rect 8485 13397 8518 13443
rect 8564 13397 8645 13443
rect 8485 13349 8645 13397
rect 8485 13303 8518 13349
rect 8564 13303 8645 13349
rect 8485 13255 8645 13303
rect 8485 13209 8518 13255
rect 8564 13209 8645 13255
rect 8485 13161 8645 13209
rect 8485 13115 8518 13161
rect 8564 13115 8645 13161
rect 8485 13077 8645 13115
rect 9153 13077 9313 13557
rect 9858 13077 10018 13557
rect 10672 13077 10832 13557
rect 18055 13534 18136 13557
rect 18182 13557 21144 13580
rect 18182 13534 18375 13557
rect 18055 13486 18375 13534
rect 18055 13440 18136 13486
rect 18182 13440 18375 13486
rect 18055 13392 18375 13440
rect 18055 13346 18136 13392
rect 18182 13346 18375 13392
rect 18055 13298 18375 13346
rect 18055 13252 18136 13298
rect 18182 13252 18375 13298
rect 18055 13204 18375 13252
rect 18055 13158 18136 13204
rect 18182 13158 18375 13204
rect 18055 13110 18375 13158
rect 18055 13077 18136 13110
rect 8485 13067 18136 13077
rect 8485 13021 8518 13067
rect 8564 13064 18136 13067
rect 18182 13064 18375 13110
rect 8564 13021 18375 13064
rect 8485 13016 18375 13021
rect 8485 12973 18136 13016
rect 8485 12927 8518 12973
rect 8564 12970 18136 12973
rect 18182 12970 18375 13016
rect 8564 12927 18375 12970
rect 8485 12922 18375 12927
rect 8485 12879 18136 12922
rect 8485 12833 8518 12879
rect 8564 12876 18136 12879
rect 18182 12876 18375 12922
rect 8564 12833 18375 12876
rect 8485 12828 18375 12833
rect 8485 12785 18136 12828
rect 8485 12739 8518 12785
rect 8564 12782 18136 12785
rect 18182 12782 18375 12828
rect 8564 12757 18375 12782
rect 8564 12739 8645 12757
rect 8485 12691 8645 12739
rect 8485 12645 8518 12691
rect 8564 12645 8645 12691
rect 8485 12597 8645 12645
rect 8485 12551 8518 12597
rect 8564 12551 8645 12597
rect 8485 12503 8645 12551
rect 8485 12448 8518 12503
rect 8564 12448 8645 12503
rect 8485 12400 8645 12448
rect 8485 12354 8518 12400
rect 8564 12354 8645 12400
rect 8485 12306 8645 12354
rect 8485 12260 8518 12306
rect 8564 12260 8645 12306
rect 8485 12212 8645 12260
rect 8485 12166 8518 12212
rect 8564 12166 8645 12212
rect 8485 12118 8645 12166
rect 8485 12072 8518 12118
rect 8564 12072 8645 12118
rect 8485 12024 8645 12072
rect 8485 11978 8518 12024
rect 8564 11978 8645 12024
rect 8485 11930 8645 11978
rect 8485 11884 8518 11930
rect 8564 11884 8645 11930
rect 8485 11836 8645 11884
rect 8485 11790 8518 11836
rect 8564 11790 8645 11836
rect 8485 11742 8645 11790
rect 8485 11696 8518 11742
rect 8564 11696 8645 11742
rect 8485 11648 8645 11696
rect 8485 11602 8518 11648
rect 8564 11602 8645 11648
rect 8485 11554 8645 11602
rect 8485 11508 8518 11554
rect 8564 11508 8645 11554
rect 8485 11460 8645 11508
rect 8485 11414 8518 11460
rect 8564 11414 8645 11460
rect 8485 11366 8645 11414
rect 8485 11320 8518 11366
rect 8564 11320 8645 11366
rect 8485 11272 8645 11320
rect 8485 11226 8518 11272
rect 8564 11235 8645 11272
rect 9153 11235 9313 12757
rect 9858 11235 10018 12757
rect 10672 11235 10832 12757
rect 18055 12734 18375 12757
rect 18055 12688 18136 12734
rect 18182 12688 18375 12734
rect 18055 12640 18375 12688
rect 18055 12594 18136 12640
rect 18182 12594 18375 12640
rect 18055 12546 18375 12594
rect 18055 12500 18136 12546
rect 18182 12500 18375 12546
rect 18055 12452 18375 12500
rect 18055 12406 18136 12452
rect 18182 12406 18375 12452
rect 18055 12358 18375 12406
rect 18055 12312 18136 12358
rect 18182 12312 18375 12358
rect 18055 12264 18375 12312
rect 18055 12218 18136 12264
rect 18182 12218 18375 12264
rect 18055 12170 18375 12218
rect 18055 12124 18136 12170
rect 18182 12124 18375 12170
rect 18055 12076 18375 12124
rect 18055 12030 18136 12076
rect 18182 12030 18375 12076
rect 18055 11982 18375 12030
rect 18055 11936 18136 11982
rect 18182 11936 18375 11982
rect 18055 11888 18375 11936
rect 18055 11842 18136 11888
rect 18182 11842 18375 11888
rect 11867 11742 17055 11799
rect 11867 11696 11900 11742
rect 11946 11696 11994 11742
rect 12040 11696 12088 11742
rect 12134 11696 12182 11742
rect 12228 11696 12276 11742
rect 12322 11696 12370 11742
rect 12416 11696 12464 11742
rect 12510 11696 12558 11742
rect 12604 11696 12652 11742
rect 12698 11696 12746 11742
rect 12792 11696 12840 11742
rect 12886 11696 12934 11742
rect 12980 11696 13028 11742
rect 13074 11696 13122 11742
rect 13168 11696 13216 11742
rect 13262 11696 13310 11742
rect 13356 11696 13404 11742
rect 13450 11696 13498 11742
rect 13544 11696 13592 11742
rect 13638 11696 13686 11742
rect 13732 11696 13780 11742
rect 13826 11696 13874 11742
rect 13920 11696 13968 11742
rect 14014 11696 14062 11742
rect 14108 11696 14156 11742
rect 14202 11696 14250 11742
rect 14296 11696 14344 11742
rect 14390 11696 14438 11742
rect 14484 11696 14532 11742
rect 14578 11696 14626 11742
rect 14672 11696 14720 11742
rect 14766 11696 14814 11742
rect 14860 11696 14908 11742
rect 14954 11696 15002 11742
rect 15048 11696 15096 11742
rect 15142 11696 15190 11742
rect 15236 11696 15284 11742
rect 15330 11696 15378 11742
rect 15424 11696 15472 11742
rect 15518 11696 15566 11742
rect 15612 11696 15660 11742
rect 15706 11696 15754 11742
rect 15800 11696 15848 11742
rect 15894 11696 15942 11742
rect 15988 11696 16036 11742
rect 16082 11696 16130 11742
rect 16176 11696 16224 11742
rect 16270 11696 16318 11742
rect 16364 11696 16412 11742
rect 16458 11696 16506 11742
rect 16552 11696 16600 11742
rect 16646 11696 16694 11742
rect 16740 11696 16788 11742
rect 16834 11696 16882 11742
rect 16928 11696 16976 11742
rect 17022 11696 17055 11742
rect 11381 11385 11541 11675
rect 11371 11373 11551 11385
rect 11371 11321 11383 11373
rect 11435 11321 11487 11373
rect 11539 11321 11551 11373
rect 11371 11269 11551 11321
rect 8564 11226 11323 11235
rect 8485 11178 11323 11226
rect 11371 11217 11383 11269
rect 11435 11217 11487 11269
rect 11539 11217 11551 11269
rect 11371 11205 11551 11217
rect 8485 11132 8518 11178
rect 8564 11132 8612 11178
rect 8658 11132 8706 11178
rect 8752 11132 8800 11178
rect 8846 11132 8894 11178
rect 8940 11132 8988 11178
rect 9034 11132 9082 11178
rect 9128 11132 9176 11178
rect 9222 11132 9270 11178
rect 9316 11132 9364 11178
rect 9410 11132 9458 11178
rect 9504 11132 9552 11178
rect 9598 11132 9646 11178
rect 9692 11132 9740 11178
rect 9786 11132 9834 11178
rect 9880 11132 9928 11178
rect 9974 11132 10022 11178
rect 10068 11132 10116 11178
rect 10162 11132 10210 11178
rect 10256 11132 10304 11178
rect 10350 11132 10398 11178
rect 10444 11132 10492 11178
rect 10538 11132 10586 11178
rect 10632 11132 10680 11178
rect 10726 11132 10774 11178
rect 10820 11132 10868 11178
rect 10914 11132 10962 11178
rect 11008 11132 11056 11178
rect 11102 11132 11150 11178
rect 11196 11132 11244 11178
rect 11290 11132 11323 11178
rect 8485 11084 11323 11132
rect 8485 11038 8518 11084
rect 8564 11075 11244 11084
rect 8564 11038 8597 11075
rect 8485 10990 8597 11038
rect 8485 10944 8518 10990
rect 8564 10944 8597 10990
rect 8485 10896 8597 10944
rect 8485 10850 8518 10896
rect 8564 10850 8597 10896
rect 8485 10802 8597 10850
rect 8485 10756 8518 10802
rect 8564 10756 8597 10802
rect 8485 10708 8597 10756
rect 8485 10662 8518 10708
rect 8564 10662 8597 10708
rect 8485 10614 8597 10662
rect 8485 10568 8518 10614
rect 8564 10568 8597 10614
rect 8485 10520 8597 10568
rect 8485 10474 8518 10520
rect 8564 10474 8597 10520
rect 8485 10426 8597 10474
rect 8485 10380 8518 10426
rect 8564 10380 8597 10426
rect 8485 10332 8597 10380
rect 8485 10286 8518 10332
rect 8564 10286 8597 10332
rect 8485 10238 8597 10286
rect 8485 10192 8518 10238
rect 8564 10192 8597 10238
rect 8485 10144 8597 10192
rect 8485 10098 8518 10144
rect 8564 10098 8597 10144
rect 8485 10050 8597 10098
rect 8485 10004 8518 10050
rect 8564 10004 8597 10050
rect 8485 9956 8597 10004
rect 8485 9910 8518 9956
rect 8564 9910 8597 9956
rect 8485 9862 8597 9910
rect 8485 9816 8518 9862
rect 8564 9816 8597 9862
rect 8485 9768 8597 9816
rect 8485 9722 8518 9768
rect 8564 9722 8597 9768
rect 8485 9674 8597 9722
rect 8485 9628 8518 9674
rect 8564 9628 8597 9674
rect 8485 9580 8597 9628
rect 8485 9534 8518 9580
rect 8564 9534 8597 9580
rect 8485 9486 8597 9534
rect 8485 9440 8518 9486
rect 8564 9440 8597 9486
rect 8485 9392 8597 9440
rect 8485 9346 8518 9392
rect 8564 9346 8597 9392
rect 8485 9298 8597 9346
rect 8485 9252 8518 9298
rect 8564 9252 8597 9298
rect 8485 9204 8597 9252
rect 8485 9158 8518 9204
rect 8564 9158 8597 9204
rect 8485 9110 8597 9158
rect 8485 9064 8518 9110
rect 8564 9064 8597 9110
rect 8485 9016 8597 9064
rect 8485 8970 8518 9016
rect 8564 8970 8597 9016
rect 8485 8922 8597 8970
rect 8485 8876 8518 8922
rect 8564 8876 8597 8922
rect 8485 8828 8597 8876
rect 8485 8782 8518 8828
rect 8564 8782 8597 8828
rect 8485 8734 8597 8782
rect 8485 8688 8518 8734
rect 8564 8688 8597 8734
rect 8485 8640 8597 8688
rect 8485 8594 8518 8640
rect 8564 8594 8597 8640
rect 8485 8546 8597 8594
rect 8485 8500 8518 8546
rect 8564 8500 8597 8546
rect 8485 8452 8597 8500
rect 8485 8406 8518 8452
rect 8564 8406 8597 8452
rect 8485 8358 8597 8406
rect 8485 8312 8518 8358
rect 8564 8312 8597 8358
rect 8485 8264 8597 8312
rect 8485 8218 8518 8264
rect 8564 8218 8597 8264
rect 8485 8170 8597 8218
rect 8485 8124 8518 8170
rect 8564 8124 8597 8170
rect 8485 8076 8597 8124
rect 8485 8030 8518 8076
rect 8564 8030 8597 8076
rect 8485 7982 8597 8030
rect 8485 7936 8518 7982
rect 8564 7936 8597 7982
rect 8485 7888 8597 7936
rect 8485 7842 8518 7888
rect 8564 7842 8597 7888
rect 8485 7794 8597 7842
rect 8485 7748 8518 7794
rect 8564 7748 8597 7794
rect 8485 7700 8597 7748
rect 8485 7654 8518 7700
rect 8564 7654 8597 7700
rect 8485 7606 8597 7654
rect 8485 7560 8518 7606
rect 8564 7560 8597 7606
rect 8485 7512 8597 7560
rect 8485 7466 8518 7512
rect 8564 7466 8597 7512
rect 8485 7418 8597 7466
rect 8485 7381 8518 7418
rect 6308 7379 8518 7381
rect 6308 7372 6879 7379
rect 6229 7327 6879 7372
rect 6931 7327 6983 7379
rect 7035 7372 8518 7379
rect 8564 7381 8597 7418
rect 8697 10796 8743 11075
rect 8697 9934 8743 10246
rect 8697 9072 8743 9384
rect 8697 8389 8743 8522
rect 8857 10796 8903 11075
rect 9145 10853 10663 10899
rect 8985 10806 9031 10807
rect 8970 10796 9046 10806
rect 8970 10794 8985 10796
rect 9031 10794 9046 10796
rect 8970 10742 8982 10794
rect 9034 10742 9046 10794
rect 8970 10690 8985 10742
rect 9031 10690 9046 10742
rect 8970 10638 8982 10690
rect 9034 10638 9046 10690
rect 8970 10626 8985 10638
rect 8857 9934 8903 10246
rect 9031 10626 9046 10638
rect 9145 10796 9191 10853
rect 8985 10235 9031 10246
rect 9145 10235 9191 10246
rect 9273 10796 9319 10807
rect 9433 10796 9479 10807
rect 9418 10423 9433 10435
rect 9593 10796 9639 10807
rect 9479 10423 9494 10435
rect 9418 10371 9430 10423
rect 9482 10371 9494 10423
rect 9418 10319 9433 10371
rect 9479 10319 9494 10371
rect 9418 10267 9430 10319
rect 9482 10267 9494 10319
rect 9418 10255 9433 10267
rect 9273 10189 9319 10246
rect 9479 10255 9494 10267
rect 9433 10235 9479 10246
rect 9593 10189 9639 10246
rect 9721 10796 9767 10853
rect 9881 10806 9927 10807
rect 9866 10796 9942 10806
rect 9866 10794 9881 10796
rect 9927 10794 9942 10796
rect 9866 10742 9878 10794
rect 9930 10742 9942 10794
rect 9866 10690 9881 10742
rect 9927 10690 9942 10742
rect 9866 10638 9878 10690
rect 9930 10638 9942 10690
rect 9866 10626 9881 10638
rect 9721 10235 9767 10246
rect 9927 10626 9942 10638
rect 10041 10796 10087 10853
rect 9881 10235 9927 10246
rect 10041 10235 10087 10246
rect 10169 10796 10215 10807
rect 10329 10796 10375 10807
rect 10314 10423 10329 10435
rect 10489 10796 10535 10807
rect 10375 10423 10390 10435
rect 10314 10371 10326 10423
rect 10378 10371 10390 10423
rect 10314 10319 10329 10371
rect 10375 10319 10390 10371
rect 10314 10267 10326 10319
rect 10378 10267 10390 10319
rect 10314 10255 10329 10267
rect 10169 10189 10215 10246
rect 10375 10255 10390 10267
rect 10329 10235 10375 10246
rect 10617 10796 10663 10853
rect 10777 10806 10823 10807
rect 10602 10423 10617 10435
rect 10762 10796 10838 10806
rect 10762 10794 10777 10796
rect 10823 10794 10838 10796
rect 10762 10742 10774 10794
rect 10826 10742 10838 10794
rect 10762 10690 10777 10742
rect 10823 10690 10838 10742
rect 10762 10638 10774 10690
rect 10826 10638 10838 10690
rect 10762 10626 10777 10638
rect 10663 10423 10678 10435
rect 10602 10371 10614 10423
rect 10666 10371 10678 10423
rect 10602 10319 10617 10371
rect 10663 10319 10678 10371
rect 10602 10267 10614 10319
rect 10666 10267 10678 10319
rect 10602 10255 10617 10267
rect 10489 10189 10535 10246
rect 10663 10255 10678 10267
rect 10617 10235 10663 10246
rect 10823 10626 10838 10638
rect 10905 10796 10951 11075
rect 10777 10235 10823 10246
rect 9273 10143 10535 10189
rect 10489 10037 10535 10143
rect 9145 9991 10663 10037
rect 8857 9072 8903 9384
rect 8985 9934 9031 9945
rect 8985 9072 9031 9384
rect 8970 8961 8985 8973
rect 9145 9934 9191 9991
rect 9145 9072 9191 9384
rect 9031 8961 9046 8973
rect 8970 8909 8982 8961
rect 9034 8909 9046 8961
rect 8970 8857 8985 8909
rect 9031 8857 9046 8909
rect 8970 8805 8982 8857
rect 9034 8805 9046 8857
rect 8970 8793 8985 8805
rect 8857 8389 8903 8522
rect 9031 8793 9046 8805
rect 8985 8511 9031 8522
rect 9145 8511 9191 8522
rect 9273 9934 9319 9945
rect 9433 9934 9479 9945
rect 9418 9561 9433 9573
rect 9593 9934 9639 9945
rect 9479 9561 9494 9573
rect 9418 9509 9430 9561
rect 9482 9509 9494 9561
rect 9418 9457 9433 9509
rect 9479 9457 9494 9509
rect 9418 9405 9430 9457
rect 9482 9405 9494 9457
rect 9418 9393 9433 9405
rect 9273 9072 9319 9384
rect 9273 8465 9319 8522
rect 9479 9393 9494 9405
rect 9433 9072 9479 9384
rect 9433 8511 9479 8522
rect 9593 9072 9639 9384
rect 9593 8465 9639 8522
rect 9721 9934 9767 9991
rect 9721 9072 9767 9384
rect 9881 9934 9927 9945
rect 9881 9072 9927 9384
rect 9866 8961 9881 8973
rect 10041 9934 10087 9991
rect 10041 9072 10087 9384
rect 9927 8961 9942 8973
rect 9866 8909 9878 8961
rect 9930 8909 9942 8961
rect 9866 8857 9881 8909
rect 9927 8857 9942 8909
rect 9866 8805 9878 8857
rect 9930 8805 9942 8857
rect 9866 8793 9881 8805
rect 9721 8511 9767 8522
rect 9927 8793 9942 8805
rect 9881 8511 9927 8522
rect 10041 8511 10087 8522
rect 10169 9934 10215 9945
rect 10329 9934 10375 9945
rect 10314 9561 10329 9573
rect 10489 9934 10535 9945
rect 10375 9561 10390 9573
rect 10314 9509 10326 9561
rect 10378 9509 10390 9561
rect 10314 9457 10329 9509
rect 10375 9457 10390 9509
rect 10314 9405 10326 9457
rect 10378 9405 10390 9457
rect 10314 9393 10329 9405
rect 10169 9072 10215 9384
rect 10169 8465 10215 8522
rect 10375 9393 10390 9405
rect 10329 9072 10375 9384
rect 10617 9934 10663 9991
rect 10602 9761 10617 9773
rect 10777 9934 10823 9945
rect 10663 9761 10678 9773
rect 10602 9709 10614 9761
rect 10666 9709 10678 9761
rect 10602 9657 10617 9709
rect 10663 9657 10678 9709
rect 10602 9605 10614 9657
rect 10666 9605 10678 9657
rect 10602 9593 10617 9605
rect 10489 9072 10535 9384
rect 10474 8703 10489 8715
rect 10663 9593 10678 9605
rect 10617 9072 10663 9384
rect 10535 8703 10550 8715
rect 10474 8651 10486 8703
rect 10538 8651 10550 8703
rect 10474 8599 10489 8651
rect 10535 8599 10550 8651
rect 10474 8547 10486 8599
rect 10538 8547 10550 8599
rect 10474 8535 10489 8547
rect 10329 8511 10375 8522
rect 10535 8535 10550 8547
rect 10489 8465 10535 8522
rect 10777 9072 10823 9384
rect 10762 8961 10777 8973
rect 10905 9934 10951 10246
rect 10905 9072 10951 9384
rect 10823 8961 10838 8973
rect 10762 8909 10774 8961
rect 10826 8909 10838 8961
rect 10762 8857 10777 8909
rect 10823 8857 10838 8909
rect 10762 8805 10774 8857
rect 10826 8805 10838 8857
rect 10762 8793 10777 8805
rect 10617 8511 10663 8522
rect 10823 8793 10838 8805
rect 10777 8511 10823 8522
rect 9273 8419 10535 8465
rect 8697 8343 8777 8389
rect 8823 8343 8903 8389
rect 8697 8210 8743 8343
rect 8697 7381 8743 7660
rect 8857 8210 8903 8343
rect 10489 8327 10535 8419
rect 10722 8453 10798 8465
rect 10722 8401 10734 8453
rect 10786 8401 10798 8453
rect 10722 8349 10798 8401
rect 9145 8281 10663 8327
rect 10722 8297 10734 8349
rect 10786 8297 10798 8349
rect 10722 8285 10798 8297
rect 10905 8389 10951 8522
rect 11065 10796 11111 11075
rect 11065 9934 11111 10246
rect 11065 9072 11111 9384
rect 11065 8389 11111 8522
rect 10905 8343 10985 8389
rect 11031 8343 11111 8389
rect 8985 8210 9031 8221
rect 8970 7831 8985 7843
rect 9145 8210 9191 8281
rect 9418 8223 9494 8235
rect 9031 7831 9046 7843
rect 8970 7779 8982 7831
rect 9034 7779 9046 7831
rect 8970 7727 8985 7779
rect 9031 7727 9046 7779
rect 8970 7675 8982 7727
rect 9034 7675 9046 7727
rect 8970 7663 8985 7675
rect 8857 7381 8903 7660
rect 9031 7663 9046 7675
rect 8985 7649 9031 7660
rect 9145 7649 9191 7660
rect 9273 8210 9319 8221
rect 9418 8171 9430 8223
rect 9482 8171 9494 8223
rect 9418 8119 9433 8171
rect 9479 8119 9494 8171
rect 9418 8067 9430 8119
rect 9482 8067 9494 8119
rect 9418 8055 9433 8067
rect 9273 7603 9319 7660
rect 9479 8055 9494 8067
rect 9593 8210 9639 8221
rect 9433 7649 9479 7660
rect 9593 7603 9639 7660
rect 9721 8210 9767 8281
rect 9881 8210 9927 8221
rect 9866 7831 9881 7843
rect 10041 8210 10087 8281
rect 10314 8223 10390 8235
rect 9927 7831 9942 7843
rect 9866 7779 9878 7831
rect 9930 7779 9942 7831
rect 9866 7727 9881 7779
rect 9927 7727 9942 7779
rect 9866 7675 9878 7727
rect 9930 7675 9942 7727
rect 9866 7663 9881 7675
rect 9721 7649 9767 7660
rect 9927 7663 9942 7675
rect 9881 7649 9927 7660
rect 10041 7649 10087 7660
rect 10169 8210 10215 8221
rect 10314 8171 10326 8223
rect 10378 8171 10390 8223
rect 10314 8119 10329 8171
rect 10375 8119 10390 8171
rect 10314 8067 10326 8119
rect 10378 8067 10390 8119
rect 10314 8055 10329 8067
rect 10169 7603 10215 7660
rect 10375 8055 10390 8067
rect 10474 8223 10550 8235
rect 10474 8171 10486 8223
rect 10538 8171 10550 8223
rect 10474 8119 10489 8171
rect 10535 8119 10550 8171
rect 10474 8067 10486 8119
rect 10538 8067 10550 8119
rect 10474 8055 10489 8067
rect 10329 7649 10375 7660
rect 10535 8055 10550 8067
rect 10617 8210 10663 8281
rect 10489 7603 10535 7660
rect 10777 8210 10823 8221
rect 10762 7831 10777 7843
rect 10905 8210 10951 8343
rect 10823 7831 10838 7843
rect 10762 7779 10774 7831
rect 10826 7779 10838 7831
rect 10762 7727 10777 7779
rect 10823 7727 10838 7779
rect 10762 7675 10774 7727
rect 10826 7675 10838 7727
rect 10762 7663 10777 7675
rect 10617 7649 10663 7660
rect 10823 7663 10838 7675
rect 10777 7649 10823 7660
rect 9273 7557 10535 7603
rect 9969 7381 10149 7391
rect 10905 7381 10951 7660
rect 11065 8210 11111 8343
rect 11065 7381 11111 7660
rect 11211 11038 11244 11075
rect 11290 11038 11323 11084
rect 11211 10990 11323 11038
rect 11211 10944 11244 10990
rect 11290 10944 11323 10990
rect 11649 10965 11809 11675
rect 11867 11648 17055 11696
rect 18055 11794 18375 11842
rect 18055 11748 18136 11794
rect 18182 11748 18375 11794
rect 18055 11700 18375 11748
rect 11867 11602 11900 11648
rect 11946 11639 14626 11648
rect 11946 11602 11979 11639
rect 11867 11554 11979 11602
rect 11867 11508 11900 11554
rect 11946 11508 11979 11554
rect 11867 11460 11979 11508
rect 11867 11414 11900 11460
rect 11946 11414 11979 11460
rect 11867 11366 11979 11414
rect 11867 11320 11900 11366
rect 11946 11320 11979 11366
rect 11867 11272 11979 11320
rect 11867 11226 11900 11272
rect 11946 11226 11979 11272
rect 11867 11178 11979 11226
rect 11867 11132 11900 11178
rect 11946 11132 11979 11178
rect 11867 11084 11979 11132
rect 11867 11038 11900 11084
rect 11946 11038 11979 11084
rect 11867 10990 11979 11038
rect 11211 10896 11323 10944
rect 11211 10850 11244 10896
rect 11290 10850 11323 10896
rect 11211 10802 11323 10850
rect 11211 10756 11244 10802
rect 11290 10756 11323 10802
rect 11639 10953 11819 10965
rect 11639 10901 11651 10953
rect 11703 10901 11755 10953
rect 11807 10901 11819 10953
rect 11639 10849 11819 10901
rect 11639 10797 11651 10849
rect 11703 10797 11755 10849
rect 11807 10797 11819 10849
rect 11639 10785 11819 10797
rect 11867 10944 11900 10990
rect 11946 10944 11979 10990
rect 11867 10896 11979 10944
rect 11867 10850 11900 10896
rect 11946 10850 11979 10896
rect 11867 10802 11979 10850
rect 11211 10708 11323 10756
rect 11211 10662 11244 10708
rect 11290 10662 11323 10708
rect 11211 10614 11323 10662
rect 11211 10568 11244 10614
rect 11290 10568 11323 10614
rect 11211 10520 11323 10568
rect 11211 10474 11244 10520
rect 11290 10474 11323 10520
rect 11211 10426 11323 10474
rect 11211 10380 11244 10426
rect 11290 10380 11323 10426
rect 11211 10332 11323 10380
rect 11211 10286 11244 10332
rect 11290 10286 11323 10332
rect 11211 10238 11323 10286
rect 11211 10192 11244 10238
rect 11290 10192 11323 10238
rect 11211 10144 11323 10192
rect 11211 10098 11244 10144
rect 11290 10098 11323 10144
rect 11211 10050 11323 10098
rect 11211 10004 11244 10050
rect 11290 10004 11323 10050
rect 11211 9956 11323 10004
rect 11211 9910 11244 9956
rect 11290 9910 11323 9956
rect 11211 9862 11323 9910
rect 11211 9816 11244 9862
rect 11290 9816 11323 9862
rect 11211 9768 11323 9816
rect 11211 9722 11244 9768
rect 11290 9722 11323 9768
rect 11211 9674 11323 9722
rect 11211 9628 11244 9674
rect 11290 9628 11323 9674
rect 11211 9580 11323 9628
rect 11211 9534 11244 9580
rect 11290 9534 11323 9580
rect 11211 9486 11323 9534
rect 11211 9440 11244 9486
rect 11290 9440 11323 9486
rect 11211 9392 11323 9440
rect 11211 9346 11244 9392
rect 11290 9346 11323 9392
rect 11211 9298 11323 9346
rect 11211 9252 11244 9298
rect 11290 9252 11323 9298
rect 11211 9204 11323 9252
rect 11211 9158 11244 9204
rect 11290 9158 11323 9204
rect 11211 9110 11323 9158
rect 11211 9064 11244 9110
rect 11290 9064 11323 9110
rect 11211 9016 11323 9064
rect 11211 8970 11244 9016
rect 11290 8970 11323 9016
rect 11211 8922 11323 8970
rect 11211 8876 11244 8922
rect 11290 8876 11323 8922
rect 11211 8828 11323 8876
rect 11211 8782 11244 8828
rect 11290 8782 11323 8828
rect 11211 8734 11323 8782
rect 11211 8688 11244 8734
rect 11290 8688 11323 8734
rect 11211 8640 11323 8688
rect 11211 8594 11244 8640
rect 11290 8594 11323 8640
rect 11211 8546 11323 8594
rect 11211 8500 11244 8546
rect 11290 8500 11323 8546
rect 11211 8452 11323 8500
rect 11211 8406 11244 8452
rect 11290 8406 11323 8452
rect 11211 8358 11323 8406
rect 11211 8312 11244 8358
rect 11290 8312 11323 8358
rect 11211 8264 11323 8312
rect 11211 8218 11244 8264
rect 11290 8218 11323 8264
rect 11211 8170 11323 8218
rect 11211 8124 11244 8170
rect 11290 8124 11323 8170
rect 11211 8076 11323 8124
rect 11211 8030 11244 8076
rect 11290 8030 11323 8076
rect 11211 7982 11323 8030
rect 11211 7936 11244 7982
rect 11290 7936 11323 7982
rect 11211 7888 11323 7936
rect 11211 7842 11244 7888
rect 11290 7842 11323 7888
rect 11211 7794 11323 7842
rect 11211 7748 11244 7794
rect 11290 7748 11323 7794
rect 11211 7700 11323 7748
rect 11211 7654 11244 7700
rect 11290 7654 11323 7700
rect 11211 7606 11323 7654
rect 11211 7560 11244 7606
rect 11290 7560 11323 7606
rect 11211 7512 11323 7560
rect 11211 7466 11244 7512
rect 11290 7466 11323 7512
rect 11211 7418 11323 7466
rect 11211 7381 11244 7418
rect 8564 7379 11244 7381
rect 8564 7372 9981 7379
rect 7035 7327 9981 7372
rect 10033 7327 10085 7379
rect 10137 7372 11244 7379
rect 11290 7372 11323 7418
rect 10137 7327 11323 7372
rect 6229 7324 11323 7327
rect 6229 7278 6262 7324
rect 6308 7278 6356 7324
rect 6402 7278 6450 7324
rect 6496 7278 6544 7324
rect 6590 7278 6638 7324
rect 6684 7278 6732 7324
rect 6778 7278 6826 7324
rect 6872 7278 6920 7324
rect 6966 7278 7014 7324
rect 7060 7278 7108 7324
rect 7154 7278 7202 7324
rect 7248 7278 7296 7324
rect 7342 7278 7390 7324
rect 7436 7278 7484 7324
rect 7530 7278 7578 7324
rect 7624 7278 7672 7324
rect 7718 7278 7766 7324
rect 7812 7278 7860 7324
rect 7906 7278 7954 7324
rect 8000 7278 8048 7324
rect 8094 7278 8142 7324
rect 8188 7278 8236 7324
rect 8282 7278 8330 7324
rect 8376 7278 8424 7324
rect 8470 7278 8518 7324
rect 8564 7278 8612 7324
rect 8658 7278 8706 7324
rect 8752 7278 8800 7324
rect 8846 7278 8894 7324
rect 8940 7278 8988 7324
rect 9034 7278 9082 7324
rect 9128 7278 9176 7324
rect 9222 7278 9270 7324
rect 9316 7278 9364 7324
rect 9410 7278 9458 7324
rect 9504 7278 9552 7324
rect 9598 7278 9646 7324
rect 9692 7278 9740 7324
rect 9786 7278 9834 7324
rect 9880 7278 9928 7324
rect 9974 7278 10022 7324
rect 10068 7278 10116 7324
rect 10162 7278 10210 7324
rect 10256 7278 10304 7324
rect 10350 7278 10398 7324
rect 10444 7278 10492 7324
rect 10538 7278 10586 7324
rect 10632 7278 10680 7324
rect 10726 7278 10774 7324
rect 10820 7278 10868 7324
rect 10914 7278 10962 7324
rect 11008 7278 11056 7324
rect 11102 7278 11150 7324
rect 11196 7278 11244 7324
rect 11290 7278 11323 7324
rect 6229 7275 11323 7278
rect 6229 7223 6879 7275
rect 6931 7223 6983 7275
rect 7035 7223 9981 7275
rect 10033 7223 10085 7275
rect 10137 7223 11323 7275
rect 6229 7221 11323 7223
rect 11867 10756 11900 10802
rect 11946 10756 11979 10802
rect 11867 10708 11979 10756
rect 11867 10662 11900 10708
rect 11946 10662 11979 10708
rect 11867 10614 11979 10662
rect 11867 10568 11900 10614
rect 11946 10568 11979 10614
rect 11867 10520 11979 10568
rect 11867 10474 11900 10520
rect 11946 10474 11979 10520
rect 11867 10426 11979 10474
rect 11867 10380 11900 10426
rect 11946 10380 11979 10426
rect 11867 10332 11979 10380
rect 11867 10286 11900 10332
rect 11946 10286 11979 10332
rect 11867 10238 11979 10286
rect 11867 10192 11900 10238
rect 11946 10192 11979 10238
rect 11867 10144 11979 10192
rect 11867 10098 11900 10144
rect 11946 10098 11979 10144
rect 11867 10050 11979 10098
rect 11867 10004 11900 10050
rect 11946 10004 11979 10050
rect 11867 9956 11979 10004
rect 11867 9910 11900 9956
rect 11946 9910 11979 9956
rect 11867 9862 11979 9910
rect 11867 9816 11900 9862
rect 11946 9816 11979 9862
rect 11867 9768 11979 9816
rect 11867 9722 11900 9768
rect 11946 9722 11979 9768
rect 11867 9674 11979 9722
rect 11867 9628 11900 9674
rect 11946 9628 11979 9674
rect 11867 9580 11979 9628
rect 11867 9534 11900 9580
rect 11946 9534 11979 9580
rect 11867 9486 11979 9534
rect 11867 9440 11900 9486
rect 11946 9440 11979 9486
rect 11867 9392 11979 9440
rect 11867 9346 11900 9392
rect 11946 9346 11979 9392
rect 11867 9298 11979 9346
rect 11867 9252 11900 9298
rect 11946 9252 11979 9298
rect 11867 9204 11979 9252
rect 11867 9158 11900 9204
rect 11946 9158 11979 9204
rect 11867 9110 11979 9158
rect 11867 9064 11900 9110
rect 11946 9064 11979 9110
rect 11867 9016 11979 9064
rect 11867 8970 11900 9016
rect 11946 8970 11979 9016
rect 11867 8922 11979 8970
rect 11867 8876 11900 8922
rect 11946 8876 11979 8922
rect 11867 8828 11979 8876
rect 11867 8782 11900 8828
rect 11946 8782 11979 8828
rect 11867 8734 11979 8782
rect 11867 8688 11900 8734
rect 11946 8688 11979 8734
rect 11867 8640 11979 8688
rect 11867 8594 11900 8640
rect 11946 8594 11979 8640
rect 11867 8546 11979 8594
rect 11867 8500 11900 8546
rect 11946 8500 11979 8546
rect 11867 8452 11979 8500
rect 11867 8406 11900 8452
rect 11946 8406 11979 8452
rect 11867 8358 11979 8406
rect 11867 8312 11900 8358
rect 11946 8312 11979 8358
rect 11867 8264 11979 8312
rect 11867 8218 11900 8264
rect 11946 8218 11979 8264
rect 11867 8170 11979 8218
rect 11867 8124 11900 8170
rect 11946 8124 11979 8170
rect 11867 8076 11979 8124
rect 11867 8030 11900 8076
rect 11946 8030 11979 8076
rect 11867 7982 11979 8030
rect 11867 7936 11900 7982
rect 11946 7936 11979 7982
rect 11867 7888 11979 7936
rect 11867 7842 11900 7888
rect 11946 7842 11979 7888
rect 11867 7794 11979 7842
rect 11867 7748 11900 7794
rect 11946 7748 11979 7794
rect 11867 7700 11979 7748
rect 11867 7654 11900 7700
rect 11946 7654 11979 7700
rect 11867 7606 11979 7654
rect 11867 7560 11900 7606
rect 11946 7560 11979 7606
rect 11867 7512 11979 7560
rect 11867 7466 11900 7512
rect 11946 7466 11979 7512
rect 11867 7418 11979 7466
rect 11867 7372 11900 7418
rect 11946 7381 11979 7418
rect 12079 11364 12125 11639
rect 12079 10328 12125 10764
rect 12079 9292 12125 9728
rect 12079 8435 12125 8692
rect 12239 11364 12285 11639
rect 12527 11444 14045 11490
rect 12367 11364 12413 11375
rect 12352 10953 12367 10965
rect 12527 11364 12573 11444
rect 12413 10953 12428 10965
rect 12352 10901 12364 10953
rect 12416 10901 12428 10953
rect 12352 10849 12367 10901
rect 12413 10849 12428 10901
rect 12352 10797 12364 10849
rect 12416 10797 12428 10849
rect 12352 10785 12367 10797
rect 12239 10328 12285 10764
rect 12413 10785 12428 10797
rect 12367 10753 12413 10764
rect 12527 10753 12573 10764
rect 12655 11364 12701 11375
rect 12800 11373 12876 11385
rect 12800 11321 12812 11373
rect 12864 11321 12876 11373
rect 12800 11269 12815 11321
rect 12861 11269 12876 11321
rect 12800 11217 12812 11269
rect 12864 11217 12876 11269
rect 12800 11205 12815 11217
rect 12655 10684 12701 10764
rect 12861 11205 12876 11217
rect 12975 11364 13021 11375
rect 12815 10753 12861 10764
rect 12975 10684 13021 10764
rect 13103 11364 13149 11444
rect 13263 11364 13309 11375
rect 13248 10953 13263 10965
rect 13423 11364 13469 11444
rect 13999 11385 14045 11444
rect 13309 10953 13324 10965
rect 13248 10901 13260 10953
rect 13312 10901 13324 10953
rect 13248 10849 13263 10901
rect 13309 10849 13324 10901
rect 13248 10797 13260 10849
rect 13312 10797 13324 10849
rect 13248 10785 13263 10797
rect 13103 10753 13149 10764
rect 13309 10785 13324 10797
rect 13263 10753 13309 10764
rect 13423 10753 13469 10764
rect 13551 11364 13597 11375
rect 13696 11373 13772 11385
rect 13696 11321 13708 11373
rect 13760 11321 13772 11373
rect 13696 11269 13711 11321
rect 13757 11269 13772 11321
rect 13696 11217 13708 11269
rect 13760 11217 13772 11269
rect 13696 11205 13711 11217
rect 13551 10684 13597 10764
rect 13757 11205 13772 11217
rect 13871 11364 13917 11375
rect 13711 10753 13757 10764
rect 13984 11373 14060 11385
rect 13984 11321 13996 11373
rect 14048 11321 14060 11373
rect 13984 11269 13999 11321
rect 14045 11269 14060 11321
rect 13984 11217 13996 11269
rect 14048 11217 14060 11269
rect 13984 11205 13999 11217
rect 13871 10684 13917 10764
rect 14045 11205 14060 11217
rect 14159 11364 14205 11375
rect 14144 10953 14159 10965
rect 14287 11364 14333 11639
rect 14205 10953 14220 10965
rect 14144 10901 14156 10953
rect 14208 10901 14220 10953
rect 14144 10849 14159 10901
rect 14205 10849 14220 10901
rect 14144 10797 14156 10849
rect 14208 10797 14220 10849
rect 14144 10785 14159 10797
rect 13999 10753 14045 10764
rect 14205 10785 14220 10797
rect 14159 10753 14205 10764
rect 12655 10638 13917 10684
rect 13871 10454 13917 10638
rect 12527 10408 14045 10454
rect 12239 9292 12285 9728
rect 12367 10328 12413 10339
rect 12367 9292 12413 9728
rect 12352 9273 12367 9285
rect 12527 10328 12573 10408
rect 12527 9292 12573 9728
rect 12413 9273 12428 9285
rect 12352 9221 12364 9273
rect 12416 9221 12428 9273
rect 12352 9169 12367 9221
rect 12413 9169 12428 9221
rect 12352 9117 12364 9169
rect 12416 9117 12428 9169
rect 12352 9105 12367 9117
rect 12239 8435 12285 8692
rect 12413 9105 12428 9117
rect 12367 8681 12413 8692
rect 12527 8681 12573 8692
rect 12655 10328 12701 10339
rect 12815 10331 12861 10339
rect 12800 10328 12876 10331
rect 12800 10319 12815 10328
rect 12861 10319 12876 10328
rect 12800 10267 12812 10319
rect 12864 10267 12876 10319
rect 12800 10215 12815 10267
rect 12861 10215 12876 10267
rect 12800 10163 12812 10215
rect 12864 10163 12876 10215
rect 12800 10151 12815 10163
rect 12655 9292 12701 9728
rect 12655 8612 12701 8692
rect 12861 10151 12876 10163
rect 12975 10328 13021 10339
rect 12815 9292 12861 9728
rect 12815 8681 12861 8692
rect 12975 9292 13021 9728
rect 12975 8612 13021 8692
rect 13103 10328 13149 10408
rect 13103 9292 13149 9728
rect 13263 10328 13309 10339
rect 13263 9292 13309 9728
rect 13248 9273 13263 9285
rect 13423 10328 13469 10408
rect 13423 9292 13469 9728
rect 13309 9273 13324 9285
rect 13248 9221 13260 9273
rect 13312 9221 13324 9273
rect 13248 9169 13263 9221
rect 13309 9169 13324 9221
rect 13248 9117 13260 9169
rect 13312 9117 13324 9169
rect 13248 9105 13263 9117
rect 13103 8681 13149 8692
rect 13309 9105 13324 9117
rect 13263 8681 13309 8692
rect 13423 8681 13469 8692
rect 13551 10328 13597 10339
rect 13711 10331 13757 10339
rect 13696 10328 13772 10331
rect 13696 10319 13711 10328
rect 13757 10319 13772 10328
rect 13696 10267 13708 10319
rect 13760 10267 13772 10319
rect 13696 10215 13711 10267
rect 13757 10215 13772 10267
rect 13696 10163 13708 10215
rect 13760 10163 13772 10215
rect 13696 10151 13711 10163
rect 13551 9292 13597 9728
rect 13551 8612 13597 8692
rect 13757 10151 13772 10163
rect 13871 10328 13917 10339
rect 13711 9292 13757 9728
rect 13999 10328 14045 10408
rect 13984 10293 13999 10305
rect 14159 10328 14205 10339
rect 14045 10293 14060 10305
rect 13984 10241 13996 10293
rect 14048 10241 14060 10293
rect 13984 10189 13999 10241
rect 14045 10189 14060 10241
rect 13984 10137 13996 10189
rect 14048 10137 14060 10189
rect 13984 10125 13999 10137
rect 13871 9292 13917 9728
rect 13856 8873 13871 8885
rect 14045 10125 14060 10137
rect 13999 9292 14045 9728
rect 13917 8873 13932 8885
rect 13856 8821 13868 8873
rect 13920 8821 13932 8873
rect 13856 8769 13871 8821
rect 13917 8769 13932 8821
rect 13856 8717 13868 8769
rect 13920 8717 13932 8769
rect 13856 8705 13871 8717
rect 13711 8681 13757 8692
rect 13917 8705 13932 8717
rect 13871 8612 13917 8692
rect 14159 9292 14205 9728
rect 14144 9273 14159 9285
rect 14287 10328 14333 10764
rect 14287 9292 14333 9728
rect 14205 9273 14220 9285
rect 14144 9221 14156 9273
rect 14208 9221 14220 9273
rect 14144 9169 14159 9221
rect 14205 9169 14220 9221
rect 14144 9117 14156 9169
rect 14208 9117 14220 9169
rect 14144 9105 14159 9117
rect 13999 8681 14045 8692
rect 14205 9105 14220 9117
rect 14159 8681 14205 8692
rect 12079 8389 12159 8435
rect 12205 8389 12285 8435
rect 12388 8563 12464 8575
rect 12655 8566 13917 8612
rect 12388 8511 12400 8563
rect 12452 8511 12464 8563
rect 12388 8459 12464 8511
rect 12388 8407 12400 8459
rect 12452 8407 12464 8459
rect 12388 8395 12464 8407
rect 12079 8256 12125 8389
rect 12079 7381 12125 7656
rect 12239 8256 12285 8389
rect 13871 8382 13917 8566
rect 14287 8435 14333 8692
rect 14447 11364 14493 11639
rect 14447 10328 14493 10764
rect 14447 9292 14493 9728
rect 14447 8435 14493 8692
rect 14287 8389 14367 8435
rect 14413 8389 14493 8435
rect 12527 8336 14045 8382
rect 12367 8256 12413 8267
rect 12239 7381 12285 7656
rect 12352 7823 12367 7835
rect 12527 8256 12573 8336
rect 12413 7823 12428 7835
rect 12352 7771 12364 7823
rect 12416 7771 12428 7823
rect 12352 7719 12367 7771
rect 12413 7719 12428 7771
rect 12352 7667 12364 7719
rect 12416 7667 12428 7719
rect 12352 7656 12367 7667
rect 12413 7656 12428 7667
rect 12352 7655 12428 7656
rect 12367 7645 12413 7655
rect 12527 7645 12573 7656
rect 12655 8256 12701 8267
rect 12815 8256 12861 8267
rect 12800 8223 12815 8235
rect 12975 8256 13021 8267
rect 12861 8223 12876 8235
rect 12800 8171 12812 8223
rect 12864 8171 12876 8223
rect 12800 8119 12815 8171
rect 12861 8119 12876 8171
rect 12800 8067 12812 8119
rect 12864 8067 12876 8119
rect 12800 8055 12815 8067
rect 12655 7576 12701 7656
rect 12861 8055 12876 8067
rect 12815 7645 12861 7656
rect 12975 7576 13021 7656
rect 13103 8256 13149 8336
rect 13263 8256 13309 8267
rect 13103 7645 13149 7656
rect 13248 7823 13263 7835
rect 13423 8256 13469 8336
rect 13309 7823 13324 7835
rect 13248 7771 13260 7823
rect 13312 7771 13324 7823
rect 13248 7719 13263 7771
rect 13309 7719 13324 7771
rect 13248 7667 13260 7719
rect 13312 7667 13324 7719
rect 13248 7656 13263 7667
rect 13309 7656 13324 7667
rect 13248 7655 13324 7656
rect 13263 7645 13309 7655
rect 13423 7645 13469 7656
rect 13551 8256 13597 8267
rect 13711 8256 13757 8267
rect 13696 8223 13711 8235
rect 13871 8256 13917 8267
rect 13757 8223 13772 8235
rect 13696 8171 13708 8223
rect 13760 8171 13772 8223
rect 13696 8119 13711 8171
rect 13757 8119 13772 8171
rect 13696 8067 13708 8119
rect 13760 8067 13772 8119
rect 13696 8055 13711 8067
rect 13551 7576 13597 7656
rect 13757 8055 13772 8067
rect 13856 8223 13871 8235
rect 13999 8256 14045 8336
rect 13917 8223 13932 8235
rect 13856 8171 13868 8223
rect 13920 8171 13932 8223
rect 13856 8119 13871 8171
rect 13917 8119 13932 8171
rect 13856 8067 13868 8119
rect 13920 8067 13932 8119
rect 13856 8055 13871 8067
rect 13711 7645 13757 7656
rect 13917 8055 13932 8067
rect 13871 7576 13917 7656
rect 14159 8256 14205 8267
rect 13999 7645 14045 7656
rect 14144 7823 14159 7835
rect 14287 8256 14333 8389
rect 14205 7823 14220 7835
rect 14144 7771 14156 7823
rect 14208 7771 14220 7823
rect 14144 7719 14159 7771
rect 14205 7719 14220 7771
rect 14144 7667 14156 7719
rect 14208 7667 14220 7719
rect 14144 7656 14159 7667
rect 14205 7656 14220 7667
rect 14144 7655 14220 7656
rect 14159 7645 14205 7655
rect 12655 7530 13917 7576
rect 14287 7381 14333 7656
rect 14447 8256 14493 8389
rect 14447 7381 14493 7656
rect 14593 11602 14626 11639
rect 14672 11639 16976 11648
rect 14672 11602 14705 11639
rect 14593 11554 14705 11602
rect 14593 11508 14626 11554
rect 14672 11508 14705 11554
rect 14593 11460 14705 11508
rect 14593 11414 14626 11460
rect 14672 11414 14705 11460
rect 14593 11366 14705 11414
rect 14593 11320 14626 11366
rect 14672 11320 14705 11366
rect 14593 11272 14705 11320
rect 14593 11226 14626 11272
rect 14672 11226 14705 11272
rect 14593 11178 14705 11226
rect 14593 11132 14626 11178
rect 14672 11132 14705 11178
rect 14593 11084 14705 11132
rect 14593 11038 14626 11084
rect 14672 11038 14705 11084
rect 14593 10990 14705 11038
rect 14593 10944 14626 10990
rect 14672 10944 14705 10990
rect 14593 10896 14705 10944
rect 14593 10850 14626 10896
rect 14672 10850 14705 10896
rect 14593 10802 14705 10850
rect 14593 10756 14626 10802
rect 14672 10756 14705 10802
rect 14593 10708 14705 10756
rect 14593 10662 14626 10708
rect 14672 10662 14705 10708
rect 14593 10614 14705 10662
rect 14593 10568 14626 10614
rect 14672 10568 14705 10614
rect 14593 10520 14705 10568
rect 14593 10474 14626 10520
rect 14672 10474 14705 10520
rect 14593 10426 14705 10474
rect 14593 10380 14626 10426
rect 14672 10380 14705 10426
rect 14593 10332 14705 10380
rect 14593 10286 14626 10332
rect 14672 10286 14705 10332
rect 14593 10238 14705 10286
rect 14593 10192 14626 10238
rect 14672 10192 14705 10238
rect 14593 10144 14705 10192
rect 14593 10098 14626 10144
rect 14672 10098 14705 10144
rect 14593 10050 14705 10098
rect 14593 10004 14626 10050
rect 14672 10004 14705 10050
rect 14593 9956 14705 10004
rect 14593 9910 14626 9956
rect 14672 9910 14705 9956
rect 14593 9862 14705 9910
rect 14593 9816 14626 9862
rect 14672 9816 14705 9862
rect 14593 9768 14705 9816
rect 14593 9722 14626 9768
rect 14672 9722 14705 9768
rect 14593 9674 14705 9722
rect 14593 9628 14626 9674
rect 14672 9628 14705 9674
rect 14593 9580 14705 9628
rect 14593 9534 14626 9580
rect 14672 9534 14705 9580
rect 14593 9486 14705 9534
rect 14593 9440 14626 9486
rect 14672 9440 14705 9486
rect 14593 9392 14705 9440
rect 14593 9346 14626 9392
rect 14672 9346 14705 9392
rect 14593 9298 14705 9346
rect 14593 9252 14626 9298
rect 14672 9252 14705 9298
rect 14593 9204 14705 9252
rect 14593 9158 14626 9204
rect 14672 9158 14705 9204
rect 14593 9110 14705 9158
rect 14593 9064 14626 9110
rect 14672 9064 14705 9110
rect 14593 9016 14705 9064
rect 14593 8970 14626 9016
rect 14672 8970 14705 9016
rect 14593 8922 14705 8970
rect 14593 8876 14626 8922
rect 14672 8876 14705 8922
rect 14593 8828 14705 8876
rect 14593 8782 14626 8828
rect 14672 8782 14705 8828
rect 14593 8734 14705 8782
rect 14593 8688 14626 8734
rect 14672 8688 14705 8734
rect 14593 8640 14705 8688
rect 14593 8594 14626 8640
rect 14672 8594 14705 8640
rect 14593 8546 14705 8594
rect 14593 8500 14626 8546
rect 14672 8500 14705 8546
rect 14593 8452 14705 8500
rect 14593 8406 14626 8452
rect 14672 8406 14705 8452
rect 14593 8358 14705 8406
rect 14593 8312 14626 8358
rect 14672 8312 14705 8358
rect 14593 8264 14705 8312
rect 14593 8218 14626 8264
rect 14672 8218 14705 8264
rect 14593 8170 14705 8218
rect 14593 8124 14626 8170
rect 14672 8124 14705 8170
rect 14593 8076 14705 8124
rect 14593 8030 14626 8076
rect 14672 8030 14705 8076
rect 14593 7982 14705 8030
rect 14593 7936 14626 7982
rect 14672 7936 14705 7982
rect 14593 7888 14705 7936
rect 14593 7842 14626 7888
rect 14672 7842 14705 7888
rect 14593 7794 14705 7842
rect 14593 7748 14626 7794
rect 14672 7748 14705 7794
rect 14593 7700 14705 7748
rect 14593 7654 14626 7700
rect 14672 7654 14705 7700
rect 14593 7606 14705 7654
rect 14873 11364 14919 11639
rect 14873 10328 14919 10764
rect 14873 9292 14919 9728
rect 14873 8435 14919 8692
rect 15033 11364 15079 11639
rect 15146 11373 15222 11385
rect 15146 11321 15158 11373
rect 15210 11321 15222 11373
rect 15146 11269 15161 11321
rect 15207 11269 15222 11321
rect 15146 11217 15158 11269
rect 15210 11217 15222 11269
rect 15146 11205 15161 11217
rect 15033 10328 15079 10764
rect 15207 11205 15222 11217
rect 15321 11364 15367 11639
rect 15161 10753 15207 10764
rect 15481 11364 15527 11375
rect 15466 10953 15481 10965
rect 15641 11364 15687 11639
rect 15527 10953 15542 10965
rect 15466 10901 15478 10953
rect 15530 10901 15542 10953
rect 15466 10849 15481 10901
rect 15527 10849 15542 10901
rect 15466 10797 15478 10849
rect 15530 10797 15542 10849
rect 15466 10785 15481 10797
rect 15161 10328 15207 10339
rect 15146 10293 15161 10305
rect 15321 10328 15367 10764
rect 15527 10785 15542 10797
rect 15481 10753 15527 10764
rect 15786 11373 15862 11385
rect 15786 11321 15798 11373
rect 15850 11321 15862 11373
rect 15786 11269 15801 11321
rect 15847 11269 15862 11321
rect 15786 11217 15798 11269
rect 15850 11217 15862 11269
rect 15786 11205 15801 11217
rect 15207 10293 15222 10305
rect 15146 10241 15158 10293
rect 15210 10241 15222 10293
rect 15146 10189 15161 10241
rect 15207 10189 15222 10241
rect 15146 10137 15158 10189
rect 15210 10137 15222 10189
rect 15146 10125 15161 10137
rect 15033 9292 15079 9728
rect 15033 8435 15079 8692
rect 15207 10125 15222 10137
rect 15161 9292 15207 9728
rect 15161 8681 15207 8692
rect 15321 9292 15367 9728
rect 15481 10328 15527 10339
rect 15481 9292 15527 9728
rect 15466 8873 15481 8885
rect 15641 10328 15687 10764
rect 15847 11205 15862 11217
rect 15961 11364 16007 11639
rect 15801 10753 15847 10764
rect 16121 11364 16167 11375
rect 16106 10953 16121 10965
rect 16281 11364 16327 11639
rect 16167 10953 16182 10965
rect 16106 10901 16118 10953
rect 16170 10901 16182 10953
rect 16106 10849 16121 10901
rect 16167 10849 16182 10901
rect 16106 10797 16118 10849
rect 16170 10797 16182 10849
rect 16106 10785 16121 10797
rect 15801 10328 15847 10339
rect 15786 10293 15801 10305
rect 15961 10328 16007 10764
rect 16167 10785 16182 10797
rect 16121 10753 16167 10764
rect 16426 11373 16502 11385
rect 16426 11321 16438 11373
rect 16490 11321 16502 11373
rect 16426 11269 16441 11321
rect 16487 11269 16502 11321
rect 16426 11217 16438 11269
rect 16490 11217 16502 11269
rect 16426 11205 16441 11217
rect 15847 10293 15862 10305
rect 15786 10241 15798 10293
rect 15850 10241 15862 10293
rect 15786 10189 15801 10241
rect 15847 10189 15862 10241
rect 15786 10137 15798 10189
rect 15850 10137 15862 10189
rect 15786 10125 15801 10137
rect 15641 9292 15687 9728
rect 15527 8873 15542 8885
rect 15466 8821 15478 8873
rect 15530 8821 15542 8873
rect 15466 8769 15481 8821
rect 15527 8769 15542 8821
rect 15466 8717 15478 8769
rect 15530 8717 15542 8769
rect 15466 8705 15481 8717
rect 14873 8389 14953 8435
rect 14999 8389 15079 8435
rect 15174 8568 15250 8580
rect 15174 8516 15186 8568
rect 15238 8516 15250 8568
rect 15174 8464 15250 8516
rect 15174 8412 15186 8464
rect 15238 8412 15250 8464
rect 15174 8400 15250 8412
rect 14873 8256 14919 8389
rect 14873 7645 14919 7656
rect 15033 8256 15079 8389
rect 15161 8256 15207 8267
rect 15146 7833 15161 7845
rect 15321 8256 15367 8692
rect 15527 8705 15542 8717
rect 15481 8681 15527 8692
rect 15207 7833 15222 7845
rect 15146 7781 15158 7833
rect 15210 7781 15222 7833
rect 15146 7729 15161 7781
rect 15207 7729 15222 7781
rect 15146 7677 15158 7729
rect 15210 7677 15222 7729
rect 15146 7665 15161 7677
rect 15033 7645 15079 7656
rect 15207 7665 15222 7677
rect 15161 7645 15207 7656
rect 15481 8256 15527 8267
rect 15466 8223 15481 8235
rect 15641 8256 15687 8692
rect 15847 10125 15862 10137
rect 15801 9292 15847 9728
rect 15801 8681 15847 8692
rect 15961 9292 16007 9728
rect 16121 10328 16167 10339
rect 16121 9292 16167 9728
rect 16106 8873 16121 8885
rect 16281 10328 16327 10764
rect 16487 11205 16502 11217
rect 16569 11364 16615 11639
rect 16441 10753 16487 10764
rect 16441 10328 16487 10339
rect 16426 10293 16441 10305
rect 16569 10328 16615 10764
rect 16487 10293 16502 10305
rect 16426 10241 16438 10293
rect 16490 10241 16502 10293
rect 16426 10189 16441 10241
rect 16487 10189 16502 10241
rect 16426 10137 16438 10189
rect 16490 10137 16502 10189
rect 16426 10125 16441 10137
rect 16281 9292 16327 9728
rect 16167 8873 16182 8885
rect 16106 8821 16118 8873
rect 16170 8821 16182 8873
rect 16106 8769 16121 8821
rect 16167 8769 16182 8821
rect 16106 8717 16118 8769
rect 16170 8717 16182 8769
rect 16106 8705 16121 8717
rect 15527 8223 15542 8235
rect 15466 8171 15478 8223
rect 15530 8171 15542 8223
rect 15466 8119 15481 8171
rect 15527 8119 15542 8171
rect 15466 8067 15478 8119
rect 15530 8067 15542 8119
rect 15466 8055 15481 8067
rect 14593 7560 14626 7606
rect 14672 7560 14705 7606
rect 14593 7512 14705 7560
rect 14593 7466 14626 7512
rect 14672 7466 14705 7512
rect 14593 7418 14705 7466
rect 14593 7381 14626 7418
rect 11946 7372 14626 7381
rect 14672 7381 14705 7418
rect 15321 7381 15367 7656
rect 15527 8055 15542 8067
rect 15481 7645 15527 7656
rect 15801 8256 15847 8267
rect 15786 7833 15801 7845
rect 15961 8256 16007 8692
rect 16167 8705 16182 8717
rect 16121 8681 16167 8692
rect 15847 7833 15862 7845
rect 15786 7781 15798 7833
rect 15850 7781 15862 7833
rect 15786 7729 15801 7781
rect 15847 7729 15862 7781
rect 15786 7677 15798 7729
rect 15850 7677 15862 7729
rect 15786 7665 15801 7677
rect 15641 7381 15687 7656
rect 15847 7665 15862 7677
rect 15801 7645 15847 7656
rect 16121 8256 16167 8267
rect 16106 8223 16121 8235
rect 16281 8256 16327 8692
rect 16487 10125 16502 10137
rect 16441 9292 16487 9728
rect 16441 8681 16487 8692
rect 16569 9292 16615 9728
rect 16569 8435 16615 8692
rect 16729 11364 16775 11639
rect 16729 10328 16775 10764
rect 16729 9292 16775 9728
rect 16729 8435 16775 8692
rect 16569 8389 16649 8435
rect 16695 8389 16775 8435
rect 16167 8223 16182 8235
rect 16106 8171 16118 8223
rect 16170 8171 16182 8223
rect 16106 8119 16121 8171
rect 16167 8119 16182 8171
rect 16106 8067 16118 8119
rect 16170 8067 16182 8119
rect 16106 8055 16121 8067
rect 15961 7381 16007 7656
rect 16167 8055 16182 8067
rect 16121 7645 16167 7656
rect 16441 8256 16487 8267
rect 16426 7833 16441 7845
rect 16569 8256 16615 8389
rect 16487 7833 16502 7845
rect 16426 7781 16438 7833
rect 16490 7781 16502 7833
rect 16426 7729 16441 7781
rect 16487 7729 16502 7781
rect 16426 7677 16438 7729
rect 16490 7677 16502 7729
rect 16426 7665 16441 7677
rect 16281 7381 16327 7656
rect 16487 7665 16502 7677
rect 16441 7645 16487 7656
rect 16569 7381 16615 7656
rect 16729 8256 16775 8389
rect 16729 7381 16775 7656
rect 16943 11602 16976 11639
rect 17022 11602 17055 11648
rect 16943 11554 17055 11602
rect 16943 11508 16976 11554
rect 17022 11508 17055 11554
rect 16943 11460 17055 11508
rect 16943 11414 16976 11460
rect 17022 11414 17055 11460
rect 16943 11366 17055 11414
rect 16943 11320 16976 11366
rect 17022 11320 17055 11366
rect 16943 11272 17055 11320
rect 16943 11226 16976 11272
rect 17022 11226 17055 11272
rect 16943 11178 17055 11226
rect 16943 11132 16976 11178
rect 17022 11132 17055 11178
rect 16943 11084 17055 11132
rect 16943 11038 16976 11084
rect 17022 11038 17055 11084
rect 16943 10990 17055 11038
rect 16943 10944 16976 10990
rect 17022 10944 17055 10990
rect 17113 10965 17273 11627
rect 17375 11385 17535 11675
rect 18055 11654 18136 11700
rect 18182 11654 18375 11700
rect 18055 11606 18375 11654
rect 18055 11560 18136 11606
rect 18182 11560 18375 11606
rect 18055 11512 18375 11560
rect 18055 11466 18136 11512
rect 18182 11466 18375 11512
rect 18055 11418 18375 11466
rect 17365 11373 17545 11385
rect 17365 11321 17377 11373
rect 17429 11321 17481 11373
rect 17533 11321 17545 11373
rect 17365 11269 17545 11321
rect 17365 11217 17377 11269
rect 17429 11217 17481 11269
rect 17533 11217 17545 11269
rect 17365 11205 17545 11217
rect 18055 11372 18136 11418
rect 18182 11372 18375 11418
rect 18055 11324 18375 11372
rect 18055 11278 18136 11324
rect 18182 11278 18375 11324
rect 18055 11230 18375 11278
rect 18055 11184 18136 11230
rect 18182 11184 18375 11230
rect 18055 11136 18375 11184
rect 18055 11090 18136 11136
rect 18182 11090 18375 11136
rect 18055 11042 18375 11090
rect 18055 10996 18136 11042
rect 18182 10996 18375 11042
rect 16943 10896 17055 10944
rect 16943 10850 16976 10896
rect 17022 10850 17055 10896
rect 16943 10802 17055 10850
rect 16943 10756 16976 10802
rect 17022 10756 17055 10802
rect 17103 10953 17283 10965
rect 17103 10901 17115 10953
rect 17167 10901 17219 10953
rect 17271 10901 17283 10953
rect 17103 10849 17283 10901
rect 17103 10797 17115 10849
rect 17167 10797 17219 10849
rect 17271 10797 17283 10849
rect 17103 10785 17283 10797
rect 18055 10948 18375 10996
rect 18055 10902 18136 10948
rect 18182 10902 18375 10948
rect 18055 10854 18375 10902
rect 18055 10808 18136 10854
rect 18182 10808 18375 10854
rect 16943 10708 17055 10756
rect 16943 10662 16976 10708
rect 17022 10662 17055 10708
rect 16943 10614 17055 10662
rect 16943 10568 16976 10614
rect 17022 10568 17055 10614
rect 16943 10520 17055 10568
rect 16943 10474 16976 10520
rect 17022 10474 17055 10520
rect 16943 10426 17055 10474
rect 16943 10380 16976 10426
rect 17022 10380 17055 10426
rect 16943 10332 17055 10380
rect 16943 10286 16976 10332
rect 17022 10286 17055 10332
rect 16943 10238 17055 10286
rect 16943 10192 16976 10238
rect 17022 10192 17055 10238
rect 16943 10144 17055 10192
rect 16943 10098 16976 10144
rect 17022 10098 17055 10144
rect 16943 10050 17055 10098
rect 16943 10004 16976 10050
rect 17022 10004 17055 10050
rect 16943 9956 17055 10004
rect 16943 9910 16976 9956
rect 17022 9910 17055 9956
rect 16943 9862 17055 9910
rect 16943 9816 16976 9862
rect 17022 9816 17055 9862
rect 16943 9768 17055 9816
rect 16943 9722 16976 9768
rect 17022 9722 17055 9768
rect 16943 9674 17055 9722
rect 16943 9628 16976 9674
rect 17022 9628 17055 9674
rect 16943 9580 17055 9628
rect 16943 9534 16976 9580
rect 17022 9534 17055 9580
rect 16943 9486 17055 9534
rect 16943 9440 16976 9486
rect 17022 9440 17055 9486
rect 16943 9392 17055 9440
rect 16943 9346 16976 9392
rect 17022 9346 17055 9392
rect 16943 9298 17055 9346
rect 16943 9252 16976 9298
rect 17022 9252 17055 9298
rect 16943 9204 17055 9252
rect 16943 9158 16976 9204
rect 17022 9158 17055 9204
rect 16943 9110 17055 9158
rect 16943 9064 16976 9110
rect 17022 9064 17055 9110
rect 16943 9016 17055 9064
rect 16943 8970 16976 9016
rect 17022 8970 17055 9016
rect 16943 8922 17055 8970
rect 16943 8876 16976 8922
rect 17022 8876 17055 8922
rect 16943 8828 17055 8876
rect 16943 8782 16976 8828
rect 17022 8782 17055 8828
rect 16943 8734 17055 8782
rect 16943 8688 16976 8734
rect 17022 8688 17055 8734
rect 16943 8640 17055 8688
rect 16943 8594 16976 8640
rect 17022 8594 17055 8640
rect 16943 8546 17055 8594
rect 16943 8500 16976 8546
rect 17022 8500 17055 8546
rect 16943 8452 17055 8500
rect 16943 8406 16976 8452
rect 17022 8406 17055 8452
rect 16943 8358 17055 8406
rect 16943 8312 16976 8358
rect 17022 8312 17055 8358
rect 16943 8264 17055 8312
rect 16943 8218 16976 8264
rect 17022 8218 17055 8264
rect 16943 8170 17055 8218
rect 16943 8124 16976 8170
rect 17022 8124 17055 8170
rect 16943 8076 17055 8124
rect 16943 8030 16976 8076
rect 17022 8030 17055 8076
rect 16943 7982 17055 8030
rect 16943 7936 16976 7982
rect 17022 7936 17055 7982
rect 16943 7888 17055 7936
rect 16943 7842 16976 7888
rect 17022 7842 17055 7888
rect 16943 7794 17055 7842
rect 16943 7748 16976 7794
rect 17022 7748 17055 7794
rect 16943 7700 17055 7748
rect 16943 7654 16976 7700
rect 17022 7654 17055 7700
rect 16943 7606 17055 7654
rect 16943 7560 16976 7606
rect 17022 7560 17055 7606
rect 16943 7541 17055 7560
rect 18055 10760 18375 10808
rect 18055 10714 18136 10760
rect 18182 10714 18375 10760
rect 18055 10666 18375 10714
rect 18055 10620 18136 10666
rect 18182 10620 18375 10666
rect 18055 10572 18375 10620
rect 18055 10526 18136 10572
rect 18182 10526 18375 10572
rect 18055 10478 18375 10526
rect 18055 10432 18136 10478
rect 18182 10432 18375 10478
rect 18055 10384 18375 10432
rect 18055 10338 18136 10384
rect 18182 10338 18375 10384
rect 18055 10290 18375 10338
rect 18055 10244 18136 10290
rect 18182 10244 18375 10290
rect 18055 10196 18375 10244
rect 18055 10150 18136 10196
rect 18182 10150 18375 10196
rect 18055 10102 18375 10150
rect 18055 10056 18136 10102
rect 18182 10056 18375 10102
rect 18055 10008 18375 10056
rect 18055 9962 18136 10008
rect 18182 9962 18375 10008
rect 18055 9914 18375 9962
rect 18055 9868 18136 9914
rect 18182 9868 18375 9914
rect 18055 9820 18375 9868
rect 18055 9774 18136 9820
rect 18182 9774 18375 9820
rect 18055 9726 18375 9774
rect 18055 9680 18136 9726
rect 18182 9680 18375 9726
rect 18055 9632 18375 9680
rect 18055 9586 18136 9632
rect 18182 9586 18375 9632
rect 18055 9538 18375 9586
rect 18055 9492 18136 9538
rect 18182 9492 18375 9538
rect 18055 9444 18375 9492
rect 18055 9398 18136 9444
rect 18182 9398 18375 9444
rect 18055 9350 18375 9398
rect 18055 9304 18136 9350
rect 18182 9304 18375 9350
rect 18055 9256 18375 9304
rect 18055 9210 18136 9256
rect 18182 9210 18375 9256
rect 18055 9162 18375 9210
rect 18055 9116 18136 9162
rect 18182 9116 18375 9162
rect 18055 9068 18375 9116
rect 18055 9022 18136 9068
rect 18182 9022 18375 9068
rect 18055 8974 18375 9022
rect 18055 8928 18136 8974
rect 18182 8928 18375 8974
rect 18055 8880 18375 8928
rect 18055 8834 18136 8880
rect 18182 8834 18375 8880
rect 18055 8786 18375 8834
rect 18055 8740 18136 8786
rect 18182 8740 18375 8786
rect 18055 8692 18375 8740
rect 18055 8646 18136 8692
rect 18182 8646 18375 8692
rect 18055 8598 18375 8646
rect 18055 8552 18136 8598
rect 18182 8552 18375 8598
rect 18055 8504 18375 8552
rect 18055 8458 18136 8504
rect 18182 8458 18375 8504
rect 18055 8410 18375 8458
rect 18055 8364 18136 8410
rect 18182 8364 18375 8410
rect 18055 8316 18375 8364
rect 18055 8270 18136 8316
rect 18182 8270 18375 8316
rect 18055 8222 18375 8270
rect 18055 8176 18136 8222
rect 18182 8176 18375 8222
rect 18055 8128 18375 8176
rect 18055 8082 18136 8128
rect 18182 8082 18375 8128
rect 18055 8034 18375 8082
rect 18055 7988 18136 8034
rect 18182 7988 18375 8034
rect 18055 7940 18375 7988
rect 18055 7894 18136 7940
rect 18182 7894 18375 7940
rect 18055 7846 18375 7894
rect 18055 7800 18136 7846
rect 18182 7800 18375 7846
rect 18055 7752 18375 7800
rect 18055 7706 18136 7752
rect 18182 7706 18375 7752
rect 18055 7658 18375 7706
rect 18055 7612 18136 7658
rect 18182 7612 18375 7658
rect 18055 7564 18375 7612
rect 16943 7512 17059 7541
rect 16943 7466 16976 7512
rect 17022 7466 17059 7512
rect 16943 7418 17059 7466
rect 16943 7381 16976 7418
rect 14672 7372 16976 7381
rect 17022 7372 17059 7418
rect 11867 7324 17059 7372
rect 11867 7278 11900 7324
rect 11946 7278 11994 7324
rect 12040 7278 12088 7324
rect 12134 7278 12182 7324
rect 12228 7278 12276 7324
rect 12322 7278 12370 7324
rect 12416 7278 12464 7324
rect 12510 7278 12558 7324
rect 12604 7278 12652 7324
rect 12698 7278 12746 7324
rect 12792 7278 12840 7324
rect 12886 7278 12934 7324
rect 12980 7278 13028 7324
rect 13074 7278 13122 7324
rect 13168 7278 13216 7324
rect 13262 7278 13310 7324
rect 13356 7278 13404 7324
rect 13450 7278 13498 7324
rect 13544 7278 13592 7324
rect 13638 7278 13686 7324
rect 13732 7278 13780 7324
rect 13826 7278 13874 7324
rect 13920 7278 13968 7324
rect 14014 7278 14062 7324
rect 14108 7278 14156 7324
rect 14202 7278 14250 7324
rect 14296 7278 14344 7324
rect 14390 7278 14438 7324
rect 14484 7278 14532 7324
rect 14578 7278 14626 7324
rect 14672 7278 14720 7324
rect 14766 7278 14814 7324
rect 14860 7278 14908 7324
rect 14954 7278 15002 7324
rect 15048 7278 15096 7324
rect 15142 7278 15190 7324
rect 15236 7278 15284 7324
rect 15330 7278 15378 7324
rect 15424 7278 15472 7324
rect 15518 7278 15566 7324
rect 15612 7278 15660 7324
rect 15706 7278 15754 7324
rect 15800 7278 15848 7324
rect 15894 7278 15942 7324
rect 15988 7278 16036 7324
rect 16082 7278 16130 7324
rect 16176 7278 16224 7324
rect 16270 7278 16318 7324
rect 16364 7278 16412 7324
rect 16458 7278 16506 7324
rect 16552 7278 16600 7324
rect 16646 7278 16694 7324
rect 16740 7278 16788 7324
rect 16834 7278 16882 7324
rect 16928 7278 16976 7324
rect 17022 7278 17059 7324
rect 11867 7221 17059 7278
rect 18055 7518 18136 7564
rect 18182 7541 18375 7564
rect 18712 13176 18758 13557
rect 18712 12444 18758 12602
rect 18872 13176 18918 13557
rect 19065 13405 19141 13417
rect 19065 13353 19077 13405
rect 19129 13402 19141 13405
rect 20185 13405 20261 13417
rect 20185 13402 20197 13405
rect 19129 13356 19560 13402
rect 19606 13356 20197 13402
rect 19129 13353 19141 13356
rect 19065 13341 19141 13353
rect 20185 13353 20197 13356
rect 20249 13353 20261 13405
rect 20185 13341 20261 13353
rect 19000 13176 19046 13187
rect 18985 12770 19000 12782
rect 19160 13176 19206 13187
rect 19320 13176 19366 13187
rect 19480 13176 19526 13187
rect 19046 12770 19061 12782
rect 18985 12718 18997 12770
rect 19049 12718 19061 12770
rect 18985 12666 19000 12718
rect 19046 12666 19061 12718
rect 18985 12614 18997 12666
rect 19049 12614 19061 12666
rect 18985 12602 19000 12614
rect 19046 12602 19061 12614
rect 19145 12770 19160 12782
rect 19305 13164 19320 13176
rect 19366 13164 19381 13176
rect 19305 13112 19317 13164
rect 19369 13112 19381 13164
rect 19305 13060 19320 13112
rect 19366 13060 19381 13112
rect 19305 13008 19317 13060
rect 19369 13008 19381 13060
rect 19305 12996 19320 13008
rect 19206 12770 19221 12782
rect 19145 12718 19157 12770
rect 19209 12718 19221 12770
rect 19145 12666 19160 12718
rect 19206 12666 19221 12718
rect 19145 12614 19157 12666
rect 19209 12614 19221 12666
rect 19145 12602 19160 12614
rect 19206 12602 19221 12614
rect 19366 12996 19381 13008
rect 19465 12770 19480 12782
rect 19640 13176 19686 13187
rect 19526 12770 19541 12782
rect 19465 12718 19477 12770
rect 19529 12718 19541 12770
rect 19465 12666 19480 12718
rect 19526 12666 19541 12718
rect 19465 12614 19477 12666
rect 19529 12614 19541 12666
rect 19465 12602 19480 12614
rect 19526 12602 19541 12614
rect 19625 12770 19640 12782
rect 19800 13176 19846 13187
rect 19960 13176 20006 13187
rect 20120 13176 20166 13187
rect 19686 12770 19701 12782
rect 19625 12718 19637 12770
rect 19689 12718 19701 12770
rect 19625 12666 19640 12718
rect 19686 12666 19701 12718
rect 19625 12614 19637 12666
rect 19689 12614 19701 12666
rect 19625 12602 19640 12614
rect 19686 12602 19701 12614
rect 19785 12770 19800 12782
rect 19945 13164 19960 13176
rect 20006 13164 20021 13176
rect 19945 13112 19957 13164
rect 20009 13112 20021 13164
rect 19945 13060 19960 13112
rect 20006 13060 20021 13112
rect 19945 13008 19957 13060
rect 20009 13008 20021 13060
rect 19945 12996 19960 13008
rect 19846 12770 19861 12782
rect 19785 12718 19797 12770
rect 19849 12718 19861 12770
rect 19785 12666 19800 12718
rect 19846 12666 19861 12718
rect 19785 12614 19797 12666
rect 19849 12614 19861 12666
rect 19785 12602 19800 12614
rect 19846 12602 19861 12614
rect 20006 12996 20021 13008
rect 20105 12770 20120 12782
rect 20280 13176 20326 13187
rect 20166 12770 20181 12782
rect 20105 12718 20117 12770
rect 20169 12718 20181 12770
rect 20105 12666 20120 12718
rect 20166 12666 20181 12718
rect 20105 12614 20117 12666
rect 20169 12614 20181 12666
rect 20105 12602 20120 12614
rect 20166 12602 20181 12614
rect 20265 12770 20280 12782
rect 20408 13176 20454 13557
rect 20326 12770 20341 12782
rect 20265 12718 20277 12770
rect 20329 12718 20341 12770
rect 20265 12666 20280 12718
rect 20326 12666 20341 12718
rect 20265 12614 20277 12666
rect 20329 12614 20341 12666
rect 20265 12602 20280 12614
rect 20326 12602 20341 12614
rect 18872 12444 18918 12602
rect 19000 12591 19046 12602
rect 19160 12543 19206 12602
rect 19320 12591 19366 12602
rect 19480 12543 19526 12602
rect 19640 12591 19686 12602
rect 19800 12591 19846 12602
rect 19960 12591 20006 12602
rect 20120 12591 20166 12602
rect 20280 12591 20326 12602
rect 19160 12497 19526 12543
rect 18712 12398 18792 12444
rect 18838 12398 18918 12444
rect 18712 12240 18758 12398
rect 18712 11304 18758 11666
rect 18712 10368 18758 10730
rect 18712 9432 18758 9794
rect 18712 8700 18758 8858
rect 18872 12240 18918 12398
rect 19065 12439 19141 12451
rect 19065 12387 19077 12439
rect 19129 12436 19141 12439
rect 20408 12444 20454 12602
rect 20568 13176 20614 13557
rect 20568 12444 20614 12602
rect 19129 12390 19240 12436
rect 19286 12390 19560 12436
rect 19606 12390 19880 12436
rect 19926 12390 20200 12436
rect 20246 12390 20257 12436
rect 20408 12398 20488 12444
rect 20534 12398 20614 12444
rect 19129 12387 19141 12390
rect 19065 12375 19141 12387
rect 19000 12240 19046 12251
rect 18985 11834 19000 11846
rect 19160 12240 19206 12251
rect 19320 12240 19366 12251
rect 19480 12240 19526 12251
rect 19046 11834 19061 11846
rect 18985 11782 18997 11834
rect 19049 11782 19061 11834
rect 18985 11730 19000 11782
rect 19046 11730 19061 11782
rect 18985 11678 18997 11730
rect 19049 11678 19061 11730
rect 18985 11666 19000 11678
rect 19046 11666 19061 11678
rect 19145 11834 19160 11846
rect 19305 12228 19320 12240
rect 19366 12228 19381 12240
rect 19305 12176 19317 12228
rect 19369 12176 19381 12228
rect 19305 12124 19320 12176
rect 19366 12124 19381 12176
rect 19305 12072 19317 12124
rect 19369 12072 19381 12124
rect 19305 12060 19320 12072
rect 19206 11834 19221 11846
rect 19145 11782 19157 11834
rect 19209 11782 19221 11834
rect 19145 11730 19160 11782
rect 19206 11730 19221 11782
rect 19145 11678 19157 11730
rect 19209 11678 19221 11730
rect 19145 11666 19160 11678
rect 19206 11666 19221 11678
rect 19366 12060 19381 12072
rect 19465 11834 19480 11846
rect 19640 12240 19686 12251
rect 19526 11834 19541 11846
rect 19465 11782 19477 11834
rect 19529 11782 19541 11834
rect 19465 11730 19480 11782
rect 19526 11730 19541 11782
rect 19465 11678 19477 11730
rect 19529 11678 19541 11730
rect 19465 11666 19480 11678
rect 19526 11666 19541 11678
rect 19625 11834 19640 11846
rect 19800 12240 19846 12251
rect 19960 12240 20006 12251
rect 20120 12240 20166 12251
rect 19686 11834 19701 11846
rect 19625 11782 19637 11834
rect 19689 11782 19701 11834
rect 19625 11730 19640 11782
rect 19686 11730 19701 11782
rect 19625 11678 19637 11730
rect 19689 11678 19701 11730
rect 19625 11666 19640 11678
rect 19686 11666 19701 11678
rect 19785 11834 19800 11846
rect 19945 12228 19960 12240
rect 20006 12228 20021 12240
rect 19945 12176 19957 12228
rect 20009 12176 20021 12228
rect 19945 12124 19960 12176
rect 20006 12124 20021 12176
rect 19945 12072 19957 12124
rect 20009 12072 20021 12124
rect 19945 12060 19960 12072
rect 19846 11834 19861 11846
rect 19785 11782 19797 11834
rect 19849 11782 19861 11834
rect 19785 11730 19800 11782
rect 19846 11730 19861 11782
rect 19785 11678 19797 11730
rect 19849 11678 19861 11730
rect 19785 11666 19800 11678
rect 19846 11666 19861 11678
rect 20006 12060 20021 12072
rect 20105 11834 20120 11846
rect 20280 12240 20326 12251
rect 20166 11834 20181 11846
rect 20105 11782 20117 11834
rect 20169 11782 20181 11834
rect 20105 11730 20120 11782
rect 20166 11730 20181 11782
rect 20105 11678 20117 11730
rect 20169 11678 20181 11730
rect 20105 11666 20120 11678
rect 20166 11666 20181 11678
rect 20265 11834 20280 11846
rect 20408 12240 20454 12398
rect 20326 11834 20341 11846
rect 20265 11782 20277 11834
rect 20329 11782 20341 11834
rect 20265 11730 20280 11782
rect 20326 11730 20341 11782
rect 20265 11678 20277 11730
rect 20329 11678 20341 11730
rect 20265 11666 20280 11678
rect 20326 11666 20341 11678
rect 18872 11304 18918 11666
rect 19000 11655 19046 11666
rect 19160 11607 19206 11666
rect 19320 11655 19366 11666
rect 19480 11607 19526 11666
rect 19640 11655 19686 11666
rect 19800 11655 19846 11666
rect 19960 11655 20006 11666
rect 20120 11655 20166 11666
rect 20280 11655 20326 11666
rect 19160 11561 19526 11607
rect 19065 11503 19141 11515
rect 19065 11451 19077 11503
rect 19129 11500 19141 11503
rect 19129 11454 19240 11500
rect 19286 11454 19560 11500
rect 19606 11454 19880 11500
rect 19926 11454 20200 11500
rect 20246 11454 20257 11500
rect 19129 11451 19141 11454
rect 19065 11439 19141 11451
rect 19000 11304 19046 11315
rect 18985 10898 19000 10910
rect 19160 11304 19206 11315
rect 19320 11304 19366 11315
rect 19480 11304 19526 11315
rect 19046 10898 19061 10910
rect 18985 10846 18997 10898
rect 19049 10846 19061 10898
rect 18985 10794 19000 10846
rect 19046 10794 19061 10846
rect 18985 10742 18997 10794
rect 19049 10742 19061 10794
rect 18985 10730 19000 10742
rect 19046 10730 19061 10742
rect 19145 10898 19160 10910
rect 19305 11292 19320 11304
rect 19366 11292 19381 11304
rect 19305 11240 19317 11292
rect 19369 11240 19381 11292
rect 19305 11188 19320 11240
rect 19366 11188 19381 11240
rect 19305 11136 19317 11188
rect 19369 11136 19381 11188
rect 19305 11124 19320 11136
rect 19206 10898 19221 10910
rect 19145 10846 19157 10898
rect 19209 10846 19221 10898
rect 19145 10794 19160 10846
rect 19206 10794 19221 10846
rect 19145 10742 19157 10794
rect 19209 10742 19221 10794
rect 19145 10730 19160 10742
rect 19206 10730 19221 10742
rect 19366 11124 19381 11136
rect 19465 10898 19480 10910
rect 19640 11304 19686 11315
rect 19526 10898 19541 10910
rect 19465 10846 19477 10898
rect 19529 10846 19541 10898
rect 19465 10794 19480 10846
rect 19526 10794 19541 10846
rect 19465 10742 19477 10794
rect 19529 10742 19541 10794
rect 19465 10730 19480 10742
rect 19526 10730 19541 10742
rect 19625 10898 19640 10910
rect 19800 11304 19846 11315
rect 19960 11304 20006 11315
rect 20120 11304 20166 11315
rect 19686 10898 19701 10910
rect 19625 10846 19637 10898
rect 19689 10846 19701 10898
rect 19625 10794 19640 10846
rect 19686 10794 19701 10846
rect 19625 10742 19637 10794
rect 19689 10742 19701 10794
rect 19625 10730 19640 10742
rect 19686 10730 19701 10742
rect 19785 10898 19800 10910
rect 19945 11292 19960 11304
rect 20006 11292 20021 11304
rect 19945 11240 19957 11292
rect 20009 11240 20021 11292
rect 19945 11188 19960 11240
rect 20006 11188 20021 11240
rect 19945 11136 19957 11188
rect 20009 11136 20021 11188
rect 19945 11124 19960 11136
rect 19846 10898 19861 10910
rect 19785 10846 19797 10898
rect 19849 10846 19861 10898
rect 19785 10794 19800 10846
rect 19846 10794 19861 10846
rect 19785 10742 19797 10794
rect 19849 10742 19861 10794
rect 19785 10730 19800 10742
rect 19846 10730 19861 10742
rect 20006 11124 20021 11136
rect 20105 10898 20120 10910
rect 20280 11304 20326 11315
rect 20166 10898 20181 10910
rect 20105 10846 20117 10898
rect 20169 10846 20181 10898
rect 20105 10794 20120 10846
rect 20166 10794 20181 10846
rect 20105 10742 20117 10794
rect 20169 10742 20181 10794
rect 20105 10730 20120 10742
rect 20166 10730 20181 10742
rect 20265 10898 20280 10910
rect 20408 11304 20454 11666
rect 20326 10898 20341 10910
rect 20265 10846 20277 10898
rect 20329 10846 20341 10898
rect 20265 10794 20280 10846
rect 20326 10794 20341 10846
rect 20265 10742 20277 10794
rect 20329 10742 20341 10794
rect 20265 10730 20280 10742
rect 20326 10730 20341 10742
rect 18872 10368 18918 10730
rect 19000 10368 19046 10730
rect 18985 9962 19000 9974
rect 19160 10368 19206 10730
rect 19320 10368 19366 10730
rect 19480 10368 19526 10730
rect 19046 9962 19061 9974
rect 18985 9910 18997 9962
rect 19049 9910 19061 9962
rect 18985 9858 19000 9910
rect 19046 9858 19061 9910
rect 18985 9806 18997 9858
rect 19049 9806 19061 9858
rect 18985 9794 19000 9806
rect 19046 9794 19061 9806
rect 19305 10356 19320 10368
rect 19366 10356 19381 10368
rect 19305 10304 19317 10356
rect 19369 10304 19381 10356
rect 19305 10252 19320 10304
rect 19366 10252 19381 10304
rect 19305 10200 19317 10252
rect 19369 10200 19381 10252
rect 19305 10188 19320 10200
rect 18872 9432 18918 9794
rect 19000 9783 19046 9794
rect 19160 9735 19206 9794
rect 19366 10188 19381 10200
rect 19320 9783 19366 9794
rect 19640 10368 19686 10730
rect 19625 9962 19640 9974
rect 19800 10368 19846 10730
rect 19960 10368 20006 10730
rect 20120 10368 20166 10730
rect 19686 9962 19701 9974
rect 19625 9910 19637 9962
rect 19689 9910 19701 9962
rect 19625 9858 19640 9910
rect 19686 9858 19701 9910
rect 19625 9806 19637 9858
rect 19689 9806 19701 9858
rect 19625 9794 19640 9806
rect 19686 9794 19701 9806
rect 19945 10356 19960 10368
rect 20006 10356 20021 10368
rect 19945 10304 19957 10356
rect 20009 10304 20021 10356
rect 19945 10252 19960 10304
rect 20006 10252 20021 10304
rect 19945 10200 19957 10252
rect 20009 10200 20021 10252
rect 19945 10188 19960 10200
rect 19480 9735 19526 9794
rect 19640 9783 19686 9794
rect 19800 9783 19846 9794
rect 20006 10188 20021 10200
rect 19960 9783 20006 9794
rect 20280 10368 20326 10730
rect 20265 9962 20280 9974
rect 20408 10368 20454 10730
rect 20326 9962 20341 9974
rect 20265 9910 20277 9962
rect 20329 9910 20341 9962
rect 20265 9858 20280 9910
rect 20326 9858 20341 9910
rect 20265 9806 20277 9858
rect 20329 9806 20341 9858
rect 20265 9794 20280 9806
rect 20326 9794 20341 9806
rect 20120 9783 20166 9794
rect 20280 9783 20326 9794
rect 19160 9689 19526 9735
rect 19065 9631 19141 9643
rect 19065 9579 19077 9631
rect 19129 9628 19141 9631
rect 19129 9582 19240 9628
rect 19286 9582 19560 9628
rect 19606 9582 19880 9628
rect 19926 9582 20200 9628
rect 20246 9582 20257 9628
rect 19129 9579 19141 9582
rect 19065 9567 19141 9579
rect 19000 9432 19046 9443
rect 18985 9026 19000 9038
rect 19160 9432 19206 9443
rect 19320 9432 19366 9443
rect 19480 9432 19526 9443
rect 19046 9026 19061 9038
rect 18985 8974 18997 9026
rect 19049 8974 19061 9026
rect 18985 8922 19000 8974
rect 19046 8922 19061 8974
rect 18985 8870 18997 8922
rect 19049 8870 19061 8922
rect 18985 8858 19000 8870
rect 19046 8858 19061 8870
rect 19145 9026 19160 9038
rect 19305 9420 19320 9432
rect 19366 9420 19381 9432
rect 19305 9368 19317 9420
rect 19369 9368 19381 9420
rect 19305 9316 19320 9368
rect 19366 9316 19381 9368
rect 19305 9264 19317 9316
rect 19369 9264 19381 9316
rect 19305 9252 19320 9264
rect 19206 9026 19221 9038
rect 19145 8974 19157 9026
rect 19209 8974 19221 9026
rect 19145 8922 19160 8974
rect 19206 8922 19221 8974
rect 19145 8870 19157 8922
rect 19209 8870 19221 8922
rect 19145 8858 19160 8870
rect 19206 8858 19221 8870
rect 19366 9252 19381 9264
rect 19465 9026 19480 9038
rect 19640 9432 19686 9443
rect 19526 9026 19541 9038
rect 19465 8974 19477 9026
rect 19529 8974 19541 9026
rect 19465 8922 19480 8974
rect 19526 8922 19541 8974
rect 19465 8870 19477 8922
rect 19529 8870 19541 8922
rect 19465 8858 19480 8870
rect 19526 8858 19541 8870
rect 19625 9026 19640 9038
rect 19800 9432 19846 9443
rect 19960 9432 20006 9443
rect 20120 9432 20166 9443
rect 19686 9026 19701 9038
rect 19625 8974 19637 9026
rect 19689 8974 19701 9026
rect 19625 8922 19640 8974
rect 19686 8922 19701 8974
rect 19625 8870 19637 8922
rect 19689 8870 19701 8922
rect 19625 8858 19640 8870
rect 19686 8858 19701 8870
rect 19785 9026 19800 9038
rect 19945 9420 19960 9432
rect 20006 9420 20021 9432
rect 19945 9368 19957 9420
rect 20009 9368 20021 9420
rect 19945 9316 19960 9368
rect 20006 9316 20021 9368
rect 19945 9264 19957 9316
rect 20009 9264 20021 9316
rect 19945 9252 19960 9264
rect 19846 9026 19861 9038
rect 19785 8974 19797 9026
rect 19849 8974 19861 9026
rect 19785 8922 19800 8974
rect 19846 8922 19861 8974
rect 19785 8870 19797 8922
rect 19849 8870 19861 8922
rect 19785 8858 19800 8870
rect 19846 8858 19861 8870
rect 20006 9252 20021 9264
rect 20105 9026 20120 9038
rect 20280 9432 20326 9443
rect 20166 9026 20181 9038
rect 20105 8974 20117 9026
rect 20169 8974 20181 9026
rect 20105 8922 20120 8974
rect 20166 8922 20181 8974
rect 20105 8870 20117 8922
rect 20169 8870 20181 8922
rect 20105 8858 20120 8870
rect 20166 8858 20181 8870
rect 20265 9026 20280 9038
rect 20408 9432 20454 9794
rect 20326 9026 20341 9038
rect 20265 8974 20277 9026
rect 20329 8974 20341 9026
rect 20265 8922 20280 8974
rect 20326 8922 20341 8974
rect 20265 8870 20277 8922
rect 20329 8870 20341 8922
rect 20265 8858 20280 8870
rect 20326 8858 20341 8870
rect 18872 8700 18918 8858
rect 19000 8847 19046 8858
rect 19160 8799 19206 8858
rect 19320 8847 19366 8858
rect 19480 8799 19526 8858
rect 19640 8847 19686 8858
rect 19800 8847 19846 8858
rect 19960 8847 20006 8858
rect 20120 8847 20166 8858
rect 20280 8847 20326 8858
rect 19160 8753 19526 8799
rect 18712 8654 18792 8700
rect 18838 8654 18918 8700
rect 18712 8496 18758 8654
rect 18712 7541 18758 7922
rect 18872 8496 18918 8654
rect 19065 8695 19141 8707
rect 19065 8643 19077 8695
rect 19129 8692 19141 8695
rect 20408 8700 20454 8858
rect 20568 12240 20614 12398
rect 20568 11304 20614 11666
rect 20568 10368 20614 10730
rect 20568 9432 20614 9794
rect 20568 8700 20614 8858
rect 19129 8646 19240 8692
rect 19286 8646 19560 8692
rect 19606 8646 19880 8692
rect 19926 8646 20200 8692
rect 20246 8646 20257 8692
rect 20408 8654 20488 8700
rect 20534 8654 20614 8700
rect 19129 8643 19141 8646
rect 19065 8631 19141 8643
rect 19000 8496 19046 8507
rect 18985 8090 19000 8102
rect 19160 8496 19206 8507
rect 19320 8496 19366 8507
rect 19480 8496 19526 8507
rect 19046 8090 19061 8102
rect 18985 8038 18997 8090
rect 19049 8038 19061 8090
rect 18985 7986 19000 8038
rect 19046 7986 19061 8038
rect 18985 7934 18997 7986
rect 19049 7934 19061 7986
rect 18985 7922 19000 7934
rect 19046 7922 19061 7934
rect 19145 8090 19160 8102
rect 19305 8484 19320 8496
rect 19366 8484 19381 8496
rect 19305 8432 19317 8484
rect 19369 8432 19381 8484
rect 19305 8380 19320 8432
rect 19366 8380 19381 8432
rect 19305 8328 19317 8380
rect 19369 8328 19381 8380
rect 19305 8316 19320 8328
rect 19206 8090 19221 8102
rect 19145 8038 19157 8090
rect 19209 8038 19221 8090
rect 19145 7986 19160 8038
rect 19206 7986 19221 8038
rect 19145 7934 19157 7986
rect 19209 7934 19221 7986
rect 19145 7922 19160 7934
rect 19206 7922 19221 7934
rect 19366 8316 19381 8328
rect 19465 8090 19480 8102
rect 19640 8496 19686 8507
rect 19526 8090 19541 8102
rect 19465 8038 19477 8090
rect 19529 8038 19541 8090
rect 19465 7986 19480 8038
rect 19526 7986 19541 8038
rect 19465 7934 19477 7986
rect 19529 7934 19541 7986
rect 19465 7922 19480 7934
rect 19526 7922 19541 7934
rect 19625 8090 19640 8102
rect 19800 8496 19846 8507
rect 19960 8496 20006 8507
rect 20120 8496 20166 8507
rect 19686 8090 19701 8102
rect 19625 8038 19637 8090
rect 19689 8038 19701 8090
rect 19625 7986 19640 8038
rect 19686 7986 19701 8038
rect 19625 7934 19637 7986
rect 19689 7934 19701 7986
rect 19625 7922 19640 7934
rect 19686 7922 19701 7934
rect 19785 8090 19800 8102
rect 19945 8484 19960 8496
rect 20006 8484 20021 8496
rect 19945 8432 19957 8484
rect 20009 8432 20021 8484
rect 19945 8380 19960 8432
rect 20006 8380 20021 8432
rect 19945 8328 19957 8380
rect 20009 8328 20021 8380
rect 19945 8316 19960 8328
rect 19846 8090 19861 8102
rect 19785 8038 19797 8090
rect 19849 8038 19861 8090
rect 19785 7986 19800 8038
rect 19846 7986 19861 8038
rect 19785 7934 19797 7986
rect 19849 7934 19861 7986
rect 19785 7922 19800 7934
rect 19846 7922 19861 7934
rect 20006 8316 20021 8328
rect 20105 8090 20120 8102
rect 20280 8496 20326 8507
rect 20166 8090 20181 8102
rect 20105 8038 20117 8090
rect 20169 8038 20181 8090
rect 20105 7986 20120 8038
rect 20166 7986 20181 8038
rect 20105 7934 20117 7986
rect 20169 7934 20181 7986
rect 20105 7922 20120 7934
rect 20166 7922 20181 7934
rect 20265 8090 20280 8102
rect 20408 8496 20454 8654
rect 20326 8090 20341 8102
rect 20265 8038 20277 8090
rect 20329 8038 20341 8090
rect 20265 7986 20280 8038
rect 20326 7986 20341 8038
rect 20265 7934 20277 7986
rect 20329 7934 20341 7986
rect 20265 7922 20280 7934
rect 20326 7922 20341 7934
rect 18872 7541 18918 7922
rect 19000 7911 19046 7922
rect 19160 7863 19206 7922
rect 19320 7911 19366 7922
rect 19480 7863 19526 7922
rect 19640 7911 19686 7922
rect 19800 7863 19846 7922
rect 19960 7911 20006 7922
rect 20120 7863 20166 7922
rect 20280 7911 20326 7922
rect 19160 7817 20166 7863
rect 19225 7759 19301 7771
rect 19225 7707 19237 7759
rect 19289 7756 19301 7759
rect 19865 7759 19941 7771
rect 19865 7756 19877 7759
rect 19289 7710 19877 7756
rect 19289 7707 19301 7710
rect 19225 7695 19301 7707
rect 19865 7707 19877 7710
rect 19929 7707 19941 7759
rect 19865 7695 19941 7707
rect 20120 7541 20166 7817
rect 20408 7541 20454 7922
rect 20568 8496 20614 8654
rect 20568 7541 20614 7922
rect 20951 13534 21144 13557
rect 21190 13557 23288 13580
rect 21190 13534 21271 13557
rect 20951 13486 21271 13534
rect 20951 13440 21144 13486
rect 21190 13440 21271 13486
rect 20951 13392 21271 13440
rect 20951 13346 21144 13392
rect 21190 13346 21271 13392
rect 20951 13298 21271 13346
rect 20951 13252 21144 13298
rect 21190 13252 21271 13298
rect 20951 13204 21271 13252
rect 20951 13158 21144 13204
rect 21190 13158 21271 13204
rect 20951 13110 21271 13158
rect 20951 13064 21144 13110
rect 21190 13064 21271 13110
rect 20951 13016 21271 13064
rect 20951 12970 21144 13016
rect 21190 12970 21271 13016
rect 20951 12922 21271 12970
rect 20951 12876 21144 12922
rect 21190 12876 21271 12922
rect 20951 12828 21271 12876
rect 20951 12782 21144 12828
rect 21190 12782 21271 12828
rect 20951 12734 21271 12782
rect 20951 12688 21144 12734
rect 21190 12688 21271 12734
rect 20951 12640 21271 12688
rect 20951 12594 21144 12640
rect 21190 12594 21271 12640
rect 20951 12546 21271 12594
rect 20951 12500 21144 12546
rect 21190 12500 21271 12546
rect 20951 12452 21271 12500
rect 20951 12406 21144 12452
rect 21190 12406 21271 12452
rect 20951 12358 21271 12406
rect 20951 12312 21144 12358
rect 21190 12312 21271 12358
rect 20951 12264 21271 12312
rect 20951 12218 21144 12264
rect 21190 12218 21271 12264
rect 20951 12170 21271 12218
rect 20951 12124 21144 12170
rect 21190 12124 21271 12170
rect 20951 12076 21271 12124
rect 20951 12030 21144 12076
rect 21190 12030 21271 12076
rect 20951 11982 21271 12030
rect 20951 11936 21144 11982
rect 21190 11936 21271 11982
rect 20951 11888 21271 11936
rect 20951 11842 21144 11888
rect 21190 11842 21271 11888
rect 20951 11794 21271 11842
rect 20951 11748 21144 11794
rect 21190 11748 21271 11794
rect 20951 11700 21271 11748
rect 20951 11654 21144 11700
rect 21190 11654 21271 11700
rect 20951 11606 21271 11654
rect 20951 11560 21144 11606
rect 21190 11560 21271 11606
rect 20951 11512 21271 11560
rect 20951 11466 21144 11512
rect 21190 11466 21271 11512
rect 20951 11418 21271 11466
rect 20951 11372 21144 11418
rect 21190 11372 21271 11418
rect 20951 11324 21271 11372
rect 20951 11278 21144 11324
rect 21190 11278 21271 11324
rect 20951 11230 21271 11278
rect 20951 11184 21144 11230
rect 21190 11184 21271 11230
rect 20951 11136 21271 11184
rect 20951 11090 21144 11136
rect 21190 11090 21271 11136
rect 20951 11042 21271 11090
rect 20951 10996 21144 11042
rect 21190 10996 21271 11042
rect 20951 10948 21271 10996
rect 20951 10902 21144 10948
rect 21190 10902 21271 10948
rect 20951 10854 21271 10902
rect 20951 10808 21144 10854
rect 21190 10808 21271 10854
rect 20951 10760 21271 10808
rect 20951 10714 21144 10760
rect 21190 10714 21271 10760
rect 20951 10666 21271 10714
rect 20951 10620 21144 10666
rect 21190 10620 21271 10666
rect 20951 10572 21271 10620
rect 20951 10526 21144 10572
rect 21190 10526 21271 10572
rect 20951 10478 21271 10526
rect 20951 10432 21144 10478
rect 21190 10432 21271 10478
rect 20951 10384 21271 10432
rect 20951 10338 21144 10384
rect 21190 10338 21271 10384
rect 20951 10290 21271 10338
rect 20951 10244 21144 10290
rect 21190 10244 21271 10290
rect 20951 10196 21271 10244
rect 20951 10150 21144 10196
rect 21190 10150 21271 10196
rect 20951 10102 21271 10150
rect 20951 10056 21144 10102
rect 21190 10056 21271 10102
rect 20951 10008 21271 10056
rect 20951 9962 21144 10008
rect 21190 9962 21271 10008
rect 20951 9914 21271 9962
rect 20951 9868 21144 9914
rect 21190 9868 21271 9914
rect 20951 9820 21271 9868
rect 20951 9774 21144 9820
rect 21190 9774 21271 9820
rect 20951 9726 21271 9774
rect 20951 9680 21144 9726
rect 21190 9680 21271 9726
rect 20951 9632 21271 9680
rect 20951 9586 21144 9632
rect 21190 9586 21271 9632
rect 20951 9538 21271 9586
rect 20951 9492 21144 9538
rect 21190 9492 21271 9538
rect 20951 9444 21271 9492
rect 20951 9398 21144 9444
rect 21190 9398 21271 9444
rect 20951 9350 21271 9398
rect 20951 9304 21144 9350
rect 21190 9304 21271 9350
rect 20951 9256 21271 9304
rect 20951 9210 21144 9256
rect 21190 9210 21271 9256
rect 20951 9162 21271 9210
rect 20951 9116 21144 9162
rect 21190 9116 21271 9162
rect 20951 9068 21271 9116
rect 20951 9022 21144 9068
rect 21190 9022 21271 9068
rect 20951 8974 21271 9022
rect 20951 8928 21144 8974
rect 21190 8928 21271 8974
rect 20951 8880 21271 8928
rect 20951 8834 21144 8880
rect 21190 8834 21271 8880
rect 20951 8786 21271 8834
rect 20951 8740 21144 8786
rect 21190 8740 21271 8786
rect 20951 8692 21271 8740
rect 20951 8646 21144 8692
rect 21190 8646 21271 8692
rect 20951 8598 21271 8646
rect 20951 8552 21144 8598
rect 21190 8552 21271 8598
rect 20951 8504 21271 8552
rect 20951 8458 21144 8504
rect 21190 8458 21271 8504
rect 20951 8410 21271 8458
rect 20951 8364 21144 8410
rect 21190 8364 21271 8410
rect 20951 8316 21271 8364
rect 20951 8270 21144 8316
rect 21190 8270 21271 8316
rect 20951 8222 21271 8270
rect 20951 8176 21144 8222
rect 21190 8176 21271 8222
rect 20951 8128 21271 8176
rect 20951 8082 21144 8128
rect 21190 8082 21271 8128
rect 20951 8034 21271 8082
rect 20951 7988 21144 8034
rect 21190 7988 21271 8034
rect 20951 7940 21271 7988
rect 20951 7894 21144 7940
rect 21190 7894 21271 7940
rect 20951 7846 21271 7894
rect 20951 7800 21144 7846
rect 21190 7800 21271 7846
rect 20951 7752 21271 7800
rect 20951 7706 21144 7752
rect 21190 7706 21271 7752
rect 20951 7658 21271 7706
rect 20951 7612 21144 7658
rect 21190 7612 21271 7658
rect 20951 7564 21271 7612
rect 20951 7541 21144 7564
rect 18182 7518 21144 7541
rect 21190 7541 21271 7564
rect 23207 13534 23288 13557
rect 23334 13557 26296 13580
rect 23334 13534 23527 13557
rect 23207 13486 23527 13534
rect 23207 13440 23288 13486
rect 23334 13440 23527 13486
rect 23207 13392 23527 13440
rect 23207 13346 23288 13392
rect 23334 13346 23527 13392
rect 23207 13298 23527 13346
rect 23207 13252 23288 13298
rect 23334 13252 23527 13298
rect 23207 13204 23527 13252
rect 23207 13158 23288 13204
rect 23334 13158 23527 13204
rect 23207 13110 23527 13158
rect 23207 13064 23288 13110
rect 23334 13064 23527 13110
rect 23207 13016 23527 13064
rect 23207 12970 23288 13016
rect 23334 12970 23527 13016
rect 23207 12922 23527 12970
rect 23207 12876 23288 12922
rect 23334 12876 23527 12922
rect 23207 12828 23527 12876
rect 23207 12782 23288 12828
rect 23334 12782 23527 12828
rect 23207 12734 23527 12782
rect 23207 12688 23288 12734
rect 23334 12688 23527 12734
rect 23207 12640 23527 12688
rect 23207 12594 23288 12640
rect 23334 12594 23527 12640
rect 23207 12546 23527 12594
rect 23207 12500 23288 12546
rect 23334 12500 23527 12546
rect 23207 12452 23527 12500
rect 23207 12406 23288 12452
rect 23334 12406 23527 12452
rect 23207 12358 23527 12406
rect 23207 12312 23288 12358
rect 23334 12312 23527 12358
rect 23207 12264 23527 12312
rect 23207 12218 23288 12264
rect 23334 12218 23527 12264
rect 23207 12170 23527 12218
rect 23207 12124 23288 12170
rect 23334 12124 23527 12170
rect 23207 12076 23527 12124
rect 23207 12030 23288 12076
rect 23334 12030 23527 12076
rect 23207 11982 23527 12030
rect 23207 11936 23288 11982
rect 23334 11936 23527 11982
rect 23207 11888 23527 11936
rect 23207 11842 23288 11888
rect 23334 11842 23527 11888
rect 23207 11794 23527 11842
rect 23207 11748 23288 11794
rect 23334 11748 23527 11794
rect 23207 11700 23527 11748
rect 23207 11654 23288 11700
rect 23334 11654 23527 11700
rect 23207 11606 23527 11654
rect 23207 11560 23288 11606
rect 23334 11560 23527 11606
rect 23207 11512 23527 11560
rect 23207 11466 23288 11512
rect 23334 11466 23527 11512
rect 23207 11418 23527 11466
rect 23207 11372 23288 11418
rect 23334 11372 23527 11418
rect 23207 11324 23527 11372
rect 23207 11278 23288 11324
rect 23334 11278 23527 11324
rect 23207 11230 23527 11278
rect 23207 11184 23288 11230
rect 23334 11184 23527 11230
rect 23207 11136 23527 11184
rect 23207 11090 23288 11136
rect 23334 11090 23527 11136
rect 23207 11042 23527 11090
rect 23207 10996 23288 11042
rect 23334 10996 23527 11042
rect 23207 10948 23527 10996
rect 23207 10902 23288 10948
rect 23334 10902 23527 10948
rect 23207 10854 23527 10902
rect 23207 10808 23288 10854
rect 23334 10808 23527 10854
rect 23207 10760 23527 10808
rect 23207 10714 23288 10760
rect 23334 10714 23527 10760
rect 23207 10666 23527 10714
rect 23207 10620 23288 10666
rect 23334 10620 23527 10666
rect 23207 10572 23527 10620
rect 23207 10526 23288 10572
rect 23334 10526 23527 10572
rect 23207 10478 23527 10526
rect 23207 10432 23288 10478
rect 23334 10432 23527 10478
rect 23207 10384 23527 10432
rect 23207 10338 23288 10384
rect 23334 10338 23527 10384
rect 23207 10290 23527 10338
rect 23207 10244 23288 10290
rect 23334 10244 23527 10290
rect 23207 10196 23527 10244
rect 23207 10150 23288 10196
rect 23334 10150 23527 10196
rect 23207 10102 23527 10150
rect 23207 10056 23288 10102
rect 23334 10056 23527 10102
rect 23207 10008 23527 10056
rect 23207 9962 23288 10008
rect 23334 9962 23527 10008
rect 23207 9914 23527 9962
rect 23207 9868 23288 9914
rect 23334 9868 23527 9914
rect 23207 9820 23527 9868
rect 23207 9774 23288 9820
rect 23334 9774 23527 9820
rect 23207 9726 23527 9774
rect 23207 9680 23288 9726
rect 23334 9680 23527 9726
rect 23207 9632 23527 9680
rect 23207 9586 23288 9632
rect 23334 9586 23527 9632
rect 23207 9538 23527 9586
rect 23207 9492 23288 9538
rect 23334 9492 23527 9538
rect 23207 9444 23527 9492
rect 23207 9398 23288 9444
rect 23334 9398 23527 9444
rect 23207 9350 23527 9398
rect 23207 9304 23288 9350
rect 23334 9304 23527 9350
rect 23207 9256 23527 9304
rect 23207 9210 23288 9256
rect 23334 9210 23527 9256
rect 23207 9162 23527 9210
rect 23207 9116 23288 9162
rect 23334 9116 23527 9162
rect 23207 9068 23527 9116
rect 23207 9022 23288 9068
rect 23334 9022 23527 9068
rect 23207 8974 23527 9022
rect 23207 8928 23288 8974
rect 23334 8928 23527 8974
rect 23207 8880 23527 8928
rect 23207 8834 23288 8880
rect 23334 8834 23527 8880
rect 23207 8786 23527 8834
rect 23207 8740 23288 8786
rect 23334 8740 23527 8786
rect 23207 8692 23527 8740
rect 23207 8646 23288 8692
rect 23334 8646 23527 8692
rect 23207 8598 23527 8646
rect 23207 8552 23288 8598
rect 23334 8552 23527 8598
rect 23207 8504 23527 8552
rect 23207 8458 23288 8504
rect 23334 8458 23527 8504
rect 23207 8410 23527 8458
rect 23207 8364 23288 8410
rect 23334 8364 23527 8410
rect 23207 8316 23527 8364
rect 23207 8270 23288 8316
rect 23334 8270 23527 8316
rect 23207 8222 23527 8270
rect 23207 8176 23288 8222
rect 23334 8176 23527 8222
rect 23207 8128 23527 8176
rect 23207 8082 23288 8128
rect 23334 8082 23527 8128
rect 23207 8034 23527 8082
rect 23207 7988 23288 8034
rect 23334 7988 23527 8034
rect 23207 7940 23527 7988
rect 23207 7894 23288 7940
rect 23334 7894 23527 7940
rect 23207 7846 23527 7894
rect 23207 7800 23288 7846
rect 23334 7800 23527 7846
rect 23207 7752 23527 7800
rect 23207 7706 23288 7752
rect 23334 7706 23527 7752
rect 23207 7658 23527 7706
rect 23207 7612 23288 7658
rect 23334 7612 23527 7658
rect 23207 7564 23527 7612
rect 23207 7541 23288 7564
rect 21190 7518 23288 7541
rect 23334 7541 23527 7564
rect 23864 13176 23910 13557
rect 23864 12444 23910 12602
rect 24024 13176 24070 13557
rect 24217 13405 24293 13417
rect 24217 13353 24229 13405
rect 24281 13402 24293 13405
rect 25337 13405 25413 13417
rect 25337 13402 25349 13405
rect 24281 13356 24872 13402
rect 24918 13356 25349 13402
rect 24281 13353 24293 13356
rect 24217 13341 24293 13353
rect 25337 13353 25349 13356
rect 25401 13353 25413 13405
rect 25337 13341 25413 13353
rect 24152 13176 24198 13187
rect 24137 12770 24152 12782
rect 24312 13176 24358 13187
rect 24472 13176 24518 13187
rect 24632 13176 24678 13187
rect 24198 12770 24213 12782
rect 24137 12718 24149 12770
rect 24201 12718 24213 12770
rect 24137 12666 24152 12718
rect 24198 12666 24213 12718
rect 24137 12614 24149 12666
rect 24201 12614 24213 12666
rect 24137 12602 24152 12614
rect 24198 12602 24213 12614
rect 24297 12770 24312 12782
rect 24457 13164 24472 13176
rect 24518 13164 24533 13176
rect 24457 13112 24469 13164
rect 24521 13112 24533 13164
rect 24457 13060 24472 13112
rect 24518 13060 24533 13112
rect 24457 13008 24469 13060
rect 24521 13008 24533 13060
rect 24457 12996 24472 13008
rect 24358 12770 24373 12782
rect 24297 12718 24309 12770
rect 24361 12718 24373 12770
rect 24297 12666 24312 12718
rect 24358 12666 24373 12718
rect 24297 12614 24309 12666
rect 24361 12614 24373 12666
rect 24297 12602 24312 12614
rect 24358 12602 24373 12614
rect 24518 12996 24533 13008
rect 24617 12770 24632 12782
rect 24792 13176 24838 13187
rect 24678 12770 24693 12782
rect 24617 12718 24629 12770
rect 24681 12718 24693 12770
rect 24617 12666 24632 12718
rect 24678 12666 24693 12718
rect 24617 12614 24629 12666
rect 24681 12614 24693 12666
rect 24617 12602 24632 12614
rect 24678 12602 24693 12614
rect 24777 12770 24792 12782
rect 24952 13176 24998 13187
rect 25112 13176 25158 13187
rect 25272 13176 25318 13187
rect 24838 12770 24853 12782
rect 24777 12718 24789 12770
rect 24841 12718 24853 12770
rect 24777 12666 24792 12718
rect 24838 12666 24853 12718
rect 24777 12614 24789 12666
rect 24841 12614 24853 12666
rect 24777 12602 24792 12614
rect 24838 12602 24853 12614
rect 24937 12770 24952 12782
rect 25097 13164 25112 13176
rect 25158 13164 25173 13176
rect 25097 13112 25109 13164
rect 25161 13112 25173 13164
rect 25097 13060 25112 13112
rect 25158 13060 25173 13112
rect 25097 13008 25109 13060
rect 25161 13008 25173 13060
rect 25097 12996 25112 13008
rect 24998 12770 25013 12782
rect 24937 12718 24949 12770
rect 25001 12718 25013 12770
rect 24937 12666 24952 12718
rect 24998 12666 25013 12718
rect 24937 12614 24949 12666
rect 25001 12614 25013 12666
rect 24937 12602 24952 12614
rect 24998 12602 25013 12614
rect 25158 12996 25173 13008
rect 25257 12770 25272 12782
rect 25432 13176 25478 13187
rect 25318 12770 25333 12782
rect 25257 12718 25269 12770
rect 25321 12718 25333 12770
rect 25257 12666 25272 12718
rect 25318 12666 25333 12718
rect 25257 12614 25269 12666
rect 25321 12614 25333 12666
rect 25257 12602 25272 12614
rect 25318 12602 25333 12614
rect 25417 12770 25432 12782
rect 25560 13176 25606 13557
rect 25478 12770 25493 12782
rect 25417 12718 25429 12770
rect 25481 12718 25493 12770
rect 25417 12666 25432 12718
rect 25478 12666 25493 12718
rect 25417 12614 25429 12666
rect 25481 12614 25493 12666
rect 25417 12602 25432 12614
rect 25478 12602 25493 12614
rect 24024 12444 24070 12602
rect 24152 12591 24198 12602
rect 24312 12591 24358 12602
rect 24472 12591 24518 12602
rect 24632 12591 24678 12602
rect 24792 12591 24838 12602
rect 24952 12543 24998 12602
rect 25112 12591 25158 12602
rect 25272 12543 25318 12602
rect 25432 12591 25478 12602
rect 24952 12497 25318 12543
rect 23864 12398 23944 12444
rect 23990 12398 24070 12444
rect 25337 12439 25413 12451
rect 25337 12436 25349 12439
rect 23864 12240 23910 12398
rect 23864 11304 23910 11666
rect 23864 10368 23910 10730
rect 23864 9432 23910 9794
rect 23864 8700 23910 8858
rect 24024 12240 24070 12398
rect 24221 12390 24232 12436
rect 24278 12390 24552 12436
rect 24598 12390 24872 12436
rect 24918 12390 25192 12436
rect 25238 12390 25349 12436
rect 25337 12387 25349 12390
rect 25401 12387 25413 12439
rect 25337 12375 25413 12387
rect 25560 12444 25606 12602
rect 25720 13176 25766 13557
rect 25720 12444 25766 12602
rect 25560 12398 25640 12444
rect 25686 12398 25766 12444
rect 24152 12240 24198 12251
rect 24137 11834 24152 11846
rect 24312 12240 24358 12251
rect 24472 12240 24518 12251
rect 24632 12240 24678 12251
rect 24198 11834 24213 11846
rect 24137 11782 24149 11834
rect 24201 11782 24213 11834
rect 24137 11730 24152 11782
rect 24198 11730 24213 11782
rect 24137 11678 24149 11730
rect 24201 11678 24213 11730
rect 24137 11666 24152 11678
rect 24198 11666 24213 11678
rect 24297 11834 24312 11846
rect 24457 12228 24472 12240
rect 24518 12228 24533 12240
rect 24457 12176 24469 12228
rect 24521 12176 24533 12228
rect 24457 12124 24472 12176
rect 24518 12124 24533 12176
rect 24457 12072 24469 12124
rect 24521 12072 24533 12124
rect 24457 12060 24472 12072
rect 24358 11834 24373 11846
rect 24297 11782 24309 11834
rect 24361 11782 24373 11834
rect 24297 11730 24312 11782
rect 24358 11730 24373 11782
rect 24297 11678 24309 11730
rect 24361 11678 24373 11730
rect 24297 11666 24312 11678
rect 24358 11666 24373 11678
rect 24518 12060 24533 12072
rect 24617 11834 24632 11846
rect 24792 12240 24838 12251
rect 24678 11834 24693 11846
rect 24617 11782 24629 11834
rect 24681 11782 24693 11834
rect 24617 11730 24632 11782
rect 24678 11730 24693 11782
rect 24617 11678 24629 11730
rect 24681 11678 24693 11730
rect 24617 11666 24632 11678
rect 24678 11666 24693 11678
rect 24777 11834 24792 11846
rect 24952 12240 24998 12251
rect 25112 12240 25158 12251
rect 25272 12240 25318 12251
rect 24838 11834 24853 11846
rect 24777 11782 24789 11834
rect 24841 11782 24853 11834
rect 24777 11730 24792 11782
rect 24838 11730 24853 11782
rect 24777 11678 24789 11730
rect 24841 11678 24853 11730
rect 24777 11666 24792 11678
rect 24838 11666 24853 11678
rect 24937 11834 24952 11846
rect 25097 12228 25112 12240
rect 25158 12228 25173 12240
rect 25097 12176 25109 12228
rect 25161 12176 25173 12228
rect 25097 12124 25112 12176
rect 25158 12124 25173 12176
rect 25097 12072 25109 12124
rect 25161 12072 25173 12124
rect 25097 12060 25112 12072
rect 24998 11834 25013 11846
rect 24937 11782 24949 11834
rect 25001 11782 25013 11834
rect 24937 11730 24952 11782
rect 24998 11730 25013 11782
rect 24937 11678 24949 11730
rect 25001 11678 25013 11730
rect 24937 11666 24952 11678
rect 24998 11666 25013 11678
rect 25158 12060 25173 12072
rect 25257 11834 25272 11846
rect 25432 12240 25478 12251
rect 25318 11834 25333 11846
rect 25257 11782 25269 11834
rect 25321 11782 25333 11834
rect 25257 11730 25272 11782
rect 25318 11730 25333 11782
rect 25257 11678 25269 11730
rect 25321 11678 25333 11730
rect 25257 11666 25272 11678
rect 25318 11666 25333 11678
rect 25417 11834 25432 11846
rect 25560 12240 25606 12398
rect 25478 11834 25493 11846
rect 25417 11782 25429 11834
rect 25481 11782 25493 11834
rect 25417 11730 25432 11782
rect 25478 11730 25493 11782
rect 25417 11678 25429 11730
rect 25481 11678 25493 11730
rect 25417 11666 25432 11678
rect 25478 11666 25493 11678
rect 24024 11304 24070 11666
rect 24152 11655 24198 11666
rect 24312 11655 24358 11666
rect 24472 11655 24518 11666
rect 24632 11655 24678 11666
rect 24792 11655 24838 11666
rect 24952 11607 24998 11666
rect 25112 11655 25158 11666
rect 25272 11607 25318 11666
rect 25432 11655 25478 11666
rect 24952 11561 25318 11607
rect 25337 11503 25413 11515
rect 25337 11500 25349 11503
rect 24221 11454 24232 11500
rect 24278 11454 24552 11500
rect 24598 11454 24872 11500
rect 24918 11454 25192 11500
rect 25238 11454 25349 11500
rect 25337 11451 25349 11454
rect 25401 11451 25413 11503
rect 25337 11439 25413 11451
rect 24152 11304 24198 11315
rect 24137 10898 24152 10910
rect 24312 11304 24358 11315
rect 24472 11304 24518 11315
rect 24632 11304 24678 11315
rect 24198 10898 24213 10910
rect 24137 10846 24149 10898
rect 24201 10846 24213 10898
rect 24137 10794 24152 10846
rect 24198 10794 24213 10846
rect 24137 10742 24149 10794
rect 24201 10742 24213 10794
rect 24137 10730 24152 10742
rect 24198 10730 24213 10742
rect 24297 10898 24312 10910
rect 24457 11292 24472 11304
rect 24518 11292 24533 11304
rect 24457 11240 24469 11292
rect 24521 11240 24533 11292
rect 24457 11188 24472 11240
rect 24518 11188 24533 11240
rect 24457 11136 24469 11188
rect 24521 11136 24533 11188
rect 24457 11124 24472 11136
rect 24358 10898 24373 10910
rect 24297 10846 24309 10898
rect 24361 10846 24373 10898
rect 24297 10794 24312 10846
rect 24358 10794 24373 10846
rect 24297 10742 24309 10794
rect 24361 10742 24373 10794
rect 24297 10730 24312 10742
rect 24358 10730 24373 10742
rect 24518 11124 24533 11136
rect 24617 10898 24632 10910
rect 24792 11304 24838 11315
rect 24678 10898 24693 10910
rect 24617 10846 24629 10898
rect 24681 10846 24693 10898
rect 24617 10794 24632 10846
rect 24678 10794 24693 10846
rect 24617 10742 24629 10794
rect 24681 10742 24693 10794
rect 24617 10730 24632 10742
rect 24678 10730 24693 10742
rect 24777 10898 24792 10910
rect 24952 11304 24998 11315
rect 25112 11304 25158 11315
rect 25272 11304 25318 11315
rect 24838 10898 24853 10910
rect 24777 10846 24789 10898
rect 24841 10846 24853 10898
rect 24777 10794 24792 10846
rect 24838 10794 24853 10846
rect 24777 10742 24789 10794
rect 24841 10742 24853 10794
rect 24777 10730 24792 10742
rect 24838 10730 24853 10742
rect 24937 10898 24952 10910
rect 25097 11292 25112 11304
rect 25158 11292 25173 11304
rect 25097 11240 25109 11292
rect 25161 11240 25173 11292
rect 25097 11188 25112 11240
rect 25158 11188 25173 11240
rect 25097 11136 25109 11188
rect 25161 11136 25173 11188
rect 25097 11124 25112 11136
rect 24998 10898 25013 10910
rect 24937 10846 24949 10898
rect 25001 10846 25013 10898
rect 24937 10794 24952 10846
rect 24998 10794 25013 10846
rect 24937 10742 24949 10794
rect 25001 10742 25013 10794
rect 24937 10730 24952 10742
rect 24998 10730 25013 10742
rect 25158 11124 25173 11136
rect 25257 10898 25272 10910
rect 25432 11304 25478 11315
rect 25318 10898 25333 10910
rect 25257 10846 25269 10898
rect 25321 10846 25333 10898
rect 25257 10794 25272 10846
rect 25318 10794 25333 10846
rect 25257 10742 25269 10794
rect 25321 10742 25333 10794
rect 25257 10730 25272 10742
rect 25318 10730 25333 10742
rect 25417 10898 25432 10910
rect 25560 11304 25606 11666
rect 25478 10898 25493 10910
rect 25417 10846 25429 10898
rect 25481 10846 25493 10898
rect 25417 10794 25432 10846
rect 25478 10794 25493 10846
rect 25417 10742 25429 10794
rect 25481 10742 25493 10794
rect 25417 10730 25432 10742
rect 25478 10730 25493 10742
rect 24024 10368 24070 10730
rect 24152 10368 24198 10730
rect 24137 9962 24152 9974
rect 24312 10368 24358 10730
rect 24472 10368 24518 10730
rect 24632 10368 24678 10730
rect 24198 9962 24213 9974
rect 24137 9910 24149 9962
rect 24201 9910 24213 9962
rect 24137 9858 24152 9910
rect 24198 9858 24213 9910
rect 24137 9806 24149 9858
rect 24201 9806 24213 9858
rect 24137 9794 24152 9806
rect 24198 9794 24213 9806
rect 24457 10356 24472 10368
rect 24518 10356 24533 10368
rect 24457 10304 24469 10356
rect 24521 10304 24533 10356
rect 24457 10252 24472 10304
rect 24518 10252 24533 10304
rect 24457 10200 24469 10252
rect 24521 10200 24533 10252
rect 24457 10188 24472 10200
rect 24024 9432 24070 9794
rect 24152 9783 24198 9794
rect 24312 9783 24358 9794
rect 24518 10188 24533 10200
rect 24472 9783 24518 9794
rect 24792 10368 24838 10730
rect 24777 9962 24792 9974
rect 24952 10368 24998 10730
rect 25112 10368 25158 10730
rect 25272 10368 25318 10730
rect 24838 9962 24853 9974
rect 24777 9910 24789 9962
rect 24841 9910 24853 9962
rect 24777 9858 24792 9910
rect 24838 9858 24853 9910
rect 24777 9806 24789 9858
rect 24841 9806 24853 9858
rect 24777 9794 24792 9806
rect 24838 9794 24853 9806
rect 25097 10356 25112 10368
rect 25158 10356 25173 10368
rect 25097 10304 25109 10356
rect 25161 10304 25173 10356
rect 25097 10252 25112 10304
rect 25158 10252 25173 10304
rect 25097 10200 25109 10252
rect 25161 10200 25173 10252
rect 25097 10188 25112 10200
rect 24632 9783 24678 9794
rect 24792 9783 24838 9794
rect 24952 9735 24998 9794
rect 25158 10188 25173 10200
rect 25112 9783 25158 9794
rect 25432 10368 25478 10730
rect 25417 9962 25432 9974
rect 25560 10368 25606 10730
rect 25478 9962 25493 9974
rect 25417 9910 25429 9962
rect 25481 9910 25493 9962
rect 25417 9858 25432 9910
rect 25478 9858 25493 9910
rect 25417 9806 25429 9858
rect 25481 9806 25493 9858
rect 25417 9794 25432 9806
rect 25478 9794 25493 9806
rect 25272 9735 25318 9794
rect 25432 9783 25478 9794
rect 24952 9689 25318 9735
rect 25337 9631 25413 9643
rect 25337 9628 25349 9631
rect 24221 9582 24232 9628
rect 24278 9582 24552 9628
rect 24598 9582 24872 9628
rect 24918 9582 25192 9628
rect 25238 9582 25349 9628
rect 25337 9579 25349 9582
rect 25401 9579 25413 9631
rect 25337 9567 25413 9579
rect 24152 9432 24198 9443
rect 24137 9026 24152 9038
rect 24312 9432 24358 9443
rect 24472 9432 24518 9443
rect 24632 9432 24678 9443
rect 24198 9026 24213 9038
rect 24137 8974 24149 9026
rect 24201 8974 24213 9026
rect 24137 8922 24152 8974
rect 24198 8922 24213 8974
rect 24137 8870 24149 8922
rect 24201 8870 24213 8922
rect 24137 8858 24152 8870
rect 24198 8858 24213 8870
rect 24297 9026 24312 9038
rect 24457 9420 24472 9432
rect 24518 9420 24533 9432
rect 24457 9368 24469 9420
rect 24521 9368 24533 9420
rect 24457 9316 24472 9368
rect 24518 9316 24533 9368
rect 24457 9264 24469 9316
rect 24521 9264 24533 9316
rect 24457 9252 24472 9264
rect 24358 9026 24373 9038
rect 24297 8974 24309 9026
rect 24361 8974 24373 9026
rect 24297 8922 24312 8974
rect 24358 8922 24373 8974
rect 24297 8870 24309 8922
rect 24361 8870 24373 8922
rect 24297 8858 24312 8870
rect 24358 8858 24373 8870
rect 24518 9252 24533 9264
rect 24617 9026 24632 9038
rect 24792 9432 24838 9443
rect 24678 9026 24693 9038
rect 24617 8974 24629 9026
rect 24681 8974 24693 9026
rect 24617 8922 24632 8974
rect 24678 8922 24693 8974
rect 24617 8870 24629 8922
rect 24681 8870 24693 8922
rect 24617 8858 24632 8870
rect 24678 8858 24693 8870
rect 24777 9026 24792 9038
rect 24952 9432 24998 9443
rect 25112 9432 25158 9443
rect 25272 9432 25318 9443
rect 24838 9026 24853 9038
rect 24777 8974 24789 9026
rect 24841 8974 24853 9026
rect 24777 8922 24792 8974
rect 24838 8922 24853 8974
rect 24777 8870 24789 8922
rect 24841 8870 24853 8922
rect 24777 8858 24792 8870
rect 24838 8858 24853 8870
rect 24937 9026 24952 9038
rect 25097 9420 25112 9432
rect 25158 9420 25173 9432
rect 25097 9368 25109 9420
rect 25161 9368 25173 9420
rect 25097 9316 25112 9368
rect 25158 9316 25173 9368
rect 25097 9264 25109 9316
rect 25161 9264 25173 9316
rect 25097 9252 25112 9264
rect 24998 9026 25013 9038
rect 24937 8974 24949 9026
rect 25001 8974 25013 9026
rect 24937 8922 24952 8974
rect 24998 8922 25013 8974
rect 24937 8870 24949 8922
rect 25001 8870 25013 8922
rect 24937 8858 24952 8870
rect 24998 8858 25013 8870
rect 25158 9252 25173 9264
rect 25257 9026 25272 9038
rect 25432 9432 25478 9443
rect 25318 9026 25333 9038
rect 25257 8974 25269 9026
rect 25321 8974 25333 9026
rect 25257 8922 25272 8974
rect 25318 8922 25333 8974
rect 25257 8870 25269 8922
rect 25321 8870 25333 8922
rect 25257 8858 25272 8870
rect 25318 8858 25333 8870
rect 25417 9026 25432 9038
rect 25560 9432 25606 9794
rect 25478 9026 25493 9038
rect 25417 8974 25429 9026
rect 25481 8974 25493 9026
rect 25417 8922 25432 8974
rect 25478 8922 25493 8974
rect 25417 8870 25429 8922
rect 25481 8870 25493 8922
rect 25417 8858 25432 8870
rect 25478 8858 25493 8870
rect 24024 8700 24070 8858
rect 24152 8847 24198 8858
rect 24312 8847 24358 8858
rect 24472 8847 24518 8858
rect 24632 8847 24678 8858
rect 24792 8847 24838 8858
rect 24952 8799 24998 8858
rect 25112 8847 25158 8858
rect 25272 8799 25318 8858
rect 25432 8847 25478 8858
rect 24952 8753 25318 8799
rect 23864 8654 23944 8700
rect 23990 8654 24070 8700
rect 25337 8695 25413 8707
rect 25337 8692 25349 8695
rect 23864 8496 23910 8654
rect 23864 7541 23910 7922
rect 24024 8496 24070 8654
rect 24221 8646 24232 8692
rect 24278 8646 24552 8692
rect 24598 8646 24872 8692
rect 24918 8646 25192 8692
rect 25238 8646 25349 8692
rect 25337 8643 25349 8646
rect 25401 8643 25413 8695
rect 25337 8631 25413 8643
rect 25560 8700 25606 8858
rect 25720 12240 25766 12398
rect 25720 11304 25766 11666
rect 25720 10368 25766 10730
rect 25720 9432 25766 9794
rect 25720 8700 25766 8858
rect 25560 8654 25640 8700
rect 25686 8654 25766 8700
rect 24152 8496 24198 8507
rect 24137 8090 24152 8102
rect 24312 8496 24358 8507
rect 24472 8496 24518 8507
rect 24632 8496 24678 8507
rect 24198 8090 24213 8102
rect 24137 8038 24149 8090
rect 24201 8038 24213 8090
rect 24137 7986 24152 8038
rect 24198 7986 24213 8038
rect 24137 7934 24149 7986
rect 24201 7934 24213 7986
rect 24137 7922 24152 7934
rect 24198 7922 24213 7934
rect 24297 8090 24312 8102
rect 24457 8484 24472 8496
rect 24518 8484 24533 8496
rect 24457 8432 24469 8484
rect 24521 8432 24533 8484
rect 24457 8380 24472 8432
rect 24518 8380 24533 8432
rect 24457 8328 24469 8380
rect 24521 8328 24533 8380
rect 24457 8316 24472 8328
rect 24358 8090 24373 8102
rect 24297 8038 24309 8090
rect 24361 8038 24373 8090
rect 24297 7986 24312 8038
rect 24358 7986 24373 8038
rect 24297 7934 24309 7986
rect 24361 7934 24373 7986
rect 24297 7922 24312 7934
rect 24358 7922 24373 7934
rect 24518 8316 24533 8328
rect 24617 8090 24632 8102
rect 24792 8496 24838 8507
rect 24678 8090 24693 8102
rect 24617 8038 24629 8090
rect 24681 8038 24693 8090
rect 24617 7986 24632 8038
rect 24678 7986 24693 8038
rect 24617 7934 24629 7986
rect 24681 7934 24693 7986
rect 24617 7922 24632 7934
rect 24678 7922 24693 7934
rect 24777 8090 24792 8102
rect 24952 8496 24998 8507
rect 25112 8496 25158 8507
rect 25272 8496 25318 8507
rect 24838 8090 24853 8102
rect 24777 8038 24789 8090
rect 24841 8038 24853 8090
rect 24777 7986 24792 8038
rect 24838 7986 24853 8038
rect 24777 7934 24789 7986
rect 24841 7934 24853 7986
rect 24777 7922 24792 7934
rect 24838 7922 24853 7934
rect 24937 8090 24952 8102
rect 25097 8484 25112 8496
rect 25158 8484 25173 8496
rect 25097 8432 25109 8484
rect 25161 8432 25173 8484
rect 25097 8380 25112 8432
rect 25158 8380 25173 8432
rect 25097 8328 25109 8380
rect 25161 8328 25173 8380
rect 25097 8316 25112 8328
rect 24998 8090 25013 8102
rect 24937 8038 24949 8090
rect 25001 8038 25013 8090
rect 24937 7986 24952 8038
rect 24998 7986 25013 8038
rect 24937 7934 24949 7986
rect 25001 7934 25013 7986
rect 24937 7922 24952 7934
rect 24998 7922 25013 7934
rect 25158 8316 25173 8328
rect 25257 8090 25272 8102
rect 25432 8496 25478 8507
rect 25318 8090 25333 8102
rect 25257 8038 25269 8090
rect 25321 8038 25333 8090
rect 25257 7986 25272 8038
rect 25318 7986 25333 8038
rect 25257 7934 25269 7986
rect 25321 7934 25333 7986
rect 25257 7922 25272 7934
rect 25318 7922 25333 7934
rect 25417 8090 25432 8102
rect 25560 8496 25606 8654
rect 25478 8090 25493 8102
rect 25417 8038 25429 8090
rect 25481 8038 25493 8090
rect 25417 7986 25432 8038
rect 25478 7986 25493 8038
rect 25417 7934 25429 7986
rect 25481 7934 25493 7986
rect 25417 7922 25432 7934
rect 25478 7922 25493 7934
rect 24024 7541 24070 7922
rect 24152 7911 24198 7922
rect 24312 7863 24358 7922
rect 24472 7911 24518 7922
rect 24632 7863 24678 7922
rect 24792 7911 24838 7922
rect 24952 7863 24998 7922
rect 25112 7911 25158 7922
rect 25272 7863 25318 7922
rect 25432 7911 25478 7922
rect 24312 7817 25318 7863
rect 24312 7541 24358 7817
rect 24537 7759 24613 7771
rect 24537 7707 24549 7759
rect 24601 7756 24613 7759
rect 25177 7759 25253 7771
rect 25177 7756 25189 7759
rect 24601 7710 25189 7756
rect 24601 7707 24613 7710
rect 24537 7695 24613 7707
rect 25177 7707 25189 7710
rect 25241 7707 25253 7759
rect 25177 7695 25253 7707
rect 25560 7541 25606 7922
rect 25720 8496 25766 8654
rect 25720 7541 25766 7922
rect 26103 13534 26296 13557
rect 26342 13557 27257 13580
rect 26342 13534 26423 13557
rect 26103 13486 26423 13534
rect 26103 13440 26296 13486
rect 26342 13440 26423 13486
rect 26103 13392 26423 13440
rect 26103 13346 26296 13392
rect 26342 13346 26423 13392
rect 26103 13298 26423 13346
rect 26103 13252 26296 13298
rect 26342 13252 26423 13298
rect 26103 13204 26423 13252
rect 26103 13158 26296 13204
rect 26342 13158 26423 13204
rect 26103 13110 26423 13158
rect 26103 13064 26296 13110
rect 26342 13064 26423 13110
rect 26103 13016 26423 13064
rect 26103 12970 26296 13016
rect 26342 12970 26423 13016
rect 26103 12922 26423 12970
rect 26103 12876 26296 12922
rect 26342 12876 26423 12922
rect 26103 12828 26423 12876
rect 26103 12782 26296 12828
rect 26342 12782 26423 12828
rect 26103 12734 26423 12782
rect 26103 12688 26296 12734
rect 26342 12688 26423 12734
rect 26103 12640 26423 12688
rect 26103 12594 26296 12640
rect 26342 12594 26423 12640
rect 26103 12546 26423 12594
rect 26103 12500 26296 12546
rect 26342 12500 26423 12546
rect 26103 12452 26423 12500
rect 26103 12406 26296 12452
rect 26342 12406 26423 12452
rect 26103 12358 26423 12406
rect 26103 12312 26296 12358
rect 26342 12312 26423 12358
rect 26103 12264 26423 12312
rect 26103 12218 26296 12264
rect 26342 12218 26423 12264
rect 26103 12170 26423 12218
rect 26103 12124 26296 12170
rect 26342 12124 26423 12170
rect 26103 12076 26423 12124
rect 26103 12030 26296 12076
rect 26342 12030 26423 12076
rect 26103 11982 26423 12030
rect 26103 11936 26296 11982
rect 26342 11936 26423 11982
rect 26103 11888 26423 11936
rect 26103 11842 26296 11888
rect 26342 11842 26423 11888
rect 26103 11794 26423 11842
rect 26103 11748 26296 11794
rect 26342 11748 26423 11794
rect 26103 11700 26423 11748
rect 26103 11654 26296 11700
rect 26342 11654 26423 11700
rect 26103 11606 26423 11654
rect 26103 11560 26296 11606
rect 26342 11560 26423 11606
rect 26103 11512 26423 11560
rect 26103 11466 26296 11512
rect 26342 11466 26423 11512
rect 26103 11418 26423 11466
rect 26103 11372 26296 11418
rect 26342 11372 26423 11418
rect 26103 11324 26423 11372
rect 26103 11278 26296 11324
rect 26342 11278 26423 11324
rect 26103 11230 26423 11278
rect 26103 11184 26296 11230
rect 26342 11184 26423 11230
rect 26103 11136 26423 11184
rect 26103 11090 26296 11136
rect 26342 11090 26423 11136
rect 26103 11042 26423 11090
rect 26103 10996 26296 11042
rect 26342 10996 26423 11042
rect 26103 10948 26423 10996
rect 26103 10902 26296 10948
rect 26342 10902 26423 10948
rect 26103 10854 26423 10902
rect 26103 10808 26296 10854
rect 26342 10808 26423 10854
rect 26103 10760 26423 10808
rect 26103 10714 26296 10760
rect 26342 10714 26423 10760
rect 26103 10666 26423 10714
rect 26103 10620 26296 10666
rect 26342 10620 26423 10666
rect 26103 10572 26423 10620
rect 26103 10526 26296 10572
rect 26342 10526 26423 10572
rect 26103 10478 26423 10526
rect 26103 10432 26296 10478
rect 26342 10432 26423 10478
rect 26103 10384 26423 10432
rect 26103 10338 26296 10384
rect 26342 10338 26423 10384
rect 26103 10290 26423 10338
rect 26103 10244 26296 10290
rect 26342 10244 26423 10290
rect 26103 10196 26423 10244
rect 26103 10150 26296 10196
rect 26342 10150 26423 10196
rect 26103 10102 26423 10150
rect 26103 10056 26296 10102
rect 26342 10056 26423 10102
rect 26103 10008 26423 10056
rect 26103 9962 26296 10008
rect 26342 9962 26423 10008
rect 26103 9914 26423 9962
rect 26103 9868 26296 9914
rect 26342 9868 26423 9914
rect 26103 9820 26423 9868
rect 26103 9774 26296 9820
rect 26342 9774 26423 9820
rect 26103 9726 26423 9774
rect 26103 9680 26296 9726
rect 26342 9680 26423 9726
rect 26103 9632 26423 9680
rect 26103 9586 26296 9632
rect 26342 9586 26423 9632
rect 26103 9538 26423 9586
rect 26103 9492 26296 9538
rect 26342 9492 26423 9538
rect 26103 9444 26423 9492
rect 26103 9398 26296 9444
rect 26342 9398 26423 9444
rect 26103 9350 26423 9398
rect 26103 9304 26296 9350
rect 26342 9304 26423 9350
rect 26103 9256 26423 9304
rect 26103 9210 26296 9256
rect 26342 9210 26423 9256
rect 26103 9162 26423 9210
rect 26103 9116 26296 9162
rect 26342 9116 26423 9162
rect 26103 9068 26423 9116
rect 26103 9022 26296 9068
rect 26342 9022 26423 9068
rect 26103 8974 26423 9022
rect 26103 8928 26296 8974
rect 26342 8928 26423 8974
rect 26103 8880 26423 8928
rect 26103 8834 26296 8880
rect 26342 8834 26423 8880
rect 26103 8786 26423 8834
rect 26103 8740 26296 8786
rect 26342 8740 26423 8786
rect 26103 8692 26423 8740
rect 26103 8646 26296 8692
rect 26342 8646 26423 8692
rect 26103 8598 26423 8646
rect 26103 8552 26296 8598
rect 26342 8552 26423 8598
rect 26103 8504 26423 8552
rect 26103 8458 26296 8504
rect 26342 8458 26423 8504
rect 26103 8410 26423 8458
rect 26103 8364 26296 8410
rect 26342 8364 26423 8410
rect 26103 8316 26423 8364
rect 26103 8270 26296 8316
rect 26342 8270 26423 8316
rect 26103 8222 26423 8270
rect 26103 8176 26296 8222
rect 26342 8176 26423 8222
rect 26103 8128 26423 8176
rect 26103 8082 26296 8128
rect 26342 8082 26423 8128
rect 26103 8034 26423 8082
rect 26103 7988 26296 8034
rect 26342 7988 26423 8034
rect 26103 7940 26423 7988
rect 26103 7894 26296 7940
rect 26342 7894 26423 7940
rect 26103 7846 26423 7894
rect 26103 7800 26296 7846
rect 26342 7800 26423 7846
rect 26103 7752 26423 7800
rect 26103 7706 26296 7752
rect 26342 7706 26423 7752
rect 26103 7658 26423 7706
rect 26103 7612 26296 7658
rect 26342 7612 26423 7658
rect 26103 7564 26423 7612
rect 26103 7541 26296 7564
rect 23334 7518 26296 7541
rect 26342 7541 26423 7564
rect 27176 13534 27257 13557
rect 27303 13557 30265 13580
rect 27303 13534 27496 13557
rect 27176 13486 27496 13534
rect 27176 13440 27257 13486
rect 27303 13440 27496 13486
rect 27176 13392 27496 13440
rect 27176 13346 27257 13392
rect 27303 13346 27496 13392
rect 27176 13298 27496 13346
rect 27176 13252 27257 13298
rect 27303 13252 27496 13298
rect 27176 13204 27496 13252
rect 27176 13158 27257 13204
rect 27303 13158 27496 13204
rect 27176 13110 27496 13158
rect 27176 13064 27257 13110
rect 27303 13064 27496 13110
rect 27176 13016 27496 13064
rect 27176 12970 27257 13016
rect 27303 12970 27496 13016
rect 27176 12922 27496 12970
rect 27176 12876 27257 12922
rect 27303 12876 27496 12922
rect 27176 12828 27496 12876
rect 27176 12782 27257 12828
rect 27303 12782 27496 12828
rect 27176 12734 27496 12782
rect 27176 12688 27257 12734
rect 27303 12688 27496 12734
rect 27176 12640 27496 12688
rect 27176 12594 27257 12640
rect 27303 12594 27496 12640
rect 27176 12546 27496 12594
rect 27176 12500 27257 12546
rect 27303 12500 27496 12546
rect 27176 12452 27496 12500
rect 27176 12406 27257 12452
rect 27303 12406 27496 12452
rect 27176 12358 27496 12406
rect 27176 12312 27257 12358
rect 27303 12312 27496 12358
rect 27176 12264 27496 12312
rect 27176 12218 27257 12264
rect 27303 12218 27496 12264
rect 27176 12170 27496 12218
rect 27176 12124 27257 12170
rect 27303 12124 27496 12170
rect 27176 12076 27496 12124
rect 27176 12030 27257 12076
rect 27303 12030 27496 12076
rect 27176 11982 27496 12030
rect 27176 11936 27257 11982
rect 27303 11936 27496 11982
rect 27176 11888 27496 11936
rect 27176 11842 27257 11888
rect 27303 11842 27496 11888
rect 27176 11794 27496 11842
rect 27176 11748 27257 11794
rect 27303 11748 27496 11794
rect 27176 11700 27496 11748
rect 27176 11654 27257 11700
rect 27303 11654 27496 11700
rect 27176 11606 27496 11654
rect 27176 11560 27257 11606
rect 27303 11560 27496 11606
rect 27176 11512 27496 11560
rect 27176 11466 27257 11512
rect 27303 11466 27496 11512
rect 27176 11418 27496 11466
rect 27176 11372 27257 11418
rect 27303 11372 27496 11418
rect 27176 11324 27496 11372
rect 27176 11278 27257 11324
rect 27303 11278 27496 11324
rect 27176 11230 27496 11278
rect 27176 11184 27257 11230
rect 27303 11184 27496 11230
rect 27176 11136 27496 11184
rect 27176 11090 27257 11136
rect 27303 11090 27496 11136
rect 27176 11042 27496 11090
rect 27176 10996 27257 11042
rect 27303 10996 27496 11042
rect 27176 10948 27496 10996
rect 27176 10902 27257 10948
rect 27303 10902 27496 10948
rect 27176 10854 27496 10902
rect 27176 10808 27257 10854
rect 27303 10808 27496 10854
rect 27176 10760 27496 10808
rect 27176 10714 27257 10760
rect 27303 10714 27496 10760
rect 27176 10666 27496 10714
rect 27176 10620 27257 10666
rect 27303 10620 27496 10666
rect 27176 10572 27496 10620
rect 27176 10526 27257 10572
rect 27303 10526 27496 10572
rect 27176 10478 27496 10526
rect 27176 10432 27257 10478
rect 27303 10432 27496 10478
rect 27176 10384 27496 10432
rect 27176 10338 27257 10384
rect 27303 10338 27496 10384
rect 27176 10290 27496 10338
rect 27176 10244 27257 10290
rect 27303 10244 27496 10290
rect 27176 10196 27496 10244
rect 27176 10150 27257 10196
rect 27303 10150 27496 10196
rect 27176 10102 27496 10150
rect 27176 10056 27257 10102
rect 27303 10056 27496 10102
rect 27176 10008 27496 10056
rect 27176 9962 27257 10008
rect 27303 9962 27496 10008
rect 27176 9914 27496 9962
rect 27176 9868 27257 9914
rect 27303 9868 27496 9914
rect 27176 9820 27496 9868
rect 27176 9774 27257 9820
rect 27303 9774 27496 9820
rect 27176 9726 27496 9774
rect 27176 9680 27257 9726
rect 27303 9680 27496 9726
rect 27176 9632 27496 9680
rect 27176 9586 27257 9632
rect 27303 9586 27496 9632
rect 27176 9538 27496 9586
rect 27176 9492 27257 9538
rect 27303 9492 27496 9538
rect 27176 9444 27496 9492
rect 27176 9398 27257 9444
rect 27303 9398 27496 9444
rect 27176 9350 27496 9398
rect 27176 9304 27257 9350
rect 27303 9304 27496 9350
rect 27176 9256 27496 9304
rect 27176 9210 27257 9256
rect 27303 9210 27496 9256
rect 27176 9162 27496 9210
rect 27176 9116 27257 9162
rect 27303 9116 27496 9162
rect 27176 9068 27496 9116
rect 27176 9022 27257 9068
rect 27303 9022 27496 9068
rect 27176 8974 27496 9022
rect 27176 8928 27257 8974
rect 27303 8928 27496 8974
rect 27176 8880 27496 8928
rect 27176 8834 27257 8880
rect 27303 8834 27496 8880
rect 27176 8786 27496 8834
rect 27176 8740 27257 8786
rect 27303 8740 27496 8786
rect 27176 8692 27496 8740
rect 27176 8646 27257 8692
rect 27303 8646 27496 8692
rect 27176 8598 27496 8646
rect 27176 8552 27257 8598
rect 27303 8552 27496 8598
rect 27176 8504 27496 8552
rect 27176 8458 27257 8504
rect 27303 8458 27496 8504
rect 27176 8410 27496 8458
rect 27176 8364 27257 8410
rect 27303 8364 27496 8410
rect 27176 8316 27496 8364
rect 27176 8270 27257 8316
rect 27303 8270 27496 8316
rect 27176 8222 27496 8270
rect 27176 8176 27257 8222
rect 27303 8176 27496 8222
rect 27176 8128 27496 8176
rect 27176 8082 27257 8128
rect 27303 8082 27496 8128
rect 27176 8034 27496 8082
rect 27176 7988 27257 8034
rect 27303 7988 27496 8034
rect 27176 7940 27496 7988
rect 27176 7894 27257 7940
rect 27303 7894 27496 7940
rect 27176 7846 27496 7894
rect 27176 7800 27257 7846
rect 27303 7800 27496 7846
rect 27176 7752 27496 7800
rect 27176 7706 27257 7752
rect 27303 7706 27496 7752
rect 27176 7658 27496 7706
rect 27176 7612 27257 7658
rect 27303 7612 27496 7658
rect 27176 7564 27496 7612
rect 27176 7541 27257 7564
rect 26342 7518 27257 7541
rect 27303 7541 27496 7564
rect 27833 13176 27879 13557
rect 27833 12444 27879 12602
rect 27993 13176 28039 13557
rect 28186 13405 28262 13417
rect 28186 13353 28198 13405
rect 28250 13402 28262 13405
rect 28250 13356 28681 13402
rect 28727 13356 29321 13402
rect 29367 13356 29378 13402
rect 28250 13353 28262 13356
rect 28186 13341 28262 13353
rect 28121 13176 28167 13187
rect 28106 12770 28121 12782
rect 28281 13176 28327 13187
rect 28441 13176 28487 13187
rect 28601 13176 28647 13187
rect 28167 12770 28182 12782
rect 28106 12718 28118 12770
rect 28170 12718 28182 12770
rect 28106 12666 28121 12718
rect 28167 12666 28182 12718
rect 28106 12614 28118 12666
rect 28170 12614 28182 12666
rect 28106 12602 28121 12614
rect 28167 12602 28182 12614
rect 28266 12770 28281 12782
rect 28426 13164 28441 13176
rect 28487 13164 28502 13176
rect 28426 13112 28438 13164
rect 28490 13112 28502 13164
rect 28426 13060 28441 13112
rect 28487 13060 28502 13112
rect 28426 13008 28438 13060
rect 28490 13008 28502 13060
rect 28426 12996 28441 13008
rect 28327 12770 28342 12782
rect 28266 12718 28278 12770
rect 28330 12718 28342 12770
rect 28266 12666 28281 12718
rect 28327 12666 28342 12718
rect 28266 12614 28278 12666
rect 28330 12614 28342 12666
rect 28266 12602 28281 12614
rect 28327 12602 28342 12614
rect 28487 12996 28502 13008
rect 28586 12770 28601 12782
rect 28761 13176 28807 13187
rect 28647 12770 28662 12782
rect 28586 12718 28598 12770
rect 28650 12718 28662 12770
rect 28586 12666 28601 12718
rect 28647 12666 28662 12718
rect 28586 12614 28598 12666
rect 28650 12614 28662 12666
rect 28586 12602 28601 12614
rect 28647 12602 28662 12614
rect 28746 12770 28761 12782
rect 28921 13176 28967 13187
rect 29081 13176 29127 13187
rect 29241 13176 29287 13187
rect 28807 12770 28822 12782
rect 28746 12718 28758 12770
rect 28810 12718 28822 12770
rect 28746 12666 28761 12718
rect 28807 12666 28822 12718
rect 28746 12614 28758 12666
rect 28810 12614 28822 12666
rect 28746 12602 28761 12614
rect 28807 12602 28822 12614
rect 28906 12770 28921 12782
rect 29066 13164 29081 13176
rect 29127 13164 29142 13176
rect 29066 13112 29078 13164
rect 29130 13112 29142 13164
rect 29066 13060 29081 13112
rect 29127 13060 29142 13112
rect 29066 13008 29078 13060
rect 29130 13008 29142 13060
rect 29066 12996 29081 13008
rect 28967 12770 28982 12782
rect 28906 12718 28918 12770
rect 28970 12718 28982 12770
rect 28906 12666 28921 12718
rect 28967 12666 28982 12718
rect 28906 12614 28918 12666
rect 28970 12614 28982 12666
rect 28906 12602 28921 12614
rect 28967 12602 28982 12614
rect 29127 12996 29142 13008
rect 29226 12770 29241 12782
rect 29401 13176 29447 13187
rect 29287 12770 29302 12782
rect 29226 12718 29238 12770
rect 29290 12718 29302 12770
rect 29226 12666 29241 12718
rect 29287 12666 29302 12718
rect 29226 12614 29238 12666
rect 29290 12614 29302 12666
rect 29226 12602 29241 12614
rect 29287 12602 29302 12614
rect 29386 12770 29401 12782
rect 29529 13176 29575 13557
rect 29447 12770 29462 12782
rect 29386 12718 29398 12770
rect 29450 12718 29462 12770
rect 29386 12666 29401 12718
rect 29447 12666 29462 12718
rect 29386 12614 29398 12666
rect 29450 12614 29462 12666
rect 29386 12602 29401 12614
rect 29447 12602 29462 12614
rect 27993 12444 28039 12602
rect 28121 12591 28167 12602
rect 28281 12543 28327 12602
rect 28441 12591 28487 12602
rect 28601 12543 28647 12602
rect 28761 12591 28807 12602
rect 28921 12591 28967 12602
rect 29081 12591 29127 12602
rect 29241 12591 29287 12602
rect 29401 12591 29447 12602
rect 28281 12497 28647 12543
rect 27833 12398 27913 12444
rect 27959 12398 28039 12444
rect 27833 12240 27879 12398
rect 27833 11304 27879 11666
rect 27833 10368 27879 10730
rect 27833 9432 27879 9794
rect 27833 8700 27879 8858
rect 27993 12240 28039 12398
rect 28186 12439 28262 12451
rect 28186 12387 28198 12439
rect 28250 12436 28262 12439
rect 29529 12444 29575 12602
rect 29689 13176 29735 13557
rect 29689 12444 29735 12602
rect 28250 12390 28361 12436
rect 28407 12390 28681 12436
rect 28727 12390 29001 12436
rect 29047 12390 29321 12436
rect 29367 12390 29378 12436
rect 29529 12398 29609 12444
rect 29655 12398 29735 12444
rect 28250 12387 28262 12390
rect 28186 12375 28262 12387
rect 28121 12240 28167 12251
rect 28106 11834 28121 11846
rect 28281 12240 28327 12251
rect 28441 12240 28487 12251
rect 28601 12240 28647 12251
rect 28167 11834 28182 11846
rect 28106 11782 28118 11834
rect 28170 11782 28182 11834
rect 28106 11730 28121 11782
rect 28167 11730 28182 11782
rect 28106 11678 28118 11730
rect 28170 11678 28182 11730
rect 28106 11666 28121 11678
rect 28167 11666 28182 11678
rect 28266 11834 28281 11846
rect 28426 12228 28441 12240
rect 28487 12228 28502 12240
rect 28426 12176 28438 12228
rect 28490 12176 28502 12228
rect 28426 12124 28441 12176
rect 28487 12124 28502 12176
rect 28426 12072 28438 12124
rect 28490 12072 28502 12124
rect 28426 12060 28441 12072
rect 28327 11834 28342 11846
rect 28266 11782 28278 11834
rect 28330 11782 28342 11834
rect 28266 11730 28281 11782
rect 28327 11730 28342 11782
rect 28266 11678 28278 11730
rect 28330 11678 28342 11730
rect 28266 11666 28281 11678
rect 28327 11666 28342 11678
rect 28487 12060 28502 12072
rect 28586 11834 28601 11846
rect 28761 12240 28807 12251
rect 28647 11834 28662 11846
rect 28586 11782 28598 11834
rect 28650 11782 28662 11834
rect 28586 11730 28601 11782
rect 28647 11730 28662 11782
rect 28586 11678 28598 11730
rect 28650 11678 28662 11730
rect 28586 11666 28601 11678
rect 28647 11666 28662 11678
rect 28746 11834 28761 11846
rect 28921 12240 28967 12251
rect 29081 12240 29127 12251
rect 29241 12240 29287 12251
rect 28807 11834 28822 11846
rect 28746 11782 28758 11834
rect 28810 11782 28822 11834
rect 28746 11730 28761 11782
rect 28807 11730 28822 11782
rect 28746 11678 28758 11730
rect 28810 11678 28822 11730
rect 28746 11666 28761 11678
rect 28807 11666 28822 11678
rect 28906 11834 28921 11846
rect 29066 12228 29081 12240
rect 29127 12228 29142 12240
rect 29066 12176 29078 12228
rect 29130 12176 29142 12228
rect 29066 12124 29081 12176
rect 29127 12124 29142 12176
rect 29066 12072 29078 12124
rect 29130 12072 29142 12124
rect 29066 12060 29081 12072
rect 28967 11834 28982 11846
rect 28906 11782 28918 11834
rect 28970 11782 28982 11834
rect 28906 11730 28921 11782
rect 28967 11730 28982 11782
rect 28906 11678 28918 11730
rect 28970 11678 28982 11730
rect 28906 11666 28921 11678
rect 28967 11666 28982 11678
rect 29127 12060 29142 12072
rect 29226 11834 29241 11846
rect 29401 12240 29447 12251
rect 29287 11834 29302 11846
rect 29226 11782 29238 11834
rect 29290 11782 29302 11834
rect 29226 11730 29241 11782
rect 29287 11730 29302 11782
rect 29226 11678 29238 11730
rect 29290 11678 29302 11730
rect 29226 11666 29241 11678
rect 29287 11666 29302 11678
rect 29386 11834 29401 11846
rect 29529 12240 29575 12398
rect 29447 11834 29462 11846
rect 29386 11782 29398 11834
rect 29450 11782 29462 11834
rect 29386 11730 29401 11782
rect 29447 11730 29462 11782
rect 29386 11678 29398 11730
rect 29450 11678 29462 11730
rect 29386 11666 29401 11678
rect 29447 11666 29462 11678
rect 27993 11304 28039 11666
rect 28121 11655 28167 11666
rect 28281 11607 28327 11666
rect 28441 11655 28487 11666
rect 28601 11607 28647 11666
rect 28761 11655 28807 11666
rect 28921 11655 28967 11666
rect 29081 11655 29127 11666
rect 29241 11655 29287 11666
rect 29401 11655 29447 11666
rect 28281 11561 28647 11607
rect 28186 11503 28262 11515
rect 28186 11451 28198 11503
rect 28250 11500 28262 11503
rect 28250 11454 28361 11500
rect 28407 11454 28681 11500
rect 28727 11454 29001 11500
rect 29047 11454 29321 11500
rect 29367 11454 29378 11500
rect 28250 11451 28262 11454
rect 28186 11439 28262 11451
rect 28121 11304 28167 11315
rect 28106 10898 28121 10910
rect 28281 11304 28327 11315
rect 28441 11304 28487 11315
rect 28601 11304 28647 11315
rect 28167 10898 28182 10910
rect 28106 10846 28118 10898
rect 28170 10846 28182 10898
rect 28106 10794 28121 10846
rect 28167 10794 28182 10846
rect 28106 10742 28118 10794
rect 28170 10742 28182 10794
rect 28106 10730 28121 10742
rect 28167 10730 28182 10742
rect 28266 10898 28281 10910
rect 28426 11292 28441 11304
rect 28487 11292 28502 11304
rect 28426 11240 28438 11292
rect 28490 11240 28502 11292
rect 28426 11188 28441 11240
rect 28487 11188 28502 11240
rect 28426 11136 28438 11188
rect 28490 11136 28502 11188
rect 28426 11124 28441 11136
rect 28327 10898 28342 10910
rect 28266 10846 28278 10898
rect 28330 10846 28342 10898
rect 28266 10794 28281 10846
rect 28327 10794 28342 10846
rect 28266 10742 28278 10794
rect 28330 10742 28342 10794
rect 28266 10730 28281 10742
rect 28327 10730 28342 10742
rect 28487 11124 28502 11136
rect 28586 10898 28601 10910
rect 28761 11304 28807 11315
rect 28647 10898 28662 10910
rect 28586 10846 28598 10898
rect 28650 10846 28662 10898
rect 28586 10794 28601 10846
rect 28647 10794 28662 10846
rect 28586 10742 28598 10794
rect 28650 10742 28662 10794
rect 28586 10730 28601 10742
rect 28647 10730 28662 10742
rect 28746 10898 28761 10910
rect 28921 11304 28967 11315
rect 29081 11304 29127 11315
rect 29241 11304 29287 11315
rect 28807 10898 28822 10910
rect 28746 10846 28758 10898
rect 28810 10846 28822 10898
rect 28746 10794 28761 10846
rect 28807 10794 28822 10846
rect 28746 10742 28758 10794
rect 28810 10742 28822 10794
rect 28746 10730 28761 10742
rect 28807 10730 28822 10742
rect 28906 10898 28921 10910
rect 29066 11292 29081 11304
rect 29127 11292 29142 11304
rect 29066 11240 29078 11292
rect 29130 11240 29142 11292
rect 29066 11188 29081 11240
rect 29127 11188 29142 11240
rect 29066 11136 29078 11188
rect 29130 11136 29142 11188
rect 29066 11124 29081 11136
rect 28967 10898 28982 10910
rect 28906 10846 28918 10898
rect 28970 10846 28982 10898
rect 28906 10794 28921 10846
rect 28967 10794 28982 10846
rect 28906 10742 28918 10794
rect 28970 10742 28982 10794
rect 28906 10730 28921 10742
rect 28967 10730 28982 10742
rect 29127 11124 29142 11136
rect 29226 10898 29241 10910
rect 29401 11304 29447 11315
rect 29287 10898 29302 10910
rect 29226 10846 29238 10898
rect 29290 10846 29302 10898
rect 29226 10794 29241 10846
rect 29287 10794 29302 10846
rect 29226 10742 29238 10794
rect 29290 10742 29302 10794
rect 29226 10730 29241 10742
rect 29287 10730 29302 10742
rect 29386 10898 29401 10910
rect 29529 11304 29575 11666
rect 29447 10898 29462 10910
rect 29386 10846 29398 10898
rect 29450 10846 29462 10898
rect 29386 10794 29401 10846
rect 29447 10794 29462 10846
rect 29386 10742 29398 10794
rect 29450 10742 29462 10794
rect 29386 10730 29401 10742
rect 29447 10730 29462 10742
rect 27993 10368 28039 10730
rect 28121 10368 28167 10730
rect 28106 9962 28121 9974
rect 28281 10368 28327 10730
rect 28441 10368 28487 10730
rect 28601 10368 28647 10730
rect 28167 9962 28182 9974
rect 28106 9910 28118 9962
rect 28170 9910 28182 9962
rect 28106 9858 28121 9910
rect 28167 9858 28182 9910
rect 28106 9806 28118 9858
rect 28170 9806 28182 9858
rect 28106 9794 28121 9806
rect 28167 9794 28182 9806
rect 28426 10356 28441 10368
rect 28487 10356 28502 10368
rect 28426 10304 28438 10356
rect 28490 10304 28502 10356
rect 28426 10252 28441 10304
rect 28487 10252 28502 10304
rect 28426 10200 28438 10252
rect 28490 10200 28502 10252
rect 28426 10188 28441 10200
rect 27993 9432 28039 9794
rect 28121 9783 28167 9794
rect 28281 9735 28327 9794
rect 28487 10188 28502 10200
rect 28441 9783 28487 9794
rect 28761 10368 28807 10730
rect 28746 9962 28761 9974
rect 28921 10368 28967 10730
rect 29081 10368 29127 10730
rect 29241 10368 29287 10730
rect 28807 9962 28822 9974
rect 28746 9910 28758 9962
rect 28810 9910 28822 9962
rect 28746 9858 28761 9910
rect 28807 9858 28822 9910
rect 28746 9806 28758 9858
rect 28810 9806 28822 9858
rect 28746 9794 28761 9806
rect 28807 9794 28822 9806
rect 29066 10356 29081 10368
rect 29127 10356 29142 10368
rect 29066 10304 29078 10356
rect 29130 10304 29142 10356
rect 29066 10252 29081 10304
rect 29127 10252 29142 10304
rect 29066 10200 29078 10252
rect 29130 10200 29142 10252
rect 29066 10188 29081 10200
rect 28601 9735 28647 9794
rect 28761 9783 28807 9794
rect 28921 9783 28967 9794
rect 29127 10188 29142 10200
rect 29081 9783 29127 9794
rect 29401 10368 29447 10730
rect 29386 9962 29401 9974
rect 29529 10368 29575 10730
rect 29447 9962 29462 9974
rect 29386 9910 29398 9962
rect 29450 9910 29462 9962
rect 29386 9858 29401 9910
rect 29447 9858 29462 9910
rect 29386 9806 29398 9858
rect 29450 9806 29462 9858
rect 29386 9794 29401 9806
rect 29447 9794 29462 9806
rect 29241 9783 29287 9794
rect 29401 9783 29447 9794
rect 28281 9689 28647 9735
rect 28186 9631 28262 9643
rect 28186 9579 28198 9631
rect 28250 9628 28262 9631
rect 28250 9582 28361 9628
rect 28407 9582 28681 9628
rect 28727 9582 29001 9628
rect 29047 9582 29321 9628
rect 29367 9582 29378 9628
rect 28250 9579 28262 9582
rect 28186 9567 28262 9579
rect 28121 9432 28167 9443
rect 28106 9026 28121 9038
rect 28281 9432 28327 9443
rect 28441 9432 28487 9443
rect 28601 9432 28647 9443
rect 28167 9026 28182 9038
rect 28106 8974 28118 9026
rect 28170 8974 28182 9026
rect 28106 8922 28121 8974
rect 28167 8922 28182 8974
rect 28106 8870 28118 8922
rect 28170 8870 28182 8922
rect 28106 8858 28121 8870
rect 28167 8858 28182 8870
rect 28266 9026 28281 9038
rect 28426 9420 28441 9432
rect 28487 9420 28502 9432
rect 28426 9368 28438 9420
rect 28490 9368 28502 9420
rect 28426 9316 28441 9368
rect 28487 9316 28502 9368
rect 28426 9264 28438 9316
rect 28490 9264 28502 9316
rect 28426 9252 28441 9264
rect 28327 9026 28342 9038
rect 28266 8974 28278 9026
rect 28330 8974 28342 9026
rect 28266 8922 28281 8974
rect 28327 8922 28342 8974
rect 28266 8870 28278 8922
rect 28330 8870 28342 8922
rect 28266 8858 28281 8870
rect 28327 8858 28342 8870
rect 28487 9252 28502 9264
rect 28586 9026 28601 9038
rect 28761 9432 28807 9443
rect 28647 9026 28662 9038
rect 28586 8974 28598 9026
rect 28650 8974 28662 9026
rect 28586 8922 28601 8974
rect 28647 8922 28662 8974
rect 28586 8870 28598 8922
rect 28650 8870 28662 8922
rect 28586 8858 28601 8870
rect 28647 8858 28662 8870
rect 28746 9026 28761 9038
rect 28921 9432 28967 9443
rect 29081 9432 29127 9443
rect 29241 9432 29287 9443
rect 28807 9026 28822 9038
rect 28746 8974 28758 9026
rect 28810 8974 28822 9026
rect 28746 8922 28761 8974
rect 28807 8922 28822 8974
rect 28746 8870 28758 8922
rect 28810 8870 28822 8922
rect 28746 8858 28761 8870
rect 28807 8858 28822 8870
rect 28906 9026 28921 9038
rect 29066 9420 29081 9432
rect 29127 9420 29142 9432
rect 29066 9368 29078 9420
rect 29130 9368 29142 9420
rect 29066 9316 29081 9368
rect 29127 9316 29142 9368
rect 29066 9264 29078 9316
rect 29130 9264 29142 9316
rect 29066 9252 29081 9264
rect 28967 9026 28982 9038
rect 28906 8974 28918 9026
rect 28970 8974 28982 9026
rect 28906 8922 28921 8974
rect 28967 8922 28982 8974
rect 28906 8870 28918 8922
rect 28970 8870 28982 8922
rect 28906 8858 28921 8870
rect 28967 8858 28982 8870
rect 29127 9252 29142 9264
rect 29226 9026 29241 9038
rect 29401 9432 29447 9443
rect 29287 9026 29302 9038
rect 29226 8974 29238 9026
rect 29290 8974 29302 9026
rect 29226 8922 29241 8974
rect 29287 8922 29302 8974
rect 29226 8870 29238 8922
rect 29290 8870 29302 8922
rect 29226 8858 29241 8870
rect 29287 8858 29302 8870
rect 29386 9026 29401 9038
rect 29529 9432 29575 9794
rect 29447 9026 29462 9038
rect 29386 8974 29398 9026
rect 29450 8974 29462 9026
rect 29386 8922 29401 8974
rect 29447 8922 29462 8974
rect 29386 8870 29398 8922
rect 29450 8870 29462 8922
rect 29386 8858 29401 8870
rect 29447 8858 29462 8870
rect 27993 8700 28039 8858
rect 28121 8847 28167 8858
rect 28281 8799 28327 8858
rect 28441 8847 28487 8858
rect 28601 8799 28647 8858
rect 28761 8847 28807 8858
rect 28921 8847 28967 8858
rect 29081 8847 29127 8858
rect 29241 8847 29287 8858
rect 29401 8847 29447 8858
rect 28281 8753 28647 8799
rect 27833 8654 27913 8700
rect 27959 8654 28039 8700
rect 27833 8496 27879 8654
rect 27833 7541 27879 7922
rect 27993 8496 28039 8654
rect 28186 8695 28262 8707
rect 28186 8643 28198 8695
rect 28250 8692 28262 8695
rect 29529 8700 29575 8858
rect 29689 12240 29735 12398
rect 29689 11304 29735 11666
rect 29689 10368 29735 10730
rect 29689 9432 29735 9794
rect 29689 8700 29735 8858
rect 28250 8646 28361 8692
rect 28407 8646 28681 8692
rect 28727 8646 29001 8692
rect 29047 8646 29321 8692
rect 29367 8646 29378 8692
rect 29529 8654 29609 8700
rect 29655 8654 29735 8700
rect 28250 8643 28262 8646
rect 28186 8631 28262 8643
rect 28121 8496 28167 8507
rect 28106 8090 28121 8102
rect 28281 8496 28327 8507
rect 28441 8496 28487 8507
rect 28601 8496 28647 8507
rect 28167 8090 28182 8102
rect 28106 8038 28118 8090
rect 28170 8038 28182 8090
rect 28106 7986 28121 8038
rect 28167 7986 28182 8038
rect 28106 7934 28118 7986
rect 28170 7934 28182 7986
rect 28106 7922 28121 7934
rect 28167 7922 28182 7934
rect 28266 8090 28281 8102
rect 28426 8484 28441 8496
rect 28487 8484 28502 8496
rect 28426 8432 28438 8484
rect 28490 8432 28502 8484
rect 28426 8380 28441 8432
rect 28487 8380 28502 8432
rect 28426 8328 28438 8380
rect 28490 8328 28502 8380
rect 28426 8316 28441 8328
rect 28327 8090 28342 8102
rect 28266 8038 28278 8090
rect 28330 8038 28342 8090
rect 28266 7986 28281 8038
rect 28327 7986 28342 8038
rect 28266 7934 28278 7986
rect 28330 7934 28342 7986
rect 28266 7922 28281 7934
rect 28327 7922 28342 7934
rect 28487 8316 28502 8328
rect 28586 8090 28601 8102
rect 28761 8496 28807 8507
rect 28647 8090 28662 8102
rect 28586 8038 28598 8090
rect 28650 8038 28662 8090
rect 28586 7986 28601 8038
rect 28647 7986 28662 8038
rect 28586 7934 28598 7986
rect 28650 7934 28662 7986
rect 28586 7922 28601 7934
rect 28647 7922 28662 7934
rect 28746 8090 28761 8102
rect 28921 8496 28967 8507
rect 29081 8496 29127 8507
rect 29241 8496 29287 8507
rect 28807 8090 28822 8102
rect 28746 8038 28758 8090
rect 28810 8038 28822 8090
rect 28746 7986 28761 8038
rect 28807 7986 28822 8038
rect 28746 7934 28758 7986
rect 28810 7934 28822 7986
rect 28746 7922 28761 7934
rect 28807 7922 28822 7934
rect 28906 8090 28921 8102
rect 29066 8484 29081 8496
rect 29127 8484 29142 8496
rect 29066 8432 29078 8484
rect 29130 8432 29142 8484
rect 29066 8380 29081 8432
rect 29127 8380 29142 8432
rect 29066 8328 29078 8380
rect 29130 8328 29142 8380
rect 29066 8316 29081 8328
rect 28967 8090 28982 8102
rect 28906 8038 28918 8090
rect 28970 8038 28982 8090
rect 28906 7986 28921 8038
rect 28967 7986 28982 8038
rect 28906 7934 28918 7986
rect 28970 7934 28982 7986
rect 28906 7922 28921 7934
rect 28967 7922 28982 7934
rect 29127 8316 29142 8328
rect 29226 8090 29241 8102
rect 29401 8496 29447 8507
rect 29287 8090 29302 8102
rect 29226 8038 29238 8090
rect 29290 8038 29302 8090
rect 29226 7986 29241 8038
rect 29287 7986 29302 8038
rect 29226 7934 29238 7986
rect 29290 7934 29302 7986
rect 29226 7922 29241 7934
rect 29287 7922 29302 7934
rect 29386 8090 29401 8102
rect 29529 8496 29575 8654
rect 29447 8090 29462 8102
rect 29386 8038 29398 8090
rect 29450 8038 29462 8090
rect 29386 7986 29401 8038
rect 29447 7986 29462 8038
rect 29386 7934 29398 7986
rect 29450 7934 29462 7986
rect 29386 7922 29401 7934
rect 29447 7922 29462 7934
rect 27993 7541 28039 7922
rect 28121 7911 28167 7922
rect 28281 7863 28327 7922
rect 28441 7911 28487 7922
rect 28601 7863 28647 7922
rect 28761 7911 28807 7922
rect 28921 7863 28967 7922
rect 29081 7911 29127 7922
rect 29241 7863 29287 7922
rect 29401 7911 29447 7922
rect 28281 7817 29287 7863
rect 28346 7759 28422 7771
rect 28346 7707 28358 7759
rect 28410 7756 28422 7759
rect 28410 7710 29001 7756
rect 29047 7710 29058 7756
rect 28410 7707 28422 7710
rect 28346 7695 28422 7707
rect 29241 7541 29287 7817
rect 29529 7541 29575 7922
rect 29689 8496 29735 8654
rect 29689 7541 29735 7922
rect 30072 13534 30265 13557
rect 30311 13534 30392 13580
rect 30072 13486 30392 13534
rect 30072 13440 30265 13486
rect 30311 13440 30392 13486
rect 30072 13392 30392 13440
rect 30072 13346 30265 13392
rect 30311 13346 30392 13392
rect 30072 13298 30392 13346
rect 30072 13252 30265 13298
rect 30311 13252 30392 13298
rect 30072 13204 30392 13252
rect 30072 13158 30265 13204
rect 30311 13158 30392 13204
rect 30072 13110 30392 13158
rect 30072 13064 30265 13110
rect 30311 13064 30392 13110
rect 30072 13016 30392 13064
rect 30072 12970 30265 13016
rect 30311 12970 30392 13016
rect 30072 12922 30392 12970
rect 30072 12876 30265 12922
rect 30311 12876 30392 12922
rect 30072 12828 30392 12876
rect 30072 12782 30265 12828
rect 30311 12782 30392 12828
rect 30072 12734 30392 12782
rect 30072 12688 30265 12734
rect 30311 12688 30392 12734
rect 30072 12640 30392 12688
rect 30072 12594 30265 12640
rect 30311 12594 30392 12640
rect 30072 12546 30392 12594
rect 30072 12500 30265 12546
rect 30311 12500 30392 12546
rect 30072 12452 30392 12500
rect 30072 12406 30265 12452
rect 30311 12406 30392 12452
rect 30072 12358 30392 12406
rect 30072 12312 30265 12358
rect 30311 12312 30392 12358
rect 30072 12264 30392 12312
rect 30072 12218 30265 12264
rect 30311 12218 30392 12264
rect 30072 12170 30392 12218
rect 30072 12124 30265 12170
rect 30311 12124 30392 12170
rect 30072 12076 30392 12124
rect 30072 12030 30265 12076
rect 30311 12030 30392 12076
rect 30072 11982 30392 12030
rect 30072 11936 30265 11982
rect 30311 11936 30392 11982
rect 30072 11888 30392 11936
rect 30072 11842 30265 11888
rect 30311 11842 30392 11888
rect 30072 11794 30392 11842
rect 30072 11748 30265 11794
rect 30311 11748 30392 11794
rect 30072 11700 30392 11748
rect 30072 11654 30265 11700
rect 30311 11654 30392 11700
rect 30072 11606 30392 11654
rect 30072 11560 30265 11606
rect 30311 11560 30392 11606
rect 30072 11512 30392 11560
rect 30072 11466 30265 11512
rect 30311 11466 30392 11512
rect 30072 11418 30392 11466
rect 30072 11372 30265 11418
rect 30311 11372 30392 11418
rect 30072 11324 30392 11372
rect 30072 11278 30265 11324
rect 30311 11278 30392 11324
rect 30072 11230 30392 11278
rect 30072 11184 30265 11230
rect 30311 11184 30392 11230
rect 30072 11136 30392 11184
rect 30072 11090 30265 11136
rect 30311 11090 30392 11136
rect 30072 11042 30392 11090
rect 30072 10996 30265 11042
rect 30311 10996 30392 11042
rect 30072 10948 30392 10996
rect 30072 10902 30265 10948
rect 30311 10902 30392 10948
rect 30072 10854 30392 10902
rect 30072 10808 30265 10854
rect 30311 10808 30392 10854
rect 30072 10760 30392 10808
rect 30072 10714 30265 10760
rect 30311 10714 30392 10760
rect 30072 10666 30392 10714
rect 30072 10620 30265 10666
rect 30311 10620 30392 10666
rect 30072 10572 30392 10620
rect 30072 10526 30265 10572
rect 30311 10526 30392 10572
rect 30072 10478 30392 10526
rect 30072 10432 30265 10478
rect 30311 10432 30392 10478
rect 30072 10384 30392 10432
rect 30072 10338 30265 10384
rect 30311 10338 30392 10384
rect 30072 10290 30392 10338
rect 30072 10244 30265 10290
rect 30311 10244 30392 10290
rect 30072 10196 30392 10244
rect 30072 10150 30265 10196
rect 30311 10150 30392 10196
rect 30072 10102 30392 10150
rect 30072 10056 30265 10102
rect 30311 10056 30392 10102
rect 30072 10008 30392 10056
rect 30072 9962 30265 10008
rect 30311 9962 30392 10008
rect 30072 9914 30392 9962
rect 30072 9868 30265 9914
rect 30311 9868 30392 9914
rect 30072 9820 30392 9868
rect 30072 9774 30265 9820
rect 30311 9774 30392 9820
rect 30072 9726 30392 9774
rect 30072 9680 30265 9726
rect 30311 9680 30392 9726
rect 30072 9632 30392 9680
rect 30072 9586 30265 9632
rect 30311 9586 30392 9632
rect 30072 9538 30392 9586
rect 30072 9492 30265 9538
rect 30311 9492 30392 9538
rect 30072 9444 30392 9492
rect 30072 9398 30265 9444
rect 30311 9398 30392 9444
rect 30072 9350 30392 9398
rect 30072 9304 30265 9350
rect 30311 9304 30392 9350
rect 30072 9256 30392 9304
rect 30072 9210 30265 9256
rect 30311 9210 30392 9256
rect 30072 9162 30392 9210
rect 30072 9116 30265 9162
rect 30311 9116 30392 9162
rect 30072 9068 30392 9116
rect 30072 9022 30265 9068
rect 30311 9022 30392 9068
rect 30072 8974 30392 9022
rect 30072 8928 30265 8974
rect 30311 8928 30392 8974
rect 30072 8880 30392 8928
rect 30072 8834 30265 8880
rect 30311 8834 30392 8880
rect 30072 8786 30392 8834
rect 30072 8740 30265 8786
rect 30311 8740 30392 8786
rect 30072 8692 30392 8740
rect 30072 8646 30265 8692
rect 30311 8646 30392 8692
rect 30072 8598 30392 8646
rect 30072 8552 30265 8598
rect 30311 8552 30392 8598
rect 30072 8504 30392 8552
rect 30072 8458 30265 8504
rect 30311 8458 30392 8504
rect 30072 8410 30392 8458
rect 30072 8364 30265 8410
rect 30311 8364 30392 8410
rect 30072 8316 30392 8364
rect 30072 8270 30265 8316
rect 30311 8270 30392 8316
rect 30072 8222 30392 8270
rect 30072 8176 30265 8222
rect 30311 8176 30392 8222
rect 30072 8128 30392 8176
rect 30072 8082 30265 8128
rect 30311 8082 30392 8128
rect 30072 8034 30392 8082
rect 30072 7988 30265 8034
rect 30311 7988 30392 8034
rect 30072 7940 30392 7988
rect 30072 7894 30265 7940
rect 30311 7894 30392 7940
rect 30072 7846 30392 7894
rect 30072 7800 30265 7846
rect 30311 7800 30392 7846
rect 30072 7752 30392 7800
rect 30072 7706 30265 7752
rect 30311 7706 30392 7752
rect 30072 7658 30392 7706
rect 30072 7612 30265 7658
rect 30311 7612 30392 7658
rect 30072 7564 30392 7612
rect 30072 7541 30265 7564
rect 27303 7518 30265 7541
rect 30311 7518 30392 7564
rect 18055 7470 30392 7518
rect 18055 7424 18136 7470
rect 18182 7424 21144 7470
rect 21190 7424 23288 7470
rect 23334 7424 26296 7470
rect 26342 7424 27257 7470
rect 27303 7424 30265 7470
rect 30311 7424 30392 7470
rect 18055 7376 30392 7424
rect 18055 7330 18136 7376
rect 18182 7330 18230 7376
rect 18276 7330 18324 7376
rect 18370 7330 18418 7376
rect 18464 7330 18512 7376
rect 18558 7330 18606 7376
rect 18652 7330 18700 7376
rect 18746 7330 18794 7376
rect 18840 7330 18888 7376
rect 18934 7330 18982 7376
rect 19028 7330 19076 7376
rect 19122 7330 19170 7376
rect 19216 7330 19264 7376
rect 19310 7330 19358 7376
rect 19404 7330 19452 7376
rect 19498 7330 19546 7376
rect 19592 7330 19640 7376
rect 19686 7330 19734 7376
rect 19780 7330 19828 7376
rect 19874 7330 19922 7376
rect 19968 7330 20016 7376
rect 20062 7330 20110 7376
rect 20156 7330 20204 7376
rect 20250 7330 20298 7376
rect 20344 7330 20392 7376
rect 20438 7330 20486 7376
rect 20532 7330 20580 7376
rect 20626 7330 20674 7376
rect 20720 7330 20768 7376
rect 20814 7330 20862 7376
rect 20908 7330 20956 7376
rect 21002 7330 21050 7376
rect 21096 7330 21144 7376
rect 21190 7330 23288 7376
rect 23334 7330 23382 7376
rect 23428 7330 23476 7376
rect 23522 7330 23570 7376
rect 23616 7330 23664 7376
rect 23710 7330 23758 7376
rect 23804 7330 23852 7376
rect 23898 7330 23946 7376
rect 23992 7330 24040 7376
rect 24086 7330 24134 7376
rect 24180 7330 24228 7376
rect 24274 7330 24322 7376
rect 24368 7330 24416 7376
rect 24462 7330 24510 7376
rect 24556 7330 24604 7376
rect 24650 7330 24698 7376
rect 24744 7330 24792 7376
rect 24838 7330 24886 7376
rect 24932 7330 24980 7376
rect 25026 7330 25074 7376
rect 25120 7330 25168 7376
rect 25214 7330 25262 7376
rect 25308 7330 25356 7376
rect 25402 7330 25450 7376
rect 25496 7330 25544 7376
rect 25590 7330 25638 7376
rect 25684 7330 25732 7376
rect 25778 7330 25826 7376
rect 25872 7330 25920 7376
rect 25966 7330 26014 7376
rect 26060 7330 26108 7376
rect 26154 7330 26202 7376
rect 26248 7330 26296 7376
rect 26342 7330 27257 7376
rect 27303 7330 27351 7376
rect 27397 7330 27445 7376
rect 27491 7330 27539 7376
rect 27585 7330 27633 7376
rect 27679 7330 27727 7376
rect 27773 7330 27821 7376
rect 27867 7330 27915 7376
rect 27961 7330 28009 7376
rect 28055 7330 28103 7376
rect 28149 7330 28197 7376
rect 28243 7330 28291 7376
rect 28337 7330 28385 7376
rect 28431 7330 28479 7376
rect 28525 7330 28573 7376
rect 28619 7330 28667 7376
rect 28713 7330 28761 7376
rect 28807 7330 28855 7376
rect 28901 7330 28949 7376
rect 28995 7330 29043 7376
rect 29089 7330 29137 7376
rect 29183 7330 29231 7376
rect 29277 7330 29325 7376
rect 29371 7330 29419 7376
rect 29465 7330 29513 7376
rect 29559 7330 29607 7376
rect 29653 7330 29701 7376
rect 29747 7330 29795 7376
rect 29841 7330 29889 7376
rect 29935 7330 29983 7376
rect 30029 7330 30077 7376
rect 30123 7330 30171 7376
rect 30217 7330 30265 7376
rect 30311 7330 30392 7376
rect 18055 7221 30392 7330
rect 32510 13917 66018 14237
rect 32510 12339 32830 13917
rect 36646 12339 36966 13917
rect 37919 13913 39343 13917
rect 40746 12339 41066 13917
rect 42206 12339 42526 13917
rect 46342 12339 46662 13917
rect 50442 12339 50762 13917
rect 51938 12339 52258 13917
rect 56038 12339 56358 13917
rect 60138 12339 60458 13917
rect 61598 12339 61918 13917
rect 65698 12339 66018 13917
rect 66914 13048 67702 13060
rect 66914 12996 66926 13048
rect 66978 12996 67030 13048
rect 67082 12996 67134 13048
rect 67186 12996 67702 13048
rect 66914 12944 67702 12996
rect 66914 12892 66926 12944
rect 66978 12892 67030 12944
rect 67082 12892 67134 12944
rect 67186 12892 67702 12944
rect 66914 12840 67702 12892
rect 66914 12788 66926 12840
rect 66978 12788 67030 12840
rect 67082 12788 67134 12840
rect 67186 12788 67702 12840
rect 66914 12776 67702 12788
rect 32510 12219 66018 12339
rect 32510 12173 32629 12219
rect 32675 12173 32723 12219
rect 32769 12173 32817 12219
rect 32863 12173 32911 12219
rect 32957 12173 33005 12219
rect 33051 12173 33099 12219
rect 33145 12173 33193 12219
rect 33239 12173 33287 12219
rect 33333 12173 33381 12219
rect 33427 12173 33475 12219
rect 33521 12173 33569 12219
rect 33615 12173 33663 12219
rect 33709 12173 33757 12219
rect 33803 12173 33851 12219
rect 33897 12173 33945 12219
rect 33991 12173 34039 12219
rect 34085 12173 34133 12219
rect 34179 12173 34227 12219
rect 34273 12173 34321 12219
rect 34367 12173 34415 12219
rect 34461 12173 34509 12219
rect 34555 12173 34603 12219
rect 34649 12173 34697 12219
rect 34743 12173 34791 12219
rect 34837 12173 34885 12219
rect 34931 12173 34979 12219
rect 35025 12173 35073 12219
rect 35119 12173 35167 12219
rect 35213 12173 35261 12219
rect 35307 12173 35355 12219
rect 35401 12173 35449 12219
rect 35495 12173 35543 12219
rect 35589 12173 35637 12219
rect 35683 12173 35731 12219
rect 35777 12173 35825 12219
rect 35871 12173 35919 12219
rect 35965 12173 36013 12219
rect 36059 12173 36107 12219
rect 36153 12173 36201 12219
rect 36247 12173 36295 12219
rect 36341 12173 36389 12219
rect 36435 12173 36483 12219
rect 36529 12173 36577 12219
rect 36623 12173 36671 12219
rect 36717 12173 36765 12219
rect 36811 12173 36859 12219
rect 36905 12173 36953 12219
rect 36999 12173 37047 12219
rect 37093 12173 37141 12219
rect 37187 12173 37235 12219
rect 37281 12173 37329 12219
rect 37375 12173 37423 12219
rect 37469 12173 37517 12219
rect 37563 12173 37611 12219
rect 37657 12173 37705 12219
rect 37751 12173 37799 12219
rect 37845 12173 37893 12219
rect 37939 12173 37987 12219
rect 38033 12173 38081 12219
rect 38127 12173 38175 12219
rect 38221 12173 38269 12219
rect 38315 12173 38363 12219
rect 38409 12173 38457 12219
rect 38503 12173 38551 12219
rect 38597 12173 38645 12219
rect 38691 12173 38739 12219
rect 38785 12173 38833 12219
rect 38879 12173 38927 12219
rect 38973 12173 39021 12219
rect 39067 12173 39115 12219
rect 39161 12173 39209 12219
rect 39255 12173 39303 12219
rect 39349 12173 39397 12219
rect 39443 12173 39491 12219
rect 39537 12173 39585 12219
rect 39631 12173 39679 12219
rect 39725 12173 39773 12219
rect 39819 12173 39867 12219
rect 39913 12173 39961 12219
rect 40007 12173 40055 12219
rect 40101 12173 40149 12219
rect 40195 12173 40243 12219
rect 40289 12173 40337 12219
rect 40383 12173 40431 12219
rect 40477 12173 40525 12219
rect 40571 12173 40619 12219
rect 40665 12173 40713 12219
rect 40759 12173 40807 12219
rect 40853 12173 40901 12219
rect 40947 12173 42325 12219
rect 42371 12173 42419 12219
rect 42465 12173 42513 12219
rect 42559 12173 42607 12219
rect 42653 12173 42701 12219
rect 42747 12173 42795 12219
rect 42841 12173 42889 12219
rect 42935 12173 42983 12219
rect 43029 12173 43077 12219
rect 43123 12173 43171 12219
rect 43217 12173 43265 12219
rect 43311 12173 43359 12219
rect 43405 12173 43453 12219
rect 43499 12173 43547 12219
rect 43593 12173 43641 12219
rect 43687 12173 43735 12219
rect 43781 12173 43829 12219
rect 43875 12173 43923 12219
rect 43969 12173 44017 12219
rect 44063 12173 44111 12219
rect 44157 12173 44205 12219
rect 44251 12173 44299 12219
rect 44345 12173 44393 12219
rect 44439 12173 44487 12219
rect 44533 12173 44581 12219
rect 44627 12173 44675 12219
rect 44721 12173 44769 12219
rect 44815 12173 44863 12219
rect 44909 12173 44957 12219
rect 45003 12173 45051 12219
rect 45097 12173 45145 12219
rect 45191 12173 45239 12219
rect 45285 12173 45333 12219
rect 45379 12173 45427 12219
rect 45473 12173 45521 12219
rect 45567 12173 45615 12219
rect 45661 12173 45709 12219
rect 45755 12173 45803 12219
rect 45849 12173 45897 12219
rect 45943 12173 45991 12219
rect 46037 12173 46085 12219
rect 46131 12173 46179 12219
rect 46225 12173 46273 12219
rect 46319 12173 46367 12219
rect 46413 12173 46461 12219
rect 46507 12173 46555 12219
rect 46601 12173 46649 12219
rect 46695 12173 46743 12219
rect 46789 12173 46837 12219
rect 46883 12173 46931 12219
rect 46977 12173 47025 12219
rect 47071 12173 47119 12219
rect 47165 12173 47213 12219
rect 47259 12173 47307 12219
rect 47353 12173 47401 12219
rect 47447 12173 47495 12219
rect 47541 12173 47589 12219
rect 47635 12173 47683 12219
rect 47729 12173 47777 12219
rect 47823 12173 47871 12219
rect 47917 12173 47965 12219
rect 48011 12173 48059 12219
rect 48105 12173 48153 12219
rect 48199 12173 48247 12219
rect 48293 12173 48341 12219
rect 48387 12173 48435 12219
rect 48481 12173 48529 12219
rect 48575 12173 48623 12219
rect 48669 12173 48717 12219
rect 48763 12173 48811 12219
rect 48857 12173 48905 12219
rect 48951 12173 48999 12219
rect 49045 12173 49093 12219
rect 49139 12173 49187 12219
rect 49233 12173 49281 12219
rect 49327 12173 49375 12219
rect 49421 12173 49469 12219
rect 49515 12173 49563 12219
rect 49609 12173 49657 12219
rect 49703 12173 49751 12219
rect 49797 12173 49845 12219
rect 49891 12173 49939 12219
rect 49985 12173 50033 12219
rect 50079 12173 50127 12219
rect 50173 12173 50221 12219
rect 50267 12173 50315 12219
rect 50361 12173 50409 12219
rect 50455 12173 50503 12219
rect 50549 12173 50597 12219
rect 50643 12173 52021 12219
rect 52067 12173 52115 12219
rect 52161 12173 52209 12219
rect 52255 12173 52303 12219
rect 52349 12173 52397 12219
rect 52443 12173 52491 12219
rect 52537 12173 52585 12219
rect 52631 12173 52679 12219
rect 52725 12173 52773 12219
rect 52819 12173 52867 12219
rect 52913 12173 52961 12219
rect 53007 12173 53055 12219
rect 53101 12173 53149 12219
rect 53195 12173 53243 12219
rect 53289 12173 53337 12219
rect 53383 12173 53431 12219
rect 53477 12173 53525 12219
rect 53571 12173 53619 12219
rect 53665 12173 53713 12219
rect 53759 12173 53807 12219
rect 53853 12173 53901 12219
rect 53947 12173 53995 12219
rect 54041 12173 54089 12219
rect 54135 12173 54183 12219
rect 54229 12173 54277 12219
rect 54323 12173 54371 12219
rect 54417 12173 54465 12219
rect 54511 12173 54559 12219
rect 54605 12173 54653 12219
rect 54699 12173 54747 12219
rect 54793 12173 54841 12219
rect 54887 12173 54935 12219
rect 54981 12173 55029 12219
rect 55075 12173 55123 12219
rect 55169 12173 55217 12219
rect 55263 12173 55311 12219
rect 55357 12173 55405 12219
rect 55451 12173 55499 12219
rect 55545 12173 55593 12219
rect 55639 12173 55687 12219
rect 55733 12173 55781 12219
rect 55827 12173 55875 12219
rect 55921 12173 55969 12219
rect 56015 12173 56063 12219
rect 56109 12173 56157 12219
rect 56203 12173 56251 12219
rect 56297 12173 56345 12219
rect 56391 12173 56439 12219
rect 56485 12173 56533 12219
rect 56579 12173 56627 12219
rect 56673 12173 56721 12219
rect 56767 12173 56815 12219
rect 56861 12173 56909 12219
rect 56955 12173 57003 12219
rect 57049 12173 57097 12219
rect 57143 12173 57191 12219
rect 57237 12173 57285 12219
rect 57331 12173 57379 12219
rect 57425 12173 57473 12219
rect 57519 12173 57567 12219
rect 57613 12173 57661 12219
rect 57707 12173 57755 12219
rect 57801 12173 57849 12219
rect 57895 12173 57943 12219
rect 57989 12173 58037 12219
rect 58083 12173 58131 12219
rect 58177 12173 58225 12219
rect 58271 12173 58319 12219
rect 58365 12173 58413 12219
rect 58459 12173 58507 12219
rect 58553 12173 58601 12219
rect 58647 12173 58695 12219
rect 58741 12173 58789 12219
rect 58835 12173 58883 12219
rect 58929 12173 58977 12219
rect 59023 12173 59071 12219
rect 59117 12173 59165 12219
rect 59211 12173 59259 12219
rect 59305 12173 59353 12219
rect 59399 12173 59447 12219
rect 59493 12173 59541 12219
rect 59587 12173 59635 12219
rect 59681 12173 59729 12219
rect 59775 12173 59823 12219
rect 59869 12173 59917 12219
rect 59963 12173 60011 12219
rect 60057 12173 60105 12219
rect 60151 12173 60199 12219
rect 60245 12173 60293 12219
rect 60339 12173 61717 12219
rect 61763 12173 61811 12219
rect 61857 12173 61905 12219
rect 61951 12173 61999 12219
rect 62045 12173 62093 12219
rect 62139 12173 62187 12219
rect 62233 12173 62281 12219
rect 62327 12173 62375 12219
rect 62421 12173 62469 12219
rect 62515 12173 62563 12219
rect 62609 12173 62657 12219
rect 62703 12173 62751 12219
rect 62797 12173 62845 12219
rect 62891 12173 62939 12219
rect 62985 12173 63033 12219
rect 63079 12173 63127 12219
rect 63173 12173 63221 12219
rect 63267 12173 63315 12219
rect 63361 12173 63409 12219
rect 63455 12173 63503 12219
rect 63549 12173 63597 12219
rect 63643 12173 63691 12219
rect 63737 12173 63785 12219
rect 63831 12173 63879 12219
rect 63925 12173 63973 12219
rect 64019 12173 64067 12219
rect 64113 12173 64161 12219
rect 64207 12173 64255 12219
rect 64301 12173 64349 12219
rect 64395 12173 64443 12219
rect 64489 12173 64537 12219
rect 64583 12173 64631 12219
rect 64677 12173 64725 12219
rect 64771 12173 64819 12219
rect 64865 12173 64913 12219
rect 64959 12173 65007 12219
rect 65053 12173 65101 12219
rect 65147 12173 65195 12219
rect 65241 12173 65289 12219
rect 65335 12173 65383 12219
rect 65429 12173 65477 12219
rect 65523 12173 65571 12219
rect 65617 12173 65665 12219
rect 65711 12173 65759 12219
rect 65805 12173 65853 12219
rect 65899 12173 66018 12219
rect 32510 12125 66018 12173
rect 32510 12079 32629 12125
rect 32675 12079 36765 12125
rect 36811 12079 40901 12125
rect 40947 12079 42325 12125
rect 42371 12079 46461 12125
rect 46507 12079 50597 12125
rect 50643 12079 52021 12125
rect 52067 12079 56157 12125
rect 56203 12079 60293 12125
rect 60339 12079 61717 12125
rect 61763 12079 65853 12125
rect 65899 12079 66018 12125
rect 32510 12031 66018 12079
rect 32510 11985 32629 12031
rect 32675 12019 36765 12031
rect 32675 11985 32830 12019
rect 32510 11937 32830 11985
rect 32510 11891 32629 11937
rect 32675 11891 32830 11937
rect 32510 11843 32830 11891
rect 32510 11797 32629 11843
rect 32675 11797 32830 11843
rect 32510 11749 32830 11797
rect 32510 11703 32629 11749
rect 32675 11703 32830 11749
rect 32510 11655 32830 11703
rect 32510 11609 32629 11655
rect 32675 11609 32830 11655
rect 32510 11561 32830 11609
rect 32510 11515 32629 11561
rect 32675 11515 32830 11561
rect 32510 11467 32830 11515
rect 32510 11421 32629 11467
rect 32675 11421 32830 11467
rect 32510 11373 32830 11421
rect 32510 11327 32629 11373
rect 32675 11327 32830 11373
rect 32510 11279 32830 11327
rect 32510 11233 32629 11279
rect 32675 11233 32830 11279
rect 32510 11185 32830 11233
rect 32510 11139 32629 11185
rect 32675 11139 32830 11185
rect 32510 11091 32830 11139
rect 32510 11045 32629 11091
rect 32675 11045 32830 11091
rect 32510 10997 32830 11045
rect 32510 10951 32629 10997
rect 32675 10951 32830 10997
rect 32510 10903 32830 10951
rect 32510 10857 32629 10903
rect 32675 10857 32830 10903
rect 32510 10809 32830 10857
rect 32510 10763 32629 10809
rect 32675 10763 32830 10809
rect 32510 10715 32830 10763
rect 32510 10669 32629 10715
rect 32675 10669 32830 10715
rect 32510 10621 32830 10669
rect 32510 10575 32629 10621
rect 32675 10575 32830 10621
rect 32510 10527 32830 10575
rect 32510 10481 32629 10527
rect 32675 10481 32830 10527
rect 32510 10433 32830 10481
rect 32510 10387 32629 10433
rect 32675 10387 32830 10433
rect 32510 10339 32830 10387
rect 32510 10293 32629 10339
rect 32675 10293 32830 10339
rect 32510 10245 32830 10293
rect 32510 10199 32629 10245
rect 32675 10199 32830 10245
rect 32510 10151 32830 10199
rect 32510 10105 32629 10151
rect 32675 10105 32830 10151
rect 32510 10057 32830 10105
rect 32510 10011 32629 10057
rect 32675 10011 32830 10057
rect 32510 9963 32830 10011
rect 32510 9917 32629 9963
rect 32675 9917 32830 9963
rect 32510 9869 32830 9917
rect 32510 9823 32629 9869
rect 32675 9823 32830 9869
rect 32510 9775 32830 9823
rect 32510 9729 32629 9775
rect 32675 9729 32830 9775
rect 32510 9681 32830 9729
rect 32510 9635 32629 9681
rect 32675 9635 32830 9681
rect 32510 9587 32830 9635
rect 32510 9541 32629 9587
rect 32675 9541 32830 9587
rect 32510 9493 32830 9541
rect 32510 9447 32629 9493
rect 32675 9447 32830 9493
rect 32510 9399 32830 9447
rect 32510 9353 32629 9399
rect 32675 9353 32830 9399
rect 32510 9305 32830 9353
rect 32510 9259 32629 9305
rect 32675 9259 32830 9305
rect 32510 9211 32830 9259
rect 32510 9165 32629 9211
rect 32675 9165 32830 9211
rect 32510 9117 32830 9165
rect 32510 9071 32629 9117
rect 32675 9071 32830 9117
rect 32510 9023 32830 9071
rect 32510 8977 32629 9023
rect 32675 8977 32830 9023
rect 32510 8929 32830 8977
rect 32510 8883 32629 8929
rect 32675 8883 32830 8929
rect 32510 8835 32830 8883
rect 32510 8789 32629 8835
rect 32675 8789 32830 8835
rect 32510 8741 32830 8789
rect 32510 8695 32629 8741
rect 32675 8695 32830 8741
rect 32510 8647 32830 8695
rect 32510 8601 32629 8647
rect 32675 8601 32830 8647
rect 32510 8553 32830 8601
rect 32510 8507 32629 8553
rect 32675 8507 32830 8553
rect 32510 8459 32830 8507
rect 32510 8413 32629 8459
rect 32675 8413 32830 8459
rect 32510 8365 32830 8413
rect 32510 8319 32629 8365
rect 32675 8319 32830 8365
rect 32510 8271 32830 8319
rect 32510 8225 32629 8271
rect 32675 8225 32830 8271
rect 32510 8177 32830 8225
rect 32510 8131 32629 8177
rect 32675 8131 32830 8177
rect 32510 8083 32830 8131
rect 32510 8037 32629 8083
rect 32675 8037 32830 8083
rect 32510 7989 32830 8037
rect 32510 7943 32629 7989
rect 32675 7943 32830 7989
rect 32510 7895 32830 7943
rect 32510 7849 32629 7895
rect 32675 7849 32830 7895
rect 32510 7801 32830 7849
rect 32510 7755 32629 7801
rect 32675 7755 32830 7801
rect 32510 7707 32830 7755
rect 32510 7661 32629 7707
rect 32675 7661 32830 7707
rect 32510 7613 32830 7661
rect 32510 7567 32629 7613
rect 32675 7579 32830 7613
rect 33129 11676 33175 12019
rect 33129 10882 33175 11102
rect 33289 11676 33335 12019
rect 33417 11676 33463 11687
rect 33402 11270 33417 11282
rect 33577 11676 33623 12019
rect 33737 11676 33783 11687
rect 33897 11676 33943 12019
rect 33463 11270 33478 11282
rect 33402 11218 33414 11270
rect 33466 11218 33478 11270
rect 33402 11166 33417 11218
rect 33463 11166 33478 11218
rect 33402 11114 33414 11166
rect 33466 11114 33478 11166
rect 33402 11102 33417 11114
rect 33463 11102 33478 11114
rect 33723 11664 33737 11676
rect 33783 11664 33799 11676
rect 33723 11612 33735 11664
rect 33787 11612 33799 11664
rect 33723 11560 33737 11612
rect 33783 11560 33799 11612
rect 33723 11508 33735 11560
rect 33787 11508 33799 11560
rect 33723 11496 33737 11508
rect 33289 10882 33335 11102
rect 33417 11091 33463 11102
rect 33129 10836 33209 10882
rect 33255 10836 33335 10882
rect 33129 10616 33175 10836
rect 33129 9556 33175 10042
rect 33129 8762 33175 8982
rect 33289 10616 33335 10836
rect 33417 10616 33463 10627
rect 33402 10210 33417 10222
rect 33577 10616 33623 11102
rect 33783 11496 33799 11508
rect 33737 11091 33783 11102
rect 34057 11676 34103 11687
rect 34042 11270 34057 11282
rect 34217 11676 34263 12019
rect 34602 11812 34678 11824
rect 34602 11760 34614 11812
rect 34666 11809 34678 11812
rect 34762 11812 34838 11824
rect 34762 11809 34774 11812
rect 34666 11760 34774 11809
rect 34826 11760 34838 11812
rect 34602 11748 34838 11760
rect 34377 11676 34423 11687
rect 34537 11676 34583 11687
rect 34103 11270 34118 11282
rect 34042 11218 34054 11270
rect 34106 11218 34118 11270
rect 34042 11166 34057 11218
rect 34103 11166 34118 11218
rect 34042 11114 34054 11166
rect 34106 11114 34118 11166
rect 34042 11102 34057 11114
rect 34103 11102 34118 11114
rect 34363 11664 34377 11676
rect 34423 11664 34439 11676
rect 34363 11612 34375 11664
rect 34427 11612 34439 11664
rect 34363 11560 34377 11612
rect 34423 11560 34439 11612
rect 34363 11508 34375 11560
rect 34427 11508 34439 11560
rect 34363 11496 34377 11508
rect 33737 10616 33783 10627
rect 33897 10616 33943 11102
rect 34057 11091 34103 11102
rect 34217 11045 34263 11102
rect 34423 11496 34439 11508
rect 34377 11091 34423 11102
rect 34537 11045 34583 11102
rect 34697 11676 34743 11748
rect 34697 11091 34743 11102
rect 34857 11676 34903 11687
rect 35017 11676 35063 11687
rect 35177 11676 35223 12019
rect 35003 11664 35017 11676
rect 35063 11664 35079 11676
rect 35003 11612 35015 11664
rect 35067 11612 35079 11664
rect 35003 11560 35017 11612
rect 35063 11560 35079 11612
rect 35003 11508 35015 11560
rect 35067 11508 35079 11560
rect 35003 11496 35017 11508
rect 34857 11045 34903 11102
rect 35063 11496 35079 11508
rect 35017 11091 35063 11102
rect 35337 11676 35383 11687
rect 35322 11270 35337 11282
rect 35497 11676 35543 12019
rect 35657 11676 35703 11687
rect 35817 11676 35863 12019
rect 35383 11270 35398 11282
rect 35322 11218 35334 11270
rect 35386 11218 35398 11270
rect 35322 11166 35337 11218
rect 35383 11166 35398 11218
rect 35322 11114 35334 11166
rect 35386 11114 35398 11166
rect 35322 11102 35337 11114
rect 35383 11102 35398 11114
rect 35643 11664 35657 11676
rect 35703 11664 35719 11676
rect 35643 11612 35655 11664
rect 35707 11612 35719 11664
rect 35643 11560 35657 11612
rect 35703 11560 35719 11612
rect 35643 11508 35655 11560
rect 35707 11508 35719 11560
rect 35643 11496 35657 11508
rect 34217 10999 34903 11045
rect 33463 10210 33478 10222
rect 33402 10158 33414 10210
rect 33466 10158 33478 10210
rect 33402 10106 33417 10158
rect 33463 10106 33478 10158
rect 33402 10054 33414 10106
rect 33466 10054 33478 10106
rect 33402 10042 33417 10054
rect 33463 10042 33478 10054
rect 33723 10604 33737 10616
rect 33783 10604 33799 10616
rect 33723 10552 33735 10604
rect 33787 10552 33799 10604
rect 33723 10500 33737 10552
rect 33783 10500 33799 10552
rect 33723 10448 33735 10500
rect 33787 10448 33799 10500
rect 33723 10436 33737 10448
rect 33289 9556 33335 10042
rect 33417 10031 33463 10042
rect 33417 9556 33463 9567
rect 33402 9150 33417 9162
rect 33577 9556 33623 10042
rect 33783 10436 33799 10448
rect 33737 10031 33783 10042
rect 34057 10616 34103 10627
rect 34042 10210 34057 10222
rect 34217 10616 34263 10999
rect 34602 10752 34678 10764
rect 34602 10700 34614 10752
rect 34666 10749 34678 10752
rect 34762 10752 34838 10764
rect 34762 10749 34774 10752
rect 34666 10700 34774 10749
rect 34826 10700 34838 10752
rect 34602 10688 34838 10700
rect 34377 10616 34423 10627
rect 34537 10616 34583 10627
rect 34103 10210 34118 10222
rect 34042 10158 34054 10210
rect 34106 10158 34118 10210
rect 34042 10106 34057 10158
rect 34103 10106 34118 10158
rect 34042 10054 34054 10106
rect 34106 10054 34118 10106
rect 34042 10042 34057 10054
rect 34103 10042 34118 10054
rect 34363 10604 34377 10616
rect 34423 10604 34439 10616
rect 34363 10552 34375 10604
rect 34427 10552 34439 10604
rect 34363 10500 34377 10552
rect 34423 10500 34439 10552
rect 34363 10448 34375 10500
rect 34427 10448 34439 10500
rect 34363 10436 34377 10448
rect 33737 9556 33783 9567
rect 33897 9556 33943 10042
rect 34057 10031 34103 10042
rect 34217 9985 34263 10042
rect 34423 10436 34439 10448
rect 34377 10031 34423 10042
rect 34537 9985 34583 10042
rect 34697 10616 34743 10688
rect 34697 10031 34743 10042
rect 34857 10616 34903 10627
rect 35017 10616 35063 10627
rect 35177 10616 35223 11102
rect 35337 11091 35383 11102
rect 35003 10604 35017 10616
rect 35063 10604 35079 10616
rect 35003 10552 35015 10604
rect 35067 10552 35079 10604
rect 35003 10500 35017 10552
rect 35063 10500 35079 10552
rect 35003 10448 35015 10500
rect 35067 10448 35079 10500
rect 35003 10436 35017 10448
rect 34857 9985 34903 10042
rect 35063 10436 35079 10448
rect 35017 10031 35063 10042
rect 35337 10616 35383 10627
rect 35322 10210 35337 10222
rect 35497 10616 35543 11102
rect 35703 11496 35719 11508
rect 35657 11091 35703 11102
rect 35977 11676 36023 11687
rect 35962 11270 35977 11282
rect 36105 11676 36151 12019
rect 36023 11270 36038 11282
rect 35962 11218 35974 11270
rect 36026 11218 36038 11270
rect 35962 11166 35977 11218
rect 36023 11166 36038 11218
rect 35962 11114 35974 11166
rect 36026 11114 36038 11166
rect 35962 11102 35977 11114
rect 36023 11102 36038 11114
rect 35657 10616 35703 10627
rect 35817 10616 35863 11102
rect 35977 11091 36023 11102
rect 36105 10882 36151 11102
rect 36265 11676 36311 12019
rect 36265 10882 36311 11102
rect 36105 10836 36185 10882
rect 36231 10836 36311 10882
rect 35383 10210 35398 10222
rect 35322 10158 35334 10210
rect 35386 10158 35398 10210
rect 35322 10106 35337 10158
rect 35383 10106 35398 10158
rect 35322 10054 35334 10106
rect 35386 10054 35398 10106
rect 35322 10042 35337 10054
rect 35383 10042 35398 10054
rect 35643 10604 35657 10616
rect 35703 10604 35719 10616
rect 35643 10552 35655 10604
rect 35707 10552 35719 10604
rect 35643 10500 35657 10552
rect 35703 10500 35719 10552
rect 35643 10448 35655 10500
rect 35707 10448 35719 10500
rect 35643 10436 35657 10448
rect 34217 9939 34903 9985
rect 33463 9150 33478 9162
rect 33402 9098 33414 9150
rect 33466 9098 33478 9150
rect 33402 9046 33417 9098
rect 33463 9046 33478 9098
rect 33402 8994 33414 9046
rect 33466 8994 33478 9046
rect 33402 8982 33417 8994
rect 33463 8982 33478 8994
rect 33723 9544 33737 9556
rect 33783 9544 33799 9556
rect 33723 9492 33735 9544
rect 33787 9492 33799 9544
rect 33723 9440 33737 9492
rect 33783 9440 33799 9492
rect 33723 9388 33735 9440
rect 33787 9388 33799 9440
rect 33723 9376 33737 9388
rect 33289 8762 33335 8982
rect 33417 8971 33463 8982
rect 33129 8716 33209 8762
rect 33255 8716 33335 8762
rect 33129 8496 33175 8716
rect 33129 7579 33175 7922
rect 33289 8496 33335 8716
rect 33417 8496 33463 8507
rect 33402 8090 33417 8102
rect 33577 8496 33623 8982
rect 33783 9376 33799 9388
rect 33737 8971 33783 8982
rect 34057 9556 34103 9567
rect 34042 9150 34057 9162
rect 34217 9556 34263 9939
rect 34602 9692 34678 9704
rect 34602 9640 34614 9692
rect 34666 9689 34678 9692
rect 34762 9692 34838 9704
rect 34762 9689 34774 9692
rect 34666 9640 34774 9689
rect 34826 9640 34838 9692
rect 34602 9628 34838 9640
rect 34377 9556 34423 9567
rect 34537 9556 34583 9567
rect 34103 9150 34118 9162
rect 34042 9098 34054 9150
rect 34106 9098 34118 9150
rect 34042 9046 34057 9098
rect 34103 9046 34118 9098
rect 34042 8994 34054 9046
rect 34106 8994 34118 9046
rect 34042 8982 34057 8994
rect 34103 8982 34118 8994
rect 34363 9544 34377 9556
rect 34423 9544 34439 9556
rect 34363 9492 34375 9544
rect 34427 9492 34439 9544
rect 34363 9440 34377 9492
rect 34423 9440 34439 9492
rect 34363 9388 34375 9440
rect 34427 9388 34439 9440
rect 34363 9376 34377 9388
rect 33737 8496 33783 8507
rect 33897 8496 33943 8982
rect 34057 8971 34103 8982
rect 34217 8925 34263 8982
rect 34423 9376 34439 9388
rect 34377 8971 34423 8982
rect 34537 8925 34583 8982
rect 34697 9556 34743 9628
rect 34697 8971 34743 8982
rect 34857 9556 34903 9567
rect 35017 9556 35063 9567
rect 35177 9556 35223 10042
rect 35337 10031 35383 10042
rect 35003 9544 35017 9556
rect 35063 9544 35079 9556
rect 35003 9492 35015 9544
rect 35067 9492 35079 9544
rect 35003 9440 35017 9492
rect 35063 9440 35079 9492
rect 35003 9388 35015 9440
rect 35067 9388 35079 9440
rect 35003 9376 35017 9388
rect 34857 8925 34903 8982
rect 35063 9376 35079 9388
rect 35017 8971 35063 8982
rect 35337 9556 35383 9567
rect 35322 9150 35337 9162
rect 35497 9556 35543 10042
rect 35703 10436 35719 10448
rect 35657 10031 35703 10042
rect 35977 10616 36023 10627
rect 35962 10210 35977 10222
rect 36105 10616 36151 10836
rect 36023 10210 36038 10222
rect 35962 10158 35974 10210
rect 36026 10158 36038 10210
rect 35962 10106 35977 10158
rect 36023 10106 36038 10158
rect 35962 10054 35974 10106
rect 36026 10054 36038 10106
rect 35962 10042 35977 10054
rect 36023 10042 36038 10054
rect 35657 9556 35703 9567
rect 35817 9556 35863 10042
rect 35977 10031 36023 10042
rect 35383 9150 35398 9162
rect 35322 9098 35334 9150
rect 35386 9098 35398 9150
rect 35322 9046 35337 9098
rect 35383 9046 35398 9098
rect 35322 8994 35334 9046
rect 35386 8994 35398 9046
rect 35322 8982 35337 8994
rect 35383 8982 35398 8994
rect 35643 9544 35657 9556
rect 35703 9544 35719 9556
rect 35643 9492 35655 9544
rect 35707 9492 35719 9544
rect 35643 9440 35657 9492
rect 35703 9440 35719 9492
rect 35643 9388 35655 9440
rect 35707 9388 35719 9440
rect 35643 9376 35657 9388
rect 34217 8879 34903 8925
rect 33463 8090 33478 8102
rect 33402 8038 33414 8090
rect 33466 8038 33478 8090
rect 33402 7986 33417 8038
rect 33463 7986 33478 8038
rect 33402 7934 33414 7986
rect 33466 7934 33478 7986
rect 33402 7922 33417 7934
rect 33463 7922 33478 7934
rect 33723 8484 33737 8496
rect 33783 8484 33799 8496
rect 33723 8432 33735 8484
rect 33787 8432 33799 8484
rect 33723 8380 33737 8432
rect 33783 8380 33799 8432
rect 33723 8328 33735 8380
rect 33787 8328 33799 8380
rect 33723 8316 33737 8328
rect 33289 7579 33335 7922
rect 33417 7911 33463 7922
rect 33577 7579 33623 7922
rect 33783 8316 33799 8328
rect 33737 7911 33783 7922
rect 34057 8496 34103 8507
rect 34042 8090 34057 8102
rect 34217 8496 34263 8879
rect 34602 8632 34678 8644
rect 34602 8580 34614 8632
rect 34666 8629 34678 8632
rect 34762 8632 34838 8644
rect 34762 8629 34774 8632
rect 34666 8580 34774 8629
rect 34826 8580 34838 8632
rect 34602 8568 34838 8580
rect 34377 8496 34423 8507
rect 34537 8496 34583 8507
rect 34103 8090 34118 8102
rect 34042 8038 34054 8090
rect 34106 8038 34118 8090
rect 34042 7986 34057 8038
rect 34103 7986 34118 8038
rect 34042 7934 34054 7986
rect 34106 7934 34118 7986
rect 34042 7922 34057 7934
rect 34103 7922 34118 7934
rect 34363 8484 34377 8496
rect 34423 8484 34439 8496
rect 34363 8432 34375 8484
rect 34427 8432 34439 8484
rect 34363 8380 34377 8432
rect 34423 8380 34439 8432
rect 34363 8328 34375 8380
rect 34427 8328 34439 8380
rect 34363 8316 34377 8328
rect 33897 7579 33943 7922
rect 34057 7911 34103 7922
rect 34217 7579 34263 7922
rect 34423 8316 34439 8328
rect 34377 7911 34423 7922
rect 34537 7579 34583 7922
rect 34697 8496 34743 8568
rect 34697 7911 34743 7922
rect 34857 8496 34903 8507
rect 35017 8496 35063 8507
rect 35177 8496 35223 8982
rect 35337 8971 35383 8982
rect 35003 8484 35017 8496
rect 35063 8484 35079 8496
rect 35003 8432 35015 8484
rect 35067 8432 35079 8484
rect 35003 8380 35017 8432
rect 35063 8380 35079 8432
rect 35003 8328 35015 8380
rect 35067 8328 35079 8380
rect 35003 8316 35017 8328
rect 34857 7579 34903 7922
rect 35063 8316 35079 8328
rect 35017 7911 35063 7922
rect 35337 8496 35383 8507
rect 35322 8090 35337 8102
rect 35497 8496 35543 8982
rect 35703 9376 35719 9388
rect 35657 8971 35703 8982
rect 35977 9556 36023 9567
rect 35962 9150 35977 9162
rect 36105 9556 36151 10042
rect 36023 9150 36038 9162
rect 35962 9098 35974 9150
rect 36026 9098 36038 9150
rect 35962 9046 35977 9098
rect 36023 9046 36038 9098
rect 35962 8994 35974 9046
rect 36026 8994 36038 9046
rect 35962 8982 35977 8994
rect 36023 8982 36038 8994
rect 35657 8496 35703 8507
rect 35817 8496 35863 8982
rect 35977 8971 36023 8982
rect 36105 8762 36151 8982
rect 36265 10616 36311 10836
rect 36265 9556 36311 10042
rect 36265 8762 36311 8982
rect 36105 8716 36185 8762
rect 36231 8716 36311 8762
rect 35383 8090 35398 8102
rect 35322 8038 35334 8090
rect 35386 8038 35398 8090
rect 35322 7986 35337 8038
rect 35383 7986 35398 8038
rect 35322 7934 35334 7986
rect 35386 7934 35398 7986
rect 35322 7922 35337 7934
rect 35383 7922 35398 7934
rect 35643 8484 35657 8496
rect 35703 8484 35719 8496
rect 35643 8432 35655 8484
rect 35707 8432 35719 8484
rect 35643 8380 35657 8432
rect 35703 8380 35719 8432
rect 35643 8328 35655 8380
rect 35707 8328 35719 8380
rect 35643 8316 35657 8328
rect 35177 7579 35223 7922
rect 35337 7911 35383 7922
rect 35497 7579 35543 7922
rect 35703 8316 35719 8328
rect 35657 7911 35703 7922
rect 35977 8496 36023 8507
rect 35962 8090 35977 8102
rect 36105 8496 36151 8716
rect 36023 8090 36038 8102
rect 35962 8038 35974 8090
rect 36026 8038 36038 8090
rect 35962 7986 35977 8038
rect 36023 7986 36038 8038
rect 35962 7934 35974 7986
rect 36026 7934 36038 7986
rect 35962 7922 35977 7934
rect 36023 7922 36038 7934
rect 35817 7579 35863 7922
rect 35977 7911 36023 7922
rect 36105 7579 36151 7922
rect 36265 8496 36311 8716
rect 36265 7579 36311 7922
rect 36610 11985 36765 12019
rect 36811 12019 40901 12031
rect 36811 11985 36966 12019
rect 36610 11937 36966 11985
rect 36610 11891 36765 11937
rect 36811 11891 36966 11937
rect 36610 11843 36966 11891
rect 36610 11797 36765 11843
rect 36811 11797 36966 11843
rect 36610 11749 36966 11797
rect 36610 11703 36765 11749
rect 36811 11703 36966 11749
rect 36610 11655 36966 11703
rect 36610 11609 36765 11655
rect 36811 11609 36966 11655
rect 36610 11561 36966 11609
rect 36610 11515 36765 11561
rect 36811 11515 36966 11561
rect 36610 11467 36966 11515
rect 36610 11421 36765 11467
rect 36811 11421 36966 11467
rect 36610 11373 36966 11421
rect 36610 11327 36765 11373
rect 36811 11327 36966 11373
rect 36610 11279 36966 11327
rect 36610 11233 36765 11279
rect 36811 11233 36966 11279
rect 36610 11185 36966 11233
rect 36610 11139 36765 11185
rect 36811 11139 36966 11185
rect 36610 11091 36966 11139
rect 36610 11045 36765 11091
rect 36811 11045 36966 11091
rect 36610 10997 36966 11045
rect 36610 10951 36765 10997
rect 36811 10951 36966 10997
rect 36610 10903 36966 10951
rect 36610 10857 36765 10903
rect 36811 10857 36966 10903
rect 36610 10809 36966 10857
rect 36610 10763 36765 10809
rect 36811 10763 36966 10809
rect 36610 10715 36966 10763
rect 36610 10669 36765 10715
rect 36811 10669 36966 10715
rect 36610 10621 36966 10669
rect 36610 10575 36765 10621
rect 36811 10575 36966 10621
rect 36610 10527 36966 10575
rect 36610 10481 36765 10527
rect 36811 10481 36966 10527
rect 36610 10433 36966 10481
rect 36610 10387 36765 10433
rect 36811 10387 36966 10433
rect 36610 10339 36966 10387
rect 36610 10293 36765 10339
rect 36811 10293 36966 10339
rect 36610 10245 36966 10293
rect 36610 10199 36765 10245
rect 36811 10199 36966 10245
rect 36610 10151 36966 10199
rect 36610 10105 36765 10151
rect 36811 10105 36966 10151
rect 36610 10057 36966 10105
rect 36610 10011 36765 10057
rect 36811 10011 36966 10057
rect 36610 9963 36966 10011
rect 36610 9917 36765 9963
rect 36811 9917 36966 9963
rect 36610 9869 36966 9917
rect 36610 9823 36765 9869
rect 36811 9823 36966 9869
rect 36610 9775 36966 9823
rect 36610 9729 36765 9775
rect 36811 9729 36966 9775
rect 36610 9681 36966 9729
rect 36610 9635 36765 9681
rect 36811 9635 36966 9681
rect 36610 9587 36966 9635
rect 36610 9541 36765 9587
rect 36811 9541 36966 9587
rect 36610 9493 36966 9541
rect 36610 9447 36765 9493
rect 36811 9447 36966 9493
rect 36610 9399 36966 9447
rect 36610 9353 36765 9399
rect 36811 9353 36966 9399
rect 36610 9305 36966 9353
rect 36610 9259 36765 9305
rect 36811 9259 36966 9305
rect 36610 9211 36966 9259
rect 36610 9165 36765 9211
rect 36811 9165 36966 9211
rect 36610 9117 36966 9165
rect 36610 9071 36765 9117
rect 36811 9071 36966 9117
rect 36610 9023 36966 9071
rect 36610 8977 36765 9023
rect 36811 8977 36966 9023
rect 36610 8929 36966 8977
rect 36610 8883 36765 8929
rect 36811 8883 36966 8929
rect 36610 8835 36966 8883
rect 36610 8789 36765 8835
rect 36811 8789 36966 8835
rect 36610 8741 36966 8789
rect 36610 8695 36765 8741
rect 36811 8695 36966 8741
rect 36610 8647 36966 8695
rect 36610 8601 36765 8647
rect 36811 8601 36966 8647
rect 36610 8553 36966 8601
rect 36610 8507 36765 8553
rect 36811 8507 36966 8553
rect 36610 8459 36966 8507
rect 36610 8413 36765 8459
rect 36811 8413 36966 8459
rect 36610 8365 36966 8413
rect 36610 8319 36765 8365
rect 36811 8319 36966 8365
rect 36610 8271 36966 8319
rect 36610 8225 36765 8271
rect 36811 8225 36966 8271
rect 36610 8177 36966 8225
rect 36610 8131 36765 8177
rect 36811 8131 36966 8177
rect 36610 8083 36966 8131
rect 36610 8037 36765 8083
rect 36811 8037 36966 8083
rect 36610 7989 36966 8037
rect 36610 7943 36765 7989
rect 36811 7943 36966 7989
rect 36610 7895 36966 7943
rect 36610 7849 36765 7895
rect 36811 7849 36966 7895
rect 36610 7801 36966 7849
rect 36610 7755 36765 7801
rect 36811 7755 36966 7801
rect 36610 7707 36966 7755
rect 36610 7661 36765 7707
rect 36811 7661 36966 7707
rect 36610 7613 36966 7661
rect 36610 7579 36765 7613
rect 32675 7567 36765 7579
rect 36811 7579 36966 7613
rect 37265 11676 37311 12019
rect 37265 10882 37311 11102
rect 37425 11676 37471 12019
rect 37553 11676 37599 11687
rect 37538 11270 37553 11282
rect 37713 11676 37759 12019
rect 37873 11676 37919 11687
rect 38033 11676 38079 12019
rect 37599 11270 37614 11282
rect 37538 11218 37550 11270
rect 37602 11218 37614 11270
rect 37538 11166 37553 11218
rect 37599 11166 37614 11218
rect 37538 11114 37550 11166
rect 37602 11114 37614 11166
rect 37538 11102 37553 11114
rect 37599 11102 37614 11114
rect 37857 11664 37873 11676
rect 37919 11664 37933 11676
rect 37857 11612 37869 11664
rect 37921 11612 37933 11664
rect 37857 11560 37873 11612
rect 37919 11560 37933 11612
rect 37857 11508 37869 11560
rect 37921 11508 37933 11560
rect 37857 11496 37873 11508
rect 37425 10882 37471 11102
rect 37553 11091 37599 11102
rect 37265 10836 37345 10882
rect 37391 10836 37471 10882
rect 37265 10616 37311 10836
rect 37265 9556 37311 10042
rect 37265 8762 37311 8982
rect 37425 10616 37471 10836
rect 37553 10616 37599 10627
rect 37538 10210 37553 10222
rect 37713 10616 37759 11102
rect 37919 11496 37933 11508
rect 37873 11091 37919 11102
rect 38193 11676 38239 11687
rect 38178 11270 38193 11282
rect 38353 11676 38399 12019
rect 38738 11812 38814 11824
rect 38738 11760 38750 11812
rect 38802 11809 38814 11812
rect 38898 11812 38974 11824
rect 38898 11809 38910 11812
rect 38802 11760 38910 11809
rect 38962 11760 38974 11812
rect 38738 11748 38974 11760
rect 38513 11676 38559 11687
rect 38673 11676 38719 11687
rect 38239 11270 38254 11282
rect 38178 11218 38190 11270
rect 38242 11218 38254 11270
rect 38178 11166 38193 11218
rect 38239 11166 38254 11218
rect 38178 11114 38190 11166
rect 38242 11114 38254 11166
rect 38178 11102 38193 11114
rect 38239 11102 38254 11114
rect 38497 11664 38513 11676
rect 38559 11664 38573 11676
rect 38497 11612 38509 11664
rect 38561 11612 38573 11664
rect 38497 11560 38513 11612
rect 38559 11560 38573 11612
rect 38497 11508 38509 11560
rect 38561 11508 38573 11560
rect 38497 11496 38513 11508
rect 37873 10616 37919 10627
rect 38033 10616 38079 11102
rect 38193 11091 38239 11102
rect 37599 10210 37614 10222
rect 37538 10158 37550 10210
rect 37602 10158 37614 10210
rect 37538 10106 37553 10158
rect 37599 10106 37614 10158
rect 37538 10054 37550 10106
rect 37602 10054 37614 10106
rect 37538 10042 37553 10054
rect 37599 10042 37614 10054
rect 37857 10604 37873 10616
rect 37919 10604 37933 10616
rect 37857 10552 37869 10604
rect 37921 10552 37933 10604
rect 37857 10500 37873 10552
rect 37919 10500 37933 10552
rect 37857 10448 37869 10500
rect 37921 10448 37933 10500
rect 37857 10436 37873 10448
rect 37425 9556 37471 10042
rect 37553 10031 37599 10042
rect 37553 9556 37599 9567
rect 37538 9150 37553 9162
rect 37713 9556 37759 10042
rect 37919 10436 37933 10448
rect 37873 10031 37919 10042
rect 38193 10616 38239 10627
rect 38178 10210 38193 10222
rect 38353 10616 38399 11102
rect 38559 11496 38573 11508
rect 38513 11091 38559 11102
rect 38673 11045 38719 11102
rect 38833 11676 38879 11748
rect 38833 11091 38879 11102
rect 38993 11676 39039 11687
rect 39153 11676 39199 11687
rect 39313 11676 39359 12019
rect 39137 11664 39153 11676
rect 39199 11664 39213 11676
rect 39137 11612 39149 11664
rect 39201 11612 39213 11664
rect 39137 11560 39153 11612
rect 39199 11560 39213 11612
rect 39137 11508 39149 11560
rect 39201 11508 39213 11560
rect 39137 11496 39153 11508
rect 38993 11045 39039 11102
rect 39199 11496 39213 11508
rect 39153 11091 39199 11102
rect 39473 11676 39519 11687
rect 39458 11270 39473 11282
rect 39633 11676 39679 12019
rect 39793 11676 39839 11687
rect 39953 11676 39999 12019
rect 39519 11270 39534 11282
rect 39458 11218 39470 11270
rect 39522 11218 39534 11270
rect 39458 11166 39473 11218
rect 39519 11166 39534 11218
rect 39458 11114 39470 11166
rect 39522 11114 39534 11166
rect 39458 11102 39473 11114
rect 39519 11102 39534 11114
rect 39777 11664 39793 11676
rect 39839 11664 39853 11676
rect 39777 11612 39789 11664
rect 39841 11612 39853 11664
rect 39777 11560 39793 11612
rect 39839 11560 39853 11612
rect 39777 11508 39789 11560
rect 39841 11508 39853 11560
rect 39777 11496 39793 11508
rect 39313 11045 39359 11102
rect 39473 11091 39519 11102
rect 38673 10999 39359 11045
rect 38738 10752 38814 10764
rect 38738 10700 38750 10752
rect 38802 10749 38814 10752
rect 38898 10752 38974 10764
rect 38898 10749 38910 10752
rect 38802 10700 38910 10749
rect 38962 10700 38974 10752
rect 38738 10688 38974 10700
rect 38513 10616 38559 10627
rect 38673 10616 38719 10627
rect 38239 10210 38254 10222
rect 38178 10158 38190 10210
rect 38242 10158 38254 10210
rect 38178 10106 38193 10158
rect 38239 10106 38254 10158
rect 38178 10054 38190 10106
rect 38242 10054 38254 10106
rect 38178 10042 38193 10054
rect 38239 10042 38254 10054
rect 38497 10604 38513 10616
rect 38559 10604 38573 10616
rect 38497 10552 38509 10604
rect 38561 10552 38573 10604
rect 38497 10500 38513 10552
rect 38559 10500 38573 10552
rect 38497 10448 38509 10500
rect 38561 10448 38573 10500
rect 38497 10436 38513 10448
rect 37873 9556 37919 9567
rect 38033 9556 38079 10042
rect 38193 10031 38239 10042
rect 37599 9150 37614 9162
rect 37538 9098 37550 9150
rect 37602 9098 37614 9150
rect 37538 9046 37553 9098
rect 37599 9046 37614 9098
rect 37538 8994 37550 9046
rect 37602 8994 37614 9046
rect 37538 8982 37553 8994
rect 37599 8982 37614 8994
rect 37857 9544 37873 9556
rect 37919 9544 37933 9556
rect 37857 9492 37869 9544
rect 37921 9492 37933 9544
rect 37857 9440 37873 9492
rect 37919 9440 37933 9492
rect 37857 9388 37869 9440
rect 37921 9388 37933 9440
rect 37857 9376 37873 9388
rect 37425 8762 37471 8982
rect 37553 8971 37599 8982
rect 37265 8716 37345 8762
rect 37391 8716 37471 8762
rect 37265 8496 37311 8716
rect 37265 7579 37311 7922
rect 37425 8496 37471 8716
rect 37553 8496 37599 8507
rect 37538 8090 37553 8102
rect 37713 8496 37759 8982
rect 37919 9376 37933 9388
rect 37873 8971 37919 8982
rect 38193 9556 38239 9567
rect 38178 9150 38193 9162
rect 38353 9556 38399 10042
rect 38559 10436 38573 10448
rect 38513 10031 38559 10042
rect 38673 9985 38719 10042
rect 38833 10616 38879 10688
rect 38833 10031 38879 10042
rect 38993 10616 39039 10627
rect 39153 10616 39199 10627
rect 39313 10616 39359 10999
rect 39137 10604 39153 10616
rect 39199 10604 39213 10616
rect 39137 10552 39149 10604
rect 39201 10552 39213 10604
rect 39137 10500 39153 10552
rect 39199 10500 39213 10552
rect 39137 10448 39149 10500
rect 39201 10448 39213 10500
rect 39137 10436 39153 10448
rect 38993 9985 39039 10042
rect 39199 10436 39213 10448
rect 39153 10031 39199 10042
rect 39473 10616 39519 10627
rect 39458 10210 39473 10222
rect 39633 10616 39679 11102
rect 39839 11496 39853 11508
rect 39793 11091 39839 11102
rect 40113 11676 40159 11687
rect 40098 11270 40113 11282
rect 40241 11676 40287 12019
rect 40159 11270 40174 11282
rect 40098 11218 40110 11270
rect 40162 11218 40174 11270
rect 40098 11166 40113 11218
rect 40159 11166 40174 11218
rect 40098 11114 40110 11166
rect 40162 11114 40174 11166
rect 40098 11102 40113 11114
rect 40159 11102 40174 11114
rect 39793 10616 39839 10627
rect 39953 10616 39999 11102
rect 40113 11091 40159 11102
rect 40241 10882 40287 11102
rect 40401 11676 40447 12019
rect 40401 10882 40447 11102
rect 40241 10836 40321 10882
rect 40367 10836 40447 10882
rect 39519 10210 39534 10222
rect 39458 10158 39470 10210
rect 39522 10158 39534 10210
rect 39458 10106 39473 10158
rect 39519 10106 39534 10158
rect 39458 10054 39470 10106
rect 39522 10054 39534 10106
rect 39458 10042 39473 10054
rect 39519 10042 39534 10054
rect 39777 10604 39793 10616
rect 39839 10604 39853 10616
rect 39777 10552 39789 10604
rect 39841 10552 39853 10604
rect 39777 10500 39793 10552
rect 39839 10500 39853 10552
rect 39777 10448 39789 10500
rect 39841 10448 39853 10500
rect 39777 10436 39793 10448
rect 39313 9985 39359 10042
rect 39473 10031 39519 10042
rect 38673 9939 39359 9985
rect 38738 9692 38814 9704
rect 38738 9640 38750 9692
rect 38802 9689 38814 9692
rect 38898 9692 38974 9704
rect 38898 9689 38910 9692
rect 38802 9640 38910 9689
rect 38962 9640 38974 9692
rect 38738 9628 38974 9640
rect 38513 9556 38559 9567
rect 38673 9556 38719 9567
rect 38239 9150 38254 9162
rect 38178 9098 38190 9150
rect 38242 9098 38254 9150
rect 38178 9046 38193 9098
rect 38239 9046 38254 9098
rect 38178 8994 38190 9046
rect 38242 8994 38254 9046
rect 38178 8982 38193 8994
rect 38239 8982 38254 8994
rect 38497 9544 38513 9556
rect 38559 9544 38573 9556
rect 38497 9492 38509 9544
rect 38561 9492 38573 9544
rect 38497 9440 38513 9492
rect 38559 9440 38573 9492
rect 38497 9388 38509 9440
rect 38561 9388 38573 9440
rect 38497 9376 38513 9388
rect 37873 8496 37919 8507
rect 38033 8496 38079 8982
rect 38193 8971 38239 8982
rect 37599 8090 37614 8102
rect 37538 8038 37550 8090
rect 37602 8038 37614 8090
rect 37538 7986 37553 8038
rect 37599 7986 37614 8038
rect 37538 7934 37550 7986
rect 37602 7934 37614 7986
rect 37538 7922 37553 7934
rect 37599 7922 37614 7934
rect 37857 8484 37873 8496
rect 37919 8484 37933 8496
rect 37857 8432 37869 8484
rect 37921 8432 37933 8484
rect 37857 8380 37873 8432
rect 37919 8380 37933 8432
rect 37857 8328 37869 8380
rect 37921 8328 37933 8380
rect 37857 8316 37873 8328
rect 37425 7579 37471 7922
rect 37553 7911 37599 7922
rect 37713 7579 37759 7922
rect 37919 8316 37933 8328
rect 37873 7911 37919 7922
rect 38193 8496 38239 8507
rect 38178 8090 38193 8102
rect 38353 8496 38399 8982
rect 38559 9376 38573 9388
rect 38513 8971 38559 8982
rect 38673 8925 38719 8982
rect 38833 9556 38879 9628
rect 38833 8971 38879 8982
rect 38993 9556 39039 9567
rect 39153 9556 39199 9567
rect 39313 9556 39359 9939
rect 39137 9544 39153 9556
rect 39199 9544 39213 9556
rect 39137 9492 39149 9544
rect 39201 9492 39213 9544
rect 39137 9440 39153 9492
rect 39199 9440 39213 9492
rect 39137 9388 39149 9440
rect 39201 9388 39213 9440
rect 39137 9376 39153 9388
rect 38993 8925 39039 8982
rect 39199 9376 39213 9388
rect 39153 8971 39199 8982
rect 39473 9556 39519 9567
rect 39458 9150 39473 9162
rect 39633 9556 39679 10042
rect 39839 10436 39853 10448
rect 39793 10031 39839 10042
rect 40113 10616 40159 10627
rect 40098 10210 40113 10222
rect 40241 10616 40287 10836
rect 40159 10210 40174 10222
rect 40098 10158 40110 10210
rect 40162 10158 40174 10210
rect 40098 10106 40113 10158
rect 40159 10106 40174 10158
rect 40098 10054 40110 10106
rect 40162 10054 40174 10106
rect 40098 10042 40113 10054
rect 40159 10042 40174 10054
rect 39793 9556 39839 9567
rect 39953 9556 39999 10042
rect 40113 10031 40159 10042
rect 39519 9150 39534 9162
rect 39458 9098 39470 9150
rect 39522 9098 39534 9150
rect 39458 9046 39473 9098
rect 39519 9046 39534 9098
rect 39458 8994 39470 9046
rect 39522 8994 39534 9046
rect 39458 8982 39473 8994
rect 39519 8982 39534 8994
rect 39777 9544 39793 9556
rect 39839 9544 39853 9556
rect 39777 9492 39789 9544
rect 39841 9492 39853 9544
rect 39777 9440 39793 9492
rect 39839 9440 39853 9492
rect 39777 9388 39789 9440
rect 39841 9388 39853 9440
rect 39777 9376 39793 9388
rect 39313 8925 39359 8982
rect 39473 8971 39519 8982
rect 38673 8879 39359 8925
rect 38738 8632 38814 8644
rect 38738 8580 38750 8632
rect 38802 8629 38814 8632
rect 38898 8632 38974 8644
rect 38898 8629 38910 8632
rect 38802 8580 38910 8629
rect 38962 8580 38974 8632
rect 38738 8568 38974 8580
rect 38513 8496 38559 8507
rect 38673 8496 38719 8507
rect 38239 8090 38254 8102
rect 38178 8038 38190 8090
rect 38242 8038 38254 8090
rect 38178 7986 38193 8038
rect 38239 7986 38254 8038
rect 38178 7934 38190 7986
rect 38242 7934 38254 7986
rect 38178 7922 38193 7934
rect 38239 7922 38254 7934
rect 38497 8484 38513 8496
rect 38559 8484 38573 8496
rect 38497 8432 38509 8484
rect 38561 8432 38573 8484
rect 38497 8380 38513 8432
rect 38559 8380 38573 8432
rect 38497 8328 38509 8380
rect 38561 8328 38573 8380
rect 38497 8316 38513 8328
rect 38033 7579 38079 7922
rect 38193 7911 38239 7922
rect 38353 7579 38399 7922
rect 38559 8316 38573 8328
rect 38513 7911 38559 7922
rect 38673 7579 38719 7922
rect 38833 8496 38879 8568
rect 38833 7911 38879 7922
rect 38993 8496 39039 8507
rect 39153 8496 39199 8507
rect 39313 8496 39359 8879
rect 39137 8484 39153 8496
rect 39199 8484 39213 8496
rect 39137 8432 39149 8484
rect 39201 8432 39213 8484
rect 39137 8380 39153 8432
rect 39199 8380 39213 8432
rect 39137 8328 39149 8380
rect 39201 8328 39213 8380
rect 39137 8316 39153 8328
rect 38993 7579 39039 7922
rect 39199 8316 39213 8328
rect 39153 7911 39199 7922
rect 39473 8496 39519 8507
rect 39458 8090 39473 8102
rect 39633 8496 39679 8982
rect 39839 9376 39853 9388
rect 39793 8971 39839 8982
rect 40113 9556 40159 9567
rect 40098 9150 40113 9162
rect 40241 9556 40287 10042
rect 40159 9150 40174 9162
rect 40098 9098 40110 9150
rect 40162 9098 40174 9150
rect 40098 9046 40113 9098
rect 40159 9046 40174 9098
rect 40098 8994 40110 9046
rect 40162 8994 40174 9046
rect 40098 8982 40113 8994
rect 40159 8982 40174 8994
rect 39793 8496 39839 8507
rect 39953 8496 39999 8982
rect 40113 8971 40159 8982
rect 40241 8762 40287 8982
rect 40401 10616 40447 10836
rect 40401 9556 40447 10042
rect 40401 8762 40447 8982
rect 40241 8716 40321 8762
rect 40367 8716 40447 8762
rect 39519 8090 39534 8102
rect 39458 8038 39470 8090
rect 39522 8038 39534 8090
rect 39458 7986 39473 8038
rect 39519 7986 39534 8038
rect 39458 7934 39470 7986
rect 39522 7934 39534 7986
rect 39458 7922 39473 7934
rect 39519 7922 39534 7934
rect 39777 8484 39793 8496
rect 39839 8484 39853 8496
rect 39777 8432 39789 8484
rect 39841 8432 39853 8484
rect 39777 8380 39793 8432
rect 39839 8380 39853 8432
rect 39777 8328 39789 8380
rect 39841 8328 39853 8380
rect 39777 8316 39793 8328
rect 39313 7579 39359 7922
rect 39473 7911 39519 7922
rect 39633 7579 39679 7922
rect 39839 8316 39853 8328
rect 39793 7911 39839 7922
rect 40113 8496 40159 8507
rect 40098 8090 40113 8102
rect 40241 8496 40287 8716
rect 40159 8090 40174 8102
rect 40098 8038 40110 8090
rect 40162 8038 40174 8090
rect 40098 7986 40113 8038
rect 40159 7986 40174 8038
rect 40098 7934 40110 7986
rect 40162 7934 40174 7986
rect 40098 7922 40113 7934
rect 40159 7922 40174 7934
rect 39953 7579 39999 7922
rect 40113 7911 40159 7922
rect 40241 7579 40287 7922
rect 40401 8496 40447 8716
rect 40401 7579 40447 7922
rect 40746 11985 40901 12019
rect 40947 12019 42325 12031
rect 40947 11985 41066 12019
rect 40746 11937 41066 11985
rect 40746 11891 40901 11937
rect 40947 11891 41066 11937
rect 40746 11843 41066 11891
rect 40746 11797 40901 11843
rect 40947 11797 41066 11843
rect 40746 11749 41066 11797
rect 40746 11703 40901 11749
rect 40947 11703 41066 11749
rect 40746 11655 41066 11703
rect 40746 11609 40901 11655
rect 40947 11609 41066 11655
rect 40746 11561 41066 11609
rect 40746 11515 40901 11561
rect 40947 11515 41066 11561
rect 40746 11467 41066 11515
rect 40746 11421 40901 11467
rect 40947 11421 41066 11467
rect 40746 11373 41066 11421
rect 40746 11327 40901 11373
rect 40947 11327 41066 11373
rect 40746 11279 41066 11327
rect 40746 11233 40901 11279
rect 40947 11233 41066 11279
rect 40746 11185 41066 11233
rect 40746 11139 40901 11185
rect 40947 11139 41066 11185
rect 40746 11091 41066 11139
rect 40746 11045 40901 11091
rect 40947 11045 41066 11091
rect 40746 10997 41066 11045
rect 40746 10951 40901 10997
rect 40947 10951 41066 10997
rect 40746 10903 41066 10951
rect 40746 10857 40901 10903
rect 40947 10857 41066 10903
rect 40746 10809 41066 10857
rect 40746 10763 40901 10809
rect 40947 10763 41066 10809
rect 40746 10715 41066 10763
rect 40746 10669 40901 10715
rect 40947 10669 41066 10715
rect 40746 10621 41066 10669
rect 40746 10575 40901 10621
rect 40947 10575 41066 10621
rect 40746 10527 41066 10575
rect 40746 10481 40901 10527
rect 40947 10481 41066 10527
rect 40746 10433 41066 10481
rect 40746 10387 40901 10433
rect 40947 10387 41066 10433
rect 40746 10339 41066 10387
rect 40746 10293 40901 10339
rect 40947 10293 41066 10339
rect 40746 10245 41066 10293
rect 40746 10199 40901 10245
rect 40947 10199 41066 10245
rect 40746 10151 41066 10199
rect 40746 10105 40901 10151
rect 40947 10105 41066 10151
rect 40746 10057 41066 10105
rect 40746 10011 40901 10057
rect 40947 10011 41066 10057
rect 40746 9963 41066 10011
rect 40746 9917 40901 9963
rect 40947 9917 41066 9963
rect 40746 9869 41066 9917
rect 40746 9823 40901 9869
rect 40947 9823 41066 9869
rect 40746 9775 41066 9823
rect 40746 9729 40901 9775
rect 40947 9729 41066 9775
rect 40746 9681 41066 9729
rect 40746 9635 40901 9681
rect 40947 9635 41066 9681
rect 40746 9587 41066 9635
rect 40746 9541 40901 9587
rect 40947 9541 41066 9587
rect 40746 9493 41066 9541
rect 40746 9447 40901 9493
rect 40947 9447 41066 9493
rect 40746 9399 41066 9447
rect 40746 9353 40901 9399
rect 40947 9353 41066 9399
rect 40746 9305 41066 9353
rect 40746 9259 40901 9305
rect 40947 9259 41066 9305
rect 40746 9211 41066 9259
rect 40746 9165 40901 9211
rect 40947 9165 41066 9211
rect 40746 9117 41066 9165
rect 40746 9071 40901 9117
rect 40947 9071 41066 9117
rect 40746 9023 41066 9071
rect 40746 8977 40901 9023
rect 40947 8977 41066 9023
rect 40746 8929 41066 8977
rect 40746 8883 40901 8929
rect 40947 8883 41066 8929
rect 40746 8835 41066 8883
rect 40746 8789 40901 8835
rect 40947 8789 41066 8835
rect 40746 8741 41066 8789
rect 40746 8695 40901 8741
rect 40947 8695 41066 8741
rect 40746 8647 41066 8695
rect 40746 8601 40901 8647
rect 40947 8601 41066 8647
rect 40746 8553 41066 8601
rect 40746 8507 40901 8553
rect 40947 8507 41066 8553
rect 40746 8459 41066 8507
rect 40746 8413 40901 8459
rect 40947 8413 41066 8459
rect 40746 8365 41066 8413
rect 40746 8319 40901 8365
rect 40947 8319 41066 8365
rect 40746 8271 41066 8319
rect 40746 8225 40901 8271
rect 40947 8225 41066 8271
rect 40746 8177 41066 8225
rect 40746 8131 40901 8177
rect 40947 8131 41066 8177
rect 40746 8083 41066 8131
rect 40746 8037 40901 8083
rect 40947 8037 41066 8083
rect 40746 7989 41066 8037
rect 40746 7943 40901 7989
rect 40947 7943 41066 7989
rect 40746 7895 41066 7943
rect 40746 7849 40901 7895
rect 40947 7849 41066 7895
rect 40746 7801 41066 7849
rect 40746 7755 40901 7801
rect 40947 7755 41066 7801
rect 40746 7707 41066 7755
rect 40746 7661 40901 7707
rect 40947 7661 41066 7707
rect 40746 7613 41066 7661
rect 40746 7579 40901 7613
rect 36811 7567 40901 7579
rect 40947 7579 41066 7613
rect 42206 11985 42325 12019
rect 42371 12019 46461 12031
rect 42371 11985 42526 12019
rect 42206 11937 42526 11985
rect 42206 11891 42325 11937
rect 42371 11891 42526 11937
rect 42206 11843 42526 11891
rect 42206 11797 42325 11843
rect 42371 11797 42526 11843
rect 42206 11749 42526 11797
rect 42206 11703 42325 11749
rect 42371 11703 42526 11749
rect 42206 11655 42526 11703
rect 42206 11609 42325 11655
rect 42371 11609 42526 11655
rect 42206 11561 42526 11609
rect 42206 11515 42325 11561
rect 42371 11515 42526 11561
rect 42206 11467 42526 11515
rect 42206 11421 42325 11467
rect 42371 11421 42526 11467
rect 42206 11373 42526 11421
rect 42206 11327 42325 11373
rect 42371 11327 42526 11373
rect 42206 11279 42526 11327
rect 42206 11233 42325 11279
rect 42371 11233 42526 11279
rect 42206 11185 42526 11233
rect 42206 11139 42325 11185
rect 42371 11139 42526 11185
rect 42206 11091 42526 11139
rect 42206 11045 42325 11091
rect 42371 11045 42526 11091
rect 42206 10997 42526 11045
rect 42206 10951 42325 10997
rect 42371 10951 42526 10997
rect 42206 10903 42526 10951
rect 42206 10857 42325 10903
rect 42371 10857 42526 10903
rect 42206 10809 42526 10857
rect 42206 10763 42325 10809
rect 42371 10763 42526 10809
rect 42206 10715 42526 10763
rect 42206 10669 42325 10715
rect 42371 10669 42526 10715
rect 42206 10621 42526 10669
rect 42206 10575 42325 10621
rect 42371 10575 42526 10621
rect 42206 10527 42526 10575
rect 42206 10481 42325 10527
rect 42371 10481 42526 10527
rect 42206 10433 42526 10481
rect 42206 10387 42325 10433
rect 42371 10387 42526 10433
rect 42206 10339 42526 10387
rect 42206 10293 42325 10339
rect 42371 10293 42526 10339
rect 42206 10245 42526 10293
rect 42206 10199 42325 10245
rect 42371 10199 42526 10245
rect 42206 10151 42526 10199
rect 42206 10105 42325 10151
rect 42371 10105 42526 10151
rect 42206 10057 42526 10105
rect 42206 10011 42325 10057
rect 42371 10011 42526 10057
rect 42206 9963 42526 10011
rect 42206 9917 42325 9963
rect 42371 9917 42526 9963
rect 42206 9869 42526 9917
rect 42206 9823 42325 9869
rect 42371 9823 42526 9869
rect 42206 9775 42526 9823
rect 42206 9729 42325 9775
rect 42371 9729 42526 9775
rect 42206 9681 42526 9729
rect 42206 9635 42325 9681
rect 42371 9635 42526 9681
rect 42206 9587 42526 9635
rect 42206 9541 42325 9587
rect 42371 9541 42526 9587
rect 42206 9493 42526 9541
rect 42206 9447 42325 9493
rect 42371 9447 42526 9493
rect 42206 9399 42526 9447
rect 42206 9353 42325 9399
rect 42371 9353 42526 9399
rect 42206 9305 42526 9353
rect 42206 9259 42325 9305
rect 42371 9259 42526 9305
rect 42206 9211 42526 9259
rect 42206 9165 42325 9211
rect 42371 9165 42526 9211
rect 42206 9117 42526 9165
rect 42206 9071 42325 9117
rect 42371 9071 42526 9117
rect 42206 9023 42526 9071
rect 42206 8977 42325 9023
rect 42371 8977 42526 9023
rect 42206 8929 42526 8977
rect 42206 8883 42325 8929
rect 42371 8883 42526 8929
rect 42206 8835 42526 8883
rect 42206 8789 42325 8835
rect 42371 8789 42526 8835
rect 42206 8741 42526 8789
rect 42206 8695 42325 8741
rect 42371 8695 42526 8741
rect 42206 8647 42526 8695
rect 42206 8601 42325 8647
rect 42371 8601 42526 8647
rect 42206 8553 42526 8601
rect 42206 8507 42325 8553
rect 42371 8507 42526 8553
rect 42206 8459 42526 8507
rect 42206 8413 42325 8459
rect 42371 8413 42526 8459
rect 42206 8365 42526 8413
rect 42206 8319 42325 8365
rect 42371 8319 42526 8365
rect 42206 8271 42526 8319
rect 42206 8225 42325 8271
rect 42371 8225 42526 8271
rect 42206 8177 42526 8225
rect 42206 8131 42325 8177
rect 42371 8131 42526 8177
rect 42206 8083 42526 8131
rect 42206 8037 42325 8083
rect 42371 8037 42526 8083
rect 42206 7989 42526 8037
rect 42206 7943 42325 7989
rect 42371 7943 42526 7989
rect 42206 7895 42526 7943
rect 42206 7849 42325 7895
rect 42371 7849 42526 7895
rect 42206 7801 42526 7849
rect 42206 7755 42325 7801
rect 42371 7755 42526 7801
rect 42206 7707 42526 7755
rect 42206 7661 42325 7707
rect 42371 7661 42526 7707
rect 42206 7613 42526 7661
rect 42206 7579 42325 7613
rect 40947 7567 42325 7579
rect 42371 7579 42526 7613
rect 42825 11676 42871 12019
rect 42825 10882 42871 11102
rect 42985 11676 43031 12019
rect 43113 11676 43159 11687
rect 43098 11270 43113 11282
rect 43273 11676 43319 12019
rect 43433 11676 43479 11687
rect 43593 11676 43639 12019
rect 43159 11270 43174 11282
rect 43098 11218 43110 11270
rect 43162 11218 43174 11270
rect 43098 11166 43113 11218
rect 43159 11166 43174 11218
rect 43098 11114 43110 11166
rect 43162 11114 43174 11166
rect 43098 11102 43113 11114
rect 43159 11102 43174 11114
rect 43419 11664 43433 11676
rect 43479 11664 43495 11676
rect 43419 11612 43431 11664
rect 43483 11612 43495 11664
rect 43419 11560 43433 11612
rect 43479 11560 43495 11612
rect 43419 11508 43431 11560
rect 43483 11508 43495 11560
rect 43419 11496 43433 11508
rect 42985 10882 43031 11102
rect 43113 11091 43159 11102
rect 42825 10836 42905 10882
rect 42951 10836 43031 10882
rect 42825 10616 42871 10836
rect 42825 9556 42871 10042
rect 42825 8762 42871 8982
rect 42985 10616 43031 10836
rect 43113 10616 43159 10627
rect 43098 10210 43113 10222
rect 43273 10616 43319 11102
rect 43479 11496 43495 11508
rect 43433 11091 43479 11102
rect 43753 11676 43799 11687
rect 43738 11270 43753 11282
rect 43913 11676 43959 12019
rect 44298 11812 44374 11824
rect 44298 11760 44310 11812
rect 44362 11809 44374 11812
rect 44458 11812 44534 11824
rect 44458 11809 44470 11812
rect 44362 11760 44470 11809
rect 44522 11760 44534 11812
rect 44298 11748 44534 11760
rect 44073 11676 44119 11687
rect 44233 11676 44279 11687
rect 43799 11270 43814 11282
rect 43738 11218 43750 11270
rect 43802 11218 43814 11270
rect 43738 11166 43753 11218
rect 43799 11166 43814 11218
rect 43738 11114 43750 11166
rect 43802 11114 43814 11166
rect 43738 11102 43753 11114
rect 43799 11102 43814 11114
rect 44059 11664 44073 11676
rect 44119 11664 44135 11676
rect 44059 11612 44071 11664
rect 44123 11612 44135 11664
rect 44059 11560 44073 11612
rect 44119 11560 44135 11612
rect 44059 11508 44071 11560
rect 44123 11508 44135 11560
rect 44059 11496 44073 11508
rect 43433 10616 43479 10627
rect 43593 10616 43639 11102
rect 43753 11091 43799 11102
rect 43913 11045 43959 11102
rect 44119 11496 44135 11508
rect 44073 11091 44119 11102
rect 44233 11045 44279 11102
rect 44393 11676 44439 11748
rect 44393 11091 44439 11102
rect 44553 11676 44599 11687
rect 44713 11676 44759 11687
rect 44873 11676 44919 12019
rect 44699 11664 44713 11676
rect 44759 11664 44775 11676
rect 44699 11612 44711 11664
rect 44763 11612 44775 11664
rect 44699 11560 44713 11612
rect 44759 11560 44775 11612
rect 44699 11508 44711 11560
rect 44763 11508 44775 11560
rect 44699 11496 44713 11508
rect 44553 11045 44599 11102
rect 44759 11496 44775 11508
rect 44713 11091 44759 11102
rect 45033 11676 45079 11687
rect 45018 11270 45033 11282
rect 45193 11676 45239 12019
rect 45353 11676 45399 11687
rect 45513 11676 45559 12019
rect 45079 11270 45094 11282
rect 45018 11218 45030 11270
rect 45082 11218 45094 11270
rect 45018 11166 45033 11218
rect 45079 11166 45094 11218
rect 45018 11114 45030 11166
rect 45082 11114 45094 11166
rect 45018 11102 45033 11114
rect 45079 11102 45094 11114
rect 45339 11664 45353 11676
rect 45399 11664 45415 11676
rect 45339 11612 45351 11664
rect 45403 11612 45415 11664
rect 45339 11560 45353 11612
rect 45399 11560 45415 11612
rect 45339 11508 45351 11560
rect 45403 11508 45415 11560
rect 45339 11496 45353 11508
rect 43913 10999 44599 11045
rect 43159 10210 43174 10222
rect 43098 10158 43110 10210
rect 43162 10158 43174 10210
rect 43098 10106 43113 10158
rect 43159 10106 43174 10158
rect 43098 10054 43110 10106
rect 43162 10054 43174 10106
rect 43098 10042 43113 10054
rect 43159 10042 43174 10054
rect 43419 10604 43433 10616
rect 43479 10604 43495 10616
rect 43419 10552 43431 10604
rect 43483 10552 43495 10604
rect 43419 10500 43433 10552
rect 43479 10500 43495 10552
rect 43419 10448 43431 10500
rect 43483 10448 43495 10500
rect 43419 10436 43433 10448
rect 42985 9556 43031 10042
rect 43113 10031 43159 10042
rect 43113 9556 43159 9567
rect 43098 9150 43113 9162
rect 43273 9556 43319 10042
rect 43479 10436 43495 10448
rect 43433 10031 43479 10042
rect 43753 10616 43799 10627
rect 43738 10210 43753 10222
rect 43913 10616 43959 10999
rect 44298 10752 44374 10764
rect 44298 10700 44310 10752
rect 44362 10749 44374 10752
rect 44458 10752 44534 10764
rect 44458 10749 44470 10752
rect 44362 10700 44470 10749
rect 44522 10700 44534 10752
rect 44298 10688 44534 10700
rect 44073 10616 44119 10627
rect 44233 10616 44279 10627
rect 43799 10210 43814 10222
rect 43738 10158 43750 10210
rect 43802 10158 43814 10210
rect 43738 10106 43753 10158
rect 43799 10106 43814 10158
rect 43738 10054 43750 10106
rect 43802 10054 43814 10106
rect 43738 10042 43753 10054
rect 43799 10042 43814 10054
rect 44059 10604 44073 10616
rect 44119 10604 44135 10616
rect 44059 10552 44071 10604
rect 44123 10552 44135 10604
rect 44059 10500 44073 10552
rect 44119 10500 44135 10552
rect 44059 10448 44071 10500
rect 44123 10448 44135 10500
rect 44059 10436 44073 10448
rect 43433 9556 43479 9567
rect 43593 9556 43639 10042
rect 43753 10031 43799 10042
rect 43913 9985 43959 10042
rect 44119 10436 44135 10448
rect 44073 10031 44119 10042
rect 44233 9985 44279 10042
rect 44393 10616 44439 10688
rect 44393 10031 44439 10042
rect 44553 10616 44599 10627
rect 44713 10616 44759 10627
rect 44873 10616 44919 11102
rect 45033 11091 45079 11102
rect 44699 10604 44713 10616
rect 44759 10604 44775 10616
rect 44699 10552 44711 10604
rect 44763 10552 44775 10604
rect 44699 10500 44713 10552
rect 44759 10500 44775 10552
rect 44699 10448 44711 10500
rect 44763 10448 44775 10500
rect 44699 10436 44713 10448
rect 44553 9985 44599 10042
rect 44759 10436 44775 10448
rect 44713 10031 44759 10042
rect 45033 10616 45079 10627
rect 45018 10210 45033 10222
rect 45193 10616 45239 11102
rect 45399 11496 45415 11508
rect 45353 11091 45399 11102
rect 45673 11676 45719 11687
rect 45658 11270 45673 11282
rect 45801 11676 45847 12019
rect 45719 11270 45734 11282
rect 45658 11218 45670 11270
rect 45722 11218 45734 11270
rect 45658 11166 45673 11218
rect 45719 11166 45734 11218
rect 45658 11114 45670 11166
rect 45722 11114 45734 11166
rect 45658 11102 45673 11114
rect 45719 11102 45734 11114
rect 45353 10616 45399 10627
rect 45513 10616 45559 11102
rect 45673 11091 45719 11102
rect 45801 10882 45847 11102
rect 45961 11676 46007 12019
rect 45961 10882 46007 11102
rect 45801 10836 45881 10882
rect 45927 10836 46007 10882
rect 45079 10210 45094 10222
rect 45018 10158 45030 10210
rect 45082 10158 45094 10210
rect 45018 10106 45033 10158
rect 45079 10106 45094 10158
rect 45018 10054 45030 10106
rect 45082 10054 45094 10106
rect 45018 10042 45033 10054
rect 45079 10042 45094 10054
rect 45339 10604 45353 10616
rect 45399 10604 45415 10616
rect 45339 10552 45351 10604
rect 45403 10552 45415 10604
rect 45339 10500 45353 10552
rect 45399 10500 45415 10552
rect 45339 10448 45351 10500
rect 45403 10448 45415 10500
rect 45339 10436 45353 10448
rect 43913 9939 44599 9985
rect 43159 9150 43174 9162
rect 43098 9098 43110 9150
rect 43162 9098 43174 9150
rect 43098 9046 43113 9098
rect 43159 9046 43174 9098
rect 43098 8994 43110 9046
rect 43162 8994 43174 9046
rect 43098 8982 43113 8994
rect 43159 8982 43174 8994
rect 43419 9544 43433 9556
rect 43479 9544 43495 9556
rect 43419 9492 43431 9544
rect 43483 9492 43495 9544
rect 43419 9440 43433 9492
rect 43479 9440 43495 9492
rect 43419 9388 43431 9440
rect 43483 9388 43495 9440
rect 43419 9376 43433 9388
rect 42985 8762 43031 8982
rect 43113 8971 43159 8982
rect 42825 8716 42905 8762
rect 42951 8716 43031 8762
rect 42825 8496 42871 8716
rect 42825 7579 42871 7922
rect 42985 8496 43031 8716
rect 43113 8496 43159 8507
rect 43098 8090 43113 8102
rect 43273 8496 43319 8982
rect 43479 9376 43495 9388
rect 43433 8971 43479 8982
rect 43753 9556 43799 9567
rect 43738 9150 43753 9162
rect 43913 9556 43959 9939
rect 44298 9692 44374 9704
rect 44298 9640 44310 9692
rect 44362 9689 44374 9692
rect 44458 9692 44534 9704
rect 44458 9689 44470 9692
rect 44362 9640 44470 9689
rect 44522 9640 44534 9692
rect 44298 9628 44534 9640
rect 44073 9556 44119 9567
rect 44233 9556 44279 9567
rect 43799 9150 43814 9162
rect 43738 9098 43750 9150
rect 43802 9098 43814 9150
rect 43738 9046 43753 9098
rect 43799 9046 43814 9098
rect 43738 8994 43750 9046
rect 43802 8994 43814 9046
rect 43738 8982 43753 8994
rect 43799 8982 43814 8994
rect 44059 9544 44073 9556
rect 44119 9544 44135 9556
rect 44059 9492 44071 9544
rect 44123 9492 44135 9544
rect 44059 9440 44073 9492
rect 44119 9440 44135 9492
rect 44059 9388 44071 9440
rect 44123 9388 44135 9440
rect 44059 9376 44073 9388
rect 43433 8496 43479 8507
rect 43593 8496 43639 8982
rect 43753 8971 43799 8982
rect 43913 8925 43959 8982
rect 44119 9376 44135 9388
rect 44073 8971 44119 8982
rect 44233 8925 44279 8982
rect 44393 9556 44439 9628
rect 44393 8971 44439 8982
rect 44553 9556 44599 9567
rect 44713 9556 44759 9567
rect 44873 9556 44919 10042
rect 45033 10031 45079 10042
rect 44699 9544 44713 9556
rect 44759 9544 44775 9556
rect 44699 9492 44711 9544
rect 44763 9492 44775 9544
rect 44699 9440 44713 9492
rect 44759 9440 44775 9492
rect 44699 9388 44711 9440
rect 44763 9388 44775 9440
rect 44699 9376 44713 9388
rect 44553 8925 44599 8982
rect 44759 9376 44775 9388
rect 44713 8971 44759 8982
rect 45033 9556 45079 9567
rect 45018 9150 45033 9162
rect 45193 9556 45239 10042
rect 45399 10436 45415 10448
rect 45353 10031 45399 10042
rect 45673 10616 45719 10627
rect 45658 10210 45673 10222
rect 45801 10616 45847 10836
rect 45719 10210 45734 10222
rect 45658 10158 45670 10210
rect 45722 10158 45734 10210
rect 45658 10106 45673 10158
rect 45719 10106 45734 10158
rect 45658 10054 45670 10106
rect 45722 10054 45734 10106
rect 45658 10042 45673 10054
rect 45719 10042 45734 10054
rect 45353 9556 45399 9567
rect 45513 9556 45559 10042
rect 45673 10031 45719 10042
rect 45079 9150 45094 9162
rect 45018 9098 45030 9150
rect 45082 9098 45094 9150
rect 45018 9046 45033 9098
rect 45079 9046 45094 9098
rect 45018 8994 45030 9046
rect 45082 8994 45094 9046
rect 45018 8982 45033 8994
rect 45079 8982 45094 8994
rect 45339 9544 45353 9556
rect 45399 9544 45415 9556
rect 45339 9492 45351 9544
rect 45403 9492 45415 9544
rect 45339 9440 45353 9492
rect 45399 9440 45415 9492
rect 45339 9388 45351 9440
rect 45403 9388 45415 9440
rect 45339 9376 45353 9388
rect 43913 8879 44599 8925
rect 43159 8090 43174 8102
rect 43098 8038 43110 8090
rect 43162 8038 43174 8090
rect 43098 7986 43113 8038
rect 43159 7986 43174 8038
rect 43098 7934 43110 7986
rect 43162 7934 43174 7986
rect 43098 7922 43113 7934
rect 43159 7922 43174 7934
rect 43419 8484 43433 8496
rect 43479 8484 43495 8496
rect 43419 8432 43431 8484
rect 43483 8432 43495 8484
rect 43419 8380 43433 8432
rect 43479 8380 43495 8432
rect 43419 8328 43431 8380
rect 43483 8328 43495 8380
rect 43419 8316 43433 8328
rect 42985 7579 43031 7922
rect 43113 7911 43159 7922
rect 43273 7579 43319 7922
rect 43479 8316 43495 8328
rect 43433 7911 43479 7922
rect 43753 8496 43799 8507
rect 43738 8090 43753 8102
rect 43913 8496 43959 8879
rect 44298 8632 44374 8644
rect 44298 8580 44310 8632
rect 44362 8629 44374 8632
rect 44458 8632 44534 8644
rect 44458 8629 44470 8632
rect 44362 8580 44470 8629
rect 44522 8580 44534 8632
rect 44298 8568 44534 8580
rect 44073 8496 44119 8507
rect 44233 8496 44279 8507
rect 43799 8090 43814 8102
rect 43738 8038 43750 8090
rect 43802 8038 43814 8090
rect 43738 7986 43753 8038
rect 43799 7986 43814 8038
rect 43738 7934 43750 7986
rect 43802 7934 43814 7986
rect 43738 7922 43753 7934
rect 43799 7922 43814 7934
rect 44059 8484 44073 8496
rect 44119 8484 44135 8496
rect 44059 8432 44071 8484
rect 44123 8432 44135 8484
rect 44059 8380 44073 8432
rect 44119 8380 44135 8432
rect 44059 8328 44071 8380
rect 44123 8328 44135 8380
rect 44059 8316 44073 8328
rect 43593 7579 43639 7922
rect 43753 7911 43799 7922
rect 43913 7579 43959 7922
rect 44119 8316 44135 8328
rect 44073 7911 44119 7922
rect 44233 7579 44279 7922
rect 44393 8496 44439 8568
rect 44393 7911 44439 7922
rect 44553 8496 44599 8507
rect 44713 8496 44759 8507
rect 44873 8496 44919 8982
rect 45033 8971 45079 8982
rect 44699 8484 44713 8496
rect 44759 8484 44775 8496
rect 44699 8432 44711 8484
rect 44763 8432 44775 8484
rect 44699 8380 44713 8432
rect 44759 8380 44775 8432
rect 44699 8328 44711 8380
rect 44763 8328 44775 8380
rect 44699 8316 44713 8328
rect 44553 7579 44599 7922
rect 44759 8316 44775 8328
rect 44713 7911 44759 7922
rect 45033 8496 45079 8507
rect 45018 8090 45033 8102
rect 45193 8496 45239 8982
rect 45399 9376 45415 9388
rect 45353 8971 45399 8982
rect 45673 9556 45719 9567
rect 45658 9150 45673 9162
rect 45801 9556 45847 10042
rect 45719 9150 45734 9162
rect 45658 9098 45670 9150
rect 45722 9098 45734 9150
rect 45658 9046 45673 9098
rect 45719 9046 45734 9098
rect 45658 8994 45670 9046
rect 45722 8994 45734 9046
rect 45658 8982 45673 8994
rect 45719 8982 45734 8994
rect 45353 8496 45399 8507
rect 45513 8496 45559 8982
rect 45673 8971 45719 8982
rect 45801 8762 45847 8982
rect 45961 10616 46007 10836
rect 45961 9556 46007 10042
rect 45961 8762 46007 8982
rect 45801 8716 45881 8762
rect 45927 8716 46007 8762
rect 45079 8090 45094 8102
rect 45018 8038 45030 8090
rect 45082 8038 45094 8090
rect 45018 7986 45033 8038
rect 45079 7986 45094 8038
rect 45018 7934 45030 7986
rect 45082 7934 45094 7986
rect 45018 7922 45033 7934
rect 45079 7922 45094 7934
rect 45339 8484 45353 8496
rect 45399 8484 45415 8496
rect 45339 8432 45351 8484
rect 45403 8432 45415 8484
rect 45339 8380 45353 8432
rect 45399 8380 45415 8432
rect 45339 8328 45351 8380
rect 45403 8328 45415 8380
rect 45339 8316 45353 8328
rect 44873 7579 44919 7922
rect 45033 7911 45079 7922
rect 45193 7579 45239 7922
rect 45399 8316 45415 8328
rect 45353 7911 45399 7922
rect 45673 8496 45719 8507
rect 45658 8090 45673 8102
rect 45801 8496 45847 8716
rect 45719 8090 45734 8102
rect 45658 8038 45670 8090
rect 45722 8038 45734 8090
rect 45658 7986 45673 8038
rect 45719 7986 45734 8038
rect 45658 7934 45670 7986
rect 45722 7934 45734 7986
rect 45658 7922 45673 7934
rect 45719 7922 45734 7934
rect 45513 7579 45559 7922
rect 45673 7911 45719 7922
rect 45801 7579 45847 7922
rect 45961 8496 46007 8716
rect 45961 7579 46007 7922
rect 46306 11985 46461 12019
rect 46507 12019 50597 12031
rect 46507 11985 46662 12019
rect 46306 11937 46662 11985
rect 46306 11891 46461 11937
rect 46507 11891 46662 11937
rect 46306 11843 46662 11891
rect 46306 11797 46461 11843
rect 46507 11797 46662 11843
rect 46306 11749 46662 11797
rect 46306 11703 46461 11749
rect 46507 11703 46662 11749
rect 46306 11655 46662 11703
rect 46306 11609 46461 11655
rect 46507 11609 46662 11655
rect 46306 11561 46662 11609
rect 46306 11515 46461 11561
rect 46507 11515 46662 11561
rect 46306 11467 46662 11515
rect 46306 11421 46461 11467
rect 46507 11421 46662 11467
rect 46306 11373 46662 11421
rect 46306 11327 46461 11373
rect 46507 11327 46662 11373
rect 46306 11279 46662 11327
rect 46306 11233 46461 11279
rect 46507 11233 46662 11279
rect 46306 11185 46662 11233
rect 46306 11139 46461 11185
rect 46507 11139 46662 11185
rect 46306 11091 46662 11139
rect 46306 11045 46461 11091
rect 46507 11045 46662 11091
rect 46306 10997 46662 11045
rect 46306 10951 46461 10997
rect 46507 10951 46662 10997
rect 46306 10903 46662 10951
rect 46306 10857 46461 10903
rect 46507 10857 46662 10903
rect 46306 10809 46662 10857
rect 46306 10763 46461 10809
rect 46507 10763 46662 10809
rect 46306 10715 46662 10763
rect 46306 10669 46461 10715
rect 46507 10669 46662 10715
rect 46306 10621 46662 10669
rect 46306 10575 46461 10621
rect 46507 10575 46662 10621
rect 46306 10527 46662 10575
rect 46306 10481 46461 10527
rect 46507 10481 46662 10527
rect 46306 10433 46662 10481
rect 46306 10387 46461 10433
rect 46507 10387 46662 10433
rect 46306 10339 46662 10387
rect 46306 10293 46461 10339
rect 46507 10293 46662 10339
rect 46306 10245 46662 10293
rect 46306 10199 46461 10245
rect 46507 10199 46662 10245
rect 46306 10151 46662 10199
rect 46306 10105 46461 10151
rect 46507 10105 46662 10151
rect 46306 10057 46662 10105
rect 46306 10011 46461 10057
rect 46507 10011 46662 10057
rect 46306 9963 46662 10011
rect 46306 9917 46461 9963
rect 46507 9917 46662 9963
rect 46306 9869 46662 9917
rect 46306 9823 46461 9869
rect 46507 9823 46662 9869
rect 46306 9775 46662 9823
rect 46306 9729 46461 9775
rect 46507 9729 46662 9775
rect 46306 9681 46662 9729
rect 46306 9635 46461 9681
rect 46507 9635 46662 9681
rect 46306 9587 46662 9635
rect 46306 9541 46461 9587
rect 46507 9541 46662 9587
rect 46306 9493 46662 9541
rect 46306 9447 46461 9493
rect 46507 9447 46662 9493
rect 46306 9399 46662 9447
rect 46306 9353 46461 9399
rect 46507 9353 46662 9399
rect 46306 9305 46662 9353
rect 46306 9259 46461 9305
rect 46507 9259 46662 9305
rect 46306 9211 46662 9259
rect 46306 9165 46461 9211
rect 46507 9165 46662 9211
rect 46306 9117 46662 9165
rect 46306 9071 46461 9117
rect 46507 9071 46662 9117
rect 46306 9023 46662 9071
rect 46306 8977 46461 9023
rect 46507 8977 46662 9023
rect 46306 8929 46662 8977
rect 46306 8883 46461 8929
rect 46507 8883 46662 8929
rect 46306 8835 46662 8883
rect 46306 8789 46461 8835
rect 46507 8789 46662 8835
rect 46306 8741 46662 8789
rect 46306 8695 46461 8741
rect 46507 8695 46662 8741
rect 46306 8647 46662 8695
rect 46306 8601 46461 8647
rect 46507 8601 46662 8647
rect 46306 8553 46662 8601
rect 46306 8507 46461 8553
rect 46507 8507 46662 8553
rect 46306 8459 46662 8507
rect 46306 8413 46461 8459
rect 46507 8413 46662 8459
rect 46306 8365 46662 8413
rect 46306 8319 46461 8365
rect 46507 8319 46662 8365
rect 46306 8271 46662 8319
rect 46306 8225 46461 8271
rect 46507 8225 46662 8271
rect 46306 8177 46662 8225
rect 46306 8131 46461 8177
rect 46507 8131 46662 8177
rect 46306 8083 46662 8131
rect 46306 8037 46461 8083
rect 46507 8037 46662 8083
rect 46306 7989 46662 8037
rect 46306 7943 46461 7989
rect 46507 7943 46662 7989
rect 46306 7895 46662 7943
rect 46306 7849 46461 7895
rect 46507 7849 46662 7895
rect 46306 7801 46662 7849
rect 46306 7755 46461 7801
rect 46507 7755 46662 7801
rect 46306 7707 46662 7755
rect 46306 7661 46461 7707
rect 46507 7661 46662 7707
rect 46306 7613 46662 7661
rect 46306 7579 46461 7613
rect 42371 7567 46461 7579
rect 46507 7579 46662 7613
rect 46961 11676 47007 12019
rect 46961 10882 47007 11102
rect 47121 11676 47167 12019
rect 47249 11676 47295 11687
rect 47234 11270 47249 11282
rect 47409 11676 47455 12019
rect 47569 11676 47615 11687
rect 47729 11676 47775 12019
rect 47295 11270 47310 11282
rect 47234 11218 47246 11270
rect 47298 11218 47310 11270
rect 47234 11166 47249 11218
rect 47295 11166 47310 11218
rect 47234 11114 47246 11166
rect 47298 11114 47310 11166
rect 47234 11102 47249 11114
rect 47295 11102 47310 11114
rect 47553 11664 47569 11676
rect 47615 11664 47629 11676
rect 47553 11612 47565 11664
rect 47617 11612 47629 11664
rect 47553 11560 47569 11612
rect 47615 11560 47629 11612
rect 47553 11508 47565 11560
rect 47617 11508 47629 11560
rect 47553 11496 47569 11508
rect 47121 10882 47167 11102
rect 47249 11091 47295 11102
rect 46961 10836 47041 10882
rect 47087 10836 47167 10882
rect 46961 10616 47007 10836
rect 46961 9556 47007 10042
rect 46961 8762 47007 8982
rect 47121 10616 47167 10836
rect 47249 10616 47295 10627
rect 47234 10210 47249 10222
rect 47409 10616 47455 11102
rect 47615 11496 47629 11508
rect 47569 11091 47615 11102
rect 47889 11676 47935 11687
rect 47874 11270 47889 11282
rect 48049 11676 48095 12019
rect 48434 11812 48510 11824
rect 48434 11760 48446 11812
rect 48498 11809 48510 11812
rect 48594 11812 48670 11824
rect 48594 11809 48606 11812
rect 48498 11760 48606 11809
rect 48658 11760 48670 11812
rect 48434 11748 48670 11760
rect 48209 11676 48255 11687
rect 48369 11676 48415 11687
rect 47935 11270 47950 11282
rect 47874 11218 47886 11270
rect 47938 11218 47950 11270
rect 47874 11166 47889 11218
rect 47935 11166 47950 11218
rect 47874 11114 47886 11166
rect 47938 11114 47950 11166
rect 47874 11102 47889 11114
rect 47935 11102 47950 11114
rect 48193 11664 48209 11676
rect 48255 11664 48269 11676
rect 48193 11612 48205 11664
rect 48257 11612 48269 11664
rect 48193 11560 48209 11612
rect 48255 11560 48269 11612
rect 48193 11508 48205 11560
rect 48257 11508 48269 11560
rect 48193 11496 48209 11508
rect 47569 10616 47615 10627
rect 47729 10616 47775 11102
rect 47889 11091 47935 11102
rect 47295 10210 47310 10222
rect 47234 10158 47246 10210
rect 47298 10158 47310 10210
rect 47234 10106 47249 10158
rect 47295 10106 47310 10158
rect 47234 10054 47246 10106
rect 47298 10054 47310 10106
rect 47234 10042 47249 10054
rect 47295 10042 47310 10054
rect 47553 10604 47569 10616
rect 47615 10604 47629 10616
rect 47553 10552 47565 10604
rect 47617 10552 47629 10604
rect 47553 10500 47569 10552
rect 47615 10500 47629 10552
rect 47553 10448 47565 10500
rect 47617 10448 47629 10500
rect 47553 10436 47569 10448
rect 47121 9556 47167 10042
rect 47249 10031 47295 10042
rect 47249 9556 47295 9567
rect 47234 9150 47249 9162
rect 47409 9556 47455 10042
rect 47615 10436 47629 10448
rect 47569 10031 47615 10042
rect 47889 10616 47935 10627
rect 47874 10210 47889 10222
rect 48049 10616 48095 11102
rect 48255 11496 48269 11508
rect 48209 11091 48255 11102
rect 48369 11045 48415 11102
rect 48529 11676 48575 11748
rect 48529 11091 48575 11102
rect 48689 11676 48735 11687
rect 48849 11676 48895 11687
rect 49009 11676 49055 12019
rect 48833 11664 48849 11676
rect 48895 11664 48909 11676
rect 48833 11612 48845 11664
rect 48897 11612 48909 11664
rect 48833 11560 48849 11612
rect 48895 11560 48909 11612
rect 48833 11508 48845 11560
rect 48897 11508 48909 11560
rect 48833 11496 48849 11508
rect 48689 11045 48735 11102
rect 48895 11496 48909 11508
rect 48849 11091 48895 11102
rect 49169 11676 49215 11687
rect 49154 11270 49169 11282
rect 49329 11676 49375 12019
rect 49489 11676 49535 11687
rect 49649 11676 49695 12019
rect 49215 11270 49230 11282
rect 49154 11218 49166 11270
rect 49218 11218 49230 11270
rect 49154 11166 49169 11218
rect 49215 11166 49230 11218
rect 49154 11114 49166 11166
rect 49218 11114 49230 11166
rect 49154 11102 49169 11114
rect 49215 11102 49230 11114
rect 49473 11664 49489 11676
rect 49535 11664 49549 11676
rect 49473 11612 49485 11664
rect 49537 11612 49549 11664
rect 49473 11560 49489 11612
rect 49535 11560 49549 11612
rect 49473 11508 49485 11560
rect 49537 11508 49549 11560
rect 49473 11496 49489 11508
rect 49009 11045 49055 11102
rect 49169 11091 49215 11102
rect 48369 10999 49055 11045
rect 48434 10752 48510 10764
rect 48434 10700 48446 10752
rect 48498 10749 48510 10752
rect 48594 10752 48670 10764
rect 48594 10749 48606 10752
rect 48498 10700 48606 10749
rect 48658 10700 48670 10752
rect 48434 10688 48670 10700
rect 48209 10616 48255 10627
rect 48369 10616 48415 10627
rect 47935 10210 47950 10222
rect 47874 10158 47886 10210
rect 47938 10158 47950 10210
rect 47874 10106 47889 10158
rect 47935 10106 47950 10158
rect 47874 10054 47886 10106
rect 47938 10054 47950 10106
rect 47874 10042 47889 10054
rect 47935 10042 47950 10054
rect 48193 10604 48209 10616
rect 48255 10604 48269 10616
rect 48193 10552 48205 10604
rect 48257 10552 48269 10604
rect 48193 10500 48209 10552
rect 48255 10500 48269 10552
rect 48193 10448 48205 10500
rect 48257 10448 48269 10500
rect 48193 10436 48209 10448
rect 47569 9556 47615 9567
rect 47729 9556 47775 10042
rect 47889 10031 47935 10042
rect 47295 9150 47310 9162
rect 47234 9098 47246 9150
rect 47298 9098 47310 9150
rect 47234 9046 47249 9098
rect 47295 9046 47310 9098
rect 47234 8994 47246 9046
rect 47298 8994 47310 9046
rect 47234 8982 47249 8994
rect 47295 8982 47310 8994
rect 47553 9544 47569 9556
rect 47615 9544 47629 9556
rect 47553 9492 47565 9544
rect 47617 9492 47629 9544
rect 47553 9440 47569 9492
rect 47615 9440 47629 9492
rect 47553 9388 47565 9440
rect 47617 9388 47629 9440
rect 47553 9376 47569 9388
rect 47121 8762 47167 8982
rect 47249 8971 47295 8982
rect 46961 8716 47041 8762
rect 47087 8716 47167 8762
rect 46961 8496 47007 8716
rect 46961 7579 47007 7922
rect 47121 8496 47167 8716
rect 47249 8496 47295 8507
rect 47234 8090 47249 8102
rect 47409 8496 47455 8982
rect 47615 9376 47629 9388
rect 47569 8971 47615 8982
rect 47889 9556 47935 9567
rect 47874 9150 47889 9162
rect 48049 9556 48095 10042
rect 48255 10436 48269 10448
rect 48209 10031 48255 10042
rect 48369 9985 48415 10042
rect 48529 10616 48575 10688
rect 48529 10031 48575 10042
rect 48689 10616 48735 10627
rect 48849 10616 48895 10627
rect 49009 10616 49055 10999
rect 48833 10604 48849 10616
rect 48895 10604 48909 10616
rect 48833 10552 48845 10604
rect 48897 10552 48909 10604
rect 48833 10500 48849 10552
rect 48895 10500 48909 10552
rect 48833 10448 48845 10500
rect 48897 10448 48909 10500
rect 48833 10436 48849 10448
rect 48689 9985 48735 10042
rect 48895 10436 48909 10448
rect 48849 10031 48895 10042
rect 49169 10616 49215 10627
rect 49154 10210 49169 10222
rect 49329 10616 49375 11102
rect 49535 11496 49549 11508
rect 49489 11091 49535 11102
rect 49809 11676 49855 11687
rect 49794 11270 49809 11282
rect 49937 11676 49983 12019
rect 49855 11270 49870 11282
rect 49794 11218 49806 11270
rect 49858 11218 49870 11270
rect 49794 11166 49809 11218
rect 49855 11166 49870 11218
rect 49794 11114 49806 11166
rect 49858 11114 49870 11166
rect 49794 11102 49809 11114
rect 49855 11102 49870 11114
rect 49489 10616 49535 10627
rect 49649 10616 49695 11102
rect 49809 11091 49855 11102
rect 49937 10882 49983 11102
rect 50097 11676 50143 12019
rect 50097 10882 50143 11102
rect 49937 10836 50017 10882
rect 50063 10836 50143 10882
rect 49215 10210 49230 10222
rect 49154 10158 49166 10210
rect 49218 10158 49230 10210
rect 49154 10106 49169 10158
rect 49215 10106 49230 10158
rect 49154 10054 49166 10106
rect 49218 10054 49230 10106
rect 49154 10042 49169 10054
rect 49215 10042 49230 10054
rect 49473 10604 49489 10616
rect 49535 10604 49549 10616
rect 49473 10552 49485 10604
rect 49537 10552 49549 10604
rect 49473 10500 49489 10552
rect 49535 10500 49549 10552
rect 49473 10448 49485 10500
rect 49537 10448 49549 10500
rect 49473 10436 49489 10448
rect 49009 9985 49055 10042
rect 49169 10031 49215 10042
rect 48369 9939 49055 9985
rect 48434 9692 48510 9704
rect 48434 9640 48446 9692
rect 48498 9689 48510 9692
rect 48594 9692 48670 9704
rect 48594 9689 48606 9692
rect 48498 9640 48606 9689
rect 48658 9640 48670 9692
rect 48434 9628 48670 9640
rect 48209 9556 48255 9567
rect 48369 9556 48415 9567
rect 47935 9150 47950 9162
rect 47874 9098 47886 9150
rect 47938 9098 47950 9150
rect 47874 9046 47889 9098
rect 47935 9046 47950 9098
rect 47874 8994 47886 9046
rect 47938 8994 47950 9046
rect 47874 8982 47889 8994
rect 47935 8982 47950 8994
rect 48193 9544 48209 9556
rect 48255 9544 48269 9556
rect 48193 9492 48205 9544
rect 48257 9492 48269 9544
rect 48193 9440 48209 9492
rect 48255 9440 48269 9492
rect 48193 9388 48205 9440
rect 48257 9388 48269 9440
rect 48193 9376 48209 9388
rect 47569 8496 47615 8507
rect 47729 8496 47775 8982
rect 47889 8971 47935 8982
rect 47295 8090 47310 8102
rect 47234 8038 47246 8090
rect 47298 8038 47310 8090
rect 47234 7986 47249 8038
rect 47295 7986 47310 8038
rect 47234 7934 47246 7986
rect 47298 7934 47310 7986
rect 47234 7922 47249 7934
rect 47295 7922 47310 7934
rect 47553 8484 47569 8496
rect 47615 8484 47629 8496
rect 47553 8432 47565 8484
rect 47617 8432 47629 8484
rect 47553 8380 47569 8432
rect 47615 8380 47629 8432
rect 47553 8328 47565 8380
rect 47617 8328 47629 8380
rect 47553 8316 47569 8328
rect 47121 7579 47167 7922
rect 47249 7911 47295 7922
rect 47409 7579 47455 7922
rect 47615 8316 47629 8328
rect 47569 7911 47615 7922
rect 47889 8496 47935 8507
rect 47874 8090 47889 8102
rect 48049 8496 48095 8982
rect 48255 9376 48269 9388
rect 48209 8971 48255 8982
rect 48369 8925 48415 8982
rect 48529 9556 48575 9628
rect 48529 8971 48575 8982
rect 48689 9556 48735 9567
rect 48849 9556 48895 9567
rect 49009 9556 49055 9939
rect 48833 9544 48849 9556
rect 48895 9544 48909 9556
rect 48833 9492 48845 9544
rect 48897 9492 48909 9544
rect 48833 9440 48849 9492
rect 48895 9440 48909 9492
rect 48833 9388 48845 9440
rect 48897 9388 48909 9440
rect 48833 9376 48849 9388
rect 48689 8925 48735 8982
rect 48895 9376 48909 9388
rect 48849 8971 48895 8982
rect 49169 9556 49215 9567
rect 49154 9150 49169 9162
rect 49329 9556 49375 10042
rect 49535 10436 49549 10448
rect 49489 10031 49535 10042
rect 49809 10616 49855 10627
rect 49794 10210 49809 10222
rect 49937 10616 49983 10836
rect 49855 10210 49870 10222
rect 49794 10158 49806 10210
rect 49858 10158 49870 10210
rect 49794 10106 49809 10158
rect 49855 10106 49870 10158
rect 49794 10054 49806 10106
rect 49858 10054 49870 10106
rect 49794 10042 49809 10054
rect 49855 10042 49870 10054
rect 49489 9556 49535 9567
rect 49649 9556 49695 10042
rect 49809 10031 49855 10042
rect 49215 9150 49230 9162
rect 49154 9098 49166 9150
rect 49218 9098 49230 9150
rect 49154 9046 49169 9098
rect 49215 9046 49230 9098
rect 49154 8994 49166 9046
rect 49218 8994 49230 9046
rect 49154 8982 49169 8994
rect 49215 8982 49230 8994
rect 49473 9544 49489 9556
rect 49535 9544 49549 9556
rect 49473 9492 49485 9544
rect 49537 9492 49549 9544
rect 49473 9440 49489 9492
rect 49535 9440 49549 9492
rect 49473 9388 49485 9440
rect 49537 9388 49549 9440
rect 49473 9376 49489 9388
rect 49009 8925 49055 8982
rect 49169 8971 49215 8982
rect 48369 8879 49055 8925
rect 48434 8632 48510 8644
rect 48434 8580 48446 8632
rect 48498 8629 48510 8632
rect 48594 8632 48670 8644
rect 48594 8629 48606 8632
rect 48498 8580 48606 8629
rect 48658 8580 48670 8632
rect 48434 8568 48670 8580
rect 48209 8496 48255 8507
rect 48369 8496 48415 8507
rect 47935 8090 47950 8102
rect 47874 8038 47886 8090
rect 47938 8038 47950 8090
rect 47874 7986 47889 8038
rect 47935 7986 47950 8038
rect 47874 7934 47886 7986
rect 47938 7934 47950 7986
rect 47874 7922 47889 7934
rect 47935 7922 47950 7934
rect 48193 8484 48209 8496
rect 48255 8484 48269 8496
rect 48193 8432 48205 8484
rect 48257 8432 48269 8484
rect 48193 8380 48209 8432
rect 48255 8380 48269 8432
rect 48193 8328 48205 8380
rect 48257 8328 48269 8380
rect 48193 8316 48209 8328
rect 47729 7579 47775 7922
rect 47889 7911 47935 7922
rect 48049 7579 48095 7922
rect 48255 8316 48269 8328
rect 48209 7911 48255 7922
rect 48369 7579 48415 7922
rect 48529 8496 48575 8568
rect 48529 7911 48575 7922
rect 48689 8496 48735 8507
rect 48849 8496 48895 8507
rect 49009 8496 49055 8879
rect 48833 8484 48849 8496
rect 48895 8484 48909 8496
rect 48833 8432 48845 8484
rect 48897 8432 48909 8484
rect 48833 8380 48849 8432
rect 48895 8380 48909 8432
rect 48833 8328 48845 8380
rect 48897 8328 48909 8380
rect 48833 8316 48849 8328
rect 48689 7579 48735 7922
rect 48895 8316 48909 8328
rect 48849 7911 48895 7922
rect 49169 8496 49215 8507
rect 49154 8090 49169 8102
rect 49329 8496 49375 8982
rect 49535 9376 49549 9388
rect 49489 8971 49535 8982
rect 49809 9556 49855 9567
rect 49794 9150 49809 9162
rect 49937 9556 49983 10042
rect 49855 9150 49870 9162
rect 49794 9098 49806 9150
rect 49858 9098 49870 9150
rect 49794 9046 49809 9098
rect 49855 9046 49870 9098
rect 49794 8994 49806 9046
rect 49858 8994 49870 9046
rect 49794 8982 49809 8994
rect 49855 8982 49870 8994
rect 49489 8496 49535 8507
rect 49649 8496 49695 8982
rect 49809 8971 49855 8982
rect 49937 8762 49983 8982
rect 50097 10616 50143 10836
rect 50097 9556 50143 10042
rect 50097 8762 50143 8982
rect 49937 8716 50017 8762
rect 50063 8716 50143 8762
rect 49215 8090 49230 8102
rect 49154 8038 49166 8090
rect 49218 8038 49230 8090
rect 49154 7986 49169 8038
rect 49215 7986 49230 8038
rect 49154 7934 49166 7986
rect 49218 7934 49230 7986
rect 49154 7922 49169 7934
rect 49215 7922 49230 7934
rect 49473 8484 49489 8496
rect 49535 8484 49549 8496
rect 49473 8432 49485 8484
rect 49537 8432 49549 8484
rect 49473 8380 49489 8432
rect 49535 8380 49549 8432
rect 49473 8328 49485 8380
rect 49537 8328 49549 8380
rect 49473 8316 49489 8328
rect 49009 7579 49055 7922
rect 49169 7911 49215 7922
rect 49329 7579 49375 7922
rect 49535 8316 49549 8328
rect 49489 7911 49535 7922
rect 49809 8496 49855 8507
rect 49794 8090 49809 8102
rect 49937 8496 49983 8716
rect 49855 8090 49870 8102
rect 49794 8038 49806 8090
rect 49858 8038 49870 8090
rect 49794 7986 49809 8038
rect 49855 7986 49870 8038
rect 49794 7934 49806 7986
rect 49858 7934 49870 7986
rect 49794 7922 49809 7934
rect 49855 7922 49870 7934
rect 49649 7579 49695 7922
rect 49809 7911 49855 7922
rect 49937 7579 49983 7922
rect 50097 8496 50143 8716
rect 50097 7579 50143 7922
rect 50442 11985 50597 12019
rect 50643 12019 52021 12031
rect 50643 11985 50762 12019
rect 50442 11937 50762 11985
rect 50442 11891 50597 11937
rect 50643 11891 50762 11937
rect 50442 11843 50762 11891
rect 50442 11797 50597 11843
rect 50643 11797 50762 11843
rect 50442 11749 50762 11797
rect 50442 11703 50597 11749
rect 50643 11703 50762 11749
rect 50442 11655 50762 11703
rect 50442 11609 50597 11655
rect 50643 11609 50762 11655
rect 50442 11561 50762 11609
rect 50442 11515 50597 11561
rect 50643 11515 50762 11561
rect 50442 11467 50762 11515
rect 50442 11421 50597 11467
rect 50643 11421 50762 11467
rect 50442 11373 50762 11421
rect 50442 11327 50597 11373
rect 50643 11327 50762 11373
rect 50442 11279 50762 11327
rect 50442 11233 50597 11279
rect 50643 11233 50762 11279
rect 50442 11185 50762 11233
rect 50442 11139 50597 11185
rect 50643 11139 50762 11185
rect 50442 11091 50762 11139
rect 50442 11045 50597 11091
rect 50643 11045 50762 11091
rect 50442 10997 50762 11045
rect 50442 10951 50597 10997
rect 50643 10951 50762 10997
rect 50442 10903 50762 10951
rect 50442 10857 50597 10903
rect 50643 10857 50762 10903
rect 50442 10809 50762 10857
rect 50442 10763 50597 10809
rect 50643 10763 50762 10809
rect 50442 10715 50762 10763
rect 50442 10669 50597 10715
rect 50643 10669 50762 10715
rect 50442 10621 50762 10669
rect 50442 10575 50597 10621
rect 50643 10575 50762 10621
rect 50442 10527 50762 10575
rect 50442 10481 50597 10527
rect 50643 10481 50762 10527
rect 50442 10433 50762 10481
rect 50442 10387 50597 10433
rect 50643 10387 50762 10433
rect 50442 10339 50762 10387
rect 50442 10293 50597 10339
rect 50643 10293 50762 10339
rect 50442 10245 50762 10293
rect 50442 10199 50597 10245
rect 50643 10199 50762 10245
rect 50442 10151 50762 10199
rect 50442 10105 50597 10151
rect 50643 10105 50762 10151
rect 50442 10057 50762 10105
rect 50442 10011 50597 10057
rect 50643 10011 50762 10057
rect 50442 9963 50762 10011
rect 50442 9917 50597 9963
rect 50643 9917 50762 9963
rect 50442 9869 50762 9917
rect 50442 9823 50597 9869
rect 50643 9823 50762 9869
rect 50442 9775 50762 9823
rect 50442 9729 50597 9775
rect 50643 9729 50762 9775
rect 50442 9681 50762 9729
rect 50442 9635 50597 9681
rect 50643 9635 50762 9681
rect 50442 9587 50762 9635
rect 50442 9541 50597 9587
rect 50643 9541 50762 9587
rect 50442 9493 50762 9541
rect 50442 9447 50597 9493
rect 50643 9447 50762 9493
rect 50442 9399 50762 9447
rect 50442 9353 50597 9399
rect 50643 9353 50762 9399
rect 50442 9305 50762 9353
rect 50442 9259 50597 9305
rect 50643 9259 50762 9305
rect 50442 9211 50762 9259
rect 50442 9165 50597 9211
rect 50643 9165 50762 9211
rect 50442 9117 50762 9165
rect 50442 9071 50597 9117
rect 50643 9071 50762 9117
rect 50442 9023 50762 9071
rect 50442 8977 50597 9023
rect 50643 8977 50762 9023
rect 50442 8929 50762 8977
rect 50442 8883 50597 8929
rect 50643 8883 50762 8929
rect 50442 8835 50762 8883
rect 50442 8789 50597 8835
rect 50643 8789 50762 8835
rect 50442 8741 50762 8789
rect 50442 8695 50597 8741
rect 50643 8695 50762 8741
rect 50442 8647 50762 8695
rect 50442 8601 50597 8647
rect 50643 8601 50762 8647
rect 50442 8553 50762 8601
rect 50442 8507 50597 8553
rect 50643 8507 50762 8553
rect 50442 8459 50762 8507
rect 50442 8413 50597 8459
rect 50643 8413 50762 8459
rect 50442 8365 50762 8413
rect 50442 8319 50597 8365
rect 50643 8319 50762 8365
rect 50442 8271 50762 8319
rect 50442 8225 50597 8271
rect 50643 8225 50762 8271
rect 50442 8177 50762 8225
rect 50442 8131 50597 8177
rect 50643 8131 50762 8177
rect 50442 8083 50762 8131
rect 50442 8037 50597 8083
rect 50643 8037 50762 8083
rect 50442 7989 50762 8037
rect 50442 7943 50597 7989
rect 50643 7943 50762 7989
rect 50442 7895 50762 7943
rect 50442 7849 50597 7895
rect 50643 7849 50762 7895
rect 50442 7801 50762 7849
rect 50442 7755 50597 7801
rect 50643 7755 50762 7801
rect 50442 7707 50762 7755
rect 50442 7661 50597 7707
rect 50643 7661 50762 7707
rect 50442 7613 50762 7661
rect 50442 7579 50597 7613
rect 46507 7567 50597 7579
rect 50643 7579 50762 7613
rect 51902 11985 52021 12019
rect 52067 12019 56157 12031
rect 52067 11985 52222 12019
rect 51902 11937 52222 11985
rect 51902 11891 52021 11937
rect 52067 11891 52222 11937
rect 51902 11843 52222 11891
rect 51902 11797 52021 11843
rect 52067 11797 52222 11843
rect 51902 11749 52222 11797
rect 51902 11703 52021 11749
rect 52067 11703 52222 11749
rect 51902 11655 52222 11703
rect 51902 11609 52021 11655
rect 52067 11609 52222 11655
rect 51902 11561 52222 11609
rect 51902 11515 52021 11561
rect 52067 11515 52222 11561
rect 51902 11467 52222 11515
rect 51902 11421 52021 11467
rect 52067 11421 52222 11467
rect 51902 11373 52222 11421
rect 51902 11327 52021 11373
rect 52067 11327 52222 11373
rect 51902 11279 52222 11327
rect 51902 11233 52021 11279
rect 52067 11233 52222 11279
rect 51902 11185 52222 11233
rect 51902 11139 52021 11185
rect 52067 11139 52222 11185
rect 51902 11091 52222 11139
rect 51902 11045 52021 11091
rect 52067 11045 52222 11091
rect 51902 10997 52222 11045
rect 51902 10951 52021 10997
rect 52067 10951 52222 10997
rect 51902 10903 52222 10951
rect 51902 10857 52021 10903
rect 52067 10857 52222 10903
rect 51902 10809 52222 10857
rect 51902 10763 52021 10809
rect 52067 10763 52222 10809
rect 51902 10715 52222 10763
rect 51902 10669 52021 10715
rect 52067 10669 52222 10715
rect 51902 10621 52222 10669
rect 51902 10575 52021 10621
rect 52067 10575 52222 10621
rect 51902 10527 52222 10575
rect 51902 10481 52021 10527
rect 52067 10481 52222 10527
rect 51902 10433 52222 10481
rect 51902 10387 52021 10433
rect 52067 10387 52222 10433
rect 51902 10339 52222 10387
rect 51902 10293 52021 10339
rect 52067 10293 52222 10339
rect 51902 10245 52222 10293
rect 51902 10199 52021 10245
rect 52067 10199 52222 10245
rect 51902 10151 52222 10199
rect 51902 10105 52021 10151
rect 52067 10105 52222 10151
rect 51902 10057 52222 10105
rect 51902 10011 52021 10057
rect 52067 10011 52222 10057
rect 51902 9963 52222 10011
rect 51902 9917 52021 9963
rect 52067 9917 52222 9963
rect 51902 9869 52222 9917
rect 51902 9823 52021 9869
rect 52067 9823 52222 9869
rect 51902 9775 52222 9823
rect 51902 9729 52021 9775
rect 52067 9729 52222 9775
rect 51902 9681 52222 9729
rect 51902 9635 52021 9681
rect 52067 9635 52222 9681
rect 51902 9587 52222 9635
rect 51902 9541 52021 9587
rect 52067 9541 52222 9587
rect 51902 9493 52222 9541
rect 51902 9447 52021 9493
rect 52067 9447 52222 9493
rect 51902 9399 52222 9447
rect 51902 9353 52021 9399
rect 52067 9353 52222 9399
rect 51902 9305 52222 9353
rect 51902 9259 52021 9305
rect 52067 9259 52222 9305
rect 51902 9211 52222 9259
rect 51902 9165 52021 9211
rect 52067 9165 52222 9211
rect 51902 9117 52222 9165
rect 51902 9071 52021 9117
rect 52067 9071 52222 9117
rect 51902 9023 52222 9071
rect 51902 8977 52021 9023
rect 52067 8977 52222 9023
rect 51902 8929 52222 8977
rect 51902 8883 52021 8929
rect 52067 8883 52222 8929
rect 51902 8835 52222 8883
rect 51902 8789 52021 8835
rect 52067 8789 52222 8835
rect 51902 8741 52222 8789
rect 51902 8695 52021 8741
rect 52067 8695 52222 8741
rect 51902 8647 52222 8695
rect 51902 8601 52021 8647
rect 52067 8601 52222 8647
rect 51902 8553 52222 8601
rect 51902 8507 52021 8553
rect 52067 8507 52222 8553
rect 51902 8459 52222 8507
rect 51902 8413 52021 8459
rect 52067 8413 52222 8459
rect 51902 8365 52222 8413
rect 51902 8319 52021 8365
rect 52067 8319 52222 8365
rect 51902 8271 52222 8319
rect 51902 8225 52021 8271
rect 52067 8225 52222 8271
rect 51902 8177 52222 8225
rect 51902 8131 52021 8177
rect 52067 8131 52222 8177
rect 51902 8083 52222 8131
rect 51902 8037 52021 8083
rect 52067 8037 52222 8083
rect 51902 7989 52222 8037
rect 51902 7943 52021 7989
rect 52067 7943 52222 7989
rect 51902 7895 52222 7943
rect 51902 7849 52021 7895
rect 52067 7849 52222 7895
rect 51902 7801 52222 7849
rect 51902 7755 52021 7801
rect 52067 7755 52222 7801
rect 51902 7707 52222 7755
rect 51902 7661 52021 7707
rect 52067 7661 52222 7707
rect 51902 7613 52222 7661
rect 51902 7579 52021 7613
rect 50643 7567 52021 7579
rect 52067 7579 52222 7613
rect 52521 11676 52567 12019
rect 52521 10882 52567 11102
rect 52681 11676 52727 12019
rect 52809 11676 52855 11687
rect 52794 11270 52809 11282
rect 52969 11676 53015 12019
rect 53129 11676 53175 11687
rect 53289 11676 53335 12019
rect 52855 11270 52870 11282
rect 52794 11218 52806 11270
rect 52858 11218 52870 11270
rect 52794 11166 52809 11218
rect 52855 11166 52870 11218
rect 52794 11114 52806 11166
rect 52858 11114 52870 11166
rect 52794 11102 52809 11114
rect 52855 11102 52870 11114
rect 53115 11664 53129 11676
rect 53175 11664 53191 11676
rect 53115 11612 53127 11664
rect 53179 11612 53191 11664
rect 53115 11560 53129 11612
rect 53175 11560 53191 11612
rect 53115 11508 53127 11560
rect 53179 11508 53191 11560
rect 53115 11496 53129 11508
rect 52681 10882 52727 11102
rect 52809 11091 52855 11102
rect 52521 10836 52601 10882
rect 52647 10836 52727 10882
rect 52521 10616 52567 10836
rect 52521 9556 52567 10042
rect 52521 8762 52567 8982
rect 52681 10616 52727 10836
rect 52809 10616 52855 10627
rect 52794 10210 52809 10222
rect 52969 10616 53015 11102
rect 53175 11496 53191 11508
rect 53129 11091 53175 11102
rect 53449 11676 53495 11687
rect 53434 11270 53449 11282
rect 53609 11676 53655 12019
rect 53994 11812 54070 11824
rect 53994 11760 54006 11812
rect 54058 11809 54070 11812
rect 54154 11812 54230 11824
rect 54154 11809 54166 11812
rect 54058 11760 54166 11809
rect 54218 11760 54230 11812
rect 53994 11748 54230 11760
rect 53769 11676 53815 11687
rect 53929 11676 53975 11687
rect 53495 11270 53510 11282
rect 53434 11218 53446 11270
rect 53498 11218 53510 11270
rect 53434 11166 53449 11218
rect 53495 11166 53510 11218
rect 53434 11114 53446 11166
rect 53498 11114 53510 11166
rect 53434 11102 53449 11114
rect 53495 11102 53510 11114
rect 53755 11664 53769 11676
rect 53815 11664 53831 11676
rect 53755 11612 53767 11664
rect 53819 11612 53831 11664
rect 53755 11560 53769 11612
rect 53815 11560 53831 11612
rect 53755 11508 53767 11560
rect 53819 11508 53831 11560
rect 53755 11496 53769 11508
rect 53129 10616 53175 10627
rect 53289 10616 53335 11102
rect 53449 11091 53495 11102
rect 53609 11045 53655 11102
rect 53815 11496 53831 11508
rect 53769 11091 53815 11102
rect 53929 11045 53975 11102
rect 54089 11676 54135 11748
rect 54089 11091 54135 11102
rect 54249 11676 54295 11687
rect 54409 11676 54455 11687
rect 54569 11676 54615 12019
rect 54395 11664 54409 11676
rect 54455 11664 54471 11676
rect 54395 11612 54407 11664
rect 54459 11612 54471 11664
rect 54395 11560 54409 11612
rect 54455 11560 54471 11612
rect 54395 11508 54407 11560
rect 54459 11508 54471 11560
rect 54395 11496 54409 11508
rect 54249 11045 54295 11102
rect 54455 11496 54471 11508
rect 54409 11091 54455 11102
rect 54729 11676 54775 11687
rect 54714 11270 54729 11282
rect 54889 11676 54935 12019
rect 55049 11676 55095 11687
rect 55209 11676 55255 12019
rect 54775 11270 54790 11282
rect 54714 11218 54726 11270
rect 54778 11218 54790 11270
rect 54714 11166 54729 11218
rect 54775 11166 54790 11218
rect 54714 11114 54726 11166
rect 54778 11114 54790 11166
rect 54714 11102 54729 11114
rect 54775 11102 54790 11114
rect 55035 11664 55049 11676
rect 55095 11664 55111 11676
rect 55035 11612 55047 11664
rect 55099 11612 55111 11664
rect 55035 11560 55049 11612
rect 55095 11560 55111 11612
rect 55035 11508 55047 11560
rect 55099 11508 55111 11560
rect 55035 11496 55049 11508
rect 53609 10999 54295 11045
rect 52855 10210 52870 10222
rect 52794 10158 52806 10210
rect 52858 10158 52870 10210
rect 52794 10106 52809 10158
rect 52855 10106 52870 10158
rect 52794 10054 52806 10106
rect 52858 10054 52870 10106
rect 52794 10042 52809 10054
rect 52855 10042 52870 10054
rect 53115 10604 53129 10616
rect 53175 10604 53191 10616
rect 53115 10552 53127 10604
rect 53179 10552 53191 10604
rect 53115 10500 53129 10552
rect 53175 10500 53191 10552
rect 53115 10448 53127 10500
rect 53179 10448 53191 10500
rect 53115 10436 53129 10448
rect 52681 9556 52727 10042
rect 52809 10031 52855 10042
rect 52809 9556 52855 9567
rect 52794 9150 52809 9162
rect 52969 9556 53015 10042
rect 53175 10436 53191 10448
rect 53129 10031 53175 10042
rect 53449 10616 53495 10627
rect 53434 10210 53449 10222
rect 53609 10616 53655 10999
rect 53994 10752 54070 10764
rect 53994 10700 54006 10752
rect 54058 10749 54070 10752
rect 54154 10752 54230 10764
rect 54154 10749 54166 10752
rect 54058 10700 54166 10749
rect 54218 10700 54230 10752
rect 53994 10688 54230 10700
rect 53769 10616 53815 10627
rect 53929 10616 53975 10627
rect 53495 10210 53510 10222
rect 53434 10158 53446 10210
rect 53498 10158 53510 10210
rect 53434 10106 53449 10158
rect 53495 10106 53510 10158
rect 53434 10054 53446 10106
rect 53498 10054 53510 10106
rect 53434 10042 53449 10054
rect 53495 10042 53510 10054
rect 53755 10604 53769 10616
rect 53815 10604 53831 10616
rect 53755 10552 53767 10604
rect 53819 10552 53831 10604
rect 53755 10500 53769 10552
rect 53815 10500 53831 10552
rect 53755 10448 53767 10500
rect 53819 10448 53831 10500
rect 53755 10436 53769 10448
rect 53129 9556 53175 9567
rect 53289 9556 53335 10042
rect 53449 10031 53495 10042
rect 53609 9985 53655 10042
rect 53815 10436 53831 10448
rect 53769 10031 53815 10042
rect 53929 9985 53975 10042
rect 54089 10616 54135 10688
rect 54089 10031 54135 10042
rect 54249 10616 54295 10627
rect 54409 10616 54455 10627
rect 54569 10616 54615 11102
rect 54729 11091 54775 11102
rect 54395 10604 54409 10616
rect 54455 10604 54471 10616
rect 54395 10552 54407 10604
rect 54459 10552 54471 10604
rect 54395 10500 54409 10552
rect 54455 10500 54471 10552
rect 54395 10448 54407 10500
rect 54459 10448 54471 10500
rect 54395 10436 54409 10448
rect 54249 9985 54295 10042
rect 54455 10436 54471 10448
rect 54409 10031 54455 10042
rect 54729 10616 54775 10627
rect 54714 10210 54729 10222
rect 54889 10616 54935 11102
rect 55095 11496 55111 11508
rect 55049 11091 55095 11102
rect 55369 11676 55415 11687
rect 55354 11270 55369 11282
rect 55497 11676 55543 12019
rect 55415 11270 55430 11282
rect 55354 11218 55366 11270
rect 55418 11218 55430 11270
rect 55354 11166 55369 11218
rect 55415 11166 55430 11218
rect 55354 11114 55366 11166
rect 55418 11114 55430 11166
rect 55354 11102 55369 11114
rect 55415 11102 55430 11114
rect 55049 10616 55095 10627
rect 55209 10616 55255 11102
rect 55369 11091 55415 11102
rect 55497 10882 55543 11102
rect 55657 11676 55703 12019
rect 55657 10882 55703 11102
rect 55497 10836 55577 10882
rect 55623 10836 55703 10882
rect 54775 10210 54790 10222
rect 54714 10158 54726 10210
rect 54778 10158 54790 10210
rect 54714 10106 54729 10158
rect 54775 10106 54790 10158
rect 54714 10054 54726 10106
rect 54778 10054 54790 10106
rect 54714 10042 54729 10054
rect 54775 10042 54790 10054
rect 55035 10604 55049 10616
rect 55095 10604 55111 10616
rect 55035 10552 55047 10604
rect 55099 10552 55111 10604
rect 55035 10500 55049 10552
rect 55095 10500 55111 10552
rect 55035 10448 55047 10500
rect 55099 10448 55111 10500
rect 55035 10436 55049 10448
rect 53609 9939 54295 9985
rect 52855 9150 52870 9162
rect 52794 9098 52806 9150
rect 52858 9098 52870 9150
rect 52794 9046 52809 9098
rect 52855 9046 52870 9098
rect 52794 8994 52806 9046
rect 52858 8994 52870 9046
rect 52794 8982 52809 8994
rect 52855 8982 52870 8994
rect 53115 9544 53129 9556
rect 53175 9544 53191 9556
rect 53115 9492 53127 9544
rect 53179 9492 53191 9544
rect 53115 9440 53129 9492
rect 53175 9440 53191 9492
rect 53115 9388 53127 9440
rect 53179 9388 53191 9440
rect 53115 9376 53129 9388
rect 52681 8762 52727 8982
rect 52809 8971 52855 8982
rect 52521 8716 52601 8762
rect 52647 8716 52727 8762
rect 52521 8496 52567 8716
rect 52521 7579 52567 7922
rect 52681 8496 52727 8716
rect 52809 8496 52855 8507
rect 52794 8090 52809 8102
rect 52969 8496 53015 8982
rect 53175 9376 53191 9388
rect 53129 8971 53175 8982
rect 53449 9556 53495 9567
rect 53434 9150 53449 9162
rect 53609 9556 53655 9939
rect 53994 9692 54070 9704
rect 53994 9640 54006 9692
rect 54058 9689 54070 9692
rect 54154 9692 54230 9704
rect 54154 9689 54166 9692
rect 54058 9640 54166 9689
rect 54218 9640 54230 9692
rect 53994 9628 54230 9640
rect 53769 9556 53815 9567
rect 53929 9556 53975 9567
rect 53495 9150 53510 9162
rect 53434 9098 53446 9150
rect 53498 9098 53510 9150
rect 53434 9046 53449 9098
rect 53495 9046 53510 9098
rect 53434 8994 53446 9046
rect 53498 8994 53510 9046
rect 53434 8982 53449 8994
rect 53495 8982 53510 8994
rect 53755 9544 53769 9556
rect 53815 9544 53831 9556
rect 53755 9492 53767 9544
rect 53819 9492 53831 9544
rect 53755 9440 53769 9492
rect 53815 9440 53831 9492
rect 53755 9388 53767 9440
rect 53819 9388 53831 9440
rect 53755 9376 53769 9388
rect 53129 8496 53175 8507
rect 53289 8496 53335 8982
rect 53449 8971 53495 8982
rect 53609 8925 53655 8982
rect 53815 9376 53831 9388
rect 53769 8971 53815 8982
rect 53929 8925 53975 8982
rect 54089 9556 54135 9628
rect 54089 8971 54135 8982
rect 54249 9556 54295 9567
rect 54409 9556 54455 9567
rect 54569 9556 54615 10042
rect 54729 10031 54775 10042
rect 54395 9544 54409 9556
rect 54455 9544 54471 9556
rect 54395 9492 54407 9544
rect 54459 9492 54471 9544
rect 54395 9440 54409 9492
rect 54455 9440 54471 9492
rect 54395 9388 54407 9440
rect 54459 9388 54471 9440
rect 54395 9376 54409 9388
rect 54249 8925 54295 8982
rect 54455 9376 54471 9388
rect 54409 8971 54455 8982
rect 54729 9556 54775 9567
rect 54714 9150 54729 9162
rect 54889 9556 54935 10042
rect 55095 10436 55111 10448
rect 55049 10031 55095 10042
rect 55369 10616 55415 10627
rect 55354 10210 55369 10222
rect 55497 10616 55543 10836
rect 55415 10210 55430 10222
rect 55354 10158 55366 10210
rect 55418 10158 55430 10210
rect 55354 10106 55369 10158
rect 55415 10106 55430 10158
rect 55354 10054 55366 10106
rect 55418 10054 55430 10106
rect 55354 10042 55369 10054
rect 55415 10042 55430 10054
rect 55049 9556 55095 9567
rect 55209 9556 55255 10042
rect 55369 10031 55415 10042
rect 54775 9150 54790 9162
rect 54714 9098 54726 9150
rect 54778 9098 54790 9150
rect 54714 9046 54729 9098
rect 54775 9046 54790 9098
rect 54714 8994 54726 9046
rect 54778 8994 54790 9046
rect 54714 8982 54729 8994
rect 54775 8982 54790 8994
rect 55035 9544 55049 9556
rect 55095 9544 55111 9556
rect 55035 9492 55047 9544
rect 55099 9492 55111 9544
rect 55035 9440 55049 9492
rect 55095 9440 55111 9492
rect 55035 9388 55047 9440
rect 55099 9388 55111 9440
rect 55035 9376 55049 9388
rect 53609 8879 54295 8925
rect 52855 8090 52870 8102
rect 52794 8038 52806 8090
rect 52858 8038 52870 8090
rect 52794 7986 52809 8038
rect 52855 7986 52870 8038
rect 52794 7934 52806 7986
rect 52858 7934 52870 7986
rect 52794 7922 52809 7934
rect 52855 7922 52870 7934
rect 53115 8484 53129 8496
rect 53175 8484 53191 8496
rect 53115 8432 53127 8484
rect 53179 8432 53191 8484
rect 53115 8380 53129 8432
rect 53175 8380 53191 8432
rect 53115 8328 53127 8380
rect 53179 8328 53191 8380
rect 53115 8316 53129 8328
rect 52681 7579 52727 7922
rect 52809 7911 52855 7922
rect 52969 7579 53015 7922
rect 53175 8316 53191 8328
rect 53129 7911 53175 7922
rect 53449 8496 53495 8507
rect 53434 8090 53449 8102
rect 53609 8496 53655 8879
rect 53994 8632 54070 8644
rect 53994 8580 54006 8632
rect 54058 8629 54070 8632
rect 54154 8632 54230 8644
rect 54154 8629 54166 8632
rect 54058 8580 54166 8629
rect 54218 8580 54230 8632
rect 53994 8568 54230 8580
rect 53769 8496 53815 8507
rect 53929 8496 53975 8507
rect 53495 8090 53510 8102
rect 53434 8038 53446 8090
rect 53498 8038 53510 8090
rect 53434 7986 53449 8038
rect 53495 7986 53510 8038
rect 53434 7934 53446 7986
rect 53498 7934 53510 7986
rect 53434 7922 53449 7934
rect 53495 7922 53510 7934
rect 53755 8484 53769 8496
rect 53815 8484 53831 8496
rect 53755 8432 53767 8484
rect 53819 8432 53831 8484
rect 53755 8380 53769 8432
rect 53815 8380 53831 8432
rect 53755 8328 53767 8380
rect 53819 8328 53831 8380
rect 53755 8316 53769 8328
rect 53289 7579 53335 7922
rect 53449 7911 53495 7922
rect 53609 7579 53655 7922
rect 53815 8316 53831 8328
rect 53769 7911 53815 7922
rect 53929 7579 53975 7922
rect 54089 8496 54135 8568
rect 54089 7911 54135 7922
rect 54249 8496 54295 8507
rect 54409 8496 54455 8507
rect 54569 8496 54615 8982
rect 54729 8971 54775 8982
rect 54395 8484 54409 8496
rect 54455 8484 54471 8496
rect 54395 8432 54407 8484
rect 54459 8432 54471 8484
rect 54395 8380 54409 8432
rect 54455 8380 54471 8432
rect 54395 8328 54407 8380
rect 54459 8328 54471 8380
rect 54395 8316 54409 8328
rect 54249 7579 54295 7922
rect 54455 8316 54471 8328
rect 54409 7911 54455 7922
rect 54729 8496 54775 8507
rect 54714 8090 54729 8102
rect 54889 8496 54935 8982
rect 55095 9376 55111 9388
rect 55049 8971 55095 8982
rect 55369 9556 55415 9567
rect 55354 9150 55369 9162
rect 55497 9556 55543 10042
rect 55415 9150 55430 9162
rect 55354 9098 55366 9150
rect 55418 9098 55430 9150
rect 55354 9046 55369 9098
rect 55415 9046 55430 9098
rect 55354 8994 55366 9046
rect 55418 8994 55430 9046
rect 55354 8982 55369 8994
rect 55415 8982 55430 8994
rect 55049 8496 55095 8507
rect 55209 8496 55255 8982
rect 55369 8971 55415 8982
rect 55497 8762 55543 8982
rect 55657 10616 55703 10836
rect 55657 9556 55703 10042
rect 55657 8762 55703 8982
rect 55497 8716 55577 8762
rect 55623 8716 55703 8762
rect 54775 8090 54790 8102
rect 54714 8038 54726 8090
rect 54778 8038 54790 8090
rect 54714 7986 54729 8038
rect 54775 7986 54790 8038
rect 54714 7934 54726 7986
rect 54778 7934 54790 7986
rect 54714 7922 54729 7934
rect 54775 7922 54790 7934
rect 55035 8484 55049 8496
rect 55095 8484 55111 8496
rect 55035 8432 55047 8484
rect 55099 8432 55111 8484
rect 55035 8380 55049 8432
rect 55095 8380 55111 8432
rect 55035 8328 55047 8380
rect 55099 8328 55111 8380
rect 55035 8316 55049 8328
rect 54569 7579 54615 7922
rect 54729 7911 54775 7922
rect 54889 7579 54935 7922
rect 55095 8316 55111 8328
rect 55049 7911 55095 7922
rect 55369 8496 55415 8507
rect 55354 8090 55369 8102
rect 55497 8496 55543 8716
rect 55415 8090 55430 8102
rect 55354 8038 55366 8090
rect 55418 8038 55430 8090
rect 55354 7986 55369 8038
rect 55415 7986 55430 8038
rect 55354 7934 55366 7986
rect 55418 7934 55430 7986
rect 55354 7922 55369 7934
rect 55415 7922 55430 7934
rect 55209 7579 55255 7922
rect 55369 7911 55415 7922
rect 55497 7579 55543 7922
rect 55657 8496 55703 8716
rect 55657 7579 55703 7922
rect 56002 11985 56157 12019
rect 56203 12019 60293 12031
rect 56203 11985 56358 12019
rect 56002 11937 56358 11985
rect 56002 11891 56157 11937
rect 56203 11891 56358 11937
rect 56002 11843 56358 11891
rect 56002 11797 56157 11843
rect 56203 11797 56358 11843
rect 56002 11749 56358 11797
rect 56002 11703 56157 11749
rect 56203 11703 56358 11749
rect 56002 11655 56358 11703
rect 56002 11609 56157 11655
rect 56203 11609 56358 11655
rect 56002 11561 56358 11609
rect 56002 11515 56157 11561
rect 56203 11515 56358 11561
rect 56002 11467 56358 11515
rect 56002 11421 56157 11467
rect 56203 11421 56358 11467
rect 56002 11373 56358 11421
rect 56002 11327 56157 11373
rect 56203 11327 56358 11373
rect 56002 11279 56358 11327
rect 56002 11233 56157 11279
rect 56203 11233 56358 11279
rect 56002 11185 56358 11233
rect 56002 11139 56157 11185
rect 56203 11139 56358 11185
rect 56002 11091 56358 11139
rect 56002 11045 56157 11091
rect 56203 11045 56358 11091
rect 56002 10997 56358 11045
rect 56002 10951 56157 10997
rect 56203 10951 56358 10997
rect 56002 10903 56358 10951
rect 56002 10857 56157 10903
rect 56203 10857 56358 10903
rect 56002 10809 56358 10857
rect 56002 10763 56157 10809
rect 56203 10763 56358 10809
rect 56002 10715 56358 10763
rect 56002 10669 56157 10715
rect 56203 10669 56358 10715
rect 56002 10621 56358 10669
rect 56002 10575 56157 10621
rect 56203 10575 56358 10621
rect 56002 10527 56358 10575
rect 56002 10481 56157 10527
rect 56203 10481 56358 10527
rect 56002 10433 56358 10481
rect 56002 10387 56157 10433
rect 56203 10387 56358 10433
rect 56002 10339 56358 10387
rect 56002 10293 56157 10339
rect 56203 10293 56358 10339
rect 56002 10245 56358 10293
rect 56002 10199 56157 10245
rect 56203 10199 56358 10245
rect 56002 10151 56358 10199
rect 56002 10105 56157 10151
rect 56203 10105 56358 10151
rect 56002 10057 56358 10105
rect 56002 10011 56157 10057
rect 56203 10011 56358 10057
rect 56002 9963 56358 10011
rect 56002 9917 56157 9963
rect 56203 9917 56358 9963
rect 56002 9869 56358 9917
rect 56002 9823 56157 9869
rect 56203 9823 56358 9869
rect 56002 9775 56358 9823
rect 56002 9729 56157 9775
rect 56203 9729 56358 9775
rect 56002 9681 56358 9729
rect 56002 9635 56157 9681
rect 56203 9635 56358 9681
rect 56002 9587 56358 9635
rect 56002 9541 56157 9587
rect 56203 9541 56358 9587
rect 56002 9493 56358 9541
rect 56002 9447 56157 9493
rect 56203 9447 56358 9493
rect 56002 9399 56358 9447
rect 56002 9353 56157 9399
rect 56203 9353 56358 9399
rect 56002 9305 56358 9353
rect 56002 9259 56157 9305
rect 56203 9259 56358 9305
rect 56002 9211 56358 9259
rect 56002 9165 56157 9211
rect 56203 9165 56358 9211
rect 56002 9117 56358 9165
rect 56002 9071 56157 9117
rect 56203 9071 56358 9117
rect 56002 9023 56358 9071
rect 56002 8977 56157 9023
rect 56203 8977 56358 9023
rect 56002 8929 56358 8977
rect 56002 8883 56157 8929
rect 56203 8883 56358 8929
rect 56002 8835 56358 8883
rect 56002 8789 56157 8835
rect 56203 8789 56358 8835
rect 56002 8741 56358 8789
rect 56002 8695 56157 8741
rect 56203 8695 56358 8741
rect 56002 8647 56358 8695
rect 56002 8601 56157 8647
rect 56203 8601 56358 8647
rect 56002 8553 56358 8601
rect 56002 8507 56157 8553
rect 56203 8507 56358 8553
rect 56002 8459 56358 8507
rect 56002 8413 56157 8459
rect 56203 8413 56358 8459
rect 56002 8365 56358 8413
rect 56002 8319 56157 8365
rect 56203 8319 56358 8365
rect 56002 8271 56358 8319
rect 56002 8225 56157 8271
rect 56203 8225 56358 8271
rect 56002 8177 56358 8225
rect 56002 8131 56157 8177
rect 56203 8131 56358 8177
rect 56002 8083 56358 8131
rect 56002 8037 56157 8083
rect 56203 8037 56358 8083
rect 56002 7989 56358 8037
rect 56002 7943 56157 7989
rect 56203 7943 56358 7989
rect 56002 7895 56358 7943
rect 56002 7849 56157 7895
rect 56203 7849 56358 7895
rect 56002 7801 56358 7849
rect 56002 7755 56157 7801
rect 56203 7755 56358 7801
rect 56002 7707 56358 7755
rect 56002 7661 56157 7707
rect 56203 7661 56358 7707
rect 56002 7613 56358 7661
rect 56002 7579 56157 7613
rect 52067 7567 56157 7579
rect 56203 7579 56358 7613
rect 56657 11676 56703 12019
rect 56657 10882 56703 11102
rect 56817 11676 56863 12019
rect 56945 11676 56991 11687
rect 56930 11270 56945 11282
rect 57105 11676 57151 12019
rect 57265 11676 57311 11687
rect 57425 11676 57471 12019
rect 56991 11270 57006 11282
rect 56930 11218 56942 11270
rect 56994 11218 57006 11270
rect 56930 11166 56945 11218
rect 56991 11166 57006 11218
rect 56930 11114 56942 11166
rect 56994 11114 57006 11166
rect 56930 11102 56945 11114
rect 56991 11102 57006 11114
rect 57249 11664 57265 11676
rect 57311 11664 57325 11676
rect 57249 11612 57261 11664
rect 57313 11612 57325 11664
rect 57249 11560 57265 11612
rect 57311 11560 57325 11612
rect 57249 11508 57261 11560
rect 57313 11508 57325 11560
rect 57249 11496 57265 11508
rect 56817 10882 56863 11102
rect 56945 11091 56991 11102
rect 56657 10836 56737 10882
rect 56783 10836 56863 10882
rect 56657 10616 56703 10836
rect 56657 9556 56703 10042
rect 56657 8762 56703 8982
rect 56817 10616 56863 10836
rect 56945 10616 56991 10627
rect 56930 10210 56945 10222
rect 57105 10616 57151 11102
rect 57311 11496 57325 11508
rect 57265 11091 57311 11102
rect 57585 11676 57631 11687
rect 57570 11270 57585 11282
rect 57745 11676 57791 12019
rect 58130 11812 58206 11824
rect 58130 11760 58142 11812
rect 58194 11809 58206 11812
rect 58290 11812 58366 11824
rect 58290 11809 58302 11812
rect 58194 11760 58302 11809
rect 58354 11760 58366 11812
rect 58130 11748 58366 11760
rect 57905 11676 57951 11687
rect 58065 11676 58111 11687
rect 57631 11270 57646 11282
rect 57570 11218 57582 11270
rect 57634 11218 57646 11270
rect 57570 11166 57585 11218
rect 57631 11166 57646 11218
rect 57570 11114 57582 11166
rect 57634 11114 57646 11166
rect 57570 11102 57585 11114
rect 57631 11102 57646 11114
rect 57889 11664 57905 11676
rect 57951 11664 57965 11676
rect 57889 11612 57901 11664
rect 57953 11612 57965 11664
rect 57889 11560 57905 11612
rect 57951 11560 57965 11612
rect 57889 11508 57901 11560
rect 57953 11508 57965 11560
rect 57889 11496 57905 11508
rect 57265 10616 57311 10627
rect 57425 10616 57471 11102
rect 57585 11091 57631 11102
rect 56991 10210 57006 10222
rect 56930 10158 56942 10210
rect 56994 10158 57006 10210
rect 56930 10106 56945 10158
rect 56991 10106 57006 10158
rect 56930 10054 56942 10106
rect 56994 10054 57006 10106
rect 56930 10042 56945 10054
rect 56991 10042 57006 10054
rect 57249 10604 57265 10616
rect 57311 10604 57325 10616
rect 57249 10552 57261 10604
rect 57313 10552 57325 10604
rect 57249 10500 57265 10552
rect 57311 10500 57325 10552
rect 57249 10448 57261 10500
rect 57313 10448 57325 10500
rect 57249 10436 57265 10448
rect 56817 9556 56863 10042
rect 56945 10031 56991 10042
rect 56945 9556 56991 9567
rect 56930 9150 56945 9162
rect 57105 9556 57151 10042
rect 57311 10436 57325 10448
rect 57265 10031 57311 10042
rect 57585 10616 57631 10627
rect 57570 10210 57585 10222
rect 57745 10616 57791 11102
rect 57951 11496 57965 11508
rect 57905 11091 57951 11102
rect 58065 11045 58111 11102
rect 58225 11676 58271 11748
rect 58225 11091 58271 11102
rect 58385 11676 58431 11687
rect 58545 11676 58591 11687
rect 58705 11676 58751 12019
rect 58529 11664 58545 11676
rect 58591 11664 58605 11676
rect 58529 11612 58541 11664
rect 58593 11612 58605 11664
rect 58529 11560 58545 11612
rect 58591 11560 58605 11612
rect 58529 11508 58541 11560
rect 58593 11508 58605 11560
rect 58529 11496 58545 11508
rect 58385 11045 58431 11102
rect 58591 11496 58605 11508
rect 58545 11091 58591 11102
rect 58865 11676 58911 11687
rect 58850 11270 58865 11282
rect 59025 11676 59071 12019
rect 59185 11676 59231 11687
rect 59345 11676 59391 12019
rect 58911 11270 58926 11282
rect 58850 11218 58862 11270
rect 58914 11218 58926 11270
rect 58850 11166 58865 11218
rect 58911 11166 58926 11218
rect 58850 11114 58862 11166
rect 58914 11114 58926 11166
rect 58850 11102 58865 11114
rect 58911 11102 58926 11114
rect 59169 11664 59185 11676
rect 59231 11664 59245 11676
rect 59169 11612 59181 11664
rect 59233 11612 59245 11664
rect 59169 11560 59185 11612
rect 59231 11560 59245 11612
rect 59169 11508 59181 11560
rect 59233 11508 59245 11560
rect 59169 11496 59185 11508
rect 58705 11045 58751 11102
rect 58865 11091 58911 11102
rect 58065 10999 58751 11045
rect 58130 10752 58206 10764
rect 58130 10700 58142 10752
rect 58194 10749 58206 10752
rect 58290 10752 58366 10764
rect 58290 10749 58302 10752
rect 58194 10700 58302 10749
rect 58354 10700 58366 10752
rect 58130 10688 58366 10700
rect 57905 10616 57951 10627
rect 58065 10616 58111 10627
rect 57631 10210 57646 10222
rect 57570 10158 57582 10210
rect 57634 10158 57646 10210
rect 57570 10106 57585 10158
rect 57631 10106 57646 10158
rect 57570 10054 57582 10106
rect 57634 10054 57646 10106
rect 57570 10042 57585 10054
rect 57631 10042 57646 10054
rect 57889 10604 57905 10616
rect 57951 10604 57965 10616
rect 57889 10552 57901 10604
rect 57953 10552 57965 10604
rect 57889 10500 57905 10552
rect 57951 10500 57965 10552
rect 57889 10448 57901 10500
rect 57953 10448 57965 10500
rect 57889 10436 57905 10448
rect 57265 9556 57311 9567
rect 57425 9556 57471 10042
rect 57585 10031 57631 10042
rect 56991 9150 57006 9162
rect 56930 9098 56942 9150
rect 56994 9098 57006 9150
rect 56930 9046 56945 9098
rect 56991 9046 57006 9098
rect 56930 8994 56942 9046
rect 56994 8994 57006 9046
rect 56930 8982 56945 8994
rect 56991 8982 57006 8994
rect 57249 9544 57265 9556
rect 57311 9544 57325 9556
rect 57249 9492 57261 9544
rect 57313 9492 57325 9544
rect 57249 9440 57265 9492
rect 57311 9440 57325 9492
rect 57249 9388 57261 9440
rect 57313 9388 57325 9440
rect 57249 9376 57265 9388
rect 56817 8762 56863 8982
rect 56945 8971 56991 8982
rect 56657 8716 56737 8762
rect 56783 8716 56863 8762
rect 56657 8496 56703 8716
rect 56657 7579 56703 7922
rect 56817 8496 56863 8716
rect 56945 8496 56991 8507
rect 56930 8090 56945 8102
rect 57105 8496 57151 8982
rect 57311 9376 57325 9388
rect 57265 8971 57311 8982
rect 57585 9556 57631 9567
rect 57570 9150 57585 9162
rect 57745 9556 57791 10042
rect 57951 10436 57965 10448
rect 57905 10031 57951 10042
rect 58065 9985 58111 10042
rect 58225 10616 58271 10688
rect 58225 10031 58271 10042
rect 58385 10616 58431 10627
rect 58545 10616 58591 10627
rect 58705 10616 58751 10999
rect 58529 10604 58545 10616
rect 58591 10604 58605 10616
rect 58529 10552 58541 10604
rect 58593 10552 58605 10604
rect 58529 10500 58545 10552
rect 58591 10500 58605 10552
rect 58529 10448 58541 10500
rect 58593 10448 58605 10500
rect 58529 10436 58545 10448
rect 58385 9985 58431 10042
rect 58591 10436 58605 10448
rect 58545 10031 58591 10042
rect 58865 10616 58911 10627
rect 58850 10210 58865 10222
rect 59025 10616 59071 11102
rect 59231 11496 59245 11508
rect 59185 11091 59231 11102
rect 59505 11676 59551 11687
rect 59490 11270 59505 11282
rect 59633 11676 59679 12019
rect 59551 11270 59566 11282
rect 59490 11218 59502 11270
rect 59554 11218 59566 11270
rect 59490 11166 59505 11218
rect 59551 11166 59566 11218
rect 59490 11114 59502 11166
rect 59554 11114 59566 11166
rect 59490 11102 59505 11114
rect 59551 11102 59566 11114
rect 59185 10616 59231 10627
rect 59345 10616 59391 11102
rect 59505 11091 59551 11102
rect 59633 10882 59679 11102
rect 59793 11676 59839 12019
rect 59793 10882 59839 11102
rect 59633 10836 59713 10882
rect 59759 10836 59839 10882
rect 58911 10210 58926 10222
rect 58850 10158 58862 10210
rect 58914 10158 58926 10210
rect 58850 10106 58865 10158
rect 58911 10106 58926 10158
rect 58850 10054 58862 10106
rect 58914 10054 58926 10106
rect 58850 10042 58865 10054
rect 58911 10042 58926 10054
rect 59169 10604 59185 10616
rect 59231 10604 59245 10616
rect 59169 10552 59181 10604
rect 59233 10552 59245 10604
rect 59169 10500 59185 10552
rect 59231 10500 59245 10552
rect 59169 10448 59181 10500
rect 59233 10448 59245 10500
rect 59169 10436 59185 10448
rect 58705 9985 58751 10042
rect 58865 10031 58911 10042
rect 58065 9939 58751 9985
rect 58130 9692 58206 9704
rect 58130 9640 58142 9692
rect 58194 9689 58206 9692
rect 58290 9692 58366 9704
rect 58290 9689 58302 9692
rect 58194 9640 58302 9689
rect 58354 9640 58366 9692
rect 58130 9628 58366 9640
rect 57905 9556 57951 9567
rect 58065 9556 58111 9567
rect 57631 9150 57646 9162
rect 57570 9098 57582 9150
rect 57634 9098 57646 9150
rect 57570 9046 57585 9098
rect 57631 9046 57646 9098
rect 57570 8994 57582 9046
rect 57634 8994 57646 9046
rect 57570 8982 57585 8994
rect 57631 8982 57646 8994
rect 57889 9544 57905 9556
rect 57951 9544 57965 9556
rect 57889 9492 57901 9544
rect 57953 9492 57965 9544
rect 57889 9440 57905 9492
rect 57951 9440 57965 9492
rect 57889 9388 57901 9440
rect 57953 9388 57965 9440
rect 57889 9376 57905 9388
rect 57265 8496 57311 8507
rect 57425 8496 57471 8982
rect 57585 8971 57631 8982
rect 56991 8090 57006 8102
rect 56930 8038 56942 8090
rect 56994 8038 57006 8090
rect 56930 7986 56945 8038
rect 56991 7986 57006 8038
rect 56930 7934 56942 7986
rect 56994 7934 57006 7986
rect 56930 7922 56945 7934
rect 56991 7922 57006 7934
rect 57249 8484 57265 8496
rect 57311 8484 57325 8496
rect 57249 8432 57261 8484
rect 57313 8432 57325 8484
rect 57249 8380 57265 8432
rect 57311 8380 57325 8432
rect 57249 8328 57261 8380
rect 57313 8328 57325 8380
rect 57249 8316 57265 8328
rect 56817 7579 56863 7922
rect 56945 7911 56991 7922
rect 57105 7579 57151 7922
rect 57311 8316 57325 8328
rect 57265 7911 57311 7922
rect 57585 8496 57631 8507
rect 57570 8090 57585 8102
rect 57745 8496 57791 8982
rect 57951 9376 57965 9388
rect 57905 8971 57951 8982
rect 58065 8925 58111 8982
rect 58225 9556 58271 9628
rect 58225 8971 58271 8982
rect 58385 9556 58431 9567
rect 58545 9556 58591 9567
rect 58705 9556 58751 9939
rect 58529 9544 58545 9556
rect 58591 9544 58605 9556
rect 58529 9492 58541 9544
rect 58593 9492 58605 9544
rect 58529 9440 58545 9492
rect 58591 9440 58605 9492
rect 58529 9388 58541 9440
rect 58593 9388 58605 9440
rect 58529 9376 58545 9388
rect 58385 8925 58431 8982
rect 58591 9376 58605 9388
rect 58545 8971 58591 8982
rect 58865 9556 58911 9567
rect 58850 9150 58865 9162
rect 59025 9556 59071 10042
rect 59231 10436 59245 10448
rect 59185 10031 59231 10042
rect 59505 10616 59551 10627
rect 59490 10210 59505 10222
rect 59633 10616 59679 10836
rect 59551 10210 59566 10222
rect 59490 10158 59502 10210
rect 59554 10158 59566 10210
rect 59490 10106 59505 10158
rect 59551 10106 59566 10158
rect 59490 10054 59502 10106
rect 59554 10054 59566 10106
rect 59490 10042 59505 10054
rect 59551 10042 59566 10054
rect 59185 9556 59231 9567
rect 59345 9556 59391 10042
rect 59505 10031 59551 10042
rect 58911 9150 58926 9162
rect 58850 9098 58862 9150
rect 58914 9098 58926 9150
rect 58850 9046 58865 9098
rect 58911 9046 58926 9098
rect 58850 8994 58862 9046
rect 58914 8994 58926 9046
rect 58850 8982 58865 8994
rect 58911 8982 58926 8994
rect 59169 9544 59185 9556
rect 59231 9544 59245 9556
rect 59169 9492 59181 9544
rect 59233 9492 59245 9544
rect 59169 9440 59185 9492
rect 59231 9440 59245 9492
rect 59169 9388 59181 9440
rect 59233 9388 59245 9440
rect 59169 9376 59185 9388
rect 58705 8925 58751 8982
rect 58865 8971 58911 8982
rect 58065 8879 58751 8925
rect 58130 8632 58206 8644
rect 58130 8580 58142 8632
rect 58194 8629 58206 8632
rect 58290 8632 58366 8644
rect 58290 8629 58302 8632
rect 58194 8580 58302 8629
rect 58354 8580 58366 8632
rect 58130 8568 58366 8580
rect 57905 8496 57951 8507
rect 58065 8496 58111 8507
rect 57631 8090 57646 8102
rect 57570 8038 57582 8090
rect 57634 8038 57646 8090
rect 57570 7986 57585 8038
rect 57631 7986 57646 8038
rect 57570 7934 57582 7986
rect 57634 7934 57646 7986
rect 57570 7922 57585 7934
rect 57631 7922 57646 7934
rect 57889 8484 57905 8496
rect 57951 8484 57965 8496
rect 57889 8432 57901 8484
rect 57953 8432 57965 8484
rect 57889 8380 57905 8432
rect 57951 8380 57965 8432
rect 57889 8328 57901 8380
rect 57953 8328 57965 8380
rect 57889 8316 57905 8328
rect 57425 7579 57471 7922
rect 57585 7911 57631 7922
rect 57745 7579 57791 7922
rect 57951 8316 57965 8328
rect 57905 7911 57951 7922
rect 58065 7579 58111 7922
rect 58225 8496 58271 8568
rect 58225 7911 58271 7922
rect 58385 8496 58431 8507
rect 58545 8496 58591 8507
rect 58705 8496 58751 8879
rect 58529 8484 58545 8496
rect 58591 8484 58605 8496
rect 58529 8432 58541 8484
rect 58593 8432 58605 8484
rect 58529 8380 58545 8432
rect 58591 8380 58605 8432
rect 58529 8328 58541 8380
rect 58593 8328 58605 8380
rect 58529 8316 58545 8328
rect 58385 7579 58431 7922
rect 58591 8316 58605 8328
rect 58545 7911 58591 7922
rect 58865 8496 58911 8507
rect 58850 8090 58865 8102
rect 59025 8496 59071 8982
rect 59231 9376 59245 9388
rect 59185 8971 59231 8982
rect 59505 9556 59551 9567
rect 59490 9150 59505 9162
rect 59633 9556 59679 10042
rect 59551 9150 59566 9162
rect 59490 9098 59502 9150
rect 59554 9098 59566 9150
rect 59490 9046 59505 9098
rect 59551 9046 59566 9098
rect 59490 8994 59502 9046
rect 59554 8994 59566 9046
rect 59490 8982 59505 8994
rect 59551 8982 59566 8994
rect 59185 8496 59231 8507
rect 59345 8496 59391 8982
rect 59505 8971 59551 8982
rect 59633 8762 59679 8982
rect 59793 10616 59839 10836
rect 59793 9556 59839 10042
rect 59793 8762 59839 8982
rect 59633 8716 59713 8762
rect 59759 8716 59839 8762
rect 58911 8090 58926 8102
rect 58850 8038 58862 8090
rect 58914 8038 58926 8090
rect 58850 7986 58865 8038
rect 58911 7986 58926 8038
rect 58850 7934 58862 7986
rect 58914 7934 58926 7986
rect 58850 7922 58865 7934
rect 58911 7922 58926 7934
rect 59169 8484 59185 8496
rect 59231 8484 59245 8496
rect 59169 8432 59181 8484
rect 59233 8432 59245 8484
rect 59169 8380 59185 8432
rect 59231 8380 59245 8432
rect 59169 8328 59181 8380
rect 59233 8328 59245 8380
rect 59169 8316 59185 8328
rect 58705 7579 58751 7922
rect 58865 7911 58911 7922
rect 59025 7579 59071 7922
rect 59231 8316 59245 8328
rect 59185 7911 59231 7922
rect 59505 8496 59551 8507
rect 59490 8090 59505 8102
rect 59633 8496 59679 8716
rect 59551 8090 59566 8102
rect 59490 8038 59502 8090
rect 59554 8038 59566 8090
rect 59490 7986 59505 8038
rect 59551 7986 59566 8038
rect 59490 7934 59502 7986
rect 59554 7934 59566 7986
rect 59490 7922 59505 7934
rect 59551 7922 59566 7934
rect 59345 7579 59391 7922
rect 59505 7911 59551 7922
rect 59633 7579 59679 7922
rect 59793 8496 59839 8716
rect 59793 7579 59839 7922
rect 60138 11985 60293 12019
rect 60339 12019 61717 12031
rect 60339 11985 60458 12019
rect 60138 11937 60458 11985
rect 60138 11891 60293 11937
rect 60339 11891 60458 11937
rect 60138 11843 60458 11891
rect 60138 11797 60293 11843
rect 60339 11797 60458 11843
rect 60138 11749 60458 11797
rect 60138 11703 60293 11749
rect 60339 11703 60458 11749
rect 60138 11655 60458 11703
rect 60138 11609 60293 11655
rect 60339 11609 60458 11655
rect 60138 11561 60458 11609
rect 60138 11515 60293 11561
rect 60339 11515 60458 11561
rect 60138 11467 60458 11515
rect 60138 11421 60293 11467
rect 60339 11421 60458 11467
rect 60138 11373 60458 11421
rect 60138 11327 60293 11373
rect 60339 11327 60458 11373
rect 60138 11279 60458 11327
rect 60138 11233 60293 11279
rect 60339 11233 60458 11279
rect 60138 11185 60458 11233
rect 60138 11139 60293 11185
rect 60339 11139 60458 11185
rect 60138 11091 60458 11139
rect 60138 11045 60293 11091
rect 60339 11045 60458 11091
rect 60138 10997 60458 11045
rect 60138 10951 60293 10997
rect 60339 10951 60458 10997
rect 60138 10903 60458 10951
rect 60138 10857 60293 10903
rect 60339 10857 60458 10903
rect 60138 10809 60458 10857
rect 60138 10763 60293 10809
rect 60339 10763 60458 10809
rect 60138 10715 60458 10763
rect 60138 10669 60293 10715
rect 60339 10669 60458 10715
rect 60138 10621 60458 10669
rect 60138 10575 60293 10621
rect 60339 10575 60458 10621
rect 60138 10527 60458 10575
rect 60138 10481 60293 10527
rect 60339 10481 60458 10527
rect 60138 10433 60458 10481
rect 60138 10387 60293 10433
rect 60339 10387 60458 10433
rect 60138 10339 60458 10387
rect 60138 10293 60293 10339
rect 60339 10293 60458 10339
rect 60138 10245 60458 10293
rect 60138 10199 60293 10245
rect 60339 10199 60458 10245
rect 60138 10151 60458 10199
rect 60138 10105 60293 10151
rect 60339 10105 60458 10151
rect 60138 10057 60458 10105
rect 60138 10011 60293 10057
rect 60339 10011 60458 10057
rect 60138 9963 60458 10011
rect 60138 9917 60293 9963
rect 60339 9917 60458 9963
rect 60138 9869 60458 9917
rect 60138 9823 60293 9869
rect 60339 9823 60458 9869
rect 60138 9775 60458 9823
rect 60138 9729 60293 9775
rect 60339 9729 60458 9775
rect 60138 9681 60458 9729
rect 60138 9635 60293 9681
rect 60339 9635 60458 9681
rect 60138 9587 60458 9635
rect 60138 9541 60293 9587
rect 60339 9541 60458 9587
rect 60138 9493 60458 9541
rect 60138 9447 60293 9493
rect 60339 9447 60458 9493
rect 60138 9399 60458 9447
rect 60138 9353 60293 9399
rect 60339 9353 60458 9399
rect 60138 9305 60458 9353
rect 60138 9259 60293 9305
rect 60339 9259 60458 9305
rect 60138 9211 60458 9259
rect 60138 9165 60293 9211
rect 60339 9165 60458 9211
rect 60138 9117 60458 9165
rect 60138 9071 60293 9117
rect 60339 9071 60458 9117
rect 60138 9023 60458 9071
rect 60138 8977 60293 9023
rect 60339 8977 60458 9023
rect 60138 8929 60458 8977
rect 60138 8883 60293 8929
rect 60339 8883 60458 8929
rect 60138 8835 60458 8883
rect 60138 8789 60293 8835
rect 60339 8789 60458 8835
rect 60138 8741 60458 8789
rect 60138 8695 60293 8741
rect 60339 8695 60458 8741
rect 60138 8647 60458 8695
rect 60138 8601 60293 8647
rect 60339 8601 60458 8647
rect 60138 8553 60458 8601
rect 60138 8507 60293 8553
rect 60339 8507 60458 8553
rect 60138 8459 60458 8507
rect 60138 8413 60293 8459
rect 60339 8413 60458 8459
rect 60138 8365 60458 8413
rect 60138 8319 60293 8365
rect 60339 8319 60458 8365
rect 60138 8271 60458 8319
rect 60138 8225 60293 8271
rect 60339 8225 60458 8271
rect 60138 8177 60458 8225
rect 60138 8131 60293 8177
rect 60339 8131 60458 8177
rect 60138 8083 60458 8131
rect 60138 8037 60293 8083
rect 60339 8037 60458 8083
rect 60138 7989 60458 8037
rect 60138 7943 60293 7989
rect 60339 7943 60458 7989
rect 60138 7895 60458 7943
rect 60138 7849 60293 7895
rect 60339 7849 60458 7895
rect 60138 7801 60458 7849
rect 60138 7755 60293 7801
rect 60339 7755 60458 7801
rect 60138 7707 60458 7755
rect 60138 7661 60293 7707
rect 60339 7661 60458 7707
rect 60138 7613 60458 7661
rect 60138 7579 60293 7613
rect 56203 7567 60293 7579
rect 60339 7579 60458 7613
rect 61598 11985 61717 12019
rect 61763 12019 65853 12031
rect 61763 11985 61918 12019
rect 61598 11937 61918 11985
rect 61598 11891 61717 11937
rect 61763 11891 61918 11937
rect 61598 11843 61918 11891
rect 61598 11797 61717 11843
rect 61763 11797 61918 11843
rect 61598 11749 61918 11797
rect 61598 11703 61717 11749
rect 61763 11703 61918 11749
rect 61598 11655 61918 11703
rect 61598 11609 61717 11655
rect 61763 11609 61918 11655
rect 61598 11561 61918 11609
rect 61598 11515 61717 11561
rect 61763 11515 61918 11561
rect 61598 11467 61918 11515
rect 61598 11421 61717 11467
rect 61763 11421 61918 11467
rect 61598 11373 61918 11421
rect 61598 11327 61717 11373
rect 61763 11327 61918 11373
rect 61598 11279 61918 11327
rect 61598 11233 61717 11279
rect 61763 11233 61918 11279
rect 61598 11185 61918 11233
rect 61598 11139 61717 11185
rect 61763 11139 61918 11185
rect 61598 11091 61918 11139
rect 61598 11045 61717 11091
rect 61763 11045 61918 11091
rect 61598 10997 61918 11045
rect 61598 10951 61717 10997
rect 61763 10951 61918 10997
rect 61598 10903 61918 10951
rect 61598 10857 61717 10903
rect 61763 10857 61918 10903
rect 61598 10809 61918 10857
rect 61598 10763 61717 10809
rect 61763 10763 61918 10809
rect 61598 10715 61918 10763
rect 61598 10669 61717 10715
rect 61763 10669 61918 10715
rect 61598 10621 61918 10669
rect 61598 10575 61717 10621
rect 61763 10575 61918 10621
rect 61598 10527 61918 10575
rect 61598 10481 61717 10527
rect 61763 10481 61918 10527
rect 61598 10433 61918 10481
rect 61598 10387 61717 10433
rect 61763 10387 61918 10433
rect 61598 10339 61918 10387
rect 61598 10293 61717 10339
rect 61763 10293 61918 10339
rect 61598 10245 61918 10293
rect 61598 10199 61717 10245
rect 61763 10199 61918 10245
rect 61598 10151 61918 10199
rect 61598 10105 61717 10151
rect 61763 10105 61918 10151
rect 61598 10057 61918 10105
rect 61598 10011 61717 10057
rect 61763 10011 61918 10057
rect 61598 9963 61918 10011
rect 61598 9917 61717 9963
rect 61763 9917 61918 9963
rect 61598 9869 61918 9917
rect 61598 9823 61717 9869
rect 61763 9823 61918 9869
rect 61598 9775 61918 9823
rect 61598 9729 61717 9775
rect 61763 9729 61918 9775
rect 61598 9681 61918 9729
rect 61598 9635 61717 9681
rect 61763 9635 61918 9681
rect 61598 9587 61918 9635
rect 61598 9541 61717 9587
rect 61763 9541 61918 9587
rect 61598 9493 61918 9541
rect 61598 9447 61717 9493
rect 61763 9447 61918 9493
rect 61598 9399 61918 9447
rect 61598 9353 61717 9399
rect 61763 9353 61918 9399
rect 61598 9305 61918 9353
rect 61598 9259 61717 9305
rect 61763 9259 61918 9305
rect 61598 9211 61918 9259
rect 61598 9165 61717 9211
rect 61763 9165 61918 9211
rect 61598 9117 61918 9165
rect 61598 9071 61717 9117
rect 61763 9071 61918 9117
rect 61598 9023 61918 9071
rect 61598 8977 61717 9023
rect 61763 8977 61918 9023
rect 61598 8929 61918 8977
rect 61598 8883 61717 8929
rect 61763 8883 61918 8929
rect 61598 8835 61918 8883
rect 61598 8789 61717 8835
rect 61763 8789 61918 8835
rect 61598 8741 61918 8789
rect 61598 8695 61717 8741
rect 61763 8695 61918 8741
rect 61598 8647 61918 8695
rect 61598 8601 61717 8647
rect 61763 8601 61918 8647
rect 61598 8553 61918 8601
rect 61598 8507 61717 8553
rect 61763 8507 61918 8553
rect 61598 8459 61918 8507
rect 61598 8413 61717 8459
rect 61763 8413 61918 8459
rect 61598 8365 61918 8413
rect 61598 8319 61717 8365
rect 61763 8319 61918 8365
rect 61598 8271 61918 8319
rect 61598 8225 61717 8271
rect 61763 8225 61918 8271
rect 61598 8177 61918 8225
rect 61598 8131 61717 8177
rect 61763 8131 61918 8177
rect 61598 8083 61918 8131
rect 61598 8037 61717 8083
rect 61763 8037 61918 8083
rect 61598 7989 61918 8037
rect 61598 7943 61717 7989
rect 61763 7943 61918 7989
rect 61598 7895 61918 7943
rect 61598 7849 61717 7895
rect 61763 7849 61918 7895
rect 61598 7801 61918 7849
rect 61598 7755 61717 7801
rect 61763 7755 61918 7801
rect 61598 7707 61918 7755
rect 61598 7661 61717 7707
rect 61763 7661 61918 7707
rect 61598 7613 61918 7661
rect 61598 7579 61717 7613
rect 60339 7567 61717 7579
rect 61763 7579 61918 7613
rect 62217 11676 62263 12019
rect 62217 10882 62263 11102
rect 62377 11676 62423 12019
rect 62505 11676 62551 11687
rect 62490 11270 62505 11282
rect 62665 11676 62711 12019
rect 62825 11676 62871 11687
rect 62985 11676 63031 12019
rect 62551 11270 62566 11282
rect 62490 11218 62502 11270
rect 62554 11218 62566 11270
rect 62490 11166 62505 11218
rect 62551 11166 62566 11218
rect 62490 11114 62502 11166
rect 62554 11114 62566 11166
rect 62490 11102 62505 11114
rect 62551 11102 62566 11114
rect 62811 11664 62825 11676
rect 62871 11664 62887 11676
rect 62811 11612 62823 11664
rect 62875 11612 62887 11664
rect 62811 11560 62825 11612
rect 62871 11560 62887 11612
rect 62811 11508 62823 11560
rect 62875 11508 62887 11560
rect 62811 11496 62825 11508
rect 62377 10882 62423 11102
rect 62505 11091 62551 11102
rect 62217 10836 62297 10882
rect 62343 10836 62423 10882
rect 62217 10616 62263 10836
rect 62217 9556 62263 10042
rect 62217 8762 62263 8982
rect 62377 10616 62423 10836
rect 62505 10616 62551 10627
rect 62490 10210 62505 10222
rect 62665 10616 62711 11102
rect 62871 11496 62887 11508
rect 62825 11091 62871 11102
rect 63145 11676 63191 11687
rect 63130 11270 63145 11282
rect 63305 11676 63351 12019
rect 63690 11812 63766 11824
rect 63690 11760 63702 11812
rect 63754 11809 63766 11812
rect 63850 11812 63926 11824
rect 63850 11809 63862 11812
rect 63754 11760 63862 11809
rect 63914 11760 63926 11812
rect 63690 11748 63926 11760
rect 63465 11676 63511 11687
rect 63625 11676 63671 11687
rect 63191 11270 63206 11282
rect 63130 11218 63142 11270
rect 63194 11218 63206 11270
rect 63130 11166 63145 11218
rect 63191 11166 63206 11218
rect 63130 11114 63142 11166
rect 63194 11114 63206 11166
rect 63130 11102 63145 11114
rect 63191 11102 63206 11114
rect 63451 11664 63465 11676
rect 63511 11664 63527 11676
rect 63451 11612 63463 11664
rect 63515 11612 63527 11664
rect 63451 11560 63465 11612
rect 63511 11560 63527 11612
rect 63451 11508 63463 11560
rect 63515 11508 63527 11560
rect 63451 11496 63465 11508
rect 62825 10616 62871 10627
rect 62985 10616 63031 11102
rect 63145 11091 63191 11102
rect 63305 11045 63351 11102
rect 63511 11496 63527 11508
rect 63465 11091 63511 11102
rect 63625 11045 63671 11102
rect 63785 11676 63831 11748
rect 63785 11091 63831 11102
rect 63945 11676 63991 11687
rect 64105 11676 64151 11687
rect 64265 11676 64311 12019
rect 64091 11664 64105 11676
rect 64151 11664 64167 11676
rect 64091 11612 64103 11664
rect 64155 11612 64167 11664
rect 64091 11560 64105 11612
rect 64151 11560 64167 11612
rect 64091 11508 64103 11560
rect 64155 11508 64167 11560
rect 64091 11496 64105 11508
rect 63945 11045 63991 11102
rect 64151 11496 64167 11508
rect 64105 11091 64151 11102
rect 64425 11676 64471 11687
rect 64410 11270 64425 11282
rect 64585 11676 64631 12019
rect 64745 11676 64791 11687
rect 64905 11676 64951 12019
rect 64471 11270 64486 11282
rect 64410 11218 64422 11270
rect 64474 11218 64486 11270
rect 64410 11166 64425 11218
rect 64471 11166 64486 11218
rect 64410 11114 64422 11166
rect 64474 11114 64486 11166
rect 64410 11102 64425 11114
rect 64471 11102 64486 11114
rect 64731 11664 64745 11676
rect 64791 11664 64807 11676
rect 64731 11612 64743 11664
rect 64795 11612 64807 11664
rect 64731 11560 64745 11612
rect 64791 11560 64807 11612
rect 64731 11508 64743 11560
rect 64795 11508 64807 11560
rect 64731 11496 64745 11508
rect 63305 10999 63991 11045
rect 62551 10210 62566 10222
rect 62490 10158 62502 10210
rect 62554 10158 62566 10210
rect 62490 10106 62505 10158
rect 62551 10106 62566 10158
rect 62490 10054 62502 10106
rect 62554 10054 62566 10106
rect 62490 10042 62505 10054
rect 62551 10042 62566 10054
rect 62811 10604 62825 10616
rect 62871 10604 62887 10616
rect 62811 10552 62823 10604
rect 62875 10552 62887 10604
rect 62811 10500 62825 10552
rect 62871 10500 62887 10552
rect 62811 10448 62823 10500
rect 62875 10448 62887 10500
rect 62811 10436 62825 10448
rect 62377 9556 62423 10042
rect 62505 10031 62551 10042
rect 62505 9556 62551 9567
rect 62490 9150 62505 9162
rect 62665 9556 62711 10042
rect 62871 10436 62887 10448
rect 62825 10031 62871 10042
rect 63145 10616 63191 10627
rect 63130 10210 63145 10222
rect 63305 10616 63351 10999
rect 63690 10752 63766 10764
rect 63690 10700 63702 10752
rect 63754 10749 63766 10752
rect 63850 10752 63926 10764
rect 63850 10749 63862 10752
rect 63754 10700 63862 10749
rect 63914 10700 63926 10752
rect 63690 10688 63926 10700
rect 63465 10616 63511 10627
rect 63625 10616 63671 10627
rect 63191 10210 63206 10222
rect 63130 10158 63142 10210
rect 63194 10158 63206 10210
rect 63130 10106 63145 10158
rect 63191 10106 63206 10158
rect 63130 10054 63142 10106
rect 63194 10054 63206 10106
rect 63130 10042 63145 10054
rect 63191 10042 63206 10054
rect 63451 10604 63465 10616
rect 63511 10604 63527 10616
rect 63451 10552 63463 10604
rect 63515 10552 63527 10604
rect 63451 10500 63465 10552
rect 63511 10500 63527 10552
rect 63451 10448 63463 10500
rect 63515 10448 63527 10500
rect 63451 10436 63465 10448
rect 62825 9556 62871 9567
rect 62985 9556 63031 10042
rect 63145 10031 63191 10042
rect 63305 9985 63351 10042
rect 63511 10436 63527 10448
rect 63465 10031 63511 10042
rect 63625 9985 63671 10042
rect 63785 10616 63831 10688
rect 63785 10031 63831 10042
rect 63945 10616 63991 10627
rect 64105 10616 64151 10627
rect 64265 10616 64311 11102
rect 64425 11091 64471 11102
rect 64091 10604 64105 10616
rect 64151 10604 64167 10616
rect 64091 10552 64103 10604
rect 64155 10552 64167 10604
rect 64091 10500 64105 10552
rect 64151 10500 64167 10552
rect 64091 10448 64103 10500
rect 64155 10448 64167 10500
rect 64091 10436 64105 10448
rect 63945 9985 63991 10042
rect 64151 10436 64167 10448
rect 64105 10031 64151 10042
rect 64425 10616 64471 10627
rect 64410 10210 64425 10222
rect 64585 10616 64631 11102
rect 64791 11496 64807 11508
rect 64745 11091 64791 11102
rect 65065 11676 65111 11687
rect 65050 11270 65065 11282
rect 65193 11676 65239 12019
rect 65111 11270 65126 11282
rect 65050 11218 65062 11270
rect 65114 11218 65126 11270
rect 65050 11166 65065 11218
rect 65111 11166 65126 11218
rect 65050 11114 65062 11166
rect 65114 11114 65126 11166
rect 65050 11102 65065 11114
rect 65111 11102 65126 11114
rect 64745 10616 64791 10627
rect 64905 10616 64951 11102
rect 65065 11091 65111 11102
rect 65193 10882 65239 11102
rect 65353 11676 65399 12019
rect 65353 10882 65399 11102
rect 65193 10836 65273 10882
rect 65319 10836 65399 10882
rect 64471 10210 64486 10222
rect 64410 10158 64422 10210
rect 64474 10158 64486 10210
rect 64410 10106 64425 10158
rect 64471 10106 64486 10158
rect 64410 10054 64422 10106
rect 64474 10054 64486 10106
rect 64410 10042 64425 10054
rect 64471 10042 64486 10054
rect 64731 10604 64745 10616
rect 64791 10604 64807 10616
rect 64731 10552 64743 10604
rect 64795 10552 64807 10604
rect 64731 10500 64745 10552
rect 64791 10500 64807 10552
rect 64731 10448 64743 10500
rect 64795 10448 64807 10500
rect 64731 10436 64745 10448
rect 63305 9939 63991 9985
rect 62551 9150 62566 9162
rect 62490 9098 62502 9150
rect 62554 9098 62566 9150
rect 62490 9046 62505 9098
rect 62551 9046 62566 9098
rect 62490 8994 62502 9046
rect 62554 8994 62566 9046
rect 62490 8982 62505 8994
rect 62551 8982 62566 8994
rect 62811 9544 62825 9556
rect 62871 9544 62887 9556
rect 62811 9492 62823 9544
rect 62875 9492 62887 9544
rect 62811 9440 62825 9492
rect 62871 9440 62887 9492
rect 62811 9388 62823 9440
rect 62875 9388 62887 9440
rect 62811 9376 62825 9388
rect 62377 8762 62423 8982
rect 62505 8971 62551 8982
rect 62217 8716 62297 8762
rect 62343 8716 62423 8762
rect 62217 8496 62263 8716
rect 62217 7579 62263 7922
rect 62377 8496 62423 8716
rect 62505 8496 62551 8507
rect 62490 8090 62505 8102
rect 62665 8496 62711 8982
rect 62871 9376 62887 9388
rect 62825 8971 62871 8982
rect 63145 9556 63191 9567
rect 63130 9150 63145 9162
rect 63305 9556 63351 9939
rect 63690 9692 63766 9704
rect 63690 9640 63702 9692
rect 63754 9689 63766 9692
rect 63850 9692 63926 9704
rect 63850 9689 63862 9692
rect 63754 9640 63862 9689
rect 63914 9640 63926 9692
rect 63690 9628 63926 9640
rect 63465 9556 63511 9567
rect 63625 9556 63671 9567
rect 63191 9150 63206 9162
rect 63130 9098 63142 9150
rect 63194 9098 63206 9150
rect 63130 9046 63145 9098
rect 63191 9046 63206 9098
rect 63130 8994 63142 9046
rect 63194 8994 63206 9046
rect 63130 8982 63145 8994
rect 63191 8982 63206 8994
rect 63451 9544 63465 9556
rect 63511 9544 63527 9556
rect 63451 9492 63463 9544
rect 63515 9492 63527 9544
rect 63451 9440 63465 9492
rect 63511 9440 63527 9492
rect 63451 9388 63463 9440
rect 63515 9388 63527 9440
rect 63451 9376 63465 9388
rect 62825 8496 62871 8507
rect 62985 8496 63031 8982
rect 63145 8971 63191 8982
rect 63305 8925 63351 8982
rect 63511 9376 63527 9388
rect 63465 8971 63511 8982
rect 63625 8925 63671 8982
rect 63785 9556 63831 9628
rect 63785 8971 63831 8982
rect 63945 9556 63991 9567
rect 64105 9556 64151 9567
rect 64265 9556 64311 10042
rect 64425 10031 64471 10042
rect 64091 9544 64105 9556
rect 64151 9544 64167 9556
rect 64091 9492 64103 9544
rect 64155 9492 64167 9544
rect 64091 9440 64105 9492
rect 64151 9440 64167 9492
rect 64091 9388 64103 9440
rect 64155 9388 64167 9440
rect 64091 9376 64105 9388
rect 63945 8925 63991 8982
rect 64151 9376 64167 9388
rect 64105 8971 64151 8982
rect 64425 9556 64471 9567
rect 64410 9150 64425 9162
rect 64585 9556 64631 10042
rect 64791 10436 64807 10448
rect 64745 10031 64791 10042
rect 65065 10616 65111 10627
rect 65050 10210 65065 10222
rect 65193 10616 65239 10836
rect 65111 10210 65126 10222
rect 65050 10158 65062 10210
rect 65114 10158 65126 10210
rect 65050 10106 65065 10158
rect 65111 10106 65126 10158
rect 65050 10054 65062 10106
rect 65114 10054 65126 10106
rect 65050 10042 65065 10054
rect 65111 10042 65126 10054
rect 64745 9556 64791 9567
rect 64905 9556 64951 10042
rect 65065 10031 65111 10042
rect 64471 9150 64486 9162
rect 64410 9098 64422 9150
rect 64474 9098 64486 9150
rect 64410 9046 64425 9098
rect 64471 9046 64486 9098
rect 64410 8994 64422 9046
rect 64474 8994 64486 9046
rect 64410 8982 64425 8994
rect 64471 8982 64486 8994
rect 64731 9544 64745 9556
rect 64791 9544 64807 9556
rect 64731 9492 64743 9544
rect 64795 9492 64807 9544
rect 64731 9440 64745 9492
rect 64791 9440 64807 9492
rect 64731 9388 64743 9440
rect 64795 9388 64807 9440
rect 64731 9376 64745 9388
rect 63305 8879 63991 8925
rect 62551 8090 62566 8102
rect 62490 8038 62502 8090
rect 62554 8038 62566 8090
rect 62490 7986 62505 8038
rect 62551 7986 62566 8038
rect 62490 7934 62502 7986
rect 62554 7934 62566 7986
rect 62490 7922 62505 7934
rect 62551 7922 62566 7934
rect 62811 8484 62825 8496
rect 62871 8484 62887 8496
rect 62811 8432 62823 8484
rect 62875 8432 62887 8484
rect 62811 8380 62825 8432
rect 62871 8380 62887 8432
rect 62811 8328 62823 8380
rect 62875 8328 62887 8380
rect 62811 8316 62825 8328
rect 62377 7579 62423 7922
rect 62505 7911 62551 7922
rect 62665 7579 62711 7922
rect 62871 8316 62887 8328
rect 62825 7911 62871 7922
rect 63145 8496 63191 8507
rect 63130 8090 63145 8102
rect 63305 8496 63351 8879
rect 63690 8632 63766 8644
rect 63690 8580 63702 8632
rect 63754 8629 63766 8632
rect 63850 8632 63926 8644
rect 63850 8629 63862 8632
rect 63754 8580 63862 8629
rect 63914 8580 63926 8632
rect 63690 8568 63926 8580
rect 63465 8496 63511 8507
rect 63625 8496 63671 8507
rect 63191 8090 63206 8102
rect 63130 8038 63142 8090
rect 63194 8038 63206 8090
rect 63130 7986 63145 8038
rect 63191 7986 63206 8038
rect 63130 7934 63142 7986
rect 63194 7934 63206 7986
rect 63130 7922 63145 7934
rect 63191 7922 63206 7934
rect 63451 8484 63465 8496
rect 63511 8484 63527 8496
rect 63451 8432 63463 8484
rect 63515 8432 63527 8484
rect 63451 8380 63465 8432
rect 63511 8380 63527 8432
rect 63451 8328 63463 8380
rect 63515 8328 63527 8380
rect 63451 8316 63465 8328
rect 62985 7579 63031 7922
rect 63145 7911 63191 7922
rect 63305 7579 63351 7922
rect 63511 8316 63527 8328
rect 63465 7911 63511 7922
rect 63625 7579 63671 7922
rect 63785 8496 63831 8568
rect 63785 7911 63831 7922
rect 63945 8496 63991 8507
rect 64105 8496 64151 8507
rect 64265 8496 64311 8982
rect 64425 8971 64471 8982
rect 64091 8484 64105 8496
rect 64151 8484 64167 8496
rect 64091 8432 64103 8484
rect 64155 8432 64167 8484
rect 64091 8380 64105 8432
rect 64151 8380 64167 8432
rect 64091 8328 64103 8380
rect 64155 8328 64167 8380
rect 64091 8316 64105 8328
rect 63945 7579 63991 7922
rect 64151 8316 64167 8328
rect 64105 7911 64151 7922
rect 64425 8496 64471 8507
rect 64410 8090 64425 8102
rect 64585 8496 64631 8982
rect 64791 9376 64807 9388
rect 64745 8971 64791 8982
rect 65065 9556 65111 9567
rect 65050 9150 65065 9162
rect 65193 9556 65239 10042
rect 65111 9150 65126 9162
rect 65050 9098 65062 9150
rect 65114 9098 65126 9150
rect 65050 9046 65065 9098
rect 65111 9046 65126 9098
rect 65050 8994 65062 9046
rect 65114 8994 65126 9046
rect 65050 8982 65065 8994
rect 65111 8982 65126 8994
rect 64745 8496 64791 8507
rect 64905 8496 64951 8982
rect 65065 8971 65111 8982
rect 65193 8762 65239 8982
rect 65353 10616 65399 10836
rect 65353 9556 65399 10042
rect 65353 8762 65399 8982
rect 65193 8716 65273 8762
rect 65319 8716 65399 8762
rect 64471 8090 64486 8102
rect 64410 8038 64422 8090
rect 64474 8038 64486 8090
rect 64410 7986 64425 8038
rect 64471 7986 64486 8038
rect 64410 7934 64422 7986
rect 64474 7934 64486 7986
rect 64410 7922 64425 7934
rect 64471 7922 64486 7934
rect 64731 8484 64745 8496
rect 64791 8484 64807 8496
rect 64731 8432 64743 8484
rect 64795 8432 64807 8484
rect 64731 8380 64745 8432
rect 64791 8380 64807 8432
rect 64731 8328 64743 8380
rect 64795 8328 64807 8380
rect 64731 8316 64745 8328
rect 64265 7579 64311 7922
rect 64425 7911 64471 7922
rect 64585 7579 64631 7922
rect 64791 8316 64807 8328
rect 64745 7911 64791 7922
rect 65065 8496 65111 8507
rect 65050 8090 65065 8102
rect 65193 8496 65239 8716
rect 65111 8090 65126 8102
rect 65050 8038 65062 8090
rect 65114 8038 65126 8090
rect 65050 7986 65065 8038
rect 65111 7986 65126 8038
rect 65050 7934 65062 7986
rect 65114 7934 65126 7986
rect 65050 7922 65065 7934
rect 65111 7922 65126 7934
rect 64905 7579 64951 7922
rect 65065 7911 65111 7922
rect 65193 7579 65239 7922
rect 65353 8496 65399 8716
rect 65353 7579 65399 7922
rect 65698 11985 65853 12019
rect 65899 11985 66018 12031
rect 65698 11937 66018 11985
rect 65698 11891 65853 11937
rect 65899 11891 66018 11937
rect 65698 11843 66018 11891
rect 65698 11797 65853 11843
rect 65899 11797 66018 11843
rect 65698 11749 66018 11797
rect 65698 11703 65853 11749
rect 65899 11703 66018 11749
rect 65698 11655 66018 11703
rect 65698 11609 65853 11655
rect 65899 11609 66018 11655
rect 65698 11561 66018 11609
rect 65698 11515 65853 11561
rect 65899 11515 66018 11561
rect 65698 11467 66018 11515
rect 65698 11421 65853 11467
rect 65899 11421 66018 11467
rect 65698 11373 66018 11421
rect 65698 11327 65853 11373
rect 65899 11327 66018 11373
rect 65698 11279 66018 11327
rect 65698 11233 65853 11279
rect 65899 11233 66018 11279
rect 65698 11185 66018 11233
rect 65698 11139 65853 11185
rect 65899 11139 66018 11185
rect 65698 11091 66018 11139
rect 65698 11045 65853 11091
rect 65899 11045 66018 11091
rect 65698 10997 66018 11045
rect 65698 10951 65853 10997
rect 65899 10951 66018 10997
rect 65698 10903 66018 10951
rect 65698 10857 65853 10903
rect 65899 10857 66018 10903
rect 65698 10809 66018 10857
rect 65698 10763 65853 10809
rect 65899 10763 66018 10809
rect 65698 10715 66018 10763
rect 65698 10669 65853 10715
rect 65899 10669 66018 10715
rect 65698 10621 66018 10669
rect 65698 10575 65853 10621
rect 65899 10575 66018 10621
rect 65698 10527 66018 10575
rect 65698 10481 65853 10527
rect 65899 10481 66018 10527
rect 65698 10433 66018 10481
rect 65698 10387 65853 10433
rect 65899 10387 66018 10433
rect 65698 10339 66018 10387
rect 65698 10293 65853 10339
rect 65899 10293 66018 10339
rect 65698 10245 66018 10293
rect 65698 10199 65853 10245
rect 65899 10199 66018 10245
rect 65698 10151 66018 10199
rect 65698 10105 65853 10151
rect 65899 10105 66018 10151
rect 65698 10057 66018 10105
rect 65698 10011 65853 10057
rect 65899 10011 66018 10057
rect 65698 9963 66018 10011
rect 65698 9917 65853 9963
rect 65899 9917 66018 9963
rect 65698 9869 66018 9917
rect 65698 9823 65853 9869
rect 65899 9823 66018 9869
rect 65698 9775 66018 9823
rect 65698 9729 65853 9775
rect 65899 9729 66018 9775
rect 65698 9681 66018 9729
rect 65698 9635 65853 9681
rect 65899 9635 66018 9681
rect 65698 9587 66018 9635
rect 65698 9541 65853 9587
rect 65899 9541 66018 9587
rect 65698 9493 66018 9541
rect 65698 9447 65853 9493
rect 65899 9447 66018 9493
rect 65698 9399 66018 9447
rect 65698 9353 65853 9399
rect 65899 9353 66018 9399
rect 65698 9305 66018 9353
rect 65698 9259 65853 9305
rect 65899 9259 66018 9305
rect 65698 9211 66018 9259
rect 65698 9165 65853 9211
rect 65899 9165 66018 9211
rect 65698 9117 66018 9165
rect 65698 9071 65853 9117
rect 65899 9071 66018 9117
rect 65698 9023 66018 9071
rect 65698 8977 65853 9023
rect 65899 8977 66018 9023
rect 65698 8929 66018 8977
rect 65698 8883 65853 8929
rect 65899 8883 66018 8929
rect 65698 8835 66018 8883
rect 65698 8789 65853 8835
rect 65899 8789 66018 8835
rect 65698 8741 66018 8789
rect 65698 8695 65853 8741
rect 65899 8695 66018 8741
rect 65698 8647 66018 8695
rect 65698 8601 65853 8647
rect 65899 8601 66018 8647
rect 65698 8553 66018 8601
rect 65698 8507 65853 8553
rect 65899 8507 66018 8553
rect 65698 8459 66018 8507
rect 65698 8413 65853 8459
rect 65899 8413 66018 8459
rect 65698 8365 66018 8413
rect 65698 8319 65853 8365
rect 65899 8319 66018 8365
rect 65698 8271 66018 8319
rect 65698 8225 65853 8271
rect 65899 8225 66018 8271
rect 65698 8177 66018 8225
rect 65698 8131 65853 8177
rect 65899 8131 66018 8177
rect 65698 8083 66018 8131
rect 65698 8037 65853 8083
rect 65899 8037 66018 8083
rect 65698 7989 66018 8037
rect 65698 7943 65853 7989
rect 65899 7943 66018 7989
rect 65698 7895 66018 7943
rect 65698 7849 65853 7895
rect 65899 7849 66018 7895
rect 65698 7801 66018 7849
rect 65698 7755 65853 7801
rect 65899 7755 66018 7801
rect 65698 7707 66018 7755
rect 65698 7661 65853 7707
rect 65899 7661 66018 7707
rect 65698 7613 66018 7661
rect 65698 7579 65853 7613
rect 61763 7567 65853 7579
rect 65899 7567 66018 7613
rect 32510 7519 66018 7567
rect 32510 7473 32629 7519
rect 32675 7473 36765 7519
rect 36811 7473 40901 7519
rect 40947 7473 42325 7519
rect 42371 7473 46461 7519
rect 46507 7473 50597 7519
rect 50643 7473 52021 7519
rect 52067 7473 56157 7519
rect 56203 7473 60293 7519
rect 60339 7473 61717 7519
rect 61763 7473 65853 7519
rect 65899 7473 66018 7519
rect 32510 7425 66018 7473
rect 32510 7379 32629 7425
rect 32675 7379 32723 7425
rect 32769 7379 32817 7425
rect 32863 7379 32911 7425
rect 32957 7379 33005 7425
rect 33051 7379 33099 7425
rect 33145 7379 33193 7425
rect 33239 7379 33287 7425
rect 33333 7379 33381 7425
rect 33427 7379 33475 7425
rect 33521 7379 33569 7425
rect 33615 7379 33663 7425
rect 33709 7379 33757 7425
rect 33803 7379 33851 7425
rect 33897 7379 33945 7425
rect 33991 7379 34039 7425
rect 34085 7379 34133 7425
rect 34179 7379 34227 7425
rect 34273 7379 34321 7425
rect 34367 7379 34415 7425
rect 34461 7379 34509 7425
rect 34555 7379 34603 7425
rect 34649 7379 34697 7425
rect 34743 7379 34791 7425
rect 34837 7379 34885 7425
rect 34931 7379 34979 7425
rect 35025 7379 35073 7425
rect 35119 7379 35167 7425
rect 35213 7379 35261 7425
rect 35307 7379 35355 7425
rect 35401 7379 35449 7425
rect 35495 7379 35543 7425
rect 35589 7379 35637 7425
rect 35683 7379 35731 7425
rect 35777 7379 35825 7425
rect 35871 7379 35919 7425
rect 35965 7379 36013 7425
rect 36059 7379 36107 7425
rect 36153 7379 36201 7425
rect 36247 7379 36295 7425
rect 36341 7379 36389 7425
rect 36435 7379 36483 7425
rect 36529 7379 36577 7425
rect 36623 7379 36671 7425
rect 36717 7379 36765 7425
rect 36811 7379 36859 7425
rect 36905 7379 36953 7425
rect 36999 7379 37047 7425
rect 37093 7379 37141 7425
rect 37187 7379 37235 7425
rect 37281 7379 37329 7425
rect 37375 7379 37423 7425
rect 37469 7379 37517 7425
rect 37563 7379 37611 7425
rect 37657 7379 37705 7425
rect 37751 7379 37799 7425
rect 37845 7379 37893 7425
rect 37939 7379 37987 7425
rect 38033 7379 38081 7425
rect 38127 7379 38175 7425
rect 38221 7379 38269 7425
rect 38315 7379 38363 7425
rect 38409 7379 38457 7425
rect 38503 7379 38551 7425
rect 38597 7379 38645 7425
rect 38691 7379 38739 7425
rect 38785 7379 38833 7425
rect 38879 7379 38927 7425
rect 38973 7379 39021 7425
rect 39067 7379 39115 7425
rect 39161 7379 39209 7425
rect 39255 7379 39303 7425
rect 39349 7379 39397 7425
rect 39443 7379 39491 7425
rect 39537 7379 39585 7425
rect 39631 7379 39679 7425
rect 39725 7379 39773 7425
rect 39819 7379 39867 7425
rect 39913 7379 39961 7425
rect 40007 7379 40055 7425
rect 40101 7379 40149 7425
rect 40195 7379 40243 7425
rect 40289 7379 40337 7425
rect 40383 7379 40431 7425
rect 40477 7379 40525 7425
rect 40571 7379 40619 7425
rect 40665 7379 40713 7425
rect 40759 7379 40807 7425
rect 40853 7379 40901 7425
rect 40947 7379 42325 7425
rect 42371 7379 42419 7425
rect 42465 7379 42513 7425
rect 42559 7379 42607 7425
rect 42653 7379 42701 7425
rect 42747 7379 42795 7425
rect 42841 7379 42889 7425
rect 42935 7379 42983 7425
rect 43029 7379 43077 7425
rect 43123 7379 43171 7425
rect 43217 7379 43265 7425
rect 43311 7379 43359 7425
rect 43405 7379 43453 7425
rect 43499 7379 43547 7425
rect 43593 7379 43641 7425
rect 43687 7379 43735 7425
rect 43781 7379 43829 7425
rect 43875 7379 43923 7425
rect 43969 7379 44017 7425
rect 44063 7379 44111 7425
rect 44157 7379 44205 7425
rect 44251 7379 44299 7425
rect 44345 7379 44393 7425
rect 44439 7379 44487 7425
rect 44533 7379 44581 7425
rect 44627 7379 44675 7425
rect 44721 7379 44769 7425
rect 44815 7379 44863 7425
rect 44909 7379 44957 7425
rect 45003 7379 45051 7425
rect 45097 7379 45145 7425
rect 45191 7379 45239 7425
rect 45285 7379 45333 7425
rect 45379 7379 45427 7425
rect 45473 7379 45521 7425
rect 45567 7379 45615 7425
rect 45661 7379 45709 7425
rect 45755 7379 45803 7425
rect 45849 7379 45897 7425
rect 45943 7379 45991 7425
rect 46037 7379 46085 7425
rect 46131 7379 46179 7425
rect 46225 7379 46273 7425
rect 46319 7379 46367 7425
rect 46413 7379 46461 7425
rect 46507 7379 46555 7425
rect 46601 7379 46649 7425
rect 46695 7379 46743 7425
rect 46789 7379 46837 7425
rect 46883 7379 46931 7425
rect 46977 7379 47025 7425
rect 47071 7379 47119 7425
rect 47165 7379 47213 7425
rect 47259 7379 47307 7425
rect 47353 7379 47401 7425
rect 47447 7379 47495 7425
rect 47541 7379 47589 7425
rect 47635 7379 47683 7425
rect 47729 7379 47777 7425
rect 47823 7379 47871 7425
rect 47917 7379 47965 7425
rect 48011 7379 48059 7425
rect 48105 7379 48153 7425
rect 48199 7379 48247 7425
rect 48293 7379 48341 7425
rect 48387 7379 48435 7425
rect 48481 7379 48529 7425
rect 48575 7379 48623 7425
rect 48669 7379 48717 7425
rect 48763 7379 48811 7425
rect 48857 7379 48905 7425
rect 48951 7379 48999 7425
rect 49045 7379 49093 7425
rect 49139 7379 49187 7425
rect 49233 7379 49281 7425
rect 49327 7379 49375 7425
rect 49421 7379 49469 7425
rect 49515 7379 49563 7425
rect 49609 7379 49657 7425
rect 49703 7379 49751 7425
rect 49797 7379 49845 7425
rect 49891 7379 49939 7425
rect 49985 7379 50033 7425
rect 50079 7379 50127 7425
rect 50173 7379 50221 7425
rect 50267 7379 50315 7425
rect 50361 7379 50409 7425
rect 50455 7379 50503 7425
rect 50549 7379 50597 7425
rect 50643 7379 52021 7425
rect 52067 7379 52115 7425
rect 52161 7379 52209 7425
rect 52255 7379 52303 7425
rect 52349 7379 52397 7425
rect 52443 7379 52491 7425
rect 52537 7379 52585 7425
rect 52631 7379 52679 7425
rect 52725 7379 52773 7425
rect 52819 7379 52867 7425
rect 52913 7379 52961 7425
rect 53007 7379 53055 7425
rect 53101 7379 53149 7425
rect 53195 7379 53243 7425
rect 53289 7379 53337 7425
rect 53383 7379 53431 7425
rect 53477 7379 53525 7425
rect 53571 7379 53619 7425
rect 53665 7379 53713 7425
rect 53759 7379 53807 7425
rect 53853 7379 53901 7425
rect 53947 7379 53995 7425
rect 54041 7379 54089 7425
rect 54135 7379 54183 7425
rect 54229 7379 54277 7425
rect 54323 7379 54371 7425
rect 54417 7379 54465 7425
rect 54511 7379 54559 7425
rect 54605 7379 54653 7425
rect 54699 7379 54747 7425
rect 54793 7379 54841 7425
rect 54887 7379 54935 7425
rect 54981 7379 55029 7425
rect 55075 7379 55123 7425
rect 55169 7379 55217 7425
rect 55263 7379 55311 7425
rect 55357 7379 55405 7425
rect 55451 7379 55499 7425
rect 55545 7379 55593 7425
rect 55639 7379 55687 7425
rect 55733 7379 55781 7425
rect 55827 7379 55875 7425
rect 55921 7379 55969 7425
rect 56015 7379 56063 7425
rect 56109 7379 56157 7425
rect 56203 7379 56251 7425
rect 56297 7379 56345 7425
rect 56391 7379 56439 7425
rect 56485 7379 56533 7425
rect 56579 7379 56627 7425
rect 56673 7379 56721 7425
rect 56767 7379 56815 7425
rect 56861 7379 56909 7425
rect 56955 7379 57003 7425
rect 57049 7379 57097 7425
rect 57143 7379 57191 7425
rect 57237 7379 57285 7425
rect 57331 7379 57379 7425
rect 57425 7379 57473 7425
rect 57519 7379 57567 7425
rect 57613 7379 57661 7425
rect 57707 7379 57755 7425
rect 57801 7379 57849 7425
rect 57895 7379 57943 7425
rect 57989 7379 58037 7425
rect 58083 7379 58131 7425
rect 58177 7379 58225 7425
rect 58271 7379 58319 7425
rect 58365 7379 58413 7425
rect 58459 7379 58507 7425
rect 58553 7379 58601 7425
rect 58647 7379 58695 7425
rect 58741 7379 58789 7425
rect 58835 7379 58883 7425
rect 58929 7379 58977 7425
rect 59023 7379 59071 7425
rect 59117 7379 59165 7425
rect 59211 7379 59259 7425
rect 59305 7379 59353 7425
rect 59399 7379 59447 7425
rect 59493 7379 59541 7425
rect 59587 7379 59635 7425
rect 59681 7379 59729 7425
rect 59775 7379 59823 7425
rect 59869 7379 59917 7425
rect 59963 7379 60011 7425
rect 60057 7379 60105 7425
rect 60151 7379 60199 7425
rect 60245 7379 60293 7425
rect 60339 7379 61717 7425
rect 61763 7379 61811 7425
rect 61857 7379 61905 7425
rect 61951 7379 61999 7425
rect 62045 7379 62093 7425
rect 62139 7379 62187 7425
rect 62233 7379 62281 7425
rect 62327 7379 62375 7425
rect 62421 7379 62469 7425
rect 62515 7379 62563 7425
rect 62609 7379 62657 7425
rect 62703 7379 62751 7425
rect 62797 7379 62845 7425
rect 62891 7379 62939 7425
rect 62985 7379 63033 7425
rect 63079 7379 63127 7425
rect 63173 7379 63221 7425
rect 63267 7379 63315 7425
rect 63361 7379 63409 7425
rect 63455 7379 63503 7425
rect 63549 7379 63597 7425
rect 63643 7379 63691 7425
rect 63737 7379 63785 7425
rect 63831 7379 63879 7425
rect 63925 7379 63973 7425
rect 64019 7379 64067 7425
rect 64113 7379 64161 7425
rect 64207 7379 64255 7425
rect 64301 7379 64349 7425
rect 64395 7379 64443 7425
rect 64489 7379 64537 7425
rect 64583 7379 64631 7425
rect 64677 7379 64725 7425
rect 64771 7379 64819 7425
rect 64865 7379 64913 7425
rect 64959 7379 65007 7425
rect 65053 7379 65101 7425
rect 65147 7379 65195 7425
rect 65241 7379 65289 7425
rect 65335 7379 65383 7425
rect 65429 7379 65477 7425
rect 65523 7379 65571 7425
rect 65617 7379 65665 7425
rect 65711 7379 65759 7425
rect 65805 7379 65853 7425
rect 65899 7379 66018 7425
rect 32510 7259 66018 7379
rect 1623 4849 1783 7221
rect 2175 5312 2355 5320
rect 2175 5308 2643 5312
rect 2175 5256 2187 5308
rect 2239 5256 2291 5308
rect 2343 5256 2643 5308
rect 2175 5204 2643 5256
rect 2175 5152 2187 5204
rect 2239 5152 2291 5204
rect 2343 5152 2643 5204
rect 3057 5185 3217 5475
rect 3047 5173 3227 5185
rect 2175 5140 2355 5152
rect 3047 5121 3059 5173
rect 3111 5121 3163 5173
rect 3215 5121 3227 5173
rect 3047 5069 3227 5121
rect 3047 5017 3059 5069
rect 3111 5017 3163 5069
rect 3215 5017 3227 5069
rect 3047 5005 3227 5017
rect 3925 4849 4085 7221
rect 4914 6860 5074 7221
rect 5525 7004 5685 7221
rect 6867 7211 6934 7221
rect 6980 7211 7047 7221
rect 9969 7211 10149 7221
rect 11867 7004 12027 7221
rect 5525 6860 12027 7004
rect 4914 6826 12027 6860
rect 12267 6826 12427 7221
rect 16899 6826 17059 7221
rect 32510 6826 32830 7259
rect 36610 6826 36930 7259
rect 40710 6826 41030 7259
rect 42170 6826 42490 7259
rect 46270 6826 46590 7259
rect 50370 6826 50690 7259
rect 51830 6826 52150 7259
rect 55930 6826 56250 7259
rect 60030 6826 60350 7259
rect 61490 6826 61810 7259
rect 65698 6826 66018 7259
rect 4914 6506 66018 6826
rect 4914 4849 5074 6506
rect 11371 6436 17403 6448
rect 8275 6411 8455 6421
rect 8275 6409 8745 6411
rect 8275 6357 8287 6409
rect 8339 6357 8391 6409
rect 8443 6357 8745 6409
rect 8275 6305 8745 6357
rect 8275 6253 8287 6305
rect 8339 6253 8391 6305
rect 8443 6253 8745 6305
rect 8275 6251 8745 6253
rect 11371 6384 11383 6436
rect 11435 6384 11487 6436
rect 11539 6384 17131 6436
rect 17183 6384 17235 6436
rect 17287 6384 17339 6436
rect 17391 6384 17403 6436
rect 11371 6332 17403 6384
rect 11371 6280 11383 6332
rect 11435 6280 11487 6332
rect 11539 6280 17131 6332
rect 17183 6280 17235 6332
rect 17287 6280 17339 6332
rect 17391 6280 17403 6332
rect 8275 6241 8455 6251
rect 11371 6228 17403 6280
rect 6867 6175 7047 6185
rect 9969 6175 10149 6185
rect 6867 6173 10149 6175
rect 6867 6121 6879 6173
rect 6931 6121 6983 6173
rect 7035 6121 9981 6173
rect 10033 6121 10085 6173
rect 10137 6121 10149 6173
rect 11371 6176 11383 6228
rect 11435 6176 11487 6228
rect 11539 6176 17131 6228
rect 17183 6176 17235 6228
rect 17287 6176 17339 6228
rect 17391 6176 17403 6228
rect 11371 6164 17403 6176
rect 6867 6118 10149 6121
rect 6877 6072 6934 6118
rect 6980 6072 7028 6118
rect 7074 6072 7122 6118
rect 7168 6072 7216 6118
rect 7262 6072 7310 6118
rect 7356 6072 7404 6118
rect 7450 6072 7498 6118
rect 7544 6072 7592 6118
rect 7638 6072 7686 6118
rect 7732 6072 7780 6118
rect 7826 6072 7874 6118
rect 7920 6072 7968 6118
rect 8014 6072 8062 6118
rect 8108 6072 8156 6118
rect 8202 6072 8250 6118
rect 8296 6072 8344 6118
rect 8390 6072 8438 6118
rect 8484 6072 8532 6118
rect 8578 6072 8626 6118
rect 8672 6072 8720 6118
rect 8766 6072 8814 6118
rect 8860 6072 8908 6118
rect 8954 6072 9002 6118
rect 9048 6072 9096 6118
rect 9142 6072 9190 6118
rect 9236 6072 9284 6118
rect 9330 6072 9378 6118
rect 9424 6072 9472 6118
rect 9518 6072 9566 6118
rect 9612 6072 9660 6118
rect 9706 6072 9754 6118
rect 9800 6072 9848 6118
rect 9894 6072 9942 6118
rect 9988 6072 10036 6118
rect 10082 6072 10149 6118
rect 6867 6069 10149 6072
rect 6867 6017 6879 6069
rect 6931 6024 6983 6069
rect 6931 6017 6934 6024
rect 6867 6005 6934 6017
rect 6877 5978 6934 6005
rect 6980 6017 6983 6024
rect 7035 6017 9981 6069
rect 10033 6024 10085 6069
rect 10033 6017 10036 6024
rect 6980 6015 10036 6017
rect 6980 6005 7047 6015
rect 6980 5978 7037 6005
rect 6877 5930 7037 5978
rect 6877 5884 6934 5930
rect 6980 5884 7037 5930
rect 6877 5836 7037 5884
rect 6877 5790 6934 5836
rect 6980 5790 7037 5836
rect 6877 5742 7037 5790
rect 6877 5696 6934 5742
rect 6980 5696 7037 5742
rect 6877 5648 7037 5696
rect 6877 5602 6934 5648
rect 6980 5602 7037 5648
rect 6877 5554 7037 5602
rect 6877 5508 6934 5554
rect 6980 5508 7037 5554
rect 5144 5463 5324 5471
rect 5144 5459 5624 5463
rect 5144 5407 5156 5459
rect 5208 5407 5260 5459
rect 5312 5407 5624 5459
rect 5144 5355 5624 5407
rect 5144 5303 5156 5355
rect 5208 5303 5260 5355
rect 5312 5303 5624 5355
rect 6877 5460 7037 5508
rect 6877 5414 6934 5460
rect 6980 5414 7037 5460
rect 6877 5366 7037 5414
rect 6877 5320 6934 5366
rect 6980 5320 7037 5366
rect 5144 5291 5324 5303
rect 872 4792 5074 4849
rect 872 4746 929 4792
rect 975 4746 1023 4792
rect 1069 4746 1117 4792
rect 1163 4746 1211 4792
rect 1257 4746 1305 4792
rect 1351 4746 1399 4792
rect 1445 4746 1493 4792
rect 1539 4746 1587 4792
rect 1633 4746 1681 4792
rect 1727 4746 1775 4792
rect 1821 4746 1869 4792
rect 1915 4746 1963 4792
rect 2009 4746 2057 4792
rect 2103 4746 2151 4792
rect 2197 4746 2245 4792
rect 2291 4746 2339 4792
rect 2385 4746 2433 4792
rect 2479 4746 2527 4792
rect 2573 4746 2621 4792
rect 2667 4746 2715 4792
rect 2761 4746 2809 4792
rect 2855 4746 2903 4792
rect 2949 4746 2997 4792
rect 3043 4746 3091 4792
rect 3137 4746 3185 4792
rect 3231 4746 3279 4792
rect 3325 4746 3373 4792
rect 3419 4746 3467 4792
rect 3513 4746 3561 4792
rect 3607 4746 3655 4792
rect 3701 4746 3749 4792
rect 3795 4746 3843 4792
rect 3889 4746 3937 4792
rect 3983 4746 4031 4792
rect 4077 4746 4125 4792
rect 4171 4746 4219 4792
rect 4265 4746 4313 4792
rect 4359 4746 4407 4792
rect 4453 4746 4501 4792
rect 4547 4746 4595 4792
rect 4641 4746 4689 4792
rect 4735 4746 4783 4792
rect 4829 4746 4877 4792
rect 4923 4746 4971 4792
rect 5017 4746 5074 4792
rect 872 4698 5074 4746
rect 872 4652 929 4698
rect 975 4689 4971 4698
rect 975 4652 1032 4689
rect 872 4604 1032 4652
rect 872 4558 929 4604
rect 975 4558 1032 4604
rect 872 4510 1032 4558
rect 872 4464 929 4510
rect 975 4464 1032 4510
rect 872 4416 1032 4464
rect 872 4370 929 4416
rect 975 4370 1032 4416
rect 872 4322 1032 4370
rect 872 4276 929 4322
rect 975 4276 1032 4322
rect 872 4228 1032 4276
rect 872 4182 929 4228
rect 975 4182 1032 4228
rect 872 4134 1032 4182
rect 872 4088 929 4134
rect 975 4088 1032 4134
rect 872 4040 1032 4088
rect 872 3994 929 4040
rect 975 3994 1032 4040
rect 872 3946 1032 3994
rect 872 3900 929 3946
rect 975 3900 1032 3946
rect 872 3852 1032 3900
rect 872 3806 929 3852
rect 975 3806 1032 3852
rect 872 3758 1032 3806
rect 872 3712 929 3758
rect 975 3712 1032 3758
rect 872 3664 1032 3712
rect 872 3618 929 3664
rect 975 3618 1032 3664
rect 872 3570 1032 3618
rect 872 3524 929 3570
rect 975 3524 1032 3570
rect 872 3476 1032 3524
rect 872 3430 929 3476
rect 975 3430 1032 3476
rect 872 3382 1032 3430
rect 872 3336 929 3382
rect 975 3336 1032 3382
rect 872 3288 1032 3336
rect 872 3242 929 3288
rect 975 3242 1032 3288
rect 872 3194 1032 3242
rect 872 3148 929 3194
rect 975 3148 1032 3194
rect 872 3100 1032 3148
rect 872 3054 929 3100
rect 975 3054 1032 3100
rect 872 3006 1032 3054
rect 872 2960 929 3006
rect 975 2960 1032 3006
rect 872 2912 1032 2960
rect 872 2866 929 2912
rect 975 2866 1032 2912
rect 872 2818 1032 2866
rect 872 2772 929 2818
rect 975 2772 1032 2818
rect 872 2724 1032 2772
rect 872 2678 929 2724
rect 975 2678 1032 2724
rect 872 2630 1032 2678
rect 872 2584 929 2630
rect 975 2584 1032 2630
rect 872 2536 1032 2584
rect 872 2490 929 2536
rect 975 2490 1032 2536
rect 872 2442 1032 2490
rect 872 2396 929 2442
rect 975 2396 1032 2442
rect 872 2348 1032 2396
rect 872 2302 929 2348
rect 975 2302 1032 2348
rect 872 2254 1032 2302
rect 872 2208 929 2254
rect 975 2208 1032 2254
rect 872 2160 1032 2208
rect 872 2114 929 2160
rect 975 2114 1032 2160
rect 872 2066 1032 2114
rect 872 2020 929 2066
rect 975 2020 1032 2066
rect 872 1972 1032 2020
rect 872 1926 929 1972
rect 975 1926 1032 1972
rect 872 1878 1032 1926
rect 872 1832 929 1878
rect 975 1832 1032 1878
rect 872 1784 1032 1832
rect 872 1738 929 1784
rect 975 1738 1032 1784
rect 872 1690 1032 1738
rect 872 1644 929 1690
rect 975 1644 1032 1690
rect 872 1596 1032 1644
rect 872 1550 929 1596
rect 975 1559 1032 1596
rect 1290 4515 1336 4689
rect 1450 4515 1496 4689
rect 1578 4515 1624 4689
rect 1738 4515 1784 4689
rect 1290 4469 1658 4515
rect 1704 4469 1784 4515
rect 1290 4421 1336 4469
rect 1290 3255 1336 3647
rect 1450 4421 1496 4469
rect 1450 3255 1496 3647
rect 1578 4421 1624 4469
rect 1578 3636 1624 3647
rect 1738 4421 1784 4469
rect 1738 3636 1784 3647
rect 1866 4421 1912 4432
rect 1866 3590 1912 3647
rect 2082 4421 2128 4689
rect 2175 4556 2355 4568
rect 2175 4504 2187 4556
rect 2239 4504 2291 4556
rect 2343 4504 2355 4556
rect 2175 4492 2355 4504
rect 2082 3636 2128 3647
rect 2298 4421 2344 4432
rect 2298 3590 2344 3647
rect 2514 4421 2560 4689
rect 2730 4431 2776 4432
rect 2715 4421 2791 4431
rect 2715 4419 2730 4421
rect 2776 4419 2791 4421
rect 2715 4367 2727 4419
rect 2779 4367 2791 4419
rect 2715 4315 2730 4367
rect 2776 4315 2791 4367
rect 2715 4263 2727 4315
rect 2779 4263 2791 4315
rect 2715 4251 2730 4263
rect 2514 3636 2560 3647
rect 2776 4251 2791 4263
rect 2946 4421 2992 4689
rect 2730 3590 2776 3647
rect 2946 3636 2992 3647
rect 3162 4421 3208 4432
rect 1866 3544 2776 3590
rect 3162 3590 3208 3647
rect 3378 4421 3424 4689
rect 3594 4421 3640 4432
rect 3378 3636 3424 3647
rect 3579 3805 3594 3817
rect 3810 4421 3856 4689
rect 4242 4513 4288 4689
rect 4402 4513 4448 4689
rect 4562 4513 4608 4689
rect 4242 4467 4322 4513
rect 4368 4467 4482 4513
rect 4528 4467 4608 4513
rect 3640 3805 3655 3817
rect 3579 3753 3591 3805
rect 3643 3753 3655 3805
rect 3579 3701 3594 3753
rect 3640 3701 3655 3753
rect 3579 3649 3591 3701
rect 3643 3649 3655 3701
rect 3579 3647 3594 3649
rect 3640 3647 3655 3649
rect 3579 3637 3655 3647
rect 4026 4421 4072 4432
rect 4011 4129 4026 4141
rect 4242 4421 4288 4467
rect 4072 4129 4087 4141
rect 4011 4077 4023 4129
rect 4075 4077 4087 4129
rect 4011 4025 4026 4077
rect 4072 4025 4087 4077
rect 4011 3973 4023 4025
rect 4075 3973 4087 4025
rect 4011 3961 4026 3973
rect 3594 3590 3640 3637
rect 3810 3636 3856 3647
rect 4072 3961 4087 3973
rect 4026 3636 4072 3647
rect 4242 3636 4288 3647
rect 4402 4421 4448 4467
rect 4402 3636 4448 3647
rect 4562 4421 4608 4467
rect 4562 3636 4608 3647
rect 4914 4652 4971 4689
rect 5017 4652 5074 4698
rect 4914 4604 5074 4652
rect 4914 4558 4971 4604
rect 5017 4558 5074 4604
rect 4914 4510 5074 4558
rect 4914 4464 4971 4510
rect 5017 4464 5074 4510
rect 4914 4416 5074 4464
rect 4914 4370 4971 4416
rect 5017 4370 5074 4416
rect 6877 5272 7037 5320
rect 6877 5226 6934 5272
rect 6980 5226 7037 5272
rect 6877 5178 7037 5226
rect 6877 5132 6934 5178
rect 6980 5132 7037 5178
rect 6877 5084 7037 5132
rect 6877 5038 6934 5084
rect 6980 5038 7037 5084
rect 6877 4990 7037 5038
rect 6877 4944 6934 4990
rect 6980 4944 7037 4990
rect 6877 4896 7037 4944
rect 6877 4850 6934 4896
rect 6980 4850 7037 4896
rect 6877 4802 7037 4850
rect 6877 4756 6934 4802
rect 6980 4756 7037 4802
rect 6877 4708 7037 4756
rect 6877 4662 6934 4708
rect 6980 4662 7037 4708
rect 6877 4614 7037 4662
rect 6877 4568 6934 4614
rect 6980 4568 7037 4614
rect 6877 4520 7037 4568
rect 6877 4474 6934 4520
rect 6980 4474 7037 4520
rect 6877 4426 7037 4474
rect 4914 4322 5074 4370
rect 4914 4276 4971 4322
rect 5017 4276 5074 4322
rect 4914 4228 5074 4276
rect 4914 4182 4971 4228
rect 5017 4182 5074 4228
rect 4914 4134 5074 4182
rect 4914 4088 4971 4134
rect 5017 4088 5074 4134
rect 6554 4113 6714 4403
rect 6877 4380 6934 4426
rect 6980 4380 7037 4426
rect 6877 4332 7037 4380
rect 6877 4286 6934 4332
rect 6980 4286 7037 4332
rect 6877 4238 7037 4286
rect 6877 4192 6934 4238
rect 6980 4192 7037 4238
rect 6877 4144 7037 4192
rect 4914 4040 5074 4088
rect 4914 3994 4971 4040
rect 5017 3994 5074 4040
rect 4914 3946 5074 3994
rect 4914 3900 4971 3946
rect 5017 3900 5074 3946
rect 6544 4101 6724 4113
rect 6544 4049 6556 4101
rect 6608 4049 6660 4101
rect 6712 4049 6724 4101
rect 6544 3997 6724 4049
rect 6544 3945 6556 3997
rect 6608 3945 6660 3997
rect 6712 3945 6724 3997
rect 6544 3933 6724 3945
rect 6877 4098 6934 4144
rect 6980 4098 7037 4144
rect 6877 4050 7037 4098
rect 6877 4004 6934 4050
rect 6980 4004 7037 4050
rect 6877 3956 7037 4004
rect 4914 3852 5074 3900
rect 4914 3806 4971 3852
rect 5017 3806 5074 3852
rect 4914 3758 5074 3806
rect 4914 3712 4971 3758
rect 5017 3712 5074 3758
rect 4914 3664 5074 3712
rect 3162 3544 3640 3590
rect 4914 3618 4971 3664
rect 5017 3618 5074 3664
rect 4914 3570 5074 3618
rect 4914 3524 4971 3570
rect 5017 3524 5074 3570
rect 4914 3476 5074 3524
rect 4914 3430 4971 3476
rect 5017 3430 5074 3476
rect 4914 3382 5074 3430
rect 1874 3295 2102 3341
rect 2148 3295 2206 3341
rect 2252 3295 2310 3341
rect 2356 3295 2414 3341
rect 2460 3295 2518 3341
rect 2564 3295 2622 3341
rect 2668 3295 2784 3341
rect 1290 3209 1370 3255
rect 1416 3209 1666 3255
rect 1712 3209 1792 3255
rect 1290 3161 1336 3209
rect 1290 1901 1336 2387
rect 1290 1559 1336 1827
rect 1450 3161 1496 3209
rect 1450 1901 1496 2387
rect 1586 3161 1632 3209
rect 1586 2376 1632 2387
rect 1746 3161 1792 3209
rect 1746 2330 1792 2387
rect 1874 3161 1920 3295
rect 1874 2376 1920 2387
rect 2090 3161 2136 3172
rect 2090 2330 2136 2387
rect 2306 3161 2352 3295
rect 2306 2376 2352 2387
rect 2522 3161 2568 3172
rect 2738 3171 2784 3295
rect 4914 3336 4971 3382
rect 5017 3336 5074 3382
rect 4914 3288 5074 3336
rect 3274 3218 4234 3264
rect 4280 3218 4530 3264
rect 4576 3218 4656 3264
rect 2725 3161 2801 3171
rect 2725 3159 2738 3161
rect 2784 3159 2801 3161
rect 2725 3107 2737 3159
rect 2789 3107 2801 3159
rect 2725 3055 2738 3107
rect 2784 3055 2801 3107
rect 2725 3003 2737 3055
rect 2789 3003 2801 3055
rect 2725 2991 2738 3003
rect 2522 2330 2568 2387
rect 2784 2991 2801 3003
rect 2954 3161 3000 3172
rect 3114 3171 3160 3172
rect 2738 2376 2784 2387
rect 3099 3161 3175 3171
rect 3099 3159 3114 3161
rect 3160 3159 3175 3161
rect 3099 3107 3111 3159
rect 3163 3107 3175 3159
rect 3099 3055 3114 3107
rect 3160 3055 3175 3107
rect 3099 3003 3111 3055
rect 3163 3003 3175 3055
rect 3099 2991 3114 3003
rect 2954 2330 3000 2387
rect 3160 2991 3175 3003
rect 3274 3161 3320 3218
rect 3434 3171 3480 3172
rect 3114 2350 3160 2387
rect 3419 3161 3495 3171
rect 3419 3159 3434 3161
rect 3480 3159 3495 3161
rect 3419 3107 3431 3159
rect 3483 3107 3495 3159
rect 3419 3055 3434 3107
rect 3480 3055 3495 3107
rect 3419 3003 3431 3055
rect 3483 3003 3495 3055
rect 3419 2991 3434 3003
rect 3274 2376 3320 2387
rect 3480 2991 3495 3003
rect 3594 3161 3640 3218
rect 3434 2350 3480 2387
rect 3594 2376 3640 2387
rect 3810 3161 3856 3172
rect 3938 3161 3984 3172
rect 1746 2284 3000 2330
rect 3103 2339 3171 2350
rect 3103 2293 3114 2339
rect 3160 2293 3171 2339
rect 3103 2282 3171 2293
rect 3423 2339 3491 2350
rect 3423 2293 3434 2339
rect 3480 2293 3491 2339
rect 3423 2282 3491 2293
rect 3691 2341 3759 2352
rect 3810 2341 3856 2387
rect 3923 2543 3938 2555
rect 4154 3161 4200 3218
rect 3984 2543 3999 2555
rect 3923 2491 3935 2543
rect 3987 2491 3999 2543
rect 3923 2439 3938 2491
rect 3984 2439 3999 2491
rect 3923 2387 3935 2439
rect 3987 2387 3999 2439
rect 3923 2375 3999 2387
rect 4154 2376 4200 2387
rect 4314 3161 4360 3218
rect 4314 2376 4360 2387
rect 4450 3161 4496 3218
rect 3691 2295 3702 2341
rect 3748 2295 3856 2341
rect 3691 2284 3759 2295
rect 1450 1559 1496 1827
rect 1586 1958 4192 2004
rect 1586 1901 1632 1958
rect 1586 1816 1632 1827
rect 1746 1901 1792 1912
rect 1746 1770 1792 1827
rect 1906 1901 1952 1958
rect 1906 1816 1952 1827
rect 2066 1901 2112 1912
rect 2066 1770 2112 1827
rect 2226 1901 2272 1958
rect 2226 1816 2272 1827
rect 2386 1901 2432 1912
rect 2386 1770 2432 1827
rect 2546 1901 2592 1958
rect 2546 1816 2592 1827
rect 2706 1901 2752 1912
rect 2706 1770 2752 1827
rect 2866 1901 2912 1958
rect 2866 1816 2912 1827
rect 3026 1901 3072 1912
rect 3026 1770 3072 1827
rect 3186 1901 3232 1958
rect 3186 1816 3232 1827
rect 3346 1901 3392 1912
rect 3346 1770 3392 1827
rect 3506 1901 3552 1958
rect 3506 1816 3552 1827
rect 3666 1901 3712 1912
rect 3666 1770 3712 1827
rect 3826 1901 3872 1958
rect 3826 1816 3872 1827
rect 3986 1901 4032 1912
rect 3986 1785 4032 1827
rect 4146 1901 4192 1958
rect 4146 1816 4192 1827
rect 4450 1901 4496 2387
rect 3971 1773 4047 1785
rect 3971 1770 3983 1773
rect 1746 1724 1826 1770
rect 1872 1724 1986 1770
rect 2032 1724 2466 1770
rect 2512 1724 3106 1770
rect 3152 1724 3983 1770
rect 3346 1723 3392 1724
rect 3971 1721 3983 1724
rect 4035 1721 4047 1773
rect 3971 1669 4047 1721
rect 3971 1617 3983 1669
rect 4035 1617 4047 1669
rect 3971 1605 4047 1617
rect 4450 1559 4496 1827
rect 4610 3161 4656 3218
rect 4610 1901 4656 2387
rect 4610 1559 4656 1827
rect 4914 3242 4971 3288
rect 5017 3242 5074 3288
rect 4914 3194 5074 3242
rect 4914 3148 4971 3194
rect 5017 3148 5074 3194
rect 4914 3100 5074 3148
rect 4914 3054 4971 3100
rect 5017 3054 5074 3100
rect 4914 3006 5074 3054
rect 4914 2960 4971 3006
rect 5017 2960 5074 3006
rect 4914 2912 5074 2960
rect 4914 2866 4971 2912
rect 5017 2866 5074 2912
rect 6877 3910 6934 3956
rect 6980 3910 7037 3956
rect 6877 3862 7037 3910
rect 6877 3816 6934 3862
rect 6980 3816 7037 3862
rect 6877 3768 7037 3816
rect 6877 3722 6934 3768
rect 6980 3722 7037 3768
rect 6877 3674 7037 3722
rect 6877 3628 6934 3674
rect 6980 3628 7037 3674
rect 6877 3580 7037 3628
rect 6877 3534 6934 3580
rect 6980 3534 7037 3580
rect 6877 3486 7037 3534
rect 6877 3440 6934 3486
rect 6980 3440 7037 3486
rect 6877 3392 7037 3440
rect 6877 3346 6934 3392
rect 6980 3346 7037 3392
rect 6877 3298 7037 3346
rect 6877 3252 6934 3298
rect 6980 3252 7037 3298
rect 6877 3204 7037 3252
rect 6877 3158 6934 3204
rect 6980 3158 7037 3204
rect 6877 3110 7037 3158
rect 6877 3064 6934 3110
rect 6980 3064 7037 3110
rect 6877 3016 7037 3064
rect 6877 2970 6934 3016
rect 6980 2970 7037 3016
rect 6877 2922 7037 2970
rect 6877 2885 6934 2922
rect 4914 2818 5074 2866
rect 4914 2772 4971 2818
rect 5017 2772 5074 2818
rect 4914 2724 5074 2772
rect 4914 2678 4971 2724
rect 5017 2678 5074 2724
rect 4914 2630 5074 2678
rect 4914 2584 4971 2630
rect 5017 2584 5074 2630
rect 4914 2536 5074 2584
rect 4914 2490 4971 2536
rect 5017 2490 5074 2536
rect 4914 2442 5074 2490
rect 4914 2396 4971 2442
rect 5017 2396 5074 2442
rect 4914 2348 5074 2396
rect 4914 2302 4971 2348
rect 5017 2302 5074 2348
rect 4914 2254 5074 2302
rect 4914 2208 4971 2254
rect 5017 2208 5074 2254
rect 4914 2160 5074 2208
rect 4914 2114 4971 2160
rect 5017 2114 5074 2160
rect 4914 2066 5074 2114
rect 4914 2020 4971 2066
rect 5017 2020 5074 2066
rect 4914 1972 5074 2020
rect 4914 1926 4971 1972
rect 5017 1926 5074 1972
rect 4914 1878 5074 1926
rect 4914 1832 4971 1878
rect 5017 1832 5074 1878
rect 4914 1784 5074 1832
rect 4914 1738 4971 1784
rect 5017 1738 5074 1784
rect 4914 1690 5074 1738
rect 4914 1644 4971 1690
rect 5017 1644 5074 1690
rect 4914 1596 5074 1644
rect 4914 1559 4971 1596
rect 975 1550 4971 1559
rect 5017 1550 5074 1596
rect 872 1502 5074 1550
rect 872 1456 929 1502
rect 975 1456 1023 1502
rect 1069 1456 1117 1502
rect 1163 1456 1211 1502
rect 1257 1456 1305 1502
rect 1351 1456 1399 1502
rect 1445 1456 1493 1502
rect 1539 1456 1587 1502
rect 1633 1456 1681 1502
rect 1727 1456 1775 1502
rect 1821 1456 1869 1502
rect 1915 1456 1963 1502
rect 2009 1456 2057 1502
rect 2103 1456 2151 1502
rect 2197 1456 2245 1502
rect 2291 1456 2339 1502
rect 2385 1456 2433 1502
rect 2479 1456 2527 1502
rect 2573 1456 2621 1502
rect 2667 1456 2715 1502
rect 2761 1456 2809 1502
rect 2855 1456 2903 1502
rect 2949 1456 2997 1502
rect 3043 1456 3091 1502
rect 3137 1456 3185 1502
rect 3231 1456 3279 1502
rect 3325 1456 3373 1502
rect 3419 1456 3467 1502
rect 3513 1456 3561 1502
rect 3607 1456 3655 1502
rect 3701 1456 3749 1502
rect 3795 1456 3843 1502
rect 3889 1456 3937 1502
rect 3983 1456 4031 1502
rect 4077 1456 4125 1502
rect 4171 1456 4219 1502
rect 4265 1456 4313 1502
rect 4359 1456 4407 1502
rect 4453 1456 4501 1502
rect 4547 1456 4595 1502
rect 4641 1456 4689 1502
rect 4735 1456 4783 1502
rect 4829 1456 4877 1502
rect 4923 1456 4971 1502
rect 5017 1456 5074 1502
rect 872 1399 5074 1456
rect 5843 2876 6934 2885
rect 6980 2876 7037 2922
rect 5843 2828 7037 2876
rect 7396 5725 7442 6015
rect 7396 5189 7442 5551
rect 7396 4653 7442 5015
rect 7396 4117 7442 4479
rect 7396 3785 7442 3943
rect 7556 5725 7602 6015
rect 9189 5938 9265 5950
rect 9189 5935 9201 5938
rect 7753 5934 8301 5935
rect 7753 5888 7764 5934
rect 7810 5888 8244 5934
rect 8290 5888 8301 5934
rect 8713 5934 9201 5935
rect 8713 5888 8724 5934
rect 8770 5888 9201 5934
rect 9253 5886 9265 5938
rect 9201 5874 9265 5886
rect 7684 5782 9330 5828
rect 7684 5725 7730 5782
rect 7556 5189 7602 5551
rect 7669 5709 7684 5721
rect 7844 5725 7890 5736
rect 7730 5709 7745 5721
rect 7669 5657 7681 5709
rect 7733 5657 7745 5709
rect 7669 5605 7684 5657
rect 7730 5605 7745 5657
rect 7669 5553 7681 5605
rect 7733 5553 7745 5605
rect 7669 5551 7684 5553
rect 7730 5551 7745 5553
rect 7669 5541 7745 5551
rect 7829 5709 7844 5721
rect 8004 5725 8050 5736
rect 7890 5709 7905 5721
rect 7829 5657 7841 5709
rect 7893 5657 7905 5709
rect 7829 5605 7844 5657
rect 7890 5605 7905 5657
rect 7829 5553 7841 5605
rect 7893 5553 7905 5605
rect 7829 5551 7844 5553
rect 7890 5551 7905 5553
rect 7829 5541 7905 5551
rect 8164 5725 8210 5736
rect 7684 5540 7730 5541
rect 7844 5540 7890 5541
rect 8004 5494 8050 5551
rect 8149 5709 8164 5721
rect 8324 5725 8370 5782
rect 8210 5709 8225 5721
rect 8149 5657 8161 5709
rect 8213 5657 8225 5709
rect 8149 5605 8164 5657
rect 8210 5605 8225 5657
rect 8149 5553 8161 5605
rect 8213 5553 8225 5605
rect 8149 5551 8164 5553
rect 8210 5551 8225 5553
rect 8149 5541 8225 5551
rect 8484 5725 8530 5736
rect 8164 5540 8210 5541
rect 8324 5540 8370 5551
rect 8469 5709 8484 5721
rect 8644 5725 8690 5782
rect 8530 5709 8545 5721
rect 8469 5657 8481 5709
rect 8533 5657 8545 5709
rect 8469 5605 8484 5657
rect 8530 5605 8545 5657
rect 8469 5553 8481 5605
rect 8533 5553 8545 5605
rect 8469 5551 8484 5553
rect 8530 5551 8545 5553
rect 8469 5541 8545 5551
rect 8804 5725 8850 5736
rect 8484 5540 8530 5541
rect 8644 5540 8690 5551
rect 8789 5709 8804 5721
rect 8964 5725 9010 5736
rect 8850 5709 8865 5721
rect 8789 5657 8801 5709
rect 8853 5657 8865 5709
rect 8789 5605 8804 5657
rect 8850 5605 8865 5657
rect 8789 5553 8801 5605
rect 8853 5553 8865 5605
rect 8789 5551 8804 5553
rect 8850 5551 8865 5553
rect 8789 5541 8865 5551
rect 8949 5709 8964 5720
rect 9124 5725 9170 5736
rect 9010 5709 9025 5720
rect 8949 5657 8961 5709
rect 9013 5657 9025 5709
rect 8949 5605 8964 5657
rect 9010 5605 9025 5657
rect 8949 5553 8961 5605
rect 9013 5553 9025 5605
rect 8949 5551 8964 5553
rect 9010 5551 9025 5553
rect 8804 5540 8850 5541
rect 8949 5540 9025 5551
rect 9109 5709 9124 5721
rect 9284 5725 9330 5782
rect 9170 5709 9185 5721
rect 9109 5657 9121 5709
rect 9173 5657 9185 5709
rect 9109 5605 9124 5657
rect 9170 5605 9185 5657
rect 9109 5553 9121 5605
rect 9173 5553 9185 5605
rect 9109 5551 9124 5553
rect 9170 5551 9185 5553
rect 9109 5541 9185 5551
rect 9124 5540 9170 5541
rect 9284 5540 9330 5551
rect 9412 5725 9458 6015
rect 8964 5494 9010 5540
rect 8004 5448 9010 5494
rect 7753 5338 7764 5384
rect 7810 5338 7924 5384
rect 7970 5338 8244 5384
rect 8290 5338 8301 5384
rect 8496 5292 8542 5448
rect 9268 5402 9344 5414
rect 9268 5384 9280 5402
rect 8713 5338 8724 5384
rect 8770 5338 8884 5384
rect 8930 5338 9204 5384
rect 9250 5350 9280 5384
rect 9332 5350 9344 5402
rect 9250 5338 9344 5350
rect 7556 4653 7602 5015
rect 7684 5246 9330 5292
rect 7684 5189 7730 5246
rect 7844 5189 7890 5200
rect 7684 5004 7730 5015
rect 7829 5173 7844 5185
rect 8004 5189 8050 5200
rect 7890 5173 7905 5185
rect 7829 5121 7841 5173
rect 7893 5121 7905 5173
rect 7829 5069 7844 5121
rect 7890 5069 7905 5121
rect 7829 5017 7841 5069
rect 7893 5017 7905 5069
rect 7829 5015 7844 5017
rect 7890 5015 7905 5017
rect 7829 5005 7905 5015
rect 7989 5173 8004 5184
rect 8164 5189 8210 5200
rect 8050 5173 8065 5184
rect 7989 5121 8001 5173
rect 8053 5121 8065 5173
rect 7989 5069 8004 5121
rect 8050 5069 8065 5121
rect 7989 5017 8001 5069
rect 8053 5017 8065 5069
rect 7989 5015 8004 5017
rect 8050 5015 8065 5017
rect 7844 5004 7890 5005
rect 7989 5004 8065 5015
rect 8149 5173 8164 5185
rect 8324 5189 8370 5246
rect 8210 5173 8225 5185
rect 8149 5121 8161 5173
rect 8213 5121 8225 5173
rect 8149 5069 8164 5121
rect 8210 5069 8225 5121
rect 8149 5017 8161 5069
rect 8213 5017 8225 5069
rect 8149 5015 8164 5017
rect 8210 5015 8225 5017
rect 8149 5005 8225 5015
rect 8484 5189 8530 5200
rect 8164 5004 8210 5005
rect 8324 5004 8370 5015
rect 8469 5173 8484 5185
rect 8644 5189 8690 5246
rect 8530 5173 8545 5185
rect 8469 5121 8481 5173
rect 8533 5121 8545 5173
rect 8469 5069 8484 5121
rect 8530 5069 8545 5121
rect 8469 5017 8481 5069
rect 8533 5017 8545 5069
rect 8469 5015 8484 5017
rect 8530 5015 8545 5017
rect 8469 5005 8545 5015
rect 8804 5189 8850 5200
rect 8484 5004 8530 5005
rect 8644 5004 8690 5015
rect 8789 5173 8804 5185
rect 8964 5189 9010 5200
rect 8850 5173 8865 5185
rect 8789 5121 8801 5173
rect 8853 5121 8865 5173
rect 8789 5069 8804 5121
rect 8850 5069 8865 5121
rect 8789 5017 8801 5069
rect 8853 5017 8865 5069
rect 8789 5015 8804 5017
rect 8850 5015 8865 5017
rect 8789 5005 8865 5015
rect 9124 5189 9170 5200
rect 8804 5004 8850 5005
rect 8004 4958 8050 5004
rect 8964 4958 9010 5015
rect 9109 5173 9124 5185
rect 9284 5189 9330 5246
rect 9170 5173 9185 5185
rect 9109 5121 9121 5173
rect 9173 5121 9185 5173
rect 9109 5069 9124 5121
rect 9170 5069 9185 5121
rect 9109 5017 9121 5069
rect 9173 5017 9185 5069
rect 9109 5015 9124 5017
rect 9170 5015 9185 5017
rect 9109 5005 9185 5015
rect 9124 5004 9170 5005
rect 9284 5004 9330 5015
rect 9412 5189 9458 5551
rect 8004 4912 9010 4958
rect 7753 4817 7764 4863
rect 7810 4817 7924 4863
rect 7970 4817 8244 4863
rect 8290 4817 8301 4863
rect 8479 4756 8525 4912
rect 9071 4866 9147 4878
rect 9071 4863 9083 4866
rect 8713 4817 8724 4863
rect 8770 4817 8884 4863
rect 8930 4817 9083 4863
rect 9071 4814 9083 4817
rect 9135 4863 9147 4866
rect 9135 4817 9204 4863
rect 9250 4817 9261 4863
rect 9135 4814 9147 4817
rect 9071 4802 9147 4814
rect 7684 4710 9330 4756
rect 7684 4653 7730 4710
rect 7556 4117 7602 4479
rect 7669 4637 7684 4649
rect 7844 4653 7890 4664
rect 7730 4637 7745 4649
rect 7669 4585 7681 4637
rect 7733 4585 7745 4637
rect 7669 4533 7684 4585
rect 7730 4533 7745 4585
rect 7669 4481 7681 4533
rect 7733 4481 7745 4533
rect 7669 4479 7684 4481
rect 7730 4479 7745 4481
rect 7669 4469 7745 4479
rect 7829 4637 7844 4649
rect 8004 4653 8050 4664
rect 7890 4637 7905 4649
rect 7829 4585 7841 4637
rect 7893 4585 7905 4637
rect 7829 4533 7844 4585
rect 7890 4533 7905 4585
rect 7829 4481 7841 4533
rect 7893 4481 7905 4533
rect 7829 4479 7844 4481
rect 7890 4479 7905 4481
rect 7829 4469 7905 4479
rect 8164 4653 8210 4664
rect 7684 4468 7730 4469
rect 7844 4468 7890 4469
rect 8004 4422 8050 4479
rect 8149 4637 8164 4649
rect 8324 4653 8370 4710
rect 8210 4637 8225 4649
rect 8149 4585 8161 4637
rect 8213 4585 8225 4637
rect 8149 4533 8164 4585
rect 8210 4533 8225 4585
rect 8149 4481 8161 4533
rect 8213 4481 8225 4533
rect 8149 4479 8164 4481
rect 8210 4479 8225 4481
rect 8149 4469 8225 4479
rect 8484 4653 8530 4664
rect 8164 4468 8210 4469
rect 8324 4468 8370 4479
rect 8469 4637 8484 4649
rect 8644 4653 8690 4710
rect 8530 4637 8545 4649
rect 8469 4585 8481 4637
rect 8533 4585 8545 4637
rect 8469 4533 8484 4585
rect 8530 4533 8545 4585
rect 8469 4481 8481 4533
rect 8533 4481 8545 4533
rect 8469 4479 8484 4481
rect 8530 4479 8545 4481
rect 8469 4469 8545 4479
rect 8804 4653 8850 4664
rect 8484 4468 8530 4469
rect 8644 4468 8690 4479
rect 8789 4637 8804 4649
rect 8964 4653 9010 4664
rect 8850 4637 8865 4649
rect 8789 4585 8801 4637
rect 8853 4585 8865 4637
rect 8789 4533 8804 4585
rect 8850 4533 8865 4585
rect 8789 4481 8801 4533
rect 8853 4481 8865 4533
rect 8789 4479 8804 4481
rect 8850 4479 8865 4481
rect 8789 4469 8865 4479
rect 8949 4637 8964 4649
rect 9124 4653 9170 4664
rect 9010 4637 9025 4649
rect 8949 4585 8961 4637
rect 9013 4585 9025 4637
rect 8949 4533 8964 4585
rect 9010 4533 9025 4585
rect 8949 4481 8961 4533
rect 9013 4481 9025 4533
rect 8949 4479 8964 4481
rect 9010 4479 9025 4481
rect 8804 4468 8850 4469
rect 8949 4468 9025 4479
rect 9109 4637 9124 4649
rect 9284 4653 9330 4710
rect 9170 4637 9185 4649
rect 9109 4585 9121 4637
rect 9173 4585 9185 4637
rect 9109 4533 9124 4585
rect 9170 4533 9185 4585
rect 9109 4481 9121 4533
rect 9173 4481 9185 4533
rect 9109 4479 9124 4481
rect 9170 4479 9185 4481
rect 9109 4469 9185 4479
rect 9124 4468 9170 4469
rect 9284 4468 9330 4479
rect 9412 4653 9458 5015
rect 8964 4422 9010 4468
rect 8004 4376 9010 4422
rect 7753 4283 7764 4329
rect 7810 4283 7924 4329
rect 7970 4283 8244 4329
rect 8290 4283 8301 4329
rect 8479 4220 8525 4376
rect 9189 4332 9265 4344
rect 9189 4329 9201 4332
rect 8713 4283 8724 4329
rect 8770 4283 8884 4329
rect 8930 4283 9201 4329
rect 9189 4280 9201 4283
rect 9253 4280 9265 4332
rect 9189 4268 9265 4280
rect 7556 3785 7602 3943
rect 7684 4174 9330 4220
rect 7684 4117 7730 4174
rect 7844 4117 7890 4128
rect 7684 3932 7730 3943
rect 7829 4101 7844 4113
rect 8004 4117 8050 4128
rect 7890 4101 7905 4113
rect 7829 4049 7841 4101
rect 7893 4049 7905 4101
rect 7829 3997 7844 4049
rect 7890 3997 7905 4049
rect 7829 3945 7841 3997
rect 7893 3945 7905 3997
rect 7829 3943 7844 3945
rect 7890 3943 7905 3945
rect 7829 3933 7905 3943
rect 7989 4101 8004 4112
rect 8164 4117 8210 4128
rect 8050 4101 8065 4112
rect 7989 4049 8001 4101
rect 8053 4049 8065 4101
rect 7989 3997 8004 4049
rect 8050 3997 8065 4049
rect 7989 3945 8001 3997
rect 8053 3945 8065 3997
rect 7989 3943 8004 3945
rect 8050 3943 8065 3945
rect 7844 3932 7890 3933
rect 7989 3932 8065 3943
rect 8149 4101 8164 4113
rect 8324 4117 8370 4174
rect 8210 4101 8225 4113
rect 8149 4049 8161 4101
rect 8213 4049 8225 4101
rect 8149 3997 8164 4049
rect 8210 3997 8225 4049
rect 8149 3945 8161 3997
rect 8213 3945 8225 3997
rect 8149 3943 8164 3945
rect 8210 3943 8225 3945
rect 8149 3933 8225 3943
rect 8484 4117 8530 4128
rect 8164 3932 8210 3933
rect 8324 3932 8370 3943
rect 8469 4101 8484 4113
rect 8644 4117 8690 4174
rect 8530 4101 8545 4113
rect 8469 4049 8481 4101
rect 8533 4049 8545 4101
rect 8469 3997 8484 4049
rect 8530 3997 8545 4049
rect 8469 3945 8481 3997
rect 8533 3945 8545 3997
rect 8469 3943 8484 3945
rect 8530 3943 8545 3945
rect 8469 3933 8545 3943
rect 8804 4117 8850 4128
rect 8484 3932 8530 3933
rect 8644 3932 8690 3943
rect 8789 4101 8804 4113
rect 8964 4117 9010 4128
rect 8850 4101 8865 4113
rect 8789 4049 8801 4101
rect 8853 4049 8865 4101
rect 8789 3997 8804 4049
rect 8850 3997 8865 4049
rect 8789 3945 8801 3997
rect 8853 3945 8865 3997
rect 8789 3943 8804 3945
rect 8850 3943 8865 3945
rect 8789 3933 8865 3943
rect 9124 4117 9170 4128
rect 8804 3932 8850 3933
rect 8004 3886 8050 3932
rect 8964 3886 9010 3943
rect 9109 4101 9124 4113
rect 9284 4117 9330 4174
rect 9170 4101 9185 4113
rect 9109 4049 9121 4101
rect 9173 4049 9185 4101
rect 9109 3997 9124 4049
rect 9170 3997 9185 4049
rect 9109 3945 9121 3997
rect 9173 3945 9185 3997
rect 9109 3943 9124 3945
rect 9170 3943 9185 3945
rect 9109 3933 9185 3943
rect 9124 3932 9170 3933
rect 9284 3932 9330 3943
rect 9412 4117 9458 4479
rect 8004 3840 9010 3886
rect 7396 3739 7476 3785
rect 7522 3739 7602 3785
rect 7753 3747 7764 3793
rect 7810 3747 7924 3793
rect 7970 3747 8244 3793
rect 8290 3747 8301 3793
rect 7396 3581 7442 3739
rect 7396 3045 7442 3407
rect 7396 2860 7442 2871
rect 7556 3581 7602 3739
rect 8479 3684 8525 3840
rect 9268 3796 9344 3808
rect 9268 3793 9280 3796
rect 8713 3747 8724 3793
rect 8770 3747 8884 3793
rect 8930 3791 9280 3793
rect 8930 3747 9204 3791
rect 9191 3745 9204 3747
rect 9250 3745 9280 3791
rect 9268 3744 9280 3745
rect 9332 3744 9344 3796
rect 9268 3732 9344 3744
rect 9412 3785 9458 3943
rect 9572 5725 9618 6015
rect 9969 6005 10036 6015
rect 9572 5189 9618 5551
rect 9572 4653 9618 5015
rect 9572 4117 9618 4479
rect 9572 3785 9618 3943
rect 9412 3739 9492 3785
rect 9538 3739 9618 3785
rect 7556 3045 7602 3407
rect 7684 3638 9330 3684
rect 7684 3581 7730 3638
rect 7844 3585 7890 3592
rect 7684 3396 7730 3407
rect 7829 3581 7905 3585
rect 7829 3573 7844 3581
rect 7890 3573 7905 3581
rect 7829 3521 7841 3573
rect 7893 3521 7905 3573
rect 7829 3469 7844 3521
rect 7890 3469 7905 3521
rect 7829 3417 7841 3469
rect 7893 3417 7905 3469
rect 7829 3407 7844 3417
rect 7890 3407 7905 3417
rect 7829 3405 7905 3407
rect 8004 3581 8050 3592
rect 8164 3585 8210 3592
rect 7844 3396 7890 3405
rect 8004 3350 8050 3407
rect 8149 3581 8225 3585
rect 8149 3573 8164 3581
rect 8210 3573 8225 3581
rect 8149 3521 8161 3573
rect 8213 3521 8225 3573
rect 8149 3469 8164 3521
rect 8210 3469 8225 3521
rect 8149 3417 8161 3469
rect 8213 3417 8225 3469
rect 8149 3407 8164 3417
rect 8210 3407 8225 3417
rect 8149 3405 8225 3407
rect 8324 3581 8370 3638
rect 8484 3585 8530 3592
rect 8164 3396 8210 3405
rect 8324 3396 8370 3407
rect 8469 3581 8545 3585
rect 8469 3573 8484 3581
rect 8530 3573 8545 3581
rect 8469 3521 8481 3573
rect 8533 3521 8545 3573
rect 8469 3469 8484 3521
rect 8530 3469 8545 3521
rect 8469 3417 8481 3469
rect 8533 3417 8545 3469
rect 8469 3407 8484 3417
rect 8530 3407 8545 3417
rect 8469 3405 8545 3407
rect 8644 3581 8690 3638
rect 8804 3585 8850 3592
rect 8484 3396 8530 3405
rect 8644 3396 8690 3407
rect 8789 3581 8865 3585
rect 8789 3573 8804 3581
rect 8850 3573 8865 3581
rect 8964 3581 9010 3592
rect 9124 3585 9170 3592
rect 8789 3521 8801 3573
rect 8853 3521 8865 3573
rect 8789 3469 8804 3521
rect 8850 3469 8865 3521
rect 8789 3417 8801 3469
rect 8853 3417 8865 3469
rect 8789 3407 8804 3417
rect 8850 3407 8865 3417
rect 8789 3405 8865 3407
rect 8949 3565 8964 3577
rect 9109 3581 9185 3585
rect 9010 3565 9025 3577
rect 8949 3513 8961 3565
rect 9013 3513 9025 3565
rect 8949 3461 8964 3513
rect 9010 3461 9025 3513
rect 8949 3409 8961 3461
rect 9013 3409 9025 3461
rect 8949 3407 8964 3409
rect 9010 3407 9025 3409
rect 8804 3396 8850 3405
rect 8949 3396 9025 3407
rect 9109 3573 9124 3581
rect 9170 3573 9185 3581
rect 9109 3521 9121 3573
rect 9173 3521 9185 3573
rect 9109 3469 9124 3521
rect 9170 3469 9185 3521
rect 9109 3417 9121 3469
rect 9173 3417 9185 3469
rect 9109 3407 9124 3417
rect 9170 3407 9185 3417
rect 9109 3405 9185 3407
rect 9284 3581 9330 3638
rect 9124 3396 9170 3405
rect 9284 3396 9330 3407
rect 9412 3581 9458 3739
rect 8964 3350 9010 3396
rect 8004 3304 9010 3350
rect 7753 3211 7764 3257
rect 7810 3211 7924 3257
rect 7970 3211 8244 3257
rect 8290 3211 8301 3257
rect 8479 3148 8525 3304
rect 9268 3281 9344 3293
rect 9268 3257 9280 3281
rect 8713 3211 8724 3257
rect 8770 3211 8884 3257
rect 8930 3255 9280 3257
rect 8930 3211 9204 3255
rect 9193 3209 9204 3211
rect 9250 3229 9280 3255
rect 9332 3229 9344 3281
rect 9250 3211 9344 3229
rect 9250 3209 9261 3211
rect 7556 2860 7602 2871
rect 7684 3102 9330 3148
rect 7684 3045 7730 3102
rect 7844 3049 7890 3056
rect 7684 2860 7730 2871
rect 7829 3045 7905 3049
rect 7829 3037 7844 3045
rect 7890 3037 7905 3045
rect 8004 3045 8050 3056
rect 8164 3049 8210 3056
rect 7829 2985 7841 3037
rect 7893 2985 7905 3037
rect 7829 2933 7844 2985
rect 7890 2933 7905 2985
rect 7829 2881 7841 2933
rect 7893 2881 7905 2933
rect 7829 2871 7844 2881
rect 7890 2871 7905 2881
rect 7829 2869 7905 2871
rect 7989 3029 8004 3040
rect 8149 3045 8225 3049
rect 8050 3029 8065 3040
rect 7989 2977 8001 3029
rect 8053 2977 8065 3029
rect 7989 2925 8004 2977
rect 8050 2925 8065 2977
rect 7989 2873 8001 2925
rect 8053 2873 8065 2925
rect 7989 2871 8004 2873
rect 8050 2871 8065 2873
rect 7844 2860 7890 2869
rect 7989 2860 8065 2871
rect 8149 3037 8164 3045
rect 8210 3037 8225 3045
rect 8149 2985 8161 3037
rect 8213 2985 8225 3037
rect 8149 2933 8164 2985
rect 8210 2933 8225 2985
rect 8149 2881 8161 2933
rect 8213 2881 8225 2933
rect 8149 2871 8164 2881
rect 8210 2871 8225 2881
rect 8149 2869 8225 2871
rect 8324 3045 8370 3102
rect 8484 3049 8530 3056
rect 8164 2860 8210 2869
rect 8324 2860 8370 2871
rect 8469 3045 8545 3049
rect 8469 3037 8484 3045
rect 8530 3037 8545 3045
rect 8469 2985 8481 3037
rect 8533 2985 8545 3037
rect 8469 2933 8484 2985
rect 8530 2933 8545 2985
rect 8469 2881 8481 2933
rect 8533 2881 8545 2933
rect 8469 2871 8484 2881
rect 8530 2871 8545 2881
rect 8469 2869 8545 2871
rect 8644 3045 8690 3102
rect 8804 3049 8850 3056
rect 8484 2860 8530 2869
rect 8644 2860 8690 2871
rect 8789 3045 8865 3049
rect 8789 3037 8804 3045
rect 8850 3037 8865 3045
rect 8789 2985 8801 3037
rect 8853 2985 8865 3037
rect 8789 2933 8804 2985
rect 8850 2933 8865 2985
rect 8789 2881 8801 2933
rect 8853 2881 8865 2933
rect 8789 2871 8804 2881
rect 8850 2871 8865 2881
rect 8789 2869 8865 2871
rect 8964 3045 9010 3056
rect 9124 3049 9170 3056
rect 8804 2860 8850 2869
rect 5843 2782 5900 2828
rect 5946 2782 5994 2828
rect 6040 2782 6088 2828
rect 6134 2782 6182 2828
rect 6228 2782 6276 2828
rect 6322 2782 6370 2828
rect 6416 2782 6464 2828
rect 6510 2782 6558 2828
rect 6604 2782 6652 2828
rect 6698 2782 6746 2828
rect 6792 2782 6840 2828
rect 6886 2782 6934 2828
rect 6980 2782 7037 2828
rect 5843 2734 7037 2782
rect 8004 2814 8050 2860
rect 8964 2814 9010 2871
rect 9109 3045 9185 3049
rect 9109 3037 9124 3045
rect 9170 3037 9185 3045
rect 9109 2985 9121 3037
rect 9173 2985 9185 3037
rect 9109 2933 9124 2985
rect 9170 2933 9185 2985
rect 9109 2881 9121 2933
rect 9173 2881 9185 2933
rect 9109 2871 9124 2881
rect 9170 2871 9185 2881
rect 9109 2869 9185 2871
rect 9284 3045 9330 3102
rect 9124 2860 9170 2869
rect 9284 2860 9330 2871
rect 9412 3045 9458 3407
rect 9412 2860 9458 2871
rect 9572 3581 9618 3739
rect 9572 3045 9618 3407
rect 9572 2860 9618 2871
rect 9979 5978 10036 6005
rect 10082 6017 10085 6024
rect 10137 6017 10149 6069
rect 11639 6094 17840 6106
rect 10082 6005 10149 6017
rect 10278 6044 10458 6054
rect 10278 6042 10748 6044
rect 10082 5978 10139 6005
rect 9979 5930 10139 5978
rect 9979 5884 10036 5930
rect 10082 5884 10139 5930
rect 9979 5836 10139 5884
rect 10278 5990 10290 6042
rect 10342 5990 10394 6042
rect 10446 5990 10748 6042
rect 10278 5938 10748 5990
rect 10278 5886 10290 5938
rect 10342 5886 10394 5938
rect 10446 5886 10748 5938
rect 10278 5884 10748 5886
rect 11639 6042 11651 6094
rect 11703 6042 11755 6094
rect 11807 6042 17568 6094
rect 17620 6042 17672 6094
rect 17724 6042 17776 6094
rect 17828 6042 17840 6094
rect 11639 5990 17840 6042
rect 11639 5938 11651 5990
rect 11703 5938 11755 5990
rect 11807 5938 17568 5990
rect 17620 5938 17672 5990
rect 17724 5938 17776 5990
rect 17828 5938 17840 5990
rect 11639 5886 17840 5938
rect 10278 5874 10458 5884
rect 9979 5790 10036 5836
rect 10082 5790 10139 5836
rect 11639 5834 11651 5886
rect 11703 5834 11755 5886
rect 11807 5834 17568 5886
rect 17620 5834 17672 5886
rect 17724 5834 17776 5886
rect 17828 5834 17840 5886
rect 11639 5822 17840 5834
rect 9979 5742 10139 5790
rect 9979 5696 10036 5742
rect 10082 5696 10139 5742
rect 18076 5811 18396 6506
rect 18576 5811 18896 6506
rect 19076 5811 19396 6506
rect 19576 5811 19896 6506
rect 20076 5811 20396 6506
rect 20576 5811 20896 6506
rect 21076 5811 21396 6506
rect 21576 5811 21896 6506
rect 22076 5811 22396 6506
rect 22856 5811 23176 6506
rect 28590 5811 28910 6506
rect 31598 5811 31918 6506
rect 9979 5648 10139 5696
rect 9979 5602 10036 5648
rect 10082 5602 10139 5648
rect 9979 5554 10139 5602
rect 9979 5508 10036 5554
rect 10082 5508 10139 5554
rect 14686 5713 14866 5721
rect 14686 5709 15154 5713
rect 14686 5657 14698 5709
rect 14750 5657 14802 5709
rect 14854 5657 15154 5709
rect 14686 5605 15154 5657
rect 14686 5553 14698 5605
rect 14750 5553 14802 5605
rect 14854 5553 15154 5605
rect 18076 5701 31918 5811
rect 18076 5655 18206 5701
rect 18252 5655 18300 5701
rect 18346 5655 18394 5701
rect 18440 5655 18488 5701
rect 18534 5655 18582 5701
rect 18628 5655 18676 5701
rect 18722 5655 18770 5701
rect 18816 5655 18864 5701
rect 18910 5655 18958 5701
rect 19004 5655 19052 5701
rect 19098 5655 19146 5701
rect 19192 5655 19240 5701
rect 19286 5655 19334 5701
rect 19380 5655 19428 5701
rect 19474 5655 19522 5701
rect 19568 5655 19616 5701
rect 19662 5655 19710 5701
rect 19756 5655 19804 5701
rect 19850 5655 19898 5701
rect 19944 5655 19992 5701
rect 20038 5655 20086 5701
rect 20132 5655 20180 5701
rect 20226 5655 20274 5701
rect 20320 5655 20368 5701
rect 20414 5655 20462 5701
rect 20508 5655 20556 5701
rect 20602 5655 20650 5701
rect 20696 5655 20744 5701
rect 20790 5655 20838 5701
rect 20884 5655 20932 5701
rect 20978 5655 21026 5701
rect 21072 5655 21120 5701
rect 21166 5655 21214 5701
rect 21260 5655 21308 5701
rect 21354 5655 21402 5701
rect 21448 5655 21496 5701
rect 21542 5655 21590 5701
rect 21636 5655 21684 5701
rect 21730 5655 21778 5701
rect 21824 5655 21872 5701
rect 21918 5655 21966 5701
rect 22012 5655 22060 5701
rect 22106 5655 22154 5701
rect 22200 5655 22248 5701
rect 22294 5655 22342 5701
rect 22388 5655 22436 5701
rect 22482 5655 22530 5701
rect 22576 5655 22624 5701
rect 22670 5655 22718 5701
rect 22764 5655 22812 5701
rect 22858 5655 22906 5701
rect 22952 5655 23000 5701
rect 23046 5655 23094 5701
rect 23140 5655 23188 5701
rect 23234 5655 23282 5701
rect 23328 5655 23376 5701
rect 23422 5655 23470 5701
rect 23516 5655 23564 5701
rect 23610 5655 23658 5701
rect 23704 5655 23752 5701
rect 23798 5655 23846 5701
rect 23892 5655 23940 5701
rect 23986 5655 24034 5701
rect 24080 5655 24128 5701
rect 24174 5655 24222 5701
rect 24268 5655 24316 5701
rect 24362 5655 24410 5701
rect 24456 5655 24504 5701
rect 24550 5655 24598 5701
rect 24644 5655 24692 5701
rect 24738 5655 24786 5701
rect 24832 5655 24880 5701
rect 24926 5655 24974 5701
rect 25020 5655 25068 5701
rect 25114 5655 25162 5701
rect 25208 5655 25256 5701
rect 25302 5655 25350 5701
rect 25396 5655 25444 5701
rect 25490 5655 25538 5701
rect 25584 5655 25632 5701
rect 25678 5655 25726 5701
rect 25772 5655 25820 5701
rect 25866 5655 25914 5701
rect 25960 5655 26008 5701
rect 26054 5655 26102 5701
rect 26148 5655 26196 5701
rect 26242 5655 26290 5701
rect 26336 5655 26384 5701
rect 26430 5655 26478 5701
rect 26524 5655 26572 5701
rect 26618 5655 26666 5701
rect 26712 5655 26760 5701
rect 26806 5655 26854 5701
rect 26900 5655 26948 5701
rect 26994 5655 27042 5701
rect 27088 5655 27136 5701
rect 27182 5655 27230 5701
rect 27276 5655 27324 5701
rect 27370 5655 27418 5701
rect 27464 5655 27512 5701
rect 27558 5655 27606 5701
rect 27652 5655 27700 5701
rect 27746 5655 27794 5701
rect 27840 5655 27888 5701
rect 27934 5655 27982 5701
rect 28028 5655 28076 5701
rect 28122 5655 28170 5701
rect 28216 5655 28264 5701
rect 28310 5655 28358 5701
rect 28404 5655 28452 5701
rect 28498 5655 28546 5701
rect 28592 5655 28640 5701
rect 28686 5655 28734 5701
rect 28780 5655 28828 5701
rect 28874 5655 28922 5701
rect 28968 5655 29016 5701
rect 29062 5655 29110 5701
rect 29156 5655 29204 5701
rect 29250 5655 29298 5701
rect 29344 5655 29392 5701
rect 29438 5655 29486 5701
rect 29532 5655 29580 5701
rect 29626 5655 29674 5701
rect 29720 5655 29768 5701
rect 29814 5655 29862 5701
rect 29908 5655 29956 5701
rect 30002 5655 30050 5701
rect 30096 5655 30144 5701
rect 30190 5655 30238 5701
rect 30284 5655 30332 5701
rect 30378 5655 30426 5701
rect 30472 5655 30520 5701
rect 30566 5655 30614 5701
rect 30660 5655 30708 5701
rect 30754 5655 30802 5701
rect 30848 5655 30896 5701
rect 30942 5655 30990 5701
rect 31036 5655 31084 5701
rect 31130 5655 31178 5701
rect 31224 5655 31272 5701
rect 31318 5655 31366 5701
rect 31412 5655 31460 5701
rect 31506 5655 31554 5701
rect 31600 5655 31648 5701
rect 31694 5655 31742 5701
rect 31788 5655 31918 5701
rect 18076 5607 31918 5655
rect 18076 5561 18206 5607
rect 18252 5561 23000 5607
rect 23046 5561 28734 5607
rect 28780 5561 31742 5607
rect 31788 5561 31918 5607
rect 14686 5541 14866 5553
rect 9979 5460 10139 5508
rect 9979 5414 10036 5460
rect 10082 5414 10139 5460
rect 18076 5513 31918 5561
rect 18076 5467 18206 5513
rect 18252 5491 23000 5513
rect 18252 5467 18396 5491
rect 9979 5366 10139 5414
rect 9979 5320 10036 5366
rect 10082 5320 10139 5366
rect 9979 5272 10139 5320
rect 10544 5446 10724 5456
rect 17334 5446 17514 5456
rect 10544 5444 17514 5446
rect 10544 5392 10556 5444
rect 10608 5392 10660 5444
rect 10712 5392 17346 5444
rect 17398 5392 17450 5444
rect 17502 5392 17514 5444
rect 10544 5340 17514 5392
rect 10544 5288 10556 5340
rect 10608 5288 10660 5340
rect 10712 5288 17346 5340
rect 17398 5288 17450 5340
rect 17502 5288 17514 5340
rect 10544 5286 17514 5288
rect 10544 5276 10724 5286
rect 17334 5276 17514 5286
rect 18076 5419 18396 5467
rect 18076 5373 18206 5419
rect 18252 5373 18396 5419
rect 18076 5325 18396 5373
rect 18076 5279 18206 5325
rect 18252 5279 18396 5325
rect 9979 5226 10036 5272
rect 10082 5226 10139 5272
rect 9979 5178 10139 5226
rect 9979 5132 10036 5178
rect 10082 5132 10139 5178
rect 9979 5084 10139 5132
rect 9979 5038 10036 5084
rect 10082 5038 10139 5084
rect 9979 4990 10139 5038
rect 9979 4944 10036 4990
rect 10082 4944 10139 4990
rect 9979 4896 10139 4944
rect 9979 4850 10036 4896
rect 10082 4850 10139 4896
rect 9979 4802 10139 4850
rect 9979 4756 10036 4802
rect 10082 4756 10139 4802
rect 9979 4708 10139 4756
rect 9979 4662 10036 4708
rect 10082 4662 10139 4708
rect 9979 4614 10139 4662
rect 9979 4568 10036 4614
rect 10082 4569 10139 4614
rect 18076 5231 18396 5279
rect 18076 5185 18206 5231
rect 18252 5185 18396 5231
rect 18076 5137 18396 5185
rect 18076 5091 18206 5137
rect 18252 5091 18396 5137
rect 18076 5043 18396 5091
rect 18076 4997 18206 5043
rect 18252 4997 18396 5043
rect 18076 4949 18396 4997
rect 18076 4903 18206 4949
rect 18252 4903 18396 4949
rect 18076 4855 18396 4903
rect 18076 4809 18206 4855
rect 18252 4809 18396 4855
rect 18076 4761 18396 4809
rect 18076 4715 18206 4761
rect 18252 4715 18396 4761
rect 18076 4667 18396 4715
rect 18076 4621 18206 4667
rect 18252 4621 18396 4667
rect 18076 4573 18396 4621
rect 10082 4568 17694 4569
rect 9979 4520 17694 4568
rect 9979 4474 10036 4520
rect 10082 4474 17694 4520
rect 9979 4469 17694 4474
rect 9979 4426 12014 4469
rect 9979 4380 10036 4426
rect 10082 4423 12014 4426
rect 12060 4423 12108 4469
rect 12154 4423 12202 4469
rect 12248 4423 12296 4469
rect 12342 4423 12390 4469
rect 12436 4423 12484 4469
rect 12530 4423 12578 4469
rect 12624 4423 12672 4469
rect 12718 4423 12766 4469
rect 12812 4423 12860 4469
rect 12906 4423 12954 4469
rect 13000 4423 13048 4469
rect 13094 4423 13142 4469
rect 13188 4423 13236 4469
rect 13282 4423 13330 4469
rect 13376 4423 13424 4469
rect 13470 4423 13518 4469
rect 13564 4423 13612 4469
rect 13658 4423 13706 4469
rect 13752 4423 13800 4469
rect 13846 4423 13894 4469
rect 13940 4423 13988 4469
rect 14034 4423 14082 4469
rect 14128 4423 14176 4469
rect 14222 4423 14270 4469
rect 14316 4423 14364 4469
rect 14410 4423 14458 4469
rect 14504 4423 14552 4469
rect 14598 4423 14646 4469
rect 14692 4423 14740 4469
rect 14786 4423 14834 4469
rect 14880 4423 14928 4469
rect 14974 4423 15022 4469
rect 15068 4423 15116 4469
rect 15162 4423 15210 4469
rect 15256 4423 15304 4469
rect 15350 4423 15398 4469
rect 15444 4423 15492 4469
rect 15538 4423 15586 4469
rect 15632 4423 15680 4469
rect 15726 4423 15774 4469
rect 15820 4423 15868 4469
rect 15914 4423 15962 4469
rect 16008 4423 16056 4469
rect 16102 4423 16150 4469
rect 16196 4423 16244 4469
rect 16290 4423 16338 4469
rect 16384 4423 16432 4469
rect 16478 4423 16526 4469
rect 16572 4423 16620 4469
rect 16666 4423 16714 4469
rect 16760 4423 16808 4469
rect 16854 4423 16902 4469
rect 16948 4423 16996 4469
rect 17042 4423 17090 4469
rect 17136 4423 17184 4469
rect 17230 4423 17278 4469
rect 17324 4423 17372 4469
rect 17418 4423 17466 4469
rect 17512 4423 17560 4469
rect 17606 4423 17694 4469
rect 10082 4380 17694 4423
rect 9979 4375 17694 4380
rect 9979 4332 12014 4375
rect 9979 4286 10036 4332
rect 10082 4329 12014 4332
rect 12060 4329 17560 4375
rect 17606 4329 17694 4375
rect 10082 4286 17694 4329
rect 9979 4281 17694 4286
rect 9979 4249 12014 4281
rect 9979 4238 10139 4249
rect 9979 4192 10036 4238
rect 10082 4192 10139 4238
rect 9979 4144 10139 4192
rect 9979 4098 10036 4144
rect 10082 4098 10139 4144
rect 9979 4050 10139 4098
rect 9979 4004 10036 4050
rect 10082 4004 10139 4050
rect 9979 3956 10139 4004
rect 9979 3910 10036 3956
rect 10082 3910 10139 3956
rect 9979 3862 10139 3910
rect 9979 3816 10036 3862
rect 10082 3816 10139 3862
rect 9979 3768 10139 3816
rect 9979 3722 10036 3768
rect 10082 3722 10139 3768
rect 9979 3674 10139 3722
rect 9979 3628 10036 3674
rect 10082 3628 10139 3674
rect 9979 3580 10139 3628
rect 9979 3534 10036 3580
rect 10082 3541 10139 3580
rect 11926 4235 12014 4249
rect 12060 4249 17560 4281
rect 12060 4235 12246 4249
rect 11926 4187 12246 4235
rect 11926 4141 12014 4187
rect 12060 4141 12246 4187
rect 11926 4093 12246 4141
rect 11926 4047 12014 4093
rect 12060 4047 12246 4093
rect 11926 3999 12246 4047
rect 11926 3953 12014 3999
rect 12060 3953 12246 3999
rect 11926 3905 12246 3953
rect 11926 3859 12014 3905
rect 12060 3859 12246 3905
rect 11926 3811 12246 3859
rect 11926 3765 12014 3811
rect 12060 3765 12246 3811
rect 11926 3717 12246 3765
rect 11926 3671 12014 3717
rect 12060 3671 12246 3717
rect 11926 3623 12246 3671
rect 11926 3577 12014 3623
rect 12060 3577 12246 3623
rect 11926 3541 12246 3577
rect 10082 3534 12246 3541
rect 9979 3529 12246 3534
rect 9979 3486 12014 3529
rect 9979 3440 10036 3486
rect 10082 3483 12014 3486
rect 12060 3483 12246 3529
rect 10082 3440 12246 3483
rect 9979 3435 12246 3440
rect 9979 3392 12014 3435
rect 9979 3346 10036 3392
rect 10082 3389 12014 3392
rect 12060 3389 12246 3435
rect 10082 3346 12246 3389
rect 9979 3341 12246 3346
rect 9979 3298 12014 3341
rect 9979 3252 10036 3298
rect 10082 3295 12014 3298
rect 12060 3295 12246 3341
rect 10082 3252 12246 3295
rect 9979 3247 12246 3252
rect 9979 3221 12014 3247
rect 9979 3204 10139 3221
rect 9979 3158 10036 3204
rect 10082 3158 10139 3204
rect 9979 3110 10139 3158
rect 9979 3064 10036 3110
rect 10082 3064 10139 3110
rect 9979 3016 10139 3064
rect 9979 2970 10036 3016
rect 10082 2970 10139 3016
rect 9979 2922 10139 2970
rect 9979 2876 10036 2922
rect 10082 2885 10139 2922
rect 11926 3201 12014 3221
rect 12060 3201 12246 3247
rect 11926 3153 12246 3201
rect 11926 3107 12014 3153
rect 12060 3107 12246 3153
rect 11926 3059 12246 3107
rect 11926 3013 12014 3059
rect 12060 3013 12246 3059
rect 11926 2965 12246 3013
rect 11926 2919 12014 2965
rect 12060 2919 12246 2965
rect 11926 2885 12246 2919
rect 10082 2876 12246 2885
rect 9979 2871 12246 2876
rect 8004 2768 9010 2814
rect 9979 2828 12014 2871
rect 9979 2782 10036 2828
rect 10082 2782 10130 2828
rect 10176 2782 10224 2828
rect 10270 2782 10318 2828
rect 10364 2782 10412 2828
rect 10458 2782 10506 2828
rect 10552 2782 10600 2828
rect 10646 2782 10694 2828
rect 10740 2782 10788 2828
rect 10834 2782 10882 2828
rect 10928 2782 10976 2828
rect 11022 2782 11070 2828
rect 11116 2825 12014 2828
rect 12060 2825 12246 2871
rect 11116 2782 12246 2825
rect 9979 2777 12246 2782
rect 5843 2688 5900 2734
rect 5946 2725 7037 2734
rect 9979 2734 12014 2777
rect 9979 2725 11070 2734
rect 5946 2688 6003 2725
rect 5843 2640 6003 2688
rect 5843 2594 5900 2640
rect 5946 2594 6003 2640
rect 5843 2546 6003 2594
rect 5843 2500 5900 2546
rect 5946 2500 6003 2546
rect 5843 2452 6003 2500
rect 5843 2406 5900 2452
rect 5946 2406 6003 2452
rect 5843 2358 6003 2406
rect 5843 2312 5900 2358
rect 5946 2312 6003 2358
rect 5843 2264 6003 2312
rect 5843 2218 5900 2264
rect 5946 2218 6003 2264
rect 5843 2170 6003 2218
rect 5843 2124 5900 2170
rect 5946 2124 6003 2170
rect 5843 2076 6003 2124
rect 5843 2030 5900 2076
rect 5946 2030 6003 2076
rect 5843 1982 6003 2030
rect 5843 1936 5900 1982
rect 5946 1936 6003 1982
rect 5843 1888 6003 1936
rect 5843 1842 5900 1888
rect 5946 1842 6003 1888
rect 5843 1794 6003 1842
rect 5843 1748 5900 1794
rect 5946 1748 6003 1794
rect 5843 1700 6003 1748
rect 5843 1654 5900 1700
rect 5946 1654 6003 1700
rect 5843 1606 6003 1654
rect 5843 1560 5900 1606
rect 5946 1560 6003 1606
rect 5843 1512 6003 1560
rect 5843 1466 5900 1512
rect 5946 1466 6003 1512
rect 5843 1418 6003 1466
rect 5843 1372 5900 1418
rect 5946 1381 6003 1418
rect 6149 2416 6195 2725
rect 6149 2033 6195 2242
rect 6309 2416 6355 2725
rect 7913 2675 7924 2721
rect 7970 2709 8884 2721
rect 8930 2709 8945 2721
rect 7970 2675 8881 2709
rect 8869 2657 8881 2675
rect 8933 2657 8945 2709
rect 7384 2639 7564 2653
rect 8869 2645 8945 2657
rect 7384 2587 7394 2639
rect 7446 2587 7498 2639
rect 7550 2587 7564 2639
rect 7384 2535 7564 2587
rect 7384 2519 7394 2535
rect 6597 2473 6677 2519
rect 6723 2473 6837 2519
rect 6883 2473 6963 2519
rect 6309 2033 6355 2242
rect 6437 2416 6483 2427
rect 6597 2416 6643 2473
rect 6437 2185 6483 2242
rect 6582 2400 6597 2412
rect 6757 2416 6803 2427
rect 6643 2400 6658 2412
rect 6582 2348 6594 2400
rect 6646 2348 6658 2400
rect 6582 2296 6597 2348
rect 6643 2296 6658 2348
rect 6582 2244 6594 2296
rect 6646 2244 6658 2296
rect 6582 2242 6597 2244
rect 6643 2242 6658 2244
rect 6582 2232 6658 2242
rect 6597 2231 6643 2232
rect 6757 2185 6803 2242
rect 6917 2416 6963 2473
rect 6917 2231 6963 2242
rect 7077 2473 7157 2519
rect 7203 2473 7317 2519
rect 7363 2483 7394 2519
rect 7446 2519 7498 2535
rect 7550 2519 7564 2535
rect 10313 2636 10493 2648
rect 10313 2584 10325 2636
rect 10377 2584 10429 2636
rect 10481 2584 10493 2636
rect 10313 2532 10493 2584
rect 7446 2483 7477 2519
rect 7550 2483 7637 2519
rect 7363 2473 7477 2483
rect 7523 2473 7637 2483
rect 7683 2473 7797 2519
rect 7843 2473 7957 2519
rect 8003 2473 8117 2519
rect 8163 2473 8277 2519
rect 8323 2473 8437 2519
rect 8483 2473 8597 2519
rect 8643 2473 8757 2519
rect 8803 2473 8917 2519
rect 8963 2473 9077 2519
rect 9123 2473 9237 2519
rect 9283 2473 9363 2519
rect 7077 2416 7123 2473
rect 7077 2185 7123 2242
rect 6437 2139 7123 2185
rect 7237 2416 7283 2427
rect 7237 2185 7283 2242
rect 7397 2416 7443 2473
rect 7397 2231 7443 2242
rect 7557 2416 7603 2427
rect 7557 2185 7603 2242
rect 7717 2416 7763 2473
rect 7717 2231 7763 2242
rect 7877 2416 7923 2427
rect 7877 2185 7923 2242
rect 8037 2416 8083 2473
rect 8037 2231 8083 2242
rect 8197 2416 8243 2427
rect 8197 2185 8243 2242
rect 8357 2416 8403 2473
rect 8357 2231 8403 2242
rect 8517 2416 8563 2427
rect 8517 2185 8563 2242
rect 8677 2416 8723 2473
rect 8677 2231 8723 2242
rect 8837 2416 8883 2427
rect 8837 2185 8883 2242
rect 8997 2416 9043 2473
rect 8997 2231 9043 2242
rect 9157 2416 9203 2427
rect 9157 2185 9203 2242
rect 9317 2416 9363 2473
rect 10313 2480 10325 2532
rect 10377 2480 10429 2532
rect 10481 2480 10493 2532
rect 10313 2468 10493 2480
rect 9317 2231 9363 2242
rect 9445 2416 9491 2427
rect 9749 2416 9795 2427
rect 10053 2416 10099 2427
rect 9445 2185 9491 2242
rect 9737 2242 9749 2416
rect 9795 2404 9917 2416
rect 9801 2352 9853 2404
rect 9905 2352 9917 2404
rect 9795 2300 9917 2352
rect 9801 2248 9853 2300
rect 9905 2248 9917 2300
rect 9795 2242 9917 2248
rect 9737 2236 9917 2242
rect 9749 2231 9795 2236
rect 10053 2185 10099 2242
rect 10357 2416 10403 2468
rect 10357 2231 10403 2242
rect 10661 2416 10707 2725
rect 10661 2185 10707 2242
rect 7237 2139 10707 2185
rect 6149 1987 6229 2033
rect 6275 1987 6355 2033
rect 10661 2033 10707 2139
rect 10821 2416 10867 2725
rect 10821 2033 10867 2242
rect 6149 1779 6195 1987
rect 6149 1381 6195 1605
rect 6309 1779 6355 1987
rect 9396 2004 9576 2016
rect 9396 1952 9408 2004
rect 9460 1952 9512 2004
rect 9564 1952 9576 2004
rect 6512 1910 6692 1924
rect 6512 1858 6524 1910
rect 6576 1858 6628 1910
rect 6680 1858 6692 1910
rect 9396 1900 9576 1952
rect 9396 1893 9408 1900
rect 6512 1846 6692 1858
rect 6869 1836 7779 1882
rect 8060 1845 8071 1891
rect 8117 1845 8165 1891
rect 8211 1845 8259 1891
rect 8305 1845 8316 1891
rect 8757 1882 9408 1893
rect 6437 1783 6483 1790
rect 6309 1381 6355 1605
rect 6422 1779 6498 1783
rect 6422 1771 6437 1779
rect 6483 1771 6498 1779
rect 6422 1719 6434 1771
rect 6486 1719 6498 1771
rect 6422 1667 6437 1719
rect 6483 1667 6498 1719
rect 6422 1615 6434 1667
rect 6486 1615 6498 1667
rect 6422 1605 6437 1615
rect 6483 1605 6498 1615
rect 6422 1603 6498 1605
rect 6653 1779 6699 1790
rect 6869 1779 6915 1836
rect 6437 1594 6483 1603
rect 6653 1381 6699 1605
rect 6854 1765 6869 1777
rect 7085 1779 7131 1790
rect 6915 1765 6930 1777
rect 6854 1713 6866 1765
rect 6918 1713 6930 1765
rect 6854 1661 6869 1713
rect 6915 1661 6930 1713
rect 6854 1609 6866 1661
rect 6918 1609 6930 1661
rect 6854 1605 6869 1609
rect 6915 1605 6930 1609
rect 6854 1597 6930 1605
rect 6869 1594 6915 1597
rect 7085 1381 7131 1605
rect 7301 1779 7347 1836
rect 7301 1594 7347 1605
rect 7517 1779 7563 1790
rect 7517 1381 7563 1605
rect 7733 1779 7779 1836
rect 7733 1594 7779 1605
rect 7949 1779 7995 1790
rect 7949 1381 7995 1605
rect 8165 1779 8211 1845
rect 8803 1836 8917 1882
rect 8963 1836 9077 1882
rect 9123 1836 9237 1882
rect 9283 1836 9397 1882
rect 9460 1848 9512 1900
rect 9564 1893 9576 1900
rect 10661 1987 10741 2033
rect 10787 1987 10867 2033
rect 9564 1882 9763 1893
rect 9443 1836 9557 1848
rect 9603 1836 9763 1882
rect 8165 1594 8211 1605
rect 8381 1779 8427 1790
rect 8381 1381 8427 1605
rect 8597 1779 8643 1790
rect 8597 1548 8643 1605
rect 8757 1779 8803 1836
rect 8757 1594 8803 1605
rect 8917 1779 8963 1790
rect 8917 1548 8963 1605
rect 9077 1779 9123 1836
rect 9077 1594 9123 1605
rect 9237 1779 9283 1790
rect 9237 1548 9283 1605
rect 9397 1779 9443 1836
rect 9397 1594 9443 1605
rect 9557 1779 9603 1790
rect 9557 1548 9603 1605
rect 9717 1779 9763 1836
rect 9717 1594 9763 1605
rect 9861 1779 9907 1790
rect 8597 1502 9603 1548
rect 9861 1381 9907 1605
rect 10021 1779 10067 1790
rect 10021 1381 10067 1605
rect 10181 1779 10227 1790
rect 10181 1381 10227 1605
rect 10341 1779 10387 1790
rect 10341 1381 10387 1605
rect 10501 1779 10547 1790
rect 10501 1381 10547 1605
rect 10661 1779 10707 1987
rect 10661 1381 10707 1605
rect 10821 1779 10867 1987
rect 10821 1381 10867 1605
rect 11013 2688 11070 2725
rect 11116 2731 12014 2734
rect 12060 2731 12246 2777
rect 11116 2688 12246 2731
rect 11013 2683 12246 2688
rect 11013 2640 12014 2683
rect 11013 2594 11070 2640
rect 11116 2637 12014 2640
rect 12060 2637 12246 2683
rect 11116 2594 12246 2637
rect 11013 2589 12246 2594
rect 11013 2565 12014 2589
rect 11013 2546 11173 2565
rect 11013 2500 11070 2546
rect 11116 2500 11173 2546
rect 11013 2452 11173 2500
rect 11013 2406 11070 2452
rect 11116 2406 11173 2452
rect 11013 2358 11173 2406
rect 11013 2312 11070 2358
rect 11116 2312 11173 2358
rect 11013 2264 11173 2312
rect 11013 2218 11070 2264
rect 11116 2218 11173 2264
rect 11013 2170 11173 2218
rect 11013 2124 11070 2170
rect 11116 2124 11173 2170
rect 11013 2076 11173 2124
rect 11013 2030 11070 2076
rect 11116 2030 11173 2076
rect 11013 1982 11173 2030
rect 11926 2543 12014 2565
rect 12060 2543 12246 2589
rect 11926 2495 12246 2543
rect 11926 2449 12014 2495
rect 12060 2449 12246 2495
rect 11926 2401 12246 2449
rect 11926 2355 12014 2401
rect 12060 2355 12246 2401
rect 11926 2307 12246 2355
rect 11926 2261 12014 2307
rect 12060 2261 12246 2307
rect 11926 2213 12246 2261
rect 11926 2167 12014 2213
rect 12060 2167 12246 2213
rect 11926 2119 12246 2167
rect 11926 2073 12014 2119
rect 12060 2073 12246 2119
rect 11926 2025 12246 2073
rect 11013 1936 11070 1982
rect 11116 1936 11173 1982
rect 11013 1888 11173 1936
rect 11013 1842 11070 1888
rect 11116 1842 11173 1888
rect 11013 1794 11173 1842
rect 11305 2006 11485 2016
rect 11305 2004 11780 2006
rect 11305 1952 11317 2004
rect 11369 1952 11421 2004
rect 11473 1952 11780 2004
rect 11305 1900 11780 1952
rect 11305 1848 11317 1900
rect 11369 1848 11421 1900
rect 11473 1848 11780 1900
rect 11305 1846 11780 1848
rect 11926 1979 12014 2025
rect 12060 1979 12246 2025
rect 11926 1931 12246 1979
rect 11926 1885 12014 1931
rect 12060 1885 12246 1931
rect 11305 1836 11485 1846
rect 11926 1837 12246 1885
rect 11013 1748 11070 1794
rect 11116 1748 11173 1794
rect 11013 1700 11173 1748
rect 11013 1654 11070 1700
rect 11116 1654 11173 1700
rect 11013 1606 11173 1654
rect 11013 1560 11070 1606
rect 11116 1560 11173 1606
rect 11013 1541 11173 1560
rect 11926 1791 12014 1837
rect 12060 1791 12246 1837
rect 11926 1743 12246 1791
rect 11926 1697 12014 1743
rect 12060 1697 12246 1743
rect 11926 1649 12246 1697
rect 11926 1603 12014 1649
rect 12060 1603 12246 1649
rect 11926 1555 12246 1603
rect 11926 1541 12014 1555
rect 11013 1512 12014 1541
rect 11013 1466 11070 1512
rect 11116 1509 12014 1512
rect 12060 1541 12246 1555
rect 12683 3768 12729 4249
rect 12683 3232 12729 3394
rect 12683 2697 12729 2858
rect 12987 3768 13033 4249
rect 12987 3232 13033 3394
rect 12987 2697 13033 2858
rect 13115 3768 13161 4249
rect 13209 4001 13371 4249
rect 13209 3955 13220 4001
rect 13266 3955 13314 4001
rect 13360 3955 13371 4001
rect 13209 3907 13371 3955
rect 13209 3861 13220 3907
rect 13266 3861 13314 3907
rect 13360 3861 13371 3907
rect 13209 3850 13371 3861
rect 13115 3232 13161 3394
rect 13115 2847 13161 2858
rect 13419 3768 13465 4249
rect 13419 3232 13465 3394
rect 12683 2651 12788 2697
rect 12834 2651 12882 2697
rect 12928 2651 13033 2697
rect 12683 2603 13033 2651
rect 12683 2557 12788 2603
rect 12834 2557 12882 2603
rect 12928 2557 13033 2603
rect 12683 2396 12729 2557
rect 12683 1541 12729 2022
rect 12987 2396 13033 2557
rect 13115 2396 13161 2407
rect 13100 2294 13115 2306
rect 13419 2396 13465 2858
rect 13723 3768 13769 3779
rect 13723 3232 13769 3394
rect 13723 2708 13769 2858
rect 14027 3768 14073 4249
rect 14027 3232 14073 3394
rect 13618 2662 13629 2708
rect 13675 2662 13723 2708
rect 13769 2662 13817 2708
rect 13863 2662 13874 2708
rect 13161 2294 13176 2306
rect 13100 2242 13112 2294
rect 13164 2242 13176 2294
rect 13100 2190 13115 2242
rect 13161 2190 13176 2242
rect 13100 2138 13112 2190
rect 13164 2138 13176 2190
rect 13100 2086 13115 2138
rect 13161 2086 13176 2138
rect 13100 2034 13112 2086
rect 13164 2034 13176 2086
rect 13100 2022 13115 2034
rect 13161 2022 13176 2034
rect 12987 1541 13033 2022
rect 13115 2011 13161 2022
rect 13419 2011 13465 2022
rect 13723 2396 13769 2407
rect 13723 1832 13769 2022
rect 14027 2396 14073 2858
rect 14331 3768 14377 3779
rect 14331 3232 14377 3394
rect 14331 2708 14377 2858
rect 14635 3768 14681 4249
rect 14635 3232 14681 3394
rect 14226 2662 14237 2708
rect 14283 2662 14331 2708
rect 14377 2662 14425 2708
rect 14471 2662 14482 2708
rect 13200 1815 13380 1827
rect 13200 1763 13212 1815
rect 13264 1763 13316 1815
rect 13368 1763 13380 1815
rect 13618 1786 13629 1832
rect 13675 1786 13723 1832
rect 13769 1786 13817 1832
rect 13863 1786 13874 1832
rect 13200 1711 13380 1763
rect 13200 1659 13212 1711
rect 13264 1659 13316 1711
rect 13368 1659 13380 1711
rect 13200 1647 13380 1659
rect 14027 1541 14073 2022
rect 14331 2396 14377 2407
rect 14331 1847 14377 2022
rect 14635 2396 14681 2858
rect 14939 3768 14985 3779
rect 15067 3768 15113 3779
rect 15052 3562 15067 3574
rect 15371 3768 15417 4249
rect 15113 3562 15128 3574
rect 15052 3510 15064 3562
rect 15116 3510 15128 3562
rect 15052 3458 15067 3510
rect 15113 3458 15128 3510
rect 15052 3406 15064 3458
rect 15116 3406 15128 3458
rect 15052 3394 15067 3406
rect 15113 3394 15128 3406
rect 15675 3768 15721 3779
rect 15660 3562 15675 3574
rect 15979 3768 16025 4249
rect 15721 3562 15736 3574
rect 15660 3510 15672 3562
rect 15724 3510 15736 3562
rect 15660 3458 15675 3510
rect 15721 3458 15736 3510
rect 15660 3406 15672 3458
rect 15724 3406 15736 3458
rect 15660 3394 15675 3406
rect 15721 3394 15736 3406
rect 16283 3768 16329 3779
rect 16268 3562 16283 3574
rect 16587 3768 16633 4249
rect 16329 3562 16344 3574
rect 16268 3510 16280 3562
rect 16332 3510 16344 3562
rect 16268 3458 16283 3510
rect 16329 3458 16344 3510
rect 16268 3406 16280 3458
rect 16332 3406 16344 3458
rect 16268 3394 16283 3406
rect 16329 3394 16344 3406
rect 14939 3232 14985 3394
rect 14939 2708 14985 2858
rect 15067 3232 15113 3394
rect 15067 2847 15113 2858
rect 15371 3232 15417 3394
rect 15371 2847 15417 2858
rect 15675 3232 15721 3394
rect 15675 2847 15721 2858
rect 15979 3232 16025 3394
rect 15979 2847 16025 2858
rect 16283 3232 16329 3394
rect 16283 2847 16329 2858
rect 16587 3232 16633 3394
rect 16171 2763 16455 2785
rect 16171 2711 16183 2763
rect 16235 2711 16287 2763
rect 16339 2711 16391 2763
rect 16443 2711 16455 2763
rect 14834 2662 14845 2708
rect 14891 2662 14939 2708
rect 14985 2662 15033 2708
rect 15079 2662 15090 2708
rect 16171 2659 16455 2711
rect 16171 2607 16183 2659
rect 16235 2607 16287 2659
rect 16339 2607 16391 2659
rect 16443 2607 16455 2659
rect 16171 2585 16455 2607
rect 16587 2697 16633 2858
rect 16891 3768 16937 4249
rect 16891 3232 16937 3394
rect 16891 2697 16937 2858
rect 16587 2651 16692 2697
rect 16738 2651 16786 2697
rect 16832 2651 16937 2697
rect 16587 2603 16937 2651
rect 16587 2557 16692 2603
rect 16738 2557 16786 2603
rect 16832 2557 16937 2603
rect 15067 2453 16329 2499
rect 14212 1835 14496 1847
rect 14212 1783 14224 1835
rect 14276 1783 14328 1835
rect 14380 1783 14432 1835
rect 14484 1783 14496 1835
rect 14212 1771 14496 1783
rect 14635 1541 14681 2022
rect 14939 2396 14985 2407
rect 14939 1832 14985 2022
rect 15067 2396 15113 2453
rect 15067 2011 15113 2022
rect 15371 2396 15417 2407
rect 15675 2396 15721 2453
rect 15660 2294 15675 2306
rect 15979 2396 16025 2407
rect 15721 2294 15736 2306
rect 15660 2242 15672 2294
rect 15724 2242 15736 2294
rect 15660 2190 15675 2242
rect 15721 2190 15736 2242
rect 15660 2138 15672 2190
rect 15724 2138 15736 2190
rect 15660 2086 15675 2138
rect 15721 2086 15736 2138
rect 15660 2034 15672 2086
rect 15724 2034 15736 2086
rect 15660 2022 15675 2034
rect 15721 2022 15736 2034
rect 14834 1786 14845 1832
rect 14891 1786 14939 1832
rect 14985 1786 15033 1832
rect 15079 1786 15090 1832
rect 15371 1541 15417 2022
rect 15675 2011 15721 2022
rect 15979 1541 16025 2022
rect 16283 2396 16329 2453
rect 16283 2011 16329 2022
rect 16587 2396 16633 2557
rect 16587 1541 16633 2022
rect 16891 2396 16937 2557
rect 16891 1541 16937 2022
rect 17374 4235 17560 4249
rect 17606 4235 17694 4281
rect 17374 4187 17694 4235
rect 17374 4141 17560 4187
rect 17606 4141 17694 4187
rect 17374 4093 17694 4141
rect 17374 4047 17560 4093
rect 17606 4047 17694 4093
rect 17374 3999 17694 4047
rect 17374 3953 17560 3999
rect 17606 3953 17694 3999
rect 17374 3905 17694 3953
rect 17374 3859 17560 3905
rect 17606 3859 17694 3905
rect 17374 3811 17694 3859
rect 17374 3765 17560 3811
rect 17606 3765 17694 3811
rect 17374 3717 17694 3765
rect 17374 3671 17560 3717
rect 17606 3671 17694 3717
rect 17374 3623 17694 3671
rect 17374 3577 17560 3623
rect 17606 3577 17694 3623
rect 17374 3529 17694 3577
rect 17374 3483 17560 3529
rect 17606 3483 17694 3529
rect 17374 3435 17694 3483
rect 17374 3389 17560 3435
rect 17606 3389 17694 3435
rect 17374 3341 17694 3389
rect 17374 3295 17560 3341
rect 17606 3295 17694 3341
rect 17374 3247 17694 3295
rect 17374 3201 17560 3247
rect 17606 3201 17694 3247
rect 17374 3153 17694 3201
rect 17374 3107 17560 3153
rect 17606 3107 17694 3153
rect 17374 3059 17694 3107
rect 17374 3013 17560 3059
rect 17606 3013 17694 3059
rect 17374 2965 17694 3013
rect 17374 2919 17560 2965
rect 17606 2919 17694 2965
rect 17374 2871 17694 2919
rect 17374 2825 17560 2871
rect 17606 2825 17694 2871
rect 17374 2777 17694 2825
rect 17374 2731 17560 2777
rect 17606 2731 17694 2777
rect 17374 2683 17694 2731
rect 17374 2637 17560 2683
rect 17606 2637 17694 2683
rect 17374 2589 17694 2637
rect 17374 2543 17560 2589
rect 17606 2543 17694 2589
rect 17374 2495 17694 2543
rect 17374 2449 17560 2495
rect 17606 2449 17694 2495
rect 17374 2401 17694 2449
rect 17374 2355 17560 2401
rect 17606 2355 17694 2401
rect 17374 2307 17694 2355
rect 17374 2261 17560 2307
rect 17606 2261 17694 2307
rect 17374 2213 17694 2261
rect 17374 2167 17560 2213
rect 17606 2167 17694 2213
rect 17374 2119 17694 2167
rect 17374 2073 17560 2119
rect 17606 2073 17694 2119
rect 17374 2025 17694 2073
rect 17374 1979 17560 2025
rect 17606 1979 17694 2025
rect 17374 1931 17694 1979
rect 17374 1885 17560 1931
rect 17606 1885 17694 1931
rect 17374 1837 17694 1885
rect 17374 1791 17560 1837
rect 17606 1791 17694 1837
rect 17374 1743 17694 1791
rect 17374 1697 17560 1743
rect 17606 1697 17694 1743
rect 17374 1649 17694 1697
rect 17374 1603 17560 1649
rect 17606 1603 17694 1649
rect 17374 1555 17694 1603
rect 17374 1541 17560 1555
rect 12060 1509 17560 1541
rect 17606 1509 17694 1555
rect 11116 1466 17694 1509
rect 11013 1461 17694 1466
rect 11013 1418 12014 1461
rect 11013 1381 11070 1418
rect 5946 1372 11070 1381
rect 11116 1415 12014 1418
rect 12060 1415 17560 1461
rect 17606 1415 17694 1461
rect 11116 1372 17694 1415
rect 5843 1367 17694 1372
rect 5843 1324 12014 1367
rect 5843 1278 5900 1324
rect 5946 1278 5994 1324
rect 6040 1278 6088 1324
rect 6134 1278 6182 1324
rect 6228 1278 6276 1324
rect 6322 1278 6370 1324
rect 6416 1278 6464 1324
rect 6510 1278 6558 1324
rect 6604 1278 6652 1324
rect 6698 1278 6746 1324
rect 6792 1278 6840 1324
rect 6886 1278 6934 1324
rect 6980 1278 7028 1324
rect 7074 1278 7122 1324
rect 7168 1278 7216 1324
rect 7262 1278 7310 1324
rect 7356 1278 7404 1324
rect 7450 1278 7498 1324
rect 7544 1278 7592 1324
rect 7638 1278 7686 1324
rect 7732 1278 7780 1324
rect 7826 1278 7874 1324
rect 7920 1278 7968 1324
rect 8014 1278 8062 1324
rect 8108 1278 8156 1324
rect 8202 1278 8250 1324
rect 8296 1278 8344 1324
rect 8390 1278 8438 1324
rect 8484 1278 8532 1324
rect 8578 1278 8626 1324
rect 8672 1278 8720 1324
rect 8766 1278 8814 1324
rect 8860 1278 8908 1324
rect 8954 1278 9002 1324
rect 9048 1278 9096 1324
rect 9142 1278 9190 1324
rect 9236 1278 9284 1324
rect 9330 1278 9378 1324
rect 9424 1278 9472 1324
rect 9518 1278 9566 1324
rect 9612 1278 9660 1324
rect 9706 1278 9754 1324
rect 9800 1278 9848 1324
rect 9894 1278 9942 1324
rect 9988 1278 10036 1324
rect 10082 1278 10130 1324
rect 10176 1278 10224 1324
rect 10270 1278 10318 1324
rect 10364 1278 10412 1324
rect 10458 1278 10506 1324
rect 10552 1278 10600 1324
rect 10646 1278 10694 1324
rect 10740 1278 10788 1324
rect 10834 1278 10882 1324
rect 10928 1278 10976 1324
rect 11022 1278 11070 1324
rect 11116 1321 12014 1324
rect 12060 1321 12108 1367
rect 12154 1321 12202 1367
rect 12248 1321 12296 1367
rect 12342 1321 12390 1367
rect 12436 1321 12484 1367
rect 12530 1321 12578 1367
rect 12624 1321 12672 1367
rect 12718 1321 12766 1367
rect 12812 1321 12860 1367
rect 12906 1321 12954 1367
rect 13000 1321 13048 1367
rect 13094 1321 13142 1367
rect 13188 1321 13236 1367
rect 13282 1321 13330 1367
rect 13376 1321 13424 1367
rect 13470 1321 13518 1367
rect 13564 1321 13612 1367
rect 13658 1321 13706 1367
rect 13752 1321 13800 1367
rect 13846 1321 13894 1367
rect 13940 1321 13988 1367
rect 14034 1321 14082 1367
rect 14128 1321 14176 1367
rect 14222 1321 14270 1367
rect 14316 1321 14364 1367
rect 14410 1321 14458 1367
rect 14504 1321 14552 1367
rect 14598 1321 14646 1367
rect 14692 1321 14740 1367
rect 14786 1321 14834 1367
rect 14880 1321 14928 1367
rect 14974 1321 15022 1367
rect 15068 1321 15116 1367
rect 15162 1321 15210 1367
rect 15256 1321 15304 1367
rect 15350 1321 15398 1367
rect 15444 1321 15492 1367
rect 15538 1321 15586 1367
rect 15632 1321 15680 1367
rect 15726 1321 15774 1367
rect 15820 1321 15868 1367
rect 15914 1321 15962 1367
rect 16008 1321 16056 1367
rect 16102 1321 16150 1367
rect 16196 1321 16244 1367
rect 16290 1321 16338 1367
rect 16384 1321 16432 1367
rect 16478 1321 16526 1367
rect 16572 1321 16620 1367
rect 16666 1321 16714 1367
rect 16760 1321 16808 1367
rect 16854 1321 16902 1367
rect 16948 1321 16996 1367
rect 17042 1321 17090 1367
rect 17136 1321 17184 1367
rect 17230 1321 17278 1367
rect 17324 1321 17372 1367
rect 17418 1321 17466 1367
rect 17512 1321 17560 1367
rect 17606 1321 17694 1367
rect 11116 1278 17694 1321
rect 5843 1221 17694 1278
rect 18076 4527 18206 4573
rect 18252 4527 18396 4573
rect 18076 4479 18396 4527
rect 18076 4433 18206 4479
rect 18252 4433 18396 4479
rect 18076 4385 18396 4433
rect 18076 4339 18206 4385
rect 18252 4339 18396 4385
rect 18076 4291 18396 4339
rect 18076 4245 18206 4291
rect 18252 4245 18396 4291
rect 18076 4197 18396 4245
rect 18076 4151 18206 4197
rect 18252 4151 18396 4197
rect 18076 4103 18396 4151
rect 18076 4057 18206 4103
rect 18252 4057 18396 4103
rect 18076 4009 18396 4057
rect 18076 3963 18206 4009
rect 18252 3963 18396 4009
rect 18076 3915 18396 3963
rect 18076 3869 18206 3915
rect 18252 3869 18396 3915
rect 18076 3821 18396 3869
rect 18076 3775 18206 3821
rect 18252 3775 18396 3821
rect 18076 3727 18396 3775
rect 18076 3681 18206 3727
rect 18252 3681 18396 3727
rect 18076 3633 18396 3681
rect 18076 3587 18206 3633
rect 18252 3587 18396 3633
rect 18076 3539 18396 3587
rect 18076 3493 18206 3539
rect 18252 3493 18396 3539
rect 18076 3445 18396 3493
rect 18076 3399 18206 3445
rect 18252 3399 18396 3445
rect 18076 3351 18396 3399
rect 18076 3305 18206 3351
rect 18252 3305 18396 3351
rect 18076 3257 18396 3305
rect 18076 3211 18206 3257
rect 18252 3211 18396 3257
rect 18076 3163 18396 3211
rect 18076 3117 18206 3163
rect 18252 3117 18396 3163
rect 18076 3069 18396 3117
rect 18076 3023 18206 3069
rect 18252 3023 18396 3069
rect 18076 2975 18396 3023
rect 18076 2929 18206 2975
rect 18252 2929 18396 2975
rect 18076 2881 18396 2929
rect 18076 2835 18206 2881
rect 18252 2835 18396 2881
rect 18076 2787 18396 2835
rect 18076 2741 18206 2787
rect 18252 2741 18396 2787
rect 18076 2693 18396 2741
rect 18076 2647 18206 2693
rect 18252 2647 18396 2693
rect 18076 2599 18396 2647
rect 18076 2553 18206 2599
rect 18252 2553 18396 2599
rect 18076 2505 18396 2553
rect 18076 2459 18206 2505
rect 18252 2459 18396 2505
rect 18076 2411 18396 2459
rect 18076 2365 18206 2411
rect 18252 2365 18396 2411
rect 18076 2317 18396 2365
rect 18076 2271 18206 2317
rect 18252 2271 18396 2317
rect 18076 2223 18396 2271
rect 18076 2177 18206 2223
rect 18252 2177 18396 2223
rect 18076 2129 18396 2177
rect 18076 2083 18206 2129
rect 18252 2083 18396 2129
rect 18076 2035 18396 2083
rect 18076 1989 18206 2035
rect 18252 1989 18396 2035
rect 18076 1941 18396 1989
rect 18076 1895 18206 1941
rect 18252 1895 18396 1941
rect 18076 1847 18396 1895
rect 18076 1801 18206 1847
rect 18252 1801 18396 1847
rect 18076 1753 18396 1801
rect 18076 1707 18206 1753
rect 18252 1707 18396 1753
rect 18076 1659 18396 1707
rect 18076 1613 18206 1659
rect 18252 1613 18396 1659
rect 18076 1565 18396 1613
rect 18076 1519 18206 1565
rect 18252 1519 18396 1565
rect 18076 1471 18396 1519
rect 18076 1425 18206 1471
rect 18252 1425 18396 1471
rect 18076 1377 18396 1425
rect 18076 1331 18206 1377
rect 18252 1331 18396 1377
rect 18076 1283 18396 1331
rect 18076 1237 18206 1283
rect 18252 1259 18396 1283
rect 18795 4766 18841 5491
rect 18795 4134 18841 4192
rect 18955 4766 19001 5491
rect 18955 4134 19001 4192
rect 18795 4088 18875 4134
rect 18921 4088 19001 4134
rect 18795 4030 18841 4088
rect 18795 3294 18841 3456
rect 18795 2662 18841 2720
rect 18955 4030 19001 4088
rect 18955 3294 19001 3456
rect 18955 2662 19001 2720
rect 18795 2616 18875 2662
rect 18921 2616 19001 2662
rect 18795 2558 18841 2616
rect 18795 1259 18841 1984
rect 18955 2558 19001 2616
rect 19115 4766 19161 4777
rect 19115 4030 19161 4192
rect 19115 3294 19161 3456
rect 19115 2558 19161 2720
rect 19100 2256 19115 2268
rect 19275 4766 19321 5491
rect 19275 4030 19321 4192
rect 19275 3294 19321 3456
rect 19275 2558 19321 2720
rect 19161 2256 19176 2268
rect 19100 2204 19112 2256
rect 19164 2204 19176 2256
rect 19100 2152 19115 2204
rect 19161 2152 19176 2204
rect 19100 2100 19112 2152
rect 19164 2100 19176 2152
rect 19100 2048 19115 2100
rect 19161 2048 19176 2100
rect 19100 1996 19112 2048
rect 19164 1996 19176 2048
rect 19100 1984 19115 1996
rect 19161 1984 19176 1996
rect 19435 4766 19481 4777
rect 19435 4030 19481 4192
rect 19435 3294 19481 3456
rect 19435 2558 19481 2720
rect 19420 2256 19435 2268
rect 19595 4766 19641 5491
rect 19595 4030 19641 4192
rect 19595 3294 19641 3456
rect 19595 2558 19641 2720
rect 19481 2256 19496 2268
rect 19420 2204 19432 2256
rect 19484 2204 19496 2256
rect 19420 2152 19435 2204
rect 19481 2152 19496 2204
rect 19420 2100 19432 2152
rect 19484 2100 19496 2152
rect 19420 2048 19435 2100
rect 19481 2048 19496 2100
rect 19420 1996 19432 2048
rect 19484 1996 19496 2048
rect 19420 1984 19435 1996
rect 19481 1984 19496 1996
rect 19755 4766 19801 4777
rect 19755 4030 19801 4192
rect 19755 3294 19801 3456
rect 19755 2558 19801 2720
rect 19740 2256 19755 2268
rect 19915 4766 19961 5491
rect 19915 4030 19961 4192
rect 19915 3294 19961 3456
rect 19915 2558 19961 2720
rect 19801 2256 19816 2268
rect 19740 2204 19752 2256
rect 19804 2204 19816 2256
rect 19740 2152 19755 2204
rect 19801 2152 19816 2204
rect 19740 2100 19752 2152
rect 19804 2100 19816 2152
rect 19740 2048 19755 2100
rect 19801 2048 19816 2100
rect 19740 1996 19752 2048
rect 19804 1996 19816 2048
rect 19740 1984 19755 1996
rect 19801 1984 19816 1996
rect 20075 4766 20121 4777
rect 20075 4030 20121 4192
rect 20075 3294 20121 3456
rect 20075 2558 20121 2720
rect 20060 2256 20075 2268
rect 20235 4766 20281 5491
rect 20235 4030 20281 4192
rect 20235 3294 20281 3456
rect 20235 2558 20281 2720
rect 20121 2256 20136 2268
rect 20060 2204 20072 2256
rect 20124 2204 20136 2256
rect 20060 2152 20075 2204
rect 20121 2152 20136 2204
rect 20060 2100 20072 2152
rect 20124 2100 20136 2152
rect 20060 2048 20075 2100
rect 20121 2048 20136 2100
rect 20060 1996 20072 2048
rect 20124 1996 20136 2048
rect 20060 1984 20075 1996
rect 20121 1984 20136 1996
rect 20395 4766 20441 4777
rect 20395 4030 20441 4192
rect 20395 3294 20441 3456
rect 20395 2558 20441 2720
rect 20380 2256 20395 2268
rect 20555 4766 20601 5491
rect 20647 4918 20827 4930
rect 20647 4866 20659 4918
rect 20711 4866 20763 4918
rect 20815 4866 20827 4918
rect 20647 4854 20827 4866
rect 20555 4030 20601 4192
rect 20555 3294 20601 3456
rect 20555 2558 20601 2720
rect 20441 2256 20456 2268
rect 20380 2204 20392 2256
rect 20444 2204 20456 2256
rect 20380 2152 20395 2204
rect 20441 2152 20456 2204
rect 20380 2100 20392 2152
rect 20444 2100 20456 2152
rect 20380 2048 20395 2100
rect 20441 2048 20456 2100
rect 20380 1996 20392 2048
rect 20444 1996 20456 2048
rect 20380 1984 20395 1996
rect 20441 1984 20456 1996
rect 20715 4766 20761 4777
rect 20715 4030 20761 4192
rect 20715 3294 20761 3456
rect 20715 2558 20761 2720
rect 20700 2256 20715 2268
rect 20875 4766 20921 5491
rect 20875 4030 20921 4192
rect 20875 3294 20921 3456
rect 20875 2558 20921 2720
rect 20761 2256 20776 2268
rect 20700 2204 20712 2256
rect 20764 2204 20776 2256
rect 20700 2152 20715 2204
rect 20761 2152 20776 2204
rect 20700 2100 20712 2152
rect 20764 2100 20776 2152
rect 20700 2048 20715 2100
rect 20761 2048 20776 2100
rect 20700 1996 20712 2048
rect 20764 1996 20776 2048
rect 20700 1984 20715 1996
rect 20761 1984 20776 1996
rect 21035 4766 21081 4777
rect 21035 4030 21081 4192
rect 21035 3294 21081 3456
rect 21035 2558 21081 2720
rect 21020 2256 21035 2268
rect 21195 4766 21241 5491
rect 21195 4030 21241 4192
rect 21195 3294 21241 3456
rect 21195 2558 21241 2720
rect 21081 2256 21096 2268
rect 21020 2204 21032 2256
rect 21084 2204 21096 2256
rect 21020 2152 21035 2204
rect 21081 2152 21096 2204
rect 21020 2100 21032 2152
rect 21084 2100 21096 2152
rect 21020 2048 21035 2100
rect 21081 2048 21096 2100
rect 21020 1996 21032 2048
rect 21084 1996 21096 2048
rect 21020 1984 21035 1996
rect 21081 1984 21096 1996
rect 18955 1259 19001 1984
rect 19115 1897 19161 1984
rect 19275 1973 19321 1984
rect 19435 1897 19481 1984
rect 19595 1973 19641 1984
rect 19755 1897 19801 1984
rect 19915 1973 19961 1984
rect 20075 1897 20121 1984
rect 20235 1973 20281 1984
rect 20395 1897 20441 1984
rect 20555 1973 20601 1984
rect 20715 1897 20761 1984
rect 20875 1973 20921 1984
rect 21035 1897 21081 1984
rect 19115 1851 21081 1897
rect 21195 1259 21241 1984
rect 21355 4915 21401 4926
rect 21355 4766 21401 4869
rect 21355 4030 21401 4192
rect 21355 3294 21401 3456
rect 21355 2558 21401 2720
rect 21355 1973 21401 1984
rect 21515 4766 21561 5491
rect 21675 4766 21721 4777
rect 21660 4464 21675 4476
rect 21835 4766 21881 5491
rect 21721 4464 21736 4476
rect 21660 4412 21672 4464
rect 21724 4412 21736 4464
rect 21660 4360 21675 4412
rect 21721 4360 21736 4412
rect 21660 4308 21672 4360
rect 21724 4308 21736 4360
rect 21660 4256 21675 4308
rect 21721 4256 21736 4308
rect 21660 4204 21672 4256
rect 21724 4204 21736 4256
rect 21660 4192 21675 4204
rect 21721 4192 21736 4204
rect 21515 4030 21561 4192
rect 21515 3294 21561 3456
rect 21515 2558 21561 2720
rect 21515 1259 21561 1984
rect 21675 4030 21721 4192
rect 21675 3294 21721 3456
rect 21675 2558 21721 2720
rect 21675 1973 21721 1984
rect 21835 4030 21881 4192
rect 21835 3294 21881 3456
rect 21963 4766 22009 5491
rect 21963 4134 22009 4192
rect 22123 4766 22169 5491
rect 22123 4134 22169 4192
rect 21963 4088 22043 4134
rect 22089 4088 22169 4134
rect 21963 4030 22009 4088
rect 21963 3445 22009 3456
rect 22123 4030 22169 4088
rect 21835 2558 21881 2720
rect 21835 1973 21881 1984
rect 21963 3194 22009 3205
rect 21963 2458 22009 2720
rect 21631 1904 21915 1916
rect 21631 1852 21643 1904
rect 21695 1852 21747 1904
rect 21799 1852 21851 1904
rect 21903 1852 21915 1904
rect 21631 1842 21915 1852
rect 21963 1901 22009 1984
rect 21963 1844 22009 1855
rect 22123 3194 22169 3456
rect 22123 2458 22169 2720
rect 22123 1259 22169 1984
rect 22251 4766 22297 5491
rect 22251 4134 22297 4192
rect 22411 4766 22457 5491
rect 22411 4134 22457 4192
rect 22251 4088 22331 4134
rect 22377 4088 22457 4134
rect 22251 4030 22297 4088
rect 22251 3294 22297 3456
rect 22251 2662 22297 2720
rect 22411 4030 22457 4088
rect 22411 3294 22457 3456
rect 22411 2662 22457 2720
rect 22251 2616 22331 2662
rect 22377 2616 22457 2662
rect 22251 2558 22297 2616
rect 22251 1259 22297 1984
rect 22411 2558 22457 2616
rect 22411 1259 22457 1984
rect 22856 5467 23000 5491
rect 23046 5491 28734 5513
rect 23046 5467 23176 5491
rect 22856 5419 23176 5467
rect 22856 5373 23000 5419
rect 23046 5373 23176 5419
rect 22856 5325 23176 5373
rect 22856 5279 23000 5325
rect 23046 5279 23176 5325
rect 22856 5231 23176 5279
rect 22856 5185 23000 5231
rect 23046 5185 23176 5231
rect 22856 5137 23176 5185
rect 22856 5091 23000 5137
rect 23046 5091 23176 5137
rect 22856 5043 23176 5091
rect 22856 4997 23000 5043
rect 23046 4997 23176 5043
rect 22856 4949 23176 4997
rect 22856 4903 23000 4949
rect 23046 4903 23176 4949
rect 22856 4855 23176 4903
rect 22856 4809 23000 4855
rect 23046 4809 23176 4855
rect 22856 4761 23176 4809
rect 22856 4715 23000 4761
rect 23046 4715 23176 4761
rect 22856 4667 23176 4715
rect 22856 4621 23000 4667
rect 23046 4621 23176 4667
rect 22856 4573 23176 4621
rect 22856 4527 23000 4573
rect 23046 4527 23176 4573
rect 22856 4479 23176 4527
rect 22856 4433 23000 4479
rect 23046 4433 23176 4479
rect 22856 4385 23176 4433
rect 22856 4339 23000 4385
rect 23046 4339 23176 4385
rect 22856 4291 23176 4339
rect 22856 4245 23000 4291
rect 23046 4245 23176 4291
rect 22856 4197 23176 4245
rect 22856 4151 23000 4197
rect 23046 4151 23176 4197
rect 22856 4103 23176 4151
rect 22856 4057 23000 4103
rect 23046 4057 23176 4103
rect 22856 4009 23176 4057
rect 22856 3963 23000 4009
rect 23046 3963 23176 4009
rect 22856 3915 23176 3963
rect 22856 3869 23000 3915
rect 23046 3869 23176 3915
rect 22856 3821 23176 3869
rect 22856 3775 23000 3821
rect 23046 3775 23176 3821
rect 22856 3727 23176 3775
rect 22856 3681 23000 3727
rect 23046 3681 23176 3727
rect 22856 3633 23176 3681
rect 22856 3587 23000 3633
rect 23046 3587 23176 3633
rect 22856 3539 23176 3587
rect 22856 3493 23000 3539
rect 23046 3493 23176 3539
rect 22856 3445 23176 3493
rect 22856 3399 23000 3445
rect 23046 3399 23176 3445
rect 22856 3351 23176 3399
rect 22856 3305 23000 3351
rect 23046 3305 23176 3351
rect 22856 3257 23176 3305
rect 22856 3211 23000 3257
rect 23046 3211 23176 3257
rect 22856 3163 23176 3211
rect 22856 3117 23000 3163
rect 23046 3117 23176 3163
rect 22856 3069 23176 3117
rect 22856 3023 23000 3069
rect 23046 3023 23176 3069
rect 22856 2975 23176 3023
rect 22856 2929 23000 2975
rect 23046 2929 23176 2975
rect 22856 2881 23176 2929
rect 22856 2835 23000 2881
rect 23046 2835 23176 2881
rect 22856 2787 23176 2835
rect 22856 2741 23000 2787
rect 23046 2741 23176 2787
rect 22856 2693 23176 2741
rect 22856 2647 23000 2693
rect 23046 2647 23176 2693
rect 22856 2599 23176 2647
rect 22856 2553 23000 2599
rect 23046 2553 23176 2599
rect 22856 2505 23176 2553
rect 22856 2459 23000 2505
rect 23046 2459 23176 2505
rect 22856 2411 23176 2459
rect 22856 2365 23000 2411
rect 23046 2365 23176 2411
rect 22856 2317 23176 2365
rect 22856 2271 23000 2317
rect 23046 2271 23176 2317
rect 22856 2223 23176 2271
rect 22856 2177 23000 2223
rect 23046 2177 23176 2223
rect 22856 2129 23176 2177
rect 22856 2083 23000 2129
rect 23046 2083 23176 2129
rect 22856 2035 23176 2083
rect 22856 1989 23000 2035
rect 23046 1989 23176 2035
rect 22856 1941 23176 1989
rect 22856 1895 23000 1941
rect 23046 1895 23176 1941
rect 22856 1847 23176 1895
rect 22856 1801 23000 1847
rect 23046 1801 23176 1847
rect 22856 1753 23176 1801
rect 22856 1707 23000 1753
rect 23046 1707 23176 1753
rect 22856 1659 23176 1707
rect 22856 1613 23000 1659
rect 23046 1613 23176 1659
rect 22856 1565 23176 1613
rect 22856 1519 23000 1565
rect 23046 1519 23176 1565
rect 22856 1471 23176 1519
rect 22856 1425 23000 1471
rect 23046 1425 23176 1471
rect 22856 1377 23176 1425
rect 22856 1331 23000 1377
rect 23046 1331 23176 1377
rect 22856 1283 23176 1331
rect 22856 1259 23000 1283
rect 18252 1237 23000 1259
rect 23046 1259 23176 1283
rect 23662 4906 23858 5491
rect 24118 5013 24298 5025
rect 24118 4961 24130 5013
rect 24182 4961 24234 5013
rect 24286 4961 24298 5013
rect 24118 4909 24298 4961
rect 24118 4906 24130 4909
rect 24182 4906 24234 4909
rect 24286 4906 24298 4909
rect 24838 4997 26210 5193
rect 24838 4906 25034 4997
rect 26014 4906 26210 4997
rect 23662 4860 23673 4906
rect 23847 4860 23858 4906
rect 24110 4860 24121 4906
rect 24295 4860 24569 4906
rect 24743 4860 24754 4906
rect 24838 4860 24849 4906
rect 25023 4860 25034 4906
rect 25286 4860 25297 4906
rect 25471 4860 25577 4906
rect 25751 4860 25762 4906
rect 26014 4860 26025 4906
rect 26199 4860 26210 4906
rect 26294 4997 27666 5193
rect 26294 4906 26490 4997
rect 27470 4906 27666 4997
rect 26294 4860 26305 4906
rect 26479 4860 26490 4906
rect 26742 4860 26753 4906
rect 26927 4860 27033 4906
rect 27207 4860 27218 4906
rect 27470 4860 27481 4906
rect 27655 4860 27666 4906
rect 27942 4906 28138 5491
rect 27942 4860 27953 4906
rect 28127 4860 28138 4906
rect 23662 3774 23858 4860
rect 24118 4857 24130 4860
rect 24182 4857 24234 4860
rect 24286 4857 24298 4860
rect 24118 4845 24298 4857
rect 27480 4305 27660 4317
rect 27042 4253 27492 4305
rect 27544 4253 27596 4305
rect 27648 4253 27660 4305
rect 27042 4201 27660 4253
rect 27042 4149 27492 4201
rect 27544 4149 27596 4201
rect 27648 4149 27660 4201
rect 27042 3774 27202 4149
rect 27480 4137 27660 4149
rect 27942 3774 28138 4860
rect 23662 3728 23673 3774
rect 23847 3728 23858 3774
rect 23662 2934 23858 3728
rect 24110 3728 24121 3774
rect 24295 3728 24306 3774
rect 24558 3728 24569 3774
rect 24743 3728 24849 3774
rect 25023 3728 25034 3774
rect 25286 3728 25297 3774
rect 25471 3728 25482 3774
rect 24110 3637 24306 3728
rect 25286 3637 25482 3728
rect 24110 3441 25482 3637
rect 25566 3728 25577 3774
rect 25751 3728 25762 3774
rect 26014 3728 26025 3774
rect 26199 3728 26305 3774
rect 26479 3728 26490 3774
rect 26742 3728 26753 3774
rect 26927 3728 26938 3774
rect 27022 3728 27033 3774
rect 27207 3728 27218 3774
rect 27470 3728 27481 3774
rect 27655 3728 27666 3774
rect 25566 3637 25762 3728
rect 26742 3637 26938 3728
rect 25566 3441 26938 3637
rect 27470 3421 27666 3728
rect 27022 3225 27666 3421
rect 27942 3728 27953 3774
rect 28127 3728 28138 3774
rect 23662 2888 23673 2934
rect 23847 2888 23858 2934
rect 24110 3025 25482 3221
rect 24110 2934 24306 3025
rect 25286 2934 25482 3025
rect 24110 2888 24121 2934
rect 24295 2888 24306 2934
rect 24558 2888 24569 2934
rect 24743 2888 24849 2934
rect 25023 2888 25034 2934
rect 25286 2888 25297 2934
rect 25471 2888 25482 2934
rect 25566 3025 26938 3221
rect 25566 2934 25762 3025
rect 26742 2934 26938 3025
rect 25566 2888 25577 2934
rect 25751 2888 25762 2934
rect 26014 2888 26025 2934
rect 26199 2888 26305 2934
rect 26479 2888 26490 2934
rect 26742 2888 26753 2934
rect 26927 2888 26938 2934
rect 27022 2934 27218 3225
rect 27478 2937 27658 2949
rect 27478 2934 27490 2937
rect 27542 2934 27594 2937
rect 27646 2934 27658 2937
rect 27942 2934 28138 3728
rect 27022 2888 27033 2934
rect 27207 2888 27218 2934
rect 27470 2888 27481 2934
rect 27655 2888 27666 2934
rect 27942 2888 27953 2934
rect 28127 2888 28138 2934
rect 23662 1802 23858 2888
rect 27478 2885 27490 2888
rect 27542 2885 27594 2888
rect 27646 2885 27658 2888
rect 27478 2833 27658 2885
rect 27478 2781 27490 2833
rect 27542 2781 27594 2833
rect 27646 2781 27658 2833
rect 27478 2769 27658 2781
rect 24118 1805 24298 1817
rect 24118 1802 24130 1805
rect 24182 1802 24234 1805
rect 24286 1802 24298 1805
rect 24568 1805 24748 1819
rect 24568 1802 24578 1805
rect 24630 1802 24682 1805
rect 24734 1802 24748 1805
rect 27942 1802 28138 2888
rect 23662 1756 23673 1802
rect 23847 1756 23858 1802
rect 24110 1756 24121 1802
rect 24295 1756 24306 1802
rect 24558 1756 24569 1802
rect 24743 1756 24754 1802
rect 24838 1756 24849 1802
rect 25023 1756 25034 1802
rect 25286 1756 25297 1802
rect 25471 1756 25577 1802
rect 25751 1756 25762 1802
rect 26014 1756 26025 1802
rect 26199 1756 26210 1802
rect 23662 1259 23858 1756
rect 24118 1753 24130 1756
rect 24182 1753 24234 1756
rect 24286 1753 24298 1756
rect 24118 1701 24298 1753
rect 24118 1649 24130 1701
rect 24182 1649 24234 1701
rect 24286 1649 24298 1701
rect 24118 1637 24298 1649
rect 24568 1753 24578 1756
rect 24630 1753 24682 1756
rect 24734 1753 24748 1756
rect 24568 1701 24748 1753
rect 24568 1649 24578 1701
rect 24630 1649 24682 1701
rect 24734 1649 24748 1701
rect 24568 1639 24748 1649
rect 24838 1665 25034 1756
rect 26014 1665 26210 1756
rect 24838 1469 26210 1665
rect 26294 1756 26305 1802
rect 26479 1756 26490 1802
rect 26742 1756 26753 1802
rect 26927 1756 27033 1802
rect 27207 1756 27218 1802
rect 27470 1756 27481 1802
rect 27655 1756 27666 1802
rect 26294 1665 26490 1756
rect 27470 1665 27666 1756
rect 26294 1469 27666 1665
rect 27942 1756 27953 1802
rect 28127 1756 28138 1802
rect 27942 1259 28138 1756
rect 28590 5467 28734 5491
rect 28780 5491 31742 5513
rect 28780 5467 28910 5491
rect 28590 5419 28910 5467
rect 28590 5373 28734 5419
rect 28780 5373 28910 5419
rect 28590 5325 28910 5373
rect 28590 5279 28734 5325
rect 28780 5279 28910 5325
rect 28590 5231 28910 5279
rect 28590 5185 28734 5231
rect 28780 5185 28910 5231
rect 28590 5137 28910 5185
rect 28590 5091 28734 5137
rect 28780 5091 28910 5137
rect 28590 5043 28910 5091
rect 28590 4997 28734 5043
rect 28780 4997 28910 5043
rect 28590 4949 28910 4997
rect 28590 4903 28734 4949
rect 28780 4903 28910 4949
rect 28590 4855 28910 4903
rect 28590 4809 28734 4855
rect 28780 4809 28910 4855
rect 28590 4761 28910 4809
rect 28590 4715 28734 4761
rect 28780 4715 28910 4761
rect 28590 4667 28910 4715
rect 28590 4621 28734 4667
rect 28780 4621 28910 4667
rect 28590 4573 28910 4621
rect 28590 4527 28734 4573
rect 28780 4527 28910 4573
rect 28590 4479 28910 4527
rect 28590 4433 28734 4479
rect 28780 4433 28910 4479
rect 28590 4385 28910 4433
rect 28590 4339 28734 4385
rect 28780 4339 28910 4385
rect 28590 4291 28910 4339
rect 28590 4245 28734 4291
rect 28780 4245 28910 4291
rect 28590 4197 28910 4245
rect 28590 4151 28734 4197
rect 28780 4151 28910 4197
rect 28590 4103 28910 4151
rect 28590 4057 28734 4103
rect 28780 4057 28910 4103
rect 28590 4009 28910 4057
rect 28590 3963 28734 4009
rect 28780 3963 28910 4009
rect 28590 3915 28910 3963
rect 28590 3869 28734 3915
rect 28780 3869 28910 3915
rect 28590 3821 28910 3869
rect 28590 3775 28734 3821
rect 28780 3775 28910 3821
rect 28590 3727 28910 3775
rect 28590 3681 28734 3727
rect 28780 3681 28910 3727
rect 28590 3633 28910 3681
rect 29288 5090 29484 5491
rect 29288 5044 29299 5090
rect 29473 5044 29484 5090
rect 29288 3718 29484 5044
rect 29736 5093 30780 5105
rect 29736 5090 30300 5093
rect 30352 5090 30404 5093
rect 30456 5090 30508 5093
rect 29736 5044 29747 5090
rect 29921 5044 30027 5090
rect 30201 5044 30300 5090
rect 30481 5044 30508 5090
rect 29736 5041 30300 5044
rect 30352 5041 30404 5044
rect 30456 5041 30508 5044
rect 30560 5090 30612 5093
rect 30664 5090 30716 5093
rect 30560 5044 30587 5090
rect 30560 5041 30612 5044
rect 30664 5041 30716 5044
rect 30768 5041 30780 5093
rect 29736 4989 30780 5041
rect 29736 4937 30300 4989
rect 30352 4937 30404 4989
rect 30456 4937 30508 4989
rect 30560 4937 30612 4989
rect 30664 4937 30716 4989
rect 30768 4937 30780 4989
rect 29736 4885 30780 4937
rect 29736 4833 30300 4885
rect 30352 4833 30404 4885
rect 30456 4833 30508 4885
rect 30560 4833 30612 4885
rect 30664 4833 30716 4885
rect 30768 4833 30780 4885
rect 29736 4821 30780 4833
rect 31024 5090 31220 5491
rect 31024 5044 31035 5090
rect 31209 5044 31220 5090
rect 29288 3672 29299 3718
rect 29473 3672 29484 3718
rect 29736 4137 30780 4149
rect 29736 4085 30300 4137
rect 30352 4085 30404 4137
rect 30456 4085 30508 4137
rect 30560 4085 30612 4137
rect 30664 4085 30716 4137
rect 30768 4085 30780 4137
rect 29736 4033 30780 4085
rect 29736 3981 30300 4033
rect 30352 3981 30404 4033
rect 30456 3981 30508 4033
rect 30560 3981 30612 4033
rect 30664 3981 30716 4033
rect 30768 3981 30780 4033
rect 29736 3929 30780 3981
rect 29736 3877 30300 3929
rect 30352 3877 30404 3929
rect 30456 3877 30508 3929
rect 30560 3877 30612 3929
rect 30664 3877 30716 3929
rect 30768 3877 30780 3929
rect 29736 3825 30780 3877
rect 29736 3773 30300 3825
rect 30352 3773 30404 3825
rect 30456 3773 30508 3825
rect 30560 3773 30612 3825
rect 30664 3773 30716 3825
rect 30768 3773 30780 3825
rect 29736 3721 30780 3773
rect 29736 3718 30300 3721
rect 30352 3718 30404 3721
rect 30456 3718 30508 3721
rect 29736 3672 29747 3718
rect 29921 3672 30027 3718
rect 30201 3672 30300 3718
rect 30481 3672 30508 3718
rect 29736 3669 30300 3672
rect 30352 3669 30404 3672
rect 30456 3669 30508 3672
rect 30560 3718 30612 3721
rect 30664 3718 30716 3721
rect 30560 3672 30587 3718
rect 30560 3669 30612 3672
rect 30664 3669 30716 3672
rect 30768 3669 30780 3721
rect 31024 3718 31220 5044
rect 31024 3672 31035 3718
rect 31209 3672 31220 3718
rect 31598 5467 31742 5491
rect 31788 5467 31918 5513
rect 31598 5419 31918 5467
rect 31598 5373 31742 5419
rect 31788 5373 31918 5419
rect 31598 5325 31918 5373
rect 31598 5279 31742 5325
rect 31788 5279 31918 5325
rect 31598 5231 31918 5279
rect 31598 5185 31742 5231
rect 31788 5185 31918 5231
rect 31598 5137 31918 5185
rect 31598 5091 31742 5137
rect 31788 5091 31918 5137
rect 31598 5043 31918 5091
rect 31598 4997 31742 5043
rect 31788 4997 31918 5043
rect 31598 4949 31918 4997
rect 31598 4903 31742 4949
rect 31788 4903 31918 4949
rect 31598 4855 31918 4903
rect 31598 4809 31742 4855
rect 31788 4809 31918 4855
rect 31598 4761 31918 4809
rect 31598 4715 31742 4761
rect 31788 4715 31918 4761
rect 31598 4667 31918 4715
rect 31598 4621 31742 4667
rect 31788 4621 31918 4667
rect 31598 4573 31918 4621
rect 31598 4527 31742 4573
rect 31788 4527 31918 4573
rect 31598 4479 31918 4527
rect 31598 4433 31742 4479
rect 31788 4433 31918 4479
rect 31598 4385 31918 4433
rect 31598 4339 31742 4385
rect 31788 4339 31918 4385
rect 31598 4291 31918 4339
rect 31598 4245 31742 4291
rect 31788 4245 31918 4291
rect 31598 4197 31918 4245
rect 31598 4151 31742 4197
rect 31788 4151 31918 4197
rect 31598 4103 31918 4151
rect 31598 4057 31742 4103
rect 31788 4057 31918 4103
rect 31598 4009 31918 4057
rect 31598 3963 31742 4009
rect 31788 3963 31918 4009
rect 31598 3915 31918 3963
rect 31598 3869 31742 3915
rect 31788 3869 31918 3915
rect 31598 3821 31918 3869
rect 31598 3775 31742 3821
rect 31788 3775 31918 3821
rect 31598 3727 31918 3775
rect 31598 3681 31742 3727
rect 31788 3681 31918 3727
rect 29736 3657 30780 3669
rect 28590 3587 28734 3633
rect 28780 3587 28910 3633
rect 28590 3539 28910 3587
rect 28590 3493 28734 3539
rect 28780 3493 28910 3539
rect 28590 3445 28910 3493
rect 28590 3399 28734 3445
rect 28780 3399 28910 3445
rect 28590 3351 28910 3399
rect 28590 3305 28734 3351
rect 28780 3305 28910 3351
rect 28590 3257 28910 3305
rect 28590 3211 28734 3257
rect 28780 3211 28910 3257
rect 28590 3163 28910 3211
rect 28590 3117 28734 3163
rect 28780 3117 28910 3163
rect 28590 3069 28910 3117
rect 31598 3633 31918 3681
rect 31598 3587 31742 3633
rect 31788 3587 31918 3633
rect 31598 3539 31918 3587
rect 31598 3493 31742 3539
rect 31788 3493 31918 3539
rect 31598 3445 31918 3493
rect 31598 3399 31742 3445
rect 31788 3399 31918 3445
rect 31598 3351 31918 3399
rect 31598 3305 31742 3351
rect 31788 3305 31918 3351
rect 31598 3257 31918 3305
rect 31598 3211 31742 3257
rect 31788 3211 31918 3257
rect 31598 3163 31918 3211
rect 31598 3117 31742 3163
rect 31788 3117 31918 3163
rect 29728 3081 30772 3093
rect 28590 3023 28734 3069
rect 28780 3023 28910 3069
rect 28590 2975 28910 3023
rect 28590 2929 28734 2975
rect 28780 2929 28910 2975
rect 28590 2881 28910 2929
rect 28590 2835 28734 2881
rect 28780 2835 28910 2881
rect 28590 2787 28910 2835
rect 28590 2741 28734 2787
rect 28780 2741 28910 2787
rect 28590 2693 28910 2741
rect 28590 2647 28734 2693
rect 28780 2647 28910 2693
rect 28590 2599 28910 2647
rect 28590 2553 28734 2599
rect 28780 2553 28910 2599
rect 28590 2505 28910 2553
rect 28590 2459 28734 2505
rect 28780 2459 28910 2505
rect 28590 2411 28910 2459
rect 28590 2365 28734 2411
rect 28780 2365 28910 2411
rect 28590 2317 28910 2365
rect 28590 2271 28734 2317
rect 28780 2271 28910 2317
rect 28590 2223 28910 2271
rect 28590 2177 28734 2223
rect 28780 2177 28910 2223
rect 28590 2129 28910 2177
rect 28590 2083 28734 2129
rect 28780 2083 28910 2129
rect 28590 2035 28910 2083
rect 28590 1989 28734 2035
rect 28780 1989 28910 2035
rect 28590 1941 28910 1989
rect 28590 1895 28734 1941
rect 28780 1895 28910 1941
rect 28590 1847 28910 1895
rect 28590 1801 28734 1847
rect 28780 1801 28910 1847
rect 28590 1753 28910 1801
rect 28590 1707 28734 1753
rect 28780 1707 28910 1753
rect 28590 1659 28910 1707
rect 28590 1613 28734 1659
rect 28780 1613 28910 1659
rect 28590 1565 28910 1613
rect 28590 1519 28734 1565
rect 28780 1519 28910 1565
rect 28590 1471 28910 1519
rect 28590 1425 28734 1471
rect 28780 1425 28910 1471
rect 28590 1377 28910 1425
rect 28590 1331 28734 1377
rect 28780 1331 28910 1377
rect 28590 1283 28910 1331
rect 28590 1259 28734 1283
rect 23046 1237 28734 1259
rect 28780 1259 28910 1283
rect 29288 3032 29299 3078
rect 29473 3032 29484 3078
rect 29288 1706 29484 3032
rect 29728 3029 29740 3081
rect 29792 3078 29844 3081
rect 29896 3078 29948 3081
rect 29921 3032 29948 3078
rect 29792 3029 29844 3032
rect 29896 3029 29948 3032
rect 30000 3078 30052 3081
rect 30104 3078 30156 3081
rect 30208 3078 30772 3081
rect 30000 3032 30027 3078
rect 30208 3032 30307 3078
rect 30481 3032 30587 3078
rect 30761 3032 30772 3078
rect 30000 3029 30052 3032
rect 30104 3029 30156 3032
rect 30208 3029 30772 3032
rect 29728 2977 30772 3029
rect 29728 2925 29740 2977
rect 29792 2925 29844 2977
rect 29896 2925 29948 2977
rect 30000 2925 30052 2977
rect 30104 2925 30156 2977
rect 30208 2925 30772 2977
rect 29728 2873 30772 2925
rect 29728 2821 29740 2873
rect 29792 2821 29844 2873
rect 29896 2821 29948 2873
rect 30000 2821 30052 2873
rect 30104 2821 30156 2873
rect 30208 2821 30772 2873
rect 29728 2809 30772 2821
rect 31024 3032 31035 3078
rect 31209 3032 31220 3078
rect 29288 1660 29299 1706
rect 29473 1660 29484 1706
rect 29288 1259 29484 1660
rect 29736 2125 30780 2137
rect 29736 2073 30300 2125
rect 30352 2073 30404 2125
rect 30456 2073 30508 2125
rect 30560 2073 30612 2125
rect 30664 2073 30716 2125
rect 30768 2073 30780 2125
rect 29736 2021 30780 2073
rect 29736 1969 30300 2021
rect 30352 1969 30404 2021
rect 30456 1969 30508 2021
rect 30560 1969 30612 2021
rect 30664 1969 30716 2021
rect 30768 1969 30780 2021
rect 29736 1917 30780 1969
rect 29736 1865 30300 1917
rect 30352 1865 30404 1917
rect 30456 1865 30508 1917
rect 30560 1865 30612 1917
rect 30664 1865 30716 1917
rect 30768 1865 30780 1917
rect 29736 1813 30780 1865
rect 29736 1761 30300 1813
rect 30352 1761 30404 1813
rect 30456 1761 30508 1813
rect 30560 1761 30612 1813
rect 30664 1761 30716 1813
rect 30768 1761 30780 1813
rect 29736 1709 30780 1761
rect 29736 1706 30300 1709
rect 30352 1706 30404 1709
rect 30456 1706 30508 1709
rect 29736 1660 29747 1706
rect 29921 1660 30027 1706
rect 30201 1660 30300 1706
rect 30481 1660 30508 1706
rect 29736 1657 30300 1660
rect 30352 1657 30404 1660
rect 30456 1657 30508 1660
rect 30560 1706 30612 1709
rect 30664 1706 30716 1709
rect 30560 1660 30587 1706
rect 30560 1657 30612 1660
rect 30664 1657 30716 1660
rect 30768 1657 30780 1709
rect 29736 1645 30780 1657
rect 31024 1706 31220 3032
rect 31024 1660 31035 1706
rect 31209 1660 31220 1706
rect 31024 1259 31220 1660
rect 31598 3069 31918 3117
rect 31598 3023 31742 3069
rect 31788 3023 31918 3069
rect 31598 2975 31918 3023
rect 31598 2929 31742 2975
rect 31788 2929 31918 2975
rect 31598 2881 31918 2929
rect 31598 2835 31742 2881
rect 31788 2835 31918 2881
rect 31598 2787 31918 2835
rect 31598 2741 31742 2787
rect 31788 2741 31918 2787
rect 31598 2693 31918 2741
rect 31598 2647 31742 2693
rect 31788 2647 31918 2693
rect 31598 2599 31918 2647
rect 31598 2553 31742 2599
rect 31788 2553 31918 2599
rect 31598 2505 31918 2553
rect 31598 2459 31742 2505
rect 31788 2459 31918 2505
rect 31598 2411 31918 2459
rect 31598 2365 31742 2411
rect 31788 2365 31918 2411
rect 31598 2317 31918 2365
rect 31598 2271 31742 2317
rect 31788 2271 31918 2317
rect 31598 2223 31918 2271
rect 31598 2177 31742 2223
rect 31788 2177 31918 2223
rect 31598 2129 31918 2177
rect 31598 2083 31742 2129
rect 31788 2083 31918 2129
rect 31598 2035 31918 2083
rect 31598 1989 31742 2035
rect 31788 1989 31918 2035
rect 31598 1941 31918 1989
rect 31598 1895 31742 1941
rect 31788 1895 31918 1941
rect 31598 1847 31918 1895
rect 31598 1801 31742 1847
rect 31788 1801 31918 1847
rect 31598 1753 31918 1801
rect 31598 1707 31742 1753
rect 31788 1707 31918 1753
rect 31598 1659 31918 1707
rect 31598 1613 31742 1659
rect 31788 1613 31918 1659
rect 31598 1565 31918 1613
rect 31598 1519 31742 1565
rect 31788 1519 31918 1565
rect 31598 1471 31918 1519
rect 31598 1425 31742 1471
rect 31788 1425 31918 1471
rect 31598 1377 31918 1425
rect 31598 1331 31742 1377
rect 31788 1331 31918 1377
rect 31598 1283 31918 1331
rect 31598 1259 31742 1283
rect 28780 1237 31742 1259
rect 31788 1237 31918 1283
rect 18076 1189 31918 1237
rect 18076 1143 18206 1189
rect 18252 1143 23000 1189
rect 23046 1143 28734 1189
rect 28780 1143 31742 1189
rect 31788 1143 31918 1189
rect 12018 1131 12198 1139
rect 12018 1127 12486 1131
rect 12018 1075 12030 1127
rect 12082 1075 12134 1127
rect 12186 1075 12486 1127
rect 12018 1023 12486 1075
rect 12018 971 12030 1023
rect 12082 971 12134 1023
rect 12186 971 12486 1023
rect 18076 1095 31918 1143
rect 45022 1201 50632 1213
rect 45022 1149 45034 1201
rect 45086 1149 45138 1201
rect 45190 1149 45242 1201
rect 45294 1149 45346 1201
rect 45398 1149 45450 1201
rect 45502 1149 49474 1201
rect 49526 1149 49578 1201
rect 49630 1149 49682 1201
rect 49734 1149 49786 1201
rect 49838 1149 49890 1201
rect 49942 1149 50632 1201
rect 18076 1049 18206 1095
rect 18252 1049 18300 1095
rect 18346 1049 18394 1095
rect 18440 1049 18488 1095
rect 18534 1049 18582 1095
rect 18628 1049 18676 1095
rect 18722 1049 18770 1095
rect 18816 1049 18864 1095
rect 18910 1049 18958 1095
rect 19004 1049 19052 1095
rect 19098 1049 19146 1095
rect 19192 1049 19240 1095
rect 19286 1049 19334 1095
rect 19380 1049 19428 1095
rect 19474 1049 19522 1095
rect 19568 1049 19616 1095
rect 19662 1049 19710 1095
rect 19756 1049 19804 1095
rect 19850 1049 19898 1095
rect 19944 1049 19992 1095
rect 20038 1049 20086 1095
rect 20132 1049 20180 1095
rect 20226 1049 20274 1095
rect 20320 1049 20368 1095
rect 20414 1049 20462 1095
rect 20508 1049 20556 1095
rect 20602 1049 20650 1095
rect 20696 1049 20744 1095
rect 20790 1049 20838 1095
rect 20884 1049 20932 1095
rect 20978 1049 21026 1095
rect 21072 1049 21120 1095
rect 21166 1049 21214 1095
rect 21260 1049 21308 1095
rect 21354 1049 21402 1095
rect 21448 1049 21496 1095
rect 21542 1049 21590 1095
rect 21636 1049 21684 1095
rect 21730 1049 21778 1095
rect 21824 1049 21872 1095
rect 21918 1049 21966 1095
rect 22012 1049 22060 1095
rect 22106 1049 22154 1095
rect 22200 1049 22248 1095
rect 22294 1049 22342 1095
rect 22388 1049 22436 1095
rect 22482 1049 22530 1095
rect 22576 1049 22624 1095
rect 22670 1049 22718 1095
rect 22764 1049 22812 1095
rect 22858 1049 22906 1095
rect 22952 1049 23000 1095
rect 23046 1049 23094 1095
rect 23140 1049 23188 1095
rect 23234 1049 23282 1095
rect 23328 1049 23376 1095
rect 23422 1049 23470 1095
rect 23516 1049 23564 1095
rect 23610 1049 23658 1095
rect 23704 1049 23752 1095
rect 23798 1049 23846 1095
rect 23892 1049 23940 1095
rect 23986 1049 24034 1095
rect 24080 1049 24128 1095
rect 24174 1049 24222 1095
rect 24268 1049 24316 1095
rect 24362 1049 24410 1095
rect 24456 1049 24504 1095
rect 24550 1049 24598 1095
rect 24644 1049 24692 1095
rect 24738 1049 24786 1095
rect 24832 1049 24880 1095
rect 24926 1049 24974 1095
rect 25020 1049 25068 1095
rect 25114 1049 25162 1095
rect 25208 1049 25256 1095
rect 25302 1049 25350 1095
rect 25396 1049 25444 1095
rect 25490 1049 25538 1095
rect 25584 1049 25632 1095
rect 25678 1049 25726 1095
rect 25772 1049 25820 1095
rect 25866 1049 25914 1095
rect 25960 1049 26008 1095
rect 26054 1049 26102 1095
rect 26148 1049 26196 1095
rect 26242 1049 26290 1095
rect 26336 1049 26384 1095
rect 26430 1049 26478 1095
rect 26524 1049 26572 1095
rect 26618 1049 26666 1095
rect 26712 1049 26760 1095
rect 26806 1049 26854 1095
rect 26900 1049 26948 1095
rect 26994 1049 27042 1095
rect 27088 1049 27136 1095
rect 27182 1049 27230 1095
rect 27276 1049 27324 1095
rect 27370 1049 27418 1095
rect 27464 1049 27512 1095
rect 27558 1049 27606 1095
rect 27652 1049 27700 1095
rect 27746 1049 27794 1095
rect 27840 1049 27888 1095
rect 27934 1049 27982 1095
rect 28028 1049 28076 1095
rect 28122 1049 28170 1095
rect 28216 1049 28264 1095
rect 28310 1049 28358 1095
rect 28404 1049 28452 1095
rect 28498 1049 28546 1095
rect 28592 1049 28640 1095
rect 28686 1049 28734 1095
rect 28780 1049 28828 1095
rect 28874 1049 28922 1095
rect 28968 1049 29016 1095
rect 29062 1049 29110 1095
rect 29156 1049 29204 1095
rect 29250 1049 29298 1095
rect 29344 1049 29392 1095
rect 29438 1049 29486 1095
rect 29532 1049 29580 1095
rect 29626 1049 29674 1095
rect 29720 1049 29768 1095
rect 29814 1049 29862 1095
rect 29908 1049 29956 1095
rect 30002 1049 30050 1095
rect 30096 1049 30144 1095
rect 30190 1049 30238 1095
rect 30284 1049 30332 1095
rect 30378 1049 30426 1095
rect 30472 1049 30520 1095
rect 30566 1049 30614 1095
rect 30660 1049 30708 1095
rect 30754 1049 30802 1095
rect 30848 1049 30896 1095
rect 30942 1049 30990 1095
rect 31036 1049 31084 1095
rect 31130 1049 31178 1095
rect 31224 1049 31272 1095
rect 31318 1049 31366 1095
rect 31412 1049 31460 1095
rect 31506 1049 31554 1095
rect 31600 1049 31648 1095
rect 31694 1049 31742 1095
rect 31788 1049 31918 1095
rect 12018 959 12198 971
rect 18076 939 31918 1049
rect 35192 1101 40802 1113
rect 35192 1049 35204 1101
rect 35256 1049 35308 1101
rect 35360 1049 35412 1101
rect 35464 1049 35516 1101
rect 35568 1049 35620 1101
rect 35672 1049 39644 1101
rect 39696 1049 39748 1101
rect 39800 1049 39852 1101
rect 39904 1049 39956 1101
rect 40008 1049 40060 1101
rect 40112 1049 40802 1101
rect 35192 997 40802 1049
rect 35192 945 35204 997
rect 35256 945 35308 997
rect 35360 945 35412 997
rect 35464 945 35516 997
rect 35568 945 35620 997
rect 35672 945 39644 997
rect 39696 945 39748 997
rect 39800 945 39852 997
rect 39904 945 39956 997
rect 40008 945 40060 997
rect 40112 945 40802 997
rect 35192 893 40802 945
rect 35192 841 35204 893
rect 35256 841 35308 893
rect 35360 841 35412 893
rect 35464 841 35516 893
rect 35568 841 35620 893
rect 35672 841 39644 893
rect 39696 841 39748 893
rect 39800 841 39852 893
rect 39904 841 39956 893
rect 40008 841 40060 893
rect 40112 841 40802 893
rect 35192 789 40802 841
rect 21631 772 22475 784
rect 21631 720 21643 772
rect 21695 720 21747 772
rect 21799 720 21851 772
rect 21903 720 22475 772
rect 21631 668 22475 720
rect 21631 616 21643 668
rect 21695 616 21747 668
rect 21799 616 21851 668
rect 21903 616 22475 668
rect 35192 737 35204 789
rect 35256 737 35308 789
rect 35360 737 35412 789
rect 35464 737 35516 789
rect 35568 737 35620 789
rect 35672 737 39644 789
rect 39696 737 39748 789
rect 39800 737 39852 789
rect 39904 737 39956 789
rect 40008 737 40060 789
rect 40112 737 40802 789
rect 35192 685 40802 737
rect 45022 1097 50632 1149
rect 45022 1045 45034 1097
rect 45086 1045 45138 1097
rect 45190 1045 45242 1097
rect 45294 1045 45346 1097
rect 45398 1045 45450 1097
rect 45502 1045 49474 1097
rect 49526 1045 49578 1097
rect 49630 1045 49682 1097
rect 49734 1045 49786 1097
rect 49838 1045 49890 1097
rect 49942 1045 50632 1097
rect 45022 993 50632 1045
rect 45022 941 45034 993
rect 45086 941 45138 993
rect 45190 941 45242 993
rect 45294 941 45346 993
rect 45398 941 45450 993
rect 45502 941 49474 993
rect 49526 941 49578 993
rect 49630 941 49682 993
rect 49734 941 49786 993
rect 49838 941 49890 993
rect 49942 941 50632 993
rect 45022 889 50632 941
rect 45022 837 45034 889
rect 45086 837 45138 889
rect 45190 837 45242 889
rect 45294 837 45346 889
rect 45398 837 45450 889
rect 45502 837 49474 889
rect 49526 837 49578 889
rect 49630 837 49682 889
rect 49734 837 49786 889
rect 49838 837 49890 889
rect 49942 837 50632 889
rect 45022 785 50632 837
rect 45022 733 45034 785
rect 45086 733 45138 785
rect 45190 733 45242 785
rect 45294 733 45346 785
rect 45398 733 45450 785
rect 45502 733 49474 785
rect 49526 733 49578 785
rect 49630 733 49682 785
rect 49734 733 49786 785
rect 49838 733 49890 785
rect 49942 733 50632 785
rect 45022 721 50632 733
rect 35192 633 35204 685
rect 35256 633 35308 685
rect 35360 633 35412 685
rect 35464 633 35516 685
rect 35568 633 35620 685
rect 35672 633 39644 685
rect 39696 633 39748 685
rect 39800 633 39852 685
rect 39904 633 39956 685
rect 40008 633 40060 685
rect 40112 633 40802 685
rect 35192 621 40802 633
rect 21631 564 22475 616
rect 21631 512 21643 564
rect 21695 512 21747 564
rect 21799 512 21851 564
rect 21903 512 22475 564
rect 21631 500 22475 512
rect 15556 272 16342 284
rect 15556 220 15568 272
rect 15620 220 15672 272
rect 15724 220 15776 272
rect 15828 220 16342 272
rect 15556 168 16342 220
rect 15556 116 15568 168
rect 15620 116 15672 168
rect 15724 116 15776 168
rect 15828 116 16342 168
rect 15556 64 16342 116
rect 15556 12 15568 64
rect 15620 12 15672 64
rect 15724 12 15776 64
rect 15828 12 16342 64
rect 15556 0 16342 12
rect -17226 -227 292 -83
rect -17258 -387 292 -227
<< via1 >>
rect 31230 15653 31282 15705
rect 31334 15653 31386 15705
rect 31438 15653 31490 15705
rect 31230 15549 31282 15601
rect 31334 15549 31386 15601
rect 31438 15549 31490 15601
rect 31230 15445 31282 15497
rect 31334 15445 31386 15497
rect 31438 15445 31490 15497
rect 32144 15067 32196 15119
rect 32248 15067 32300 15119
rect 32352 15067 32404 15119
rect 32144 14963 32196 15015
rect 32248 14963 32300 15015
rect 32352 14963 32404 15015
rect 32144 14859 32196 14911
rect 32248 14859 32300 14911
rect 32352 14859 32404 14911
rect 1812 14265 1868 14321
rect 1922 14265 1978 14321
rect 2032 14265 2088 14321
rect 2142 14265 2198 14321
rect 3173 14274 3225 14326
rect 3277 14274 3329 14326
rect 1812 14155 1868 14211
rect 1922 14155 1978 14211
rect 2032 14155 2088 14211
rect 2142 14155 2198 14211
rect 3173 14170 3225 14222
rect 3277 14170 3329 14222
rect 1812 14045 1868 14101
rect 1922 14045 1978 14101
rect 2032 14045 2088 14101
rect 2142 14045 2198 14101
rect 2532 13925 2584 13977
rect 2636 13925 2688 13977
rect 2532 13821 2584 13873
rect 2636 13821 2688 13873
rect 2893 13146 2945 13198
rect 2997 13146 3049 13198
rect 2893 13042 2945 13094
rect 2997 13042 3049 13094
rect -3594 10371 -3538 10427
rect -3484 10371 -3428 10427
rect -7089 10310 -7033 10345
rect -6979 10310 -6923 10345
rect -7089 10289 -7033 10310
rect -6979 10289 -6923 10310
rect -6809 10310 -6753 10345
rect -6699 10310 -6643 10345
rect -6809 10289 -6753 10310
rect -6699 10289 -6643 10310
rect -3594 10261 -3538 10317
rect -3484 10261 -3428 10317
rect -3594 10151 -3538 10207
rect -3484 10151 -3428 10207
rect -3594 10041 -3538 10097
rect -3484 10041 -3428 10097
rect -3594 9931 -3538 9987
rect -3484 9931 -3428 9987
rect -4569 9764 -4513 9780
rect -4459 9764 -4403 9780
rect -4569 9724 -4513 9764
rect -4459 9724 -4403 9764
rect -7089 9393 -7033 9428
rect -6979 9393 -6923 9428
rect -5409 9393 -5353 9428
rect -5299 9393 -5243 9428
rect -4569 9393 -4513 9428
rect -4459 9393 -4403 9428
rect -7089 9372 -7033 9393
rect -6979 9372 -6923 9393
rect -5409 9372 -5353 9393
rect -5299 9372 -5243 9393
rect -4569 9372 -4513 9393
rect -4459 9372 -4403 9393
rect -6809 8847 -6753 8863
rect -6699 8847 -6643 8863
rect -4849 8847 -4793 8863
rect -4739 8847 -4683 8863
rect -6809 8807 -6753 8847
rect -6699 8807 -6643 8847
rect -4849 8807 -4793 8847
rect -4739 8807 -4683 8847
rect -7089 8476 -7033 8511
rect -6979 8476 -6923 8511
rect -7089 8455 -7033 8476
rect -6979 8455 -6923 8476
rect -4569 8476 -4513 8511
rect -4459 8476 -4403 8511
rect -4569 8455 -4513 8476
rect -4459 8455 -4403 8476
rect 238 7531 290 7583
rect 342 7531 394 7583
rect -7089 6516 -7033 6537
rect -6979 6516 -6923 6537
rect -7089 6481 -7033 6516
rect -6979 6481 -6923 6516
rect -4569 6516 -4513 6537
rect -4459 6516 -4403 6537
rect -4569 6481 -4513 6516
rect -4459 6481 -4403 6516
rect -6809 6145 -6753 6185
rect -6699 6145 -6643 6185
rect -4849 6145 -4793 6185
rect -4739 6145 -4683 6185
rect -6809 6129 -6753 6145
rect -6699 6129 -6643 6145
rect -4849 6129 -4793 6145
rect -4739 6129 -4683 6145
rect -7089 5599 -7033 5620
rect -6979 5599 -6923 5620
rect -5409 5599 -5353 5620
rect -5299 5599 -5243 5620
rect -4569 5599 -4513 5620
rect -4459 5599 -4403 5620
rect -7089 5564 -7033 5599
rect -6979 5564 -6923 5599
rect -5409 5564 -5353 5599
rect -5299 5564 -5243 5599
rect -4569 5564 -4513 5599
rect -4459 5564 -4403 5599
rect -4569 5228 -4513 5268
rect -4459 5228 -4403 5268
rect -4569 5212 -4513 5228
rect -4459 5212 -4403 5228
rect -7089 4682 -7033 4703
rect -6979 4682 -6923 4703
rect -7089 4647 -7033 4682
rect -6979 4647 -6923 4682
rect -6809 4682 -6753 4703
rect -6699 4682 -6643 4703
rect -6809 4647 -6753 4682
rect -6699 4647 -6643 4682
rect 238 7427 290 7479
rect 342 7427 394 7479
rect 1239 7580 1291 7583
rect 1239 7534 1242 7580
rect 1242 7534 1288 7580
rect 1288 7534 1291 7580
rect 1239 7531 1291 7534
rect 1343 7580 1395 7583
rect 1343 7534 1346 7580
rect 1346 7534 1392 7580
rect 1392 7534 1395 7580
rect 1343 7531 1395 7534
rect 2532 10271 2584 10323
rect 2636 10271 2639 10323
rect 2639 10271 2685 10323
rect 2685 10271 2688 10323
rect 2532 10167 2584 10219
rect 2636 10167 2639 10219
rect 2639 10167 2685 10219
rect 2685 10167 2688 10219
rect 2636 9405 2639 9457
rect 2639 9405 2685 9457
rect 2685 9405 2688 9457
rect 2636 9301 2639 9353
rect 2639 9301 2685 9353
rect 2685 9301 2688 9353
rect 2636 8075 2639 8127
rect 2639 8075 2685 8127
rect 2685 8075 2688 8127
rect 2636 7971 2639 8023
rect 2639 7971 2685 8023
rect 2685 7971 2688 8023
rect 3962 14219 4014 14222
rect 3962 14173 3965 14219
rect 3965 14173 4011 14219
rect 4011 14173 4014 14219
rect 3962 14170 4014 14173
rect 4042 13925 4045 13977
rect 4045 13925 4091 13977
rect 4091 13925 4094 13977
rect 4042 13821 4045 13873
rect 4045 13821 4091 13873
rect 4091 13821 4094 13873
rect 3882 13429 3885 13481
rect 3885 13429 3931 13481
rect 3931 13429 3934 13481
rect 3882 13325 3885 13377
rect 3885 13325 3931 13377
rect 3931 13325 3934 13377
rect 4202 13925 4205 13977
rect 4205 13925 4251 13977
rect 4251 13925 4254 13977
rect 4202 13821 4205 13873
rect 4205 13821 4251 13873
rect 4251 13821 4254 13873
rect 4522 13429 4525 13481
rect 4525 13429 4571 13481
rect 4571 13429 4574 13481
rect 4522 13325 4525 13377
rect 4525 13325 4571 13377
rect 4571 13325 4574 13377
rect 4843 13925 4845 13977
rect 4845 13925 4891 13977
rect 4891 13925 4895 13977
rect 4843 13821 4845 13873
rect 4845 13821 4891 13873
rect 4891 13821 4895 13873
rect 5162 13429 5165 13481
rect 5165 13429 5211 13481
rect 5211 13429 5214 13481
rect 5162 13325 5165 13377
rect 5165 13325 5211 13377
rect 5211 13325 5214 13377
rect 3962 13146 4014 13198
rect 3962 13091 4014 13094
rect 3962 13045 3965 13091
rect 3965 13045 4011 13091
rect 4011 13045 4014 13091
rect 3962 13042 4014 13045
rect 4042 12795 4045 12847
rect 4045 12795 4091 12847
rect 4091 12795 4094 12847
rect 4042 12691 4045 12743
rect 4045 12691 4091 12743
rect 4091 12691 4094 12743
rect 3882 12403 3885 12455
rect 3885 12403 3931 12455
rect 3931 12403 3934 12455
rect 3882 12299 3885 12351
rect 3885 12299 3931 12351
rect 3931 12299 3934 12351
rect 4202 12795 4205 12847
rect 4205 12795 4251 12847
rect 4251 12795 4254 12847
rect 4202 12691 4205 12743
rect 4205 12691 4251 12743
rect 4251 12691 4254 12743
rect 4522 12403 4525 12455
rect 4525 12403 4571 12455
rect 4571 12403 4574 12455
rect 4522 12299 4525 12351
rect 4525 12299 4571 12351
rect 4571 12299 4574 12351
rect 4843 12795 4845 12847
rect 4845 12795 4891 12847
rect 4891 12795 4895 12847
rect 4843 12691 4845 12743
rect 4845 12691 4891 12743
rect 4891 12691 4895 12743
rect 5162 12403 5165 12455
rect 5165 12403 5211 12455
rect 5211 12403 5214 12455
rect 5162 12299 5165 12351
rect 5165 12299 5211 12351
rect 5211 12299 5214 12351
rect 3962 12016 4014 12068
rect 3962 11963 4014 11964
rect 3962 11917 3965 11963
rect 3965 11917 4011 11963
rect 4011 11917 4014 11963
rect 3962 11912 4014 11917
rect 3882 11169 3885 11221
rect 3885 11169 3931 11221
rect 3931 11169 3934 11221
rect 3882 11065 3885 11117
rect 3885 11065 3931 11117
rect 3931 11065 3934 11117
rect 4202 11665 4205 11717
rect 4205 11665 4251 11717
rect 4251 11665 4254 11717
rect 4202 11561 4205 11613
rect 4205 11561 4251 11613
rect 4251 11561 4254 11613
rect 4042 10271 4045 10323
rect 4045 10271 4091 10323
rect 4091 10271 4094 10323
rect 4042 10167 4045 10219
rect 4045 10167 4091 10219
rect 4091 10167 4094 10219
rect 4522 11169 4525 11221
rect 4525 11169 4571 11221
rect 4571 11169 4574 11221
rect 4522 11065 4525 11117
rect 4525 11065 4571 11117
rect 4571 11065 4574 11117
rect 4843 11665 4845 11717
rect 4845 11665 4891 11717
rect 4891 11665 4895 11717
rect 4843 11561 4845 11613
rect 4845 11561 4891 11613
rect 4891 11561 4895 11613
rect 5162 11169 5165 11221
rect 5165 11169 5211 11221
rect 5211 11169 5214 11221
rect 5162 11065 5165 11117
rect 5165 11065 5211 11117
rect 5211 11065 5214 11117
rect 3962 9758 4014 9810
rect 3962 9703 4014 9706
rect 3962 9657 3965 9703
rect 3965 9657 4011 9703
rect 4011 9657 4014 9703
rect 3962 9654 4014 9657
rect 4042 9405 4045 9457
rect 4045 9405 4091 9457
rect 4091 9405 4094 9457
rect 4042 9301 4045 9353
rect 4045 9301 4091 9353
rect 4091 9301 4094 9353
rect 3882 8909 3885 8961
rect 3885 8909 3931 8961
rect 3931 8909 3934 8961
rect 3882 8805 3885 8857
rect 3885 8805 3931 8857
rect 3931 8805 3934 8857
rect 4202 9405 4205 9457
rect 4205 9405 4251 9457
rect 4251 9405 4254 9457
rect 4202 9301 4205 9353
rect 4205 9301 4251 9353
rect 4251 9301 4254 9353
rect 4522 8909 4525 8961
rect 4525 8909 4571 8961
rect 4571 8909 4574 8961
rect 4522 8805 4525 8857
rect 4525 8805 4571 8857
rect 4571 8805 4574 8857
rect 4843 9405 4845 9457
rect 4845 9405 4891 9457
rect 4891 9405 4895 9457
rect 4843 9301 4845 9353
rect 4845 9301 4891 9353
rect 4891 9301 4895 9353
rect 5162 8909 5165 8961
rect 5165 8909 5211 8961
rect 5211 8909 5214 8961
rect 5162 8805 5165 8857
rect 5165 8805 5211 8857
rect 5211 8805 5214 8857
rect 3962 8628 4014 8680
rect 3962 8573 4014 8576
rect 3962 8527 3965 8573
rect 3965 8527 4011 8573
rect 4011 8527 4014 8573
rect 3962 8524 4014 8527
rect 4202 8275 4205 8327
rect 4205 8275 4251 8327
rect 4251 8275 4254 8327
rect 4202 8171 4205 8223
rect 4205 8171 4251 8223
rect 4251 8171 4254 8223
rect 4042 8075 4045 8127
rect 4045 8075 4091 8127
rect 4091 8075 4094 8127
rect 4042 7971 4045 8023
rect 4045 7971 4091 8023
rect 4091 7971 4094 8023
rect 3882 7779 3885 7831
rect 3885 7779 3931 7831
rect 3931 7779 3934 7831
rect 3882 7675 3885 7727
rect 3885 7675 3931 7727
rect 3931 7675 3934 7727
rect 4522 7779 4525 7831
rect 4525 7779 4571 7831
rect 4571 7779 4574 7831
rect 4522 7675 4525 7727
rect 4525 7675 4571 7727
rect 4571 7675 4574 7727
rect 4843 8275 4845 8327
rect 4845 8275 4891 8327
rect 4891 8275 4895 8327
rect 4843 8171 4845 8223
rect 4845 8171 4891 8223
rect 4891 8171 4895 8223
rect 5162 7779 5165 7831
rect 5165 7779 5211 7831
rect 5211 7779 5214 7831
rect 5162 7675 5165 7727
rect 5165 7675 5211 7727
rect 5211 7675 5214 7727
rect 4122 7489 4174 7492
rect 4122 7443 4125 7489
rect 4125 7443 4171 7489
rect 4171 7443 4174 7489
rect 4122 7440 4174 7443
rect 5743 14220 5795 14272
rect 5847 14220 5899 14272
rect 5743 14116 5795 14168
rect 5847 14116 5899 14168
rect 6015 13925 6067 13977
rect 6119 13925 6171 13977
rect 6015 13821 6067 13873
rect 6119 13821 6171 13873
rect 6747 14263 6799 14272
rect 6747 14220 6750 14263
rect 6750 14220 6796 14263
rect 6796 14220 6799 14263
rect 6747 14116 6750 14168
rect 6750 14116 6796 14168
rect 6796 14116 6799 14168
rect 7067 13925 7070 13977
rect 7070 13925 7116 13977
rect 7116 13925 7119 13977
rect 7067 13821 7070 13873
rect 7070 13821 7116 13873
rect 7116 13821 7119 13873
rect 7387 14263 7439 14272
rect 7387 14220 7390 14263
rect 7390 14220 7436 14263
rect 7436 14220 7439 14263
rect 7387 14116 7390 14168
rect 7390 14116 7436 14168
rect 7436 14116 7439 14168
rect 6747 12946 6750 12998
rect 6750 12946 6796 12998
rect 6796 12946 6799 12998
rect 6747 12851 6750 12894
rect 6750 12851 6796 12894
rect 6796 12851 6799 12894
rect 6747 12842 6799 12851
rect 7707 13925 7710 13977
rect 7710 13925 7756 13977
rect 7756 13925 7759 13977
rect 7707 13821 7710 13873
rect 7710 13821 7756 13873
rect 7756 13821 7759 13873
rect 7067 13325 7070 13377
rect 7070 13325 7116 13377
rect 7116 13325 7119 13377
rect 7067 13221 7070 13273
rect 7070 13221 7116 13273
rect 7116 13221 7119 13273
rect 6747 12084 6750 12136
rect 6750 12084 6796 12136
rect 6796 12084 6799 12136
rect 6747 11989 6750 12032
rect 6750 11989 6796 12032
rect 6796 11989 6799 12032
rect 6747 11980 6799 11989
rect 8027 14263 8079 14272
rect 8027 14220 8030 14263
rect 8030 14220 8076 14263
rect 8076 14220 8079 14263
rect 8027 14116 8030 14168
rect 8030 14116 8076 14168
rect 8076 14116 8079 14168
rect 7387 12946 7390 12998
rect 7390 12946 7436 12998
rect 7436 12946 7439 12998
rect 7387 12851 7390 12894
rect 7390 12851 7436 12894
rect 7436 12851 7439 12894
rect 7387 12842 7439 12851
rect 7707 13325 7710 13377
rect 7710 13325 7756 13377
rect 7756 13325 7759 13377
rect 7707 13221 7710 13273
rect 7710 13221 7756 13273
rect 7756 13221 7759 13273
rect 7067 12403 7070 12455
rect 7070 12403 7116 12455
rect 7116 12403 7119 12455
rect 7067 12299 7070 12351
rect 7070 12299 7116 12351
rect 7116 12299 7119 12351
rect 6747 11561 6750 11613
rect 6750 11561 6796 11613
rect 6796 11561 6799 11613
rect 6747 11457 6750 11509
rect 6750 11457 6796 11509
rect 6796 11457 6799 11509
rect 7387 12084 7390 12136
rect 7390 12084 7436 12136
rect 7436 12084 7439 12136
rect 7387 11989 7390 12032
rect 7390 11989 7436 12032
rect 7436 11989 7439 12032
rect 7387 11980 7439 11989
rect 8027 12946 8030 12998
rect 8030 12946 8076 12998
rect 8076 12946 8079 12998
rect 8027 12851 8030 12894
rect 8030 12851 8076 12894
rect 8076 12851 8079 12894
rect 8027 12842 8079 12851
rect 7707 12403 7710 12455
rect 7710 12403 7756 12455
rect 7756 12403 7759 12455
rect 7707 12299 7710 12351
rect 7710 12299 7756 12351
rect 7756 12299 7759 12351
rect 7067 11273 7070 11325
rect 7070 11273 7116 11325
rect 7116 11273 7119 11325
rect 7067 11169 7070 11221
rect 7070 11169 7116 11221
rect 7116 11169 7119 11221
rect 7387 11561 7390 11613
rect 7390 11561 7436 11613
rect 7436 11561 7439 11613
rect 7387 11457 7390 11509
rect 7390 11457 7436 11509
rect 7436 11457 7439 11509
rect 6747 9509 6750 9561
rect 6750 9509 6796 9561
rect 6796 9509 6799 9561
rect 6747 9405 6750 9457
rect 6750 9405 6796 9457
rect 6796 9405 6799 9457
rect 7067 9953 7119 9962
rect 7067 9910 7070 9953
rect 7070 9910 7116 9953
rect 7116 9910 7119 9953
rect 7067 9806 7070 9858
rect 7070 9806 7116 9858
rect 7116 9806 7119 9858
rect 8027 12084 8030 12136
rect 8030 12084 8076 12136
rect 8076 12084 8079 12136
rect 8027 11989 8030 12032
rect 8030 11989 8076 12032
rect 8076 11989 8079 12032
rect 8027 11980 8079 11989
rect 7707 11273 7710 11325
rect 7710 11273 7756 11325
rect 7756 11273 7759 11325
rect 7707 11169 7710 11221
rect 7710 11169 7756 11221
rect 7756 11169 7759 11221
rect 6747 8909 6750 8961
rect 6750 8909 6796 8961
rect 6796 8909 6799 8961
rect 6747 8805 6750 8857
rect 6750 8805 6796 8857
rect 6796 8805 6799 8857
rect 8027 11561 8030 11613
rect 8030 11561 8076 11613
rect 8076 11561 8079 11613
rect 8027 11457 8030 11509
rect 8030 11457 8076 11509
rect 8076 11457 8079 11509
rect 7387 9509 7390 9561
rect 7390 9509 7436 9561
rect 7436 9509 7439 9561
rect 7387 9405 7390 9457
rect 7390 9405 7436 9457
rect 7436 9405 7439 9457
rect 7707 9953 7759 9962
rect 7707 9910 7710 9953
rect 7710 9910 7756 9953
rect 7756 9910 7759 9953
rect 7707 9806 7710 9858
rect 7710 9806 7756 9858
rect 7756 9806 7759 9858
rect 7067 8636 7070 8688
rect 7070 8636 7116 8688
rect 7116 8636 7119 8688
rect 7067 8541 7070 8584
rect 7070 8541 7116 8584
rect 7116 8541 7119 8584
rect 7067 8532 7119 8541
rect 7387 8909 7390 8961
rect 7390 8909 7436 8961
rect 7436 8909 7439 8961
rect 7387 8805 7390 8857
rect 7390 8805 7436 8857
rect 7436 8805 7439 8857
rect 6747 7779 6750 7831
rect 6750 7779 6796 7831
rect 6796 7779 6799 7831
rect 6747 7679 6750 7727
rect 6750 7679 6796 7727
rect 6796 7679 6799 7727
rect 6747 7675 6799 7679
rect 7067 8171 7070 8223
rect 7070 8171 7116 8223
rect 7116 8171 7119 8223
rect 7067 8067 7070 8119
rect 7070 8067 7116 8119
rect 7116 8067 7119 8119
rect 8027 9509 8030 9561
rect 8030 9509 8076 9561
rect 8076 9509 8079 9561
rect 8027 9405 8030 9457
rect 8030 9405 8076 9457
rect 8076 9405 8079 9457
rect 7707 8636 7710 8688
rect 7710 8636 7756 8688
rect 7756 8636 7759 8688
rect 7707 8541 7710 8584
rect 7710 8541 7756 8584
rect 7756 8541 7759 8584
rect 7707 8532 7759 8541
rect 8027 8909 8030 8961
rect 8030 8909 8076 8961
rect 8076 8909 8079 8961
rect 8027 8805 8030 8857
rect 8030 8805 8076 8857
rect 8076 8805 8079 8857
rect 7387 7779 7390 7831
rect 7390 7779 7436 7831
rect 7436 7779 7439 7831
rect 7387 7679 7390 7727
rect 7390 7679 7436 7727
rect 7436 7679 7439 7727
rect 7387 7675 7439 7679
rect 7707 8171 7710 8223
rect 7710 8171 7756 8223
rect 7756 8171 7759 8223
rect 7707 8067 7710 8119
rect 7710 8067 7756 8119
rect 7756 8067 7759 8119
rect 8001 8461 8053 8464
rect 8001 8415 8004 8461
rect 8004 8415 8050 8461
rect 8050 8415 8053 8461
rect 8001 8412 8053 8415
rect 8001 8357 8053 8360
rect 8001 8311 8004 8357
rect 8004 8311 8050 8357
rect 8050 8311 8053 8357
rect 8001 8308 8053 8311
rect 8027 7779 8030 7831
rect 8030 7779 8076 7831
rect 8076 7779 8079 7831
rect 8027 7679 8030 7727
rect 8030 7679 8076 7727
rect 8076 7679 8079 7727
rect 8027 7675 8079 7679
rect 11383 11321 11435 11373
rect 11487 11321 11539 11373
rect 11383 11217 11435 11269
rect 11487 11217 11539 11269
rect 6879 7327 6931 7379
rect 6983 7327 7035 7379
rect 8982 10742 8985 10794
rect 8985 10742 9031 10794
rect 9031 10742 9034 10794
rect 8982 10638 8985 10690
rect 8985 10638 9031 10690
rect 9031 10638 9034 10690
rect 9430 10371 9433 10423
rect 9433 10371 9479 10423
rect 9479 10371 9482 10423
rect 9430 10267 9433 10319
rect 9433 10267 9479 10319
rect 9479 10267 9482 10319
rect 9878 10742 9881 10794
rect 9881 10742 9927 10794
rect 9927 10742 9930 10794
rect 9878 10638 9881 10690
rect 9881 10638 9927 10690
rect 9927 10638 9930 10690
rect 10326 10371 10329 10423
rect 10329 10371 10375 10423
rect 10375 10371 10378 10423
rect 10326 10267 10329 10319
rect 10329 10267 10375 10319
rect 10375 10267 10378 10319
rect 10774 10742 10777 10794
rect 10777 10742 10823 10794
rect 10823 10742 10826 10794
rect 10774 10638 10777 10690
rect 10777 10638 10823 10690
rect 10823 10638 10826 10690
rect 10614 10371 10617 10423
rect 10617 10371 10663 10423
rect 10663 10371 10666 10423
rect 10614 10267 10617 10319
rect 10617 10267 10663 10319
rect 10663 10267 10666 10319
rect 8982 8909 8985 8961
rect 8985 8909 9031 8961
rect 9031 8909 9034 8961
rect 8982 8805 8985 8857
rect 8985 8805 9031 8857
rect 9031 8805 9034 8857
rect 9430 9509 9433 9561
rect 9433 9509 9479 9561
rect 9479 9509 9482 9561
rect 9430 9405 9433 9457
rect 9433 9405 9479 9457
rect 9479 9405 9482 9457
rect 9878 8909 9881 8961
rect 9881 8909 9927 8961
rect 9927 8909 9930 8961
rect 9878 8805 9881 8857
rect 9881 8805 9927 8857
rect 9927 8805 9930 8857
rect 10326 9509 10329 9561
rect 10329 9509 10375 9561
rect 10375 9509 10378 9561
rect 10326 9405 10329 9457
rect 10329 9405 10375 9457
rect 10375 9405 10378 9457
rect 10614 9709 10617 9761
rect 10617 9709 10663 9761
rect 10663 9709 10666 9761
rect 10614 9605 10617 9657
rect 10617 9605 10663 9657
rect 10663 9605 10666 9657
rect 10486 8651 10489 8703
rect 10489 8651 10535 8703
rect 10535 8651 10538 8703
rect 10486 8547 10489 8599
rect 10489 8547 10535 8599
rect 10535 8547 10538 8599
rect 10774 8909 10777 8961
rect 10777 8909 10823 8961
rect 10823 8909 10826 8961
rect 10774 8805 10777 8857
rect 10777 8805 10823 8857
rect 10823 8805 10826 8857
rect 10734 8450 10786 8453
rect 10734 8404 10737 8450
rect 10737 8404 10783 8450
rect 10783 8404 10786 8450
rect 10734 8401 10786 8404
rect 10734 8346 10786 8349
rect 10734 8300 10737 8346
rect 10737 8300 10783 8346
rect 10783 8300 10786 8346
rect 10734 8297 10786 8300
rect 8982 7779 8985 7831
rect 8985 7779 9031 7831
rect 9031 7779 9034 7831
rect 8982 7675 8985 7727
rect 8985 7675 9031 7727
rect 9031 7675 9034 7727
rect 9430 8210 9482 8223
rect 9430 8171 9433 8210
rect 9433 8171 9479 8210
rect 9479 8171 9482 8210
rect 9430 8067 9433 8119
rect 9433 8067 9479 8119
rect 9479 8067 9482 8119
rect 9878 7779 9881 7831
rect 9881 7779 9927 7831
rect 9927 7779 9930 7831
rect 9878 7675 9881 7727
rect 9881 7675 9927 7727
rect 9927 7675 9930 7727
rect 10326 8210 10378 8223
rect 10326 8171 10329 8210
rect 10329 8171 10375 8210
rect 10375 8171 10378 8210
rect 10326 8067 10329 8119
rect 10329 8067 10375 8119
rect 10375 8067 10378 8119
rect 10486 8210 10538 8223
rect 10486 8171 10489 8210
rect 10489 8171 10535 8210
rect 10535 8171 10538 8210
rect 10486 8067 10489 8119
rect 10489 8067 10535 8119
rect 10535 8067 10538 8119
rect 10774 7779 10777 7831
rect 10777 7779 10823 7831
rect 10823 7779 10826 7831
rect 10774 7675 10777 7727
rect 10777 7675 10823 7727
rect 10823 7675 10826 7727
rect 11651 10901 11703 10953
rect 11755 10901 11807 10953
rect 11651 10797 11703 10849
rect 11755 10797 11807 10849
rect 9981 7327 10033 7379
rect 10085 7327 10137 7379
rect 6879 7223 6931 7275
rect 6983 7223 7035 7275
rect 9981 7223 10033 7275
rect 10085 7223 10137 7275
rect 12364 10901 12367 10953
rect 12367 10901 12413 10953
rect 12413 10901 12416 10953
rect 12364 10797 12367 10849
rect 12367 10797 12413 10849
rect 12413 10797 12416 10849
rect 12812 11364 12864 11373
rect 12812 11321 12815 11364
rect 12815 11321 12861 11364
rect 12861 11321 12864 11364
rect 12812 11217 12815 11269
rect 12815 11217 12861 11269
rect 12861 11217 12864 11269
rect 13260 10901 13263 10953
rect 13263 10901 13309 10953
rect 13309 10901 13312 10953
rect 13260 10797 13263 10849
rect 13263 10797 13309 10849
rect 13309 10797 13312 10849
rect 13708 11364 13760 11373
rect 13708 11321 13711 11364
rect 13711 11321 13757 11364
rect 13757 11321 13760 11364
rect 13708 11217 13711 11269
rect 13711 11217 13757 11269
rect 13757 11217 13760 11269
rect 13996 11364 14048 11373
rect 13996 11321 13999 11364
rect 13999 11321 14045 11364
rect 14045 11321 14048 11364
rect 13996 11217 13999 11269
rect 13999 11217 14045 11269
rect 14045 11217 14048 11269
rect 14156 10901 14159 10953
rect 14159 10901 14205 10953
rect 14205 10901 14208 10953
rect 14156 10797 14159 10849
rect 14159 10797 14205 10849
rect 14205 10797 14208 10849
rect 12364 9221 12367 9273
rect 12367 9221 12413 9273
rect 12413 9221 12416 9273
rect 12364 9117 12367 9169
rect 12367 9117 12413 9169
rect 12413 9117 12416 9169
rect 12812 10267 12815 10319
rect 12815 10267 12861 10319
rect 12861 10267 12864 10319
rect 12812 10163 12815 10215
rect 12815 10163 12861 10215
rect 12861 10163 12864 10215
rect 13260 9221 13263 9273
rect 13263 9221 13309 9273
rect 13309 9221 13312 9273
rect 13260 9117 13263 9169
rect 13263 9117 13309 9169
rect 13309 9117 13312 9169
rect 13708 10267 13711 10319
rect 13711 10267 13757 10319
rect 13757 10267 13760 10319
rect 13708 10163 13711 10215
rect 13711 10163 13757 10215
rect 13757 10163 13760 10215
rect 13996 10241 13999 10293
rect 13999 10241 14045 10293
rect 14045 10241 14048 10293
rect 13996 10137 13999 10189
rect 13999 10137 14045 10189
rect 14045 10137 14048 10189
rect 13868 8821 13871 8873
rect 13871 8821 13917 8873
rect 13917 8821 13920 8873
rect 13868 8717 13871 8769
rect 13871 8717 13917 8769
rect 13917 8717 13920 8769
rect 14156 9221 14159 9273
rect 14159 9221 14205 9273
rect 14205 9221 14208 9273
rect 14156 9117 14159 9169
rect 14159 9117 14205 9169
rect 14205 9117 14208 9169
rect 12400 8560 12452 8563
rect 12400 8514 12403 8560
rect 12403 8514 12449 8560
rect 12449 8514 12452 8560
rect 12400 8511 12452 8514
rect 12400 8456 12452 8459
rect 12400 8410 12403 8456
rect 12403 8410 12449 8456
rect 12449 8410 12452 8456
rect 12400 8407 12452 8410
rect 12364 7771 12367 7823
rect 12367 7771 12413 7823
rect 12413 7771 12416 7823
rect 12364 7667 12367 7719
rect 12367 7667 12413 7719
rect 12413 7667 12416 7719
rect 12812 8171 12815 8223
rect 12815 8171 12861 8223
rect 12861 8171 12864 8223
rect 12812 8067 12815 8119
rect 12815 8067 12861 8119
rect 12861 8067 12864 8119
rect 13260 7771 13263 7823
rect 13263 7771 13309 7823
rect 13309 7771 13312 7823
rect 13260 7667 13263 7719
rect 13263 7667 13309 7719
rect 13309 7667 13312 7719
rect 13708 8171 13711 8223
rect 13711 8171 13757 8223
rect 13757 8171 13760 8223
rect 13708 8067 13711 8119
rect 13711 8067 13757 8119
rect 13757 8067 13760 8119
rect 13868 8171 13871 8223
rect 13871 8171 13917 8223
rect 13917 8171 13920 8223
rect 13868 8067 13871 8119
rect 13871 8067 13917 8119
rect 13917 8067 13920 8119
rect 14156 7771 14159 7823
rect 14159 7771 14205 7823
rect 14205 7771 14208 7823
rect 14156 7667 14159 7719
rect 14159 7667 14205 7719
rect 14205 7667 14208 7719
rect 15158 11364 15210 11373
rect 15158 11321 15161 11364
rect 15161 11321 15207 11364
rect 15207 11321 15210 11364
rect 15158 11217 15161 11269
rect 15161 11217 15207 11269
rect 15207 11217 15210 11269
rect 15478 10901 15481 10953
rect 15481 10901 15527 10953
rect 15527 10901 15530 10953
rect 15478 10797 15481 10849
rect 15481 10797 15527 10849
rect 15527 10797 15530 10849
rect 15798 11364 15850 11373
rect 15798 11321 15801 11364
rect 15801 11321 15847 11364
rect 15847 11321 15850 11364
rect 15798 11217 15801 11269
rect 15801 11217 15847 11269
rect 15847 11217 15850 11269
rect 15158 10241 15161 10293
rect 15161 10241 15207 10293
rect 15207 10241 15210 10293
rect 15158 10137 15161 10189
rect 15161 10137 15207 10189
rect 15207 10137 15210 10189
rect 16118 10901 16121 10953
rect 16121 10901 16167 10953
rect 16167 10901 16170 10953
rect 16118 10797 16121 10849
rect 16121 10797 16167 10849
rect 16167 10797 16170 10849
rect 16438 11364 16490 11373
rect 16438 11321 16441 11364
rect 16441 11321 16487 11364
rect 16487 11321 16490 11364
rect 16438 11217 16441 11269
rect 16441 11217 16487 11269
rect 16487 11217 16490 11269
rect 15798 10241 15801 10293
rect 15801 10241 15847 10293
rect 15847 10241 15850 10293
rect 15798 10137 15801 10189
rect 15801 10137 15847 10189
rect 15847 10137 15850 10189
rect 15478 8821 15481 8873
rect 15481 8821 15527 8873
rect 15527 8821 15530 8873
rect 15478 8717 15481 8769
rect 15481 8717 15527 8769
rect 15527 8717 15530 8769
rect 15186 8565 15238 8568
rect 15186 8519 15189 8565
rect 15189 8519 15235 8565
rect 15235 8519 15238 8565
rect 15186 8516 15238 8519
rect 15186 8461 15238 8464
rect 15186 8415 15189 8461
rect 15189 8415 15235 8461
rect 15235 8415 15238 8461
rect 15186 8412 15238 8415
rect 15158 7781 15161 7833
rect 15161 7781 15207 7833
rect 15207 7781 15210 7833
rect 15158 7677 15161 7729
rect 15161 7677 15207 7729
rect 15207 7677 15210 7729
rect 16438 10241 16441 10293
rect 16441 10241 16487 10293
rect 16487 10241 16490 10293
rect 16438 10137 16441 10189
rect 16441 10137 16487 10189
rect 16487 10137 16490 10189
rect 16118 8821 16121 8873
rect 16121 8821 16167 8873
rect 16167 8821 16170 8873
rect 16118 8717 16121 8769
rect 16121 8717 16167 8769
rect 16167 8717 16170 8769
rect 15478 8171 15481 8223
rect 15481 8171 15527 8223
rect 15527 8171 15530 8223
rect 15478 8067 15481 8119
rect 15481 8067 15527 8119
rect 15527 8067 15530 8119
rect 15798 7781 15801 7833
rect 15801 7781 15847 7833
rect 15847 7781 15850 7833
rect 15798 7677 15801 7729
rect 15801 7677 15847 7729
rect 15847 7677 15850 7729
rect 16118 8171 16121 8223
rect 16121 8171 16167 8223
rect 16167 8171 16170 8223
rect 16118 8067 16121 8119
rect 16121 8067 16167 8119
rect 16167 8067 16170 8119
rect 16438 7781 16441 7833
rect 16441 7781 16487 7833
rect 16487 7781 16490 7833
rect 16438 7677 16441 7729
rect 16441 7677 16487 7729
rect 16487 7677 16490 7729
rect 17377 11321 17429 11373
rect 17481 11321 17533 11373
rect 17377 11217 17429 11269
rect 17481 11217 17533 11269
rect 17115 10901 17167 10953
rect 17219 10901 17271 10953
rect 17115 10797 17167 10849
rect 17219 10797 17271 10849
rect 19077 13402 19129 13405
rect 20197 13402 20249 13405
rect 19077 13356 19080 13402
rect 19080 13356 19126 13402
rect 19126 13356 19129 13402
rect 20197 13356 20200 13402
rect 20200 13356 20246 13402
rect 20246 13356 20249 13402
rect 19077 13353 19129 13356
rect 20197 13353 20249 13356
rect 18997 12718 19000 12770
rect 19000 12718 19046 12770
rect 19046 12718 19049 12770
rect 18997 12614 19000 12666
rect 19000 12614 19046 12666
rect 19046 12614 19049 12666
rect 19317 13112 19320 13164
rect 19320 13112 19366 13164
rect 19366 13112 19369 13164
rect 19317 13008 19320 13060
rect 19320 13008 19366 13060
rect 19366 13008 19369 13060
rect 19157 12718 19160 12770
rect 19160 12718 19206 12770
rect 19206 12718 19209 12770
rect 19157 12614 19160 12666
rect 19160 12614 19206 12666
rect 19206 12614 19209 12666
rect 19477 12718 19480 12770
rect 19480 12718 19526 12770
rect 19526 12718 19529 12770
rect 19477 12614 19480 12666
rect 19480 12614 19526 12666
rect 19526 12614 19529 12666
rect 19637 12718 19640 12770
rect 19640 12718 19686 12770
rect 19686 12718 19689 12770
rect 19637 12614 19640 12666
rect 19640 12614 19686 12666
rect 19686 12614 19689 12666
rect 19957 13112 19960 13164
rect 19960 13112 20006 13164
rect 20006 13112 20009 13164
rect 19957 13008 19960 13060
rect 19960 13008 20006 13060
rect 20006 13008 20009 13060
rect 19797 12718 19800 12770
rect 19800 12718 19846 12770
rect 19846 12718 19849 12770
rect 19797 12614 19800 12666
rect 19800 12614 19846 12666
rect 19846 12614 19849 12666
rect 20117 12718 20120 12770
rect 20120 12718 20166 12770
rect 20166 12718 20169 12770
rect 20117 12614 20120 12666
rect 20120 12614 20166 12666
rect 20166 12614 20169 12666
rect 20277 12718 20280 12770
rect 20280 12718 20326 12770
rect 20326 12718 20329 12770
rect 20277 12614 20280 12666
rect 20280 12614 20326 12666
rect 20326 12614 20329 12666
rect 19077 12436 19129 12439
rect 19077 12390 19080 12436
rect 19080 12390 19126 12436
rect 19126 12390 19129 12436
rect 19077 12387 19129 12390
rect 18997 11782 19000 11834
rect 19000 11782 19046 11834
rect 19046 11782 19049 11834
rect 18997 11678 19000 11730
rect 19000 11678 19046 11730
rect 19046 11678 19049 11730
rect 19317 12176 19320 12228
rect 19320 12176 19366 12228
rect 19366 12176 19369 12228
rect 19317 12072 19320 12124
rect 19320 12072 19366 12124
rect 19366 12072 19369 12124
rect 19157 11782 19160 11834
rect 19160 11782 19206 11834
rect 19206 11782 19209 11834
rect 19157 11678 19160 11730
rect 19160 11678 19206 11730
rect 19206 11678 19209 11730
rect 19477 11782 19480 11834
rect 19480 11782 19526 11834
rect 19526 11782 19529 11834
rect 19477 11678 19480 11730
rect 19480 11678 19526 11730
rect 19526 11678 19529 11730
rect 19637 11782 19640 11834
rect 19640 11782 19686 11834
rect 19686 11782 19689 11834
rect 19637 11678 19640 11730
rect 19640 11678 19686 11730
rect 19686 11678 19689 11730
rect 19957 12176 19960 12228
rect 19960 12176 20006 12228
rect 20006 12176 20009 12228
rect 19957 12072 19960 12124
rect 19960 12072 20006 12124
rect 20006 12072 20009 12124
rect 19797 11782 19800 11834
rect 19800 11782 19846 11834
rect 19846 11782 19849 11834
rect 19797 11678 19800 11730
rect 19800 11678 19846 11730
rect 19846 11678 19849 11730
rect 20117 11782 20120 11834
rect 20120 11782 20166 11834
rect 20166 11782 20169 11834
rect 20117 11678 20120 11730
rect 20120 11678 20166 11730
rect 20166 11678 20169 11730
rect 20277 11782 20280 11834
rect 20280 11782 20326 11834
rect 20326 11782 20329 11834
rect 20277 11678 20280 11730
rect 20280 11678 20326 11730
rect 20326 11678 20329 11730
rect 19077 11500 19129 11503
rect 19077 11454 19080 11500
rect 19080 11454 19126 11500
rect 19126 11454 19129 11500
rect 19077 11451 19129 11454
rect 18997 10846 19000 10898
rect 19000 10846 19046 10898
rect 19046 10846 19049 10898
rect 18997 10742 19000 10794
rect 19000 10742 19046 10794
rect 19046 10742 19049 10794
rect 19317 11240 19320 11292
rect 19320 11240 19366 11292
rect 19366 11240 19369 11292
rect 19317 11136 19320 11188
rect 19320 11136 19366 11188
rect 19366 11136 19369 11188
rect 19157 10846 19160 10898
rect 19160 10846 19206 10898
rect 19206 10846 19209 10898
rect 19157 10742 19160 10794
rect 19160 10742 19206 10794
rect 19206 10742 19209 10794
rect 19477 10846 19480 10898
rect 19480 10846 19526 10898
rect 19526 10846 19529 10898
rect 19477 10742 19480 10794
rect 19480 10742 19526 10794
rect 19526 10742 19529 10794
rect 19637 10846 19640 10898
rect 19640 10846 19686 10898
rect 19686 10846 19689 10898
rect 19637 10742 19640 10794
rect 19640 10742 19686 10794
rect 19686 10742 19689 10794
rect 19957 11240 19960 11292
rect 19960 11240 20006 11292
rect 20006 11240 20009 11292
rect 19957 11136 19960 11188
rect 19960 11136 20006 11188
rect 20006 11136 20009 11188
rect 19797 10846 19800 10898
rect 19800 10846 19846 10898
rect 19846 10846 19849 10898
rect 19797 10742 19800 10794
rect 19800 10742 19846 10794
rect 19846 10742 19849 10794
rect 20117 10846 20120 10898
rect 20120 10846 20166 10898
rect 20166 10846 20169 10898
rect 20117 10742 20120 10794
rect 20120 10742 20166 10794
rect 20166 10742 20169 10794
rect 20277 10846 20280 10898
rect 20280 10846 20326 10898
rect 20326 10846 20329 10898
rect 20277 10742 20280 10794
rect 20280 10742 20326 10794
rect 20326 10742 20329 10794
rect 18997 9910 19000 9962
rect 19000 9910 19046 9962
rect 19046 9910 19049 9962
rect 18997 9806 19000 9858
rect 19000 9806 19046 9858
rect 19046 9806 19049 9858
rect 19317 10304 19320 10356
rect 19320 10304 19366 10356
rect 19366 10304 19369 10356
rect 19317 10200 19320 10252
rect 19320 10200 19366 10252
rect 19366 10200 19369 10252
rect 19637 9910 19640 9962
rect 19640 9910 19686 9962
rect 19686 9910 19689 9962
rect 19637 9806 19640 9858
rect 19640 9806 19686 9858
rect 19686 9806 19689 9858
rect 19957 10304 19960 10356
rect 19960 10304 20006 10356
rect 20006 10304 20009 10356
rect 19957 10200 19960 10252
rect 19960 10200 20006 10252
rect 20006 10200 20009 10252
rect 20277 9910 20280 9962
rect 20280 9910 20326 9962
rect 20326 9910 20329 9962
rect 20277 9806 20280 9858
rect 20280 9806 20326 9858
rect 20326 9806 20329 9858
rect 19077 9628 19129 9631
rect 19077 9582 19080 9628
rect 19080 9582 19126 9628
rect 19126 9582 19129 9628
rect 19077 9579 19129 9582
rect 18997 8974 19000 9026
rect 19000 8974 19046 9026
rect 19046 8974 19049 9026
rect 18997 8870 19000 8922
rect 19000 8870 19046 8922
rect 19046 8870 19049 8922
rect 19317 9368 19320 9420
rect 19320 9368 19366 9420
rect 19366 9368 19369 9420
rect 19317 9264 19320 9316
rect 19320 9264 19366 9316
rect 19366 9264 19369 9316
rect 19157 8974 19160 9026
rect 19160 8974 19206 9026
rect 19206 8974 19209 9026
rect 19157 8870 19160 8922
rect 19160 8870 19206 8922
rect 19206 8870 19209 8922
rect 19477 8974 19480 9026
rect 19480 8974 19526 9026
rect 19526 8974 19529 9026
rect 19477 8870 19480 8922
rect 19480 8870 19526 8922
rect 19526 8870 19529 8922
rect 19637 8974 19640 9026
rect 19640 8974 19686 9026
rect 19686 8974 19689 9026
rect 19637 8870 19640 8922
rect 19640 8870 19686 8922
rect 19686 8870 19689 8922
rect 19957 9368 19960 9420
rect 19960 9368 20006 9420
rect 20006 9368 20009 9420
rect 19957 9264 19960 9316
rect 19960 9264 20006 9316
rect 20006 9264 20009 9316
rect 19797 8974 19800 9026
rect 19800 8974 19846 9026
rect 19846 8974 19849 9026
rect 19797 8870 19800 8922
rect 19800 8870 19846 8922
rect 19846 8870 19849 8922
rect 20117 8974 20120 9026
rect 20120 8974 20166 9026
rect 20166 8974 20169 9026
rect 20117 8870 20120 8922
rect 20120 8870 20166 8922
rect 20166 8870 20169 8922
rect 20277 8974 20280 9026
rect 20280 8974 20326 9026
rect 20326 8974 20329 9026
rect 20277 8870 20280 8922
rect 20280 8870 20326 8922
rect 20326 8870 20329 8922
rect 19077 8692 19129 8695
rect 19077 8646 19080 8692
rect 19080 8646 19126 8692
rect 19126 8646 19129 8692
rect 19077 8643 19129 8646
rect 18997 8038 19000 8090
rect 19000 8038 19046 8090
rect 19046 8038 19049 8090
rect 18997 7934 19000 7986
rect 19000 7934 19046 7986
rect 19046 7934 19049 7986
rect 19317 8432 19320 8484
rect 19320 8432 19366 8484
rect 19366 8432 19369 8484
rect 19317 8328 19320 8380
rect 19320 8328 19366 8380
rect 19366 8328 19369 8380
rect 19157 8038 19160 8090
rect 19160 8038 19206 8090
rect 19206 8038 19209 8090
rect 19157 7934 19160 7986
rect 19160 7934 19206 7986
rect 19206 7934 19209 7986
rect 19477 8038 19480 8090
rect 19480 8038 19526 8090
rect 19526 8038 19529 8090
rect 19477 7934 19480 7986
rect 19480 7934 19526 7986
rect 19526 7934 19529 7986
rect 19637 8038 19640 8090
rect 19640 8038 19686 8090
rect 19686 8038 19689 8090
rect 19637 7934 19640 7986
rect 19640 7934 19686 7986
rect 19686 7934 19689 7986
rect 19957 8432 19960 8484
rect 19960 8432 20006 8484
rect 20006 8432 20009 8484
rect 19957 8328 19960 8380
rect 19960 8328 20006 8380
rect 20006 8328 20009 8380
rect 19797 8038 19800 8090
rect 19800 8038 19846 8090
rect 19846 8038 19849 8090
rect 19797 7934 19800 7986
rect 19800 7934 19846 7986
rect 19846 7934 19849 7986
rect 20117 8038 20120 8090
rect 20120 8038 20166 8090
rect 20166 8038 20169 8090
rect 20117 7934 20120 7986
rect 20120 7934 20166 7986
rect 20166 7934 20169 7986
rect 20277 8038 20280 8090
rect 20280 8038 20326 8090
rect 20326 8038 20329 8090
rect 20277 7934 20280 7986
rect 20280 7934 20326 7986
rect 20326 7934 20329 7986
rect 19237 7756 19289 7759
rect 19877 7756 19929 7759
rect 19237 7710 19240 7756
rect 19240 7710 19286 7756
rect 19286 7710 19289 7756
rect 19877 7710 19880 7756
rect 19880 7710 19926 7756
rect 19926 7710 19929 7756
rect 19237 7707 19289 7710
rect 19877 7707 19929 7710
rect 24229 13402 24281 13405
rect 25349 13402 25401 13405
rect 24229 13356 24232 13402
rect 24232 13356 24278 13402
rect 24278 13356 24281 13402
rect 25349 13356 25352 13402
rect 25352 13356 25398 13402
rect 25398 13356 25401 13402
rect 24229 13353 24281 13356
rect 25349 13353 25401 13356
rect 24149 12718 24152 12770
rect 24152 12718 24198 12770
rect 24198 12718 24201 12770
rect 24149 12614 24152 12666
rect 24152 12614 24198 12666
rect 24198 12614 24201 12666
rect 24469 13112 24472 13164
rect 24472 13112 24518 13164
rect 24518 13112 24521 13164
rect 24469 13008 24472 13060
rect 24472 13008 24518 13060
rect 24518 13008 24521 13060
rect 24309 12718 24312 12770
rect 24312 12718 24358 12770
rect 24358 12718 24361 12770
rect 24309 12614 24312 12666
rect 24312 12614 24358 12666
rect 24358 12614 24361 12666
rect 24629 12718 24632 12770
rect 24632 12718 24678 12770
rect 24678 12718 24681 12770
rect 24629 12614 24632 12666
rect 24632 12614 24678 12666
rect 24678 12614 24681 12666
rect 24789 12718 24792 12770
rect 24792 12718 24838 12770
rect 24838 12718 24841 12770
rect 24789 12614 24792 12666
rect 24792 12614 24838 12666
rect 24838 12614 24841 12666
rect 25109 13112 25112 13164
rect 25112 13112 25158 13164
rect 25158 13112 25161 13164
rect 25109 13008 25112 13060
rect 25112 13008 25158 13060
rect 25158 13008 25161 13060
rect 24949 12718 24952 12770
rect 24952 12718 24998 12770
rect 24998 12718 25001 12770
rect 24949 12614 24952 12666
rect 24952 12614 24998 12666
rect 24998 12614 25001 12666
rect 25269 12718 25272 12770
rect 25272 12718 25318 12770
rect 25318 12718 25321 12770
rect 25269 12614 25272 12666
rect 25272 12614 25318 12666
rect 25318 12614 25321 12666
rect 25429 12718 25432 12770
rect 25432 12718 25478 12770
rect 25478 12718 25481 12770
rect 25429 12614 25432 12666
rect 25432 12614 25478 12666
rect 25478 12614 25481 12666
rect 25349 12436 25401 12439
rect 25349 12390 25352 12436
rect 25352 12390 25398 12436
rect 25398 12390 25401 12436
rect 25349 12387 25401 12390
rect 24149 11782 24152 11834
rect 24152 11782 24198 11834
rect 24198 11782 24201 11834
rect 24149 11678 24152 11730
rect 24152 11678 24198 11730
rect 24198 11678 24201 11730
rect 24469 12176 24472 12228
rect 24472 12176 24518 12228
rect 24518 12176 24521 12228
rect 24469 12072 24472 12124
rect 24472 12072 24518 12124
rect 24518 12072 24521 12124
rect 24309 11782 24312 11834
rect 24312 11782 24358 11834
rect 24358 11782 24361 11834
rect 24309 11678 24312 11730
rect 24312 11678 24358 11730
rect 24358 11678 24361 11730
rect 24629 11782 24632 11834
rect 24632 11782 24678 11834
rect 24678 11782 24681 11834
rect 24629 11678 24632 11730
rect 24632 11678 24678 11730
rect 24678 11678 24681 11730
rect 24789 11782 24792 11834
rect 24792 11782 24838 11834
rect 24838 11782 24841 11834
rect 24789 11678 24792 11730
rect 24792 11678 24838 11730
rect 24838 11678 24841 11730
rect 25109 12176 25112 12228
rect 25112 12176 25158 12228
rect 25158 12176 25161 12228
rect 25109 12072 25112 12124
rect 25112 12072 25158 12124
rect 25158 12072 25161 12124
rect 24949 11782 24952 11834
rect 24952 11782 24998 11834
rect 24998 11782 25001 11834
rect 24949 11678 24952 11730
rect 24952 11678 24998 11730
rect 24998 11678 25001 11730
rect 25269 11782 25272 11834
rect 25272 11782 25318 11834
rect 25318 11782 25321 11834
rect 25269 11678 25272 11730
rect 25272 11678 25318 11730
rect 25318 11678 25321 11730
rect 25429 11782 25432 11834
rect 25432 11782 25478 11834
rect 25478 11782 25481 11834
rect 25429 11678 25432 11730
rect 25432 11678 25478 11730
rect 25478 11678 25481 11730
rect 25349 11500 25401 11503
rect 25349 11454 25352 11500
rect 25352 11454 25398 11500
rect 25398 11454 25401 11500
rect 25349 11451 25401 11454
rect 24149 10846 24152 10898
rect 24152 10846 24198 10898
rect 24198 10846 24201 10898
rect 24149 10742 24152 10794
rect 24152 10742 24198 10794
rect 24198 10742 24201 10794
rect 24469 11240 24472 11292
rect 24472 11240 24518 11292
rect 24518 11240 24521 11292
rect 24469 11136 24472 11188
rect 24472 11136 24518 11188
rect 24518 11136 24521 11188
rect 24309 10846 24312 10898
rect 24312 10846 24358 10898
rect 24358 10846 24361 10898
rect 24309 10742 24312 10794
rect 24312 10742 24358 10794
rect 24358 10742 24361 10794
rect 24629 10846 24632 10898
rect 24632 10846 24678 10898
rect 24678 10846 24681 10898
rect 24629 10742 24632 10794
rect 24632 10742 24678 10794
rect 24678 10742 24681 10794
rect 24789 10846 24792 10898
rect 24792 10846 24838 10898
rect 24838 10846 24841 10898
rect 24789 10742 24792 10794
rect 24792 10742 24838 10794
rect 24838 10742 24841 10794
rect 25109 11240 25112 11292
rect 25112 11240 25158 11292
rect 25158 11240 25161 11292
rect 25109 11136 25112 11188
rect 25112 11136 25158 11188
rect 25158 11136 25161 11188
rect 24949 10846 24952 10898
rect 24952 10846 24998 10898
rect 24998 10846 25001 10898
rect 24949 10742 24952 10794
rect 24952 10742 24998 10794
rect 24998 10742 25001 10794
rect 25269 10846 25272 10898
rect 25272 10846 25318 10898
rect 25318 10846 25321 10898
rect 25269 10742 25272 10794
rect 25272 10742 25318 10794
rect 25318 10742 25321 10794
rect 25429 10846 25432 10898
rect 25432 10846 25478 10898
rect 25478 10846 25481 10898
rect 25429 10742 25432 10794
rect 25432 10742 25478 10794
rect 25478 10742 25481 10794
rect 24149 9910 24152 9962
rect 24152 9910 24198 9962
rect 24198 9910 24201 9962
rect 24149 9806 24152 9858
rect 24152 9806 24198 9858
rect 24198 9806 24201 9858
rect 24469 10304 24472 10356
rect 24472 10304 24518 10356
rect 24518 10304 24521 10356
rect 24469 10200 24472 10252
rect 24472 10200 24518 10252
rect 24518 10200 24521 10252
rect 24789 9910 24792 9962
rect 24792 9910 24838 9962
rect 24838 9910 24841 9962
rect 24789 9806 24792 9858
rect 24792 9806 24838 9858
rect 24838 9806 24841 9858
rect 25109 10304 25112 10356
rect 25112 10304 25158 10356
rect 25158 10304 25161 10356
rect 25109 10200 25112 10252
rect 25112 10200 25158 10252
rect 25158 10200 25161 10252
rect 25429 9910 25432 9962
rect 25432 9910 25478 9962
rect 25478 9910 25481 9962
rect 25429 9806 25432 9858
rect 25432 9806 25478 9858
rect 25478 9806 25481 9858
rect 25349 9628 25401 9631
rect 25349 9582 25352 9628
rect 25352 9582 25398 9628
rect 25398 9582 25401 9628
rect 25349 9579 25401 9582
rect 24149 8974 24152 9026
rect 24152 8974 24198 9026
rect 24198 8974 24201 9026
rect 24149 8870 24152 8922
rect 24152 8870 24198 8922
rect 24198 8870 24201 8922
rect 24469 9368 24472 9420
rect 24472 9368 24518 9420
rect 24518 9368 24521 9420
rect 24469 9264 24472 9316
rect 24472 9264 24518 9316
rect 24518 9264 24521 9316
rect 24309 8974 24312 9026
rect 24312 8974 24358 9026
rect 24358 8974 24361 9026
rect 24309 8870 24312 8922
rect 24312 8870 24358 8922
rect 24358 8870 24361 8922
rect 24629 8974 24632 9026
rect 24632 8974 24678 9026
rect 24678 8974 24681 9026
rect 24629 8870 24632 8922
rect 24632 8870 24678 8922
rect 24678 8870 24681 8922
rect 24789 8974 24792 9026
rect 24792 8974 24838 9026
rect 24838 8974 24841 9026
rect 24789 8870 24792 8922
rect 24792 8870 24838 8922
rect 24838 8870 24841 8922
rect 25109 9368 25112 9420
rect 25112 9368 25158 9420
rect 25158 9368 25161 9420
rect 25109 9264 25112 9316
rect 25112 9264 25158 9316
rect 25158 9264 25161 9316
rect 24949 8974 24952 9026
rect 24952 8974 24998 9026
rect 24998 8974 25001 9026
rect 24949 8870 24952 8922
rect 24952 8870 24998 8922
rect 24998 8870 25001 8922
rect 25269 8974 25272 9026
rect 25272 8974 25318 9026
rect 25318 8974 25321 9026
rect 25269 8870 25272 8922
rect 25272 8870 25318 8922
rect 25318 8870 25321 8922
rect 25429 8974 25432 9026
rect 25432 8974 25478 9026
rect 25478 8974 25481 9026
rect 25429 8870 25432 8922
rect 25432 8870 25478 8922
rect 25478 8870 25481 8922
rect 25349 8692 25401 8695
rect 25349 8646 25352 8692
rect 25352 8646 25398 8692
rect 25398 8646 25401 8692
rect 25349 8643 25401 8646
rect 24149 8038 24152 8090
rect 24152 8038 24198 8090
rect 24198 8038 24201 8090
rect 24149 7934 24152 7986
rect 24152 7934 24198 7986
rect 24198 7934 24201 7986
rect 24469 8432 24472 8484
rect 24472 8432 24518 8484
rect 24518 8432 24521 8484
rect 24469 8328 24472 8380
rect 24472 8328 24518 8380
rect 24518 8328 24521 8380
rect 24309 8038 24312 8090
rect 24312 8038 24358 8090
rect 24358 8038 24361 8090
rect 24309 7934 24312 7986
rect 24312 7934 24358 7986
rect 24358 7934 24361 7986
rect 24629 8038 24632 8090
rect 24632 8038 24678 8090
rect 24678 8038 24681 8090
rect 24629 7934 24632 7986
rect 24632 7934 24678 7986
rect 24678 7934 24681 7986
rect 24789 8038 24792 8090
rect 24792 8038 24838 8090
rect 24838 8038 24841 8090
rect 24789 7934 24792 7986
rect 24792 7934 24838 7986
rect 24838 7934 24841 7986
rect 25109 8432 25112 8484
rect 25112 8432 25158 8484
rect 25158 8432 25161 8484
rect 25109 8328 25112 8380
rect 25112 8328 25158 8380
rect 25158 8328 25161 8380
rect 24949 8038 24952 8090
rect 24952 8038 24998 8090
rect 24998 8038 25001 8090
rect 24949 7934 24952 7986
rect 24952 7934 24998 7986
rect 24998 7934 25001 7986
rect 25269 8038 25272 8090
rect 25272 8038 25318 8090
rect 25318 8038 25321 8090
rect 25269 7934 25272 7986
rect 25272 7934 25318 7986
rect 25318 7934 25321 7986
rect 25429 8038 25432 8090
rect 25432 8038 25478 8090
rect 25478 8038 25481 8090
rect 25429 7934 25432 7986
rect 25432 7934 25478 7986
rect 25478 7934 25481 7986
rect 24549 7756 24601 7759
rect 25189 7756 25241 7759
rect 24549 7710 24552 7756
rect 24552 7710 24598 7756
rect 24598 7710 24601 7756
rect 25189 7710 25192 7756
rect 25192 7710 25238 7756
rect 25238 7710 25241 7756
rect 24549 7707 24601 7710
rect 25189 7707 25241 7710
rect 28198 13402 28250 13405
rect 28198 13356 28201 13402
rect 28201 13356 28247 13402
rect 28247 13356 28250 13402
rect 28198 13353 28250 13356
rect 28118 12718 28121 12770
rect 28121 12718 28167 12770
rect 28167 12718 28170 12770
rect 28118 12614 28121 12666
rect 28121 12614 28167 12666
rect 28167 12614 28170 12666
rect 28438 13112 28441 13164
rect 28441 13112 28487 13164
rect 28487 13112 28490 13164
rect 28438 13008 28441 13060
rect 28441 13008 28487 13060
rect 28487 13008 28490 13060
rect 28278 12718 28281 12770
rect 28281 12718 28327 12770
rect 28327 12718 28330 12770
rect 28278 12614 28281 12666
rect 28281 12614 28327 12666
rect 28327 12614 28330 12666
rect 28598 12718 28601 12770
rect 28601 12718 28647 12770
rect 28647 12718 28650 12770
rect 28598 12614 28601 12666
rect 28601 12614 28647 12666
rect 28647 12614 28650 12666
rect 28758 12718 28761 12770
rect 28761 12718 28807 12770
rect 28807 12718 28810 12770
rect 28758 12614 28761 12666
rect 28761 12614 28807 12666
rect 28807 12614 28810 12666
rect 29078 13112 29081 13164
rect 29081 13112 29127 13164
rect 29127 13112 29130 13164
rect 29078 13008 29081 13060
rect 29081 13008 29127 13060
rect 29127 13008 29130 13060
rect 28918 12718 28921 12770
rect 28921 12718 28967 12770
rect 28967 12718 28970 12770
rect 28918 12614 28921 12666
rect 28921 12614 28967 12666
rect 28967 12614 28970 12666
rect 29238 12718 29241 12770
rect 29241 12718 29287 12770
rect 29287 12718 29290 12770
rect 29238 12614 29241 12666
rect 29241 12614 29287 12666
rect 29287 12614 29290 12666
rect 29398 12718 29401 12770
rect 29401 12718 29447 12770
rect 29447 12718 29450 12770
rect 29398 12614 29401 12666
rect 29401 12614 29447 12666
rect 29447 12614 29450 12666
rect 28198 12436 28250 12439
rect 28198 12390 28201 12436
rect 28201 12390 28247 12436
rect 28247 12390 28250 12436
rect 28198 12387 28250 12390
rect 28118 11782 28121 11834
rect 28121 11782 28167 11834
rect 28167 11782 28170 11834
rect 28118 11678 28121 11730
rect 28121 11678 28167 11730
rect 28167 11678 28170 11730
rect 28438 12176 28441 12228
rect 28441 12176 28487 12228
rect 28487 12176 28490 12228
rect 28438 12072 28441 12124
rect 28441 12072 28487 12124
rect 28487 12072 28490 12124
rect 28278 11782 28281 11834
rect 28281 11782 28327 11834
rect 28327 11782 28330 11834
rect 28278 11678 28281 11730
rect 28281 11678 28327 11730
rect 28327 11678 28330 11730
rect 28598 11782 28601 11834
rect 28601 11782 28647 11834
rect 28647 11782 28650 11834
rect 28598 11678 28601 11730
rect 28601 11678 28647 11730
rect 28647 11678 28650 11730
rect 28758 11782 28761 11834
rect 28761 11782 28807 11834
rect 28807 11782 28810 11834
rect 28758 11678 28761 11730
rect 28761 11678 28807 11730
rect 28807 11678 28810 11730
rect 29078 12176 29081 12228
rect 29081 12176 29127 12228
rect 29127 12176 29130 12228
rect 29078 12072 29081 12124
rect 29081 12072 29127 12124
rect 29127 12072 29130 12124
rect 28918 11782 28921 11834
rect 28921 11782 28967 11834
rect 28967 11782 28970 11834
rect 28918 11678 28921 11730
rect 28921 11678 28967 11730
rect 28967 11678 28970 11730
rect 29238 11782 29241 11834
rect 29241 11782 29287 11834
rect 29287 11782 29290 11834
rect 29238 11678 29241 11730
rect 29241 11678 29287 11730
rect 29287 11678 29290 11730
rect 29398 11782 29401 11834
rect 29401 11782 29447 11834
rect 29447 11782 29450 11834
rect 29398 11678 29401 11730
rect 29401 11678 29447 11730
rect 29447 11678 29450 11730
rect 28198 11500 28250 11503
rect 28198 11454 28201 11500
rect 28201 11454 28247 11500
rect 28247 11454 28250 11500
rect 28198 11451 28250 11454
rect 28118 10846 28121 10898
rect 28121 10846 28167 10898
rect 28167 10846 28170 10898
rect 28118 10742 28121 10794
rect 28121 10742 28167 10794
rect 28167 10742 28170 10794
rect 28438 11240 28441 11292
rect 28441 11240 28487 11292
rect 28487 11240 28490 11292
rect 28438 11136 28441 11188
rect 28441 11136 28487 11188
rect 28487 11136 28490 11188
rect 28278 10846 28281 10898
rect 28281 10846 28327 10898
rect 28327 10846 28330 10898
rect 28278 10742 28281 10794
rect 28281 10742 28327 10794
rect 28327 10742 28330 10794
rect 28598 10846 28601 10898
rect 28601 10846 28647 10898
rect 28647 10846 28650 10898
rect 28598 10742 28601 10794
rect 28601 10742 28647 10794
rect 28647 10742 28650 10794
rect 28758 10846 28761 10898
rect 28761 10846 28807 10898
rect 28807 10846 28810 10898
rect 28758 10742 28761 10794
rect 28761 10742 28807 10794
rect 28807 10742 28810 10794
rect 29078 11240 29081 11292
rect 29081 11240 29127 11292
rect 29127 11240 29130 11292
rect 29078 11136 29081 11188
rect 29081 11136 29127 11188
rect 29127 11136 29130 11188
rect 28918 10846 28921 10898
rect 28921 10846 28967 10898
rect 28967 10846 28970 10898
rect 28918 10742 28921 10794
rect 28921 10742 28967 10794
rect 28967 10742 28970 10794
rect 29238 10846 29241 10898
rect 29241 10846 29287 10898
rect 29287 10846 29290 10898
rect 29238 10742 29241 10794
rect 29241 10742 29287 10794
rect 29287 10742 29290 10794
rect 29398 10846 29401 10898
rect 29401 10846 29447 10898
rect 29447 10846 29450 10898
rect 29398 10742 29401 10794
rect 29401 10742 29447 10794
rect 29447 10742 29450 10794
rect 28118 9910 28121 9962
rect 28121 9910 28167 9962
rect 28167 9910 28170 9962
rect 28118 9806 28121 9858
rect 28121 9806 28167 9858
rect 28167 9806 28170 9858
rect 28438 10304 28441 10356
rect 28441 10304 28487 10356
rect 28487 10304 28490 10356
rect 28438 10200 28441 10252
rect 28441 10200 28487 10252
rect 28487 10200 28490 10252
rect 28758 9910 28761 9962
rect 28761 9910 28807 9962
rect 28807 9910 28810 9962
rect 28758 9806 28761 9858
rect 28761 9806 28807 9858
rect 28807 9806 28810 9858
rect 29078 10304 29081 10356
rect 29081 10304 29127 10356
rect 29127 10304 29130 10356
rect 29078 10200 29081 10252
rect 29081 10200 29127 10252
rect 29127 10200 29130 10252
rect 29398 9910 29401 9962
rect 29401 9910 29447 9962
rect 29447 9910 29450 9962
rect 29398 9806 29401 9858
rect 29401 9806 29447 9858
rect 29447 9806 29450 9858
rect 28198 9628 28250 9631
rect 28198 9582 28201 9628
rect 28201 9582 28247 9628
rect 28247 9582 28250 9628
rect 28198 9579 28250 9582
rect 28118 8974 28121 9026
rect 28121 8974 28167 9026
rect 28167 8974 28170 9026
rect 28118 8870 28121 8922
rect 28121 8870 28167 8922
rect 28167 8870 28170 8922
rect 28438 9368 28441 9420
rect 28441 9368 28487 9420
rect 28487 9368 28490 9420
rect 28438 9264 28441 9316
rect 28441 9264 28487 9316
rect 28487 9264 28490 9316
rect 28278 8974 28281 9026
rect 28281 8974 28327 9026
rect 28327 8974 28330 9026
rect 28278 8870 28281 8922
rect 28281 8870 28327 8922
rect 28327 8870 28330 8922
rect 28598 8974 28601 9026
rect 28601 8974 28647 9026
rect 28647 8974 28650 9026
rect 28598 8870 28601 8922
rect 28601 8870 28647 8922
rect 28647 8870 28650 8922
rect 28758 8974 28761 9026
rect 28761 8974 28807 9026
rect 28807 8974 28810 9026
rect 28758 8870 28761 8922
rect 28761 8870 28807 8922
rect 28807 8870 28810 8922
rect 29078 9368 29081 9420
rect 29081 9368 29127 9420
rect 29127 9368 29130 9420
rect 29078 9264 29081 9316
rect 29081 9264 29127 9316
rect 29127 9264 29130 9316
rect 28918 8974 28921 9026
rect 28921 8974 28967 9026
rect 28967 8974 28970 9026
rect 28918 8870 28921 8922
rect 28921 8870 28967 8922
rect 28967 8870 28970 8922
rect 29238 8974 29241 9026
rect 29241 8974 29287 9026
rect 29287 8974 29290 9026
rect 29238 8870 29241 8922
rect 29241 8870 29287 8922
rect 29287 8870 29290 8922
rect 29398 8974 29401 9026
rect 29401 8974 29447 9026
rect 29447 8974 29450 9026
rect 29398 8870 29401 8922
rect 29401 8870 29447 8922
rect 29447 8870 29450 8922
rect 28198 8692 28250 8695
rect 28198 8646 28201 8692
rect 28201 8646 28247 8692
rect 28247 8646 28250 8692
rect 28198 8643 28250 8646
rect 28118 8038 28121 8090
rect 28121 8038 28167 8090
rect 28167 8038 28170 8090
rect 28118 7934 28121 7986
rect 28121 7934 28167 7986
rect 28167 7934 28170 7986
rect 28438 8432 28441 8484
rect 28441 8432 28487 8484
rect 28487 8432 28490 8484
rect 28438 8328 28441 8380
rect 28441 8328 28487 8380
rect 28487 8328 28490 8380
rect 28278 8038 28281 8090
rect 28281 8038 28327 8090
rect 28327 8038 28330 8090
rect 28278 7934 28281 7986
rect 28281 7934 28327 7986
rect 28327 7934 28330 7986
rect 28598 8038 28601 8090
rect 28601 8038 28647 8090
rect 28647 8038 28650 8090
rect 28598 7934 28601 7986
rect 28601 7934 28647 7986
rect 28647 7934 28650 7986
rect 28758 8038 28761 8090
rect 28761 8038 28807 8090
rect 28807 8038 28810 8090
rect 28758 7934 28761 7986
rect 28761 7934 28807 7986
rect 28807 7934 28810 7986
rect 29078 8432 29081 8484
rect 29081 8432 29127 8484
rect 29127 8432 29130 8484
rect 29078 8328 29081 8380
rect 29081 8328 29127 8380
rect 29127 8328 29130 8380
rect 28918 8038 28921 8090
rect 28921 8038 28967 8090
rect 28967 8038 28970 8090
rect 28918 7934 28921 7986
rect 28921 7934 28967 7986
rect 28967 7934 28970 7986
rect 29238 8038 29241 8090
rect 29241 8038 29287 8090
rect 29287 8038 29290 8090
rect 29238 7934 29241 7986
rect 29241 7934 29287 7986
rect 29287 7934 29290 7986
rect 29398 8038 29401 8090
rect 29401 8038 29447 8090
rect 29447 8038 29450 8090
rect 29398 7934 29401 7986
rect 29401 7934 29447 7986
rect 29447 7934 29450 7986
rect 28358 7756 28410 7759
rect 28358 7710 28361 7756
rect 28361 7710 28407 7756
rect 28407 7710 28410 7756
rect 28358 7707 28410 7710
rect 66926 12996 66978 13048
rect 67030 12996 67082 13048
rect 67134 12996 67186 13048
rect 66926 12892 66978 12944
rect 67030 12892 67082 12944
rect 67134 12892 67186 12944
rect 66926 12788 66978 12840
rect 67030 12788 67082 12840
rect 67134 12788 67186 12840
rect 33414 11218 33417 11270
rect 33417 11218 33463 11270
rect 33463 11218 33466 11270
rect 33414 11114 33417 11166
rect 33417 11114 33463 11166
rect 33463 11114 33466 11166
rect 33735 11612 33737 11664
rect 33737 11612 33783 11664
rect 33783 11612 33787 11664
rect 33735 11508 33737 11560
rect 33737 11508 33783 11560
rect 33783 11508 33787 11560
rect 34614 11809 34666 11812
rect 34774 11809 34826 11812
rect 34614 11763 34617 11809
rect 34617 11763 34663 11809
rect 34663 11763 34666 11809
rect 34614 11760 34666 11763
rect 34774 11763 34777 11809
rect 34777 11763 34823 11809
rect 34823 11763 34826 11809
rect 34774 11760 34826 11763
rect 34054 11218 34057 11270
rect 34057 11218 34103 11270
rect 34103 11218 34106 11270
rect 34054 11114 34057 11166
rect 34057 11114 34103 11166
rect 34103 11114 34106 11166
rect 34375 11612 34377 11664
rect 34377 11612 34423 11664
rect 34423 11612 34427 11664
rect 34375 11508 34377 11560
rect 34377 11508 34423 11560
rect 34423 11508 34427 11560
rect 35015 11612 35017 11664
rect 35017 11612 35063 11664
rect 35063 11612 35067 11664
rect 35015 11508 35017 11560
rect 35017 11508 35063 11560
rect 35063 11508 35067 11560
rect 35334 11218 35337 11270
rect 35337 11218 35383 11270
rect 35383 11218 35386 11270
rect 35334 11114 35337 11166
rect 35337 11114 35383 11166
rect 35383 11114 35386 11166
rect 35655 11612 35657 11664
rect 35657 11612 35703 11664
rect 35703 11612 35707 11664
rect 35655 11508 35657 11560
rect 35657 11508 35703 11560
rect 35703 11508 35707 11560
rect 33414 10158 33417 10210
rect 33417 10158 33463 10210
rect 33463 10158 33466 10210
rect 33414 10054 33417 10106
rect 33417 10054 33463 10106
rect 33463 10054 33466 10106
rect 33735 10552 33737 10604
rect 33737 10552 33783 10604
rect 33783 10552 33787 10604
rect 33735 10448 33737 10500
rect 33737 10448 33783 10500
rect 33783 10448 33787 10500
rect 34614 10749 34666 10752
rect 34774 10749 34826 10752
rect 34614 10703 34617 10749
rect 34617 10703 34663 10749
rect 34663 10703 34666 10749
rect 34614 10700 34666 10703
rect 34774 10703 34777 10749
rect 34777 10703 34823 10749
rect 34823 10703 34826 10749
rect 34774 10700 34826 10703
rect 34054 10158 34057 10210
rect 34057 10158 34103 10210
rect 34103 10158 34106 10210
rect 34054 10054 34057 10106
rect 34057 10054 34103 10106
rect 34103 10054 34106 10106
rect 34375 10552 34377 10604
rect 34377 10552 34423 10604
rect 34423 10552 34427 10604
rect 34375 10448 34377 10500
rect 34377 10448 34423 10500
rect 34423 10448 34427 10500
rect 35015 10552 35017 10604
rect 35017 10552 35063 10604
rect 35063 10552 35067 10604
rect 35015 10448 35017 10500
rect 35017 10448 35063 10500
rect 35063 10448 35067 10500
rect 35974 11218 35977 11270
rect 35977 11218 36023 11270
rect 36023 11218 36026 11270
rect 35974 11114 35977 11166
rect 35977 11114 36023 11166
rect 36023 11114 36026 11166
rect 35334 10158 35337 10210
rect 35337 10158 35383 10210
rect 35383 10158 35386 10210
rect 35334 10054 35337 10106
rect 35337 10054 35383 10106
rect 35383 10054 35386 10106
rect 35655 10552 35657 10604
rect 35657 10552 35703 10604
rect 35703 10552 35707 10604
rect 35655 10448 35657 10500
rect 35657 10448 35703 10500
rect 35703 10448 35707 10500
rect 33414 9098 33417 9150
rect 33417 9098 33463 9150
rect 33463 9098 33466 9150
rect 33414 8994 33417 9046
rect 33417 8994 33463 9046
rect 33463 8994 33466 9046
rect 33735 9492 33737 9544
rect 33737 9492 33783 9544
rect 33783 9492 33787 9544
rect 33735 9388 33737 9440
rect 33737 9388 33783 9440
rect 33783 9388 33787 9440
rect 34614 9689 34666 9692
rect 34774 9689 34826 9692
rect 34614 9643 34617 9689
rect 34617 9643 34663 9689
rect 34663 9643 34666 9689
rect 34614 9640 34666 9643
rect 34774 9643 34777 9689
rect 34777 9643 34823 9689
rect 34823 9643 34826 9689
rect 34774 9640 34826 9643
rect 34054 9098 34057 9150
rect 34057 9098 34103 9150
rect 34103 9098 34106 9150
rect 34054 8994 34057 9046
rect 34057 8994 34103 9046
rect 34103 8994 34106 9046
rect 34375 9492 34377 9544
rect 34377 9492 34423 9544
rect 34423 9492 34427 9544
rect 34375 9388 34377 9440
rect 34377 9388 34423 9440
rect 34423 9388 34427 9440
rect 35015 9492 35017 9544
rect 35017 9492 35063 9544
rect 35063 9492 35067 9544
rect 35015 9388 35017 9440
rect 35017 9388 35063 9440
rect 35063 9388 35067 9440
rect 35974 10158 35977 10210
rect 35977 10158 36023 10210
rect 36023 10158 36026 10210
rect 35974 10054 35977 10106
rect 35977 10054 36023 10106
rect 36023 10054 36026 10106
rect 35334 9098 35337 9150
rect 35337 9098 35383 9150
rect 35383 9098 35386 9150
rect 35334 8994 35337 9046
rect 35337 8994 35383 9046
rect 35383 8994 35386 9046
rect 35655 9492 35657 9544
rect 35657 9492 35703 9544
rect 35703 9492 35707 9544
rect 35655 9388 35657 9440
rect 35657 9388 35703 9440
rect 35703 9388 35707 9440
rect 33414 8038 33417 8090
rect 33417 8038 33463 8090
rect 33463 8038 33466 8090
rect 33414 7934 33417 7986
rect 33417 7934 33463 7986
rect 33463 7934 33466 7986
rect 33735 8432 33737 8484
rect 33737 8432 33783 8484
rect 33783 8432 33787 8484
rect 33735 8328 33737 8380
rect 33737 8328 33783 8380
rect 33783 8328 33787 8380
rect 34614 8629 34666 8632
rect 34774 8629 34826 8632
rect 34614 8583 34617 8629
rect 34617 8583 34663 8629
rect 34663 8583 34666 8629
rect 34614 8580 34666 8583
rect 34774 8583 34777 8629
rect 34777 8583 34823 8629
rect 34823 8583 34826 8629
rect 34774 8580 34826 8583
rect 34054 8038 34057 8090
rect 34057 8038 34103 8090
rect 34103 8038 34106 8090
rect 34054 7934 34057 7986
rect 34057 7934 34103 7986
rect 34103 7934 34106 7986
rect 34375 8432 34377 8484
rect 34377 8432 34423 8484
rect 34423 8432 34427 8484
rect 34375 8328 34377 8380
rect 34377 8328 34423 8380
rect 34423 8328 34427 8380
rect 35015 8432 35017 8484
rect 35017 8432 35063 8484
rect 35063 8432 35067 8484
rect 35015 8328 35017 8380
rect 35017 8328 35063 8380
rect 35063 8328 35067 8380
rect 35974 9098 35977 9150
rect 35977 9098 36023 9150
rect 36023 9098 36026 9150
rect 35974 8994 35977 9046
rect 35977 8994 36023 9046
rect 36023 8994 36026 9046
rect 35334 8038 35337 8090
rect 35337 8038 35383 8090
rect 35383 8038 35386 8090
rect 35334 7934 35337 7986
rect 35337 7934 35383 7986
rect 35383 7934 35386 7986
rect 35655 8432 35657 8484
rect 35657 8432 35703 8484
rect 35703 8432 35707 8484
rect 35655 8328 35657 8380
rect 35657 8328 35703 8380
rect 35703 8328 35707 8380
rect 35974 8038 35977 8090
rect 35977 8038 36023 8090
rect 36023 8038 36026 8090
rect 35974 7934 35977 7986
rect 35977 7934 36023 7986
rect 36023 7934 36026 7986
rect 37550 11218 37553 11270
rect 37553 11218 37599 11270
rect 37599 11218 37602 11270
rect 37550 11114 37553 11166
rect 37553 11114 37599 11166
rect 37599 11114 37602 11166
rect 37869 11612 37873 11664
rect 37873 11612 37919 11664
rect 37919 11612 37921 11664
rect 37869 11508 37873 11560
rect 37873 11508 37919 11560
rect 37919 11508 37921 11560
rect 38750 11809 38802 11812
rect 38910 11809 38962 11812
rect 38750 11763 38753 11809
rect 38753 11763 38799 11809
rect 38799 11763 38802 11809
rect 38750 11760 38802 11763
rect 38910 11763 38913 11809
rect 38913 11763 38959 11809
rect 38959 11763 38962 11809
rect 38910 11760 38962 11763
rect 38190 11218 38193 11270
rect 38193 11218 38239 11270
rect 38239 11218 38242 11270
rect 38190 11114 38193 11166
rect 38193 11114 38239 11166
rect 38239 11114 38242 11166
rect 38509 11612 38513 11664
rect 38513 11612 38559 11664
rect 38559 11612 38561 11664
rect 38509 11508 38513 11560
rect 38513 11508 38559 11560
rect 38559 11508 38561 11560
rect 37550 10158 37553 10210
rect 37553 10158 37599 10210
rect 37599 10158 37602 10210
rect 37550 10054 37553 10106
rect 37553 10054 37599 10106
rect 37599 10054 37602 10106
rect 37869 10552 37873 10604
rect 37873 10552 37919 10604
rect 37919 10552 37921 10604
rect 37869 10448 37873 10500
rect 37873 10448 37919 10500
rect 37919 10448 37921 10500
rect 39149 11612 39153 11664
rect 39153 11612 39199 11664
rect 39199 11612 39201 11664
rect 39149 11508 39153 11560
rect 39153 11508 39199 11560
rect 39199 11508 39201 11560
rect 39470 11218 39473 11270
rect 39473 11218 39519 11270
rect 39519 11218 39522 11270
rect 39470 11114 39473 11166
rect 39473 11114 39519 11166
rect 39519 11114 39522 11166
rect 39789 11612 39793 11664
rect 39793 11612 39839 11664
rect 39839 11612 39841 11664
rect 39789 11508 39793 11560
rect 39793 11508 39839 11560
rect 39839 11508 39841 11560
rect 38750 10749 38802 10752
rect 38910 10749 38962 10752
rect 38750 10703 38753 10749
rect 38753 10703 38799 10749
rect 38799 10703 38802 10749
rect 38750 10700 38802 10703
rect 38910 10703 38913 10749
rect 38913 10703 38959 10749
rect 38959 10703 38962 10749
rect 38910 10700 38962 10703
rect 38190 10158 38193 10210
rect 38193 10158 38239 10210
rect 38239 10158 38242 10210
rect 38190 10054 38193 10106
rect 38193 10054 38239 10106
rect 38239 10054 38242 10106
rect 38509 10552 38513 10604
rect 38513 10552 38559 10604
rect 38559 10552 38561 10604
rect 38509 10448 38513 10500
rect 38513 10448 38559 10500
rect 38559 10448 38561 10500
rect 37550 9098 37553 9150
rect 37553 9098 37599 9150
rect 37599 9098 37602 9150
rect 37550 8994 37553 9046
rect 37553 8994 37599 9046
rect 37599 8994 37602 9046
rect 37869 9492 37873 9544
rect 37873 9492 37919 9544
rect 37919 9492 37921 9544
rect 37869 9388 37873 9440
rect 37873 9388 37919 9440
rect 37919 9388 37921 9440
rect 39149 10552 39153 10604
rect 39153 10552 39199 10604
rect 39199 10552 39201 10604
rect 39149 10448 39153 10500
rect 39153 10448 39199 10500
rect 39199 10448 39201 10500
rect 40110 11218 40113 11270
rect 40113 11218 40159 11270
rect 40159 11218 40162 11270
rect 40110 11114 40113 11166
rect 40113 11114 40159 11166
rect 40159 11114 40162 11166
rect 39470 10158 39473 10210
rect 39473 10158 39519 10210
rect 39519 10158 39522 10210
rect 39470 10054 39473 10106
rect 39473 10054 39519 10106
rect 39519 10054 39522 10106
rect 39789 10552 39793 10604
rect 39793 10552 39839 10604
rect 39839 10552 39841 10604
rect 39789 10448 39793 10500
rect 39793 10448 39839 10500
rect 39839 10448 39841 10500
rect 38750 9689 38802 9692
rect 38910 9689 38962 9692
rect 38750 9643 38753 9689
rect 38753 9643 38799 9689
rect 38799 9643 38802 9689
rect 38750 9640 38802 9643
rect 38910 9643 38913 9689
rect 38913 9643 38959 9689
rect 38959 9643 38962 9689
rect 38910 9640 38962 9643
rect 38190 9098 38193 9150
rect 38193 9098 38239 9150
rect 38239 9098 38242 9150
rect 38190 8994 38193 9046
rect 38193 8994 38239 9046
rect 38239 8994 38242 9046
rect 38509 9492 38513 9544
rect 38513 9492 38559 9544
rect 38559 9492 38561 9544
rect 38509 9388 38513 9440
rect 38513 9388 38559 9440
rect 38559 9388 38561 9440
rect 37550 8038 37553 8090
rect 37553 8038 37599 8090
rect 37599 8038 37602 8090
rect 37550 7934 37553 7986
rect 37553 7934 37599 7986
rect 37599 7934 37602 7986
rect 37869 8432 37873 8484
rect 37873 8432 37919 8484
rect 37919 8432 37921 8484
rect 37869 8328 37873 8380
rect 37873 8328 37919 8380
rect 37919 8328 37921 8380
rect 39149 9492 39153 9544
rect 39153 9492 39199 9544
rect 39199 9492 39201 9544
rect 39149 9388 39153 9440
rect 39153 9388 39199 9440
rect 39199 9388 39201 9440
rect 40110 10158 40113 10210
rect 40113 10158 40159 10210
rect 40159 10158 40162 10210
rect 40110 10054 40113 10106
rect 40113 10054 40159 10106
rect 40159 10054 40162 10106
rect 39470 9098 39473 9150
rect 39473 9098 39519 9150
rect 39519 9098 39522 9150
rect 39470 8994 39473 9046
rect 39473 8994 39519 9046
rect 39519 8994 39522 9046
rect 39789 9492 39793 9544
rect 39793 9492 39839 9544
rect 39839 9492 39841 9544
rect 39789 9388 39793 9440
rect 39793 9388 39839 9440
rect 39839 9388 39841 9440
rect 38750 8629 38802 8632
rect 38910 8629 38962 8632
rect 38750 8583 38753 8629
rect 38753 8583 38799 8629
rect 38799 8583 38802 8629
rect 38750 8580 38802 8583
rect 38910 8583 38913 8629
rect 38913 8583 38959 8629
rect 38959 8583 38962 8629
rect 38910 8580 38962 8583
rect 38190 8038 38193 8090
rect 38193 8038 38239 8090
rect 38239 8038 38242 8090
rect 38190 7934 38193 7986
rect 38193 7934 38239 7986
rect 38239 7934 38242 7986
rect 38509 8432 38513 8484
rect 38513 8432 38559 8484
rect 38559 8432 38561 8484
rect 38509 8328 38513 8380
rect 38513 8328 38559 8380
rect 38559 8328 38561 8380
rect 39149 8432 39153 8484
rect 39153 8432 39199 8484
rect 39199 8432 39201 8484
rect 39149 8328 39153 8380
rect 39153 8328 39199 8380
rect 39199 8328 39201 8380
rect 40110 9098 40113 9150
rect 40113 9098 40159 9150
rect 40159 9098 40162 9150
rect 40110 8994 40113 9046
rect 40113 8994 40159 9046
rect 40159 8994 40162 9046
rect 39470 8038 39473 8090
rect 39473 8038 39519 8090
rect 39519 8038 39522 8090
rect 39470 7934 39473 7986
rect 39473 7934 39519 7986
rect 39519 7934 39522 7986
rect 39789 8432 39793 8484
rect 39793 8432 39839 8484
rect 39839 8432 39841 8484
rect 39789 8328 39793 8380
rect 39793 8328 39839 8380
rect 39839 8328 39841 8380
rect 40110 8038 40113 8090
rect 40113 8038 40159 8090
rect 40159 8038 40162 8090
rect 40110 7934 40113 7986
rect 40113 7934 40159 7986
rect 40159 7934 40162 7986
rect 43110 11218 43113 11270
rect 43113 11218 43159 11270
rect 43159 11218 43162 11270
rect 43110 11114 43113 11166
rect 43113 11114 43159 11166
rect 43159 11114 43162 11166
rect 43431 11612 43433 11664
rect 43433 11612 43479 11664
rect 43479 11612 43483 11664
rect 43431 11508 43433 11560
rect 43433 11508 43479 11560
rect 43479 11508 43483 11560
rect 44310 11809 44362 11812
rect 44470 11809 44522 11812
rect 44310 11763 44313 11809
rect 44313 11763 44359 11809
rect 44359 11763 44362 11809
rect 44310 11760 44362 11763
rect 44470 11763 44473 11809
rect 44473 11763 44519 11809
rect 44519 11763 44522 11809
rect 44470 11760 44522 11763
rect 43750 11218 43753 11270
rect 43753 11218 43799 11270
rect 43799 11218 43802 11270
rect 43750 11114 43753 11166
rect 43753 11114 43799 11166
rect 43799 11114 43802 11166
rect 44071 11612 44073 11664
rect 44073 11612 44119 11664
rect 44119 11612 44123 11664
rect 44071 11508 44073 11560
rect 44073 11508 44119 11560
rect 44119 11508 44123 11560
rect 44711 11612 44713 11664
rect 44713 11612 44759 11664
rect 44759 11612 44763 11664
rect 44711 11508 44713 11560
rect 44713 11508 44759 11560
rect 44759 11508 44763 11560
rect 45030 11218 45033 11270
rect 45033 11218 45079 11270
rect 45079 11218 45082 11270
rect 45030 11114 45033 11166
rect 45033 11114 45079 11166
rect 45079 11114 45082 11166
rect 45351 11612 45353 11664
rect 45353 11612 45399 11664
rect 45399 11612 45403 11664
rect 45351 11508 45353 11560
rect 45353 11508 45399 11560
rect 45399 11508 45403 11560
rect 43110 10158 43113 10210
rect 43113 10158 43159 10210
rect 43159 10158 43162 10210
rect 43110 10054 43113 10106
rect 43113 10054 43159 10106
rect 43159 10054 43162 10106
rect 43431 10552 43433 10604
rect 43433 10552 43479 10604
rect 43479 10552 43483 10604
rect 43431 10448 43433 10500
rect 43433 10448 43479 10500
rect 43479 10448 43483 10500
rect 44310 10749 44362 10752
rect 44470 10749 44522 10752
rect 44310 10703 44313 10749
rect 44313 10703 44359 10749
rect 44359 10703 44362 10749
rect 44310 10700 44362 10703
rect 44470 10703 44473 10749
rect 44473 10703 44519 10749
rect 44519 10703 44522 10749
rect 44470 10700 44522 10703
rect 43750 10158 43753 10210
rect 43753 10158 43799 10210
rect 43799 10158 43802 10210
rect 43750 10054 43753 10106
rect 43753 10054 43799 10106
rect 43799 10054 43802 10106
rect 44071 10552 44073 10604
rect 44073 10552 44119 10604
rect 44119 10552 44123 10604
rect 44071 10448 44073 10500
rect 44073 10448 44119 10500
rect 44119 10448 44123 10500
rect 44711 10552 44713 10604
rect 44713 10552 44759 10604
rect 44759 10552 44763 10604
rect 44711 10448 44713 10500
rect 44713 10448 44759 10500
rect 44759 10448 44763 10500
rect 45670 11218 45673 11270
rect 45673 11218 45719 11270
rect 45719 11218 45722 11270
rect 45670 11114 45673 11166
rect 45673 11114 45719 11166
rect 45719 11114 45722 11166
rect 45030 10158 45033 10210
rect 45033 10158 45079 10210
rect 45079 10158 45082 10210
rect 45030 10054 45033 10106
rect 45033 10054 45079 10106
rect 45079 10054 45082 10106
rect 45351 10552 45353 10604
rect 45353 10552 45399 10604
rect 45399 10552 45403 10604
rect 45351 10448 45353 10500
rect 45353 10448 45399 10500
rect 45399 10448 45403 10500
rect 43110 9098 43113 9150
rect 43113 9098 43159 9150
rect 43159 9098 43162 9150
rect 43110 8994 43113 9046
rect 43113 8994 43159 9046
rect 43159 8994 43162 9046
rect 43431 9492 43433 9544
rect 43433 9492 43479 9544
rect 43479 9492 43483 9544
rect 43431 9388 43433 9440
rect 43433 9388 43479 9440
rect 43479 9388 43483 9440
rect 44310 9689 44362 9692
rect 44470 9689 44522 9692
rect 44310 9643 44313 9689
rect 44313 9643 44359 9689
rect 44359 9643 44362 9689
rect 44310 9640 44362 9643
rect 44470 9643 44473 9689
rect 44473 9643 44519 9689
rect 44519 9643 44522 9689
rect 44470 9640 44522 9643
rect 43750 9098 43753 9150
rect 43753 9098 43799 9150
rect 43799 9098 43802 9150
rect 43750 8994 43753 9046
rect 43753 8994 43799 9046
rect 43799 8994 43802 9046
rect 44071 9492 44073 9544
rect 44073 9492 44119 9544
rect 44119 9492 44123 9544
rect 44071 9388 44073 9440
rect 44073 9388 44119 9440
rect 44119 9388 44123 9440
rect 44711 9492 44713 9544
rect 44713 9492 44759 9544
rect 44759 9492 44763 9544
rect 44711 9388 44713 9440
rect 44713 9388 44759 9440
rect 44759 9388 44763 9440
rect 45670 10158 45673 10210
rect 45673 10158 45719 10210
rect 45719 10158 45722 10210
rect 45670 10054 45673 10106
rect 45673 10054 45719 10106
rect 45719 10054 45722 10106
rect 45030 9098 45033 9150
rect 45033 9098 45079 9150
rect 45079 9098 45082 9150
rect 45030 8994 45033 9046
rect 45033 8994 45079 9046
rect 45079 8994 45082 9046
rect 45351 9492 45353 9544
rect 45353 9492 45399 9544
rect 45399 9492 45403 9544
rect 45351 9388 45353 9440
rect 45353 9388 45399 9440
rect 45399 9388 45403 9440
rect 43110 8038 43113 8090
rect 43113 8038 43159 8090
rect 43159 8038 43162 8090
rect 43110 7934 43113 7986
rect 43113 7934 43159 7986
rect 43159 7934 43162 7986
rect 43431 8432 43433 8484
rect 43433 8432 43479 8484
rect 43479 8432 43483 8484
rect 43431 8328 43433 8380
rect 43433 8328 43479 8380
rect 43479 8328 43483 8380
rect 44310 8629 44362 8632
rect 44470 8629 44522 8632
rect 44310 8583 44313 8629
rect 44313 8583 44359 8629
rect 44359 8583 44362 8629
rect 44310 8580 44362 8583
rect 44470 8583 44473 8629
rect 44473 8583 44519 8629
rect 44519 8583 44522 8629
rect 44470 8580 44522 8583
rect 43750 8038 43753 8090
rect 43753 8038 43799 8090
rect 43799 8038 43802 8090
rect 43750 7934 43753 7986
rect 43753 7934 43799 7986
rect 43799 7934 43802 7986
rect 44071 8432 44073 8484
rect 44073 8432 44119 8484
rect 44119 8432 44123 8484
rect 44071 8328 44073 8380
rect 44073 8328 44119 8380
rect 44119 8328 44123 8380
rect 44711 8432 44713 8484
rect 44713 8432 44759 8484
rect 44759 8432 44763 8484
rect 44711 8328 44713 8380
rect 44713 8328 44759 8380
rect 44759 8328 44763 8380
rect 45670 9098 45673 9150
rect 45673 9098 45719 9150
rect 45719 9098 45722 9150
rect 45670 8994 45673 9046
rect 45673 8994 45719 9046
rect 45719 8994 45722 9046
rect 45030 8038 45033 8090
rect 45033 8038 45079 8090
rect 45079 8038 45082 8090
rect 45030 7934 45033 7986
rect 45033 7934 45079 7986
rect 45079 7934 45082 7986
rect 45351 8432 45353 8484
rect 45353 8432 45399 8484
rect 45399 8432 45403 8484
rect 45351 8328 45353 8380
rect 45353 8328 45399 8380
rect 45399 8328 45403 8380
rect 45670 8038 45673 8090
rect 45673 8038 45719 8090
rect 45719 8038 45722 8090
rect 45670 7934 45673 7986
rect 45673 7934 45719 7986
rect 45719 7934 45722 7986
rect 47246 11218 47249 11270
rect 47249 11218 47295 11270
rect 47295 11218 47298 11270
rect 47246 11114 47249 11166
rect 47249 11114 47295 11166
rect 47295 11114 47298 11166
rect 47565 11612 47569 11664
rect 47569 11612 47615 11664
rect 47615 11612 47617 11664
rect 47565 11508 47569 11560
rect 47569 11508 47615 11560
rect 47615 11508 47617 11560
rect 48446 11809 48498 11812
rect 48606 11809 48658 11812
rect 48446 11763 48449 11809
rect 48449 11763 48495 11809
rect 48495 11763 48498 11809
rect 48446 11760 48498 11763
rect 48606 11763 48609 11809
rect 48609 11763 48655 11809
rect 48655 11763 48658 11809
rect 48606 11760 48658 11763
rect 47886 11218 47889 11270
rect 47889 11218 47935 11270
rect 47935 11218 47938 11270
rect 47886 11114 47889 11166
rect 47889 11114 47935 11166
rect 47935 11114 47938 11166
rect 48205 11612 48209 11664
rect 48209 11612 48255 11664
rect 48255 11612 48257 11664
rect 48205 11508 48209 11560
rect 48209 11508 48255 11560
rect 48255 11508 48257 11560
rect 47246 10158 47249 10210
rect 47249 10158 47295 10210
rect 47295 10158 47298 10210
rect 47246 10054 47249 10106
rect 47249 10054 47295 10106
rect 47295 10054 47298 10106
rect 47565 10552 47569 10604
rect 47569 10552 47615 10604
rect 47615 10552 47617 10604
rect 47565 10448 47569 10500
rect 47569 10448 47615 10500
rect 47615 10448 47617 10500
rect 48845 11612 48849 11664
rect 48849 11612 48895 11664
rect 48895 11612 48897 11664
rect 48845 11508 48849 11560
rect 48849 11508 48895 11560
rect 48895 11508 48897 11560
rect 49166 11218 49169 11270
rect 49169 11218 49215 11270
rect 49215 11218 49218 11270
rect 49166 11114 49169 11166
rect 49169 11114 49215 11166
rect 49215 11114 49218 11166
rect 49485 11612 49489 11664
rect 49489 11612 49535 11664
rect 49535 11612 49537 11664
rect 49485 11508 49489 11560
rect 49489 11508 49535 11560
rect 49535 11508 49537 11560
rect 48446 10749 48498 10752
rect 48606 10749 48658 10752
rect 48446 10703 48449 10749
rect 48449 10703 48495 10749
rect 48495 10703 48498 10749
rect 48446 10700 48498 10703
rect 48606 10703 48609 10749
rect 48609 10703 48655 10749
rect 48655 10703 48658 10749
rect 48606 10700 48658 10703
rect 47886 10158 47889 10210
rect 47889 10158 47935 10210
rect 47935 10158 47938 10210
rect 47886 10054 47889 10106
rect 47889 10054 47935 10106
rect 47935 10054 47938 10106
rect 48205 10552 48209 10604
rect 48209 10552 48255 10604
rect 48255 10552 48257 10604
rect 48205 10448 48209 10500
rect 48209 10448 48255 10500
rect 48255 10448 48257 10500
rect 47246 9098 47249 9150
rect 47249 9098 47295 9150
rect 47295 9098 47298 9150
rect 47246 8994 47249 9046
rect 47249 8994 47295 9046
rect 47295 8994 47298 9046
rect 47565 9492 47569 9544
rect 47569 9492 47615 9544
rect 47615 9492 47617 9544
rect 47565 9388 47569 9440
rect 47569 9388 47615 9440
rect 47615 9388 47617 9440
rect 48845 10552 48849 10604
rect 48849 10552 48895 10604
rect 48895 10552 48897 10604
rect 48845 10448 48849 10500
rect 48849 10448 48895 10500
rect 48895 10448 48897 10500
rect 49806 11218 49809 11270
rect 49809 11218 49855 11270
rect 49855 11218 49858 11270
rect 49806 11114 49809 11166
rect 49809 11114 49855 11166
rect 49855 11114 49858 11166
rect 49166 10158 49169 10210
rect 49169 10158 49215 10210
rect 49215 10158 49218 10210
rect 49166 10054 49169 10106
rect 49169 10054 49215 10106
rect 49215 10054 49218 10106
rect 49485 10552 49489 10604
rect 49489 10552 49535 10604
rect 49535 10552 49537 10604
rect 49485 10448 49489 10500
rect 49489 10448 49535 10500
rect 49535 10448 49537 10500
rect 48446 9689 48498 9692
rect 48606 9689 48658 9692
rect 48446 9643 48449 9689
rect 48449 9643 48495 9689
rect 48495 9643 48498 9689
rect 48446 9640 48498 9643
rect 48606 9643 48609 9689
rect 48609 9643 48655 9689
rect 48655 9643 48658 9689
rect 48606 9640 48658 9643
rect 47886 9098 47889 9150
rect 47889 9098 47935 9150
rect 47935 9098 47938 9150
rect 47886 8994 47889 9046
rect 47889 8994 47935 9046
rect 47935 8994 47938 9046
rect 48205 9492 48209 9544
rect 48209 9492 48255 9544
rect 48255 9492 48257 9544
rect 48205 9388 48209 9440
rect 48209 9388 48255 9440
rect 48255 9388 48257 9440
rect 47246 8038 47249 8090
rect 47249 8038 47295 8090
rect 47295 8038 47298 8090
rect 47246 7934 47249 7986
rect 47249 7934 47295 7986
rect 47295 7934 47298 7986
rect 47565 8432 47569 8484
rect 47569 8432 47615 8484
rect 47615 8432 47617 8484
rect 47565 8328 47569 8380
rect 47569 8328 47615 8380
rect 47615 8328 47617 8380
rect 48845 9492 48849 9544
rect 48849 9492 48895 9544
rect 48895 9492 48897 9544
rect 48845 9388 48849 9440
rect 48849 9388 48895 9440
rect 48895 9388 48897 9440
rect 49806 10158 49809 10210
rect 49809 10158 49855 10210
rect 49855 10158 49858 10210
rect 49806 10054 49809 10106
rect 49809 10054 49855 10106
rect 49855 10054 49858 10106
rect 49166 9098 49169 9150
rect 49169 9098 49215 9150
rect 49215 9098 49218 9150
rect 49166 8994 49169 9046
rect 49169 8994 49215 9046
rect 49215 8994 49218 9046
rect 49485 9492 49489 9544
rect 49489 9492 49535 9544
rect 49535 9492 49537 9544
rect 49485 9388 49489 9440
rect 49489 9388 49535 9440
rect 49535 9388 49537 9440
rect 48446 8629 48498 8632
rect 48606 8629 48658 8632
rect 48446 8583 48449 8629
rect 48449 8583 48495 8629
rect 48495 8583 48498 8629
rect 48446 8580 48498 8583
rect 48606 8583 48609 8629
rect 48609 8583 48655 8629
rect 48655 8583 48658 8629
rect 48606 8580 48658 8583
rect 47886 8038 47889 8090
rect 47889 8038 47935 8090
rect 47935 8038 47938 8090
rect 47886 7934 47889 7986
rect 47889 7934 47935 7986
rect 47935 7934 47938 7986
rect 48205 8432 48209 8484
rect 48209 8432 48255 8484
rect 48255 8432 48257 8484
rect 48205 8328 48209 8380
rect 48209 8328 48255 8380
rect 48255 8328 48257 8380
rect 48845 8432 48849 8484
rect 48849 8432 48895 8484
rect 48895 8432 48897 8484
rect 48845 8328 48849 8380
rect 48849 8328 48895 8380
rect 48895 8328 48897 8380
rect 49806 9098 49809 9150
rect 49809 9098 49855 9150
rect 49855 9098 49858 9150
rect 49806 8994 49809 9046
rect 49809 8994 49855 9046
rect 49855 8994 49858 9046
rect 49166 8038 49169 8090
rect 49169 8038 49215 8090
rect 49215 8038 49218 8090
rect 49166 7934 49169 7986
rect 49169 7934 49215 7986
rect 49215 7934 49218 7986
rect 49485 8432 49489 8484
rect 49489 8432 49535 8484
rect 49535 8432 49537 8484
rect 49485 8328 49489 8380
rect 49489 8328 49535 8380
rect 49535 8328 49537 8380
rect 49806 8038 49809 8090
rect 49809 8038 49855 8090
rect 49855 8038 49858 8090
rect 49806 7934 49809 7986
rect 49809 7934 49855 7986
rect 49855 7934 49858 7986
rect 52806 11218 52809 11270
rect 52809 11218 52855 11270
rect 52855 11218 52858 11270
rect 52806 11114 52809 11166
rect 52809 11114 52855 11166
rect 52855 11114 52858 11166
rect 53127 11612 53129 11664
rect 53129 11612 53175 11664
rect 53175 11612 53179 11664
rect 53127 11508 53129 11560
rect 53129 11508 53175 11560
rect 53175 11508 53179 11560
rect 54006 11809 54058 11812
rect 54166 11809 54218 11812
rect 54006 11763 54009 11809
rect 54009 11763 54055 11809
rect 54055 11763 54058 11809
rect 54006 11760 54058 11763
rect 54166 11763 54169 11809
rect 54169 11763 54215 11809
rect 54215 11763 54218 11809
rect 54166 11760 54218 11763
rect 53446 11218 53449 11270
rect 53449 11218 53495 11270
rect 53495 11218 53498 11270
rect 53446 11114 53449 11166
rect 53449 11114 53495 11166
rect 53495 11114 53498 11166
rect 53767 11612 53769 11664
rect 53769 11612 53815 11664
rect 53815 11612 53819 11664
rect 53767 11508 53769 11560
rect 53769 11508 53815 11560
rect 53815 11508 53819 11560
rect 54407 11612 54409 11664
rect 54409 11612 54455 11664
rect 54455 11612 54459 11664
rect 54407 11508 54409 11560
rect 54409 11508 54455 11560
rect 54455 11508 54459 11560
rect 54726 11218 54729 11270
rect 54729 11218 54775 11270
rect 54775 11218 54778 11270
rect 54726 11114 54729 11166
rect 54729 11114 54775 11166
rect 54775 11114 54778 11166
rect 55047 11612 55049 11664
rect 55049 11612 55095 11664
rect 55095 11612 55099 11664
rect 55047 11508 55049 11560
rect 55049 11508 55095 11560
rect 55095 11508 55099 11560
rect 52806 10158 52809 10210
rect 52809 10158 52855 10210
rect 52855 10158 52858 10210
rect 52806 10054 52809 10106
rect 52809 10054 52855 10106
rect 52855 10054 52858 10106
rect 53127 10552 53129 10604
rect 53129 10552 53175 10604
rect 53175 10552 53179 10604
rect 53127 10448 53129 10500
rect 53129 10448 53175 10500
rect 53175 10448 53179 10500
rect 54006 10749 54058 10752
rect 54166 10749 54218 10752
rect 54006 10703 54009 10749
rect 54009 10703 54055 10749
rect 54055 10703 54058 10749
rect 54006 10700 54058 10703
rect 54166 10703 54169 10749
rect 54169 10703 54215 10749
rect 54215 10703 54218 10749
rect 54166 10700 54218 10703
rect 53446 10158 53449 10210
rect 53449 10158 53495 10210
rect 53495 10158 53498 10210
rect 53446 10054 53449 10106
rect 53449 10054 53495 10106
rect 53495 10054 53498 10106
rect 53767 10552 53769 10604
rect 53769 10552 53815 10604
rect 53815 10552 53819 10604
rect 53767 10448 53769 10500
rect 53769 10448 53815 10500
rect 53815 10448 53819 10500
rect 54407 10552 54409 10604
rect 54409 10552 54455 10604
rect 54455 10552 54459 10604
rect 54407 10448 54409 10500
rect 54409 10448 54455 10500
rect 54455 10448 54459 10500
rect 55366 11218 55369 11270
rect 55369 11218 55415 11270
rect 55415 11218 55418 11270
rect 55366 11114 55369 11166
rect 55369 11114 55415 11166
rect 55415 11114 55418 11166
rect 54726 10158 54729 10210
rect 54729 10158 54775 10210
rect 54775 10158 54778 10210
rect 54726 10054 54729 10106
rect 54729 10054 54775 10106
rect 54775 10054 54778 10106
rect 55047 10552 55049 10604
rect 55049 10552 55095 10604
rect 55095 10552 55099 10604
rect 55047 10448 55049 10500
rect 55049 10448 55095 10500
rect 55095 10448 55099 10500
rect 52806 9098 52809 9150
rect 52809 9098 52855 9150
rect 52855 9098 52858 9150
rect 52806 8994 52809 9046
rect 52809 8994 52855 9046
rect 52855 8994 52858 9046
rect 53127 9492 53129 9544
rect 53129 9492 53175 9544
rect 53175 9492 53179 9544
rect 53127 9388 53129 9440
rect 53129 9388 53175 9440
rect 53175 9388 53179 9440
rect 54006 9689 54058 9692
rect 54166 9689 54218 9692
rect 54006 9643 54009 9689
rect 54009 9643 54055 9689
rect 54055 9643 54058 9689
rect 54006 9640 54058 9643
rect 54166 9643 54169 9689
rect 54169 9643 54215 9689
rect 54215 9643 54218 9689
rect 54166 9640 54218 9643
rect 53446 9098 53449 9150
rect 53449 9098 53495 9150
rect 53495 9098 53498 9150
rect 53446 8994 53449 9046
rect 53449 8994 53495 9046
rect 53495 8994 53498 9046
rect 53767 9492 53769 9544
rect 53769 9492 53815 9544
rect 53815 9492 53819 9544
rect 53767 9388 53769 9440
rect 53769 9388 53815 9440
rect 53815 9388 53819 9440
rect 54407 9492 54409 9544
rect 54409 9492 54455 9544
rect 54455 9492 54459 9544
rect 54407 9388 54409 9440
rect 54409 9388 54455 9440
rect 54455 9388 54459 9440
rect 55366 10158 55369 10210
rect 55369 10158 55415 10210
rect 55415 10158 55418 10210
rect 55366 10054 55369 10106
rect 55369 10054 55415 10106
rect 55415 10054 55418 10106
rect 54726 9098 54729 9150
rect 54729 9098 54775 9150
rect 54775 9098 54778 9150
rect 54726 8994 54729 9046
rect 54729 8994 54775 9046
rect 54775 8994 54778 9046
rect 55047 9492 55049 9544
rect 55049 9492 55095 9544
rect 55095 9492 55099 9544
rect 55047 9388 55049 9440
rect 55049 9388 55095 9440
rect 55095 9388 55099 9440
rect 52806 8038 52809 8090
rect 52809 8038 52855 8090
rect 52855 8038 52858 8090
rect 52806 7934 52809 7986
rect 52809 7934 52855 7986
rect 52855 7934 52858 7986
rect 53127 8432 53129 8484
rect 53129 8432 53175 8484
rect 53175 8432 53179 8484
rect 53127 8328 53129 8380
rect 53129 8328 53175 8380
rect 53175 8328 53179 8380
rect 54006 8629 54058 8632
rect 54166 8629 54218 8632
rect 54006 8583 54009 8629
rect 54009 8583 54055 8629
rect 54055 8583 54058 8629
rect 54006 8580 54058 8583
rect 54166 8583 54169 8629
rect 54169 8583 54215 8629
rect 54215 8583 54218 8629
rect 54166 8580 54218 8583
rect 53446 8038 53449 8090
rect 53449 8038 53495 8090
rect 53495 8038 53498 8090
rect 53446 7934 53449 7986
rect 53449 7934 53495 7986
rect 53495 7934 53498 7986
rect 53767 8432 53769 8484
rect 53769 8432 53815 8484
rect 53815 8432 53819 8484
rect 53767 8328 53769 8380
rect 53769 8328 53815 8380
rect 53815 8328 53819 8380
rect 54407 8432 54409 8484
rect 54409 8432 54455 8484
rect 54455 8432 54459 8484
rect 54407 8328 54409 8380
rect 54409 8328 54455 8380
rect 54455 8328 54459 8380
rect 55366 9098 55369 9150
rect 55369 9098 55415 9150
rect 55415 9098 55418 9150
rect 55366 8994 55369 9046
rect 55369 8994 55415 9046
rect 55415 8994 55418 9046
rect 54726 8038 54729 8090
rect 54729 8038 54775 8090
rect 54775 8038 54778 8090
rect 54726 7934 54729 7986
rect 54729 7934 54775 7986
rect 54775 7934 54778 7986
rect 55047 8432 55049 8484
rect 55049 8432 55095 8484
rect 55095 8432 55099 8484
rect 55047 8328 55049 8380
rect 55049 8328 55095 8380
rect 55095 8328 55099 8380
rect 55366 8038 55369 8090
rect 55369 8038 55415 8090
rect 55415 8038 55418 8090
rect 55366 7934 55369 7986
rect 55369 7934 55415 7986
rect 55415 7934 55418 7986
rect 56942 11218 56945 11270
rect 56945 11218 56991 11270
rect 56991 11218 56994 11270
rect 56942 11114 56945 11166
rect 56945 11114 56991 11166
rect 56991 11114 56994 11166
rect 57261 11612 57265 11664
rect 57265 11612 57311 11664
rect 57311 11612 57313 11664
rect 57261 11508 57265 11560
rect 57265 11508 57311 11560
rect 57311 11508 57313 11560
rect 58142 11809 58194 11812
rect 58302 11809 58354 11812
rect 58142 11763 58145 11809
rect 58145 11763 58191 11809
rect 58191 11763 58194 11809
rect 58142 11760 58194 11763
rect 58302 11763 58305 11809
rect 58305 11763 58351 11809
rect 58351 11763 58354 11809
rect 58302 11760 58354 11763
rect 57582 11218 57585 11270
rect 57585 11218 57631 11270
rect 57631 11218 57634 11270
rect 57582 11114 57585 11166
rect 57585 11114 57631 11166
rect 57631 11114 57634 11166
rect 57901 11612 57905 11664
rect 57905 11612 57951 11664
rect 57951 11612 57953 11664
rect 57901 11508 57905 11560
rect 57905 11508 57951 11560
rect 57951 11508 57953 11560
rect 56942 10158 56945 10210
rect 56945 10158 56991 10210
rect 56991 10158 56994 10210
rect 56942 10054 56945 10106
rect 56945 10054 56991 10106
rect 56991 10054 56994 10106
rect 57261 10552 57265 10604
rect 57265 10552 57311 10604
rect 57311 10552 57313 10604
rect 57261 10448 57265 10500
rect 57265 10448 57311 10500
rect 57311 10448 57313 10500
rect 58541 11612 58545 11664
rect 58545 11612 58591 11664
rect 58591 11612 58593 11664
rect 58541 11508 58545 11560
rect 58545 11508 58591 11560
rect 58591 11508 58593 11560
rect 58862 11218 58865 11270
rect 58865 11218 58911 11270
rect 58911 11218 58914 11270
rect 58862 11114 58865 11166
rect 58865 11114 58911 11166
rect 58911 11114 58914 11166
rect 59181 11612 59185 11664
rect 59185 11612 59231 11664
rect 59231 11612 59233 11664
rect 59181 11508 59185 11560
rect 59185 11508 59231 11560
rect 59231 11508 59233 11560
rect 58142 10749 58194 10752
rect 58302 10749 58354 10752
rect 58142 10703 58145 10749
rect 58145 10703 58191 10749
rect 58191 10703 58194 10749
rect 58142 10700 58194 10703
rect 58302 10703 58305 10749
rect 58305 10703 58351 10749
rect 58351 10703 58354 10749
rect 58302 10700 58354 10703
rect 57582 10158 57585 10210
rect 57585 10158 57631 10210
rect 57631 10158 57634 10210
rect 57582 10054 57585 10106
rect 57585 10054 57631 10106
rect 57631 10054 57634 10106
rect 57901 10552 57905 10604
rect 57905 10552 57951 10604
rect 57951 10552 57953 10604
rect 57901 10448 57905 10500
rect 57905 10448 57951 10500
rect 57951 10448 57953 10500
rect 56942 9098 56945 9150
rect 56945 9098 56991 9150
rect 56991 9098 56994 9150
rect 56942 8994 56945 9046
rect 56945 8994 56991 9046
rect 56991 8994 56994 9046
rect 57261 9492 57265 9544
rect 57265 9492 57311 9544
rect 57311 9492 57313 9544
rect 57261 9388 57265 9440
rect 57265 9388 57311 9440
rect 57311 9388 57313 9440
rect 58541 10552 58545 10604
rect 58545 10552 58591 10604
rect 58591 10552 58593 10604
rect 58541 10448 58545 10500
rect 58545 10448 58591 10500
rect 58591 10448 58593 10500
rect 59502 11218 59505 11270
rect 59505 11218 59551 11270
rect 59551 11218 59554 11270
rect 59502 11114 59505 11166
rect 59505 11114 59551 11166
rect 59551 11114 59554 11166
rect 58862 10158 58865 10210
rect 58865 10158 58911 10210
rect 58911 10158 58914 10210
rect 58862 10054 58865 10106
rect 58865 10054 58911 10106
rect 58911 10054 58914 10106
rect 59181 10552 59185 10604
rect 59185 10552 59231 10604
rect 59231 10552 59233 10604
rect 59181 10448 59185 10500
rect 59185 10448 59231 10500
rect 59231 10448 59233 10500
rect 58142 9689 58194 9692
rect 58302 9689 58354 9692
rect 58142 9643 58145 9689
rect 58145 9643 58191 9689
rect 58191 9643 58194 9689
rect 58142 9640 58194 9643
rect 58302 9643 58305 9689
rect 58305 9643 58351 9689
rect 58351 9643 58354 9689
rect 58302 9640 58354 9643
rect 57582 9098 57585 9150
rect 57585 9098 57631 9150
rect 57631 9098 57634 9150
rect 57582 8994 57585 9046
rect 57585 8994 57631 9046
rect 57631 8994 57634 9046
rect 57901 9492 57905 9544
rect 57905 9492 57951 9544
rect 57951 9492 57953 9544
rect 57901 9388 57905 9440
rect 57905 9388 57951 9440
rect 57951 9388 57953 9440
rect 56942 8038 56945 8090
rect 56945 8038 56991 8090
rect 56991 8038 56994 8090
rect 56942 7934 56945 7986
rect 56945 7934 56991 7986
rect 56991 7934 56994 7986
rect 57261 8432 57265 8484
rect 57265 8432 57311 8484
rect 57311 8432 57313 8484
rect 57261 8328 57265 8380
rect 57265 8328 57311 8380
rect 57311 8328 57313 8380
rect 58541 9492 58545 9544
rect 58545 9492 58591 9544
rect 58591 9492 58593 9544
rect 58541 9388 58545 9440
rect 58545 9388 58591 9440
rect 58591 9388 58593 9440
rect 59502 10158 59505 10210
rect 59505 10158 59551 10210
rect 59551 10158 59554 10210
rect 59502 10054 59505 10106
rect 59505 10054 59551 10106
rect 59551 10054 59554 10106
rect 58862 9098 58865 9150
rect 58865 9098 58911 9150
rect 58911 9098 58914 9150
rect 58862 8994 58865 9046
rect 58865 8994 58911 9046
rect 58911 8994 58914 9046
rect 59181 9492 59185 9544
rect 59185 9492 59231 9544
rect 59231 9492 59233 9544
rect 59181 9388 59185 9440
rect 59185 9388 59231 9440
rect 59231 9388 59233 9440
rect 58142 8629 58194 8632
rect 58302 8629 58354 8632
rect 58142 8583 58145 8629
rect 58145 8583 58191 8629
rect 58191 8583 58194 8629
rect 58142 8580 58194 8583
rect 58302 8583 58305 8629
rect 58305 8583 58351 8629
rect 58351 8583 58354 8629
rect 58302 8580 58354 8583
rect 57582 8038 57585 8090
rect 57585 8038 57631 8090
rect 57631 8038 57634 8090
rect 57582 7934 57585 7986
rect 57585 7934 57631 7986
rect 57631 7934 57634 7986
rect 57901 8432 57905 8484
rect 57905 8432 57951 8484
rect 57951 8432 57953 8484
rect 57901 8328 57905 8380
rect 57905 8328 57951 8380
rect 57951 8328 57953 8380
rect 58541 8432 58545 8484
rect 58545 8432 58591 8484
rect 58591 8432 58593 8484
rect 58541 8328 58545 8380
rect 58545 8328 58591 8380
rect 58591 8328 58593 8380
rect 59502 9098 59505 9150
rect 59505 9098 59551 9150
rect 59551 9098 59554 9150
rect 59502 8994 59505 9046
rect 59505 8994 59551 9046
rect 59551 8994 59554 9046
rect 58862 8038 58865 8090
rect 58865 8038 58911 8090
rect 58911 8038 58914 8090
rect 58862 7934 58865 7986
rect 58865 7934 58911 7986
rect 58911 7934 58914 7986
rect 59181 8432 59185 8484
rect 59185 8432 59231 8484
rect 59231 8432 59233 8484
rect 59181 8328 59185 8380
rect 59185 8328 59231 8380
rect 59231 8328 59233 8380
rect 59502 8038 59505 8090
rect 59505 8038 59551 8090
rect 59551 8038 59554 8090
rect 59502 7934 59505 7986
rect 59505 7934 59551 7986
rect 59551 7934 59554 7986
rect 62502 11218 62505 11270
rect 62505 11218 62551 11270
rect 62551 11218 62554 11270
rect 62502 11114 62505 11166
rect 62505 11114 62551 11166
rect 62551 11114 62554 11166
rect 62823 11612 62825 11664
rect 62825 11612 62871 11664
rect 62871 11612 62875 11664
rect 62823 11508 62825 11560
rect 62825 11508 62871 11560
rect 62871 11508 62875 11560
rect 63702 11809 63754 11812
rect 63862 11809 63914 11812
rect 63702 11763 63705 11809
rect 63705 11763 63751 11809
rect 63751 11763 63754 11809
rect 63702 11760 63754 11763
rect 63862 11763 63865 11809
rect 63865 11763 63911 11809
rect 63911 11763 63914 11809
rect 63862 11760 63914 11763
rect 63142 11218 63145 11270
rect 63145 11218 63191 11270
rect 63191 11218 63194 11270
rect 63142 11114 63145 11166
rect 63145 11114 63191 11166
rect 63191 11114 63194 11166
rect 63463 11612 63465 11664
rect 63465 11612 63511 11664
rect 63511 11612 63515 11664
rect 63463 11508 63465 11560
rect 63465 11508 63511 11560
rect 63511 11508 63515 11560
rect 64103 11612 64105 11664
rect 64105 11612 64151 11664
rect 64151 11612 64155 11664
rect 64103 11508 64105 11560
rect 64105 11508 64151 11560
rect 64151 11508 64155 11560
rect 64422 11218 64425 11270
rect 64425 11218 64471 11270
rect 64471 11218 64474 11270
rect 64422 11114 64425 11166
rect 64425 11114 64471 11166
rect 64471 11114 64474 11166
rect 64743 11612 64745 11664
rect 64745 11612 64791 11664
rect 64791 11612 64795 11664
rect 64743 11508 64745 11560
rect 64745 11508 64791 11560
rect 64791 11508 64795 11560
rect 62502 10158 62505 10210
rect 62505 10158 62551 10210
rect 62551 10158 62554 10210
rect 62502 10054 62505 10106
rect 62505 10054 62551 10106
rect 62551 10054 62554 10106
rect 62823 10552 62825 10604
rect 62825 10552 62871 10604
rect 62871 10552 62875 10604
rect 62823 10448 62825 10500
rect 62825 10448 62871 10500
rect 62871 10448 62875 10500
rect 63702 10749 63754 10752
rect 63862 10749 63914 10752
rect 63702 10703 63705 10749
rect 63705 10703 63751 10749
rect 63751 10703 63754 10749
rect 63702 10700 63754 10703
rect 63862 10703 63865 10749
rect 63865 10703 63911 10749
rect 63911 10703 63914 10749
rect 63862 10700 63914 10703
rect 63142 10158 63145 10210
rect 63145 10158 63191 10210
rect 63191 10158 63194 10210
rect 63142 10054 63145 10106
rect 63145 10054 63191 10106
rect 63191 10054 63194 10106
rect 63463 10552 63465 10604
rect 63465 10552 63511 10604
rect 63511 10552 63515 10604
rect 63463 10448 63465 10500
rect 63465 10448 63511 10500
rect 63511 10448 63515 10500
rect 64103 10552 64105 10604
rect 64105 10552 64151 10604
rect 64151 10552 64155 10604
rect 64103 10448 64105 10500
rect 64105 10448 64151 10500
rect 64151 10448 64155 10500
rect 65062 11218 65065 11270
rect 65065 11218 65111 11270
rect 65111 11218 65114 11270
rect 65062 11114 65065 11166
rect 65065 11114 65111 11166
rect 65111 11114 65114 11166
rect 64422 10158 64425 10210
rect 64425 10158 64471 10210
rect 64471 10158 64474 10210
rect 64422 10054 64425 10106
rect 64425 10054 64471 10106
rect 64471 10054 64474 10106
rect 64743 10552 64745 10604
rect 64745 10552 64791 10604
rect 64791 10552 64795 10604
rect 64743 10448 64745 10500
rect 64745 10448 64791 10500
rect 64791 10448 64795 10500
rect 62502 9098 62505 9150
rect 62505 9098 62551 9150
rect 62551 9098 62554 9150
rect 62502 8994 62505 9046
rect 62505 8994 62551 9046
rect 62551 8994 62554 9046
rect 62823 9492 62825 9544
rect 62825 9492 62871 9544
rect 62871 9492 62875 9544
rect 62823 9388 62825 9440
rect 62825 9388 62871 9440
rect 62871 9388 62875 9440
rect 63702 9689 63754 9692
rect 63862 9689 63914 9692
rect 63702 9643 63705 9689
rect 63705 9643 63751 9689
rect 63751 9643 63754 9689
rect 63702 9640 63754 9643
rect 63862 9643 63865 9689
rect 63865 9643 63911 9689
rect 63911 9643 63914 9689
rect 63862 9640 63914 9643
rect 63142 9098 63145 9150
rect 63145 9098 63191 9150
rect 63191 9098 63194 9150
rect 63142 8994 63145 9046
rect 63145 8994 63191 9046
rect 63191 8994 63194 9046
rect 63463 9492 63465 9544
rect 63465 9492 63511 9544
rect 63511 9492 63515 9544
rect 63463 9388 63465 9440
rect 63465 9388 63511 9440
rect 63511 9388 63515 9440
rect 64103 9492 64105 9544
rect 64105 9492 64151 9544
rect 64151 9492 64155 9544
rect 64103 9388 64105 9440
rect 64105 9388 64151 9440
rect 64151 9388 64155 9440
rect 65062 10158 65065 10210
rect 65065 10158 65111 10210
rect 65111 10158 65114 10210
rect 65062 10054 65065 10106
rect 65065 10054 65111 10106
rect 65111 10054 65114 10106
rect 64422 9098 64425 9150
rect 64425 9098 64471 9150
rect 64471 9098 64474 9150
rect 64422 8994 64425 9046
rect 64425 8994 64471 9046
rect 64471 8994 64474 9046
rect 64743 9492 64745 9544
rect 64745 9492 64791 9544
rect 64791 9492 64795 9544
rect 64743 9388 64745 9440
rect 64745 9388 64791 9440
rect 64791 9388 64795 9440
rect 62502 8038 62505 8090
rect 62505 8038 62551 8090
rect 62551 8038 62554 8090
rect 62502 7934 62505 7986
rect 62505 7934 62551 7986
rect 62551 7934 62554 7986
rect 62823 8432 62825 8484
rect 62825 8432 62871 8484
rect 62871 8432 62875 8484
rect 62823 8328 62825 8380
rect 62825 8328 62871 8380
rect 62871 8328 62875 8380
rect 63702 8629 63754 8632
rect 63862 8629 63914 8632
rect 63702 8583 63705 8629
rect 63705 8583 63751 8629
rect 63751 8583 63754 8629
rect 63702 8580 63754 8583
rect 63862 8583 63865 8629
rect 63865 8583 63911 8629
rect 63911 8583 63914 8629
rect 63862 8580 63914 8583
rect 63142 8038 63145 8090
rect 63145 8038 63191 8090
rect 63191 8038 63194 8090
rect 63142 7934 63145 7986
rect 63145 7934 63191 7986
rect 63191 7934 63194 7986
rect 63463 8432 63465 8484
rect 63465 8432 63511 8484
rect 63511 8432 63515 8484
rect 63463 8328 63465 8380
rect 63465 8328 63511 8380
rect 63511 8328 63515 8380
rect 64103 8432 64105 8484
rect 64105 8432 64151 8484
rect 64151 8432 64155 8484
rect 64103 8328 64105 8380
rect 64105 8328 64151 8380
rect 64151 8328 64155 8380
rect 65062 9098 65065 9150
rect 65065 9098 65111 9150
rect 65111 9098 65114 9150
rect 65062 8994 65065 9046
rect 65065 8994 65111 9046
rect 65111 8994 65114 9046
rect 64422 8038 64425 8090
rect 64425 8038 64471 8090
rect 64471 8038 64474 8090
rect 64422 7934 64425 7986
rect 64425 7934 64471 7986
rect 64471 7934 64474 7986
rect 64743 8432 64745 8484
rect 64745 8432 64791 8484
rect 64791 8432 64795 8484
rect 64743 8328 64745 8380
rect 64745 8328 64791 8380
rect 64791 8328 64795 8380
rect 65062 8038 65065 8090
rect 65065 8038 65111 8090
rect 65111 8038 65114 8090
rect 65062 7934 65065 7986
rect 65065 7934 65111 7986
rect 65111 7934 65114 7986
rect 2187 5256 2239 5308
rect 2291 5256 2343 5308
rect 2187 5152 2239 5204
rect 2291 5152 2343 5204
rect 3059 5121 3111 5173
rect 3163 5121 3215 5173
rect 3059 5017 3111 5069
rect 3163 5017 3215 5069
rect 8287 6357 8339 6409
rect 8391 6357 8443 6409
rect 8287 6253 8339 6305
rect 8391 6253 8443 6305
rect 11383 6384 11435 6436
rect 11487 6384 11539 6436
rect 17131 6384 17183 6436
rect 17235 6384 17287 6436
rect 17339 6384 17391 6436
rect 11383 6280 11435 6332
rect 11487 6280 11539 6332
rect 17131 6280 17183 6332
rect 17235 6280 17287 6332
rect 17339 6280 17391 6332
rect 6879 6121 6931 6173
rect 6983 6121 7035 6173
rect 9981 6121 10033 6173
rect 10085 6121 10137 6173
rect 11383 6176 11435 6228
rect 11487 6176 11539 6228
rect 17131 6176 17183 6228
rect 17235 6176 17287 6228
rect 17339 6176 17391 6228
rect 6879 6017 6931 6069
rect 6983 6017 7035 6069
rect 9981 6017 10033 6069
rect 5156 5407 5208 5459
rect 5260 5407 5312 5459
rect 5156 5303 5208 5355
rect 5260 5303 5312 5355
rect 2187 4553 2239 4556
rect 2187 4507 2190 4553
rect 2190 4507 2236 4553
rect 2236 4507 2239 4553
rect 2187 4504 2239 4507
rect 2291 4553 2343 4556
rect 2291 4507 2294 4553
rect 2294 4507 2340 4553
rect 2340 4507 2343 4553
rect 2291 4504 2343 4507
rect 2727 4367 2730 4419
rect 2730 4367 2776 4419
rect 2776 4367 2779 4419
rect 2727 4263 2730 4315
rect 2730 4263 2776 4315
rect 2776 4263 2779 4315
rect 3591 3753 3594 3805
rect 3594 3753 3640 3805
rect 3640 3753 3643 3805
rect 3591 3649 3594 3701
rect 3594 3649 3640 3701
rect 3640 3649 3643 3701
rect 4023 4077 4026 4129
rect 4026 4077 4072 4129
rect 4072 4077 4075 4129
rect 4023 3973 4026 4025
rect 4026 3973 4072 4025
rect 4072 3973 4075 4025
rect 6556 4049 6608 4101
rect 6660 4049 6712 4101
rect 6556 3945 6608 3997
rect 6660 3945 6712 3997
rect 2737 3107 2738 3159
rect 2738 3107 2784 3159
rect 2784 3107 2789 3159
rect 2737 3003 2738 3055
rect 2738 3003 2784 3055
rect 2784 3003 2789 3055
rect 3111 3107 3114 3159
rect 3114 3107 3160 3159
rect 3160 3107 3163 3159
rect 3111 3003 3114 3055
rect 3114 3003 3160 3055
rect 3160 3003 3163 3055
rect 3431 3107 3434 3159
rect 3434 3107 3480 3159
rect 3480 3107 3483 3159
rect 3431 3003 3434 3055
rect 3434 3003 3480 3055
rect 3480 3003 3483 3055
rect 3935 2491 3938 2543
rect 3938 2491 3984 2543
rect 3984 2491 3987 2543
rect 3935 2387 3938 2439
rect 3938 2387 3984 2439
rect 3984 2387 3987 2439
rect 3983 1721 4035 1773
rect 3983 1617 4035 1669
rect 9201 5935 9253 5938
rect 9201 5889 9204 5935
rect 9204 5889 9250 5935
rect 9250 5889 9253 5935
rect 9201 5886 9253 5889
rect 7681 5657 7684 5709
rect 7684 5657 7730 5709
rect 7730 5657 7733 5709
rect 7681 5553 7684 5605
rect 7684 5553 7730 5605
rect 7730 5553 7733 5605
rect 7841 5657 7844 5709
rect 7844 5657 7890 5709
rect 7890 5657 7893 5709
rect 7841 5553 7844 5605
rect 7844 5553 7890 5605
rect 7890 5553 7893 5605
rect 8161 5657 8164 5709
rect 8164 5657 8210 5709
rect 8210 5657 8213 5709
rect 8161 5553 8164 5605
rect 8164 5553 8210 5605
rect 8210 5553 8213 5605
rect 8481 5657 8484 5709
rect 8484 5657 8530 5709
rect 8530 5657 8533 5709
rect 8481 5553 8484 5605
rect 8484 5553 8530 5605
rect 8530 5553 8533 5605
rect 8801 5657 8804 5709
rect 8804 5657 8850 5709
rect 8850 5657 8853 5709
rect 8801 5553 8804 5605
rect 8804 5553 8850 5605
rect 8850 5553 8853 5605
rect 8961 5657 8964 5709
rect 8964 5657 9010 5709
rect 9010 5657 9013 5709
rect 8961 5553 8964 5605
rect 8964 5553 9010 5605
rect 9010 5553 9013 5605
rect 9121 5657 9124 5709
rect 9124 5657 9170 5709
rect 9170 5657 9173 5709
rect 9121 5553 9124 5605
rect 9124 5553 9170 5605
rect 9170 5553 9173 5605
rect 9280 5350 9332 5402
rect 7841 5121 7844 5173
rect 7844 5121 7890 5173
rect 7890 5121 7893 5173
rect 7841 5017 7844 5069
rect 7844 5017 7890 5069
rect 7890 5017 7893 5069
rect 8001 5121 8004 5173
rect 8004 5121 8050 5173
rect 8050 5121 8053 5173
rect 8001 5017 8004 5069
rect 8004 5017 8050 5069
rect 8050 5017 8053 5069
rect 8161 5121 8164 5173
rect 8164 5121 8210 5173
rect 8210 5121 8213 5173
rect 8161 5017 8164 5069
rect 8164 5017 8210 5069
rect 8210 5017 8213 5069
rect 8481 5121 8484 5173
rect 8484 5121 8530 5173
rect 8530 5121 8533 5173
rect 8481 5017 8484 5069
rect 8484 5017 8530 5069
rect 8530 5017 8533 5069
rect 8801 5121 8804 5173
rect 8804 5121 8850 5173
rect 8850 5121 8853 5173
rect 8801 5017 8804 5069
rect 8804 5017 8850 5069
rect 8850 5017 8853 5069
rect 9121 5121 9124 5173
rect 9124 5121 9170 5173
rect 9170 5121 9173 5173
rect 9121 5017 9124 5069
rect 9124 5017 9170 5069
rect 9170 5017 9173 5069
rect 9083 4814 9135 4866
rect 7681 4585 7684 4637
rect 7684 4585 7730 4637
rect 7730 4585 7733 4637
rect 7681 4481 7684 4533
rect 7684 4481 7730 4533
rect 7730 4481 7733 4533
rect 7841 4585 7844 4637
rect 7844 4585 7890 4637
rect 7890 4585 7893 4637
rect 7841 4481 7844 4533
rect 7844 4481 7890 4533
rect 7890 4481 7893 4533
rect 8161 4585 8164 4637
rect 8164 4585 8210 4637
rect 8210 4585 8213 4637
rect 8161 4481 8164 4533
rect 8164 4481 8210 4533
rect 8210 4481 8213 4533
rect 8481 4585 8484 4637
rect 8484 4585 8530 4637
rect 8530 4585 8533 4637
rect 8481 4481 8484 4533
rect 8484 4481 8530 4533
rect 8530 4481 8533 4533
rect 8801 4585 8804 4637
rect 8804 4585 8850 4637
rect 8850 4585 8853 4637
rect 8801 4481 8804 4533
rect 8804 4481 8850 4533
rect 8850 4481 8853 4533
rect 8961 4585 8964 4637
rect 8964 4585 9010 4637
rect 9010 4585 9013 4637
rect 8961 4481 8964 4533
rect 8964 4481 9010 4533
rect 9010 4481 9013 4533
rect 9121 4585 9124 4637
rect 9124 4585 9170 4637
rect 9170 4585 9173 4637
rect 9121 4481 9124 4533
rect 9124 4481 9170 4533
rect 9170 4481 9173 4533
rect 9201 4329 9253 4332
rect 9201 4283 9204 4329
rect 9204 4283 9250 4329
rect 9250 4283 9253 4329
rect 9201 4280 9253 4283
rect 7841 4049 7844 4101
rect 7844 4049 7890 4101
rect 7890 4049 7893 4101
rect 7841 3945 7844 3997
rect 7844 3945 7890 3997
rect 7890 3945 7893 3997
rect 8001 4049 8004 4101
rect 8004 4049 8050 4101
rect 8050 4049 8053 4101
rect 8001 3945 8004 3997
rect 8004 3945 8050 3997
rect 8050 3945 8053 3997
rect 8161 4049 8164 4101
rect 8164 4049 8210 4101
rect 8210 4049 8213 4101
rect 8161 3945 8164 3997
rect 8164 3945 8210 3997
rect 8210 3945 8213 3997
rect 8481 4049 8484 4101
rect 8484 4049 8530 4101
rect 8530 4049 8533 4101
rect 8481 3945 8484 3997
rect 8484 3945 8530 3997
rect 8530 3945 8533 3997
rect 8801 4049 8804 4101
rect 8804 4049 8850 4101
rect 8850 4049 8853 4101
rect 8801 3945 8804 3997
rect 8804 3945 8850 3997
rect 8850 3945 8853 3997
rect 9121 4049 9124 4101
rect 9124 4049 9170 4101
rect 9170 4049 9173 4101
rect 9121 3945 9124 3997
rect 9124 3945 9170 3997
rect 9170 3945 9173 3997
rect 9280 3744 9332 3796
rect 7841 3521 7844 3573
rect 7844 3521 7890 3573
rect 7890 3521 7893 3573
rect 7841 3417 7844 3469
rect 7844 3417 7890 3469
rect 7890 3417 7893 3469
rect 8161 3521 8164 3573
rect 8164 3521 8210 3573
rect 8210 3521 8213 3573
rect 8161 3417 8164 3469
rect 8164 3417 8210 3469
rect 8210 3417 8213 3469
rect 8481 3521 8484 3573
rect 8484 3521 8530 3573
rect 8530 3521 8533 3573
rect 8481 3417 8484 3469
rect 8484 3417 8530 3469
rect 8530 3417 8533 3469
rect 8801 3521 8804 3573
rect 8804 3521 8850 3573
rect 8850 3521 8853 3573
rect 8801 3417 8804 3469
rect 8804 3417 8850 3469
rect 8850 3417 8853 3469
rect 8961 3513 8964 3565
rect 8964 3513 9010 3565
rect 9010 3513 9013 3565
rect 8961 3409 8964 3461
rect 8964 3409 9010 3461
rect 9010 3409 9013 3461
rect 9121 3521 9124 3573
rect 9124 3521 9170 3573
rect 9170 3521 9173 3573
rect 9121 3417 9124 3469
rect 9124 3417 9170 3469
rect 9170 3417 9173 3469
rect 9280 3229 9332 3281
rect 7841 2985 7844 3037
rect 7844 2985 7890 3037
rect 7890 2985 7893 3037
rect 7841 2881 7844 2933
rect 7844 2881 7890 2933
rect 7890 2881 7893 2933
rect 8001 2977 8004 3029
rect 8004 2977 8050 3029
rect 8050 2977 8053 3029
rect 8001 2873 8004 2925
rect 8004 2873 8050 2925
rect 8050 2873 8053 2925
rect 8161 2985 8164 3037
rect 8164 2985 8210 3037
rect 8210 2985 8213 3037
rect 8161 2881 8164 2933
rect 8164 2881 8210 2933
rect 8210 2881 8213 2933
rect 8481 2985 8484 3037
rect 8484 2985 8530 3037
rect 8530 2985 8533 3037
rect 8481 2881 8484 2933
rect 8484 2881 8530 2933
rect 8530 2881 8533 2933
rect 8801 2985 8804 3037
rect 8804 2985 8850 3037
rect 8850 2985 8853 3037
rect 8801 2881 8804 2933
rect 8804 2881 8850 2933
rect 8850 2881 8853 2933
rect 9121 2985 9124 3037
rect 9124 2985 9170 3037
rect 9170 2985 9173 3037
rect 9121 2881 9124 2933
rect 9124 2881 9170 2933
rect 9170 2881 9173 2933
rect 10085 6017 10137 6069
rect 10290 5990 10342 6042
rect 10394 5990 10446 6042
rect 10290 5886 10342 5938
rect 10394 5886 10446 5938
rect 11651 6042 11703 6094
rect 11755 6042 11807 6094
rect 17568 6042 17620 6094
rect 17672 6042 17724 6094
rect 17776 6042 17828 6094
rect 11651 5938 11703 5990
rect 11755 5938 11807 5990
rect 17568 5938 17620 5990
rect 17672 5938 17724 5990
rect 17776 5938 17828 5990
rect 11651 5834 11703 5886
rect 11755 5834 11807 5886
rect 17568 5834 17620 5886
rect 17672 5834 17724 5886
rect 17776 5834 17828 5886
rect 14698 5657 14750 5709
rect 14802 5657 14854 5709
rect 14698 5553 14750 5605
rect 14802 5553 14854 5605
rect 10556 5392 10608 5444
rect 10660 5392 10712 5444
rect 17346 5392 17398 5444
rect 17450 5392 17502 5444
rect 10556 5288 10608 5340
rect 10660 5288 10712 5340
rect 17346 5288 17398 5340
rect 17450 5288 17502 5340
rect 8881 2675 8884 2709
rect 8884 2675 8930 2709
rect 8930 2675 8933 2709
rect 8881 2657 8933 2675
rect 7394 2587 7446 2639
rect 7498 2587 7550 2639
rect 6594 2348 6597 2400
rect 6597 2348 6643 2400
rect 6643 2348 6646 2400
rect 6594 2244 6597 2296
rect 6597 2244 6643 2296
rect 6643 2244 6646 2296
rect 7394 2483 7446 2535
rect 7498 2519 7550 2535
rect 10325 2633 10377 2636
rect 10325 2587 10328 2633
rect 10328 2587 10374 2633
rect 10374 2587 10377 2633
rect 10325 2584 10377 2587
rect 10429 2633 10481 2636
rect 10429 2587 10432 2633
rect 10432 2587 10478 2633
rect 10478 2587 10481 2633
rect 10429 2584 10481 2587
rect 7498 2483 7523 2519
rect 7523 2483 7550 2519
rect 10325 2529 10377 2532
rect 10325 2483 10328 2529
rect 10328 2483 10374 2529
rect 10374 2483 10377 2529
rect 10325 2480 10377 2483
rect 10429 2529 10481 2532
rect 10429 2483 10432 2529
rect 10432 2483 10478 2529
rect 10478 2483 10481 2529
rect 10429 2480 10481 2483
rect 9749 2352 9795 2404
rect 9795 2352 9801 2404
rect 9853 2352 9905 2404
rect 9749 2248 9795 2300
rect 9795 2248 9801 2300
rect 9853 2248 9905 2300
rect 9408 1952 9460 2004
rect 9512 1952 9564 2004
rect 6524 1907 6576 1910
rect 6524 1861 6527 1907
rect 6527 1861 6573 1907
rect 6573 1861 6576 1907
rect 6524 1858 6576 1861
rect 6628 1907 6680 1910
rect 6628 1861 6631 1907
rect 6631 1861 6677 1907
rect 6677 1861 6680 1907
rect 6628 1858 6680 1861
rect 9408 1882 9460 1900
rect 6434 1719 6437 1771
rect 6437 1719 6483 1771
rect 6483 1719 6486 1771
rect 6434 1615 6437 1667
rect 6437 1615 6483 1667
rect 6483 1615 6486 1667
rect 6866 1713 6869 1765
rect 6869 1713 6915 1765
rect 6915 1713 6918 1765
rect 6866 1609 6869 1661
rect 6869 1609 6915 1661
rect 6915 1609 6918 1661
rect 9408 1848 9443 1882
rect 9443 1848 9460 1882
rect 9512 1882 9564 1900
rect 9512 1848 9557 1882
rect 9557 1848 9564 1882
rect 11317 1952 11369 2004
rect 11421 1952 11473 2004
rect 11317 1848 11369 1900
rect 11421 1848 11473 1900
rect 13112 2242 13115 2294
rect 13115 2242 13161 2294
rect 13161 2242 13164 2294
rect 13112 2138 13115 2190
rect 13115 2138 13161 2190
rect 13161 2138 13164 2190
rect 13112 2034 13115 2086
rect 13115 2034 13161 2086
rect 13161 2034 13164 2086
rect 13212 1812 13264 1815
rect 13212 1766 13215 1812
rect 13215 1766 13261 1812
rect 13261 1766 13264 1812
rect 13212 1763 13264 1766
rect 13316 1812 13368 1815
rect 13316 1766 13319 1812
rect 13319 1766 13365 1812
rect 13365 1766 13368 1812
rect 13316 1763 13368 1766
rect 13212 1708 13264 1711
rect 13212 1662 13215 1708
rect 13215 1662 13261 1708
rect 13261 1662 13264 1708
rect 13212 1659 13264 1662
rect 13316 1708 13368 1711
rect 13316 1662 13319 1708
rect 13319 1662 13365 1708
rect 13365 1662 13368 1708
rect 13316 1659 13368 1662
rect 15064 3510 15067 3562
rect 15067 3510 15113 3562
rect 15113 3510 15116 3562
rect 15064 3406 15067 3458
rect 15067 3406 15113 3458
rect 15113 3406 15116 3458
rect 15672 3510 15675 3562
rect 15675 3510 15721 3562
rect 15721 3510 15724 3562
rect 15672 3406 15675 3458
rect 15675 3406 15721 3458
rect 15721 3406 15724 3458
rect 16280 3510 16283 3562
rect 16283 3510 16329 3562
rect 16329 3510 16332 3562
rect 16280 3406 16283 3458
rect 16283 3406 16329 3458
rect 16329 3406 16332 3458
rect 16183 2760 16235 2763
rect 16183 2714 16186 2760
rect 16186 2714 16232 2760
rect 16232 2714 16235 2760
rect 16183 2711 16235 2714
rect 16287 2760 16339 2763
rect 16287 2714 16290 2760
rect 16290 2714 16336 2760
rect 16336 2714 16339 2760
rect 16287 2711 16339 2714
rect 16391 2760 16443 2763
rect 16391 2714 16394 2760
rect 16394 2714 16440 2760
rect 16440 2714 16443 2760
rect 16391 2711 16443 2714
rect 16183 2656 16235 2659
rect 16183 2610 16186 2656
rect 16186 2610 16232 2656
rect 16232 2610 16235 2656
rect 16183 2607 16235 2610
rect 16287 2656 16339 2659
rect 16287 2610 16290 2656
rect 16290 2610 16336 2656
rect 16336 2610 16339 2656
rect 16287 2607 16339 2610
rect 16391 2656 16443 2659
rect 16391 2610 16394 2656
rect 16394 2610 16440 2656
rect 16440 2610 16443 2656
rect 16391 2607 16443 2610
rect 14224 1832 14276 1835
rect 14224 1786 14227 1832
rect 14227 1786 14273 1832
rect 14273 1786 14276 1832
rect 14224 1783 14276 1786
rect 14328 1832 14380 1835
rect 14328 1786 14331 1832
rect 14331 1786 14377 1832
rect 14377 1786 14380 1832
rect 14328 1783 14380 1786
rect 14432 1832 14484 1835
rect 14432 1786 14435 1832
rect 14435 1786 14481 1832
rect 14481 1786 14484 1832
rect 14432 1783 14484 1786
rect 15672 2242 15675 2294
rect 15675 2242 15721 2294
rect 15721 2242 15724 2294
rect 15672 2138 15675 2190
rect 15675 2138 15721 2190
rect 15721 2138 15724 2190
rect 15672 2034 15675 2086
rect 15675 2034 15721 2086
rect 15721 2034 15724 2086
rect 19112 2204 19115 2256
rect 19115 2204 19161 2256
rect 19161 2204 19164 2256
rect 19112 2100 19115 2152
rect 19115 2100 19161 2152
rect 19161 2100 19164 2152
rect 19112 1996 19115 2048
rect 19115 1996 19161 2048
rect 19161 1996 19164 2048
rect 19432 2204 19435 2256
rect 19435 2204 19481 2256
rect 19481 2204 19484 2256
rect 19432 2100 19435 2152
rect 19435 2100 19481 2152
rect 19481 2100 19484 2152
rect 19432 1996 19435 2048
rect 19435 1996 19481 2048
rect 19481 1996 19484 2048
rect 19752 2204 19755 2256
rect 19755 2204 19801 2256
rect 19801 2204 19804 2256
rect 19752 2100 19755 2152
rect 19755 2100 19801 2152
rect 19801 2100 19804 2152
rect 19752 1996 19755 2048
rect 19755 1996 19801 2048
rect 19801 1996 19804 2048
rect 20072 2204 20075 2256
rect 20075 2204 20121 2256
rect 20121 2204 20124 2256
rect 20072 2100 20075 2152
rect 20075 2100 20121 2152
rect 20121 2100 20124 2152
rect 20072 1996 20075 2048
rect 20075 1996 20121 2048
rect 20121 1996 20124 2048
rect 20659 4915 20711 4918
rect 20659 4869 20662 4915
rect 20662 4869 20708 4915
rect 20708 4869 20711 4915
rect 20659 4866 20711 4869
rect 20763 4915 20815 4918
rect 20763 4869 20766 4915
rect 20766 4869 20812 4915
rect 20812 4869 20815 4915
rect 20763 4866 20815 4869
rect 20392 2204 20395 2256
rect 20395 2204 20441 2256
rect 20441 2204 20444 2256
rect 20392 2100 20395 2152
rect 20395 2100 20441 2152
rect 20441 2100 20444 2152
rect 20392 1996 20395 2048
rect 20395 1996 20441 2048
rect 20441 1996 20444 2048
rect 20712 2204 20715 2256
rect 20715 2204 20761 2256
rect 20761 2204 20764 2256
rect 20712 2100 20715 2152
rect 20715 2100 20761 2152
rect 20761 2100 20764 2152
rect 20712 1996 20715 2048
rect 20715 1996 20761 2048
rect 20761 1996 20764 2048
rect 21032 2204 21035 2256
rect 21035 2204 21081 2256
rect 21081 2204 21084 2256
rect 21032 2100 21035 2152
rect 21035 2100 21081 2152
rect 21081 2100 21084 2152
rect 21032 1996 21035 2048
rect 21035 1996 21081 2048
rect 21081 1996 21084 2048
rect 21672 4412 21675 4464
rect 21675 4412 21721 4464
rect 21721 4412 21724 4464
rect 21672 4308 21675 4360
rect 21675 4308 21721 4360
rect 21721 4308 21724 4360
rect 21672 4204 21675 4256
rect 21675 4204 21721 4256
rect 21721 4204 21724 4256
rect 21643 1901 21695 1904
rect 21643 1855 21646 1901
rect 21646 1855 21692 1901
rect 21692 1855 21695 1901
rect 21643 1852 21695 1855
rect 21747 1901 21799 1904
rect 21747 1855 21750 1901
rect 21750 1855 21796 1901
rect 21796 1855 21799 1901
rect 21747 1852 21799 1855
rect 21851 1901 21903 1904
rect 21851 1855 21854 1901
rect 21854 1855 21900 1901
rect 21900 1855 21903 1901
rect 21851 1852 21903 1855
rect 24130 4961 24182 5013
rect 24234 4961 24286 5013
rect 24130 4906 24182 4909
rect 24234 4906 24286 4909
rect 24130 4860 24182 4906
rect 24234 4860 24286 4906
rect 24130 4857 24182 4860
rect 24234 4857 24286 4860
rect 27492 4253 27544 4305
rect 27596 4253 27648 4305
rect 27492 4149 27544 4201
rect 27596 4149 27648 4201
rect 27490 2934 27542 2937
rect 27594 2934 27646 2937
rect 27490 2888 27542 2934
rect 27594 2888 27646 2934
rect 27490 2885 27542 2888
rect 27594 2885 27646 2888
rect 27490 2781 27542 2833
rect 27594 2781 27646 2833
rect 24130 1802 24182 1805
rect 24234 1802 24286 1805
rect 24578 1802 24630 1805
rect 24682 1802 24734 1805
rect 24130 1756 24182 1802
rect 24234 1756 24286 1802
rect 24578 1756 24630 1802
rect 24682 1756 24734 1802
rect 24130 1753 24182 1756
rect 24234 1753 24286 1756
rect 24130 1649 24182 1701
rect 24234 1649 24286 1701
rect 24578 1753 24630 1756
rect 24682 1753 24734 1756
rect 24578 1649 24630 1701
rect 24682 1649 24734 1701
rect 30300 5090 30352 5093
rect 30404 5090 30456 5093
rect 30300 5044 30307 5090
rect 30307 5044 30352 5090
rect 30404 5044 30456 5090
rect 30300 5041 30352 5044
rect 30404 5041 30456 5044
rect 30508 5041 30560 5093
rect 30612 5090 30664 5093
rect 30716 5090 30768 5093
rect 30612 5044 30664 5090
rect 30716 5044 30761 5090
rect 30761 5044 30768 5090
rect 30612 5041 30664 5044
rect 30716 5041 30768 5044
rect 30300 4937 30352 4989
rect 30404 4937 30456 4989
rect 30508 4937 30560 4989
rect 30612 4937 30664 4989
rect 30716 4937 30768 4989
rect 30300 4833 30352 4885
rect 30404 4833 30456 4885
rect 30508 4833 30560 4885
rect 30612 4833 30664 4885
rect 30716 4833 30768 4885
rect 30300 4085 30352 4137
rect 30404 4085 30456 4137
rect 30508 4085 30560 4137
rect 30612 4085 30664 4137
rect 30716 4085 30768 4137
rect 30300 3981 30352 4033
rect 30404 3981 30456 4033
rect 30508 3981 30560 4033
rect 30612 3981 30664 4033
rect 30716 3981 30768 4033
rect 30300 3877 30352 3929
rect 30404 3877 30456 3929
rect 30508 3877 30560 3929
rect 30612 3877 30664 3929
rect 30716 3877 30768 3929
rect 30300 3773 30352 3825
rect 30404 3773 30456 3825
rect 30508 3773 30560 3825
rect 30612 3773 30664 3825
rect 30716 3773 30768 3825
rect 30300 3718 30352 3721
rect 30404 3718 30456 3721
rect 30300 3672 30307 3718
rect 30307 3672 30352 3718
rect 30404 3672 30456 3718
rect 30300 3669 30352 3672
rect 30404 3669 30456 3672
rect 30508 3669 30560 3721
rect 30612 3718 30664 3721
rect 30716 3718 30768 3721
rect 30612 3672 30664 3718
rect 30716 3672 30761 3718
rect 30761 3672 30768 3718
rect 30612 3669 30664 3672
rect 30716 3669 30768 3672
rect 29740 3078 29792 3081
rect 29844 3078 29896 3081
rect 29740 3032 29747 3078
rect 29747 3032 29792 3078
rect 29844 3032 29896 3078
rect 29740 3029 29792 3032
rect 29844 3029 29896 3032
rect 29948 3029 30000 3081
rect 30052 3078 30104 3081
rect 30156 3078 30208 3081
rect 30052 3032 30104 3078
rect 30156 3032 30201 3078
rect 30201 3032 30208 3078
rect 30052 3029 30104 3032
rect 30156 3029 30208 3032
rect 29740 2925 29792 2977
rect 29844 2925 29896 2977
rect 29948 2925 30000 2977
rect 30052 2925 30104 2977
rect 30156 2925 30208 2977
rect 29740 2821 29792 2873
rect 29844 2821 29896 2873
rect 29948 2821 30000 2873
rect 30052 2821 30104 2873
rect 30156 2821 30208 2873
rect 30300 2073 30352 2125
rect 30404 2073 30456 2125
rect 30508 2073 30560 2125
rect 30612 2073 30664 2125
rect 30716 2073 30768 2125
rect 30300 1969 30352 2021
rect 30404 1969 30456 2021
rect 30508 1969 30560 2021
rect 30612 1969 30664 2021
rect 30716 1969 30768 2021
rect 30300 1865 30352 1917
rect 30404 1865 30456 1917
rect 30508 1865 30560 1917
rect 30612 1865 30664 1917
rect 30716 1865 30768 1917
rect 30300 1761 30352 1813
rect 30404 1761 30456 1813
rect 30508 1761 30560 1813
rect 30612 1761 30664 1813
rect 30716 1761 30768 1813
rect 30300 1706 30352 1709
rect 30404 1706 30456 1709
rect 30300 1660 30307 1706
rect 30307 1660 30352 1706
rect 30404 1660 30456 1706
rect 30300 1657 30352 1660
rect 30404 1657 30456 1660
rect 30508 1657 30560 1709
rect 30612 1706 30664 1709
rect 30716 1706 30768 1709
rect 30612 1660 30664 1706
rect 30716 1660 30761 1706
rect 30761 1660 30768 1706
rect 30612 1657 30664 1660
rect 30716 1657 30768 1660
rect 12030 1075 12082 1127
rect 12134 1075 12186 1127
rect 12030 971 12082 1023
rect 12134 971 12186 1023
rect 45034 1149 45086 1201
rect 45138 1149 45190 1201
rect 45242 1149 45294 1201
rect 45346 1149 45398 1201
rect 45450 1149 45502 1201
rect 49474 1149 49526 1201
rect 49578 1149 49630 1201
rect 49682 1149 49734 1201
rect 49786 1149 49838 1201
rect 49890 1149 49942 1201
rect 35204 1049 35256 1101
rect 35308 1049 35360 1101
rect 35412 1049 35464 1101
rect 35516 1049 35568 1101
rect 35620 1049 35672 1101
rect 39644 1049 39696 1101
rect 39748 1049 39800 1101
rect 39852 1049 39904 1101
rect 39956 1049 40008 1101
rect 40060 1049 40112 1101
rect 35204 945 35256 997
rect 35308 945 35360 997
rect 35412 945 35464 997
rect 35516 945 35568 997
rect 35620 945 35672 997
rect 39644 945 39696 997
rect 39748 945 39800 997
rect 39852 945 39904 997
rect 39956 945 40008 997
rect 40060 945 40112 997
rect 35204 841 35256 893
rect 35308 841 35360 893
rect 35412 841 35464 893
rect 35516 841 35568 893
rect 35620 841 35672 893
rect 39644 841 39696 893
rect 39748 841 39800 893
rect 39852 841 39904 893
rect 39956 841 40008 893
rect 40060 841 40112 893
rect 21643 720 21695 772
rect 21747 720 21799 772
rect 21851 720 21903 772
rect 21643 616 21695 668
rect 21747 616 21799 668
rect 21851 616 21903 668
rect 35204 737 35256 789
rect 35308 737 35360 789
rect 35412 737 35464 789
rect 35516 737 35568 789
rect 35620 737 35672 789
rect 39644 737 39696 789
rect 39748 737 39800 789
rect 39852 737 39904 789
rect 39956 737 40008 789
rect 40060 737 40112 789
rect 45034 1045 45086 1097
rect 45138 1045 45190 1097
rect 45242 1045 45294 1097
rect 45346 1045 45398 1097
rect 45450 1045 45502 1097
rect 49474 1045 49526 1097
rect 49578 1045 49630 1097
rect 49682 1045 49734 1097
rect 49786 1045 49838 1097
rect 49890 1045 49942 1097
rect 45034 941 45086 993
rect 45138 941 45190 993
rect 45242 941 45294 993
rect 45346 941 45398 993
rect 45450 941 45502 993
rect 49474 941 49526 993
rect 49578 941 49630 993
rect 49682 941 49734 993
rect 49786 941 49838 993
rect 49890 941 49942 993
rect 45034 837 45086 889
rect 45138 837 45190 889
rect 45242 837 45294 889
rect 45346 837 45398 889
rect 45450 837 45502 889
rect 49474 837 49526 889
rect 49578 837 49630 889
rect 49682 837 49734 889
rect 49786 837 49838 889
rect 49890 837 49942 889
rect 45034 733 45086 785
rect 45138 733 45190 785
rect 45242 733 45294 785
rect 45346 733 45398 785
rect 45450 733 45502 785
rect 49474 733 49526 785
rect 49578 733 49630 785
rect 49682 733 49734 785
rect 49786 733 49838 785
rect 49890 733 49942 785
rect 35204 633 35256 685
rect 35308 633 35360 685
rect 35412 633 35464 685
rect 35516 633 35568 685
rect 35620 633 35672 685
rect 39644 633 39696 685
rect 39748 633 39800 685
rect 39852 633 39904 685
rect 39956 633 40008 685
rect 40060 633 40112 685
rect 21643 512 21695 564
rect 21747 512 21799 564
rect 21851 512 21903 564
rect 15568 220 15620 272
rect 15672 220 15724 272
rect 15776 220 15828 272
rect 15568 116 15620 168
rect 15672 116 15724 168
rect 15776 116 15828 168
rect 15568 12 15620 64
rect 15672 12 15724 64
rect 15776 12 15828 64
<< metal2 >>
rect 31218 15706 31505 15718
rect 31218 15650 31226 15706
rect 31282 15705 31336 15706
rect 31392 15705 31446 15706
rect 31282 15653 31334 15705
rect 31392 15653 31438 15705
rect 31282 15650 31336 15653
rect 31392 15650 31446 15653
rect 31502 15650 31505 15706
rect 31218 15601 31505 15650
rect 31218 15596 31230 15601
rect 31218 15540 31226 15596
rect 31282 15549 31334 15601
rect 31386 15596 31438 15601
rect 31490 15596 31505 15601
rect 31392 15549 31438 15596
rect 31282 15540 31336 15549
rect 31392 15540 31446 15549
rect 31502 15540 31505 15596
rect 31218 15497 31505 15540
rect 31218 15486 31230 15497
rect 31218 15430 31226 15486
rect 31282 15445 31334 15497
rect 31386 15486 31438 15497
rect 31490 15486 31505 15497
rect 31392 15445 31438 15486
rect 31282 15430 31336 15445
rect 31392 15430 31446 15445
rect 31502 15430 31505 15486
rect 31218 15420 31505 15430
rect 826 14773 1083 14774
rect -7190 14772 1260 14773
rect -7190 14742 1700 14772
rect -7190 14686 1233 14742
rect 1289 14686 1343 14742
rect 1399 14686 1453 14742
rect 1509 14686 1563 14742
rect 1619 14686 1700 14742
rect -7190 14632 1700 14686
rect -7190 14576 1233 14632
rect 1289 14576 1343 14632
rect 1399 14576 1453 14632
rect 1509 14576 1563 14632
rect 1619 14576 1700 14632
rect -7190 14490 1700 14576
rect -8178 13055 -7966 13067
rect -8178 12999 -8163 13055
rect -8107 12999 -8053 13055
rect -7997 13045 -7966 13055
rect -7190 13045 -6907 14490
rect 976 14489 1700 14490
rect 1224 14488 1700 14489
rect 1803 14325 2238 14334
rect -3119 14321 2238 14325
rect -3119 14265 1812 14321
rect 1868 14265 1922 14321
rect 1978 14265 2032 14321
rect 2088 14265 2142 14321
rect 2198 14265 2238 14321
rect -3119 14211 2238 14265
rect -3119 14206 1812 14211
rect -3120 14155 1812 14206
rect 1868 14155 1922 14211
rect 1978 14155 2032 14211
rect 2088 14155 2142 14211
rect 2198 14155 2238 14211
rect 3161 14328 3341 14338
rect 3161 14272 3171 14328
rect 3227 14272 3275 14328
rect 3331 14272 3341 14328
rect 3161 14224 3341 14272
rect 3161 14168 3171 14224
rect 3227 14168 3275 14224
rect 3331 14168 3341 14224
rect 3161 14158 3341 14168
rect 3950 14328 4026 14338
rect 3950 14272 3960 14328
rect 4016 14272 4026 14328
rect 3950 14224 4026 14272
rect 3950 14168 3960 14224
rect 4016 14168 4026 14224
rect 3950 14158 4026 14168
rect 5731 14274 5911 14284
rect 5731 14218 5741 14274
rect 5797 14218 5845 14274
rect 5901 14218 5911 14274
rect 5731 14170 5911 14218
rect -3120 14101 2238 14155
rect -3120 14049 1812 14101
rect -7997 12999 -6907 13045
rect -8178 12945 -6907 12999
rect -8178 12889 -8163 12945
rect -8107 12889 -8053 12945
rect -7997 12889 -6907 12945
rect -8178 12888 -6907 12889
rect -8178 12855 -7966 12888
rect -7190 12588 -6907 12888
rect -7088 10356 -6931 12588
rect -3626 10729 -3414 10752
rect -3626 10673 -3604 10729
rect -3548 10673 -3494 10729
rect -3438 10673 -3414 10729
rect -3626 10619 -3414 10673
rect -3626 10563 -3604 10619
rect -3548 10563 -3494 10619
rect -3438 10563 -3414 10619
rect -3626 10540 -3414 10563
rect -3601 10435 -3444 10540
rect -3602 10427 -3416 10435
rect -3602 10371 -3594 10427
rect -3538 10371 -3484 10427
rect -3428 10371 -3416 10427
rect -7106 10345 -6906 10356
rect -7106 10289 -7089 10345
rect -7033 10289 -6979 10345
rect -6923 10289 -6906 10345
rect -7106 10283 -6906 10289
rect -6826 10345 -6626 10356
rect -6826 10289 -6809 10345
rect -6753 10289 -6699 10345
rect -6643 10289 -6626 10345
rect -6826 10283 -6626 10289
rect -3602 10317 -3416 10371
rect -8154 9711 -7942 9721
rect -8154 9655 -8141 9711
rect -8085 9655 -8031 9711
rect -7975 9655 -7942 9711
rect -8154 9646 -7942 9655
rect -6796 9646 -6685 10283
rect -3602 10261 -3594 10317
rect -3538 10261 -3484 10317
rect -3428 10261 -3416 10317
rect -3602 10207 -3416 10261
rect -3602 10151 -3594 10207
rect -3538 10151 -3484 10207
rect -3428 10151 -3416 10207
rect -3602 10097 -3416 10151
rect -3602 10041 -3594 10097
rect -3538 10041 -3484 10097
rect -3428 10041 -3416 10097
rect -3602 9987 -3416 10041
rect -3602 9931 -3594 9987
rect -3538 9931 -3484 9987
rect -3428 9931 -3416 9987
rect -3602 9916 -3416 9931
rect -4586 9780 -4386 9791
rect -4586 9724 -4569 9780
rect -4513 9724 -4459 9780
rect -4403 9724 -4386 9780
rect -4586 9718 -4386 9724
rect -4525 9658 -4425 9718
rect -8154 9606 -6685 9646
rect -8154 9550 -8141 9606
rect -8085 9550 -8031 9606
rect -7975 9550 -6685 9606
rect -8154 9501 -6685 9550
rect -8154 9445 -8141 9501
rect -8085 9445 -8031 9501
rect -7975 9493 -6685 9501
rect -5348 9558 -4425 9658
rect -7975 9445 -7942 9493
rect -8154 9430 -7942 9445
rect -7106 9428 -6906 9493
rect -5348 9439 -5248 9558
rect -7106 9372 -7089 9428
rect -7033 9372 -6979 9428
rect -6923 9372 -6906 9428
rect -7106 9366 -6906 9372
rect -5426 9428 -5226 9439
rect -5426 9372 -5409 9428
rect -5353 9372 -5299 9428
rect -5243 9372 -5226 9428
rect -5426 9366 -5226 9372
rect -4586 9428 -4386 9439
rect -4586 9372 -4569 9428
rect -4513 9372 -4459 9428
rect -4403 9372 -4386 9428
rect -4586 9366 -4386 9372
rect -16674 8972 -4666 9200
rect -6826 8863 -6626 8874
rect -6826 8807 -6809 8863
rect -6753 8807 -6699 8863
rect -6643 8807 -6626 8863
rect -8513 8782 -8303 8794
rect -8513 8726 -8491 8782
rect -8435 8726 -8381 8782
rect -8325 8749 -8303 8782
rect -6826 8749 -6626 8807
rect -4868 8863 -4666 8972
rect -4868 8807 -4849 8863
rect -4793 8807 -4739 8863
rect -4683 8807 -4666 8863
rect -4868 8803 -4666 8807
rect -4866 8801 -4666 8803
rect -8325 8726 -6626 8749
rect -8513 8672 -6626 8726
rect -8513 8616 -8491 8672
rect -8435 8616 -8381 8672
rect -8325 8616 -6626 8672
rect -8513 8578 -6626 8616
rect -8513 8577 -6669 8578
rect -8513 8562 -8303 8577
rect -8513 8506 -8491 8562
rect -8435 8506 -8381 8562
rect -8325 8506 -8303 8562
rect -8513 8452 -8303 8506
rect -8513 8396 -8491 8452
rect -8435 8396 -8381 8452
rect -8325 8396 -8303 8452
rect -7106 8511 -6906 8577
rect -7106 8455 -7089 8511
rect -7033 8455 -6979 8511
rect -6923 8455 -6906 8511
rect -7106 8449 -6906 8455
rect -4586 8511 -4386 8522
rect -4586 8455 -4569 8511
rect -4513 8455 -4459 8511
rect -4403 8455 -4386 8511
rect -4586 8449 -4386 8455
rect -8513 8368 -8303 8396
rect -4564 8289 -4407 8449
rect -3601 8289 -3444 9916
rect -4564 8132 -3444 8289
rect -10593 7925 -10178 7946
rect -10593 7920 -8256 7925
rect -10593 7864 -10576 7920
rect -10520 7864 -10466 7920
rect -10410 7864 -10356 7920
rect -10300 7864 -10246 7920
rect -10190 7864 -8256 7920
rect -10593 7810 -8256 7864
rect -10593 7754 -10576 7810
rect -10520 7754 -10466 7810
rect -10410 7754 -10356 7810
rect -10300 7754 -10246 7810
rect -10190 7754 -8256 7810
rect -10593 7753 -8256 7754
rect -10593 7721 -10178 7753
rect -8428 6415 -8256 7753
rect -3119 6955 -2860 14049
rect 1805 14045 1812 14049
rect 1868 14045 1922 14101
rect 1978 14045 2032 14101
rect 2088 14045 2142 14101
rect 2198 14045 2238 14101
rect 1805 14031 2238 14045
rect 2520 13979 2700 13989
rect 2520 13923 2530 13979
rect 2586 13923 2634 13979
rect 2690 13923 2700 13979
rect 2520 13875 2700 13923
rect 2520 13819 2530 13875
rect 2586 13819 2634 13875
rect 2690 13819 2700 13875
rect 2520 13809 2700 13819
rect 527 13794 1084 13795
rect -1867 13763 1084 13794
rect -1867 13707 554 13763
rect 610 13707 664 13763
rect 720 13707 774 13763
rect 830 13707 884 13763
rect 940 13707 994 13763
rect 1050 13707 1084 13763
rect -1867 13653 1084 13707
rect -1869 13597 554 13653
rect 610 13597 664 13653
rect 720 13597 774 13653
rect 830 13597 884 13653
rect 940 13597 994 13653
rect 1050 13597 1084 13653
rect -1869 13496 1084 13597
rect -4565 6798 -2860 6955
rect -4564 6703 -2860 6798
rect -4564 6543 -4407 6703
rect -7106 6537 -6906 6543
rect -7106 6481 -7089 6537
rect -7033 6481 -6979 6537
rect -6923 6481 -6906 6537
rect -7106 6474 -6906 6481
rect -7107 6415 -6906 6474
rect -4586 6537 -4386 6543
rect -4586 6481 -4569 6537
rect -4513 6481 -4459 6537
rect -4403 6481 -4386 6537
rect -4586 6470 -4386 6481
rect -8428 6243 -6626 6415
rect -6826 6185 -6626 6243
rect -6826 6129 -6809 6185
rect -6753 6129 -6699 6185
rect -6643 6129 -6626 6185
rect -6826 6118 -6626 6129
rect -4866 6185 -4666 6191
rect -4866 6129 -4849 6185
rect -4793 6129 -4739 6185
rect -4683 6129 -4666 6185
rect -4866 6020 -4666 6129
rect -16479 5778 -4666 6020
rect -16479 5777 -4712 5778
rect -7106 5620 -6906 5626
rect -7106 5564 -7089 5620
rect -7033 5564 -6979 5620
rect -6923 5564 -6906 5620
rect -7106 5553 -6906 5564
rect -5426 5620 -5226 5626
rect -5426 5564 -5409 5620
rect -5353 5564 -5299 5620
rect -5243 5564 -5226 5620
rect -5426 5553 -5226 5564
rect -4586 5620 -4386 5626
rect -4586 5564 -4569 5620
rect -4513 5564 -4459 5620
rect -4403 5564 -4386 5620
rect -4586 5553 -4386 5564
rect -8159 5532 -7863 5550
rect -7106 5532 -6989 5553
rect -8215 5476 -8146 5532
rect -8090 5476 -8041 5532
rect -7985 5476 -7936 5532
rect -7880 5476 -6989 5532
rect -8215 5475 -6989 5476
rect -8215 5422 -6685 5475
rect -8215 5366 -8146 5422
rect -8090 5366 -8041 5422
rect -7985 5366 -7936 5422
rect -7880 5366 -6685 5422
rect -8215 5364 -6685 5366
rect -8215 5362 -7108 5364
rect -8159 5338 -7863 5362
rect -6796 4709 -6685 5364
rect -5348 5434 -5248 5553
rect -5348 5334 -4425 5434
rect -4525 5274 -4425 5334
rect -4586 5268 -4386 5274
rect -4586 5212 -4569 5268
rect -4513 5212 -4459 5268
rect -4403 5212 -4386 5268
rect -4586 5201 -4386 5212
rect -7106 4703 -6906 4709
rect -7106 4647 -7089 4703
rect -7033 4647 -6979 4703
rect -6923 4647 -6906 4703
rect -7106 4636 -6906 4647
rect -6826 4703 -6626 4709
rect -6826 4647 -6809 4703
rect -6753 4647 -6699 4703
rect -6643 4647 -6626 4703
rect -6826 4636 -6626 4647
rect -7088 2259 -6931 4636
rect -3601 4452 -3444 6703
rect -3626 4429 -3414 4452
rect -3626 4373 -3604 4429
rect -3548 4373 -3494 4429
rect -3438 4373 -3414 4429
rect -3626 4319 -3414 4373
rect -3626 4263 -3604 4319
rect -3548 4263 -3494 4319
rect -3438 4263 -3414 4319
rect -3626 4240 -3414 4263
rect -1867 2259 -1568 13496
rect 2530 12859 2690 13809
rect 2881 13200 3061 13210
rect 2881 13144 2891 13200
rect 2947 13144 2995 13200
rect 3051 13144 3061 13200
rect 2881 13096 3061 13144
rect 2881 13040 2891 13096
rect 2947 13040 2995 13096
rect 3051 13040 3061 13096
rect 2881 13030 3061 13040
rect 2520 12849 2700 12859
rect 2520 12793 2530 12849
rect 2586 12793 2634 12849
rect 2690 12793 2700 12849
rect 2520 12745 2700 12793
rect 2520 12689 2530 12745
rect 2586 12689 2634 12745
rect 2690 12689 2700 12745
rect 2520 12679 2700 12689
rect 2530 10335 2690 12679
rect 2520 10325 2700 10335
rect 2520 10269 2530 10325
rect 2586 10269 2634 10325
rect 2690 10269 2700 10325
rect 2520 10221 2700 10269
rect 2520 10165 2530 10221
rect 2586 10165 2634 10221
rect 2690 10165 2700 10221
rect 2520 10155 2700 10165
rect 2891 9822 3051 13030
rect 3171 12080 3331 14158
rect 5731 14114 5741 14170
rect 5797 14114 5845 14170
rect 5901 14114 5911 14170
rect 5731 14104 5911 14114
rect 6735 14274 6811 14284
rect 6735 14218 6745 14274
rect 6801 14218 6811 14274
rect 6735 14170 6811 14218
rect 6735 14114 6745 14170
rect 6801 14114 6811 14170
rect 6735 14104 6811 14114
rect 7375 14274 7451 14284
rect 7375 14218 7385 14274
rect 7441 14218 7451 14274
rect 7375 14170 7451 14218
rect 7375 14114 7385 14170
rect 7441 14114 7451 14170
rect 7375 14104 7451 14114
rect 8015 14274 8091 14284
rect 8015 14218 8025 14274
rect 8081 14218 8091 14274
rect 8015 14170 8091 14218
rect 8015 14114 8025 14170
rect 8081 14114 8091 14170
rect 8015 14104 8091 14114
rect 4030 13979 4106 13989
rect 4030 13923 4040 13979
rect 4096 13923 4106 13979
rect 4030 13875 4106 13923
rect 4030 13819 4040 13875
rect 4096 13819 4106 13875
rect 4030 13809 4106 13819
rect 4190 13979 4266 13989
rect 4190 13923 4200 13979
rect 4256 13923 4266 13979
rect 4190 13875 4266 13923
rect 4190 13819 4200 13875
rect 4256 13819 4266 13875
rect 4190 13809 4266 13819
rect 4831 13979 4907 13989
rect 4831 13923 4841 13979
rect 4897 13923 4907 13979
rect 4831 13875 4907 13923
rect 4831 13819 4841 13875
rect 4897 13819 4907 13875
rect 4831 13809 4907 13819
rect 5741 13493 5901 14104
rect 6003 13979 6183 13989
rect 6003 13923 6013 13979
rect 6069 13923 6117 13979
rect 6173 13923 6183 13979
rect 6003 13875 6183 13923
rect 6003 13819 6013 13875
rect 6069 13819 6117 13875
rect 6173 13819 6183 13875
rect 6003 13809 6183 13819
rect 7055 13979 7131 13989
rect 7055 13923 7065 13979
rect 7121 13923 7131 13979
rect 7055 13875 7131 13923
rect 7055 13819 7065 13875
rect 7121 13819 7131 13875
rect 7055 13809 7131 13819
rect 7695 13979 7771 13989
rect 7695 13923 7705 13979
rect 7761 13923 7771 13979
rect 7695 13875 7771 13923
rect 7695 13819 7705 13875
rect 7761 13819 7771 13875
rect 7695 13809 7771 13819
rect 3870 13483 3946 13493
rect 3870 13427 3880 13483
rect 3936 13427 3946 13483
rect 3870 13379 3946 13427
rect 3870 13323 3880 13379
rect 3936 13323 3946 13379
rect 3870 13313 3946 13323
rect 4510 13483 4586 13493
rect 4510 13427 4520 13483
rect 4576 13427 4586 13483
rect 4510 13379 4586 13427
rect 4510 13323 4520 13379
rect 4576 13323 4586 13379
rect 4510 13313 4586 13323
rect 5150 13483 5226 13493
rect 5150 13427 5160 13483
rect 5216 13427 5226 13483
rect 5150 13379 5226 13427
rect 5150 13323 5160 13379
rect 5216 13323 5226 13379
rect 5150 13313 5226 13323
rect 5731 13483 5911 13493
rect 5731 13427 5741 13483
rect 5797 13427 5845 13483
rect 5901 13427 5911 13483
rect 5731 13379 5911 13427
rect 5731 13323 5741 13379
rect 5797 13323 5845 13379
rect 5901 13323 5911 13379
rect 5731 13275 5911 13323
rect 5731 13219 5741 13275
rect 5797 13219 5845 13275
rect 5901 13219 5911 13275
rect 3950 13200 4026 13210
rect 5731 13209 5911 13219
rect 3950 13144 3960 13200
rect 4016 13144 4026 13200
rect 3950 13096 4026 13144
rect 3950 13040 3960 13096
rect 4016 13040 4026 13096
rect 3950 13030 4026 13040
rect 5741 12859 5901 13209
rect 6013 13010 6173 13809
rect 11639 13459 11819 13469
rect 11639 13403 11649 13459
rect 11705 13403 11753 13459
rect 11809 13403 11819 13459
rect 7055 13379 7131 13389
rect 7055 13323 7065 13379
rect 7121 13323 7131 13379
rect 7055 13275 7131 13323
rect 7055 13219 7065 13275
rect 7121 13219 7131 13275
rect 7055 13209 7131 13219
rect 7695 13379 7771 13389
rect 7695 13323 7705 13379
rect 7761 13323 7771 13379
rect 7695 13275 7771 13323
rect 11639 13355 11819 13403
rect 11639 13299 11649 13355
rect 11705 13299 11753 13355
rect 11809 13299 11819 13355
rect 11639 13289 11819 13299
rect 17641 13407 17716 13417
rect 17641 13351 17651 13407
rect 17707 13351 17716 13407
rect 7695 13219 7705 13275
rect 7761 13219 7771 13275
rect 7695 13209 7771 13219
rect 6003 13000 6183 13010
rect 6003 12944 6013 13000
rect 6069 12944 6117 13000
rect 6173 12944 6183 13000
rect 6003 12896 6183 12944
rect 4030 12849 4106 12859
rect 4030 12793 4040 12849
rect 4096 12793 4106 12849
rect 4030 12745 4106 12793
rect 4030 12689 4040 12745
rect 4096 12689 4106 12745
rect 4030 12679 4106 12689
rect 4190 12849 4266 12859
rect 4190 12793 4200 12849
rect 4256 12793 4266 12849
rect 4190 12745 4266 12793
rect 4190 12689 4200 12745
rect 4256 12689 4266 12745
rect 4190 12679 4266 12689
rect 4831 12849 4907 12859
rect 4831 12793 4841 12849
rect 4897 12793 4907 12849
rect 4831 12745 4907 12793
rect 4831 12689 4841 12745
rect 4897 12689 4907 12745
rect 4831 12679 4907 12689
rect 5731 12849 5911 12859
rect 5731 12793 5741 12849
rect 5797 12793 5845 12849
rect 5901 12793 5911 12849
rect 6003 12840 6013 12896
rect 6069 12840 6117 12896
rect 6173 12840 6183 12896
rect 6003 12830 6183 12840
rect 6735 13000 6811 13010
rect 6735 12944 6745 13000
rect 6801 12944 6811 13000
rect 6735 12896 6811 12944
rect 6735 12840 6745 12896
rect 6801 12840 6811 12896
rect 6735 12830 6811 12840
rect 7375 13000 7451 13010
rect 7375 12944 7385 13000
rect 7441 12944 7451 13000
rect 7375 12896 7451 12944
rect 7375 12840 7385 12896
rect 7441 12840 7451 12896
rect 7375 12830 7451 12840
rect 8015 13000 8091 13010
rect 8015 12944 8025 13000
rect 8081 12944 8091 13000
rect 8015 12896 8091 12944
rect 8015 12840 8025 12896
rect 8081 12840 8091 12896
rect 8015 12830 8091 12840
rect 5731 12745 5911 12793
rect 5731 12689 5741 12745
rect 5797 12689 5845 12745
rect 5901 12689 5911 12745
rect 5731 12679 5911 12689
rect 3870 12457 3946 12467
rect 3870 12401 3880 12457
rect 3936 12401 3946 12457
rect 3870 12353 3946 12401
rect 3870 12297 3880 12353
rect 3936 12297 3946 12353
rect 3870 12287 3946 12297
rect 4510 12457 4586 12467
rect 4510 12401 4520 12457
rect 4576 12401 4586 12457
rect 4510 12353 4586 12401
rect 4510 12297 4520 12353
rect 4576 12297 4586 12353
rect 4510 12287 4586 12297
rect 5150 12457 5226 12467
rect 5150 12401 5160 12457
rect 5216 12401 5226 12457
rect 5150 12353 5226 12401
rect 5150 12297 5160 12353
rect 5216 12297 5226 12353
rect 5150 12287 5226 12297
rect 5741 12148 5901 12679
rect 6013 12467 6173 12830
rect 11371 12493 11551 12503
rect 6003 12457 6183 12467
rect 6003 12401 6013 12457
rect 6069 12401 6117 12457
rect 6173 12401 6183 12457
rect 6003 12353 6183 12401
rect 6003 12297 6013 12353
rect 6069 12297 6117 12353
rect 6173 12297 6183 12353
rect 6003 12287 6183 12297
rect 7055 12457 7131 12467
rect 7055 12401 7065 12457
rect 7121 12401 7131 12457
rect 7055 12353 7131 12401
rect 7055 12297 7065 12353
rect 7121 12297 7131 12353
rect 7055 12287 7131 12297
rect 7695 12457 7771 12467
rect 7695 12401 7705 12457
rect 7761 12401 7771 12457
rect 7695 12353 7771 12401
rect 7695 12297 7705 12353
rect 7761 12297 7771 12353
rect 11371 12437 11381 12493
rect 11437 12437 11485 12493
rect 11541 12437 11551 12493
rect 11371 12389 11551 12437
rect 11371 12333 11381 12389
rect 11437 12333 11485 12389
rect 11541 12333 11551 12389
rect 11371 12323 11551 12333
rect 7695 12287 7771 12297
rect 5731 12138 5911 12148
rect 5731 12082 5741 12138
rect 5797 12082 5845 12138
rect 5901 12082 5911 12138
rect 3161 12070 3341 12080
rect 3161 12014 3171 12070
rect 3227 12014 3275 12070
rect 3331 12014 3341 12070
rect 3161 11966 3341 12014
rect 3161 11910 3171 11966
rect 3227 11910 3275 11966
rect 3331 11910 3341 11966
rect 3161 11900 3341 11910
rect 3950 12070 4026 12080
rect 3950 12014 3960 12070
rect 4016 12014 4026 12070
rect 3950 11966 4026 12014
rect 5731 12034 5911 12082
rect 5731 11978 5741 12034
rect 5797 11978 5845 12034
rect 5901 11978 5911 12034
rect 5731 11968 5911 11978
rect 3950 11910 3960 11966
rect 4016 11910 4026 11966
rect 3950 11900 4026 11910
rect 2881 9812 3061 9822
rect 2881 9756 2891 9812
rect 2947 9756 2995 9812
rect 3051 9756 3061 9812
rect 2881 9708 3061 9756
rect 2881 9652 2891 9708
rect 2947 9652 2995 9708
rect 3051 9652 3061 9708
rect 2881 9642 3061 9652
rect 2624 9459 2700 9469
rect 2624 9403 2634 9459
rect 2690 9403 2700 9459
rect 2624 9355 2700 9403
rect 2624 9299 2634 9355
rect 2690 9299 2700 9355
rect 2624 9289 2700 9299
rect 2624 8129 2700 8139
rect 2624 8073 2634 8129
rect 2690 8073 2700 8129
rect 2624 8025 2700 8073
rect 2624 7969 2634 8025
rect 2690 7969 2700 8025
rect 2624 7959 2700 7969
rect 226 7585 406 7595
rect 226 7529 236 7585
rect 292 7529 340 7585
rect 396 7529 406 7585
rect 226 7481 406 7529
rect 226 7425 236 7481
rect 292 7425 340 7481
rect 396 7425 406 7481
rect 226 7415 406 7425
rect 1227 7585 1407 7595
rect 1227 7529 1237 7585
rect 1293 7529 1341 7585
rect 1397 7529 1407 7585
rect 1227 7481 1407 7529
rect 2891 7504 3051 9642
rect 3171 8692 3331 11900
rect 4190 11719 4266 11729
rect 4190 11663 4200 11719
rect 4256 11663 4266 11719
rect 4190 11615 4266 11663
rect 4190 11559 4200 11615
rect 4256 11559 4266 11615
rect 4190 11549 4266 11559
rect 4831 11719 4907 11729
rect 4831 11663 4841 11719
rect 4897 11663 4907 11719
rect 4831 11615 4907 11663
rect 4831 11559 4841 11615
rect 4897 11559 4907 11615
rect 4831 11549 4907 11559
rect 5741 11337 5901 11968
rect 6013 11729 6173 12287
rect 6735 12138 6811 12148
rect 6735 12082 6745 12138
rect 6801 12082 6811 12138
rect 6735 12034 6811 12082
rect 6735 11978 6745 12034
rect 6801 11978 6811 12034
rect 6735 11968 6811 11978
rect 7375 12138 7451 12148
rect 7375 12082 7385 12138
rect 7441 12082 7451 12138
rect 7375 12034 7451 12082
rect 7375 11978 7385 12034
rect 7441 11978 7451 12034
rect 7375 11968 7451 11978
rect 8015 12138 8091 12148
rect 8015 12082 8025 12138
rect 8081 12082 8091 12138
rect 8015 12034 8091 12082
rect 8015 11978 8025 12034
rect 8081 11978 8091 12034
rect 8015 11968 8091 11978
rect 6003 11719 6183 11729
rect 6003 11663 6013 11719
rect 6069 11663 6117 11719
rect 6173 11663 6183 11719
rect 6003 11615 6183 11663
rect 6003 11559 6013 11615
rect 6069 11559 6117 11615
rect 6173 11559 6183 11615
rect 6003 11511 6183 11559
rect 6003 11455 6013 11511
rect 6069 11455 6117 11511
rect 6173 11455 6183 11511
rect 6003 11445 6183 11455
rect 6735 11615 6811 11625
rect 6735 11559 6745 11615
rect 6801 11559 6811 11615
rect 6735 11511 6811 11559
rect 6735 11455 6745 11511
rect 6801 11455 6811 11511
rect 6735 11445 6811 11455
rect 7375 11615 7451 11625
rect 7375 11559 7385 11615
rect 7441 11559 7451 11615
rect 7375 11511 7451 11559
rect 7375 11455 7385 11511
rect 7441 11455 7451 11511
rect 7375 11445 7451 11455
rect 8015 11615 8091 11625
rect 8015 11559 8025 11615
rect 8081 11559 8091 11615
rect 8015 11511 8091 11559
rect 8015 11455 8025 11511
rect 8081 11455 8091 11511
rect 8015 11445 8091 11455
rect 5731 11327 5911 11337
rect 5731 11271 5741 11327
rect 5797 11271 5845 11327
rect 5901 11271 5911 11327
rect 3870 11223 3946 11233
rect 3870 11167 3880 11223
rect 3936 11167 3946 11223
rect 3870 11119 3946 11167
rect 3870 11063 3880 11119
rect 3936 11063 3946 11119
rect 3870 11053 3946 11063
rect 4510 11223 4586 11233
rect 4510 11167 4520 11223
rect 4576 11167 4586 11223
rect 4510 11119 4586 11167
rect 4510 11063 4520 11119
rect 4576 11063 4586 11119
rect 4510 11053 4586 11063
rect 5150 11223 5226 11233
rect 5150 11167 5160 11223
rect 5216 11167 5226 11223
rect 5150 11119 5226 11167
rect 5150 11063 5160 11119
rect 5216 11063 5226 11119
rect 5150 11053 5226 11063
rect 5731 11223 5911 11271
rect 5731 11167 5741 11223
rect 5797 11167 5845 11223
rect 5901 11167 5911 11223
rect 5731 11119 5911 11167
rect 5731 11063 5741 11119
rect 5797 11063 5845 11119
rect 5901 11063 5911 11119
rect 5731 11053 5911 11063
rect 5741 10806 5901 11053
rect 5731 10796 5911 10806
rect 5731 10740 5741 10796
rect 5797 10740 5845 10796
rect 5901 10740 5911 10796
rect 5731 10692 5911 10740
rect 5731 10636 5741 10692
rect 5797 10636 5845 10692
rect 5901 10636 5911 10692
rect 5731 10626 5911 10636
rect 4030 10325 4106 10335
rect 4030 10269 4040 10325
rect 4096 10269 4106 10325
rect 4030 10221 4106 10269
rect 4030 10165 4040 10221
rect 4096 10165 4106 10221
rect 4030 10155 4106 10165
rect 3950 9812 4026 9822
rect 3950 9756 3960 9812
rect 4016 9756 4026 9812
rect 3950 9708 4026 9756
rect 3950 9652 3960 9708
rect 4016 9652 4026 9708
rect 3950 9640 4026 9652
rect 5741 9573 5901 10626
rect 6013 10435 6173 11445
rect 11381 11385 11541 12323
rect 11371 11375 11551 11385
rect 7055 11327 7131 11337
rect 7055 11271 7065 11327
rect 7121 11271 7131 11327
rect 7055 11223 7131 11271
rect 7055 11167 7065 11223
rect 7121 11167 7131 11223
rect 7055 11157 7131 11167
rect 7695 11327 7771 11337
rect 7695 11271 7705 11327
rect 7761 11271 7771 11327
rect 7695 11223 7771 11271
rect 7695 11167 7705 11223
rect 7761 11167 7771 11223
rect 11371 11319 11381 11375
rect 11437 11319 11485 11375
rect 11541 11319 11551 11375
rect 11371 11271 11551 11319
rect 11371 11215 11381 11271
rect 11437 11215 11485 11271
rect 11541 11215 11551 11271
rect 11371 11205 11551 11215
rect 7695 11157 7771 11167
rect 8970 10796 9046 10806
rect 8970 10740 8980 10796
rect 9036 10740 9046 10796
rect 8970 10692 9046 10740
rect 8970 10636 8980 10692
rect 9036 10636 9046 10692
rect 8970 10626 9046 10636
rect 9866 10796 9942 10806
rect 9866 10740 9876 10796
rect 9932 10740 9942 10796
rect 9866 10692 9942 10740
rect 9866 10636 9876 10692
rect 9932 10636 9942 10692
rect 9866 10626 9942 10636
rect 10762 10796 10838 10806
rect 10762 10740 10772 10796
rect 10828 10740 10838 10796
rect 10762 10692 10838 10740
rect 10762 10636 10772 10692
rect 10828 10636 10838 10692
rect 10762 10626 10838 10636
rect 6003 10425 6183 10435
rect 6003 10369 6013 10425
rect 6069 10369 6117 10425
rect 6173 10369 6183 10425
rect 6003 10321 6183 10369
rect 6003 10265 6013 10321
rect 6069 10265 6117 10321
rect 6173 10265 6183 10321
rect 6003 10255 6183 10265
rect 9418 10425 9494 10435
rect 9418 10369 9428 10425
rect 9484 10369 9494 10425
rect 9418 10321 9494 10369
rect 9418 10265 9428 10321
rect 9484 10265 9494 10321
rect 9418 10255 9494 10265
rect 10314 10425 10390 10435
rect 10314 10369 10324 10425
rect 10380 10369 10390 10425
rect 10314 10321 10390 10369
rect 10314 10265 10324 10321
rect 10380 10265 10390 10321
rect 10314 10255 10390 10265
rect 10602 10425 10678 10435
rect 10602 10369 10612 10425
rect 10668 10369 10678 10425
rect 10602 10321 10678 10369
rect 10602 10265 10612 10321
rect 10668 10265 10678 10321
rect 10602 10255 10678 10265
rect 6013 9974 6173 10255
rect 6003 9964 6183 9974
rect 6003 9908 6013 9964
rect 6069 9908 6117 9964
rect 6173 9908 6183 9964
rect 6003 9860 6183 9908
rect 6003 9804 6013 9860
rect 6069 9804 6117 9860
rect 6173 9804 6183 9860
rect 6003 9794 6183 9804
rect 7055 9964 7131 9974
rect 7055 9908 7065 9964
rect 7121 9908 7131 9964
rect 7055 9860 7131 9908
rect 7055 9804 7065 9860
rect 7121 9804 7131 9860
rect 7055 9794 7131 9804
rect 7695 9964 7771 9974
rect 7695 9908 7705 9964
rect 7761 9908 7771 9964
rect 7695 9860 7771 9908
rect 7695 9804 7705 9860
rect 7761 9804 7771 9860
rect 7695 9794 7771 9804
rect 5731 9563 5911 9573
rect 5731 9507 5741 9563
rect 5797 9507 5845 9563
rect 5901 9507 5911 9563
rect 4030 9459 4106 9469
rect 4030 9403 4040 9459
rect 4096 9403 4106 9459
rect 4030 9355 4106 9403
rect 4030 9299 4040 9355
rect 4096 9299 4106 9355
rect 4030 9289 4106 9299
rect 4190 9459 4266 9469
rect 4190 9403 4200 9459
rect 4256 9403 4266 9459
rect 4190 9355 4266 9403
rect 4190 9299 4200 9355
rect 4256 9299 4266 9355
rect 4190 9289 4266 9299
rect 4831 9459 4907 9469
rect 4831 9403 4841 9459
rect 4897 9403 4907 9459
rect 4831 9355 4907 9403
rect 4831 9299 4841 9355
rect 4897 9299 4907 9355
rect 4831 9289 4907 9299
rect 5731 9459 5911 9507
rect 5731 9403 5741 9459
rect 5797 9403 5845 9459
rect 5901 9403 5911 9459
rect 5731 9355 5911 9403
rect 5731 9299 5741 9355
rect 5797 9299 5845 9355
rect 5901 9299 5911 9355
rect 5731 9289 5911 9299
rect 3870 8963 3946 8973
rect 3870 8907 3880 8963
rect 3936 8907 3946 8963
rect 3870 8859 3946 8907
rect 3870 8803 3880 8859
rect 3936 8803 3946 8859
rect 3870 8793 3946 8803
rect 4510 8963 4586 8973
rect 4510 8907 4520 8963
rect 4576 8907 4586 8963
rect 4510 8859 4586 8907
rect 4510 8803 4520 8859
rect 4576 8803 4586 8859
rect 4510 8793 4586 8803
rect 5150 8963 5226 8973
rect 5150 8907 5160 8963
rect 5216 8907 5226 8963
rect 5150 8859 5226 8907
rect 5150 8803 5160 8859
rect 5216 8803 5226 8859
rect 5150 8793 5226 8803
rect 5741 8700 5901 9289
rect 6013 8973 6173 9794
rect 11381 9773 11541 11205
rect 11649 10965 11809 13289
rect 17641 11505 17716 13351
rect 19065 13407 19141 13417
rect 19065 13351 19075 13407
rect 19131 13351 19141 13407
rect 19065 13341 19141 13351
rect 20185 13407 20261 13417
rect 20185 13351 20195 13407
rect 20251 13351 20261 13407
rect 20185 13341 20261 13351
rect 24217 13407 24293 13417
rect 24217 13351 24227 13407
rect 24283 13351 24293 13407
rect 24217 13341 24293 13351
rect 25337 13407 25413 13417
rect 25337 13351 25347 13407
rect 25403 13351 25413 13407
rect 25337 13341 25413 13351
rect 26762 13407 26837 13417
rect 26762 13351 26771 13407
rect 26828 13351 26837 13407
rect 22097 13270 22381 13280
rect 22097 13214 22107 13270
rect 22163 13214 22211 13270
rect 22267 13214 22315 13270
rect 22371 13214 22381 13270
rect 19305 13166 19381 13176
rect 19305 13110 19315 13166
rect 19371 13110 19381 13166
rect 19305 13062 19381 13110
rect 19305 13006 19315 13062
rect 19371 13006 19381 13062
rect 19305 12996 19381 13006
rect 19945 13166 20021 13176
rect 19945 13110 19955 13166
rect 20011 13110 20021 13166
rect 19945 13062 20021 13110
rect 19945 13006 19955 13062
rect 20011 13006 20021 13062
rect 19945 12996 20021 13006
rect 22097 13166 22381 13214
rect 22097 13110 22107 13166
rect 22163 13110 22211 13166
rect 22267 13110 22315 13166
rect 22371 13110 22381 13166
rect 22097 13062 22381 13110
rect 22097 13006 22107 13062
rect 22163 13006 22211 13062
rect 22267 13006 22315 13062
rect 22371 13006 22381 13062
rect 21448 12876 21732 12886
rect 21448 12820 21458 12876
rect 21514 12820 21562 12876
rect 21618 12820 21666 12876
rect 21722 12820 21732 12876
rect 18985 12772 19061 12782
rect 18985 12716 18995 12772
rect 19051 12716 19061 12772
rect 18985 12668 19061 12716
rect 18985 12612 18995 12668
rect 19051 12612 19061 12668
rect 18985 12602 19061 12612
rect 19145 12770 19221 12782
rect 19145 12718 19157 12770
rect 19209 12718 19221 12770
rect 19145 12666 19221 12718
rect 19145 12614 19157 12666
rect 19209 12614 19221 12666
rect 19145 12602 19221 12614
rect 19465 12770 19541 12782
rect 19465 12718 19477 12770
rect 19529 12718 19541 12770
rect 19465 12666 19541 12718
rect 19465 12614 19477 12666
rect 19529 12614 19541 12666
rect 19465 12602 19541 12614
rect 19625 12772 19701 12782
rect 19625 12716 19635 12772
rect 19691 12716 19701 12772
rect 19625 12668 19701 12716
rect 19625 12612 19635 12668
rect 19691 12612 19701 12668
rect 19625 12602 19701 12612
rect 19785 12770 19861 12782
rect 19785 12718 19797 12770
rect 19849 12718 19861 12770
rect 19785 12666 19861 12718
rect 19785 12614 19797 12666
rect 19849 12614 19861 12666
rect 19785 12602 19861 12614
rect 20105 12770 20181 12782
rect 20105 12718 20117 12770
rect 20169 12718 20181 12770
rect 20105 12666 20181 12718
rect 20105 12614 20117 12666
rect 20169 12614 20181 12666
rect 20105 12602 20181 12614
rect 20265 12772 20341 12782
rect 20265 12716 20275 12772
rect 20331 12716 20341 12772
rect 20265 12668 20341 12716
rect 20265 12612 20275 12668
rect 20331 12612 20341 12668
rect 20265 12602 20341 12612
rect 21448 12772 21732 12820
rect 21448 12716 21458 12772
rect 21514 12716 21562 12772
rect 21618 12716 21666 12772
rect 21722 12716 21732 12772
rect 21448 12668 21732 12716
rect 21448 12612 21458 12668
rect 21514 12612 21562 12668
rect 21618 12612 21666 12668
rect 21722 12612 21732 12668
rect 17641 11449 17651 11505
rect 17707 11449 17716 11505
rect 12800 11375 12876 11385
rect 12800 11319 12810 11375
rect 12866 11319 12876 11375
rect 12800 11271 12876 11319
rect 12800 11215 12810 11271
rect 12866 11215 12876 11271
rect 12800 11205 12876 11215
rect 13696 11375 13772 11385
rect 13696 11319 13706 11375
rect 13762 11319 13772 11375
rect 13696 11271 13772 11319
rect 13696 11215 13706 11271
rect 13762 11215 13772 11271
rect 13696 11205 13772 11215
rect 13984 11375 14060 11385
rect 13984 11319 13994 11375
rect 14050 11319 14060 11375
rect 13984 11271 14060 11319
rect 13984 11215 13994 11271
rect 14050 11215 14060 11271
rect 13984 11205 14060 11215
rect 15146 11375 15222 11385
rect 15146 11319 15156 11375
rect 15212 11319 15222 11375
rect 15146 11271 15222 11319
rect 15146 11215 15156 11271
rect 15212 11215 15222 11271
rect 15146 11205 15222 11215
rect 15786 11375 15862 11385
rect 15786 11319 15796 11375
rect 15852 11319 15862 11375
rect 15786 11271 15862 11319
rect 15786 11215 15796 11271
rect 15852 11215 15862 11271
rect 15786 11205 15862 11215
rect 16426 11375 16502 11385
rect 16426 11319 16436 11375
rect 16492 11319 16502 11375
rect 16426 11271 16502 11319
rect 16426 11215 16436 11271
rect 16492 11215 16502 11271
rect 16426 11205 16502 11215
rect 17365 11375 17545 11385
rect 17365 11319 17375 11375
rect 17431 11319 17479 11375
rect 17535 11319 17545 11375
rect 17365 11271 17545 11319
rect 17365 11215 17375 11271
rect 17431 11215 17479 11271
rect 17535 11215 17545 11271
rect 17365 11205 17545 11215
rect 11639 10955 11819 10965
rect 11639 10899 11649 10955
rect 11705 10899 11753 10955
rect 11809 10899 11819 10955
rect 11639 10851 11819 10899
rect 11639 10795 11649 10851
rect 11705 10795 11753 10851
rect 11809 10795 11819 10851
rect 11639 10785 11819 10795
rect 12352 10955 12428 10965
rect 12352 10899 12362 10955
rect 12418 10899 12428 10955
rect 12352 10851 12428 10899
rect 12352 10795 12362 10851
rect 12418 10795 12428 10851
rect 12352 10785 12428 10795
rect 13248 10955 13324 10965
rect 13248 10899 13258 10955
rect 13314 10899 13324 10955
rect 13248 10851 13324 10899
rect 13248 10795 13258 10851
rect 13314 10795 13324 10851
rect 13248 10785 13324 10795
rect 14144 10955 14220 10965
rect 14144 10899 14154 10955
rect 14210 10899 14220 10955
rect 14144 10851 14220 10899
rect 14144 10795 14154 10851
rect 14210 10795 14220 10851
rect 14144 10785 14220 10795
rect 15466 10955 15542 10965
rect 15466 10899 15476 10955
rect 15532 10899 15542 10955
rect 15466 10851 15542 10899
rect 15466 10795 15476 10851
rect 15532 10795 15542 10851
rect 15466 10785 15542 10795
rect 16106 10955 16182 10965
rect 16106 10899 16116 10955
rect 16172 10899 16182 10955
rect 16106 10851 16182 10899
rect 16106 10795 16116 10851
rect 16172 10795 16182 10851
rect 16106 10785 16182 10795
rect 17103 10955 17283 10965
rect 17103 10899 17113 10955
rect 17169 10899 17217 10955
rect 17273 10899 17283 10955
rect 17103 10851 17283 10899
rect 17103 10795 17113 10851
rect 17169 10795 17217 10851
rect 17273 10795 17283 10851
rect 17103 10785 17283 10795
rect 11649 10435 11809 10785
rect 11639 10425 11819 10435
rect 11639 10369 11649 10425
rect 11705 10369 11753 10425
rect 11809 10369 11819 10425
rect 11639 10321 11819 10369
rect 11639 10265 11649 10321
rect 11705 10265 11753 10321
rect 11809 10265 11819 10321
rect 11639 10217 11819 10265
rect 11639 10161 11649 10217
rect 11705 10161 11753 10217
rect 11809 10161 11819 10217
rect 11639 10151 11819 10161
rect 12800 10321 12876 10331
rect 12800 10265 12810 10321
rect 12866 10265 12876 10321
rect 12800 10217 12876 10265
rect 12800 10161 12810 10217
rect 12866 10161 12876 10217
rect 12800 10151 12876 10161
rect 13696 10321 13772 10331
rect 13696 10265 13706 10321
rect 13762 10265 13772 10321
rect 17113 10305 17273 10785
rect 13696 10217 13772 10265
rect 13696 10161 13706 10217
rect 13762 10161 13772 10217
rect 13696 10151 13772 10161
rect 13984 10295 14060 10305
rect 13984 10239 13994 10295
rect 14050 10239 14060 10295
rect 13984 10191 14060 10239
rect 10602 9763 10678 9773
rect 10602 9707 10612 9763
rect 10668 9707 10678 9763
rect 10602 9659 10678 9707
rect 10602 9603 10612 9659
rect 10668 9603 10678 9659
rect 10602 9593 10678 9603
rect 11371 9763 11551 9773
rect 11371 9707 11381 9763
rect 11437 9707 11485 9763
rect 11541 9707 11551 9763
rect 11371 9659 11551 9707
rect 11371 9603 11381 9659
rect 11437 9603 11485 9659
rect 11541 9603 11551 9659
rect 11371 9593 11551 9603
rect 6735 9563 6811 9573
rect 6735 9507 6745 9563
rect 6801 9507 6811 9563
rect 6735 9459 6811 9507
rect 6735 9403 6745 9459
rect 6801 9403 6811 9459
rect 6735 9393 6811 9403
rect 7375 9563 7451 9573
rect 7375 9507 7385 9563
rect 7441 9507 7451 9563
rect 7375 9459 7451 9507
rect 7375 9403 7385 9459
rect 7441 9403 7451 9459
rect 7375 9393 7451 9403
rect 8015 9563 8091 9573
rect 8015 9507 8025 9563
rect 8081 9507 8091 9563
rect 8015 9459 8091 9507
rect 8015 9403 8025 9459
rect 8081 9403 8091 9459
rect 8015 9393 8091 9403
rect 9418 9563 9494 9573
rect 9418 9507 9428 9563
rect 9484 9507 9494 9563
rect 9418 9459 9494 9507
rect 9418 9403 9428 9459
rect 9484 9403 9494 9459
rect 9418 9393 9494 9403
rect 10314 9563 10390 9573
rect 10314 9507 10324 9563
rect 10380 9507 10390 9563
rect 10314 9459 10390 9507
rect 10314 9403 10324 9459
rect 10380 9403 10390 9459
rect 10314 9393 10390 9403
rect 11381 9285 11541 9593
rect 11371 9275 11551 9285
rect 11371 9219 11381 9275
rect 11437 9219 11485 9275
rect 11541 9219 11551 9275
rect 11371 9171 11551 9219
rect 11371 9115 11381 9171
rect 11437 9115 11485 9171
rect 11541 9115 11551 9171
rect 11371 9105 11551 9115
rect 6003 8963 6183 8973
rect 6003 8907 6013 8963
rect 6069 8907 6117 8963
rect 6173 8907 6183 8963
rect 6003 8859 6183 8907
rect 6003 8803 6013 8859
rect 6069 8803 6117 8859
rect 6173 8803 6183 8859
rect 6003 8793 6183 8803
rect 6735 8963 6811 8973
rect 6735 8907 6745 8963
rect 6801 8907 6811 8963
rect 6735 8859 6811 8907
rect 6735 8803 6745 8859
rect 6801 8803 6811 8859
rect 6735 8793 6811 8803
rect 7375 8963 7451 8973
rect 7375 8907 7385 8963
rect 7441 8907 7451 8963
rect 7375 8859 7451 8907
rect 7375 8803 7385 8859
rect 7441 8803 7451 8859
rect 7375 8793 7451 8803
rect 8015 8963 8091 8973
rect 8015 8907 8025 8963
rect 8081 8907 8091 8963
rect 8015 8859 8091 8907
rect 8015 8803 8025 8859
rect 8081 8803 8091 8859
rect 8015 8793 8091 8803
rect 8970 8963 9046 8973
rect 8970 8907 8980 8963
rect 9036 8907 9046 8963
rect 8970 8859 9046 8907
rect 8970 8803 8980 8859
rect 9036 8803 9046 8859
rect 8970 8793 9046 8803
rect 9866 8963 9942 8973
rect 9866 8907 9876 8963
rect 9932 8907 9942 8963
rect 9866 8859 9942 8907
rect 9866 8803 9876 8859
rect 9932 8803 9942 8859
rect 9866 8793 9942 8803
rect 10762 8963 10838 8973
rect 10762 8907 10772 8963
rect 10828 8907 10838 8963
rect 10762 8859 10838 8907
rect 10762 8803 10772 8859
rect 10828 8803 10838 8859
rect 10762 8793 10838 8803
rect 3161 8682 3341 8692
rect 3161 8626 3171 8682
rect 3227 8626 3275 8682
rect 3331 8626 3341 8682
rect 3161 8578 3341 8626
rect 3161 8522 3171 8578
rect 3227 8522 3275 8578
rect 3331 8522 3341 8578
rect 3161 8512 3341 8522
rect 3950 8682 4026 8692
rect 3950 8626 3960 8682
rect 4016 8626 4026 8682
rect 3950 8578 4026 8626
rect 3950 8522 3960 8578
rect 4016 8522 4026 8578
rect 3950 8512 4026 8522
rect 5731 8690 5911 8700
rect 5731 8634 5741 8690
rect 5797 8634 5845 8690
rect 5901 8634 5911 8690
rect 5731 8586 5911 8634
rect 5731 8530 5741 8586
rect 5797 8530 5845 8586
rect 5901 8530 5911 8586
rect 5731 8520 5911 8530
rect 4190 8329 4266 8339
rect 4190 8273 4200 8329
rect 4256 8273 4266 8329
rect 4190 8225 4266 8273
rect 4190 8169 4200 8225
rect 4256 8169 4266 8225
rect 4190 8159 4266 8169
rect 4831 8329 4907 8339
rect 4831 8273 4841 8329
rect 4897 8273 4907 8329
rect 4831 8225 4907 8273
rect 4831 8169 4841 8225
rect 4897 8169 4907 8225
rect 4831 8159 4907 8169
rect 4030 8129 4106 8139
rect 4030 8073 4040 8129
rect 4096 8073 4106 8129
rect 4030 8025 4106 8073
rect 4030 7969 4040 8025
rect 4096 7969 4106 8025
rect 4030 7959 4106 7969
rect 5741 7843 5901 8520
rect 6013 8339 6173 8793
rect 10474 8705 10550 8715
rect 7055 8690 7131 8700
rect 7055 8634 7065 8690
rect 7121 8634 7131 8690
rect 7055 8586 7131 8634
rect 7055 8530 7065 8586
rect 7121 8530 7131 8586
rect 7055 8520 7131 8530
rect 7695 8690 7771 8700
rect 7695 8634 7705 8690
rect 7761 8634 7771 8690
rect 7695 8586 7771 8634
rect 7695 8530 7705 8586
rect 7761 8530 7771 8586
rect 10474 8649 10484 8705
rect 10540 8649 10550 8705
rect 10474 8601 10550 8649
rect 10474 8545 10484 8601
rect 10540 8545 10550 8601
rect 10474 8535 10550 8545
rect 7695 8520 7771 8530
rect 7989 8466 8065 8476
rect 7989 8410 7999 8466
rect 8055 8410 8065 8466
rect 7989 8362 8065 8410
rect 6003 8329 6183 8339
rect 6003 8273 6013 8329
rect 6069 8273 6117 8329
rect 6173 8273 6183 8329
rect 7989 8306 7999 8362
rect 8055 8306 8065 8362
rect 7989 8296 8065 8306
rect 8275 8466 8455 8476
rect 8275 8410 8285 8466
rect 8341 8410 8389 8466
rect 8445 8410 8455 8466
rect 8275 8362 8455 8410
rect 8275 8306 8285 8362
rect 8341 8306 8389 8362
rect 8445 8306 8455 8362
rect 8275 8296 8455 8306
rect 10722 8455 10798 8465
rect 10722 8399 10732 8455
rect 10788 8399 10798 8455
rect 10722 8351 10798 8399
rect 6003 8225 6183 8273
rect 6003 8169 6013 8225
rect 6069 8169 6117 8225
rect 6173 8169 6183 8225
rect 6003 8121 6183 8169
rect 6003 8065 6013 8121
rect 6069 8065 6117 8121
rect 6173 8065 6183 8121
rect 6003 8055 6183 8065
rect 7055 8225 7131 8235
rect 7055 8169 7065 8225
rect 7121 8169 7131 8225
rect 7055 8121 7131 8169
rect 7055 8065 7065 8121
rect 7121 8065 7131 8121
rect 7055 8055 7131 8065
rect 7695 8225 7771 8235
rect 7695 8169 7705 8225
rect 7761 8169 7771 8225
rect 7695 8121 7771 8169
rect 7695 8065 7705 8121
rect 7761 8065 7771 8121
rect 7695 8055 7771 8065
rect 3870 7833 3946 7843
rect 3870 7777 3880 7833
rect 3936 7777 3946 7833
rect 3870 7729 3946 7777
rect 3870 7673 3880 7729
rect 3936 7673 3946 7729
rect 3870 7663 3946 7673
rect 4510 7833 4586 7843
rect 4510 7777 4520 7833
rect 4576 7777 4586 7833
rect 4510 7729 4586 7777
rect 4510 7673 4520 7729
rect 4576 7673 4586 7729
rect 4510 7663 4586 7673
rect 5150 7833 5226 7843
rect 5150 7777 5160 7833
rect 5216 7777 5226 7833
rect 5150 7729 5226 7777
rect 5150 7673 5160 7729
rect 5216 7673 5226 7729
rect 5150 7663 5226 7673
rect 5731 7833 5911 7843
rect 5731 7777 5741 7833
rect 5797 7777 5845 7833
rect 5901 7777 5911 7833
rect 5731 7729 5911 7777
rect 5731 7673 5741 7729
rect 5797 7673 5845 7729
rect 5901 7673 5911 7729
rect 5731 7663 5911 7673
rect 6735 7833 6811 7843
rect 6735 7777 6745 7833
rect 6801 7777 6811 7833
rect 6735 7729 6811 7777
rect 6735 7673 6745 7729
rect 6801 7673 6811 7729
rect 6735 7663 6811 7673
rect 7375 7833 7451 7843
rect 7375 7777 7385 7833
rect 7441 7777 7451 7833
rect 7375 7729 7451 7777
rect 7375 7673 7385 7729
rect 7441 7673 7451 7729
rect 7375 7663 7451 7673
rect 8015 7833 8091 7843
rect 8015 7777 8025 7833
rect 8081 7777 8091 7833
rect 8015 7729 8091 7777
rect 8015 7673 8025 7729
rect 8081 7673 8091 7729
rect 8015 7663 8091 7673
rect 1227 7425 1237 7481
rect 1293 7425 1341 7481
rect 1397 7425 1407 7481
rect 1227 7415 1407 7425
rect 2881 7494 3061 7504
rect 2881 7438 2891 7494
rect 2947 7438 2995 7494
rect 3051 7438 3061 7494
rect 1237 3171 1397 7415
rect 2881 7390 3061 7438
rect 2881 7334 2891 7390
rect 2947 7334 2995 7390
rect 3051 7334 3061 7390
rect 2881 7324 3061 7334
rect 4110 7494 4186 7504
rect 4110 7438 4120 7494
rect 4176 7438 4186 7494
rect 4110 7390 4186 7438
rect 4110 7334 4120 7390
rect 4176 7334 4186 7390
rect 4110 7324 4186 7334
rect 6867 7379 7047 7391
rect 6867 7327 6879 7379
rect 6931 7327 6983 7379
rect 7035 7327 7047 7379
rect 6867 7275 7047 7327
rect 6867 7223 6879 7275
rect 6931 7223 6983 7275
rect 7035 7223 7047 7275
rect 6867 7211 7047 7223
rect 6879 6185 7039 7211
rect 8285 6421 8445 8296
rect 10722 8295 10732 8351
rect 10788 8295 10798 8351
rect 10722 8285 10798 8295
rect 10918 8455 11098 8465
rect 10918 8399 10928 8455
rect 10984 8399 11032 8455
rect 11088 8399 11098 8455
rect 10918 8351 11098 8399
rect 10918 8295 10928 8351
rect 10984 8295 11032 8351
rect 11088 8295 11098 8351
rect 10918 8285 11098 8295
rect 9418 8225 9494 8235
rect 9418 8169 9428 8225
rect 9484 8169 9494 8225
rect 9418 8121 9494 8169
rect 9418 8065 9428 8121
rect 9484 8065 9494 8121
rect 9418 8055 9494 8065
rect 10314 8225 10390 8235
rect 10314 8169 10324 8225
rect 10380 8169 10390 8225
rect 10314 8121 10390 8169
rect 10314 8065 10324 8121
rect 10380 8065 10390 8121
rect 10314 8055 10390 8065
rect 10474 8225 10550 8235
rect 10474 8169 10484 8225
rect 10540 8169 10550 8225
rect 10474 8121 10550 8169
rect 10474 8065 10484 8121
rect 10540 8065 10550 8121
rect 10474 8055 10550 8065
rect 8970 7833 9046 7843
rect 8970 7777 8980 7833
rect 9036 7777 9046 7833
rect 8970 7729 9046 7777
rect 8970 7673 8980 7729
rect 9036 7673 9046 7729
rect 8970 7663 9046 7673
rect 9866 7833 9942 7843
rect 9866 7777 9876 7833
rect 9932 7777 9942 7833
rect 9866 7729 9942 7777
rect 9866 7673 9876 7729
rect 9932 7673 9942 7729
rect 9866 7663 9942 7673
rect 10762 7833 10838 7843
rect 10762 7777 10772 7833
rect 10828 7777 10838 7833
rect 10762 7729 10838 7777
rect 10762 7673 10772 7729
rect 10828 7673 10838 7729
rect 10762 7663 10838 7673
rect 9969 7379 10149 7391
rect 9969 7327 9981 7379
rect 10033 7327 10085 7379
rect 10137 7327 10149 7379
rect 9969 7275 10149 7327
rect 9969 7223 9981 7275
rect 10033 7223 10085 7275
rect 10137 7223 10149 7275
rect 9969 7211 10149 7223
rect 7382 6411 7562 6421
rect 7382 6355 7392 6411
rect 7448 6355 7496 6411
rect 7552 6355 7562 6411
rect 7382 6307 7562 6355
rect 7382 6251 7392 6307
rect 7448 6251 7496 6307
rect 7552 6251 7562 6307
rect 7382 6241 7562 6251
rect 8275 6411 8455 6421
rect 8275 6355 8285 6411
rect 8341 6355 8389 6411
rect 8445 6355 8455 6411
rect 8275 6307 8455 6355
rect 8275 6251 8285 6307
rect 8341 6251 8389 6307
rect 8445 6251 8455 6307
rect 8275 6241 8455 6251
rect 6867 6173 7047 6185
rect 6867 6121 6879 6173
rect 6931 6121 6983 6173
rect 7035 6121 7047 6173
rect 6867 6069 7047 6121
rect 6867 6017 6879 6069
rect 6931 6017 6983 6069
rect 7035 6017 7047 6069
rect 6867 6005 7047 6017
rect 5144 5459 5324 5471
rect 5144 5407 5156 5459
rect 5208 5407 5260 5459
rect 5312 5407 5324 5459
rect 5144 5355 5324 5407
rect 2175 5308 2355 5320
rect 2175 5256 2187 5308
rect 2239 5256 2291 5308
rect 2343 5256 2355 5308
rect 5144 5303 5156 5355
rect 5208 5303 5260 5355
rect 5312 5303 5324 5355
rect 5144 5291 5324 5303
rect 2175 5204 2355 5256
rect 2175 5152 2187 5204
rect 2239 5152 2291 5204
rect 2343 5152 2355 5204
rect 2175 5140 2355 5152
rect 3047 5175 3227 5185
rect 2185 4568 2345 5140
rect 3047 5119 3057 5175
rect 3113 5119 3161 5175
rect 3217 5119 3227 5175
rect 3047 5071 3227 5119
rect 3047 5015 3057 5071
rect 3113 5015 3161 5071
rect 3217 5015 3227 5071
rect 3047 5005 3227 5015
rect 2175 4556 2355 4568
rect 2175 4504 2187 4556
rect 2239 4504 2291 4556
rect 2343 4504 2355 4556
rect 2175 4492 2355 4504
rect 2715 4421 2791 4431
rect 2715 4365 2725 4421
rect 2781 4365 2791 4421
rect 2715 4317 2791 4365
rect 2715 4261 2725 4317
rect 2781 4261 2791 4317
rect 2715 4251 2791 4261
rect 3109 3171 3165 5005
rect 4011 4131 4087 4141
rect 4011 4075 4021 4131
rect 4077 4075 4087 4131
rect 4011 4027 4087 4075
rect 4011 3971 4021 4027
rect 4077 3971 4087 4027
rect 4011 3961 4087 3971
rect 3579 3807 3655 3817
rect 3579 3751 3589 3807
rect 3645 3751 3655 3807
rect 3579 3703 3655 3751
rect 3579 3647 3589 3703
rect 3645 3647 3655 3703
rect 3579 3637 3655 3647
rect 3419 3405 3599 3415
rect 3419 3349 3429 3405
rect 3485 3349 3533 3405
rect 3589 3349 3599 3405
rect 3419 3301 3599 3349
rect 3419 3245 3429 3301
rect 3485 3245 3533 3301
rect 3589 3245 3599 3301
rect 3419 3235 3599 3245
rect 3429 3171 3485 3235
rect 1227 3161 1407 3171
rect 1227 3105 1237 3161
rect 1293 3105 1341 3161
rect 1397 3105 1407 3161
rect 1227 3057 1407 3105
rect 1227 3001 1237 3057
rect 1293 3001 1341 3057
rect 1397 3001 1407 3057
rect 1227 2991 1407 3001
rect 2725 3161 2801 3171
rect 2725 3105 2735 3161
rect 2791 3105 2801 3161
rect 2725 3057 2801 3105
rect 2725 3001 2735 3057
rect 2791 3001 2801 3057
rect 2725 2991 2801 3001
rect 3099 3159 3175 3171
rect 3099 3107 3111 3159
rect 3163 3107 3175 3159
rect 3099 3055 3175 3107
rect 3099 3003 3111 3055
rect 3163 3003 3175 3055
rect 3099 2991 3175 3003
rect 3419 3159 3495 3171
rect 3419 3107 3431 3159
rect 3483 3107 3495 3159
rect 3419 3055 3495 3107
rect 3419 3003 3431 3055
rect 3483 3003 3495 3055
rect 3419 2991 3495 3003
rect 5154 2555 5314 5291
rect 5620 4421 5800 4431
rect 5620 4365 5630 4421
rect 5686 4365 5734 4421
rect 5790 4365 5800 4421
rect 5620 4317 5800 4365
rect 5620 4261 5630 4317
rect 5686 4261 5734 4317
rect 5790 4261 5800 4317
rect 5620 4251 5800 4261
rect 5384 3807 5564 3817
rect 5384 3751 5394 3807
rect 5450 3751 5498 3807
rect 5554 3751 5564 3807
rect 5384 3703 5564 3751
rect 5384 3647 5394 3703
rect 5450 3647 5498 3703
rect 5554 3647 5564 3703
rect 5384 3637 5564 3647
rect 3923 2545 3999 2555
rect 3923 2489 3933 2545
rect 3989 2489 3999 2545
rect 3923 2441 3999 2489
rect 3923 2385 3933 2441
rect 3989 2385 3999 2441
rect 3923 2375 3999 2385
rect 5144 2545 5324 2555
rect 5144 2489 5154 2545
rect 5210 2489 5258 2545
rect 5314 2489 5324 2545
rect 5144 2441 5324 2489
rect 5144 2385 5154 2441
rect 5210 2385 5258 2441
rect 5314 2385 5324 2441
rect 5394 2412 5554 3637
rect 5144 2375 5324 2385
rect 5384 2402 5564 2412
rect -8069 2137 -1434 2259
rect -8178 2103 -1434 2137
rect -8178 2047 -8163 2103
rect -8107 2047 -8053 2103
rect -7997 2047 -1434 2103
rect -8178 1993 -1434 2047
rect 5154 2026 5314 2375
rect 5384 2346 5394 2402
rect 5450 2346 5498 2402
rect 5554 2346 5564 2402
rect 5384 2298 5564 2346
rect 5384 2242 5394 2298
rect 5450 2242 5498 2298
rect 5554 2242 5564 2298
rect 5384 2232 5564 2242
rect -8178 1937 -8163 1993
rect -8107 1937 -8053 1993
rect -7997 1978 -1434 1993
rect 5144 2016 5324 2026
rect -7997 1947 -6931 1978
rect 5144 1960 5154 2016
rect 5210 1960 5258 2016
rect 5314 1960 5324 2016
rect -7997 1937 -7966 1947
rect -8178 1925 -7966 1937
rect 5144 1912 5324 1960
rect 5144 1856 5154 1912
rect 5210 1856 5258 1912
rect 5314 1856 5324 1912
rect 5144 1846 5324 1856
rect 3971 1775 4047 1785
rect 3971 1719 3981 1775
rect 4037 1719 4047 1775
rect 3971 1671 4047 1719
rect 3971 1615 3981 1671
rect 4037 1615 4047 1671
rect 3971 1605 4047 1615
rect 5154 567 5314 1846
rect 5630 887 5790 4251
rect 6093 4131 6273 4141
rect 6093 4075 6103 4131
rect 6159 4075 6207 4131
rect 6263 4075 6273 4131
rect 6093 4027 6273 4075
rect 6093 3971 6103 4027
rect 6159 3971 6207 4027
rect 6263 3971 6273 4027
rect 6093 3961 6273 3971
rect 6544 4103 6724 4113
rect 6544 4047 6554 4103
rect 6610 4047 6658 4103
rect 6714 4047 6724 4103
rect 6544 3999 6724 4047
rect 5851 3613 6031 3623
rect 5851 3557 5861 3613
rect 5917 3557 5965 3613
rect 6021 3557 6031 3613
rect 5851 3509 6031 3557
rect 5851 3453 5861 3509
rect 5917 3453 5965 3509
rect 6021 3453 6031 3509
rect 5851 3405 6031 3453
rect 5851 3349 5861 3405
rect 5917 3349 5965 3405
rect 6021 3349 6031 3405
rect 5851 3301 6031 3349
rect 5851 3245 5861 3301
rect 5917 3245 5965 3301
rect 6021 3245 6031 3301
rect 5851 3235 6031 3245
rect 6103 2899 6263 3961
rect 6544 3943 6554 3999
rect 6610 3943 6658 3999
rect 6714 3943 6724 3999
rect 6544 3933 6724 3943
rect 6854 4103 7034 4113
rect 6854 4047 6864 4103
rect 6920 4047 6968 4103
rect 7024 4047 7034 4103
rect 6854 3999 7034 4047
rect 6854 3943 6864 3999
rect 6920 3943 6968 3999
rect 7024 3943 7034 3999
rect 6854 3933 7034 3943
rect 6093 2889 6273 2899
rect 6093 2833 6103 2889
rect 6159 2833 6207 2889
rect 6263 2833 6273 2889
rect 6093 2785 6273 2833
rect 6093 2729 6103 2785
rect 6159 2729 6207 2785
rect 6263 2729 6273 2785
rect 6093 2719 6273 2729
rect 6582 2402 6658 2412
rect 6582 2346 6592 2402
rect 6648 2346 6658 2402
rect 6582 2298 6658 2346
rect 6582 2242 6592 2298
rect 6648 2242 6658 2298
rect 6582 2232 6658 2242
rect 6512 2016 6692 2026
rect 6512 1960 6522 2016
rect 6578 1960 6626 2016
rect 6682 1960 6692 2016
rect 6512 1912 6692 1960
rect 6512 1856 6522 1912
rect 6578 1856 6626 1912
rect 6682 1856 6692 1912
rect 6512 1846 6692 1856
rect 6422 1773 6498 1783
rect 6864 1777 7024 3933
rect 7118 2889 7298 2899
rect 7118 2833 7128 2889
rect 7184 2833 7232 2889
rect 7288 2833 7298 2889
rect 7118 2785 7298 2833
rect 7118 2729 7128 2785
rect 7184 2729 7232 2785
rect 7288 2729 7298 2785
rect 7118 2719 7298 2729
rect 7128 2016 7288 2719
rect 7392 2653 7552 6241
rect 9979 6185 10139 7211
rect 9969 6173 10149 6185
rect 9969 6121 9981 6173
rect 10033 6121 10085 6173
rect 10137 6121 10149 6173
rect 9969 6069 10149 6121
rect 9189 6044 9265 6054
rect 9189 5988 9199 6044
rect 9255 5988 9265 6044
rect 9969 6017 9981 6069
rect 10033 6017 10085 6069
rect 10137 6017 10149 6069
rect 9969 6005 10149 6017
rect 10278 6044 10458 6054
rect 9189 5940 9265 5988
rect 9189 5884 9199 5940
rect 9255 5884 9265 5940
rect 9189 5874 9265 5884
rect 10278 5988 10288 6044
rect 10344 5988 10392 6044
rect 10448 5988 10458 6044
rect 10278 5940 10458 5988
rect 10278 5884 10288 5940
rect 10344 5884 10392 5940
rect 10448 5884 10458 5940
rect 10278 5874 10458 5884
rect 7669 5709 7745 5721
rect 7669 5657 7681 5709
rect 7733 5657 7745 5709
rect 7669 5605 7745 5657
rect 7669 5553 7681 5605
rect 7733 5553 7745 5605
rect 7669 5541 7745 5553
rect 7829 5711 7905 5721
rect 7829 5655 7839 5711
rect 7895 5655 7905 5711
rect 7829 5607 7905 5655
rect 7829 5551 7839 5607
rect 7895 5551 7905 5607
rect 7829 5541 7905 5551
rect 8149 5711 8225 5721
rect 8149 5655 8159 5711
rect 8215 5655 8225 5711
rect 8149 5607 8225 5655
rect 8149 5551 8159 5607
rect 8215 5551 8225 5607
rect 8149 5541 8225 5551
rect 8469 5711 8545 5721
rect 8469 5655 8479 5711
rect 8535 5655 8545 5711
rect 8469 5607 8545 5655
rect 8469 5551 8479 5607
rect 8535 5551 8545 5607
rect 8469 5541 8545 5551
rect 8789 5711 8865 5721
rect 8789 5655 8799 5711
rect 8855 5655 8865 5711
rect 8789 5607 8865 5655
rect 8789 5551 8799 5607
rect 8855 5551 8865 5607
rect 8789 5541 8865 5551
rect 8949 5711 9025 5720
rect 8949 5655 8959 5711
rect 9015 5655 9025 5711
rect 8949 5607 9025 5655
rect 8949 5551 8959 5607
rect 9015 5551 9025 5607
rect 7679 4649 7735 5541
rect 7839 5185 7895 5541
rect 8949 5540 9025 5551
rect 9109 5709 9185 5721
rect 9109 5657 9121 5709
rect 9173 5657 9185 5709
rect 9109 5605 9185 5657
rect 9109 5553 9121 5605
rect 9173 5553 9185 5605
rect 9109 5541 9185 5553
rect 7829 5173 7905 5185
rect 7829 5121 7841 5173
rect 7893 5121 7905 5173
rect 7829 5069 7905 5121
rect 7829 5017 7841 5069
rect 7893 5017 7905 5069
rect 7829 5005 7905 5017
rect 7989 5175 8065 5184
rect 7989 5119 7999 5175
rect 8055 5119 8065 5175
rect 7989 5071 8065 5119
rect 7989 5015 7999 5071
rect 8055 5015 8065 5071
rect 7839 4649 7895 5005
rect 7989 5004 8065 5015
rect 8149 5175 8225 5185
rect 8149 5119 8159 5175
rect 8215 5119 8225 5175
rect 8149 5071 8225 5119
rect 8149 5015 8159 5071
rect 8215 5015 8225 5071
rect 8149 5005 8225 5015
rect 8469 5175 8545 5185
rect 8469 5119 8479 5175
rect 8535 5119 8545 5175
rect 8469 5071 8545 5119
rect 8469 5015 8479 5071
rect 8535 5015 8545 5071
rect 8469 5005 8545 5015
rect 8789 5175 8865 5185
rect 8789 5119 8799 5175
rect 8855 5119 8865 5175
rect 8789 5071 8865 5119
rect 8789 5015 8799 5071
rect 8855 5015 8865 5071
rect 8789 5005 8865 5015
rect 7669 4637 7745 4649
rect 7669 4585 7681 4637
rect 7733 4585 7745 4637
rect 7669 4533 7745 4585
rect 7669 4481 7681 4533
rect 7733 4481 7745 4533
rect 7669 4469 7745 4481
rect 7829 4639 7905 4649
rect 7829 4583 7839 4639
rect 7895 4583 7905 4639
rect 7829 4535 7905 4583
rect 7829 4479 7839 4535
rect 7895 4479 7905 4535
rect 7829 4469 7905 4479
rect 7839 4113 7895 4469
rect 7829 4103 7905 4113
rect 7999 4112 8055 5004
rect 8159 4649 8215 5005
rect 8959 4649 9015 5540
rect 9119 5185 9175 5541
rect 9268 5404 9344 5414
rect 9268 5348 9278 5404
rect 9334 5348 9344 5404
rect 9268 5338 9344 5348
rect 9109 5175 9185 5185
rect 9109 5119 9119 5175
rect 9175 5119 9185 5175
rect 9109 5071 9185 5119
rect 9109 5015 9119 5071
rect 9175 5015 9185 5071
rect 9109 5005 9185 5015
rect 10288 4930 10448 5874
rect 10544 5446 10724 5456
rect 10544 5390 10554 5446
rect 10610 5390 10658 5446
rect 10714 5390 10724 5446
rect 10544 5342 10724 5390
rect 10544 5286 10554 5342
rect 10610 5286 10658 5342
rect 10714 5286 10724 5342
rect 10544 5276 10724 5286
rect 10278 4920 10458 4930
rect 9071 4868 9147 4878
rect 9071 4812 9081 4868
rect 9137 4812 9147 4868
rect 9071 4802 9147 4812
rect 10278 4864 10288 4920
rect 10344 4864 10392 4920
rect 10448 4864 10458 4920
rect 10278 4816 10458 4864
rect 10278 4760 10288 4816
rect 10344 4760 10392 4816
rect 10448 4760 10458 4816
rect 10278 4750 10458 4760
rect 8149 4639 8225 4649
rect 8149 4583 8159 4639
rect 8215 4583 8225 4639
rect 8149 4535 8225 4583
rect 8149 4479 8159 4535
rect 8215 4479 8225 4535
rect 8149 4469 8225 4479
rect 8469 4639 8545 4649
rect 8469 4583 8479 4639
rect 8535 4583 8545 4639
rect 8469 4535 8545 4583
rect 8469 4479 8479 4535
rect 8535 4479 8545 4535
rect 8469 4469 8545 4479
rect 8789 4639 8865 4649
rect 8789 4583 8799 4639
rect 8855 4583 8865 4639
rect 8789 4535 8865 4583
rect 8789 4479 8799 4535
rect 8855 4479 8865 4535
rect 8789 4469 8865 4479
rect 8949 4637 9025 4649
rect 8949 4585 8961 4637
rect 9013 4585 9025 4637
rect 8949 4533 9025 4585
rect 8949 4481 8961 4533
rect 9013 4481 9025 4533
rect 8949 4468 9025 4481
rect 9109 4639 9185 4649
rect 9109 4583 9119 4639
rect 9175 4583 9185 4639
rect 9109 4535 9185 4583
rect 9109 4479 9119 4535
rect 9175 4479 9185 4535
rect 9109 4469 9185 4479
rect 7829 4047 7839 4103
rect 7895 4047 7905 4103
rect 7829 3999 7905 4047
rect 7829 3943 7839 3999
rect 7895 3943 7905 3999
rect 7829 3933 7905 3943
rect 7989 4101 8065 4112
rect 7989 4049 8001 4101
rect 8053 4049 8065 4101
rect 7989 3997 8065 4049
rect 7989 3945 8001 3997
rect 8053 3945 8065 3997
rect 7839 3585 7895 3933
rect 7989 3932 8065 3945
rect 8149 4103 8225 4113
rect 8149 4047 8159 4103
rect 8215 4047 8225 4103
rect 8149 3999 8225 4047
rect 8149 3943 8159 3999
rect 8215 3943 8225 3999
rect 8149 3933 8225 3943
rect 8469 4103 8545 4113
rect 8469 4047 8479 4103
rect 8535 4047 8545 4103
rect 8469 3999 8545 4047
rect 8469 3943 8479 3999
rect 8535 3943 8545 3999
rect 8469 3933 8545 3943
rect 8789 4103 8865 4113
rect 8789 4047 8799 4103
rect 8855 4047 8865 4103
rect 8789 3999 8865 4047
rect 8789 3943 8799 3999
rect 8855 3943 8865 3999
rect 8789 3933 8865 3943
rect 7829 3573 7905 3585
rect 7829 3521 7841 3573
rect 7893 3521 7905 3573
rect 7829 3469 7905 3521
rect 7829 3417 7841 3469
rect 7893 3417 7905 3469
rect 7829 3405 7905 3417
rect 7839 3049 7895 3405
rect 7829 3037 7905 3049
rect 7999 3040 8055 3932
rect 8159 3585 8215 3933
rect 8479 3585 8535 3933
rect 8799 3585 8855 3933
rect 8149 3573 8225 3585
rect 8149 3521 8161 3573
rect 8213 3521 8225 3573
rect 8149 3469 8225 3521
rect 8149 3417 8161 3469
rect 8213 3417 8225 3469
rect 8149 3405 8225 3417
rect 8469 3573 8545 3585
rect 8469 3521 8481 3573
rect 8533 3521 8545 3573
rect 8469 3469 8545 3521
rect 8469 3417 8481 3469
rect 8533 3417 8545 3469
rect 8469 3405 8545 3417
rect 8789 3573 8865 3585
rect 8959 3577 9015 4468
rect 9189 4334 9265 4344
rect 9189 4278 9199 4334
rect 9255 4278 9265 4334
rect 9189 4268 9265 4278
rect 9109 4103 9185 4113
rect 9109 4047 9119 4103
rect 9175 4047 9185 4103
rect 9109 3999 9185 4047
rect 9109 3943 9119 3999
rect 9175 3943 9185 3999
rect 9109 3933 9185 3943
rect 9119 3585 9175 3933
rect 9268 3902 9344 3912
rect 9268 3846 9278 3902
rect 9334 3846 9344 3902
rect 9268 3798 9344 3846
rect 9268 3742 9278 3798
rect 9334 3742 9344 3798
rect 9268 3732 9344 3742
rect 10006 3902 10186 3912
rect 10288 3910 10448 4750
rect 10554 4396 10714 5276
rect 10544 4386 10724 4396
rect 10544 4330 10554 4386
rect 10610 4330 10658 4386
rect 10714 4330 10724 4386
rect 10544 4282 10724 4330
rect 10544 4226 10554 4282
rect 10610 4226 10658 4282
rect 10714 4226 10724 4282
rect 10544 4216 10724 4226
rect 10006 3846 10016 3902
rect 10072 3846 10120 3902
rect 10176 3846 10186 3902
rect 10006 3798 10186 3846
rect 10006 3742 10016 3798
rect 10072 3742 10120 3798
rect 10176 3742 10186 3798
rect 10006 3732 10186 3742
rect 10278 3900 10458 3910
rect 10278 3844 10288 3900
rect 10344 3844 10392 3900
rect 10448 3844 10458 3900
rect 10278 3796 10458 3844
rect 10278 3740 10288 3796
rect 10344 3740 10392 3796
rect 10448 3740 10458 3796
rect 8789 3521 8801 3573
rect 8853 3521 8865 3573
rect 8789 3469 8865 3521
rect 8789 3417 8801 3469
rect 8853 3417 8865 3469
rect 8789 3405 8865 3417
rect 8949 3567 9025 3577
rect 8949 3511 8959 3567
rect 9015 3511 9025 3567
rect 8949 3463 9025 3511
rect 8949 3407 8959 3463
rect 9015 3407 9025 3463
rect 8159 3049 8215 3405
rect 8479 3049 8535 3405
rect 8799 3049 8855 3405
rect 8949 3396 9025 3407
rect 9109 3573 9185 3585
rect 9109 3521 9121 3573
rect 9173 3521 9185 3573
rect 9109 3469 9185 3521
rect 9109 3417 9121 3469
rect 9173 3417 9185 3469
rect 9109 3405 9185 3417
rect 9119 3049 9175 3405
rect 9268 3387 9344 3397
rect 9268 3331 9278 3387
rect 9334 3331 9344 3387
rect 9268 3283 9344 3331
rect 9268 3227 9278 3283
rect 9334 3227 9344 3283
rect 9268 3217 9344 3227
rect 9739 3161 9919 3171
rect 9739 3105 9749 3161
rect 9805 3105 9853 3161
rect 9909 3105 9919 3161
rect 9739 3057 9919 3105
rect 7829 2985 7841 3037
rect 7893 2985 7905 3037
rect 7829 2933 7905 2985
rect 7829 2881 7841 2933
rect 7893 2881 7905 2933
rect 7829 2869 7905 2881
rect 7989 3029 8065 3040
rect 7989 2977 8001 3029
rect 8053 2977 8065 3029
rect 7989 2925 8065 2977
rect 7989 2873 8001 2925
rect 8053 2873 8065 2925
rect 7989 2860 8065 2873
rect 8149 3037 8225 3049
rect 8149 2985 8161 3037
rect 8213 2985 8225 3037
rect 8149 2933 8225 2985
rect 8149 2881 8161 2933
rect 8213 2881 8225 2933
rect 8149 2869 8225 2881
rect 8469 3037 8545 3049
rect 8469 2985 8481 3037
rect 8533 2985 8545 3037
rect 8469 2933 8545 2985
rect 8469 2881 8481 2933
rect 8533 2881 8545 2933
rect 8469 2869 8545 2881
rect 8789 3037 8865 3049
rect 8789 2985 8801 3037
rect 8853 2985 8865 3037
rect 8789 2933 8865 2985
rect 8789 2881 8801 2933
rect 8853 2881 8865 2933
rect 8789 2869 8865 2881
rect 9109 3037 9185 3049
rect 9109 2985 9121 3037
rect 9173 2985 9185 3037
rect 9739 3001 9749 3057
rect 9805 3001 9853 3057
rect 9909 3001 9919 3057
rect 9739 2991 9919 3001
rect 9109 2933 9185 2985
rect 9109 2881 9121 2933
rect 9173 2881 9185 2933
rect 9109 2869 9185 2881
rect 8869 2711 8945 2721
rect 8869 2655 8879 2711
rect 8935 2655 8945 2711
rect 7384 2639 7564 2653
rect 7384 2587 7394 2639
rect 7446 2587 7498 2639
rect 7550 2587 7564 2639
rect 7384 2535 7564 2587
rect 8869 2607 8945 2655
rect 8869 2551 8879 2607
rect 8935 2551 8945 2607
rect 8869 2541 8945 2551
rect 7384 2483 7394 2535
rect 7446 2483 7498 2535
rect 7550 2483 7564 2535
rect 7384 2473 7564 2483
rect 9749 2416 9909 2991
rect 10016 2721 10176 3732
rect 10278 3730 10458 3740
rect 10554 3397 10714 4216
rect 10544 3387 10724 3397
rect 10544 3331 10554 3387
rect 10610 3331 10658 3387
rect 10714 3331 10724 3387
rect 10544 3283 10724 3331
rect 10544 3227 10554 3283
rect 10610 3227 10658 3283
rect 10714 3227 10724 3283
rect 10544 3217 10724 3227
rect 10006 2711 10186 2721
rect 10006 2655 10016 2711
rect 10072 2655 10120 2711
rect 10176 2655 10186 2711
rect 10006 2607 10186 2655
rect 10006 2551 10016 2607
rect 10072 2551 10120 2607
rect 10176 2551 10186 2607
rect 10006 2541 10186 2551
rect 10313 2636 10493 2648
rect 10313 2584 10325 2636
rect 10377 2584 10429 2636
rect 10481 2584 10493 2636
rect 10313 2532 10493 2584
rect 10313 2480 10325 2532
rect 10377 2480 10429 2532
rect 10481 2480 10493 2532
rect 10313 2468 10493 2480
rect 9737 2404 9917 2416
rect 9737 2352 9749 2404
rect 9801 2352 9853 2404
rect 9905 2352 9917 2404
rect 9737 2300 9917 2352
rect 9737 2248 9749 2300
rect 9801 2248 9853 2300
rect 9905 2248 9917 2300
rect 9737 2236 9917 2248
rect 7118 2006 7298 2016
rect 7118 1950 7128 2006
rect 7184 1950 7232 2006
rect 7288 1950 7298 2006
rect 7118 1902 7298 1950
rect 7118 1846 7128 1902
rect 7184 1846 7232 1902
rect 7288 1846 7298 1902
rect 7118 1836 7298 1846
rect 9396 2006 9576 2016
rect 9396 1950 9406 2006
rect 9462 1950 9510 2006
rect 9566 1950 9576 2006
rect 9396 1902 9576 1950
rect 9396 1846 9406 1902
rect 9462 1846 9510 1902
rect 9566 1846 9576 1902
rect 9396 1836 9576 1846
rect 6422 1717 6432 1773
rect 6488 1717 6498 1773
rect 6422 1669 6498 1717
rect 6422 1613 6432 1669
rect 6488 1613 6498 1669
rect 6422 1603 6498 1613
rect 6854 1767 7034 1777
rect 6854 1711 6864 1767
rect 6920 1711 6968 1767
rect 7024 1711 7034 1767
rect 6854 1663 7034 1711
rect 6854 1607 6864 1663
rect 6920 1607 6968 1663
rect 7024 1607 7034 1663
rect 6432 1139 6488 1603
rect 6854 1597 7034 1607
rect 6370 1129 6550 1139
rect 6370 1073 6380 1129
rect 6436 1073 6484 1129
rect 6540 1073 6550 1129
rect 6370 1025 6550 1073
rect 6370 969 6380 1025
rect 6436 969 6484 1025
rect 6540 969 6550 1025
rect 6370 959 6550 969
rect 10323 887 10483 2468
rect 10928 2016 11088 8285
rect 11381 8235 11541 9105
rect 11649 8715 11809 10151
rect 13984 10135 13994 10191
rect 14050 10135 14060 10191
rect 13984 10125 14060 10135
rect 15146 10295 15222 10305
rect 15146 10239 15156 10295
rect 15212 10239 15222 10295
rect 15146 10191 15222 10239
rect 15146 10135 15156 10191
rect 15212 10135 15222 10191
rect 15146 10125 15222 10135
rect 15786 10295 15862 10305
rect 15786 10239 15796 10295
rect 15852 10239 15862 10295
rect 15786 10191 15862 10239
rect 15786 10135 15796 10191
rect 15852 10135 15862 10191
rect 15786 10125 15862 10135
rect 16426 10295 16502 10305
rect 16426 10239 16436 10295
rect 16492 10239 16502 10295
rect 16426 10191 16502 10239
rect 16426 10135 16436 10191
rect 16492 10135 16502 10191
rect 16426 10125 16502 10135
rect 17103 10295 17283 10305
rect 17103 10239 17113 10295
rect 17169 10239 17217 10295
rect 17273 10239 17283 10295
rect 17103 10191 17283 10239
rect 17103 10135 17113 10191
rect 17169 10135 17217 10191
rect 17273 10135 17283 10191
rect 17103 10125 17283 10135
rect 12352 9275 12428 9285
rect 12352 9219 12362 9275
rect 12418 9219 12428 9275
rect 12352 9171 12428 9219
rect 12352 9115 12362 9171
rect 12418 9115 12428 9171
rect 12352 9105 12428 9115
rect 13248 9275 13324 9285
rect 13248 9219 13258 9275
rect 13314 9219 13324 9275
rect 13248 9171 13324 9219
rect 13248 9115 13258 9171
rect 13314 9115 13324 9171
rect 13248 9105 13324 9115
rect 14144 9275 14220 9285
rect 14144 9219 14154 9275
rect 14210 9219 14220 9275
rect 14144 9171 14220 9219
rect 14144 9115 14154 9171
rect 14210 9115 14220 9171
rect 14144 9105 14220 9115
rect 13856 8875 13932 8885
rect 13856 8819 13866 8875
rect 13922 8819 13932 8875
rect 13856 8771 13932 8819
rect 13856 8715 13866 8771
rect 13922 8715 13932 8771
rect 11639 8705 11819 8715
rect 13856 8705 13932 8715
rect 15466 8875 15542 8885
rect 15466 8819 15476 8875
rect 15532 8819 15542 8875
rect 15466 8771 15542 8819
rect 15466 8715 15476 8771
rect 15532 8715 15542 8771
rect 15466 8705 15542 8715
rect 16106 8875 16182 8885
rect 16106 8819 16116 8875
rect 16172 8819 16182 8875
rect 16106 8771 16182 8819
rect 16106 8715 16116 8771
rect 16172 8715 16182 8771
rect 16106 8705 16182 8715
rect 11639 8649 11649 8705
rect 11705 8649 11753 8705
rect 11809 8649 11819 8705
rect 11639 8601 11819 8649
rect 11639 8545 11649 8601
rect 11705 8545 11753 8601
rect 11809 8545 11819 8601
rect 11639 8535 11819 8545
rect 12018 8565 12198 8575
rect 11371 8225 11551 8235
rect 11371 8169 11381 8225
rect 11437 8169 11485 8225
rect 11541 8169 11551 8225
rect 11371 8121 11551 8169
rect 11371 8065 11381 8121
rect 11437 8065 11485 8121
rect 11541 8065 11551 8121
rect 11371 8055 11551 8065
rect 11381 6448 11541 8055
rect 11649 7835 11809 8535
rect 12018 8509 12028 8565
rect 12084 8509 12132 8565
rect 12188 8509 12198 8565
rect 12018 8461 12198 8509
rect 12018 8405 12028 8461
rect 12084 8405 12132 8461
rect 12188 8405 12198 8461
rect 12018 8395 12198 8405
rect 12388 8565 12464 8575
rect 12388 8509 12398 8565
rect 12454 8509 12464 8565
rect 12388 8461 12464 8509
rect 12388 8405 12398 8461
rect 12454 8405 12464 8461
rect 12388 8395 12464 8405
rect 14686 8570 14866 8580
rect 14686 8514 14696 8570
rect 14752 8514 14800 8570
rect 14856 8514 14866 8570
rect 14686 8466 14866 8514
rect 14686 8410 14696 8466
rect 14752 8410 14800 8466
rect 14856 8410 14866 8466
rect 14686 8400 14866 8410
rect 15174 8570 15250 8580
rect 15174 8514 15184 8570
rect 15240 8514 15250 8570
rect 15174 8466 15250 8514
rect 15174 8410 15184 8466
rect 15240 8410 15250 8466
rect 15174 8400 15250 8410
rect 11639 7825 11819 7835
rect 11639 7769 11649 7825
rect 11705 7769 11753 7825
rect 11809 7769 11819 7825
rect 11639 7721 11819 7769
rect 11639 7665 11649 7721
rect 11705 7665 11753 7721
rect 11809 7665 11819 7721
rect 11639 7655 11819 7665
rect 11371 6436 11551 6448
rect 11371 6384 11383 6436
rect 11435 6384 11487 6436
rect 11539 6384 11551 6436
rect 11371 6332 11551 6384
rect 11371 6280 11383 6332
rect 11435 6280 11487 6332
rect 11539 6280 11551 6332
rect 11371 6228 11551 6280
rect 11371 6176 11383 6228
rect 11435 6176 11487 6228
rect 11539 6176 11551 6228
rect 11371 6164 11551 6176
rect 11649 6106 11809 7655
rect 11639 6094 11819 6106
rect 11639 6042 11651 6094
rect 11703 6042 11755 6094
rect 11807 6042 11819 6094
rect 11639 5990 11819 6042
rect 11639 5938 11651 5990
rect 11703 5938 11755 5990
rect 11807 5938 11819 5990
rect 11639 5886 11819 5938
rect 11639 5834 11651 5886
rect 11703 5834 11755 5886
rect 11807 5834 11819 5886
rect 11639 5822 11819 5834
rect 10918 2006 11098 2016
rect 10918 1950 10928 2006
rect 10984 1950 11032 2006
rect 11088 1950 11098 2006
rect 10918 1902 11098 1950
rect 10918 1846 10928 1902
rect 10984 1846 11032 1902
rect 11088 1846 11098 1902
rect 10918 1836 11098 1846
rect 11305 2006 11485 2016
rect 11305 1950 11315 2006
rect 11371 1950 11419 2006
rect 11475 1950 11485 2006
rect 11305 1902 11485 1950
rect 11305 1846 11315 1902
rect 11371 1846 11419 1902
rect 11475 1846 11485 1902
rect 11305 1836 11485 1846
rect 12028 1139 12188 8395
rect 12800 8225 12876 8235
rect 12800 8169 12810 8225
rect 12866 8169 12876 8225
rect 12800 8121 12876 8169
rect 12800 8065 12810 8121
rect 12866 8065 12876 8121
rect 12800 8055 12876 8065
rect 13696 8225 13772 8235
rect 13696 8169 13706 8225
rect 13762 8169 13772 8225
rect 13696 8121 13772 8169
rect 13696 8065 13706 8121
rect 13762 8065 13772 8121
rect 13696 8055 13772 8065
rect 13856 8225 13932 8235
rect 13856 8169 13866 8225
rect 13922 8169 13932 8225
rect 13856 8121 13932 8169
rect 13856 8065 13866 8121
rect 13922 8065 13932 8121
rect 13856 8055 13932 8065
rect 12352 7825 12428 7835
rect 12352 7769 12362 7825
rect 12418 7769 12428 7825
rect 12352 7721 12428 7769
rect 12352 7665 12362 7721
rect 12418 7665 12428 7721
rect 12352 7655 12428 7665
rect 13248 7825 13324 7835
rect 13248 7769 13258 7825
rect 13314 7769 13324 7825
rect 13248 7721 13324 7769
rect 13248 7665 13258 7721
rect 13314 7665 13324 7721
rect 13248 7655 13324 7665
rect 14144 7825 14220 7835
rect 14144 7769 14154 7825
rect 14210 7769 14220 7825
rect 14144 7721 14220 7769
rect 14144 7665 14154 7721
rect 14210 7665 14220 7721
rect 14144 7655 14220 7665
rect 14696 5721 14856 8400
rect 17113 8235 17273 10125
rect 17375 8885 17535 11205
rect 17365 8875 17545 8885
rect 17365 8819 17375 8875
rect 17431 8819 17479 8875
rect 17535 8819 17545 8875
rect 17365 8771 17545 8819
rect 17365 8715 17375 8771
rect 17431 8715 17479 8771
rect 17535 8715 17545 8771
rect 17365 8705 17545 8715
rect 15466 8225 15542 8235
rect 15466 8169 15476 8225
rect 15532 8169 15542 8225
rect 15466 8121 15542 8169
rect 15466 8065 15476 8121
rect 15532 8065 15542 8121
rect 15466 8055 15542 8065
rect 16106 8225 16182 8235
rect 16106 8169 16116 8225
rect 16172 8169 16182 8225
rect 16106 8121 16182 8169
rect 16106 8065 16116 8121
rect 16172 8065 16182 8121
rect 16106 8055 16182 8065
rect 17103 8225 17283 8235
rect 17103 8169 17113 8225
rect 17169 8169 17217 8225
rect 17273 8169 17283 8225
rect 17103 8121 17283 8169
rect 17103 8065 17113 8121
rect 17169 8065 17217 8121
rect 17273 8065 17283 8121
rect 17103 8055 17283 8065
rect 17375 7845 17535 8705
rect 17641 8697 17716 11449
rect 17641 8641 17651 8697
rect 17707 8641 17716 8697
rect 17641 8631 17716 8641
rect 17841 12441 17917 12451
rect 17841 12385 17851 12441
rect 17907 12385 17917 12441
rect 17841 9633 17917 12385
rect 19065 12441 19141 12451
rect 19065 12385 19075 12441
rect 19131 12385 19141 12441
rect 19065 12375 19141 12385
rect 19305 12230 19381 12240
rect 19305 12174 19315 12230
rect 19371 12174 19381 12230
rect 19305 12126 19381 12174
rect 19305 12070 19315 12126
rect 19371 12070 19381 12126
rect 19305 12060 19381 12070
rect 19475 11846 19531 12602
rect 19795 11846 19851 12602
rect 19945 12230 20021 12240
rect 19945 12174 19955 12230
rect 20011 12174 20021 12230
rect 19945 12126 20021 12174
rect 19945 12070 19955 12126
rect 20011 12070 20021 12126
rect 19945 12060 20021 12070
rect 20115 11846 20171 12602
rect 21448 12334 21732 12612
rect 21448 12278 21458 12334
rect 21514 12278 21562 12334
rect 21618 12278 21666 12334
rect 21722 12278 21732 12334
rect 21448 12230 21732 12278
rect 21448 12174 21458 12230
rect 21514 12174 21562 12230
rect 21618 12174 21666 12230
rect 21722 12174 21732 12230
rect 21448 12126 21732 12174
rect 21448 12070 21458 12126
rect 21514 12070 21562 12126
rect 21618 12070 21666 12126
rect 21722 12070 21732 12126
rect 18985 11836 19061 11846
rect 18985 11780 18995 11836
rect 19051 11780 19061 11836
rect 18985 11732 19061 11780
rect 18985 11676 18995 11732
rect 19051 11676 19061 11732
rect 18985 11666 19061 11676
rect 19145 11834 19221 11846
rect 19145 11782 19157 11834
rect 19209 11782 19221 11834
rect 19145 11730 19221 11782
rect 19145 11678 19157 11730
rect 19209 11678 19221 11730
rect 19145 11666 19221 11678
rect 19465 11834 19541 11846
rect 19465 11782 19477 11834
rect 19529 11782 19541 11834
rect 19465 11730 19541 11782
rect 19465 11678 19477 11730
rect 19529 11678 19541 11730
rect 19465 11666 19541 11678
rect 19625 11836 19701 11846
rect 19625 11780 19635 11836
rect 19691 11780 19701 11836
rect 19625 11732 19701 11780
rect 19625 11676 19635 11732
rect 19691 11676 19701 11732
rect 19625 11666 19701 11676
rect 19785 11834 19861 11846
rect 19785 11782 19797 11834
rect 19849 11782 19861 11834
rect 19785 11730 19861 11782
rect 19785 11678 19797 11730
rect 19849 11678 19861 11730
rect 19785 11666 19861 11678
rect 20105 11834 20181 11846
rect 20105 11782 20117 11834
rect 20169 11782 20181 11834
rect 20105 11730 20181 11782
rect 20105 11678 20117 11730
rect 20169 11678 20181 11730
rect 20105 11666 20181 11678
rect 20265 11836 20341 11846
rect 20265 11780 20275 11836
rect 20331 11780 20341 11836
rect 20265 11732 20341 11780
rect 20265 11676 20275 11732
rect 20331 11676 20341 11732
rect 20265 11666 20341 11676
rect 19065 11505 19141 11515
rect 19065 11449 19075 11505
rect 19131 11449 19141 11505
rect 19065 11439 19141 11449
rect 19305 11294 19381 11304
rect 19305 11238 19315 11294
rect 19371 11238 19381 11294
rect 19305 11190 19381 11238
rect 19305 11134 19315 11190
rect 19371 11134 19381 11190
rect 19305 11124 19381 11134
rect 19475 10910 19531 11666
rect 19795 10910 19851 11666
rect 19945 11294 20021 11304
rect 19945 11238 19955 11294
rect 20011 11238 20021 11294
rect 19945 11190 20021 11238
rect 19945 11134 19955 11190
rect 20011 11134 20021 11190
rect 19945 11124 20021 11134
rect 20115 10910 20171 11666
rect 21448 11004 21732 12070
rect 21448 10948 21458 11004
rect 21514 10948 21562 11004
rect 21618 10948 21666 11004
rect 21722 10948 21732 11004
rect 18985 10900 19061 10910
rect 18985 10844 18995 10900
rect 19051 10844 19061 10900
rect 18985 10796 19061 10844
rect 18985 10740 18995 10796
rect 19051 10740 19061 10796
rect 18985 10730 19061 10740
rect 19145 10898 19221 10910
rect 19145 10846 19157 10898
rect 19209 10846 19221 10898
rect 19145 10794 19221 10846
rect 19145 10742 19157 10794
rect 19209 10742 19221 10794
rect 19145 10730 19221 10742
rect 19465 10898 19541 10910
rect 19465 10846 19477 10898
rect 19529 10846 19541 10898
rect 19465 10794 19541 10846
rect 19465 10742 19477 10794
rect 19529 10742 19541 10794
rect 19465 10730 19541 10742
rect 19625 10900 19701 10910
rect 19625 10844 19635 10900
rect 19691 10844 19701 10900
rect 19625 10796 19701 10844
rect 19625 10740 19635 10796
rect 19691 10740 19701 10796
rect 19625 10730 19701 10740
rect 19785 10898 19861 10910
rect 19785 10846 19797 10898
rect 19849 10846 19861 10898
rect 19785 10794 19861 10846
rect 19785 10742 19797 10794
rect 19849 10742 19861 10794
rect 19785 10730 19861 10742
rect 20105 10898 20181 10910
rect 20105 10846 20117 10898
rect 20169 10846 20181 10898
rect 20105 10794 20181 10846
rect 20105 10742 20117 10794
rect 20169 10742 20181 10794
rect 20105 10730 20181 10742
rect 20265 10900 20341 10910
rect 20265 10844 20275 10900
rect 20331 10844 20341 10900
rect 20265 10796 20341 10844
rect 20265 10740 20275 10796
rect 20331 10740 20341 10796
rect 20265 10730 20341 10740
rect 21448 10900 21732 10948
rect 21448 10844 21458 10900
rect 21514 10844 21562 10900
rect 21618 10844 21666 10900
rect 21722 10844 21732 10900
rect 21448 10796 21732 10844
rect 21448 10740 21458 10796
rect 21514 10740 21562 10796
rect 21618 10740 21666 10796
rect 21722 10740 21732 10796
rect 19305 10358 19381 10368
rect 19305 10302 19315 10358
rect 19371 10302 19381 10358
rect 19305 10254 19381 10302
rect 19305 10198 19315 10254
rect 19371 10198 19381 10254
rect 19305 10188 19381 10198
rect 18985 9964 19061 9974
rect 18985 9908 18995 9964
rect 19051 9908 19061 9964
rect 18985 9860 19061 9908
rect 18985 9804 18995 9860
rect 19051 9804 19061 9860
rect 18985 9794 19061 9804
rect 17841 9577 17851 9633
rect 17907 9577 17917 9633
rect 15146 7835 15222 7845
rect 15146 7779 15156 7835
rect 15212 7779 15222 7835
rect 15146 7731 15222 7779
rect 15146 7675 15156 7731
rect 15212 7675 15222 7731
rect 15146 7665 15222 7675
rect 15786 7835 15862 7845
rect 15786 7779 15796 7835
rect 15852 7779 15862 7835
rect 15786 7731 15862 7779
rect 15786 7675 15796 7731
rect 15852 7675 15862 7731
rect 15786 7665 15862 7675
rect 16426 7835 16502 7845
rect 16426 7779 16436 7835
rect 16492 7779 16502 7835
rect 16426 7731 16502 7779
rect 16426 7675 16436 7731
rect 16492 7675 16502 7731
rect 16426 7665 16502 7675
rect 17365 7835 17545 7845
rect 17365 7779 17375 7835
rect 17431 7779 17479 7835
rect 17535 7779 17545 7835
rect 17365 7731 17545 7779
rect 17365 7675 17375 7731
rect 17431 7675 17479 7731
rect 17535 7675 17545 7731
rect 17841 7761 17917 9577
rect 19065 9633 19141 9643
rect 19065 9577 19075 9633
rect 19131 9577 19141 9633
rect 19065 9567 19141 9577
rect 19305 9422 19381 9432
rect 19305 9366 19315 9422
rect 19371 9366 19381 9422
rect 19305 9318 19381 9366
rect 19305 9262 19315 9318
rect 19371 9262 19381 9318
rect 19305 9252 19381 9262
rect 19475 9038 19531 10730
rect 19625 9964 19701 9974
rect 19625 9908 19635 9964
rect 19691 9908 19701 9964
rect 19625 9860 19701 9908
rect 19625 9804 19635 9860
rect 19691 9804 19701 9860
rect 19625 9794 19701 9804
rect 19795 9038 19851 10730
rect 19945 10358 20021 10368
rect 19945 10302 19955 10358
rect 20011 10302 20021 10358
rect 19945 10254 20021 10302
rect 19945 10198 19955 10254
rect 20011 10198 20021 10254
rect 19945 10188 20021 10198
rect 19945 9422 20021 9432
rect 19945 9366 19955 9422
rect 20011 9366 20021 9422
rect 19945 9318 20021 9366
rect 19945 9262 19955 9318
rect 20011 9262 20021 9318
rect 19945 9252 20021 9262
rect 20115 9038 20171 10730
rect 21448 10068 21732 10740
rect 21448 10012 21458 10068
rect 21514 10012 21562 10068
rect 21618 10012 21666 10068
rect 21722 10012 21732 10068
rect 20265 9964 20341 9974
rect 20265 9908 20275 9964
rect 20331 9908 20341 9964
rect 20265 9860 20341 9908
rect 20265 9804 20275 9860
rect 20331 9804 20341 9860
rect 20265 9794 20341 9804
rect 21448 9964 21732 10012
rect 21448 9908 21458 9964
rect 21514 9908 21562 9964
rect 21618 9908 21666 9964
rect 21722 9908 21732 9964
rect 21448 9860 21732 9908
rect 21448 9804 21458 9860
rect 21514 9804 21562 9860
rect 21618 9804 21666 9860
rect 21722 9804 21732 9860
rect 21448 9526 21732 9804
rect 21448 9470 21458 9526
rect 21514 9470 21562 9526
rect 21618 9470 21666 9526
rect 21722 9470 21732 9526
rect 21448 9422 21732 9470
rect 21448 9366 21458 9422
rect 21514 9366 21562 9422
rect 21618 9366 21666 9422
rect 21722 9366 21732 9422
rect 21448 9318 21732 9366
rect 21448 9262 21458 9318
rect 21514 9262 21562 9318
rect 21618 9262 21666 9318
rect 21722 9262 21732 9318
rect 18985 9028 19061 9038
rect 18985 8972 18995 9028
rect 19051 8972 19061 9028
rect 18985 8924 19061 8972
rect 18985 8868 18995 8924
rect 19051 8868 19061 8924
rect 18985 8858 19061 8868
rect 19145 9026 19221 9038
rect 19145 8974 19157 9026
rect 19209 8974 19221 9026
rect 19145 8922 19221 8974
rect 19145 8870 19157 8922
rect 19209 8870 19221 8922
rect 19145 8858 19221 8870
rect 19465 9026 19541 9038
rect 19465 8974 19477 9026
rect 19529 8974 19541 9026
rect 19465 8922 19541 8974
rect 19465 8870 19477 8922
rect 19529 8870 19541 8922
rect 19465 8858 19541 8870
rect 19625 9028 19701 9038
rect 19625 8972 19635 9028
rect 19691 8972 19701 9028
rect 19625 8924 19701 8972
rect 19625 8868 19635 8924
rect 19691 8868 19701 8924
rect 19625 8858 19701 8868
rect 19785 9026 19861 9038
rect 19785 8974 19797 9026
rect 19849 8974 19861 9026
rect 19785 8922 19861 8974
rect 19785 8870 19797 8922
rect 19849 8870 19861 8922
rect 19785 8858 19861 8870
rect 20105 9026 20181 9038
rect 20105 8974 20117 9026
rect 20169 8974 20181 9026
rect 20105 8922 20181 8974
rect 20105 8870 20117 8922
rect 20169 8870 20181 8922
rect 20105 8858 20181 8870
rect 20265 9028 20341 9038
rect 20265 8972 20275 9028
rect 20331 8972 20341 9028
rect 20265 8924 20341 8972
rect 20265 8868 20275 8924
rect 20331 8868 20341 8924
rect 20265 8858 20341 8868
rect 19065 8697 19141 8707
rect 19065 8641 19075 8697
rect 19131 8641 19141 8697
rect 19065 8631 19141 8641
rect 19305 8486 19381 8496
rect 19305 8430 19315 8486
rect 19371 8430 19381 8486
rect 19305 8382 19381 8430
rect 19305 8326 19315 8382
rect 19371 8326 19381 8382
rect 19305 8316 19381 8326
rect 19475 8102 19531 8858
rect 19795 8102 19851 8858
rect 19945 8486 20021 8496
rect 19945 8430 19955 8486
rect 20011 8430 20021 8486
rect 19945 8382 20021 8430
rect 19945 8326 19955 8382
rect 20011 8326 20021 8382
rect 19945 8316 20021 8326
rect 20115 8102 20171 8858
rect 21448 8196 21732 9262
rect 22097 11940 22381 13006
rect 24457 13166 24533 13176
rect 24457 13110 24467 13166
rect 24523 13110 24533 13166
rect 24457 13062 24533 13110
rect 24457 13006 24467 13062
rect 24523 13006 24533 13062
rect 24457 12996 24533 13006
rect 25097 13166 25173 13176
rect 25097 13110 25107 13166
rect 25163 13110 25173 13166
rect 25097 13062 25173 13110
rect 25097 13006 25107 13062
rect 25163 13006 25173 13062
rect 25097 12996 25173 13006
rect 22097 11884 22107 11940
rect 22163 11884 22211 11940
rect 22267 11884 22315 11940
rect 22371 11884 22381 11940
rect 22097 11836 22381 11884
rect 22097 11780 22107 11836
rect 22163 11780 22211 11836
rect 22267 11780 22315 11836
rect 22371 11780 22381 11836
rect 22097 11732 22381 11780
rect 22097 11676 22107 11732
rect 22163 11676 22211 11732
rect 22267 11676 22315 11732
rect 22371 11676 22381 11732
rect 22097 11398 22381 11676
rect 22097 11342 22107 11398
rect 22163 11342 22211 11398
rect 22267 11342 22315 11398
rect 22371 11342 22381 11398
rect 22097 11294 22381 11342
rect 22097 11238 22107 11294
rect 22163 11238 22211 11294
rect 22267 11238 22315 11294
rect 22371 11238 22381 11294
rect 22097 11190 22381 11238
rect 22097 11134 22107 11190
rect 22163 11134 22211 11190
rect 22267 11134 22315 11190
rect 22371 11134 22381 11190
rect 22097 10462 22381 11134
rect 22097 10406 22107 10462
rect 22163 10406 22211 10462
rect 22267 10406 22315 10462
rect 22371 10406 22381 10462
rect 22097 10358 22381 10406
rect 22097 10302 22107 10358
rect 22163 10302 22211 10358
rect 22267 10302 22315 10358
rect 22371 10302 22381 10358
rect 22097 10254 22381 10302
rect 22097 10198 22107 10254
rect 22163 10198 22211 10254
rect 22267 10198 22315 10254
rect 22371 10198 22381 10254
rect 22097 9132 22381 10198
rect 22097 9076 22107 9132
rect 22163 9076 22211 9132
rect 22267 9076 22315 9132
rect 22371 9076 22381 9132
rect 22097 9028 22381 9076
rect 22097 8972 22107 9028
rect 22163 8972 22211 9028
rect 22267 8972 22315 9028
rect 22371 8972 22381 9028
rect 22097 8924 22381 8972
rect 22097 8868 22107 8924
rect 22163 8868 22211 8924
rect 22267 8868 22315 8924
rect 22371 8868 22381 8924
rect 22097 8590 22381 8868
rect 22097 8534 22107 8590
rect 22163 8534 22211 8590
rect 22267 8534 22315 8590
rect 22371 8534 22381 8590
rect 22097 8486 22381 8534
rect 22097 8430 22107 8486
rect 22163 8430 22211 8486
rect 22267 8430 22315 8486
rect 22371 8430 22381 8486
rect 22097 8382 22381 8430
rect 22097 8326 22107 8382
rect 22163 8326 22211 8382
rect 22267 8326 22315 8382
rect 22371 8326 22381 8382
rect 22097 8316 22381 8326
rect 22746 12876 23030 12886
rect 22746 12820 22756 12876
rect 22812 12820 22860 12876
rect 22916 12820 22964 12876
rect 23020 12820 23030 12876
rect 22746 12772 23030 12820
rect 22746 12716 22756 12772
rect 22812 12716 22860 12772
rect 22916 12716 22964 12772
rect 23020 12716 23030 12772
rect 22746 12668 23030 12716
rect 22746 12612 22756 12668
rect 22812 12612 22860 12668
rect 22916 12612 22964 12668
rect 23020 12612 23030 12668
rect 22746 12334 23030 12612
rect 24137 12772 24213 12782
rect 24137 12716 24147 12772
rect 24203 12716 24213 12772
rect 24137 12668 24213 12716
rect 24137 12612 24147 12668
rect 24203 12612 24213 12668
rect 24137 12602 24213 12612
rect 24297 12770 24373 12782
rect 24297 12718 24309 12770
rect 24361 12718 24373 12770
rect 24297 12666 24373 12718
rect 24297 12614 24309 12666
rect 24361 12614 24373 12666
rect 24297 12602 24373 12614
rect 24617 12770 24693 12782
rect 24617 12718 24629 12770
rect 24681 12718 24693 12770
rect 24617 12666 24693 12718
rect 24617 12614 24629 12666
rect 24681 12614 24693 12666
rect 24617 12602 24693 12614
rect 24777 12772 24853 12782
rect 24777 12716 24787 12772
rect 24843 12716 24853 12772
rect 24777 12668 24853 12716
rect 24777 12612 24787 12668
rect 24843 12612 24853 12668
rect 24777 12602 24853 12612
rect 24937 12770 25013 12782
rect 24937 12718 24949 12770
rect 25001 12718 25013 12770
rect 24937 12666 25013 12718
rect 24937 12614 24949 12666
rect 25001 12614 25013 12666
rect 24937 12602 25013 12614
rect 25257 12770 25333 12782
rect 25257 12718 25269 12770
rect 25321 12718 25333 12770
rect 25257 12666 25333 12718
rect 25257 12614 25269 12666
rect 25321 12614 25333 12666
rect 25257 12602 25333 12614
rect 25417 12772 25493 12782
rect 25417 12716 25427 12772
rect 25483 12716 25493 12772
rect 25417 12668 25493 12716
rect 25417 12612 25427 12668
rect 25483 12612 25493 12668
rect 25417 12602 25493 12612
rect 22746 12278 22756 12334
rect 22812 12278 22860 12334
rect 22916 12278 22964 12334
rect 23020 12278 23030 12334
rect 22746 12230 23030 12278
rect 22746 12174 22756 12230
rect 22812 12174 22860 12230
rect 22916 12174 22964 12230
rect 23020 12174 23030 12230
rect 22746 12126 23030 12174
rect 22746 12070 22756 12126
rect 22812 12070 22860 12126
rect 22916 12070 22964 12126
rect 23020 12070 23030 12126
rect 22746 11004 23030 12070
rect 24307 11846 24363 12602
rect 24457 12230 24533 12240
rect 24457 12174 24467 12230
rect 24523 12174 24533 12230
rect 24457 12126 24533 12174
rect 24457 12070 24467 12126
rect 24523 12070 24533 12126
rect 24457 12060 24533 12070
rect 24627 11846 24683 12602
rect 24947 11846 25003 12602
rect 25337 12441 25413 12451
rect 25337 12385 25347 12441
rect 25403 12385 25413 12441
rect 25337 12375 25413 12385
rect 26561 12441 26637 12451
rect 26561 12385 26571 12441
rect 26627 12385 26637 12441
rect 25097 12230 25173 12240
rect 25097 12174 25107 12230
rect 25163 12174 25173 12230
rect 25097 12126 25173 12174
rect 25097 12070 25107 12126
rect 25163 12070 25173 12126
rect 25097 12060 25173 12070
rect 24137 11836 24213 11846
rect 24137 11780 24147 11836
rect 24203 11780 24213 11836
rect 24137 11732 24213 11780
rect 24137 11676 24147 11732
rect 24203 11676 24213 11732
rect 24137 11666 24213 11676
rect 24297 11834 24373 11846
rect 24297 11782 24309 11834
rect 24361 11782 24373 11834
rect 24297 11730 24373 11782
rect 24297 11678 24309 11730
rect 24361 11678 24373 11730
rect 24297 11666 24373 11678
rect 24617 11834 24693 11846
rect 24617 11782 24629 11834
rect 24681 11782 24693 11834
rect 24617 11730 24693 11782
rect 24617 11678 24629 11730
rect 24681 11678 24693 11730
rect 24617 11666 24693 11678
rect 24777 11836 24853 11846
rect 24777 11780 24787 11836
rect 24843 11780 24853 11836
rect 24777 11732 24853 11780
rect 24777 11676 24787 11732
rect 24843 11676 24853 11732
rect 24777 11666 24853 11676
rect 24937 11834 25013 11846
rect 24937 11782 24949 11834
rect 25001 11782 25013 11834
rect 24937 11730 25013 11782
rect 24937 11678 24949 11730
rect 25001 11678 25013 11730
rect 24937 11666 25013 11678
rect 25257 11834 25333 11846
rect 25257 11782 25269 11834
rect 25321 11782 25333 11834
rect 25257 11730 25333 11782
rect 25257 11678 25269 11730
rect 25321 11678 25333 11730
rect 25257 11666 25333 11678
rect 25417 11836 25493 11846
rect 25417 11780 25427 11836
rect 25483 11780 25493 11836
rect 25417 11732 25493 11780
rect 25417 11676 25427 11732
rect 25483 11676 25493 11732
rect 25417 11666 25493 11676
rect 22746 10948 22756 11004
rect 22812 10948 22860 11004
rect 22916 10948 22964 11004
rect 23020 10948 23030 11004
rect 22746 10900 23030 10948
rect 24307 10910 24363 11666
rect 24457 11294 24533 11304
rect 24457 11238 24467 11294
rect 24523 11238 24533 11294
rect 24457 11190 24533 11238
rect 24457 11134 24467 11190
rect 24523 11134 24533 11190
rect 24457 11124 24533 11134
rect 24627 10910 24683 11666
rect 24947 10910 25003 11666
rect 25337 11505 25413 11515
rect 25337 11449 25347 11505
rect 25403 11449 25413 11505
rect 25337 11439 25413 11449
rect 25097 11294 25173 11304
rect 25097 11238 25107 11294
rect 25163 11238 25173 11294
rect 25097 11190 25173 11238
rect 25097 11134 25107 11190
rect 25163 11134 25173 11190
rect 25097 11124 25173 11134
rect 22746 10844 22756 10900
rect 22812 10844 22860 10900
rect 22916 10844 22964 10900
rect 23020 10844 23030 10900
rect 22746 10796 23030 10844
rect 22746 10740 22756 10796
rect 22812 10740 22860 10796
rect 22916 10740 22964 10796
rect 23020 10740 23030 10796
rect 22746 10068 23030 10740
rect 24137 10900 24213 10910
rect 24137 10844 24147 10900
rect 24203 10844 24213 10900
rect 24137 10796 24213 10844
rect 24137 10740 24147 10796
rect 24203 10740 24213 10796
rect 24137 10730 24213 10740
rect 24297 10898 24373 10910
rect 24297 10846 24309 10898
rect 24361 10846 24373 10898
rect 24297 10794 24373 10846
rect 24297 10742 24309 10794
rect 24361 10742 24373 10794
rect 24297 10730 24373 10742
rect 24617 10898 24693 10910
rect 24617 10846 24629 10898
rect 24681 10846 24693 10898
rect 24617 10794 24693 10846
rect 24617 10742 24629 10794
rect 24681 10742 24693 10794
rect 24617 10730 24693 10742
rect 24777 10900 24853 10910
rect 24777 10844 24787 10900
rect 24843 10844 24853 10900
rect 24777 10796 24853 10844
rect 24777 10740 24787 10796
rect 24843 10740 24853 10796
rect 24777 10730 24853 10740
rect 24937 10898 25013 10910
rect 24937 10846 24949 10898
rect 25001 10846 25013 10898
rect 24937 10794 25013 10846
rect 24937 10742 24949 10794
rect 25001 10742 25013 10794
rect 24937 10730 25013 10742
rect 25257 10898 25333 10910
rect 25257 10846 25269 10898
rect 25321 10846 25333 10898
rect 25257 10794 25333 10846
rect 25257 10742 25269 10794
rect 25321 10742 25333 10794
rect 25257 10730 25333 10742
rect 25417 10900 25493 10910
rect 25417 10844 25427 10900
rect 25483 10844 25493 10900
rect 25417 10796 25493 10844
rect 25417 10740 25427 10796
rect 25483 10740 25493 10796
rect 25417 10730 25493 10740
rect 22746 10012 22756 10068
rect 22812 10012 22860 10068
rect 22916 10012 22964 10068
rect 23020 10012 23030 10068
rect 22746 9964 23030 10012
rect 22746 9908 22756 9964
rect 22812 9908 22860 9964
rect 22916 9908 22964 9964
rect 23020 9908 23030 9964
rect 22746 9860 23030 9908
rect 22746 9804 22756 9860
rect 22812 9804 22860 9860
rect 22916 9804 22964 9860
rect 23020 9804 23030 9860
rect 22746 9526 23030 9804
rect 24137 9964 24213 9974
rect 24137 9908 24147 9964
rect 24203 9908 24213 9964
rect 24137 9860 24213 9908
rect 24137 9804 24147 9860
rect 24203 9804 24213 9860
rect 24137 9794 24213 9804
rect 22746 9470 22756 9526
rect 22812 9470 22860 9526
rect 22916 9470 22964 9526
rect 23020 9470 23030 9526
rect 22746 9422 23030 9470
rect 22746 9366 22756 9422
rect 22812 9366 22860 9422
rect 22916 9366 22964 9422
rect 23020 9366 23030 9422
rect 22746 9318 23030 9366
rect 22746 9262 22756 9318
rect 22812 9262 22860 9318
rect 22916 9262 22964 9318
rect 23020 9262 23030 9318
rect 21448 8140 21458 8196
rect 21514 8140 21562 8196
rect 21618 8140 21666 8196
rect 21722 8140 21732 8196
rect 18985 8092 19061 8102
rect 18985 8036 18995 8092
rect 19051 8036 19061 8092
rect 18985 7988 19061 8036
rect 18985 7932 18995 7988
rect 19051 7932 19061 7988
rect 18985 7922 19061 7932
rect 19145 8090 19221 8102
rect 19145 8038 19157 8090
rect 19209 8038 19221 8090
rect 19145 7986 19221 8038
rect 19145 7934 19157 7986
rect 19209 7934 19221 7986
rect 19145 7922 19221 7934
rect 19465 8090 19541 8102
rect 19465 8038 19477 8090
rect 19529 8038 19541 8090
rect 19465 7986 19541 8038
rect 19465 7934 19477 7986
rect 19529 7934 19541 7986
rect 19465 7922 19541 7934
rect 19625 8092 19701 8102
rect 19625 8036 19635 8092
rect 19691 8036 19701 8092
rect 19625 7988 19701 8036
rect 19625 7932 19635 7988
rect 19691 7932 19701 7988
rect 19625 7922 19701 7932
rect 19785 8090 19861 8102
rect 19785 8038 19797 8090
rect 19849 8038 19861 8090
rect 19785 7986 19861 8038
rect 19785 7934 19797 7986
rect 19849 7934 19861 7986
rect 19785 7922 19861 7934
rect 20105 8090 20181 8102
rect 20105 8038 20117 8090
rect 20169 8038 20181 8090
rect 20105 7986 20181 8038
rect 20105 7934 20117 7986
rect 20169 7934 20181 7986
rect 20105 7922 20181 7934
rect 20265 8092 20341 8102
rect 20265 8036 20275 8092
rect 20331 8036 20341 8092
rect 20265 7988 20341 8036
rect 20265 7932 20275 7988
rect 20331 7932 20341 7988
rect 20265 7922 20341 7932
rect 21448 8092 21732 8140
rect 21448 8036 21458 8092
rect 21514 8036 21562 8092
rect 21618 8036 21666 8092
rect 21722 8036 21732 8092
rect 21448 7988 21732 8036
rect 21448 7932 21458 7988
rect 21514 7932 21562 7988
rect 21618 7932 21666 7988
rect 21722 7932 21732 7988
rect 21448 7922 21732 7932
rect 22746 8196 23030 9262
rect 24307 9038 24363 10730
rect 24457 10358 24533 10368
rect 24457 10302 24467 10358
rect 24523 10302 24533 10358
rect 24457 10254 24533 10302
rect 24457 10198 24467 10254
rect 24523 10198 24533 10254
rect 24457 10188 24533 10198
rect 24457 9422 24533 9432
rect 24457 9366 24467 9422
rect 24523 9366 24533 9422
rect 24457 9318 24533 9366
rect 24457 9262 24467 9318
rect 24523 9262 24533 9318
rect 24457 9252 24533 9262
rect 24627 9038 24683 10730
rect 24777 9964 24853 9974
rect 24777 9908 24787 9964
rect 24843 9908 24853 9964
rect 24777 9860 24853 9908
rect 24777 9804 24787 9860
rect 24843 9804 24853 9860
rect 24777 9794 24853 9804
rect 24947 9038 25003 10730
rect 25097 10358 25173 10368
rect 25097 10302 25107 10358
rect 25163 10302 25173 10358
rect 25097 10254 25173 10302
rect 25097 10198 25107 10254
rect 25163 10198 25173 10254
rect 25097 10188 25173 10198
rect 25417 9964 25493 9974
rect 25417 9908 25427 9964
rect 25483 9908 25493 9964
rect 25417 9860 25493 9908
rect 25417 9804 25427 9860
rect 25483 9804 25493 9860
rect 25417 9794 25493 9804
rect 25337 9633 25413 9643
rect 25337 9577 25347 9633
rect 25403 9577 25413 9633
rect 25337 9567 25413 9577
rect 26561 9633 26637 12385
rect 26561 9577 26571 9633
rect 26627 9577 26637 9633
rect 25097 9422 25173 9432
rect 25097 9366 25107 9422
rect 25163 9366 25173 9422
rect 25097 9318 25173 9366
rect 25097 9262 25107 9318
rect 25163 9262 25173 9318
rect 25097 9252 25173 9262
rect 24137 9028 24213 9038
rect 24137 8972 24147 9028
rect 24203 8972 24213 9028
rect 24137 8924 24213 8972
rect 24137 8868 24147 8924
rect 24203 8868 24213 8924
rect 24137 8858 24213 8868
rect 24297 9026 24373 9038
rect 24297 8974 24309 9026
rect 24361 8974 24373 9026
rect 24297 8922 24373 8974
rect 24297 8870 24309 8922
rect 24361 8870 24373 8922
rect 24297 8858 24373 8870
rect 24617 9026 24693 9038
rect 24617 8974 24629 9026
rect 24681 8974 24693 9026
rect 24617 8922 24693 8974
rect 24617 8870 24629 8922
rect 24681 8870 24693 8922
rect 24617 8858 24693 8870
rect 24777 9028 24853 9038
rect 24777 8972 24787 9028
rect 24843 8972 24853 9028
rect 24777 8924 24853 8972
rect 24777 8868 24787 8924
rect 24843 8868 24853 8924
rect 24777 8858 24853 8868
rect 24937 9026 25013 9038
rect 24937 8974 24949 9026
rect 25001 8974 25013 9026
rect 24937 8922 25013 8974
rect 24937 8870 24949 8922
rect 25001 8870 25013 8922
rect 24937 8858 25013 8870
rect 25257 9026 25333 9038
rect 25257 8974 25269 9026
rect 25321 8974 25333 9026
rect 25257 8922 25333 8974
rect 25257 8870 25269 8922
rect 25321 8870 25333 8922
rect 25257 8858 25333 8870
rect 25417 9028 25493 9038
rect 25417 8972 25427 9028
rect 25483 8972 25493 9028
rect 25417 8924 25493 8972
rect 25417 8868 25427 8924
rect 25483 8868 25493 8924
rect 25417 8858 25493 8868
rect 22746 8140 22756 8196
rect 22812 8140 22860 8196
rect 22916 8140 22964 8196
rect 23020 8140 23030 8196
rect 22746 8092 23030 8140
rect 24307 8102 24363 8858
rect 24457 8486 24533 8496
rect 24457 8430 24467 8486
rect 24523 8430 24533 8486
rect 24457 8382 24533 8430
rect 24457 8326 24467 8382
rect 24523 8326 24533 8382
rect 24457 8316 24533 8326
rect 24627 8102 24683 8858
rect 24947 8102 25003 8858
rect 25337 8697 25413 8707
rect 25337 8641 25347 8697
rect 25403 8641 25413 8697
rect 25337 8631 25413 8641
rect 25097 8486 25173 8496
rect 25097 8430 25107 8486
rect 25163 8430 25173 8486
rect 25097 8382 25173 8430
rect 25097 8326 25107 8382
rect 25163 8326 25173 8382
rect 25097 8316 25173 8326
rect 22746 8036 22756 8092
rect 22812 8036 22860 8092
rect 22916 8036 22964 8092
rect 23020 8036 23030 8092
rect 22746 7988 23030 8036
rect 22746 7932 22756 7988
rect 22812 7932 22860 7988
rect 22916 7932 22964 7988
rect 23020 7932 23030 7988
rect 22746 7922 23030 7932
rect 24137 8092 24213 8102
rect 24137 8036 24147 8092
rect 24203 8036 24213 8092
rect 24137 7988 24213 8036
rect 24137 7932 24147 7988
rect 24203 7932 24213 7988
rect 24137 7922 24213 7932
rect 24297 8090 24373 8102
rect 24297 8038 24309 8090
rect 24361 8038 24373 8090
rect 24297 7986 24373 8038
rect 24297 7934 24309 7986
rect 24361 7934 24373 7986
rect 24297 7922 24373 7934
rect 24617 8090 24693 8102
rect 24617 8038 24629 8090
rect 24681 8038 24693 8090
rect 24617 7986 24693 8038
rect 24617 7934 24629 7986
rect 24681 7934 24693 7986
rect 24617 7922 24693 7934
rect 24777 8092 24853 8102
rect 24777 8036 24787 8092
rect 24843 8036 24853 8092
rect 24777 7988 24853 8036
rect 24777 7932 24787 7988
rect 24843 7932 24853 7988
rect 24777 7922 24853 7932
rect 24937 8090 25013 8102
rect 24937 8038 24949 8090
rect 25001 8038 25013 8090
rect 24937 7986 25013 8038
rect 24937 7934 24949 7986
rect 25001 7934 25013 7986
rect 24937 7922 25013 7934
rect 25257 8090 25333 8102
rect 25257 8038 25269 8090
rect 25321 8038 25333 8090
rect 25257 7986 25333 8038
rect 25257 7934 25269 7986
rect 25321 7934 25333 7986
rect 25257 7922 25333 7934
rect 25417 8092 25493 8102
rect 25417 8036 25427 8092
rect 25483 8036 25493 8092
rect 25417 7988 25493 8036
rect 25417 7932 25427 7988
rect 25483 7932 25493 7988
rect 25417 7922 25493 7932
rect 17841 7705 17851 7761
rect 17907 7705 17917 7761
rect 17841 7695 17917 7705
rect 19225 7761 19301 7771
rect 19225 7705 19235 7761
rect 19291 7705 19301 7761
rect 19225 7695 19301 7705
rect 19865 7761 19941 7771
rect 19865 7705 19875 7761
rect 19931 7705 19941 7761
rect 19865 7695 19941 7705
rect 24537 7761 24613 7771
rect 24537 7705 24547 7761
rect 24603 7705 24613 7761
rect 24537 7695 24613 7705
rect 25177 7761 25253 7771
rect 25177 7705 25187 7761
rect 25243 7705 25253 7761
rect 25177 7695 25253 7705
rect 26561 7761 26637 9577
rect 26762 11505 26837 13351
rect 28186 13407 28262 13417
rect 28186 13351 28196 13407
rect 28252 13351 28262 13407
rect 28186 13341 28262 13351
rect 31218 13270 31502 15420
rect 31218 13214 31228 13270
rect 31284 13214 31332 13270
rect 31388 13214 31436 13270
rect 31492 13214 31502 13270
rect 28426 13166 28502 13176
rect 28426 13110 28436 13166
rect 28492 13110 28502 13166
rect 28426 13062 28502 13110
rect 28426 13006 28436 13062
rect 28492 13006 28502 13062
rect 28426 12996 28502 13006
rect 29066 13166 29142 13176
rect 29066 13110 29076 13166
rect 29132 13110 29142 13166
rect 29066 13062 29142 13110
rect 29066 13006 29076 13062
rect 29132 13006 29142 13062
rect 29066 12996 29142 13006
rect 31218 13166 31502 13214
rect 31218 13110 31228 13166
rect 31284 13110 31332 13166
rect 31388 13110 31436 13166
rect 31492 13110 31502 13166
rect 31218 13062 31502 13110
rect 31218 13006 31228 13062
rect 31284 13006 31332 13062
rect 31388 13006 31436 13062
rect 31492 13006 31502 13062
rect 30569 12876 30853 12886
rect 30569 12820 30579 12876
rect 30635 12820 30683 12876
rect 30739 12820 30787 12876
rect 30843 12820 30853 12876
rect 28106 12772 28182 12782
rect 28106 12716 28116 12772
rect 28172 12716 28182 12772
rect 28106 12668 28182 12716
rect 28106 12612 28116 12668
rect 28172 12612 28182 12668
rect 28106 12602 28182 12612
rect 28266 12770 28342 12782
rect 28266 12718 28278 12770
rect 28330 12718 28342 12770
rect 28266 12666 28342 12718
rect 28266 12614 28278 12666
rect 28330 12614 28342 12666
rect 28266 12602 28342 12614
rect 28586 12770 28662 12782
rect 28586 12718 28598 12770
rect 28650 12718 28662 12770
rect 28586 12666 28662 12718
rect 28586 12614 28598 12666
rect 28650 12614 28662 12666
rect 28586 12602 28662 12614
rect 28746 12772 28822 12782
rect 28746 12716 28756 12772
rect 28812 12716 28822 12772
rect 28746 12668 28822 12716
rect 28746 12612 28756 12668
rect 28812 12612 28822 12668
rect 28746 12602 28822 12612
rect 28906 12770 28982 12782
rect 28906 12718 28918 12770
rect 28970 12718 28982 12770
rect 28906 12666 28982 12718
rect 28906 12614 28918 12666
rect 28970 12614 28982 12666
rect 28906 12602 28982 12614
rect 29226 12770 29302 12782
rect 29226 12718 29238 12770
rect 29290 12718 29302 12770
rect 29226 12666 29302 12718
rect 29226 12614 29238 12666
rect 29290 12614 29302 12666
rect 29226 12602 29302 12614
rect 29386 12772 29462 12782
rect 29386 12716 29396 12772
rect 29452 12716 29462 12772
rect 29386 12668 29462 12716
rect 29386 12612 29396 12668
rect 29452 12612 29462 12668
rect 29386 12602 29462 12612
rect 30569 12772 30853 12820
rect 30569 12716 30579 12772
rect 30635 12716 30683 12772
rect 30739 12716 30787 12772
rect 30843 12716 30853 12772
rect 30569 12668 30853 12716
rect 30569 12612 30579 12668
rect 30635 12612 30683 12668
rect 30739 12612 30787 12668
rect 30843 12612 30853 12668
rect 26762 11449 26771 11505
rect 26828 11449 26837 11505
rect 26762 8697 26837 11449
rect 26762 8641 26771 8697
rect 26828 8641 26837 8697
rect 26762 8631 26837 8641
rect 26962 12441 27038 12451
rect 26962 12385 26972 12441
rect 27028 12385 27038 12441
rect 26962 9633 27038 12385
rect 28186 12441 28262 12451
rect 28186 12385 28196 12441
rect 28252 12385 28262 12441
rect 28186 12375 28262 12385
rect 28426 12230 28502 12240
rect 28426 12174 28436 12230
rect 28492 12174 28502 12230
rect 28426 12126 28502 12174
rect 28426 12070 28436 12126
rect 28492 12070 28502 12126
rect 28426 12060 28502 12070
rect 28596 11846 28652 12602
rect 28916 11846 28972 12602
rect 29066 12230 29142 12240
rect 29066 12174 29076 12230
rect 29132 12174 29142 12230
rect 29066 12126 29142 12174
rect 29066 12070 29076 12126
rect 29132 12070 29142 12126
rect 29066 12060 29142 12070
rect 29236 11846 29292 12602
rect 30569 12334 30853 12612
rect 30569 12278 30579 12334
rect 30635 12278 30683 12334
rect 30739 12278 30787 12334
rect 30843 12278 30853 12334
rect 30569 12230 30853 12278
rect 30569 12174 30579 12230
rect 30635 12174 30683 12230
rect 30739 12174 30787 12230
rect 30843 12174 30853 12230
rect 30569 12126 30853 12174
rect 30569 12070 30579 12126
rect 30635 12070 30683 12126
rect 30739 12070 30787 12126
rect 30843 12070 30853 12126
rect 28106 11836 28182 11846
rect 28106 11780 28116 11836
rect 28172 11780 28182 11836
rect 28106 11732 28182 11780
rect 28106 11676 28116 11732
rect 28172 11676 28182 11732
rect 28106 11666 28182 11676
rect 28266 11834 28342 11846
rect 28266 11782 28278 11834
rect 28330 11782 28342 11834
rect 28266 11730 28342 11782
rect 28266 11678 28278 11730
rect 28330 11678 28342 11730
rect 28266 11666 28342 11678
rect 28586 11834 28662 11846
rect 28586 11782 28598 11834
rect 28650 11782 28662 11834
rect 28586 11730 28662 11782
rect 28586 11678 28598 11730
rect 28650 11678 28662 11730
rect 28586 11666 28662 11678
rect 28746 11836 28822 11846
rect 28746 11780 28756 11836
rect 28812 11780 28822 11836
rect 28746 11732 28822 11780
rect 28746 11676 28756 11732
rect 28812 11676 28822 11732
rect 28746 11666 28822 11676
rect 28906 11834 28982 11846
rect 28906 11782 28918 11834
rect 28970 11782 28982 11834
rect 28906 11730 28982 11782
rect 28906 11678 28918 11730
rect 28970 11678 28982 11730
rect 28906 11666 28982 11678
rect 29226 11834 29302 11846
rect 29226 11782 29238 11834
rect 29290 11782 29302 11834
rect 29226 11730 29302 11782
rect 29226 11678 29238 11730
rect 29290 11678 29302 11730
rect 29226 11666 29302 11678
rect 29386 11836 29462 11846
rect 29386 11780 29396 11836
rect 29452 11780 29462 11836
rect 29386 11732 29462 11780
rect 29386 11676 29396 11732
rect 29452 11676 29462 11732
rect 29386 11666 29462 11676
rect 28186 11505 28262 11515
rect 28186 11449 28196 11505
rect 28252 11449 28262 11505
rect 28186 11439 28262 11449
rect 28426 11294 28502 11304
rect 28426 11238 28436 11294
rect 28492 11238 28502 11294
rect 28426 11190 28502 11238
rect 28426 11134 28436 11190
rect 28492 11134 28502 11190
rect 28426 11124 28502 11134
rect 28596 10910 28652 11666
rect 28916 10910 28972 11666
rect 29066 11294 29142 11304
rect 29066 11238 29076 11294
rect 29132 11238 29142 11294
rect 29066 11190 29142 11238
rect 29066 11134 29076 11190
rect 29132 11134 29142 11190
rect 29066 11124 29142 11134
rect 29236 10910 29292 11666
rect 30569 11004 30853 12070
rect 30569 10948 30579 11004
rect 30635 10948 30683 11004
rect 30739 10948 30787 11004
rect 30843 10948 30853 11004
rect 28106 10900 28182 10910
rect 28106 10844 28116 10900
rect 28172 10844 28182 10900
rect 28106 10796 28182 10844
rect 28106 10740 28116 10796
rect 28172 10740 28182 10796
rect 28106 10730 28182 10740
rect 28266 10898 28342 10910
rect 28266 10846 28278 10898
rect 28330 10846 28342 10898
rect 28266 10794 28342 10846
rect 28266 10742 28278 10794
rect 28330 10742 28342 10794
rect 28266 10730 28342 10742
rect 28586 10898 28662 10910
rect 28586 10846 28598 10898
rect 28650 10846 28662 10898
rect 28586 10794 28662 10846
rect 28586 10742 28598 10794
rect 28650 10742 28662 10794
rect 28586 10730 28662 10742
rect 28746 10900 28822 10910
rect 28746 10844 28756 10900
rect 28812 10844 28822 10900
rect 28746 10796 28822 10844
rect 28746 10740 28756 10796
rect 28812 10740 28822 10796
rect 28746 10730 28822 10740
rect 28906 10898 28982 10910
rect 28906 10846 28918 10898
rect 28970 10846 28982 10898
rect 28906 10794 28982 10846
rect 28906 10742 28918 10794
rect 28970 10742 28982 10794
rect 28906 10730 28982 10742
rect 29226 10898 29302 10910
rect 29226 10846 29238 10898
rect 29290 10846 29302 10898
rect 29226 10794 29302 10846
rect 29226 10742 29238 10794
rect 29290 10742 29302 10794
rect 29226 10730 29302 10742
rect 29386 10900 29462 10910
rect 29386 10844 29396 10900
rect 29452 10844 29462 10900
rect 29386 10796 29462 10844
rect 29386 10740 29396 10796
rect 29452 10740 29462 10796
rect 29386 10730 29462 10740
rect 30569 10900 30853 10948
rect 30569 10844 30579 10900
rect 30635 10844 30683 10900
rect 30739 10844 30787 10900
rect 30843 10844 30853 10900
rect 30569 10796 30853 10844
rect 30569 10740 30579 10796
rect 30635 10740 30683 10796
rect 30739 10740 30787 10796
rect 30843 10740 30853 10796
rect 28426 10358 28502 10368
rect 28426 10302 28436 10358
rect 28492 10302 28502 10358
rect 28426 10254 28502 10302
rect 28426 10198 28436 10254
rect 28492 10198 28502 10254
rect 28426 10188 28502 10198
rect 28106 9964 28182 9974
rect 28106 9908 28116 9964
rect 28172 9908 28182 9964
rect 28106 9860 28182 9908
rect 28106 9804 28116 9860
rect 28172 9804 28182 9860
rect 28106 9794 28182 9804
rect 26962 9577 26972 9633
rect 27028 9577 27038 9633
rect 26561 7705 26571 7761
rect 26627 7705 26637 7761
rect 26561 7695 26637 7705
rect 26962 7761 27038 9577
rect 28186 9633 28262 9643
rect 28186 9577 28196 9633
rect 28252 9577 28262 9633
rect 28186 9567 28262 9577
rect 28426 9422 28502 9432
rect 28426 9366 28436 9422
rect 28492 9366 28502 9422
rect 28426 9318 28502 9366
rect 28426 9262 28436 9318
rect 28492 9262 28502 9318
rect 28426 9252 28502 9262
rect 28596 9038 28652 10730
rect 28746 9964 28822 9974
rect 28746 9908 28756 9964
rect 28812 9908 28822 9964
rect 28746 9860 28822 9908
rect 28746 9804 28756 9860
rect 28812 9804 28822 9860
rect 28746 9794 28822 9804
rect 28916 9038 28972 10730
rect 29066 10358 29142 10368
rect 29066 10302 29076 10358
rect 29132 10302 29142 10358
rect 29066 10254 29142 10302
rect 29066 10198 29076 10254
rect 29132 10198 29142 10254
rect 29066 10188 29142 10198
rect 29066 9422 29142 9432
rect 29066 9366 29076 9422
rect 29132 9366 29142 9422
rect 29066 9318 29142 9366
rect 29066 9262 29076 9318
rect 29132 9262 29142 9318
rect 29066 9252 29142 9262
rect 29236 9038 29292 10730
rect 30569 10068 30853 10740
rect 30569 10012 30579 10068
rect 30635 10012 30683 10068
rect 30739 10012 30787 10068
rect 30843 10012 30853 10068
rect 29386 9964 29462 9974
rect 29386 9908 29396 9964
rect 29452 9908 29462 9964
rect 29386 9860 29462 9908
rect 29386 9804 29396 9860
rect 29452 9804 29462 9860
rect 29386 9794 29462 9804
rect 30569 9964 30853 10012
rect 30569 9908 30579 9964
rect 30635 9908 30683 9964
rect 30739 9908 30787 9964
rect 30843 9908 30853 9964
rect 30569 9860 30853 9908
rect 30569 9804 30579 9860
rect 30635 9804 30683 9860
rect 30739 9804 30787 9860
rect 30843 9804 30853 9860
rect 30569 9526 30853 9804
rect 30569 9470 30579 9526
rect 30635 9470 30683 9526
rect 30739 9470 30787 9526
rect 30843 9470 30853 9526
rect 30569 9422 30853 9470
rect 30569 9366 30579 9422
rect 30635 9366 30683 9422
rect 30739 9366 30787 9422
rect 30843 9366 30853 9422
rect 30569 9318 30853 9366
rect 30569 9262 30579 9318
rect 30635 9262 30683 9318
rect 30739 9262 30787 9318
rect 30843 9262 30853 9318
rect 28106 9028 28182 9038
rect 28106 8972 28116 9028
rect 28172 8972 28182 9028
rect 28106 8924 28182 8972
rect 28106 8868 28116 8924
rect 28172 8868 28182 8924
rect 28106 8858 28182 8868
rect 28266 9026 28342 9038
rect 28266 8974 28278 9026
rect 28330 8974 28342 9026
rect 28266 8922 28342 8974
rect 28266 8870 28278 8922
rect 28330 8870 28342 8922
rect 28266 8858 28342 8870
rect 28586 9026 28662 9038
rect 28586 8974 28598 9026
rect 28650 8974 28662 9026
rect 28586 8922 28662 8974
rect 28586 8870 28598 8922
rect 28650 8870 28662 8922
rect 28586 8858 28662 8870
rect 28746 9028 28822 9038
rect 28746 8972 28756 9028
rect 28812 8972 28822 9028
rect 28746 8924 28822 8972
rect 28746 8868 28756 8924
rect 28812 8868 28822 8924
rect 28746 8858 28822 8868
rect 28906 9026 28982 9038
rect 28906 8974 28918 9026
rect 28970 8974 28982 9026
rect 28906 8922 28982 8974
rect 28906 8870 28918 8922
rect 28970 8870 28982 8922
rect 28906 8858 28982 8870
rect 29226 9026 29302 9038
rect 29226 8974 29238 9026
rect 29290 8974 29302 9026
rect 29226 8922 29302 8974
rect 29226 8870 29238 8922
rect 29290 8870 29302 8922
rect 29226 8858 29302 8870
rect 29386 9028 29462 9038
rect 29386 8972 29396 9028
rect 29452 8972 29462 9028
rect 29386 8924 29462 8972
rect 29386 8868 29396 8924
rect 29452 8868 29462 8924
rect 29386 8858 29462 8868
rect 28186 8697 28262 8707
rect 28186 8641 28196 8697
rect 28252 8641 28262 8697
rect 28186 8631 28262 8641
rect 28426 8486 28502 8496
rect 28426 8430 28436 8486
rect 28492 8430 28502 8486
rect 28426 8382 28502 8430
rect 28426 8326 28436 8382
rect 28492 8326 28502 8382
rect 28426 8316 28502 8326
rect 28596 8102 28652 8858
rect 28916 8102 28972 8858
rect 29066 8486 29142 8496
rect 29066 8430 29076 8486
rect 29132 8430 29142 8486
rect 29066 8382 29142 8430
rect 29066 8326 29076 8382
rect 29132 8326 29142 8382
rect 29066 8316 29142 8326
rect 29236 8102 29292 8858
rect 30569 8196 30853 9262
rect 30569 8140 30579 8196
rect 30635 8140 30683 8196
rect 30739 8140 30787 8196
rect 30843 8140 30853 8196
rect 28106 8092 28182 8102
rect 28106 8036 28116 8092
rect 28172 8036 28182 8092
rect 28106 7988 28182 8036
rect 28106 7932 28116 7988
rect 28172 7932 28182 7988
rect 28106 7922 28182 7932
rect 28266 8090 28342 8102
rect 28266 8038 28278 8090
rect 28330 8038 28342 8090
rect 28266 7986 28342 8038
rect 28266 7934 28278 7986
rect 28330 7934 28342 7986
rect 28266 7922 28342 7934
rect 28586 8090 28662 8102
rect 28586 8038 28598 8090
rect 28650 8038 28662 8090
rect 28586 7986 28662 8038
rect 28586 7934 28598 7986
rect 28650 7934 28662 7986
rect 28586 7922 28662 7934
rect 28746 8092 28822 8102
rect 28746 8036 28756 8092
rect 28812 8036 28822 8092
rect 28746 7988 28822 8036
rect 28746 7932 28756 7988
rect 28812 7932 28822 7988
rect 28746 7922 28822 7932
rect 28906 8090 28982 8102
rect 28906 8038 28918 8090
rect 28970 8038 28982 8090
rect 28906 7986 28982 8038
rect 28906 7934 28918 7986
rect 28970 7934 28982 7986
rect 28906 7922 28982 7934
rect 29226 8090 29302 8102
rect 29226 8038 29238 8090
rect 29290 8038 29302 8090
rect 29226 7986 29302 8038
rect 29226 7934 29238 7986
rect 29290 7934 29302 7986
rect 29226 7922 29302 7934
rect 29386 8092 29462 8102
rect 29386 8036 29396 8092
rect 29452 8036 29462 8092
rect 29386 7988 29462 8036
rect 29386 7932 29396 7988
rect 29452 7932 29462 7988
rect 29386 7922 29462 7932
rect 30569 8092 30853 8140
rect 30569 8036 30579 8092
rect 30635 8036 30683 8092
rect 30739 8036 30787 8092
rect 30843 8036 30853 8092
rect 30569 7988 30853 8036
rect 30569 7932 30579 7988
rect 30635 7932 30683 7988
rect 30739 7932 30787 7988
rect 30843 7932 30853 7988
rect 30569 7922 30853 7932
rect 31218 11940 31502 13006
rect 32132 15119 32416 15131
rect 32132 15067 32144 15119
rect 32196 15067 32248 15119
rect 32300 15067 32352 15119
rect 32404 15067 32416 15119
rect 32132 15015 32416 15067
rect 32132 14963 32144 15015
rect 32196 14963 32248 15015
rect 32300 14963 32352 15015
rect 32404 14963 32416 15015
rect 32132 14911 32416 14963
rect 32132 14859 32144 14911
rect 32196 14859 32248 14911
rect 32300 14859 32352 14911
rect 32404 14859 32416 14911
rect 32132 14847 32416 14859
rect 32132 12886 32410 14847
rect 31218 11884 31228 11940
rect 31284 11884 31332 11940
rect 31388 11884 31436 11940
rect 31492 11884 31502 11940
rect 31218 11836 31502 11884
rect 31218 11780 31228 11836
rect 31284 11780 31332 11836
rect 31388 11780 31436 11836
rect 31492 11780 31502 11836
rect 32126 12876 32410 12886
rect 32126 12820 32136 12876
rect 32192 12820 32240 12876
rect 32296 12820 32344 12876
rect 32400 12820 32410 12876
rect 32126 12772 32410 12820
rect 34578 13050 34862 13060
rect 34578 12994 34588 13050
rect 34644 12994 34692 13050
rect 34748 12994 34796 13050
rect 34852 12994 34862 13050
rect 34578 12946 34862 12994
rect 34578 12890 34588 12946
rect 34644 12890 34692 12946
rect 34748 12890 34796 12946
rect 34852 12890 34862 12946
rect 34578 12842 34862 12890
rect 34578 12786 34588 12842
rect 34644 12786 34692 12842
rect 34748 12786 34796 12842
rect 34852 12786 34862 12842
rect 34578 12776 34862 12786
rect 38714 13050 38998 13060
rect 38714 12994 38724 13050
rect 38780 12994 38828 13050
rect 38884 12994 38932 13050
rect 38988 12994 38998 13050
rect 38714 12946 38998 12994
rect 38714 12890 38724 12946
rect 38780 12890 38828 12946
rect 38884 12890 38932 12946
rect 38988 12890 38998 12946
rect 38714 12842 38998 12890
rect 38714 12786 38724 12842
rect 38780 12786 38828 12842
rect 38884 12786 38932 12842
rect 38988 12786 38998 12842
rect 38714 12776 38998 12786
rect 44274 13050 44558 13060
rect 44274 12994 44284 13050
rect 44340 12994 44388 13050
rect 44444 12994 44492 13050
rect 44548 12994 44558 13050
rect 44274 12946 44558 12994
rect 44274 12890 44284 12946
rect 44340 12890 44388 12946
rect 44444 12890 44492 12946
rect 44548 12890 44558 12946
rect 44274 12842 44558 12890
rect 44274 12786 44284 12842
rect 44340 12786 44388 12842
rect 44444 12786 44492 12842
rect 44548 12786 44558 12842
rect 44274 12776 44558 12786
rect 48410 13050 48694 13060
rect 48410 12994 48420 13050
rect 48476 12994 48524 13050
rect 48580 12994 48628 13050
rect 48684 12994 48694 13050
rect 48410 12946 48694 12994
rect 48410 12890 48420 12946
rect 48476 12890 48524 12946
rect 48580 12890 48628 12946
rect 48684 12890 48694 12946
rect 48410 12842 48694 12890
rect 48410 12786 48420 12842
rect 48476 12786 48524 12842
rect 48580 12786 48628 12842
rect 48684 12786 48694 12842
rect 48410 12776 48694 12786
rect 53970 13050 54254 13060
rect 53970 12994 53980 13050
rect 54036 12994 54084 13050
rect 54140 12994 54188 13050
rect 54244 12994 54254 13050
rect 53970 12946 54254 12994
rect 53970 12890 53980 12946
rect 54036 12890 54084 12946
rect 54140 12890 54188 12946
rect 54244 12890 54254 12946
rect 53970 12842 54254 12890
rect 53970 12786 53980 12842
rect 54036 12786 54084 12842
rect 54140 12786 54188 12842
rect 54244 12786 54254 12842
rect 53970 12776 54254 12786
rect 58106 13050 58390 13060
rect 58106 12994 58116 13050
rect 58172 12994 58220 13050
rect 58276 12994 58324 13050
rect 58380 12994 58390 13050
rect 58106 12946 58390 12994
rect 58106 12890 58116 12946
rect 58172 12890 58220 12946
rect 58276 12890 58324 12946
rect 58380 12890 58390 12946
rect 58106 12842 58390 12890
rect 58106 12786 58116 12842
rect 58172 12786 58220 12842
rect 58276 12786 58324 12842
rect 58380 12786 58390 12842
rect 58106 12776 58390 12786
rect 63666 13050 63950 13060
rect 63666 12994 63676 13050
rect 63732 12994 63780 13050
rect 63836 12994 63884 13050
rect 63940 12994 63950 13050
rect 63666 12946 63950 12994
rect 63666 12890 63676 12946
rect 63732 12890 63780 12946
rect 63836 12890 63884 12946
rect 63940 12890 63950 12946
rect 63666 12842 63950 12890
rect 63666 12786 63676 12842
rect 63732 12786 63780 12842
rect 63836 12786 63884 12842
rect 63940 12786 63950 12842
rect 63666 12776 63950 12786
rect 66914 13050 67198 13060
rect 66914 12994 66924 13050
rect 66980 12994 67028 13050
rect 67084 12994 67132 13050
rect 67188 12994 67198 13050
rect 66914 12946 67198 12994
rect 66914 12890 66924 12946
rect 66980 12890 67028 12946
rect 67084 12890 67132 12946
rect 67188 12890 67198 12946
rect 66914 12842 67198 12890
rect 66914 12786 66924 12842
rect 66980 12786 67028 12842
rect 67084 12786 67132 12842
rect 67188 12786 67198 12842
rect 66914 12776 67198 12786
rect 32126 12716 32136 12772
rect 32192 12716 32240 12772
rect 32296 12716 32344 12772
rect 32400 12716 32410 12772
rect 32126 12668 32410 12716
rect 32126 12612 32136 12668
rect 32192 12612 32240 12668
rect 32296 12612 32344 12668
rect 32400 12612 32410 12668
rect 32126 12334 32410 12612
rect 32126 12278 32136 12334
rect 32192 12278 32240 12334
rect 32296 12278 32344 12334
rect 32400 12278 32410 12334
rect 32126 12230 32410 12278
rect 32126 12174 32136 12230
rect 32192 12174 32240 12230
rect 32296 12174 32344 12230
rect 32400 12174 32410 12230
rect 32126 12126 32410 12174
rect 32126 12070 32136 12126
rect 32192 12070 32240 12126
rect 32296 12070 32344 12126
rect 32400 12070 32410 12126
rect 31218 11732 31502 11780
rect 31218 11676 31228 11732
rect 31284 11676 31332 11732
rect 31388 11676 31436 11732
rect 31492 11676 31502 11732
rect 31218 11398 31502 11676
rect 31218 11342 31228 11398
rect 31284 11342 31332 11398
rect 31388 11342 31436 11398
rect 31492 11342 31502 11398
rect 31218 11294 31502 11342
rect 31218 11238 31228 11294
rect 31284 11238 31332 11294
rect 31388 11238 31436 11294
rect 31492 11238 31502 11294
rect 31218 11190 31502 11238
rect 31218 11134 31228 11190
rect 31284 11134 31332 11190
rect 31388 11134 31436 11190
rect 31492 11134 31502 11190
rect 31218 10462 31502 11134
rect 31218 10406 31228 10462
rect 31284 10406 31332 10462
rect 31388 10406 31436 10462
rect 31492 10406 31502 10462
rect 31218 10358 31502 10406
rect 31218 10302 31228 10358
rect 31284 10302 31332 10358
rect 31388 10302 31436 10358
rect 31492 10302 31502 10358
rect 31218 10254 31502 10302
rect 31218 10198 31228 10254
rect 31284 10198 31332 10254
rect 31388 10198 31436 10254
rect 31492 10198 31502 10254
rect 31218 9132 31502 10198
rect 31218 9076 31228 9132
rect 31284 9076 31332 9132
rect 31388 9076 31436 9132
rect 31492 9076 31502 9132
rect 31218 9028 31502 9076
rect 31218 8972 31228 9028
rect 31284 8972 31332 9028
rect 31388 8972 31436 9028
rect 31492 8972 31502 9028
rect 31218 8924 31502 8972
rect 31218 8868 31228 8924
rect 31284 8868 31332 8924
rect 31388 8868 31436 8924
rect 31492 8868 31502 8924
rect 31218 8590 31502 8868
rect 31218 8534 31228 8590
rect 31284 8534 31332 8590
rect 31388 8534 31436 8590
rect 31492 8534 31502 8590
rect 31218 8486 31502 8534
rect 31218 8430 31228 8486
rect 31284 8430 31332 8486
rect 31388 8430 31436 8486
rect 31492 8430 31502 8486
rect 31218 8382 31502 8430
rect 31218 8326 31228 8382
rect 31284 8326 31332 8382
rect 31388 8326 31436 8382
rect 31492 8326 31502 8382
rect 26962 7705 26972 7761
rect 27028 7705 27038 7761
rect 26962 7695 27038 7705
rect 28346 7761 28422 7771
rect 28346 7705 28356 7761
rect 28412 7705 28422 7761
rect 28346 7695 28422 7705
rect 17365 7665 17545 7675
rect 17119 6438 17403 6448
rect 17119 6382 17129 6438
rect 17185 6382 17233 6438
rect 17289 6382 17337 6438
rect 17393 6382 17403 6438
rect 17119 6334 17403 6382
rect 17119 6278 17129 6334
rect 17185 6278 17233 6334
rect 17289 6278 17337 6334
rect 17393 6278 17403 6334
rect 17119 6230 17403 6278
rect 17119 6174 17129 6230
rect 17185 6174 17233 6230
rect 17289 6174 17337 6230
rect 17393 6174 17403 6230
rect 17119 6164 17403 6174
rect 30288 6438 30780 6448
rect 30288 6382 30298 6438
rect 30354 6382 30402 6438
rect 30458 6382 30506 6438
rect 30562 6382 30610 6438
rect 30666 6382 30714 6438
rect 30770 6382 30780 6438
rect 30288 6334 30780 6382
rect 30288 6278 30298 6334
rect 30354 6278 30402 6334
rect 30458 6278 30506 6334
rect 30562 6278 30610 6334
rect 30666 6278 30714 6334
rect 30770 6278 30780 6334
rect 30288 6230 30780 6278
rect 30288 6174 30298 6230
rect 30354 6174 30402 6230
rect 30458 6174 30506 6230
rect 30562 6174 30610 6230
rect 30666 6174 30714 6230
rect 30770 6174 30780 6230
rect 17556 6096 17840 6106
rect 17556 6040 17566 6096
rect 17622 6040 17670 6096
rect 17726 6040 17774 6096
rect 17830 6040 17840 6096
rect 17556 5992 17840 6040
rect 17556 5936 17566 5992
rect 17622 5936 17670 5992
rect 17726 5936 17774 5992
rect 17830 5936 17840 5992
rect 17556 5888 17840 5936
rect 17556 5832 17566 5888
rect 17622 5832 17670 5888
rect 17726 5832 17774 5888
rect 17830 5832 17840 5888
rect 17556 5822 17840 5832
rect 29728 6096 30220 6106
rect 29728 6040 29738 6096
rect 29794 6040 29842 6096
rect 29898 6040 29946 6096
rect 30002 6040 30050 6096
rect 30106 6040 30154 6096
rect 30210 6040 30220 6096
rect 29728 5992 30220 6040
rect 29728 5936 29738 5992
rect 29794 5936 29842 5992
rect 29898 5936 29946 5992
rect 30002 5936 30050 5992
rect 30106 5936 30154 5992
rect 30210 5936 30220 5992
rect 29728 5888 30220 5936
rect 29728 5832 29738 5888
rect 29794 5832 29842 5888
rect 29898 5832 29946 5888
rect 30002 5832 30050 5888
rect 30106 5832 30154 5888
rect 30210 5832 30220 5888
rect 14686 5711 14866 5721
rect 14686 5655 14696 5711
rect 14752 5655 14800 5711
rect 14856 5655 14866 5711
rect 14686 5607 14866 5655
rect 14686 5551 14696 5607
rect 14752 5551 14800 5607
rect 14856 5551 14866 5607
rect 14686 5541 14866 5551
rect 17334 5446 17514 5456
rect 17334 5390 17344 5446
rect 17400 5390 17448 5446
rect 17504 5390 17514 5446
rect 17334 5342 17514 5390
rect 17334 5286 17344 5342
rect 17400 5286 17448 5342
rect 17504 5286 17514 5342
rect 17334 5276 17514 5286
rect 24120 5446 24300 5456
rect 24120 5390 24130 5446
rect 24186 5390 24234 5446
rect 24290 5390 24300 5446
rect 24120 5342 24300 5390
rect 24120 5286 24130 5342
rect 24186 5286 24234 5342
rect 24290 5286 24300 5342
rect 24120 5276 24300 5286
rect 24130 5025 24290 5276
rect 24118 5013 24298 5025
rect 24118 4961 24130 5013
rect 24182 4961 24234 5013
rect 24286 4961 24298 5013
rect 20570 4918 20854 4930
rect 20570 4866 20659 4918
rect 20711 4866 20763 4918
rect 20815 4866 20854 4918
rect 14212 4466 14496 4476
rect 14212 4410 14222 4466
rect 14278 4410 14326 4466
rect 14382 4410 14430 4466
rect 14486 4410 14496 4466
rect 14212 4362 14496 4410
rect 14212 4306 14222 4362
rect 14278 4306 14326 4362
rect 14382 4306 14430 4362
rect 14486 4306 14496 4362
rect 14212 4258 14496 4306
rect 14212 4202 14222 4258
rect 14278 4202 14326 4258
rect 14382 4202 14430 4258
rect 14486 4202 14496 4258
rect 13100 2296 13176 2306
rect 13100 2240 13110 2296
rect 13166 2240 13176 2296
rect 13100 2192 13176 2240
rect 13100 2136 13110 2192
rect 13166 2136 13176 2192
rect 13100 2088 13176 2136
rect 13100 2032 13110 2088
rect 13166 2032 13176 2088
rect 13100 2022 13176 2032
rect 14212 1835 14496 4202
rect 15052 3564 15128 3574
rect 15052 3508 15062 3564
rect 15118 3508 15128 3564
rect 15052 3460 15128 3508
rect 15052 3404 15062 3460
rect 15118 3404 15128 3460
rect 15052 3394 15128 3404
rect 15660 3564 15736 3574
rect 15660 3508 15670 3564
rect 15726 3508 15736 3564
rect 15660 3460 15736 3508
rect 15660 3404 15670 3460
rect 15726 3404 15736 3460
rect 15660 3394 15736 3404
rect 16268 3564 16344 3574
rect 16268 3508 16278 3564
rect 16334 3508 16344 3564
rect 16268 3460 16344 3508
rect 16268 3404 16278 3460
rect 16334 3404 16344 3460
rect 16268 3394 16344 3404
rect 15556 3164 15840 3174
rect 15556 3108 15566 3164
rect 15622 3108 15670 3164
rect 15726 3108 15774 3164
rect 15830 3108 15840 3164
rect 15556 3060 15840 3108
rect 15556 3004 15566 3060
rect 15622 3004 15670 3060
rect 15726 3004 15774 3060
rect 15830 3004 15840 3060
rect 15556 2956 15840 3004
rect 15556 2900 15566 2956
rect 15622 2900 15670 2956
rect 15726 2900 15774 2956
rect 15830 2900 15840 2956
rect 13200 1815 13380 1827
rect 13200 1763 13212 1815
rect 13264 1763 13316 1815
rect 13368 1763 13380 1815
rect 14212 1783 14224 1835
rect 14276 1783 14328 1835
rect 14380 1783 14432 1835
rect 14484 1783 14496 1835
rect 14212 1771 14496 1783
rect 14889 2296 15173 2306
rect 14889 2240 14899 2296
rect 14955 2240 15003 2296
rect 15059 2240 15107 2296
rect 15163 2240 15173 2296
rect 14889 2192 15173 2240
rect 14889 2136 14899 2192
rect 14955 2136 15003 2192
rect 15059 2136 15107 2192
rect 15163 2136 15173 2192
rect 14889 2088 15173 2136
rect 14889 2032 14899 2088
rect 14955 2032 15003 2088
rect 15059 2032 15107 2088
rect 15163 2032 15173 2088
rect 13200 1711 13380 1763
rect 13200 1659 13212 1711
rect 13264 1659 13316 1711
rect 13368 1659 13380 1711
rect 12018 1129 12198 1139
rect 12018 1073 12028 1129
rect 12084 1073 12132 1129
rect 12188 1073 12198 1129
rect 12018 1025 12198 1073
rect 12018 969 12028 1025
rect 12084 969 12132 1025
rect 12188 969 12198 1025
rect 12018 959 12198 969
rect 5620 877 5800 887
rect 5620 821 5630 877
rect 5686 821 5734 877
rect 5790 821 5800 877
rect 5620 773 5800 821
rect 5620 717 5630 773
rect 5686 717 5734 773
rect 5790 717 5800 773
rect 5620 707 5800 717
rect 10313 877 10493 887
rect 10313 821 10323 877
rect 10379 821 10427 877
rect 10483 821 10493 877
rect 10313 773 10493 821
rect 10313 717 10323 773
rect 10379 717 10427 773
rect 10483 717 10493 773
rect 10313 707 10493 717
rect 5144 557 5324 567
rect 5144 501 5154 557
rect 5210 501 5258 557
rect 5314 501 5324 557
rect 5144 453 5324 501
rect 5144 397 5154 453
rect 5210 397 5258 453
rect 5314 397 5324 453
rect 5144 387 5324 397
rect 13200 557 13380 1659
rect 13200 501 13210 557
rect 13266 501 13314 557
rect 13370 501 13380 557
rect 13200 453 13380 501
rect 14889 774 15173 2032
rect 14889 718 14899 774
rect 14955 718 15003 774
rect 15059 718 15107 774
rect 15163 718 15173 774
rect 14889 670 15173 718
rect 14889 614 14899 670
rect 14955 614 15003 670
rect 15059 614 15107 670
rect 15163 614 15173 670
rect 14889 566 15173 614
rect 14889 510 14899 566
rect 14955 510 15003 566
rect 15059 510 15107 566
rect 15163 510 15173 566
rect 14889 500 15173 510
rect 15556 2296 15840 2900
rect 20570 3164 20854 4866
rect 24118 4909 24298 4961
rect 24118 4857 24130 4909
rect 24182 4857 24234 4909
rect 24286 4857 24298 4909
rect 24118 4845 24298 4857
rect 21660 4466 21736 4476
rect 21660 4410 21670 4466
rect 21726 4410 21736 4466
rect 21660 4362 21736 4410
rect 21660 4306 21670 4362
rect 21726 4306 21736 4362
rect 21660 4258 21736 4306
rect 21660 4202 21670 4258
rect 21726 4202 21736 4258
rect 21660 4192 21736 4202
rect 27480 4305 27660 4317
rect 27480 4253 27492 4305
rect 27544 4253 27596 4305
rect 27648 4253 27660 4305
rect 27480 4201 27660 4253
rect 27480 4149 27492 4201
rect 27544 4149 27596 4201
rect 27648 4149 27660 4201
rect 20570 3108 20580 3164
rect 20636 3108 20684 3164
rect 20740 3108 20788 3164
rect 20844 3108 20854 3164
rect 20570 3060 20854 3108
rect 20570 3004 20580 3060
rect 20636 3004 20684 3060
rect 20740 3004 20788 3060
rect 20844 3004 20854 3060
rect 20570 2956 20854 3004
rect 20570 2900 20580 2956
rect 20636 2900 20684 2956
rect 20740 2900 20788 2956
rect 20844 2900 20854 2956
rect 20570 2890 20854 2900
rect 27478 2937 27660 4149
rect 27478 2885 27490 2937
rect 27542 2885 27594 2937
rect 27646 2935 27660 2937
rect 29728 3081 30220 5832
rect 30288 5093 30780 6174
rect 30288 5041 30300 5093
rect 30352 5041 30404 5093
rect 30456 5041 30508 5093
rect 30560 5041 30612 5093
rect 30664 5041 30716 5093
rect 30768 5041 30780 5093
rect 30288 4989 30780 5041
rect 30288 4937 30300 4989
rect 30352 4937 30404 4989
rect 30456 4937 30508 4989
rect 30560 4937 30612 4989
rect 30664 4937 30716 4989
rect 30768 4937 30780 4989
rect 30288 4885 30780 4937
rect 30288 4833 30300 4885
rect 30352 4833 30404 4885
rect 30456 4833 30508 4885
rect 30560 4833 30612 4885
rect 30664 4833 30716 4885
rect 30768 4833 30780 4885
rect 30288 4821 30780 4833
rect 30288 4139 30780 4149
rect 30288 4083 30298 4139
rect 30354 4083 30402 4139
rect 30458 4083 30506 4139
rect 30562 4083 30610 4139
rect 30666 4083 30714 4139
rect 30770 4083 30780 4139
rect 30288 4035 30780 4083
rect 30288 3979 30298 4035
rect 30354 3979 30402 4035
rect 30458 3979 30506 4035
rect 30562 3979 30610 4035
rect 30666 3979 30714 4035
rect 30770 3979 30780 4035
rect 30288 3931 30780 3979
rect 30288 3875 30298 3931
rect 30354 3875 30402 3931
rect 30458 3875 30506 3931
rect 30562 3875 30610 3931
rect 30666 3875 30714 3931
rect 30770 3875 30780 3931
rect 30288 3827 30780 3875
rect 30288 3771 30298 3827
rect 30354 3771 30402 3827
rect 30458 3771 30506 3827
rect 30562 3771 30610 3827
rect 30666 3771 30714 3827
rect 30770 3771 30780 3827
rect 30288 3723 30780 3771
rect 30288 3667 30298 3723
rect 30354 3667 30402 3723
rect 30458 3667 30506 3723
rect 30562 3667 30610 3723
rect 30666 3667 30714 3723
rect 30770 3667 30780 3723
rect 30288 3657 30780 3667
rect 29728 3029 29740 3081
rect 29792 3029 29844 3081
rect 29896 3029 29948 3081
rect 30000 3029 30052 3081
rect 30104 3029 30156 3081
rect 30208 3029 30220 3081
rect 29728 2977 30220 3029
rect 27646 2885 27658 2935
rect 27478 2833 27658 2885
rect 15556 2240 15566 2296
rect 15622 2240 15670 2296
rect 15726 2240 15774 2296
rect 15830 2240 15840 2296
rect 15556 2192 15840 2240
rect 15556 2136 15566 2192
rect 15622 2136 15670 2192
rect 15726 2136 15774 2192
rect 15830 2136 15840 2192
rect 15556 2088 15840 2136
rect 15556 2032 15566 2088
rect 15622 2032 15670 2088
rect 15726 2032 15774 2088
rect 15830 2032 15840 2088
rect 13200 397 13210 453
rect 13266 397 13314 453
rect 13370 397 13380 453
rect 13200 387 13380 397
rect 15556 272 15840 2032
rect 16171 2763 16455 2785
rect 27478 2781 27490 2833
rect 27542 2781 27594 2833
rect 27646 2781 27658 2833
rect 29728 2925 29740 2977
rect 29792 2925 29844 2977
rect 29896 2925 29948 2977
rect 30000 2925 30052 2977
rect 30104 2925 30156 2977
rect 30208 2925 30220 2977
rect 29728 2873 30220 2925
rect 29728 2821 29740 2873
rect 29792 2821 29844 2873
rect 29896 2821 29948 2873
rect 30000 2821 30052 2873
rect 30104 2821 30156 2873
rect 30208 2821 30220 2873
rect 29728 2809 30220 2821
rect 27478 2769 27658 2781
rect 16171 2711 16183 2763
rect 16235 2711 16287 2763
rect 16339 2711 16391 2763
rect 16443 2711 16455 2763
rect 16171 2659 16455 2711
rect 16171 2607 16183 2659
rect 16235 2607 16287 2659
rect 16339 2607 16391 2659
rect 16443 2607 16455 2659
rect 16171 2258 16455 2607
rect 16171 2202 16181 2258
rect 16237 2202 16285 2258
rect 16341 2202 16389 2258
rect 16445 2202 16455 2258
rect 16171 2154 16455 2202
rect 16171 2098 16181 2154
rect 16237 2098 16285 2154
rect 16341 2098 16389 2154
rect 16445 2098 16455 2154
rect 16171 2050 16455 2098
rect 16171 1994 16181 2050
rect 16237 1994 16285 2050
rect 16341 1994 16389 2050
rect 16445 1994 16455 2050
rect 16171 1984 16455 1994
rect 19100 2258 19176 2268
rect 19100 2202 19110 2258
rect 19166 2202 19176 2258
rect 19100 2154 19176 2202
rect 19100 2098 19110 2154
rect 19166 2098 19176 2154
rect 19100 2050 19176 2098
rect 19100 1994 19110 2050
rect 19166 1994 19176 2050
rect 19100 1984 19176 1994
rect 19420 2258 19496 2268
rect 19420 2202 19430 2258
rect 19486 2202 19496 2258
rect 19420 2154 19496 2202
rect 19420 2098 19430 2154
rect 19486 2098 19496 2154
rect 19420 2050 19496 2098
rect 19420 1994 19430 2050
rect 19486 1994 19496 2050
rect 19420 1984 19496 1994
rect 19740 2258 19816 2268
rect 19740 2202 19750 2258
rect 19806 2202 19816 2258
rect 19740 2154 19816 2202
rect 19740 2098 19750 2154
rect 19806 2098 19816 2154
rect 19740 2050 19816 2098
rect 19740 1994 19750 2050
rect 19806 1994 19816 2050
rect 19740 1984 19816 1994
rect 20060 2258 20136 2268
rect 20060 2202 20070 2258
rect 20126 2202 20136 2258
rect 20060 2154 20136 2202
rect 20060 2098 20070 2154
rect 20126 2098 20136 2154
rect 20060 2050 20136 2098
rect 20060 1994 20070 2050
rect 20126 1994 20136 2050
rect 20060 1984 20136 1994
rect 20380 2258 20456 2268
rect 20380 2202 20390 2258
rect 20446 2202 20456 2258
rect 20380 2154 20456 2202
rect 20380 2098 20390 2154
rect 20446 2098 20456 2154
rect 20380 2050 20456 2098
rect 20380 1994 20390 2050
rect 20446 1994 20456 2050
rect 20380 1984 20456 1994
rect 20700 2258 20776 2268
rect 20700 2202 20710 2258
rect 20766 2202 20776 2258
rect 20700 2154 20776 2202
rect 20700 2098 20710 2154
rect 20766 2098 20776 2154
rect 20700 2050 20776 2098
rect 20700 1994 20710 2050
rect 20766 1994 20776 2050
rect 20700 1984 20776 1994
rect 21020 2258 21096 2268
rect 21020 2202 21030 2258
rect 21086 2202 21096 2258
rect 21020 2154 21096 2202
rect 21020 2098 21030 2154
rect 21086 2098 21096 2154
rect 21020 2050 21096 2098
rect 21020 1994 21030 2050
rect 21086 1994 21096 2050
rect 21020 1984 21096 1994
rect 30288 2127 30780 2137
rect 30288 2071 30298 2127
rect 30354 2071 30402 2127
rect 30458 2071 30506 2127
rect 30562 2071 30610 2127
rect 30666 2071 30714 2127
rect 30770 2071 30780 2127
rect 30288 2023 30780 2071
rect 30288 1967 30298 2023
rect 30354 1967 30402 2023
rect 30458 1967 30506 2023
rect 30562 1967 30610 2023
rect 30666 1967 30714 2023
rect 30770 1967 30780 2023
rect 30288 1919 30780 1967
rect 21631 1904 21915 1916
rect 21631 1852 21643 1904
rect 21695 1852 21747 1904
rect 21799 1852 21851 1904
rect 21903 1852 21915 1904
rect 21631 774 21915 1852
rect 30288 1863 30298 1919
rect 30354 1863 30402 1919
rect 30458 1863 30506 1919
rect 30562 1863 30610 1919
rect 30666 1863 30714 1919
rect 30770 1863 30780 1919
rect 21631 718 21641 774
rect 21697 718 21745 774
rect 21801 718 21849 774
rect 21905 718 21915 774
rect 21631 670 21915 718
rect 21631 614 21641 670
rect 21697 614 21745 670
rect 21801 614 21849 670
rect 21905 614 21915 670
rect 21631 566 21915 614
rect 21631 510 21641 566
rect 21697 510 21745 566
rect 21801 510 21849 566
rect 21905 510 21915 566
rect 24118 1805 24298 1817
rect 24118 1753 24130 1805
rect 24182 1753 24234 1805
rect 24286 1753 24298 1805
rect 24118 1701 24298 1753
rect 24118 1649 24130 1701
rect 24182 1649 24234 1701
rect 24286 1649 24298 1701
rect 24118 787 24298 1649
rect 24118 731 24128 787
rect 24184 731 24232 787
rect 24288 731 24298 787
rect 24118 683 24298 731
rect 24118 627 24128 683
rect 24184 627 24232 683
rect 24288 627 24298 683
rect 24118 579 24298 627
rect 24118 523 24128 579
rect 24184 523 24232 579
rect 24288 523 24298 579
rect 24118 513 24298 523
rect 24568 1805 24748 1819
rect 24568 1753 24578 1805
rect 24630 1753 24682 1805
rect 24734 1753 24748 1805
rect 24568 1701 24748 1753
rect 24568 1649 24578 1701
rect 24630 1649 24682 1701
rect 24734 1649 24748 1701
rect 21631 500 21915 510
rect 15556 220 15568 272
rect 15620 220 15672 272
rect 15724 220 15776 272
rect 15828 220 15840 272
rect 15556 168 15840 220
rect 15556 116 15568 168
rect 15620 116 15672 168
rect 15724 116 15776 168
rect 15828 116 15840 168
rect 15556 64 15840 116
rect 24568 386 24748 1649
rect 30288 1815 30780 1863
rect 30288 1759 30298 1815
rect 30354 1759 30402 1815
rect 30458 1759 30506 1815
rect 30562 1759 30610 1815
rect 30666 1759 30714 1815
rect 30770 1759 30780 1815
rect 30288 1711 30780 1759
rect 30288 1655 30298 1711
rect 30354 1655 30402 1711
rect 30458 1655 30506 1711
rect 30562 1655 30610 1711
rect 30666 1655 30714 1711
rect 30770 1655 30780 1711
rect 30288 1645 30780 1655
rect 31218 787 31502 8326
rect 31746 11770 32030 11780
rect 31746 11714 31756 11770
rect 31812 11714 31860 11770
rect 31916 11714 31964 11770
rect 32020 11714 32030 11770
rect 31746 11666 32030 11714
rect 31746 11610 31756 11666
rect 31812 11610 31860 11666
rect 31916 11610 31964 11666
rect 32020 11610 32030 11666
rect 31746 11562 32030 11610
rect 31746 11506 31756 11562
rect 31812 11506 31860 11562
rect 31916 11506 31964 11562
rect 32020 11506 32030 11562
rect 31746 10316 32030 11506
rect 31746 10260 31756 10316
rect 31812 10260 31860 10316
rect 31916 10260 31964 10316
rect 32020 10260 32030 10316
rect 31746 10212 32030 10260
rect 31746 10156 31756 10212
rect 31812 10156 31860 10212
rect 31916 10156 31964 10212
rect 32020 10156 32030 10212
rect 31746 10108 32030 10156
rect 31746 10052 31756 10108
rect 31812 10052 31860 10108
rect 31916 10052 31964 10108
rect 32020 10052 32030 10108
rect 31746 9256 32030 10052
rect 31746 9200 31756 9256
rect 31812 9200 31860 9256
rect 31916 9200 31964 9256
rect 32020 9200 32030 9256
rect 31746 9152 32030 9200
rect 31746 9096 31756 9152
rect 31812 9096 31860 9152
rect 31916 9096 31964 9152
rect 32020 9096 32030 9152
rect 31746 9048 32030 9096
rect 31746 8992 31756 9048
rect 31812 8992 31860 9048
rect 31916 8992 31964 9048
rect 32020 8992 32030 9048
rect 31746 8590 32030 8992
rect 31746 8534 31756 8590
rect 31812 8534 31860 8590
rect 31916 8534 31964 8590
rect 32020 8534 32030 8590
rect 31746 8486 32030 8534
rect 31746 8430 31756 8486
rect 31812 8430 31860 8486
rect 31916 8430 31964 8486
rect 32020 8430 32030 8486
rect 31746 8382 32030 8430
rect 31746 8326 31756 8382
rect 31812 8326 31860 8382
rect 31916 8326 31964 8382
rect 32020 8326 32030 8382
rect 31746 8316 32030 8326
rect 32126 11376 32410 12070
rect 34602 11812 34838 12776
rect 34602 11760 34614 11812
rect 34666 11760 34774 11812
rect 34826 11760 34838 11812
rect 33723 11666 33799 11676
rect 33723 11610 33733 11666
rect 33789 11610 33799 11666
rect 33723 11562 33799 11610
rect 33723 11506 33733 11562
rect 33789 11506 33799 11562
rect 33723 11496 33799 11506
rect 34363 11666 34439 11676
rect 34363 11610 34373 11666
rect 34429 11610 34439 11666
rect 34363 11562 34439 11610
rect 34363 11506 34373 11562
rect 34429 11506 34439 11562
rect 34363 11496 34439 11506
rect 32126 11320 32136 11376
rect 32192 11320 32240 11376
rect 32296 11320 32344 11376
rect 32400 11320 32410 11376
rect 32126 11272 32410 11320
rect 32126 11216 32136 11272
rect 32192 11216 32240 11272
rect 32296 11216 32344 11272
rect 32400 11216 32410 11272
rect 32126 11168 32410 11216
rect 32126 11112 32136 11168
rect 32192 11112 32240 11168
rect 32296 11112 32344 11168
rect 32400 11112 32410 11168
rect 32126 10710 32410 11112
rect 33402 11272 33478 11282
rect 33402 11216 33412 11272
rect 33468 11216 33478 11272
rect 33402 11168 33478 11216
rect 33402 11112 33412 11168
rect 33468 11112 33478 11168
rect 33402 11102 33478 11112
rect 34042 11272 34118 11282
rect 34042 11216 34052 11272
rect 34108 11216 34118 11272
rect 34042 11168 34118 11216
rect 34042 11112 34052 11168
rect 34108 11112 34118 11168
rect 34042 11102 34118 11112
rect 32126 10654 32136 10710
rect 32192 10654 32240 10710
rect 32296 10654 32344 10710
rect 32400 10654 32410 10710
rect 32126 10606 32410 10654
rect 34602 10752 34838 11760
rect 38738 11812 38974 12776
rect 38738 11760 38750 11812
rect 38802 11760 38910 11812
rect 38962 11760 38974 11812
rect 44298 11812 44534 12776
rect 35003 11666 35079 11676
rect 35003 11610 35013 11666
rect 35069 11610 35079 11666
rect 35003 11562 35079 11610
rect 35003 11506 35013 11562
rect 35069 11506 35079 11562
rect 35003 11496 35079 11506
rect 35643 11666 35719 11676
rect 35643 11610 35653 11666
rect 35709 11610 35719 11666
rect 35643 11562 35719 11610
rect 35643 11506 35653 11562
rect 35709 11506 35719 11562
rect 35643 11496 35719 11506
rect 37857 11666 37933 11676
rect 37857 11610 37867 11666
rect 37923 11610 37933 11666
rect 37857 11562 37933 11610
rect 37857 11506 37867 11562
rect 37923 11506 37933 11562
rect 37857 11496 37933 11506
rect 38497 11666 38573 11676
rect 38497 11610 38507 11666
rect 38563 11610 38573 11666
rect 38497 11562 38573 11610
rect 38497 11506 38507 11562
rect 38563 11506 38573 11562
rect 38497 11496 38573 11506
rect 35322 11272 35398 11282
rect 35322 11216 35332 11272
rect 35388 11216 35398 11272
rect 35322 11168 35398 11216
rect 35322 11112 35332 11168
rect 35388 11112 35398 11168
rect 35322 11102 35398 11112
rect 35962 11272 36038 11282
rect 35962 11216 35972 11272
rect 36028 11216 36038 11272
rect 35962 11168 36038 11216
rect 35962 11112 35972 11168
rect 36028 11112 36038 11168
rect 35962 11102 36038 11112
rect 37538 11272 37614 11282
rect 37538 11216 37548 11272
rect 37604 11216 37614 11272
rect 37538 11168 37614 11216
rect 37538 11112 37548 11168
rect 37604 11112 37614 11168
rect 37538 11102 37614 11112
rect 38178 11272 38254 11282
rect 38178 11216 38188 11272
rect 38244 11216 38254 11272
rect 38178 11168 38254 11216
rect 38178 11112 38188 11168
rect 38244 11112 38254 11168
rect 38178 11102 38254 11112
rect 34602 10700 34614 10752
rect 34666 10700 34774 10752
rect 34826 10700 34838 10752
rect 32126 10550 32136 10606
rect 32192 10550 32240 10606
rect 32296 10550 32344 10606
rect 32400 10550 32410 10606
rect 32126 10502 32410 10550
rect 32126 10446 32136 10502
rect 32192 10446 32240 10502
rect 32296 10446 32344 10502
rect 32400 10446 32410 10502
rect 32126 9650 32410 10446
rect 33723 10606 33799 10616
rect 33723 10550 33733 10606
rect 33789 10550 33799 10606
rect 33723 10502 33799 10550
rect 33723 10446 33733 10502
rect 33789 10446 33799 10502
rect 33723 10436 33799 10446
rect 34363 10606 34439 10616
rect 34363 10550 34373 10606
rect 34429 10550 34439 10606
rect 34363 10502 34439 10550
rect 34363 10446 34373 10502
rect 34429 10446 34439 10502
rect 34363 10436 34439 10446
rect 33402 10212 33478 10222
rect 33402 10156 33412 10212
rect 33468 10156 33478 10212
rect 33402 10108 33478 10156
rect 33402 10052 33412 10108
rect 33468 10052 33478 10108
rect 33402 10042 33478 10052
rect 34042 10212 34118 10222
rect 34042 10156 34052 10212
rect 34108 10156 34118 10212
rect 34042 10108 34118 10156
rect 34042 10052 34052 10108
rect 34108 10052 34118 10108
rect 34042 10042 34118 10052
rect 32126 9594 32136 9650
rect 32192 9594 32240 9650
rect 32296 9594 32344 9650
rect 32400 9594 32410 9650
rect 32126 9546 32410 9594
rect 34602 9692 34838 10700
rect 38738 10752 38974 11760
rect 41473 11770 41757 11780
rect 41473 11714 41483 11770
rect 41539 11714 41587 11770
rect 41643 11714 41691 11770
rect 41747 11714 41757 11770
rect 39137 11666 39213 11676
rect 39137 11610 39147 11666
rect 39203 11610 39213 11666
rect 39137 11562 39213 11610
rect 39137 11506 39147 11562
rect 39203 11506 39213 11562
rect 39137 11496 39213 11506
rect 39777 11666 39853 11676
rect 39777 11610 39787 11666
rect 39843 11610 39853 11666
rect 39777 11562 39853 11610
rect 39777 11506 39787 11562
rect 39843 11506 39853 11562
rect 39777 11496 39853 11506
rect 41473 11666 41757 11714
rect 44298 11760 44310 11812
rect 44362 11760 44470 11812
rect 44522 11760 44534 11812
rect 41473 11610 41483 11666
rect 41539 11610 41587 11666
rect 41643 11610 41691 11666
rect 41747 11610 41757 11666
rect 41473 11562 41757 11610
rect 41473 11506 41483 11562
rect 41539 11506 41587 11562
rect 41643 11506 41691 11562
rect 41747 11506 41757 11562
rect 41112 11376 41396 11386
rect 41112 11320 41122 11376
rect 41178 11320 41226 11376
rect 41282 11320 41330 11376
rect 41386 11320 41396 11376
rect 39458 11272 39534 11282
rect 39458 11216 39468 11272
rect 39524 11216 39534 11272
rect 39458 11168 39534 11216
rect 39458 11112 39468 11168
rect 39524 11112 39534 11168
rect 39458 11102 39534 11112
rect 40098 11272 40174 11282
rect 40098 11216 40108 11272
rect 40164 11216 40174 11272
rect 40098 11168 40174 11216
rect 40098 11112 40108 11168
rect 40164 11112 40174 11168
rect 40098 11102 40174 11112
rect 41112 11272 41396 11320
rect 41112 11216 41122 11272
rect 41178 11216 41226 11272
rect 41282 11216 41330 11272
rect 41386 11216 41396 11272
rect 41112 11168 41396 11216
rect 41112 11112 41122 11168
rect 41178 11112 41226 11168
rect 41282 11112 41330 11168
rect 41386 11112 41396 11168
rect 38738 10700 38750 10752
rect 38802 10700 38910 10752
rect 38962 10700 38974 10752
rect 35003 10606 35079 10616
rect 35003 10550 35013 10606
rect 35069 10550 35079 10606
rect 35003 10502 35079 10550
rect 35003 10446 35013 10502
rect 35069 10446 35079 10502
rect 35003 10436 35079 10446
rect 35643 10606 35719 10616
rect 35643 10550 35653 10606
rect 35709 10550 35719 10606
rect 35643 10502 35719 10550
rect 35643 10446 35653 10502
rect 35709 10446 35719 10502
rect 35643 10436 35719 10446
rect 37857 10606 37933 10616
rect 37857 10550 37867 10606
rect 37923 10550 37933 10606
rect 37857 10502 37933 10550
rect 37857 10446 37867 10502
rect 37923 10446 37933 10502
rect 37857 10436 37933 10446
rect 38497 10606 38573 10616
rect 38497 10550 38507 10606
rect 38563 10550 38573 10606
rect 38497 10502 38573 10550
rect 38497 10446 38507 10502
rect 38563 10446 38573 10502
rect 38497 10436 38573 10446
rect 35322 10212 35398 10222
rect 35322 10156 35332 10212
rect 35388 10156 35398 10212
rect 35322 10108 35398 10156
rect 35322 10052 35332 10108
rect 35388 10052 35398 10108
rect 35322 10042 35398 10052
rect 35962 10212 36038 10222
rect 35962 10156 35972 10212
rect 36028 10156 36038 10212
rect 35962 10108 36038 10156
rect 35962 10052 35972 10108
rect 36028 10052 36038 10108
rect 35962 10042 36038 10052
rect 37538 10212 37614 10222
rect 37538 10156 37548 10212
rect 37604 10156 37614 10212
rect 37538 10108 37614 10156
rect 37538 10052 37548 10108
rect 37604 10052 37614 10108
rect 37538 10042 37614 10052
rect 38178 10212 38254 10222
rect 38178 10156 38188 10212
rect 38244 10156 38254 10212
rect 38178 10108 38254 10156
rect 38178 10052 38188 10108
rect 38244 10052 38254 10108
rect 38178 10042 38254 10052
rect 34602 9640 34614 9692
rect 34666 9640 34774 9692
rect 34826 9640 34838 9692
rect 32126 9490 32136 9546
rect 32192 9490 32240 9546
rect 32296 9490 32344 9546
rect 32400 9490 32410 9546
rect 32126 9442 32410 9490
rect 32126 9386 32136 9442
rect 32192 9386 32240 9442
rect 32296 9386 32344 9442
rect 32400 9386 32410 9442
rect 31218 731 31228 787
rect 31284 731 31332 787
rect 31388 731 31436 787
rect 31492 731 31502 787
rect 31218 683 31502 731
rect 31218 627 31228 683
rect 31284 627 31332 683
rect 31388 627 31436 683
rect 31492 627 31502 683
rect 31218 579 31502 627
rect 31218 523 31228 579
rect 31284 523 31332 579
rect 31388 523 31436 579
rect 31492 523 31502 579
rect 31218 513 31502 523
rect 32126 8196 32410 9386
rect 33723 9546 33799 9556
rect 33723 9490 33733 9546
rect 33789 9490 33799 9546
rect 33723 9442 33799 9490
rect 33723 9386 33733 9442
rect 33789 9386 33799 9442
rect 33723 9376 33799 9386
rect 34363 9546 34439 9556
rect 34363 9490 34373 9546
rect 34429 9490 34439 9546
rect 34363 9442 34439 9490
rect 34363 9386 34373 9442
rect 34429 9386 34439 9442
rect 34363 9376 34439 9386
rect 33402 9152 33478 9162
rect 33402 9096 33412 9152
rect 33468 9096 33478 9152
rect 33402 9048 33478 9096
rect 33402 8992 33412 9048
rect 33468 8992 33478 9048
rect 33402 8982 33478 8992
rect 34042 9152 34118 9162
rect 34042 9096 34052 9152
rect 34108 9096 34118 9152
rect 34042 9048 34118 9096
rect 34042 8992 34052 9048
rect 34108 8992 34118 9048
rect 34042 8982 34118 8992
rect 34602 8632 34838 9640
rect 38738 9692 38974 10700
rect 41112 10710 41396 11112
rect 41112 10654 41122 10710
rect 41178 10654 41226 10710
rect 41282 10654 41330 10710
rect 41386 10654 41396 10710
rect 39137 10606 39213 10616
rect 39137 10550 39147 10606
rect 39203 10550 39213 10606
rect 39137 10502 39213 10550
rect 39137 10446 39147 10502
rect 39203 10446 39213 10502
rect 39137 10436 39213 10446
rect 39777 10606 39853 10616
rect 39777 10550 39787 10606
rect 39843 10550 39853 10606
rect 39777 10502 39853 10550
rect 39777 10446 39787 10502
rect 39843 10446 39853 10502
rect 39777 10436 39853 10446
rect 41112 10606 41396 10654
rect 41112 10550 41122 10606
rect 41178 10550 41226 10606
rect 41282 10550 41330 10606
rect 41386 10550 41396 10606
rect 41112 10502 41396 10550
rect 41112 10446 41122 10502
rect 41178 10446 41226 10502
rect 41282 10446 41330 10502
rect 41386 10446 41396 10502
rect 39458 10212 39534 10222
rect 39458 10156 39468 10212
rect 39524 10156 39534 10212
rect 39458 10108 39534 10156
rect 39458 10052 39468 10108
rect 39524 10052 39534 10108
rect 39458 10042 39534 10052
rect 40098 10212 40174 10222
rect 40098 10156 40108 10212
rect 40164 10156 40174 10212
rect 40098 10108 40174 10156
rect 40098 10052 40108 10108
rect 40164 10052 40174 10108
rect 40098 10042 40174 10052
rect 38738 9640 38750 9692
rect 38802 9640 38910 9692
rect 38962 9640 38974 9692
rect 35003 9546 35079 9556
rect 35003 9490 35013 9546
rect 35069 9490 35079 9546
rect 35003 9442 35079 9490
rect 35003 9386 35013 9442
rect 35069 9386 35079 9442
rect 35003 9376 35079 9386
rect 35643 9546 35719 9556
rect 35643 9490 35653 9546
rect 35709 9490 35719 9546
rect 35643 9442 35719 9490
rect 35643 9386 35653 9442
rect 35709 9386 35719 9442
rect 35643 9376 35719 9386
rect 37857 9546 37933 9556
rect 37857 9490 37867 9546
rect 37923 9490 37933 9546
rect 37857 9442 37933 9490
rect 37857 9386 37867 9442
rect 37923 9386 37933 9442
rect 37857 9376 37933 9386
rect 38497 9546 38573 9556
rect 38497 9490 38507 9546
rect 38563 9490 38573 9546
rect 38497 9442 38573 9490
rect 38497 9386 38507 9442
rect 38563 9386 38573 9442
rect 38497 9376 38573 9386
rect 35322 9152 35398 9162
rect 35322 9096 35332 9152
rect 35388 9096 35398 9152
rect 35322 9048 35398 9096
rect 35322 8992 35332 9048
rect 35388 8992 35398 9048
rect 35322 8982 35398 8992
rect 35962 9152 36038 9162
rect 35962 9096 35972 9152
rect 36028 9096 36038 9152
rect 35962 9048 36038 9096
rect 35962 8992 35972 9048
rect 36028 8992 36038 9048
rect 35962 8982 36038 8992
rect 37538 9152 37614 9162
rect 37538 9096 37548 9152
rect 37604 9096 37614 9152
rect 37538 9048 37614 9096
rect 37538 8992 37548 9048
rect 37604 8992 37614 9048
rect 37538 8982 37614 8992
rect 38178 9152 38254 9162
rect 38178 9096 38188 9152
rect 38244 9096 38254 9152
rect 38178 9048 38254 9096
rect 38178 8992 38188 9048
rect 38244 8992 38254 9048
rect 38178 8982 38254 8992
rect 34602 8580 34614 8632
rect 34666 8580 34774 8632
rect 34826 8580 34838 8632
rect 33723 8486 33799 8496
rect 33723 8430 33733 8486
rect 33789 8430 33799 8486
rect 33723 8382 33799 8430
rect 33723 8326 33733 8382
rect 33789 8326 33799 8382
rect 33723 8316 33799 8326
rect 34363 8486 34439 8496
rect 34363 8430 34373 8486
rect 34429 8430 34439 8486
rect 34363 8382 34439 8430
rect 34363 8326 34373 8382
rect 34429 8326 34439 8382
rect 34363 8316 34439 8326
rect 32126 8140 32136 8196
rect 32192 8140 32240 8196
rect 32296 8140 32344 8196
rect 32400 8140 32410 8196
rect 32126 8092 32410 8140
rect 32126 8036 32136 8092
rect 32192 8036 32240 8092
rect 32296 8036 32344 8092
rect 32400 8036 32410 8092
rect 32126 7988 32410 8036
rect 32126 7932 32136 7988
rect 32192 7932 32240 7988
rect 32296 7932 32344 7988
rect 32400 7932 32410 7988
rect 24568 330 24578 386
rect 24634 330 24682 386
rect 24738 330 24748 386
rect 24568 282 24748 330
rect 24568 226 24578 282
rect 24634 226 24682 282
rect 24738 226 24748 282
rect 24568 178 24748 226
rect 24568 122 24578 178
rect 24634 122 24682 178
rect 24738 122 24748 178
rect 24568 112 24748 122
rect 32126 386 32410 7932
rect 33402 8092 33478 8102
rect 33402 8036 33412 8092
rect 33468 8036 33478 8092
rect 33402 7988 33478 8036
rect 33402 7932 33412 7988
rect 33468 7932 33478 7988
rect 33402 7922 33478 7932
rect 34042 8092 34118 8102
rect 34042 8036 34052 8092
rect 34108 8036 34118 8092
rect 34042 7988 34118 8036
rect 34042 7932 34052 7988
rect 34108 7932 34118 7988
rect 34042 7922 34118 7932
rect 34602 3564 34838 8580
rect 38738 8632 38974 9640
rect 41112 9650 41396 10446
rect 41112 9594 41122 9650
rect 41178 9594 41226 9650
rect 41282 9594 41330 9650
rect 41386 9594 41396 9650
rect 39137 9546 39213 9556
rect 39137 9490 39147 9546
rect 39203 9490 39213 9546
rect 39137 9442 39213 9490
rect 39137 9386 39147 9442
rect 39203 9386 39213 9442
rect 39137 9376 39213 9386
rect 39777 9546 39853 9556
rect 39777 9490 39787 9546
rect 39843 9490 39853 9546
rect 39777 9442 39853 9490
rect 39777 9386 39787 9442
rect 39843 9386 39853 9442
rect 39777 9376 39853 9386
rect 41112 9546 41396 9594
rect 41112 9490 41122 9546
rect 41178 9490 41226 9546
rect 41282 9490 41330 9546
rect 41386 9490 41396 9546
rect 41112 9442 41396 9490
rect 41112 9386 41122 9442
rect 41178 9386 41226 9442
rect 41282 9386 41330 9442
rect 41386 9386 41396 9442
rect 39458 9152 39534 9162
rect 39458 9096 39468 9152
rect 39524 9096 39534 9152
rect 39458 9048 39534 9096
rect 39458 8992 39468 9048
rect 39524 8992 39534 9048
rect 39458 8982 39534 8992
rect 40098 9152 40174 9162
rect 40098 9096 40108 9152
rect 40164 9096 40174 9152
rect 40098 9048 40174 9096
rect 40098 8992 40108 9048
rect 40164 8992 40174 9048
rect 40098 8982 40174 8992
rect 38738 8580 38750 8632
rect 38802 8580 38910 8632
rect 38962 8580 38974 8632
rect 38738 8568 38974 8580
rect 35003 8486 35079 8496
rect 35003 8430 35013 8486
rect 35069 8430 35079 8486
rect 35003 8382 35079 8430
rect 35003 8326 35013 8382
rect 35069 8326 35079 8382
rect 35003 8316 35079 8326
rect 35643 8486 35719 8496
rect 35643 8430 35653 8486
rect 35709 8430 35719 8486
rect 35643 8382 35719 8430
rect 35643 8326 35653 8382
rect 35709 8326 35719 8382
rect 35643 8316 35719 8326
rect 37857 8486 37933 8496
rect 37857 8430 37867 8486
rect 37923 8430 37933 8486
rect 37857 8382 37933 8430
rect 37857 8326 37867 8382
rect 37923 8326 37933 8382
rect 37857 8316 37933 8326
rect 38497 8486 38573 8496
rect 38497 8430 38507 8486
rect 38563 8430 38573 8486
rect 38497 8382 38573 8430
rect 38497 8326 38507 8382
rect 38563 8326 38573 8382
rect 38497 8316 38573 8326
rect 39137 8486 39213 8496
rect 39137 8430 39147 8486
rect 39203 8430 39213 8486
rect 39137 8382 39213 8430
rect 39137 8326 39147 8382
rect 39203 8326 39213 8382
rect 39137 8316 39213 8326
rect 39777 8486 39853 8496
rect 39777 8430 39787 8486
rect 39843 8430 39853 8486
rect 39777 8382 39853 8430
rect 39777 8326 39787 8382
rect 39843 8326 39853 8382
rect 39777 8316 39853 8326
rect 41112 8196 41396 9386
rect 41473 10316 41757 11506
rect 43419 11666 43495 11676
rect 43419 11610 43429 11666
rect 43485 11610 43495 11666
rect 43419 11562 43495 11610
rect 43419 11506 43429 11562
rect 43485 11506 43495 11562
rect 43419 11496 43495 11506
rect 44059 11666 44135 11676
rect 44059 11610 44069 11666
rect 44125 11610 44135 11666
rect 44059 11562 44135 11610
rect 44059 11506 44069 11562
rect 44125 11506 44135 11562
rect 44059 11496 44135 11506
rect 41473 10260 41483 10316
rect 41539 10260 41587 10316
rect 41643 10260 41691 10316
rect 41747 10260 41757 10316
rect 41473 10212 41757 10260
rect 41473 10156 41483 10212
rect 41539 10156 41587 10212
rect 41643 10156 41691 10212
rect 41747 10156 41757 10212
rect 41473 10108 41757 10156
rect 41473 10052 41483 10108
rect 41539 10052 41587 10108
rect 41643 10052 41691 10108
rect 41747 10052 41757 10108
rect 41473 9256 41757 10052
rect 41473 9200 41483 9256
rect 41539 9200 41587 9256
rect 41643 9200 41691 9256
rect 41747 9200 41757 9256
rect 41473 9152 41757 9200
rect 41473 9096 41483 9152
rect 41539 9096 41587 9152
rect 41643 9096 41691 9152
rect 41747 9096 41757 9152
rect 41473 9048 41757 9096
rect 41473 8992 41483 9048
rect 41539 8992 41587 9048
rect 41643 8992 41691 9048
rect 41747 8992 41757 9048
rect 41473 8590 41757 8992
rect 41473 8534 41483 8590
rect 41539 8534 41587 8590
rect 41643 8534 41691 8590
rect 41747 8534 41757 8590
rect 41473 8486 41757 8534
rect 41473 8430 41483 8486
rect 41539 8430 41587 8486
rect 41643 8430 41691 8486
rect 41747 8430 41757 8486
rect 41473 8382 41757 8430
rect 41473 8326 41483 8382
rect 41539 8326 41587 8382
rect 41643 8326 41691 8382
rect 41747 8326 41757 8382
rect 41473 8316 41757 8326
rect 41832 11376 42116 11386
rect 41832 11320 41842 11376
rect 41898 11320 41946 11376
rect 42002 11320 42050 11376
rect 42106 11320 42116 11376
rect 41832 11272 42116 11320
rect 41832 11216 41842 11272
rect 41898 11216 41946 11272
rect 42002 11216 42050 11272
rect 42106 11216 42116 11272
rect 41832 11168 42116 11216
rect 41832 11112 41842 11168
rect 41898 11112 41946 11168
rect 42002 11112 42050 11168
rect 42106 11112 42116 11168
rect 41832 10710 42116 11112
rect 43098 11272 43174 11282
rect 43098 11216 43108 11272
rect 43164 11216 43174 11272
rect 43098 11168 43174 11216
rect 43098 11112 43108 11168
rect 43164 11112 43174 11168
rect 43098 11102 43174 11112
rect 43738 11272 43814 11282
rect 43738 11216 43748 11272
rect 43804 11216 43814 11272
rect 43738 11168 43814 11216
rect 43738 11112 43748 11168
rect 43804 11112 43814 11168
rect 43738 11102 43814 11112
rect 41832 10654 41842 10710
rect 41898 10654 41946 10710
rect 42002 10654 42050 10710
rect 42106 10654 42116 10710
rect 41832 10606 42116 10654
rect 44298 10752 44534 11760
rect 48434 11812 48670 12776
rect 48434 11760 48446 11812
rect 48498 11760 48606 11812
rect 48658 11760 48670 11812
rect 53994 11812 54230 12776
rect 44699 11666 44775 11676
rect 44699 11610 44709 11666
rect 44765 11610 44775 11666
rect 44699 11562 44775 11610
rect 44699 11506 44709 11562
rect 44765 11506 44775 11562
rect 44699 11496 44775 11506
rect 45339 11666 45415 11676
rect 45339 11610 45349 11666
rect 45405 11610 45415 11666
rect 45339 11562 45415 11610
rect 45339 11506 45349 11562
rect 45405 11506 45415 11562
rect 45339 11496 45415 11506
rect 47553 11666 47629 11676
rect 47553 11610 47563 11666
rect 47619 11610 47629 11666
rect 47553 11562 47629 11610
rect 47553 11506 47563 11562
rect 47619 11506 47629 11562
rect 47553 11496 47629 11506
rect 48193 11666 48269 11676
rect 48193 11610 48203 11666
rect 48259 11610 48269 11666
rect 48193 11562 48269 11610
rect 48193 11506 48203 11562
rect 48259 11506 48269 11562
rect 48193 11496 48269 11506
rect 45018 11272 45094 11282
rect 45018 11216 45028 11272
rect 45084 11216 45094 11272
rect 45018 11168 45094 11216
rect 45018 11112 45028 11168
rect 45084 11112 45094 11168
rect 45018 11102 45094 11112
rect 45658 11272 45734 11282
rect 45658 11216 45668 11272
rect 45724 11216 45734 11272
rect 45658 11168 45734 11216
rect 45658 11112 45668 11168
rect 45724 11112 45734 11168
rect 45658 11102 45734 11112
rect 47234 11272 47310 11282
rect 47234 11216 47244 11272
rect 47300 11216 47310 11272
rect 47234 11168 47310 11216
rect 47234 11112 47244 11168
rect 47300 11112 47310 11168
rect 47234 11102 47310 11112
rect 47874 11272 47950 11282
rect 47874 11216 47884 11272
rect 47940 11216 47950 11272
rect 47874 11168 47950 11216
rect 47874 11112 47884 11168
rect 47940 11112 47950 11168
rect 47874 11102 47950 11112
rect 44298 10700 44310 10752
rect 44362 10700 44470 10752
rect 44522 10700 44534 10752
rect 41832 10550 41842 10606
rect 41898 10550 41946 10606
rect 42002 10550 42050 10606
rect 42106 10550 42116 10606
rect 41832 10502 42116 10550
rect 41832 10446 41842 10502
rect 41898 10446 41946 10502
rect 42002 10446 42050 10502
rect 42106 10446 42116 10502
rect 41832 9650 42116 10446
rect 43419 10606 43495 10616
rect 43419 10550 43429 10606
rect 43485 10550 43495 10606
rect 43419 10502 43495 10550
rect 43419 10446 43429 10502
rect 43485 10446 43495 10502
rect 43419 10436 43495 10446
rect 44059 10606 44135 10616
rect 44059 10550 44069 10606
rect 44125 10550 44135 10606
rect 44059 10502 44135 10550
rect 44059 10446 44069 10502
rect 44125 10446 44135 10502
rect 44059 10436 44135 10446
rect 43098 10212 43174 10222
rect 43098 10156 43108 10212
rect 43164 10156 43174 10212
rect 43098 10108 43174 10156
rect 43098 10052 43108 10108
rect 43164 10052 43174 10108
rect 43098 10042 43174 10052
rect 43738 10212 43814 10222
rect 43738 10156 43748 10212
rect 43804 10156 43814 10212
rect 43738 10108 43814 10156
rect 43738 10052 43748 10108
rect 43804 10052 43814 10108
rect 43738 10042 43814 10052
rect 41832 9594 41842 9650
rect 41898 9594 41946 9650
rect 42002 9594 42050 9650
rect 42106 9594 42116 9650
rect 41832 9546 42116 9594
rect 44298 9692 44534 10700
rect 48434 10752 48670 11760
rect 51128 11770 51412 11780
rect 51128 11714 51138 11770
rect 51194 11714 51242 11770
rect 51298 11714 51346 11770
rect 51402 11714 51412 11770
rect 48833 11666 48909 11676
rect 48833 11610 48843 11666
rect 48899 11610 48909 11666
rect 48833 11562 48909 11610
rect 48833 11506 48843 11562
rect 48899 11506 48909 11562
rect 48833 11496 48909 11506
rect 49473 11666 49549 11676
rect 49473 11610 49483 11666
rect 49539 11610 49549 11666
rect 49473 11562 49549 11610
rect 49473 11506 49483 11562
rect 49539 11506 49549 11562
rect 49473 11496 49549 11506
rect 51128 11666 51412 11714
rect 53994 11760 54006 11812
rect 54058 11760 54166 11812
rect 54218 11760 54230 11812
rect 51128 11610 51138 11666
rect 51194 11610 51242 11666
rect 51298 11610 51346 11666
rect 51402 11610 51412 11666
rect 51128 11562 51412 11610
rect 51128 11506 51138 11562
rect 51194 11506 51242 11562
rect 51298 11506 51346 11562
rect 51402 11506 51412 11562
rect 50788 11376 51072 11386
rect 50788 11320 50798 11376
rect 50854 11320 50902 11376
rect 50958 11320 51006 11376
rect 51062 11320 51072 11376
rect 49154 11272 49230 11282
rect 49154 11216 49164 11272
rect 49220 11216 49230 11272
rect 49154 11168 49230 11216
rect 49154 11112 49164 11168
rect 49220 11112 49230 11168
rect 49154 11102 49230 11112
rect 49794 11272 49870 11282
rect 49794 11216 49804 11272
rect 49860 11216 49870 11272
rect 49794 11168 49870 11216
rect 49794 11112 49804 11168
rect 49860 11112 49870 11168
rect 49794 11102 49870 11112
rect 50788 11272 51072 11320
rect 50788 11216 50798 11272
rect 50854 11216 50902 11272
rect 50958 11216 51006 11272
rect 51062 11216 51072 11272
rect 50788 11168 51072 11216
rect 50788 11112 50798 11168
rect 50854 11112 50902 11168
rect 50958 11112 51006 11168
rect 51062 11112 51072 11168
rect 48434 10700 48446 10752
rect 48498 10700 48606 10752
rect 48658 10700 48670 10752
rect 44699 10606 44775 10616
rect 44699 10550 44709 10606
rect 44765 10550 44775 10606
rect 44699 10502 44775 10550
rect 44699 10446 44709 10502
rect 44765 10446 44775 10502
rect 44699 10436 44775 10446
rect 45339 10606 45415 10616
rect 45339 10550 45349 10606
rect 45405 10550 45415 10606
rect 45339 10502 45415 10550
rect 45339 10446 45349 10502
rect 45405 10446 45415 10502
rect 45339 10436 45415 10446
rect 47553 10606 47629 10616
rect 47553 10550 47563 10606
rect 47619 10550 47629 10606
rect 47553 10502 47629 10550
rect 47553 10446 47563 10502
rect 47619 10446 47629 10502
rect 47553 10436 47629 10446
rect 48193 10606 48269 10616
rect 48193 10550 48203 10606
rect 48259 10550 48269 10606
rect 48193 10502 48269 10550
rect 48193 10446 48203 10502
rect 48259 10446 48269 10502
rect 48193 10436 48269 10446
rect 45018 10212 45094 10222
rect 45018 10156 45028 10212
rect 45084 10156 45094 10212
rect 45018 10108 45094 10156
rect 45018 10052 45028 10108
rect 45084 10052 45094 10108
rect 45018 10042 45094 10052
rect 45658 10212 45734 10222
rect 45658 10156 45668 10212
rect 45724 10156 45734 10212
rect 45658 10108 45734 10156
rect 45658 10052 45668 10108
rect 45724 10052 45734 10108
rect 45658 10042 45734 10052
rect 47234 10212 47310 10222
rect 47234 10156 47244 10212
rect 47300 10156 47310 10212
rect 47234 10108 47310 10156
rect 47234 10052 47244 10108
rect 47300 10052 47310 10108
rect 47234 10042 47310 10052
rect 47874 10212 47950 10222
rect 47874 10156 47884 10212
rect 47940 10156 47950 10212
rect 47874 10108 47950 10156
rect 47874 10052 47884 10108
rect 47940 10052 47950 10108
rect 47874 10042 47950 10052
rect 44298 9640 44310 9692
rect 44362 9640 44470 9692
rect 44522 9640 44534 9692
rect 41832 9490 41842 9546
rect 41898 9490 41946 9546
rect 42002 9490 42050 9546
rect 42106 9490 42116 9546
rect 41832 9442 42116 9490
rect 41832 9386 41842 9442
rect 41898 9386 41946 9442
rect 42002 9386 42050 9442
rect 42106 9386 42116 9442
rect 41112 8140 41122 8196
rect 41178 8140 41226 8196
rect 41282 8140 41330 8196
rect 41386 8140 41396 8196
rect 35322 8092 35398 8102
rect 35322 8036 35332 8092
rect 35388 8036 35398 8092
rect 35322 7988 35398 8036
rect 35322 7932 35332 7988
rect 35388 7932 35398 7988
rect 35322 7922 35398 7932
rect 35962 8092 36038 8102
rect 35962 8036 35972 8092
rect 36028 8036 36038 8092
rect 35962 7988 36038 8036
rect 35962 7932 35972 7988
rect 36028 7932 36038 7988
rect 35962 7922 36038 7932
rect 37538 8092 37614 8102
rect 37538 8036 37548 8092
rect 37604 8036 37614 8092
rect 37538 7988 37614 8036
rect 37538 7932 37548 7988
rect 37604 7932 37614 7988
rect 37538 7922 37614 7932
rect 38178 8092 38254 8102
rect 38178 8036 38188 8092
rect 38244 8036 38254 8092
rect 38178 7988 38254 8036
rect 38178 7932 38188 7988
rect 38244 7932 38254 7988
rect 38178 7922 38254 7932
rect 39458 8092 39534 8102
rect 39458 8036 39468 8092
rect 39524 8036 39534 8092
rect 39458 7988 39534 8036
rect 39458 7932 39468 7988
rect 39524 7932 39534 7988
rect 39458 7922 39534 7932
rect 40098 8092 40174 8102
rect 40098 8036 40108 8092
rect 40164 8036 40174 8092
rect 40098 7988 40174 8036
rect 40098 7932 40108 7988
rect 40164 7932 40174 7988
rect 40098 7922 40174 7932
rect 41112 8092 41396 8140
rect 41112 8036 41122 8092
rect 41178 8036 41226 8092
rect 41282 8036 41330 8092
rect 41386 8036 41396 8092
rect 41112 7988 41396 8036
rect 41112 7932 41122 7988
rect 41178 7932 41226 7988
rect 41282 7932 41330 7988
rect 41386 7932 41396 7988
rect 41112 7922 41396 7932
rect 41832 8196 42116 9386
rect 43419 9546 43495 9556
rect 43419 9490 43429 9546
rect 43485 9490 43495 9546
rect 43419 9442 43495 9490
rect 43419 9386 43429 9442
rect 43485 9386 43495 9442
rect 43419 9376 43495 9386
rect 44059 9546 44135 9556
rect 44059 9490 44069 9546
rect 44125 9490 44135 9546
rect 44059 9442 44135 9490
rect 44059 9386 44069 9442
rect 44125 9386 44135 9442
rect 44059 9376 44135 9386
rect 43098 9152 43174 9162
rect 43098 9096 43108 9152
rect 43164 9096 43174 9152
rect 43098 9048 43174 9096
rect 43098 8992 43108 9048
rect 43164 8992 43174 9048
rect 43098 8982 43174 8992
rect 43738 9152 43814 9162
rect 43738 9096 43748 9152
rect 43804 9096 43814 9152
rect 43738 9048 43814 9096
rect 43738 8992 43748 9048
rect 43804 8992 43814 9048
rect 43738 8982 43814 8992
rect 44298 8632 44534 9640
rect 48434 9692 48670 10700
rect 50788 10710 51072 11112
rect 50788 10654 50798 10710
rect 50854 10654 50902 10710
rect 50958 10654 51006 10710
rect 51062 10654 51072 10710
rect 48833 10606 48909 10616
rect 48833 10550 48843 10606
rect 48899 10550 48909 10606
rect 48833 10502 48909 10550
rect 48833 10446 48843 10502
rect 48899 10446 48909 10502
rect 48833 10436 48909 10446
rect 49473 10606 49549 10616
rect 49473 10550 49483 10606
rect 49539 10550 49549 10606
rect 49473 10502 49549 10550
rect 49473 10446 49483 10502
rect 49539 10446 49549 10502
rect 49473 10436 49549 10446
rect 50788 10606 51072 10654
rect 50788 10550 50798 10606
rect 50854 10550 50902 10606
rect 50958 10550 51006 10606
rect 51062 10550 51072 10606
rect 50788 10502 51072 10550
rect 50788 10446 50798 10502
rect 50854 10446 50902 10502
rect 50958 10446 51006 10502
rect 51062 10446 51072 10502
rect 49154 10212 49230 10222
rect 49154 10156 49164 10212
rect 49220 10156 49230 10212
rect 49154 10108 49230 10156
rect 49154 10052 49164 10108
rect 49220 10052 49230 10108
rect 49154 10042 49230 10052
rect 49794 10212 49870 10222
rect 49794 10156 49804 10212
rect 49860 10156 49870 10212
rect 49794 10108 49870 10156
rect 49794 10052 49804 10108
rect 49860 10052 49870 10108
rect 49794 10042 49870 10052
rect 48434 9640 48446 9692
rect 48498 9640 48606 9692
rect 48658 9640 48670 9692
rect 44699 9546 44775 9556
rect 44699 9490 44709 9546
rect 44765 9490 44775 9546
rect 44699 9442 44775 9490
rect 44699 9386 44709 9442
rect 44765 9386 44775 9442
rect 44699 9376 44775 9386
rect 45339 9546 45415 9556
rect 45339 9490 45349 9546
rect 45405 9490 45415 9546
rect 45339 9442 45415 9490
rect 45339 9386 45349 9442
rect 45405 9386 45415 9442
rect 45339 9376 45415 9386
rect 47553 9546 47629 9556
rect 47553 9490 47563 9546
rect 47619 9490 47629 9546
rect 47553 9442 47629 9490
rect 47553 9386 47563 9442
rect 47619 9386 47629 9442
rect 47553 9376 47629 9386
rect 48193 9546 48269 9556
rect 48193 9490 48203 9546
rect 48259 9490 48269 9546
rect 48193 9442 48269 9490
rect 48193 9386 48203 9442
rect 48259 9386 48269 9442
rect 48193 9376 48269 9386
rect 45018 9152 45094 9162
rect 45018 9096 45028 9152
rect 45084 9096 45094 9152
rect 45018 9048 45094 9096
rect 45018 8992 45028 9048
rect 45084 8992 45094 9048
rect 45018 8982 45094 8992
rect 45658 9152 45734 9162
rect 45658 9096 45668 9152
rect 45724 9096 45734 9152
rect 45658 9048 45734 9096
rect 45658 8992 45668 9048
rect 45724 8992 45734 9048
rect 45658 8982 45734 8992
rect 47234 9152 47310 9162
rect 47234 9096 47244 9152
rect 47300 9096 47310 9152
rect 47234 9048 47310 9096
rect 47234 8992 47244 9048
rect 47300 8992 47310 9048
rect 47234 8982 47310 8992
rect 47874 9152 47950 9162
rect 47874 9096 47884 9152
rect 47940 9096 47950 9152
rect 47874 9048 47950 9096
rect 47874 8992 47884 9048
rect 47940 8992 47950 9048
rect 47874 8982 47950 8992
rect 44298 8580 44310 8632
rect 44362 8580 44470 8632
rect 44522 8580 44534 8632
rect 44298 8568 44534 8580
rect 48434 8632 48670 9640
rect 50788 9650 51072 10446
rect 50788 9594 50798 9650
rect 50854 9594 50902 9650
rect 50958 9594 51006 9650
rect 51062 9594 51072 9650
rect 48833 9546 48909 9556
rect 48833 9490 48843 9546
rect 48899 9490 48909 9546
rect 48833 9442 48909 9490
rect 48833 9386 48843 9442
rect 48899 9386 48909 9442
rect 48833 9376 48909 9386
rect 49473 9546 49549 9556
rect 49473 9490 49483 9546
rect 49539 9490 49549 9546
rect 49473 9442 49549 9490
rect 49473 9386 49483 9442
rect 49539 9386 49549 9442
rect 49473 9376 49549 9386
rect 50788 9546 51072 9594
rect 50788 9490 50798 9546
rect 50854 9490 50902 9546
rect 50958 9490 51006 9546
rect 51062 9490 51072 9546
rect 50788 9442 51072 9490
rect 50788 9386 50798 9442
rect 50854 9386 50902 9442
rect 50958 9386 51006 9442
rect 51062 9386 51072 9442
rect 49154 9152 49230 9162
rect 49154 9096 49164 9152
rect 49220 9096 49230 9152
rect 49154 9048 49230 9096
rect 49154 8992 49164 9048
rect 49220 8992 49230 9048
rect 49154 8982 49230 8992
rect 49794 9152 49870 9162
rect 49794 9096 49804 9152
rect 49860 9096 49870 9152
rect 49794 9048 49870 9096
rect 49794 8992 49804 9048
rect 49860 8992 49870 9048
rect 49794 8982 49870 8992
rect 48434 8580 48446 8632
rect 48498 8580 48606 8632
rect 48658 8580 48670 8632
rect 48434 8568 48670 8580
rect 43419 8486 43495 8496
rect 43419 8430 43429 8486
rect 43485 8430 43495 8486
rect 43419 8382 43495 8430
rect 43419 8326 43429 8382
rect 43485 8326 43495 8382
rect 43419 8316 43495 8326
rect 44059 8486 44135 8496
rect 44059 8430 44069 8486
rect 44125 8430 44135 8486
rect 44059 8382 44135 8430
rect 44059 8326 44069 8382
rect 44125 8326 44135 8382
rect 44059 8316 44135 8326
rect 44699 8486 44775 8496
rect 44699 8430 44709 8486
rect 44765 8430 44775 8486
rect 44699 8382 44775 8430
rect 44699 8326 44709 8382
rect 44765 8326 44775 8382
rect 44699 8316 44775 8326
rect 45339 8486 45415 8496
rect 45339 8430 45349 8486
rect 45405 8430 45415 8486
rect 45339 8382 45415 8430
rect 45339 8326 45349 8382
rect 45405 8326 45415 8382
rect 45339 8316 45415 8326
rect 47553 8486 47629 8496
rect 47553 8430 47563 8486
rect 47619 8430 47629 8486
rect 47553 8382 47629 8430
rect 47553 8326 47563 8382
rect 47619 8326 47629 8382
rect 47553 8316 47629 8326
rect 48193 8486 48269 8496
rect 48193 8430 48203 8486
rect 48259 8430 48269 8486
rect 48193 8382 48269 8430
rect 48193 8326 48203 8382
rect 48259 8326 48269 8382
rect 48193 8316 48269 8326
rect 48833 8486 48909 8496
rect 48833 8430 48843 8486
rect 48899 8430 48909 8486
rect 48833 8382 48909 8430
rect 48833 8326 48843 8382
rect 48899 8326 48909 8382
rect 48833 8316 48909 8326
rect 49473 8486 49549 8496
rect 49473 8430 49483 8486
rect 49539 8430 49549 8486
rect 49473 8382 49549 8430
rect 49473 8326 49483 8382
rect 49539 8326 49549 8382
rect 49473 8316 49549 8326
rect 41832 8140 41842 8196
rect 41898 8140 41946 8196
rect 42002 8140 42050 8196
rect 42106 8140 42116 8196
rect 41832 8092 42116 8140
rect 50788 8196 51072 9386
rect 51128 10316 51412 11506
rect 53115 11666 53191 11676
rect 53115 11610 53125 11666
rect 53181 11610 53191 11666
rect 53115 11562 53191 11610
rect 53115 11506 53125 11562
rect 53181 11506 53191 11562
rect 53115 11496 53191 11506
rect 53755 11666 53831 11676
rect 53755 11610 53765 11666
rect 53821 11610 53831 11666
rect 53755 11562 53831 11610
rect 53755 11506 53765 11562
rect 53821 11506 53831 11562
rect 53755 11496 53831 11506
rect 51128 10260 51138 10316
rect 51194 10260 51242 10316
rect 51298 10260 51346 10316
rect 51402 10260 51412 10316
rect 51128 10212 51412 10260
rect 51128 10156 51138 10212
rect 51194 10156 51242 10212
rect 51298 10156 51346 10212
rect 51402 10156 51412 10212
rect 51128 10108 51412 10156
rect 51128 10052 51138 10108
rect 51194 10052 51242 10108
rect 51298 10052 51346 10108
rect 51402 10052 51412 10108
rect 51128 9256 51412 10052
rect 51128 9200 51138 9256
rect 51194 9200 51242 9256
rect 51298 9200 51346 9256
rect 51402 9200 51412 9256
rect 51128 9152 51412 9200
rect 51128 9096 51138 9152
rect 51194 9096 51242 9152
rect 51298 9096 51346 9152
rect 51402 9096 51412 9152
rect 51128 9048 51412 9096
rect 51128 8992 51138 9048
rect 51194 8992 51242 9048
rect 51298 8992 51346 9048
rect 51402 8992 51412 9048
rect 51128 8590 51412 8992
rect 51128 8534 51138 8590
rect 51194 8534 51242 8590
rect 51298 8534 51346 8590
rect 51402 8534 51412 8590
rect 51128 8486 51412 8534
rect 51128 8430 51138 8486
rect 51194 8430 51242 8486
rect 51298 8430 51346 8486
rect 51402 8430 51412 8486
rect 51128 8382 51412 8430
rect 51128 8326 51138 8382
rect 51194 8326 51242 8382
rect 51298 8326 51346 8382
rect 51402 8326 51412 8382
rect 51128 8316 51412 8326
rect 51520 11376 51804 11386
rect 51520 11320 51530 11376
rect 51586 11320 51634 11376
rect 51690 11320 51738 11376
rect 51794 11320 51804 11376
rect 51520 11272 51804 11320
rect 51520 11216 51530 11272
rect 51586 11216 51634 11272
rect 51690 11216 51738 11272
rect 51794 11216 51804 11272
rect 51520 11168 51804 11216
rect 51520 11112 51530 11168
rect 51586 11112 51634 11168
rect 51690 11112 51738 11168
rect 51794 11112 51804 11168
rect 51520 10710 51804 11112
rect 52794 11272 52870 11282
rect 52794 11216 52804 11272
rect 52860 11216 52870 11272
rect 52794 11168 52870 11216
rect 52794 11112 52804 11168
rect 52860 11112 52870 11168
rect 52794 11102 52870 11112
rect 53434 11272 53510 11282
rect 53434 11216 53444 11272
rect 53500 11216 53510 11272
rect 53434 11168 53510 11216
rect 53434 11112 53444 11168
rect 53500 11112 53510 11168
rect 53434 11102 53510 11112
rect 51520 10654 51530 10710
rect 51586 10654 51634 10710
rect 51690 10654 51738 10710
rect 51794 10654 51804 10710
rect 51520 10606 51804 10654
rect 53994 10752 54230 11760
rect 58130 11812 58366 12776
rect 58130 11760 58142 11812
rect 58194 11760 58302 11812
rect 58354 11760 58366 11812
rect 63690 11812 63926 12776
rect 54395 11666 54471 11676
rect 54395 11610 54405 11666
rect 54461 11610 54471 11666
rect 54395 11562 54471 11610
rect 54395 11506 54405 11562
rect 54461 11506 54471 11562
rect 54395 11496 54471 11506
rect 55035 11666 55111 11676
rect 55035 11610 55045 11666
rect 55101 11610 55111 11666
rect 55035 11562 55111 11610
rect 55035 11506 55045 11562
rect 55101 11506 55111 11562
rect 55035 11496 55111 11506
rect 57249 11666 57325 11676
rect 57249 11610 57259 11666
rect 57315 11610 57325 11666
rect 57249 11562 57325 11610
rect 57249 11506 57259 11562
rect 57315 11506 57325 11562
rect 57249 11496 57325 11506
rect 57889 11666 57965 11676
rect 57889 11610 57899 11666
rect 57955 11610 57965 11666
rect 57889 11562 57965 11610
rect 57889 11506 57899 11562
rect 57955 11506 57965 11562
rect 57889 11496 57965 11506
rect 54714 11272 54790 11282
rect 54714 11216 54724 11272
rect 54780 11216 54790 11272
rect 54714 11168 54790 11216
rect 54714 11112 54724 11168
rect 54780 11112 54790 11168
rect 54714 11102 54790 11112
rect 55354 11272 55430 11282
rect 55354 11216 55364 11272
rect 55420 11216 55430 11272
rect 55354 11168 55430 11216
rect 55354 11112 55364 11168
rect 55420 11112 55430 11168
rect 55354 11102 55430 11112
rect 56930 11272 57006 11282
rect 56930 11216 56940 11272
rect 56996 11216 57006 11272
rect 56930 11168 57006 11216
rect 56930 11112 56940 11168
rect 56996 11112 57006 11168
rect 56930 11102 57006 11112
rect 57570 11272 57646 11282
rect 57570 11216 57580 11272
rect 57636 11216 57646 11272
rect 57570 11168 57646 11216
rect 57570 11112 57580 11168
rect 57636 11112 57646 11168
rect 57570 11102 57646 11112
rect 53994 10700 54006 10752
rect 54058 10700 54166 10752
rect 54218 10700 54230 10752
rect 51520 10550 51530 10606
rect 51586 10550 51634 10606
rect 51690 10550 51738 10606
rect 51794 10550 51804 10606
rect 51520 10502 51804 10550
rect 51520 10446 51530 10502
rect 51586 10446 51634 10502
rect 51690 10446 51738 10502
rect 51794 10446 51804 10502
rect 51520 9650 51804 10446
rect 53115 10606 53191 10616
rect 53115 10550 53125 10606
rect 53181 10550 53191 10606
rect 53115 10502 53191 10550
rect 53115 10446 53125 10502
rect 53181 10446 53191 10502
rect 53115 10436 53191 10446
rect 53755 10606 53831 10616
rect 53755 10550 53765 10606
rect 53821 10550 53831 10606
rect 53755 10502 53831 10550
rect 53755 10446 53765 10502
rect 53821 10446 53831 10502
rect 53755 10436 53831 10446
rect 52794 10212 52870 10222
rect 52794 10156 52804 10212
rect 52860 10156 52870 10212
rect 52794 10108 52870 10156
rect 52794 10052 52804 10108
rect 52860 10052 52870 10108
rect 52794 10042 52870 10052
rect 53434 10212 53510 10222
rect 53434 10156 53444 10212
rect 53500 10156 53510 10212
rect 53434 10108 53510 10156
rect 53434 10052 53444 10108
rect 53500 10052 53510 10108
rect 53434 10042 53510 10052
rect 51520 9594 51530 9650
rect 51586 9594 51634 9650
rect 51690 9594 51738 9650
rect 51794 9594 51804 9650
rect 51520 9546 51804 9594
rect 53994 9692 54230 10700
rect 58130 10752 58366 11760
rect 60909 11770 61193 11780
rect 60909 11714 60919 11770
rect 60975 11714 61023 11770
rect 61079 11714 61127 11770
rect 61183 11714 61193 11770
rect 58529 11666 58605 11676
rect 58529 11610 58539 11666
rect 58595 11610 58605 11666
rect 58529 11562 58605 11610
rect 58529 11506 58539 11562
rect 58595 11506 58605 11562
rect 58529 11496 58605 11506
rect 59169 11666 59245 11676
rect 59169 11610 59179 11666
rect 59235 11610 59245 11666
rect 59169 11562 59245 11610
rect 59169 11506 59179 11562
rect 59235 11506 59245 11562
rect 59169 11496 59245 11506
rect 60909 11666 61193 11714
rect 63690 11760 63702 11812
rect 63754 11760 63862 11812
rect 63914 11760 63926 11812
rect 60909 11610 60919 11666
rect 60975 11610 61023 11666
rect 61079 11610 61127 11666
rect 61183 11610 61193 11666
rect 60909 11562 61193 11610
rect 60909 11506 60919 11562
rect 60975 11506 61023 11562
rect 61079 11506 61127 11562
rect 61183 11506 61193 11562
rect 60504 11376 60788 11386
rect 60504 11320 60514 11376
rect 60570 11320 60618 11376
rect 60674 11320 60722 11376
rect 60778 11320 60788 11376
rect 58850 11272 58926 11282
rect 58850 11216 58860 11272
rect 58916 11216 58926 11272
rect 58850 11168 58926 11216
rect 58850 11112 58860 11168
rect 58916 11112 58926 11168
rect 58850 11102 58926 11112
rect 59490 11272 59566 11282
rect 59490 11216 59500 11272
rect 59556 11216 59566 11272
rect 59490 11168 59566 11216
rect 59490 11112 59500 11168
rect 59556 11112 59566 11168
rect 59490 11102 59566 11112
rect 60504 11272 60788 11320
rect 60504 11216 60514 11272
rect 60570 11216 60618 11272
rect 60674 11216 60722 11272
rect 60778 11216 60788 11272
rect 60504 11168 60788 11216
rect 60504 11112 60514 11168
rect 60570 11112 60618 11168
rect 60674 11112 60722 11168
rect 60778 11112 60788 11168
rect 58130 10700 58142 10752
rect 58194 10700 58302 10752
rect 58354 10700 58366 10752
rect 54395 10606 54471 10616
rect 54395 10550 54405 10606
rect 54461 10550 54471 10606
rect 54395 10502 54471 10550
rect 54395 10446 54405 10502
rect 54461 10446 54471 10502
rect 54395 10436 54471 10446
rect 55035 10606 55111 10616
rect 55035 10550 55045 10606
rect 55101 10550 55111 10606
rect 55035 10502 55111 10550
rect 55035 10446 55045 10502
rect 55101 10446 55111 10502
rect 55035 10436 55111 10446
rect 57249 10606 57325 10616
rect 57249 10550 57259 10606
rect 57315 10550 57325 10606
rect 57249 10502 57325 10550
rect 57249 10446 57259 10502
rect 57315 10446 57325 10502
rect 57249 10436 57325 10446
rect 57889 10606 57965 10616
rect 57889 10550 57899 10606
rect 57955 10550 57965 10606
rect 57889 10502 57965 10550
rect 57889 10446 57899 10502
rect 57955 10446 57965 10502
rect 57889 10436 57965 10446
rect 54714 10212 54790 10222
rect 54714 10156 54724 10212
rect 54780 10156 54790 10212
rect 54714 10108 54790 10156
rect 54714 10052 54724 10108
rect 54780 10052 54790 10108
rect 54714 10042 54790 10052
rect 55354 10212 55430 10222
rect 55354 10156 55364 10212
rect 55420 10156 55430 10212
rect 55354 10108 55430 10156
rect 55354 10052 55364 10108
rect 55420 10052 55430 10108
rect 55354 10042 55430 10052
rect 56930 10212 57006 10222
rect 56930 10156 56940 10212
rect 56996 10156 57006 10212
rect 56930 10108 57006 10156
rect 56930 10052 56940 10108
rect 56996 10052 57006 10108
rect 56930 10042 57006 10052
rect 57570 10212 57646 10222
rect 57570 10156 57580 10212
rect 57636 10156 57646 10212
rect 57570 10108 57646 10156
rect 57570 10052 57580 10108
rect 57636 10052 57646 10108
rect 57570 10042 57646 10052
rect 53994 9640 54006 9692
rect 54058 9640 54166 9692
rect 54218 9640 54230 9692
rect 51520 9490 51530 9546
rect 51586 9490 51634 9546
rect 51690 9490 51738 9546
rect 51794 9490 51804 9546
rect 51520 9442 51804 9490
rect 51520 9386 51530 9442
rect 51586 9386 51634 9442
rect 51690 9386 51738 9442
rect 51794 9386 51804 9442
rect 50788 8140 50798 8196
rect 50854 8140 50902 8196
rect 50958 8140 51006 8196
rect 51062 8140 51072 8196
rect 41832 8036 41842 8092
rect 41898 8036 41946 8092
rect 42002 8036 42050 8092
rect 42106 8036 42116 8092
rect 41832 7988 42116 8036
rect 41832 7932 41842 7988
rect 41898 7932 41946 7988
rect 42002 7932 42050 7988
rect 42106 7932 42116 7988
rect 41832 7922 42116 7932
rect 43098 8092 43174 8102
rect 43098 8036 43108 8092
rect 43164 8036 43174 8092
rect 43098 7988 43174 8036
rect 43098 7932 43108 7988
rect 43164 7932 43174 7988
rect 43098 7922 43174 7932
rect 43738 8092 43814 8102
rect 43738 8036 43748 8092
rect 43804 8036 43814 8092
rect 43738 7988 43814 8036
rect 43738 7932 43748 7988
rect 43804 7932 43814 7988
rect 43738 7922 43814 7932
rect 45018 8092 45094 8102
rect 45018 8036 45028 8092
rect 45084 8036 45094 8092
rect 45018 7988 45094 8036
rect 45018 7932 45028 7988
rect 45084 7932 45094 7988
rect 45018 7922 45094 7932
rect 45658 8092 45734 8102
rect 45658 8036 45668 8092
rect 45724 8036 45734 8092
rect 45658 7988 45734 8036
rect 45658 7932 45668 7988
rect 45724 7932 45734 7988
rect 45658 7922 45734 7932
rect 47234 8092 47310 8102
rect 47234 8036 47244 8092
rect 47300 8036 47310 8092
rect 47234 7988 47310 8036
rect 47234 7932 47244 7988
rect 47300 7932 47310 7988
rect 47234 7922 47310 7932
rect 47874 8092 47950 8102
rect 47874 8036 47884 8092
rect 47940 8036 47950 8092
rect 47874 7988 47950 8036
rect 47874 7932 47884 7988
rect 47940 7932 47950 7988
rect 47874 7922 47950 7932
rect 49154 8092 49230 8102
rect 49154 8036 49164 8092
rect 49220 8036 49230 8092
rect 49154 7988 49230 8036
rect 49154 7932 49164 7988
rect 49220 7932 49230 7988
rect 49154 7922 49230 7932
rect 49794 8092 49870 8102
rect 49794 8036 49804 8092
rect 49860 8036 49870 8092
rect 49794 7988 49870 8036
rect 49794 7932 49804 7988
rect 49860 7932 49870 7988
rect 49794 7922 49870 7932
rect 50788 8092 51072 8140
rect 50788 8036 50798 8092
rect 50854 8036 50902 8092
rect 50958 8036 51006 8092
rect 51062 8036 51072 8092
rect 50788 7988 51072 8036
rect 50788 7932 50798 7988
rect 50854 7932 50902 7988
rect 50958 7932 51006 7988
rect 51062 7932 51072 7988
rect 50788 7922 51072 7932
rect 51520 8196 51804 9386
rect 53115 9546 53191 9556
rect 53115 9490 53125 9546
rect 53181 9490 53191 9546
rect 53115 9442 53191 9490
rect 53115 9386 53125 9442
rect 53181 9386 53191 9442
rect 53115 9376 53191 9386
rect 53755 9546 53831 9556
rect 53755 9490 53765 9546
rect 53821 9490 53831 9546
rect 53755 9442 53831 9490
rect 53755 9386 53765 9442
rect 53821 9386 53831 9442
rect 53755 9376 53831 9386
rect 52794 9152 52870 9162
rect 52794 9096 52804 9152
rect 52860 9096 52870 9152
rect 52794 9048 52870 9096
rect 52794 8992 52804 9048
rect 52860 8992 52870 9048
rect 52794 8982 52870 8992
rect 53434 9152 53510 9162
rect 53434 9096 53444 9152
rect 53500 9096 53510 9152
rect 53434 9048 53510 9096
rect 53434 8992 53444 9048
rect 53500 8992 53510 9048
rect 53434 8982 53510 8992
rect 53994 8632 54230 9640
rect 58130 9692 58366 10700
rect 60504 10710 60788 11112
rect 60504 10654 60514 10710
rect 60570 10654 60618 10710
rect 60674 10654 60722 10710
rect 60778 10654 60788 10710
rect 58529 10606 58605 10616
rect 58529 10550 58539 10606
rect 58595 10550 58605 10606
rect 58529 10502 58605 10550
rect 58529 10446 58539 10502
rect 58595 10446 58605 10502
rect 58529 10436 58605 10446
rect 59169 10606 59245 10616
rect 59169 10550 59179 10606
rect 59235 10550 59245 10606
rect 59169 10502 59245 10550
rect 59169 10446 59179 10502
rect 59235 10446 59245 10502
rect 59169 10436 59245 10446
rect 60504 10606 60788 10654
rect 60504 10550 60514 10606
rect 60570 10550 60618 10606
rect 60674 10550 60722 10606
rect 60778 10550 60788 10606
rect 60504 10502 60788 10550
rect 60504 10446 60514 10502
rect 60570 10446 60618 10502
rect 60674 10446 60722 10502
rect 60778 10446 60788 10502
rect 58850 10212 58926 10222
rect 58850 10156 58860 10212
rect 58916 10156 58926 10212
rect 58850 10108 58926 10156
rect 58850 10052 58860 10108
rect 58916 10052 58926 10108
rect 58850 10042 58926 10052
rect 59490 10212 59566 10222
rect 59490 10156 59500 10212
rect 59556 10156 59566 10212
rect 59490 10108 59566 10156
rect 59490 10052 59500 10108
rect 59556 10052 59566 10108
rect 59490 10042 59566 10052
rect 58130 9640 58142 9692
rect 58194 9640 58302 9692
rect 58354 9640 58366 9692
rect 54395 9546 54471 9556
rect 54395 9490 54405 9546
rect 54461 9490 54471 9546
rect 54395 9442 54471 9490
rect 54395 9386 54405 9442
rect 54461 9386 54471 9442
rect 54395 9376 54471 9386
rect 55035 9546 55111 9556
rect 55035 9490 55045 9546
rect 55101 9490 55111 9546
rect 55035 9442 55111 9490
rect 55035 9386 55045 9442
rect 55101 9386 55111 9442
rect 55035 9376 55111 9386
rect 57249 9546 57325 9556
rect 57249 9490 57259 9546
rect 57315 9490 57325 9546
rect 57249 9442 57325 9490
rect 57249 9386 57259 9442
rect 57315 9386 57325 9442
rect 57249 9376 57325 9386
rect 57889 9546 57965 9556
rect 57889 9490 57899 9546
rect 57955 9490 57965 9546
rect 57889 9442 57965 9490
rect 57889 9386 57899 9442
rect 57955 9386 57965 9442
rect 57889 9376 57965 9386
rect 54714 9152 54790 9162
rect 54714 9096 54724 9152
rect 54780 9096 54790 9152
rect 54714 9048 54790 9096
rect 54714 8992 54724 9048
rect 54780 8992 54790 9048
rect 54714 8982 54790 8992
rect 55354 9152 55430 9162
rect 55354 9096 55364 9152
rect 55420 9096 55430 9152
rect 55354 9048 55430 9096
rect 55354 8992 55364 9048
rect 55420 8992 55430 9048
rect 55354 8982 55430 8992
rect 56930 9152 57006 9162
rect 56930 9096 56940 9152
rect 56996 9096 57006 9152
rect 56930 9048 57006 9096
rect 56930 8992 56940 9048
rect 56996 8992 57006 9048
rect 56930 8982 57006 8992
rect 57570 9152 57646 9162
rect 57570 9096 57580 9152
rect 57636 9096 57646 9152
rect 57570 9048 57646 9096
rect 57570 8992 57580 9048
rect 57636 8992 57646 9048
rect 57570 8982 57646 8992
rect 53994 8580 54006 8632
rect 54058 8580 54166 8632
rect 54218 8580 54230 8632
rect 53994 8568 54230 8580
rect 58130 8632 58366 9640
rect 60504 9650 60788 10446
rect 60504 9594 60514 9650
rect 60570 9594 60618 9650
rect 60674 9594 60722 9650
rect 60778 9594 60788 9650
rect 58529 9546 58605 9556
rect 58529 9490 58539 9546
rect 58595 9490 58605 9546
rect 58529 9442 58605 9490
rect 58529 9386 58539 9442
rect 58595 9386 58605 9442
rect 58529 9376 58605 9386
rect 59169 9546 59245 9556
rect 59169 9490 59179 9546
rect 59235 9490 59245 9546
rect 59169 9442 59245 9490
rect 59169 9386 59179 9442
rect 59235 9386 59245 9442
rect 59169 9376 59245 9386
rect 60504 9546 60788 9594
rect 60504 9490 60514 9546
rect 60570 9490 60618 9546
rect 60674 9490 60722 9546
rect 60778 9490 60788 9546
rect 60504 9442 60788 9490
rect 60504 9386 60514 9442
rect 60570 9386 60618 9442
rect 60674 9386 60722 9442
rect 60778 9386 60788 9442
rect 58850 9152 58926 9162
rect 58850 9096 58860 9152
rect 58916 9096 58926 9152
rect 58850 9048 58926 9096
rect 58850 8992 58860 9048
rect 58916 8992 58926 9048
rect 58850 8982 58926 8992
rect 59490 9152 59566 9162
rect 59490 9096 59500 9152
rect 59556 9096 59566 9152
rect 59490 9048 59566 9096
rect 59490 8992 59500 9048
rect 59556 8992 59566 9048
rect 59490 8982 59566 8992
rect 58130 8580 58142 8632
rect 58194 8580 58302 8632
rect 58354 8580 58366 8632
rect 58130 8568 58366 8580
rect 53115 8486 53191 8496
rect 53115 8430 53125 8486
rect 53181 8430 53191 8486
rect 53115 8382 53191 8430
rect 53115 8326 53125 8382
rect 53181 8326 53191 8382
rect 53115 8316 53191 8326
rect 53755 8486 53831 8496
rect 53755 8430 53765 8486
rect 53821 8430 53831 8486
rect 53755 8382 53831 8430
rect 53755 8326 53765 8382
rect 53821 8326 53831 8382
rect 53755 8316 53831 8326
rect 54395 8486 54471 8496
rect 54395 8430 54405 8486
rect 54461 8430 54471 8486
rect 54395 8382 54471 8430
rect 54395 8326 54405 8382
rect 54461 8326 54471 8382
rect 54395 8316 54471 8326
rect 55035 8486 55111 8496
rect 55035 8430 55045 8486
rect 55101 8430 55111 8486
rect 55035 8382 55111 8430
rect 55035 8326 55045 8382
rect 55101 8326 55111 8382
rect 55035 8316 55111 8326
rect 57249 8486 57325 8496
rect 57249 8430 57259 8486
rect 57315 8430 57325 8486
rect 57249 8382 57325 8430
rect 57249 8326 57259 8382
rect 57315 8326 57325 8382
rect 57249 8316 57325 8326
rect 57889 8486 57965 8496
rect 57889 8430 57899 8486
rect 57955 8430 57965 8486
rect 57889 8382 57965 8430
rect 57889 8326 57899 8382
rect 57955 8326 57965 8382
rect 57889 8316 57965 8326
rect 58529 8486 58605 8496
rect 58529 8430 58539 8486
rect 58595 8430 58605 8486
rect 58529 8382 58605 8430
rect 58529 8326 58539 8382
rect 58595 8326 58605 8382
rect 58529 8316 58605 8326
rect 59169 8486 59245 8496
rect 59169 8430 59179 8486
rect 59235 8430 59245 8486
rect 59169 8382 59245 8430
rect 59169 8326 59179 8382
rect 59235 8326 59245 8382
rect 59169 8316 59245 8326
rect 51520 8140 51530 8196
rect 51586 8140 51634 8196
rect 51690 8140 51738 8196
rect 51794 8140 51804 8196
rect 51520 8092 51804 8140
rect 60504 8196 60788 9386
rect 60909 10316 61193 11506
rect 62811 11666 62887 11676
rect 62811 11610 62821 11666
rect 62877 11610 62887 11666
rect 62811 11562 62887 11610
rect 62811 11506 62821 11562
rect 62877 11506 62887 11562
rect 62811 11496 62887 11506
rect 63451 11666 63527 11676
rect 63451 11610 63461 11666
rect 63517 11610 63527 11666
rect 63451 11562 63527 11610
rect 63451 11506 63461 11562
rect 63517 11506 63527 11562
rect 63451 11496 63527 11506
rect 60909 10260 60919 10316
rect 60975 10260 61023 10316
rect 61079 10260 61127 10316
rect 61183 10260 61193 10316
rect 60909 10212 61193 10260
rect 60909 10156 60919 10212
rect 60975 10156 61023 10212
rect 61079 10156 61127 10212
rect 61183 10156 61193 10212
rect 60909 10108 61193 10156
rect 60909 10052 60919 10108
rect 60975 10052 61023 10108
rect 61079 10052 61127 10108
rect 61183 10052 61193 10108
rect 60909 9256 61193 10052
rect 60909 9200 60919 9256
rect 60975 9200 61023 9256
rect 61079 9200 61127 9256
rect 61183 9200 61193 9256
rect 60909 9152 61193 9200
rect 60909 9096 60919 9152
rect 60975 9096 61023 9152
rect 61079 9096 61127 9152
rect 61183 9096 61193 9152
rect 60909 9048 61193 9096
rect 60909 8992 60919 9048
rect 60975 8992 61023 9048
rect 61079 8992 61127 9048
rect 61183 8992 61193 9048
rect 60909 8590 61193 8992
rect 60909 8534 60919 8590
rect 60975 8534 61023 8590
rect 61079 8534 61127 8590
rect 61183 8534 61193 8590
rect 60909 8486 61193 8534
rect 60909 8430 60919 8486
rect 60975 8430 61023 8486
rect 61079 8430 61127 8486
rect 61183 8430 61193 8486
rect 60909 8382 61193 8430
rect 60909 8326 60919 8382
rect 60975 8326 61023 8382
rect 61079 8326 61127 8382
rect 61183 8326 61193 8382
rect 60909 8316 61193 8326
rect 61268 11376 61552 11386
rect 61268 11320 61278 11376
rect 61334 11320 61382 11376
rect 61438 11320 61486 11376
rect 61542 11320 61552 11376
rect 61268 11272 61552 11320
rect 61268 11216 61278 11272
rect 61334 11216 61382 11272
rect 61438 11216 61486 11272
rect 61542 11216 61552 11272
rect 61268 11168 61552 11216
rect 61268 11112 61278 11168
rect 61334 11112 61382 11168
rect 61438 11112 61486 11168
rect 61542 11112 61552 11168
rect 61268 10710 61552 11112
rect 62490 11272 62566 11282
rect 62490 11216 62500 11272
rect 62556 11216 62566 11272
rect 62490 11168 62566 11216
rect 62490 11112 62500 11168
rect 62556 11112 62566 11168
rect 62490 11102 62566 11112
rect 63130 11272 63206 11282
rect 63130 11216 63140 11272
rect 63196 11216 63206 11272
rect 63130 11168 63206 11216
rect 63130 11112 63140 11168
rect 63196 11112 63206 11168
rect 63130 11102 63206 11112
rect 61268 10654 61278 10710
rect 61334 10654 61382 10710
rect 61438 10654 61486 10710
rect 61542 10654 61552 10710
rect 61268 10606 61552 10654
rect 63690 10752 63926 11760
rect 64091 11666 64167 11676
rect 64091 11610 64101 11666
rect 64157 11610 64167 11666
rect 64091 11562 64167 11610
rect 64091 11506 64101 11562
rect 64157 11506 64167 11562
rect 64091 11496 64167 11506
rect 64731 11666 64807 11676
rect 64731 11610 64741 11666
rect 64797 11610 64807 11666
rect 64731 11562 64807 11610
rect 64731 11506 64741 11562
rect 64797 11506 64807 11562
rect 64731 11496 64807 11506
rect 64410 11272 64486 11282
rect 64410 11216 64420 11272
rect 64476 11216 64486 11272
rect 64410 11168 64486 11216
rect 64410 11112 64420 11168
rect 64476 11112 64486 11168
rect 64410 11102 64486 11112
rect 65050 11272 65126 11282
rect 65050 11216 65060 11272
rect 65116 11216 65126 11272
rect 65050 11168 65126 11216
rect 65050 11112 65060 11168
rect 65116 11112 65126 11168
rect 65050 11102 65126 11112
rect 63690 10700 63702 10752
rect 63754 10700 63862 10752
rect 63914 10700 63926 10752
rect 61268 10550 61278 10606
rect 61334 10550 61382 10606
rect 61438 10550 61486 10606
rect 61542 10550 61552 10606
rect 61268 10502 61552 10550
rect 61268 10446 61278 10502
rect 61334 10446 61382 10502
rect 61438 10446 61486 10502
rect 61542 10446 61552 10502
rect 61268 9650 61552 10446
rect 62811 10606 62887 10616
rect 62811 10550 62821 10606
rect 62877 10550 62887 10606
rect 62811 10502 62887 10550
rect 62811 10446 62821 10502
rect 62877 10446 62887 10502
rect 62811 10436 62887 10446
rect 63451 10606 63527 10616
rect 63451 10550 63461 10606
rect 63517 10550 63527 10606
rect 63451 10502 63527 10550
rect 63451 10446 63461 10502
rect 63517 10446 63527 10502
rect 63451 10436 63527 10446
rect 62490 10212 62566 10222
rect 62490 10156 62500 10212
rect 62556 10156 62566 10212
rect 62490 10108 62566 10156
rect 62490 10052 62500 10108
rect 62556 10052 62566 10108
rect 62490 10042 62566 10052
rect 63130 10212 63206 10222
rect 63130 10156 63140 10212
rect 63196 10156 63206 10212
rect 63130 10108 63206 10156
rect 63130 10052 63140 10108
rect 63196 10052 63206 10108
rect 63130 10042 63206 10052
rect 61268 9594 61278 9650
rect 61334 9594 61382 9650
rect 61438 9594 61486 9650
rect 61542 9594 61552 9650
rect 61268 9546 61552 9594
rect 63690 9692 63926 10700
rect 64091 10606 64167 10616
rect 64091 10550 64101 10606
rect 64157 10550 64167 10606
rect 64091 10502 64167 10550
rect 64091 10446 64101 10502
rect 64157 10446 64167 10502
rect 64091 10436 64167 10446
rect 64731 10606 64807 10616
rect 64731 10550 64741 10606
rect 64797 10550 64807 10606
rect 64731 10502 64807 10550
rect 64731 10446 64741 10502
rect 64797 10446 64807 10502
rect 64731 10436 64807 10446
rect 64410 10212 64486 10222
rect 64410 10156 64420 10212
rect 64476 10156 64486 10212
rect 64410 10108 64486 10156
rect 64410 10052 64420 10108
rect 64476 10052 64486 10108
rect 64410 10042 64486 10052
rect 65050 10212 65126 10222
rect 65050 10156 65060 10212
rect 65116 10156 65126 10212
rect 65050 10108 65126 10156
rect 65050 10052 65060 10108
rect 65116 10052 65126 10108
rect 65050 10042 65126 10052
rect 63690 9640 63702 9692
rect 63754 9640 63862 9692
rect 63914 9640 63926 9692
rect 61268 9490 61278 9546
rect 61334 9490 61382 9546
rect 61438 9490 61486 9546
rect 61542 9490 61552 9546
rect 61268 9442 61552 9490
rect 61268 9386 61278 9442
rect 61334 9386 61382 9442
rect 61438 9386 61486 9442
rect 61542 9386 61552 9442
rect 60504 8140 60514 8196
rect 60570 8140 60618 8196
rect 60674 8140 60722 8196
rect 60778 8140 60788 8196
rect 51520 8036 51530 8092
rect 51586 8036 51634 8092
rect 51690 8036 51738 8092
rect 51794 8036 51804 8092
rect 51520 7988 51804 8036
rect 51520 7932 51530 7988
rect 51586 7932 51634 7988
rect 51690 7932 51738 7988
rect 51794 7932 51804 7988
rect 51520 7922 51804 7932
rect 52794 8092 52870 8102
rect 52794 8036 52804 8092
rect 52860 8036 52870 8092
rect 52794 7988 52870 8036
rect 52794 7932 52804 7988
rect 52860 7932 52870 7988
rect 52794 7922 52870 7932
rect 53434 8092 53510 8102
rect 53434 8036 53444 8092
rect 53500 8036 53510 8092
rect 53434 7988 53510 8036
rect 53434 7932 53444 7988
rect 53500 7932 53510 7988
rect 53434 7922 53510 7932
rect 54714 8092 54790 8102
rect 54714 8036 54724 8092
rect 54780 8036 54790 8092
rect 54714 7988 54790 8036
rect 54714 7932 54724 7988
rect 54780 7932 54790 7988
rect 54714 7922 54790 7932
rect 55354 8092 55430 8102
rect 55354 8036 55364 8092
rect 55420 8036 55430 8092
rect 55354 7988 55430 8036
rect 55354 7932 55364 7988
rect 55420 7932 55430 7988
rect 55354 7922 55430 7932
rect 56930 8092 57006 8102
rect 56930 8036 56940 8092
rect 56996 8036 57006 8092
rect 56930 7988 57006 8036
rect 56930 7932 56940 7988
rect 56996 7932 57006 7988
rect 56930 7922 57006 7932
rect 57570 8092 57646 8102
rect 57570 8036 57580 8092
rect 57636 8036 57646 8092
rect 57570 7988 57646 8036
rect 57570 7932 57580 7988
rect 57636 7932 57646 7988
rect 57570 7922 57646 7932
rect 58850 8092 58926 8102
rect 58850 8036 58860 8092
rect 58916 8036 58926 8092
rect 58850 7988 58926 8036
rect 58850 7932 58860 7988
rect 58916 7932 58926 7988
rect 58850 7922 58926 7932
rect 59490 8092 59566 8102
rect 59490 8036 59500 8092
rect 59556 8036 59566 8092
rect 59490 7988 59566 8036
rect 59490 7932 59500 7988
rect 59556 7932 59566 7988
rect 59490 7922 59566 7932
rect 60504 8092 60788 8140
rect 60504 8036 60514 8092
rect 60570 8036 60618 8092
rect 60674 8036 60722 8092
rect 60778 8036 60788 8092
rect 60504 7988 60788 8036
rect 60504 7932 60514 7988
rect 60570 7932 60618 7988
rect 60674 7932 60722 7988
rect 60778 7932 60788 7988
rect 60504 7922 60788 7932
rect 61268 8196 61552 9386
rect 62811 9546 62887 9556
rect 62811 9490 62821 9546
rect 62877 9490 62887 9546
rect 62811 9442 62887 9490
rect 62811 9386 62821 9442
rect 62877 9386 62887 9442
rect 62811 9376 62887 9386
rect 63451 9546 63527 9556
rect 63451 9490 63461 9546
rect 63517 9490 63527 9546
rect 63451 9442 63527 9490
rect 63451 9386 63461 9442
rect 63517 9386 63527 9442
rect 63451 9376 63527 9386
rect 62490 9152 62566 9162
rect 62490 9096 62500 9152
rect 62556 9096 62566 9152
rect 62490 9048 62566 9096
rect 62490 8992 62500 9048
rect 62556 8992 62566 9048
rect 62490 8982 62566 8992
rect 63130 9152 63206 9162
rect 63130 9096 63140 9152
rect 63196 9096 63206 9152
rect 63130 9048 63206 9096
rect 63130 8992 63140 9048
rect 63196 8992 63206 9048
rect 63130 8982 63206 8992
rect 63690 8632 63926 9640
rect 64091 9546 64167 9556
rect 64091 9490 64101 9546
rect 64157 9490 64167 9546
rect 64091 9442 64167 9490
rect 64091 9386 64101 9442
rect 64157 9386 64167 9442
rect 64091 9376 64167 9386
rect 64731 9546 64807 9556
rect 64731 9490 64741 9546
rect 64797 9490 64807 9546
rect 64731 9442 64807 9490
rect 64731 9386 64741 9442
rect 64797 9386 64807 9442
rect 64731 9376 64807 9386
rect 64410 9152 64486 9162
rect 64410 9096 64420 9152
rect 64476 9096 64486 9152
rect 64410 9048 64486 9096
rect 64410 8992 64420 9048
rect 64476 8992 64486 9048
rect 64410 8982 64486 8992
rect 65050 9152 65126 9162
rect 65050 9096 65060 9152
rect 65116 9096 65126 9152
rect 65050 9048 65126 9096
rect 65050 8992 65060 9048
rect 65116 8992 65126 9048
rect 65050 8982 65126 8992
rect 63690 8580 63702 8632
rect 63754 8580 63862 8632
rect 63914 8580 63926 8632
rect 63690 8568 63926 8580
rect 62811 8486 62887 8496
rect 62811 8430 62821 8486
rect 62877 8430 62887 8486
rect 62811 8382 62887 8430
rect 62811 8326 62821 8382
rect 62877 8326 62887 8382
rect 62811 8316 62887 8326
rect 63451 8486 63527 8496
rect 63451 8430 63461 8486
rect 63517 8430 63527 8486
rect 63451 8382 63527 8430
rect 63451 8326 63461 8382
rect 63517 8326 63527 8382
rect 63451 8316 63527 8326
rect 64091 8486 64167 8496
rect 64091 8430 64101 8486
rect 64157 8430 64167 8486
rect 64091 8382 64167 8430
rect 64091 8326 64101 8382
rect 64157 8326 64167 8382
rect 64091 8316 64167 8326
rect 64731 8486 64807 8496
rect 64731 8430 64741 8486
rect 64797 8430 64807 8486
rect 64731 8382 64807 8430
rect 64731 8326 64741 8382
rect 64797 8326 64807 8382
rect 64731 8316 64807 8326
rect 61268 8140 61278 8196
rect 61334 8140 61382 8196
rect 61438 8140 61486 8196
rect 61542 8140 61552 8196
rect 61268 8092 61552 8140
rect 61268 8036 61278 8092
rect 61334 8036 61382 8092
rect 61438 8036 61486 8092
rect 61542 8036 61552 8092
rect 61268 7988 61552 8036
rect 61268 7932 61278 7988
rect 61334 7932 61382 7988
rect 61438 7932 61486 7988
rect 61542 7932 61552 7988
rect 61268 7922 61552 7932
rect 62490 8092 62566 8102
rect 62490 8036 62500 8092
rect 62556 8036 62566 8092
rect 62490 7988 62566 8036
rect 62490 7932 62500 7988
rect 62556 7932 62566 7988
rect 62490 7922 62566 7932
rect 63130 8092 63206 8102
rect 63130 8036 63140 8092
rect 63196 8036 63206 8092
rect 63130 7988 63206 8036
rect 63130 7932 63140 7988
rect 63196 7932 63206 7988
rect 63130 7922 63206 7932
rect 64410 8092 64486 8102
rect 64410 8036 64420 8092
rect 64476 8036 64486 8092
rect 64410 7988 64486 8036
rect 64410 7932 64420 7988
rect 64476 7932 64486 7988
rect 64410 7922 64486 7932
rect 65050 8092 65126 8102
rect 65050 8036 65060 8092
rect 65116 8036 65126 8092
rect 65050 7988 65126 8036
rect 65050 7932 65060 7988
rect 65116 7932 65126 7988
rect 65050 7922 65126 7932
rect 34602 3508 34640 3564
rect 34696 3508 34744 3564
rect 34800 3508 34838 3564
rect 34602 3460 34838 3508
rect 34602 3404 34640 3460
rect 34696 3404 34744 3460
rect 34800 3404 34838 3460
rect 34602 3394 34838 3404
rect 45022 1203 45514 1213
rect 45022 1147 45032 1203
rect 45088 1147 45136 1203
rect 45192 1147 45240 1203
rect 45296 1147 45344 1203
rect 45400 1147 45448 1203
rect 45504 1147 45514 1203
rect 35192 1103 35684 1113
rect 35192 1047 35202 1103
rect 35258 1047 35306 1103
rect 35362 1047 35410 1103
rect 35466 1047 35514 1103
rect 35570 1047 35618 1103
rect 35674 1047 35684 1103
rect 35192 999 35684 1047
rect 35192 943 35202 999
rect 35258 943 35306 999
rect 35362 943 35410 999
rect 35466 943 35514 999
rect 35570 943 35618 999
rect 35674 943 35684 999
rect 35192 895 35684 943
rect 35192 839 35202 895
rect 35258 839 35306 895
rect 35362 839 35410 895
rect 35466 839 35514 895
rect 35570 839 35618 895
rect 35674 839 35684 895
rect 35192 791 35684 839
rect 35192 735 35202 791
rect 35258 735 35306 791
rect 35362 735 35410 791
rect 35466 735 35514 791
rect 35570 735 35618 791
rect 35674 735 35684 791
rect 35192 687 35684 735
rect 35192 631 35202 687
rect 35258 631 35306 687
rect 35362 631 35410 687
rect 35466 631 35514 687
rect 35570 631 35618 687
rect 35674 631 35684 687
rect 35192 621 35684 631
rect 39632 1103 40124 1113
rect 39632 1047 39642 1103
rect 39698 1047 39746 1103
rect 39802 1047 39850 1103
rect 39906 1047 39954 1103
rect 40010 1047 40058 1103
rect 40114 1047 40124 1103
rect 39632 999 40124 1047
rect 39632 943 39642 999
rect 39698 943 39746 999
rect 39802 943 39850 999
rect 39906 943 39954 999
rect 40010 943 40058 999
rect 40114 943 40124 999
rect 39632 895 40124 943
rect 39632 839 39642 895
rect 39698 839 39746 895
rect 39802 839 39850 895
rect 39906 839 39954 895
rect 40010 839 40058 895
rect 40114 839 40124 895
rect 39632 791 40124 839
rect 39632 735 39642 791
rect 39698 735 39746 791
rect 39802 735 39850 791
rect 39906 735 39954 791
rect 40010 735 40058 791
rect 40114 735 40124 791
rect 39632 687 40124 735
rect 45022 1099 45514 1147
rect 45022 1043 45032 1099
rect 45088 1043 45136 1099
rect 45192 1043 45240 1099
rect 45296 1043 45344 1099
rect 45400 1043 45448 1099
rect 45504 1043 45514 1099
rect 45022 995 45514 1043
rect 45022 939 45032 995
rect 45088 939 45136 995
rect 45192 939 45240 995
rect 45296 939 45344 995
rect 45400 939 45448 995
rect 45504 939 45514 995
rect 45022 891 45514 939
rect 45022 835 45032 891
rect 45088 835 45136 891
rect 45192 835 45240 891
rect 45296 835 45344 891
rect 45400 835 45448 891
rect 45504 835 45514 891
rect 45022 787 45514 835
rect 45022 731 45032 787
rect 45088 731 45136 787
rect 45192 731 45240 787
rect 45296 731 45344 787
rect 45400 731 45448 787
rect 45504 731 45514 787
rect 45022 721 45514 731
rect 49462 1203 49954 1213
rect 49462 1147 49472 1203
rect 49528 1147 49576 1203
rect 49632 1147 49680 1203
rect 49736 1147 49784 1203
rect 49840 1147 49888 1203
rect 49944 1147 49954 1203
rect 49462 1099 49954 1147
rect 49462 1043 49472 1099
rect 49528 1043 49576 1099
rect 49632 1043 49680 1099
rect 49736 1043 49784 1099
rect 49840 1043 49888 1099
rect 49944 1043 49954 1099
rect 49462 995 49954 1043
rect 49462 939 49472 995
rect 49528 939 49576 995
rect 49632 939 49680 995
rect 49736 939 49784 995
rect 49840 939 49888 995
rect 49944 939 49954 995
rect 49462 891 49954 939
rect 49462 835 49472 891
rect 49528 835 49576 891
rect 49632 835 49680 891
rect 49736 835 49784 891
rect 49840 835 49888 891
rect 49944 835 49954 891
rect 49462 787 49954 835
rect 49462 731 49472 787
rect 49528 731 49576 787
rect 49632 731 49680 787
rect 49736 731 49784 787
rect 49840 731 49888 787
rect 49944 731 49954 787
rect 49462 721 49954 731
rect 39632 631 39642 687
rect 39698 631 39746 687
rect 39802 631 39850 687
rect 39906 631 39954 687
rect 40010 631 40058 687
rect 40114 631 40124 687
rect 39632 621 40124 631
rect 32126 330 32136 386
rect 32192 330 32240 386
rect 32296 330 32344 386
rect 32400 330 32410 386
rect 32126 282 32410 330
rect 32126 226 32136 282
rect 32192 226 32240 282
rect 32296 226 32344 282
rect 32400 226 32410 282
rect 32126 178 32410 226
rect 32126 122 32136 178
rect 32192 122 32240 178
rect 32296 122 32344 178
rect 32400 122 32410 178
rect 32126 112 32410 122
rect 15556 12 15568 64
rect 15620 12 15672 64
rect 15724 12 15776 64
rect 15828 12 15840 64
rect 15556 0 15840 12
<< via2 >>
rect 31226 15705 31282 15706
rect 31336 15705 31392 15706
rect 31446 15705 31502 15706
rect 31226 15653 31230 15705
rect 31230 15653 31282 15705
rect 31336 15653 31386 15705
rect 31386 15653 31392 15705
rect 31446 15653 31490 15705
rect 31490 15653 31502 15705
rect 31226 15650 31282 15653
rect 31336 15650 31392 15653
rect 31446 15650 31502 15653
rect 31226 15549 31230 15596
rect 31230 15549 31282 15596
rect 31336 15549 31386 15596
rect 31386 15549 31392 15596
rect 31446 15549 31490 15596
rect 31490 15549 31502 15596
rect 31226 15540 31282 15549
rect 31336 15540 31392 15549
rect 31446 15540 31502 15549
rect 31226 15445 31230 15486
rect 31230 15445 31282 15486
rect 31336 15445 31386 15486
rect 31386 15445 31392 15486
rect 31446 15445 31490 15486
rect 31490 15445 31502 15486
rect 31226 15430 31282 15445
rect 31336 15430 31392 15445
rect 31446 15430 31502 15445
rect 1233 14686 1289 14742
rect 1343 14686 1399 14742
rect 1453 14686 1509 14742
rect 1563 14686 1619 14742
rect 1233 14576 1289 14632
rect 1343 14576 1399 14632
rect 1453 14576 1509 14632
rect 1563 14576 1619 14632
rect -8163 12999 -8107 13055
rect -8053 12999 -7997 13055
rect 3171 14326 3227 14328
rect 3171 14274 3173 14326
rect 3173 14274 3225 14326
rect 3225 14274 3227 14326
rect 3171 14272 3227 14274
rect 3275 14326 3331 14328
rect 3275 14274 3277 14326
rect 3277 14274 3329 14326
rect 3329 14274 3331 14326
rect 3275 14272 3331 14274
rect 3171 14222 3227 14224
rect 3171 14170 3173 14222
rect 3173 14170 3225 14222
rect 3225 14170 3227 14222
rect 3171 14168 3227 14170
rect 3275 14222 3331 14224
rect 3275 14170 3277 14222
rect 3277 14170 3329 14222
rect 3329 14170 3331 14222
rect 3275 14168 3331 14170
rect 3960 14272 4016 14328
rect 3960 14222 4016 14224
rect 3960 14170 3962 14222
rect 3962 14170 4014 14222
rect 4014 14170 4016 14222
rect 3960 14168 4016 14170
rect 5741 14272 5797 14274
rect 5741 14220 5743 14272
rect 5743 14220 5795 14272
rect 5795 14220 5797 14272
rect 5741 14218 5797 14220
rect 5845 14272 5901 14274
rect 5845 14220 5847 14272
rect 5847 14220 5899 14272
rect 5899 14220 5901 14272
rect 5845 14218 5901 14220
rect -8163 12889 -8107 12945
rect -8053 12889 -7997 12945
rect -3604 10673 -3548 10729
rect -3494 10673 -3438 10729
rect -3604 10563 -3548 10619
rect -3494 10563 -3438 10619
rect -8141 9655 -8085 9711
rect -8031 9655 -7975 9711
rect -8141 9550 -8085 9606
rect -8031 9550 -7975 9606
rect -8141 9445 -8085 9501
rect -8031 9445 -7975 9501
rect -8491 8726 -8435 8782
rect -8381 8726 -8325 8782
rect -8491 8616 -8435 8672
rect -8381 8616 -8325 8672
rect -8491 8506 -8435 8562
rect -8381 8506 -8325 8562
rect -8491 8396 -8435 8452
rect -8381 8396 -8325 8452
rect -10576 7864 -10520 7920
rect -10466 7864 -10410 7920
rect -10356 7864 -10300 7920
rect -10246 7864 -10190 7920
rect -10576 7754 -10520 7810
rect -10466 7754 -10410 7810
rect -10356 7754 -10300 7810
rect -10246 7754 -10190 7810
rect 2530 13977 2586 13979
rect 2530 13925 2532 13977
rect 2532 13925 2584 13977
rect 2584 13925 2586 13977
rect 2530 13923 2586 13925
rect 2634 13977 2690 13979
rect 2634 13925 2636 13977
rect 2636 13925 2688 13977
rect 2688 13925 2690 13977
rect 2634 13923 2690 13925
rect 2530 13873 2586 13875
rect 2530 13821 2532 13873
rect 2532 13821 2584 13873
rect 2584 13821 2586 13873
rect 2530 13819 2586 13821
rect 2634 13873 2690 13875
rect 2634 13821 2636 13873
rect 2636 13821 2688 13873
rect 2688 13821 2690 13873
rect 2634 13819 2690 13821
rect 554 13707 610 13763
rect 664 13707 720 13763
rect 774 13707 830 13763
rect 884 13707 940 13763
rect 994 13707 1050 13763
rect 554 13597 610 13653
rect 664 13597 720 13653
rect 774 13597 830 13653
rect 884 13597 940 13653
rect 994 13597 1050 13653
rect -8146 5476 -8090 5532
rect -8041 5476 -7985 5532
rect -7936 5476 -7880 5532
rect -8146 5366 -8090 5422
rect -8041 5366 -7985 5422
rect -7936 5366 -7880 5422
rect -3604 4373 -3548 4429
rect -3494 4373 -3438 4429
rect -3604 4263 -3548 4319
rect -3494 4263 -3438 4319
rect 2891 13198 2947 13200
rect 2891 13146 2893 13198
rect 2893 13146 2945 13198
rect 2945 13146 2947 13198
rect 2891 13144 2947 13146
rect 2995 13198 3051 13200
rect 2995 13146 2997 13198
rect 2997 13146 3049 13198
rect 3049 13146 3051 13198
rect 2995 13144 3051 13146
rect 2891 13094 2947 13096
rect 2891 13042 2893 13094
rect 2893 13042 2945 13094
rect 2945 13042 2947 13094
rect 2891 13040 2947 13042
rect 2995 13094 3051 13096
rect 2995 13042 2997 13094
rect 2997 13042 3049 13094
rect 3049 13042 3051 13094
rect 2995 13040 3051 13042
rect 2530 12793 2586 12849
rect 2634 12793 2690 12849
rect 2530 12689 2586 12745
rect 2634 12689 2690 12745
rect 2530 10323 2586 10325
rect 2530 10271 2532 10323
rect 2532 10271 2584 10323
rect 2584 10271 2586 10323
rect 2530 10269 2586 10271
rect 2634 10323 2690 10325
rect 2634 10271 2636 10323
rect 2636 10271 2688 10323
rect 2688 10271 2690 10323
rect 2634 10269 2690 10271
rect 2530 10219 2586 10221
rect 2530 10167 2532 10219
rect 2532 10167 2584 10219
rect 2584 10167 2586 10219
rect 2530 10165 2586 10167
rect 2634 10219 2690 10221
rect 2634 10167 2636 10219
rect 2636 10167 2688 10219
rect 2688 10167 2690 10219
rect 2634 10165 2690 10167
rect 5741 14168 5797 14170
rect 5741 14116 5743 14168
rect 5743 14116 5795 14168
rect 5795 14116 5797 14168
rect 5741 14114 5797 14116
rect 5845 14168 5901 14170
rect 5845 14116 5847 14168
rect 5847 14116 5899 14168
rect 5899 14116 5901 14168
rect 5845 14114 5901 14116
rect 6745 14272 6801 14274
rect 6745 14220 6747 14272
rect 6747 14220 6799 14272
rect 6799 14220 6801 14272
rect 6745 14218 6801 14220
rect 6745 14168 6801 14170
rect 6745 14116 6747 14168
rect 6747 14116 6799 14168
rect 6799 14116 6801 14168
rect 6745 14114 6801 14116
rect 7385 14272 7441 14274
rect 7385 14220 7387 14272
rect 7387 14220 7439 14272
rect 7439 14220 7441 14272
rect 7385 14218 7441 14220
rect 7385 14168 7441 14170
rect 7385 14116 7387 14168
rect 7387 14116 7439 14168
rect 7439 14116 7441 14168
rect 7385 14114 7441 14116
rect 8025 14272 8081 14274
rect 8025 14220 8027 14272
rect 8027 14220 8079 14272
rect 8079 14220 8081 14272
rect 8025 14218 8081 14220
rect 8025 14168 8081 14170
rect 8025 14116 8027 14168
rect 8027 14116 8079 14168
rect 8079 14116 8081 14168
rect 8025 14114 8081 14116
rect 4040 13977 4096 13979
rect 4040 13925 4042 13977
rect 4042 13925 4094 13977
rect 4094 13925 4096 13977
rect 4040 13923 4096 13925
rect 4040 13873 4096 13875
rect 4040 13821 4042 13873
rect 4042 13821 4094 13873
rect 4094 13821 4096 13873
rect 4040 13819 4096 13821
rect 4200 13977 4256 13979
rect 4200 13925 4202 13977
rect 4202 13925 4254 13977
rect 4254 13925 4256 13977
rect 4200 13923 4256 13925
rect 4200 13873 4256 13875
rect 4200 13821 4202 13873
rect 4202 13821 4254 13873
rect 4254 13821 4256 13873
rect 4200 13819 4256 13821
rect 4841 13977 4897 13979
rect 4841 13925 4843 13977
rect 4843 13925 4895 13977
rect 4895 13925 4897 13977
rect 4841 13923 4897 13925
rect 4841 13873 4897 13875
rect 4841 13821 4843 13873
rect 4843 13821 4895 13873
rect 4895 13821 4897 13873
rect 4841 13819 4897 13821
rect 6013 13977 6069 13979
rect 6013 13925 6015 13977
rect 6015 13925 6067 13977
rect 6067 13925 6069 13977
rect 6013 13923 6069 13925
rect 6117 13977 6173 13979
rect 6117 13925 6119 13977
rect 6119 13925 6171 13977
rect 6171 13925 6173 13977
rect 6117 13923 6173 13925
rect 6013 13873 6069 13875
rect 6013 13821 6015 13873
rect 6015 13821 6067 13873
rect 6067 13821 6069 13873
rect 6013 13819 6069 13821
rect 6117 13873 6173 13875
rect 6117 13821 6119 13873
rect 6119 13821 6171 13873
rect 6171 13821 6173 13873
rect 6117 13819 6173 13821
rect 7065 13977 7121 13979
rect 7065 13925 7067 13977
rect 7067 13925 7119 13977
rect 7119 13925 7121 13977
rect 7065 13923 7121 13925
rect 7065 13873 7121 13875
rect 7065 13821 7067 13873
rect 7067 13821 7119 13873
rect 7119 13821 7121 13873
rect 7065 13819 7121 13821
rect 7705 13977 7761 13979
rect 7705 13925 7707 13977
rect 7707 13925 7759 13977
rect 7759 13925 7761 13977
rect 7705 13923 7761 13925
rect 7705 13873 7761 13875
rect 7705 13821 7707 13873
rect 7707 13821 7759 13873
rect 7759 13821 7761 13873
rect 7705 13819 7761 13821
rect 3880 13481 3936 13483
rect 3880 13429 3882 13481
rect 3882 13429 3934 13481
rect 3934 13429 3936 13481
rect 3880 13427 3936 13429
rect 3880 13377 3936 13379
rect 3880 13325 3882 13377
rect 3882 13325 3934 13377
rect 3934 13325 3936 13377
rect 3880 13323 3936 13325
rect 4520 13481 4576 13483
rect 4520 13429 4522 13481
rect 4522 13429 4574 13481
rect 4574 13429 4576 13481
rect 4520 13427 4576 13429
rect 4520 13377 4576 13379
rect 4520 13325 4522 13377
rect 4522 13325 4574 13377
rect 4574 13325 4576 13377
rect 4520 13323 4576 13325
rect 5160 13481 5216 13483
rect 5160 13429 5162 13481
rect 5162 13429 5214 13481
rect 5214 13429 5216 13481
rect 5160 13427 5216 13429
rect 5160 13377 5216 13379
rect 5160 13325 5162 13377
rect 5162 13325 5214 13377
rect 5214 13325 5216 13377
rect 5160 13323 5216 13325
rect 5741 13427 5797 13483
rect 5845 13427 5901 13483
rect 5741 13323 5797 13379
rect 5845 13323 5901 13379
rect 5741 13219 5797 13275
rect 5845 13219 5901 13275
rect 3960 13198 4016 13200
rect 3960 13146 3962 13198
rect 3962 13146 4014 13198
rect 4014 13146 4016 13198
rect 3960 13144 4016 13146
rect 3960 13094 4016 13096
rect 3960 13042 3962 13094
rect 3962 13042 4014 13094
rect 4014 13042 4016 13094
rect 3960 13040 4016 13042
rect 11649 13403 11705 13459
rect 11753 13403 11809 13459
rect 7065 13377 7121 13379
rect 7065 13325 7067 13377
rect 7067 13325 7119 13377
rect 7119 13325 7121 13377
rect 7065 13323 7121 13325
rect 7065 13273 7121 13275
rect 7065 13221 7067 13273
rect 7067 13221 7119 13273
rect 7119 13221 7121 13273
rect 7065 13219 7121 13221
rect 7705 13377 7761 13379
rect 7705 13325 7707 13377
rect 7707 13325 7759 13377
rect 7759 13325 7761 13377
rect 7705 13323 7761 13325
rect 11649 13299 11705 13355
rect 11753 13299 11809 13355
rect 17651 13351 17707 13407
rect 7705 13273 7761 13275
rect 7705 13221 7707 13273
rect 7707 13221 7759 13273
rect 7759 13221 7761 13273
rect 7705 13219 7761 13221
rect 6013 12944 6069 13000
rect 6117 12944 6173 13000
rect 4040 12847 4096 12849
rect 4040 12795 4042 12847
rect 4042 12795 4094 12847
rect 4094 12795 4096 12847
rect 4040 12793 4096 12795
rect 4040 12743 4096 12745
rect 4040 12691 4042 12743
rect 4042 12691 4094 12743
rect 4094 12691 4096 12743
rect 4040 12689 4096 12691
rect 4200 12847 4256 12849
rect 4200 12795 4202 12847
rect 4202 12795 4254 12847
rect 4254 12795 4256 12847
rect 4200 12793 4256 12795
rect 4200 12743 4256 12745
rect 4200 12691 4202 12743
rect 4202 12691 4254 12743
rect 4254 12691 4256 12743
rect 4200 12689 4256 12691
rect 4841 12847 4897 12849
rect 4841 12795 4843 12847
rect 4843 12795 4895 12847
rect 4895 12795 4897 12847
rect 4841 12793 4897 12795
rect 4841 12743 4897 12745
rect 4841 12691 4843 12743
rect 4843 12691 4895 12743
rect 4895 12691 4897 12743
rect 4841 12689 4897 12691
rect 5741 12793 5797 12849
rect 5845 12793 5901 12849
rect 6013 12840 6069 12896
rect 6117 12840 6173 12896
rect 6745 12998 6801 13000
rect 6745 12946 6747 12998
rect 6747 12946 6799 12998
rect 6799 12946 6801 12998
rect 6745 12944 6801 12946
rect 6745 12894 6801 12896
rect 6745 12842 6747 12894
rect 6747 12842 6799 12894
rect 6799 12842 6801 12894
rect 6745 12840 6801 12842
rect 7385 12998 7441 13000
rect 7385 12946 7387 12998
rect 7387 12946 7439 12998
rect 7439 12946 7441 12998
rect 7385 12944 7441 12946
rect 7385 12894 7441 12896
rect 7385 12842 7387 12894
rect 7387 12842 7439 12894
rect 7439 12842 7441 12894
rect 7385 12840 7441 12842
rect 8025 12998 8081 13000
rect 8025 12946 8027 12998
rect 8027 12946 8079 12998
rect 8079 12946 8081 12998
rect 8025 12944 8081 12946
rect 8025 12894 8081 12896
rect 8025 12842 8027 12894
rect 8027 12842 8079 12894
rect 8079 12842 8081 12894
rect 8025 12840 8081 12842
rect 5741 12689 5797 12745
rect 5845 12689 5901 12745
rect 3880 12455 3936 12457
rect 3880 12403 3882 12455
rect 3882 12403 3934 12455
rect 3934 12403 3936 12455
rect 3880 12401 3936 12403
rect 3880 12351 3936 12353
rect 3880 12299 3882 12351
rect 3882 12299 3934 12351
rect 3934 12299 3936 12351
rect 3880 12297 3936 12299
rect 4520 12455 4576 12457
rect 4520 12403 4522 12455
rect 4522 12403 4574 12455
rect 4574 12403 4576 12455
rect 4520 12401 4576 12403
rect 4520 12351 4576 12353
rect 4520 12299 4522 12351
rect 4522 12299 4574 12351
rect 4574 12299 4576 12351
rect 4520 12297 4576 12299
rect 5160 12455 5216 12457
rect 5160 12403 5162 12455
rect 5162 12403 5214 12455
rect 5214 12403 5216 12455
rect 5160 12401 5216 12403
rect 5160 12351 5216 12353
rect 5160 12299 5162 12351
rect 5162 12299 5214 12351
rect 5214 12299 5216 12351
rect 5160 12297 5216 12299
rect 6013 12401 6069 12457
rect 6117 12401 6173 12457
rect 6013 12297 6069 12353
rect 6117 12297 6173 12353
rect 7065 12455 7121 12457
rect 7065 12403 7067 12455
rect 7067 12403 7119 12455
rect 7119 12403 7121 12455
rect 7065 12401 7121 12403
rect 7065 12351 7121 12353
rect 7065 12299 7067 12351
rect 7067 12299 7119 12351
rect 7119 12299 7121 12351
rect 7065 12297 7121 12299
rect 7705 12455 7761 12457
rect 7705 12403 7707 12455
rect 7707 12403 7759 12455
rect 7759 12403 7761 12455
rect 7705 12401 7761 12403
rect 7705 12351 7761 12353
rect 7705 12299 7707 12351
rect 7707 12299 7759 12351
rect 7759 12299 7761 12351
rect 7705 12297 7761 12299
rect 11381 12437 11437 12493
rect 11485 12437 11541 12493
rect 11381 12333 11437 12389
rect 11485 12333 11541 12389
rect 5741 12082 5797 12138
rect 5845 12082 5901 12138
rect 3171 12014 3227 12070
rect 3275 12014 3331 12070
rect 3171 11910 3227 11966
rect 3275 11910 3331 11966
rect 3960 12068 4016 12070
rect 3960 12016 3962 12068
rect 3962 12016 4014 12068
rect 4014 12016 4016 12068
rect 3960 12014 4016 12016
rect 5741 11978 5797 12034
rect 5845 11978 5901 12034
rect 3960 11964 4016 11966
rect 3960 11912 3962 11964
rect 3962 11912 4014 11964
rect 4014 11912 4016 11964
rect 3960 11910 4016 11912
rect 2891 9756 2947 9812
rect 2995 9756 3051 9812
rect 2891 9652 2947 9708
rect 2995 9652 3051 9708
rect 2634 9457 2690 9459
rect 2634 9405 2636 9457
rect 2636 9405 2688 9457
rect 2688 9405 2690 9457
rect 2634 9403 2690 9405
rect 2634 9353 2690 9355
rect 2634 9301 2636 9353
rect 2636 9301 2688 9353
rect 2688 9301 2690 9353
rect 2634 9299 2690 9301
rect 2634 8127 2690 8129
rect 2634 8075 2636 8127
rect 2636 8075 2688 8127
rect 2688 8075 2690 8127
rect 2634 8073 2690 8075
rect 2634 8023 2690 8025
rect 2634 7971 2636 8023
rect 2636 7971 2688 8023
rect 2688 7971 2690 8023
rect 2634 7969 2690 7971
rect 236 7583 292 7585
rect 236 7531 238 7583
rect 238 7531 290 7583
rect 290 7531 292 7583
rect 236 7529 292 7531
rect 340 7583 396 7585
rect 340 7531 342 7583
rect 342 7531 394 7583
rect 394 7531 396 7583
rect 340 7529 396 7531
rect 236 7479 292 7481
rect 236 7427 238 7479
rect 238 7427 290 7479
rect 290 7427 292 7479
rect 236 7425 292 7427
rect 340 7479 396 7481
rect 340 7427 342 7479
rect 342 7427 394 7479
rect 394 7427 396 7479
rect 340 7425 396 7427
rect 1237 7583 1293 7585
rect 1237 7531 1239 7583
rect 1239 7531 1291 7583
rect 1291 7531 1293 7583
rect 1237 7529 1293 7531
rect 1341 7583 1397 7585
rect 1341 7531 1343 7583
rect 1343 7531 1395 7583
rect 1395 7531 1397 7583
rect 1341 7529 1397 7531
rect 4200 11717 4256 11719
rect 4200 11665 4202 11717
rect 4202 11665 4254 11717
rect 4254 11665 4256 11717
rect 4200 11663 4256 11665
rect 4200 11613 4256 11615
rect 4200 11561 4202 11613
rect 4202 11561 4254 11613
rect 4254 11561 4256 11613
rect 4200 11559 4256 11561
rect 4841 11717 4897 11719
rect 4841 11665 4843 11717
rect 4843 11665 4895 11717
rect 4895 11665 4897 11717
rect 4841 11663 4897 11665
rect 4841 11613 4897 11615
rect 4841 11561 4843 11613
rect 4843 11561 4895 11613
rect 4895 11561 4897 11613
rect 4841 11559 4897 11561
rect 6745 12136 6801 12138
rect 6745 12084 6747 12136
rect 6747 12084 6799 12136
rect 6799 12084 6801 12136
rect 6745 12082 6801 12084
rect 6745 12032 6801 12034
rect 6745 11980 6747 12032
rect 6747 11980 6799 12032
rect 6799 11980 6801 12032
rect 6745 11978 6801 11980
rect 7385 12136 7441 12138
rect 7385 12084 7387 12136
rect 7387 12084 7439 12136
rect 7439 12084 7441 12136
rect 7385 12082 7441 12084
rect 7385 12032 7441 12034
rect 7385 11980 7387 12032
rect 7387 11980 7439 12032
rect 7439 11980 7441 12032
rect 7385 11978 7441 11980
rect 8025 12136 8081 12138
rect 8025 12084 8027 12136
rect 8027 12084 8079 12136
rect 8079 12084 8081 12136
rect 8025 12082 8081 12084
rect 8025 12032 8081 12034
rect 8025 11980 8027 12032
rect 8027 11980 8079 12032
rect 8079 11980 8081 12032
rect 8025 11978 8081 11980
rect 6013 11663 6069 11719
rect 6117 11663 6173 11719
rect 6013 11559 6069 11615
rect 6117 11559 6173 11615
rect 6013 11455 6069 11511
rect 6117 11455 6173 11511
rect 6745 11613 6801 11615
rect 6745 11561 6747 11613
rect 6747 11561 6799 11613
rect 6799 11561 6801 11613
rect 6745 11559 6801 11561
rect 6745 11509 6801 11511
rect 6745 11457 6747 11509
rect 6747 11457 6799 11509
rect 6799 11457 6801 11509
rect 6745 11455 6801 11457
rect 7385 11613 7441 11615
rect 7385 11561 7387 11613
rect 7387 11561 7439 11613
rect 7439 11561 7441 11613
rect 7385 11559 7441 11561
rect 7385 11509 7441 11511
rect 7385 11457 7387 11509
rect 7387 11457 7439 11509
rect 7439 11457 7441 11509
rect 7385 11455 7441 11457
rect 8025 11613 8081 11615
rect 8025 11561 8027 11613
rect 8027 11561 8079 11613
rect 8079 11561 8081 11613
rect 8025 11559 8081 11561
rect 8025 11509 8081 11511
rect 8025 11457 8027 11509
rect 8027 11457 8079 11509
rect 8079 11457 8081 11509
rect 8025 11455 8081 11457
rect 5741 11271 5797 11327
rect 5845 11271 5901 11327
rect 3880 11221 3936 11223
rect 3880 11169 3882 11221
rect 3882 11169 3934 11221
rect 3934 11169 3936 11221
rect 3880 11167 3936 11169
rect 3880 11117 3936 11119
rect 3880 11065 3882 11117
rect 3882 11065 3934 11117
rect 3934 11065 3936 11117
rect 3880 11063 3936 11065
rect 4520 11221 4576 11223
rect 4520 11169 4522 11221
rect 4522 11169 4574 11221
rect 4574 11169 4576 11221
rect 4520 11167 4576 11169
rect 4520 11117 4576 11119
rect 4520 11065 4522 11117
rect 4522 11065 4574 11117
rect 4574 11065 4576 11117
rect 4520 11063 4576 11065
rect 5160 11221 5216 11223
rect 5160 11169 5162 11221
rect 5162 11169 5214 11221
rect 5214 11169 5216 11221
rect 5160 11167 5216 11169
rect 5160 11117 5216 11119
rect 5160 11065 5162 11117
rect 5162 11065 5214 11117
rect 5214 11065 5216 11117
rect 5160 11063 5216 11065
rect 5741 11167 5797 11223
rect 5845 11167 5901 11223
rect 5741 11063 5797 11119
rect 5845 11063 5901 11119
rect 5741 10740 5797 10796
rect 5845 10740 5901 10796
rect 5741 10636 5797 10692
rect 5845 10636 5901 10692
rect 4040 10323 4096 10325
rect 4040 10271 4042 10323
rect 4042 10271 4094 10323
rect 4094 10271 4096 10323
rect 4040 10269 4096 10271
rect 4040 10219 4096 10221
rect 4040 10167 4042 10219
rect 4042 10167 4094 10219
rect 4094 10167 4096 10219
rect 4040 10165 4096 10167
rect 3960 9810 4016 9812
rect 3960 9758 3962 9810
rect 3962 9758 4014 9810
rect 4014 9758 4016 9810
rect 3960 9756 4016 9758
rect 3960 9706 4016 9708
rect 3960 9654 3962 9706
rect 3962 9654 4014 9706
rect 4014 9654 4016 9706
rect 3960 9652 4016 9654
rect 7065 11325 7121 11327
rect 7065 11273 7067 11325
rect 7067 11273 7119 11325
rect 7119 11273 7121 11325
rect 7065 11271 7121 11273
rect 7065 11221 7121 11223
rect 7065 11169 7067 11221
rect 7067 11169 7119 11221
rect 7119 11169 7121 11221
rect 7065 11167 7121 11169
rect 7705 11325 7761 11327
rect 7705 11273 7707 11325
rect 7707 11273 7759 11325
rect 7759 11273 7761 11325
rect 7705 11271 7761 11273
rect 7705 11221 7761 11223
rect 7705 11169 7707 11221
rect 7707 11169 7759 11221
rect 7759 11169 7761 11221
rect 7705 11167 7761 11169
rect 11381 11373 11437 11375
rect 11381 11321 11383 11373
rect 11383 11321 11435 11373
rect 11435 11321 11437 11373
rect 11381 11319 11437 11321
rect 11485 11373 11541 11375
rect 11485 11321 11487 11373
rect 11487 11321 11539 11373
rect 11539 11321 11541 11373
rect 11485 11319 11541 11321
rect 11381 11269 11437 11271
rect 11381 11217 11383 11269
rect 11383 11217 11435 11269
rect 11435 11217 11437 11269
rect 11381 11215 11437 11217
rect 11485 11269 11541 11271
rect 11485 11217 11487 11269
rect 11487 11217 11539 11269
rect 11539 11217 11541 11269
rect 11485 11215 11541 11217
rect 8980 10794 9036 10796
rect 8980 10742 8982 10794
rect 8982 10742 9034 10794
rect 9034 10742 9036 10794
rect 8980 10740 9036 10742
rect 8980 10690 9036 10692
rect 8980 10638 8982 10690
rect 8982 10638 9034 10690
rect 9034 10638 9036 10690
rect 8980 10636 9036 10638
rect 9876 10794 9932 10796
rect 9876 10742 9878 10794
rect 9878 10742 9930 10794
rect 9930 10742 9932 10794
rect 9876 10740 9932 10742
rect 9876 10690 9932 10692
rect 9876 10638 9878 10690
rect 9878 10638 9930 10690
rect 9930 10638 9932 10690
rect 9876 10636 9932 10638
rect 10772 10794 10828 10796
rect 10772 10742 10774 10794
rect 10774 10742 10826 10794
rect 10826 10742 10828 10794
rect 10772 10740 10828 10742
rect 10772 10690 10828 10692
rect 10772 10638 10774 10690
rect 10774 10638 10826 10690
rect 10826 10638 10828 10690
rect 10772 10636 10828 10638
rect 6013 10369 6069 10425
rect 6117 10369 6173 10425
rect 6013 10265 6069 10321
rect 6117 10265 6173 10321
rect 9428 10423 9484 10425
rect 9428 10371 9430 10423
rect 9430 10371 9482 10423
rect 9482 10371 9484 10423
rect 9428 10369 9484 10371
rect 9428 10319 9484 10321
rect 9428 10267 9430 10319
rect 9430 10267 9482 10319
rect 9482 10267 9484 10319
rect 9428 10265 9484 10267
rect 10324 10423 10380 10425
rect 10324 10371 10326 10423
rect 10326 10371 10378 10423
rect 10378 10371 10380 10423
rect 10324 10369 10380 10371
rect 10324 10319 10380 10321
rect 10324 10267 10326 10319
rect 10326 10267 10378 10319
rect 10378 10267 10380 10319
rect 10324 10265 10380 10267
rect 10612 10423 10668 10425
rect 10612 10371 10614 10423
rect 10614 10371 10666 10423
rect 10666 10371 10668 10423
rect 10612 10369 10668 10371
rect 10612 10319 10668 10321
rect 10612 10267 10614 10319
rect 10614 10267 10666 10319
rect 10666 10267 10668 10319
rect 10612 10265 10668 10267
rect 6013 9908 6069 9964
rect 6117 9908 6173 9964
rect 6013 9804 6069 9860
rect 6117 9804 6173 9860
rect 7065 9962 7121 9964
rect 7065 9910 7067 9962
rect 7067 9910 7119 9962
rect 7119 9910 7121 9962
rect 7065 9908 7121 9910
rect 7065 9858 7121 9860
rect 7065 9806 7067 9858
rect 7067 9806 7119 9858
rect 7119 9806 7121 9858
rect 7065 9804 7121 9806
rect 7705 9962 7761 9964
rect 7705 9910 7707 9962
rect 7707 9910 7759 9962
rect 7759 9910 7761 9962
rect 7705 9908 7761 9910
rect 7705 9858 7761 9860
rect 7705 9806 7707 9858
rect 7707 9806 7759 9858
rect 7759 9806 7761 9858
rect 7705 9804 7761 9806
rect 5741 9507 5797 9563
rect 5845 9507 5901 9563
rect 4040 9457 4096 9459
rect 4040 9405 4042 9457
rect 4042 9405 4094 9457
rect 4094 9405 4096 9457
rect 4040 9403 4096 9405
rect 4040 9353 4096 9355
rect 4040 9301 4042 9353
rect 4042 9301 4094 9353
rect 4094 9301 4096 9353
rect 4040 9299 4096 9301
rect 4200 9457 4256 9459
rect 4200 9405 4202 9457
rect 4202 9405 4254 9457
rect 4254 9405 4256 9457
rect 4200 9403 4256 9405
rect 4200 9353 4256 9355
rect 4200 9301 4202 9353
rect 4202 9301 4254 9353
rect 4254 9301 4256 9353
rect 4200 9299 4256 9301
rect 4841 9457 4897 9459
rect 4841 9405 4843 9457
rect 4843 9405 4895 9457
rect 4895 9405 4897 9457
rect 4841 9403 4897 9405
rect 4841 9353 4897 9355
rect 4841 9301 4843 9353
rect 4843 9301 4895 9353
rect 4895 9301 4897 9353
rect 4841 9299 4897 9301
rect 5741 9403 5797 9459
rect 5845 9403 5901 9459
rect 5741 9299 5797 9355
rect 5845 9299 5901 9355
rect 3880 8961 3936 8963
rect 3880 8909 3882 8961
rect 3882 8909 3934 8961
rect 3934 8909 3936 8961
rect 3880 8907 3936 8909
rect 3880 8857 3936 8859
rect 3880 8805 3882 8857
rect 3882 8805 3934 8857
rect 3934 8805 3936 8857
rect 3880 8803 3936 8805
rect 4520 8961 4576 8963
rect 4520 8909 4522 8961
rect 4522 8909 4574 8961
rect 4574 8909 4576 8961
rect 4520 8907 4576 8909
rect 4520 8857 4576 8859
rect 4520 8805 4522 8857
rect 4522 8805 4574 8857
rect 4574 8805 4576 8857
rect 4520 8803 4576 8805
rect 5160 8961 5216 8963
rect 5160 8909 5162 8961
rect 5162 8909 5214 8961
rect 5214 8909 5216 8961
rect 5160 8907 5216 8909
rect 5160 8857 5216 8859
rect 5160 8805 5162 8857
rect 5162 8805 5214 8857
rect 5214 8805 5216 8857
rect 5160 8803 5216 8805
rect 19075 13405 19131 13407
rect 19075 13353 19077 13405
rect 19077 13353 19129 13405
rect 19129 13353 19131 13405
rect 19075 13351 19131 13353
rect 20195 13405 20251 13407
rect 20195 13353 20197 13405
rect 20197 13353 20249 13405
rect 20249 13353 20251 13405
rect 20195 13351 20251 13353
rect 24227 13405 24283 13407
rect 24227 13353 24229 13405
rect 24229 13353 24281 13405
rect 24281 13353 24283 13405
rect 24227 13351 24283 13353
rect 25347 13405 25403 13407
rect 25347 13353 25349 13405
rect 25349 13353 25401 13405
rect 25401 13353 25403 13405
rect 25347 13351 25403 13353
rect 26771 13351 26828 13407
rect 22107 13214 22163 13270
rect 22211 13214 22267 13270
rect 22315 13214 22371 13270
rect 19315 13164 19371 13166
rect 19315 13112 19317 13164
rect 19317 13112 19369 13164
rect 19369 13112 19371 13164
rect 19315 13110 19371 13112
rect 19315 13060 19371 13062
rect 19315 13008 19317 13060
rect 19317 13008 19369 13060
rect 19369 13008 19371 13060
rect 19315 13006 19371 13008
rect 19955 13164 20011 13166
rect 19955 13112 19957 13164
rect 19957 13112 20009 13164
rect 20009 13112 20011 13164
rect 19955 13110 20011 13112
rect 19955 13060 20011 13062
rect 19955 13008 19957 13060
rect 19957 13008 20009 13060
rect 20009 13008 20011 13060
rect 19955 13006 20011 13008
rect 22107 13110 22163 13166
rect 22211 13110 22267 13166
rect 22315 13110 22371 13166
rect 22107 13006 22163 13062
rect 22211 13006 22267 13062
rect 22315 13006 22371 13062
rect 21458 12820 21514 12876
rect 21562 12820 21618 12876
rect 21666 12820 21722 12876
rect 18995 12770 19051 12772
rect 18995 12718 18997 12770
rect 18997 12718 19049 12770
rect 19049 12718 19051 12770
rect 18995 12716 19051 12718
rect 18995 12666 19051 12668
rect 18995 12614 18997 12666
rect 18997 12614 19049 12666
rect 19049 12614 19051 12666
rect 18995 12612 19051 12614
rect 19635 12770 19691 12772
rect 19635 12718 19637 12770
rect 19637 12718 19689 12770
rect 19689 12718 19691 12770
rect 19635 12716 19691 12718
rect 19635 12666 19691 12668
rect 19635 12614 19637 12666
rect 19637 12614 19689 12666
rect 19689 12614 19691 12666
rect 19635 12612 19691 12614
rect 20275 12770 20331 12772
rect 20275 12718 20277 12770
rect 20277 12718 20329 12770
rect 20329 12718 20331 12770
rect 20275 12716 20331 12718
rect 20275 12666 20331 12668
rect 20275 12614 20277 12666
rect 20277 12614 20329 12666
rect 20329 12614 20331 12666
rect 20275 12612 20331 12614
rect 21458 12716 21514 12772
rect 21562 12716 21618 12772
rect 21666 12716 21722 12772
rect 21458 12612 21514 12668
rect 21562 12612 21618 12668
rect 21666 12612 21722 12668
rect 17651 11449 17707 11505
rect 12810 11373 12866 11375
rect 12810 11321 12812 11373
rect 12812 11321 12864 11373
rect 12864 11321 12866 11373
rect 12810 11319 12866 11321
rect 12810 11269 12866 11271
rect 12810 11217 12812 11269
rect 12812 11217 12864 11269
rect 12864 11217 12866 11269
rect 12810 11215 12866 11217
rect 13706 11373 13762 11375
rect 13706 11321 13708 11373
rect 13708 11321 13760 11373
rect 13760 11321 13762 11373
rect 13706 11319 13762 11321
rect 13706 11269 13762 11271
rect 13706 11217 13708 11269
rect 13708 11217 13760 11269
rect 13760 11217 13762 11269
rect 13706 11215 13762 11217
rect 13994 11373 14050 11375
rect 13994 11321 13996 11373
rect 13996 11321 14048 11373
rect 14048 11321 14050 11373
rect 13994 11319 14050 11321
rect 13994 11269 14050 11271
rect 13994 11217 13996 11269
rect 13996 11217 14048 11269
rect 14048 11217 14050 11269
rect 13994 11215 14050 11217
rect 15156 11373 15212 11375
rect 15156 11321 15158 11373
rect 15158 11321 15210 11373
rect 15210 11321 15212 11373
rect 15156 11319 15212 11321
rect 15156 11269 15212 11271
rect 15156 11217 15158 11269
rect 15158 11217 15210 11269
rect 15210 11217 15212 11269
rect 15156 11215 15212 11217
rect 15796 11373 15852 11375
rect 15796 11321 15798 11373
rect 15798 11321 15850 11373
rect 15850 11321 15852 11373
rect 15796 11319 15852 11321
rect 15796 11269 15852 11271
rect 15796 11217 15798 11269
rect 15798 11217 15850 11269
rect 15850 11217 15852 11269
rect 15796 11215 15852 11217
rect 16436 11373 16492 11375
rect 16436 11321 16438 11373
rect 16438 11321 16490 11373
rect 16490 11321 16492 11373
rect 16436 11319 16492 11321
rect 16436 11269 16492 11271
rect 16436 11217 16438 11269
rect 16438 11217 16490 11269
rect 16490 11217 16492 11269
rect 16436 11215 16492 11217
rect 17375 11373 17431 11375
rect 17375 11321 17377 11373
rect 17377 11321 17429 11373
rect 17429 11321 17431 11373
rect 17375 11319 17431 11321
rect 17479 11373 17535 11375
rect 17479 11321 17481 11373
rect 17481 11321 17533 11373
rect 17533 11321 17535 11373
rect 17479 11319 17535 11321
rect 17375 11269 17431 11271
rect 17375 11217 17377 11269
rect 17377 11217 17429 11269
rect 17429 11217 17431 11269
rect 17375 11215 17431 11217
rect 17479 11269 17535 11271
rect 17479 11217 17481 11269
rect 17481 11217 17533 11269
rect 17533 11217 17535 11269
rect 17479 11215 17535 11217
rect 11649 10953 11705 10955
rect 11649 10901 11651 10953
rect 11651 10901 11703 10953
rect 11703 10901 11705 10953
rect 11649 10899 11705 10901
rect 11753 10953 11809 10955
rect 11753 10901 11755 10953
rect 11755 10901 11807 10953
rect 11807 10901 11809 10953
rect 11753 10899 11809 10901
rect 11649 10849 11705 10851
rect 11649 10797 11651 10849
rect 11651 10797 11703 10849
rect 11703 10797 11705 10849
rect 11649 10795 11705 10797
rect 11753 10849 11809 10851
rect 11753 10797 11755 10849
rect 11755 10797 11807 10849
rect 11807 10797 11809 10849
rect 11753 10795 11809 10797
rect 12362 10953 12418 10955
rect 12362 10901 12364 10953
rect 12364 10901 12416 10953
rect 12416 10901 12418 10953
rect 12362 10899 12418 10901
rect 12362 10849 12418 10851
rect 12362 10797 12364 10849
rect 12364 10797 12416 10849
rect 12416 10797 12418 10849
rect 12362 10795 12418 10797
rect 13258 10953 13314 10955
rect 13258 10901 13260 10953
rect 13260 10901 13312 10953
rect 13312 10901 13314 10953
rect 13258 10899 13314 10901
rect 13258 10849 13314 10851
rect 13258 10797 13260 10849
rect 13260 10797 13312 10849
rect 13312 10797 13314 10849
rect 13258 10795 13314 10797
rect 14154 10953 14210 10955
rect 14154 10901 14156 10953
rect 14156 10901 14208 10953
rect 14208 10901 14210 10953
rect 14154 10899 14210 10901
rect 14154 10849 14210 10851
rect 14154 10797 14156 10849
rect 14156 10797 14208 10849
rect 14208 10797 14210 10849
rect 14154 10795 14210 10797
rect 15476 10953 15532 10955
rect 15476 10901 15478 10953
rect 15478 10901 15530 10953
rect 15530 10901 15532 10953
rect 15476 10899 15532 10901
rect 15476 10849 15532 10851
rect 15476 10797 15478 10849
rect 15478 10797 15530 10849
rect 15530 10797 15532 10849
rect 15476 10795 15532 10797
rect 16116 10953 16172 10955
rect 16116 10901 16118 10953
rect 16118 10901 16170 10953
rect 16170 10901 16172 10953
rect 16116 10899 16172 10901
rect 16116 10849 16172 10851
rect 16116 10797 16118 10849
rect 16118 10797 16170 10849
rect 16170 10797 16172 10849
rect 16116 10795 16172 10797
rect 17113 10953 17169 10955
rect 17113 10901 17115 10953
rect 17115 10901 17167 10953
rect 17167 10901 17169 10953
rect 17113 10899 17169 10901
rect 17217 10953 17273 10955
rect 17217 10901 17219 10953
rect 17219 10901 17271 10953
rect 17271 10901 17273 10953
rect 17217 10899 17273 10901
rect 17113 10849 17169 10851
rect 17113 10797 17115 10849
rect 17115 10797 17167 10849
rect 17167 10797 17169 10849
rect 17113 10795 17169 10797
rect 17217 10849 17273 10851
rect 17217 10797 17219 10849
rect 17219 10797 17271 10849
rect 17271 10797 17273 10849
rect 17217 10795 17273 10797
rect 11649 10369 11705 10425
rect 11753 10369 11809 10425
rect 11649 10265 11705 10321
rect 11753 10265 11809 10321
rect 11649 10161 11705 10217
rect 11753 10161 11809 10217
rect 12810 10319 12866 10321
rect 12810 10267 12812 10319
rect 12812 10267 12864 10319
rect 12864 10267 12866 10319
rect 12810 10265 12866 10267
rect 12810 10215 12866 10217
rect 12810 10163 12812 10215
rect 12812 10163 12864 10215
rect 12864 10163 12866 10215
rect 12810 10161 12866 10163
rect 13706 10319 13762 10321
rect 13706 10267 13708 10319
rect 13708 10267 13760 10319
rect 13760 10267 13762 10319
rect 13706 10265 13762 10267
rect 13706 10215 13762 10217
rect 13706 10163 13708 10215
rect 13708 10163 13760 10215
rect 13760 10163 13762 10215
rect 13706 10161 13762 10163
rect 13994 10293 14050 10295
rect 13994 10241 13996 10293
rect 13996 10241 14048 10293
rect 14048 10241 14050 10293
rect 13994 10239 14050 10241
rect 10612 9761 10668 9763
rect 10612 9709 10614 9761
rect 10614 9709 10666 9761
rect 10666 9709 10668 9761
rect 10612 9707 10668 9709
rect 10612 9657 10668 9659
rect 10612 9605 10614 9657
rect 10614 9605 10666 9657
rect 10666 9605 10668 9657
rect 10612 9603 10668 9605
rect 11381 9707 11437 9763
rect 11485 9707 11541 9763
rect 11381 9603 11437 9659
rect 11485 9603 11541 9659
rect 6745 9561 6801 9563
rect 6745 9509 6747 9561
rect 6747 9509 6799 9561
rect 6799 9509 6801 9561
rect 6745 9507 6801 9509
rect 6745 9457 6801 9459
rect 6745 9405 6747 9457
rect 6747 9405 6799 9457
rect 6799 9405 6801 9457
rect 6745 9403 6801 9405
rect 7385 9561 7441 9563
rect 7385 9509 7387 9561
rect 7387 9509 7439 9561
rect 7439 9509 7441 9561
rect 7385 9507 7441 9509
rect 7385 9457 7441 9459
rect 7385 9405 7387 9457
rect 7387 9405 7439 9457
rect 7439 9405 7441 9457
rect 7385 9403 7441 9405
rect 8025 9561 8081 9563
rect 8025 9509 8027 9561
rect 8027 9509 8079 9561
rect 8079 9509 8081 9561
rect 8025 9507 8081 9509
rect 8025 9457 8081 9459
rect 8025 9405 8027 9457
rect 8027 9405 8079 9457
rect 8079 9405 8081 9457
rect 8025 9403 8081 9405
rect 9428 9561 9484 9563
rect 9428 9509 9430 9561
rect 9430 9509 9482 9561
rect 9482 9509 9484 9561
rect 9428 9507 9484 9509
rect 9428 9457 9484 9459
rect 9428 9405 9430 9457
rect 9430 9405 9482 9457
rect 9482 9405 9484 9457
rect 9428 9403 9484 9405
rect 10324 9561 10380 9563
rect 10324 9509 10326 9561
rect 10326 9509 10378 9561
rect 10378 9509 10380 9561
rect 10324 9507 10380 9509
rect 10324 9457 10380 9459
rect 10324 9405 10326 9457
rect 10326 9405 10378 9457
rect 10378 9405 10380 9457
rect 10324 9403 10380 9405
rect 11381 9219 11437 9275
rect 11485 9219 11541 9275
rect 11381 9115 11437 9171
rect 11485 9115 11541 9171
rect 6013 8907 6069 8963
rect 6117 8907 6173 8963
rect 6013 8803 6069 8859
rect 6117 8803 6173 8859
rect 6745 8961 6801 8963
rect 6745 8909 6747 8961
rect 6747 8909 6799 8961
rect 6799 8909 6801 8961
rect 6745 8907 6801 8909
rect 6745 8857 6801 8859
rect 6745 8805 6747 8857
rect 6747 8805 6799 8857
rect 6799 8805 6801 8857
rect 6745 8803 6801 8805
rect 7385 8961 7441 8963
rect 7385 8909 7387 8961
rect 7387 8909 7439 8961
rect 7439 8909 7441 8961
rect 7385 8907 7441 8909
rect 7385 8857 7441 8859
rect 7385 8805 7387 8857
rect 7387 8805 7439 8857
rect 7439 8805 7441 8857
rect 7385 8803 7441 8805
rect 8025 8961 8081 8963
rect 8025 8909 8027 8961
rect 8027 8909 8079 8961
rect 8079 8909 8081 8961
rect 8025 8907 8081 8909
rect 8025 8857 8081 8859
rect 8025 8805 8027 8857
rect 8027 8805 8079 8857
rect 8079 8805 8081 8857
rect 8025 8803 8081 8805
rect 8980 8961 9036 8963
rect 8980 8909 8982 8961
rect 8982 8909 9034 8961
rect 9034 8909 9036 8961
rect 8980 8907 9036 8909
rect 8980 8857 9036 8859
rect 8980 8805 8982 8857
rect 8982 8805 9034 8857
rect 9034 8805 9036 8857
rect 8980 8803 9036 8805
rect 9876 8961 9932 8963
rect 9876 8909 9878 8961
rect 9878 8909 9930 8961
rect 9930 8909 9932 8961
rect 9876 8907 9932 8909
rect 9876 8857 9932 8859
rect 9876 8805 9878 8857
rect 9878 8805 9930 8857
rect 9930 8805 9932 8857
rect 9876 8803 9932 8805
rect 10772 8961 10828 8963
rect 10772 8909 10774 8961
rect 10774 8909 10826 8961
rect 10826 8909 10828 8961
rect 10772 8907 10828 8909
rect 10772 8857 10828 8859
rect 10772 8805 10774 8857
rect 10774 8805 10826 8857
rect 10826 8805 10828 8857
rect 10772 8803 10828 8805
rect 3171 8626 3227 8682
rect 3275 8626 3331 8682
rect 3171 8522 3227 8578
rect 3275 8522 3331 8578
rect 3960 8680 4016 8682
rect 3960 8628 3962 8680
rect 3962 8628 4014 8680
rect 4014 8628 4016 8680
rect 3960 8626 4016 8628
rect 3960 8576 4016 8578
rect 3960 8524 3962 8576
rect 3962 8524 4014 8576
rect 4014 8524 4016 8576
rect 3960 8522 4016 8524
rect 5741 8634 5797 8690
rect 5845 8634 5901 8690
rect 5741 8530 5797 8586
rect 5845 8530 5901 8586
rect 4200 8327 4256 8329
rect 4200 8275 4202 8327
rect 4202 8275 4254 8327
rect 4254 8275 4256 8327
rect 4200 8273 4256 8275
rect 4200 8223 4256 8225
rect 4200 8171 4202 8223
rect 4202 8171 4254 8223
rect 4254 8171 4256 8223
rect 4200 8169 4256 8171
rect 4841 8327 4897 8329
rect 4841 8275 4843 8327
rect 4843 8275 4895 8327
rect 4895 8275 4897 8327
rect 4841 8273 4897 8275
rect 4841 8223 4897 8225
rect 4841 8171 4843 8223
rect 4843 8171 4895 8223
rect 4895 8171 4897 8223
rect 4841 8169 4897 8171
rect 4040 8127 4096 8129
rect 4040 8075 4042 8127
rect 4042 8075 4094 8127
rect 4094 8075 4096 8127
rect 4040 8073 4096 8075
rect 4040 8023 4096 8025
rect 4040 7971 4042 8023
rect 4042 7971 4094 8023
rect 4094 7971 4096 8023
rect 4040 7969 4096 7971
rect 7065 8688 7121 8690
rect 7065 8636 7067 8688
rect 7067 8636 7119 8688
rect 7119 8636 7121 8688
rect 7065 8634 7121 8636
rect 7065 8584 7121 8586
rect 7065 8532 7067 8584
rect 7067 8532 7119 8584
rect 7119 8532 7121 8584
rect 7065 8530 7121 8532
rect 7705 8688 7761 8690
rect 7705 8636 7707 8688
rect 7707 8636 7759 8688
rect 7759 8636 7761 8688
rect 7705 8634 7761 8636
rect 7705 8584 7761 8586
rect 7705 8532 7707 8584
rect 7707 8532 7759 8584
rect 7759 8532 7761 8584
rect 7705 8530 7761 8532
rect 10484 8703 10540 8705
rect 10484 8651 10486 8703
rect 10486 8651 10538 8703
rect 10538 8651 10540 8703
rect 10484 8649 10540 8651
rect 10484 8599 10540 8601
rect 10484 8547 10486 8599
rect 10486 8547 10538 8599
rect 10538 8547 10540 8599
rect 10484 8545 10540 8547
rect 7999 8464 8055 8466
rect 7999 8412 8001 8464
rect 8001 8412 8053 8464
rect 8053 8412 8055 8464
rect 7999 8410 8055 8412
rect 6013 8273 6069 8329
rect 6117 8273 6173 8329
rect 7999 8360 8055 8362
rect 7999 8308 8001 8360
rect 8001 8308 8053 8360
rect 8053 8308 8055 8360
rect 7999 8306 8055 8308
rect 8285 8410 8341 8466
rect 8389 8410 8445 8466
rect 8285 8306 8341 8362
rect 8389 8306 8445 8362
rect 10732 8453 10788 8455
rect 10732 8401 10734 8453
rect 10734 8401 10786 8453
rect 10786 8401 10788 8453
rect 10732 8399 10788 8401
rect 6013 8169 6069 8225
rect 6117 8169 6173 8225
rect 6013 8065 6069 8121
rect 6117 8065 6173 8121
rect 7065 8223 7121 8225
rect 7065 8171 7067 8223
rect 7067 8171 7119 8223
rect 7119 8171 7121 8223
rect 7065 8169 7121 8171
rect 7065 8119 7121 8121
rect 7065 8067 7067 8119
rect 7067 8067 7119 8119
rect 7119 8067 7121 8119
rect 7065 8065 7121 8067
rect 7705 8223 7761 8225
rect 7705 8171 7707 8223
rect 7707 8171 7759 8223
rect 7759 8171 7761 8223
rect 7705 8169 7761 8171
rect 7705 8119 7761 8121
rect 7705 8067 7707 8119
rect 7707 8067 7759 8119
rect 7759 8067 7761 8119
rect 7705 8065 7761 8067
rect 3880 7831 3936 7833
rect 3880 7779 3882 7831
rect 3882 7779 3934 7831
rect 3934 7779 3936 7831
rect 3880 7777 3936 7779
rect 3880 7727 3936 7729
rect 3880 7675 3882 7727
rect 3882 7675 3934 7727
rect 3934 7675 3936 7727
rect 3880 7673 3936 7675
rect 4520 7831 4576 7833
rect 4520 7779 4522 7831
rect 4522 7779 4574 7831
rect 4574 7779 4576 7831
rect 4520 7777 4576 7779
rect 4520 7727 4576 7729
rect 4520 7675 4522 7727
rect 4522 7675 4574 7727
rect 4574 7675 4576 7727
rect 4520 7673 4576 7675
rect 5160 7831 5216 7833
rect 5160 7779 5162 7831
rect 5162 7779 5214 7831
rect 5214 7779 5216 7831
rect 5160 7777 5216 7779
rect 5160 7727 5216 7729
rect 5160 7675 5162 7727
rect 5162 7675 5214 7727
rect 5214 7675 5216 7727
rect 5160 7673 5216 7675
rect 5741 7777 5797 7833
rect 5845 7777 5901 7833
rect 5741 7673 5797 7729
rect 5845 7673 5901 7729
rect 6745 7831 6801 7833
rect 6745 7779 6747 7831
rect 6747 7779 6799 7831
rect 6799 7779 6801 7831
rect 6745 7777 6801 7779
rect 6745 7727 6801 7729
rect 6745 7675 6747 7727
rect 6747 7675 6799 7727
rect 6799 7675 6801 7727
rect 6745 7673 6801 7675
rect 7385 7831 7441 7833
rect 7385 7779 7387 7831
rect 7387 7779 7439 7831
rect 7439 7779 7441 7831
rect 7385 7777 7441 7779
rect 7385 7727 7441 7729
rect 7385 7675 7387 7727
rect 7387 7675 7439 7727
rect 7439 7675 7441 7727
rect 7385 7673 7441 7675
rect 8025 7831 8081 7833
rect 8025 7779 8027 7831
rect 8027 7779 8079 7831
rect 8079 7779 8081 7831
rect 8025 7777 8081 7779
rect 8025 7727 8081 7729
rect 8025 7675 8027 7727
rect 8027 7675 8079 7727
rect 8079 7675 8081 7727
rect 8025 7673 8081 7675
rect 1237 7425 1293 7481
rect 1341 7425 1397 7481
rect 2891 7438 2947 7494
rect 2995 7438 3051 7494
rect 2891 7334 2947 7390
rect 2995 7334 3051 7390
rect 4120 7492 4176 7494
rect 4120 7440 4122 7492
rect 4122 7440 4174 7492
rect 4174 7440 4176 7492
rect 4120 7438 4176 7440
rect 4120 7334 4176 7390
rect 10732 8349 10788 8351
rect 10732 8297 10734 8349
rect 10734 8297 10786 8349
rect 10786 8297 10788 8349
rect 10732 8295 10788 8297
rect 10928 8399 10984 8455
rect 11032 8399 11088 8455
rect 10928 8295 10984 8351
rect 11032 8295 11088 8351
rect 9428 8223 9484 8225
rect 9428 8171 9430 8223
rect 9430 8171 9482 8223
rect 9482 8171 9484 8223
rect 9428 8169 9484 8171
rect 9428 8119 9484 8121
rect 9428 8067 9430 8119
rect 9430 8067 9482 8119
rect 9482 8067 9484 8119
rect 9428 8065 9484 8067
rect 10324 8223 10380 8225
rect 10324 8171 10326 8223
rect 10326 8171 10378 8223
rect 10378 8171 10380 8223
rect 10324 8169 10380 8171
rect 10324 8119 10380 8121
rect 10324 8067 10326 8119
rect 10326 8067 10378 8119
rect 10378 8067 10380 8119
rect 10324 8065 10380 8067
rect 10484 8223 10540 8225
rect 10484 8171 10486 8223
rect 10486 8171 10538 8223
rect 10538 8171 10540 8223
rect 10484 8169 10540 8171
rect 10484 8119 10540 8121
rect 10484 8067 10486 8119
rect 10486 8067 10538 8119
rect 10538 8067 10540 8119
rect 10484 8065 10540 8067
rect 8980 7831 9036 7833
rect 8980 7779 8982 7831
rect 8982 7779 9034 7831
rect 9034 7779 9036 7831
rect 8980 7777 9036 7779
rect 8980 7727 9036 7729
rect 8980 7675 8982 7727
rect 8982 7675 9034 7727
rect 9034 7675 9036 7727
rect 8980 7673 9036 7675
rect 9876 7831 9932 7833
rect 9876 7779 9878 7831
rect 9878 7779 9930 7831
rect 9930 7779 9932 7831
rect 9876 7777 9932 7779
rect 9876 7727 9932 7729
rect 9876 7675 9878 7727
rect 9878 7675 9930 7727
rect 9930 7675 9932 7727
rect 9876 7673 9932 7675
rect 10772 7831 10828 7833
rect 10772 7779 10774 7831
rect 10774 7779 10826 7831
rect 10826 7779 10828 7831
rect 10772 7777 10828 7779
rect 10772 7727 10828 7729
rect 10772 7675 10774 7727
rect 10774 7675 10826 7727
rect 10826 7675 10828 7727
rect 10772 7673 10828 7675
rect 7392 6355 7448 6411
rect 7496 6355 7552 6411
rect 7392 6251 7448 6307
rect 7496 6251 7552 6307
rect 8285 6409 8341 6411
rect 8285 6357 8287 6409
rect 8287 6357 8339 6409
rect 8339 6357 8341 6409
rect 8285 6355 8341 6357
rect 8389 6409 8445 6411
rect 8389 6357 8391 6409
rect 8391 6357 8443 6409
rect 8443 6357 8445 6409
rect 8389 6355 8445 6357
rect 8285 6305 8341 6307
rect 8285 6253 8287 6305
rect 8287 6253 8339 6305
rect 8339 6253 8341 6305
rect 8285 6251 8341 6253
rect 8389 6305 8445 6307
rect 8389 6253 8391 6305
rect 8391 6253 8443 6305
rect 8443 6253 8445 6305
rect 8389 6251 8445 6253
rect 3057 5173 3113 5175
rect 3057 5121 3059 5173
rect 3059 5121 3111 5173
rect 3111 5121 3113 5173
rect 3057 5119 3113 5121
rect 3161 5173 3217 5175
rect 3161 5121 3163 5173
rect 3163 5121 3215 5173
rect 3215 5121 3217 5173
rect 3161 5119 3217 5121
rect 3057 5069 3113 5071
rect 3057 5017 3059 5069
rect 3059 5017 3111 5069
rect 3111 5017 3113 5069
rect 3057 5015 3113 5017
rect 3161 5069 3217 5071
rect 3161 5017 3163 5069
rect 3163 5017 3215 5069
rect 3215 5017 3217 5069
rect 3161 5015 3217 5017
rect 2725 4419 2781 4421
rect 2725 4367 2727 4419
rect 2727 4367 2779 4419
rect 2779 4367 2781 4419
rect 2725 4365 2781 4367
rect 2725 4315 2781 4317
rect 2725 4263 2727 4315
rect 2727 4263 2779 4315
rect 2779 4263 2781 4315
rect 2725 4261 2781 4263
rect 4021 4129 4077 4131
rect 4021 4077 4023 4129
rect 4023 4077 4075 4129
rect 4075 4077 4077 4129
rect 4021 4075 4077 4077
rect 4021 4025 4077 4027
rect 4021 3973 4023 4025
rect 4023 3973 4075 4025
rect 4075 3973 4077 4025
rect 4021 3971 4077 3973
rect 3589 3805 3645 3807
rect 3589 3753 3591 3805
rect 3591 3753 3643 3805
rect 3643 3753 3645 3805
rect 3589 3751 3645 3753
rect 3589 3701 3645 3703
rect 3589 3649 3591 3701
rect 3591 3649 3643 3701
rect 3643 3649 3645 3701
rect 3589 3647 3645 3649
rect 3429 3349 3485 3405
rect 3533 3349 3589 3405
rect 3429 3245 3485 3301
rect 3533 3245 3589 3301
rect 1237 3105 1293 3161
rect 1341 3105 1397 3161
rect 1237 3001 1293 3057
rect 1341 3001 1397 3057
rect 2735 3159 2791 3161
rect 2735 3107 2737 3159
rect 2737 3107 2789 3159
rect 2789 3107 2791 3159
rect 2735 3105 2791 3107
rect 2735 3055 2791 3057
rect 2735 3003 2737 3055
rect 2737 3003 2789 3055
rect 2789 3003 2791 3055
rect 2735 3001 2791 3003
rect 5630 4365 5686 4421
rect 5734 4365 5790 4421
rect 5630 4261 5686 4317
rect 5734 4261 5790 4317
rect 5394 3751 5450 3807
rect 5498 3751 5554 3807
rect 5394 3647 5450 3703
rect 5498 3647 5554 3703
rect 3933 2543 3989 2545
rect 3933 2491 3935 2543
rect 3935 2491 3987 2543
rect 3987 2491 3989 2543
rect 3933 2489 3989 2491
rect 3933 2439 3989 2441
rect 3933 2387 3935 2439
rect 3935 2387 3987 2439
rect 3987 2387 3989 2439
rect 3933 2385 3989 2387
rect 5154 2489 5210 2545
rect 5258 2489 5314 2545
rect 5154 2385 5210 2441
rect 5258 2385 5314 2441
rect -8163 2047 -8107 2103
rect -8053 2047 -7997 2103
rect 5394 2346 5450 2402
rect 5498 2346 5554 2402
rect 5394 2242 5450 2298
rect 5498 2242 5554 2298
rect -8163 1937 -8107 1993
rect -8053 1937 -7997 1993
rect 5154 1960 5210 2016
rect 5258 1960 5314 2016
rect 5154 1856 5210 1912
rect 5258 1856 5314 1912
rect 3981 1773 4037 1775
rect 3981 1721 3983 1773
rect 3983 1721 4035 1773
rect 4035 1721 4037 1773
rect 3981 1719 4037 1721
rect 3981 1669 4037 1671
rect 3981 1617 3983 1669
rect 3983 1617 4035 1669
rect 4035 1617 4037 1669
rect 3981 1615 4037 1617
rect 6103 4075 6159 4131
rect 6207 4075 6263 4131
rect 6103 3971 6159 4027
rect 6207 3971 6263 4027
rect 6554 4101 6610 4103
rect 6554 4049 6556 4101
rect 6556 4049 6608 4101
rect 6608 4049 6610 4101
rect 6554 4047 6610 4049
rect 6658 4101 6714 4103
rect 6658 4049 6660 4101
rect 6660 4049 6712 4101
rect 6712 4049 6714 4101
rect 6658 4047 6714 4049
rect 5861 3557 5917 3613
rect 5965 3557 6021 3613
rect 5861 3453 5917 3509
rect 5965 3453 6021 3509
rect 5861 3349 5917 3405
rect 5965 3349 6021 3405
rect 5861 3245 5917 3301
rect 5965 3245 6021 3301
rect 6554 3997 6610 3999
rect 6554 3945 6556 3997
rect 6556 3945 6608 3997
rect 6608 3945 6610 3997
rect 6554 3943 6610 3945
rect 6658 3997 6714 3999
rect 6658 3945 6660 3997
rect 6660 3945 6712 3997
rect 6712 3945 6714 3997
rect 6658 3943 6714 3945
rect 6864 4047 6920 4103
rect 6968 4047 7024 4103
rect 6864 3943 6920 3999
rect 6968 3943 7024 3999
rect 6103 2833 6159 2889
rect 6207 2833 6263 2889
rect 6103 2729 6159 2785
rect 6207 2729 6263 2785
rect 6592 2400 6648 2402
rect 6592 2348 6594 2400
rect 6594 2348 6646 2400
rect 6646 2348 6648 2400
rect 6592 2346 6648 2348
rect 6592 2296 6648 2298
rect 6592 2244 6594 2296
rect 6594 2244 6646 2296
rect 6646 2244 6648 2296
rect 6592 2242 6648 2244
rect 6522 1960 6578 2016
rect 6626 1960 6682 2016
rect 6522 1910 6578 1912
rect 6522 1858 6524 1910
rect 6524 1858 6576 1910
rect 6576 1858 6578 1910
rect 6522 1856 6578 1858
rect 6626 1910 6682 1912
rect 6626 1858 6628 1910
rect 6628 1858 6680 1910
rect 6680 1858 6682 1910
rect 6626 1856 6682 1858
rect 7128 2833 7184 2889
rect 7232 2833 7288 2889
rect 7128 2729 7184 2785
rect 7232 2729 7288 2785
rect 9199 5988 9255 6044
rect 9199 5938 9255 5940
rect 9199 5886 9201 5938
rect 9201 5886 9253 5938
rect 9253 5886 9255 5938
rect 9199 5884 9255 5886
rect 10288 6042 10344 6044
rect 10288 5990 10290 6042
rect 10290 5990 10342 6042
rect 10342 5990 10344 6042
rect 10288 5988 10344 5990
rect 10392 6042 10448 6044
rect 10392 5990 10394 6042
rect 10394 5990 10446 6042
rect 10446 5990 10448 6042
rect 10392 5988 10448 5990
rect 10288 5938 10344 5940
rect 10288 5886 10290 5938
rect 10290 5886 10342 5938
rect 10342 5886 10344 5938
rect 10288 5884 10344 5886
rect 10392 5938 10448 5940
rect 10392 5886 10394 5938
rect 10394 5886 10446 5938
rect 10446 5886 10448 5938
rect 10392 5884 10448 5886
rect 7839 5709 7895 5711
rect 7839 5657 7841 5709
rect 7841 5657 7893 5709
rect 7893 5657 7895 5709
rect 7839 5655 7895 5657
rect 7839 5605 7895 5607
rect 7839 5553 7841 5605
rect 7841 5553 7893 5605
rect 7893 5553 7895 5605
rect 7839 5551 7895 5553
rect 8159 5709 8215 5711
rect 8159 5657 8161 5709
rect 8161 5657 8213 5709
rect 8213 5657 8215 5709
rect 8159 5655 8215 5657
rect 8159 5605 8215 5607
rect 8159 5553 8161 5605
rect 8161 5553 8213 5605
rect 8213 5553 8215 5605
rect 8159 5551 8215 5553
rect 8479 5709 8535 5711
rect 8479 5657 8481 5709
rect 8481 5657 8533 5709
rect 8533 5657 8535 5709
rect 8479 5655 8535 5657
rect 8479 5605 8535 5607
rect 8479 5553 8481 5605
rect 8481 5553 8533 5605
rect 8533 5553 8535 5605
rect 8479 5551 8535 5553
rect 8799 5709 8855 5711
rect 8799 5657 8801 5709
rect 8801 5657 8853 5709
rect 8853 5657 8855 5709
rect 8799 5655 8855 5657
rect 8799 5605 8855 5607
rect 8799 5553 8801 5605
rect 8801 5553 8853 5605
rect 8853 5553 8855 5605
rect 8799 5551 8855 5553
rect 8959 5709 9015 5711
rect 8959 5657 8961 5709
rect 8961 5657 9013 5709
rect 9013 5657 9015 5709
rect 8959 5655 9015 5657
rect 8959 5605 9015 5607
rect 8959 5553 8961 5605
rect 8961 5553 9013 5605
rect 9013 5553 9015 5605
rect 8959 5551 9015 5553
rect 7999 5173 8055 5175
rect 7999 5121 8001 5173
rect 8001 5121 8053 5173
rect 8053 5121 8055 5173
rect 7999 5119 8055 5121
rect 7999 5069 8055 5071
rect 7999 5017 8001 5069
rect 8001 5017 8053 5069
rect 8053 5017 8055 5069
rect 7999 5015 8055 5017
rect 8159 5173 8215 5175
rect 8159 5121 8161 5173
rect 8161 5121 8213 5173
rect 8213 5121 8215 5173
rect 8159 5119 8215 5121
rect 8159 5069 8215 5071
rect 8159 5017 8161 5069
rect 8161 5017 8213 5069
rect 8213 5017 8215 5069
rect 8159 5015 8215 5017
rect 8479 5173 8535 5175
rect 8479 5121 8481 5173
rect 8481 5121 8533 5173
rect 8533 5121 8535 5173
rect 8479 5119 8535 5121
rect 8479 5069 8535 5071
rect 8479 5017 8481 5069
rect 8481 5017 8533 5069
rect 8533 5017 8535 5069
rect 8479 5015 8535 5017
rect 8799 5173 8855 5175
rect 8799 5121 8801 5173
rect 8801 5121 8853 5173
rect 8853 5121 8855 5173
rect 8799 5119 8855 5121
rect 8799 5069 8855 5071
rect 8799 5017 8801 5069
rect 8801 5017 8853 5069
rect 8853 5017 8855 5069
rect 8799 5015 8855 5017
rect 7839 4637 7895 4639
rect 7839 4585 7841 4637
rect 7841 4585 7893 4637
rect 7893 4585 7895 4637
rect 7839 4583 7895 4585
rect 7839 4533 7895 4535
rect 7839 4481 7841 4533
rect 7841 4481 7893 4533
rect 7893 4481 7895 4533
rect 7839 4479 7895 4481
rect 9278 5402 9334 5404
rect 9278 5350 9280 5402
rect 9280 5350 9332 5402
rect 9332 5350 9334 5402
rect 9278 5348 9334 5350
rect 9119 5173 9175 5175
rect 9119 5121 9121 5173
rect 9121 5121 9173 5173
rect 9173 5121 9175 5173
rect 9119 5119 9175 5121
rect 9119 5069 9175 5071
rect 9119 5017 9121 5069
rect 9121 5017 9173 5069
rect 9173 5017 9175 5069
rect 9119 5015 9175 5017
rect 10554 5444 10610 5446
rect 10554 5392 10556 5444
rect 10556 5392 10608 5444
rect 10608 5392 10610 5444
rect 10554 5390 10610 5392
rect 10658 5444 10714 5446
rect 10658 5392 10660 5444
rect 10660 5392 10712 5444
rect 10712 5392 10714 5444
rect 10658 5390 10714 5392
rect 10554 5340 10610 5342
rect 10554 5288 10556 5340
rect 10556 5288 10608 5340
rect 10608 5288 10610 5340
rect 10554 5286 10610 5288
rect 10658 5340 10714 5342
rect 10658 5288 10660 5340
rect 10660 5288 10712 5340
rect 10712 5288 10714 5340
rect 10658 5286 10714 5288
rect 9081 4866 9137 4868
rect 9081 4814 9083 4866
rect 9083 4814 9135 4866
rect 9135 4814 9137 4866
rect 9081 4812 9137 4814
rect 10288 4864 10344 4920
rect 10392 4864 10448 4920
rect 10288 4760 10344 4816
rect 10392 4760 10448 4816
rect 8159 4637 8215 4639
rect 8159 4585 8161 4637
rect 8161 4585 8213 4637
rect 8213 4585 8215 4637
rect 8159 4583 8215 4585
rect 8159 4533 8215 4535
rect 8159 4481 8161 4533
rect 8161 4481 8213 4533
rect 8213 4481 8215 4533
rect 8159 4479 8215 4481
rect 8479 4637 8535 4639
rect 8479 4585 8481 4637
rect 8481 4585 8533 4637
rect 8533 4585 8535 4637
rect 8479 4583 8535 4585
rect 8479 4533 8535 4535
rect 8479 4481 8481 4533
rect 8481 4481 8533 4533
rect 8533 4481 8535 4533
rect 8479 4479 8535 4481
rect 8799 4637 8855 4639
rect 8799 4585 8801 4637
rect 8801 4585 8853 4637
rect 8853 4585 8855 4637
rect 8799 4583 8855 4585
rect 8799 4533 8855 4535
rect 8799 4481 8801 4533
rect 8801 4481 8853 4533
rect 8853 4481 8855 4533
rect 8799 4479 8855 4481
rect 9119 4637 9175 4639
rect 9119 4585 9121 4637
rect 9121 4585 9173 4637
rect 9173 4585 9175 4637
rect 9119 4583 9175 4585
rect 9119 4533 9175 4535
rect 9119 4481 9121 4533
rect 9121 4481 9173 4533
rect 9173 4481 9175 4533
rect 9119 4479 9175 4481
rect 7839 4101 7895 4103
rect 7839 4049 7841 4101
rect 7841 4049 7893 4101
rect 7893 4049 7895 4101
rect 7839 4047 7895 4049
rect 7839 3997 7895 3999
rect 7839 3945 7841 3997
rect 7841 3945 7893 3997
rect 7893 3945 7895 3997
rect 7839 3943 7895 3945
rect 8159 4101 8215 4103
rect 8159 4049 8161 4101
rect 8161 4049 8213 4101
rect 8213 4049 8215 4101
rect 8159 4047 8215 4049
rect 8159 3997 8215 3999
rect 8159 3945 8161 3997
rect 8161 3945 8213 3997
rect 8213 3945 8215 3997
rect 8159 3943 8215 3945
rect 8479 4101 8535 4103
rect 8479 4049 8481 4101
rect 8481 4049 8533 4101
rect 8533 4049 8535 4101
rect 8479 4047 8535 4049
rect 8479 3997 8535 3999
rect 8479 3945 8481 3997
rect 8481 3945 8533 3997
rect 8533 3945 8535 3997
rect 8479 3943 8535 3945
rect 8799 4101 8855 4103
rect 8799 4049 8801 4101
rect 8801 4049 8853 4101
rect 8853 4049 8855 4101
rect 8799 4047 8855 4049
rect 8799 3997 8855 3999
rect 8799 3945 8801 3997
rect 8801 3945 8853 3997
rect 8853 3945 8855 3997
rect 8799 3943 8855 3945
rect 9199 4332 9255 4334
rect 9199 4280 9201 4332
rect 9201 4280 9253 4332
rect 9253 4280 9255 4332
rect 9199 4278 9255 4280
rect 9119 4101 9175 4103
rect 9119 4049 9121 4101
rect 9121 4049 9173 4101
rect 9173 4049 9175 4101
rect 9119 4047 9175 4049
rect 9119 3997 9175 3999
rect 9119 3945 9121 3997
rect 9121 3945 9173 3997
rect 9173 3945 9175 3997
rect 9119 3943 9175 3945
rect 9278 3846 9334 3902
rect 9278 3796 9334 3798
rect 9278 3744 9280 3796
rect 9280 3744 9332 3796
rect 9332 3744 9334 3796
rect 9278 3742 9334 3744
rect 10554 4330 10610 4386
rect 10658 4330 10714 4386
rect 10554 4226 10610 4282
rect 10658 4226 10714 4282
rect 10016 3846 10072 3902
rect 10120 3846 10176 3902
rect 10016 3742 10072 3798
rect 10120 3742 10176 3798
rect 10288 3844 10344 3900
rect 10392 3844 10448 3900
rect 10288 3740 10344 3796
rect 10392 3740 10448 3796
rect 8959 3565 9015 3567
rect 8959 3513 8961 3565
rect 8961 3513 9013 3565
rect 9013 3513 9015 3565
rect 8959 3511 9015 3513
rect 8959 3461 9015 3463
rect 8959 3409 8961 3461
rect 8961 3409 9013 3461
rect 9013 3409 9015 3461
rect 8959 3407 9015 3409
rect 9278 3331 9334 3387
rect 9278 3281 9334 3283
rect 9278 3229 9280 3281
rect 9280 3229 9332 3281
rect 9332 3229 9334 3281
rect 9278 3227 9334 3229
rect 9749 3105 9805 3161
rect 9853 3105 9909 3161
rect 9749 3001 9805 3057
rect 9853 3001 9909 3057
rect 8879 2709 8935 2711
rect 8879 2657 8881 2709
rect 8881 2657 8933 2709
rect 8933 2657 8935 2709
rect 8879 2655 8935 2657
rect 8879 2551 8935 2607
rect 10554 3331 10610 3387
rect 10658 3331 10714 3387
rect 10554 3227 10610 3283
rect 10658 3227 10714 3283
rect 10016 2655 10072 2711
rect 10120 2655 10176 2711
rect 10016 2551 10072 2607
rect 10120 2551 10176 2607
rect 7128 1950 7184 2006
rect 7232 1950 7288 2006
rect 7128 1846 7184 1902
rect 7232 1846 7288 1902
rect 9406 2004 9462 2006
rect 9406 1952 9408 2004
rect 9408 1952 9460 2004
rect 9460 1952 9462 2004
rect 9406 1950 9462 1952
rect 9510 2004 9566 2006
rect 9510 1952 9512 2004
rect 9512 1952 9564 2004
rect 9564 1952 9566 2004
rect 9510 1950 9566 1952
rect 9406 1900 9462 1902
rect 9406 1848 9408 1900
rect 9408 1848 9460 1900
rect 9460 1848 9462 1900
rect 9406 1846 9462 1848
rect 9510 1900 9566 1902
rect 9510 1848 9512 1900
rect 9512 1848 9564 1900
rect 9564 1848 9566 1900
rect 9510 1846 9566 1848
rect 6432 1771 6488 1773
rect 6432 1719 6434 1771
rect 6434 1719 6486 1771
rect 6486 1719 6488 1771
rect 6432 1717 6488 1719
rect 6432 1667 6488 1669
rect 6432 1615 6434 1667
rect 6434 1615 6486 1667
rect 6486 1615 6488 1667
rect 6432 1613 6488 1615
rect 6864 1765 6920 1767
rect 6864 1713 6866 1765
rect 6866 1713 6918 1765
rect 6918 1713 6920 1765
rect 6864 1711 6920 1713
rect 6968 1711 7024 1767
rect 6864 1661 6920 1663
rect 6864 1609 6866 1661
rect 6866 1609 6918 1661
rect 6918 1609 6920 1661
rect 6864 1607 6920 1609
rect 6968 1607 7024 1663
rect 6380 1073 6436 1129
rect 6484 1073 6540 1129
rect 6380 969 6436 1025
rect 6484 969 6540 1025
rect 13994 10189 14050 10191
rect 13994 10137 13996 10189
rect 13996 10137 14048 10189
rect 14048 10137 14050 10189
rect 13994 10135 14050 10137
rect 15156 10293 15212 10295
rect 15156 10241 15158 10293
rect 15158 10241 15210 10293
rect 15210 10241 15212 10293
rect 15156 10239 15212 10241
rect 15156 10189 15212 10191
rect 15156 10137 15158 10189
rect 15158 10137 15210 10189
rect 15210 10137 15212 10189
rect 15156 10135 15212 10137
rect 15796 10293 15852 10295
rect 15796 10241 15798 10293
rect 15798 10241 15850 10293
rect 15850 10241 15852 10293
rect 15796 10239 15852 10241
rect 15796 10189 15852 10191
rect 15796 10137 15798 10189
rect 15798 10137 15850 10189
rect 15850 10137 15852 10189
rect 15796 10135 15852 10137
rect 16436 10293 16492 10295
rect 16436 10241 16438 10293
rect 16438 10241 16490 10293
rect 16490 10241 16492 10293
rect 16436 10239 16492 10241
rect 16436 10189 16492 10191
rect 16436 10137 16438 10189
rect 16438 10137 16490 10189
rect 16490 10137 16492 10189
rect 16436 10135 16492 10137
rect 17113 10239 17169 10295
rect 17217 10239 17273 10295
rect 17113 10135 17169 10191
rect 17217 10135 17273 10191
rect 12362 9273 12418 9275
rect 12362 9221 12364 9273
rect 12364 9221 12416 9273
rect 12416 9221 12418 9273
rect 12362 9219 12418 9221
rect 12362 9169 12418 9171
rect 12362 9117 12364 9169
rect 12364 9117 12416 9169
rect 12416 9117 12418 9169
rect 12362 9115 12418 9117
rect 13258 9273 13314 9275
rect 13258 9221 13260 9273
rect 13260 9221 13312 9273
rect 13312 9221 13314 9273
rect 13258 9219 13314 9221
rect 13258 9169 13314 9171
rect 13258 9117 13260 9169
rect 13260 9117 13312 9169
rect 13312 9117 13314 9169
rect 13258 9115 13314 9117
rect 14154 9273 14210 9275
rect 14154 9221 14156 9273
rect 14156 9221 14208 9273
rect 14208 9221 14210 9273
rect 14154 9219 14210 9221
rect 14154 9169 14210 9171
rect 14154 9117 14156 9169
rect 14156 9117 14208 9169
rect 14208 9117 14210 9169
rect 14154 9115 14210 9117
rect 13866 8873 13922 8875
rect 13866 8821 13868 8873
rect 13868 8821 13920 8873
rect 13920 8821 13922 8873
rect 13866 8819 13922 8821
rect 13866 8769 13922 8771
rect 13866 8717 13868 8769
rect 13868 8717 13920 8769
rect 13920 8717 13922 8769
rect 13866 8715 13922 8717
rect 15476 8873 15532 8875
rect 15476 8821 15478 8873
rect 15478 8821 15530 8873
rect 15530 8821 15532 8873
rect 15476 8819 15532 8821
rect 15476 8769 15532 8771
rect 15476 8717 15478 8769
rect 15478 8717 15530 8769
rect 15530 8717 15532 8769
rect 15476 8715 15532 8717
rect 16116 8873 16172 8875
rect 16116 8821 16118 8873
rect 16118 8821 16170 8873
rect 16170 8821 16172 8873
rect 16116 8819 16172 8821
rect 16116 8769 16172 8771
rect 16116 8717 16118 8769
rect 16118 8717 16170 8769
rect 16170 8717 16172 8769
rect 16116 8715 16172 8717
rect 11649 8649 11705 8705
rect 11753 8649 11809 8705
rect 11649 8545 11705 8601
rect 11753 8545 11809 8601
rect 11381 8169 11437 8225
rect 11485 8169 11541 8225
rect 11381 8065 11437 8121
rect 11485 8065 11541 8121
rect 12028 8509 12084 8565
rect 12132 8509 12188 8565
rect 12028 8405 12084 8461
rect 12132 8405 12188 8461
rect 12398 8563 12454 8565
rect 12398 8511 12400 8563
rect 12400 8511 12452 8563
rect 12452 8511 12454 8563
rect 12398 8509 12454 8511
rect 12398 8459 12454 8461
rect 12398 8407 12400 8459
rect 12400 8407 12452 8459
rect 12452 8407 12454 8459
rect 12398 8405 12454 8407
rect 14696 8514 14752 8570
rect 14800 8514 14856 8570
rect 14696 8410 14752 8466
rect 14800 8410 14856 8466
rect 15184 8568 15240 8570
rect 15184 8516 15186 8568
rect 15186 8516 15238 8568
rect 15238 8516 15240 8568
rect 15184 8514 15240 8516
rect 15184 8464 15240 8466
rect 15184 8412 15186 8464
rect 15186 8412 15238 8464
rect 15238 8412 15240 8464
rect 15184 8410 15240 8412
rect 11649 7769 11705 7825
rect 11753 7769 11809 7825
rect 11649 7665 11705 7721
rect 11753 7665 11809 7721
rect 10928 1950 10984 2006
rect 11032 1950 11088 2006
rect 10928 1846 10984 1902
rect 11032 1846 11088 1902
rect 11315 2004 11371 2006
rect 11315 1952 11317 2004
rect 11317 1952 11369 2004
rect 11369 1952 11371 2004
rect 11315 1950 11371 1952
rect 11419 2004 11475 2006
rect 11419 1952 11421 2004
rect 11421 1952 11473 2004
rect 11473 1952 11475 2004
rect 11419 1950 11475 1952
rect 11315 1900 11371 1902
rect 11315 1848 11317 1900
rect 11317 1848 11369 1900
rect 11369 1848 11371 1900
rect 11315 1846 11371 1848
rect 11419 1900 11475 1902
rect 11419 1848 11421 1900
rect 11421 1848 11473 1900
rect 11473 1848 11475 1900
rect 11419 1846 11475 1848
rect 12810 8223 12866 8225
rect 12810 8171 12812 8223
rect 12812 8171 12864 8223
rect 12864 8171 12866 8223
rect 12810 8169 12866 8171
rect 12810 8119 12866 8121
rect 12810 8067 12812 8119
rect 12812 8067 12864 8119
rect 12864 8067 12866 8119
rect 12810 8065 12866 8067
rect 13706 8223 13762 8225
rect 13706 8171 13708 8223
rect 13708 8171 13760 8223
rect 13760 8171 13762 8223
rect 13706 8169 13762 8171
rect 13706 8119 13762 8121
rect 13706 8067 13708 8119
rect 13708 8067 13760 8119
rect 13760 8067 13762 8119
rect 13706 8065 13762 8067
rect 13866 8223 13922 8225
rect 13866 8171 13868 8223
rect 13868 8171 13920 8223
rect 13920 8171 13922 8223
rect 13866 8169 13922 8171
rect 13866 8119 13922 8121
rect 13866 8067 13868 8119
rect 13868 8067 13920 8119
rect 13920 8067 13922 8119
rect 13866 8065 13922 8067
rect 12362 7823 12418 7825
rect 12362 7771 12364 7823
rect 12364 7771 12416 7823
rect 12416 7771 12418 7823
rect 12362 7769 12418 7771
rect 12362 7719 12418 7721
rect 12362 7667 12364 7719
rect 12364 7667 12416 7719
rect 12416 7667 12418 7719
rect 12362 7665 12418 7667
rect 13258 7823 13314 7825
rect 13258 7771 13260 7823
rect 13260 7771 13312 7823
rect 13312 7771 13314 7823
rect 13258 7769 13314 7771
rect 13258 7719 13314 7721
rect 13258 7667 13260 7719
rect 13260 7667 13312 7719
rect 13312 7667 13314 7719
rect 13258 7665 13314 7667
rect 14154 7823 14210 7825
rect 14154 7771 14156 7823
rect 14156 7771 14208 7823
rect 14208 7771 14210 7823
rect 14154 7769 14210 7771
rect 14154 7719 14210 7721
rect 14154 7667 14156 7719
rect 14156 7667 14208 7719
rect 14208 7667 14210 7719
rect 14154 7665 14210 7667
rect 17375 8819 17431 8875
rect 17479 8819 17535 8875
rect 17375 8715 17431 8771
rect 17479 8715 17535 8771
rect 15476 8223 15532 8225
rect 15476 8171 15478 8223
rect 15478 8171 15530 8223
rect 15530 8171 15532 8223
rect 15476 8169 15532 8171
rect 15476 8119 15532 8121
rect 15476 8067 15478 8119
rect 15478 8067 15530 8119
rect 15530 8067 15532 8119
rect 15476 8065 15532 8067
rect 16116 8223 16172 8225
rect 16116 8171 16118 8223
rect 16118 8171 16170 8223
rect 16170 8171 16172 8223
rect 16116 8169 16172 8171
rect 16116 8119 16172 8121
rect 16116 8067 16118 8119
rect 16118 8067 16170 8119
rect 16170 8067 16172 8119
rect 16116 8065 16172 8067
rect 17113 8169 17169 8225
rect 17217 8169 17273 8225
rect 17113 8065 17169 8121
rect 17217 8065 17273 8121
rect 17651 8641 17707 8697
rect 17851 12385 17907 12441
rect 19075 12439 19131 12441
rect 19075 12387 19077 12439
rect 19077 12387 19129 12439
rect 19129 12387 19131 12439
rect 19075 12385 19131 12387
rect 19315 12228 19371 12230
rect 19315 12176 19317 12228
rect 19317 12176 19369 12228
rect 19369 12176 19371 12228
rect 19315 12174 19371 12176
rect 19315 12124 19371 12126
rect 19315 12072 19317 12124
rect 19317 12072 19369 12124
rect 19369 12072 19371 12124
rect 19315 12070 19371 12072
rect 19955 12228 20011 12230
rect 19955 12176 19957 12228
rect 19957 12176 20009 12228
rect 20009 12176 20011 12228
rect 19955 12174 20011 12176
rect 19955 12124 20011 12126
rect 19955 12072 19957 12124
rect 19957 12072 20009 12124
rect 20009 12072 20011 12124
rect 19955 12070 20011 12072
rect 21458 12278 21514 12334
rect 21562 12278 21618 12334
rect 21666 12278 21722 12334
rect 21458 12174 21514 12230
rect 21562 12174 21618 12230
rect 21666 12174 21722 12230
rect 21458 12070 21514 12126
rect 21562 12070 21618 12126
rect 21666 12070 21722 12126
rect 18995 11834 19051 11836
rect 18995 11782 18997 11834
rect 18997 11782 19049 11834
rect 19049 11782 19051 11834
rect 18995 11780 19051 11782
rect 18995 11730 19051 11732
rect 18995 11678 18997 11730
rect 18997 11678 19049 11730
rect 19049 11678 19051 11730
rect 18995 11676 19051 11678
rect 19635 11834 19691 11836
rect 19635 11782 19637 11834
rect 19637 11782 19689 11834
rect 19689 11782 19691 11834
rect 19635 11780 19691 11782
rect 19635 11730 19691 11732
rect 19635 11678 19637 11730
rect 19637 11678 19689 11730
rect 19689 11678 19691 11730
rect 19635 11676 19691 11678
rect 20275 11834 20331 11836
rect 20275 11782 20277 11834
rect 20277 11782 20329 11834
rect 20329 11782 20331 11834
rect 20275 11780 20331 11782
rect 20275 11730 20331 11732
rect 20275 11678 20277 11730
rect 20277 11678 20329 11730
rect 20329 11678 20331 11730
rect 20275 11676 20331 11678
rect 19075 11503 19131 11505
rect 19075 11451 19077 11503
rect 19077 11451 19129 11503
rect 19129 11451 19131 11503
rect 19075 11449 19131 11451
rect 19315 11292 19371 11294
rect 19315 11240 19317 11292
rect 19317 11240 19369 11292
rect 19369 11240 19371 11292
rect 19315 11238 19371 11240
rect 19315 11188 19371 11190
rect 19315 11136 19317 11188
rect 19317 11136 19369 11188
rect 19369 11136 19371 11188
rect 19315 11134 19371 11136
rect 19955 11292 20011 11294
rect 19955 11240 19957 11292
rect 19957 11240 20009 11292
rect 20009 11240 20011 11292
rect 19955 11238 20011 11240
rect 19955 11188 20011 11190
rect 19955 11136 19957 11188
rect 19957 11136 20009 11188
rect 20009 11136 20011 11188
rect 19955 11134 20011 11136
rect 21458 10948 21514 11004
rect 21562 10948 21618 11004
rect 21666 10948 21722 11004
rect 18995 10898 19051 10900
rect 18995 10846 18997 10898
rect 18997 10846 19049 10898
rect 19049 10846 19051 10898
rect 18995 10844 19051 10846
rect 18995 10794 19051 10796
rect 18995 10742 18997 10794
rect 18997 10742 19049 10794
rect 19049 10742 19051 10794
rect 18995 10740 19051 10742
rect 19635 10898 19691 10900
rect 19635 10846 19637 10898
rect 19637 10846 19689 10898
rect 19689 10846 19691 10898
rect 19635 10844 19691 10846
rect 19635 10794 19691 10796
rect 19635 10742 19637 10794
rect 19637 10742 19689 10794
rect 19689 10742 19691 10794
rect 19635 10740 19691 10742
rect 20275 10898 20331 10900
rect 20275 10846 20277 10898
rect 20277 10846 20329 10898
rect 20329 10846 20331 10898
rect 20275 10844 20331 10846
rect 20275 10794 20331 10796
rect 20275 10742 20277 10794
rect 20277 10742 20329 10794
rect 20329 10742 20331 10794
rect 20275 10740 20331 10742
rect 21458 10844 21514 10900
rect 21562 10844 21618 10900
rect 21666 10844 21722 10900
rect 21458 10740 21514 10796
rect 21562 10740 21618 10796
rect 21666 10740 21722 10796
rect 19315 10356 19371 10358
rect 19315 10304 19317 10356
rect 19317 10304 19369 10356
rect 19369 10304 19371 10356
rect 19315 10302 19371 10304
rect 19315 10252 19371 10254
rect 19315 10200 19317 10252
rect 19317 10200 19369 10252
rect 19369 10200 19371 10252
rect 19315 10198 19371 10200
rect 18995 9962 19051 9964
rect 18995 9910 18997 9962
rect 18997 9910 19049 9962
rect 19049 9910 19051 9962
rect 18995 9908 19051 9910
rect 18995 9858 19051 9860
rect 18995 9806 18997 9858
rect 18997 9806 19049 9858
rect 19049 9806 19051 9858
rect 18995 9804 19051 9806
rect 17851 9577 17907 9633
rect 15156 7833 15212 7835
rect 15156 7781 15158 7833
rect 15158 7781 15210 7833
rect 15210 7781 15212 7833
rect 15156 7779 15212 7781
rect 15156 7729 15212 7731
rect 15156 7677 15158 7729
rect 15158 7677 15210 7729
rect 15210 7677 15212 7729
rect 15156 7675 15212 7677
rect 15796 7833 15852 7835
rect 15796 7781 15798 7833
rect 15798 7781 15850 7833
rect 15850 7781 15852 7833
rect 15796 7779 15852 7781
rect 15796 7729 15852 7731
rect 15796 7677 15798 7729
rect 15798 7677 15850 7729
rect 15850 7677 15852 7729
rect 15796 7675 15852 7677
rect 16436 7833 16492 7835
rect 16436 7781 16438 7833
rect 16438 7781 16490 7833
rect 16490 7781 16492 7833
rect 16436 7779 16492 7781
rect 16436 7729 16492 7731
rect 16436 7677 16438 7729
rect 16438 7677 16490 7729
rect 16490 7677 16492 7729
rect 16436 7675 16492 7677
rect 17375 7779 17431 7835
rect 17479 7779 17535 7835
rect 17375 7675 17431 7731
rect 17479 7675 17535 7731
rect 19075 9631 19131 9633
rect 19075 9579 19077 9631
rect 19077 9579 19129 9631
rect 19129 9579 19131 9631
rect 19075 9577 19131 9579
rect 19315 9420 19371 9422
rect 19315 9368 19317 9420
rect 19317 9368 19369 9420
rect 19369 9368 19371 9420
rect 19315 9366 19371 9368
rect 19315 9316 19371 9318
rect 19315 9264 19317 9316
rect 19317 9264 19369 9316
rect 19369 9264 19371 9316
rect 19315 9262 19371 9264
rect 19635 9962 19691 9964
rect 19635 9910 19637 9962
rect 19637 9910 19689 9962
rect 19689 9910 19691 9962
rect 19635 9908 19691 9910
rect 19635 9858 19691 9860
rect 19635 9806 19637 9858
rect 19637 9806 19689 9858
rect 19689 9806 19691 9858
rect 19635 9804 19691 9806
rect 19955 10356 20011 10358
rect 19955 10304 19957 10356
rect 19957 10304 20009 10356
rect 20009 10304 20011 10356
rect 19955 10302 20011 10304
rect 19955 10252 20011 10254
rect 19955 10200 19957 10252
rect 19957 10200 20009 10252
rect 20009 10200 20011 10252
rect 19955 10198 20011 10200
rect 19955 9420 20011 9422
rect 19955 9368 19957 9420
rect 19957 9368 20009 9420
rect 20009 9368 20011 9420
rect 19955 9366 20011 9368
rect 19955 9316 20011 9318
rect 19955 9264 19957 9316
rect 19957 9264 20009 9316
rect 20009 9264 20011 9316
rect 19955 9262 20011 9264
rect 21458 10012 21514 10068
rect 21562 10012 21618 10068
rect 21666 10012 21722 10068
rect 20275 9962 20331 9964
rect 20275 9910 20277 9962
rect 20277 9910 20329 9962
rect 20329 9910 20331 9962
rect 20275 9908 20331 9910
rect 20275 9858 20331 9860
rect 20275 9806 20277 9858
rect 20277 9806 20329 9858
rect 20329 9806 20331 9858
rect 20275 9804 20331 9806
rect 21458 9908 21514 9964
rect 21562 9908 21618 9964
rect 21666 9908 21722 9964
rect 21458 9804 21514 9860
rect 21562 9804 21618 9860
rect 21666 9804 21722 9860
rect 21458 9470 21514 9526
rect 21562 9470 21618 9526
rect 21666 9470 21722 9526
rect 21458 9366 21514 9422
rect 21562 9366 21618 9422
rect 21666 9366 21722 9422
rect 21458 9262 21514 9318
rect 21562 9262 21618 9318
rect 21666 9262 21722 9318
rect 18995 9026 19051 9028
rect 18995 8974 18997 9026
rect 18997 8974 19049 9026
rect 19049 8974 19051 9026
rect 18995 8972 19051 8974
rect 18995 8922 19051 8924
rect 18995 8870 18997 8922
rect 18997 8870 19049 8922
rect 19049 8870 19051 8922
rect 18995 8868 19051 8870
rect 19635 9026 19691 9028
rect 19635 8974 19637 9026
rect 19637 8974 19689 9026
rect 19689 8974 19691 9026
rect 19635 8972 19691 8974
rect 19635 8922 19691 8924
rect 19635 8870 19637 8922
rect 19637 8870 19689 8922
rect 19689 8870 19691 8922
rect 19635 8868 19691 8870
rect 20275 9026 20331 9028
rect 20275 8974 20277 9026
rect 20277 8974 20329 9026
rect 20329 8974 20331 9026
rect 20275 8972 20331 8974
rect 20275 8922 20331 8924
rect 20275 8870 20277 8922
rect 20277 8870 20329 8922
rect 20329 8870 20331 8922
rect 20275 8868 20331 8870
rect 19075 8695 19131 8697
rect 19075 8643 19077 8695
rect 19077 8643 19129 8695
rect 19129 8643 19131 8695
rect 19075 8641 19131 8643
rect 19315 8484 19371 8486
rect 19315 8432 19317 8484
rect 19317 8432 19369 8484
rect 19369 8432 19371 8484
rect 19315 8430 19371 8432
rect 19315 8380 19371 8382
rect 19315 8328 19317 8380
rect 19317 8328 19369 8380
rect 19369 8328 19371 8380
rect 19315 8326 19371 8328
rect 19955 8484 20011 8486
rect 19955 8432 19957 8484
rect 19957 8432 20009 8484
rect 20009 8432 20011 8484
rect 19955 8430 20011 8432
rect 19955 8380 20011 8382
rect 19955 8328 19957 8380
rect 19957 8328 20009 8380
rect 20009 8328 20011 8380
rect 19955 8326 20011 8328
rect 24467 13164 24523 13166
rect 24467 13112 24469 13164
rect 24469 13112 24521 13164
rect 24521 13112 24523 13164
rect 24467 13110 24523 13112
rect 24467 13060 24523 13062
rect 24467 13008 24469 13060
rect 24469 13008 24521 13060
rect 24521 13008 24523 13060
rect 24467 13006 24523 13008
rect 25107 13164 25163 13166
rect 25107 13112 25109 13164
rect 25109 13112 25161 13164
rect 25161 13112 25163 13164
rect 25107 13110 25163 13112
rect 25107 13060 25163 13062
rect 25107 13008 25109 13060
rect 25109 13008 25161 13060
rect 25161 13008 25163 13060
rect 25107 13006 25163 13008
rect 22107 11884 22163 11940
rect 22211 11884 22267 11940
rect 22315 11884 22371 11940
rect 22107 11780 22163 11836
rect 22211 11780 22267 11836
rect 22315 11780 22371 11836
rect 22107 11676 22163 11732
rect 22211 11676 22267 11732
rect 22315 11676 22371 11732
rect 22107 11342 22163 11398
rect 22211 11342 22267 11398
rect 22315 11342 22371 11398
rect 22107 11238 22163 11294
rect 22211 11238 22267 11294
rect 22315 11238 22371 11294
rect 22107 11134 22163 11190
rect 22211 11134 22267 11190
rect 22315 11134 22371 11190
rect 22107 10406 22163 10462
rect 22211 10406 22267 10462
rect 22315 10406 22371 10462
rect 22107 10302 22163 10358
rect 22211 10302 22267 10358
rect 22315 10302 22371 10358
rect 22107 10198 22163 10254
rect 22211 10198 22267 10254
rect 22315 10198 22371 10254
rect 22107 9076 22163 9132
rect 22211 9076 22267 9132
rect 22315 9076 22371 9132
rect 22107 8972 22163 9028
rect 22211 8972 22267 9028
rect 22315 8972 22371 9028
rect 22107 8868 22163 8924
rect 22211 8868 22267 8924
rect 22315 8868 22371 8924
rect 22107 8534 22163 8590
rect 22211 8534 22267 8590
rect 22315 8534 22371 8590
rect 22107 8430 22163 8486
rect 22211 8430 22267 8486
rect 22315 8430 22371 8486
rect 22107 8326 22163 8382
rect 22211 8326 22267 8382
rect 22315 8326 22371 8382
rect 22756 12820 22812 12876
rect 22860 12820 22916 12876
rect 22964 12820 23020 12876
rect 22756 12716 22812 12772
rect 22860 12716 22916 12772
rect 22964 12716 23020 12772
rect 22756 12612 22812 12668
rect 22860 12612 22916 12668
rect 22964 12612 23020 12668
rect 24147 12770 24203 12772
rect 24147 12718 24149 12770
rect 24149 12718 24201 12770
rect 24201 12718 24203 12770
rect 24147 12716 24203 12718
rect 24147 12666 24203 12668
rect 24147 12614 24149 12666
rect 24149 12614 24201 12666
rect 24201 12614 24203 12666
rect 24147 12612 24203 12614
rect 24787 12770 24843 12772
rect 24787 12718 24789 12770
rect 24789 12718 24841 12770
rect 24841 12718 24843 12770
rect 24787 12716 24843 12718
rect 24787 12666 24843 12668
rect 24787 12614 24789 12666
rect 24789 12614 24841 12666
rect 24841 12614 24843 12666
rect 24787 12612 24843 12614
rect 25427 12770 25483 12772
rect 25427 12718 25429 12770
rect 25429 12718 25481 12770
rect 25481 12718 25483 12770
rect 25427 12716 25483 12718
rect 25427 12666 25483 12668
rect 25427 12614 25429 12666
rect 25429 12614 25481 12666
rect 25481 12614 25483 12666
rect 25427 12612 25483 12614
rect 22756 12278 22812 12334
rect 22860 12278 22916 12334
rect 22964 12278 23020 12334
rect 22756 12174 22812 12230
rect 22860 12174 22916 12230
rect 22964 12174 23020 12230
rect 22756 12070 22812 12126
rect 22860 12070 22916 12126
rect 22964 12070 23020 12126
rect 24467 12228 24523 12230
rect 24467 12176 24469 12228
rect 24469 12176 24521 12228
rect 24521 12176 24523 12228
rect 24467 12174 24523 12176
rect 24467 12124 24523 12126
rect 24467 12072 24469 12124
rect 24469 12072 24521 12124
rect 24521 12072 24523 12124
rect 24467 12070 24523 12072
rect 25347 12439 25403 12441
rect 25347 12387 25349 12439
rect 25349 12387 25401 12439
rect 25401 12387 25403 12439
rect 25347 12385 25403 12387
rect 26571 12385 26627 12441
rect 25107 12228 25163 12230
rect 25107 12176 25109 12228
rect 25109 12176 25161 12228
rect 25161 12176 25163 12228
rect 25107 12174 25163 12176
rect 25107 12124 25163 12126
rect 25107 12072 25109 12124
rect 25109 12072 25161 12124
rect 25161 12072 25163 12124
rect 25107 12070 25163 12072
rect 24147 11834 24203 11836
rect 24147 11782 24149 11834
rect 24149 11782 24201 11834
rect 24201 11782 24203 11834
rect 24147 11780 24203 11782
rect 24147 11730 24203 11732
rect 24147 11678 24149 11730
rect 24149 11678 24201 11730
rect 24201 11678 24203 11730
rect 24147 11676 24203 11678
rect 24787 11834 24843 11836
rect 24787 11782 24789 11834
rect 24789 11782 24841 11834
rect 24841 11782 24843 11834
rect 24787 11780 24843 11782
rect 24787 11730 24843 11732
rect 24787 11678 24789 11730
rect 24789 11678 24841 11730
rect 24841 11678 24843 11730
rect 24787 11676 24843 11678
rect 25427 11834 25483 11836
rect 25427 11782 25429 11834
rect 25429 11782 25481 11834
rect 25481 11782 25483 11834
rect 25427 11780 25483 11782
rect 25427 11730 25483 11732
rect 25427 11678 25429 11730
rect 25429 11678 25481 11730
rect 25481 11678 25483 11730
rect 25427 11676 25483 11678
rect 22756 10948 22812 11004
rect 22860 10948 22916 11004
rect 22964 10948 23020 11004
rect 24467 11292 24523 11294
rect 24467 11240 24469 11292
rect 24469 11240 24521 11292
rect 24521 11240 24523 11292
rect 24467 11238 24523 11240
rect 24467 11188 24523 11190
rect 24467 11136 24469 11188
rect 24469 11136 24521 11188
rect 24521 11136 24523 11188
rect 24467 11134 24523 11136
rect 25347 11503 25403 11505
rect 25347 11451 25349 11503
rect 25349 11451 25401 11503
rect 25401 11451 25403 11503
rect 25347 11449 25403 11451
rect 25107 11292 25163 11294
rect 25107 11240 25109 11292
rect 25109 11240 25161 11292
rect 25161 11240 25163 11292
rect 25107 11238 25163 11240
rect 25107 11188 25163 11190
rect 25107 11136 25109 11188
rect 25109 11136 25161 11188
rect 25161 11136 25163 11188
rect 25107 11134 25163 11136
rect 22756 10844 22812 10900
rect 22860 10844 22916 10900
rect 22964 10844 23020 10900
rect 22756 10740 22812 10796
rect 22860 10740 22916 10796
rect 22964 10740 23020 10796
rect 24147 10898 24203 10900
rect 24147 10846 24149 10898
rect 24149 10846 24201 10898
rect 24201 10846 24203 10898
rect 24147 10844 24203 10846
rect 24147 10794 24203 10796
rect 24147 10742 24149 10794
rect 24149 10742 24201 10794
rect 24201 10742 24203 10794
rect 24147 10740 24203 10742
rect 24787 10898 24843 10900
rect 24787 10846 24789 10898
rect 24789 10846 24841 10898
rect 24841 10846 24843 10898
rect 24787 10844 24843 10846
rect 24787 10794 24843 10796
rect 24787 10742 24789 10794
rect 24789 10742 24841 10794
rect 24841 10742 24843 10794
rect 24787 10740 24843 10742
rect 25427 10898 25483 10900
rect 25427 10846 25429 10898
rect 25429 10846 25481 10898
rect 25481 10846 25483 10898
rect 25427 10844 25483 10846
rect 25427 10794 25483 10796
rect 25427 10742 25429 10794
rect 25429 10742 25481 10794
rect 25481 10742 25483 10794
rect 25427 10740 25483 10742
rect 22756 10012 22812 10068
rect 22860 10012 22916 10068
rect 22964 10012 23020 10068
rect 22756 9908 22812 9964
rect 22860 9908 22916 9964
rect 22964 9908 23020 9964
rect 22756 9804 22812 9860
rect 22860 9804 22916 9860
rect 22964 9804 23020 9860
rect 24147 9962 24203 9964
rect 24147 9910 24149 9962
rect 24149 9910 24201 9962
rect 24201 9910 24203 9962
rect 24147 9908 24203 9910
rect 24147 9858 24203 9860
rect 24147 9806 24149 9858
rect 24149 9806 24201 9858
rect 24201 9806 24203 9858
rect 24147 9804 24203 9806
rect 22756 9470 22812 9526
rect 22860 9470 22916 9526
rect 22964 9470 23020 9526
rect 22756 9366 22812 9422
rect 22860 9366 22916 9422
rect 22964 9366 23020 9422
rect 22756 9262 22812 9318
rect 22860 9262 22916 9318
rect 22964 9262 23020 9318
rect 21458 8140 21514 8196
rect 21562 8140 21618 8196
rect 21666 8140 21722 8196
rect 18995 8090 19051 8092
rect 18995 8038 18997 8090
rect 18997 8038 19049 8090
rect 19049 8038 19051 8090
rect 18995 8036 19051 8038
rect 18995 7986 19051 7988
rect 18995 7934 18997 7986
rect 18997 7934 19049 7986
rect 19049 7934 19051 7986
rect 18995 7932 19051 7934
rect 19635 8090 19691 8092
rect 19635 8038 19637 8090
rect 19637 8038 19689 8090
rect 19689 8038 19691 8090
rect 19635 8036 19691 8038
rect 19635 7986 19691 7988
rect 19635 7934 19637 7986
rect 19637 7934 19689 7986
rect 19689 7934 19691 7986
rect 19635 7932 19691 7934
rect 20275 8090 20331 8092
rect 20275 8038 20277 8090
rect 20277 8038 20329 8090
rect 20329 8038 20331 8090
rect 20275 8036 20331 8038
rect 20275 7986 20331 7988
rect 20275 7934 20277 7986
rect 20277 7934 20329 7986
rect 20329 7934 20331 7986
rect 20275 7932 20331 7934
rect 21458 8036 21514 8092
rect 21562 8036 21618 8092
rect 21666 8036 21722 8092
rect 21458 7932 21514 7988
rect 21562 7932 21618 7988
rect 21666 7932 21722 7988
rect 24467 10356 24523 10358
rect 24467 10304 24469 10356
rect 24469 10304 24521 10356
rect 24521 10304 24523 10356
rect 24467 10302 24523 10304
rect 24467 10252 24523 10254
rect 24467 10200 24469 10252
rect 24469 10200 24521 10252
rect 24521 10200 24523 10252
rect 24467 10198 24523 10200
rect 24467 9420 24523 9422
rect 24467 9368 24469 9420
rect 24469 9368 24521 9420
rect 24521 9368 24523 9420
rect 24467 9366 24523 9368
rect 24467 9316 24523 9318
rect 24467 9264 24469 9316
rect 24469 9264 24521 9316
rect 24521 9264 24523 9316
rect 24467 9262 24523 9264
rect 24787 9962 24843 9964
rect 24787 9910 24789 9962
rect 24789 9910 24841 9962
rect 24841 9910 24843 9962
rect 24787 9908 24843 9910
rect 24787 9858 24843 9860
rect 24787 9806 24789 9858
rect 24789 9806 24841 9858
rect 24841 9806 24843 9858
rect 24787 9804 24843 9806
rect 25107 10356 25163 10358
rect 25107 10304 25109 10356
rect 25109 10304 25161 10356
rect 25161 10304 25163 10356
rect 25107 10302 25163 10304
rect 25107 10252 25163 10254
rect 25107 10200 25109 10252
rect 25109 10200 25161 10252
rect 25161 10200 25163 10252
rect 25107 10198 25163 10200
rect 25427 9962 25483 9964
rect 25427 9910 25429 9962
rect 25429 9910 25481 9962
rect 25481 9910 25483 9962
rect 25427 9908 25483 9910
rect 25427 9858 25483 9860
rect 25427 9806 25429 9858
rect 25429 9806 25481 9858
rect 25481 9806 25483 9858
rect 25427 9804 25483 9806
rect 25347 9631 25403 9633
rect 25347 9579 25349 9631
rect 25349 9579 25401 9631
rect 25401 9579 25403 9631
rect 25347 9577 25403 9579
rect 26571 9577 26627 9633
rect 25107 9420 25163 9422
rect 25107 9368 25109 9420
rect 25109 9368 25161 9420
rect 25161 9368 25163 9420
rect 25107 9366 25163 9368
rect 25107 9316 25163 9318
rect 25107 9264 25109 9316
rect 25109 9264 25161 9316
rect 25161 9264 25163 9316
rect 25107 9262 25163 9264
rect 24147 9026 24203 9028
rect 24147 8974 24149 9026
rect 24149 8974 24201 9026
rect 24201 8974 24203 9026
rect 24147 8972 24203 8974
rect 24147 8922 24203 8924
rect 24147 8870 24149 8922
rect 24149 8870 24201 8922
rect 24201 8870 24203 8922
rect 24147 8868 24203 8870
rect 24787 9026 24843 9028
rect 24787 8974 24789 9026
rect 24789 8974 24841 9026
rect 24841 8974 24843 9026
rect 24787 8972 24843 8974
rect 24787 8922 24843 8924
rect 24787 8870 24789 8922
rect 24789 8870 24841 8922
rect 24841 8870 24843 8922
rect 24787 8868 24843 8870
rect 25427 9026 25483 9028
rect 25427 8974 25429 9026
rect 25429 8974 25481 9026
rect 25481 8974 25483 9026
rect 25427 8972 25483 8974
rect 25427 8922 25483 8924
rect 25427 8870 25429 8922
rect 25429 8870 25481 8922
rect 25481 8870 25483 8922
rect 25427 8868 25483 8870
rect 22756 8140 22812 8196
rect 22860 8140 22916 8196
rect 22964 8140 23020 8196
rect 24467 8484 24523 8486
rect 24467 8432 24469 8484
rect 24469 8432 24521 8484
rect 24521 8432 24523 8484
rect 24467 8430 24523 8432
rect 24467 8380 24523 8382
rect 24467 8328 24469 8380
rect 24469 8328 24521 8380
rect 24521 8328 24523 8380
rect 24467 8326 24523 8328
rect 25347 8695 25403 8697
rect 25347 8643 25349 8695
rect 25349 8643 25401 8695
rect 25401 8643 25403 8695
rect 25347 8641 25403 8643
rect 25107 8484 25163 8486
rect 25107 8432 25109 8484
rect 25109 8432 25161 8484
rect 25161 8432 25163 8484
rect 25107 8430 25163 8432
rect 25107 8380 25163 8382
rect 25107 8328 25109 8380
rect 25109 8328 25161 8380
rect 25161 8328 25163 8380
rect 25107 8326 25163 8328
rect 22756 8036 22812 8092
rect 22860 8036 22916 8092
rect 22964 8036 23020 8092
rect 22756 7932 22812 7988
rect 22860 7932 22916 7988
rect 22964 7932 23020 7988
rect 24147 8090 24203 8092
rect 24147 8038 24149 8090
rect 24149 8038 24201 8090
rect 24201 8038 24203 8090
rect 24147 8036 24203 8038
rect 24147 7986 24203 7988
rect 24147 7934 24149 7986
rect 24149 7934 24201 7986
rect 24201 7934 24203 7986
rect 24147 7932 24203 7934
rect 24787 8090 24843 8092
rect 24787 8038 24789 8090
rect 24789 8038 24841 8090
rect 24841 8038 24843 8090
rect 24787 8036 24843 8038
rect 24787 7986 24843 7988
rect 24787 7934 24789 7986
rect 24789 7934 24841 7986
rect 24841 7934 24843 7986
rect 24787 7932 24843 7934
rect 25427 8090 25483 8092
rect 25427 8038 25429 8090
rect 25429 8038 25481 8090
rect 25481 8038 25483 8090
rect 25427 8036 25483 8038
rect 25427 7986 25483 7988
rect 25427 7934 25429 7986
rect 25429 7934 25481 7986
rect 25481 7934 25483 7986
rect 25427 7932 25483 7934
rect 17851 7705 17907 7761
rect 19235 7759 19291 7761
rect 19235 7707 19237 7759
rect 19237 7707 19289 7759
rect 19289 7707 19291 7759
rect 19235 7705 19291 7707
rect 19875 7759 19931 7761
rect 19875 7707 19877 7759
rect 19877 7707 19929 7759
rect 19929 7707 19931 7759
rect 19875 7705 19931 7707
rect 24547 7759 24603 7761
rect 24547 7707 24549 7759
rect 24549 7707 24601 7759
rect 24601 7707 24603 7759
rect 24547 7705 24603 7707
rect 25187 7759 25243 7761
rect 25187 7707 25189 7759
rect 25189 7707 25241 7759
rect 25241 7707 25243 7759
rect 25187 7705 25243 7707
rect 28196 13405 28252 13407
rect 28196 13353 28198 13405
rect 28198 13353 28250 13405
rect 28250 13353 28252 13405
rect 28196 13351 28252 13353
rect 31228 13214 31284 13270
rect 31332 13214 31388 13270
rect 31436 13214 31492 13270
rect 28436 13164 28492 13166
rect 28436 13112 28438 13164
rect 28438 13112 28490 13164
rect 28490 13112 28492 13164
rect 28436 13110 28492 13112
rect 28436 13060 28492 13062
rect 28436 13008 28438 13060
rect 28438 13008 28490 13060
rect 28490 13008 28492 13060
rect 28436 13006 28492 13008
rect 29076 13164 29132 13166
rect 29076 13112 29078 13164
rect 29078 13112 29130 13164
rect 29130 13112 29132 13164
rect 29076 13110 29132 13112
rect 29076 13060 29132 13062
rect 29076 13008 29078 13060
rect 29078 13008 29130 13060
rect 29130 13008 29132 13060
rect 29076 13006 29132 13008
rect 31228 13110 31284 13166
rect 31332 13110 31388 13166
rect 31436 13110 31492 13166
rect 31228 13006 31284 13062
rect 31332 13006 31388 13062
rect 31436 13006 31492 13062
rect 30579 12820 30635 12876
rect 30683 12820 30739 12876
rect 30787 12820 30843 12876
rect 28116 12770 28172 12772
rect 28116 12718 28118 12770
rect 28118 12718 28170 12770
rect 28170 12718 28172 12770
rect 28116 12716 28172 12718
rect 28116 12666 28172 12668
rect 28116 12614 28118 12666
rect 28118 12614 28170 12666
rect 28170 12614 28172 12666
rect 28116 12612 28172 12614
rect 28756 12770 28812 12772
rect 28756 12718 28758 12770
rect 28758 12718 28810 12770
rect 28810 12718 28812 12770
rect 28756 12716 28812 12718
rect 28756 12666 28812 12668
rect 28756 12614 28758 12666
rect 28758 12614 28810 12666
rect 28810 12614 28812 12666
rect 28756 12612 28812 12614
rect 29396 12770 29452 12772
rect 29396 12718 29398 12770
rect 29398 12718 29450 12770
rect 29450 12718 29452 12770
rect 29396 12716 29452 12718
rect 29396 12666 29452 12668
rect 29396 12614 29398 12666
rect 29398 12614 29450 12666
rect 29450 12614 29452 12666
rect 29396 12612 29452 12614
rect 30579 12716 30635 12772
rect 30683 12716 30739 12772
rect 30787 12716 30843 12772
rect 30579 12612 30635 12668
rect 30683 12612 30739 12668
rect 30787 12612 30843 12668
rect 26771 11449 26828 11505
rect 26771 8641 26828 8697
rect 26972 12385 27028 12441
rect 28196 12439 28252 12441
rect 28196 12387 28198 12439
rect 28198 12387 28250 12439
rect 28250 12387 28252 12439
rect 28196 12385 28252 12387
rect 28436 12228 28492 12230
rect 28436 12176 28438 12228
rect 28438 12176 28490 12228
rect 28490 12176 28492 12228
rect 28436 12174 28492 12176
rect 28436 12124 28492 12126
rect 28436 12072 28438 12124
rect 28438 12072 28490 12124
rect 28490 12072 28492 12124
rect 28436 12070 28492 12072
rect 29076 12228 29132 12230
rect 29076 12176 29078 12228
rect 29078 12176 29130 12228
rect 29130 12176 29132 12228
rect 29076 12174 29132 12176
rect 29076 12124 29132 12126
rect 29076 12072 29078 12124
rect 29078 12072 29130 12124
rect 29130 12072 29132 12124
rect 29076 12070 29132 12072
rect 30579 12278 30635 12334
rect 30683 12278 30739 12334
rect 30787 12278 30843 12334
rect 30579 12174 30635 12230
rect 30683 12174 30739 12230
rect 30787 12174 30843 12230
rect 30579 12070 30635 12126
rect 30683 12070 30739 12126
rect 30787 12070 30843 12126
rect 28116 11834 28172 11836
rect 28116 11782 28118 11834
rect 28118 11782 28170 11834
rect 28170 11782 28172 11834
rect 28116 11780 28172 11782
rect 28116 11730 28172 11732
rect 28116 11678 28118 11730
rect 28118 11678 28170 11730
rect 28170 11678 28172 11730
rect 28116 11676 28172 11678
rect 28756 11834 28812 11836
rect 28756 11782 28758 11834
rect 28758 11782 28810 11834
rect 28810 11782 28812 11834
rect 28756 11780 28812 11782
rect 28756 11730 28812 11732
rect 28756 11678 28758 11730
rect 28758 11678 28810 11730
rect 28810 11678 28812 11730
rect 28756 11676 28812 11678
rect 29396 11834 29452 11836
rect 29396 11782 29398 11834
rect 29398 11782 29450 11834
rect 29450 11782 29452 11834
rect 29396 11780 29452 11782
rect 29396 11730 29452 11732
rect 29396 11678 29398 11730
rect 29398 11678 29450 11730
rect 29450 11678 29452 11730
rect 29396 11676 29452 11678
rect 28196 11503 28252 11505
rect 28196 11451 28198 11503
rect 28198 11451 28250 11503
rect 28250 11451 28252 11503
rect 28196 11449 28252 11451
rect 28436 11292 28492 11294
rect 28436 11240 28438 11292
rect 28438 11240 28490 11292
rect 28490 11240 28492 11292
rect 28436 11238 28492 11240
rect 28436 11188 28492 11190
rect 28436 11136 28438 11188
rect 28438 11136 28490 11188
rect 28490 11136 28492 11188
rect 28436 11134 28492 11136
rect 29076 11292 29132 11294
rect 29076 11240 29078 11292
rect 29078 11240 29130 11292
rect 29130 11240 29132 11292
rect 29076 11238 29132 11240
rect 29076 11188 29132 11190
rect 29076 11136 29078 11188
rect 29078 11136 29130 11188
rect 29130 11136 29132 11188
rect 29076 11134 29132 11136
rect 30579 10948 30635 11004
rect 30683 10948 30739 11004
rect 30787 10948 30843 11004
rect 28116 10898 28172 10900
rect 28116 10846 28118 10898
rect 28118 10846 28170 10898
rect 28170 10846 28172 10898
rect 28116 10844 28172 10846
rect 28116 10794 28172 10796
rect 28116 10742 28118 10794
rect 28118 10742 28170 10794
rect 28170 10742 28172 10794
rect 28116 10740 28172 10742
rect 28756 10898 28812 10900
rect 28756 10846 28758 10898
rect 28758 10846 28810 10898
rect 28810 10846 28812 10898
rect 28756 10844 28812 10846
rect 28756 10794 28812 10796
rect 28756 10742 28758 10794
rect 28758 10742 28810 10794
rect 28810 10742 28812 10794
rect 28756 10740 28812 10742
rect 29396 10898 29452 10900
rect 29396 10846 29398 10898
rect 29398 10846 29450 10898
rect 29450 10846 29452 10898
rect 29396 10844 29452 10846
rect 29396 10794 29452 10796
rect 29396 10742 29398 10794
rect 29398 10742 29450 10794
rect 29450 10742 29452 10794
rect 29396 10740 29452 10742
rect 30579 10844 30635 10900
rect 30683 10844 30739 10900
rect 30787 10844 30843 10900
rect 30579 10740 30635 10796
rect 30683 10740 30739 10796
rect 30787 10740 30843 10796
rect 28436 10356 28492 10358
rect 28436 10304 28438 10356
rect 28438 10304 28490 10356
rect 28490 10304 28492 10356
rect 28436 10302 28492 10304
rect 28436 10252 28492 10254
rect 28436 10200 28438 10252
rect 28438 10200 28490 10252
rect 28490 10200 28492 10252
rect 28436 10198 28492 10200
rect 28116 9962 28172 9964
rect 28116 9910 28118 9962
rect 28118 9910 28170 9962
rect 28170 9910 28172 9962
rect 28116 9908 28172 9910
rect 28116 9858 28172 9860
rect 28116 9806 28118 9858
rect 28118 9806 28170 9858
rect 28170 9806 28172 9858
rect 28116 9804 28172 9806
rect 26972 9577 27028 9633
rect 26571 7705 26627 7761
rect 28196 9631 28252 9633
rect 28196 9579 28198 9631
rect 28198 9579 28250 9631
rect 28250 9579 28252 9631
rect 28196 9577 28252 9579
rect 28436 9420 28492 9422
rect 28436 9368 28438 9420
rect 28438 9368 28490 9420
rect 28490 9368 28492 9420
rect 28436 9366 28492 9368
rect 28436 9316 28492 9318
rect 28436 9264 28438 9316
rect 28438 9264 28490 9316
rect 28490 9264 28492 9316
rect 28436 9262 28492 9264
rect 28756 9962 28812 9964
rect 28756 9910 28758 9962
rect 28758 9910 28810 9962
rect 28810 9910 28812 9962
rect 28756 9908 28812 9910
rect 28756 9858 28812 9860
rect 28756 9806 28758 9858
rect 28758 9806 28810 9858
rect 28810 9806 28812 9858
rect 28756 9804 28812 9806
rect 29076 10356 29132 10358
rect 29076 10304 29078 10356
rect 29078 10304 29130 10356
rect 29130 10304 29132 10356
rect 29076 10302 29132 10304
rect 29076 10252 29132 10254
rect 29076 10200 29078 10252
rect 29078 10200 29130 10252
rect 29130 10200 29132 10252
rect 29076 10198 29132 10200
rect 29076 9420 29132 9422
rect 29076 9368 29078 9420
rect 29078 9368 29130 9420
rect 29130 9368 29132 9420
rect 29076 9366 29132 9368
rect 29076 9316 29132 9318
rect 29076 9264 29078 9316
rect 29078 9264 29130 9316
rect 29130 9264 29132 9316
rect 29076 9262 29132 9264
rect 30579 10012 30635 10068
rect 30683 10012 30739 10068
rect 30787 10012 30843 10068
rect 29396 9962 29452 9964
rect 29396 9910 29398 9962
rect 29398 9910 29450 9962
rect 29450 9910 29452 9962
rect 29396 9908 29452 9910
rect 29396 9858 29452 9860
rect 29396 9806 29398 9858
rect 29398 9806 29450 9858
rect 29450 9806 29452 9858
rect 29396 9804 29452 9806
rect 30579 9908 30635 9964
rect 30683 9908 30739 9964
rect 30787 9908 30843 9964
rect 30579 9804 30635 9860
rect 30683 9804 30739 9860
rect 30787 9804 30843 9860
rect 30579 9470 30635 9526
rect 30683 9470 30739 9526
rect 30787 9470 30843 9526
rect 30579 9366 30635 9422
rect 30683 9366 30739 9422
rect 30787 9366 30843 9422
rect 30579 9262 30635 9318
rect 30683 9262 30739 9318
rect 30787 9262 30843 9318
rect 28116 9026 28172 9028
rect 28116 8974 28118 9026
rect 28118 8974 28170 9026
rect 28170 8974 28172 9026
rect 28116 8972 28172 8974
rect 28116 8922 28172 8924
rect 28116 8870 28118 8922
rect 28118 8870 28170 8922
rect 28170 8870 28172 8922
rect 28116 8868 28172 8870
rect 28756 9026 28812 9028
rect 28756 8974 28758 9026
rect 28758 8974 28810 9026
rect 28810 8974 28812 9026
rect 28756 8972 28812 8974
rect 28756 8922 28812 8924
rect 28756 8870 28758 8922
rect 28758 8870 28810 8922
rect 28810 8870 28812 8922
rect 28756 8868 28812 8870
rect 29396 9026 29452 9028
rect 29396 8974 29398 9026
rect 29398 8974 29450 9026
rect 29450 8974 29452 9026
rect 29396 8972 29452 8974
rect 29396 8922 29452 8924
rect 29396 8870 29398 8922
rect 29398 8870 29450 8922
rect 29450 8870 29452 8922
rect 29396 8868 29452 8870
rect 28196 8695 28252 8697
rect 28196 8643 28198 8695
rect 28198 8643 28250 8695
rect 28250 8643 28252 8695
rect 28196 8641 28252 8643
rect 28436 8484 28492 8486
rect 28436 8432 28438 8484
rect 28438 8432 28490 8484
rect 28490 8432 28492 8484
rect 28436 8430 28492 8432
rect 28436 8380 28492 8382
rect 28436 8328 28438 8380
rect 28438 8328 28490 8380
rect 28490 8328 28492 8380
rect 28436 8326 28492 8328
rect 29076 8484 29132 8486
rect 29076 8432 29078 8484
rect 29078 8432 29130 8484
rect 29130 8432 29132 8484
rect 29076 8430 29132 8432
rect 29076 8380 29132 8382
rect 29076 8328 29078 8380
rect 29078 8328 29130 8380
rect 29130 8328 29132 8380
rect 29076 8326 29132 8328
rect 30579 8140 30635 8196
rect 30683 8140 30739 8196
rect 30787 8140 30843 8196
rect 28116 8090 28172 8092
rect 28116 8038 28118 8090
rect 28118 8038 28170 8090
rect 28170 8038 28172 8090
rect 28116 8036 28172 8038
rect 28116 7986 28172 7988
rect 28116 7934 28118 7986
rect 28118 7934 28170 7986
rect 28170 7934 28172 7986
rect 28116 7932 28172 7934
rect 28756 8090 28812 8092
rect 28756 8038 28758 8090
rect 28758 8038 28810 8090
rect 28810 8038 28812 8090
rect 28756 8036 28812 8038
rect 28756 7986 28812 7988
rect 28756 7934 28758 7986
rect 28758 7934 28810 7986
rect 28810 7934 28812 7986
rect 28756 7932 28812 7934
rect 29396 8090 29452 8092
rect 29396 8038 29398 8090
rect 29398 8038 29450 8090
rect 29450 8038 29452 8090
rect 29396 8036 29452 8038
rect 29396 7986 29452 7988
rect 29396 7934 29398 7986
rect 29398 7934 29450 7986
rect 29450 7934 29452 7986
rect 29396 7932 29452 7934
rect 30579 8036 30635 8092
rect 30683 8036 30739 8092
rect 30787 8036 30843 8092
rect 30579 7932 30635 7988
rect 30683 7932 30739 7988
rect 30787 7932 30843 7988
rect 31228 11884 31284 11940
rect 31332 11884 31388 11940
rect 31436 11884 31492 11940
rect 31228 11780 31284 11836
rect 31332 11780 31388 11836
rect 31436 11780 31492 11836
rect 32136 12820 32192 12876
rect 32240 12820 32296 12876
rect 32344 12820 32400 12876
rect 34588 12994 34644 13050
rect 34692 12994 34748 13050
rect 34796 12994 34852 13050
rect 34588 12890 34644 12946
rect 34692 12890 34748 12946
rect 34796 12890 34852 12946
rect 34588 12786 34644 12842
rect 34692 12786 34748 12842
rect 34796 12786 34852 12842
rect 38724 12994 38780 13050
rect 38828 12994 38884 13050
rect 38932 12994 38988 13050
rect 38724 12890 38780 12946
rect 38828 12890 38884 12946
rect 38932 12890 38988 12946
rect 38724 12786 38780 12842
rect 38828 12786 38884 12842
rect 38932 12786 38988 12842
rect 44284 12994 44340 13050
rect 44388 12994 44444 13050
rect 44492 12994 44548 13050
rect 44284 12890 44340 12946
rect 44388 12890 44444 12946
rect 44492 12890 44548 12946
rect 44284 12786 44340 12842
rect 44388 12786 44444 12842
rect 44492 12786 44548 12842
rect 48420 12994 48476 13050
rect 48524 12994 48580 13050
rect 48628 12994 48684 13050
rect 48420 12890 48476 12946
rect 48524 12890 48580 12946
rect 48628 12890 48684 12946
rect 48420 12786 48476 12842
rect 48524 12786 48580 12842
rect 48628 12786 48684 12842
rect 53980 12994 54036 13050
rect 54084 12994 54140 13050
rect 54188 12994 54244 13050
rect 53980 12890 54036 12946
rect 54084 12890 54140 12946
rect 54188 12890 54244 12946
rect 53980 12786 54036 12842
rect 54084 12786 54140 12842
rect 54188 12786 54244 12842
rect 58116 12994 58172 13050
rect 58220 12994 58276 13050
rect 58324 12994 58380 13050
rect 58116 12890 58172 12946
rect 58220 12890 58276 12946
rect 58324 12890 58380 12946
rect 58116 12786 58172 12842
rect 58220 12786 58276 12842
rect 58324 12786 58380 12842
rect 63676 12994 63732 13050
rect 63780 12994 63836 13050
rect 63884 12994 63940 13050
rect 63676 12890 63732 12946
rect 63780 12890 63836 12946
rect 63884 12890 63940 12946
rect 63676 12786 63732 12842
rect 63780 12786 63836 12842
rect 63884 12786 63940 12842
rect 66924 13048 66980 13050
rect 66924 12996 66926 13048
rect 66926 12996 66978 13048
rect 66978 12996 66980 13048
rect 66924 12994 66980 12996
rect 67028 13048 67084 13050
rect 67028 12996 67030 13048
rect 67030 12996 67082 13048
rect 67082 12996 67084 13048
rect 67028 12994 67084 12996
rect 67132 13048 67188 13050
rect 67132 12996 67134 13048
rect 67134 12996 67186 13048
rect 67186 12996 67188 13048
rect 67132 12994 67188 12996
rect 66924 12944 66980 12946
rect 66924 12892 66926 12944
rect 66926 12892 66978 12944
rect 66978 12892 66980 12944
rect 66924 12890 66980 12892
rect 67028 12944 67084 12946
rect 67028 12892 67030 12944
rect 67030 12892 67082 12944
rect 67082 12892 67084 12944
rect 67028 12890 67084 12892
rect 67132 12944 67188 12946
rect 67132 12892 67134 12944
rect 67134 12892 67186 12944
rect 67186 12892 67188 12944
rect 67132 12890 67188 12892
rect 66924 12840 66980 12842
rect 66924 12788 66926 12840
rect 66926 12788 66978 12840
rect 66978 12788 66980 12840
rect 66924 12786 66980 12788
rect 67028 12840 67084 12842
rect 67028 12788 67030 12840
rect 67030 12788 67082 12840
rect 67082 12788 67084 12840
rect 67028 12786 67084 12788
rect 67132 12840 67188 12842
rect 67132 12788 67134 12840
rect 67134 12788 67186 12840
rect 67186 12788 67188 12840
rect 67132 12786 67188 12788
rect 32136 12716 32192 12772
rect 32240 12716 32296 12772
rect 32344 12716 32400 12772
rect 32136 12612 32192 12668
rect 32240 12612 32296 12668
rect 32344 12612 32400 12668
rect 32136 12278 32192 12334
rect 32240 12278 32296 12334
rect 32344 12278 32400 12334
rect 32136 12174 32192 12230
rect 32240 12174 32296 12230
rect 32344 12174 32400 12230
rect 32136 12070 32192 12126
rect 32240 12070 32296 12126
rect 32344 12070 32400 12126
rect 31228 11676 31284 11732
rect 31332 11676 31388 11732
rect 31436 11676 31492 11732
rect 31228 11342 31284 11398
rect 31332 11342 31388 11398
rect 31436 11342 31492 11398
rect 31228 11238 31284 11294
rect 31332 11238 31388 11294
rect 31436 11238 31492 11294
rect 31228 11134 31284 11190
rect 31332 11134 31388 11190
rect 31436 11134 31492 11190
rect 31228 10406 31284 10462
rect 31332 10406 31388 10462
rect 31436 10406 31492 10462
rect 31228 10302 31284 10358
rect 31332 10302 31388 10358
rect 31436 10302 31492 10358
rect 31228 10198 31284 10254
rect 31332 10198 31388 10254
rect 31436 10198 31492 10254
rect 31228 9076 31284 9132
rect 31332 9076 31388 9132
rect 31436 9076 31492 9132
rect 31228 8972 31284 9028
rect 31332 8972 31388 9028
rect 31436 8972 31492 9028
rect 31228 8868 31284 8924
rect 31332 8868 31388 8924
rect 31436 8868 31492 8924
rect 31228 8534 31284 8590
rect 31332 8534 31388 8590
rect 31436 8534 31492 8590
rect 31228 8430 31284 8486
rect 31332 8430 31388 8486
rect 31436 8430 31492 8486
rect 31228 8326 31284 8382
rect 31332 8326 31388 8382
rect 31436 8326 31492 8382
rect 26972 7705 27028 7761
rect 28356 7759 28412 7761
rect 28356 7707 28358 7759
rect 28358 7707 28410 7759
rect 28410 7707 28412 7759
rect 28356 7705 28412 7707
rect 17129 6436 17185 6438
rect 17129 6384 17131 6436
rect 17131 6384 17183 6436
rect 17183 6384 17185 6436
rect 17129 6382 17185 6384
rect 17233 6436 17289 6438
rect 17233 6384 17235 6436
rect 17235 6384 17287 6436
rect 17287 6384 17289 6436
rect 17233 6382 17289 6384
rect 17337 6436 17393 6438
rect 17337 6384 17339 6436
rect 17339 6384 17391 6436
rect 17391 6384 17393 6436
rect 17337 6382 17393 6384
rect 17129 6332 17185 6334
rect 17129 6280 17131 6332
rect 17131 6280 17183 6332
rect 17183 6280 17185 6332
rect 17129 6278 17185 6280
rect 17233 6332 17289 6334
rect 17233 6280 17235 6332
rect 17235 6280 17287 6332
rect 17287 6280 17289 6332
rect 17233 6278 17289 6280
rect 17337 6332 17393 6334
rect 17337 6280 17339 6332
rect 17339 6280 17391 6332
rect 17391 6280 17393 6332
rect 17337 6278 17393 6280
rect 17129 6228 17185 6230
rect 17129 6176 17131 6228
rect 17131 6176 17183 6228
rect 17183 6176 17185 6228
rect 17129 6174 17185 6176
rect 17233 6228 17289 6230
rect 17233 6176 17235 6228
rect 17235 6176 17287 6228
rect 17287 6176 17289 6228
rect 17233 6174 17289 6176
rect 17337 6228 17393 6230
rect 17337 6176 17339 6228
rect 17339 6176 17391 6228
rect 17391 6176 17393 6228
rect 17337 6174 17393 6176
rect 30298 6382 30354 6438
rect 30402 6382 30458 6438
rect 30506 6382 30562 6438
rect 30610 6382 30666 6438
rect 30714 6382 30770 6438
rect 30298 6278 30354 6334
rect 30402 6278 30458 6334
rect 30506 6278 30562 6334
rect 30610 6278 30666 6334
rect 30714 6278 30770 6334
rect 30298 6174 30354 6230
rect 30402 6174 30458 6230
rect 30506 6174 30562 6230
rect 30610 6174 30666 6230
rect 30714 6174 30770 6230
rect 17566 6094 17622 6096
rect 17566 6042 17568 6094
rect 17568 6042 17620 6094
rect 17620 6042 17622 6094
rect 17566 6040 17622 6042
rect 17670 6094 17726 6096
rect 17670 6042 17672 6094
rect 17672 6042 17724 6094
rect 17724 6042 17726 6094
rect 17670 6040 17726 6042
rect 17774 6094 17830 6096
rect 17774 6042 17776 6094
rect 17776 6042 17828 6094
rect 17828 6042 17830 6094
rect 17774 6040 17830 6042
rect 17566 5990 17622 5992
rect 17566 5938 17568 5990
rect 17568 5938 17620 5990
rect 17620 5938 17622 5990
rect 17566 5936 17622 5938
rect 17670 5990 17726 5992
rect 17670 5938 17672 5990
rect 17672 5938 17724 5990
rect 17724 5938 17726 5990
rect 17670 5936 17726 5938
rect 17774 5990 17830 5992
rect 17774 5938 17776 5990
rect 17776 5938 17828 5990
rect 17828 5938 17830 5990
rect 17774 5936 17830 5938
rect 17566 5886 17622 5888
rect 17566 5834 17568 5886
rect 17568 5834 17620 5886
rect 17620 5834 17622 5886
rect 17566 5832 17622 5834
rect 17670 5886 17726 5888
rect 17670 5834 17672 5886
rect 17672 5834 17724 5886
rect 17724 5834 17726 5886
rect 17670 5832 17726 5834
rect 17774 5886 17830 5888
rect 17774 5834 17776 5886
rect 17776 5834 17828 5886
rect 17828 5834 17830 5886
rect 17774 5832 17830 5834
rect 29738 6040 29794 6096
rect 29842 6040 29898 6096
rect 29946 6040 30002 6096
rect 30050 6040 30106 6096
rect 30154 6040 30210 6096
rect 29738 5936 29794 5992
rect 29842 5936 29898 5992
rect 29946 5936 30002 5992
rect 30050 5936 30106 5992
rect 30154 5936 30210 5992
rect 29738 5832 29794 5888
rect 29842 5832 29898 5888
rect 29946 5832 30002 5888
rect 30050 5832 30106 5888
rect 30154 5832 30210 5888
rect 14696 5709 14752 5711
rect 14696 5657 14698 5709
rect 14698 5657 14750 5709
rect 14750 5657 14752 5709
rect 14696 5655 14752 5657
rect 14800 5709 14856 5711
rect 14800 5657 14802 5709
rect 14802 5657 14854 5709
rect 14854 5657 14856 5709
rect 14800 5655 14856 5657
rect 14696 5605 14752 5607
rect 14696 5553 14698 5605
rect 14698 5553 14750 5605
rect 14750 5553 14752 5605
rect 14696 5551 14752 5553
rect 14800 5605 14856 5607
rect 14800 5553 14802 5605
rect 14802 5553 14854 5605
rect 14854 5553 14856 5605
rect 14800 5551 14856 5553
rect 17344 5444 17400 5446
rect 17344 5392 17346 5444
rect 17346 5392 17398 5444
rect 17398 5392 17400 5444
rect 17344 5390 17400 5392
rect 17448 5444 17504 5446
rect 17448 5392 17450 5444
rect 17450 5392 17502 5444
rect 17502 5392 17504 5444
rect 17448 5390 17504 5392
rect 17344 5340 17400 5342
rect 17344 5288 17346 5340
rect 17346 5288 17398 5340
rect 17398 5288 17400 5340
rect 17344 5286 17400 5288
rect 17448 5340 17504 5342
rect 17448 5288 17450 5340
rect 17450 5288 17502 5340
rect 17502 5288 17504 5340
rect 17448 5286 17504 5288
rect 24130 5390 24186 5446
rect 24234 5390 24290 5446
rect 24130 5286 24186 5342
rect 24234 5286 24290 5342
rect 14222 4410 14278 4466
rect 14326 4410 14382 4466
rect 14430 4410 14486 4466
rect 14222 4306 14278 4362
rect 14326 4306 14382 4362
rect 14430 4306 14486 4362
rect 14222 4202 14278 4258
rect 14326 4202 14382 4258
rect 14430 4202 14486 4258
rect 13110 2294 13166 2296
rect 13110 2242 13112 2294
rect 13112 2242 13164 2294
rect 13164 2242 13166 2294
rect 13110 2240 13166 2242
rect 13110 2190 13166 2192
rect 13110 2138 13112 2190
rect 13112 2138 13164 2190
rect 13164 2138 13166 2190
rect 13110 2136 13166 2138
rect 13110 2086 13166 2088
rect 13110 2034 13112 2086
rect 13112 2034 13164 2086
rect 13164 2034 13166 2086
rect 13110 2032 13166 2034
rect 15062 3562 15118 3564
rect 15062 3510 15064 3562
rect 15064 3510 15116 3562
rect 15116 3510 15118 3562
rect 15062 3508 15118 3510
rect 15062 3458 15118 3460
rect 15062 3406 15064 3458
rect 15064 3406 15116 3458
rect 15116 3406 15118 3458
rect 15062 3404 15118 3406
rect 15670 3562 15726 3564
rect 15670 3510 15672 3562
rect 15672 3510 15724 3562
rect 15724 3510 15726 3562
rect 15670 3508 15726 3510
rect 15670 3458 15726 3460
rect 15670 3406 15672 3458
rect 15672 3406 15724 3458
rect 15724 3406 15726 3458
rect 15670 3404 15726 3406
rect 16278 3562 16334 3564
rect 16278 3510 16280 3562
rect 16280 3510 16332 3562
rect 16332 3510 16334 3562
rect 16278 3508 16334 3510
rect 16278 3458 16334 3460
rect 16278 3406 16280 3458
rect 16280 3406 16332 3458
rect 16332 3406 16334 3458
rect 16278 3404 16334 3406
rect 15566 3108 15622 3164
rect 15670 3108 15726 3164
rect 15774 3108 15830 3164
rect 15566 3004 15622 3060
rect 15670 3004 15726 3060
rect 15774 3004 15830 3060
rect 15566 2900 15622 2956
rect 15670 2900 15726 2956
rect 15774 2900 15830 2956
rect 14899 2240 14955 2296
rect 15003 2240 15059 2296
rect 15107 2240 15163 2296
rect 14899 2136 14955 2192
rect 15003 2136 15059 2192
rect 15107 2136 15163 2192
rect 14899 2032 14955 2088
rect 15003 2032 15059 2088
rect 15107 2032 15163 2088
rect 12028 1127 12084 1129
rect 12028 1075 12030 1127
rect 12030 1075 12082 1127
rect 12082 1075 12084 1127
rect 12028 1073 12084 1075
rect 12132 1127 12188 1129
rect 12132 1075 12134 1127
rect 12134 1075 12186 1127
rect 12186 1075 12188 1127
rect 12132 1073 12188 1075
rect 12028 1023 12084 1025
rect 12028 971 12030 1023
rect 12030 971 12082 1023
rect 12082 971 12084 1023
rect 12028 969 12084 971
rect 12132 1023 12188 1025
rect 12132 971 12134 1023
rect 12134 971 12186 1023
rect 12186 971 12188 1023
rect 12132 969 12188 971
rect 5630 821 5686 877
rect 5734 821 5790 877
rect 5630 717 5686 773
rect 5734 717 5790 773
rect 10323 821 10379 877
rect 10427 821 10483 877
rect 10323 717 10379 773
rect 10427 717 10483 773
rect 5154 501 5210 557
rect 5258 501 5314 557
rect 5154 397 5210 453
rect 5258 397 5314 453
rect 13210 501 13266 557
rect 13314 501 13370 557
rect 14899 718 14955 774
rect 15003 718 15059 774
rect 15107 718 15163 774
rect 14899 614 14955 670
rect 15003 614 15059 670
rect 15107 614 15163 670
rect 14899 510 14955 566
rect 15003 510 15059 566
rect 15107 510 15163 566
rect 21670 4464 21726 4466
rect 21670 4412 21672 4464
rect 21672 4412 21724 4464
rect 21724 4412 21726 4464
rect 21670 4410 21726 4412
rect 21670 4360 21726 4362
rect 21670 4308 21672 4360
rect 21672 4308 21724 4360
rect 21724 4308 21726 4360
rect 21670 4306 21726 4308
rect 21670 4256 21726 4258
rect 21670 4204 21672 4256
rect 21672 4204 21724 4256
rect 21724 4204 21726 4256
rect 21670 4202 21726 4204
rect 20580 3108 20636 3164
rect 20684 3108 20740 3164
rect 20788 3108 20844 3164
rect 20580 3004 20636 3060
rect 20684 3004 20740 3060
rect 20788 3004 20844 3060
rect 20580 2900 20636 2956
rect 20684 2900 20740 2956
rect 20788 2900 20844 2956
rect 30298 4137 30354 4139
rect 30298 4085 30300 4137
rect 30300 4085 30352 4137
rect 30352 4085 30354 4137
rect 30298 4083 30354 4085
rect 30402 4137 30458 4139
rect 30402 4085 30404 4137
rect 30404 4085 30456 4137
rect 30456 4085 30458 4137
rect 30402 4083 30458 4085
rect 30506 4137 30562 4139
rect 30506 4085 30508 4137
rect 30508 4085 30560 4137
rect 30560 4085 30562 4137
rect 30506 4083 30562 4085
rect 30610 4137 30666 4139
rect 30610 4085 30612 4137
rect 30612 4085 30664 4137
rect 30664 4085 30666 4137
rect 30610 4083 30666 4085
rect 30714 4137 30770 4139
rect 30714 4085 30716 4137
rect 30716 4085 30768 4137
rect 30768 4085 30770 4137
rect 30714 4083 30770 4085
rect 30298 4033 30354 4035
rect 30298 3981 30300 4033
rect 30300 3981 30352 4033
rect 30352 3981 30354 4033
rect 30298 3979 30354 3981
rect 30402 4033 30458 4035
rect 30402 3981 30404 4033
rect 30404 3981 30456 4033
rect 30456 3981 30458 4033
rect 30402 3979 30458 3981
rect 30506 4033 30562 4035
rect 30506 3981 30508 4033
rect 30508 3981 30560 4033
rect 30560 3981 30562 4033
rect 30506 3979 30562 3981
rect 30610 4033 30666 4035
rect 30610 3981 30612 4033
rect 30612 3981 30664 4033
rect 30664 3981 30666 4033
rect 30610 3979 30666 3981
rect 30714 4033 30770 4035
rect 30714 3981 30716 4033
rect 30716 3981 30768 4033
rect 30768 3981 30770 4033
rect 30714 3979 30770 3981
rect 30298 3929 30354 3931
rect 30298 3877 30300 3929
rect 30300 3877 30352 3929
rect 30352 3877 30354 3929
rect 30298 3875 30354 3877
rect 30402 3929 30458 3931
rect 30402 3877 30404 3929
rect 30404 3877 30456 3929
rect 30456 3877 30458 3929
rect 30402 3875 30458 3877
rect 30506 3929 30562 3931
rect 30506 3877 30508 3929
rect 30508 3877 30560 3929
rect 30560 3877 30562 3929
rect 30506 3875 30562 3877
rect 30610 3929 30666 3931
rect 30610 3877 30612 3929
rect 30612 3877 30664 3929
rect 30664 3877 30666 3929
rect 30610 3875 30666 3877
rect 30714 3929 30770 3931
rect 30714 3877 30716 3929
rect 30716 3877 30768 3929
rect 30768 3877 30770 3929
rect 30714 3875 30770 3877
rect 30298 3825 30354 3827
rect 30298 3773 30300 3825
rect 30300 3773 30352 3825
rect 30352 3773 30354 3825
rect 30298 3771 30354 3773
rect 30402 3825 30458 3827
rect 30402 3773 30404 3825
rect 30404 3773 30456 3825
rect 30456 3773 30458 3825
rect 30402 3771 30458 3773
rect 30506 3825 30562 3827
rect 30506 3773 30508 3825
rect 30508 3773 30560 3825
rect 30560 3773 30562 3825
rect 30506 3771 30562 3773
rect 30610 3825 30666 3827
rect 30610 3773 30612 3825
rect 30612 3773 30664 3825
rect 30664 3773 30666 3825
rect 30610 3771 30666 3773
rect 30714 3825 30770 3827
rect 30714 3773 30716 3825
rect 30716 3773 30768 3825
rect 30768 3773 30770 3825
rect 30714 3771 30770 3773
rect 30298 3721 30354 3723
rect 30298 3669 30300 3721
rect 30300 3669 30352 3721
rect 30352 3669 30354 3721
rect 30298 3667 30354 3669
rect 30402 3721 30458 3723
rect 30402 3669 30404 3721
rect 30404 3669 30456 3721
rect 30456 3669 30458 3721
rect 30402 3667 30458 3669
rect 30506 3721 30562 3723
rect 30506 3669 30508 3721
rect 30508 3669 30560 3721
rect 30560 3669 30562 3721
rect 30506 3667 30562 3669
rect 30610 3721 30666 3723
rect 30610 3669 30612 3721
rect 30612 3669 30664 3721
rect 30664 3669 30666 3721
rect 30610 3667 30666 3669
rect 30714 3721 30770 3723
rect 30714 3669 30716 3721
rect 30716 3669 30768 3721
rect 30768 3669 30770 3721
rect 30714 3667 30770 3669
rect 15566 2240 15622 2296
rect 15670 2294 15726 2296
rect 15670 2242 15672 2294
rect 15672 2242 15724 2294
rect 15724 2242 15726 2294
rect 15670 2240 15726 2242
rect 15774 2240 15830 2296
rect 15566 2136 15622 2192
rect 15670 2190 15726 2192
rect 15670 2138 15672 2190
rect 15672 2138 15724 2190
rect 15724 2138 15726 2190
rect 15670 2136 15726 2138
rect 15774 2136 15830 2192
rect 15566 2032 15622 2088
rect 15670 2086 15726 2088
rect 15670 2034 15672 2086
rect 15672 2034 15724 2086
rect 15724 2034 15726 2086
rect 15670 2032 15726 2034
rect 15774 2032 15830 2088
rect 13210 397 13266 453
rect 13314 397 13370 453
rect 16181 2202 16237 2258
rect 16285 2202 16341 2258
rect 16389 2202 16445 2258
rect 16181 2098 16237 2154
rect 16285 2098 16341 2154
rect 16389 2098 16445 2154
rect 16181 1994 16237 2050
rect 16285 1994 16341 2050
rect 16389 1994 16445 2050
rect 19110 2256 19166 2258
rect 19110 2204 19112 2256
rect 19112 2204 19164 2256
rect 19164 2204 19166 2256
rect 19110 2202 19166 2204
rect 19110 2152 19166 2154
rect 19110 2100 19112 2152
rect 19112 2100 19164 2152
rect 19164 2100 19166 2152
rect 19110 2098 19166 2100
rect 19110 2048 19166 2050
rect 19110 1996 19112 2048
rect 19112 1996 19164 2048
rect 19164 1996 19166 2048
rect 19110 1994 19166 1996
rect 19430 2256 19486 2258
rect 19430 2204 19432 2256
rect 19432 2204 19484 2256
rect 19484 2204 19486 2256
rect 19430 2202 19486 2204
rect 19430 2152 19486 2154
rect 19430 2100 19432 2152
rect 19432 2100 19484 2152
rect 19484 2100 19486 2152
rect 19430 2098 19486 2100
rect 19430 2048 19486 2050
rect 19430 1996 19432 2048
rect 19432 1996 19484 2048
rect 19484 1996 19486 2048
rect 19430 1994 19486 1996
rect 19750 2256 19806 2258
rect 19750 2204 19752 2256
rect 19752 2204 19804 2256
rect 19804 2204 19806 2256
rect 19750 2202 19806 2204
rect 19750 2152 19806 2154
rect 19750 2100 19752 2152
rect 19752 2100 19804 2152
rect 19804 2100 19806 2152
rect 19750 2098 19806 2100
rect 19750 2048 19806 2050
rect 19750 1996 19752 2048
rect 19752 1996 19804 2048
rect 19804 1996 19806 2048
rect 19750 1994 19806 1996
rect 20070 2256 20126 2258
rect 20070 2204 20072 2256
rect 20072 2204 20124 2256
rect 20124 2204 20126 2256
rect 20070 2202 20126 2204
rect 20070 2152 20126 2154
rect 20070 2100 20072 2152
rect 20072 2100 20124 2152
rect 20124 2100 20126 2152
rect 20070 2098 20126 2100
rect 20070 2048 20126 2050
rect 20070 1996 20072 2048
rect 20072 1996 20124 2048
rect 20124 1996 20126 2048
rect 20070 1994 20126 1996
rect 20390 2256 20446 2258
rect 20390 2204 20392 2256
rect 20392 2204 20444 2256
rect 20444 2204 20446 2256
rect 20390 2202 20446 2204
rect 20390 2152 20446 2154
rect 20390 2100 20392 2152
rect 20392 2100 20444 2152
rect 20444 2100 20446 2152
rect 20390 2098 20446 2100
rect 20390 2048 20446 2050
rect 20390 1996 20392 2048
rect 20392 1996 20444 2048
rect 20444 1996 20446 2048
rect 20390 1994 20446 1996
rect 20710 2256 20766 2258
rect 20710 2204 20712 2256
rect 20712 2204 20764 2256
rect 20764 2204 20766 2256
rect 20710 2202 20766 2204
rect 20710 2152 20766 2154
rect 20710 2100 20712 2152
rect 20712 2100 20764 2152
rect 20764 2100 20766 2152
rect 20710 2098 20766 2100
rect 20710 2048 20766 2050
rect 20710 1996 20712 2048
rect 20712 1996 20764 2048
rect 20764 1996 20766 2048
rect 20710 1994 20766 1996
rect 21030 2256 21086 2258
rect 21030 2204 21032 2256
rect 21032 2204 21084 2256
rect 21084 2204 21086 2256
rect 21030 2202 21086 2204
rect 21030 2152 21086 2154
rect 21030 2100 21032 2152
rect 21032 2100 21084 2152
rect 21084 2100 21086 2152
rect 21030 2098 21086 2100
rect 21030 2048 21086 2050
rect 21030 1996 21032 2048
rect 21032 1996 21084 2048
rect 21084 1996 21086 2048
rect 21030 1994 21086 1996
rect 30298 2125 30354 2127
rect 30298 2073 30300 2125
rect 30300 2073 30352 2125
rect 30352 2073 30354 2125
rect 30298 2071 30354 2073
rect 30402 2125 30458 2127
rect 30402 2073 30404 2125
rect 30404 2073 30456 2125
rect 30456 2073 30458 2125
rect 30402 2071 30458 2073
rect 30506 2125 30562 2127
rect 30506 2073 30508 2125
rect 30508 2073 30560 2125
rect 30560 2073 30562 2125
rect 30506 2071 30562 2073
rect 30610 2125 30666 2127
rect 30610 2073 30612 2125
rect 30612 2073 30664 2125
rect 30664 2073 30666 2125
rect 30610 2071 30666 2073
rect 30714 2125 30770 2127
rect 30714 2073 30716 2125
rect 30716 2073 30768 2125
rect 30768 2073 30770 2125
rect 30714 2071 30770 2073
rect 30298 2021 30354 2023
rect 30298 1969 30300 2021
rect 30300 1969 30352 2021
rect 30352 1969 30354 2021
rect 30298 1967 30354 1969
rect 30402 2021 30458 2023
rect 30402 1969 30404 2021
rect 30404 1969 30456 2021
rect 30456 1969 30458 2021
rect 30402 1967 30458 1969
rect 30506 2021 30562 2023
rect 30506 1969 30508 2021
rect 30508 1969 30560 2021
rect 30560 1969 30562 2021
rect 30506 1967 30562 1969
rect 30610 2021 30666 2023
rect 30610 1969 30612 2021
rect 30612 1969 30664 2021
rect 30664 1969 30666 2021
rect 30610 1967 30666 1969
rect 30714 2021 30770 2023
rect 30714 1969 30716 2021
rect 30716 1969 30768 2021
rect 30768 1969 30770 2021
rect 30714 1967 30770 1969
rect 30298 1917 30354 1919
rect 30298 1865 30300 1917
rect 30300 1865 30352 1917
rect 30352 1865 30354 1917
rect 30298 1863 30354 1865
rect 30402 1917 30458 1919
rect 30402 1865 30404 1917
rect 30404 1865 30456 1917
rect 30456 1865 30458 1917
rect 30402 1863 30458 1865
rect 30506 1917 30562 1919
rect 30506 1865 30508 1917
rect 30508 1865 30560 1917
rect 30560 1865 30562 1917
rect 30506 1863 30562 1865
rect 30610 1917 30666 1919
rect 30610 1865 30612 1917
rect 30612 1865 30664 1917
rect 30664 1865 30666 1917
rect 30610 1863 30666 1865
rect 30714 1917 30770 1919
rect 30714 1865 30716 1917
rect 30716 1865 30768 1917
rect 30768 1865 30770 1917
rect 30714 1863 30770 1865
rect 21641 772 21697 774
rect 21641 720 21643 772
rect 21643 720 21695 772
rect 21695 720 21697 772
rect 21641 718 21697 720
rect 21745 772 21801 774
rect 21745 720 21747 772
rect 21747 720 21799 772
rect 21799 720 21801 772
rect 21745 718 21801 720
rect 21849 772 21905 774
rect 21849 720 21851 772
rect 21851 720 21903 772
rect 21903 720 21905 772
rect 21849 718 21905 720
rect 21641 668 21697 670
rect 21641 616 21643 668
rect 21643 616 21695 668
rect 21695 616 21697 668
rect 21641 614 21697 616
rect 21745 668 21801 670
rect 21745 616 21747 668
rect 21747 616 21799 668
rect 21799 616 21801 668
rect 21745 614 21801 616
rect 21849 668 21905 670
rect 21849 616 21851 668
rect 21851 616 21903 668
rect 21903 616 21905 668
rect 21849 614 21905 616
rect 21641 564 21697 566
rect 21641 512 21643 564
rect 21643 512 21695 564
rect 21695 512 21697 564
rect 21641 510 21697 512
rect 21745 564 21801 566
rect 21745 512 21747 564
rect 21747 512 21799 564
rect 21799 512 21801 564
rect 21745 510 21801 512
rect 21849 564 21905 566
rect 21849 512 21851 564
rect 21851 512 21903 564
rect 21903 512 21905 564
rect 21849 510 21905 512
rect 24128 731 24184 787
rect 24232 731 24288 787
rect 24128 627 24184 683
rect 24232 627 24288 683
rect 24128 523 24184 579
rect 24232 523 24288 579
rect 30298 1813 30354 1815
rect 30298 1761 30300 1813
rect 30300 1761 30352 1813
rect 30352 1761 30354 1813
rect 30298 1759 30354 1761
rect 30402 1813 30458 1815
rect 30402 1761 30404 1813
rect 30404 1761 30456 1813
rect 30456 1761 30458 1813
rect 30402 1759 30458 1761
rect 30506 1813 30562 1815
rect 30506 1761 30508 1813
rect 30508 1761 30560 1813
rect 30560 1761 30562 1813
rect 30506 1759 30562 1761
rect 30610 1813 30666 1815
rect 30610 1761 30612 1813
rect 30612 1761 30664 1813
rect 30664 1761 30666 1813
rect 30610 1759 30666 1761
rect 30714 1813 30770 1815
rect 30714 1761 30716 1813
rect 30716 1761 30768 1813
rect 30768 1761 30770 1813
rect 30714 1759 30770 1761
rect 30298 1709 30354 1711
rect 30298 1657 30300 1709
rect 30300 1657 30352 1709
rect 30352 1657 30354 1709
rect 30298 1655 30354 1657
rect 30402 1709 30458 1711
rect 30402 1657 30404 1709
rect 30404 1657 30456 1709
rect 30456 1657 30458 1709
rect 30402 1655 30458 1657
rect 30506 1709 30562 1711
rect 30506 1657 30508 1709
rect 30508 1657 30560 1709
rect 30560 1657 30562 1709
rect 30506 1655 30562 1657
rect 30610 1709 30666 1711
rect 30610 1657 30612 1709
rect 30612 1657 30664 1709
rect 30664 1657 30666 1709
rect 30610 1655 30666 1657
rect 30714 1709 30770 1711
rect 30714 1657 30716 1709
rect 30716 1657 30768 1709
rect 30768 1657 30770 1709
rect 30714 1655 30770 1657
rect 31756 11714 31812 11770
rect 31860 11714 31916 11770
rect 31964 11714 32020 11770
rect 31756 11610 31812 11666
rect 31860 11610 31916 11666
rect 31964 11610 32020 11666
rect 31756 11506 31812 11562
rect 31860 11506 31916 11562
rect 31964 11506 32020 11562
rect 31756 10260 31812 10316
rect 31860 10260 31916 10316
rect 31964 10260 32020 10316
rect 31756 10156 31812 10212
rect 31860 10156 31916 10212
rect 31964 10156 32020 10212
rect 31756 10052 31812 10108
rect 31860 10052 31916 10108
rect 31964 10052 32020 10108
rect 31756 9200 31812 9256
rect 31860 9200 31916 9256
rect 31964 9200 32020 9256
rect 31756 9096 31812 9152
rect 31860 9096 31916 9152
rect 31964 9096 32020 9152
rect 31756 8992 31812 9048
rect 31860 8992 31916 9048
rect 31964 8992 32020 9048
rect 31756 8534 31812 8590
rect 31860 8534 31916 8590
rect 31964 8534 32020 8590
rect 31756 8430 31812 8486
rect 31860 8430 31916 8486
rect 31964 8430 32020 8486
rect 31756 8326 31812 8382
rect 31860 8326 31916 8382
rect 31964 8326 32020 8382
rect 33733 11664 33789 11666
rect 33733 11612 33735 11664
rect 33735 11612 33787 11664
rect 33787 11612 33789 11664
rect 33733 11610 33789 11612
rect 33733 11560 33789 11562
rect 33733 11508 33735 11560
rect 33735 11508 33787 11560
rect 33787 11508 33789 11560
rect 33733 11506 33789 11508
rect 34373 11664 34429 11666
rect 34373 11612 34375 11664
rect 34375 11612 34427 11664
rect 34427 11612 34429 11664
rect 34373 11610 34429 11612
rect 34373 11560 34429 11562
rect 34373 11508 34375 11560
rect 34375 11508 34427 11560
rect 34427 11508 34429 11560
rect 34373 11506 34429 11508
rect 32136 11320 32192 11376
rect 32240 11320 32296 11376
rect 32344 11320 32400 11376
rect 32136 11216 32192 11272
rect 32240 11216 32296 11272
rect 32344 11216 32400 11272
rect 32136 11112 32192 11168
rect 32240 11112 32296 11168
rect 32344 11112 32400 11168
rect 33412 11270 33468 11272
rect 33412 11218 33414 11270
rect 33414 11218 33466 11270
rect 33466 11218 33468 11270
rect 33412 11216 33468 11218
rect 33412 11166 33468 11168
rect 33412 11114 33414 11166
rect 33414 11114 33466 11166
rect 33466 11114 33468 11166
rect 33412 11112 33468 11114
rect 34052 11270 34108 11272
rect 34052 11218 34054 11270
rect 34054 11218 34106 11270
rect 34106 11218 34108 11270
rect 34052 11216 34108 11218
rect 34052 11166 34108 11168
rect 34052 11114 34054 11166
rect 34054 11114 34106 11166
rect 34106 11114 34108 11166
rect 34052 11112 34108 11114
rect 32136 10654 32192 10710
rect 32240 10654 32296 10710
rect 32344 10654 32400 10710
rect 35013 11664 35069 11666
rect 35013 11612 35015 11664
rect 35015 11612 35067 11664
rect 35067 11612 35069 11664
rect 35013 11610 35069 11612
rect 35013 11560 35069 11562
rect 35013 11508 35015 11560
rect 35015 11508 35067 11560
rect 35067 11508 35069 11560
rect 35013 11506 35069 11508
rect 35653 11664 35709 11666
rect 35653 11612 35655 11664
rect 35655 11612 35707 11664
rect 35707 11612 35709 11664
rect 35653 11610 35709 11612
rect 35653 11560 35709 11562
rect 35653 11508 35655 11560
rect 35655 11508 35707 11560
rect 35707 11508 35709 11560
rect 35653 11506 35709 11508
rect 37867 11664 37923 11666
rect 37867 11612 37869 11664
rect 37869 11612 37921 11664
rect 37921 11612 37923 11664
rect 37867 11610 37923 11612
rect 37867 11560 37923 11562
rect 37867 11508 37869 11560
rect 37869 11508 37921 11560
rect 37921 11508 37923 11560
rect 37867 11506 37923 11508
rect 38507 11664 38563 11666
rect 38507 11612 38509 11664
rect 38509 11612 38561 11664
rect 38561 11612 38563 11664
rect 38507 11610 38563 11612
rect 38507 11560 38563 11562
rect 38507 11508 38509 11560
rect 38509 11508 38561 11560
rect 38561 11508 38563 11560
rect 38507 11506 38563 11508
rect 35332 11270 35388 11272
rect 35332 11218 35334 11270
rect 35334 11218 35386 11270
rect 35386 11218 35388 11270
rect 35332 11216 35388 11218
rect 35332 11166 35388 11168
rect 35332 11114 35334 11166
rect 35334 11114 35386 11166
rect 35386 11114 35388 11166
rect 35332 11112 35388 11114
rect 35972 11270 36028 11272
rect 35972 11218 35974 11270
rect 35974 11218 36026 11270
rect 36026 11218 36028 11270
rect 35972 11216 36028 11218
rect 35972 11166 36028 11168
rect 35972 11114 35974 11166
rect 35974 11114 36026 11166
rect 36026 11114 36028 11166
rect 35972 11112 36028 11114
rect 37548 11270 37604 11272
rect 37548 11218 37550 11270
rect 37550 11218 37602 11270
rect 37602 11218 37604 11270
rect 37548 11216 37604 11218
rect 37548 11166 37604 11168
rect 37548 11114 37550 11166
rect 37550 11114 37602 11166
rect 37602 11114 37604 11166
rect 37548 11112 37604 11114
rect 38188 11270 38244 11272
rect 38188 11218 38190 11270
rect 38190 11218 38242 11270
rect 38242 11218 38244 11270
rect 38188 11216 38244 11218
rect 38188 11166 38244 11168
rect 38188 11114 38190 11166
rect 38190 11114 38242 11166
rect 38242 11114 38244 11166
rect 38188 11112 38244 11114
rect 32136 10550 32192 10606
rect 32240 10550 32296 10606
rect 32344 10550 32400 10606
rect 32136 10446 32192 10502
rect 32240 10446 32296 10502
rect 32344 10446 32400 10502
rect 33733 10604 33789 10606
rect 33733 10552 33735 10604
rect 33735 10552 33787 10604
rect 33787 10552 33789 10604
rect 33733 10550 33789 10552
rect 33733 10500 33789 10502
rect 33733 10448 33735 10500
rect 33735 10448 33787 10500
rect 33787 10448 33789 10500
rect 33733 10446 33789 10448
rect 34373 10604 34429 10606
rect 34373 10552 34375 10604
rect 34375 10552 34427 10604
rect 34427 10552 34429 10604
rect 34373 10550 34429 10552
rect 34373 10500 34429 10502
rect 34373 10448 34375 10500
rect 34375 10448 34427 10500
rect 34427 10448 34429 10500
rect 34373 10446 34429 10448
rect 33412 10210 33468 10212
rect 33412 10158 33414 10210
rect 33414 10158 33466 10210
rect 33466 10158 33468 10210
rect 33412 10156 33468 10158
rect 33412 10106 33468 10108
rect 33412 10054 33414 10106
rect 33414 10054 33466 10106
rect 33466 10054 33468 10106
rect 33412 10052 33468 10054
rect 34052 10210 34108 10212
rect 34052 10158 34054 10210
rect 34054 10158 34106 10210
rect 34106 10158 34108 10210
rect 34052 10156 34108 10158
rect 34052 10106 34108 10108
rect 34052 10054 34054 10106
rect 34054 10054 34106 10106
rect 34106 10054 34108 10106
rect 34052 10052 34108 10054
rect 32136 9594 32192 9650
rect 32240 9594 32296 9650
rect 32344 9594 32400 9650
rect 41483 11714 41539 11770
rect 41587 11714 41643 11770
rect 41691 11714 41747 11770
rect 39147 11664 39203 11666
rect 39147 11612 39149 11664
rect 39149 11612 39201 11664
rect 39201 11612 39203 11664
rect 39147 11610 39203 11612
rect 39147 11560 39203 11562
rect 39147 11508 39149 11560
rect 39149 11508 39201 11560
rect 39201 11508 39203 11560
rect 39147 11506 39203 11508
rect 39787 11664 39843 11666
rect 39787 11612 39789 11664
rect 39789 11612 39841 11664
rect 39841 11612 39843 11664
rect 39787 11610 39843 11612
rect 39787 11560 39843 11562
rect 39787 11508 39789 11560
rect 39789 11508 39841 11560
rect 39841 11508 39843 11560
rect 39787 11506 39843 11508
rect 41483 11610 41539 11666
rect 41587 11610 41643 11666
rect 41691 11610 41747 11666
rect 41483 11506 41539 11562
rect 41587 11506 41643 11562
rect 41691 11506 41747 11562
rect 41122 11320 41178 11376
rect 41226 11320 41282 11376
rect 41330 11320 41386 11376
rect 39468 11270 39524 11272
rect 39468 11218 39470 11270
rect 39470 11218 39522 11270
rect 39522 11218 39524 11270
rect 39468 11216 39524 11218
rect 39468 11166 39524 11168
rect 39468 11114 39470 11166
rect 39470 11114 39522 11166
rect 39522 11114 39524 11166
rect 39468 11112 39524 11114
rect 40108 11270 40164 11272
rect 40108 11218 40110 11270
rect 40110 11218 40162 11270
rect 40162 11218 40164 11270
rect 40108 11216 40164 11218
rect 40108 11166 40164 11168
rect 40108 11114 40110 11166
rect 40110 11114 40162 11166
rect 40162 11114 40164 11166
rect 40108 11112 40164 11114
rect 41122 11216 41178 11272
rect 41226 11216 41282 11272
rect 41330 11216 41386 11272
rect 41122 11112 41178 11168
rect 41226 11112 41282 11168
rect 41330 11112 41386 11168
rect 35013 10604 35069 10606
rect 35013 10552 35015 10604
rect 35015 10552 35067 10604
rect 35067 10552 35069 10604
rect 35013 10550 35069 10552
rect 35013 10500 35069 10502
rect 35013 10448 35015 10500
rect 35015 10448 35067 10500
rect 35067 10448 35069 10500
rect 35013 10446 35069 10448
rect 35653 10604 35709 10606
rect 35653 10552 35655 10604
rect 35655 10552 35707 10604
rect 35707 10552 35709 10604
rect 35653 10550 35709 10552
rect 35653 10500 35709 10502
rect 35653 10448 35655 10500
rect 35655 10448 35707 10500
rect 35707 10448 35709 10500
rect 35653 10446 35709 10448
rect 37867 10604 37923 10606
rect 37867 10552 37869 10604
rect 37869 10552 37921 10604
rect 37921 10552 37923 10604
rect 37867 10550 37923 10552
rect 37867 10500 37923 10502
rect 37867 10448 37869 10500
rect 37869 10448 37921 10500
rect 37921 10448 37923 10500
rect 37867 10446 37923 10448
rect 38507 10604 38563 10606
rect 38507 10552 38509 10604
rect 38509 10552 38561 10604
rect 38561 10552 38563 10604
rect 38507 10550 38563 10552
rect 38507 10500 38563 10502
rect 38507 10448 38509 10500
rect 38509 10448 38561 10500
rect 38561 10448 38563 10500
rect 38507 10446 38563 10448
rect 35332 10210 35388 10212
rect 35332 10158 35334 10210
rect 35334 10158 35386 10210
rect 35386 10158 35388 10210
rect 35332 10156 35388 10158
rect 35332 10106 35388 10108
rect 35332 10054 35334 10106
rect 35334 10054 35386 10106
rect 35386 10054 35388 10106
rect 35332 10052 35388 10054
rect 35972 10210 36028 10212
rect 35972 10158 35974 10210
rect 35974 10158 36026 10210
rect 36026 10158 36028 10210
rect 35972 10156 36028 10158
rect 35972 10106 36028 10108
rect 35972 10054 35974 10106
rect 35974 10054 36026 10106
rect 36026 10054 36028 10106
rect 35972 10052 36028 10054
rect 37548 10210 37604 10212
rect 37548 10158 37550 10210
rect 37550 10158 37602 10210
rect 37602 10158 37604 10210
rect 37548 10156 37604 10158
rect 37548 10106 37604 10108
rect 37548 10054 37550 10106
rect 37550 10054 37602 10106
rect 37602 10054 37604 10106
rect 37548 10052 37604 10054
rect 38188 10210 38244 10212
rect 38188 10158 38190 10210
rect 38190 10158 38242 10210
rect 38242 10158 38244 10210
rect 38188 10156 38244 10158
rect 38188 10106 38244 10108
rect 38188 10054 38190 10106
rect 38190 10054 38242 10106
rect 38242 10054 38244 10106
rect 38188 10052 38244 10054
rect 32136 9490 32192 9546
rect 32240 9490 32296 9546
rect 32344 9490 32400 9546
rect 32136 9386 32192 9442
rect 32240 9386 32296 9442
rect 32344 9386 32400 9442
rect 31228 731 31284 787
rect 31332 731 31388 787
rect 31436 731 31492 787
rect 31228 627 31284 683
rect 31332 627 31388 683
rect 31436 627 31492 683
rect 31228 523 31284 579
rect 31332 523 31388 579
rect 31436 523 31492 579
rect 33733 9544 33789 9546
rect 33733 9492 33735 9544
rect 33735 9492 33787 9544
rect 33787 9492 33789 9544
rect 33733 9490 33789 9492
rect 33733 9440 33789 9442
rect 33733 9388 33735 9440
rect 33735 9388 33787 9440
rect 33787 9388 33789 9440
rect 33733 9386 33789 9388
rect 34373 9544 34429 9546
rect 34373 9492 34375 9544
rect 34375 9492 34427 9544
rect 34427 9492 34429 9544
rect 34373 9490 34429 9492
rect 34373 9440 34429 9442
rect 34373 9388 34375 9440
rect 34375 9388 34427 9440
rect 34427 9388 34429 9440
rect 34373 9386 34429 9388
rect 33412 9150 33468 9152
rect 33412 9098 33414 9150
rect 33414 9098 33466 9150
rect 33466 9098 33468 9150
rect 33412 9096 33468 9098
rect 33412 9046 33468 9048
rect 33412 8994 33414 9046
rect 33414 8994 33466 9046
rect 33466 8994 33468 9046
rect 33412 8992 33468 8994
rect 34052 9150 34108 9152
rect 34052 9098 34054 9150
rect 34054 9098 34106 9150
rect 34106 9098 34108 9150
rect 34052 9096 34108 9098
rect 34052 9046 34108 9048
rect 34052 8994 34054 9046
rect 34054 8994 34106 9046
rect 34106 8994 34108 9046
rect 34052 8992 34108 8994
rect 41122 10654 41178 10710
rect 41226 10654 41282 10710
rect 41330 10654 41386 10710
rect 39147 10604 39203 10606
rect 39147 10552 39149 10604
rect 39149 10552 39201 10604
rect 39201 10552 39203 10604
rect 39147 10550 39203 10552
rect 39147 10500 39203 10502
rect 39147 10448 39149 10500
rect 39149 10448 39201 10500
rect 39201 10448 39203 10500
rect 39147 10446 39203 10448
rect 39787 10604 39843 10606
rect 39787 10552 39789 10604
rect 39789 10552 39841 10604
rect 39841 10552 39843 10604
rect 39787 10550 39843 10552
rect 39787 10500 39843 10502
rect 39787 10448 39789 10500
rect 39789 10448 39841 10500
rect 39841 10448 39843 10500
rect 39787 10446 39843 10448
rect 41122 10550 41178 10606
rect 41226 10550 41282 10606
rect 41330 10550 41386 10606
rect 41122 10446 41178 10502
rect 41226 10446 41282 10502
rect 41330 10446 41386 10502
rect 39468 10210 39524 10212
rect 39468 10158 39470 10210
rect 39470 10158 39522 10210
rect 39522 10158 39524 10210
rect 39468 10156 39524 10158
rect 39468 10106 39524 10108
rect 39468 10054 39470 10106
rect 39470 10054 39522 10106
rect 39522 10054 39524 10106
rect 39468 10052 39524 10054
rect 40108 10210 40164 10212
rect 40108 10158 40110 10210
rect 40110 10158 40162 10210
rect 40162 10158 40164 10210
rect 40108 10156 40164 10158
rect 40108 10106 40164 10108
rect 40108 10054 40110 10106
rect 40110 10054 40162 10106
rect 40162 10054 40164 10106
rect 40108 10052 40164 10054
rect 35013 9544 35069 9546
rect 35013 9492 35015 9544
rect 35015 9492 35067 9544
rect 35067 9492 35069 9544
rect 35013 9490 35069 9492
rect 35013 9440 35069 9442
rect 35013 9388 35015 9440
rect 35015 9388 35067 9440
rect 35067 9388 35069 9440
rect 35013 9386 35069 9388
rect 35653 9544 35709 9546
rect 35653 9492 35655 9544
rect 35655 9492 35707 9544
rect 35707 9492 35709 9544
rect 35653 9490 35709 9492
rect 35653 9440 35709 9442
rect 35653 9388 35655 9440
rect 35655 9388 35707 9440
rect 35707 9388 35709 9440
rect 35653 9386 35709 9388
rect 37867 9544 37923 9546
rect 37867 9492 37869 9544
rect 37869 9492 37921 9544
rect 37921 9492 37923 9544
rect 37867 9490 37923 9492
rect 37867 9440 37923 9442
rect 37867 9388 37869 9440
rect 37869 9388 37921 9440
rect 37921 9388 37923 9440
rect 37867 9386 37923 9388
rect 38507 9544 38563 9546
rect 38507 9492 38509 9544
rect 38509 9492 38561 9544
rect 38561 9492 38563 9544
rect 38507 9490 38563 9492
rect 38507 9440 38563 9442
rect 38507 9388 38509 9440
rect 38509 9388 38561 9440
rect 38561 9388 38563 9440
rect 38507 9386 38563 9388
rect 35332 9150 35388 9152
rect 35332 9098 35334 9150
rect 35334 9098 35386 9150
rect 35386 9098 35388 9150
rect 35332 9096 35388 9098
rect 35332 9046 35388 9048
rect 35332 8994 35334 9046
rect 35334 8994 35386 9046
rect 35386 8994 35388 9046
rect 35332 8992 35388 8994
rect 35972 9150 36028 9152
rect 35972 9098 35974 9150
rect 35974 9098 36026 9150
rect 36026 9098 36028 9150
rect 35972 9096 36028 9098
rect 35972 9046 36028 9048
rect 35972 8994 35974 9046
rect 35974 8994 36026 9046
rect 36026 8994 36028 9046
rect 35972 8992 36028 8994
rect 37548 9150 37604 9152
rect 37548 9098 37550 9150
rect 37550 9098 37602 9150
rect 37602 9098 37604 9150
rect 37548 9096 37604 9098
rect 37548 9046 37604 9048
rect 37548 8994 37550 9046
rect 37550 8994 37602 9046
rect 37602 8994 37604 9046
rect 37548 8992 37604 8994
rect 38188 9150 38244 9152
rect 38188 9098 38190 9150
rect 38190 9098 38242 9150
rect 38242 9098 38244 9150
rect 38188 9096 38244 9098
rect 38188 9046 38244 9048
rect 38188 8994 38190 9046
rect 38190 8994 38242 9046
rect 38242 8994 38244 9046
rect 38188 8992 38244 8994
rect 33733 8484 33789 8486
rect 33733 8432 33735 8484
rect 33735 8432 33787 8484
rect 33787 8432 33789 8484
rect 33733 8430 33789 8432
rect 33733 8380 33789 8382
rect 33733 8328 33735 8380
rect 33735 8328 33787 8380
rect 33787 8328 33789 8380
rect 33733 8326 33789 8328
rect 34373 8484 34429 8486
rect 34373 8432 34375 8484
rect 34375 8432 34427 8484
rect 34427 8432 34429 8484
rect 34373 8430 34429 8432
rect 34373 8380 34429 8382
rect 34373 8328 34375 8380
rect 34375 8328 34427 8380
rect 34427 8328 34429 8380
rect 34373 8326 34429 8328
rect 32136 8140 32192 8196
rect 32240 8140 32296 8196
rect 32344 8140 32400 8196
rect 32136 8036 32192 8092
rect 32240 8036 32296 8092
rect 32344 8036 32400 8092
rect 32136 7932 32192 7988
rect 32240 7932 32296 7988
rect 32344 7932 32400 7988
rect 24578 330 24634 386
rect 24682 330 24738 386
rect 24578 226 24634 282
rect 24682 226 24738 282
rect 24578 122 24634 178
rect 24682 122 24738 178
rect 33412 8090 33468 8092
rect 33412 8038 33414 8090
rect 33414 8038 33466 8090
rect 33466 8038 33468 8090
rect 33412 8036 33468 8038
rect 33412 7986 33468 7988
rect 33412 7934 33414 7986
rect 33414 7934 33466 7986
rect 33466 7934 33468 7986
rect 33412 7932 33468 7934
rect 34052 8090 34108 8092
rect 34052 8038 34054 8090
rect 34054 8038 34106 8090
rect 34106 8038 34108 8090
rect 34052 8036 34108 8038
rect 34052 7986 34108 7988
rect 34052 7934 34054 7986
rect 34054 7934 34106 7986
rect 34106 7934 34108 7986
rect 34052 7932 34108 7934
rect 41122 9594 41178 9650
rect 41226 9594 41282 9650
rect 41330 9594 41386 9650
rect 39147 9544 39203 9546
rect 39147 9492 39149 9544
rect 39149 9492 39201 9544
rect 39201 9492 39203 9544
rect 39147 9490 39203 9492
rect 39147 9440 39203 9442
rect 39147 9388 39149 9440
rect 39149 9388 39201 9440
rect 39201 9388 39203 9440
rect 39147 9386 39203 9388
rect 39787 9544 39843 9546
rect 39787 9492 39789 9544
rect 39789 9492 39841 9544
rect 39841 9492 39843 9544
rect 39787 9490 39843 9492
rect 39787 9440 39843 9442
rect 39787 9388 39789 9440
rect 39789 9388 39841 9440
rect 39841 9388 39843 9440
rect 39787 9386 39843 9388
rect 41122 9490 41178 9546
rect 41226 9490 41282 9546
rect 41330 9490 41386 9546
rect 41122 9386 41178 9442
rect 41226 9386 41282 9442
rect 41330 9386 41386 9442
rect 39468 9150 39524 9152
rect 39468 9098 39470 9150
rect 39470 9098 39522 9150
rect 39522 9098 39524 9150
rect 39468 9096 39524 9098
rect 39468 9046 39524 9048
rect 39468 8994 39470 9046
rect 39470 8994 39522 9046
rect 39522 8994 39524 9046
rect 39468 8992 39524 8994
rect 40108 9150 40164 9152
rect 40108 9098 40110 9150
rect 40110 9098 40162 9150
rect 40162 9098 40164 9150
rect 40108 9096 40164 9098
rect 40108 9046 40164 9048
rect 40108 8994 40110 9046
rect 40110 8994 40162 9046
rect 40162 8994 40164 9046
rect 40108 8992 40164 8994
rect 35013 8484 35069 8486
rect 35013 8432 35015 8484
rect 35015 8432 35067 8484
rect 35067 8432 35069 8484
rect 35013 8430 35069 8432
rect 35013 8380 35069 8382
rect 35013 8328 35015 8380
rect 35015 8328 35067 8380
rect 35067 8328 35069 8380
rect 35013 8326 35069 8328
rect 35653 8484 35709 8486
rect 35653 8432 35655 8484
rect 35655 8432 35707 8484
rect 35707 8432 35709 8484
rect 35653 8430 35709 8432
rect 35653 8380 35709 8382
rect 35653 8328 35655 8380
rect 35655 8328 35707 8380
rect 35707 8328 35709 8380
rect 35653 8326 35709 8328
rect 37867 8484 37923 8486
rect 37867 8432 37869 8484
rect 37869 8432 37921 8484
rect 37921 8432 37923 8484
rect 37867 8430 37923 8432
rect 37867 8380 37923 8382
rect 37867 8328 37869 8380
rect 37869 8328 37921 8380
rect 37921 8328 37923 8380
rect 37867 8326 37923 8328
rect 38507 8484 38563 8486
rect 38507 8432 38509 8484
rect 38509 8432 38561 8484
rect 38561 8432 38563 8484
rect 38507 8430 38563 8432
rect 38507 8380 38563 8382
rect 38507 8328 38509 8380
rect 38509 8328 38561 8380
rect 38561 8328 38563 8380
rect 38507 8326 38563 8328
rect 39147 8484 39203 8486
rect 39147 8432 39149 8484
rect 39149 8432 39201 8484
rect 39201 8432 39203 8484
rect 39147 8430 39203 8432
rect 39147 8380 39203 8382
rect 39147 8328 39149 8380
rect 39149 8328 39201 8380
rect 39201 8328 39203 8380
rect 39147 8326 39203 8328
rect 39787 8484 39843 8486
rect 39787 8432 39789 8484
rect 39789 8432 39841 8484
rect 39841 8432 39843 8484
rect 39787 8430 39843 8432
rect 39787 8380 39843 8382
rect 39787 8328 39789 8380
rect 39789 8328 39841 8380
rect 39841 8328 39843 8380
rect 39787 8326 39843 8328
rect 43429 11664 43485 11666
rect 43429 11612 43431 11664
rect 43431 11612 43483 11664
rect 43483 11612 43485 11664
rect 43429 11610 43485 11612
rect 43429 11560 43485 11562
rect 43429 11508 43431 11560
rect 43431 11508 43483 11560
rect 43483 11508 43485 11560
rect 43429 11506 43485 11508
rect 44069 11664 44125 11666
rect 44069 11612 44071 11664
rect 44071 11612 44123 11664
rect 44123 11612 44125 11664
rect 44069 11610 44125 11612
rect 44069 11560 44125 11562
rect 44069 11508 44071 11560
rect 44071 11508 44123 11560
rect 44123 11508 44125 11560
rect 44069 11506 44125 11508
rect 41483 10260 41539 10316
rect 41587 10260 41643 10316
rect 41691 10260 41747 10316
rect 41483 10156 41539 10212
rect 41587 10156 41643 10212
rect 41691 10156 41747 10212
rect 41483 10052 41539 10108
rect 41587 10052 41643 10108
rect 41691 10052 41747 10108
rect 41483 9200 41539 9256
rect 41587 9200 41643 9256
rect 41691 9200 41747 9256
rect 41483 9096 41539 9152
rect 41587 9096 41643 9152
rect 41691 9096 41747 9152
rect 41483 8992 41539 9048
rect 41587 8992 41643 9048
rect 41691 8992 41747 9048
rect 41483 8534 41539 8590
rect 41587 8534 41643 8590
rect 41691 8534 41747 8590
rect 41483 8430 41539 8486
rect 41587 8430 41643 8486
rect 41691 8430 41747 8486
rect 41483 8326 41539 8382
rect 41587 8326 41643 8382
rect 41691 8326 41747 8382
rect 41842 11320 41898 11376
rect 41946 11320 42002 11376
rect 42050 11320 42106 11376
rect 41842 11216 41898 11272
rect 41946 11216 42002 11272
rect 42050 11216 42106 11272
rect 41842 11112 41898 11168
rect 41946 11112 42002 11168
rect 42050 11112 42106 11168
rect 43108 11270 43164 11272
rect 43108 11218 43110 11270
rect 43110 11218 43162 11270
rect 43162 11218 43164 11270
rect 43108 11216 43164 11218
rect 43108 11166 43164 11168
rect 43108 11114 43110 11166
rect 43110 11114 43162 11166
rect 43162 11114 43164 11166
rect 43108 11112 43164 11114
rect 43748 11270 43804 11272
rect 43748 11218 43750 11270
rect 43750 11218 43802 11270
rect 43802 11218 43804 11270
rect 43748 11216 43804 11218
rect 43748 11166 43804 11168
rect 43748 11114 43750 11166
rect 43750 11114 43802 11166
rect 43802 11114 43804 11166
rect 43748 11112 43804 11114
rect 41842 10654 41898 10710
rect 41946 10654 42002 10710
rect 42050 10654 42106 10710
rect 44709 11664 44765 11666
rect 44709 11612 44711 11664
rect 44711 11612 44763 11664
rect 44763 11612 44765 11664
rect 44709 11610 44765 11612
rect 44709 11560 44765 11562
rect 44709 11508 44711 11560
rect 44711 11508 44763 11560
rect 44763 11508 44765 11560
rect 44709 11506 44765 11508
rect 45349 11664 45405 11666
rect 45349 11612 45351 11664
rect 45351 11612 45403 11664
rect 45403 11612 45405 11664
rect 45349 11610 45405 11612
rect 45349 11560 45405 11562
rect 45349 11508 45351 11560
rect 45351 11508 45403 11560
rect 45403 11508 45405 11560
rect 45349 11506 45405 11508
rect 47563 11664 47619 11666
rect 47563 11612 47565 11664
rect 47565 11612 47617 11664
rect 47617 11612 47619 11664
rect 47563 11610 47619 11612
rect 47563 11560 47619 11562
rect 47563 11508 47565 11560
rect 47565 11508 47617 11560
rect 47617 11508 47619 11560
rect 47563 11506 47619 11508
rect 48203 11664 48259 11666
rect 48203 11612 48205 11664
rect 48205 11612 48257 11664
rect 48257 11612 48259 11664
rect 48203 11610 48259 11612
rect 48203 11560 48259 11562
rect 48203 11508 48205 11560
rect 48205 11508 48257 11560
rect 48257 11508 48259 11560
rect 48203 11506 48259 11508
rect 45028 11270 45084 11272
rect 45028 11218 45030 11270
rect 45030 11218 45082 11270
rect 45082 11218 45084 11270
rect 45028 11216 45084 11218
rect 45028 11166 45084 11168
rect 45028 11114 45030 11166
rect 45030 11114 45082 11166
rect 45082 11114 45084 11166
rect 45028 11112 45084 11114
rect 45668 11270 45724 11272
rect 45668 11218 45670 11270
rect 45670 11218 45722 11270
rect 45722 11218 45724 11270
rect 45668 11216 45724 11218
rect 45668 11166 45724 11168
rect 45668 11114 45670 11166
rect 45670 11114 45722 11166
rect 45722 11114 45724 11166
rect 45668 11112 45724 11114
rect 47244 11270 47300 11272
rect 47244 11218 47246 11270
rect 47246 11218 47298 11270
rect 47298 11218 47300 11270
rect 47244 11216 47300 11218
rect 47244 11166 47300 11168
rect 47244 11114 47246 11166
rect 47246 11114 47298 11166
rect 47298 11114 47300 11166
rect 47244 11112 47300 11114
rect 47884 11270 47940 11272
rect 47884 11218 47886 11270
rect 47886 11218 47938 11270
rect 47938 11218 47940 11270
rect 47884 11216 47940 11218
rect 47884 11166 47940 11168
rect 47884 11114 47886 11166
rect 47886 11114 47938 11166
rect 47938 11114 47940 11166
rect 47884 11112 47940 11114
rect 41842 10550 41898 10606
rect 41946 10550 42002 10606
rect 42050 10550 42106 10606
rect 41842 10446 41898 10502
rect 41946 10446 42002 10502
rect 42050 10446 42106 10502
rect 43429 10604 43485 10606
rect 43429 10552 43431 10604
rect 43431 10552 43483 10604
rect 43483 10552 43485 10604
rect 43429 10550 43485 10552
rect 43429 10500 43485 10502
rect 43429 10448 43431 10500
rect 43431 10448 43483 10500
rect 43483 10448 43485 10500
rect 43429 10446 43485 10448
rect 44069 10604 44125 10606
rect 44069 10552 44071 10604
rect 44071 10552 44123 10604
rect 44123 10552 44125 10604
rect 44069 10550 44125 10552
rect 44069 10500 44125 10502
rect 44069 10448 44071 10500
rect 44071 10448 44123 10500
rect 44123 10448 44125 10500
rect 44069 10446 44125 10448
rect 43108 10210 43164 10212
rect 43108 10158 43110 10210
rect 43110 10158 43162 10210
rect 43162 10158 43164 10210
rect 43108 10156 43164 10158
rect 43108 10106 43164 10108
rect 43108 10054 43110 10106
rect 43110 10054 43162 10106
rect 43162 10054 43164 10106
rect 43108 10052 43164 10054
rect 43748 10210 43804 10212
rect 43748 10158 43750 10210
rect 43750 10158 43802 10210
rect 43802 10158 43804 10210
rect 43748 10156 43804 10158
rect 43748 10106 43804 10108
rect 43748 10054 43750 10106
rect 43750 10054 43802 10106
rect 43802 10054 43804 10106
rect 43748 10052 43804 10054
rect 41842 9594 41898 9650
rect 41946 9594 42002 9650
rect 42050 9594 42106 9650
rect 51138 11714 51194 11770
rect 51242 11714 51298 11770
rect 51346 11714 51402 11770
rect 48843 11664 48899 11666
rect 48843 11612 48845 11664
rect 48845 11612 48897 11664
rect 48897 11612 48899 11664
rect 48843 11610 48899 11612
rect 48843 11560 48899 11562
rect 48843 11508 48845 11560
rect 48845 11508 48897 11560
rect 48897 11508 48899 11560
rect 48843 11506 48899 11508
rect 49483 11664 49539 11666
rect 49483 11612 49485 11664
rect 49485 11612 49537 11664
rect 49537 11612 49539 11664
rect 49483 11610 49539 11612
rect 49483 11560 49539 11562
rect 49483 11508 49485 11560
rect 49485 11508 49537 11560
rect 49537 11508 49539 11560
rect 49483 11506 49539 11508
rect 51138 11610 51194 11666
rect 51242 11610 51298 11666
rect 51346 11610 51402 11666
rect 51138 11506 51194 11562
rect 51242 11506 51298 11562
rect 51346 11506 51402 11562
rect 50798 11320 50854 11376
rect 50902 11320 50958 11376
rect 51006 11320 51062 11376
rect 49164 11270 49220 11272
rect 49164 11218 49166 11270
rect 49166 11218 49218 11270
rect 49218 11218 49220 11270
rect 49164 11216 49220 11218
rect 49164 11166 49220 11168
rect 49164 11114 49166 11166
rect 49166 11114 49218 11166
rect 49218 11114 49220 11166
rect 49164 11112 49220 11114
rect 49804 11270 49860 11272
rect 49804 11218 49806 11270
rect 49806 11218 49858 11270
rect 49858 11218 49860 11270
rect 49804 11216 49860 11218
rect 49804 11166 49860 11168
rect 49804 11114 49806 11166
rect 49806 11114 49858 11166
rect 49858 11114 49860 11166
rect 49804 11112 49860 11114
rect 50798 11216 50854 11272
rect 50902 11216 50958 11272
rect 51006 11216 51062 11272
rect 50798 11112 50854 11168
rect 50902 11112 50958 11168
rect 51006 11112 51062 11168
rect 44709 10604 44765 10606
rect 44709 10552 44711 10604
rect 44711 10552 44763 10604
rect 44763 10552 44765 10604
rect 44709 10550 44765 10552
rect 44709 10500 44765 10502
rect 44709 10448 44711 10500
rect 44711 10448 44763 10500
rect 44763 10448 44765 10500
rect 44709 10446 44765 10448
rect 45349 10604 45405 10606
rect 45349 10552 45351 10604
rect 45351 10552 45403 10604
rect 45403 10552 45405 10604
rect 45349 10550 45405 10552
rect 45349 10500 45405 10502
rect 45349 10448 45351 10500
rect 45351 10448 45403 10500
rect 45403 10448 45405 10500
rect 45349 10446 45405 10448
rect 47563 10604 47619 10606
rect 47563 10552 47565 10604
rect 47565 10552 47617 10604
rect 47617 10552 47619 10604
rect 47563 10550 47619 10552
rect 47563 10500 47619 10502
rect 47563 10448 47565 10500
rect 47565 10448 47617 10500
rect 47617 10448 47619 10500
rect 47563 10446 47619 10448
rect 48203 10604 48259 10606
rect 48203 10552 48205 10604
rect 48205 10552 48257 10604
rect 48257 10552 48259 10604
rect 48203 10550 48259 10552
rect 48203 10500 48259 10502
rect 48203 10448 48205 10500
rect 48205 10448 48257 10500
rect 48257 10448 48259 10500
rect 48203 10446 48259 10448
rect 45028 10210 45084 10212
rect 45028 10158 45030 10210
rect 45030 10158 45082 10210
rect 45082 10158 45084 10210
rect 45028 10156 45084 10158
rect 45028 10106 45084 10108
rect 45028 10054 45030 10106
rect 45030 10054 45082 10106
rect 45082 10054 45084 10106
rect 45028 10052 45084 10054
rect 45668 10210 45724 10212
rect 45668 10158 45670 10210
rect 45670 10158 45722 10210
rect 45722 10158 45724 10210
rect 45668 10156 45724 10158
rect 45668 10106 45724 10108
rect 45668 10054 45670 10106
rect 45670 10054 45722 10106
rect 45722 10054 45724 10106
rect 45668 10052 45724 10054
rect 47244 10210 47300 10212
rect 47244 10158 47246 10210
rect 47246 10158 47298 10210
rect 47298 10158 47300 10210
rect 47244 10156 47300 10158
rect 47244 10106 47300 10108
rect 47244 10054 47246 10106
rect 47246 10054 47298 10106
rect 47298 10054 47300 10106
rect 47244 10052 47300 10054
rect 47884 10210 47940 10212
rect 47884 10158 47886 10210
rect 47886 10158 47938 10210
rect 47938 10158 47940 10210
rect 47884 10156 47940 10158
rect 47884 10106 47940 10108
rect 47884 10054 47886 10106
rect 47886 10054 47938 10106
rect 47938 10054 47940 10106
rect 47884 10052 47940 10054
rect 41842 9490 41898 9546
rect 41946 9490 42002 9546
rect 42050 9490 42106 9546
rect 41842 9386 41898 9442
rect 41946 9386 42002 9442
rect 42050 9386 42106 9442
rect 41122 8140 41178 8196
rect 41226 8140 41282 8196
rect 41330 8140 41386 8196
rect 35332 8090 35388 8092
rect 35332 8038 35334 8090
rect 35334 8038 35386 8090
rect 35386 8038 35388 8090
rect 35332 8036 35388 8038
rect 35332 7986 35388 7988
rect 35332 7934 35334 7986
rect 35334 7934 35386 7986
rect 35386 7934 35388 7986
rect 35332 7932 35388 7934
rect 35972 8090 36028 8092
rect 35972 8038 35974 8090
rect 35974 8038 36026 8090
rect 36026 8038 36028 8090
rect 35972 8036 36028 8038
rect 35972 7986 36028 7988
rect 35972 7934 35974 7986
rect 35974 7934 36026 7986
rect 36026 7934 36028 7986
rect 35972 7932 36028 7934
rect 37548 8090 37604 8092
rect 37548 8038 37550 8090
rect 37550 8038 37602 8090
rect 37602 8038 37604 8090
rect 37548 8036 37604 8038
rect 37548 7986 37604 7988
rect 37548 7934 37550 7986
rect 37550 7934 37602 7986
rect 37602 7934 37604 7986
rect 37548 7932 37604 7934
rect 38188 8090 38244 8092
rect 38188 8038 38190 8090
rect 38190 8038 38242 8090
rect 38242 8038 38244 8090
rect 38188 8036 38244 8038
rect 38188 7986 38244 7988
rect 38188 7934 38190 7986
rect 38190 7934 38242 7986
rect 38242 7934 38244 7986
rect 38188 7932 38244 7934
rect 39468 8090 39524 8092
rect 39468 8038 39470 8090
rect 39470 8038 39522 8090
rect 39522 8038 39524 8090
rect 39468 8036 39524 8038
rect 39468 7986 39524 7988
rect 39468 7934 39470 7986
rect 39470 7934 39522 7986
rect 39522 7934 39524 7986
rect 39468 7932 39524 7934
rect 40108 8090 40164 8092
rect 40108 8038 40110 8090
rect 40110 8038 40162 8090
rect 40162 8038 40164 8090
rect 40108 8036 40164 8038
rect 40108 7986 40164 7988
rect 40108 7934 40110 7986
rect 40110 7934 40162 7986
rect 40162 7934 40164 7986
rect 40108 7932 40164 7934
rect 41122 8036 41178 8092
rect 41226 8036 41282 8092
rect 41330 8036 41386 8092
rect 41122 7932 41178 7988
rect 41226 7932 41282 7988
rect 41330 7932 41386 7988
rect 43429 9544 43485 9546
rect 43429 9492 43431 9544
rect 43431 9492 43483 9544
rect 43483 9492 43485 9544
rect 43429 9490 43485 9492
rect 43429 9440 43485 9442
rect 43429 9388 43431 9440
rect 43431 9388 43483 9440
rect 43483 9388 43485 9440
rect 43429 9386 43485 9388
rect 44069 9544 44125 9546
rect 44069 9492 44071 9544
rect 44071 9492 44123 9544
rect 44123 9492 44125 9544
rect 44069 9490 44125 9492
rect 44069 9440 44125 9442
rect 44069 9388 44071 9440
rect 44071 9388 44123 9440
rect 44123 9388 44125 9440
rect 44069 9386 44125 9388
rect 43108 9150 43164 9152
rect 43108 9098 43110 9150
rect 43110 9098 43162 9150
rect 43162 9098 43164 9150
rect 43108 9096 43164 9098
rect 43108 9046 43164 9048
rect 43108 8994 43110 9046
rect 43110 8994 43162 9046
rect 43162 8994 43164 9046
rect 43108 8992 43164 8994
rect 43748 9150 43804 9152
rect 43748 9098 43750 9150
rect 43750 9098 43802 9150
rect 43802 9098 43804 9150
rect 43748 9096 43804 9098
rect 43748 9046 43804 9048
rect 43748 8994 43750 9046
rect 43750 8994 43802 9046
rect 43802 8994 43804 9046
rect 43748 8992 43804 8994
rect 50798 10654 50854 10710
rect 50902 10654 50958 10710
rect 51006 10654 51062 10710
rect 48843 10604 48899 10606
rect 48843 10552 48845 10604
rect 48845 10552 48897 10604
rect 48897 10552 48899 10604
rect 48843 10550 48899 10552
rect 48843 10500 48899 10502
rect 48843 10448 48845 10500
rect 48845 10448 48897 10500
rect 48897 10448 48899 10500
rect 48843 10446 48899 10448
rect 49483 10604 49539 10606
rect 49483 10552 49485 10604
rect 49485 10552 49537 10604
rect 49537 10552 49539 10604
rect 49483 10550 49539 10552
rect 49483 10500 49539 10502
rect 49483 10448 49485 10500
rect 49485 10448 49537 10500
rect 49537 10448 49539 10500
rect 49483 10446 49539 10448
rect 50798 10550 50854 10606
rect 50902 10550 50958 10606
rect 51006 10550 51062 10606
rect 50798 10446 50854 10502
rect 50902 10446 50958 10502
rect 51006 10446 51062 10502
rect 49164 10210 49220 10212
rect 49164 10158 49166 10210
rect 49166 10158 49218 10210
rect 49218 10158 49220 10210
rect 49164 10156 49220 10158
rect 49164 10106 49220 10108
rect 49164 10054 49166 10106
rect 49166 10054 49218 10106
rect 49218 10054 49220 10106
rect 49164 10052 49220 10054
rect 49804 10210 49860 10212
rect 49804 10158 49806 10210
rect 49806 10158 49858 10210
rect 49858 10158 49860 10210
rect 49804 10156 49860 10158
rect 49804 10106 49860 10108
rect 49804 10054 49806 10106
rect 49806 10054 49858 10106
rect 49858 10054 49860 10106
rect 49804 10052 49860 10054
rect 44709 9544 44765 9546
rect 44709 9492 44711 9544
rect 44711 9492 44763 9544
rect 44763 9492 44765 9544
rect 44709 9490 44765 9492
rect 44709 9440 44765 9442
rect 44709 9388 44711 9440
rect 44711 9388 44763 9440
rect 44763 9388 44765 9440
rect 44709 9386 44765 9388
rect 45349 9544 45405 9546
rect 45349 9492 45351 9544
rect 45351 9492 45403 9544
rect 45403 9492 45405 9544
rect 45349 9490 45405 9492
rect 45349 9440 45405 9442
rect 45349 9388 45351 9440
rect 45351 9388 45403 9440
rect 45403 9388 45405 9440
rect 45349 9386 45405 9388
rect 47563 9544 47619 9546
rect 47563 9492 47565 9544
rect 47565 9492 47617 9544
rect 47617 9492 47619 9544
rect 47563 9490 47619 9492
rect 47563 9440 47619 9442
rect 47563 9388 47565 9440
rect 47565 9388 47617 9440
rect 47617 9388 47619 9440
rect 47563 9386 47619 9388
rect 48203 9544 48259 9546
rect 48203 9492 48205 9544
rect 48205 9492 48257 9544
rect 48257 9492 48259 9544
rect 48203 9490 48259 9492
rect 48203 9440 48259 9442
rect 48203 9388 48205 9440
rect 48205 9388 48257 9440
rect 48257 9388 48259 9440
rect 48203 9386 48259 9388
rect 45028 9150 45084 9152
rect 45028 9098 45030 9150
rect 45030 9098 45082 9150
rect 45082 9098 45084 9150
rect 45028 9096 45084 9098
rect 45028 9046 45084 9048
rect 45028 8994 45030 9046
rect 45030 8994 45082 9046
rect 45082 8994 45084 9046
rect 45028 8992 45084 8994
rect 45668 9150 45724 9152
rect 45668 9098 45670 9150
rect 45670 9098 45722 9150
rect 45722 9098 45724 9150
rect 45668 9096 45724 9098
rect 45668 9046 45724 9048
rect 45668 8994 45670 9046
rect 45670 8994 45722 9046
rect 45722 8994 45724 9046
rect 45668 8992 45724 8994
rect 47244 9150 47300 9152
rect 47244 9098 47246 9150
rect 47246 9098 47298 9150
rect 47298 9098 47300 9150
rect 47244 9096 47300 9098
rect 47244 9046 47300 9048
rect 47244 8994 47246 9046
rect 47246 8994 47298 9046
rect 47298 8994 47300 9046
rect 47244 8992 47300 8994
rect 47884 9150 47940 9152
rect 47884 9098 47886 9150
rect 47886 9098 47938 9150
rect 47938 9098 47940 9150
rect 47884 9096 47940 9098
rect 47884 9046 47940 9048
rect 47884 8994 47886 9046
rect 47886 8994 47938 9046
rect 47938 8994 47940 9046
rect 47884 8992 47940 8994
rect 50798 9594 50854 9650
rect 50902 9594 50958 9650
rect 51006 9594 51062 9650
rect 48843 9544 48899 9546
rect 48843 9492 48845 9544
rect 48845 9492 48897 9544
rect 48897 9492 48899 9544
rect 48843 9490 48899 9492
rect 48843 9440 48899 9442
rect 48843 9388 48845 9440
rect 48845 9388 48897 9440
rect 48897 9388 48899 9440
rect 48843 9386 48899 9388
rect 49483 9544 49539 9546
rect 49483 9492 49485 9544
rect 49485 9492 49537 9544
rect 49537 9492 49539 9544
rect 49483 9490 49539 9492
rect 49483 9440 49539 9442
rect 49483 9388 49485 9440
rect 49485 9388 49537 9440
rect 49537 9388 49539 9440
rect 49483 9386 49539 9388
rect 50798 9490 50854 9546
rect 50902 9490 50958 9546
rect 51006 9490 51062 9546
rect 50798 9386 50854 9442
rect 50902 9386 50958 9442
rect 51006 9386 51062 9442
rect 49164 9150 49220 9152
rect 49164 9098 49166 9150
rect 49166 9098 49218 9150
rect 49218 9098 49220 9150
rect 49164 9096 49220 9098
rect 49164 9046 49220 9048
rect 49164 8994 49166 9046
rect 49166 8994 49218 9046
rect 49218 8994 49220 9046
rect 49164 8992 49220 8994
rect 49804 9150 49860 9152
rect 49804 9098 49806 9150
rect 49806 9098 49858 9150
rect 49858 9098 49860 9150
rect 49804 9096 49860 9098
rect 49804 9046 49860 9048
rect 49804 8994 49806 9046
rect 49806 8994 49858 9046
rect 49858 8994 49860 9046
rect 49804 8992 49860 8994
rect 43429 8484 43485 8486
rect 43429 8432 43431 8484
rect 43431 8432 43483 8484
rect 43483 8432 43485 8484
rect 43429 8430 43485 8432
rect 43429 8380 43485 8382
rect 43429 8328 43431 8380
rect 43431 8328 43483 8380
rect 43483 8328 43485 8380
rect 43429 8326 43485 8328
rect 44069 8484 44125 8486
rect 44069 8432 44071 8484
rect 44071 8432 44123 8484
rect 44123 8432 44125 8484
rect 44069 8430 44125 8432
rect 44069 8380 44125 8382
rect 44069 8328 44071 8380
rect 44071 8328 44123 8380
rect 44123 8328 44125 8380
rect 44069 8326 44125 8328
rect 44709 8484 44765 8486
rect 44709 8432 44711 8484
rect 44711 8432 44763 8484
rect 44763 8432 44765 8484
rect 44709 8430 44765 8432
rect 44709 8380 44765 8382
rect 44709 8328 44711 8380
rect 44711 8328 44763 8380
rect 44763 8328 44765 8380
rect 44709 8326 44765 8328
rect 45349 8484 45405 8486
rect 45349 8432 45351 8484
rect 45351 8432 45403 8484
rect 45403 8432 45405 8484
rect 45349 8430 45405 8432
rect 45349 8380 45405 8382
rect 45349 8328 45351 8380
rect 45351 8328 45403 8380
rect 45403 8328 45405 8380
rect 45349 8326 45405 8328
rect 47563 8484 47619 8486
rect 47563 8432 47565 8484
rect 47565 8432 47617 8484
rect 47617 8432 47619 8484
rect 47563 8430 47619 8432
rect 47563 8380 47619 8382
rect 47563 8328 47565 8380
rect 47565 8328 47617 8380
rect 47617 8328 47619 8380
rect 47563 8326 47619 8328
rect 48203 8484 48259 8486
rect 48203 8432 48205 8484
rect 48205 8432 48257 8484
rect 48257 8432 48259 8484
rect 48203 8430 48259 8432
rect 48203 8380 48259 8382
rect 48203 8328 48205 8380
rect 48205 8328 48257 8380
rect 48257 8328 48259 8380
rect 48203 8326 48259 8328
rect 48843 8484 48899 8486
rect 48843 8432 48845 8484
rect 48845 8432 48897 8484
rect 48897 8432 48899 8484
rect 48843 8430 48899 8432
rect 48843 8380 48899 8382
rect 48843 8328 48845 8380
rect 48845 8328 48897 8380
rect 48897 8328 48899 8380
rect 48843 8326 48899 8328
rect 49483 8484 49539 8486
rect 49483 8432 49485 8484
rect 49485 8432 49537 8484
rect 49537 8432 49539 8484
rect 49483 8430 49539 8432
rect 49483 8380 49539 8382
rect 49483 8328 49485 8380
rect 49485 8328 49537 8380
rect 49537 8328 49539 8380
rect 49483 8326 49539 8328
rect 41842 8140 41898 8196
rect 41946 8140 42002 8196
rect 42050 8140 42106 8196
rect 53125 11664 53181 11666
rect 53125 11612 53127 11664
rect 53127 11612 53179 11664
rect 53179 11612 53181 11664
rect 53125 11610 53181 11612
rect 53125 11560 53181 11562
rect 53125 11508 53127 11560
rect 53127 11508 53179 11560
rect 53179 11508 53181 11560
rect 53125 11506 53181 11508
rect 53765 11664 53821 11666
rect 53765 11612 53767 11664
rect 53767 11612 53819 11664
rect 53819 11612 53821 11664
rect 53765 11610 53821 11612
rect 53765 11560 53821 11562
rect 53765 11508 53767 11560
rect 53767 11508 53819 11560
rect 53819 11508 53821 11560
rect 53765 11506 53821 11508
rect 51138 10260 51194 10316
rect 51242 10260 51298 10316
rect 51346 10260 51402 10316
rect 51138 10156 51194 10212
rect 51242 10156 51298 10212
rect 51346 10156 51402 10212
rect 51138 10052 51194 10108
rect 51242 10052 51298 10108
rect 51346 10052 51402 10108
rect 51138 9200 51194 9256
rect 51242 9200 51298 9256
rect 51346 9200 51402 9256
rect 51138 9096 51194 9152
rect 51242 9096 51298 9152
rect 51346 9096 51402 9152
rect 51138 8992 51194 9048
rect 51242 8992 51298 9048
rect 51346 8992 51402 9048
rect 51138 8534 51194 8590
rect 51242 8534 51298 8590
rect 51346 8534 51402 8590
rect 51138 8430 51194 8486
rect 51242 8430 51298 8486
rect 51346 8430 51402 8486
rect 51138 8326 51194 8382
rect 51242 8326 51298 8382
rect 51346 8326 51402 8382
rect 51530 11320 51586 11376
rect 51634 11320 51690 11376
rect 51738 11320 51794 11376
rect 51530 11216 51586 11272
rect 51634 11216 51690 11272
rect 51738 11216 51794 11272
rect 51530 11112 51586 11168
rect 51634 11112 51690 11168
rect 51738 11112 51794 11168
rect 52804 11270 52860 11272
rect 52804 11218 52806 11270
rect 52806 11218 52858 11270
rect 52858 11218 52860 11270
rect 52804 11216 52860 11218
rect 52804 11166 52860 11168
rect 52804 11114 52806 11166
rect 52806 11114 52858 11166
rect 52858 11114 52860 11166
rect 52804 11112 52860 11114
rect 53444 11270 53500 11272
rect 53444 11218 53446 11270
rect 53446 11218 53498 11270
rect 53498 11218 53500 11270
rect 53444 11216 53500 11218
rect 53444 11166 53500 11168
rect 53444 11114 53446 11166
rect 53446 11114 53498 11166
rect 53498 11114 53500 11166
rect 53444 11112 53500 11114
rect 51530 10654 51586 10710
rect 51634 10654 51690 10710
rect 51738 10654 51794 10710
rect 54405 11664 54461 11666
rect 54405 11612 54407 11664
rect 54407 11612 54459 11664
rect 54459 11612 54461 11664
rect 54405 11610 54461 11612
rect 54405 11560 54461 11562
rect 54405 11508 54407 11560
rect 54407 11508 54459 11560
rect 54459 11508 54461 11560
rect 54405 11506 54461 11508
rect 55045 11664 55101 11666
rect 55045 11612 55047 11664
rect 55047 11612 55099 11664
rect 55099 11612 55101 11664
rect 55045 11610 55101 11612
rect 55045 11560 55101 11562
rect 55045 11508 55047 11560
rect 55047 11508 55099 11560
rect 55099 11508 55101 11560
rect 55045 11506 55101 11508
rect 57259 11664 57315 11666
rect 57259 11612 57261 11664
rect 57261 11612 57313 11664
rect 57313 11612 57315 11664
rect 57259 11610 57315 11612
rect 57259 11560 57315 11562
rect 57259 11508 57261 11560
rect 57261 11508 57313 11560
rect 57313 11508 57315 11560
rect 57259 11506 57315 11508
rect 57899 11664 57955 11666
rect 57899 11612 57901 11664
rect 57901 11612 57953 11664
rect 57953 11612 57955 11664
rect 57899 11610 57955 11612
rect 57899 11560 57955 11562
rect 57899 11508 57901 11560
rect 57901 11508 57953 11560
rect 57953 11508 57955 11560
rect 57899 11506 57955 11508
rect 54724 11270 54780 11272
rect 54724 11218 54726 11270
rect 54726 11218 54778 11270
rect 54778 11218 54780 11270
rect 54724 11216 54780 11218
rect 54724 11166 54780 11168
rect 54724 11114 54726 11166
rect 54726 11114 54778 11166
rect 54778 11114 54780 11166
rect 54724 11112 54780 11114
rect 55364 11270 55420 11272
rect 55364 11218 55366 11270
rect 55366 11218 55418 11270
rect 55418 11218 55420 11270
rect 55364 11216 55420 11218
rect 55364 11166 55420 11168
rect 55364 11114 55366 11166
rect 55366 11114 55418 11166
rect 55418 11114 55420 11166
rect 55364 11112 55420 11114
rect 56940 11270 56996 11272
rect 56940 11218 56942 11270
rect 56942 11218 56994 11270
rect 56994 11218 56996 11270
rect 56940 11216 56996 11218
rect 56940 11166 56996 11168
rect 56940 11114 56942 11166
rect 56942 11114 56994 11166
rect 56994 11114 56996 11166
rect 56940 11112 56996 11114
rect 57580 11270 57636 11272
rect 57580 11218 57582 11270
rect 57582 11218 57634 11270
rect 57634 11218 57636 11270
rect 57580 11216 57636 11218
rect 57580 11166 57636 11168
rect 57580 11114 57582 11166
rect 57582 11114 57634 11166
rect 57634 11114 57636 11166
rect 57580 11112 57636 11114
rect 51530 10550 51586 10606
rect 51634 10550 51690 10606
rect 51738 10550 51794 10606
rect 51530 10446 51586 10502
rect 51634 10446 51690 10502
rect 51738 10446 51794 10502
rect 53125 10604 53181 10606
rect 53125 10552 53127 10604
rect 53127 10552 53179 10604
rect 53179 10552 53181 10604
rect 53125 10550 53181 10552
rect 53125 10500 53181 10502
rect 53125 10448 53127 10500
rect 53127 10448 53179 10500
rect 53179 10448 53181 10500
rect 53125 10446 53181 10448
rect 53765 10604 53821 10606
rect 53765 10552 53767 10604
rect 53767 10552 53819 10604
rect 53819 10552 53821 10604
rect 53765 10550 53821 10552
rect 53765 10500 53821 10502
rect 53765 10448 53767 10500
rect 53767 10448 53819 10500
rect 53819 10448 53821 10500
rect 53765 10446 53821 10448
rect 52804 10210 52860 10212
rect 52804 10158 52806 10210
rect 52806 10158 52858 10210
rect 52858 10158 52860 10210
rect 52804 10156 52860 10158
rect 52804 10106 52860 10108
rect 52804 10054 52806 10106
rect 52806 10054 52858 10106
rect 52858 10054 52860 10106
rect 52804 10052 52860 10054
rect 53444 10210 53500 10212
rect 53444 10158 53446 10210
rect 53446 10158 53498 10210
rect 53498 10158 53500 10210
rect 53444 10156 53500 10158
rect 53444 10106 53500 10108
rect 53444 10054 53446 10106
rect 53446 10054 53498 10106
rect 53498 10054 53500 10106
rect 53444 10052 53500 10054
rect 51530 9594 51586 9650
rect 51634 9594 51690 9650
rect 51738 9594 51794 9650
rect 60919 11714 60975 11770
rect 61023 11714 61079 11770
rect 61127 11714 61183 11770
rect 58539 11664 58595 11666
rect 58539 11612 58541 11664
rect 58541 11612 58593 11664
rect 58593 11612 58595 11664
rect 58539 11610 58595 11612
rect 58539 11560 58595 11562
rect 58539 11508 58541 11560
rect 58541 11508 58593 11560
rect 58593 11508 58595 11560
rect 58539 11506 58595 11508
rect 59179 11664 59235 11666
rect 59179 11612 59181 11664
rect 59181 11612 59233 11664
rect 59233 11612 59235 11664
rect 59179 11610 59235 11612
rect 59179 11560 59235 11562
rect 59179 11508 59181 11560
rect 59181 11508 59233 11560
rect 59233 11508 59235 11560
rect 59179 11506 59235 11508
rect 60919 11610 60975 11666
rect 61023 11610 61079 11666
rect 61127 11610 61183 11666
rect 60919 11506 60975 11562
rect 61023 11506 61079 11562
rect 61127 11506 61183 11562
rect 60514 11320 60570 11376
rect 60618 11320 60674 11376
rect 60722 11320 60778 11376
rect 58860 11270 58916 11272
rect 58860 11218 58862 11270
rect 58862 11218 58914 11270
rect 58914 11218 58916 11270
rect 58860 11216 58916 11218
rect 58860 11166 58916 11168
rect 58860 11114 58862 11166
rect 58862 11114 58914 11166
rect 58914 11114 58916 11166
rect 58860 11112 58916 11114
rect 59500 11270 59556 11272
rect 59500 11218 59502 11270
rect 59502 11218 59554 11270
rect 59554 11218 59556 11270
rect 59500 11216 59556 11218
rect 59500 11166 59556 11168
rect 59500 11114 59502 11166
rect 59502 11114 59554 11166
rect 59554 11114 59556 11166
rect 59500 11112 59556 11114
rect 60514 11216 60570 11272
rect 60618 11216 60674 11272
rect 60722 11216 60778 11272
rect 60514 11112 60570 11168
rect 60618 11112 60674 11168
rect 60722 11112 60778 11168
rect 54405 10604 54461 10606
rect 54405 10552 54407 10604
rect 54407 10552 54459 10604
rect 54459 10552 54461 10604
rect 54405 10550 54461 10552
rect 54405 10500 54461 10502
rect 54405 10448 54407 10500
rect 54407 10448 54459 10500
rect 54459 10448 54461 10500
rect 54405 10446 54461 10448
rect 55045 10604 55101 10606
rect 55045 10552 55047 10604
rect 55047 10552 55099 10604
rect 55099 10552 55101 10604
rect 55045 10550 55101 10552
rect 55045 10500 55101 10502
rect 55045 10448 55047 10500
rect 55047 10448 55099 10500
rect 55099 10448 55101 10500
rect 55045 10446 55101 10448
rect 57259 10604 57315 10606
rect 57259 10552 57261 10604
rect 57261 10552 57313 10604
rect 57313 10552 57315 10604
rect 57259 10550 57315 10552
rect 57259 10500 57315 10502
rect 57259 10448 57261 10500
rect 57261 10448 57313 10500
rect 57313 10448 57315 10500
rect 57259 10446 57315 10448
rect 57899 10604 57955 10606
rect 57899 10552 57901 10604
rect 57901 10552 57953 10604
rect 57953 10552 57955 10604
rect 57899 10550 57955 10552
rect 57899 10500 57955 10502
rect 57899 10448 57901 10500
rect 57901 10448 57953 10500
rect 57953 10448 57955 10500
rect 57899 10446 57955 10448
rect 54724 10210 54780 10212
rect 54724 10158 54726 10210
rect 54726 10158 54778 10210
rect 54778 10158 54780 10210
rect 54724 10156 54780 10158
rect 54724 10106 54780 10108
rect 54724 10054 54726 10106
rect 54726 10054 54778 10106
rect 54778 10054 54780 10106
rect 54724 10052 54780 10054
rect 55364 10210 55420 10212
rect 55364 10158 55366 10210
rect 55366 10158 55418 10210
rect 55418 10158 55420 10210
rect 55364 10156 55420 10158
rect 55364 10106 55420 10108
rect 55364 10054 55366 10106
rect 55366 10054 55418 10106
rect 55418 10054 55420 10106
rect 55364 10052 55420 10054
rect 56940 10210 56996 10212
rect 56940 10158 56942 10210
rect 56942 10158 56994 10210
rect 56994 10158 56996 10210
rect 56940 10156 56996 10158
rect 56940 10106 56996 10108
rect 56940 10054 56942 10106
rect 56942 10054 56994 10106
rect 56994 10054 56996 10106
rect 56940 10052 56996 10054
rect 57580 10210 57636 10212
rect 57580 10158 57582 10210
rect 57582 10158 57634 10210
rect 57634 10158 57636 10210
rect 57580 10156 57636 10158
rect 57580 10106 57636 10108
rect 57580 10054 57582 10106
rect 57582 10054 57634 10106
rect 57634 10054 57636 10106
rect 57580 10052 57636 10054
rect 51530 9490 51586 9546
rect 51634 9490 51690 9546
rect 51738 9490 51794 9546
rect 51530 9386 51586 9442
rect 51634 9386 51690 9442
rect 51738 9386 51794 9442
rect 50798 8140 50854 8196
rect 50902 8140 50958 8196
rect 51006 8140 51062 8196
rect 41842 8036 41898 8092
rect 41946 8036 42002 8092
rect 42050 8036 42106 8092
rect 41842 7932 41898 7988
rect 41946 7932 42002 7988
rect 42050 7932 42106 7988
rect 43108 8090 43164 8092
rect 43108 8038 43110 8090
rect 43110 8038 43162 8090
rect 43162 8038 43164 8090
rect 43108 8036 43164 8038
rect 43108 7986 43164 7988
rect 43108 7934 43110 7986
rect 43110 7934 43162 7986
rect 43162 7934 43164 7986
rect 43108 7932 43164 7934
rect 43748 8090 43804 8092
rect 43748 8038 43750 8090
rect 43750 8038 43802 8090
rect 43802 8038 43804 8090
rect 43748 8036 43804 8038
rect 43748 7986 43804 7988
rect 43748 7934 43750 7986
rect 43750 7934 43802 7986
rect 43802 7934 43804 7986
rect 43748 7932 43804 7934
rect 45028 8090 45084 8092
rect 45028 8038 45030 8090
rect 45030 8038 45082 8090
rect 45082 8038 45084 8090
rect 45028 8036 45084 8038
rect 45028 7986 45084 7988
rect 45028 7934 45030 7986
rect 45030 7934 45082 7986
rect 45082 7934 45084 7986
rect 45028 7932 45084 7934
rect 45668 8090 45724 8092
rect 45668 8038 45670 8090
rect 45670 8038 45722 8090
rect 45722 8038 45724 8090
rect 45668 8036 45724 8038
rect 45668 7986 45724 7988
rect 45668 7934 45670 7986
rect 45670 7934 45722 7986
rect 45722 7934 45724 7986
rect 45668 7932 45724 7934
rect 47244 8090 47300 8092
rect 47244 8038 47246 8090
rect 47246 8038 47298 8090
rect 47298 8038 47300 8090
rect 47244 8036 47300 8038
rect 47244 7986 47300 7988
rect 47244 7934 47246 7986
rect 47246 7934 47298 7986
rect 47298 7934 47300 7986
rect 47244 7932 47300 7934
rect 47884 8090 47940 8092
rect 47884 8038 47886 8090
rect 47886 8038 47938 8090
rect 47938 8038 47940 8090
rect 47884 8036 47940 8038
rect 47884 7986 47940 7988
rect 47884 7934 47886 7986
rect 47886 7934 47938 7986
rect 47938 7934 47940 7986
rect 47884 7932 47940 7934
rect 49164 8090 49220 8092
rect 49164 8038 49166 8090
rect 49166 8038 49218 8090
rect 49218 8038 49220 8090
rect 49164 8036 49220 8038
rect 49164 7986 49220 7988
rect 49164 7934 49166 7986
rect 49166 7934 49218 7986
rect 49218 7934 49220 7986
rect 49164 7932 49220 7934
rect 49804 8090 49860 8092
rect 49804 8038 49806 8090
rect 49806 8038 49858 8090
rect 49858 8038 49860 8090
rect 49804 8036 49860 8038
rect 49804 7986 49860 7988
rect 49804 7934 49806 7986
rect 49806 7934 49858 7986
rect 49858 7934 49860 7986
rect 49804 7932 49860 7934
rect 50798 8036 50854 8092
rect 50902 8036 50958 8092
rect 51006 8036 51062 8092
rect 50798 7932 50854 7988
rect 50902 7932 50958 7988
rect 51006 7932 51062 7988
rect 53125 9544 53181 9546
rect 53125 9492 53127 9544
rect 53127 9492 53179 9544
rect 53179 9492 53181 9544
rect 53125 9490 53181 9492
rect 53125 9440 53181 9442
rect 53125 9388 53127 9440
rect 53127 9388 53179 9440
rect 53179 9388 53181 9440
rect 53125 9386 53181 9388
rect 53765 9544 53821 9546
rect 53765 9492 53767 9544
rect 53767 9492 53819 9544
rect 53819 9492 53821 9544
rect 53765 9490 53821 9492
rect 53765 9440 53821 9442
rect 53765 9388 53767 9440
rect 53767 9388 53819 9440
rect 53819 9388 53821 9440
rect 53765 9386 53821 9388
rect 52804 9150 52860 9152
rect 52804 9098 52806 9150
rect 52806 9098 52858 9150
rect 52858 9098 52860 9150
rect 52804 9096 52860 9098
rect 52804 9046 52860 9048
rect 52804 8994 52806 9046
rect 52806 8994 52858 9046
rect 52858 8994 52860 9046
rect 52804 8992 52860 8994
rect 53444 9150 53500 9152
rect 53444 9098 53446 9150
rect 53446 9098 53498 9150
rect 53498 9098 53500 9150
rect 53444 9096 53500 9098
rect 53444 9046 53500 9048
rect 53444 8994 53446 9046
rect 53446 8994 53498 9046
rect 53498 8994 53500 9046
rect 53444 8992 53500 8994
rect 60514 10654 60570 10710
rect 60618 10654 60674 10710
rect 60722 10654 60778 10710
rect 58539 10604 58595 10606
rect 58539 10552 58541 10604
rect 58541 10552 58593 10604
rect 58593 10552 58595 10604
rect 58539 10550 58595 10552
rect 58539 10500 58595 10502
rect 58539 10448 58541 10500
rect 58541 10448 58593 10500
rect 58593 10448 58595 10500
rect 58539 10446 58595 10448
rect 59179 10604 59235 10606
rect 59179 10552 59181 10604
rect 59181 10552 59233 10604
rect 59233 10552 59235 10604
rect 59179 10550 59235 10552
rect 59179 10500 59235 10502
rect 59179 10448 59181 10500
rect 59181 10448 59233 10500
rect 59233 10448 59235 10500
rect 59179 10446 59235 10448
rect 60514 10550 60570 10606
rect 60618 10550 60674 10606
rect 60722 10550 60778 10606
rect 60514 10446 60570 10502
rect 60618 10446 60674 10502
rect 60722 10446 60778 10502
rect 58860 10210 58916 10212
rect 58860 10158 58862 10210
rect 58862 10158 58914 10210
rect 58914 10158 58916 10210
rect 58860 10156 58916 10158
rect 58860 10106 58916 10108
rect 58860 10054 58862 10106
rect 58862 10054 58914 10106
rect 58914 10054 58916 10106
rect 58860 10052 58916 10054
rect 59500 10210 59556 10212
rect 59500 10158 59502 10210
rect 59502 10158 59554 10210
rect 59554 10158 59556 10210
rect 59500 10156 59556 10158
rect 59500 10106 59556 10108
rect 59500 10054 59502 10106
rect 59502 10054 59554 10106
rect 59554 10054 59556 10106
rect 59500 10052 59556 10054
rect 54405 9544 54461 9546
rect 54405 9492 54407 9544
rect 54407 9492 54459 9544
rect 54459 9492 54461 9544
rect 54405 9490 54461 9492
rect 54405 9440 54461 9442
rect 54405 9388 54407 9440
rect 54407 9388 54459 9440
rect 54459 9388 54461 9440
rect 54405 9386 54461 9388
rect 55045 9544 55101 9546
rect 55045 9492 55047 9544
rect 55047 9492 55099 9544
rect 55099 9492 55101 9544
rect 55045 9490 55101 9492
rect 55045 9440 55101 9442
rect 55045 9388 55047 9440
rect 55047 9388 55099 9440
rect 55099 9388 55101 9440
rect 55045 9386 55101 9388
rect 57259 9544 57315 9546
rect 57259 9492 57261 9544
rect 57261 9492 57313 9544
rect 57313 9492 57315 9544
rect 57259 9490 57315 9492
rect 57259 9440 57315 9442
rect 57259 9388 57261 9440
rect 57261 9388 57313 9440
rect 57313 9388 57315 9440
rect 57259 9386 57315 9388
rect 57899 9544 57955 9546
rect 57899 9492 57901 9544
rect 57901 9492 57953 9544
rect 57953 9492 57955 9544
rect 57899 9490 57955 9492
rect 57899 9440 57955 9442
rect 57899 9388 57901 9440
rect 57901 9388 57953 9440
rect 57953 9388 57955 9440
rect 57899 9386 57955 9388
rect 54724 9150 54780 9152
rect 54724 9098 54726 9150
rect 54726 9098 54778 9150
rect 54778 9098 54780 9150
rect 54724 9096 54780 9098
rect 54724 9046 54780 9048
rect 54724 8994 54726 9046
rect 54726 8994 54778 9046
rect 54778 8994 54780 9046
rect 54724 8992 54780 8994
rect 55364 9150 55420 9152
rect 55364 9098 55366 9150
rect 55366 9098 55418 9150
rect 55418 9098 55420 9150
rect 55364 9096 55420 9098
rect 55364 9046 55420 9048
rect 55364 8994 55366 9046
rect 55366 8994 55418 9046
rect 55418 8994 55420 9046
rect 55364 8992 55420 8994
rect 56940 9150 56996 9152
rect 56940 9098 56942 9150
rect 56942 9098 56994 9150
rect 56994 9098 56996 9150
rect 56940 9096 56996 9098
rect 56940 9046 56996 9048
rect 56940 8994 56942 9046
rect 56942 8994 56994 9046
rect 56994 8994 56996 9046
rect 56940 8992 56996 8994
rect 57580 9150 57636 9152
rect 57580 9098 57582 9150
rect 57582 9098 57634 9150
rect 57634 9098 57636 9150
rect 57580 9096 57636 9098
rect 57580 9046 57636 9048
rect 57580 8994 57582 9046
rect 57582 8994 57634 9046
rect 57634 8994 57636 9046
rect 57580 8992 57636 8994
rect 60514 9594 60570 9650
rect 60618 9594 60674 9650
rect 60722 9594 60778 9650
rect 58539 9544 58595 9546
rect 58539 9492 58541 9544
rect 58541 9492 58593 9544
rect 58593 9492 58595 9544
rect 58539 9490 58595 9492
rect 58539 9440 58595 9442
rect 58539 9388 58541 9440
rect 58541 9388 58593 9440
rect 58593 9388 58595 9440
rect 58539 9386 58595 9388
rect 59179 9544 59235 9546
rect 59179 9492 59181 9544
rect 59181 9492 59233 9544
rect 59233 9492 59235 9544
rect 59179 9490 59235 9492
rect 59179 9440 59235 9442
rect 59179 9388 59181 9440
rect 59181 9388 59233 9440
rect 59233 9388 59235 9440
rect 59179 9386 59235 9388
rect 60514 9490 60570 9546
rect 60618 9490 60674 9546
rect 60722 9490 60778 9546
rect 60514 9386 60570 9442
rect 60618 9386 60674 9442
rect 60722 9386 60778 9442
rect 58860 9150 58916 9152
rect 58860 9098 58862 9150
rect 58862 9098 58914 9150
rect 58914 9098 58916 9150
rect 58860 9096 58916 9098
rect 58860 9046 58916 9048
rect 58860 8994 58862 9046
rect 58862 8994 58914 9046
rect 58914 8994 58916 9046
rect 58860 8992 58916 8994
rect 59500 9150 59556 9152
rect 59500 9098 59502 9150
rect 59502 9098 59554 9150
rect 59554 9098 59556 9150
rect 59500 9096 59556 9098
rect 59500 9046 59556 9048
rect 59500 8994 59502 9046
rect 59502 8994 59554 9046
rect 59554 8994 59556 9046
rect 59500 8992 59556 8994
rect 53125 8484 53181 8486
rect 53125 8432 53127 8484
rect 53127 8432 53179 8484
rect 53179 8432 53181 8484
rect 53125 8430 53181 8432
rect 53125 8380 53181 8382
rect 53125 8328 53127 8380
rect 53127 8328 53179 8380
rect 53179 8328 53181 8380
rect 53125 8326 53181 8328
rect 53765 8484 53821 8486
rect 53765 8432 53767 8484
rect 53767 8432 53819 8484
rect 53819 8432 53821 8484
rect 53765 8430 53821 8432
rect 53765 8380 53821 8382
rect 53765 8328 53767 8380
rect 53767 8328 53819 8380
rect 53819 8328 53821 8380
rect 53765 8326 53821 8328
rect 54405 8484 54461 8486
rect 54405 8432 54407 8484
rect 54407 8432 54459 8484
rect 54459 8432 54461 8484
rect 54405 8430 54461 8432
rect 54405 8380 54461 8382
rect 54405 8328 54407 8380
rect 54407 8328 54459 8380
rect 54459 8328 54461 8380
rect 54405 8326 54461 8328
rect 55045 8484 55101 8486
rect 55045 8432 55047 8484
rect 55047 8432 55099 8484
rect 55099 8432 55101 8484
rect 55045 8430 55101 8432
rect 55045 8380 55101 8382
rect 55045 8328 55047 8380
rect 55047 8328 55099 8380
rect 55099 8328 55101 8380
rect 55045 8326 55101 8328
rect 57259 8484 57315 8486
rect 57259 8432 57261 8484
rect 57261 8432 57313 8484
rect 57313 8432 57315 8484
rect 57259 8430 57315 8432
rect 57259 8380 57315 8382
rect 57259 8328 57261 8380
rect 57261 8328 57313 8380
rect 57313 8328 57315 8380
rect 57259 8326 57315 8328
rect 57899 8484 57955 8486
rect 57899 8432 57901 8484
rect 57901 8432 57953 8484
rect 57953 8432 57955 8484
rect 57899 8430 57955 8432
rect 57899 8380 57955 8382
rect 57899 8328 57901 8380
rect 57901 8328 57953 8380
rect 57953 8328 57955 8380
rect 57899 8326 57955 8328
rect 58539 8484 58595 8486
rect 58539 8432 58541 8484
rect 58541 8432 58593 8484
rect 58593 8432 58595 8484
rect 58539 8430 58595 8432
rect 58539 8380 58595 8382
rect 58539 8328 58541 8380
rect 58541 8328 58593 8380
rect 58593 8328 58595 8380
rect 58539 8326 58595 8328
rect 59179 8484 59235 8486
rect 59179 8432 59181 8484
rect 59181 8432 59233 8484
rect 59233 8432 59235 8484
rect 59179 8430 59235 8432
rect 59179 8380 59235 8382
rect 59179 8328 59181 8380
rect 59181 8328 59233 8380
rect 59233 8328 59235 8380
rect 59179 8326 59235 8328
rect 51530 8140 51586 8196
rect 51634 8140 51690 8196
rect 51738 8140 51794 8196
rect 62821 11664 62877 11666
rect 62821 11612 62823 11664
rect 62823 11612 62875 11664
rect 62875 11612 62877 11664
rect 62821 11610 62877 11612
rect 62821 11560 62877 11562
rect 62821 11508 62823 11560
rect 62823 11508 62875 11560
rect 62875 11508 62877 11560
rect 62821 11506 62877 11508
rect 63461 11664 63517 11666
rect 63461 11612 63463 11664
rect 63463 11612 63515 11664
rect 63515 11612 63517 11664
rect 63461 11610 63517 11612
rect 63461 11560 63517 11562
rect 63461 11508 63463 11560
rect 63463 11508 63515 11560
rect 63515 11508 63517 11560
rect 63461 11506 63517 11508
rect 60919 10260 60975 10316
rect 61023 10260 61079 10316
rect 61127 10260 61183 10316
rect 60919 10156 60975 10212
rect 61023 10156 61079 10212
rect 61127 10156 61183 10212
rect 60919 10052 60975 10108
rect 61023 10052 61079 10108
rect 61127 10052 61183 10108
rect 60919 9200 60975 9256
rect 61023 9200 61079 9256
rect 61127 9200 61183 9256
rect 60919 9096 60975 9152
rect 61023 9096 61079 9152
rect 61127 9096 61183 9152
rect 60919 8992 60975 9048
rect 61023 8992 61079 9048
rect 61127 8992 61183 9048
rect 60919 8534 60975 8590
rect 61023 8534 61079 8590
rect 61127 8534 61183 8590
rect 60919 8430 60975 8486
rect 61023 8430 61079 8486
rect 61127 8430 61183 8486
rect 60919 8326 60975 8382
rect 61023 8326 61079 8382
rect 61127 8326 61183 8382
rect 61278 11320 61334 11376
rect 61382 11320 61438 11376
rect 61486 11320 61542 11376
rect 61278 11216 61334 11272
rect 61382 11216 61438 11272
rect 61486 11216 61542 11272
rect 61278 11112 61334 11168
rect 61382 11112 61438 11168
rect 61486 11112 61542 11168
rect 62500 11270 62556 11272
rect 62500 11218 62502 11270
rect 62502 11218 62554 11270
rect 62554 11218 62556 11270
rect 62500 11216 62556 11218
rect 62500 11166 62556 11168
rect 62500 11114 62502 11166
rect 62502 11114 62554 11166
rect 62554 11114 62556 11166
rect 62500 11112 62556 11114
rect 63140 11270 63196 11272
rect 63140 11218 63142 11270
rect 63142 11218 63194 11270
rect 63194 11218 63196 11270
rect 63140 11216 63196 11218
rect 63140 11166 63196 11168
rect 63140 11114 63142 11166
rect 63142 11114 63194 11166
rect 63194 11114 63196 11166
rect 63140 11112 63196 11114
rect 61278 10654 61334 10710
rect 61382 10654 61438 10710
rect 61486 10654 61542 10710
rect 64101 11664 64157 11666
rect 64101 11612 64103 11664
rect 64103 11612 64155 11664
rect 64155 11612 64157 11664
rect 64101 11610 64157 11612
rect 64101 11560 64157 11562
rect 64101 11508 64103 11560
rect 64103 11508 64155 11560
rect 64155 11508 64157 11560
rect 64101 11506 64157 11508
rect 64741 11664 64797 11666
rect 64741 11612 64743 11664
rect 64743 11612 64795 11664
rect 64795 11612 64797 11664
rect 64741 11610 64797 11612
rect 64741 11560 64797 11562
rect 64741 11508 64743 11560
rect 64743 11508 64795 11560
rect 64795 11508 64797 11560
rect 64741 11506 64797 11508
rect 64420 11270 64476 11272
rect 64420 11218 64422 11270
rect 64422 11218 64474 11270
rect 64474 11218 64476 11270
rect 64420 11216 64476 11218
rect 64420 11166 64476 11168
rect 64420 11114 64422 11166
rect 64422 11114 64474 11166
rect 64474 11114 64476 11166
rect 64420 11112 64476 11114
rect 65060 11270 65116 11272
rect 65060 11218 65062 11270
rect 65062 11218 65114 11270
rect 65114 11218 65116 11270
rect 65060 11216 65116 11218
rect 65060 11166 65116 11168
rect 65060 11114 65062 11166
rect 65062 11114 65114 11166
rect 65114 11114 65116 11166
rect 65060 11112 65116 11114
rect 61278 10550 61334 10606
rect 61382 10550 61438 10606
rect 61486 10550 61542 10606
rect 61278 10446 61334 10502
rect 61382 10446 61438 10502
rect 61486 10446 61542 10502
rect 62821 10604 62877 10606
rect 62821 10552 62823 10604
rect 62823 10552 62875 10604
rect 62875 10552 62877 10604
rect 62821 10550 62877 10552
rect 62821 10500 62877 10502
rect 62821 10448 62823 10500
rect 62823 10448 62875 10500
rect 62875 10448 62877 10500
rect 62821 10446 62877 10448
rect 63461 10604 63517 10606
rect 63461 10552 63463 10604
rect 63463 10552 63515 10604
rect 63515 10552 63517 10604
rect 63461 10550 63517 10552
rect 63461 10500 63517 10502
rect 63461 10448 63463 10500
rect 63463 10448 63515 10500
rect 63515 10448 63517 10500
rect 63461 10446 63517 10448
rect 62500 10210 62556 10212
rect 62500 10158 62502 10210
rect 62502 10158 62554 10210
rect 62554 10158 62556 10210
rect 62500 10156 62556 10158
rect 62500 10106 62556 10108
rect 62500 10054 62502 10106
rect 62502 10054 62554 10106
rect 62554 10054 62556 10106
rect 62500 10052 62556 10054
rect 63140 10210 63196 10212
rect 63140 10158 63142 10210
rect 63142 10158 63194 10210
rect 63194 10158 63196 10210
rect 63140 10156 63196 10158
rect 63140 10106 63196 10108
rect 63140 10054 63142 10106
rect 63142 10054 63194 10106
rect 63194 10054 63196 10106
rect 63140 10052 63196 10054
rect 61278 9594 61334 9650
rect 61382 9594 61438 9650
rect 61486 9594 61542 9650
rect 64101 10604 64157 10606
rect 64101 10552 64103 10604
rect 64103 10552 64155 10604
rect 64155 10552 64157 10604
rect 64101 10550 64157 10552
rect 64101 10500 64157 10502
rect 64101 10448 64103 10500
rect 64103 10448 64155 10500
rect 64155 10448 64157 10500
rect 64101 10446 64157 10448
rect 64741 10604 64797 10606
rect 64741 10552 64743 10604
rect 64743 10552 64795 10604
rect 64795 10552 64797 10604
rect 64741 10550 64797 10552
rect 64741 10500 64797 10502
rect 64741 10448 64743 10500
rect 64743 10448 64795 10500
rect 64795 10448 64797 10500
rect 64741 10446 64797 10448
rect 64420 10210 64476 10212
rect 64420 10158 64422 10210
rect 64422 10158 64474 10210
rect 64474 10158 64476 10210
rect 64420 10156 64476 10158
rect 64420 10106 64476 10108
rect 64420 10054 64422 10106
rect 64422 10054 64474 10106
rect 64474 10054 64476 10106
rect 64420 10052 64476 10054
rect 65060 10210 65116 10212
rect 65060 10158 65062 10210
rect 65062 10158 65114 10210
rect 65114 10158 65116 10210
rect 65060 10156 65116 10158
rect 65060 10106 65116 10108
rect 65060 10054 65062 10106
rect 65062 10054 65114 10106
rect 65114 10054 65116 10106
rect 65060 10052 65116 10054
rect 61278 9490 61334 9546
rect 61382 9490 61438 9546
rect 61486 9490 61542 9546
rect 61278 9386 61334 9442
rect 61382 9386 61438 9442
rect 61486 9386 61542 9442
rect 60514 8140 60570 8196
rect 60618 8140 60674 8196
rect 60722 8140 60778 8196
rect 51530 8036 51586 8092
rect 51634 8036 51690 8092
rect 51738 8036 51794 8092
rect 51530 7932 51586 7988
rect 51634 7932 51690 7988
rect 51738 7932 51794 7988
rect 52804 8090 52860 8092
rect 52804 8038 52806 8090
rect 52806 8038 52858 8090
rect 52858 8038 52860 8090
rect 52804 8036 52860 8038
rect 52804 7986 52860 7988
rect 52804 7934 52806 7986
rect 52806 7934 52858 7986
rect 52858 7934 52860 7986
rect 52804 7932 52860 7934
rect 53444 8090 53500 8092
rect 53444 8038 53446 8090
rect 53446 8038 53498 8090
rect 53498 8038 53500 8090
rect 53444 8036 53500 8038
rect 53444 7986 53500 7988
rect 53444 7934 53446 7986
rect 53446 7934 53498 7986
rect 53498 7934 53500 7986
rect 53444 7932 53500 7934
rect 54724 8090 54780 8092
rect 54724 8038 54726 8090
rect 54726 8038 54778 8090
rect 54778 8038 54780 8090
rect 54724 8036 54780 8038
rect 54724 7986 54780 7988
rect 54724 7934 54726 7986
rect 54726 7934 54778 7986
rect 54778 7934 54780 7986
rect 54724 7932 54780 7934
rect 55364 8090 55420 8092
rect 55364 8038 55366 8090
rect 55366 8038 55418 8090
rect 55418 8038 55420 8090
rect 55364 8036 55420 8038
rect 55364 7986 55420 7988
rect 55364 7934 55366 7986
rect 55366 7934 55418 7986
rect 55418 7934 55420 7986
rect 55364 7932 55420 7934
rect 56940 8090 56996 8092
rect 56940 8038 56942 8090
rect 56942 8038 56994 8090
rect 56994 8038 56996 8090
rect 56940 8036 56996 8038
rect 56940 7986 56996 7988
rect 56940 7934 56942 7986
rect 56942 7934 56994 7986
rect 56994 7934 56996 7986
rect 56940 7932 56996 7934
rect 57580 8090 57636 8092
rect 57580 8038 57582 8090
rect 57582 8038 57634 8090
rect 57634 8038 57636 8090
rect 57580 8036 57636 8038
rect 57580 7986 57636 7988
rect 57580 7934 57582 7986
rect 57582 7934 57634 7986
rect 57634 7934 57636 7986
rect 57580 7932 57636 7934
rect 58860 8090 58916 8092
rect 58860 8038 58862 8090
rect 58862 8038 58914 8090
rect 58914 8038 58916 8090
rect 58860 8036 58916 8038
rect 58860 7986 58916 7988
rect 58860 7934 58862 7986
rect 58862 7934 58914 7986
rect 58914 7934 58916 7986
rect 58860 7932 58916 7934
rect 59500 8090 59556 8092
rect 59500 8038 59502 8090
rect 59502 8038 59554 8090
rect 59554 8038 59556 8090
rect 59500 8036 59556 8038
rect 59500 7986 59556 7988
rect 59500 7934 59502 7986
rect 59502 7934 59554 7986
rect 59554 7934 59556 7986
rect 59500 7932 59556 7934
rect 60514 8036 60570 8092
rect 60618 8036 60674 8092
rect 60722 8036 60778 8092
rect 60514 7932 60570 7988
rect 60618 7932 60674 7988
rect 60722 7932 60778 7988
rect 62821 9544 62877 9546
rect 62821 9492 62823 9544
rect 62823 9492 62875 9544
rect 62875 9492 62877 9544
rect 62821 9490 62877 9492
rect 62821 9440 62877 9442
rect 62821 9388 62823 9440
rect 62823 9388 62875 9440
rect 62875 9388 62877 9440
rect 62821 9386 62877 9388
rect 63461 9544 63517 9546
rect 63461 9492 63463 9544
rect 63463 9492 63515 9544
rect 63515 9492 63517 9544
rect 63461 9490 63517 9492
rect 63461 9440 63517 9442
rect 63461 9388 63463 9440
rect 63463 9388 63515 9440
rect 63515 9388 63517 9440
rect 63461 9386 63517 9388
rect 62500 9150 62556 9152
rect 62500 9098 62502 9150
rect 62502 9098 62554 9150
rect 62554 9098 62556 9150
rect 62500 9096 62556 9098
rect 62500 9046 62556 9048
rect 62500 8994 62502 9046
rect 62502 8994 62554 9046
rect 62554 8994 62556 9046
rect 62500 8992 62556 8994
rect 63140 9150 63196 9152
rect 63140 9098 63142 9150
rect 63142 9098 63194 9150
rect 63194 9098 63196 9150
rect 63140 9096 63196 9098
rect 63140 9046 63196 9048
rect 63140 8994 63142 9046
rect 63142 8994 63194 9046
rect 63194 8994 63196 9046
rect 63140 8992 63196 8994
rect 64101 9544 64157 9546
rect 64101 9492 64103 9544
rect 64103 9492 64155 9544
rect 64155 9492 64157 9544
rect 64101 9490 64157 9492
rect 64101 9440 64157 9442
rect 64101 9388 64103 9440
rect 64103 9388 64155 9440
rect 64155 9388 64157 9440
rect 64101 9386 64157 9388
rect 64741 9544 64797 9546
rect 64741 9492 64743 9544
rect 64743 9492 64795 9544
rect 64795 9492 64797 9544
rect 64741 9490 64797 9492
rect 64741 9440 64797 9442
rect 64741 9388 64743 9440
rect 64743 9388 64795 9440
rect 64795 9388 64797 9440
rect 64741 9386 64797 9388
rect 64420 9150 64476 9152
rect 64420 9098 64422 9150
rect 64422 9098 64474 9150
rect 64474 9098 64476 9150
rect 64420 9096 64476 9098
rect 64420 9046 64476 9048
rect 64420 8994 64422 9046
rect 64422 8994 64474 9046
rect 64474 8994 64476 9046
rect 64420 8992 64476 8994
rect 65060 9150 65116 9152
rect 65060 9098 65062 9150
rect 65062 9098 65114 9150
rect 65114 9098 65116 9150
rect 65060 9096 65116 9098
rect 65060 9046 65116 9048
rect 65060 8994 65062 9046
rect 65062 8994 65114 9046
rect 65114 8994 65116 9046
rect 65060 8992 65116 8994
rect 62821 8484 62877 8486
rect 62821 8432 62823 8484
rect 62823 8432 62875 8484
rect 62875 8432 62877 8484
rect 62821 8430 62877 8432
rect 62821 8380 62877 8382
rect 62821 8328 62823 8380
rect 62823 8328 62875 8380
rect 62875 8328 62877 8380
rect 62821 8326 62877 8328
rect 63461 8484 63517 8486
rect 63461 8432 63463 8484
rect 63463 8432 63515 8484
rect 63515 8432 63517 8484
rect 63461 8430 63517 8432
rect 63461 8380 63517 8382
rect 63461 8328 63463 8380
rect 63463 8328 63515 8380
rect 63515 8328 63517 8380
rect 63461 8326 63517 8328
rect 64101 8484 64157 8486
rect 64101 8432 64103 8484
rect 64103 8432 64155 8484
rect 64155 8432 64157 8484
rect 64101 8430 64157 8432
rect 64101 8380 64157 8382
rect 64101 8328 64103 8380
rect 64103 8328 64155 8380
rect 64155 8328 64157 8380
rect 64101 8326 64157 8328
rect 64741 8484 64797 8486
rect 64741 8432 64743 8484
rect 64743 8432 64795 8484
rect 64795 8432 64797 8484
rect 64741 8430 64797 8432
rect 64741 8380 64797 8382
rect 64741 8328 64743 8380
rect 64743 8328 64795 8380
rect 64795 8328 64797 8380
rect 64741 8326 64797 8328
rect 61278 8140 61334 8196
rect 61382 8140 61438 8196
rect 61486 8140 61542 8196
rect 61278 8036 61334 8092
rect 61382 8036 61438 8092
rect 61486 8036 61542 8092
rect 61278 7932 61334 7988
rect 61382 7932 61438 7988
rect 61486 7932 61542 7988
rect 62500 8090 62556 8092
rect 62500 8038 62502 8090
rect 62502 8038 62554 8090
rect 62554 8038 62556 8090
rect 62500 8036 62556 8038
rect 62500 7986 62556 7988
rect 62500 7934 62502 7986
rect 62502 7934 62554 7986
rect 62554 7934 62556 7986
rect 62500 7932 62556 7934
rect 63140 8090 63196 8092
rect 63140 8038 63142 8090
rect 63142 8038 63194 8090
rect 63194 8038 63196 8090
rect 63140 8036 63196 8038
rect 63140 7986 63196 7988
rect 63140 7934 63142 7986
rect 63142 7934 63194 7986
rect 63194 7934 63196 7986
rect 63140 7932 63196 7934
rect 64420 8090 64476 8092
rect 64420 8038 64422 8090
rect 64422 8038 64474 8090
rect 64474 8038 64476 8090
rect 64420 8036 64476 8038
rect 64420 7986 64476 7988
rect 64420 7934 64422 7986
rect 64422 7934 64474 7986
rect 64474 7934 64476 7986
rect 64420 7932 64476 7934
rect 65060 8090 65116 8092
rect 65060 8038 65062 8090
rect 65062 8038 65114 8090
rect 65114 8038 65116 8090
rect 65060 8036 65116 8038
rect 65060 7986 65116 7988
rect 65060 7934 65062 7986
rect 65062 7934 65114 7986
rect 65114 7934 65116 7986
rect 65060 7932 65116 7934
rect 34640 3508 34696 3564
rect 34744 3508 34800 3564
rect 34640 3404 34696 3460
rect 34744 3404 34800 3460
rect 45032 1201 45088 1203
rect 45032 1149 45034 1201
rect 45034 1149 45086 1201
rect 45086 1149 45088 1201
rect 45032 1147 45088 1149
rect 45136 1201 45192 1203
rect 45136 1149 45138 1201
rect 45138 1149 45190 1201
rect 45190 1149 45192 1201
rect 45136 1147 45192 1149
rect 45240 1201 45296 1203
rect 45240 1149 45242 1201
rect 45242 1149 45294 1201
rect 45294 1149 45296 1201
rect 45240 1147 45296 1149
rect 45344 1201 45400 1203
rect 45344 1149 45346 1201
rect 45346 1149 45398 1201
rect 45398 1149 45400 1201
rect 45344 1147 45400 1149
rect 45448 1201 45504 1203
rect 45448 1149 45450 1201
rect 45450 1149 45502 1201
rect 45502 1149 45504 1201
rect 45448 1147 45504 1149
rect 35202 1101 35258 1103
rect 35202 1049 35204 1101
rect 35204 1049 35256 1101
rect 35256 1049 35258 1101
rect 35202 1047 35258 1049
rect 35306 1101 35362 1103
rect 35306 1049 35308 1101
rect 35308 1049 35360 1101
rect 35360 1049 35362 1101
rect 35306 1047 35362 1049
rect 35410 1101 35466 1103
rect 35410 1049 35412 1101
rect 35412 1049 35464 1101
rect 35464 1049 35466 1101
rect 35410 1047 35466 1049
rect 35514 1101 35570 1103
rect 35514 1049 35516 1101
rect 35516 1049 35568 1101
rect 35568 1049 35570 1101
rect 35514 1047 35570 1049
rect 35618 1101 35674 1103
rect 35618 1049 35620 1101
rect 35620 1049 35672 1101
rect 35672 1049 35674 1101
rect 35618 1047 35674 1049
rect 35202 997 35258 999
rect 35202 945 35204 997
rect 35204 945 35256 997
rect 35256 945 35258 997
rect 35202 943 35258 945
rect 35306 997 35362 999
rect 35306 945 35308 997
rect 35308 945 35360 997
rect 35360 945 35362 997
rect 35306 943 35362 945
rect 35410 997 35466 999
rect 35410 945 35412 997
rect 35412 945 35464 997
rect 35464 945 35466 997
rect 35410 943 35466 945
rect 35514 997 35570 999
rect 35514 945 35516 997
rect 35516 945 35568 997
rect 35568 945 35570 997
rect 35514 943 35570 945
rect 35618 997 35674 999
rect 35618 945 35620 997
rect 35620 945 35672 997
rect 35672 945 35674 997
rect 35618 943 35674 945
rect 35202 893 35258 895
rect 35202 841 35204 893
rect 35204 841 35256 893
rect 35256 841 35258 893
rect 35202 839 35258 841
rect 35306 893 35362 895
rect 35306 841 35308 893
rect 35308 841 35360 893
rect 35360 841 35362 893
rect 35306 839 35362 841
rect 35410 893 35466 895
rect 35410 841 35412 893
rect 35412 841 35464 893
rect 35464 841 35466 893
rect 35410 839 35466 841
rect 35514 893 35570 895
rect 35514 841 35516 893
rect 35516 841 35568 893
rect 35568 841 35570 893
rect 35514 839 35570 841
rect 35618 893 35674 895
rect 35618 841 35620 893
rect 35620 841 35672 893
rect 35672 841 35674 893
rect 35618 839 35674 841
rect 35202 789 35258 791
rect 35202 737 35204 789
rect 35204 737 35256 789
rect 35256 737 35258 789
rect 35202 735 35258 737
rect 35306 789 35362 791
rect 35306 737 35308 789
rect 35308 737 35360 789
rect 35360 737 35362 789
rect 35306 735 35362 737
rect 35410 789 35466 791
rect 35410 737 35412 789
rect 35412 737 35464 789
rect 35464 737 35466 789
rect 35410 735 35466 737
rect 35514 789 35570 791
rect 35514 737 35516 789
rect 35516 737 35568 789
rect 35568 737 35570 789
rect 35514 735 35570 737
rect 35618 789 35674 791
rect 35618 737 35620 789
rect 35620 737 35672 789
rect 35672 737 35674 789
rect 35618 735 35674 737
rect 35202 685 35258 687
rect 35202 633 35204 685
rect 35204 633 35256 685
rect 35256 633 35258 685
rect 35202 631 35258 633
rect 35306 685 35362 687
rect 35306 633 35308 685
rect 35308 633 35360 685
rect 35360 633 35362 685
rect 35306 631 35362 633
rect 35410 685 35466 687
rect 35410 633 35412 685
rect 35412 633 35464 685
rect 35464 633 35466 685
rect 35410 631 35466 633
rect 35514 685 35570 687
rect 35514 633 35516 685
rect 35516 633 35568 685
rect 35568 633 35570 685
rect 35514 631 35570 633
rect 35618 685 35674 687
rect 35618 633 35620 685
rect 35620 633 35672 685
rect 35672 633 35674 685
rect 35618 631 35674 633
rect 39642 1101 39698 1103
rect 39642 1049 39644 1101
rect 39644 1049 39696 1101
rect 39696 1049 39698 1101
rect 39642 1047 39698 1049
rect 39746 1101 39802 1103
rect 39746 1049 39748 1101
rect 39748 1049 39800 1101
rect 39800 1049 39802 1101
rect 39746 1047 39802 1049
rect 39850 1101 39906 1103
rect 39850 1049 39852 1101
rect 39852 1049 39904 1101
rect 39904 1049 39906 1101
rect 39850 1047 39906 1049
rect 39954 1101 40010 1103
rect 39954 1049 39956 1101
rect 39956 1049 40008 1101
rect 40008 1049 40010 1101
rect 39954 1047 40010 1049
rect 40058 1101 40114 1103
rect 40058 1049 40060 1101
rect 40060 1049 40112 1101
rect 40112 1049 40114 1101
rect 40058 1047 40114 1049
rect 39642 997 39698 999
rect 39642 945 39644 997
rect 39644 945 39696 997
rect 39696 945 39698 997
rect 39642 943 39698 945
rect 39746 997 39802 999
rect 39746 945 39748 997
rect 39748 945 39800 997
rect 39800 945 39802 997
rect 39746 943 39802 945
rect 39850 997 39906 999
rect 39850 945 39852 997
rect 39852 945 39904 997
rect 39904 945 39906 997
rect 39850 943 39906 945
rect 39954 997 40010 999
rect 39954 945 39956 997
rect 39956 945 40008 997
rect 40008 945 40010 997
rect 39954 943 40010 945
rect 40058 997 40114 999
rect 40058 945 40060 997
rect 40060 945 40112 997
rect 40112 945 40114 997
rect 40058 943 40114 945
rect 39642 893 39698 895
rect 39642 841 39644 893
rect 39644 841 39696 893
rect 39696 841 39698 893
rect 39642 839 39698 841
rect 39746 893 39802 895
rect 39746 841 39748 893
rect 39748 841 39800 893
rect 39800 841 39802 893
rect 39746 839 39802 841
rect 39850 893 39906 895
rect 39850 841 39852 893
rect 39852 841 39904 893
rect 39904 841 39906 893
rect 39850 839 39906 841
rect 39954 893 40010 895
rect 39954 841 39956 893
rect 39956 841 40008 893
rect 40008 841 40010 893
rect 39954 839 40010 841
rect 40058 893 40114 895
rect 40058 841 40060 893
rect 40060 841 40112 893
rect 40112 841 40114 893
rect 40058 839 40114 841
rect 39642 789 39698 791
rect 39642 737 39644 789
rect 39644 737 39696 789
rect 39696 737 39698 789
rect 39642 735 39698 737
rect 39746 789 39802 791
rect 39746 737 39748 789
rect 39748 737 39800 789
rect 39800 737 39802 789
rect 39746 735 39802 737
rect 39850 789 39906 791
rect 39850 737 39852 789
rect 39852 737 39904 789
rect 39904 737 39906 789
rect 39850 735 39906 737
rect 39954 789 40010 791
rect 39954 737 39956 789
rect 39956 737 40008 789
rect 40008 737 40010 789
rect 39954 735 40010 737
rect 40058 789 40114 791
rect 40058 737 40060 789
rect 40060 737 40112 789
rect 40112 737 40114 789
rect 40058 735 40114 737
rect 45032 1097 45088 1099
rect 45032 1045 45034 1097
rect 45034 1045 45086 1097
rect 45086 1045 45088 1097
rect 45032 1043 45088 1045
rect 45136 1097 45192 1099
rect 45136 1045 45138 1097
rect 45138 1045 45190 1097
rect 45190 1045 45192 1097
rect 45136 1043 45192 1045
rect 45240 1097 45296 1099
rect 45240 1045 45242 1097
rect 45242 1045 45294 1097
rect 45294 1045 45296 1097
rect 45240 1043 45296 1045
rect 45344 1097 45400 1099
rect 45344 1045 45346 1097
rect 45346 1045 45398 1097
rect 45398 1045 45400 1097
rect 45344 1043 45400 1045
rect 45448 1097 45504 1099
rect 45448 1045 45450 1097
rect 45450 1045 45502 1097
rect 45502 1045 45504 1097
rect 45448 1043 45504 1045
rect 45032 993 45088 995
rect 45032 941 45034 993
rect 45034 941 45086 993
rect 45086 941 45088 993
rect 45032 939 45088 941
rect 45136 993 45192 995
rect 45136 941 45138 993
rect 45138 941 45190 993
rect 45190 941 45192 993
rect 45136 939 45192 941
rect 45240 993 45296 995
rect 45240 941 45242 993
rect 45242 941 45294 993
rect 45294 941 45296 993
rect 45240 939 45296 941
rect 45344 993 45400 995
rect 45344 941 45346 993
rect 45346 941 45398 993
rect 45398 941 45400 993
rect 45344 939 45400 941
rect 45448 993 45504 995
rect 45448 941 45450 993
rect 45450 941 45502 993
rect 45502 941 45504 993
rect 45448 939 45504 941
rect 45032 889 45088 891
rect 45032 837 45034 889
rect 45034 837 45086 889
rect 45086 837 45088 889
rect 45032 835 45088 837
rect 45136 889 45192 891
rect 45136 837 45138 889
rect 45138 837 45190 889
rect 45190 837 45192 889
rect 45136 835 45192 837
rect 45240 889 45296 891
rect 45240 837 45242 889
rect 45242 837 45294 889
rect 45294 837 45296 889
rect 45240 835 45296 837
rect 45344 889 45400 891
rect 45344 837 45346 889
rect 45346 837 45398 889
rect 45398 837 45400 889
rect 45344 835 45400 837
rect 45448 889 45504 891
rect 45448 837 45450 889
rect 45450 837 45502 889
rect 45502 837 45504 889
rect 45448 835 45504 837
rect 45032 785 45088 787
rect 45032 733 45034 785
rect 45034 733 45086 785
rect 45086 733 45088 785
rect 45032 731 45088 733
rect 45136 785 45192 787
rect 45136 733 45138 785
rect 45138 733 45190 785
rect 45190 733 45192 785
rect 45136 731 45192 733
rect 45240 785 45296 787
rect 45240 733 45242 785
rect 45242 733 45294 785
rect 45294 733 45296 785
rect 45240 731 45296 733
rect 45344 785 45400 787
rect 45344 733 45346 785
rect 45346 733 45398 785
rect 45398 733 45400 785
rect 45344 731 45400 733
rect 45448 785 45504 787
rect 45448 733 45450 785
rect 45450 733 45502 785
rect 45502 733 45504 785
rect 45448 731 45504 733
rect 49472 1201 49528 1203
rect 49472 1149 49474 1201
rect 49474 1149 49526 1201
rect 49526 1149 49528 1201
rect 49472 1147 49528 1149
rect 49576 1201 49632 1203
rect 49576 1149 49578 1201
rect 49578 1149 49630 1201
rect 49630 1149 49632 1201
rect 49576 1147 49632 1149
rect 49680 1201 49736 1203
rect 49680 1149 49682 1201
rect 49682 1149 49734 1201
rect 49734 1149 49736 1201
rect 49680 1147 49736 1149
rect 49784 1201 49840 1203
rect 49784 1149 49786 1201
rect 49786 1149 49838 1201
rect 49838 1149 49840 1201
rect 49784 1147 49840 1149
rect 49888 1201 49944 1203
rect 49888 1149 49890 1201
rect 49890 1149 49942 1201
rect 49942 1149 49944 1201
rect 49888 1147 49944 1149
rect 49472 1097 49528 1099
rect 49472 1045 49474 1097
rect 49474 1045 49526 1097
rect 49526 1045 49528 1097
rect 49472 1043 49528 1045
rect 49576 1097 49632 1099
rect 49576 1045 49578 1097
rect 49578 1045 49630 1097
rect 49630 1045 49632 1097
rect 49576 1043 49632 1045
rect 49680 1097 49736 1099
rect 49680 1045 49682 1097
rect 49682 1045 49734 1097
rect 49734 1045 49736 1097
rect 49680 1043 49736 1045
rect 49784 1097 49840 1099
rect 49784 1045 49786 1097
rect 49786 1045 49838 1097
rect 49838 1045 49840 1097
rect 49784 1043 49840 1045
rect 49888 1097 49944 1099
rect 49888 1045 49890 1097
rect 49890 1045 49942 1097
rect 49942 1045 49944 1097
rect 49888 1043 49944 1045
rect 49472 993 49528 995
rect 49472 941 49474 993
rect 49474 941 49526 993
rect 49526 941 49528 993
rect 49472 939 49528 941
rect 49576 993 49632 995
rect 49576 941 49578 993
rect 49578 941 49630 993
rect 49630 941 49632 993
rect 49576 939 49632 941
rect 49680 993 49736 995
rect 49680 941 49682 993
rect 49682 941 49734 993
rect 49734 941 49736 993
rect 49680 939 49736 941
rect 49784 993 49840 995
rect 49784 941 49786 993
rect 49786 941 49838 993
rect 49838 941 49840 993
rect 49784 939 49840 941
rect 49888 993 49944 995
rect 49888 941 49890 993
rect 49890 941 49942 993
rect 49942 941 49944 993
rect 49888 939 49944 941
rect 49472 889 49528 891
rect 49472 837 49474 889
rect 49474 837 49526 889
rect 49526 837 49528 889
rect 49472 835 49528 837
rect 49576 889 49632 891
rect 49576 837 49578 889
rect 49578 837 49630 889
rect 49630 837 49632 889
rect 49576 835 49632 837
rect 49680 889 49736 891
rect 49680 837 49682 889
rect 49682 837 49734 889
rect 49734 837 49736 889
rect 49680 835 49736 837
rect 49784 889 49840 891
rect 49784 837 49786 889
rect 49786 837 49838 889
rect 49838 837 49840 889
rect 49784 835 49840 837
rect 49888 889 49944 891
rect 49888 837 49890 889
rect 49890 837 49942 889
rect 49942 837 49944 889
rect 49888 835 49944 837
rect 49472 785 49528 787
rect 49472 733 49474 785
rect 49474 733 49526 785
rect 49526 733 49528 785
rect 49472 731 49528 733
rect 49576 785 49632 787
rect 49576 733 49578 785
rect 49578 733 49630 785
rect 49630 733 49632 785
rect 49576 731 49632 733
rect 49680 785 49736 787
rect 49680 733 49682 785
rect 49682 733 49734 785
rect 49734 733 49736 785
rect 49680 731 49736 733
rect 49784 785 49840 787
rect 49784 733 49786 785
rect 49786 733 49838 785
rect 49838 733 49840 785
rect 49784 731 49840 733
rect 49888 785 49944 787
rect 49888 733 49890 785
rect 49890 733 49942 785
rect 49942 733 49944 785
rect 49888 731 49944 733
rect 39642 685 39698 687
rect 39642 633 39644 685
rect 39644 633 39696 685
rect 39696 633 39698 685
rect 39642 631 39698 633
rect 39746 685 39802 687
rect 39746 633 39748 685
rect 39748 633 39800 685
rect 39800 633 39802 685
rect 39746 631 39802 633
rect 39850 685 39906 687
rect 39850 633 39852 685
rect 39852 633 39904 685
rect 39904 633 39906 685
rect 39850 631 39906 633
rect 39954 685 40010 687
rect 39954 633 39956 685
rect 39956 633 40008 685
rect 40008 633 40010 685
rect 39954 631 40010 633
rect 40058 685 40114 687
rect 40058 633 40060 685
rect 40060 633 40112 685
rect 40112 633 40114 685
rect 40058 631 40114 633
rect 32136 330 32192 386
rect 32240 330 32296 386
rect 32344 330 32400 386
rect 32136 226 32192 282
rect 32240 226 32296 282
rect 32344 226 32400 282
rect 32136 122 32192 178
rect 32240 122 32296 178
rect 32344 122 32400 178
<< mimcap >>
rect -16170 14548 -12970 14628
rect -16170 11668 -16090 14548
rect -13050 11668 -12970 14548
rect -16170 11588 -12970 11668
rect -12086 14745 -8886 14825
rect -12086 11865 -12006 14745
rect -8966 11865 -8886 14745
rect -12086 11785 -8886 11865
rect -16170 11148 -12970 11228
rect -16170 8268 -16090 11148
rect -13050 8268 -12970 11148
rect -16170 8188 -12970 8268
rect -12086 11345 -8886 11425
rect -12086 8465 -12006 11345
rect -8966 8465 -8886 11345
rect -12086 8385 -8886 8465
rect -7599 14481 -4559 14561
rect -7599 11441 -7519 14481
rect -4639 11441 -4559 14481
rect -7599 11361 -4559 11441
rect -4199 14481 -1159 14561
rect -4199 11441 -4119 14481
rect -1239 11441 -1159 14481
rect -4199 11361 -1159 11441
rect -16170 7000 -12970 7080
rect -16170 4120 -16090 7000
rect -13050 4120 -12970 7000
rect -16170 4040 -12970 4120
rect -12066 7037 -8866 7117
rect -12066 4157 -11986 7037
rect -8946 4157 -8866 7037
rect -12066 4077 -8866 4157
rect -16170 3600 -12970 3680
rect -16170 720 -16090 3600
rect -13050 720 -12970 3600
rect -16170 640 -12970 720
rect -12066 3637 -8866 3717
rect -12066 757 -11986 3637
rect -8946 757 -8866 3637
rect -12066 677 -8866 757
rect -7599 3551 -4559 3631
rect -7599 511 -7519 3551
rect -4639 511 -4559 3551
rect -7599 431 -4559 511
rect -4199 3551 -1159 3631
rect -4199 511 -4119 3551
rect -1239 511 -1159 3551
rect -4199 431 -1159 511
rect 33338 5933 37538 6013
rect 33338 1893 33418 5933
rect 37458 1893 37538 5933
rect 33338 1813 37538 1893
rect 37898 5933 42098 6013
rect 37898 1893 37978 5933
rect 42018 1893 42098 5933
rect 37898 1813 42098 1893
rect 43168 5933 47368 6013
rect 43168 1893 43248 5933
rect 47288 1893 47368 5933
rect 43168 1813 47368 1893
rect 47728 5933 51928 6013
rect 47728 1893 47808 5933
rect 51848 1893 51928 5933
rect 47728 1813 51928 1893
<< mimcapcontact >>
rect -16090 11668 -13050 14548
rect -12006 11865 -8966 14745
rect -16090 8268 -13050 11148
rect -12006 8465 -8966 11345
rect -7519 11441 -4639 14481
rect -4119 11441 -1239 14481
rect -16090 4120 -13050 7000
rect -11986 4157 -8946 7037
rect -16090 720 -13050 3600
rect -11986 757 -8946 3637
rect -7519 511 -4639 3551
rect -4119 511 -1239 3551
rect 33418 1893 37458 5933
rect 37978 1893 42018 5933
rect 43248 1893 47288 5933
rect 47808 1893 51848 5933
<< metal3 >>
rect 374 15706 31505 15718
rect 374 15650 31226 15706
rect 31282 15650 31336 15706
rect 31392 15650 31446 15706
rect 31502 15650 31505 15706
rect 374 15596 31505 15650
rect 374 15540 31226 15596
rect 31282 15540 31336 15596
rect 31392 15540 31446 15596
rect 31502 15540 31505 15596
rect 374 15491 31505 15540
rect 374 15486 31509 15491
rect 374 15430 31226 15486
rect 31282 15430 31336 15486
rect 31392 15430 31446 15486
rect 31502 15430 31509 15486
rect 374 15207 31509 15430
rect 374 13795 957 15207
rect 1233 14772 9208 14935
rect 1224 14742 9208 14772
rect 1223 14686 1233 14742
rect 1289 14686 1343 14742
rect 1399 14686 1453 14742
rect 1509 14686 1563 14742
rect 1619 14686 9208 14742
rect 1224 14632 9208 14686
rect 1224 14576 1233 14632
rect 1289 14576 1343 14632
rect 1399 14576 1453 14632
rect 1509 14576 1563 14632
rect 1619 14576 9208 14632
rect 1224 14488 9208 14576
rect 3161 14328 3341 14338
rect 3950 14328 4026 14338
rect 3161 14272 3171 14328
rect 3227 14272 3275 14328
rect 3331 14272 3960 14328
rect 4016 14272 4026 14328
rect 3161 14224 4026 14272
rect 3161 14168 3171 14224
rect 3227 14168 3275 14224
rect 3331 14168 3960 14224
rect 4016 14168 4026 14224
rect 3161 14158 3341 14168
rect 3950 14158 4026 14168
rect 5731 14274 5911 14284
rect 6735 14274 6811 14284
rect 7375 14274 7451 14284
rect 8015 14274 8091 14284
rect 5731 14218 5741 14274
rect 5797 14218 5845 14274
rect 5901 14218 6745 14274
rect 6801 14218 7385 14274
rect 7441 14218 8025 14274
rect 8081 14218 8091 14274
rect 5731 14170 8091 14218
rect 5731 14114 5741 14170
rect 5797 14114 5845 14170
rect 5901 14114 6745 14170
rect 6801 14114 7385 14170
rect 7441 14114 8025 14170
rect 8081 14114 8091 14170
rect 5731 14104 5911 14114
rect 6735 14104 6811 14114
rect 7375 14104 7451 14114
rect 8015 14104 8091 14114
rect 2520 13979 2700 13989
rect 4030 13979 4106 13989
rect 2520 13923 2530 13979
rect 2586 13923 2634 13979
rect 2690 13923 4040 13979
rect 4096 13923 4106 13979
rect 2520 13875 4106 13923
rect 2520 13819 2530 13875
rect 2586 13819 2634 13875
rect 2690 13819 4040 13875
rect 4096 13819 4106 13875
rect 2520 13809 2700 13819
rect 4030 13809 4106 13819
rect 4190 13979 4266 13989
rect 4831 13979 4907 13989
rect 6003 13979 6183 13989
rect 7055 13979 7131 13989
rect 7695 13979 7771 13989
rect 4190 13923 4200 13979
rect 4256 13923 4841 13979
rect 4897 13923 6013 13979
rect 6069 13923 6117 13979
rect 6173 13923 7065 13979
rect 7121 13923 7705 13979
rect 7761 13923 7771 13979
rect 4190 13875 7771 13923
rect 4190 13819 4200 13875
rect 4256 13819 4841 13875
rect 4897 13819 6013 13875
rect 6069 13819 6117 13875
rect 6173 13819 7065 13875
rect 7121 13819 7705 13875
rect 7761 13819 7771 13875
rect 4190 13809 4266 13819
rect 4831 13809 4907 13819
rect 6003 13809 6183 13819
rect 7055 13809 7131 13819
rect 7695 13809 7771 13819
rect 374 13763 1084 13795
rect 374 13707 554 13763
rect 610 13707 664 13763
rect 720 13707 774 13763
rect 830 13707 884 13763
rect 940 13707 994 13763
rect 1050 13707 1084 13763
rect 374 13653 1084 13707
rect 374 13597 554 13653
rect 610 13597 664 13653
rect 720 13597 774 13653
rect 830 13597 884 13653
rect 940 13597 994 13653
rect 1050 13597 1084 13653
rect 374 13509 1084 13597
rect 527 13497 1084 13509
rect 3870 13483 3946 13493
rect 4510 13483 4586 13493
rect 5150 13483 5226 13493
rect 5731 13483 5911 13493
rect 3870 13427 3880 13483
rect 3936 13427 4520 13483
rect 4576 13427 5160 13483
rect 5216 13427 5741 13483
rect 5797 13427 5845 13483
rect 5901 13427 5911 13483
rect 3870 13379 5911 13427
rect 7055 13379 7131 13389
rect 7695 13379 7771 13389
rect 3870 13323 3880 13379
rect 3936 13323 4520 13379
rect 4576 13323 5160 13379
rect 5216 13323 5741 13379
rect 5797 13323 5845 13379
rect 5901 13323 7065 13379
rect 7121 13323 7705 13379
rect 7761 13323 7771 13379
rect 3870 13313 3946 13323
rect 4510 13313 4586 13323
rect 5150 13313 5226 13323
rect 5731 13275 7771 13323
rect 5731 13219 5741 13275
rect 5797 13219 5845 13275
rect 5901 13219 7065 13275
rect 7121 13219 7705 13275
rect 7761 13219 7771 13275
rect 2881 13200 3061 13210
rect 3950 13200 4026 13210
rect 5731 13209 5911 13219
rect 7055 13209 7131 13219
rect 7695 13209 7771 13219
rect 2881 13144 2891 13200
rect 2947 13144 2995 13200
rect 3051 13144 3960 13200
rect 4016 13144 4026 13200
rect 2881 13096 4026 13144
rect -8178 13055 -7966 13067
rect -8178 12999 -8163 13055
rect -8107 12999 -8053 13055
rect -7997 12999 -7966 13055
rect 2881 13040 2891 13096
rect 2947 13040 2995 13096
rect 3051 13040 3960 13096
rect 4016 13040 4026 13096
rect 2881 13030 3061 13040
rect 3950 13030 4026 13040
rect 8788 13105 9208 14488
rect 11639 13459 11819 13469
rect 11639 13403 11649 13459
rect 11705 13403 11753 13459
rect 11809 13417 11819 13459
rect 11809 13407 19141 13417
rect 11809 13403 17651 13407
rect 11639 13355 17651 13403
rect 11639 13299 11649 13355
rect 11705 13299 11753 13355
rect 11809 13351 17651 13355
rect 17707 13351 19075 13407
rect 19131 13351 19141 13407
rect 11809 13341 19141 13351
rect 20185 13407 24293 13417
rect 20185 13351 20195 13407
rect 20251 13351 24227 13407
rect 24283 13351 24293 13407
rect 20185 13341 24293 13351
rect 25337 13407 28262 13417
rect 25337 13351 25347 13407
rect 25403 13351 26771 13407
rect 26828 13351 28196 13407
rect 28252 13351 28262 13407
rect 25337 13341 28262 13351
rect 11809 13299 11819 13341
rect 11639 13289 11819 13299
rect 19305 13270 25173 13280
rect 19305 13214 22107 13270
rect 22163 13214 22211 13270
rect 22267 13214 22315 13270
rect 22371 13214 25173 13270
rect 19305 13166 25173 13214
rect 19305 13110 19315 13166
rect 19371 13110 19955 13166
rect 20011 13110 22107 13166
rect 22163 13110 22211 13166
rect 22267 13110 22315 13166
rect 22371 13110 24467 13166
rect 24523 13110 25107 13166
rect 25163 13110 25173 13166
rect -8178 12945 -7966 12999
rect -8178 12889 -8163 12945
rect -8107 12889 -8053 12945
rect -7997 12889 -7966 12945
rect -8178 12855 -7966 12889
rect 6003 13000 6183 13010
rect 6735 13000 6811 13010
rect 7375 13000 7451 13010
rect 8015 13000 8091 13010
rect 6003 12944 6013 13000
rect 6069 12944 6117 13000
rect 6173 12944 6745 13000
rect 6801 12944 7385 13000
rect 7441 12944 8025 13000
rect 8081 12944 8091 13000
rect 6003 12896 8091 12944
rect 2520 12849 2700 12859
rect 4030 12849 4106 12859
rect 2520 12793 2530 12849
rect 2586 12793 2634 12849
rect 2690 12793 4040 12849
rect 4096 12793 4106 12849
rect 2520 12745 4106 12793
rect 2520 12689 2530 12745
rect 2586 12689 2634 12745
rect 2690 12689 4040 12745
rect 4096 12689 4106 12745
rect 2520 12679 2700 12689
rect 4030 12679 4106 12689
rect 4190 12849 4266 12859
rect 4831 12849 4907 12859
rect 5731 12849 5911 12859
rect 4190 12793 4200 12849
rect 4256 12793 4841 12849
rect 4897 12793 5741 12849
rect 5797 12793 5845 12849
rect 5901 12793 5911 12849
rect 6003 12840 6013 12896
rect 6069 12840 6117 12896
rect 6173 12840 6745 12896
rect 6801 12840 7385 12896
rect 7441 12840 8025 12896
rect 8081 12840 8091 12896
rect 6003 12830 6183 12840
rect 6735 12830 6811 12840
rect 7375 12830 7451 12840
rect 8015 12830 8091 12840
rect 8788 12886 18923 13105
rect 19305 13062 25173 13110
rect 19305 13006 19315 13062
rect 19371 13006 19955 13062
rect 20011 13006 22107 13062
rect 22163 13006 22211 13062
rect 22267 13006 22315 13062
rect 22371 13006 24467 13062
rect 24523 13006 25107 13062
rect 25163 13006 25173 13062
rect 19305 12996 25173 13006
rect 28426 13270 31502 13280
rect 28426 13214 31228 13270
rect 31284 13214 31332 13270
rect 31388 13214 31436 13270
rect 31492 13214 31502 13270
rect 28426 13166 31502 13214
rect 28426 13110 28436 13166
rect 28492 13110 29076 13166
rect 29132 13110 31228 13166
rect 31284 13110 31332 13166
rect 31388 13110 31436 13166
rect 31492 13110 31502 13166
rect 28426 13062 31502 13110
rect 28426 13006 28436 13062
rect 28492 13006 29076 13062
rect 29132 13006 31228 13062
rect 31284 13006 31332 13062
rect 31388 13006 31436 13062
rect 31492 13006 31502 13062
rect 28426 12996 31502 13006
rect 34578 13050 67198 13060
rect 34578 12994 34588 13050
rect 34644 12994 34692 13050
rect 34748 12994 34796 13050
rect 34852 12994 38724 13050
rect 38780 12994 38828 13050
rect 38884 12994 38932 13050
rect 38988 12994 44284 13050
rect 44340 12994 44388 13050
rect 44444 12994 44492 13050
rect 44548 12994 48420 13050
rect 48476 12994 48524 13050
rect 48580 12994 48628 13050
rect 48684 12994 53980 13050
rect 54036 12994 54084 13050
rect 54140 12994 54188 13050
rect 54244 12994 58116 13050
rect 58172 12994 58220 13050
rect 58276 12994 58324 13050
rect 58380 12994 63676 13050
rect 63732 12994 63780 13050
rect 63836 12994 63884 13050
rect 63940 12994 66924 13050
rect 66980 12994 67028 13050
rect 67084 12994 67132 13050
rect 67188 12994 67198 13050
rect 34578 12946 67198 12994
rect 34578 12890 34588 12946
rect 34644 12890 34692 12946
rect 34748 12890 34796 12946
rect 34852 12890 38724 12946
rect 38780 12890 38828 12946
rect 38884 12890 38932 12946
rect 38988 12890 44284 12946
rect 44340 12890 44388 12946
rect 44444 12890 44492 12946
rect 44548 12890 48420 12946
rect 48476 12890 48524 12946
rect 48580 12890 48628 12946
rect 48684 12890 53980 12946
rect 54036 12890 54084 12946
rect 54140 12890 54188 12946
rect 54244 12890 58116 12946
rect 58172 12890 58220 12946
rect 58276 12890 58324 12946
rect 58380 12890 63676 12946
rect 63732 12890 63780 12946
rect 63836 12890 63884 12946
rect 63940 12890 66924 12946
rect 66980 12890 67028 12946
rect 67084 12890 67132 12946
rect 67188 12890 67198 12946
rect 8788 12876 32410 12886
rect 4190 12745 5911 12793
rect 4190 12689 4200 12745
rect 4256 12689 4841 12745
rect 4897 12689 5741 12745
rect 5797 12689 5845 12745
rect 5901 12689 5911 12745
rect 4190 12679 4266 12689
rect 4831 12679 4907 12689
rect 5731 12679 5911 12689
rect 8788 12820 21458 12876
rect 21514 12820 21562 12876
rect 21618 12820 21666 12876
rect 21722 12820 22756 12876
rect 22812 12820 22860 12876
rect 22916 12820 22964 12876
rect 23020 12820 30579 12876
rect 30635 12820 30683 12876
rect 30739 12820 30787 12876
rect 30843 12820 32136 12876
rect 32192 12820 32240 12876
rect 32296 12820 32344 12876
rect 32400 12820 32410 12876
rect 8788 12772 32410 12820
rect 34578 12842 67198 12890
rect 34578 12786 34588 12842
rect 34644 12786 34692 12842
rect 34748 12786 34796 12842
rect 34852 12786 38724 12842
rect 38780 12786 38828 12842
rect 38884 12786 38932 12842
rect 38988 12786 44284 12842
rect 44340 12786 44388 12842
rect 44444 12786 44492 12842
rect 44548 12786 48420 12842
rect 48476 12786 48524 12842
rect 48580 12786 48628 12842
rect 48684 12786 53980 12842
rect 54036 12786 54084 12842
rect 54140 12786 54188 12842
rect 54244 12786 58116 12842
rect 58172 12786 58220 12842
rect 58276 12786 58324 12842
rect 58380 12786 63676 12842
rect 63732 12786 63780 12842
rect 63836 12786 63884 12842
rect 63940 12786 66924 12842
rect 66980 12786 67028 12842
rect 67084 12786 67132 12842
rect 67188 12786 67198 12842
rect 34578 12776 67198 12786
rect 8788 12716 18995 12772
rect 19051 12716 19635 12772
rect 19691 12716 20275 12772
rect 20331 12716 21458 12772
rect 21514 12716 21562 12772
rect 21618 12716 21666 12772
rect 21722 12716 22756 12772
rect 22812 12716 22860 12772
rect 22916 12716 22964 12772
rect 23020 12716 24147 12772
rect 24203 12716 24787 12772
rect 24843 12716 25427 12772
rect 25483 12716 28116 12772
rect 28172 12716 28756 12772
rect 28812 12716 29396 12772
rect 29452 12716 30579 12772
rect 30635 12716 30683 12772
rect 30739 12716 30787 12772
rect 30843 12716 32136 12772
rect 32192 12716 32240 12772
rect 32296 12716 32344 12772
rect 32400 12716 32410 12772
rect 8788 12668 32410 12716
rect 8788 12612 18995 12668
rect 19051 12612 19635 12668
rect 19691 12612 20275 12668
rect 20331 12612 21458 12668
rect 21514 12612 21562 12668
rect 21618 12612 21666 12668
rect 21722 12612 22756 12668
rect 22812 12612 22860 12668
rect 22916 12612 22964 12668
rect 23020 12612 24147 12668
rect 24203 12612 24787 12668
rect 24843 12612 25427 12668
rect 25483 12612 28116 12668
rect 28172 12612 28756 12668
rect 28812 12612 29396 12668
rect 29452 12612 30579 12668
rect 30635 12612 30683 12668
rect 30739 12612 30787 12668
rect 30843 12612 32136 12668
rect 32192 12612 32240 12668
rect 32296 12612 32344 12668
rect 32400 12612 32410 12668
rect 8788 12602 32410 12612
rect 11371 12493 11551 12503
rect 3870 12457 3946 12467
rect 4510 12457 4586 12467
rect 5150 12457 5226 12467
rect 6003 12457 6183 12467
rect 7055 12457 7131 12467
rect 7695 12457 7771 12467
rect 3870 12401 3880 12457
rect 3936 12401 4520 12457
rect 4576 12401 5160 12457
rect 5216 12401 6013 12457
rect 6069 12401 6117 12457
rect 6173 12401 7065 12457
rect 7121 12401 7705 12457
rect 7761 12401 7771 12457
rect 3870 12353 7771 12401
rect -10442 12259 -10354 12347
rect 3870 12297 3880 12353
rect 3936 12297 4520 12353
rect 4576 12297 5160 12353
rect 5216 12297 6013 12353
rect 6069 12297 6117 12353
rect 6173 12297 7065 12353
rect 7121 12297 7705 12353
rect 7761 12297 7771 12353
rect 11371 12437 11381 12493
rect 11437 12437 11485 12493
rect 11541 12451 11551 12493
rect 11541 12441 19141 12451
rect 11541 12437 17851 12441
rect 11371 12389 17851 12437
rect 11371 12333 11381 12389
rect 11437 12333 11485 12389
rect 11541 12385 17851 12389
rect 17907 12385 19075 12441
rect 19131 12385 19141 12441
rect 11541 12375 19141 12385
rect 25337 12441 28262 12451
rect 25337 12385 25347 12441
rect 25403 12385 26571 12441
rect 26627 12385 26972 12441
rect 27028 12385 28196 12441
rect 28252 12385 28262 12441
rect 25337 12375 28262 12385
rect 11541 12333 11551 12375
rect 11371 12323 11551 12333
rect 19305 12334 25173 12344
rect 3870 12287 3946 12297
rect 4510 12287 4586 12297
rect 5150 12287 5226 12297
rect 6003 12287 6183 12297
rect 7055 12287 7131 12297
rect 7695 12287 7771 12297
rect 19305 12278 21458 12334
rect 21514 12278 21562 12334
rect 21618 12278 21666 12334
rect 21722 12278 22756 12334
rect 22812 12278 22860 12334
rect 22916 12278 22964 12334
rect 23020 12278 25173 12334
rect 19305 12230 25173 12278
rect 19305 12174 19315 12230
rect 19371 12174 19955 12230
rect 20011 12174 21458 12230
rect 21514 12174 21562 12230
rect 21618 12174 21666 12230
rect 21722 12174 22756 12230
rect 22812 12174 22860 12230
rect 22916 12174 22964 12230
rect 23020 12174 24467 12230
rect 24523 12174 25107 12230
rect 25163 12174 25173 12230
rect 5731 12138 5911 12148
rect 6735 12138 6811 12148
rect 7375 12138 7451 12148
rect 8015 12138 8091 12148
rect 5731 12082 5741 12138
rect 5797 12082 5845 12138
rect 5901 12082 6745 12138
rect 6801 12082 7385 12138
rect 7441 12082 8025 12138
rect 8081 12082 8091 12138
rect 3161 12070 3341 12080
rect 3950 12070 4026 12080
rect 3161 12014 3171 12070
rect 3227 12014 3275 12070
rect 3331 12014 3960 12070
rect 4016 12014 4026 12070
rect 3161 11966 4026 12014
rect 5731 12034 8091 12082
rect 19305 12126 25173 12174
rect 19305 12070 19315 12126
rect 19371 12070 19955 12126
rect 20011 12070 21458 12126
rect 21514 12070 21562 12126
rect 21618 12070 21666 12126
rect 21722 12070 22756 12126
rect 22812 12070 22860 12126
rect 22916 12070 22964 12126
rect 23020 12070 24467 12126
rect 24523 12070 25107 12126
rect 25163 12070 25173 12126
rect 19305 12060 25173 12070
rect 28426 12334 32410 12344
rect 28426 12278 30579 12334
rect 30635 12278 30683 12334
rect 30739 12278 30787 12334
rect 30843 12278 32136 12334
rect 32192 12278 32240 12334
rect 32296 12278 32344 12334
rect 32400 12278 32410 12334
rect 28426 12230 32410 12278
rect 28426 12174 28436 12230
rect 28492 12174 29076 12230
rect 29132 12174 30579 12230
rect 30635 12174 30683 12230
rect 30739 12174 30787 12230
rect 30843 12174 32136 12230
rect 32192 12174 32240 12230
rect 32296 12174 32344 12230
rect 32400 12174 32410 12230
rect 28426 12126 32410 12174
rect 28426 12070 28436 12126
rect 28492 12070 29076 12126
rect 29132 12070 30579 12126
rect 30635 12070 30683 12126
rect 30739 12070 30787 12126
rect 30843 12070 32136 12126
rect 32192 12070 32240 12126
rect 32296 12070 32344 12126
rect 32400 12070 32410 12126
rect 28426 12060 32410 12070
rect 5731 11978 5741 12034
rect 5797 11978 5845 12034
rect 5901 11978 6745 12034
rect 6801 11978 7385 12034
rect 7441 11978 8025 12034
rect 8081 11978 8091 12034
rect 5731 11968 5911 11978
rect 6735 11968 6811 11978
rect 7375 11968 7451 11978
rect 8015 11968 8091 11978
rect 3161 11910 3171 11966
rect 3227 11910 3275 11966
rect 3331 11910 3960 11966
rect 4016 11910 4026 11966
rect 3161 11900 3341 11910
rect 3950 11900 4026 11910
rect 18985 11940 32030 11950
rect 18985 11884 22107 11940
rect 22163 11884 22211 11940
rect 22267 11884 22315 11940
rect 22371 11884 31228 11940
rect 31284 11884 31332 11940
rect 31388 11884 31436 11940
rect 31492 11884 32030 11940
rect 18985 11836 32030 11884
rect 18985 11780 18995 11836
rect 19051 11780 19635 11836
rect 19691 11780 20275 11836
rect 20331 11780 22107 11836
rect 22163 11780 22211 11836
rect 22267 11780 22315 11836
rect 22371 11780 24147 11836
rect 24203 11780 24787 11836
rect 24843 11780 25427 11836
rect 25483 11780 28116 11836
rect 28172 11780 28756 11836
rect 28812 11780 29396 11836
rect 29452 11780 31228 11836
rect 31284 11780 31332 11836
rect 31388 11780 31436 11836
rect 31492 11780 32030 11836
rect 18985 11770 64807 11780
rect 18985 11732 31756 11770
rect 4190 11719 4266 11729
rect 4831 11719 4907 11729
rect 6003 11719 6183 11729
rect 4190 11663 4200 11719
rect 4256 11663 4841 11719
rect 4897 11663 6013 11719
rect 6069 11663 6117 11719
rect 6173 11663 6183 11719
rect 18985 11676 18995 11732
rect 19051 11676 19635 11732
rect 19691 11676 20275 11732
rect 20331 11676 22107 11732
rect 22163 11676 22211 11732
rect 22267 11676 22315 11732
rect 22371 11676 24147 11732
rect 24203 11676 24787 11732
rect 24843 11676 25427 11732
rect 25483 11676 28116 11732
rect 28172 11676 28756 11732
rect 28812 11676 29396 11732
rect 29452 11676 31228 11732
rect 31284 11676 31332 11732
rect 31388 11676 31436 11732
rect 31492 11714 31756 11732
rect 31812 11714 31860 11770
rect 31916 11714 31964 11770
rect 32020 11714 41483 11770
rect 41539 11714 41587 11770
rect 41643 11714 41691 11770
rect 41747 11714 51138 11770
rect 51194 11714 51242 11770
rect 51298 11714 51346 11770
rect 51402 11714 60919 11770
rect 60975 11714 61023 11770
rect 61079 11714 61127 11770
rect 61183 11714 64807 11770
rect 31492 11676 64807 11714
rect 18985 11666 64807 11676
rect 4190 11615 6183 11663
rect 6735 11615 6811 11625
rect 7375 11615 7451 11625
rect 8015 11615 8091 11625
rect 4190 11559 4200 11615
rect 4256 11559 4841 11615
rect 4897 11559 6013 11615
rect 6069 11559 6117 11615
rect 6173 11559 6745 11615
rect 6801 11559 7385 11615
rect 7441 11559 8025 11615
rect 8081 11559 8091 11615
rect 4190 11549 4266 11559
rect 4831 11549 4907 11559
rect 6003 11511 8091 11559
rect 31746 11610 31756 11666
rect 31812 11610 31860 11666
rect 31916 11610 31964 11666
rect 32020 11610 33733 11666
rect 33789 11610 34373 11666
rect 34429 11610 35013 11666
rect 35069 11610 35653 11666
rect 35709 11610 37867 11666
rect 37923 11610 38507 11666
rect 38563 11610 39147 11666
rect 39203 11610 39787 11666
rect 39843 11610 41483 11666
rect 41539 11610 41587 11666
rect 41643 11610 41691 11666
rect 41747 11610 43429 11666
rect 43485 11610 44069 11666
rect 44125 11610 44709 11666
rect 44765 11610 45349 11666
rect 45405 11610 47563 11666
rect 47619 11610 48203 11666
rect 48259 11610 48843 11666
rect 48899 11610 49483 11666
rect 49539 11610 51138 11666
rect 51194 11610 51242 11666
rect 51298 11610 51346 11666
rect 51402 11610 53125 11666
rect 53181 11610 53765 11666
rect 53821 11610 54405 11666
rect 54461 11610 55045 11666
rect 55101 11610 57259 11666
rect 57315 11610 57899 11666
rect 57955 11610 58539 11666
rect 58595 11610 59179 11666
rect 59235 11610 60919 11666
rect 60975 11610 61023 11666
rect 61079 11610 61127 11666
rect 61183 11610 62821 11666
rect 62877 11610 63461 11666
rect 63517 11610 64101 11666
rect 64157 11610 64741 11666
rect 64797 11610 64807 11666
rect 31746 11562 64807 11610
rect 6003 11455 6013 11511
rect 6069 11455 6117 11511
rect 6173 11455 6745 11511
rect 6801 11455 7385 11511
rect 7441 11455 8025 11511
rect 8081 11455 8091 11511
rect 6003 11445 6183 11455
rect 6735 11445 6811 11455
rect 7375 11445 7451 11455
rect 8015 11445 8091 11455
rect 17641 11505 19141 11515
rect 17641 11449 17651 11505
rect 17707 11449 19075 11505
rect 19131 11449 19141 11505
rect 17641 11439 19141 11449
rect 25337 11505 28262 11515
rect 25337 11449 25347 11505
rect 25403 11449 26771 11505
rect 26828 11449 28196 11505
rect 28252 11449 28262 11505
rect 31746 11506 31756 11562
rect 31812 11506 31860 11562
rect 31916 11506 31964 11562
rect 32020 11506 33733 11562
rect 33789 11506 34373 11562
rect 34429 11506 35013 11562
rect 35069 11506 35653 11562
rect 35709 11506 37867 11562
rect 37923 11506 38507 11562
rect 38563 11506 39147 11562
rect 39203 11506 39787 11562
rect 39843 11506 41483 11562
rect 41539 11506 41587 11562
rect 41643 11506 41691 11562
rect 41747 11506 43429 11562
rect 43485 11506 44069 11562
rect 44125 11506 44709 11562
rect 44765 11506 45349 11562
rect 45405 11506 47563 11562
rect 47619 11506 48203 11562
rect 48259 11506 48843 11562
rect 48899 11506 49483 11562
rect 49539 11506 51138 11562
rect 51194 11506 51242 11562
rect 51298 11506 51346 11562
rect 51402 11506 53125 11562
rect 53181 11506 53765 11562
rect 53821 11506 54405 11562
rect 54461 11506 55045 11562
rect 55101 11506 57259 11562
rect 57315 11506 57899 11562
rect 57955 11506 58539 11562
rect 58595 11506 59179 11562
rect 59235 11506 60919 11562
rect 60975 11506 61023 11562
rect 61079 11506 61127 11562
rect 61183 11506 62821 11562
rect 62877 11506 63461 11562
rect 63517 11506 64101 11562
rect 64157 11506 64741 11562
rect 64797 11506 64807 11562
rect 31746 11496 64807 11506
rect 25337 11439 28262 11449
rect 19305 11398 25173 11408
rect 11371 11375 11551 11385
rect 12800 11375 12876 11385
rect 13696 11375 13772 11385
rect 5731 11327 5911 11337
rect 7055 11327 7131 11337
rect 7695 11327 7771 11337
rect 5731 11271 5741 11327
rect 5797 11271 5845 11327
rect 5901 11271 7065 11327
rect 7121 11271 7705 11327
rect 7761 11271 7771 11327
rect 3870 11223 3946 11233
rect 4510 11223 4586 11233
rect 5150 11223 5226 11233
rect 5731 11223 7771 11271
rect 3870 11167 3880 11223
rect 3936 11167 4520 11223
rect 4576 11167 5160 11223
rect 5216 11167 5741 11223
rect 5797 11167 5845 11223
rect 5901 11167 7065 11223
rect 7121 11167 7705 11223
rect 7761 11167 7771 11223
rect 11371 11319 11381 11375
rect 11437 11319 11485 11375
rect 11541 11319 12810 11375
rect 12866 11319 13706 11375
rect 13762 11319 13772 11375
rect 11371 11271 13772 11319
rect 11371 11215 11381 11271
rect 11437 11215 11485 11271
rect 11541 11215 12810 11271
rect 12866 11215 13706 11271
rect 13762 11215 13772 11271
rect 11371 11205 11551 11215
rect 12800 11205 12876 11215
rect 13696 11205 13772 11215
rect 13984 11375 14060 11385
rect 15146 11375 15222 11385
rect 15786 11375 15862 11385
rect 16426 11375 16502 11385
rect 17365 11375 17545 11385
rect 13984 11319 13994 11375
rect 14050 11319 15156 11375
rect 15212 11319 15796 11375
rect 15852 11319 16436 11375
rect 16492 11319 17375 11375
rect 17431 11319 17479 11375
rect 17535 11319 17545 11375
rect 13984 11271 17545 11319
rect 13984 11215 13994 11271
rect 14050 11215 15156 11271
rect 15212 11215 15796 11271
rect 15852 11215 16436 11271
rect 16492 11215 17375 11271
rect 17431 11215 17479 11271
rect 17535 11215 17545 11271
rect 13984 11205 14060 11215
rect 15146 11205 15222 11215
rect 15786 11205 15862 11215
rect 16426 11205 16502 11215
rect 17365 11205 17545 11215
rect 19305 11342 22107 11398
rect 22163 11342 22211 11398
rect 22267 11342 22315 11398
rect 22371 11342 25173 11398
rect 19305 11294 25173 11342
rect 19305 11238 19315 11294
rect 19371 11238 19955 11294
rect 20011 11238 22107 11294
rect 22163 11238 22211 11294
rect 22267 11238 22315 11294
rect 22371 11238 24467 11294
rect 24523 11238 25107 11294
rect 25163 11238 25173 11294
rect 3870 11119 5911 11167
rect 7055 11157 7131 11167
rect 7695 11157 7771 11167
rect 19305 11190 25173 11238
rect 19305 11134 19315 11190
rect 19371 11134 19955 11190
rect 20011 11134 22107 11190
rect 22163 11134 22211 11190
rect 22267 11134 22315 11190
rect 22371 11134 24467 11190
rect 24523 11134 25107 11190
rect 25163 11134 25173 11190
rect 19305 11124 25173 11134
rect 28426 11398 31502 11408
rect 28426 11342 31228 11398
rect 31284 11342 31332 11398
rect 31388 11342 31436 11398
rect 31492 11342 31502 11398
rect 28426 11294 31502 11342
rect 28426 11238 28436 11294
rect 28492 11238 29076 11294
rect 29132 11238 31228 11294
rect 31284 11238 31332 11294
rect 31388 11238 31436 11294
rect 31492 11238 31502 11294
rect 28426 11190 31502 11238
rect 28426 11134 28436 11190
rect 28492 11134 29076 11190
rect 29132 11134 31228 11190
rect 31284 11134 31332 11190
rect 31388 11134 31436 11190
rect 31492 11134 31502 11190
rect 28426 11124 31502 11134
rect 32126 11376 65126 11386
rect 32126 11320 32136 11376
rect 32192 11320 32240 11376
rect 32296 11320 32344 11376
rect 32400 11320 41122 11376
rect 41178 11320 41226 11376
rect 41282 11320 41330 11376
rect 41386 11320 41842 11376
rect 41898 11320 41946 11376
rect 42002 11320 42050 11376
rect 42106 11320 50798 11376
rect 50854 11320 50902 11376
rect 50958 11320 51006 11376
rect 51062 11320 51530 11376
rect 51586 11320 51634 11376
rect 51690 11320 51738 11376
rect 51794 11320 60514 11376
rect 60570 11320 60618 11376
rect 60674 11320 60722 11376
rect 60778 11320 61278 11376
rect 61334 11320 61382 11376
rect 61438 11320 61486 11376
rect 61542 11320 65126 11376
rect 32126 11272 65126 11320
rect 32126 11216 32136 11272
rect 32192 11216 32240 11272
rect 32296 11216 32344 11272
rect 32400 11216 33412 11272
rect 33468 11216 34052 11272
rect 34108 11216 35332 11272
rect 35388 11216 35972 11272
rect 36028 11216 37548 11272
rect 37604 11216 38188 11272
rect 38244 11216 39468 11272
rect 39524 11216 40108 11272
rect 40164 11216 41122 11272
rect 41178 11216 41226 11272
rect 41282 11216 41330 11272
rect 41386 11216 41842 11272
rect 41898 11216 41946 11272
rect 42002 11216 42050 11272
rect 42106 11216 43108 11272
rect 43164 11216 43748 11272
rect 43804 11216 45028 11272
rect 45084 11216 45668 11272
rect 45724 11216 47244 11272
rect 47300 11216 47884 11272
rect 47940 11216 49164 11272
rect 49220 11216 49804 11272
rect 49860 11216 50798 11272
rect 50854 11216 50902 11272
rect 50958 11216 51006 11272
rect 51062 11216 51530 11272
rect 51586 11216 51634 11272
rect 51690 11216 51738 11272
rect 51794 11216 52804 11272
rect 52860 11216 53444 11272
rect 53500 11216 54724 11272
rect 54780 11216 55364 11272
rect 55420 11216 56940 11272
rect 56996 11216 57580 11272
rect 57636 11216 58860 11272
rect 58916 11216 59500 11272
rect 59556 11216 60514 11272
rect 60570 11216 60618 11272
rect 60674 11216 60722 11272
rect 60778 11216 61278 11272
rect 61334 11216 61382 11272
rect 61438 11216 61486 11272
rect 61542 11216 62500 11272
rect 62556 11216 63140 11272
rect 63196 11216 64420 11272
rect 64476 11216 65060 11272
rect 65116 11216 65126 11272
rect 32126 11168 65126 11216
rect 3870 11063 3880 11119
rect 3936 11063 4520 11119
rect 4576 11063 5160 11119
rect 5216 11063 5741 11119
rect 5797 11063 5845 11119
rect 5901 11063 5911 11119
rect 32126 11112 32136 11168
rect 32192 11112 32240 11168
rect 32296 11112 32344 11168
rect 32400 11112 33412 11168
rect 33468 11112 34052 11168
rect 34108 11112 35332 11168
rect 35388 11112 35972 11168
rect 36028 11112 37548 11168
rect 37604 11112 38188 11168
rect 38244 11112 39468 11168
rect 39524 11112 40108 11168
rect 40164 11112 41122 11168
rect 41178 11112 41226 11168
rect 41282 11112 41330 11168
rect 41386 11112 41842 11168
rect 41898 11112 41946 11168
rect 42002 11112 42050 11168
rect 42106 11112 43108 11168
rect 43164 11112 43748 11168
rect 43804 11112 45028 11168
rect 45084 11112 45668 11168
rect 45724 11112 47244 11168
rect 47300 11112 47884 11168
rect 47940 11112 49164 11168
rect 49220 11112 49804 11168
rect 49860 11112 50798 11168
rect 50854 11112 50902 11168
rect 50958 11112 51006 11168
rect 51062 11112 51530 11168
rect 51586 11112 51634 11168
rect 51690 11112 51738 11168
rect 51794 11112 52804 11168
rect 52860 11112 53444 11168
rect 53500 11112 54724 11168
rect 54780 11112 55364 11168
rect 55420 11112 56940 11168
rect 56996 11112 57580 11168
rect 57636 11112 58860 11168
rect 58916 11112 59500 11168
rect 59556 11112 60514 11168
rect 60570 11112 60618 11168
rect 60674 11112 60722 11168
rect 60778 11112 61278 11168
rect 61334 11112 61382 11168
rect 61438 11112 61486 11168
rect 61542 11112 62500 11168
rect 62556 11112 63140 11168
rect 63196 11112 64420 11168
rect 64476 11112 65060 11168
rect 65116 11112 65126 11168
rect 32126 11102 65126 11112
rect 3870 11053 3946 11063
rect 4510 11053 4586 11063
rect 5150 11053 5226 11063
rect 5731 11053 5911 11063
rect 18985 11004 25493 11014
rect 11639 10955 11819 10965
rect 12352 10955 12428 10965
rect 13248 10955 13324 10965
rect 14144 10955 14220 10965
rect 11639 10899 11649 10955
rect 11705 10899 11753 10955
rect 11809 10899 12362 10955
rect 12418 10899 13258 10955
rect 13314 10899 14154 10955
rect 14210 10899 14220 10955
rect 11639 10851 14220 10899
rect 5731 10796 5911 10806
rect 8970 10796 9046 10806
rect 9866 10796 9942 10806
rect 10762 10796 10838 10806
rect -3626 10729 -3414 10752
rect -3626 10673 -3604 10729
rect -3548 10673 -3494 10729
rect -3438 10673 -3414 10729
rect -3626 10619 -3414 10673
rect 5731 10740 5741 10796
rect 5797 10740 5845 10796
rect 5901 10740 8980 10796
rect 9036 10740 9876 10796
rect 9932 10740 10772 10796
rect 10828 10740 10838 10796
rect 11639 10795 11649 10851
rect 11705 10795 11753 10851
rect 11809 10795 12362 10851
rect 12418 10795 13258 10851
rect 13314 10795 14154 10851
rect 14210 10795 14220 10851
rect 11639 10785 11819 10795
rect 12352 10785 12428 10795
rect 13248 10785 13324 10795
rect 14144 10785 14220 10795
rect 15466 10955 15542 10965
rect 16106 10955 16182 10965
rect 17103 10955 17283 10965
rect 15466 10899 15476 10955
rect 15532 10899 16116 10955
rect 16172 10899 17113 10955
rect 17169 10899 17217 10955
rect 17273 10899 17283 10955
rect 15466 10851 17283 10899
rect 15466 10795 15476 10851
rect 15532 10795 16116 10851
rect 16172 10795 17113 10851
rect 17169 10795 17217 10851
rect 17273 10795 17283 10851
rect 15466 10785 15542 10795
rect 16106 10785 16182 10795
rect 17103 10785 17283 10795
rect 18985 10948 21458 11004
rect 21514 10948 21562 11004
rect 21618 10948 21666 11004
rect 21722 10948 22756 11004
rect 22812 10948 22860 11004
rect 22916 10948 22964 11004
rect 23020 10948 25493 11004
rect 18985 10900 25493 10948
rect 18985 10844 18995 10900
rect 19051 10844 19635 10900
rect 19691 10844 20275 10900
rect 20331 10844 21458 10900
rect 21514 10844 21562 10900
rect 21618 10844 21666 10900
rect 21722 10844 22756 10900
rect 22812 10844 22860 10900
rect 22916 10844 22964 10900
rect 23020 10844 24147 10900
rect 24203 10844 24787 10900
rect 24843 10844 25427 10900
rect 25483 10844 25493 10900
rect 18985 10796 25493 10844
rect 5731 10692 10838 10740
rect 18985 10740 18995 10796
rect 19051 10740 19635 10796
rect 19691 10740 20275 10796
rect 20331 10740 21458 10796
rect 21514 10740 21562 10796
rect 21618 10740 21666 10796
rect 21722 10740 22756 10796
rect 22812 10740 22860 10796
rect 22916 10740 22964 10796
rect 23020 10740 24147 10796
rect 24203 10740 24787 10796
rect 24843 10740 25427 10796
rect 25483 10740 25493 10796
rect 18985 10730 25493 10740
rect 28106 11004 30853 11014
rect 28106 10948 30579 11004
rect 30635 10948 30683 11004
rect 30739 10948 30787 11004
rect 30843 10948 30853 11004
rect 28106 10900 30853 10948
rect 28106 10844 28116 10900
rect 28172 10844 28756 10900
rect 28812 10844 29396 10900
rect 29452 10844 30579 10900
rect 30635 10844 30683 10900
rect 30739 10844 30787 10900
rect 30843 10844 30853 10900
rect 28106 10796 30853 10844
rect 28106 10740 28116 10796
rect 28172 10740 28756 10796
rect 28812 10740 29396 10796
rect 29452 10740 30579 10796
rect 30635 10740 30683 10796
rect 30739 10740 30787 10796
rect 30843 10740 30853 10796
rect 28106 10730 30853 10740
rect 5731 10636 5741 10692
rect 5797 10636 5845 10692
rect 5901 10636 8980 10692
rect 9036 10636 9876 10692
rect 9932 10636 10772 10692
rect 10828 10636 10838 10692
rect 5731 10626 5911 10636
rect 8970 10626 9046 10636
rect 9866 10626 9942 10636
rect 10762 10626 10838 10636
rect 32126 10710 64807 10720
rect 32126 10654 32136 10710
rect 32192 10654 32240 10710
rect 32296 10654 32344 10710
rect 32400 10654 41122 10710
rect 41178 10654 41226 10710
rect 41282 10654 41330 10710
rect 41386 10654 41842 10710
rect 41898 10654 41946 10710
rect 42002 10654 42050 10710
rect 42106 10654 50798 10710
rect 50854 10654 50902 10710
rect 50958 10654 51006 10710
rect 51062 10654 51530 10710
rect 51586 10654 51634 10710
rect 51690 10654 51738 10710
rect 51794 10654 60514 10710
rect 60570 10654 60618 10710
rect 60674 10654 60722 10710
rect 60778 10654 61278 10710
rect 61334 10654 61382 10710
rect 61438 10654 61486 10710
rect 61542 10654 64807 10710
rect -3626 10563 -3604 10619
rect -3548 10563 -3494 10619
rect -3438 10563 -3414 10619
rect -3626 10540 -3414 10563
rect 32126 10606 64807 10654
rect 32126 10550 32136 10606
rect 32192 10550 32240 10606
rect 32296 10550 32344 10606
rect 32400 10550 33733 10606
rect 33789 10550 34373 10606
rect 34429 10550 35013 10606
rect 35069 10550 35653 10606
rect 35709 10550 37867 10606
rect 37923 10550 38507 10606
rect 38563 10550 39147 10606
rect 39203 10550 39787 10606
rect 39843 10550 41122 10606
rect 41178 10550 41226 10606
rect 41282 10550 41330 10606
rect 41386 10550 41842 10606
rect 41898 10550 41946 10606
rect 42002 10550 42050 10606
rect 42106 10550 43429 10606
rect 43485 10550 44069 10606
rect 44125 10550 44709 10606
rect 44765 10550 45349 10606
rect 45405 10550 47563 10606
rect 47619 10550 48203 10606
rect 48259 10550 48843 10606
rect 48899 10550 49483 10606
rect 49539 10550 50798 10606
rect 50854 10550 50902 10606
rect 50958 10550 51006 10606
rect 51062 10550 51530 10606
rect 51586 10550 51634 10606
rect 51690 10550 51738 10606
rect 51794 10550 53125 10606
rect 53181 10550 53765 10606
rect 53821 10550 54405 10606
rect 54461 10550 55045 10606
rect 55101 10550 57259 10606
rect 57315 10550 57899 10606
rect 57955 10550 58539 10606
rect 58595 10550 59179 10606
rect 59235 10550 60514 10606
rect 60570 10550 60618 10606
rect 60674 10550 60722 10606
rect 60778 10550 61278 10606
rect 61334 10550 61382 10606
rect 61438 10550 61486 10606
rect 61542 10550 62821 10606
rect 62877 10550 63461 10606
rect 63517 10550 64101 10606
rect 64157 10550 64741 10606
rect 64797 10550 64807 10606
rect 32126 10502 64807 10550
rect 19305 10462 32030 10472
rect 6003 10425 6183 10435
rect 9418 10425 9494 10435
rect 10314 10425 10390 10435
rect 6003 10369 6013 10425
rect 6069 10369 6117 10425
rect 6173 10369 9428 10425
rect 9484 10369 10324 10425
rect 10380 10369 10390 10425
rect 2520 10325 2700 10335
rect 4030 10325 4106 10335
rect 2520 10269 2530 10325
rect 2586 10269 2634 10325
rect 2690 10269 4040 10325
rect 4096 10269 4106 10325
rect 2520 10221 4106 10269
rect 6003 10321 10390 10369
rect 6003 10265 6013 10321
rect 6069 10265 6117 10321
rect 6173 10265 9428 10321
rect 9484 10265 10324 10321
rect 10380 10265 10390 10321
rect 6003 10255 6183 10265
rect 9418 10255 9494 10265
rect 10314 10255 10390 10265
rect 10602 10425 10678 10435
rect 11639 10425 11819 10435
rect 10602 10369 10612 10425
rect 10668 10369 11649 10425
rect 11705 10369 11753 10425
rect 11809 10369 11819 10425
rect 10602 10321 11819 10369
rect 19305 10406 22107 10462
rect 22163 10406 22211 10462
rect 22267 10406 22315 10462
rect 22371 10406 31228 10462
rect 31284 10406 31332 10462
rect 31388 10406 31436 10462
rect 31492 10406 32030 10462
rect 32126 10446 32136 10502
rect 32192 10446 32240 10502
rect 32296 10446 32344 10502
rect 32400 10446 33733 10502
rect 33789 10446 34373 10502
rect 34429 10446 35013 10502
rect 35069 10446 35653 10502
rect 35709 10446 37867 10502
rect 37923 10446 38507 10502
rect 38563 10446 39147 10502
rect 39203 10446 39787 10502
rect 39843 10446 41122 10502
rect 41178 10446 41226 10502
rect 41282 10446 41330 10502
rect 41386 10446 41842 10502
rect 41898 10446 41946 10502
rect 42002 10446 42050 10502
rect 42106 10446 43429 10502
rect 43485 10446 44069 10502
rect 44125 10446 44709 10502
rect 44765 10446 45349 10502
rect 45405 10446 47563 10502
rect 47619 10446 48203 10502
rect 48259 10446 48843 10502
rect 48899 10446 49483 10502
rect 49539 10446 50798 10502
rect 50854 10446 50902 10502
rect 50958 10446 51006 10502
rect 51062 10446 51530 10502
rect 51586 10446 51634 10502
rect 51690 10446 51738 10502
rect 51794 10446 53125 10502
rect 53181 10446 53765 10502
rect 53821 10446 54405 10502
rect 54461 10446 55045 10502
rect 55101 10446 57259 10502
rect 57315 10446 57899 10502
rect 57955 10446 58539 10502
rect 58595 10446 59179 10502
rect 59235 10446 60514 10502
rect 60570 10446 60618 10502
rect 60674 10446 60722 10502
rect 60778 10446 61278 10502
rect 61334 10446 61382 10502
rect 61438 10446 61486 10502
rect 61542 10446 62821 10502
rect 62877 10446 63461 10502
rect 63517 10446 64101 10502
rect 64157 10446 64741 10502
rect 64797 10446 64807 10502
rect 32126 10436 64807 10446
rect 19305 10358 32030 10406
rect 12800 10321 12876 10331
rect 13696 10321 13772 10331
rect 10602 10265 10612 10321
rect 10668 10265 11649 10321
rect 11705 10265 11753 10321
rect 11809 10265 12810 10321
rect 12866 10265 13706 10321
rect 13762 10265 13772 10321
rect 10602 10255 10678 10265
rect 2520 10165 2530 10221
rect 2586 10165 2634 10221
rect 2690 10165 4040 10221
rect 4096 10165 4106 10221
rect 2520 10155 2700 10165
rect 4030 10155 4106 10165
rect 11639 10217 13772 10265
rect 11639 10161 11649 10217
rect 11705 10161 11753 10217
rect 11809 10161 12810 10217
rect 12866 10161 13706 10217
rect 13762 10161 13772 10217
rect 11639 10151 11819 10161
rect 12800 10151 12876 10161
rect 13696 10151 13772 10161
rect 13984 10295 14060 10305
rect 15146 10295 15222 10305
rect 15786 10295 15862 10305
rect 16426 10295 16502 10305
rect 17103 10295 17283 10305
rect 13984 10239 13994 10295
rect 14050 10239 15156 10295
rect 15212 10239 15796 10295
rect 15852 10239 16436 10295
rect 16492 10239 17113 10295
rect 17169 10239 17217 10295
rect 17273 10239 17283 10295
rect 13984 10191 17283 10239
rect 13984 10135 13994 10191
rect 14050 10135 15156 10191
rect 15212 10135 15796 10191
rect 15852 10135 16436 10191
rect 16492 10135 17113 10191
rect 17169 10135 17217 10191
rect 17273 10135 17283 10191
rect 19305 10302 19315 10358
rect 19371 10302 19955 10358
rect 20011 10302 22107 10358
rect 22163 10302 22211 10358
rect 22267 10302 22315 10358
rect 22371 10302 24467 10358
rect 24523 10302 25107 10358
rect 25163 10302 28436 10358
rect 28492 10302 29076 10358
rect 29132 10302 31228 10358
rect 31284 10302 31332 10358
rect 31388 10302 31436 10358
rect 31492 10326 32030 10358
rect 31492 10316 65126 10326
rect 31492 10302 31756 10316
rect 19305 10260 31756 10302
rect 31812 10260 31860 10316
rect 31916 10260 31964 10316
rect 32020 10260 41483 10316
rect 41539 10260 41587 10316
rect 41643 10260 41691 10316
rect 41747 10260 51138 10316
rect 51194 10260 51242 10316
rect 51298 10260 51346 10316
rect 51402 10260 60919 10316
rect 60975 10260 61023 10316
rect 61079 10260 61127 10316
rect 61183 10260 65126 10316
rect 19305 10254 65126 10260
rect 19305 10198 19315 10254
rect 19371 10198 19955 10254
rect 20011 10198 22107 10254
rect 22163 10198 22211 10254
rect 22267 10198 22315 10254
rect 22371 10198 24467 10254
rect 24523 10198 25107 10254
rect 25163 10198 28436 10254
rect 28492 10198 29076 10254
rect 29132 10198 31228 10254
rect 31284 10198 31332 10254
rect 31388 10198 31436 10254
rect 31492 10212 65126 10254
rect 31492 10198 31756 10212
rect 19305 10188 31756 10198
rect 13984 10125 14060 10135
rect 15146 10125 15222 10135
rect 15786 10125 15862 10135
rect 16426 10125 16502 10135
rect 17103 10125 17283 10135
rect 31746 10156 31756 10188
rect 31812 10156 31860 10212
rect 31916 10156 31964 10212
rect 32020 10156 33412 10212
rect 33468 10156 34052 10212
rect 34108 10156 35332 10212
rect 35388 10156 35972 10212
rect 36028 10156 37548 10212
rect 37604 10156 38188 10212
rect 38244 10156 39468 10212
rect 39524 10156 40108 10212
rect 40164 10156 41483 10212
rect 41539 10156 41587 10212
rect 41643 10156 41691 10212
rect 41747 10156 43108 10212
rect 43164 10156 43748 10212
rect 43804 10156 45028 10212
rect 45084 10156 45668 10212
rect 45724 10156 47244 10212
rect 47300 10156 47884 10212
rect 47940 10156 49164 10212
rect 49220 10156 49804 10212
rect 49860 10156 51138 10212
rect 51194 10156 51242 10212
rect 51298 10156 51346 10212
rect 51402 10156 52804 10212
rect 52860 10156 53444 10212
rect 53500 10156 54724 10212
rect 54780 10156 55364 10212
rect 55420 10156 56940 10212
rect 56996 10156 57580 10212
rect 57636 10156 58860 10212
rect 58916 10156 59500 10212
rect 59556 10156 60919 10212
rect 60975 10156 61023 10212
rect 61079 10156 61127 10212
rect 61183 10156 62500 10212
rect 62556 10156 63140 10212
rect 63196 10156 64420 10212
rect 64476 10156 65060 10212
rect 65116 10156 65126 10212
rect 31746 10108 65126 10156
rect 18985 10068 25493 10078
rect 18985 10012 21458 10068
rect 21514 10012 21562 10068
rect 21618 10012 21666 10068
rect 21722 10012 22756 10068
rect 22812 10012 22860 10068
rect 22916 10012 22964 10068
rect 23020 10012 25493 10068
rect 6003 9964 6183 9974
rect 7055 9964 7131 9974
rect 7695 9964 7771 9974
rect 6003 9908 6013 9964
rect 6069 9908 6117 9964
rect 6173 9908 7065 9964
rect 7121 9908 7705 9964
rect 7761 9908 7771 9964
rect 6003 9860 7771 9908
rect 2881 9812 3061 9822
rect 3950 9812 4026 9822
rect 2881 9756 2891 9812
rect 2947 9756 2995 9812
rect 3051 9756 3960 9812
rect 4016 9756 4026 9812
rect 6003 9804 6013 9860
rect 6069 9804 6117 9860
rect 6173 9804 7065 9860
rect 7121 9804 7705 9860
rect 7761 9804 7771 9860
rect 6003 9794 6183 9804
rect 7055 9794 7131 9804
rect 7695 9794 7771 9804
rect 18985 9964 25493 10012
rect 18985 9908 18995 9964
rect 19051 9908 19635 9964
rect 19691 9908 20275 9964
rect 20331 9908 21458 9964
rect 21514 9908 21562 9964
rect 21618 9908 21666 9964
rect 21722 9908 22756 9964
rect 22812 9908 22860 9964
rect 22916 9908 22964 9964
rect 23020 9908 24147 9964
rect 24203 9908 24787 9964
rect 24843 9908 25427 9964
rect 25483 9908 25493 9964
rect 18985 9860 25493 9908
rect 18985 9804 18995 9860
rect 19051 9804 19635 9860
rect 19691 9804 20275 9860
rect 20331 9804 21458 9860
rect 21514 9804 21562 9860
rect 21618 9804 21666 9860
rect 21722 9804 22756 9860
rect 22812 9804 22860 9860
rect 22916 9804 22964 9860
rect 23020 9804 24147 9860
rect 24203 9804 24787 9860
rect 24843 9804 25427 9860
rect 25483 9804 25493 9860
rect 18985 9794 25493 9804
rect 28106 10068 30853 10078
rect 28106 10012 30579 10068
rect 30635 10012 30683 10068
rect 30739 10012 30787 10068
rect 30843 10012 30853 10068
rect 31746 10052 31756 10108
rect 31812 10052 31860 10108
rect 31916 10052 31964 10108
rect 32020 10052 33412 10108
rect 33468 10052 34052 10108
rect 34108 10052 35332 10108
rect 35388 10052 35972 10108
rect 36028 10052 37548 10108
rect 37604 10052 38188 10108
rect 38244 10052 39468 10108
rect 39524 10052 40108 10108
rect 40164 10052 41483 10108
rect 41539 10052 41587 10108
rect 41643 10052 41691 10108
rect 41747 10052 43108 10108
rect 43164 10052 43748 10108
rect 43804 10052 45028 10108
rect 45084 10052 45668 10108
rect 45724 10052 47244 10108
rect 47300 10052 47884 10108
rect 47940 10052 49164 10108
rect 49220 10052 49804 10108
rect 49860 10052 51138 10108
rect 51194 10052 51242 10108
rect 51298 10052 51346 10108
rect 51402 10052 52804 10108
rect 52860 10052 53444 10108
rect 53500 10052 54724 10108
rect 54780 10052 55364 10108
rect 55420 10052 56940 10108
rect 56996 10052 57580 10108
rect 57636 10052 58860 10108
rect 58916 10052 59500 10108
rect 59556 10052 60919 10108
rect 60975 10052 61023 10108
rect 61079 10052 61127 10108
rect 61183 10052 62500 10108
rect 62556 10052 63140 10108
rect 63196 10052 64420 10108
rect 64476 10052 65060 10108
rect 65116 10052 65126 10108
rect 31746 10042 65126 10052
rect 28106 9964 30853 10012
rect 28106 9908 28116 9964
rect 28172 9908 28756 9964
rect 28812 9908 29396 9964
rect 29452 9908 30579 9964
rect 30635 9908 30683 9964
rect 30739 9908 30787 9964
rect 30843 9908 30853 9964
rect 28106 9860 30853 9908
rect 28106 9804 28116 9860
rect 28172 9804 28756 9860
rect 28812 9804 29396 9860
rect 29452 9804 30579 9860
rect 30635 9804 30683 9860
rect 30739 9804 30787 9860
rect 30843 9804 30853 9860
rect 28106 9794 30853 9804
rect -8154 9711 -7942 9721
rect -8154 9655 -8141 9711
rect -8085 9655 -8031 9711
rect -7975 9655 -7942 9711
rect -8154 9606 -7942 9655
rect 2881 9708 4026 9756
rect 2881 9652 2891 9708
rect 2947 9652 2995 9708
rect 3051 9652 3960 9708
rect 4016 9652 4026 9708
rect 2881 9642 3061 9652
rect 3950 9640 4026 9652
rect 10602 9763 10678 9773
rect 11371 9763 11551 9773
rect 10602 9707 10612 9763
rect 10668 9707 11381 9763
rect 11437 9707 11485 9763
rect 11541 9707 11551 9763
rect 10602 9659 11551 9707
rect -8154 9550 -8141 9606
rect -8085 9550 -8031 9606
rect -7975 9550 -7942 9606
rect 10602 9603 10612 9659
rect 10668 9603 11381 9659
rect 11437 9603 11485 9659
rect 11541 9603 11551 9659
rect 32126 9650 64807 9660
rect 10602 9593 10678 9603
rect 11371 9593 11551 9603
rect 17841 9633 19141 9643
rect 17841 9577 17851 9633
rect 17907 9577 19075 9633
rect 19131 9577 19141 9633
rect -8154 9501 -7942 9550
rect -8154 9445 -8141 9501
rect -8085 9445 -8031 9501
rect -7975 9445 -7942 9501
rect 5731 9563 5911 9573
rect 6735 9563 6811 9573
rect 7375 9563 7451 9573
rect 8015 9563 8091 9573
rect 9418 9563 9494 9573
rect 10314 9563 10390 9573
rect 17841 9567 19141 9577
rect 25337 9633 28262 9643
rect 25337 9577 25347 9633
rect 25403 9577 26571 9633
rect 26627 9577 26972 9633
rect 27028 9577 28196 9633
rect 28252 9577 28262 9633
rect 25337 9567 28262 9577
rect 32126 9594 32136 9650
rect 32192 9594 32240 9650
rect 32296 9594 32344 9650
rect 32400 9594 41122 9650
rect 41178 9594 41226 9650
rect 41282 9594 41330 9650
rect 41386 9594 41842 9650
rect 41898 9594 41946 9650
rect 42002 9594 42050 9650
rect 42106 9594 50798 9650
rect 50854 9594 50902 9650
rect 50958 9594 51006 9650
rect 51062 9594 51530 9650
rect 51586 9594 51634 9650
rect 51690 9594 51738 9650
rect 51794 9594 60514 9650
rect 60570 9594 60618 9650
rect 60674 9594 60722 9650
rect 60778 9594 61278 9650
rect 61334 9594 61382 9650
rect 61438 9594 61486 9650
rect 61542 9594 64807 9650
rect 5731 9507 5741 9563
rect 5797 9507 5845 9563
rect 5901 9507 6745 9563
rect 6801 9507 7385 9563
rect 7441 9507 8025 9563
rect 8081 9507 9428 9563
rect 9484 9507 10324 9563
rect 10380 9507 10390 9563
rect 32126 9546 64807 9594
rect -8154 9430 -7942 9445
rect 2624 9459 2700 9469
rect 4030 9459 4106 9469
rect 2624 9403 2634 9459
rect 2690 9403 4040 9459
rect 4096 9403 4106 9459
rect 2624 9355 4106 9403
rect 2624 9299 2634 9355
rect 2690 9299 4040 9355
rect 4096 9299 4106 9355
rect 2624 9289 2700 9299
rect 4030 9289 4106 9299
rect 4190 9459 4266 9469
rect 4831 9459 4907 9469
rect 5731 9459 10390 9507
rect 4190 9403 4200 9459
rect 4256 9403 4841 9459
rect 4897 9403 5741 9459
rect 5797 9403 5845 9459
rect 5901 9403 6745 9459
rect 6801 9403 7385 9459
rect 7441 9403 8025 9459
rect 8081 9403 9428 9459
rect 9484 9403 10324 9459
rect 10380 9403 10390 9459
rect 4190 9355 5911 9403
rect 6735 9393 6811 9403
rect 7375 9393 7451 9403
rect 8015 9393 8091 9403
rect 9418 9393 9494 9403
rect 10314 9393 10390 9403
rect 19305 9526 25173 9536
rect 19305 9470 21458 9526
rect 21514 9470 21562 9526
rect 21618 9470 21666 9526
rect 21722 9470 22756 9526
rect 22812 9470 22860 9526
rect 22916 9470 22964 9526
rect 23020 9470 25173 9526
rect 19305 9422 25173 9470
rect 4190 9299 4200 9355
rect 4256 9299 4841 9355
rect 4897 9299 5741 9355
rect 5797 9299 5845 9355
rect 5901 9299 5911 9355
rect 4190 9289 4266 9299
rect 4831 9289 4907 9299
rect 5731 9289 5911 9299
rect 19305 9366 19315 9422
rect 19371 9366 19955 9422
rect 20011 9366 21458 9422
rect 21514 9366 21562 9422
rect 21618 9366 21666 9422
rect 21722 9366 22756 9422
rect 22812 9366 22860 9422
rect 22916 9366 22964 9422
rect 23020 9366 24467 9422
rect 24523 9366 25107 9422
rect 25163 9366 25173 9422
rect 19305 9318 25173 9366
rect 11371 9275 11551 9285
rect 12352 9275 12428 9285
rect 13248 9275 13324 9285
rect 14144 9275 14220 9285
rect 11371 9219 11381 9275
rect 11437 9219 11485 9275
rect 11541 9219 12362 9275
rect 12418 9219 13258 9275
rect 13314 9219 14154 9275
rect 14210 9219 14220 9275
rect 19305 9262 19315 9318
rect 19371 9262 19955 9318
rect 20011 9262 21458 9318
rect 21514 9262 21562 9318
rect 21618 9262 21666 9318
rect 21722 9262 22756 9318
rect 22812 9262 22860 9318
rect 22916 9262 22964 9318
rect 23020 9262 24467 9318
rect 24523 9262 25107 9318
rect 25163 9262 25173 9318
rect 19305 9252 25173 9262
rect 28426 9526 30853 9536
rect 28426 9470 30579 9526
rect 30635 9470 30683 9526
rect 30739 9470 30787 9526
rect 30843 9470 30853 9526
rect 28426 9422 30853 9470
rect 28426 9366 28436 9422
rect 28492 9366 29076 9422
rect 29132 9366 30579 9422
rect 30635 9366 30683 9422
rect 30739 9366 30787 9422
rect 30843 9366 30853 9422
rect 32126 9490 32136 9546
rect 32192 9490 32240 9546
rect 32296 9490 32344 9546
rect 32400 9490 33733 9546
rect 33789 9490 34373 9546
rect 34429 9490 35013 9546
rect 35069 9490 35653 9546
rect 35709 9490 37867 9546
rect 37923 9490 38507 9546
rect 38563 9490 39147 9546
rect 39203 9490 39787 9546
rect 39843 9490 41122 9546
rect 41178 9490 41226 9546
rect 41282 9490 41330 9546
rect 41386 9490 41842 9546
rect 41898 9490 41946 9546
rect 42002 9490 42050 9546
rect 42106 9490 43429 9546
rect 43485 9490 44069 9546
rect 44125 9490 44709 9546
rect 44765 9490 45349 9546
rect 45405 9490 47563 9546
rect 47619 9490 48203 9546
rect 48259 9490 48843 9546
rect 48899 9490 49483 9546
rect 49539 9490 50798 9546
rect 50854 9490 50902 9546
rect 50958 9490 51006 9546
rect 51062 9490 51530 9546
rect 51586 9490 51634 9546
rect 51690 9490 51738 9546
rect 51794 9490 53125 9546
rect 53181 9490 53765 9546
rect 53821 9490 54405 9546
rect 54461 9490 55045 9546
rect 55101 9490 57259 9546
rect 57315 9490 57899 9546
rect 57955 9490 58539 9546
rect 58595 9490 59179 9546
rect 59235 9490 60514 9546
rect 60570 9490 60618 9546
rect 60674 9490 60722 9546
rect 60778 9490 61278 9546
rect 61334 9490 61382 9546
rect 61438 9490 61486 9546
rect 61542 9490 62821 9546
rect 62877 9490 63461 9546
rect 63517 9490 64101 9546
rect 64157 9490 64741 9546
rect 64797 9490 64807 9546
rect 32126 9442 64807 9490
rect 32126 9386 32136 9442
rect 32192 9386 32240 9442
rect 32296 9386 32344 9442
rect 32400 9386 33733 9442
rect 33789 9386 34373 9442
rect 34429 9386 35013 9442
rect 35069 9386 35653 9442
rect 35709 9386 37867 9442
rect 37923 9386 38507 9442
rect 38563 9386 39147 9442
rect 39203 9386 39787 9442
rect 39843 9386 41122 9442
rect 41178 9386 41226 9442
rect 41282 9386 41330 9442
rect 41386 9386 41842 9442
rect 41898 9386 41946 9442
rect 42002 9386 42050 9442
rect 42106 9386 43429 9442
rect 43485 9386 44069 9442
rect 44125 9386 44709 9442
rect 44765 9386 45349 9442
rect 45405 9386 47563 9442
rect 47619 9386 48203 9442
rect 48259 9386 48843 9442
rect 48899 9386 49483 9442
rect 49539 9386 50798 9442
rect 50854 9386 50902 9442
rect 50958 9386 51006 9442
rect 51062 9386 51530 9442
rect 51586 9386 51634 9442
rect 51690 9386 51738 9442
rect 51794 9386 53125 9442
rect 53181 9386 53765 9442
rect 53821 9386 54405 9442
rect 54461 9386 55045 9442
rect 55101 9386 57259 9442
rect 57315 9386 57899 9442
rect 57955 9386 58539 9442
rect 58595 9386 59179 9442
rect 59235 9386 60514 9442
rect 60570 9386 60618 9442
rect 60674 9386 60722 9442
rect 60778 9386 61278 9442
rect 61334 9386 61382 9442
rect 61438 9386 61486 9442
rect 61542 9386 62821 9442
rect 62877 9386 63461 9442
rect 63517 9386 64101 9442
rect 64157 9386 64741 9442
rect 64797 9386 64807 9442
rect 32126 9376 64807 9386
rect 28426 9318 30853 9366
rect 28426 9262 28436 9318
rect 28492 9262 29076 9318
rect 29132 9262 30579 9318
rect 30635 9262 30683 9318
rect 30739 9262 30787 9318
rect 30843 9262 30853 9318
rect 28426 9252 30853 9262
rect 31746 9256 65126 9266
rect 11371 9171 14220 9219
rect 11371 9115 11381 9171
rect 11437 9115 11485 9171
rect 11541 9115 12362 9171
rect 12418 9115 13258 9171
rect 13314 9115 14154 9171
rect 14210 9115 14220 9171
rect 31746 9200 31756 9256
rect 31812 9200 31860 9256
rect 31916 9200 31964 9256
rect 32020 9200 41483 9256
rect 41539 9200 41587 9256
rect 41643 9200 41691 9256
rect 41747 9200 51138 9256
rect 51194 9200 51242 9256
rect 51298 9200 51346 9256
rect 51402 9200 60919 9256
rect 60975 9200 61023 9256
rect 61079 9200 61127 9256
rect 61183 9200 65126 9256
rect 31746 9152 65126 9200
rect 31746 9142 31756 9152
rect 11371 9105 11551 9115
rect 12352 9105 12428 9115
rect 13248 9105 13324 9115
rect 14144 9105 14220 9115
rect 18985 9132 31756 9142
rect 18985 9076 22107 9132
rect 22163 9076 22211 9132
rect 22267 9076 22315 9132
rect 22371 9076 31228 9132
rect 31284 9076 31332 9132
rect 31388 9076 31436 9132
rect 31492 9096 31756 9132
rect 31812 9096 31860 9152
rect 31916 9096 31964 9152
rect 32020 9096 33412 9152
rect 33468 9096 34052 9152
rect 34108 9096 35332 9152
rect 35388 9096 35972 9152
rect 36028 9096 37548 9152
rect 37604 9096 38188 9152
rect 38244 9096 39468 9152
rect 39524 9096 40108 9152
rect 40164 9096 41483 9152
rect 41539 9096 41587 9152
rect 41643 9096 41691 9152
rect 41747 9096 43108 9152
rect 43164 9096 43748 9152
rect 43804 9096 45028 9152
rect 45084 9096 45668 9152
rect 45724 9096 47244 9152
rect 47300 9096 47884 9152
rect 47940 9096 49164 9152
rect 49220 9096 49804 9152
rect 49860 9096 51138 9152
rect 51194 9096 51242 9152
rect 51298 9096 51346 9152
rect 51402 9096 52804 9152
rect 52860 9096 53444 9152
rect 53500 9096 54724 9152
rect 54780 9096 55364 9152
rect 55420 9096 56940 9152
rect 56996 9096 57580 9152
rect 57636 9096 58860 9152
rect 58916 9096 59500 9152
rect 59556 9096 60919 9152
rect 60975 9096 61023 9152
rect 61079 9096 61127 9152
rect 61183 9096 62500 9152
rect 62556 9096 63140 9152
rect 63196 9096 64420 9152
rect 64476 9096 65060 9152
rect 65116 9096 65126 9152
rect 31492 9076 65126 9096
rect 18985 9048 65126 9076
rect 18985 9028 31756 9048
rect 3870 8963 3946 8973
rect 4510 8963 4586 8973
rect 5150 8963 5226 8973
rect 6003 8963 6183 8973
rect 6735 8963 6811 8973
rect 7375 8963 7451 8973
rect 8015 8963 8091 8973
rect 8970 8963 9046 8973
rect 9866 8963 9942 8973
rect 10762 8963 10838 8973
rect 3870 8907 3880 8963
rect 3936 8907 4520 8963
rect 4576 8907 5160 8963
rect 5216 8907 6013 8963
rect 6069 8907 6117 8963
rect 6173 8907 6745 8963
rect 6801 8907 7385 8963
rect 7441 8907 8025 8963
rect 8081 8907 8980 8963
rect 9036 8907 9876 8963
rect 9932 8907 10772 8963
rect 10828 8907 10838 8963
rect 3870 8859 10838 8907
rect 18985 8972 18995 9028
rect 19051 8972 19635 9028
rect 19691 8972 20275 9028
rect 20331 8972 22107 9028
rect 22163 8972 22211 9028
rect 22267 8972 22315 9028
rect 22371 8972 24147 9028
rect 24203 8972 24787 9028
rect 24843 8972 25427 9028
rect 25483 8972 28116 9028
rect 28172 8972 28756 9028
rect 28812 8972 29396 9028
rect 29452 8972 31228 9028
rect 31284 8972 31332 9028
rect 31388 8972 31436 9028
rect 31492 8992 31756 9028
rect 31812 8992 31860 9048
rect 31916 8992 31964 9048
rect 32020 8992 33412 9048
rect 33468 8992 34052 9048
rect 34108 8992 35332 9048
rect 35388 8992 35972 9048
rect 36028 8992 37548 9048
rect 37604 8992 38188 9048
rect 38244 8992 39468 9048
rect 39524 8992 40108 9048
rect 40164 8992 41483 9048
rect 41539 8992 41587 9048
rect 41643 8992 41691 9048
rect 41747 8992 43108 9048
rect 43164 8992 43748 9048
rect 43804 8992 45028 9048
rect 45084 8992 45668 9048
rect 45724 8992 47244 9048
rect 47300 8992 47884 9048
rect 47940 8992 49164 9048
rect 49220 8992 49804 9048
rect 49860 8992 51138 9048
rect 51194 8992 51242 9048
rect 51298 8992 51346 9048
rect 51402 8992 52804 9048
rect 52860 8992 53444 9048
rect 53500 8992 54724 9048
rect 54780 8992 55364 9048
rect 55420 8992 56940 9048
rect 56996 8992 57580 9048
rect 57636 8992 58860 9048
rect 58916 8992 59500 9048
rect 59556 8992 60919 9048
rect 60975 8992 61023 9048
rect 61079 8992 61127 9048
rect 61183 8992 62500 9048
rect 62556 8992 63140 9048
rect 63196 8992 64420 9048
rect 64476 8992 65060 9048
rect 65116 8992 65126 9048
rect 31492 8982 65126 8992
rect 31492 8972 32030 8982
rect 18985 8924 32030 8972
rect 3870 8803 3880 8859
rect 3936 8803 4520 8859
rect 4576 8803 5160 8859
rect 5216 8803 6013 8859
rect 6069 8803 6117 8859
rect 6173 8803 6745 8859
rect 6801 8803 7385 8859
rect 7441 8803 8025 8859
rect 8081 8803 8980 8859
rect 9036 8803 9876 8859
rect 9932 8803 10772 8859
rect 10828 8803 10838 8859
rect -8513 8782 -8303 8794
rect 3870 8793 3946 8803
rect 4510 8793 4586 8803
rect 5150 8793 5226 8803
rect 6003 8793 6183 8803
rect 6735 8793 6811 8803
rect 7375 8793 7451 8803
rect 8015 8793 8091 8803
rect 8970 8793 9046 8803
rect 9866 8793 9942 8803
rect 10762 8793 10838 8803
rect 13856 8875 13932 8885
rect 15466 8875 15542 8885
rect 16106 8875 16182 8885
rect 17365 8875 17545 8885
rect 13856 8819 13866 8875
rect 13922 8819 15476 8875
rect 15532 8819 16116 8875
rect 16172 8819 17375 8875
rect 17431 8819 17479 8875
rect 17535 8819 17545 8875
rect 18985 8868 18995 8924
rect 19051 8868 19635 8924
rect 19691 8868 20275 8924
rect 20331 8868 22107 8924
rect 22163 8868 22211 8924
rect 22267 8868 22315 8924
rect 22371 8868 24147 8924
rect 24203 8868 24787 8924
rect 24843 8868 25427 8924
rect 25483 8868 28116 8924
rect 28172 8868 28756 8924
rect 28812 8868 29396 8924
rect 29452 8868 31228 8924
rect 31284 8868 31332 8924
rect 31388 8868 31436 8924
rect 31492 8868 32030 8924
rect 18985 8858 32030 8868
rect -8513 8726 -8491 8782
rect -8435 8726 -8381 8782
rect -8325 8726 -8303 8782
rect -8513 8672 -8303 8726
rect 13856 8771 17545 8819
rect 13856 8715 13866 8771
rect 13922 8715 15476 8771
rect 15532 8715 16116 8771
rect 16172 8715 17375 8771
rect 17431 8715 17479 8771
rect 17535 8715 17545 8771
rect 10474 8705 10550 8715
rect 11639 8705 11819 8715
rect 13856 8705 13932 8715
rect 15466 8705 15542 8715
rect 16106 8705 16182 8715
rect 17365 8705 17545 8715
rect -8513 8616 -8491 8672
rect -8435 8616 -8381 8672
rect -8325 8616 -8303 8672
rect -8513 8562 -8303 8616
rect -8513 8506 -8491 8562
rect -8435 8506 -8381 8562
rect -8325 8506 -8303 8562
rect 3161 8682 3341 8692
rect 3950 8682 4026 8692
rect 3161 8626 3171 8682
rect 3227 8626 3275 8682
rect 3331 8626 3960 8682
rect 4016 8626 4026 8682
rect 3161 8578 4026 8626
rect 3161 8522 3171 8578
rect 3227 8522 3275 8578
rect 3331 8522 3960 8578
rect 4016 8522 4026 8578
rect 3161 8512 3341 8522
rect 3950 8512 4026 8522
rect 5731 8690 5911 8700
rect 7055 8690 7131 8700
rect 7695 8690 7771 8700
rect 5731 8634 5741 8690
rect 5797 8634 5845 8690
rect 5901 8634 7065 8690
rect 7121 8634 7705 8690
rect 7761 8634 7771 8690
rect 5731 8586 7771 8634
rect 5731 8530 5741 8586
rect 5797 8530 5845 8586
rect 5901 8530 7065 8586
rect 7121 8530 7705 8586
rect 7761 8530 7771 8586
rect 10474 8649 10484 8705
rect 10540 8649 11649 8705
rect 11705 8649 11753 8705
rect 11809 8649 11819 8705
rect 10474 8601 11819 8649
rect 17641 8697 19141 8707
rect 17641 8641 17651 8697
rect 17707 8641 19075 8697
rect 19131 8641 19141 8697
rect 17641 8631 19141 8641
rect 25337 8697 28262 8707
rect 25337 8641 25347 8697
rect 25403 8641 26771 8697
rect 26828 8641 28196 8697
rect 28252 8641 28262 8697
rect 25337 8631 28262 8641
rect 10474 8545 10484 8601
rect 10540 8545 11649 8601
rect 11705 8545 11753 8601
rect 11809 8545 11819 8601
rect 19305 8590 25173 8600
rect 10474 8535 10550 8545
rect 11639 8535 11819 8545
rect 12018 8565 12198 8575
rect 12388 8565 12464 8575
rect 5731 8520 5911 8530
rect 7055 8520 7131 8530
rect 7695 8520 7771 8530
rect -8513 8452 -8303 8506
rect 12018 8509 12028 8565
rect 12084 8509 12132 8565
rect 12188 8509 12398 8565
rect 12454 8509 12464 8565
rect -8513 8396 -8491 8452
rect -8435 8396 -8381 8452
rect -8325 8396 -8303 8452
rect -8513 8368 -8303 8396
rect 7989 8466 8065 8476
rect 8275 8466 8455 8476
rect 7989 8410 7999 8466
rect 8055 8410 8285 8466
rect 8341 8410 8389 8466
rect 8445 8410 8455 8466
rect 7989 8362 8455 8410
rect 4190 8329 4266 8339
rect 4831 8329 4907 8339
rect 6003 8329 6183 8339
rect 4190 8273 4200 8329
rect 4256 8273 4841 8329
rect 4897 8273 6013 8329
rect 6069 8273 6117 8329
rect 6173 8273 6183 8329
rect 7989 8306 7999 8362
rect 8055 8306 8285 8362
rect 8341 8306 8389 8362
rect 8445 8306 8455 8362
rect 7989 8296 8065 8306
rect 8275 8296 8455 8306
rect 10722 8455 10798 8465
rect 10918 8455 11098 8465
rect 10722 8399 10732 8455
rect 10788 8399 10928 8455
rect 10984 8399 11032 8455
rect 11088 8399 11098 8455
rect 10722 8351 11098 8399
rect 12018 8461 12464 8509
rect 12018 8405 12028 8461
rect 12084 8405 12132 8461
rect 12188 8405 12398 8461
rect 12454 8405 12464 8461
rect 12018 8395 12198 8405
rect 12388 8395 12464 8405
rect 14686 8570 14866 8580
rect 15174 8570 15250 8580
rect 14686 8514 14696 8570
rect 14752 8514 14800 8570
rect 14856 8514 15184 8570
rect 15240 8514 15250 8570
rect 14686 8466 15250 8514
rect 14686 8410 14696 8466
rect 14752 8410 14800 8466
rect 14856 8410 15184 8466
rect 15240 8410 15250 8466
rect 14686 8400 14866 8410
rect 15174 8400 15250 8410
rect 19305 8534 22107 8590
rect 22163 8534 22211 8590
rect 22267 8534 22315 8590
rect 22371 8534 25173 8590
rect 19305 8486 25173 8534
rect 19305 8430 19315 8486
rect 19371 8430 19955 8486
rect 20011 8430 22107 8486
rect 22163 8430 22211 8486
rect 22267 8430 22315 8486
rect 22371 8430 24467 8486
rect 24523 8430 25107 8486
rect 25163 8430 25173 8486
rect 10722 8295 10732 8351
rect 10788 8295 10928 8351
rect 10984 8295 11032 8351
rect 11088 8295 11098 8351
rect 19305 8382 25173 8430
rect 19305 8326 19315 8382
rect 19371 8326 19955 8382
rect 20011 8326 22107 8382
rect 22163 8326 22211 8382
rect 22267 8326 22315 8382
rect 22371 8326 24467 8382
rect 24523 8326 25107 8382
rect 25163 8326 25173 8382
rect 19305 8316 25173 8326
rect 28426 8590 64807 8600
rect 28426 8534 31228 8590
rect 31284 8534 31332 8590
rect 31388 8534 31436 8590
rect 31492 8534 31756 8590
rect 31812 8534 31860 8590
rect 31916 8534 31964 8590
rect 32020 8534 41483 8590
rect 41539 8534 41587 8590
rect 41643 8534 41691 8590
rect 41747 8534 51138 8590
rect 51194 8534 51242 8590
rect 51298 8534 51346 8590
rect 51402 8534 60919 8590
rect 60975 8534 61023 8590
rect 61079 8534 61127 8590
rect 61183 8534 64807 8590
rect 28426 8486 64807 8534
rect 28426 8430 28436 8486
rect 28492 8430 29076 8486
rect 29132 8430 31228 8486
rect 31284 8430 31332 8486
rect 31388 8430 31436 8486
rect 31492 8430 31756 8486
rect 31812 8430 31860 8486
rect 31916 8430 31964 8486
rect 32020 8430 33733 8486
rect 33789 8430 34373 8486
rect 34429 8430 35013 8486
rect 35069 8430 35653 8486
rect 35709 8430 37867 8486
rect 37923 8430 38507 8486
rect 38563 8430 39147 8486
rect 39203 8430 39787 8486
rect 39843 8430 41483 8486
rect 41539 8430 41587 8486
rect 41643 8430 41691 8486
rect 41747 8430 43429 8486
rect 43485 8430 44069 8486
rect 44125 8430 44709 8486
rect 44765 8430 45349 8486
rect 45405 8430 47563 8486
rect 47619 8430 48203 8486
rect 48259 8430 48843 8486
rect 48899 8430 49483 8486
rect 49539 8430 51138 8486
rect 51194 8430 51242 8486
rect 51298 8430 51346 8486
rect 51402 8430 53125 8486
rect 53181 8430 53765 8486
rect 53821 8430 54405 8486
rect 54461 8430 55045 8486
rect 55101 8430 57259 8486
rect 57315 8430 57899 8486
rect 57955 8430 58539 8486
rect 58595 8430 59179 8486
rect 59235 8430 60919 8486
rect 60975 8430 61023 8486
rect 61079 8430 61127 8486
rect 61183 8430 62821 8486
rect 62877 8430 63461 8486
rect 63517 8430 64101 8486
rect 64157 8430 64741 8486
rect 64797 8430 64807 8486
rect 28426 8382 64807 8430
rect 28426 8326 28436 8382
rect 28492 8326 29076 8382
rect 29132 8326 31228 8382
rect 31284 8326 31332 8382
rect 31388 8326 31436 8382
rect 31492 8326 31756 8382
rect 31812 8326 31860 8382
rect 31916 8326 31964 8382
rect 32020 8326 33733 8382
rect 33789 8326 34373 8382
rect 34429 8326 35013 8382
rect 35069 8326 35653 8382
rect 35709 8326 37867 8382
rect 37923 8326 38507 8382
rect 38563 8326 39147 8382
rect 39203 8326 39787 8382
rect 39843 8326 41483 8382
rect 41539 8326 41587 8382
rect 41643 8326 41691 8382
rect 41747 8326 43429 8382
rect 43485 8326 44069 8382
rect 44125 8326 44709 8382
rect 44765 8326 45349 8382
rect 45405 8326 47563 8382
rect 47619 8326 48203 8382
rect 48259 8326 48843 8382
rect 48899 8326 49483 8382
rect 49539 8326 51138 8382
rect 51194 8326 51242 8382
rect 51298 8326 51346 8382
rect 51402 8326 53125 8382
rect 53181 8326 53765 8382
rect 53821 8326 54405 8382
rect 54461 8326 55045 8382
rect 55101 8326 57259 8382
rect 57315 8326 57899 8382
rect 57955 8326 58539 8382
rect 58595 8326 59179 8382
rect 59235 8326 60919 8382
rect 60975 8326 61023 8382
rect 61079 8326 61127 8382
rect 61183 8326 62821 8382
rect 62877 8326 63461 8382
rect 63517 8326 64101 8382
rect 64157 8326 64741 8382
rect 64797 8326 64807 8382
rect 28426 8316 64807 8326
rect 10722 8285 10798 8295
rect 10918 8285 11098 8295
rect 4190 8225 6183 8273
rect 7055 8225 7131 8235
rect 7695 8225 7771 8235
rect 9418 8225 9494 8235
rect 10314 8225 10390 8235
rect 4190 8169 4200 8225
rect 4256 8169 4841 8225
rect 4897 8169 6013 8225
rect 6069 8169 6117 8225
rect 6173 8169 7065 8225
rect 7121 8169 7705 8225
rect 7761 8169 9428 8225
rect 9484 8169 10324 8225
rect 10380 8169 10390 8225
rect 4190 8159 4266 8169
rect 4831 8159 4907 8169
rect 2624 8129 2700 8139
rect 4030 8129 4106 8139
rect 2624 8073 2634 8129
rect 2690 8073 4040 8129
rect 4096 8073 4106 8129
rect 2624 8025 4106 8073
rect 6003 8121 10390 8169
rect 6003 8065 6013 8121
rect 6069 8065 6117 8121
rect 6173 8065 7065 8121
rect 7121 8065 7705 8121
rect 7761 8065 9428 8121
rect 9484 8065 10324 8121
rect 10380 8065 10390 8121
rect 6003 8055 6183 8065
rect 7055 8055 7131 8065
rect 7695 8055 7771 8065
rect 9418 8055 9494 8065
rect 10314 8055 10390 8065
rect 10474 8225 10550 8235
rect 11371 8225 11551 8235
rect 12800 8225 12876 8235
rect 13696 8225 13772 8235
rect 10474 8169 10484 8225
rect 10540 8169 11381 8225
rect 11437 8169 11485 8225
rect 11541 8169 12810 8225
rect 12866 8169 13706 8225
rect 13762 8169 13772 8225
rect 10474 8121 13772 8169
rect 10474 8065 10484 8121
rect 10540 8065 11381 8121
rect 11437 8065 11485 8121
rect 11541 8065 12810 8121
rect 12866 8065 13706 8121
rect 13762 8065 13772 8121
rect 10474 8055 10550 8065
rect 11371 8055 11551 8065
rect 12800 8055 12876 8065
rect 13696 8055 13772 8065
rect 13856 8225 13932 8235
rect 15466 8225 15542 8235
rect 16106 8225 16182 8235
rect 17103 8225 17283 8235
rect 13856 8169 13866 8225
rect 13922 8169 15476 8225
rect 15532 8169 16116 8225
rect 16172 8169 17113 8225
rect 17169 8169 17217 8225
rect 17273 8169 17283 8225
rect 13856 8121 17283 8169
rect 13856 8065 13866 8121
rect 13922 8065 15476 8121
rect 15532 8065 16116 8121
rect 16172 8065 17113 8121
rect 17169 8065 17217 8121
rect 17273 8065 17283 8121
rect 13856 8055 13932 8065
rect 15466 8055 15542 8065
rect 16106 8055 16182 8065
rect 17103 8055 17283 8065
rect 18985 8196 65126 8206
rect 18985 8140 21458 8196
rect 21514 8140 21562 8196
rect 21618 8140 21666 8196
rect 21722 8140 22756 8196
rect 22812 8140 22860 8196
rect 22916 8140 22964 8196
rect 23020 8140 30579 8196
rect 30635 8140 30683 8196
rect 30739 8140 30787 8196
rect 30843 8140 32136 8196
rect 32192 8140 32240 8196
rect 32296 8140 32344 8196
rect 32400 8140 41122 8196
rect 41178 8140 41226 8196
rect 41282 8140 41330 8196
rect 41386 8140 41842 8196
rect 41898 8140 41946 8196
rect 42002 8140 42050 8196
rect 42106 8140 50798 8196
rect 50854 8140 50902 8196
rect 50958 8140 51006 8196
rect 51062 8140 51530 8196
rect 51586 8140 51634 8196
rect 51690 8140 51738 8196
rect 51794 8140 60514 8196
rect 60570 8140 60618 8196
rect 60674 8140 60722 8196
rect 60778 8140 61278 8196
rect 61334 8140 61382 8196
rect 61438 8140 61486 8196
rect 61542 8140 65126 8196
rect 18985 8092 65126 8140
rect 2624 7969 2634 8025
rect 2690 7969 4040 8025
rect 4096 7969 4106 8025
rect 2624 7959 2700 7969
rect 4030 7959 4106 7969
rect 18985 8036 18995 8092
rect 19051 8036 19635 8092
rect 19691 8036 20275 8092
rect 20331 8036 21458 8092
rect 21514 8036 21562 8092
rect 21618 8036 21666 8092
rect 21722 8036 22756 8092
rect 22812 8036 22860 8092
rect 22916 8036 22964 8092
rect 23020 8036 24147 8092
rect 24203 8036 24787 8092
rect 24843 8036 25427 8092
rect 25483 8036 28116 8092
rect 28172 8036 28756 8092
rect 28812 8036 29396 8092
rect 29452 8036 30579 8092
rect 30635 8036 30683 8092
rect 30739 8036 30787 8092
rect 30843 8036 32136 8092
rect 32192 8036 32240 8092
rect 32296 8036 32344 8092
rect 32400 8036 33412 8092
rect 33468 8036 34052 8092
rect 34108 8036 35332 8092
rect 35388 8036 35972 8092
rect 36028 8036 37548 8092
rect 37604 8036 38188 8092
rect 38244 8036 39468 8092
rect 39524 8036 40108 8092
rect 40164 8036 41122 8092
rect 41178 8036 41226 8092
rect 41282 8036 41330 8092
rect 41386 8036 41842 8092
rect 41898 8036 41946 8092
rect 42002 8036 42050 8092
rect 42106 8036 43108 8092
rect 43164 8036 43748 8092
rect 43804 8036 45028 8092
rect 45084 8036 45668 8092
rect 45724 8036 47244 8092
rect 47300 8036 47884 8092
rect 47940 8036 49164 8092
rect 49220 8036 49804 8092
rect 49860 8036 50798 8092
rect 50854 8036 50902 8092
rect 50958 8036 51006 8092
rect 51062 8036 51530 8092
rect 51586 8036 51634 8092
rect 51690 8036 51738 8092
rect 51794 8036 52804 8092
rect 52860 8036 53444 8092
rect 53500 8036 54724 8092
rect 54780 8036 55364 8092
rect 55420 8036 56940 8092
rect 56996 8036 57580 8092
rect 57636 8036 58860 8092
rect 58916 8036 59500 8092
rect 59556 8036 60514 8092
rect 60570 8036 60618 8092
rect 60674 8036 60722 8092
rect 60778 8036 61278 8092
rect 61334 8036 61382 8092
rect 61438 8036 61486 8092
rect 61542 8036 62500 8092
rect 62556 8036 63140 8092
rect 63196 8036 64420 8092
rect 64476 8036 65060 8092
rect 65116 8036 65126 8092
rect 18985 7988 65126 8036
rect -10593 7920 -10178 7946
rect 18985 7932 18995 7988
rect 19051 7932 19635 7988
rect 19691 7932 20275 7988
rect 20331 7932 21458 7988
rect 21514 7932 21562 7988
rect 21618 7932 21666 7988
rect 21722 7932 22756 7988
rect 22812 7932 22860 7988
rect 22916 7932 22964 7988
rect 23020 7932 24147 7988
rect 24203 7932 24787 7988
rect 24843 7932 25427 7988
rect 25483 7932 28116 7988
rect 28172 7932 28756 7988
rect 28812 7932 29396 7988
rect 29452 7932 30579 7988
rect 30635 7932 30683 7988
rect 30739 7932 30787 7988
rect 30843 7932 32136 7988
rect 32192 7932 32240 7988
rect 32296 7932 32344 7988
rect 32400 7932 33412 7988
rect 33468 7932 34052 7988
rect 34108 7932 35332 7988
rect 35388 7932 35972 7988
rect 36028 7932 37548 7988
rect 37604 7932 38188 7988
rect 38244 7932 39468 7988
rect 39524 7932 40108 7988
rect 40164 7932 41122 7988
rect 41178 7932 41226 7988
rect 41282 7932 41330 7988
rect 41386 7932 41842 7988
rect 41898 7932 41946 7988
rect 42002 7932 42050 7988
rect 42106 7932 43108 7988
rect 43164 7932 43748 7988
rect 43804 7932 45028 7988
rect 45084 7932 45668 7988
rect 45724 7932 47244 7988
rect 47300 7932 47884 7988
rect 47940 7932 49164 7988
rect 49220 7932 49804 7988
rect 49860 7932 50798 7988
rect 50854 7932 50902 7988
rect 50958 7932 51006 7988
rect 51062 7932 51530 7988
rect 51586 7932 51634 7988
rect 51690 7932 51738 7988
rect 51794 7932 52804 7988
rect 52860 7932 53444 7988
rect 53500 7932 54724 7988
rect 54780 7932 55364 7988
rect 55420 7932 56940 7988
rect 56996 7932 57580 7988
rect 57636 7932 58860 7988
rect 58916 7932 59500 7988
rect 59556 7932 60514 7988
rect 60570 7932 60618 7988
rect 60674 7932 60722 7988
rect 60778 7932 61278 7988
rect 61334 7932 61382 7988
rect 61438 7932 61486 7988
rect 61542 7932 62500 7988
rect 62556 7932 63140 7988
rect 63196 7932 64420 7988
rect 64476 7932 65060 7988
rect 65116 7932 65126 7988
rect 18985 7922 65126 7932
rect -10593 7864 -10576 7920
rect -10520 7864 -10466 7920
rect -10410 7864 -10356 7920
rect -10300 7864 -10246 7920
rect -10190 7864 -10178 7920
rect -10593 7810 -10178 7864
rect -10593 7754 -10576 7810
rect -10520 7754 -10466 7810
rect -10410 7754 -10356 7810
rect -10300 7754 -10246 7810
rect -10190 7754 -10178 7810
rect -10593 7721 -10178 7754
rect 3870 7833 3946 7843
rect 4510 7833 4586 7843
rect 5150 7833 5226 7843
rect 5731 7833 5911 7843
rect 6735 7833 6811 7843
rect 7375 7833 7451 7843
rect 8015 7833 8091 7843
rect 8970 7833 9046 7843
rect 9866 7833 9942 7843
rect 10762 7833 10838 7843
rect 15146 7835 15222 7845
rect 15786 7835 15862 7845
rect 16426 7835 16502 7845
rect 17365 7835 17545 7845
rect 3870 7777 3880 7833
rect 3936 7777 4520 7833
rect 4576 7777 5160 7833
rect 5216 7777 5741 7833
rect 5797 7777 5845 7833
rect 5901 7777 6745 7833
rect 6801 7777 7385 7833
rect 7441 7777 8025 7833
rect 8081 7777 8980 7833
rect 9036 7777 9876 7833
rect 9932 7777 10772 7833
rect 10828 7777 10838 7833
rect 3870 7729 10838 7777
rect 3870 7673 3880 7729
rect 3936 7673 4520 7729
rect 4576 7673 5160 7729
rect 5216 7673 5741 7729
rect 5797 7673 5845 7729
rect 5901 7673 6745 7729
rect 6801 7673 7385 7729
rect 7441 7673 8025 7729
rect 8081 7673 8980 7729
rect 9036 7673 9876 7729
rect 9932 7673 10772 7729
rect 10828 7673 10838 7729
rect 3870 7663 3946 7673
rect 4510 7663 4586 7673
rect 5150 7663 5226 7673
rect 5731 7663 5911 7673
rect 6735 7663 6811 7673
rect 7375 7663 7451 7673
rect 8015 7663 8091 7673
rect 8970 7663 9046 7673
rect 9866 7663 9942 7673
rect 10762 7663 10838 7673
rect 11639 7825 11819 7835
rect 12352 7825 12428 7835
rect 13248 7825 13324 7835
rect 14144 7825 14220 7835
rect 11639 7769 11649 7825
rect 11705 7769 11753 7825
rect 11809 7769 12362 7825
rect 12418 7769 13258 7825
rect 13314 7769 14154 7825
rect 14210 7769 14220 7825
rect 11639 7721 14220 7769
rect 11639 7665 11649 7721
rect 11705 7665 11753 7721
rect 11809 7665 12362 7721
rect 12418 7665 13258 7721
rect 13314 7665 14154 7721
rect 14210 7665 14220 7721
rect 15146 7779 15156 7835
rect 15212 7779 15796 7835
rect 15852 7779 16436 7835
rect 16492 7779 17375 7835
rect 17431 7779 17479 7835
rect 17535 7779 17545 7835
rect 15146 7731 17545 7779
rect 15146 7675 15156 7731
rect 15212 7675 15796 7731
rect 15852 7675 16436 7731
rect 16492 7675 17375 7731
rect 17431 7675 17479 7731
rect 17535 7675 17545 7731
rect 17841 7761 19301 7771
rect 17841 7705 17851 7761
rect 17907 7705 19235 7761
rect 19291 7705 19301 7761
rect 17841 7695 19301 7705
rect 19865 7761 24613 7771
rect 19865 7705 19875 7761
rect 19931 7705 24547 7761
rect 24603 7705 24613 7761
rect 19865 7695 24613 7705
rect 25177 7761 28422 7771
rect 25177 7705 25187 7761
rect 25243 7705 26571 7761
rect 26627 7705 26972 7761
rect 27028 7705 28356 7761
rect 28412 7705 28422 7761
rect 25177 7695 28422 7705
rect 15146 7665 15222 7675
rect 15786 7665 15862 7675
rect 16426 7665 16502 7675
rect 17365 7665 17545 7675
rect 11639 7655 11819 7665
rect 12352 7655 12428 7665
rect 13248 7655 13324 7665
rect 14144 7655 14220 7665
rect 226 7585 406 7595
rect 1227 7585 1407 7595
rect 226 7529 236 7585
rect 292 7529 340 7585
rect 396 7529 1237 7585
rect 1293 7529 1341 7585
rect 1397 7529 1407 7585
rect 226 7481 1407 7529
rect 226 7425 236 7481
rect 292 7425 340 7481
rect 396 7425 1237 7481
rect 1293 7425 1341 7481
rect 1397 7425 1407 7481
rect 226 7415 406 7425
rect 1227 7415 1407 7425
rect 2881 7494 3061 7504
rect 4110 7494 4186 7504
rect 2881 7438 2891 7494
rect 2947 7438 2995 7494
rect 3051 7438 4120 7494
rect 4176 7438 4186 7494
rect 2881 7390 4186 7438
rect 2881 7334 2891 7390
rect 2947 7334 2995 7390
rect 3051 7334 4120 7390
rect 4176 7334 4186 7390
rect 2881 7324 3061 7334
rect 4110 7324 4186 7334
rect 17119 6438 30780 6448
rect 7382 6411 7562 6421
rect 8275 6411 8455 6421
rect 7382 6355 7392 6411
rect 7448 6355 7496 6411
rect 7552 6355 8285 6411
rect 8341 6355 8389 6411
rect 8445 6355 8455 6411
rect 7382 6307 8455 6355
rect 7382 6251 7392 6307
rect 7448 6251 7496 6307
rect 7552 6251 8285 6307
rect 8341 6251 8389 6307
rect 8445 6251 8455 6307
rect 7382 6241 7562 6251
rect 8275 6241 8455 6251
rect 17119 6382 17129 6438
rect 17185 6382 17233 6438
rect 17289 6382 17337 6438
rect 17393 6382 30298 6438
rect 30354 6382 30402 6438
rect 30458 6382 30506 6438
rect 30562 6382 30610 6438
rect 30666 6382 30714 6438
rect 30770 6382 30780 6438
rect 17119 6334 30780 6382
rect 17119 6278 17129 6334
rect 17185 6278 17233 6334
rect 17289 6278 17337 6334
rect 17393 6278 30298 6334
rect 30354 6278 30402 6334
rect 30458 6278 30506 6334
rect 30562 6278 30610 6334
rect 30666 6278 30714 6334
rect 30770 6278 30780 6334
rect 17119 6230 30780 6278
rect 17119 6174 17129 6230
rect 17185 6174 17233 6230
rect 17289 6174 17337 6230
rect 17393 6174 30298 6230
rect 30354 6174 30402 6230
rect 30458 6174 30506 6230
rect 30562 6174 30610 6230
rect 30666 6174 30714 6230
rect 30770 6174 30780 6230
rect 17119 6164 30780 6174
rect 17556 6096 30220 6106
rect 9189 6044 9265 6054
rect 10278 6044 10458 6054
rect -3303 5988 9199 6044
rect 9255 5988 10288 6044
rect 10344 5988 10392 6044
rect 10448 5988 10458 6044
rect -3303 5940 10458 5988
rect -3303 5884 9199 5940
rect 9255 5884 10288 5940
rect 10344 5884 10392 5940
rect 10448 5884 10458 5940
rect -8159 5532 -7863 5550
rect -8159 5476 -8146 5532
rect -8090 5476 -8041 5532
rect -7985 5476 -7936 5532
rect -7880 5476 -7863 5532
rect -8159 5422 -7863 5476
rect -8159 5366 -8146 5422
rect -8090 5366 -8041 5422
rect -7985 5366 -7936 5422
rect -7880 5366 -7863 5422
rect -8159 5338 -7863 5366
rect -3303 5277 -3143 5884
rect 9189 5874 9265 5884
rect 10278 5874 10458 5884
rect 17556 6040 17566 6096
rect 17622 6040 17670 6096
rect 17726 6040 17774 6096
rect 17830 6040 29738 6096
rect 29794 6040 29842 6096
rect 29898 6040 29946 6096
rect 30002 6040 30050 6096
rect 30106 6040 30154 6096
rect 30210 6040 30220 6096
rect 17556 5992 30220 6040
rect 17556 5936 17566 5992
rect 17622 5936 17670 5992
rect 17726 5936 17774 5992
rect 17830 5936 29738 5992
rect 29794 5936 29842 5992
rect 29898 5936 29946 5992
rect 30002 5936 30050 5992
rect 30106 5936 30154 5992
rect 30210 5936 30220 5992
rect 17556 5888 30220 5936
rect 17556 5832 17566 5888
rect 17622 5832 17670 5888
rect 17726 5832 17774 5888
rect 17830 5832 29738 5888
rect 29794 5832 29842 5888
rect 29898 5832 29946 5888
rect 30002 5832 30050 5888
rect 30106 5832 30154 5888
rect 30210 5832 30220 5888
rect 17556 5822 30220 5832
rect 7829 5711 7905 5721
rect 8149 5711 8225 5721
rect 8469 5711 8545 5721
rect 8789 5711 8865 5721
rect 7829 5655 7839 5711
rect 7895 5655 8159 5711
rect 8215 5655 8479 5711
rect 8535 5655 8799 5711
rect 8855 5655 8865 5711
rect 7829 5607 8865 5655
rect 7829 5551 7839 5607
rect 7895 5551 8159 5607
rect 8215 5551 8479 5607
rect 8535 5551 8799 5607
rect 8855 5551 8865 5607
rect 7829 5541 7905 5551
rect 8149 5541 8225 5551
rect 8469 5541 8545 5551
rect 8789 5541 8865 5551
rect 8949 5711 9025 5720
rect 14686 5711 14866 5721
rect 8949 5655 8959 5711
rect 9015 5655 14696 5711
rect 14752 5655 14800 5711
rect 14856 5655 14866 5711
rect 8949 5607 14866 5655
rect 8949 5551 8959 5607
rect 9015 5551 14696 5607
rect 14752 5551 14800 5607
rect 14856 5551 14866 5607
rect 8949 5540 9025 5551
rect 14686 5541 14866 5551
rect 10544 5446 10724 5456
rect 9268 5404 9344 5414
rect 10544 5404 10554 5446
rect 9268 5348 9278 5404
rect 9334 5390 10554 5404
rect 10610 5390 10658 5446
rect 10714 5390 10724 5446
rect 9334 5348 10724 5390
rect 9268 5338 9344 5348
rect 10544 5342 10724 5348
rect -16666 5117 -3143 5277
rect 10544 5286 10554 5342
rect 10610 5286 10658 5342
rect 10714 5286 10724 5342
rect 10544 5276 10724 5286
rect 17334 5446 17514 5456
rect 24120 5446 24300 5456
rect 17334 5390 17344 5446
rect 17400 5390 17448 5446
rect 17504 5390 24130 5446
rect 24186 5390 24234 5446
rect 24290 5390 24300 5446
rect 17334 5342 24300 5390
rect 17334 5286 17344 5342
rect 17400 5286 17448 5342
rect 17504 5286 24130 5342
rect 24186 5286 24234 5342
rect 24290 5286 24300 5342
rect 17334 5276 17514 5286
rect 24120 5276 24300 5286
rect 3047 5175 3227 5185
rect 7989 5175 8065 5184
rect 3047 5119 3057 5175
rect 3113 5119 3161 5175
rect 3217 5119 7999 5175
rect 8055 5119 8065 5175
rect 3047 5071 8065 5119
rect 3047 5015 3057 5071
rect 3113 5015 3161 5071
rect 3217 5015 7999 5071
rect 8055 5015 8065 5071
rect 3047 5005 3227 5015
rect 7989 5004 8065 5015
rect 8149 5175 8225 5185
rect 8469 5175 8545 5185
rect 8789 5175 8865 5185
rect 9109 5175 9185 5185
rect 8149 5119 8159 5175
rect 8215 5119 8479 5175
rect 8535 5119 8799 5175
rect 8855 5119 9119 5175
rect 9175 5119 9185 5175
rect 8149 5071 9185 5119
rect 8149 5015 8159 5071
rect 8215 5015 8479 5071
rect 8535 5015 8799 5071
rect 8855 5015 9119 5071
rect 9175 5015 9185 5071
rect 8149 5005 8225 5015
rect 8469 5005 8545 5015
rect 8789 5005 8865 5015
rect 9109 5005 9185 5015
rect 10278 4920 10458 4930
rect 9071 4868 9147 4878
rect 10278 4868 10288 4920
rect 9071 4812 9081 4868
rect 9137 4864 10288 4868
rect 10344 4864 10392 4920
rect 10448 4864 10458 4920
rect 9137 4816 10458 4864
rect 9137 4812 10288 4816
rect 9071 4802 9147 4812
rect 10278 4760 10288 4812
rect 10344 4760 10392 4816
rect 10448 4760 10458 4816
rect 10278 4750 10458 4760
rect 7829 4639 7905 4649
rect 8149 4639 8225 4649
rect 8469 4639 8545 4649
rect 8789 4639 8865 4649
rect 9109 4639 9185 4649
rect 7829 4583 7839 4639
rect 7895 4583 8159 4639
rect 8215 4583 8479 4639
rect 8535 4583 8799 4639
rect 8855 4583 9119 4639
rect 9175 4583 9185 4639
rect 7829 4535 9185 4583
rect 7829 4479 7839 4535
rect 7895 4479 8159 4535
rect 8215 4479 8479 4535
rect 8535 4479 8799 4535
rect 8855 4479 9119 4535
rect 9175 4479 9185 4535
rect 7829 4469 7905 4479
rect 8149 4469 8225 4479
rect 8469 4469 8545 4479
rect 8789 4469 8865 4479
rect 9109 4469 9185 4479
rect 14212 4466 21736 4476
rect -3626 4429 -3414 4452
rect -3626 4373 -3604 4429
rect -3548 4373 -3494 4429
rect -3438 4373 -3414 4429
rect -3626 4319 -3414 4373
rect -3626 4263 -3604 4319
rect -3548 4263 -3494 4319
rect -3438 4263 -3414 4319
rect -3626 4240 -3414 4263
rect 2715 4421 2791 4431
rect 5620 4421 5800 4431
rect 2715 4365 2725 4421
rect 2781 4365 5630 4421
rect 5686 4365 5734 4421
rect 5790 4365 5800 4421
rect 14212 4410 14222 4466
rect 14278 4410 14326 4466
rect 14382 4410 14430 4466
rect 14486 4410 21670 4466
rect 21726 4410 21736 4466
rect 2715 4317 5800 4365
rect 10544 4386 10724 4396
rect 2715 4261 2725 4317
rect 2781 4261 5630 4317
rect 5686 4261 5734 4317
rect 5790 4261 5800 4317
rect 9189 4334 9265 4344
rect 10544 4334 10554 4386
rect 9189 4278 9199 4334
rect 9255 4330 10554 4334
rect 10610 4330 10658 4386
rect 10714 4330 10724 4386
rect 9255 4282 10724 4330
rect 9255 4278 10554 4282
rect 9189 4268 9265 4278
rect 2715 4251 2791 4261
rect 5620 4251 5800 4261
rect 10544 4226 10554 4278
rect 10610 4226 10658 4282
rect 10714 4226 10724 4282
rect 10544 4216 10724 4226
rect 14212 4362 21736 4410
rect 14212 4306 14222 4362
rect 14278 4306 14326 4362
rect 14382 4306 14430 4362
rect 14486 4306 21670 4362
rect 21726 4306 21736 4362
rect 14212 4258 21736 4306
rect 14212 4202 14222 4258
rect 14278 4202 14326 4258
rect 14382 4202 14430 4258
rect 14486 4202 21670 4258
rect 21726 4202 21736 4258
rect 14212 4192 21736 4202
rect 4011 4131 4087 4141
rect 6093 4131 6273 4141
rect 4011 4075 4021 4131
rect 4077 4075 6103 4131
rect 6159 4075 6207 4131
rect 6263 4075 6273 4131
rect 30288 4139 32566 4149
rect 4011 4027 6273 4075
rect 4011 3971 4021 4027
rect 4077 3971 6103 4027
rect 6159 3971 6207 4027
rect 6263 3971 6273 4027
rect 4011 3961 4087 3971
rect 6093 3961 6273 3971
rect 6544 4103 6724 4113
rect 6854 4103 7034 4113
rect 7829 4104 7905 4113
rect 8149 4104 8225 4113
rect 8469 4104 8545 4113
rect 8789 4104 8865 4113
rect 9109 4104 9185 4113
rect 7829 4103 9185 4104
rect 6544 4047 6554 4103
rect 6610 4047 6658 4103
rect 6714 4047 6864 4103
rect 6920 4047 6968 4103
rect 7024 4047 7839 4103
rect 7895 4047 8159 4103
rect 8215 4047 8479 4103
rect 8535 4047 8799 4103
rect 8855 4047 9119 4103
rect 9175 4047 9185 4103
rect 6544 3999 9185 4047
rect 6544 3943 6554 3999
rect 6610 3943 6658 3999
rect 6714 3943 6864 3999
rect 6920 3943 6968 3999
rect 7024 3943 7839 3999
rect 7895 3943 8159 3999
rect 8215 3943 8479 3999
rect 8535 3943 8799 3999
rect 8855 3943 9119 3999
rect 9175 3943 9185 3999
rect 6544 3933 6724 3943
rect 6854 3933 7034 3943
rect 7829 3933 7905 3943
rect 8149 3933 8225 3943
rect 8469 3933 8545 3943
rect 8789 3933 8865 3943
rect 9109 3933 9185 3943
rect 30288 4083 30298 4139
rect 30354 4083 30402 4139
rect 30458 4083 30506 4139
rect 30562 4083 30610 4139
rect 30666 4083 30714 4139
rect 30770 4083 32084 4139
rect 32140 4083 32188 4139
rect 32244 4083 32292 4139
rect 32348 4083 32396 4139
rect 32452 4083 32500 4139
rect 32556 4083 32566 4139
rect 30288 4035 32566 4083
rect 30288 3979 30298 4035
rect 30354 3979 30402 4035
rect 30458 3979 30506 4035
rect 30562 3979 30610 4035
rect 30666 3979 30714 4035
rect 30770 3979 32084 4035
rect 32140 3979 32188 4035
rect 32244 3979 32292 4035
rect 32348 3979 32396 4035
rect 32452 3979 32500 4035
rect 32556 3979 32566 4035
rect 30288 3931 32566 3979
rect 9268 3902 9344 3912
rect 10006 3902 10186 3912
rect 10278 3902 10458 3910
rect 9268 3846 9278 3902
rect 9334 3846 10016 3902
rect 10072 3846 10120 3902
rect 10176 3900 10458 3902
rect 10176 3846 10288 3900
rect 9268 3844 10288 3846
rect 10344 3844 10392 3900
rect 10448 3844 10458 3900
rect 3579 3807 3655 3817
rect 5384 3807 5564 3817
rect 3579 3751 3589 3807
rect 3645 3751 5394 3807
rect 5450 3751 5498 3807
rect 5554 3751 5564 3807
rect 3579 3703 5564 3751
rect 9268 3798 10458 3844
rect 9268 3742 9278 3798
rect 9334 3742 10016 3798
rect 10072 3742 10120 3798
rect 10176 3796 10458 3798
rect 10176 3742 10288 3796
rect 9268 3732 9344 3742
rect 10006 3732 10186 3742
rect 10278 3740 10288 3742
rect 10344 3740 10392 3796
rect 10448 3740 10458 3796
rect 10278 3730 10458 3740
rect 30288 3875 30298 3931
rect 30354 3875 30402 3931
rect 30458 3875 30506 3931
rect 30562 3875 30610 3931
rect 30666 3875 30714 3931
rect 30770 3875 32084 3931
rect 32140 3875 32188 3931
rect 32244 3875 32292 3931
rect 32348 3875 32396 3931
rect 32452 3875 32500 3931
rect 32556 3875 32566 3931
rect 30288 3827 32566 3875
rect 30288 3771 30298 3827
rect 30354 3771 30402 3827
rect 30458 3771 30506 3827
rect 30562 3771 30610 3827
rect 30666 3771 30714 3827
rect 30770 3771 32084 3827
rect 32140 3771 32188 3827
rect 32244 3771 32292 3827
rect 32348 3771 32396 3827
rect 32452 3771 32500 3827
rect 32556 3771 32566 3827
rect 3579 3647 3589 3703
rect 3645 3647 5394 3703
rect 5450 3647 5498 3703
rect 5554 3647 5564 3703
rect 30288 3723 32566 3771
rect 30288 3667 30298 3723
rect 30354 3667 30402 3723
rect 30458 3667 30506 3723
rect 30562 3667 30610 3723
rect 30666 3667 30714 3723
rect 30770 3667 32084 3723
rect 32140 3667 32188 3723
rect 32244 3667 32292 3723
rect 32348 3667 32396 3723
rect 32452 3667 32500 3723
rect 32556 3667 32566 3723
rect 30288 3657 32566 3667
rect 3579 3637 3655 3647
rect 5384 3637 5564 3647
rect 5851 3613 6031 3623
rect 5851 3557 5861 3613
rect 5917 3557 5965 3613
rect 6021 3567 6031 3613
rect 8949 3567 9025 3577
rect 6021 3557 8959 3567
rect 5851 3511 8959 3557
rect 9015 3511 9025 3567
rect 5851 3509 9025 3511
rect 5851 3453 5861 3509
rect 5917 3453 5965 3509
rect 6021 3463 9025 3509
rect 6021 3453 8959 3463
rect 3419 3405 3599 3415
rect 5851 3407 8959 3453
rect 9015 3407 9025 3463
rect 5851 3405 6031 3407
rect 3419 3349 3429 3405
rect 3485 3349 3533 3405
rect 3589 3349 5861 3405
rect 5917 3349 5965 3405
rect 6021 3349 6031 3405
rect 8949 3396 9025 3407
rect 15052 3564 34838 3574
rect 15052 3508 15062 3564
rect 15118 3508 15670 3564
rect 15726 3508 16278 3564
rect 16334 3508 34640 3564
rect 34696 3508 34744 3564
rect 34800 3508 34838 3564
rect 15052 3460 34838 3508
rect 15052 3404 15062 3460
rect 15118 3404 15670 3460
rect 15726 3404 16278 3460
rect 16334 3404 34640 3460
rect 34696 3404 34744 3460
rect 34800 3404 34838 3460
rect 3419 3301 6031 3349
rect 3419 3245 3429 3301
rect 3485 3245 3533 3301
rect 3589 3245 5861 3301
rect 5917 3245 5965 3301
rect 6021 3245 6031 3301
rect 3419 3235 3599 3245
rect 5851 3235 6031 3245
rect 9268 3387 9344 3397
rect 10544 3387 10724 3397
rect 15052 3394 34838 3404
rect 9268 3331 9278 3387
rect 9334 3331 10554 3387
rect 10610 3331 10658 3387
rect 10714 3331 10724 3387
rect 9268 3283 10724 3331
rect 9268 3227 9278 3283
rect 9334 3227 10554 3283
rect 10610 3227 10658 3283
rect 10714 3227 10724 3283
rect 9268 3217 9344 3227
rect 10544 3217 10724 3227
rect 1227 3161 1407 3171
rect 2725 3161 2801 3171
rect 9739 3161 9919 3171
rect 1227 3105 1237 3161
rect 1293 3105 1341 3161
rect 1397 3105 2735 3161
rect 2791 3105 9749 3161
rect 9805 3105 9853 3161
rect 9909 3105 9919 3161
rect 1227 3057 9919 3105
rect 1227 3001 1237 3057
rect 1293 3001 1341 3057
rect 1397 3001 2735 3057
rect 2791 3001 9749 3057
rect 9805 3001 9853 3057
rect 9909 3001 9919 3057
rect 1227 2991 1407 3001
rect 2725 2991 2801 3001
rect 9739 2991 9919 3001
rect 15556 3164 20854 3174
rect 15556 3108 15566 3164
rect 15622 3108 15670 3164
rect 15726 3108 15774 3164
rect 15830 3108 20580 3164
rect 20636 3108 20684 3164
rect 20740 3108 20788 3164
rect 20844 3108 20854 3164
rect 15556 3060 20854 3108
rect 15556 3004 15566 3060
rect 15622 3004 15670 3060
rect 15726 3004 15774 3060
rect 15830 3004 20580 3060
rect 20636 3004 20684 3060
rect 20740 3004 20788 3060
rect 20844 3004 20854 3060
rect 15556 2956 20854 3004
rect 15556 2900 15566 2956
rect 15622 2900 15670 2956
rect 15726 2900 15774 2956
rect 15830 2900 20580 2956
rect 20636 2900 20684 2956
rect 20740 2900 20788 2956
rect 20844 2900 20854 2956
rect 6093 2889 6273 2899
rect 7118 2889 7298 2899
rect 15556 2890 20854 2900
rect 6093 2833 6103 2889
rect 6159 2833 6207 2889
rect 6263 2833 7128 2889
rect 7184 2833 7232 2889
rect 7288 2833 7298 2889
rect 6093 2785 7298 2833
rect 6093 2729 6103 2785
rect 6159 2729 6207 2785
rect 6263 2729 7128 2785
rect 7184 2729 7232 2785
rect 7288 2729 7298 2785
rect 6093 2719 6273 2729
rect 7118 2719 7298 2729
rect 8869 2711 8945 2721
rect 10006 2711 10186 2721
rect 8869 2655 8879 2711
rect 8935 2655 10016 2711
rect 10072 2655 10120 2711
rect 10176 2655 10186 2711
rect 8869 2607 10186 2655
rect 3923 2545 3999 2555
rect 5144 2545 5324 2555
rect 3923 2489 3933 2545
rect 3989 2489 5154 2545
rect 5210 2489 5258 2545
rect 5314 2489 5324 2545
rect 8869 2551 8879 2607
rect 8935 2551 10016 2607
rect 10072 2551 10120 2607
rect 10176 2551 10186 2607
rect 8869 2541 8945 2551
rect 10006 2541 10186 2551
rect 3923 2441 5324 2489
rect 3923 2385 3933 2441
rect 3989 2385 5154 2441
rect 5210 2385 5258 2441
rect 5314 2385 5324 2441
rect 3923 2375 3999 2385
rect 5144 2375 5324 2385
rect 5384 2402 5564 2412
rect 6582 2402 6658 2412
rect 5384 2346 5394 2402
rect 5450 2346 5498 2402
rect 5554 2346 6592 2402
rect 6648 2346 6658 2402
rect 5384 2298 6658 2346
rect 5384 2242 5394 2298
rect 5450 2242 5498 2298
rect 5554 2242 6592 2298
rect 6648 2242 6658 2298
rect 5384 2232 5564 2242
rect 6582 2232 6658 2242
rect 13100 2296 15173 2306
rect 13100 2240 13110 2296
rect 13166 2240 14899 2296
rect 14955 2240 15003 2296
rect 15059 2240 15107 2296
rect 15163 2240 15173 2296
rect 13100 2192 15173 2240
rect -8178 2103 -7966 2137
rect -8178 2047 -8163 2103
rect -8107 2047 -8053 2103
rect -7997 2047 -7966 2103
rect -8178 1993 -7966 2047
rect 13100 2136 13110 2192
rect 13166 2136 14899 2192
rect 14955 2136 15003 2192
rect 15059 2136 15107 2192
rect 15163 2136 15173 2192
rect 13100 2088 15173 2136
rect 13100 2032 13110 2088
rect 13166 2032 14899 2088
rect 14955 2032 15003 2088
rect 15059 2032 15107 2088
rect 15163 2032 15173 2088
rect -8178 1937 -8163 1993
rect -8107 1937 -8053 1993
rect -7997 1937 -7966 1993
rect -8178 1925 -7966 1937
rect 5144 2016 5324 2026
rect 6512 2016 6692 2026
rect 13100 2022 15173 2032
rect 15556 2296 15840 2306
rect 15556 2240 15566 2296
rect 15622 2240 15670 2296
rect 15726 2240 15774 2296
rect 15830 2240 15840 2296
rect 15556 2192 15840 2240
rect 15556 2136 15566 2192
rect 15622 2136 15670 2192
rect 15726 2136 15774 2192
rect 15830 2136 15840 2192
rect 15556 2088 15840 2136
rect 15556 2032 15566 2088
rect 15622 2032 15670 2088
rect 15726 2032 15774 2088
rect 15830 2032 15840 2088
rect 15556 2022 15840 2032
rect 16171 2258 21096 2268
rect 16171 2202 16181 2258
rect 16237 2202 16285 2258
rect 16341 2202 16389 2258
rect 16445 2202 19110 2258
rect 19166 2202 19430 2258
rect 19486 2202 19750 2258
rect 19806 2202 20070 2258
rect 20126 2202 20390 2258
rect 20446 2202 20710 2258
rect 20766 2202 21030 2258
rect 21086 2202 21096 2258
rect 16171 2154 21096 2202
rect 16171 2098 16181 2154
rect 16237 2098 16285 2154
rect 16341 2098 16389 2154
rect 16445 2098 19110 2154
rect 19166 2098 19430 2154
rect 19486 2098 19750 2154
rect 19806 2098 20070 2154
rect 20126 2098 20390 2154
rect 20446 2098 20710 2154
rect 20766 2098 21030 2154
rect 21086 2098 21096 2154
rect 16171 2050 21096 2098
rect 5144 1960 5154 2016
rect 5210 1960 5258 2016
rect 5314 1960 6522 2016
rect 6578 1960 6626 2016
rect 6682 1960 6692 2016
rect 5144 1912 6692 1960
rect 5144 1856 5154 1912
rect 5210 1856 5258 1912
rect 5314 1856 6522 1912
rect 6578 1856 6626 1912
rect 6682 1856 6692 1912
rect 5144 1846 5324 1856
rect 6512 1846 6692 1856
rect 7118 2006 7298 2016
rect 9396 2006 9576 2016
rect 10918 2006 11098 2016
rect 11305 2006 11485 2016
rect 7118 1950 7128 2006
rect 7184 1950 7232 2006
rect 7288 1950 9406 2006
rect 9462 1950 9510 2006
rect 9566 1950 10928 2006
rect 10984 1950 11032 2006
rect 11088 1950 11315 2006
rect 11371 1950 11419 2006
rect 11475 1950 11485 2006
rect 16171 1994 16181 2050
rect 16237 1994 16285 2050
rect 16341 1994 16389 2050
rect 16445 1994 19110 2050
rect 19166 1994 19430 2050
rect 19486 1994 19750 2050
rect 19806 1994 20070 2050
rect 20126 1994 20390 2050
rect 20446 1994 20710 2050
rect 20766 1994 21030 2050
rect 21086 1994 21096 2050
rect 16171 1984 21096 1994
rect 30288 2127 42796 2137
rect 30288 2071 30298 2127
rect 30354 2071 30402 2127
rect 30458 2071 30506 2127
rect 30562 2071 30610 2127
rect 30666 2071 30714 2127
rect 30770 2071 42508 2127
rect 42564 2071 42612 2127
rect 42668 2071 42716 2127
rect 42772 2071 42796 2127
rect 30288 2023 42796 2071
rect 7118 1902 11485 1950
rect 7118 1846 7128 1902
rect 7184 1846 7232 1902
rect 7288 1846 9406 1902
rect 9462 1846 9510 1902
rect 9566 1846 10928 1902
rect 10984 1846 11032 1902
rect 11088 1846 11315 1902
rect 11371 1846 11419 1902
rect 11475 1846 11485 1902
rect 7118 1836 7298 1846
rect 9396 1836 9576 1846
rect 10918 1836 11098 1846
rect 11305 1836 11485 1846
rect 30288 1967 30298 2023
rect 30354 1967 30402 2023
rect 30458 1967 30506 2023
rect 30562 1967 30610 2023
rect 30666 1967 30714 2023
rect 30770 1967 42508 2023
rect 42564 1967 42612 2023
rect 42668 1967 42716 2023
rect 42772 1967 42796 2023
rect 30288 1919 42796 1967
rect 30288 1863 30298 1919
rect 30354 1863 30402 1919
rect 30458 1863 30506 1919
rect 30562 1863 30610 1919
rect 30666 1863 30714 1919
rect 30770 1863 42508 1919
rect 42564 1863 42612 1919
rect 42668 1863 42716 1919
rect 42772 1863 42796 1919
rect 30288 1815 42796 1863
rect 3971 1775 4047 1785
rect 6422 1775 6498 1783
rect 3971 1719 3981 1775
rect 4037 1773 6498 1775
rect 4037 1719 6432 1773
rect 3971 1717 6432 1719
rect 6488 1717 6498 1773
rect 3971 1671 6498 1717
rect 3971 1615 3981 1671
rect 4037 1669 6498 1671
rect 4037 1615 6432 1669
rect 3971 1605 4047 1615
rect 6422 1613 6432 1615
rect 6488 1613 6498 1669
rect 6422 1603 6498 1613
rect 6854 1767 7034 1777
rect 6854 1711 6864 1767
rect 6920 1711 6968 1767
rect 7024 1711 7034 1767
rect 6854 1663 7034 1711
rect 6854 1607 6864 1663
rect 6920 1607 6968 1663
rect 7024 1607 7034 1663
rect 30288 1759 30298 1815
rect 30354 1759 30402 1815
rect 30458 1759 30506 1815
rect 30562 1759 30610 1815
rect 30666 1759 30714 1815
rect 30770 1759 42508 1815
rect 42564 1759 42612 1815
rect 42668 1759 42716 1815
rect 42772 1759 42796 1815
rect 30288 1711 42796 1759
rect 30288 1655 30298 1711
rect 30354 1655 30402 1711
rect 30458 1655 30506 1711
rect 30562 1655 30610 1711
rect 30666 1655 30714 1711
rect 30770 1655 42508 1711
rect 42564 1655 42612 1711
rect 42668 1655 42716 1711
rect 42772 1655 42796 1711
rect 30288 1645 42796 1655
rect 6854 1597 7034 1607
rect 45022 1203 45514 1213
rect 45022 1147 45032 1203
rect 45088 1147 45136 1203
rect 45192 1147 45240 1203
rect 45296 1147 45344 1203
rect 45400 1147 45448 1203
rect 45504 1147 45514 1203
rect 6370 1129 6550 1139
rect 12018 1129 12198 1139
rect 6370 1073 6380 1129
rect 6436 1073 6484 1129
rect 6540 1073 12028 1129
rect 12084 1073 12132 1129
rect 12188 1073 12198 1129
rect 6370 1025 12198 1073
rect 6370 969 6380 1025
rect 6436 969 6484 1025
rect 6540 969 12028 1025
rect 12084 969 12132 1025
rect 12188 969 12198 1025
rect 6370 959 6550 969
rect 12018 959 12198 969
rect 35192 1103 35684 1113
rect 35192 1047 35202 1103
rect 35258 1047 35306 1103
rect 35362 1047 35410 1103
rect 35466 1047 35514 1103
rect 35570 1047 35618 1103
rect 35674 1047 35684 1103
rect 35192 999 35684 1047
rect 35192 943 35202 999
rect 35258 943 35306 999
rect 35362 943 35410 999
rect 35466 943 35514 999
rect 35570 943 35618 999
rect 35674 943 35684 999
rect 35192 895 35684 943
rect 5620 877 5800 887
rect 10313 877 10493 887
rect 5620 821 5630 877
rect 5686 821 5734 877
rect 5790 821 10323 877
rect 10379 821 10427 877
rect 10483 821 10493 877
rect 5620 773 10493 821
rect 35192 839 35202 895
rect 35258 839 35306 895
rect 35362 839 35410 895
rect 35466 839 35514 895
rect 35570 839 35618 895
rect 35674 839 35684 895
rect 35192 797 35684 839
rect 39632 1103 40124 1113
rect 39632 1047 39642 1103
rect 39698 1047 39746 1103
rect 39802 1047 39850 1103
rect 39906 1047 39954 1103
rect 40010 1047 40058 1103
rect 40114 1047 40124 1103
rect 39632 999 40124 1047
rect 39632 943 39642 999
rect 39698 943 39746 999
rect 39802 943 39850 999
rect 39906 943 39954 999
rect 40010 943 40058 999
rect 40114 943 40124 999
rect 39632 895 40124 943
rect 39632 839 39642 895
rect 39698 839 39746 895
rect 39802 839 39850 895
rect 39906 839 39954 895
rect 40010 839 40058 895
rect 40114 839 40124 895
rect 39632 797 40124 839
rect 24118 791 40124 797
rect 24118 787 35202 791
rect 5620 717 5630 773
rect 5686 717 5734 773
rect 5790 717 10323 773
rect 10379 717 10427 773
rect 10483 717 10493 773
rect 5620 707 5800 717
rect 10313 707 10493 717
rect 14889 774 21915 784
rect 14889 718 14899 774
rect 14955 718 15003 774
rect 15059 718 15107 774
rect 15163 718 21641 774
rect 21697 718 21745 774
rect 21801 718 21849 774
rect 21905 718 21915 774
rect 14889 670 21915 718
rect 14889 614 14899 670
rect 14955 614 15003 670
rect 15059 614 15107 670
rect 15163 614 21641 670
rect 21697 614 21745 670
rect 21801 614 21849 670
rect 21905 614 21915 670
rect 5144 557 13380 567
rect 5144 501 5154 557
rect 5210 501 5258 557
rect 5314 501 13210 557
rect 13266 501 13314 557
rect 13370 501 13380 557
rect 5144 453 13380 501
rect 14889 566 21915 614
rect 14889 510 14899 566
rect 14955 510 15003 566
rect 15059 510 15107 566
rect 15163 510 21641 566
rect 21697 510 21745 566
rect 21801 510 21849 566
rect 21905 510 21915 566
rect 24118 731 24128 787
rect 24184 731 24232 787
rect 24288 731 31228 787
rect 31284 731 31332 787
rect 31388 731 31436 787
rect 31492 735 35202 787
rect 35258 735 35306 791
rect 35362 735 35410 791
rect 35466 735 35514 791
rect 35570 735 35618 791
rect 35674 735 39642 791
rect 39698 735 39746 791
rect 39802 735 39850 791
rect 39906 735 39954 791
rect 40010 735 40058 791
rect 40114 735 40124 791
rect 31492 731 40124 735
rect 24118 687 40124 731
rect 45022 1099 45514 1147
rect 45022 1043 45032 1099
rect 45088 1043 45136 1099
rect 45192 1043 45240 1099
rect 45296 1043 45344 1099
rect 45400 1043 45448 1099
rect 45504 1043 45514 1099
rect 45022 995 45514 1043
rect 45022 939 45032 995
rect 45088 939 45136 995
rect 45192 939 45240 995
rect 45296 939 45344 995
rect 45400 939 45448 995
rect 45504 939 45514 995
rect 45022 891 45514 939
rect 45022 835 45032 891
rect 45088 835 45136 891
rect 45192 835 45240 891
rect 45296 835 45344 891
rect 45400 835 45448 891
rect 45504 835 45514 891
rect 45022 787 45514 835
rect 45022 731 45032 787
rect 45088 731 45136 787
rect 45192 731 45240 787
rect 45296 731 45344 787
rect 45400 731 45448 787
rect 45504 731 45514 787
rect 45022 721 45514 731
rect 49462 1203 49954 1213
rect 49462 1147 49472 1203
rect 49528 1147 49576 1203
rect 49632 1147 49680 1203
rect 49736 1147 49784 1203
rect 49840 1147 49888 1203
rect 49944 1147 49954 1203
rect 49462 1099 49954 1147
rect 49462 1043 49472 1099
rect 49528 1043 49576 1099
rect 49632 1043 49680 1099
rect 49736 1043 49784 1099
rect 49840 1043 49888 1099
rect 49944 1043 49954 1099
rect 49462 995 49954 1043
rect 49462 939 49472 995
rect 49528 939 49576 995
rect 49632 939 49680 995
rect 49736 939 49784 995
rect 49840 939 49888 995
rect 49944 939 49954 995
rect 49462 891 49954 939
rect 49462 835 49472 891
rect 49528 835 49576 891
rect 49632 835 49680 891
rect 49736 835 49784 891
rect 49840 835 49888 891
rect 49944 835 49954 891
rect 49462 787 49954 835
rect 49462 731 49472 787
rect 49528 731 49576 787
rect 49632 731 49680 787
rect 49736 731 49784 787
rect 49840 731 49888 787
rect 49944 731 49954 787
rect 49462 721 49954 731
rect 24118 683 35202 687
rect 24118 627 24128 683
rect 24184 627 24232 683
rect 24288 627 31228 683
rect 31284 627 31332 683
rect 31388 627 31436 683
rect 31492 631 35202 683
rect 35258 631 35306 687
rect 35362 631 35410 687
rect 35466 631 35514 687
rect 35570 631 35618 687
rect 35674 631 39642 687
rect 39698 631 39746 687
rect 39802 631 39850 687
rect 39906 631 39954 687
rect 40010 631 40058 687
rect 40114 631 40124 687
rect 31492 627 40124 631
rect 24118 621 40124 627
rect 24118 579 40106 621
rect 24118 523 24128 579
rect 24184 523 24232 579
rect 24288 523 31228 579
rect 31284 523 31332 579
rect 31388 523 31436 579
rect 31492 523 40106 579
rect 24118 513 40106 523
rect 14889 500 21915 510
rect 5144 397 5154 453
rect 5210 397 5258 453
rect 5314 397 13210 453
rect 13266 397 13314 453
rect 13370 397 13380 453
rect 5144 387 13380 397
rect 45095 396 45379 721
rect 49576 396 49860 721
rect 24568 386 49985 396
rect 24568 330 24578 386
rect 24634 330 24682 386
rect 24738 330 32136 386
rect 32192 330 32240 386
rect 32296 330 32344 386
rect 32400 330 49985 386
rect 24568 282 49985 330
rect 24568 226 24578 282
rect 24634 226 24682 282
rect 24738 226 32136 282
rect 32192 226 32240 282
rect 32296 226 32344 282
rect 32400 226 49985 282
rect 24568 178 49985 226
rect 24568 122 24578 178
rect 24634 122 24682 178
rect 24738 122 32136 178
rect 32192 122 32240 178
rect 32296 122 32344 178
rect 32400 122 49985 178
rect 24568 112 49985 122
<< via3 >>
rect -8163 12999 -8107 13055
rect -8053 12999 -7997 13055
rect -8163 12889 -8107 12945
rect -8053 12889 -7997 12945
rect -3604 10673 -3548 10729
rect -3494 10673 -3438 10729
rect -3604 10563 -3548 10619
rect -3494 10563 -3438 10619
rect -8141 9655 -8085 9711
rect -8031 9655 -7975 9711
rect -8141 9550 -8085 9606
rect -8031 9550 -7975 9606
rect -8141 9445 -8085 9501
rect -8031 9445 -7975 9501
rect -8491 8726 -8435 8782
rect -8381 8726 -8325 8782
rect -8491 8616 -8435 8672
rect -8381 8616 -8325 8672
rect -8491 8506 -8435 8562
rect -8381 8506 -8325 8562
rect -8491 8396 -8435 8452
rect -8381 8396 -8325 8452
rect -10576 7864 -10520 7920
rect -10466 7864 -10410 7920
rect -10356 7864 -10300 7920
rect -10246 7864 -10190 7920
rect -10576 7754 -10520 7810
rect -10466 7754 -10410 7810
rect -10356 7754 -10300 7810
rect -10246 7754 -10190 7810
rect -8146 5476 -8090 5532
rect -8041 5476 -7985 5532
rect -7936 5476 -7880 5532
rect -8146 5366 -8090 5422
rect -8041 5366 -7985 5422
rect -7936 5366 -7880 5422
rect -3604 4373 -3548 4429
rect -3494 4373 -3438 4429
rect -3604 4263 -3548 4319
rect -3494 4263 -3438 4319
rect 32084 4083 32140 4139
rect 32188 4083 32244 4139
rect 32292 4083 32348 4139
rect 32396 4083 32452 4139
rect 32500 4083 32556 4139
rect 32084 3979 32140 4035
rect 32188 3979 32244 4035
rect 32292 3979 32348 4035
rect 32396 3979 32452 4035
rect 32500 3979 32556 4035
rect 32084 3875 32140 3931
rect 32188 3875 32244 3931
rect 32292 3875 32348 3931
rect 32396 3875 32452 3931
rect 32500 3875 32556 3931
rect 32084 3771 32140 3827
rect 32188 3771 32244 3827
rect 32292 3771 32348 3827
rect 32396 3771 32452 3827
rect 32500 3771 32556 3827
rect 32084 3667 32140 3723
rect 32188 3667 32244 3723
rect 32292 3667 32348 3723
rect 32396 3667 32452 3723
rect 32500 3667 32556 3723
rect -8163 2047 -8107 2103
rect -8053 2047 -7997 2103
rect -8163 1937 -8107 1993
rect -8053 1937 -7997 1993
rect 42508 2071 42564 2127
rect 42612 2071 42668 2127
rect 42716 2071 42772 2127
rect 42508 1967 42564 2023
rect 42612 1967 42668 2023
rect 42716 1967 42772 2023
rect 42508 1863 42564 1919
rect 42612 1863 42668 1919
rect 42716 1863 42772 1919
rect 42508 1759 42564 1815
rect 42612 1759 42668 1815
rect 42716 1759 42772 1815
rect 42508 1655 42564 1711
rect 42612 1655 42668 1711
rect 42716 1655 42772 1711
rect 45032 1147 45088 1203
rect 45136 1147 45192 1203
rect 45240 1147 45296 1203
rect 45344 1147 45400 1203
rect 45448 1147 45504 1203
rect 35202 1047 35258 1103
rect 35306 1047 35362 1103
rect 35410 1047 35466 1103
rect 35514 1047 35570 1103
rect 35618 1047 35674 1103
rect 35202 943 35258 999
rect 35306 943 35362 999
rect 35410 943 35466 999
rect 35514 943 35570 999
rect 35618 943 35674 999
rect 35202 839 35258 895
rect 35306 839 35362 895
rect 35410 839 35466 895
rect 35514 839 35570 895
rect 35618 839 35674 895
rect 39642 1047 39698 1103
rect 39746 1047 39802 1103
rect 39850 1047 39906 1103
rect 39954 1047 40010 1103
rect 40058 1047 40114 1103
rect 39642 943 39698 999
rect 39746 943 39802 999
rect 39850 943 39906 999
rect 39954 943 40010 999
rect 40058 943 40114 999
rect 39642 839 39698 895
rect 39746 839 39802 895
rect 39850 839 39906 895
rect 39954 839 40010 895
rect 40058 839 40114 895
rect 35202 735 35258 791
rect 35306 735 35362 791
rect 35410 735 35466 791
rect 35514 735 35570 791
rect 35618 735 35674 791
rect 39642 735 39698 791
rect 39746 735 39802 791
rect 39850 735 39906 791
rect 39954 735 40010 791
rect 40058 735 40114 791
rect 45032 1043 45088 1099
rect 45136 1043 45192 1099
rect 45240 1043 45296 1099
rect 45344 1043 45400 1099
rect 45448 1043 45504 1099
rect 45032 939 45088 995
rect 45136 939 45192 995
rect 45240 939 45296 995
rect 45344 939 45400 995
rect 45448 939 45504 995
rect 45032 835 45088 891
rect 45136 835 45192 891
rect 45240 835 45296 891
rect 45344 835 45400 891
rect 45448 835 45504 891
rect 45032 731 45088 787
rect 45136 731 45192 787
rect 45240 731 45296 787
rect 45344 731 45400 787
rect 45448 731 45504 787
rect 49472 1147 49528 1203
rect 49576 1147 49632 1203
rect 49680 1147 49736 1203
rect 49784 1147 49840 1203
rect 49888 1147 49944 1203
rect 49472 1043 49528 1099
rect 49576 1043 49632 1099
rect 49680 1043 49736 1099
rect 49784 1043 49840 1099
rect 49888 1043 49944 1099
rect 49472 939 49528 995
rect 49576 939 49632 995
rect 49680 939 49736 995
rect 49784 939 49840 995
rect 49888 939 49944 995
rect 49472 835 49528 891
rect 49576 835 49632 891
rect 49680 835 49736 891
rect 49784 835 49840 891
rect 49888 835 49944 891
rect 49472 731 49528 787
rect 49576 731 49632 787
rect 49680 731 49736 787
rect 49784 731 49840 787
rect 49888 731 49944 787
rect 35202 631 35258 687
rect 35306 631 35362 687
rect 35410 631 35466 687
rect 35514 631 35570 687
rect 35618 631 35674 687
rect 39642 631 39698 687
rect 39746 631 39802 687
rect 39850 631 39906 687
rect 39954 631 40010 687
rect 40058 631 40114 687
<< metal4 >>
rect -12206 14878 -8526 14945
rect -12206 14825 -8676 14878
rect -16290 14681 -12610 14748
rect -16290 14628 -12760 14681
rect -16290 11588 -16170 14628
rect -12970 11588 -12760 14628
rect -16290 11535 -12760 11588
rect -12672 11535 -12610 14681
rect -12206 11785 -12086 14825
rect -8886 11785 -8676 14825
rect -12206 11732 -8676 11785
rect -8588 11732 -8526 14878
rect -7719 14561 -4439 14681
rect -8178 13055 -7966 13067
rect -8178 12999 -8163 13055
rect -8107 12999 -8053 13055
rect -7997 12999 -7966 13055
rect -8178 12945 -7966 12999
rect -8178 12889 -8163 12945
rect -8107 12889 -8053 12945
rect -7997 12889 -7966 12945
rect -8178 12855 -7966 12889
rect -12206 11665 -8526 11732
rect -16290 11468 -12610 11535
rect -12206 11478 -8526 11545
rect -12206 11425 -8676 11478
rect -16290 11281 -12610 11348
rect -16290 11228 -12760 11281
rect -16290 8188 -16170 11228
rect -12970 8188 -12760 11228
rect -16290 8135 -12760 8188
rect -12672 8135 -12610 11281
rect -12206 8385 -12086 11425
rect -8886 8385 -8676 11425
rect -12206 8332 -8676 8385
rect -8588 8796 -8526 11478
rect -7719 11361 -7599 14561
rect -4559 11361 -4439 14561
rect -7719 11151 -4439 11361
rect -7719 11063 -7652 11151
rect -4506 11063 -4439 11151
rect -7719 11001 -4439 11063
rect -4319 14561 -1039 14681
rect -4319 11361 -4199 14561
rect -1159 11361 -1039 14561
rect -4319 11151 -1039 11361
rect -4319 11063 -4252 11151
rect -1106 11063 -1039 11151
rect -4319 11001 -1039 11063
rect -3626 10729 -3414 10752
rect -3626 10673 -3604 10729
rect -3548 10673 -3494 10729
rect -3438 10673 -3414 10729
rect -3626 10619 -3414 10673
rect -3626 10563 -3604 10619
rect -3548 10563 -3494 10619
rect -3438 10563 -3414 10619
rect -3626 10540 -3414 10563
rect -8154 9711 -7942 9721
rect -8154 9655 -8141 9711
rect -8085 9655 -8031 9711
rect -7975 9655 -7942 9711
rect -8154 9606 -7942 9655
rect -8154 9550 -8141 9606
rect -8085 9550 -8031 9606
rect -7975 9550 -7942 9606
rect -8154 9501 -7942 9550
rect -8154 9445 -8141 9501
rect -8085 9445 -8031 9501
rect -7975 9445 -7942 9501
rect -8154 9430 -7942 9445
rect -8588 8794 -8375 8796
rect -8588 8782 -8303 8794
rect -8588 8726 -8491 8782
rect -8435 8726 -8381 8782
rect -8325 8726 -8303 8782
rect -8588 8672 -8303 8726
rect -8588 8616 -8491 8672
rect -8435 8616 -8381 8672
rect -8325 8616 -8303 8672
rect -8588 8562 -8303 8616
rect -8588 8506 -8491 8562
rect -8435 8506 -8381 8562
rect -8325 8506 -8303 8562
rect -8588 8452 -8303 8506
rect -8588 8396 -8491 8452
rect -8435 8396 -8381 8452
rect -8325 8396 -8303 8452
rect -8588 8368 -8303 8396
rect -8588 8366 -8373 8368
rect -8588 8332 -8526 8366
rect -12206 8265 -8526 8332
rect -16290 8068 -12610 8135
rect -12822 7200 -12610 8068
rect -10593 7920 -10178 7946
rect -10593 7864 -10576 7920
rect -10520 7864 -10466 7920
rect -10410 7864 -10356 7920
rect -10300 7864 -10246 7920
rect -10190 7864 -10178 7920
rect -10593 7810 -10178 7864
rect -10593 7754 -10576 7810
rect -10520 7754 -10466 7810
rect -10410 7754 -10356 7810
rect -10300 7754 -10246 7810
rect -10190 7754 -10178 7810
rect -10593 7721 -10178 7754
rect -16290 7133 -12610 7200
rect -16290 7080 -12760 7133
rect -16290 4040 -16170 7080
rect -12970 4040 -12760 7080
rect -16290 3987 -12760 4040
rect -12672 3987 -12610 7133
rect -16290 3920 -12610 3987
rect -12186 7170 -8506 7237
rect -12186 7117 -8656 7170
rect -12186 4077 -12066 7117
rect -8866 4077 -8656 7117
rect -12186 4024 -8656 4077
rect -8568 4024 -8506 7170
rect 33218 6013 37658 6133
rect -8159 5532 -7863 5550
rect -8159 5476 -8146 5532
rect -8090 5476 -8041 5532
rect -7985 5476 -7936 5532
rect -7880 5476 -7863 5532
rect -8159 5422 -7863 5476
rect -8159 5366 -8146 5422
rect -8090 5366 -8041 5422
rect -7985 5366 -7936 5422
rect -7880 5366 -7863 5422
rect -8159 5338 -7863 5366
rect -3626 4429 -3414 4452
rect -3626 4373 -3604 4429
rect -3548 4373 -3494 4429
rect -3438 4373 -3414 4429
rect -3626 4319 -3414 4373
rect -3626 4263 -3604 4319
rect -3548 4263 -3494 4319
rect -3438 4263 -3414 4319
rect -3626 4240 -3414 4263
rect -12186 3957 -8506 4024
rect 32074 4139 32566 4149
rect 32074 4083 32084 4139
rect 32140 4083 32188 4139
rect 32244 4083 32292 4139
rect 32348 4083 32396 4139
rect 32452 4083 32500 4139
rect 32556 4083 32566 4139
rect 32074 4035 32566 4083
rect -7719 3929 -4439 3991
rect -7719 3841 -7652 3929
rect -4506 3841 -4439 3929
rect -16290 3733 -12610 3800
rect -16290 3680 -12760 3733
rect -16290 640 -16170 3680
rect -12970 640 -12760 3680
rect -16290 587 -12760 640
rect -12672 587 -12610 3733
rect -16290 520 -12610 587
rect -12186 3770 -8506 3837
rect -12186 3717 -8656 3770
rect -12186 677 -12066 3717
rect -8866 677 -8656 3717
rect -12186 624 -8656 677
rect -8568 624 -8506 3770
rect -7719 3631 -4439 3841
rect -8178 2103 -7966 2137
rect -8178 2047 -8163 2103
rect -8107 2047 -8053 2103
rect -7997 2047 -7966 2103
rect -8178 1993 -7966 2047
rect -8178 1937 -8163 1993
rect -8107 1937 -8053 1993
rect -7997 1937 -7966 1993
rect -8178 1925 -7966 1937
rect -12186 557 -8506 624
rect -7719 431 -7599 3631
rect -4559 431 -4439 3631
rect -7719 311 -4439 431
rect -4319 3929 -1039 3991
rect -4319 3841 -4252 3929
rect -1106 3841 -1039 3929
rect -4319 3631 -1039 3841
rect 32074 3979 32084 4035
rect 32140 3979 32188 4035
rect 32244 3979 32292 4035
rect 32348 3979 32396 4035
rect 32452 3979 32500 4035
rect 32556 3979 32566 4035
rect 32074 3931 32566 3979
rect 32074 3875 32084 3931
rect 32140 3875 32188 3931
rect 32244 3875 32292 3931
rect 32348 3875 32396 3931
rect 32452 3875 32500 3931
rect 32556 3875 32566 3931
rect 32074 3827 32566 3875
rect 32074 3771 32084 3827
rect 32140 3771 32188 3827
rect 32244 3771 32292 3827
rect 32348 3771 32396 3827
rect 32452 3771 32500 3827
rect 32556 3771 32566 3827
rect 32074 3723 32566 3771
rect 32074 3667 32084 3723
rect 32140 3667 32188 3723
rect 32244 3667 32292 3723
rect 32348 3667 32396 3723
rect 32452 3667 32500 3723
rect 32556 3667 32566 3723
rect 32074 3657 32566 3667
rect -4319 431 -4199 3631
rect -1159 431 -1039 3631
rect 33218 1813 33338 6013
rect 37538 1813 37658 6013
rect 33218 1603 37658 1813
rect 33218 1515 33285 1603
rect 37591 1515 37658 1603
rect 33218 1453 37658 1515
rect 37778 6013 42218 6133
rect 37778 1813 37898 6013
rect 42098 1813 42218 6013
rect 43048 6013 47488 6133
rect 37778 1603 42218 1813
rect 42462 4139 42796 4149
rect 42462 4083 42508 4139
rect 42564 4083 42612 4139
rect 42668 4083 42716 4139
rect 42772 4083 42796 4139
rect 42462 4035 42796 4083
rect 42462 3979 42508 4035
rect 42564 3979 42612 4035
rect 42668 3979 42716 4035
rect 42772 3979 42796 4035
rect 42462 3931 42796 3979
rect 42462 3875 42508 3931
rect 42564 3875 42612 3931
rect 42668 3875 42716 3931
rect 42772 3875 42796 3931
rect 42462 3827 42796 3875
rect 42462 3771 42508 3827
rect 42564 3771 42612 3827
rect 42668 3771 42716 3827
rect 42772 3771 42796 3827
rect 42462 3723 42796 3771
rect 42462 3667 42508 3723
rect 42564 3667 42612 3723
rect 42668 3667 42716 3723
rect 42772 3667 42796 3723
rect 42462 2127 42796 3667
rect 42462 2071 42508 2127
rect 42564 2071 42612 2127
rect 42668 2071 42716 2127
rect 42772 2071 42796 2127
rect 42462 2023 42796 2071
rect 42462 1967 42508 2023
rect 42564 1967 42612 2023
rect 42668 1967 42716 2023
rect 42772 1967 42796 2023
rect 42462 1919 42796 1967
rect 42462 1863 42508 1919
rect 42564 1863 42612 1919
rect 42668 1863 42716 1919
rect 42772 1863 42796 1919
rect 42462 1815 42796 1863
rect 42462 1759 42508 1815
rect 42564 1759 42612 1815
rect 42668 1759 42716 1815
rect 42772 1759 42796 1815
rect 42462 1711 42796 1759
rect 42462 1655 42508 1711
rect 42564 1655 42612 1711
rect 42668 1655 42716 1711
rect 42772 1655 42796 1711
rect 42462 1645 42796 1655
rect 43048 1813 43168 6013
rect 47368 1813 47488 6013
rect 37778 1515 37845 1603
rect 42151 1515 42218 1603
rect 37778 1453 42218 1515
rect 43048 1603 47488 1813
rect 43048 1515 43115 1603
rect 47421 1515 47488 1603
rect 43048 1453 47488 1515
rect 47608 6013 52048 6133
rect 47608 1813 47728 6013
rect 51928 1813 52048 6013
rect 47608 1603 52048 1813
rect 47608 1515 47675 1603
rect 51981 1515 52048 1603
rect 47608 1453 52048 1515
rect 35192 1103 35684 1453
rect 35192 1047 35202 1103
rect 35258 1047 35306 1103
rect 35362 1047 35410 1103
rect 35466 1047 35514 1103
rect 35570 1047 35618 1103
rect 35674 1047 35684 1103
rect 35192 999 35684 1047
rect 35192 943 35202 999
rect 35258 943 35306 999
rect 35362 943 35410 999
rect 35466 943 35514 999
rect 35570 943 35618 999
rect 35674 943 35684 999
rect 35192 895 35684 943
rect 35192 839 35202 895
rect 35258 839 35306 895
rect 35362 839 35410 895
rect 35466 839 35514 895
rect 35570 839 35618 895
rect 35674 839 35684 895
rect 35192 791 35684 839
rect 35192 735 35202 791
rect 35258 735 35306 791
rect 35362 735 35410 791
rect 35466 735 35514 791
rect 35570 735 35618 791
rect 35674 735 35684 791
rect 35192 687 35684 735
rect 35192 631 35202 687
rect 35258 631 35306 687
rect 35362 631 35410 687
rect 35466 631 35514 687
rect 35570 631 35618 687
rect 35674 631 35684 687
rect 35192 621 35684 631
rect 39632 1103 40124 1453
rect 39632 1047 39642 1103
rect 39698 1047 39746 1103
rect 39802 1047 39850 1103
rect 39906 1047 39954 1103
rect 40010 1047 40058 1103
rect 40114 1047 40124 1103
rect 39632 999 40124 1047
rect 39632 943 39642 999
rect 39698 943 39746 999
rect 39802 943 39850 999
rect 39906 943 39954 999
rect 40010 943 40058 999
rect 40114 943 40124 999
rect 39632 895 40124 943
rect 39632 839 39642 895
rect 39698 839 39746 895
rect 39802 839 39850 895
rect 39906 839 39954 895
rect 40010 839 40058 895
rect 40114 839 40124 895
rect 39632 791 40124 839
rect 39632 735 39642 791
rect 39698 735 39746 791
rect 39802 735 39850 791
rect 39906 735 39954 791
rect 40010 735 40058 791
rect 40114 735 40124 791
rect 39632 687 40124 735
rect 45022 1203 45514 1453
rect 45022 1147 45032 1203
rect 45088 1147 45136 1203
rect 45192 1147 45240 1203
rect 45296 1147 45344 1203
rect 45400 1147 45448 1203
rect 45504 1147 45514 1203
rect 45022 1099 45514 1147
rect 45022 1043 45032 1099
rect 45088 1043 45136 1099
rect 45192 1043 45240 1099
rect 45296 1043 45344 1099
rect 45400 1043 45448 1099
rect 45504 1043 45514 1099
rect 45022 995 45514 1043
rect 45022 939 45032 995
rect 45088 939 45136 995
rect 45192 939 45240 995
rect 45296 939 45344 995
rect 45400 939 45448 995
rect 45504 939 45514 995
rect 45022 891 45514 939
rect 45022 835 45032 891
rect 45088 835 45136 891
rect 45192 835 45240 891
rect 45296 835 45344 891
rect 45400 835 45448 891
rect 45504 835 45514 891
rect 45022 787 45514 835
rect 45022 731 45032 787
rect 45088 731 45136 787
rect 45192 731 45240 787
rect 45296 731 45344 787
rect 45400 731 45448 787
rect 45504 731 45514 787
rect 45022 721 45514 731
rect 49462 1203 49954 1453
rect 49462 1147 49472 1203
rect 49528 1147 49576 1203
rect 49632 1147 49680 1203
rect 49736 1147 49784 1203
rect 49840 1147 49888 1203
rect 49944 1147 49954 1203
rect 49462 1099 49954 1147
rect 49462 1043 49472 1099
rect 49528 1043 49576 1099
rect 49632 1043 49680 1099
rect 49736 1043 49784 1099
rect 49840 1043 49888 1099
rect 49944 1043 49954 1099
rect 49462 995 49954 1043
rect 49462 939 49472 995
rect 49528 939 49576 995
rect 49632 939 49680 995
rect 49736 939 49784 995
rect 49840 939 49888 995
rect 49944 939 49954 995
rect 49462 891 49954 939
rect 49462 835 49472 891
rect 49528 835 49576 891
rect 49632 835 49680 891
rect 49736 835 49784 891
rect 49840 835 49888 891
rect 49944 835 49954 891
rect 49462 787 49954 835
rect 49462 731 49472 787
rect 49528 731 49576 787
rect 49632 731 49680 787
rect 49736 731 49784 787
rect 49840 731 49888 787
rect 49944 731 49954 787
rect 49462 721 49954 731
rect 39632 631 39642 687
rect 39698 631 39746 687
rect 39802 631 39850 687
rect 39906 631 39954 687
rect 40010 631 40058 687
rect 40114 631 40124 687
rect 39632 621 40124 631
rect -4319 311 -1039 431
<< via4 >>
rect -12760 11535 -12672 14681
rect -8676 11732 -8588 14878
rect -8163 12999 -8107 13055
rect -8053 12999 -7997 13055
rect -8163 12889 -8107 12945
rect -8053 12889 -7997 12945
rect -12760 8135 -12672 11281
rect -8676 8332 -8588 11478
rect -7652 11063 -4506 11151
rect -4252 11063 -1106 11151
rect -3604 10673 -3548 10729
rect -3494 10673 -3438 10729
rect -3604 10563 -3548 10619
rect -3494 10563 -3438 10619
rect -8141 9655 -8085 9711
rect -8031 9655 -7975 9711
rect -8141 9550 -8085 9606
rect -8031 9550 -7975 9606
rect -8141 9445 -8085 9501
rect -8031 9445 -7975 9501
rect -8491 8726 -8435 8782
rect -8381 8726 -8325 8782
rect -8491 8616 -8435 8672
rect -8381 8616 -8325 8672
rect -8491 8506 -8435 8562
rect -8381 8506 -8325 8562
rect -8491 8396 -8435 8452
rect -8381 8396 -8325 8452
rect -10576 7864 -10520 7920
rect -10466 7864 -10410 7920
rect -10356 7864 -10300 7920
rect -10246 7864 -10190 7920
rect -10576 7754 -10520 7810
rect -10466 7754 -10410 7810
rect -10356 7754 -10300 7810
rect -10246 7754 -10190 7810
rect -12760 3987 -12672 7133
rect -8656 4024 -8568 7170
rect -8146 5476 -8090 5532
rect -8041 5476 -7985 5532
rect -7936 5476 -7880 5532
rect -8146 5366 -8090 5422
rect -8041 5366 -7985 5422
rect -7936 5366 -7880 5422
rect -3604 4373 -3548 4429
rect -3494 4373 -3438 4429
rect -3604 4263 -3548 4319
rect -3494 4263 -3438 4319
rect 32084 4083 32140 4139
rect 32188 4083 32244 4139
rect 32292 4083 32348 4139
rect 32396 4083 32452 4139
rect 32500 4083 32556 4139
rect -7652 3841 -4506 3929
rect -12760 587 -12672 3733
rect -8656 624 -8568 3770
rect -8163 2047 -8107 2103
rect -8053 2047 -7997 2103
rect -8163 1937 -8107 1993
rect -8053 1937 -7997 1993
rect -4252 3841 -1106 3929
rect 32084 3979 32140 4035
rect 32188 3979 32244 4035
rect 32292 3979 32348 4035
rect 32396 3979 32452 4035
rect 32500 3979 32556 4035
rect 32084 3875 32140 3931
rect 32188 3875 32244 3931
rect 32292 3875 32348 3931
rect 32396 3875 32452 3931
rect 32500 3875 32556 3931
rect 32084 3771 32140 3827
rect 32188 3771 32244 3827
rect 32292 3771 32348 3827
rect 32396 3771 32452 3827
rect 32500 3771 32556 3827
rect 32084 3667 32140 3723
rect 32188 3667 32244 3723
rect 32292 3667 32348 3723
rect 32396 3667 32452 3723
rect 32500 3667 32556 3723
rect 33285 1515 37591 1603
rect 42508 4083 42564 4139
rect 42612 4083 42668 4139
rect 42716 4083 42772 4139
rect 42508 3979 42564 4035
rect 42612 3979 42668 4035
rect 42716 3979 42772 4035
rect 42508 3875 42564 3931
rect 42612 3875 42668 3931
rect 42716 3875 42772 3931
rect 42508 3771 42564 3827
rect 42612 3771 42668 3827
rect 42716 3771 42772 3827
rect 42508 3667 42564 3723
rect 42612 3667 42668 3723
rect 42716 3667 42772 3723
rect 42508 2071 42564 2127
rect 42612 2071 42668 2127
rect 42716 2071 42772 2127
rect 42508 1967 42564 2023
rect 42612 1967 42668 2023
rect 42716 1967 42772 2023
rect 42508 1863 42564 1919
rect 42612 1863 42668 1919
rect 42716 1863 42772 1919
rect 42508 1759 42564 1815
rect 42612 1759 42668 1815
rect 42716 1759 42772 1815
rect 42508 1655 42564 1711
rect 42612 1655 42668 1711
rect 42716 1655 42772 1711
rect 37845 1515 42151 1603
rect 43115 1515 47421 1603
rect 47675 1515 51981 1603
<< metal5 >>
rect -14676 14548 -14464 14808
rect -12822 14681 -12610 14808
rect -10592 14745 -10380 15005
rect -8738 14878 -8526 15005
rect -14676 11148 -14464 11668
rect -12822 11535 -12760 14681
rect -12672 11535 -12610 14681
rect -12822 11281 -12610 11535
rect -10592 11345 -10380 11865
rect -8738 11732 -8676 14878
rect -8588 11732 -8526 14878
rect -8178 13055 -7519 13067
rect -8178 12999 -8163 13055
rect -8107 12999 -8053 13055
rect -7997 12999 -7519 13055
rect -8178 12945 -7519 12999
rect -8178 12889 -8163 12945
rect -8107 12889 -8053 12945
rect -7997 12889 -7519 12945
rect -8178 12855 -7519 12889
rect -8738 11478 -8526 11732
rect -14676 7611 -14464 8268
rect -12822 8135 -12760 11281
rect -12672 8135 -12610 11281
rect -12822 8008 -12610 8135
rect -10592 7946 -10380 8465
rect -8738 8332 -8676 11478
rect -8588 8796 -8526 11478
rect -4639 12855 -4119 13067
rect -1239 12855 -979 13067
rect -7779 11151 -979 11213
rect -7779 11063 -7652 11151
rect -4506 11063 -4252 11151
rect -1106 11063 -979 11151
rect -7779 11001 -979 11063
rect -3601 10752 -3444 11001
rect -3626 10729 -3414 10752
rect -3626 10673 -3604 10729
rect -3548 10673 -3494 10729
rect -3438 10673 -3414 10729
rect -3626 10619 -3414 10673
rect -3626 10563 -3604 10619
rect -3548 10563 -3494 10619
rect -3438 10563 -3414 10619
rect -3626 10540 -3414 10563
rect -8154 9711 -7942 9721
rect -8154 9655 -8141 9711
rect -8085 9655 -8031 9711
rect -7975 9655 -7942 9711
rect -8154 9606 -7942 9655
rect -8154 9550 -8141 9606
rect -8085 9550 -8031 9606
rect -7975 9550 -7942 9606
rect -8154 9501 -7942 9550
rect -8154 9445 -8141 9501
rect -8085 9445 -8031 9501
rect -7975 9445 -7942 9501
rect -8588 8794 -8375 8796
rect -8588 8782 -8303 8794
rect -8588 8726 -8491 8782
rect -8435 8726 -8381 8782
rect -8325 8726 -8303 8782
rect -8588 8672 -8303 8726
rect -8588 8616 -8491 8672
rect -8435 8616 -8381 8672
rect -8325 8616 -8303 8672
rect -8588 8562 -8303 8616
rect -8588 8506 -8491 8562
rect -8435 8506 -8381 8562
rect -8325 8506 -8303 8562
rect -8588 8452 -8303 8506
rect -8588 8396 -8491 8452
rect -8435 8396 -8381 8452
rect -8325 8396 -8303 8452
rect -8588 8368 -8303 8396
rect -8588 8366 -8373 8368
rect -8588 8332 -8526 8366
rect -8738 8205 -8526 8332
rect -10593 7920 -10178 7946
rect -10593 7864 -10576 7920
rect -10520 7864 -10466 7920
rect -10410 7864 -10356 7920
rect -10300 7864 -10246 7920
rect -10190 7864 -10178 7920
rect -10593 7810 -10178 7864
rect -10593 7754 -10576 7810
rect -10520 7754 -10466 7810
rect -10410 7754 -10356 7810
rect -10300 7754 -10246 7810
rect -10190 7754 -10178 7810
rect -10593 7721 -10178 7754
rect -8154 7611 -7942 9445
rect -14676 7399 -7942 7611
rect -14676 7000 -14464 7399
rect -12822 7133 -12610 7260
rect -14676 3600 -14464 4120
rect -12822 3987 -12760 7133
rect -12672 3987 -12610 7133
rect -10572 7037 -10360 7399
rect -8718 7170 -8506 7297
rect -12822 3733 -12610 3987
rect -14676 460 -14464 720
rect -12822 587 -12760 3733
rect -12672 587 -12610 3733
rect -10572 3637 -10360 4157
rect -8718 4024 -8656 7170
rect -8568 5550 -8506 7170
rect -8568 5532 -7863 5550
rect -8568 5476 -8146 5532
rect -8090 5476 -8041 5532
rect -7985 5476 -7936 5532
rect -7880 5476 -7863 5532
rect -8568 5422 -7863 5476
rect -8568 5366 -8146 5422
rect -8090 5366 -8041 5422
rect -7985 5366 -7936 5422
rect -7880 5366 -7863 5422
rect -8568 5338 -7863 5366
rect -8568 4024 -8506 5338
rect -3626 4429 -3414 4452
rect -3626 4373 -3604 4429
rect -3548 4373 -3494 4429
rect -3438 4373 -3414 4429
rect -3626 4319 -3414 4373
rect -3626 4263 -3604 4319
rect -3548 4263 -3494 4319
rect -3438 4263 -3414 4319
rect -3626 4240 -3414 4263
rect -8718 3770 -8506 4024
rect -3596 3991 -3439 4240
rect 32074 4139 33298 4149
rect 32074 4083 32084 4139
rect 32140 4083 32188 4139
rect 32244 4083 32292 4139
rect 32348 4083 32396 4139
rect 32452 4083 32500 4139
rect 32556 4083 33298 4139
rect 32074 4035 33298 4083
rect -7779 3929 -979 3991
rect -7779 3841 -7652 3929
rect -4506 3841 -4252 3929
rect -1106 3841 -979 3929
rect -7779 3779 -979 3841
rect 32074 3979 32084 4035
rect 32140 3979 32188 4035
rect 32244 3979 32292 4035
rect 32348 3979 32396 4035
rect 32452 3979 32500 4035
rect 32556 4019 33298 4035
rect 32556 3979 33418 4019
rect 32074 3931 33418 3979
rect 32074 3875 32084 3931
rect 32140 3875 32188 3931
rect 32244 3875 32292 3931
rect 32348 3875 32396 3931
rect 32452 3875 32500 3931
rect 32556 3875 33418 3931
rect 32074 3827 33418 3875
rect -12822 402 -12610 587
rect -10572 497 -10360 757
rect -8718 624 -8656 3770
rect -8568 624 -8506 3770
rect 32074 3771 32084 3827
rect 32140 3771 32188 3827
rect 32244 3771 32292 3827
rect 32348 3771 32396 3827
rect 32452 3771 32500 3827
rect 32556 3807 33418 3827
rect 32556 3771 33298 3807
rect 32074 3723 33298 3771
rect 32074 3667 32084 3723
rect 32140 3667 32188 3723
rect 32244 3667 32292 3723
rect 32348 3667 32396 3723
rect 32452 3667 32500 3723
rect 32556 3667 33298 3723
rect 32074 3657 33298 3667
rect -8178 2103 -7519 2137
rect -8178 2047 -8163 2103
rect -8107 2047 -8053 2103
rect -7997 2047 -7519 2103
rect -8178 1993 -7519 2047
rect -8178 1937 -8163 1993
rect -8107 1937 -8053 1993
rect -7997 1937 -7519 1993
rect -8178 1925 -7519 1937
rect -8718 402 -8506 624
rect -4639 1925 -4119 2137
rect -1239 1925 -979 2137
rect 37458 3807 37978 4019
rect 42462 4139 43128 4149
rect 42462 4083 42508 4139
rect 42564 4083 42612 4139
rect 42668 4083 42716 4139
rect 42772 4083 43128 4139
rect 42462 4035 43128 4083
rect 42018 3807 42278 4019
rect 42462 3979 42508 4035
rect 42564 3979 42612 4035
rect 42668 3979 42716 4035
rect 42772 4019 43128 4035
rect 42772 3979 43248 4019
rect 42462 3931 43248 3979
rect 42462 3875 42508 3931
rect 42564 3875 42612 3931
rect 42668 3875 42716 3931
rect 42772 3875 43248 3931
rect 42462 3827 43248 3875
rect 42462 3771 42508 3827
rect 42564 3771 42612 3827
rect 42668 3771 42716 3827
rect 42772 3807 43248 3827
rect 42772 3771 43128 3807
rect 42462 3723 43128 3771
rect 42462 3667 42508 3723
rect 42564 3667 42612 3723
rect 42668 3667 42716 3723
rect 42772 3667 43128 3723
rect 42462 3657 43128 3667
rect 42462 2127 42796 2137
rect 42462 2071 42508 2127
rect 42564 2071 42612 2127
rect 42668 2071 42716 2127
rect 42772 2071 42796 2127
rect 42462 2023 42796 2071
rect 42462 1967 42508 2023
rect 42564 1967 42612 2023
rect 42668 1967 42716 2023
rect 42772 1967 42796 2023
rect 42462 1919 42796 1967
rect 42462 1863 42508 1919
rect 42564 1863 42612 1919
rect 42668 1863 42716 1919
rect 42772 1863 42796 1919
rect 47288 3807 47808 4019
rect 51848 3807 52108 4019
rect 42462 1815 42796 1863
rect 42462 1759 42508 1815
rect 42564 1759 42612 1815
rect 42668 1759 42716 1815
rect 42772 1759 42796 1815
rect 42462 1711 42796 1759
rect 33158 1603 42278 1665
rect 42462 1655 42508 1711
rect 42564 1655 42612 1711
rect 42668 1655 42716 1711
rect 42772 1655 42796 1711
rect 42462 1645 42796 1655
rect 33158 1515 33285 1603
rect 37591 1515 37845 1603
rect 42151 1515 42278 1603
rect 33158 1453 42278 1515
rect 42988 1603 52108 1665
rect 42988 1515 43115 1603
rect 47421 1515 47675 1603
rect 51981 1515 52108 1603
rect 42988 1453 52108 1515
rect -12825 190 -8506 402
<< labels >>
flabel metal1 33652 15036 33652 15036 0 FreeSans 1600 0 0 0 VOUT_N
port 5 nsew
flabel metal1 32948 15654 32948 15654 0 FreeSans 1600 0 0 0 VOUT_P
port 6 nsew
flabel metal1 38509 14010 38509 14010 0 FreeSans 1600 0 0 0 VDD
port 7 nsew
flabel metal1 16460 14550 16460 14550 0 FreeSans 1600 0 0 0 VSS
port 9 nsew
flabel metal1 -1080 10090 -1080 10090 0 FreeSans 1600 0 0 0 VOUT_OPAMP_P
port 11 nsew
flabel metal2 -3040 7540 -3040 7540 0 FreeSans 1600 0 0 0 VOUT_OPAMP_N
port 12 nsew
flabel metal2 -16437 5875 -16437 5875 0 FreeSans 1600 0 0 0 VIN_N1
port 1 nsew
flabel metal2 -17125 -191 -17125 -191 0 FreeSans 1600 0 0 0 IBIAS1
port 1 nsew
flabel metal3 -16560 5220 -16560 5220 0 FreeSans 1600 0 0 0 VCM1
port 13 nsew
flabel metal2 -16600 9060 -16600 9060 0 FreeSans 1600 0 0 0 VIN_P1
port 14 nsew
flabel metal2 -7400 5460 -7400 5460 0 FreeSans 1600 0 0 0 R3_R7_1
port 15 nsew
flabel metal2 -7980 6330 -7980 6330 0 FreeSans 1600 0 0 0 R7_R8_R10_C1
port 16 nsew
flabel metal1 3160 1980 3160 1980 0 FreeSans 1600 0 0 0 IB21
port 17 nsew
flabel metal1 2440 5270 2440 5270 0 FreeSans 1600 0 0 0 IBIAS11
port 18 nsew
flabel metal1 3130 5380 3130 5380 0 FreeSans 1600 0 0 0 VBM1
port 19 nsew
flabel metal1 5490 5430 5490 5430 0 FreeSans 1600 0 0 0 VBIASN1
port 20 nsew
flabel metal1 8940 1510 8940 1510 0 FreeSans 1600 0 0 0 IB31
port 21 nsew
flabel metal3 9880 760 9880 760 0 FreeSans 1600 0 0 0 IBS1
port 22 nsew
flabel metal1 12290 1080 12290 1080 0 FreeSans 1600 0 0 0 VB21
port 23 nsew
flabel metal1 11560 1940 11560 1940 0 FreeSans 1600 0 0 0 VB31
port 24 nsew
flabel metal1 8540 6320 8540 6320 0 FreeSans 1600 0 0 0 VB41
port 25 nsew
flabel metal1 6620 4310 6620 4310 0 FreeSans 1600 0 0 0 VCD1
port 26 nsew
flabel metal1 5800 14420 5800 14420 0 FreeSans 1600 0 0 0 IND1
port 27 nsew
flabel metal1 6130 14390 6130 14390 0 FreeSans 1600 0 0 0 IPD1
port 28 nsew
flabel metal2 11480 12040 11480 12040 0 FreeSans 1600 0 0 0 OUT2_1
port 29 nsew
flabel metal1 11710 11070 11710 11070 0 FreeSans 1600 0 0 0 OUT1_1
port 30 nsew
flabel metal1 16030 180 16030 180 0 FreeSans 1600 0 0 0 IBIAS3_1
port 32 nsew
flabel metal3 17890 4430 17890 4430 0 FreeSans 1600 0 0 0 IB4_1
port 33 nsew
flabel metal1 22190 700 22190 700 0 FreeSans 1600 0 0 0 IBIAS4_1
port 34 nsew
flabel metal3 17870 2220 17870 2220 0 FreeSans 1600 0 0 0 IVS_1
port 35 nsew
flabel metal1 67400 13010 67400 13010 0 FreeSans 1600 0 0 0 IBIAS2_1
port 36 nsew
flabel metal1 14950 5670 14950 5670 0 FreeSans 1600 0 0 0 VB1_1
port 37 nsew
flabel metal1 2400 13930 2400 13930 0 FreeSans 1600 0 0 0 BD_1
port 38 nsew
flabel metal2 -7820 8650 -7820 8650 0 FreeSans 1600 0 0 0 R_1
port 39 nsew
flabel metal5 -8120 8070 -8120 8070 0 FreeSans 1600 0 0 0 R11_1
port 40 nsew
flabel metal3 32800 1940 32800 1940 0 FreeSans 1600 0 0 0 OPAMP_C_1
port 41 nsew
flabel metal3 31560 3900 31560 3900 0 FreeSans 1600 0 0 0 OPAMP_C1_1
port 42 nsew
flabel metal1 11360 5390 11360 5390 0 FreeSans 1600 0 0 0 VOUT_1_1
port 43 nsew
flabel metal1 2418 13899 2418 13899 0 FreeSans 320 0 0 0 Folded_Diff_Op_Amp_Layout_0.BD
flabel metal1 5821 14354 5821 14354 0 FreeSans 320 0 0 0 Folded_Diff_Op_Amp_Layout_0.IND
flabel metal1 6093 14384 6093 14384 0 FreeSans 320 0 0 0 Folded_Diff_Op_Amp_Layout_0.IPD
flabel psubdiffcont 8541 7301 8541 7301 0 FreeSans 320 0 0 0 Folded_Diff_Op_Amp_Layout_0.VSS
flabel metal1 17455 11525 17455 11525 0 FreeSans 320 0 0 0 Folded_Diff_Op_Amp_Layout_0.VND
flabel metal1 17193 11457 17193 11457 0 FreeSans 320 0 0 0 Folded_Diff_Op_Amp_Layout_0.VPD
flabel metal1 12336 1051 12336 1051 0 FreeSans 320 0 0 0 Folded_Diff_Op_Amp_Layout_0.VB2
flabel metal1 2493 5232 2493 5232 0 FreeSans 320 0 0 0 Folded_Diff_Op_Amp_Layout_0.IBIAS1
flabel metal1 8595 6331 8595 6331 0 FreeSans 320 0 0 0 Folded_Diff_Op_Amp_Layout_0.VB4
flabel metal1 11627 1926 11627 1926 0 FreeSans 320 0 0 0 Folded_Diff_Op_Amp_Layout_0.VB3
flabel metal1 10864 5366 10864 5366 0 FreeSans 320 0 0 0 Folded_Diff_Op_Amp_Layout_0.VOUT
flabel metal1 3137 5325 3137 5325 0 FreeSans 320 0 0 0 Folded_Diff_Op_Amp_Layout_0.VBM
flabel metal1 6634 4253 6634 4253 0 FreeSans 320 0 0 0 Folded_Diff_Op_Amp_Layout_0.VCD
flabel metal1 5484 5383 5484 5383 0 FreeSans 320 0 0 0 Folded_Diff_Op_Amp_Layout_0.VBIASN
flabel metal1 15004 5633 15004 5633 0 FreeSans 320 0 0 0 Folded_Diff_Op_Amp_Layout_0.VB1
flabel metal1 16090 142 16090 142 0 FreeSans 320 0 0 0 Folded_Diff_Op_Amp_Layout_0.IBIAS3
flabel metal1 22195 642 22195 642 0 FreeSans 320 0 0 0 Folded_Diff_Op_Amp_Layout_0.IBIAS4
flabel nsubdiffcont 1869 10873 1869 10873 0 FreeSans 320 0 0 0 Folded_Diff_Op_Amp_Layout_0.VDD
flabel metal3 10158 787 10158 787 0 FreeSans 1600 0 0 0 Folded_Diff_Op_Amp_Layout_0.IBS
flabel metal1 31678 15565 31687 15565 0 FreeSans 1600 0 0 0 Folded_Diff_Op_Amp_Layout_0.OUT_P
flabel metal1 32640 14985 32640 14985 0 FreeSans 1600 0 0 0 Folded_Diff_Op_Amp_Layout_0.OUT_N
flabel metal1 67418 12909 67418 12909 0 FreeSans 1600 0 0 0 Folded_Diff_Op_Amp_Layout_0.IBIAS2
flabel metal1 111 7498 111 7498 0 FreeSans 1600 0 0 0 Folded_Diff_Op_Amp_Layout_0.IBIAS
flabel metal1 10577 5951 10577 5951 0 FreeSans 1600 0 0 0 Folded_Diff_Op_Amp_Layout_0.VCM
flabel metal3 17841 2113 17841 2113 0 FreeSans 800 0 0 0 Folded_Diff_Op_Amp_Layout_0.IVS
flabel metal3 17858 4327 17858 4327 0 FreeSans 800 0 0 0 Folded_Diff_Op_Amp_Layout_0.IB4
flabel metal1 3272 1982 3272 1982 0 FreeSans 800 0 0 0 Folded_Diff_Op_Amp_Layout_0.IB2
flabel metal1 9100 1513 9100 1513 0 FreeSans 800 0 0 0 Folded_Diff_Op_Amp_Layout_0.IB3
flabel metal2 5467 3504 5467 3504 0 FreeSans 800 0 0 0 Folded_Diff_Op_Amp_Layout_0.IB5
flabel metal1 2712 13110 2712 13110 0 FreeSans 1600 0 0 0 Folded_Diff_Op_Amp_Layout_0.IN_P
flabel metal1 3019 14247 3019 14247 0 FreeSans 1600 0 0 0 Folded_Diff_Op_Amp_Layout_0.IN_N
flabel metal2 11448 11552 11448 11552 0 FreeSans 1600 0 0 0 Folded_Diff_Op_Amp_Layout_0.OUT2
flabel metal1 11649 10953 11809 11675 0 FreeSans 1600 0 0 0 Folded_Diff_Op_Amp_Layout_0.OUT1
flabel metal2 -7612 5400 -7612 5400 0 FreeSans 800 0 0 0 filter_res_magic_0.R3_R7
flabel metal2 -7604 6354 -7604 6354 0 FreeSans 800 0 0 0 filter_res_magic_0.R7_R8_R10_C
flabel metal1 -5775 10629 -5775 10629 0 FreeSans 1600 0 0 0 filter_res_magic_0.VDD
flabel metal2 -7393 5902 -7393 5902 0 FreeSans 1600 0 0 0 filter_res_magic_0.VIN_N
flabel metal2 -7783 9112 -7783 9112 0 FreeSans 1600 0 0 0 filter_res_magic_0.VIN_P
flabel metal2 -3523 6272 -3523 6272 0 FreeSans 1600 0 0 0 filter_res_magic_0.VOUT_OPAMP_N
flabel metal2 -3543 8682 -3543 8682 0 FreeSans 1600 0 0 0 filter_res_magic_0.VOUT_OPAMP_P
flabel metal2 -7013 10842 -7013 10842 0 FreeSans 1600 0 0 0 filter_res_magic_0.VOUT_N
flabel metal2 -7023 4112 -7023 4112 0 FreeSans 1600 0 0 0 filter_res_magic_0.VOUT_P
<< end >>
