magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1484 -1329 1484 1329
<< metal2 >>
rect -484 324 484 329
rect -484 296 -479 324
rect -451 296 -417 324
rect -389 296 -355 324
rect -327 296 -293 324
rect -265 296 -231 324
rect -203 296 -169 324
rect -141 296 -107 324
rect -79 296 -45 324
rect -17 296 17 324
rect 45 296 79 324
rect 107 296 141 324
rect 169 296 203 324
rect 231 296 265 324
rect 293 296 327 324
rect 355 296 389 324
rect 417 296 451 324
rect 479 296 484 324
rect -484 262 484 296
rect -484 234 -479 262
rect -451 234 -417 262
rect -389 234 -355 262
rect -327 234 -293 262
rect -265 234 -231 262
rect -203 234 -169 262
rect -141 234 -107 262
rect -79 234 -45 262
rect -17 234 17 262
rect 45 234 79 262
rect 107 234 141 262
rect 169 234 203 262
rect 231 234 265 262
rect 293 234 327 262
rect 355 234 389 262
rect 417 234 451 262
rect 479 234 484 262
rect -484 200 484 234
rect -484 172 -479 200
rect -451 172 -417 200
rect -389 172 -355 200
rect -327 172 -293 200
rect -265 172 -231 200
rect -203 172 -169 200
rect -141 172 -107 200
rect -79 172 -45 200
rect -17 172 17 200
rect 45 172 79 200
rect 107 172 141 200
rect 169 172 203 200
rect 231 172 265 200
rect 293 172 327 200
rect 355 172 389 200
rect 417 172 451 200
rect 479 172 484 200
rect -484 138 484 172
rect -484 110 -479 138
rect -451 110 -417 138
rect -389 110 -355 138
rect -327 110 -293 138
rect -265 110 -231 138
rect -203 110 -169 138
rect -141 110 -107 138
rect -79 110 -45 138
rect -17 110 17 138
rect 45 110 79 138
rect 107 110 141 138
rect 169 110 203 138
rect 231 110 265 138
rect 293 110 327 138
rect 355 110 389 138
rect 417 110 451 138
rect 479 110 484 138
rect -484 76 484 110
rect -484 48 -479 76
rect -451 48 -417 76
rect -389 48 -355 76
rect -327 48 -293 76
rect -265 48 -231 76
rect -203 48 -169 76
rect -141 48 -107 76
rect -79 48 -45 76
rect -17 48 17 76
rect 45 48 79 76
rect 107 48 141 76
rect 169 48 203 76
rect 231 48 265 76
rect 293 48 327 76
rect 355 48 389 76
rect 417 48 451 76
rect 479 48 484 76
rect -484 14 484 48
rect -484 -14 -479 14
rect -451 -14 -417 14
rect -389 -14 -355 14
rect -327 -14 -293 14
rect -265 -14 -231 14
rect -203 -14 -169 14
rect -141 -14 -107 14
rect -79 -14 -45 14
rect -17 -14 17 14
rect 45 -14 79 14
rect 107 -14 141 14
rect 169 -14 203 14
rect 231 -14 265 14
rect 293 -14 327 14
rect 355 -14 389 14
rect 417 -14 451 14
rect 479 -14 484 14
rect -484 -48 484 -14
rect -484 -76 -479 -48
rect -451 -76 -417 -48
rect -389 -76 -355 -48
rect -327 -76 -293 -48
rect -265 -76 -231 -48
rect -203 -76 -169 -48
rect -141 -76 -107 -48
rect -79 -76 -45 -48
rect -17 -76 17 -48
rect 45 -76 79 -48
rect 107 -76 141 -48
rect 169 -76 203 -48
rect 231 -76 265 -48
rect 293 -76 327 -48
rect 355 -76 389 -48
rect 417 -76 451 -48
rect 479 -76 484 -48
rect -484 -110 484 -76
rect -484 -138 -479 -110
rect -451 -138 -417 -110
rect -389 -138 -355 -110
rect -327 -138 -293 -110
rect -265 -138 -231 -110
rect -203 -138 -169 -110
rect -141 -138 -107 -110
rect -79 -138 -45 -110
rect -17 -138 17 -110
rect 45 -138 79 -110
rect 107 -138 141 -110
rect 169 -138 203 -110
rect 231 -138 265 -110
rect 293 -138 327 -110
rect 355 -138 389 -110
rect 417 -138 451 -110
rect 479 -138 484 -110
rect -484 -172 484 -138
rect -484 -200 -479 -172
rect -451 -200 -417 -172
rect -389 -200 -355 -172
rect -327 -200 -293 -172
rect -265 -200 -231 -172
rect -203 -200 -169 -172
rect -141 -200 -107 -172
rect -79 -200 -45 -172
rect -17 -200 17 -172
rect 45 -200 79 -172
rect 107 -200 141 -172
rect 169 -200 203 -172
rect 231 -200 265 -172
rect 293 -200 327 -172
rect 355 -200 389 -172
rect 417 -200 451 -172
rect 479 -200 484 -172
rect -484 -234 484 -200
rect -484 -262 -479 -234
rect -451 -262 -417 -234
rect -389 -262 -355 -234
rect -327 -262 -293 -234
rect -265 -262 -231 -234
rect -203 -262 -169 -234
rect -141 -262 -107 -234
rect -79 -262 -45 -234
rect -17 -262 17 -234
rect 45 -262 79 -234
rect 107 -262 141 -234
rect 169 -262 203 -234
rect 231 -262 265 -234
rect 293 -262 327 -234
rect 355 -262 389 -234
rect 417 -262 451 -234
rect 479 -262 484 -234
rect -484 -296 484 -262
rect -484 -324 -479 -296
rect -451 -324 -417 -296
rect -389 -324 -355 -296
rect -327 -324 -293 -296
rect -265 -324 -231 -296
rect -203 -324 -169 -296
rect -141 -324 -107 -296
rect -79 -324 -45 -296
rect -17 -324 17 -296
rect 45 -324 79 -296
rect 107 -324 141 -296
rect 169 -324 203 -296
rect 231 -324 265 -296
rect 293 -324 327 -296
rect 355 -324 389 -296
rect 417 -324 451 -296
rect 479 -324 484 -296
rect -484 -329 484 -324
<< via2 >>
rect -479 296 -451 324
rect -417 296 -389 324
rect -355 296 -327 324
rect -293 296 -265 324
rect -231 296 -203 324
rect -169 296 -141 324
rect -107 296 -79 324
rect -45 296 -17 324
rect 17 296 45 324
rect 79 296 107 324
rect 141 296 169 324
rect 203 296 231 324
rect 265 296 293 324
rect 327 296 355 324
rect 389 296 417 324
rect 451 296 479 324
rect -479 234 -451 262
rect -417 234 -389 262
rect -355 234 -327 262
rect -293 234 -265 262
rect -231 234 -203 262
rect -169 234 -141 262
rect -107 234 -79 262
rect -45 234 -17 262
rect 17 234 45 262
rect 79 234 107 262
rect 141 234 169 262
rect 203 234 231 262
rect 265 234 293 262
rect 327 234 355 262
rect 389 234 417 262
rect 451 234 479 262
rect -479 172 -451 200
rect -417 172 -389 200
rect -355 172 -327 200
rect -293 172 -265 200
rect -231 172 -203 200
rect -169 172 -141 200
rect -107 172 -79 200
rect -45 172 -17 200
rect 17 172 45 200
rect 79 172 107 200
rect 141 172 169 200
rect 203 172 231 200
rect 265 172 293 200
rect 327 172 355 200
rect 389 172 417 200
rect 451 172 479 200
rect -479 110 -451 138
rect -417 110 -389 138
rect -355 110 -327 138
rect -293 110 -265 138
rect -231 110 -203 138
rect -169 110 -141 138
rect -107 110 -79 138
rect -45 110 -17 138
rect 17 110 45 138
rect 79 110 107 138
rect 141 110 169 138
rect 203 110 231 138
rect 265 110 293 138
rect 327 110 355 138
rect 389 110 417 138
rect 451 110 479 138
rect -479 48 -451 76
rect -417 48 -389 76
rect -355 48 -327 76
rect -293 48 -265 76
rect -231 48 -203 76
rect -169 48 -141 76
rect -107 48 -79 76
rect -45 48 -17 76
rect 17 48 45 76
rect 79 48 107 76
rect 141 48 169 76
rect 203 48 231 76
rect 265 48 293 76
rect 327 48 355 76
rect 389 48 417 76
rect 451 48 479 76
rect -479 -14 -451 14
rect -417 -14 -389 14
rect -355 -14 -327 14
rect -293 -14 -265 14
rect -231 -14 -203 14
rect -169 -14 -141 14
rect -107 -14 -79 14
rect -45 -14 -17 14
rect 17 -14 45 14
rect 79 -14 107 14
rect 141 -14 169 14
rect 203 -14 231 14
rect 265 -14 293 14
rect 327 -14 355 14
rect 389 -14 417 14
rect 451 -14 479 14
rect -479 -76 -451 -48
rect -417 -76 -389 -48
rect -355 -76 -327 -48
rect -293 -76 -265 -48
rect -231 -76 -203 -48
rect -169 -76 -141 -48
rect -107 -76 -79 -48
rect -45 -76 -17 -48
rect 17 -76 45 -48
rect 79 -76 107 -48
rect 141 -76 169 -48
rect 203 -76 231 -48
rect 265 -76 293 -48
rect 327 -76 355 -48
rect 389 -76 417 -48
rect 451 -76 479 -48
rect -479 -138 -451 -110
rect -417 -138 -389 -110
rect -355 -138 -327 -110
rect -293 -138 -265 -110
rect -231 -138 -203 -110
rect -169 -138 -141 -110
rect -107 -138 -79 -110
rect -45 -138 -17 -110
rect 17 -138 45 -110
rect 79 -138 107 -110
rect 141 -138 169 -110
rect 203 -138 231 -110
rect 265 -138 293 -110
rect 327 -138 355 -110
rect 389 -138 417 -110
rect 451 -138 479 -110
rect -479 -200 -451 -172
rect -417 -200 -389 -172
rect -355 -200 -327 -172
rect -293 -200 -265 -172
rect -231 -200 -203 -172
rect -169 -200 -141 -172
rect -107 -200 -79 -172
rect -45 -200 -17 -172
rect 17 -200 45 -172
rect 79 -200 107 -172
rect 141 -200 169 -172
rect 203 -200 231 -172
rect 265 -200 293 -172
rect 327 -200 355 -172
rect 389 -200 417 -172
rect 451 -200 479 -172
rect -479 -262 -451 -234
rect -417 -262 -389 -234
rect -355 -262 -327 -234
rect -293 -262 -265 -234
rect -231 -262 -203 -234
rect -169 -262 -141 -234
rect -107 -262 -79 -234
rect -45 -262 -17 -234
rect 17 -262 45 -234
rect 79 -262 107 -234
rect 141 -262 169 -234
rect 203 -262 231 -234
rect 265 -262 293 -234
rect 327 -262 355 -234
rect 389 -262 417 -234
rect 451 -262 479 -234
rect -479 -324 -451 -296
rect -417 -324 -389 -296
rect -355 -324 -327 -296
rect -293 -324 -265 -296
rect -231 -324 -203 -296
rect -169 -324 -141 -296
rect -107 -324 -79 -296
rect -45 -324 -17 -296
rect 17 -324 45 -296
rect 79 -324 107 -296
rect 141 -324 169 -296
rect 203 -324 231 -296
rect 265 -324 293 -296
rect 327 -324 355 -296
rect 389 -324 417 -296
rect 451 -324 479 -296
<< metal3 >>
rect -484 324 484 329
rect -484 296 -479 324
rect -451 296 -417 324
rect -389 296 -355 324
rect -327 296 -293 324
rect -265 296 -231 324
rect -203 296 -169 324
rect -141 296 -107 324
rect -79 296 -45 324
rect -17 296 17 324
rect 45 296 79 324
rect 107 296 141 324
rect 169 296 203 324
rect 231 296 265 324
rect 293 296 327 324
rect 355 296 389 324
rect 417 296 451 324
rect 479 296 484 324
rect -484 262 484 296
rect -484 234 -479 262
rect -451 234 -417 262
rect -389 234 -355 262
rect -327 234 -293 262
rect -265 234 -231 262
rect -203 234 -169 262
rect -141 234 -107 262
rect -79 234 -45 262
rect -17 234 17 262
rect 45 234 79 262
rect 107 234 141 262
rect 169 234 203 262
rect 231 234 265 262
rect 293 234 327 262
rect 355 234 389 262
rect 417 234 451 262
rect 479 234 484 262
rect -484 200 484 234
rect -484 172 -479 200
rect -451 172 -417 200
rect -389 172 -355 200
rect -327 172 -293 200
rect -265 172 -231 200
rect -203 172 -169 200
rect -141 172 -107 200
rect -79 172 -45 200
rect -17 172 17 200
rect 45 172 79 200
rect 107 172 141 200
rect 169 172 203 200
rect 231 172 265 200
rect 293 172 327 200
rect 355 172 389 200
rect 417 172 451 200
rect 479 172 484 200
rect -484 138 484 172
rect -484 110 -479 138
rect -451 110 -417 138
rect -389 110 -355 138
rect -327 110 -293 138
rect -265 110 -231 138
rect -203 110 -169 138
rect -141 110 -107 138
rect -79 110 -45 138
rect -17 110 17 138
rect 45 110 79 138
rect 107 110 141 138
rect 169 110 203 138
rect 231 110 265 138
rect 293 110 327 138
rect 355 110 389 138
rect 417 110 451 138
rect 479 110 484 138
rect -484 76 484 110
rect -484 48 -479 76
rect -451 48 -417 76
rect -389 48 -355 76
rect -327 48 -293 76
rect -265 48 -231 76
rect -203 48 -169 76
rect -141 48 -107 76
rect -79 48 -45 76
rect -17 48 17 76
rect 45 48 79 76
rect 107 48 141 76
rect 169 48 203 76
rect 231 48 265 76
rect 293 48 327 76
rect 355 48 389 76
rect 417 48 451 76
rect 479 48 484 76
rect -484 14 484 48
rect -484 -14 -479 14
rect -451 -14 -417 14
rect -389 -14 -355 14
rect -327 -14 -293 14
rect -265 -14 -231 14
rect -203 -14 -169 14
rect -141 -14 -107 14
rect -79 -14 -45 14
rect -17 -14 17 14
rect 45 -14 79 14
rect 107 -14 141 14
rect 169 -14 203 14
rect 231 -14 265 14
rect 293 -14 327 14
rect 355 -14 389 14
rect 417 -14 451 14
rect 479 -14 484 14
rect -484 -48 484 -14
rect -484 -76 -479 -48
rect -451 -76 -417 -48
rect -389 -76 -355 -48
rect -327 -76 -293 -48
rect -265 -76 -231 -48
rect -203 -76 -169 -48
rect -141 -76 -107 -48
rect -79 -76 -45 -48
rect -17 -76 17 -48
rect 45 -76 79 -48
rect 107 -76 141 -48
rect 169 -76 203 -48
rect 231 -76 265 -48
rect 293 -76 327 -48
rect 355 -76 389 -48
rect 417 -76 451 -48
rect 479 -76 484 -48
rect -484 -110 484 -76
rect -484 -138 -479 -110
rect -451 -138 -417 -110
rect -389 -138 -355 -110
rect -327 -138 -293 -110
rect -265 -138 -231 -110
rect -203 -138 -169 -110
rect -141 -138 -107 -110
rect -79 -138 -45 -110
rect -17 -138 17 -110
rect 45 -138 79 -110
rect 107 -138 141 -110
rect 169 -138 203 -110
rect 231 -138 265 -110
rect 293 -138 327 -110
rect 355 -138 389 -110
rect 417 -138 451 -110
rect 479 -138 484 -110
rect -484 -172 484 -138
rect -484 -200 -479 -172
rect -451 -200 -417 -172
rect -389 -200 -355 -172
rect -327 -200 -293 -172
rect -265 -200 -231 -172
rect -203 -200 -169 -172
rect -141 -200 -107 -172
rect -79 -200 -45 -172
rect -17 -200 17 -172
rect 45 -200 79 -172
rect 107 -200 141 -172
rect 169 -200 203 -172
rect 231 -200 265 -172
rect 293 -200 327 -172
rect 355 -200 389 -172
rect 417 -200 451 -172
rect 479 -200 484 -172
rect -484 -234 484 -200
rect -484 -262 -479 -234
rect -451 -262 -417 -234
rect -389 -262 -355 -234
rect -327 -262 -293 -234
rect -265 -262 -231 -234
rect -203 -262 -169 -234
rect -141 -262 -107 -234
rect -79 -262 -45 -234
rect -17 -262 17 -234
rect 45 -262 79 -234
rect 107 -262 141 -234
rect 169 -262 203 -234
rect 231 -262 265 -234
rect 293 -262 327 -234
rect 355 -262 389 -234
rect 417 -262 451 -234
rect 479 -262 484 -234
rect -484 -296 484 -262
rect -484 -324 -479 -296
rect -451 -324 -417 -296
rect -389 -324 -355 -296
rect -327 -324 -293 -296
rect -265 -324 -231 -296
rect -203 -324 -169 -296
rect -141 -324 -107 -296
rect -79 -324 -45 -296
rect -17 -324 17 -296
rect 45 -324 79 -296
rect 107 -324 141 -296
rect 169 -324 203 -296
rect 231 -324 265 -296
rect 293 -324 327 -296
rect 355 -324 389 -296
rect 417 -324 451 -296
rect 479 -324 484 -296
rect -484 -329 484 -324
<< end >>
