magic
tech gf180mcuC
magscale 1 10
timestamp 1692184121
<< nwell >>
rect -350 1262 1462 3508
<< pwell >>
rect -288 0 -8 1158
rect 0 0 1400 1158
<< nmos >>
rect -176 840 -120 1090
rect 112 840 168 1090
rect 272 840 328 1090
rect 432 840 488 1090
rect 592 840 648 1090
rect 752 840 808 1090
rect 912 840 968 1090
rect 1072 840 1128 1090
rect 1232 840 1288 1090
rect -176 454 -120 704
rect 112 454 168 704
rect 272 454 328 704
rect 432 454 488 704
rect 592 454 648 704
rect 752 454 808 704
rect 912 454 968 704
rect 1072 454 1128 704
rect 1232 454 1288 704
rect -176 68 -120 318
rect 112 68 168 318
rect 272 68 328 318
rect 432 68 488 318
rect 592 68 648 318
rect 752 68 808 318
rect 912 68 968 318
rect 1072 68 1128 318
rect 1232 68 1288 318
<< pmos >>
rect -176 2664 -120 3164
rect 112 2664 168 3164
rect 272 2664 328 3164
rect 432 2664 488 3164
rect 592 2664 648 3164
rect 752 2664 808 3164
rect 912 2664 968 3164
rect 1072 2664 1128 3164
rect 1232 2664 1288 3164
rect -176 2028 -120 2528
rect 112 2028 168 2528
rect 272 2028 328 2528
rect 432 2028 488 2528
rect 592 2028 648 2528
rect 752 2028 808 2528
rect 912 2028 968 2528
rect 1072 2028 1128 2528
rect 1232 2028 1288 2528
rect -176 1392 -120 1892
rect 112 1392 168 1892
rect 272 1392 328 1892
rect 432 1392 488 1892
rect 592 1392 648 1892
rect 752 1392 808 1892
rect 912 1392 968 1892
rect 1072 1392 1128 1892
rect 1232 1392 1288 1892
<< ndiff >>
rect -264 1077 -176 1090
rect -264 853 -251 1077
rect -205 853 -176 1077
rect -264 840 -176 853
rect -120 1077 -32 1090
rect -120 853 -91 1077
rect -45 853 -32 1077
rect -120 840 -32 853
rect 24 1077 112 1090
rect 24 853 37 1077
rect 83 853 112 1077
rect 24 840 112 853
rect 168 1077 272 1090
rect 168 853 197 1077
rect 243 853 272 1077
rect 168 840 272 853
rect 328 1077 432 1090
rect 328 853 357 1077
rect 403 853 432 1077
rect 328 840 432 853
rect 488 1077 592 1090
rect 488 853 517 1077
rect 563 853 592 1077
rect 488 840 592 853
rect 648 1077 752 1090
rect 648 853 677 1077
rect 723 853 752 1077
rect 648 840 752 853
rect 808 1077 912 1090
rect 808 853 837 1077
rect 883 853 912 1077
rect 808 840 912 853
rect 968 1077 1072 1090
rect 968 853 997 1077
rect 1043 853 1072 1077
rect 968 840 1072 853
rect 1128 1077 1232 1090
rect 1128 853 1157 1077
rect 1203 853 1232 1077
rect 1128 840 1232 853
rect 1288 1077 1376 1090
rect 1288 853 1317 1077
rect 1363 853 1376 1077
rect 1288 840 1376 853
rect -264 691 -176 704
rect -264 467 -251 691
rect -205 467 -176 691
rect -264 454 -176 467
rect -120 691 -32 704
rect -120 467 -91 691
rect -45 467 -32 691
rect -120 454 -32 467
rect 24 691 112 704
rect 24 467 37 691
rect 83 467 112 691
rect 24 454 112 467
rect 168 691 272 704
rect 168 467 197 691
rect 243 467 272 691
rect 168 454 272 467
rect 328 691 432 704
rect 328 467 357 691
rect 403 467 432 691
rect 328 454 432 467
rect 488 691 592 704
rect 488 467 517 691
rect 563 467 592 691
rect 488 454 592 467
rect 648 691 752 704
rect 648 467 677 691
rect 723 467 752 691
rect 648 454 752 467
rect 808 691 912 704
rect 808 467 837 691
rect 883 467 912 691
rect 808 454 912 467
rect 968 691 1072 704
rect 968 467 997 691
rect 1043 467 1072 691
rect 968 454 1072 467
rect 1128 691 1232 704
rect 1128 467 1157 691
rect 1203 467 1232 691
rect 1128 454 1232 467
rect 1288 691 1376 704
rect 1288 467 1317 691
rect 1363 467 1376 691
rect 1288 454 1376 467
rect -264 305 -176 318
rect -264 81 -251 305
rect -205 81 -176 305
rect -264 68 -176 81
rect -120 305 -32 318
rect -120 81 -91 305
rect -45 81 -32 305
rect -120 68 -32 81
rect 24 305 112 318
rect 24 81 37 305
rect 83 81 112 305
rect 24 68 112 81
rect 168 305 272 318
rect 168 81 197 305
rect 243 81 272 305
rect 168 68 272 81
rect 328 305 432 318
rect 328 81 357 305
rect 403 81 432 305
rect 328 68 432 81
rect 488 305 592 318
rect 488 81 517 305
rect 563 81 592 305
rect 488 68 592 81
rect 648 305 752 318
rect 648 81 677 305
rect 723 81 752 305
rect 648 68 752 81
rect 808 305 912 318
rect 808 81 837 305
rect 883 81 912 305
rect 808 68 912 81
rect 968 305 1072 318
rect 968 81 997 305
rect 1043 81 1072 305
rect 968 68 1072 81
rect 1128 305 1232 318
rect 1128 81 1157 305
rect 1203 81 1232 305
rect 1128 68 1232 81
rect 1288 305 1376 318
rect 1288 81 1317 305
rect 1363 81 1376 305
rect 1288 68 1376 81
<< pdiff >>
rect -264 3151 -176 3164
rect -264 2677 -251 3151
rect -205 2677 -176 3151
rect -264 2664 -176 2677
rect -120 3151 -32 3164
rect -120 2677 -91 3151
rect -45 2677 -32 3151
rect -120 2664 -32 2677
rect 24 3151 112 3164
rect 24 2677 37 3151
rect 83 2677 112 3151
rect 24 2664 112 2677
rect 168 3151 272 3164
rect 168 2677 197 3151
rect 243 2677 272 3151
rect 168 2664 272 2677
rect 328 3151 432 3164
rect 328 2677 357 3151
rect 403 2677 432 3151
rect 328 2664 432 2677
rect 488 3151 592 3164
rect 488 2677 517 3151
rect 563 2677 592 3151
rect 488 2664 592 2677
rect 648 3151 752 3164
rect 648 2677 677 3151
rect 723 2677 752 3151
rect 648 2664 752 2677
rect 808 3151 912 3164
rect 808 2677 837 3151
rect 883 2677 912 3151
rect 808 2664 912 2677
rect 968 3151 1072 3164
rect 968 2677 997 3151
rect 1043 2677 1072 3151
rect 968 2664 1072 2677
rect 1128 3151 1232 3164
rect 1128 2677 1157 3151
rect 1203 2677 1232 3151
rect 1128 2664 1232 2677
rect 1288 3151 1376 3164
rect 1288 2677 1317 3151
rect 1363 2677 1376 3151
rect 1288 2664 1376 2677
rect -264 2515 -176 2528
rect -264 2041 -251 2515
rect -205 2041 -176 2515
rect -264 2028 -176 2041
rect -120 2515 -32 2528
rect -120 2041 -91 2515
rect -45 2041 -32 2515
rect -120 2028 -32 2041
rect 24 2515 112 2528
rect 24 2041 37 2515
rect 83 2041 112 2515
rect 24 2028 112 2041
rect 168 2515 272 2528
rect 168 2041 197 2515
rect 243 2041 272 2515
rect 168 2028 272 2041
rect 328 2515 432 2528
rect 328 2041 357 2515
rect 403 2041 432 2515
rect 328 2028 432 2041
rect 488 2515 592 2528
rect 488 2041 517 2515
rect 563 2041 592 2515
rect 488 2028 592 2041
rect 648 2515 752 2528
rect 648 2041 677 2515
rect 723 2041 752 2515
rect 648 2028 752 2041
rect 808 2515 912 2528
rect 808 2041 837 2515
rect 883 2041 912 2515
rect 808 2028 912 2041
rect 968 2515 1072 2528
rect 968 2041 997 2515
rect 1043 2041 1072 2515
rect 968 2028 1072 2041
rect 1128 2515 1232 2528
rect 1128 2041 1157 2515
rect 1203 2041 1232 2515
rect 1128 2028 1232 2041
rect 1288 2515 1376 2528
rect 1288 2041 1317 2515
rect 1363 2041 1376 2515
rect 1288 2028 1376 2041
rect -264 1879 -176 1892
rect -264 1405 -251 1879
rect -205 1405 -176 1879
rect -264 1392 -176 1405
rect -120 1879 -32 1892
rect -120 1405 -91 1879
rect -45 1405 -32 1879
rect -120 1392 -32 1405
rect 24 1879 112 1892
rect 24 1405 37 1879
rect 83 1405 112 1879
rect 24 1392 112 1405
rect 168 1879 272 1892
rect 168 1405 197 1879
rect 243 1405 272 1879
rect 168 1392 272 1405
rect 328 1879 432 1892
rect 328 1405 357 1879
rect 403 1405 432 1879
rect 328 1392 432 1405
rect 488 1879 592 1892
rect 488 1405 517 1879
rect 563 1405 592 1879
rect 488 1392 592 1405
rect 648 1879 752 1892
rect 648 1405 677 1879
rect 723 1405 752 1879
rect 648 1392 752 1405
rect 808 1879 912 1892
rect 808 1405 837 1879
rect 883 1405 912 1879
rect 808 1392 912 1405
rect 968 1879 1072 1892
rect 968 1405 997 1879
rect 1043 1405 1072 1879
rect 968 1392 1072 1405
rect 1128 1879 1232 1892
rect 1128 1405 1157 1879
rect 1203 1405 1232 1879
rect 1128 1392 1232 1405
rect 1288 1879 1376 1892
rect 1288 1405 1317 1879
rect 1363 1405 1376 1879
rect 1288 1392 1376 1405
<< ndiffc >>
rect -251 853 -205 1077
rect -91 853 -45 1077
rect 37 853 83 1077
rect 197 853 243 1077
rect 357 853 403 1077
rect 517 853 563 1077
rect 677 853 723 1077
rect 837 853 883 1077
rect 997 853 1043 1077
rect 1157 853 1203 1077
rect 1317 853 1363 1077
rect -251 467 -205 691
rect -91 467 -45 691
rect 37 467 83 691
rect 197 467 243 691
rect 357 467 403 691
rect 517 467 563 691
rect 677 467 723 691
rect 837 467 883 691
rect 997 467 1043 691
rect 1157 467 1203 691
rect 1317 467 1363 691
rect -251 81 -205 305
rect -91 81 -45 305
rect 37 81 83 305
rect 197 81 243 305
rect 357 81 403 305
rect 517 81 563 305
rect 677 81 723 305
rect 837 81 883 305
rect 997 81 1043 305
rect 1157 81 1203 305
rect 1317 81 1363 305
<< pdiffc >>
rect -251 2677 -205 3151
rect -91 2677 -45 3151
rect 37 2677 83 3151
rect 197 2677 243 3151
rect 357 2677 403 3151
rect 517 2677 563 3151
rect 677 2677 723 3151
rect 837 2677 883 3151
rect 997 2677 1043 3151
rect 1157 2677 1203 3151
rect 1317 2677 1363 3151
rect -251 2041 -205 2515
rect -91 2041 -45 2515
rect 37 2041 83 2515
rect 197 2041 243 2515
rect 357 2041 403 2515
rect 517 2041 563 2515
rect 677 2041 723 2515
rect 837 2041 883 2515
rect 997 2041 1043 2515
rect 1157 2041 1203 2515
rect 1317 2041 1363 2515
rect -251 1405 -205 1879
rect -91 1405 -45 1879
rect 37 1405 83 1879
rect 197 1405 243 1879
rect 357 1405 403 1879
rect 517 1405 563 1879
rect 677 1405 723 1879
rect 837 1405 883 1879
rect 997 1405 1043 1879
rect 1157 1405 1203 1879
rect 1317 1405 1363 1879
<< psubdiff >>
rect -279 -193 1391 -180
rect -279 -239 -266 -193
rect -220 -239 -172 -193
rect -126 -239 -78 -193
rect -32 -239 16 -193
rect 62 -239 110 -193
rect 156 -239 204 -193
rect 250 -239 298 -193
rect 344 -239 392 -193
rect 438 -239 486 -193
rect 532 -239 580 -193
rect 626 -239 674 -193
rect 720 -239 768 -193
rect 814 -239 862 -193
rect 908 -239 956 -193
rect 1002 -239 1050 -193
rect 1096 -239 1144 -193
rect 1190 -239 1238 -193
rect 1284 -239 1332 -193
rect 1378 -239 1391 -193
rect -279 -252 1391 -239
<< nsubdiff >>
rect -326 3471 1438 3484
rect -326 3425 -313 3471
rect -267 3425 -219 3471
rect -173 3425 -125 3471
rect -79 3425 -31 3471
rect 15 3425 63 3471
rect 109 3425 157 3471
rect 203 3425 251 3471
rect 297 3425 345 3471
rect 391 3425 439 3471
rect 485 3425 533 3471
rect 579 3425 627 3471
rect 673 3425 721 3471
rect 767 3425 815 3471
rect 861 3425 909 3471
rect 955 3425 1003 3471
rect 1049 3425 1097 3471
rect 1143 3425 1191 3471
rect 1237 3425 1285 3471
rect 1331 3425 1379 3471
rect 1425 3425 1438 3471
rect -326 3412 1438 3425
<< psubdiffcont >>
rect -266 -239 -220 -193
rect -172 -239 -126 -193
rect -78 -239 -32 -193
rect 16 -239 62 -193
rect 110 -239 156 -193
rect 204 -239 250 -193
rect 298 -239 344 -193
rect 392 -239 438 -193
rect 486 -239 532 -193
rect 580 -239 626 -193
rect 674 -239 720 -193
rect 768 -239 814 -193
rect 862 -239 908 -193
rect 956 -239 1002 -193
rect 1050 -239 1096 -193
rect 1144 -239 1190 -193
rect 1238 -239 1284 -193
rect 1332 -239 1378 -193
<< nsubdiffcont >>
rect -313 3425 -267 3471
rect -219 3425 -173 3471
rect -125 3425 -79 3471
rect -31 3425 15 3471
rect 63 3425 109 3471
rect 157 3425 203 3471
rect 251 3425 297 3471
rect 345 3425 391 3471
rect 439 3425 485 3471
rect 533 3425 579 3471
rect 627 3425 673 3471
rect 721 3425 767 3471
rect 815 3425 861 3471
rect 909 3425 955 3471
rect 1003 3425 1049 3471
rect 1097 3425 1143 3471
rect 1191 3425 1237 3471
rect 1285 3425 1331 3471
rect 1379 3425 1425 3471
<< polysilicon >>
rect -176 3164 -120 3208
rect 112 3184 1288 3240
rect 112 3164 168 3184
rect 272 3164 328 3184
rect 432 3164 488 3184
rect 592 3164 648 3184
rect 752 3164 808 3184
rect 912 3164 968 3184
rect 1072 3164 1128 3184
rect 1232 3164 1288 3184
rect -176 2528 -120 2664
rect 112 2528 168 2664
rect 272 2528 328 2664
rect 432 2528 488 2664
rect 592 2528 648 2664
rect 752 2528 808 2664
rect 912 2528 968 2664
rect 1072 2528 1128 2664
rect 1232 2528 1288 2664
rect -176 1892 -120 2028
rect 112 1892 168 2028
rect 272 1892 328 2028
rect 432 1892 488 2028
rect 592 1892 648 2028
rect 752 1892 808 2028
rect 912 1892 968 2028
rect 1072 1892 1128 2028
rect 1232 1892 1288 2028
rect -329 1260 -257 1268
rect -176 1260 -120 1392
rect -329 1255 -120 1260
rect -329 1209 -316 1255
rect -270 1209 -120 1255
rect -329 1204 -120 1209
rect -72 1270 0 1278
rect 112 1270 168 1392
rect 272 1348 328 1392
rect 432 1348 488 1392
rect 592 1348 648 1392
rect 752 1348 808 1392
rect 912 1348 968 1392
rect 1072 1348 1128 1392
rect 1232 1348 1288 1392
rect -72 1265 168 1270
rect -72 1219 -59 1265
rect -13 1219 168 1265
rect -72 1214 168 1219
rect -72 1206 0 1214
rect -329 1196 -257 1204
rect -176 1090 -120 1204
rect 112 1090 168 1134
rect 272 1090 328 1134
rect 432 1090 488 1134
rect 592 1090 648 1134
rect 752 1090 808 1134
rect 912 1090 968 1134
rect 1072 1090 1128 1134
rect 1232 1090 1288 1134
rect -176 704 -120 840
rect 112 704 168 840
rect 272 704 328 840
rect 432 704 488 840
rect 592 704 648 840
rect 752 704 808 840
rect 912 704 968 840
rect 1072 704 1128 840
rect 1232 704 1288 840
rect -176 318 -120 454
rect 112 318 168 454
rect 272 318 328 454
rect 432 318 488 454
rect 592 318 648 454
rect 752 318 808 454
rect 912 318 968 454
rect 1072 318 1128 454
rect 1232 318 1288 454
rect -176 48 -120 68
rect 112 48 168 68
rect 272 48 328 68
rect 432 48 488 68
rect 592 48 648 68
rect 752 48 808 68
rect 912 48 968 68
rect 1072 48 1128 68
rect 1232 48 1288 68
rect -176 -8 1288 48
<< polycontact >>
rect -316 1209 -270 1255
rect -59 1219 -13 1265
<< metal1 >>
rect -350 3471 1462 3504
rect -350 3425 -313 3471
rect -267 3425 -219 3471
rect -173 3425 -125 3471
rect -79 3425 -31 3471
rect 15 3425 63 3471
rect 109 3425 157 3471
rect 203 3425 251 3471
rect 297 3425 345 3471
rect 391 3425 439 3471
rect 485 3425 533 3471
rect 579 3425 627 3471
rect 673 3425 721 3471
rect 767 3425 815 3471
rect 861 3425 909 3471
rect 955 3425 1003 3471
rect 1049 3425 1097 3471
rect 1143 3425 1191 3471
rect 1237 3425 1285 3471
rect 1331 3425 1379 3471
rect 1425 3425 1462 3471
rect -350 3392 1462 3425
rect -251 3151 -205 3392
rect 37 3300 1043 3346
rect -251 2515 -205 2677
rect -251 1879 -205 2041
rect -251 1394 -205 1405
rect -91 3151 -45 3162
rect -91 2515 -45 2677
rect -91 1879 -45 2041
rect -91 1276 -45 1405
rect 37 3151 83 3300
rect 997 3254 1043 3300
rect 37 2515 83 2677
rect 37 1879 83 2041
rect 37 1348 83 1405
rect 197 3208 883 3254
rect 197 3151 243 3208
rect 197 2515 243 2677
rect 197 1879 243 2041
rect 197 1394 243 1405
rect 357 3151 403 3162
rect 357 2515 403 2677
rect 357 1879 403 2041
rect 357 1348 403 1405
rect 517 3151 563 3208
rect 517 2515 563 2677
rect 517 1879 563 2041
rect 517 1394 563 1405
rect 677 3151 723 3162
rect 677 2515 723 2677
rect 677 1879 723 2041
rect 677 1348 723 1405
rect 37 1302 723 1348
rect -327 1255 -259 1266
rect -372 1209 -316 1255
rect -270 1209 -259 1255
rect -327 1198 -259 1209
rect -91 1265 -2 1276
rect -91 1219 -59 1265
rect -13 1219 -2 1265
rect -91 1208 -2 1219
rect -251 1077 -205 1088
rect -251 691 -205 853
rect -251 305 -205 467
rect -251 -160 -205 81
rect -91 1077 -45 1208
rect 677 1180 723 1302
rect -91 691 -45 853
rect -91 305 -45 467
rect -91 70 -45 81
rect 37 1134 723 1180
rect 37 1077 83 1134
rect 37 691 83 853
rect 37 305 83 467
rect 37 -68 83 81
rect 197 1077 243 1088
rect 197 691 243 853
rect 197 305 243 467
rect 197 24 243 81
rect 357 1077 403 1134
rect 357 691 403 853
rect 357 305 403 467
rect 357 70 403 81
rect 517 1077 563 1088
rect 517 691 563 853
rect 517 305 563 467
rect 517 24 563 81
rect 677 1077 723 1134
rect 677 691 723 853
rect 677 305 723 467
rect 677 70 723 81
rect 837 3151 883 3208
rect 837 2515 883 2677
rect 837 1879 883 2041
rect 837 1180 883 1405
rect 997 3208 1363 3254
rect 997 3151 1043 3208
rect 997 2515 1043 2677
rect 997 1879 1043 2041
rect 997 1394 1043 1405
rect 1157 3151 1203 3162
rect 1157 2515 1203 2677
rect 1157 1879 1203 2041
rect 1157 1181 1203 1405
rect 1317 3151 1363 3208
rect 1317 2515 1363 2677
rect 1317 1879 1363 2041
rect 1317 1338 1363 1405
rect 1317 1292 1631 1338
rect 1157 1180 1637 1181
rect 837 1135 1637 1180
rect 837 1134 1203 1135
rect 837 1077 883 1134
rect 837 691 883 853
rect 837 305 883 467
rect 837 24 883 81
rect 197 -22 883 24
rect 997 1077 1043 1088
rect 997 691 1043 853
rect 997 305 1043 467
rect 997 24 1043 81
rect 1157 1077 1203 1134
rect 1157 691 1203 853
rect 1157 305 1203 467
rect 1157 70 1203 81
rect 1317 1077 1363 1088
rect 1317 691 1363 853
rect 1317 305 1363 467
rect 1317 24 1363 81
rect 997 -22 1363 24
rect 997 -68 1043 -22
rect 37 -114 1043 -68
rect -288 -193 1400 -160
rect -288 -239 -266 -193
rect -220 -239 -172 -193
rect -126 -239 -78 -193
rect -32 -239 16 -193
rect 62 -239 110 -193
rect 156 -239 204 -193
rect 250 -239 298 -193
rect 344 -239 392 -193
rect 438 -239 486 -193
rect 532 -239 580 -193
rect 626 -239 674 -193
rect 720 -239 768 -193
rect 814 -239 862 -193
rect 908 -239 956 -193
rect 1002 -239 1050 -193
rect 1096 -239 1144 -193
rect 1190 -239 1238 -193
rect 1284 -239 1332 -193
rect 1378 -239 1400 -193
rect -288 -272 1400 -239
<< labels >>
flabel metal1 561 -216 561 -216 0 FreeSans 320 0 0 0 VSS
port 1 nsew
flabel nsubdiffcont 462 3448 462 3448 0 FreeSans 320 0 0 0 VDD
port 2 nsew
flabel polycontact -293 1232 -293 1232 0 FreeSans 320 0 0 0 CLK
port 3 nsew
flabel metal1 1575 1316 1575 1316 0 FreeSans 320 0 0 0 VIN
port 4 nsew
flabel metal1 1448 1156 1448 1156 0 FreeSans 320 0 0 0 VOUT
port 5 nsew
<< end >>
