magic
tech gf180mcuC
magscale 1 10
timestamp 1697518002
<< nwell >>
rect -938 -410 938 410
<< pmos >>
rect -764 -280 -664 280
rect -560 -280 -460 280
rect -356 -280 -256 280
rect -152 -280 -52 280
rect 52 -280 152 280
rect 256 -280 356 280
rect 460 -280 560 280
rect 664 -280 764 280
<< pdiff >>
rect -852 267 -764 280
rect -852 -267 -839 267
rect -793 -267 -764 267
rect -852 -280 -764 -267
rect -664 267 -560 280
rect -664 -267 -635 267
rect -589 -267 -560 267
rect -664 -280 -560 -267
rect -460 267 -356 280
rect -460 -267 -431 267
rect -385 -267 -356 267
rect -460 -280 -356 -267
rect -256 267 -152 280
rect -256 -267 -227 267
rect -181 -267 -152 267
rect -256 -280 -152 -267
rect -52 267 52 280
rect -52 -267 -23 267
rect 23 -267 52 267
rect -52 -280 52 -267
rect 152 267 256 280
rect 152 -267 181 267
rect 227 -267 256 267
rect 152 -280 256 -267
rect 356 267 460 280
rect 356 -267 385 267
rect 431 -267 460 267
rect 356 -280 460 -267
rect 560 267 664 280
rect 560 -267 589 267
rect 635 -267 664 267
rect 560 -280 664 -267
rect 764 267 852 280
rect 764 -267 793 267
rect 839 -267 852 267
rect 764 -280 852 -267
<< pdiffc >>
rect -839 -267 -793 267
rect -635 -267 -589 267
rect -431 -267 -385 267
rect -227 -267 -181 267
rect -23 -267 23 267
rect 181 -267 227 267
rect 385 -267 431 267
rect 589 -267 635 267
rect 793 -267 839 267
<< polysilicon >>
rect -764 280 -664 324
rect -560 280 -460 324
rect -356 280 -256 324
rect -152 280 -52 324
rect 52 280 152 324
rect 256 280 356 324
rect 460 280 560 324
rect 664 280 764 324
rect -764 -324 -664 -280
rect -560 -324 -460 -280
rect -356 -324 -256 -280
rect -152 -324 -52 -280
rect 52 -324 152 -280
rect 256 -324 356 -280
rect 460 -324 560 -280
rect 664 -324 764 -280
<< metal1 >>
rect -839 267 -793 278
rect -839 -278 -793 -267
rect -635 267 -589 278
rect -635 -278 -589 -267
rect -431 267 -385 278
rect -431 -278 -385 -267
rect -227 267 -181 278
rect -227 -278 -181 -267
rect -23 267 23 278
rect -23 -278 23 -267
rect 181 267 227 278
rect 181 -278 227 -267
rect 385 267 431 278
rect 385 -278 431 -267
rect 589 267 635 278
rect 589 -278 635 -267
rect 793 267 839 278
rect 793 -278 839 -267
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 2.8 l 0.5 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
