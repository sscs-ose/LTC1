** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/DAC_12bit_TB_V2.sch
**.subckt DAC_12bit_TB_V2
V1 VSS GND 0
.save i(v1)
V2 VDD VSS 3.3
.save i(v2)
V6 net1 VSS pulse(0 3.3 0 10p 10p 20n 40n)
.save i(v6)
V7 net2 VSS pulse(0 3.3 0 10p 10p 40n 80n)
.save i(v7)
V8 net3 VSS pulse(0 3.3 0 10p 10p 80n 160n)
.save i(v8)
V10 net4 VSS pulse(0 3.3 0 10p 10p 10n 20n)
.save i(v10)
V11 net5 VSS pulse(0 3.3 0 10p 10p 5n 10n)
.save i(v11)
V12 net6 VSS pulse(0 3.3 0 10p 10p 2.5n 5n)
.save i(v12)
I0 VDD I1 20u
V3 net7 VSS pulse(0 3.3 0 10p 10p 1280n 2560n)
.save i(v3)
V4 net8 VSS pulse(0 3.3 0 10p 10p 2560n 5120n)
.save i(v4)
V5 net9 VSS pulse(0 3.3 0 10p 10p 5120n 10240n)
.save i(v5)
V9 net10 VSS pulse(0 3.3 0 10p 10p 640n 1280n)
.save i(v9)
V13 net11 VSS pulse(0 3.3 0 10p 10p 320n 640n)
.save i(v13)
V14 net12 VSS pulse(0 3.3 0 10p 10p 160n 320n)
.save i(v14)
I1 VDD I2 20u
R1 Out+ VDD 25 m=1
R2 Out- VDD 25 m=1
x1 net2 net10 VDD I2 net8 net6 net12 Out+ net4 net9 net7 net1 net11 Out- I1 net3 net5 VSS
+ DAC_12Bit_V2
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.options savecurrents
.control
save all
op

tran 1000p 10240n
plot v(Out-) v(Out+)

write DAC_12bit_TB_V2.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  DAC_12Bit_V2.sym # of pins=18
** sym_path: /home/shahid/GF180Projects/GF_INV/Xschem/DAC_12Bit_V2.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/DAC_12Bit_V2.sch
.subckt DAC_12Bit_V2 B5 B9 VDD I1 B11 B1 B7 Iout- B3 B12 B10 B4 B8 Iout+ I2 B6 B2 VSS
*.iopin VDD
*.iopin VSS
*.ipin B1
*.ipin B2
*.ipin B3
*.ipin B4
*.ipin B5
*.ipin B6
*.ipin B7
*.ipin B8
*.ipin B9
*.ipin B10
*.ipin B11
*.ipin B12
*.ipin I1
*.ipin I2
*.opin Iout-
*.opin Iout+
x1 VDD VSS B1 B2 B3 B4 B5 B6 VDD I1 Iout+ Iout- LSB
x3 VSS VDD B11 B7 B8 B12 B9 I2 B10 Iout- Iout+ MSB_6Bit
.ends


* expanding   symbol:  LSB.sym # of pins=12
** sym_path: /home/shahid/GF180Projects/GF_INV/Xschem/LSB.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/LSB.sch
.subckt LSB VDD VSS B1 B2 B3 B4 B5 B6 CLK ITAIL IOUT+ IOUT-
*.iopin VDD
*.iopin VSS
*.ipin B1
*.ipin B2
*.ipin B3
*.ipin B4
*.ipin B5
*.ipin B6
*.ipin CLK
*.ipin ITAIL
*.opin IOUT+
*.opin IOUT-
x1 VDD VSS B1 b1b b1 Balanced_Inverter
x2 VDD VSS B2 b2b b2 Balanced_Inverter
x3 VDD VSS B3 b3b b3 Balanced_Inverter
x4 VDD VSS B4 b4b b4 Balanced_Inverter
x5 VDD VSS B5 b5b b5 Balanced_Inverter
x6 VDD VSS B6 b6b b6 Balanced_Inverter
x7 VDD VSS CLK clkb clk Balanced_Inverter
XM21 IOUT+ net15 IOUT+ VSS nfet_03v3 L=0.28u W=0.25u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
x9 VDD VSS b5 b5b clk clkb net4 net3 CMLL
x10 VDD VSS b4 b4b clk clkb net6 net5 CMLL
x11 VDD VSS b3 b3b clk clkb net10 net9 CMLL
x12 VDD VSS b2 b2b clk clkb net12 net11 CMLL
x13 VDD VSS b1 b1b clk clkb net14 net15 CMLL
x14 VDD VSS b6 b6b clk clkb net1 net2 CMLL
XM23 IOUT- net14 IOUT- VSS nfet_03v3 L=0.28u W=0.25u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
x8 net13 IOUT- VSS net15 nfet_03V3_m2
x15 net13 IOUT+ VSS net14 nfet_03V3_m2
x16 net16 ITAIL VSS ITAIL nfet_03V3_m2
x17 VSS net16 VSS net16 nfet_03V3_m2
x18 net20 net13 VSS ITAIL nfet_03V3_m2
x19 VSS net20 VSS net16 nfet_03V3_m2
x20 IOUT+ IOUT+ VSS net11 nfet_03V3_m2
x21 IOUT- IOUT- VSS net12 nfet_03V3_m2
x22 net17 IOUT+ VSS net12 nfet_03V3_m4
x23 net17 IOUT- VSS net11 nfet_03V3_m4
x24 IOUT+ IOUT+ VSS net9 nfet_03V3_m4
x25 IOUT- IOUT- VSS net10 nfet_03V3_m4
x26 net21 net17 VSS ITAIL nfet_03V3_m4
x27 VSS net21 VSS net16 nfet_03V3_m4
x28 net22 net8 VSS ITAIL nfet_03V3_m8
x29 VSS net22 VSS net16 nfet_03V3_m8
x30 net8 IOUT- VSS net9 nfet_03V3_m8
x31 net8 IOUT+ VSS net10 nfet_03V3_m8
x32 IOUT- IOUT- VSS net6 nfet_03V3_m8
x33 IOUT+ IOUT+ VSS net5 nfet_03V3_m8
x34 net7 IOUT- VSS net5 nfet_03V3_m16
x35 net7 IOUT+ VSS net6 nfet_03V3_m16
x36 IOUT- IOUT- VSS net4 nfet_03V3_m16
x37 IOUT+ IOUT+ VSS net3 nfet_03V3_m16
x38 net23 net7 VSS ITAIL nfet_03V3_m16
x39 VSS net23 VSS net16 nfet_03V3_m16
x40 net24 net18 VSS ITAIL nfet_03V3_m32
x41 VSS net24 VSS net16 nfet_03V3_m32
x42 net18 IOUT- VSS net3 nfet_03V3_m32
x43 net18 IOUT+ VSS net4 nfet_03V3_m32
x44 IOUT- IOUT- VSS net1 nfet_03V3_m32
x45 IOUT+ IOUT+ VSS net2 nfet_03V3_m32
x46 net25 net19 VSS ITAIL nfet_03V3_m64
x47 VSS net25 VSS net16 nfet_03V3_m64
x48 net19 IOUT- VSS net2 nfet_03V3_m64
x49 net19 IOUT+ VSS net1 nfet_03V3_m64
.ends


* expanding   symbol:  MSB_6Bit.sym # of pins=11
** sym_path: /home/shahid/GF180Projects/GF_INV/Xschem/MSB_6Bit.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/MSB_6Bit.sch
.subckt MSB_6Bit VSS VDD B11 B7 B8 B12 B9 IM_T B10 IOUT- IOUT+
*.iopin VDD
*.iopin VSS
*.ipin B7
*.ipin B11
*.ipin B8
*.ipin B12
*.ipin B9
*.ipin IM_T
*.ipin B10
*.opin IOUT+
*.opin IOUT-
x57 IOUT+ IOUT- VDD VDD R0 C0 IM_T IM VSS MSB_UNIT_CELL
x58 IOUT+ IOUT- VDD VDD R0 C1 IM_T IM VSS MSB_UNIT_CELL
x59 IOUT+ IOUT- VDD VDD R0 C2 IM_T IM VSS MSB_UNIT_CELL
x60 IOUT+ IOUT- VDD VDD R0 C3 IM_T IM VSS MSB_UNIT_CELL
x61 IOUT+ IOUT- VDD VDD R0 C4 IM_T IM VSS MSB_UNIT_CELL
x62 IOUT+ IOUT- VDD VDD R0 C5 IM_T IM VSS MSB_UNIT_CELL
x63 IOUT+ IOUT- VDD VDD R0 C6 IM_T IM VSS MSB_UNIT_CELL
x64 IOUT+ IOUT- VDD VDD R0 VSS IM_T IM VSS MSB_UNIT_CELL
x1 IOUT+ IOUT- VDD R0 R1 C0 IM_T IM VSS MSB_UNIT_CELL
x2 IOUT+ IOUT- VDD R0 R1 C1 IM_T IM VSS MSB_UNIT_CELL
x3 IOUT+ IOUT- VDD R0 R1 C2 IM_T IM VSS MSB_UNIT_CELL
x4 IOUT+ IOUT- VDD R0 R1 C3 IM_T IM VSS MSB_UNIT_CELL
x5 IOUT+ IOUT- VDD R0 R1 C4 IM_T IM VSS MSB_UNIT_CELL
x6 IOUT+ IOUT- VDD R0 R1 C5 IM_T IM VSS MSB_UNIT_CELL
x7 IOUT+ IOUT- VDD R0 R1 C6 IM_T IM VSS MSB_UNIT_CELL
x8 IOUT+ IOUT- VDD R0 R1 VSS IM_T IM VSS MSB_UNIT_CELL
x9 IOUT+ IOUT- VDD R1 R2 C0 IM_T IM VSS MSB_UNIT_CELL
x10 IOUT+ IOUT- VDD R1 R2 C1 IM_T IM VSS MSB_UNIT_CELL
x11 IOUT+ IOUT- VDD R1 R2 C2 IM_T IM VSS MSB_UNIT_CELL
x12 IOUT+ IOUT- VDD R1 R2 C3 IM_T IM VSS MSB_UNIT_CELL
x13 IOUT+ IOUT- VDD R1 R2 C4 IM_T IM VSS MSB_UNIT_CELL
x14 IOUT+ IOUT- VDD R1 R2 C5 IM_T IM VSS MSB_UNIT_CELL
x15 IOUT+ IOUT- VDD R1 R2 C6 IM_T IM VSS MSB_UNIT_CELL
x16 IOUT+ IOUT- VDD R1 R2 R2 IM_T IM VSS MSB_UNIT_CELL
x17 IOUT+ IOUT- VDD R2 R3 C0 IM_T IM VSS MSB_UNIT_CELL
x18 IOUT+ IOUT- VDD R2 R3 C1 IM_T IM VSS MSB_UNIT_CELL
x19 IOUT+ IOUT- VDD R2 R3 C2 IM_T IM VSS MSB_UNIT_CELL
x20 IOUT+ IOUT- VDD R2 R3 C3 IM_T IM VSS MSB_UNIT_CELL
x21 IOUT+ IOUT- VDD R2 R3 C4 IM_T IM VSS MSB_UNIT_CELL
x22 IOUT+ IOUT- VDD R2 R3 C5 IM_T IM VSS MSB_UNIT_CELL
x23 IOUT+ IOUT- VDD R2 R3 C6 IM_T IM VSS MSB_UNIT_CELL
x24 IOUT+ IOUT- VDD R2 R3 VSS IM_T IM VSS MSB_UNIT_CELL
x25 IOUT+ IOUT- VDD R3 R4 C0 IM_T IM VSS MSB_UNIT_CELL
x26 IOUT+ IOUT- VDD R3 R4 C1 IM_T IM VSS MSB_UNIT_CELL
x27 IOUT+ IOUT- VDD R3 R4 C2 IM_T IM VSS MSB_UNIT_CELL
x28 IOUT+ IOUT- VDD R3 R4 C3 IM_T IM VSS MSB_UNIT_CELL
x29 IOUT+ IOUT- VDD R3 R4 C4 IM_T IM VSS MSB_UNIT_CELL
x30 IOUT+ IOUT- VDD R3 R4 C5 IM_T IM VSS MSB_UNIT_CELL
x31 IOUT+ IOUT- VDD R3 R4 C6 IM_T IM VSS MSB_UNIT_CELL
x32 IOUT+ IOUT- VDD R3 R4 VSS IM_T IM VSS MSB_UNIT_CELL
x33 IOUT+ IOUT- VDD R4 R5 C0 IM_T IM VSS MSB_UNIT_CELL
x34 IOUT+ IOUT- VDD R4 R5 C1 IM_T IM VSS MSB_UNIT_CELL
x35 IOUT+ IOUT- VDD R4 R5 C2 IM_T IM VSS MSB_UNIT_CELL
x36 IOUT+ IOUT- VDD R4 R5 C3 IM_T IM VSS MSB_UNIT_CELL
x37 IOUT+ IOUT- VDD R4 R5 C4 IM_T IM VSS MSB_UNIT_CELL
x38 IOUT+ IOUT- VDD R4 R5 C5 IM_T IM VSS MSB_UNIT_CELL
x39 IOUT+ IOUT- VDD R4 R5 C6 IM_T IM VSS MSB_UNIT_CELL
x40 IOUT+ IOUT- VDD R4 R5 VSS IM_T IM VSS MSB_UNIT_CELL
x41 IOUT+ IOUT- VDD R5 R6 C0 IM_T IM VSS MSB_UNIT_CELL
x42 IOUT+ IOUT- VDD R5 R6 C1 IM_T IM VSS MSB_UNIT_CELL
x43 IOUT+ IOUT- VDD R5 R6 C2 IM_T IM VSS MSB_UNIT_CELL
x44 IOUT+ IOUT- VDD R5 R6 C3 IM_T IM VSS MSB_UNIT_CELL
x45 IOUT+ IOUT- VDD R5 R6 C4 IM_T IM VSS MSB_UNIT_CELL
x46 IOUT+ IOUT- VDD R5 R6 C5 IM_T IM VSS MSB_UNIT_CELL
x47 IOUT+ IOUT- VDD R5 R6 C6 IM_T IM VSS MSB_UNIT_CELL
x48 IOUT+ IOUT- VDD R5 R6 VSS IM_T IM VSS MSB_UNIT_CELL
x49 IOUT+ IOUT- VDD R6 VSS C0 IM_T IM VSS MSB_UNIT_CELL
x50 IOUT+ IOUT- VDD R6 VSS C1 IM_T IM VSS MSB_UNIT_CELL
x51 IOUT+ IOUT- VDD R6 VSS C2 IM_T IM VSS MSB_UNIT_CELL
x52 IOUT+ IOUT- VDD R6 VSS C3 IM_T IM VSS MSB_UNIT_CELL
x53 IOUT+ IOUT- VDD R6 VSS C4 IM_T IM VSS MSB_UNIT_CELL
x54 IOUT+ IOUT- VDD R6 VSS C5 IM_T IM VSS MSB_UNIT_CELL
x55 IOUT+ IOUT- VDD R6 VSS C6 IM_T IM VSS MSB_UNIT_CELL
x56 C6 VDD C5 VSS C4 B9 C3 C2 B8 C1 B7 C0 Thermo_Decoder
x65 R6 VDD R5 VSS R4 B12 R3 R2 B11 R1 B10 R0 Thermo_Decoder
XM1 IM_T IM_T IM VSS nfet_03v3 L=0.28u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 IM IM VSS VSS nfet_03v3 L=0.28u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  Balanced_Inverter.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/GF_INV/Xschem/Balanced_Inverter.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/Balanced_Inverter.sch
.subckt Balanced_Inverter VDD VSS VIN OUT_B OUT
*.iopin VSS
*.ipin VIN
*.opin OUT_B
*.iopin VDD
*.opin OUT
XM1 OUT_B VIN VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT_B OUT VDD VDD pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 OUT net1 VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 OUT OUT_B VDD VDD pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
x1 VSS VDD net1 VIN GF_INV
.ends


* expanding   symbol:  CMLL.sym # of pins=8
** sym_path: /home/shahid/GF180Projects/GF_INV/Xschem/CMLL.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/CMLL.sch
.subckt CMLL VDD VSS D D_B CLK CLKB Q Q_B
*.iopin VDD
*.iopin VSS
*.ipin D
*.ipin D_B
*.ipin CLK
*.ipin CLKB
*.opin Q
*.opin Q_B
XM2 Q D_B net1 VSS nfet_03v3 L=0.28u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 Q Q_B net2 VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 Q_B Q net2 VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 net2 CLKB net3 VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM6 Q_B D net1 VSS nfet_03v3 L=0.28u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
R1 VDD Q_B 20k m=1
R2 VDD Q 20k m=1
I0 net3 VSS 50u
XM1 net1 CLK net3 VSS nfet_03v3 L=0.28u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  nfet_03V3_m2.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/GF_INV/Xschem/nfet_03V3_m2.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/nfet_03V3_m2.sch
.subckt nfet_03V3_m2 S D B G
*.iopin G
*.iopin S
*.iopin D
*.iopin B
XM1 D G S B nfet_03v3 L=0.28u W=0.25u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 D G S B nfet_03v3 L=0.28u W=0.25u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  nfet_03V3_m4.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/GF_INV/Xschem/nfet_03V3_m4.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/nfet_03V3_m4.sch
.subckt nfet_03V3_m4 S D B G
*.iopin G
*.iopin S
*.iopin D
*.iopin B
x1 S D B G nfet_03V3_m2
x2 S D B G nfet_03V3_m2
.ends


* expanding   symbol:  nfet_03V3_m8.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/GF_INV/Xschem/nfet_03V3_m8.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/nfet_03V3_m8.sch
.subckt nfet_03V3_m8 S D B G
*.iopin G
*.iopin S
*.iopin D
*.iopin B
x1 S D B G nfet_03V3_m4
x2 S D B G nfet_03V3_m4
.ends


* expanding   symbol:  nfet_03V3_m16.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/GF_INV/Xschem/nfet_03V3_m16.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/nfet_03V3_m16.sch
.subckt nfet_03V3_m16 S D B G
*.iopin G
*.iopin S
*.iopin D
*.iopin B
x1 S D B G nfet_03V3_m8
x2 S D B G nfet_03V3_m8
.ends


* expanding   symbol:  nfet_03V3_m32.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/GF_INV/Xschem/nfet_03V3_m32.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/nfet_03V3_m32.sch
.subckt nfet_03V3_m32 S D B G
*.iopin G
*.iopin S
*.iopin D
*.iopin B
x1 S D B G nfet_03V3_m16
x2 S D B G nfet_03V3_m16
.ends


* expanding   symbol:  nfet_03V3_m64.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/GF_INV/Xschem/nfet_03V3_m64.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/nfet_03V3_m64.sch
.subckt nfet_03V3_m64 S D B G
*.iopin G
*.iopin S
*.iopin D
*.iopin B
x1 S D B G nfet_03V3_m32
x2 S D B G nfet_03V3_m32
.ends


* expanding   symbol:  MSB_UNIT_CELL.sym # of pins=9
** sym_path: /home/shahid/GF180Projects/GF_INV/Xschem/MSB_UNIT_CELL.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/MSB_UNIT_CELL.sch
.subckt MSB_UNIT_CELL IOUT+ IOUT- VDD Ri-1 Ri Ci IM_T IM VSS
*.iopin VDD
*.iopin VSS
*.ipin Ri-1
*.ipin Ri
*.ipin Ci
*.ipin IM_T
*.ipin IM
*.opin IOUT+
*.opin IOUT-
x1 VDD VSS Ri-1 Ri Ci net2 net3 Local_Enc
XM1 IOUT+ net2 net1 VSS nfet_03v3 L=0.28u W=32u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 IOUT- net3 net1 VSS nfet_03v3 L=0.28u W=32u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 net1 IM_T net4 VSS nfet_03v3 L=0.28u W=32u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 net4 IM VSS VSS nfet_03v3 L=0.28u W=32u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  Thermo_Decoder.sym # of pins=12
** sym_path: /home/shahid/GF180Projects/GF_INV/Xschem/Thermo_Decoder.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/Thermo_Decoder.sch
.subckt Thermo_Decoder D1 VDD D2 VSS D3 B1 D4 D5 B2 D6 B3 D7
*.iopin VDD
*.iopin VSS
*.ipin B1
*.ipin B2
*.ipin B3
*.opin D3
*.opin D4
*.opin D1
*.opin D2
*.opin D6
*.opin D7
*.opin D5
x1 VDD VSS B1 B2 net1 AND
x2 VDD VSS net2 D1 inv
x3 VDD VSS B1 B2 net6 OR
x4 VDD VSS B2 B3 net4 OR
x5 VDD VSS B1 B2 net3 AND
x6 VDD VSS net1 B3 net2 AND
x7 VDD VSS net3 D2 inv
x8 VDD VSS net4 B1 net5 AND
x9 VDD VSS net5 D3 inv
x10 VDD VSS B1 D4 inv
x11 VDD VSS net6 D6 inv
x12 VDD VSS B2 B3 net9 AND
x13 VDD VSS B1 net9 net10 OR
x14 VDD VSS net10 D5 inv
x15 VDD VSS B1 B2 net7 OR
x16 VDD VSS net7 B3 net8 OR
x17 VDD VSS net8 D7 inv
.ends


* expanding   symbol:  GF_INV.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/GF_INV/Xschem/GF_INV.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/GF_INV.sch
.subckt GF_INV VSS VDD OUT IN
*.iopin VDD
*.iopin VSS
*.ipin IN
*.opin OUT
XM1 OUT IN VSS VSS nfet_03v3 L=0.28u W=0.25u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT IN VDD VDD pfet_03v3 L=0.28u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  Local_Enc.sym # of pins=7
** sym_path: /home/shahid/GF180Projects/GF_INV/Xschem/Local_Enc.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/Local_Enc.sch
.subckt Local_Enc VDD VSS Ri-1 Ri Ci Q QB
*.iopin VDD
*.iopin VSS
*.ipin Ri-1
*.ipin Ri
*.ipin Ci
*.opin Q
*.opin QB
x1 VDD VSS Ri-1 Ri-1 net5 NAND
x2 VDD VSS Ri Ri net6 NAND
x3 VDD VSS Ci Ci net7 NAND
x4 VDD VSS net5 net5 net3 NAND
x5 VDD VSS net6 net7 net4 NAND
x6 VDD VSS net3 net4 net2 NAND
x7 VDD VSS net2 net2 net1 NAND
x8 VDD VSS Q net1 QB NAND
x9 VDD VSS net2 QB Q NAND
.ends


* expanding   symbol:  AND.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/GF_INV/Xschem/AND.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/AND.sch
.subckt AND VDD VSS A B OUT
*.iopin VDD
*.iopin VSS
*.ipin A
*.ipin B
*.opin OUT
XM1 net2 B VSS VSS nfet_03v3 L=0.28u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 net1 A VDD VDD pfet_03v3 L=0.28u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 net1 B VDD VDD pfet_03v3 L=0.28u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 net1 A net2 VSS nfet_03v3 L=0.28u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
x1 VSS VDD OUT net1 GF_INV
.ends


* expanding   symbol:  inv.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/GF_INV/Xschem/inv.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/inv.sch
.subckt inv VDD VSS IN OUT
*.opin OUT
*.iopin VDD
*.iopin VSS
*.ipin IN
x1 VSS VDD net1 IN GF_INV
x2 VSS VDD OUT net1 GF_INV
.ends


* expanding   symbol:  OR.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/GF_INV/Xschem/OR.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/OR.sch
.subckt OR VDD VSS A B OUT
*.iopin VDD
*.iopin VSS
*.ipin A
*.ipin B
*.opin OUT
x1 VSS VDD OUT net1 GF_INV
XM1 net1 B VSS VSS nfet_03v3 L=0.28u W=0.25u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 net2 A VDD VDD pfet_03v3 L=0.28u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 net1 B net2 VDD pfet_03v3 L=0.28u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM6 net1 A VSS VSS nfet_03v3 L=0.28u W=0.25u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  NAND.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/GF_INV/Xschem/NAND.sym
** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/NAND.sch
.subckt NAND VDD VSS A B OUT
*.iopin VDD
*.iopin VSS
*.ipin A
*.ipin B
*.opin OUT
XM2 OUT A VDD VDD pfet_03v3 L=0.28u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 OUT B VDD VDD pfet_03v3 L=0.28u W=0.5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
x1 VSS net1 VSS B nfet_03V3_m2
x2 net1 OUT VSS A nfet_03V3_m2
.ends

.GLOBAL GND
.end
