magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1478 -1073 1478 1073
<< metal1 >>
rect -478 67 478 73
rect -478 41 -472 67
rect -446 41 -418 67
rect -392 41 -364 67
rect -338 41 -310 67
rect -284 41 -256 67
rect -230 41 -202 67
rect -176 41 -148 67
rect -122 41 -94 67
rect -68 41 -40 67
rect -14 41 14 67
rect 40 41 68 67
rect 94 41 122 67
rect 148 41 176 67
rect 202 41 230 67
rect 256 41 284 67
rect 310 41 338 67
rect 364 41 392 67
rect 418 41 446 67
rect 472 41 478 67
rect -478 13 478 41
rect -478 -13 -472 13
rect -446 -13 -418 13
rect -392 -13 -364 13
rect -338 -13 -310 13
rect -284 -13 -256 13
rect -230 -13 -202 13
rect -176 -13 -148 13
rect -122 -13 -94 13
rect -68 -13 -40 13
rect -14 -13 14 13
rect 40 -13 68 13
rect 94 -13 122 13
rect 148 -13 176 13
rect 202 -13 230 13
rect 256 -13 284 13
rect 310 -13 338 13
rect 364 -13 392 13
rect 418 -13 446 13
rect 472 -13 478 13
rect -478 -41 478 -13
rect -478 -67 -472 -41
rect -446 -67 -418 -41
rect -392 -67 -364 -41
rect -338 -67 -310 -41
rect -284 -67 -256 -41
rect -230 -67 -202 -41
rect -176 -67 -148 -41
rect -122 -67 -94 -41
rect -68 -67 -40 -41
rect -14 -67 14 -41
rect 40 -67 68 -41
rect 94 -67 122 -41
rect 148 -67 176 -41
rect 202 -67 230 -41
rect 256 -67 284 -41
rect 310 -67 338 -41
rect 364 -67 392 -41
rect 418 -67 446 -41
rect 472 -67 478 -41
rect -478 -73 478 -67
<< via1 >>
rect -472 41 -446 67
rect -418 41 -392 67
rect -364 41 -338 67
rect -310 41 -284 67
rect -256 41 -230 67
rect -202 41 -176 67
rect -148 41 -122 67
rect -94 41 -68 67
rect -40 41 -14 67
rect 14 41 40 67
rect 68 41 94 67
rect 122 41 148 67
rect 176 41 202 67
rect 230 41 256 67
rect 284 41 310 67
rect 338 41 364 67
rect 392 41 418 67
rect 446 41 472 67
rect -472 -13 -446 13
rect -418 -13 -392 13
rect -364 -13 -338 13
rect -310 -13 -284 13
rect -256 -13 -230 13
rect -202 -13 -176 13
rect -148 -13 -122 13
rect -94 -13 -68 13
rect -40 -13 -14 13
rect 14 -13 40 13
rect 68 -13 94 13
rect 122 -13 148 13
rect 176 -13 202 13
rect 230 -13 256 13
rect 284 -13 310 13
rect 338 -13 364 13
rect 392 -13 418 13
rect 446 -13 472 13
rect -472 -67 -446 -41
rect -418 -67 -392 -41
rect -364 -67 -338 -41
rect -310 -67 -284 -41
rect -256 -67 -230 -41
rect -202 -67 -176 -41
rect -148 -67 -122 -41
rect -94 -67 -68 -41
rect -40 -67 -14 -41
rect 14 -67 40 -41
rect 68 -67 94 -41
rect 122 -67 148 -41
rect 176 -67 202 -41
rect 230 -67 256 -41
rect 284 -67 310 -41
rect 338 -67 364 -41
rect 392 -67 418 -41
rect 446 -67 472 -41
<< metal2 >>
rect -478 67 478 73
rect -478 41 -472 67
rect -446 41 -418 67
rect -392 41 -364 67
rect -338 41 -310 67
rect -284 41 -256 67
rect -230 41 -202 67
rect -176 41 -148 67
rect -122 41 -94 67
rect -68 41 -40 67
rect -14 41 14 67
rect 40 41 68 67
rect 94 41 122 67
rect 148 41 176 67
rect 202 41 230 67
rect 256 41 284 67
rect 310 41 338 67
rect 364 41 392 67
rect 418 41 446 67
rect 472 41 478 67
rect -478 13 478 41
rect -478 -13 -472 13
rect -446 -13 -418 13
rect -392 -13 -364 13
rect -338 -13 -310 13
rect -284 -13 -256 13
rect -230 -13 -202 13
rect -176 -13 -148 13
rect -122 -13 -94 13
rect -68 -13 -40 13
rect -14 -13 14 13
rect 40 -13 68 13
rect 94 -13 122 13
rect 148 -13 176 13
rect 202 -13 230 13
rect 256 -13 284 13
rect 310 -13 338 13
rect 364 -13 392 13
rect 418 -13 446 13
rect 472 -13 478 13
rect -478 -41 478 -13
rect -478 -67 -472 -41
rect -446 -67 -418 -41
rect -392 -67 -364 -41
rect -338 -67 -310 -41
rect -284 -67 -256 -41
rect -230 -67 -202 -41
rect -176 -67 -148 -41
rect -122 -67 -94 -41
rect -68 -67 -40 -41
rect -14 -67 14 -41
rect 40 -67 68 -41
rect 94 -67 122 -41
rect 148 -67 176 -41
rect 202 -67 230 -41
rect 256 -67 284 -41
rect 310 -67 338 -41
rect 364 -67 392 -41
rect 418 -67 446 -41
rect 472 -67 478 -41
rect -478 -73 478 -67
<< end >>
