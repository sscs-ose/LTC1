magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1349 -2372 1349 2372
<< metal3 >>
rect -349 1367 349 1372
rect -349 1339 -344 1367
rect -316 1339 -278 1367
rect -250 1339 -212 1367
rect -184 1339 -146 1367
rect -118 1339 -80 1367
rect -52 1339 -14 1367
rect 14 1339 52 1367
rect 80 1339 118 1367
rect 146 1339 184 1367
rect 212 1339 250 1367
rect 278 1339 316 1367
rect 344 1339 349 1367
rect -349 1301 349 1339
rect -349 1273 -344 1301
rect -316 1273 -278 1301
rect -250 1273 -212 1301
rect -184 1273 -146 1301
rect -118 1273 -80 1301
rect -52 1273 -14 1301
rect 14 1273 52 1301
rect 80 1273 118 1301
rect 146 1273 184 1301
rect 212 1273 250 1301
rect 278 1273 316 1301
rect 344 1273 349 1301
rect -349 1235 349 1273
rect -349 1207 -344 1235
rect -316 1207 -278 1235
rect -250 1207 -212 1235
rect -184 1207 -146 1235
rect -118 1207 -80 1235
rect -52 1207 -14 1235
rect 14 1207 52 1235
rect 80 1207 118 1235
rect 146 1207 184 1235
rect 212 1207 250 1235
rect 278 1207 316 1235
rect 344 1207 349 1235
rect -349 1169 349 1207
rect -349 1141 -344 1169
rect -316 1141 -278 1169
rect -250 1141 -212 1169
rect -184 1141 -146 1169
rect -118 1141 -80 1169
rect -52 1141 -14 1169
rect 14 1141 52 1169
rect 80 1141 118 1169
rect 146 1141 184 1169
rect 212 1141 250 1169
rect 278 1141 316 1169
rect 344 1141 349 1169
rect -349 1103 349 1141
rect -349 1075 -344 1103
rect -316 1075 -278 1103
rect -250 1075 -212 1103
rect -184 1075 -146 1103
rect -118 1075 -80 1103
rect -52 1075 -14 1103
rect 14 1075 52 1103
rect 80 1075 118 1103
rect 146 1075 184 1103
rect 212 1075 250 1103
rect 278 1075 316 1103
rect 344 1075 349 1103
rect -349 1037 349 1075
rect -349 1009 -344 1037
rect -316 1009 -278 1037
rect -250 1009 -212 1037
rect -184 1009 -146 1037
rect -118 1009 -80 1037
rect -52 1009 -14 1037
rect 14 1009 52 1037
rect 80 1009 118 1037
rect 146 1009 184 1037
rect 212 1009 250 1037
rect 278 1009 316 1037
rect 344 1009 349 1037
rect -349 971 349 1009
rect -349 943 -344 971
rect -316 943 -278 971
rect -250 943 -212 971
rect -184 943 -146 971
rect -118 943 -80 971
rect -52 943 -14 971
rect 14 943 52 971
rect 80 943 118 971
rect 146 943 184 971
rect 212 943 250 971
rect 278 943 316 971
rect 344 943 349 971
rect -349 905 349 943
rect -349 877 -344 905
rect -316 877 -278 905
rect -250 877 -212 905
rect -184 877 -146 905
rect -118 877 -80 905
rect -52 877 -14 905
rect 14 877 52 905
rect 80 877 118 905
rect 146 877 184 905
rect 212 877 250 905
rect 278 877 316 905
rect 344 877 349 905
rect -349 839 349 877
rect -349 811 -344 839
rect -316 811 -278 839
rect -250 811 -212 839
rect -184 811 -146 839
rect -118 811 -80 839
rect -52 811 -14 839
rect 14 811 52 839
rect 80 811 118 839
rect 146 811 184 839
rect 212 811 250 839
rect 278 811 316 839
rect 344 811 349 839
rect -349 773 349 811
rect -349 745 -344 773
rect -316 745 -278 773
rect -250 745 -212 773
rect -184 745 -146 773
rect -118 745 -80 773
rect -52 745 -14 773
rect 14 745 52 773
rect 80 745 118 773
rect 146 745 184 773
rect 212 745 250 773
rect 278 745 316 773
rect 344 745 349 773
rect -349 707 349 745
rect -349 679 -344 707
rect -316 679 -278 707
rect -250 679 -212 707
rect -184 679 -146 707
rect -118 679 -80 707
rect -52 679 -14 707
rect 14 679 52 707
rect 80 679 118 707
rect 146 679 184 707
rect 212 679 250 707
rect 278 679 316 707
rect 344 679 349 707
rect -349 641 349 679
rect -349 613 -344 641
rect -316 613 -278 641
rect -250 613 -212 641
rect -184 613 -146 641
rect -118 613 -80 641
rect -52 613 -14 641
rect 14 613 52 641
rect 80 613 118 641
rect 146 613 184 641
rect 212 613 250 641
rect 278 613 316 641
rect 344 613 349 641
rect -349 575 349 613
rect -349 547 -344 575
rect -316 547 -278 575
rect -250 547 -212 575
rect -184 547 -146 575
rect -118 547 -80 575
rect -52 547 -14 575
rect 14 547 52 575
rect 80 547 118 575
rect 146 547 184 575
rect 212 547 250 575
rect 278 547 316 575
rect 344 547 349 575
rect -349 509 349 547
rect -349 481 -344 509
rect -316 481 -278 509
rect -250 481 -212 509
rect -184 481 -146 509
rect -118 481 -80 509
rect -52 481 -14 509
rect 14 481 52 509
rect 80 481 118 509
rect 146 481 184 509
rect 212 481 250 509
rect 278 481 316 509
rect 344 481 349 509
rect -349 443 349 481
rect -349 415 -344 443
rect -316 415 -278 443
rect -250 415 -212 443
rect -184 415 -146 443
rect -118 415 -80 443
rect -52 415 -14 443
rect 14 415 52 443
rect 80 415 118 443
rect 146 415 184 443
rect 212 415 250 443
rect 278 415 316 443
rect 344 415 349 443
rect -349 377 349 415
rect -349 349 -344 377
rect -316 349 -278 377
rect -250 349 -212 377
rect -184 349 -146 377
rect -118 349 -80 377
rect -52 349 -14 377
rect 14 349 52 377
rect 80 349 118 377
rect 146 349 184 377
rect 212 349 250 377
rect 278 349 316 377
rect 344 349 349 377
rect -349 311 349 349
rect -349 283 -344 311
rect -316 283 -278 311
rect -250 283 -212 311
rect -184 283 -146 311
rect -118 283 -80 311
rect -52 283 -14 311
rect 14 283 52 311
rect 80 283 118 311
rect 146 283 184 311
rect 212 283 250 311
rect 278 283 316 311
rect 344 283 349 311
rect -349 245 349 283
rect -349 217 -344 245
rect -316 217 -278 245
rect -250 217 -212 245
rect -184 217 -146 245
rect -118 217 -80 245
rect -52 217 -14 245
rect 14 217 52 245
rect 80 217 118 245
rect 146 217 184 245
rect 212 217 250 245
rect 278 217 316 245
rect 344 217 349 245
rect -349 179 349 217
rect -349 151 -344 179
rect -316 151 -278 179
rect -250 151 -212 179
rect -184 151 -146 179
rect -118 151 -80 179
rect -52 151 -14 179
rect 14 151 52 179
rect 80 151 118 179
rect 146 151 184 179
rect 212 151 250 179
rect 278 151 316 179
rect 344 151 349 179
rect -349 113 349 151
rect -349 85 -344 113
rect -316 85 -278 113
rect -250 85 -212 113
rect -184 85 -146 113
rect -118 85 -80 113
rect -52 85 -14 113
rect 14 85 52 113
rect 80 85 118 113
rect 146 85 184 113
rect 212 85 250 113
rect 278 85 316 113
rect 344 85 349 113
rect -349 47 349 85
rect -349 19 -344 47
rect -316 19 -278 47
rect -250 19 -212 47
rect -184 19 -146 47
rect -118 19 -80 47
rect -52 19 -14 47
rect 14 19 52 47
rect 80 19 118 47
rect 146 19 184 47
rect 212 19 250 47
rect 278 19 316 47
rect 344 19 349 47
rect -349 -19 349 19
rect -349 -47 -344 -19
rect -316 -47 -278 -19
rect -250 -47 -212 -19
rect -184 -47 -146 -19
rect -118 -47 -80 -19
rect -52 -47 -14 -19
rect 14 -47 52 -19
rect 80 -47 118 -19
rect 146 -47 184 -19
rect 212 -47 250 -19
rect 278 -47 316 -19
rect 344 -47 349 -19
rect -349 -85 349 -47
rect -349 -113 -344 -85
rect -316 -113 -278 -85
rect -250 -113 -212 -85
rect -184 -113 -146 -85
rect -118 -113 -80 -85
rect -52 -113 -14 -85
rect 14 -113 52 -85
rect 80 -113 118 -85
rect 146 -113 184 -85
rect 212 -113 250 -85
rect 278 -113 316 -85
rect 344 -113 349 -85
rect -349 -151 349 -113
rect -349 -179 -344 -151
rect -316 -179 -278 -151
rect -250 -179 -212 -151
rect -184 -179 -146 -151
rect -118 -179 -80 -151
rect -52 -179 -14 -151
rect 14 -179 52 -151
rect 80 -179 118 -151
rect 146 -179 184 -151
rect 212 -179 250 -151
rect 278 -179 316 -151
rect 344 -179 349 -151
rect -349 -217 349 -179
rect -349 -245 -344 -217
rect -316 -245 -278 -217
rect -250 -245 -212 -217
rect -184 -245 -146 -217
rect -118 -245 -80 -217
rect -52 -245 -14 -217
rect 14 -245 52 -217
rect 80 -245 118 -217
rect 146 -245 184 -217
rect 212 -245 250 -217
rect 278 -245 316 -217
rect 344 -245 349 -217
rect -349 -283 349 -245
rect -349 -311 -344 -283
rect -316 -311 -278 -283
rect -250 -311 -212 -283
rect -184 -311 -146 -283
rect -118 -311 -80 -283
rect -52 -311 -14 -283
rect 14 -311 52 -283
rect 80 -311 118 -283
rect 146 -311 184 -283
rect 212 -311 250 -283
rect 278 -311 316 -283
rect 344 -311 349 -283
rect -349 -349 349 -311
rect -349 -377 -344 -349
rect -316 -377 -278 -349
rect -250 -377 -212 -349
rect -184 -377 -146 -349
rect -118 -377 -80 -349
rect -52 -377 -14 -349
rect 14 -377 52 -349
rect 80 -377 118 -349
rect 146 -377 184 -349
rect 212 -377 250 -349
rect 278 -377 316 -349
rect 344 -377 349 -349
rect -349 -415 349 -377
rect -349 -443 -344 -415
rect -316 -443 -278 -415
rect -250 -443 -212 -415
rect -184 -443 -146 -415
rect -118 -443 -80 -415
rect -52 -443 -14 -415
rect 14 -443 52 -415
rect 80 -443 118 -415
rect 146 -443 184 -415
rect 212 -443 250 -415
rect 278 -443 316 -415
rect 344 -443 349 -415
rect -349 -481 349 -443
rect -349 -509 -344 -481
rect -316 -509 -278 -481
rect -250 -509 -212 -481
rect -184 -509 -146 -481
rect -118 -509 -80 -481
rect -52 -509 -14 -481
rect 14 -509 52 -481
rect 80 -509 118 -481
rect 146 -509 184 -481
rect 212 -509 250 -481
rect 278 -509 316 -481
rect 344 -509 349 -481
rect -349 -547 349 -509
rect -349 -575 -344 -547
rect -316 -575 -278 -547
rect -250 -575 -212 -547
rect -184 -575 -146 -547
rect -118 -575 -80 -547
rect -52 -575 -14 -547
rect 14 -575 52 -547
rect 80 -575 118 -547
rect 146 -575 184 -547
rect 212 -575 250 -547
rect 278 -575 316 -547
rect 344 -575 349 -547
rect -349 -613 349 -575
rect -349 -641 -344 -613
rect -316 -641 -278 -613
rect -250 -641 -212 -613
rect -184 -641 -146 -613
rect -118 -641 -80 -613
rect -52 -641 -14 -613
rect 14 -641 52 -613
rect 80 -641 118 -613
rect 146 -641 184 -613
rect 212 -641 250 -613
rect 278 -641 316 -613
rect 344 -641 349 -613
rect -349 -679 349 -641
rect -349 -707 -344 -679
rect -316 -707 -278 -679
rect -250 -707 -212 -679
rect -184 -707 -146 -679
rect -118 -707 -80 -679
rect -52 -707 -14 -679
rect 14 -707 52 -679
rect 80 -707 118 -679
rect 146 -707 184 -679
rect 212 -707 250 -679
rect 278 -707 316 -679
rect 344 -707 349 -679
rect -349 -745 349 -707
rect -349 -773 -344 -745
rect -316 -773 -278 -745
rect -250 -773 -212 -745
rect -184 -773 -146 -745
rect -118 -773 -80 -745
rect -52 -773 -14 -745
rect 14 -773 52 -745
rect 80 -773 118 -745
rect 146 -773 184 -745
rect 212 -773 250 -745
rect 278 -773 316 -745
rect 344 -773 349 -745
rect -349 -811 349 -773
rect -349 -839 -344 -811
rect -316 -839 -278 -811
rect -250 -839 -212 -811
rect -184 -839 -146 -811
rect -118 -839 -80 -811
rect -52 -839 -14 -811
rect 14 -839 52 -811
rect 80 -839 118 -811
rect 146 -839 184 -811
rect 212 -839 250 -811
rect 278 -839 316 -811
rect 344 -839 349 -811
rect -349 -877 349 -839
rect -349 -905 -344 -877
rect -316 -905 -278 -877
rect -250 -905 -212 -877
rect -184 -905 -146 -877
rect -118 -905 -80 -877
rect -52 -905 -14 -877
rect 14 -905 52 -877
rect 80 -905 118 -877
rect 146 -905 184 -877
rect 212 -905 250 -877
rect 278 -905 316 -877
rect 344 -905 349 -877
rect -349 -943 349 -905
rect -349 -971 -344 -943
rect -316 -971 -278 -943
rect -250 -971 -212 -943
rect -184 -971 -146 -943
rect -118 -971 -80 -943
rect -52 -971 -14 -943
rect 14 -971 52 -943
rect 80 -971 118 -943
rect 146 -971 184 -943
rect 212 -971 250 -943
rect 278 -971 316 -943
rect 344 -971 349 -943
rect -349 -1009 349 -971
rect -349 -1037 -344 -1009
rect -316 -1037 -278 -1009
rect -250 -1037 -212 -1009
rect -184 -1037 -146 -1009
rect -118 -1037 -80 -1009
rect -52 -1037 -14 -1009
rect 14 -1037 52 -1009
rect 80 -1037 118 -1009
rect 146 -1037 184 -1009
rect 212 -1037 250 -1009
rect 278 -1037 316 -1009
rect 344 -1037 349 -1009
rect -349 -1075 349 -1037
rect -349 -1103 -344 -1075
rect -316 -1103 -278 -1075
rect -250 -1103 -212 -1075
rect -184 -1103 -146 -1075
rect -118 -1103 -80 -1075
rect -52 -1103 -14 -1075
rect 14 -1103 52 -1075
rect 80 -1103 118 -1075
rect 146 -1103 184 -1075
rect 212 -1103 250 -1075
rect 278 -1103 316 -1075
rect 344 -1103 349 -1075
rect -349 -1141 349 -1103
rect -349 -1169 -344 -1141
rect -316 -1169 -278 -1141
rect -250 -1169 -212 -1141
rect -184 -1169 -146 -1141
rect -118 -1169 -80 -1141
rect -52 -1169 -14 -1141
rect 14 -1169 52 -1141
rect 80 -1169 118 -1141
rect 146 -1169 184 -1141
rect 212 -1169 250 -1141
rect 278 -1169 316 -1141
rect 344 -1169 349 -1141
rect -349 -1207 349 -1169
rect -349 -1235 -344 -1207
rect -316 -1235 -278 -1207
rect -250 -1235 -212 -1207
rect -184 -1235 -146 -1207
rect -118 -1235 -80 -1207
rect -52 -1235 -14 -1207
rect 14 -1235 52 -1207
rect 80 -1235 118 -1207
rect 146 -1235 184 -1207
rect 212 -1235 250 -1207
rect 278 -1235 316 -1207
rect 344 -1235 349 -1207
rect -349 -1273 349 -1235
rect -349 -1301 -344 -1273
rect -316 -1301 -278 -1273
rect -250 -1301 -212 -1273
rect -184 -1301 -146 -1273
rect -118 -1301 -80 -1273
rect -52 -1301 -14 -1273
rect 14 -1301 52 -1273
rect 80 -1301 118 -1273
rect 146 -1301 184 -1273
rect 212 -1301 250 -1273
rect 278 -1301 316 -1273
rect 344 -1301 349 -1273
rect -349 -1339 349 -1301
rect -349 -1367 -344 -1339
rect -316 -1367 -278 -1339
rect -250 -1367 -212 -1339
rect -184 -1367 -146 -1339
rect -118 -1367 -80 -1339
rect -52 -1367 -14 -1339
rect 14 -1367 52 -1339
rect 80 -1367 118 -1339
rect 146 -1367 184 -1339
rect 212 -1367 250 -1339
rect 278 -1367 316 -1339
rect 344 -1367 349 -1339
rect -349 -1372 349 -1367
<< via3 >>
rect -344 1339 -316 1367
rect -278 1339 -250 1367
rect -212 1339 -184 1367
rect -146 1339 -118 1367
rect -80 1339 -52 1367
rect -14 1339 14 1367
rect 52 1339 80 1367
rect 118 1339 146 1367
rect 184 1339 212 1367
rect 250 1339 278 1367
rect 316 1339 344 1367
rect -344 1273 -316 1301
rect -278 1273 -250 1301
rect -212 1273 -184 1301
rect -146 1273 -118 1301
rect -80 1273 -52 1301
rect -14 1273 14 1301
rect 52 1273 80 1301
rect 118 1273 146 1301
rect 184 1273 212 1301
rect 250 1273 278 1301
rect 316 1273 344 1301
rect -344 1207 -316 1235
rect -278 1207 -250 1235
rect -212 1207 -184 1235
rect -146 1207 -118 1235
rect -80 1207 -52 1235
rect -14 1207 14 1235
rect 52 1207 80 1235
rect 118 1207 146 1235
rect 184 1207 212 1235
rect 250 1207 278 1235
rect 316 1207 344 1235
rect -344 1141 -316 1169
rect -278 1141 -250 1169
rect -212 1141 -184 1169
rect -146 1141 -118 1169
rect -80 1141 -52 1169
rect -14 1141 14 1169
rect 52 1141 80 1169
rect 118 1141 146 1169
rect 184 1141 212 1169
rect 250 1141 278 1169
rect 316 1141 344 1169
rect -344 1075 -316 1103
rect -278 1075 -250 1103
rect -212 1075 -184 1103
rect -146 1075 -118 1103
rect -80 1075 -52 1103
rect -14 1075 14 1103
rect 52 1075 80 1103
rect 118 1075 146 1103
rect 184 1075 212 1103
rect 250 1075 278 1103
rect 316 1075 344 1103
rect -344 1009 -316 1037
rect -278 1009 -250 1037
rect -212 1009 -184 1037
rect -146 1009 -118 1037
rect -80 1009 -52 1037
rect -14 1009 14 1037
rect 52 1009 80 1037
rect 118 1009 146 1037
rect 184 1009 212 1037
rect 250 1009 278 1037
rect 316 1009 344 1037
rect -344 943 -316 971
rect -278 943 -250 971
rect -212 943 -184 971
rect -146 943 -118 971
rect -80 943 -52 971
rect -14 943 14 971
rect 52 943 80 971
rect 118 943 146 971
rect 184 943 212 971
rect 250 943 278 971
rect 316 943 344 971
rect -344 877 -316 905
rect -278 877 -250 905
rect -212 877 -184 905
rect -146 877 -118 905
rect -80 877 -52 905
rect -14 877 14 905
rect 52 877 80 905
rect 118 877 146 905
rect 184 877 212 905
rect 250 877 278 905
rect 316 877 344 905
rect -344 811 -316 839
rect -278 811 -250 839
rect -212 811 -184 839
rect -146 811 -118 839
rect -80 811 -52 839
rect -14 811 14 839
rect 52 811 80 839
rect 118 811 146 839
rect 184 811 212 839
rect 250 811 278 839
rect 316 811 344 839
rect -344 745 -316 773
rect -278 745 -250 773
rect -212 745 -184 773
rect -146 745 -118 773
rect -80 745 -52 773
rect -14 745 14 773
rect 52 745 80 773
rect 118 745 146 773
rect 184 745 212 773
rect 250 745 278 773
rect 316 745 344 773
rect -344 679 -316 707
rect -278 679 -250 707
rect -212 679 -184 707
rect -146 679 -118 707
rect -80 679 -52 707
rect -14 679 14 707
rect 52 679 80 707
rect 118 679 146 707
rect 184 679 212 707
rect 250 679 278 707
rect 316 679 344 707
rect -344 613 -316 641
rect -278 613 -250 641
rect -212 613 -184 641
rect -146 613 -118 641
rect -80 613 -52 641
rect -14 613 14 641
rect 52 613 80 641
rect 118 613 146 641
rect 184 613 212 641
rect 250 613 278 641
rect 316 613 344 641
rect -344 547 -316 575
rect -278 547 -250 575
rect -212 547 -184 575
rect -146 547 -118 575
rect -80 547 -52 575
rect -14 547 14 575
rect 52 547 80 575
rect 118 547 146 575
rect 184 547 212 575
rect 250 547 278 575
rect 316 547 344 575
rect -344 481 -316 509
rect -278 481 -250 509
rect -212 481 -184 509
rect -146 481 -118 509
rect -80 481 -52 509
rect -14 481 14 509
rect 52 481 80 509
rect 118 481 146 509
rect 184 481 212 509
rect 250 481 278 509
rect 316 481 344 509
rect -344 415 -316 443
rect -278 415 -250 443
rect -212 415 -184 443
rect -146 415 -118 443
rect -80 415 -52 443
rect -14 415 14 443
rect 52 415 80 443
rect 118 415 146 443
rect 184 415 212 443
rect 250 415 278 443
rect 316 415 344 443
rect -344 349 -316 377
rect -278 349 -250 377
rect -212 349 -184 377
rect -146 349 -118 377
rect -80 349 -52 377
rect -14 349 14 377
rect 52 349 80 377
rect 118 349 146 377
rect 184 349 212 377
rect 250 349 278 377
rect 316 349 344 377
rect -344 283 -316 311
rect -278 283 -250 311
rect -212 283 -184 311
rect -146 283 -118 311
rect -80 283 -52 311
rect -14 283 14 311
rect 52 283 80 311
rect 118 283 146 311
rect 184 283 212 311
rect 250 283 278 311
rect 316 283 344 311
rect -344 217 -316 245
rect -278 217 -250 245
rect -212 217 -184 245
rect -146 217 -118 245
rect -80 217 -52 245
rect -14 217 14 245
rect 52 217 80 245
rect 118 217 146 245
rect 184 217 212 245
rect 250 217 278 245
rect 316 217 344 245
rect -344 151 -316 179
rect -278 151 -250 179
rect -212 151 -184 179
rect -146 151 -118 179
rect -80 151 -52 179
rect -14 151 14 179
rect 52 151 80 179
rect 118 151 146 179
rect 184 151 212 179
rect 250 151 278 179
rect 316 151 344 179
rect -344 85 -316 113
rect -278 85 -250 113
rect -212 85 -184 113
rect -146 85 -118 113
rect -80 85 -52 113
rect -14 85 14 113
rect 52 85 80 113
rect 118 85 146 113
rect 184 85 212 113
rect 250 85 278 113
rect 316 85 344 113
rect -344 19 -316 47
rect -278 19 -250 47
rect -212 19 -184 47
rect -146 19 -118 47
rect -80 19 -52 47
rect -14 19 14 47
rect 52 19 80 47
rect 118 19 146 47
rect 184 19 212 47
rect 250 19 278 47
rect 316 19 344 47
rect -344 -47 -316 -19
rect -278 -47 -250 -19
rect -212 -47 -184 -19
rect -146 -47 -118 -19
rect -80 -47 -52 -19
rect -14 -47 14 -19
rect 52 -47 80 -19
rect 118 -47 146 -19
rect 184 -47 212 -19
rect 250 -47 278 -19
rect 316 -47 344 -19
rect -344 -113 -316 -85
rect -278 -113 -250 -85
rect -212 -113 -184 -85
rect -146 -113 -118 -85
rect -80 -113 -52 -85
rect -14 -113 14 -85
rect 52 -113 80 -85
rect 118 -113 146 -85
rect 184 -113 212 -85
rect 250 -113 278 -85
rect 316 -113 344 -85
rect -344 -179 -316 -151
rect -278 -179 -250 -151
rect -212 -179 -184 -151
rect -146 -179 -118 -151
rect -80 -179 -52 -151
rect -14 -179 14 -151
rect 52 -179 80 -151
rect 118 -179 146 -151
rect 184 -179 212 -151
rect 250 -179 278 -151
rect 316 -179 344 -151
rect -344 -245 -316 -217
rect -278 -245 -250 -217
rect -212 -245 -184 -217
rect -146 -245 -118 -217
rect -80 -245 -52 -217
rect -14 -245 14 -217
rect 52 -245 80 -217
rect 118 -245 146 -217
rect 184 -245 212 -217
rect 250 -245 278 -217
rect 316 -245 344 -217
rect -344 -311 -316 -283
rect -278 -311 -250 -283
rect -212 -311 -184 -283
rect -146 -311 -118 -283
rect -80 -311 -52 -283
rect -14 -311 14 -283
rect 52 -311 80 -283
rect 118 -311 146 -283
rect 184 -311 212 -283
rect 250 -311 278 -283
rect 316 -311 344 -283
rect -344 -377 -316 -349
rect -278 -377 -250 -349
rect -212 -377 -184 -349
rect -146 -377 -118 -349
rect -80 -377 -52 -349
rect -14 -377 14 -349
rect 52 -377 80 -349
rect 118 -377 146 -349
rect 184 -377 212 -349
rect 250 -377 278 -349
rect 316 -377 344 -349
rect -344 -443 -316 -415
rect -278 -443 -250 -415
rect -212 -443 -184 -415
rect -146 -443 -118 -415
rect -80 -443 -52 -415
rect -14 -443 14 -415
rect 52 -443 80 -415
rect 118 -443 146 -415
rect 184 -443 212 -415
rect 250 -443 278 -415
rect 316 -443 344 -415
rect -344 -509 -316 -481
rect -278 -509 -250 -481
rect -212 -509 -184 -481
rect -146 -509 -118 -481
rect -80 -509 -52 -481
rect -14 -509 14 -481
rect 52 -509 80 -481
rect 118 -509 146 -481
rect 184 -509 212 -481
rect 250 -509 278 -481
rect 316 -509 344 -481
rect -344 -575 -316 -547
rect -278 -575 -250 -547
rect -212 -575 -184 -547
rect -146 -575 -118 -547
rect -80 -575 -52 -547
rect -14 -575 14 -547
rect 52 -575 80 -547
rect 118 -575 146 -547
rect 184 -575 212 -547
rect 250 -575 278 -547
rect 316 -575 344 -547
rect -344 -641 -316 -613
rect -278 -641 -250 -613
rect -212 -641 -184 -613
rect -146 -641 -118 -613
rect -80 -641 -52 -613
rect -14 -641 14 -613
rect 52 -641 80 -613
rect 118 -641 146 -613
rect 184 -641 212 -613
rect 250 -641 278 -613
rect 316 -641 344 -613
rect -344 -707 -316 -679
rect -278 -707 -250 -679
rect -212 -707 -184 -679
rect -146 -707 -118 -679
rect -80 -707 -52 -679
rect -14 -707 14 -679
rect 52 -707 80 -679
rect 118 -707 146 -679
rect 184 -707 212 -679
rect 250 -707 278 -679
rect 316 -707 344 -679
rect -344 -773 -316 -745
rect -278 -773 -250 -745
rect -212 -773 -184 -745
rect -146 -773 -118 -745
rect -80 -773 -52 -745
rect -14 -773 14 -745
rect 52 -773 80 -745
rect 118 -773 146 -745
rect 184 -773 212 -745
rect 250 -773 278 -745
rect 316 -773 344 -745
rect -344 -839 -316 -811
rect -278 -839 -250 -811
rect -212 -839 -184 -811
rect -146 -839 -118 -811
rect -80 -839 -52 -811
rect -14 -839 14 -811
rect 52 -839 80 -811
rect 118 -839 146 -811
rect 184 -839 212 -811
rect 250 -839 278 -811
rect 316 -839 344 -811
rect -344 -905 -316 -877
rect -278 -905 -250 -877
rect -212 -905 -184 -877
rect -146 -905 -118 -877
rect -80 -905 -52 -877
rect -14 -905 14 -877
rect 52 -905 80 -877
rect 118 -905 146 -877
rect 184 -905 212 -877
rect 250 -905 278 -877
rect 316 -905 344 -877
rect -344 -971 -316 -943
rect -278 -971 -250 -943
rect -212 -971 -184 -943
rect -146 -971 -118 -943
rect -80 -971 -52 -943
rect -14 -971 14 -943
rect 52 -971 80 -943
rect 118 -971 146 -943
rect 184 -971 212 -943
rect 250 -971 278 -943
rect 316 -971 344 -943
rect -344 -1037 -316 -1009
rect -278 -1037 -250 -1009
rect -212 -1037 -184 -1009
rect -146 -1037 -118 -1009
rect -80 -1037 -52 -1009
rect -14 -1037 14 -1009
rect 52 -1037 80 -1009
rect 118 -1037 146 -1009
rect 184 -1037 212 -1009
rect 250 -1037 278 -1009
rect 316 -1037 344 -1009
rect -344 -1103 -316 -1075
rect -278 -1103 -250 -1075
rect -212 -1103 -184 -1075
rect -146 -1103 -118 -1075
rect -80 -1103 -52 -1075
rect -14 -1103 14 -1075
rect 52 -1103 80 -1075
rect 118 -1103 146 -1075
rect 184 -1103 212 -1075
rect 250 -1103 278 -1075
rect 316 -1103 344 -1075
rect -344 -1169 -316 -1141
rect -278 -1169 -250 -1141
rect -212 -1169 -184 -1141
rect -146 -1169 -118 -1141
rect -80 -1169 -52 -1141
rect -14 -1169 14 -1141
rect 52 -1169 80 -1141
rect 118 -1169 146 -1141
rect 184 -1169 212 -1141
rect 250 -1169 278 -1141
rect 316 -1169 344 -1141
rect -344 -1235 -316 -1207
rect -278 -1235 -250 -1207
rect -212 -1235 -184 -1207
rect -146 -1235 -118 -1207
rect -80 -1235 -52 -1207
rect -14 -1235 14 -1207
rect 52 -1235 80 -1207
rect 118 -1235 146 -1207
rect 184 -1235 212 -1207
rect 250 -1235 278 -1207
rect 316 -1235 344 -1207
rect -344 -1301 -316 -1273
rect -278 -1301 -250 -1273
rect -212 -1301 -184 -1273
rect -146 -1301 -118 -1273
rect -80 -1301 -52 -1273
rect -14 -1301 14 -1273
rect 52 -1301 80 -1273
rect 118 -1301 146 -1273
rect 184 -1301 212 -1273
rect 250 -1301 278 -1273
rect 316 -1301 344 -1273
rect -344 -1367 -316 -1339
rect -278 -1367 -250 -1339
rect -212 -1367 -184 -1339
rect -146 -1367 -118 -1339
rect -80 -1367 -52 -1339
rect -14 -1367 14 -1339
rect 52 -1367 80 -1339
rect 118 -1367 146 -1339
rect 184 -1367 212 -1339
rect 250 -1367 278 -1339
rect 316 -1367 344 -1339
<< metal4 >>
rect -349 1367 349 1372
rect -349 1339 -344 1367
rect -316 1339 -278 1367
rect -250 1339 -212 1367
rect -184 1339 -146 1367
rect -118 1339 -80 1367
rect -52 1339 -14 1367
rect 14 1339 52 1367
rect 80 1339 118 1367
rect 146 1339 184 1367
rect 212 1339 250 1367
rect 278 1339 316 1367
rect 344 1339 349 1367
rect -349 1301 349 1339
rect -349 1273 -344 1301
rect -316 1273 -278 1301
rect -250 1273 -212 1301
rect -184 1273 -146 1301
rect -118 1273 -80 1301
rect -52 1273 -14 1301
rect 14 1273 52 1301
rect 80 1273 118 1301
rect 146 1273 184 1301
rect 212 1273 250 1301
rect 278 1273 316 1301
rect 344 1273 349 1301
rect -349 1235 349 1273
rect -349 1207 -344 1235
rect -316 1207 -278 1235
rect -250 1207 -212 1235
rect -184 1207 -146 1235
rect -118 1207 -80 1235
rect -52 1207 -14 1235
rect 14 1207 52 1235
rect 80 1207 118 1235
rect 146 1207 184 1235
rect 212 1207 250 1235
rect 278 1207 316 1235
rect 344 1207 349 1235
rect -349 1169 349 1207
rect -349 1141 -344 1169
rect -316 1141 -278 1169
rect -250 1141 -212 1169
rect -184 1141 -146 1169
rect -118 1141 -80 1169
rect -52 1141 -14 1169
rect 14 1141 52 1169
rect 80 1141 118 1169
rect 146 1141 184 1169
rect 212 1141 250 1169
rect 278 1141 316 1169
rect 344 1141 349 1169
rect -349 1103 349 1141
rect -349 1075 -344 1103
rect -316 1075 -278 1103
rect -250 1075 -212 1103
rect -184 1075 -146 1103
rect -118 1075 -80 1103
rect -52 1075 -14 1103
rect 14 1075 52 1103
rect 80 1075 118 1103
rect 146 1075 184 1103
rect 212 1075 250 1103
rect 278 1075 316 1103
rect 344 1075 349 1103
rect -349 1037 349 1075
rect -349 1009 -344 1037
rect -316 1009 -278 1037
rect -250 1009 -212 1037
rect -184 1009 -146 1037
rect -118 1009 -80 1037
rect -52 1009 -14 1037
rect 14 1009 52 1037
rect 80 1009 118 1037
rect 146 1009 184 1037
rect 212 1009 250 1037
rect 278 1009 316 1037
rect 344 1009 349 1037
rect -349 971 349 1009
rect -349 943 -344 971
rect -316 943 -278 971
rect -250 943 -212 971
rect -184 943 -146 971
rect -118 943 -80 971
rect -52 943 -14 971
rect 14 943 52 971
rect 80 943 118 971
rect 146 943 184 971
rect 212 943 250 971
rect 278 943 316 971
rect 344 943 349 971
rect -349 905 349 943
rect -349 877 -344 905
rect -316 877 -278 905
rect -250 877 -212 905
rect -184 877 -146 905
rect -118 877 -80 905
rect -52 877 -14 905
rect 14 877 52 905
rect 80 877 118 905
rect 146 877 184 905
rect 212 877 250 905
rect 278 877 316 905
rect 344 877 349 905
rect -349 839 349 877
rect -349 811 -344 839
rect -316 811 -278 839
rect -250 811 -212 839
rect -184 811 -146 839
rect -118 811 -80 839
rect -52 811 -14 839
rect 14 811 52 839
rect 80 811 118 839
rect 146 811 184 839
rect 212 811 250 839
rect 278 811 316 839
rect 344 811 349 839
rect -349 773 349 811
rect -349 745 -344 773
rect -316 745 -278 773
rect -250 745 -212 773
rect -184 745 -146 773
rect -118 745 -80 773
rect -52 745 -14 773
rect 14 745 52 773
rect 80 745 118 773
rect 146 745 184 773
rect 212 745 250 773
rect 278 745 316 773
rect 344 745 349 773
rect -349 707 349 745
rect -349 679 -344 707
rect -316 679 -278 707
rect -250 679 -212 707
rect -184 679 -146 707
rect -118 679 -80 707
rect -52 679 -14 707
rect 14 679 52 707
rect 80 679 118 707
rect 146 679 184 707
rect 212 679 250 707
rect 278 679 316 707
rect 344 679 349 707
rect -349 641 349 679
rect -349 613 -344 641
rect -316 613 -278 641
rect -250 613 -212 641
rect -184 613 -146 641
rect -118 613 -80 641
rect -52 613 -14 641
rect 14 613 52 641
rect 80 613 118 641
rect 146 613 184 641
rect 212 613 250 641
rect 278 613 316 641
rect 344 613 349 641
rect -349 575 349 613
rect -349 547 -344 575
rect -316 547 -278 575
rect -250 547 -212 575
rect -184 547 -146 575
rect -118 547 -80 575
rect -52 547 -14 575
rect 14 547 52 575
rect 80 547 118 575
rect 146 547 184 575
rect 212 547 250 575
rect 278 547 316 575
rect 344 547 349 575
rect -349 509 349 547
rect -349 481 -344 509
rect -316 481 -278 509
rect -250 481 -212 509
rect -184 481 -146 509
rect -118 481 -80 509
rect -52 481 -14 509
rect 14 481 52 509
rect 80 481 118 509
rect 146 481 184 509
rect 212 481 250 509
rect 278 481 316 509
rect 344 481 349 509
rect -349 443 349 481
rect -349 415 -344 443
rect -316 415 -278 443
rect -250 415 -212 443
rect -184 415 -146 443
rect -118 415 -80 443
rect -52 415 -14 443
rect 14 415 52 443
rect 80 415 118 443
rect 146 415 184 443
rect 212 415 250 443
rect 278 415 316 443
rect 344 415 349 443
rect -349 377 349 415
rect -349 349 -344 377
rect -316 349 -278 377
rect -250 349 -212 377
rect -184 349 -146 377
rect -118 349 -80 377
rect -52 349 -14 377
rect 14 349 52 377
rect 80 349 118 377
rect 146 349 184 377
rect 212 349 250 377
rect 278 349 316 377
rect 344 349 349 377
rect -349 311 349 349
rect -349 283 -344 311
rect -316 283 -278 311
rect -250 283 -212 311
rect -184 283 -146 311
rect -118 283 -80 311
rect -52 283 -14 311
rect 14 283 52 311
rect 80 283 118 311
rect 146 283 184 311
rect 212 283 250 311
rect 278 283 316 311
rect 344 283 349 311
rect -349 245 349 283
rect -349 217 -344 245
rect -316 217 -278 245
rect -250 217 -212 245
rect -184 217 -146 245
rect -118 217 -80 245
rect -52 217 -14 245
rect 14 217 52 245
rect 80 217 118 245
rect 146 217 184 245
rect 212 217 250 245
rect 278 217 316 245
rect 344 217 349 245
rect -349 179 349 217
rect -349 151 -344 179
rect -316 151 -278 179
rect -250 151 -212 179
rect -184 151 -146 179
rect -118 151 -80 179
rect -52 151 -14 179
rect 14 151 52 179
rect 80 151 118 179
rect 146 151 184 179
rect 212 151 250 179
rect 278 151 316 179
rect 344 151 349 179
rect -349 113 349 151
rect -349 85 -344 113
rect -316 85 -278 113
rect -250 85 -212 113
rect -184 85 -146 113
rect -118 85 -80 113
rect -52 85 -14 113
rect 14 85 52 113
rect 80 85 118 113
rect 146 85 184 113
rect 212 85 250 113
rect 278 85 316 113
rect 344 85 349 113
rect -349 47 349 85
rect -349 19 -344 47
rect -316 19 -278 47
rect -250 19 -212 47
rect -184 19 -146 47
rect -118 19 -80 47
rect -52 19 -14 47
rect 14 19 52 47
rect 80 19 118 47
rect 146 19 184 47
rect 212 19 250 47
rect 278 19 316 47
rect 344 19 349 47
rect -349 -19 349 19
rect -349 -47 -344 -19
rect -316 -47 -278 -19
rect -250 -47 -212 -19
rect -184 -47 -146 -19
rect -118 -47 -80 -19
rect -52 -47 -14 -19
rect 14 -47 52 -19
rect 80 -47 118 -19
rect 146 -47 184 -19
rect 212 -47 250 -19
rect 278 -47 316 -19
rect 344 -47 349 -19
rect -349 -85 349 -47
rect -349 -113 -344 -85
rect -316 -113 -278 -85
rect -250 -113 -212 -85
rect -184 -113 -146 -85
rect -118 -113 -80 -85
rect -52 -113 -14 -85
rect 14 -113 52 -85
rect 80 -113 118 -85
rect 146 -113 184 -85
rect 212 -113 250 -85
rect 278 -113 316 -85
rect 344 -113 349 -85
rect -349 -151 349 -113
rect -349 -179 -344 -151
rect -316 -179 -278 -151
rect -250 -179 -212 -151
rect -184 -179 -146 -151
rect -118 -179 -80 -151
rect -52 -179 -14 -151
rect 14 -179 52 -151
rect 80 -179 118 -151
rect 146 -179 184 -151
rect 212 -179 250 -151
rect 278 -179 316 -151
rect 344 -179 349 -151
rect -349 -217 349 -179
rect -349 -245 -344 -217
rect -316 -245 -278 -217
rect -250 -245 -212 -217
rect -184 -245 -146 -217
rect -118 -245 -80 -217
rect -52 -245 -14 -217
rect 14 -245 52 -217
rect 80 -245 118 -217
rect 146 -245 184 -217
rect 212 -245 250 -217
rect 278 -245 316 -217
rect 344 -245 349 -217
rect -349 -283 349 -245
rect -349 -311 -344 -283
rect -316 -311 -278 -283
rect -250 -311 -212 -283
rect -184 -311 -146 -283
rect -118 -311 -80 -283
rect -52 -311 -14 -283
rect 14 -311 52 -283
rect 80 -311 118 -283
rect 146 -311 184 -283
rect 212 -311 250 -283
rect 278 -311 316 -283
rect 344 -311 349 -283
rect -349 -349 349 -311
rect -349 -377 -344 -349
rect -316 -377 -278 -349
rect -250 -377 -212 -349
rect -184 -377 -146 -349
rect -118 -377 -80 -349
rect -52 -377 -14 -349
rect 14 -377 52 -349
rect 80 -377 118 -349
rect 146 -377 184 -349
rect 212 -377 250 -349
rect 278 -377 316 -349
rect 344 -377 349 -349
rect -349 -415 349 -377
rect -349 -443 -344 -415
rect -316 -443 -278 -415
rect -250 -443 -212 -415
rect -184 -443 -146 -415
rect -118 -443 -80 -415
rect -52 -443 -14 -415
rect 14 -443 52 -415
rect 80 -443 118 -415
rect 146 -443 184 -415
rect 212 -443 250 -415
rect 278 -443 316 -415
rect 344 -443 349 -415
rect -349 -481 349 -443
rect -349 -509 -344 -481
rect -316 -509 -278 -481
rect -250 -509 -212 -481
rect -184 -509 -146 -481
rect -118 -509 -80 -481
rect -52 -509 -14 -481
rect 14 -509 52 -481
rect 80 -509 118 -481
rect 146 -509 184 -481
rect 212 -509 250 -481
rect 278 -509 316 -481
rect 344 -509 349 -481
rect -349 -547 349 -509
rect -349 -575 -344 -547
rect -316 -575 -278 -547
rect -250 -575 -212 -547
rect -184 -575 -146 -547
rect -118 -575 -80 -547
rect -52 -575 -14 -547
rect 14 -575 52 -547
rect 80 -575 118 -547
rect 146 -575 184 -547
rect 212 -575 250 -547
rect 278 -575 316 -547
rect 344 -575 349 -547
rect -349 -613 349 -575
rect -349 -641 -344 -613
rect -316 -641 -278 -613
rect -250 -641 -212 -613
rect -184 -641 -146 -613
rect -118 -641 -80 -613
rect -52 -641 -14 -613
rect 14 -641 52 -613
rect 80 -641 118 -613
rect 146 -641 184 -613
rect 212 -641 250 -613
rect 278 -641 316 -613
rect 344 -641 349 -613
rect -349 -679 349 -641
rect -349 -707 -344 -679
rect -316 -707 -278 -679
rect -250 -707 -212 -679
rect -184 -707 -146 -679
rect -118 -707 -80 -679
rect -52 -707 -14 -679
rect 14 -707 52 -679
rect 80 -707 118 -679
rect 146 -707 184 -679
rect 212 -707 250 -679
rect 278 -707 316 -679
rect 344 -707 349 -679
rect -349 -745 349 -707
rect -349 -773 -344 -745
rect -316 -773 -278 -745
rect -250 -773 -212 -745
rect -184 -773 -146 -745
rect -118 -773 -80 -745
rect -52 -773 -14 -745
rect 14 -773 52 -745
rect 80 -773 118 -745
rect 146 -773 184 -745
rect 212 -773 250 -745
rect 278 -773 316 -745
rect 344 -773 349 -745
rect -349 -811 349 -773
rect -349 -839 -344 -811
rect -316 -839 -278 -811
rect -250 -839 -212 -811
rect -184 -839 -146 -811
rect -118 -839 -80 -811
rect -52 -839 -14 -811
rect 14 -839 52 -811
rect 80 -839 118 -811
rect 146 -839 184 -811
rect 212 -839 250 -811
rect 278 -839 316 -811
rect 344 -839 349 -811
rect -349 -877 349 -839
rect -349 -905 -344 -877
rect -316 -905 -278 -877
rect -250 -905 -212 -877
rect -184 -905 -146 -877
rect -118 -905 -80 -877
rect -52 -905 -14 -877
rect 14 -905 52 -877
rect 80 -905 118 -877
rect 146 -905 184 -877
rect 212 -905 250 -877
rect 278 -905 316 -877
rect 344 -905 349 -877
rect -349 -943 349 -905
rect -349 -971 -344 -943
rect -316 -971 -278 -943
rect -250 -971 -212 -943
rect -184 -971 -146 -943
rect -118 -971 -80 -943
rect -52 -971 -14 -943
rect 14 -971 52 -943
rect 80 -971 118 -943
rect 146 -971 184 -943
rect 212 -971 250 -943
rect 278 -971 316 -943
rect 344 -971 349 -943
rect -349 -1009 349 -971
rect -349 -1037 -344 -1009
rect -316 -1037 -278 -1009
rect -250 -1037 -212 -1009
rect -184 -1037 -146 -1009
rect -118 -1037 -80 -1009
rect -52 -1037 -14 -1009
rect 14 -1037 52 -1009
rect 80 -1037 118 -1009
rect 146 -1037 184 -1009
rect 212 -1037 250 -1009
rect 278 -1037 316 -1009
rect 344 -1037 349 -1009
rect -349 -1075 349 -1037
rect -349 -1103 -344 -1075
rect -316 -1103 -278 -1075
rect -250 -1103 -212 -1075
rect -184 -1103 -146 -1075
rect -118 -1103 -80 -1075
rect -52 -1103 -14 -1075
rect 14 -1103 52 -1075
rect 80 -1103 118 -1075
rect 146 -1103 184 -1075
rect 212 -1103 250 -1075
rect 278 -1103 316 -1075
rect 344 -1103 349 -1075
rect -349 -1141 349 -1103
rect -349 -1169 -344 -1141
rect -316 -1169 -278 -1141
rect -250 -1169 -212 -1141
rect -184 -1169 -146 -1141
rect -118 -1169 -80 -1141
rect -52 -1169 -14 -1141
rect 14 -1169 52 -1141
rect 80 -1169 118 -1141
rect 146 -1169 184 -1141
rect 212 -1169 250 -1141
rect 278 -1169 316 -1141
rect 344 -1169 349 -1141
rect -349 -1207 349 -1169
rect -349 -1235 -344 -1207
rect -316 -1235 -278 -1207
rect -250 -1235 -212 -1207
rect -184 -1235 -146 -1207
rect -118 -1235 -80 -1207
rect -52 -1235 -14 -1207
rect 14 -1235 52 -1207
rect 80 -1235 118 -1207
rect 146 -1235 184 -1207
rect 212 -1235 250 -1207
rect 278 -1235 316 -1207
rect 344 -1235 349 -1207
rect -349 -1273 349 -1235
rect -349 -1301 -344 -1273
rect -316 -1301 -278 -1273
rect -250 -1301 -212 -1273
rect -184 -1301 -146 -1273
rect -118 -1301 -80 -1273
rect -52 -1301 -14 -1273
rect 14 -1301 52 -1273
rect 80 -1301 118 -1273
rect 146 -1301 184 -1273
rect 212 -1301 250 -1273
rect 278 -1301 316 -1273
rect 344 -1301 349 -1273
rect -349 -1339 349 -1301
rect -349 -1367 -344 -1339
rect -316 -1367 -278 -1339
rect -250 -1367 -212 -1339
rect -184 -1367 -146 -1339
rect -118 -1367 -80 -1339
rect -52 -1367 -14 -1339
rect 14 -1367 52 -1339
rect 80 -1367 118 -1339
rect 146 -1367 184 -1339
rect 212 -1367 250 -1339
rect 278 -1367 316 -1339
rect 344 -1367 349 -1339
rect -349 -1372 349 -1367
<< end >>
