** sch_path: /home/shahid/GF180Projects/Top_test3/Top_test/top/xschem/pex_CLK_div_96_TB.sch
**.subckt pex_CLK_div_96_TB
V1 VDD VSS 3.3
.save i(v1)
V2 VSS GND 0
.save i(v2)
V3 CLK VSS pulse(3.3 0 0 100p 100p 2.50n 5n)
.save i(v3)
C5 Vdiv96 VSS 10f m=1
V5 RST VSS PWL( 0 0 10n 0 10.001n 3)
.save i(v5)
x1 VSS VDD RST Vdiv96 CLK pex_CLK_div_96_mag
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.include pex_CLK_div_96_mag.spice
.control
save all
tran 1n 1u
plot v(CLK) v(Vdiv96)+3.5 v(RST)+7
*write pex_CLK_div_96_TB.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
