** sch_path: /home/shahid/GF180Projects/Top_test/top/xschem/pex_PFD_test.sch
**.subckt pex_PFD_test
V1 VDD VSS 3.3
.save i(v1)
V2 VSS GND 0
.save i(v2)
V3 VDIV VSS pulse(3.3 0 10n 100p 100p 50n 100n)
.save i(v3)
V4 VREF VSS pulse(3.3 0 0 100p 100p 50n 100n)
.save i(v4)
C1 PD VSS 50f m=1
C2 PU VSS 50f m=1
x1 VSS VREF VDIV PU PD VDD pex_PFD_layout
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.include pex_PFD_layout.spice
.control
save all
tran 50p 500n
plot v(VREF) V(VDIV)+5 v(PU)+10 v(PD)+15
*write test_nfet_03v3.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
