magic
tech gf180mcuC
magscale 1 10
timestamp 1692005851
<< nwell >>
rect 0 310 884 901
<< pwell >>
rect 222 0 662 236
<< nmos >>
rect 334 68 390 168
rect 494 68 550 168
<< pmos >>
rect 174 440 230 640
rect 334 440 390 640
rect 494 440 550 640
rect 654 440 710 640
<< ndiff >>
rect 246 155 334 168
rect 246 81 259 155
rect 305 81 334 155
rect 246 68 334 81
rect 390 155 494 168
rect 390 81 419 155
rect 465 81 494 155
rect 390 68 494 81
rect 550 155 638 168
rect 550 81 579 155
rect 625 81 638 155
rect 550 68 638 81
<< pdiff >>
rect 86 627 174 640
rect 86 453 99 627
rect 145 453 174 627
rect 86 440 174 453
rect 230 627 334 640
rect 230 453 259 627
rect 305 453 334 627
rect 230 440 334 453
rect 390 627 494 640
rect 390 453 419 627
rect 465 453 494 627
rect 390 440 494 453
rect 550 627 654 640
rect 550 453 579 627
rect 625 453 654 627
rect 550 440 654 453
rect 710 627 798 640
rect 710 453 739 627
rect 785 453 798 627
rect 710 440 798 453
<< ndiffc >>
rect 259 81 305 155
rect 419 81 465 155
rect 579 81 625 155
<< pdiffc >>
rect 99 453 145 627
rect 259 453 305 627
rect 419 453 465 627
rect 579 453 625 627
rect 739 453 785 627
<< psubdiff >>
rect 265 -33 619 -20
rect 265 -79 278 -33
rect 324 -79 372 -33
rect 418 -79 466 -33
rect 512 -79 560 -33
rect 606 -79 619 -33
rect 265 -92 619 -79
<< nsubdiff >>
rect 30 855 854 868
rect 30 809 43 855
rect 89 809 137 855
rect 183 809 231 855
rect 277 809 325 855
rect 371 809 419 855
rect 465 809 513 855
rect 559 809 607 855
rect 653 809 701 855
rect 747 809 795 855
rect 841 809 854 855
rect 30 796 854 809
<< psubdiffcont >>
rect 278 -79 324 -33
rect 372 -79 418 -33
rect 466 -79 512 -33
rect 560 -79 606 -33
<< nsubdiffcont >>
rect 43 809 89 855
rect 137 809 183 855
rect 231 809 277 855
rect 325 809 371 855
rect 419 809 465 855
rect 513 809 559 855
rect 607 809 653 855
rect 701 809 747 855
rect 795 809 841 855
<< polysilicon >>
rect 174 640 230 684
rect 334 640 390 684
rect 494 640 550 684
rect 654 640 710 684
rect 174 301 230 440
rect 166 293 238 301
rect 334 293 390 440
rect 166 288 390 293
rect 166 242 179 288
rect 225 242 390 288
rect 166 237 390 242
rect 166 229 238 237
rect 334 168 390 237
rect 494 376 550 440
rect 654 376 710 440
rect 758 376 830 384
rect 494 371 830 376
rect 494 324 771 371
rect 817 324 830 371
rect 494 320 830 324
rect 494 168 550 320
rect 758 311 830 320
rect 334 24 390 68
rect 494 24 550 68
<< polycontact >>
rect 179 242 225 288
rect 771 324 817 371
<< metal1 >>
rect 0 855 884 888
rect 0 809 43 855
rect 89 809 137 855
rect 183 809 231 855
rect 277 809 325 855
rect 371 809 419 855
rect 465 809 513 855
rect 559 809 607 855
rect 653 809 701 855
rect 747 809 795 855
rect 841 809 884 855
rect 0 776 884 809
rect 99 627 145 638
rect 99 396 145 453
rect 259 627 305 776
rect 259 442 305 453
rect 419 684 785 730
rect 419 627 465 684
rect 419 396 465 453
rect 99 350 465 396
rect 579 627 625 638
rect 168 288 236 299
rect 124 242 179 288
rect 225 242 236 288
rect 579 258 625 453
rect 739 627 785 684
rect 739 442 785 453
rect 760 371 828 382
rect 760 324 771 371
rect 817 324 898 371
rect 760 313 828 324
rect 168 231 236 242
rect 419 212 713 258
rect 259 155 305 166
rect 259 0 305 81
rect 419 155 465 212
rect 419 70 465 81
rect 579 155 625 166
rect 579 0 625 81
rect 222 -33 662 0
rect 222 -79 278 -33
rect 324 -79 372 -33
rect 418 -79 466 -33
rect 512 -79 560 -33
rect 606 -79 662 -33
rect 222 -112 662 -79
<< labels >>
flabel metal1 134 265 134 265 0 FreeSans 320 0 0 0 A
port 0 nsew
flabel metal1 884 348 884 348 0 FreeSans 320 0 0 0 B
port 1 nsew
flabel metal1 681 235 681 235 0 FreeSans 320 0 0 0 OUT
port 4 nsew
flabel nsubdiffcont 442 832 442 832 0 FreeSans 320 0 0 0 VDD
port 6 nsew
flabel metal1 437 -56 437 -56 0 FreeSans 320 0 0 0 VSS
port 7 nsew
<< end >>
