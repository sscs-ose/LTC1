magic
tech gf180mcuC
magscale 1 10
timestamp 1691477108
<< error_p >>
rect 83 -455 884 -394
rect 72 -468 895 -455
rect 72 -566 83 -468
rect 96 -492 871 -479
rect 96 -542 107 -492
rect 860 -542 871 -492
rect 96 -555 871 -542
rect 884 -566 895 -468
rect 72 -579 895 -566
<< nwell >>
rect 83 -566 884 -468
<< psubdiff >>
rect 94 -775 869 -760
rect 94 -821 121 -775
rect 167 -821 216 -775
rect 262 -821 314 -775
rect 360 -821 409 -775
rect 455 -821 506 -775
rect 552 -821 601 -775
rect 647 -821 699 -775
rect 745 -821 794 -775
rect 840 -821 869 -775
rect 94 -836 869 -821
<< nsubdiff >>
rect 96 -494 871 -479
rect 96 -540 125 -494
rect 171 -540 219 -494
rect 265 -540 320 -494
rect 366 -540 414 -494
rect 460 -540 510 -494
rect 556 -540 604 -494
rect 650 -540 705 -494
rect 751 -540 799 -494
rect 845 -540 871 -494
rect 96 -555 871 -540
<< psubdiffcont >>
rect 121 -821 167 -775
rect 216 -821 262 -775
rect 314 -821 360 -775
rect 409 -821 455 -775
rect 506 -821 552 -775
rect 601 -821 647 -775
rect 699 -821 745 -775
rect 794 -821 840 -775
<< nsubdiffcont >>
rect 125 -540 171 -494
rect 219 -540 265 -494
rect 320 -540 366 -494
rect 414 -540 460 -494
rect 510 -540 556 -494
rect 604 -540 650 -494
rect 705 -540 751 -494
rect 799 -540 845 -494
<< metal1 >>
rect 83 -494 884 -468
rect 83 -540 125 -494
rect 171 -540 219 -494
rect 265 -540 320 -494
rect 366 -540 414 -494
rect 460 -540 510 -494
rect 556 -540 604 -494
rect 650 -540 705 -494
rect 751 -540 799 -494
rect 845 -540 884 -494
rect 83 -566 884 -540
rect 74 -775 886 -749
rect 74 -821 121 -775
rect 167 -821 216 -775
rect 262 -821 314 -775
rect 360 -821 409 -775
rect 455 -821 506 -775
rect 552 -821 601 -775
rect 647 -821 699 -775
rect 745 -821 794 -775
rect 840 -821 886 -775
rect 74 -846 886 -821
<< end >>
