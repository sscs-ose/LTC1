magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -49022 -57377 11837 2076
<< psubdiff >>
rect -45183 -25693 -44782 -25625
rect -45083 -25871 -44714 -25693
rect -42953 -25739 -42843 -25693
rect -42953 -27561 -42736 -25739
rect -42953 -27629 -40520 -27561
rect -42843 -27682 -40520 -27629
rect -42843 -27751 -8119 -27682
rect -40588 -27881 -8119 -27751
rect -42963 -28013 -40723 -27881
rect -35307 -27949 -35226 -27881
rect -40833 -29771 -40723 -28013
rect -35307 -29831 -35226 -29703
rect -40901 -30099 -35226 -29967
rect -38771 -31635 -38536 -30099
rect -39141 -31733 -38536 -31635
rect -39041 -31903 -38536 -31733
rect -38661 -31917 -38536 -31903
rect -38704 -32241 -35215 -32109
rect -36976 -33875 -36211 -32241
rect -36844 -34059 -36211 -33875
rect -35370 -34059 -35215 -32241
rect -34330 -34240 -34190 -34176
rect -36513 -34372 -34190 -34240
rect -34409 -36413 -32150 -36281
rect -32673 -38103 -32478 -38102
rect -32673 -38217 -32150 -38103
rect -32566 -38427 -30326 -38295
rect -30436 -40185 -30326 -38427
rect -28100 -40413 -28015 -40401
rect -30340 -40545 -28015 -40413
rect -28210 -42303 -28015 -40545
rect -28236 -42586 -25996 -42454
rect -26106 -44344 -25996 -42586
rect -26393 -44600 -24082 -44468
rect -24263 -46358 -24082 -44600
rect -22901 -46562 -21868 -46528
rect -24191 -46580 -21868 -46562
rect -18070 -46580 -17926 -46528
rect -24191 -46694 -21936 -46580
rect -22455 -48498 -21936 -48384
rect -22087 -48735 -19828 -48603
rect -20351 -50539 -19828 -50425
rect -18002 -50553 -17926 -46580
rect -20244 -50749 -18004 -50617
rect -18126 -52507 -18004 -50749
rect -17973 -53022 -15733 -52888
rect -15843 -54778 -15733 -53022
<< metal1 >>
rect -44835 -13476 -8101 -12068
rect -44839 -23792 -44771 -13476
rect -47011 -23957 -44759 -23792
rect -46898 -24081 -44759 -23957
rect -46774 -24205 -44759 -24081
rect -46650 -24329 -44759 -24205
rect -46526 -24453 -44759 -24329
rect -46402 -24577 -44759 -24453
rect -46278 -24701 -44759 -24577
rect -46154 -24825 -44759 -24701
rect -46030 -24949 -44759 -24825
rect -45906 -25073 -44759 -24949
rect -45782 -25197 -44759 -25073
rect -45658 -25321 -44759 -25197
rect -45534 -25445 -44759 -25321
rect -45410 -25569 -44759 -25445
rect -45286 -25728 -44759 -25569
rect -45286 -25729 -8130 -25728
rect -45072 -25812 -8130 -25729
rect -45072 -25893 -42784 -25812
rect -44959 -26017 -42784 -25893
rect -44835 -26141 -42784 -26017
rect -44711 -26265 -42784 -26141
rect -44587 -26389 -42784 -26265
rect -44463 -26513 -42784 -26389
rect -44339 -26637 -42784 -26513
rect -44215 -26761 -42784 -26637
rect -44091 -26885 -42784 -26761
rect -43967 -27009 -42784 -26885
rect -43843 -27133 -42784 -27009
rect -43719 -27257 -42784 -27133
rect -43595 -27381 -42784 -27257
rect -43471 -27505 -42784 -27381
rect -43347 -27665 -42784 -27505
rect -42952 -28035 -35186 -27892
rect -42839 -28159 -35186 -28035
rect -42715 -28283 -35186 -28159
rect -42591 -28407 -35186 -28283
rect -42467 -28531 -35186 -28407
rect -42343 -28655 -35186 -28531
rect -42219 -28779 -35186 -28655
rect -42095 -28903 -35186 -28779
rect -41971 -29027 -35186 -28903
rect -41847 -29151 -35186 -29027
rect -41723 -29275 -35186 -29151
rect -41599 -29399 -35186 -29275
rect -41475 -29523 -35186 -29399
rect -41351 -29647 -35186 -29523
rect -41227 -29807 -35186 -29647
rect -38782 -31906 -35163 -30042
rect -36756 -34048 -35201 -32120
rect -34766 -34430 -34242 -34402
rect -35215 -35623 -34242 -34430
rect -34766 -36167 -34242 -35623
rect -30335 -36167 -30249 -34430
rect -32415 -38220 -30234 -36292
rect -30904 -40159 -30234 -38220
rect -28582 -42292 -27966 -40488
rect -26500 -44393 -22865 -42465
rect -24658 -46407 -22865 -44479
rect -22444 -48441 -21925 -46782
rect -20363 -50542 -17881 -48678
rect -18497 -52494 -17909 -50692
rect -16182 -52494 -15237 -52449
rect -18497 -52496 -15237 -52494
rect -17962 -52511 -15237 -52496
rect -17962 -52694 -4013 -52511
rect -17962 -52963 -15237 -52694
rect -16182 -54767 -15237 -52963
rect -15387 -55366 -15237 -54767
<< metal2 >>
rect -44125 -14116 -8753 -13916
rect -33258 -14199 -32390 -14116
rect -44125 -25372 -8753 -25172
rect -34569 -28546 -4665 -28346
rect -21335 -29838 -20335 -28546
rect -16462 -29838 -15462 -28546
rect -29773 -39802 -4665 -39602
rect -21950 -40898 -4494 -40698
rect -4686 -51954 -4494 -40898
rect -17281 -52154 -4494 -51954
use M1_PSUB_CDNS_69033583165389  M1_PSUB_CDNS_69033583165389_0
timestamp 1713338890
transform 1 0 -16812 0 1 -53121
box -1037 -45 1037 45
use M1_PSUB_CDNS_69033583165389  M1_PSUB_CDNS_69033583165389_1
timestamp 1713338890
transform 1 0 -19083 0 1 -50850
box -1037 -45 1037 45
use M1_PSUB_CDNS_69033583165389  M1_PSUB_CDNS_69033583165389_2
timestamp 1713338890
transform 1 0 -20926 0 1 -48836
box -1037 -45 1037 45
use M1_PSUB_CDNS_69033583165389  M1_PSUB_CDNS_69033583165389_3
timestamp 1713338890
transform 1 0 -23030 0 1 -46795
box -1037 -45 1037 45
use M1_PSUB_CDNS_69033583165389  M1_PSUB_CDNS_69033583165389_4
timestamp 1713338890
transform 1 0 -25232 0 1 -44701
box -1037 -45 1037 45
use M1_PSUB_CDNS_69033583165389  M1_PSUB_CDNS_69033583165389_5
timestamp 1713338890
transform 1 0 -29179 0 1 -40646
box -1037 -45 1037 45
use M1_PSUB_CDNS_69033583165389  M1_PSUB_CDNS_69033583165389_6
timestamp 1713338890
transform 1 0 -27075 0 1 -42687
box -1037 -45 1037 45
use M1_PSUB_CDNS_69033583165389  M1_PSUB_CDNS_69033583165389_7
timestamp 1713338890
transform 1 0 -31405 0 1 -38528
box -1037 -45 1037 45
use M1_PSUB_CDNS_69033583165389  M1_PSUB_CDNS_69033583165389_8
timestamp 1713338890
transform 1 0 -33248 0 1 -36514
box -1037 -45 1037 45
use M1_PSUB_CDNS_69033583165389  M1_PSUB_CDNS_69033583165389_9
timestamp 1713338890
transform 1 0 -35352 0 1 -34473
box -1037 -45 1037 45
use M1_PSUB_CDNS_69033583165389  M1_PSUB_CDNS_69033583165389_10
timestamp 1713338890
transform 1 0 -37543 0 1 -32342
box -1037 -45 1037 45
use M1_PSUB_CDNS_69033583165389  M1_PSUB_CDNS_69033583165389_11
timestamp 1713338890
transform 1 0 -41802 0 1 -28114
box -1037 -45 1037 45
use M1_PSUB_CDNS_69033583165389  M1_PSUB_CDNS_69033583165389_12
timestamp 1713338890
transform 1 0 -43922 0 1 -25972
box -1037 -45 1037 45
use M1_PSUB_CDNS_69033583165389  M1_PSUB_CDNS_69033583165389_13
timestamp 1713338890
transform 1 0 -45861 0 1 -24036
box -1037 -45 1037 45
use M1_PSUB_CDNS_69033583165389  M1_PSUB_CDNS_69033583165389_14
timestamp 1713338890
transform 1 0 -39740 0 1 -30200
box -1037 -45 1037 45
use M1_PSUB_CDNS_69033583165390  M1_PSUB_CDNS_69033583165390_0
timestamp 1713338890
transform 1 0 -16750 0 1 -53245
box -975 -45 975 45
use M1_PSUB_CDNS_69033583165390  M1_PSUB_CDNS_69033583165390_1
timestamp 1713338890
transform 1 0 -19021 0 1 -50974
box -975 -45 975 45
use M1_PSUB_CDNS_69033583165390  M1_PSUB_CDNS_69033583165390_2
timestamp 1713338890
transform 1 0 -20864 0 1 -48960
box -975 -45 975 45
use M1_PSUB_CDNS_69033583165390  M1_PSUB_CDNS_69033583165390_3
timestamp 1713338890
transform 1 0 -22968 0 1 -46919
box -975 -45 975 45
use M1_PSUB_CDNS_69033583165390  M1_PSUB_CDNS_69033583165390_4
timestamp 1713338890
transform 1 0 -25170 0 1 -44825
box -975 -45 975 45
use M1_PSUB_CDNS_69033583165390  M1_PSUB_CDNS_69033583165390_5
timestamp 1713338890
transform 1 0 -29117 0 1 -40770
box -975 -45 975 45
use M1_PSUB_CDNS_69033583165390  M1_PSUB_CDNS_69033583165390_6
timestamp 1713338890
transform 1 0 -27013 0 1 -42811
box -975 -45 975 45
use M1_PSUB_CDNS_69033583165390  M1_PSUB_CDNS_69033583165390_7
timestamp 1713338890
transform 1 0 -31343 0 1 -38652
box -975 -45 975 45
use M1_PSUB_CDNS_69033583165390  M1_PSUB_CDNS_69033583165390_8
timestamp 1713338890
transform 1 0 -33186 0 1 -36638
box -975 -45 975 45
use M1_PSUB_CDNS_69033583165390  M1_PSUB_CDNS_69033583165390_9
timestamp 1713338890
transform 1 0 -35290 0 1 -34597
box -975 -45 975 45
use M1_PSUB_CDNS_69033583165390  M1_PSUB_CDNS_69033583165390_10
timestamp 1713338890
transform 1 0 -37481 0 1 -32466
box -975 -45 975 45
use M1_PSUB_CDNS_69033583165390  M1_PSUB_CDNS_69033583165390_11
timestamp 1713338890
transform 1 0 -41740 0 1 -28238
box -975 -45 975 45
use M1_PSUB_CDNS_69033583165390  M1_PSUB_CDNS_69033583165390_12
timestamp 1713338890
transform 1 0 -43860 0 1 -26096
box -975 -45 975 45
use M1_PSUB_CDNS_69033583165390  M1_PSUB_CDNS_69033583165390_13
timestamp 1713338890
transform 1 0 -45799 0 1 -24160
box -975 -45 975 45
use M1_PSUB_CDNS_69033583165390  M1_PSUB_CDNS_69033583165390_14
timestamp 1713338890
transform 1 0 -39678 0 1 -30324
box -975 -45 975 45
use M1_PSUB_CDNS_69033583165391  M1_PSUB_CDNS_69033583165391_0
timestamp 1713338890
transform 1 0 -16688 0 1 -53369
box -913 -45 913 45
use M1_PSUB_CDNS_69033583165391  M1_PSUB_CDNS_69033583165391_1
timestamp 1713338890
transform 1 0 -18959 0 1 -51098
box -913 -45 913 45
use M1_PSUB_CDNS_69033583165391  M1_PSUB_CDNS_69033583165391_2
timestamp 1713338890
transform 1 0 -20802 0 1 -49084
box -913 -45 913 45
use M1_PSUB_CDNS_69033583165391  M1_PSUB_CDNS_69033583165391_3
timestamp 1713338890
transform 1 0 -22906 0 1 -47043
box -913 -45 913 45
use M1_PSUB_CDNS_69033583165391  M1_PSUB_CDNS_69033583165391_4
timestamp 1713338890
transform 1 0 -25108 0 1 -44949
box -913 -45 913 45
use M1_PSUB_CDNS_69033583165391  M1_PSUB_CDNS_69033583165391_5
timestamp 1713338890
transform 1 0 -29055 0 1 -40894
box -913 -45 913 45
use M1_PSUB_CDNS_69033583165391  M1_PSUB_CDNS_69033583165391_6
timestamp 1713338890
transform 1 0 -26951 0 1 -42935
box -913 -45 913 45
use M1_PSUB_CDNS_69033583165391  M1_PSUB_CDNS_69033583165391_7
timestamp 1713338890
transform 1 0 -31281 0 1 -38776
box -913 -45 913 45
use M1_PSUB_CDNS_69033583165391  M1_PSUB_CDNS_69033583165391_8
timestamp 1713338890
transform 1 0 -35228 0 1 -34721
box -913 -45 913 45
use M1_PSUB_CDNS_69033583165391  M1_PSUB_CDNS_69033583165391_9
timestamp 1713338890
transform 1 0 -33124 0 1 -36762
box -913 -45 913 45
use M1_PSUB_CDNS_69033583165391  M1_PSUB_CDNS_69033583165391_10
timestamp 1713338890
transform 1 0 -37419 0 1 -32590
box -913 -45 913 45
use M1_PSUB_CDNS_69033583165391  M1_PSUB_CDNS_69033583165391_11
timestamp 1713338890
transform 1 0 -41678 0 1 -28362
box -913 -45 913 45
use M1_PSUB_CDNS_69033583165391  M1_PSUB_CDNS_69033583165391_12
timestamp 1713338890
transform 1 0 -43798 0 1 -26220
box -913 -45 913 45
use M1_PSUB_CDNS_69033583165391  M1_PSUB_CDNS_69033583165391_13
timestamp 1713338890
transform 1 0 -45737 0 1 -24284
box -913 -45 913 45
use M1_PSUB_CDNS_69033583165391  M1_PSUB_CDNS_69033583165391_14
timestamp 1713338890
transform 1 0 -39616 0 1 -30448
box -913 -45 913 45
use M1_PSUB_CDNS_69033583165392  M1_PSUB_CDNS_69033583165392_0
timestamp 1713338890
transform 1 0 -16626 0 1 -53493
box -851 -45 851 45
use M1_PSUB_CDNS_69033583165392  M1_PSUB_CDNS_69033583165392_1
timestamp 1713338890
transform 1 0 -18897 0 1 -51222
box -851 -45 851 45
use M1_PSUB_CDNS_69033583165392  M1_PSUB_CDNS_69033583165392_2
timestamp 1713338890
transform 1 0 -20740 0 1 -49208
box -851 -45 851 45
use M1_PSUB_CDNS_69033583165392  M1_PSUB_CDNS_69033583165392_3
timestamp 1713338890
transform 1 0 -25046 0 1 -45073
box -851 -45 851 45
use M1_PSUB_CDNS_69033583165392  M1_PSUB_CDNS_69033583165392_4
timestamp 1713338890
transform 1 0 -22844 0 1 -47167
box -851 -45 851 45
use M1_PSUB_CDNS_69033583165392  M1_PSUB_CDNS_69033583165392_5
timestamp 1713338890
transform 1 0 -28993 0 1 -41018
box -851 -45 851 45
use M1_PSUB_CDNS_69033583165392  M1_PSUB_CDNS_69033583165392_6
timestamp 1713338890
transform 1 0 -26889 0 1 -43059
box -851 -45 851 45
use M1_PSUB_CDNS_69033583165392  M1_PSUB_CDNS_69033583165392_7
timestamp 1713338890
transform 1 0 -31219 0 1 -38900
box -851 -45 851 45
use M1_PSUB_CDNS_69033583165392  M1_PSUB_CDNS_69033583165392_8
timestamp 1713338890
transform 1 0 -35166 0 1 -34845
box -851 -45 851 45
use M1_PSUB_CDNS_69033583165392  M1_PSUB_CDNS_69033583165392_9
timestamp 1713338890
transform 1 0 -33062 0 1 -36886
box -851 -45 851 45
use M1_PSUB_CDNS_69033583165392  M1_PSUB_CDNS_69033583165392_10
timestamp 1713338890
transform 1 0 -37357 0 1 -32714
box -851 -45 851 45
use M1_PSUB_CDNS_69033583165392  M1_PSUB_CDNS_69033583165392_11
timestamp 1713338890
transform 1 0 -43736 0 1 -26344
box -851 -45 851 45
use M1_PSUB_CDNS_69033583165392  M1_PSUB_CDNS_69033583165392_12
timestamp 1713338890
transform 1 0 -45675 0 1 -24408
box -851 -45 851 45
use M1_PSUB_CDNS_69033583165392  M1_PSUB_CDNS_69033583165392_13
timestamp 1713338890
transform 1 0 -39554 0 1 -30572
box -851 -45 851 45
use M1_PSUB_CDNS_69033583165392  M1_PSUB_CDNS_69033583165392_14
timestamp 1713338890
transform 1 0 -41616 0 1 -28486
box -851 -45 851 45
use M1_PSUB_CDNS_69033583165393  M1_PSUB_CDNS_69033583165393_0
timestamp 1713338890
transform 1 0 -16564 0 1 -53617
box -789 -45 789 45
use M1_PSUB_CDNS_69033583165393  M1_PSUB_CDNS_69033583165393_1
timestamp 1713338890
transform 1 0 -18835 0 1 -51346
box -789 -45 789 45
use M1_PSUB_CDNS_69033583165393  M1_PSUB_CDNS_69033583165393_2
timestamp 1713338890
transform 1 0 -20678 0 1 -49332
box -789 -45 789 45
use M1_PSUB_CDNS_69033583165393  M1_PSUB_CDNS_69033583165393_3
timestamp 1713338890
transform 1 0 -24984 0 1 -45197
box -789 -45 789 45
use M1_PSUB_CDNS_69033583165393  M1_PSUB_CDNS_69033583165393_4
timestamp 1713338890
transform 1 0 -22782 0 1 -47291
box -789 -45 789 45
use M1_PSUB_CDNS_69033583165393  M1_PSUB_CDNS_69033583165393_5
timestamp 1713338890
transform 1 0 -28931 0 1 -41142
box -789 -45 789 45
use M1_PSUB_CDNS_69033583165393  M1_PSUB_CDNS_69033583165393_6
timestamp 1713338890
transform 1 0 -26827 0 1 -43183
box -789 -45 789 45
use M1_PSUB_CDNS_69033583165393  M1_PSUB_CDNS_69033583165393_7
timestamp 1713338890
transform 1 0 -31157 0 1 -39024
box -789 -45 789 45
use M1_PSUB_CDNS_69033583165393  M1_PSUB_CDNS_69033583165393_8
timestamp 1713338890
transform 1 0 -35104 0 1 -34969
box -789 -45 789 45
use M1_PSUB_CDNS_69033583165393  M1_PSUB_CDNS_69033583165393_9
timestamp 1713338890
transform 1 0 -33000 0 1 -37010
box -789 -45 789 45
use M1_PSUB_CDNS_69033583165393  M1_PSUB_CDNS_69033583165393_10
timestamp 1713338890
transform 1 0 -37295 0 1 -32838
box -789 -45 789 45
use M1_PSUB_CDNS_69033583165393  M1_PSUB_CDNS_69033583165393_11
timestamp 1713338890
transform 1 0 -43674 0 1 -26468
box -789 -45 789 45
use M1_PSUB_CDNS_69033583165393  M1_PSUB_CDNS_69033583165393_12
timestamp 1713338890
transform 1 0 -45613 0 1 -24532
box -789 -45 789 45
use M1_PSUB_CDNS_69033583165393  M1_PSUB_CDNS_69033583165393_13
timestamp 1713338890
transform 1 0 -39492 0 1 -30696
box -789 -45 789 45
use M1_PSUB_CDNS_69033583165393  M1_PSUB_CDNS_69033583165393_14
timestamp 1713338890
transform 1 0 -41554 0 1 -28610
box -789 -45 789 45
use M1_PSUB_CDNS_69033583165394  M1_PSUB_CDNS_69033583165394_0
timestamp 1713338890
transform 1 0 -26425 0 1 -12722
box -18335 -665 18335 665
use M1_PSUB_CDNS_69033583165395  M1_PSUB_CDNS_69033583165395_0
timestamp 1713338890
transform 1 0 -16502 0 1 -53741
box -727 -45 727 45
use M1_PSUB_CDNS_69033583165395  M1_PSUB_CDNS_69033583165395_1
timestamp 1713338890
transform 1 0 -18773 0 1 -51470
box -727 -45 727 45
use M1_PSUB_CDNS_69033583165395  M1_PSUB_CDNS_69033583165395_2
timestamp 1713338890
transform 1 0 -20616 0 1 -49456
box -727 -45 727 45
use M1_PSUB_CDNS_69033583165395  M1_PSUB_CDNS_69033583165395_3
timestamp 1713338890
transform 1 0 -24922 0 1 -45321
box -727 -45 727 45
use M1_PSUB_CDNS_69033583165395  M1_PSUB_CDNS_69033583165395_4
timestamp 1713338890
transform 1 0 -22720 0 1 -47415
box -727 -45 727 45
use M1_PSUB_CDNS_69033583165395  M1_PSUB_CDNS_69033583165395_5
timestamp 1713338890
transform 1 0 -28869 0 1 -41266
box -727 -45 727 45
use M1_PSUB_CDNS_69033583165395  M1_PSUB_CDNS_69033583165395_6
timestamp 1713338890
transform 1 0 -26765 0 1 -43307
box -727 -45 727 45
use M1_PSUB_CDNS_69033583165395  M1_PSUB_CDNS_69033583165395_7
timestamp 1713338890
transform 1 0 -31095 0 1 -39148
box -727 -45 727 45
use M1_PSUB_CDNS_69033583165395  M1_PSUB_CDNS_69033583165395_8
timestamp 1713338890
transform 1 0 -32938 0 1 -37134
box -727 -45 727 45
use M1_PSUB_CDNS_69033583165395  M1_PSUB_CDNS_69033583165395_9
timestamp 1713338890
transform 1 0 -35042 0 1 -35093
box -727 -45 727 45
use M1_PSUB_CDNS_69033583165395  M1_PSUB_CDNS_69033583165395_10
timestamp 1713338890
transform 1 0 -37233 0 1 -32962
box -727 -45 727 45
use M1_PSUB_CDNS_69033583165395  M1_PSUB_CDNS_69033583165395_11
timestamp 1713338890
transform 1 0 -43612 0 1 -26592
box -727 -45 727 45
use M1_PSUB_CDNS_69033583165395  M1_PSUB_CDNS_69033583165395_12
timestamp 1713338890
transform 1 0 -45551 0 1 -24656
box -727 -45 727 45
use M1_PSUB_CDNS_69033583165395  M1_PSUB_CDNS_69033583165395_13
timestamp 1713338890
transform 1 0 -39430 0 1 -30820
box -727 -45 727 45
use M1_PSUB_CDNS_69033583165395  M1_PSUB_CDNS_69033583165395_14
timestamp 1713338890
transform 1 0 -41492 0 1 -28734
box -727 -45 727 45
use M1_PSUB_CDNS_69033583165396  M1_PSUB_CDNS_69033583165396_0
timestamp 1713338890
transform 1 0 -16440 0 1 -53865
box -665 -45 665 45
use M1_PSUB_CDNS_69033583165396  M1_PSUB_CDNS_69033583165396_1
timestamp 1713338890
transform 1 0 -18711 0 1 -51594
box -665 -45 665 45
use M1_PSUB_CDNS_69033583165396  M1_PSUB_CDNS_69033583165396_2
timestamp 1713338890
transform 1 0 -20554 0 1 -49580
box -665 -45 665 45
use M1_PSUB_CDNS_69033583165396  M1_PSUB_CDNS_69033583165396_3
timestamp 1713338890
transform 1 0 -24860 0 1 -45445
box -665 -45 665 45
use M1_PSUB_CDNS_69033583165396  M1_PSUB_CDNS_69033583165396_4
timestamp 1713338890
transform 1 0 -22658 0 1 -47539
box -665 -45 665 45
use M1_PSUB_CDNS_69033583165396  M1_PSUB_CDNS_69033583165396_5
timestamp 1713338890
transform 1 0 -28807 0 1 -41390
box -665 -45 665 45
use M1_PSUB_CDNS_69033583165396  M1_PSUB_CDNS_69033583165396_6
timestamp 1713338890
transform 1 0 -26703 0 1 -43431
box -665 -45 665 45
use M1_PSUB_CDNS_69033583165396  M1_PSUB_CDNS_69033583165396_7
timestamp 1713338890
transform 1 0 -31033 0 1 -39272
box -665 -45 665 45
use M1_PSUB_CDNS_69033583165396  M1_PSUB_CDNS_69033583165396_8
timestamp 1713338890
transform 1 0 -32876 0 1 -37258
box -665 -45 665 45
use M1_PSUB_CDNS_69033583165396  M1_PSUB_CDNS_69033583165396_9
timestamp 1713338890
transform 1 0 -34980 0 1 -35217
box -665 -45 665 45
use M1_PSUB_CDNS_69033583165396  M1_PSUB_CDNS_69033583165396_10
timestamp 1713338890
transform 1 0 -37171 0 1 -33086
box -665 -45 665 45
use M1_PSUB_CDNS_69033583165396  M1_PSUB_CDNS_69033583165396_11
timestamp 1713338890
transform 1 0 -43550 0 1 -26716
box -665 -45 665 45
use M1_PSUB_CDNS_69033583165396  M1_PSUB_CDNS_69033583165396_12
timestamp 1713338890
transform 1 0 -45489 0 1 -24780
box -665 -45 665 45
use M1_PSUB_CDNS_69033583165396  M1_PSUB_CDNS_69033583165396_13
timestamp 1713338890
transform 1 0 -39368 0 1 -30944
box -665 -45 665 45
use M1_PSUB_CDNS_69033583165396  M1_PSUB_CDNS_69033583165396_14
timestamp 1713338890
transform 1 0 -41430 0 1 -28858
box -665 -45 665 45
use M1_PSUB_CDNS_69033583165397  M1_PSUB_CDNS_69033583165397_0
timestamp 1713338890
transform 1 0 -16378 0 1 -53989
box -603 -45 603 45
use M1_PSUB_CDNS_69033583165397  M1_PSUB_CDNS_69033583165397_1
timestamp 1713338890
transform 1 0 -18649 0 1 -51718
box -603 -45 603 45
use M1_PSUB_CDNS_69033583165397  M1_PSUB_CDNS_69033583165397_2
timestamp 1713338890
transform 1 0 -20492 0 1 -49704
box -603 -45 603 45
use M1_PSUB_CDNS_69033583165397  M1_PSUB_CDNS_69033583165397_3
timestamp 1713338890
transform 1 0 -22596 0 1 -47663
box -603 -45 603 45
use M1_PSUB_CDNS_69033583165397  M1_PSUB_CDNS_69033583165397_4
timestamp 1713338890
transform 1 0 -24798 0 1 -45569
box -603 -45 603 45
use M1_PSUB_CDNS_69033583165397  M1_PSUB_CDNS_69033583165397_5
timestamp 1713338890
transform 1 0 -28745 0 1 -41514
box -603 -45 603 45
use M1_PSUB_CDNS_69033583165397  M1_PSUB_CDNS_69033583165397_6
timestamp 1713338890
transform 1 0 -26641 0 1 -43555
box -603 -45 603 45
use M1_PSUB_CDNS_69033583165397  M1_PSUB_CDNS_69033583165397_7
timestamp 1713338890
transform 1 0 -30971 0 1 -39396
box -603 -45 603 45
use M1_PSUB_CDNS_69033583165397  M1_PSUB_CDNS_69033583165397_8
timestamp 1713338890
transform 1 0 -32814 0 1 -37382
box -603 -45 603 45
use M1_PSUB_CDNS_69033583165397  M1_PSUB_CDNS_69033583165397_9
timestamp 1713338890
transform 1 0 -34918 0 1 -35341
box -603 -45 603 45
use M1_PSUB_CDNS_69033583165397  M1_PSUB_CDNS_69033583165397_10
timestamp 1713338890
transform 1 0 -37109 0 1 -33210
box -603 -45 603 45
use M1_PSUB_CDNS_69033583165397  M1_PSUB_CDNS_69033583165397_11
timestamp 1713338890
transform 1 0 -43488 0 1 -26840
box -603 -45 603 45
use M1_PSUB_CDNS_69033583165397  M1_PSUB_CDNS_69033583165397_12
timestamp 1713338890
transform 1 0 -45427 0 1 -24904
box -603 -45 603 45
use M1_PSUB_CDNS_69033583165397  M1_PSUB_CDNS_69033583165397_13
timestamp 1713338890
transform 1 0 -39306 0 1 -31068
box -603 -45 603 45
use M1_PSUB_CDNS_69033583165397  M1_PSUB_CDNS_69033583165397_14
timestamp 1713338890
transform 1 0 -41368 0 1 -28982
box -603 -45 603 45
use M1_PSUB_CDNS_69033583165398  M1_PSUB_CDNS_69033583165398_0
timestamp 1713338890
transform 1 0 -16874 0 1 -52997
box -1099 -45 1099 45
use M1_PSUB_CDNS_69033583165398  M1_PSUB_CDNS_69033583165398_1
timestamp 1713338890
transform 1 0 -19145 0 1 -50726
box -1099 -45 1099 45
use M1_PSUB_CDNS_69033583165398  M1_PSUB_CDNS_69033583165398_2
timestamp 1713338890
transform 1 0 -20988 0 1 -48712
box -1099 -45 1099 45
use M1_PSUB_CDNS_69033583165398  M1_PSUB_CDNS_69033583165398_3
timestamp 1713338890
transform 1 0 -23092 0 1 -46671
box -1099 -45 1099 45
use M1_PSUB_CDNS_69033583165398  M1_PSUB_CDNS_69033583165398_4
timestamp 1713338890
transform 1 0 -25294 0 1 -44577
box -1099 -45 1099 45
use M1_PSUB_CDNS_69033583165398  M1_PSUB_CDNS_69033583165398_5
timestamp 1713338890
transform 1 0 -29241 0 1 -40522
box -1099 -45 1099 45
use M1_PSUB_CDNS_69033583165398  M1_PSUB_CDNS_69033583165398_6
timestamp 1713338890
transform 1 0 -27137 0 1 -42563
box -1099 -45 1099 45
use M1_PSUB_CDNS_69033583165398  M1_PSUB_CDNS_69033583165398_7
timestamp 1713338890
transform 1 0 -31467 0 1 -38404
box -1099 -45 1099 45
use M1_PSUB_CDNS_69033583165398  M1_PSUB_CDNS_69033583165398_8
timestamp 1713338890
transform 1 0 -33310 0 1 -36390
box -1099 -45 1099 45
use M1_PSUB_CDNS_69033583165398  M1_PSUB_CDNS_69033583165398_9
timestamp 1713338890
transform 1 0 -35414 0 1 -34349
box -1099 -45 1099 45
use M1_PSUB_CDNS_69033583165398  M1_PSUB_CDNS_69033583165398_10
timestamp 1713338890
transform 1 0 -37605 0 1 -32218
box -1099 -45 1099 45
use M1_PSUB_CDNS_69033583165398  M1_PSUB_CDNS_69033583165398_11
timestamp 1713338890
transform 1 0 -41864 0 1 -27990
box -1099 -45 1099 45
use M1_PSUB_CDNS_69033583165398  M1_PSUB_CDNS_69033583165398_12
timestamp 1713338890
transform 1 0 -43984 0 1 -25848
box -1099 -45 1099 45
use M1_PSUB_CDNS_69033583165398  M1_PSUB_CDNS_69033583165398_13
timestamp 1713338890
transform 1 0 -45923 0 1 -23912
box -1099 -45 1099 45
use M1_PSUB_CDNS_69033583165398  M1_PSUB_CDNS_69033583165398_14
timestamp 1713338890
transform 1 0 -39802 0 1 -30076
box -1099 -45 1099 45
use M1_PSUB_CDNS_69033583165399  M1_PSUB_CDNS_69033583165399_0
timestamp 1713338890
transform 1 0 -16316 0 1 -54113
box -541 -45 541 45
use M1_PSUB_CDNS_69033583165399  M1_PSUB_CDNS_69033583165399_1
timestamp 1713338890
transform 1 0 -18587 0 1 -51842
box -541 -45 541 45
use M1_PSUB_CDNS_69033583165399  M1_PSUB_CDNS_69033583165399_2
timestamp 1713338890
transform 1 0 -20430 0 1 -49828
box -541 -45 541 45
use M1_PSUB_CDNS_69033583165399  M1_PSUB_CDNS_69033583165399_3
timestamp 1713338890
transform 1 0 -22534 0 1 -47787
box -541 -45 541 45
use M1_PSUB_CDNS_69033583165399  M1_PSUB_CDNS_69033583165399_4
timestamp 1713338890
transform 1 0 -24736 0 1 -45693
box -541 -45 541 45
use M1_PSUB_CDNS_69033583165399  M1_PSUB_CDNS_69033583165399_5
timestamp 1713338890
transform 1 0 -26579 0 1 -43679
box -541 -45 541 45
use M1_PSUB_CDNS_69033583165399  M1_PSUB_CDNS_69033583165399_6
timestamp 1713338890
transform 1 0 -28683 0 1 -41638
box -541 -45 541 45
use M1_PSUB_CDNS_69033583165399  M1_PSUB_CDNS_69033583165399_7
timestamp 1713338890
transform 1 0 -30909 0 1 -39520
box -541 -45 541 45
use M1_PSUB_CDNS_69033583165399  M1_PSUB_CDNS_69033583165399_8
timestamp 1713338890
transform 1 0 -32752 0 1 -37506
box -541 -45 541 45
use M1_PSUB_CDNS_69033583165399  M1_PSUB_CDNS_69033583165399_9
timestamp 1713338890
transform 1 0 -34856 0 1 -35465
box -541 -45 541 45
use M1_PSUB_CDNS_69033583165399  M1_PSUB_CDNS_69033583165399_10
timestamp 1713338890
transform 1 0 -37047 0 1 -33334
box -541 -45 541 45
use M1_PSUB_CDNS_69033583165399  M1_PSUB_CDNS_69033583165399_11
timestamp 1713338890
transform 1 0 -43426 0 1 -26964
box -541 -45 541 45
use M1_PSUB_CDNS_69033583165399  M1_PSUB_CDNS_69033583165399_12
timestamp 1713338890
transform 1 0 -45365 0 1 -25028
box -541 -45 541 45
use M1_PSUB_CDNS_69033583165399  M1_PSUB_CDNS_69033583165399_13
timestamp 1713338890
transform 1 0 -39244 0 1 -31192
box -541 -45 541 45
use M1_PSUB_CDNS_69033583165399  M1_PSUB_CDNS_69033583165399_14
timestamp 1713338890
transform 1 0 -41306 0 1 -29106
box -541 -45 541 45
use M1_PSUB_CDNS_69033583165400  M1_PSUB_CDNS_69033583165400_0
timestamp 1713338890
transform 1 0 -16254 0 1 -54237
box -479 -45 479 45
use M1_PSUB_CDNS_69033583165400  M1_PSUB_CDNS_69033583165400_1
timestamp 1713338890
transform 1 0 -18525 0 1 -51966
box -479 -45 479 45
use M1_PSUB_CDNS_69033583165400  M1_PSUB_CDNS_69033583165400_2
timestamp 1713338890
transform 1 0 -20368 0 1 -49952
box -479 -45 479 45
use M1_PSUB_CDNS_69033583165400  M1_PSUB_CDNS_69033583165400_3
timestamp 1713338890
transform 1 0 -22472 0 1 -47911
box -479 -45 479 45
use M1_PSUB_CDNS_69033583165400  M1_PSUB_CDNS_69033583165400_4
timestamp 1713338890
transform 1 0 -24674 0 1 -45817
box -479 -45 479 45
use M1_PSUB_CDNS_69033583165400  M1_PSUB_CDNS_69033583165400_5
timestamp 1713338890
transform 1 0 -26517 0 1 -43803
box -479 -45 479 45
use M1_PSUB_CDNS_69033583165400  M1_PSUB_CDNS_69033583165400_6
timestamp 1713338890
transform 1 0 -28621 0 1 -41762
box -479 -45 479 45
use M1_PSUB_CDNS_69033583165400  M1_PSUB_CDNS_69033583165400_7
timestamp 1713338890
transform 1 0 -30847 0 1 -39644
box -479 -45 479 45
use M1_PSUB_CDNS_69033583165400  M1_PSUB_CDNS_69033583165400_8
timestamp 1713338890
transform 1 0 -32690 0 1 -37630
box -479 -45 479 45
use M1_PSUB_CDNS_69033583165400  M1_PSUB_CDNS_69033583165400_9
timestamp 1713338890
transform 1 0 -34794 0 1 -35589
box -479 -45 479 45
use M1_PSUB_CDNS_69033583165400  M1_PSUB_CDNS_69033583165400_10
timestamp 1713338890
transform 1 0 -36985 0 1 -33458
box -479 -45 479 45
use M1_PSUB_CDNS_69033583165400  M1_PSUB_CDNS_69033583165400_11
timestamp 1713338890
transform 1 0 -43364 0 1 -27088
box -479 -45 479 45
use M1_PSUB_CDNS_69033583165400  M1_PSUB_CDNS_69033583165400_12
timestamp 1713338890
transform 1 0 -45303 0 1 -25152
box -479 -45 479 45
use M1_PSUB_CDNS_69033583165400  M1_PSUB_CDNS_69033583165400_13
timestamp 1713338890
transform 1 0 -39182 0 1 -31316
box -479 -45 479 45
use M1_PSUB_CDNS_69033583165400  M1_PSUB_CDNS_69033583165400_14
timestamp 1713338890
transform 1 0 -41244 0 1 -29230
box -479 -45 479 45
use M1_PSUB_CDNS_69033583165401  M1_PSUB_CDNS_69033583165401_0
timestamp 1713338890
transform 1 0 -16192 0 1 -54361
box -417 -45 417 45
use M1_PSUB_CDNS_69033583165401  M1_PSUB_CDNS_69033583165401_1
timestamp 1713338890
transform 1 0 -18463 0 1 -52090
box -417 -45 417 45
use M1_PSUB_CDNS_69033583165401  M1_PSUB_CDNS_69033583165401_2
timestamp 1713338890
transform 1 0 -20306 0 1 -50076
box -417 -45 417 45
use M1_PSUB_CDNS_69033583165401  M1_PSUB_CDNS_69033583165401_3
timestamp 1713338890
transform 1 0 -22410 0 1 -48035
box -417 -45 417 45
use M1_PSUB_CDNS_69033583165401  M1_PSUB_CDNS_69033583165401_4
timestamp 1713338890
transform 1 0 -24612 0 1 -45941
box -417 -45 417 45
use M1_PSUB_CDNS_69033583165401  M1_PSUB_CDNS_69033583165401_5
timestamp 1713338890
transform 1 0 -26455 0 1 -43927
box -417 -45 417 45
use M1_PSUB_CDNS_69033583165401  M1_PSUB_CDNS_69033583165401_6
timestamp 1713338890
transform 1 0 -28559 0 1 -41886
box -417 -45 417 45
use M1_PSUB_CDNS_69033583165401  M1_PSUB_CDNS_69033583165401_7
timestamp 1713338890
transform 1 0 -30785 0 1 -39768
box -417 -45 417 45
use M1_PSUB_CDNS_69033583165401  M1_PSUB_CDNS_69033583165401_8
timestamp 1713338890
transform 1 0 -32628 0 1 -37754
box -417 -45 417 45
use M1_PSUB_CDNS_69033583165401  M1_PSUB_CDNS_69033583165401_9
timestamp 1713338890
transform 1 0 -34732 0 1 -35713
box -417 -45 417 45
use M1_PSUB_CDNS_69033583165401  M1_PSUB_CDNS_69033583165401_10
timestamp 1713338890
transform 1 0 -36923 0 1 -33582
box -417 -45 417 45
use M1_PSUB_CDNS_69033583165401  M1_PSUB_CDNS_69033583165401_11
timestamp 1713338890
transform 1 0 -43302 0 1 -27212
box -417 -45 417 45
use M1_PSUB_CDNS_69033583165401  M1_PSUB_CDNS_69033583165401_12
timestamp 1713338890
transform 1 0 -45241 0 1 -25276
box -417 -45 417 45
use M1_PSUB_CDNS_69033583165401  M1_PSUB_CDNS_69033583165401_13
timestamp 1713338890
transform 1 0 -39120 0 1 -31440
box -417 -45 417 45
use M1_PSUB_CDNS_69033583165401  M1_PSUB_CDNS_69033583165401_14
timestamp 1713338890
transform 1 0 -41182 0 1 -29354
box -417 -45 417 45
use M1_PSUB_CDNS_69033583165402  M1_PSUB_CDNS_69033583165402_0
timestamp 1713338890
transform 1 0 -16130 0 1 -54485
box -355 -45 355 45
use M1_PSUB_CDNS_69033583165402  M1_PSUB_CDNS_69033583165402_1
timestamp 1713338890
transform 1 0 -18401 0 1 -52214
box -355 -45 355 45
use M1_PSUB_CDNS_69033583165402  M1_PSUB_CDNS_69033583165402_2
timestamp 1713338890
transform 1 0 -20244 0 1 -50200
box -355 -45 355 45
use M1_PSUB_CDNS_69033583165402  M1_PSUB_CDNS_69033583165402_3
timestamp 1713338890
transform 1 0 -22348 0 1 -48159
box -355 -45 355 45
use M1_PSUB_CDNS_69033583165402  M1_PSUB_CDNS_69033583165402_4
timestamp 1713338890
transform 1 0 -24550 0 1 -46065
box -355 -45 355 45
use M1_PSUB_CDNS_69033583165402  M1_PSUB_CDNS_69033583165402_5
timestamp 1713338890
transform 1 0 -26393 0 1 -44051
box -355 -45 355 45
use M1_PSUB_CDNS_69033583165402  M1_PSUB_CDNS_69033583165402_6
timestamp 1713338890
transform 1 0 -28497 0 1 -42010
box -355 -45 355 45
use M1_PSUB_CDNS_69033583165402  M1_PSUB_CDNS_69033583165402_7
timestamp 1713338890
transform 1 0 -30723 0 1 -39892
box -355 -45 355 45
use M1_PSUB_CDNS_69033583165402  M1_PSUB_CDNS_69033583165402_8
timestamp 1713338890
transform 1 0 -32566 0 1 -37878
box -355 -45 355 45
use M1_PSUB_CDNS_69033583165402  M1_PSUB_CDNS_69033583165402_9
timestamp 1713338890
transform 1 0 -34670 0 1 -35837
box -355 -45 355 45
use M1_PSUB_CDNS_69033583165402  M1_PSUB_CDNS_69033583165402_10
timestamp 1713338890
transform 1 0 -36861 0 1 -33706
box -355 -45 355 45
use M1_PSUB_CDNS_69033583165402  M1_PSUB_CDNS_69033583165402_11
timestamp 1713338890
transform 1 0 -43240 0 1 -27336
box -355 -45 355 45
use M1_PSUB_CDNS_69033583165402  M1_PSUB_CDNS_69033583165402_12
timestamp 1713338890
transform 1 0 -45179 0 1 -25400
box -355 -45 355 45
use M1_PSUB_CDNS_69033583165402  M1_PSUB_CDNS_69033583165402_13
timestamp 1713338890
transform 1 0 -39058 0 1 -31564
box -355 -45 355 45
use M1_PSUB_CDNS_69033583165402  M1_PSUB_CDNS_69033583165402_14
timestamp 1713338890
transform 1 0 -41120 0 1 -29478
box -355 -45 355 45
use M1_PSUB_CDNS_69033583165403  M1_PSUB_CDNS_69033583165403_0
timestamp 1713338890
transform 1 0 -16068 0 1 -54609
box -293 -45 293 45
use M1_PSUB_CDNS_69033583165403  M1_PSUB_CDNS_69033583165403_1
timestamp 1713338890
transform 1 0 -18339 0 1 -52338
box -293 -45 293 45
use M1_PSUB_CDNS_69033583165403  M1_PSUB_CDNS_69033583165403_2
timestamp 1713338890
transform 1 0 -20182 0 1 -50324
box -293 -45 293 45
use M1_PSUB_CDNS_69033583165403  M1_PSUB_CDNS_69033583165403_3
timestamp 1713338890
transform 1 0 -22286 0 1 -48283
box -293 -45 293 45
use M1_PSUB_CDNS_69033583165403  M1_PSUB_CDNS_69033583165403_4
timestamp 1713338890
transform 1 0 -24488 0 1 -46189
box -293 -45 293 45
use M1_PSUB_CDNS_69033583165403  M1_PSUB_CDNS_69033583165403_5
timestamp 1713338890
transform 1 0 -26331 0 1 -44175
box -293 -45 293 45
use M1_PSUB_CDNS_69033583165403  M1_PSUB_CDNS_69033583165403_6
timestamp 1713338890
transform 1 0 -28435 0 1 -42134
box -293 -45 293 45
use M1_PSUB_CDNS_69033583165403  M1_PSUB_CDNS_69033583165403_7
timestamp 1713338890
transform 1 0 -30661 0 1 -40016
box -293 -45 293 45
use M1_PSUB_CDNS_69033583165403  M1_PSUB_CDNS_69033583165403_8
timestamp 1713338890
transform 1 0 -32504 0 1 -38002
box -293 -45 293 45
use M1_PSUB_CDNS_69033583165403  M1_PSUB_CDNS_69033583165403_9
timestamp 1713338890
transform 1 0 -34608 0 1 -35961
box -293 -45 293 45
use M1_PSUB_CDNS_69033583165403  M1_PSUB_CDNS_69033583165403_10
timestamp 1713338890
transform 1 0 -36799 0 1 -33830
box -293 -45 293 45
use M1_PSUB_CDNS_69033583165403  M1_PSUB_CDNS_69033583165403_11
timestamp 1713338890
transform 1 0 -43178 0 1 -27460
box -293 -45 293 45
use M1_PSUB_CDNS_69033583165403  M1_PSUB_CDNS_69033583165403_12
timestamp 1713338890
transform 1 0 -45117 0 1 -25524
box -293 -45 293 45
use M1_PSUB_CDNS_69033583165403  M1_PSUB_CDNS_69033583165403_13
timestamp 1713338890
transform 1 0 -38996 0 1 -31688
box -293 -45 293 45
use M1_PSUB_CDNS_69033583165403  M1_PSUB_CDNS_69033583165403_14
timestamp 1713338890
transform 1 0 -41058 0 1 -29602
box -293 -45 293 45
use M1_PSUB_CDNS_69033583165404  M1_PSUB_CDNS_69033583165404_0
timestamp 1713338890
transform 1 0 -25462 0 1 -26776
box -17343 -975 17343 975
use M1_PSUB_CDNS_69033583165405  M1_PSUB_CDNS_69033583165405_0
timestamp 1713338890
transform 1 0 -19969 0 1 -47525
box -1967 -975 1967 975
use M1_PSUB_CDNS_69033583165405  M1_PSUB_CDNS_69033583165405_1
timestamp 1713338890
transform 1 0 -32291 0 1 -35203
box -1967 -975 1967 975
use M1_PSUB_CDNS_69033583165406  M1_PSUB_CDNS_69033583165406_0
timestamp 1713338890
transform 1 0 -18915 0 1 -49578
box -913 -975 913 975
use M1_PSUB_CDNS_69033583165406  M1_PSUB_CDNS_69033583165406_1
timestamp 1713338890
transform 1 0 -31237 0 1 -37256
box -913 -975 913 975
use M1_PSUB_CDNS_69033583165435  M1_PSUB_CDNS_69033583165435_0
timestamp 1713338890
transform 1 0 -45923 0 1 -17930
box -1099 -5873 1099 5873
use M1_PSUB_CDNS_69033583165442  M1_PSUB_CDNS_69033583165442_0
timestamp 1713338890
transform 1 0 -16006 0 1 -54733
box -231 -45 231 45
use M1_PSUB_CDNS_69033583165442  M1_PSUB_CDNS_69033583165442_1
timestamp 1713338890
transform 1 0 -18277 0 1 -52462
box -231 -45 231 45
use M1_PSUB_CDNS_69033583165442  M1_PSUB_CDNS_69033583165442_2
timestamp 1713338890
transform 1 0 -20120 0 1 -50448
box -231 -45 231 45
use M1_PSUB_CDNS_69033583165442  M1_PSUB_CDNS_69033583165442_3
timestamp 1713338890
transform 1 0 -22224 0 1 -48407
box -231 -45 231 45
use M1_PSUB_CDNS_69033583165442  M1_PSUB_CDNS_69033583165442_4
timestamp 1713338890
transform 1 0 -24426 0 1 -46313
box -231 -45 231 45
use M1_PSUB_CDNS_69033583165442  M1_PSUB_CDNS_69033583165442_5
timestamp 1713338890
transform 1 0 -26269 0 1 -44299
box -231 -45 231 45
use M1_PSUB_CDNS_69033583165442  M1_PSUB_CDNS_69033583165442_6
timestamp 1713338890
transform 1 0 -28373 0 1 -42258
box -231 -45 231 45
use M1_PSUB_CDNS_69033583165442  M1_PSUB_CDNS_69033583165442_7
timestamp 1713338890
transform 1 0 -30599 0 1 -40140
box -231 -45 231 45
use M1_PSUB_CDNS_69033583165442  M1_PSUB_CDNS_69033583165442_8
timestamp 1713338890
transform 1 0 -32442 0 1 -38126
box -231 -45 231 45
use M1_PSUB_CDNS_69033583165442  M1_PSUB_CDNS_69033583165442_9
timestamp 1713338890
transform 1 0 -34546 0 1 -36085
box -231 -45 231 45
use M1_PSUB_CDNS_69033583165442  M1_PSUB_CDNS_69033583165442_10
timestamp 1713338890
transform 1 0 -43116 0 1 -27584
box -231 -45 231 45
use M1_PSUB_CDNS_69033583165442  M1_PSUB_CDNS_69033583165442_11
timestamp 1713338890
transform 1 0 -45055 0 1 -25648
box -231 -45 231 45
use M1_PSUB_CDNS_69033583165442  M1_PSUB_CDNS_69033583165442_12
timestamp 1713338890
transform 1 0 -40996 0 1 -29726
box -231 -45 231 45
use M1_PSUB_CDNS_69033583165451  M1_PSUB_CDNS_69033583165451_0
timestamp 1713338890
transform 1 0 -25490 0 1 -41376
box -2525 -975 2525 975
use M1_PSUB_CDNS_69033583165459  M1_PSUB_CDNS_69033583165459_0
timestamp 1713338890
transform 1 0 -37939 0 1 -28856
box -2649 -975 2649 975
use M1_PSUB_CDNS_69033583165460  M1_PSUB_CDNS_69033583165460_0
timestamp 1713338890
transform 1 0 -36947 0 1 -30942
box -1657 -975 1657 975
use M1_PSUB_CDNS_69033583165462  M1_PSUB_CDNS_69033583165462_0
timestamp 1713338890
transform 1 0 -23541 0 1 -45443
box -541 -975 541 975
use M1_PSUB_CDNS_69033583165462  M1_PSUB_CDNS_69033583165462_1
timestamp 1713338890
transform 1 0 -35842 0 1 -33084
box -541 -975 541 975
use M1_PSUB_CDNS_69033583165463  M1_PSUB_CDNS_69033583165463_0
timestamp 1713338890
transform 1 0 -36675 0 1 -33954
box -169 -45 169 45
use M1_PSUB_CDNS_69033583165463  M1_PSUB_CDNS_69033583165463_1
timestamp 1713338890
transform 1 0 -38872 0 1 -31812
box -169 -45 169 45
use M1_PSUB_CDNS_69033583165465  M1_PSUB_CDNS_69033583165465_0
timestamp 1713338890
transform 1 0 -24436 0 1 -43429
box -1471 -975 1471 975
use M1_PSUB_CDNS_69033583165479  M1_PSUB_CDNS_69033583165479_0
timestamp 1713338890
transform 1 0 -9468 0 1 -54092
box -5811 -1285 5811 1285
use M2_M1_CDNS_69033583165409  M2_M1_CDNS_69033583165409_0
timestamp 1713338890
transform 1 0 -12921 0 1 -36139
box -434 -1622 434 1622
use M2_M1_CDNS_69033583165409  M2_M1_CDNS_69033583165409_1
timestamp 1713338890
transform 1 0 -8078 0 1 -36503
box -434 -1622 434 1622
use M2_M1_CDNS_69033583165409  M2_M1_CDNS_69033583165409_2
timestamp 1713338890
transform 1 0 -18419 0 1 -30678
box -434 -1622 434 1622
use M2_M1_CDNS_69033583165409  M2_M1_CDNS_69033583165409_3
timestamp 1713338890
transform 1 0 -12921 0 1 -31665
box -434 -1622 434 1622
use M2_M1_CDNS_69033583165409  M2_M1_CDNS_69033583165409_4
timestamp 1713338890
transform 1 0 -8041 0 1 -31997
box -434 -1622 434 1622
use M2_M1_CDNS_69033583165410  M2_M1_CDNS_69033583165410_0
timestamp 1713338890
transform 1 0 -19727 0 1 -47419
box -1178 -570 1178 570
use M2_M1_CDNS_69033583165410  M2_M1_CDNS_69033583165410_1
timestamp 1713338890
transform 1 0 -23781 0 1 -43365
box -1178 -570 1178 570
use M2_M1_CDNS_69033583165410  M2_M1_CDNS_69033583165410_2
timestamp 1713338890
transform 1 0 -25879 0 1 -41267
box -1178 -570 1178 570
use M2_M1_CDNS_69033583165411  M2_M1_CDNS_69033583165411_0
timestamp 1713338890
transform 1 0 -9214 0 1 -52063
box -4522 -38 4522 38
use M2_M1_CDNS_69033583165411  M2_M1_CDNS_69033583165411_1
timestamp 1713338890
transform 1 0 -9214 0 1 -40765
box -4522 -38 4522 38
use M2_M1_CDNS_69033583165411  M2_M1_CDNS_69033583165411_2
timestamp 1713338890
transform 1 0 -19546 0 1 -39718
box -4522 -38 4522 38
use M2_M1_CDNS_69033583165411  M2_M1_CDNS_69033583165411_3
timestamp 1713338890
transform 1 0 -9214 0 1 -39718
box -4522 -38 4522 38
use M2_M1_CDNS_69033583165411  M2_M1_CDNS_69033583165411_4
timestamp 1713338890
transform 1 0 -34040 0 1 -25281
box -4522 -38 4522 38
use M2_M1_CDNS_69033583165411  M2_M1_CDNS_69033583165411_5
timestamp 1713338890
transform 1 0 -29996 0 1 -28425
box -4522 -38 4522 38
use M2_M1_CDNS_69033583165411  M2_M1_CDNS_69033583165411_6
timestamp 1713338890
transform 1 0 -19546 0 1 -28425
box -4522 -38 4522 38
use M2_M1_CDNS_69033583165411  M2_M1_CDNS_69033583165411_7
timestamp 1713338890
transform 1 0 -23658 0 1 -25281
box -4522 -38 4522 38
use M2_M1_CDNS_69033583165411  M2_M1_CDNS_69033583165411_8
timestamp 1713338890
transform 1 0 -13326 0 1 -25281
box -4522 -38 4522 38
use M2_M1_CDNS_69033583165411  M2_M1_CDNS_69033583165411_9
timestamp 1713338890
transform 1 0 -9214 0 1 -28425
box -4522 -38 4522 38
use M2_M1_CDNS_69033583165411  M2_M1_CDNS_69033583165411_10
timestamp 1713338890
transform 1 0 -13326 0 1 -13985
box -4522 -38 4522 38
use M2_M1_CDNS_69033583165411  M2_M1_CDNS_69033583165411_11
timestamp 1713338890
transform 1 0 -34040 0 1 -13985
box -4522 -38 4522 38
use M2_M1_CDNS_69033583165411  M2_M1_CDNS_69033583165411_12
timestamp 1713338890
transform 1 0 -23658 0 1 -13985
box -4522 -38 4522 38
use M2_M1_CDNS_69033583165412  M2_M1_CDNS_69033583165412_0
timestamp 1713338890
transform 1 0 -18490 0 1 -40765
box -3002 -38 3002 38
use M2_M1_CDNS_69033583165417  M2_M1_CDNS_69033583165417_0
timestamp 1713338890
transform 1 0 9643 0 1 -10945
box -162 -596 162 596
use M2_M1_CDNS_69033583165417  M2_M1_CDNS_69033583165417_1
timestamp 1713338890
transform 1 0 9635 0 1 -7796
box -162 -596 162 596
use M2_M1_CDNS_69033583165417  M2_M1_CDNS_69033583165417_2
timestamp 1713338890
transform 1 0 9655 0 1 -2992
box -162 -596 162 596
use M2_M1_CDNS_69033583165419  M2_M1_CDNS_69033583165419_0
timestamp 1713338890
transform 1 0 -17015 0 1 -18078
box -494 -1102 494 1102
use M2_M1_CDNS_69033583165421  M2_M1_CDNS_69033583165421_0
timestamp 1713338890
transform 1 0 8277 0 1 -1404
box -368 -632 368 632
use M2_M1_CDNS_69033583165422  M2_M1_CDNS_69033583165422_0
timestamp 1713338890
transform 1 0 542 0 1 38
box -596 -38 596 38
use M2_M1_CDNS_69033583165422  M2_M1_CDNS_69033583165422_1
timestamp 1713338890
transform 1 0 5317 0 1 38
box -596 -38 596 38
use M2_M1_CDNS_69033583165423  M2_M1_CDNS_69033583165423_0
timestamp 1713338890
transform 1 0 5824 0 1 -9409
box -410 -658 410 658
use M2_M1_CDNS_69033583165424  M2_M1_CDNS_69033583165424_0
timestamp 1713338890
transform 1 0 6950 0 1 -377
box -658 -38 658 38
use M2_M1_CDNS_69033583165425  M2_M1_CDNS_69033583165425_0
timestamp 1713338890
transform 1 0 8869 0 1 38
box -968 -38 968 38
use M2_M1_CDNS_69033583165431  M2_M1_CDNS_69033583165431_0
timestamp 1713338890
transform 1 0 -32824 0 1 -16019
box -434 -1820 434 1820
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_0
timestamp 1713338890
transform 1 0 -27597 0 1 -39718
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_1
timestamp 1713338890
transform 1 0 -32235 0 1 -35063
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_2
timestamp 1713338890
transform 1 0 -32387 0 1 -34911
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_3
timestamp 1713338890
transform 1 0 -32539 0 1 -34759
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_4
timestamp 1713338890
transform 1 0 -32691 0 1 -34607
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_5
timestamp 1713338890
transform 1 0 -32843 0 1 -34455
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_6
timestamp 1713338890
transform 1 0 -32995 0 1 -34303
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_7
timestamp 1713338890
transform 1 0 -33147 0 1 -34151
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_8
timestamp 1713338890
transform 1 0 -33299 0 1 -33999
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_9
timestamp 1713338890
transform 1 0 -32083 0 1 -35215
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_10
timestamp 1713338890
transform 1 0 -31931 0 1 -35367
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_11
timestamp 1713338890
transform 1 0 -31779 0 1 -35519
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_12
timestamp 1713338890
transform 1 0 -33451 0 1 -33847
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_13
timestamp 1713338890
transform 1 0 -40754 0 1 -26544
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_14
timestamp 1713338890
transform 1 0 -40906 0 1 -26392
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_15
timestamp 1713338890
transform 1 0 -41058 0 1 -26240
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_16
timestamp 1713338890
transform 1 0 -41210 0 1 -26088
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_17
timestamp 1713338890
transform 1 0 -41362 0 1 -25936
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_18
timestamp 1713338890
transform 1 0 -41514 0 1 -25784
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_19
timestamp 1713338890
transform 1 0 -41666 0 1 -25632
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_20
timestamp 1713338890
transform 1 0 -37602 0 1 -29696
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_21
timestamp 1713338890
transform 1 0 -37754 0 1 -29544
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_22
timestamp 1713338890
transform 1 0 -37906 0 1 -29392
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_23
timestamp 1713338890
transform 1 0 -38058 0 1 -29240
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_24
timestamp 1713338890
transform 1 0 -38210 0 1 -29088
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_25
timestamp 1713338890
transform 1 0 -38362 0 1 -28936
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_26
timestamp 1713338890
transform 1 0 -38514 0 1 -28784
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_27
timestamp 1713338890
transform 1 0 -38666 0 1 -28632
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_28
timestamp 1713338890
transform 1 0 -38818 0 1 -28480
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_29
timestamp 1713338890
transform 1 0 -38970 0 1 -28328
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_30
timestamp 1713338890
transform 1 0 -39122 0 1 -28176
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_31
timestamp 1713338890
transform 1 0 -39274 0 1 -28024
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_32
timestamp 1713338890
transform 1 0 -39690 0 1 -27608
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_33
timestamp 1713338890
transform 1 0 -39842 0 1 -27456
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_34
timestamp 1713338890
transform 1 0 -39994 0 1 -27304
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_35
timestamp 1713338890
transform 1 0 -40146 0 1 -27152
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_36
timestamp 1713338890
transform 1 0 -40298 0 1 -27000
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_37
timestamp 1713338890
transform 1 0 -40450 0 1 -26848
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_38
timestamp 1713338890
transform 1 0 -40602 0 1 -26696
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_39
timestamp 1713338890
transform 1 0 -36130 0 1 -26544
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_40
timestamp 1713338890
transform 1 0 -36282 0 1 -26392
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_41
timestamp 1713338890
transform 1 0 -36434 0 1 -26240
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_42
timestamp 1713338890
transform 1 0 -36586 0 1 -26088
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_43
timestamp 1713338890
transform 1 0 -36738 0 1 -25936
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_44
timestamp 1713338890
transform 1 0 -36890 0 1 -25784
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_45
timestamp 1713338890
transform 1 0 -37042 0 1 -25632
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_46
timestamp 1713338890
transform 1 0 -35066 0 1 -27608
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_47
timestamp 1713338890
transform 1 0 -30567 0 1 -27608
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_48
timestamp 1713338890
transform 1 0 -35218 0 1 -27456
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_49
timestamp 1713338890
transform 1 0 -30719 0 1 -27456
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_50
timestamp 1713338890
transform 1 0 -35370 0 1 -27304
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_51
timestamp 1713338890
transform 1 0 -30871 0 1 -27304
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_52
timestamp 1713338890
transform 1 0 -31023 0 1 -27152
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_53
timestamp 1713338890
transform 1 0 -35522 0 1 -27152
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_54
timestamp 1713338890
transform 1 0 -31175 0 1 -27000
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_55
timestamp 1713338890
transform 1 0 -35674 0 1 -27000
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_56
timestamp 1713338890
transform 1 0 -31327 0 1 -26848
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_57
timestamp 1713338890
transform 1 0 -35826 0 1 -26848
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_58
timestamp 1713338890
transform 1 0 -31479 0 1 -26696
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_59
timestamp 1713338890
transform 1 0 -35978 0 1 -26696
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_60
timestamp 1713338890
transform 1 0 -32087 0 1 -26088
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_61
timestamp 1713338890
transform 1 0 -31935 0 1 -26240
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_62
timestamp 1713338890
transform 1 0 -31783 0 1 -26392
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_63
timestamp 1713338890
transform 1 0 -31631 0 1 -26544
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_64
timestamp 1713338890
transform 1 0 -32391 0 1 -25784
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_65
timestamp 1713338890
transform 1 0 -32543 0 1 -25632
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165432  M2_M1_CDNS_69033583165432_66
timestamp 1713338890
transform 1 0 -32239 0 1 -25936
box -1862 -38 1862 38
use M2_M1_CDNS_69033583165433  M2_M1_CDNS_69033583165433_0
timestamp 1713338890
transform 1 0 -32827 0 1 -21936
box -494 -266 494 266
use M2_M1_CDNS_69033583165433  M2_M1_CDNS_69033583165433_1
timestamp 1713338890
transform 1 0 -32918 0 1 -19655
box -494 -266 494 266
use M2_M1_CDNS_69033583165434  M2_M1_CDNS_69033583165434_0
timestamp 1713338890
transform 1 0 -45402 0 1 -17451
box -1026 -5282 1026 5282
use M2_M1_CDNS_69033583165436  M2_M1_CDNS_69033583165436_0
timestamp 1713338890
transform 1 0 -34669 0 1 -12857
box -632 -632 632 632
use M2_M1_CDNS_69033583165438  M2_M1_CDNS_69033583165438_0
timestamp 1713338890
transform 1 0 -41853 0 1 -12857
box -1358 -632 1358 632
use M2_M1_CDNS_69033583165438  M2_M1_CDNS_69033583165438_1
timestamp 1713338890
transform 1 0 -38682 0 1 -12857
box -1358 -632 1358 632
use M2_M1_CDNS_69033583165439  M2_M1_CDNS_69033583165439_0
timestamp 1713338890
transform 1 0 -41969 0 1 -25281
box -2090 -38 2090 38
use M2_M1_CDNS_69033583165439  M2_M1_CDNS_69033583165439_1
timestamp 1713338890
transform 1 0 -41969 0 1 -13985
box -2090 -38 2090 38
use M2_M1_CDNS_69033583165441  M2_M1_CDNS_69033583165441_0
timestamp 1713338890
transform 1 0 -41853 0 1 -19655
box -1406 -266 1406 266
use M2_M1_CDNS_69033583165441  M2_M1_CDNS_69033583165441_1
timestamp 1713338890
transform 1 0 -38433 0 1 -19655
box -1406 -266 1406 266
use M2_M1_CDNS_69033583165443  M2_M1_CDNS_69033583165443_0
timestamp 1713338890
transform 1 0 -24918 0 1 -27608
box -874 -38 874 38
use M2_M1_CDNS_69033583165443  M2_M1_CDNS_69033583165443_1
timestamp 1713338890
transform 1 0 -25070 0 1 -27456
box -874 -38 874 38
use M2_M1_CDNS_69033583165443  M2_M1_CDNS_69033583165443_2
timestamp 1713338890
transform 1 0 -25222 0 1 -27304
box -874 -38 874 38
use M2_M1_CDNS_69033583165443  M2_M1_CDNS_69033583165443_3
timestamp 1713338890
transform 1 0 -25374 0 1 -27152
box -874 -38 874 38
use M2_M1_CDNS_69033583165443  M2_M1_CDNS_69033583165443_4
timestamp 1713338890
transform 1 0 -25526 0 1 -27000
box -874 -38 874 38
use M2_M1_CDNS_69033583165443  M2_M1_CDNS_69033583165443_5
timestamp 1713338890
transform 1 0 -25678 0 1 -26848
box -874 -38 874 38
use M2_M1_CDNS_69033583165443  M2_M1_CDNS_69033583165443_6
timestamp 1713338890
transform 1 0 -25830 0 1 -26696
box -874 -38 874 38
use M2_M1_CDNS_69033583165443  M2_M1_CDNS_69033583165443_7
timestamp 1713338890
transform 1 0 -25982 0 1 -26544
box -874 -38 874 38
use M2_M1_CDNS_69033583165443  M2_M1_CDNS_69033583165443_8
timestamp 1713338890
transform 1 0 -26134 0 1 -26392
box -874 -38 874 38
use M2_M1_CDNS_69033583165443  M2_M1_CDNS_69033583165443_9
timestamp 1713338890
transform 1 0 -26286 0 1 -26240
box -874 -38 874 38
use M2_M1_CDNS_69033583165443  M2_M1_CDNS_69033583165443_10
timestamp 1713338890
transform 1 0 -26438 0 1 -26088
box -874 -38 874 38
use M2_M1_CDNS_69033583165443  M2_M1_CDNS_69033583165443_11
timestamp 1713338890
transform 1 0 -26590 0 1 -25936
box -874 -38 874 38
use M2_M1_CDNS_69033583165443  M2_M1_CDNS_69033583165443_12
timestamp 1713338890
transform 1 0 -26742 0 1 -25784
box -874 -38 874 38
use M2_M1_CDNS_69033583165443  M2_M1_CDNS_69033583165443_13
timestamp 1713338890
transform 1 0 -26894 0 1 -25632
box -874 -38 874 38
use M2_M1_CDNS_69033583165445  M2_M1_CDNS_69033583165445_0
timestamp 1713338890
transform 1 0 -27366 0 1 -21818
box -494 -1482 494 1482
use M2_M1_CDNS_69033583165445  M2_M1_CDNS_69033583165445_1
timestamp 1713338890
transform 1 0 -22483 0 1 -22111
box -494 -1482 494 1482
use M2_M1_CDNS_69033583165445  M2_M1_CDNS_69033583165445_2
timestamp 1713338890
transform 1 0 -27354 0 1 -17335
box -494 -1482 494 1482
use M2_M1_CDNS_69033583165445  M2_M1_CDNS_69033583165445_3
timestamp 1713338890
transform 1 0 -22483 0 1 -17565
box -494 -1482 494 1482
use M2_M1_CDNS_69033583165449  M2_M1_CDNS_69033583165449_0
timestamp 1713338890
transform 1 0 -20046 0 1 -15668
box -494 -1330 494 1330
use M2_M1_CDNS_69033583165450  M2_M1_CDNS_69033583165450_0
timestamp 1713338890
transform 1 0 -24927 0 1 -15475
box -494 -1178 494 1178
use M2_M1_CDNS_69033583165454  M2_M1_CDNS_69033583165454_0
timestamp 1713338890
transform 1 0 -6846 0 1 -50175
box -170 -1292 170 1292
use M2_M1_CDNS_69033583165454  M2_M1_CDNS_69033583165454_1
timestamp 1713338890
transform 1 0 -9282 0 1 -50175
box -170 -1292 170 1292
use M2_M1_CDNS_69033583165454  M2_M1_CDNS_69033583165454_2
timestamp 1713338890
transform 1 0 -11708 0 1 -50175
box -170 -1292 170 1292
use M2_M1_CDNS_69033583165454  M2_M1_CDNS_69033583165454_3
timestamp 1713338890
transform 1 0 -14674 0 1 -48201
box -170 -1292 170 1292
use M2_M1_CDNS_69033583165454  M2_M1_CDNS_69033583165454_4
timestamp 1713338890
transform 1 0 -11708 0 1 -46375
box -170 -1292 170 1292
use M2_M1_CDNS_69033583165454  M2_M1_CDNS_69033583165454_5
timestamp 1713338890
transform 1 0 -17450 0 1 -44680
box -170 -1292 170 1292
use M2_M1_CDNS_69033583165454  M2_M1_CDNS_69033583165454_6
timestamp 1713338890
transform 1 0 -19888 0 1 -43196
box -170 -1292 170 1292
use M2_M1_CDNS_69033583165454  M2_M1_CDNS_69033583165454_7
timestamp 1713338890
transform 1 0 -14529 0 1 -43196
box -170 -1292 170 1292
use M2_M1_CDNS_69033583165454  M2_M1_CDNS_69033583165454_8
timestamp 1713338890
transform 1 0 -24750 0 1 -37781
box -170 -1292 170 1292
use M2_M1_CDNS_69033583165454  M2_M1_CDNS_69033583165454_9
timestamp 1713338890
transform 1 0 -22049 0 1 -35676
box -170 -1292 170 1292
use M2_M1_CDNS_69033583165454  M2_M1_CDNS_69033583165454_10
timestamp 1713338890
transform 1 0 -27517 0 1 -35676
box -170 -1292 170 1292
use M2_M1_CDNS_69033583165454  M2_M1_CDNS_69033583165454_11
timestamp 1713338890
transform 1 0 -29962 0 1 -32230
box -170 -1292 170 1292
use M2_M1_CDNS_69033583165454  M2_M1_CDNS_69033583165454_12
timestamp 1713338890
transform 1 0 -32401 0 1 -30500
box -170 -1292 170 1292
use M2_M1_CDNS_69033583165454  M2_M1_CDNS_69033583165454_13
timestamp 1713338890
transform 1 0 -27517 0 1 -30500
box -170 -1292 170 1292
use M2_M1_CDNS_69033583165455  M2_M1_CDNS_69033583165455_0
timestamp 1713338890
transform 1 0 -20832 0 1 -29202
box -434 -632 434 632
use M2_M1_CDNS_69033583165455  M2_M1_CDNS_69033583165455_1
timestamp 1713338890
transform 1 0 -15959 0 1 -29202
box -434 -632 434 632
use M2_M1_CDNS_69033583165456  M2_M1_CDNS_69033583165456_0
timestamp 1713338890
transform 1 0 -31074 0 1 -36991
box -570 -570 570 570
use M2_M1_CDNS_69033583165464  M2_M1_CDNS_69033583165464_0
timestamp 1713338890
transform 1 0 -34922 0 1 -32114
box -266 -1482 266 1482
use M2_M1_CDNS_69033583165466  M2_M1_CDNS_69033583165466_0
timestamp 1713338890
transform 1 0 -16281 0 1 -52063
box -722 -38 722 38
use M2_M1_CDNS_69033583165469  M2_M1_CDNS_69033583165469_0
timestamp 1713338890
transform 1 0 -5590 0 1 -37452
box -368 -1160 368 1160
use M2_M1_CDNS_69033583165469  M2_M1_CDNS_69033583165469_1
timestamp 1713338890
transform 1 0 -10498 0 1 -29849
box -368 -1160 368 1160
use M2_M1_CDNS_69033583165469  M2_M1_CDNS_69033583165469_2
timestamp 1713338890
transform 1 0 -5590 0 1 -29849
box -368 -1160 368 1160
use M2_M1_CDNS_69033583165470  M2_M1_CDNS_69033583165470_0
timestamp 1713338890
transform 1 0 -10498 0 1 -33018
box -368 -566 368 566
use M2_M1_CDNS_69033583165473  M2_M1_CDNS_69033583165473_0
timestamp 1713338890
transform 1 0 -9174 0 1 -53792
box -5252 -764 5252 764
use M2_M1_CDNS_69033583165474  M2_M1_CDNS_69033583165474_0
timestamp 1713338890
transform 1 0 -10487 0 1 -38325
box -434 -1292 434 1292
use M2_M1_CDNS_69033583165475  M2_M1_CDNS_69033583165475_0
timestamp 1713338890
transform 1 0 -16423 0 1 -46423
box -1292 -302 1292 302
use M2_M1_CDNS_69033583165476  M2_M1_CDNS_69033583165476_0
timestamp 1713338890
transform 1 0 -8110 0 1 -46423
box -3272 -302 3272 302
use M3_M2_CDNS_6903358316542  M3_M2_CDNS_6903358316542_0
timestamp 1713338890
transform 1 0 9643 0 1 -10945
box -162 -596 162 596
use M3_M2_CDNS_6903358316542  M3_M2_CDNS_6903358316542_1
timestamp 1713338890
transform 1 0 9635 0 1 -7796
box -162 -596 162 596
use M3_M2_CDNS_6903358316542  M3_M2_CDNS_6903358316542_2
timestamp 1713338890
transform 1 0 9655 0 1 -2992
box -162 -596 162 596
use M3_M2_CDNS_69033583165407  M3_M2_CDNS_69033583165407_0
timestamp 1713338890
transform 1 0 -19727 0 1 -47419
box -1178 -570 1178 570
use M3_M2_CDNS_69033583165407  M3_M2_CDNS_69033583165407_1
timestamp 1713338890
transform 1 0 -23781 0 1 -43365
box -1178 -570 1178 570
use M3_M2_CDNS_69033583165407  M3_M2_CDNS_69033583165407_2
timestamp 1713338890
transform 1 0 -25879 0 1 -41267
box -1178 -570 1178 570
use M3_M2_CDNS_69033583165408  M3_M2_CDNS_69033583165408_0
timestamp 1713338890
transform 1 0 -12921 0 1 -36139
box -434 -1622 434 1622
use M3_M2_CDNS_69033583165408  M3_M2_CDNS_69033583165408_1
timestamp 1713338890
transform 1 0 -8078 0 1 -36503
box -434 -1622 434 1622
use M3_M2_CDNS_69033583165408  M3_M2_CDNS_69033583165408_2
timestamp 1713338890
transform 1 0 -18419 0 1 -30678
box -434 -1622 434 1622
use M3_M2_CDNS_69033583165408  M3_M2_CDNS_69033583165408_3
timestamp 1713338890
transform 1 0 -12921 0 1 -31665
box -434 -1622 434 1622
use M3_M2_CDNS_69033583165408  M3_M2_CDNS_69033583165408_4
timestamp 1713338890
transform 1 0 -8041 0 1 -31997
box -434 -1622 434 1622
use M3_M2_CDNS_69033583165413  M3_M2_CDNS_69033583165413_0
timestamp 1713338890
transform 1 0 8277 0 1 -1404
box -368 -632 368 632
use M3_M2_CDNS_69033583165414  M3_M2_CDNS_69033583165414_0
timestamp 1713338890
transform 1 0 8869 0 1 38
box -968 -38 968 38
use M3_M2_CDNS_69033583165415  M3_M2_CDNS_69033583165415_0
timestamp 1713338890
transform 1 0 5824 0 1 -9409
box -410 -658 410 658
use M3_M2_CDNS_69033583165416  M3_M2_CDNS_69033583165416_0
timestamp 1713338890
transform 1 0 542 0 1 38
box -596 -38 596 38
use M3_M2_CDNS_69033583165416  M3_M2_CDNS_69033583165416_1
timestamp 1713338890
transform 1 0 5317 0 1 38
box -596 -38 596 38
use M3_M2_CDNS_69033583165418  M3_M2_CDNS_69033583165418_0
timestamp 1713338890
transform 1 0 -17015 0 1 -18078
box -494 -1102 494 1102
use M3_M2_CDNS_69033583165420  M3_M2_CDNS_69033583165420_0
timestamp 1713338890
transform 1 0 6950 0 1 -377
box -658 -38 658 38
use M3_M2_CDNS_69033583165426  M3_M2_CDNS_69033583165426_0
timestamp 1713338890
transform 1 0 -45402 0 1 -17451
box -1026 -5282 1026 5282
use M3_M2_CDNS_69033583165427  M3_M2_CDNS_69033583165427_0
timestamp 1713338890
transform 1 0 -32827 0 1 -21936
box -494 -266 494 266
use M3_M2_CDNS_69033583165427  M3_M2_CDNS_69033583165427_1
timestamp 1713338890
transform 1 0 -32918 0 1 -19655
box -494 -266 494 266
use M3_M2_CDNS_69033583165428  M3_M2_CDNS_69033583165428_0
timestamp 1713338890
transform 1 0 -14299 0 1 -40790
box -566 -38 566 38
use M3_M2_CDNS_69033583165428  M3_M2_CDNS_69033583165428_1
timestamp 1713338890
transform 1 0 -15374 0 1 -39715
box -566 -38 566 38
use M3_M2_CDNS_69033583165428  M3_M2_CDNS_69033583165428_2
timestamp 1713338890
transform 1 0 -32941 0 1 -13985
box -566 -38 566 38
use M3_M2_CDNS_69033583165428  M3_M2_CDNS_69033583165428_3
timestamp 1713338890
transform 1 0 -36244 0 1 -13985
box -566 -38 566 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_0
timestamp 1713338890
transform 1 0 -32235 0 1 -35063
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_1
timestamp 1713338890
transform 1 0 -32387 0 1 -34911
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_2
timestamp 1713338890
transform 1 0 -32539 0 1 -34759
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_3
timestamp 1713338890
transform 1 0 -32691 0 1 -34607
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_4
timestamp 1713338890
transform 1 0 -32843 0 1 -34455
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_5
timestamp 1713338890
transform 1 0 -32995 0 1 -34303
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_6
timestamp 1713338890
transform 1 0 -33147 0 1 -34151
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_7
timestamp 1713338890
transform 1 0 -33299 0 1 -33999
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_8
timestamp 1713338890
transform 1 0 -32083 0 1 -35215
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_9
timestamp 1713338890
transform 1 0 -31931 0 1 -35367
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_10
timestamp 1713338890
transform 1 0 -31779 0 1 -35519
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_11
timestamp 1713338890
transform 1 0 -33451 0 1 -33847
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_12
timestamp 1713338890
transform 1 0 -40754 0 1 -26544
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_13
timestamp 1713338890
transform 1 0 -41058 0 1 -26240
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_14
timestamp 1713338890
transform 1 0 -40906 0 1 -26392
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_15
timestamp 1713338890
transform 1 0 -41210 0 1 -26088
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_16
timestamp 1713338890
transform 1 0 -41362 0 1 -25936
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_17
timestamp 1713338890
transform 1 0 -41514 0 1 -25784
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_18
timestamp 1713338890
transform 1 0 -41666 0 1 -25632
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_19
timestamp 1713338890
transform 1 0 -37602 0 1 -29696
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_20
timestamp 1713338890
transform 1 0 -37754 0 1 -29544
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_21
timestamp 1713338890
transform 1 0 -37906 0 1 -29392
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_22
timestamp 1713338890
transform 1 0 -38058 0 1 -29240
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_23
timestamp 1713338890
transform 1 0 -38210 0 1 -29088
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_24
timestamp 1713338890
transform 1 0 -38362 0 1 -28936
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_25
timestamp 1713338890
transform 1 0 -38514 0 1 -28784
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_26
timestamp 1713338890
transform 1 0 -38666 0 1 -28632
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_27
timestamp 1713338890
transform 1 0 -38818 0 1 -28480
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_28
timestamp 1713338890
transform 1 0 -38970 0 1 -28328
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_29
timestamp 1713338890
transform 1 0 -39122 0 1 -28176
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_30
timestamp 1713338890
transform 1 0 -39274 0 1 -28024
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_31
timestamp 1713338890
transform 1 0 -39690 0 1 -27608
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_32
timestamp 1713338890
transform 1 0 -39842 0 1 -27456
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_33
timestamp 1713338890
transform 1 0 -39994 0 1 -27304
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_34
timestamp 1713338890
transform 1 0 -40146 0 1 -27152
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_35
timestamp 1713338890
transform 1 0 -40298 0 1 -27000
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_36
timestamp 1713338890
transform 1 0 -40450 0 1 -26848
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_37
timestamp 1713338890
transform 1 0 -40602 0 1 -26696
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_38
timestamp 1713338890
transform 1 0 -36130 0 1 -26544
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_39
timestamp 1713338890
transform 1 0 -36282 0 1 -26392
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_40
timestamp 1713338890
transform 1 0 -36434 0 1 -26240
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_41
timestamp 1713338890
transform 1 0 -36586 0 1 -26088
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_42
timestamp 1713338890
transform 1 0 -36738 0 1 -25936
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_43
timestamp 1713338890
transform 1 0 -36890 0 1 -25784
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_44
timestamp 1713338890
transform 1 0 -37042 0 1 -25632
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_45
timestamp 1713338890
transform 1 0 -35066 0 1 -27608
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_46
timestamp 1713338890
transform 1 0 -30567 0 1 -27608
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_47
timestamp 1713338890
transform 1 0 -35218 0 1 -27456
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_48
timestamp 1713338890
transform 1 0 -30719 0 1 -27456
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_49
timestamp 1713338890
transform 1 0 -35370 0 1 -27304
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_50
timestamp 1713338890
transform 1 0 -30871 0 1 -27304
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_51
timestamp 1713338890
transform 1 0 -31023 0 1 -27152
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_52
timestamp 1713338890
transform 1 0 -35522 0 1 -27152
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_53
timestamp 1713338890
transform 1 0 -31175 0 1 -27000
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_54
timestamp 1713338890
transform 1 0 -35674 0 1 -27000
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_55
timestamp 1713338890
transform 1 0 -31327 0 1 -26848
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_56
timestamp 1713338890
transform 1 0 -35826 0 1 -26848
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_57
timestamp 1713338890
transform 1 0 -31479 0 1 -26696
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_58
timestamp 1713338890
transform 1 0 -35978 0 1 -26696
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_59
timestamp 1713338890
transform 1 0 -32087 0 1 -26088
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_60
timestamp 1713338890
transform 1 0 -31783 0 1 -26392
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_61
timestamp 1713338890
transform 1 0 -31631 0 1 -26544
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_62
timestamp 1713338890
transform 1 0 -31935 0 1 -26240
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_63
timestamp 1713338890
transform 1 0 -32391 0 1 -25784
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_64
timestamp 1713338890
transform 1 0 -32543 0 1 -25632
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165429  M3_M2_CDNS_69033583165429_65
timestamp 1713338890
transform 1 0 -32239 0 1 -25936
box -1862 -38 1862 38
use M3_M2_CDNS_69033583165430  M3_M2_CDNS_69033583165430_0
timestamp 1713338890
transform 1 0 -32824 0 1 -16019
box -434 -1820 434 1820
use M3_M2_CDNS_69033583165437  M3_M2_CDNS_69033583165437_0
timestamp 1713338890
transform 1 0 -38682 0 1 -12857
box -1358 -632 1358 632
use M3_M2_CDNS_69033583165437  M3_M2_CDNS_69033583165437_1
timestamp 1713338890
transform 1 0 -41853 0 1 -12857
box -1358 -632 1358 632
use M3_M2_CDNS_69033583165440  M3_M2_CDNS_69033583165440_0
timestamp 1713338890
transform 1 0 -41853 0 1 -19655
box -1406 -266 1406 266
use M3_M2_CDNS_69033583165440  M3_M2_CDNS_69033583165440_1
timestamp 1713338890
transform 1 0 -38433 0 1 -19655
box -1406 -266 1406 266
use M3_M2_CDNS_69033583165444  M3_M2_CDNS_69033583165444_0
timestamp 1713338890
transform 1 0 -24918 0 1 -27608
box -874 -38 874 38
use M3_M2_CDNS_69033583165444  M3_M2_CDNS_69033583165444_1
timestamp 1713338890
transform 1 0 -25070 0 1 -27456
box -874 -38 874 38
use M3_M2_CDNS_69033583165444  M3_M2_CDNS_69033583165444_2
timestamp 1713338890
transform 1 0 -25222 0 1 -27304
box -874 -38 874 38
use M3_M2_CDNS_69033583165444  M3_M2_CDNS_69033583165444_3
timestamp 1713338890
transform 1 0 -25374 0 1 -27152
box -874 -38 874 38
use M3_M2_CDNS_69033583165444  M3_M2_CDNS_69033583165444_4
timestamp 1713338890
transform 1 0 -25526 0 1 -27000
box -874 -38 874 38
use M3_M2_CDNS_69033583165444  M3_M2_CDNS_69033583165444_5
timestamp 1713338890
transform 1 0 -25678 0 1 -26848
box -874 -38 874 38
use M3_M2_CDNS_69033583165444  M3_M2_CDNS_69033583165444_6
timestamp 1713338890
transform 1 0 -25830 0 1 -26696
box -874 -38 874 38
use M3_M2_CDNS_69033583165444  M3_M2_CDNS_69033583165444_7
timestamp 1713338890
transform 1 0 -25982 0 1 -26544
box -874 -38 874 38
use M3_M2_CDNS_69033583165444  M3_M2_CDNS_69033583165444_8
timestamp 1713338890
transform 1 0 -26134 0 1 -26392
box -874 -38 874 38
use M3_M2_CDNS_69033583165444  M3_M2_CDNS_69033583165444_9
timestamp 1713338890
transform 1 0 -26286 0 1 -26240
box -874 -38 874 38
use M3_M2_CDNS_69033583165444  M3_M2_CDNS_69033583165444_10
timestamp 1713338890
transform 1 0 -26438 0 1 -26088
box -874 -38 874 38
use M3_M2_CDNS_69033583165444  M3_M2_CDNS_69033583165444_11
timestamp 1713338890
transform 1 0 -26590 0 1 -25936
box -874 -38 874 38
use M3_M2_CDNS_69033583165444  M3_M2_CDNS_69033583165444_12
timestamp 1713338890
transform 1 0 -26894 0 1 -25632
box -874 -38 874 38
use M3_M2_CDNS_69033583165444  M3_M2_CDNS_69033583165444_13
timestamp 1713338890
transform 1 0 -26742 0 1 -25784
box -874 -38 874 38
use M3_M2_CDNS_69033583165446  M3_M2_CDNS_69033583165446_0
timestamp 1713338890
transform 1 0 -27366 0 1 -21818
box -494 -1482 494 1482
use M3_M2_CDNS_69033583165446  M3_M2_CDNS_69033583165446_1
timestamp 1713338890
transform 1 0 -22483 0 1 -22111
box -494 -1482 494 1482
use M3_M2_CDNS_69033583165446  M3_M2_CDNS_69033583165446_2
timestamp 1713338890
transform 1 0 -27354 0 1 -17335
box -494 -1482 494 1482
use M3_M2_CDNS_69033583165446  M3_M2_CDNS_69033583165446_3
timestamp 1713338890
transform 1 0 -22483 0 1 -17565
box -494 -1482 494 1482
use M3_M2_CDNS_69033583165447  M3_M2_CDNS_69033583165447_0
timestamp 1713338890
transform 1 0 -24927 0 1 -15475
box -494 -1178 494 1178
use M3_M2_CDNS_69033583165448  M3_M2_CDNS_69033583165448_0
timestamp 1713338890
transform 1 0 -20046 0 1 -15668
box -494 -1330 494 1330
use M3_M2_CDNS_69033583165452  M3_M2_CDNS_69033583165452_0
timestamp 1713338890
transform 1 0 -6846 0 1 -50175
box -170 -1292 170 1292
use M3_M2_CDNS_69033583165452  M3_M2_CDNS_69033583165452_1
timestamp 1713338890
transform 1 0 -9282 0 1 -50175
box -170 -1292 170 1292
use M3_M2_CDNS_69033583165452  M3_M2_CDNS_69033583165452_2
timestamp 1713338890
transform 1 0 -11708 0 1 -50175
box -170 -1292 170 1292
use M3_M2_CDNS_69033583165452  M3_M2_CDNS_69033583165452_3
timestamp 1713338890
transform 1 0 -14674 0 1 -48201
box -170 -1292 170 1292
use M3_M2_CDNS_69033583165452  M3_M2_CDNS_69033583165452_4
timestamp 1713338890
transform 1 0 -11708 0 1 -46375
box -170 -1292 170 1292
use M3_M2_CDNS_69033583165452  M3_M2_CDNS_69033583165452_5
timestamp 1713338890
transform 1 0 -17450 0 1 -44680
box -170 -1292 170 1292
use M3_M2_CDNS_69033583165452  M3_M2_CDNS_69033583165452_6
timestamp 1713338890
transform 1 0 -19888 0 1 -43196
box -170 -1292 170 1292
use M3_M2_CDNS_69033583165452  M3_M2_CDNS_69033583165452_7
timestamp 1713338890
transform 1 0 -14529 0 1 -43196
box -170 -1292 170 1292
use M3_M2_CDNS_69033583165452  M3_M2_CDNS_69033583165452_8
timestamp 1713338890
transform 1 0 -24750 0 1 -37781
box -170 -1292 170 1292
use M3_M2_CDNS_69033583165452  M3_M2_CDNS_69033583165452_9
timestamp 1713338890
transform 1 0 -22049 0 1 -35676
box -170 -1292 170 1292
use M3_M2_CDNS_69033583165452  M3_M2_CDNS_69033583165452_10
timestamp 1713338890
transform 1 0 -27517 0 1 -35676
box -170 -1292 170 1292
use M3_M2_CDNS_69033583165452  M3_M2_CDNS_69033583165452_11
timestamp 1713338890
transform 1 0 -29962 0 1 -32230
box -170 -1292 170 1292
use M3_M2_CDNS_69033583165452  M3_M2_CDNS_69033583165452_12
timestamp 1713338890
transform 1 0 -32401 0 1 -30500
box -170 -1292 170 1292
use M3_M2_CDNS_69033583165452  M3_M2_CDNS_69033583165452_13
timestamp 1713338890
transform 1 0 -27517 0 1 -30500
box -170 -1292 170 1292
use M3_M2_CDNS_69033583165453  M3_M2_CDNS_69033583165453_0
timestamp 1713338890
transform 1 0 -26321 0 1 -28433
box -830 -38 830 38
use M3_M2_CDNS_69033583165457  M3_M2_CDNS_69033583165457_0
timestamp 1713338890
transform 1 0 -31074 0 1 -36991
box -570 -570 570 570
use M3_M2_CDNS_69033583165458  M3_M2_CDNS_69033583165458_0
timestamp 1713338890
transform 1 0 -20832 0 1 -29202
box -434 -632 434 632
use M3_M2_CDNS_69033583165458  M3_M2_CDNS_69033583165458_1
timestamp 1713338890
transform 1 0 -15959 0 1 -29202
box -434 -632 434 632
use M3_M2_CDNS_69033583165461  M3_M2_CDNS_69033583165461_0
timestamp 1713338890
transform 1 0 -34922 0 1 -32114
box -266 -1482 266 1482
use M3_M2_CDNS_69033583165467  M3_M2_CDNS_69033583165467_0
timestamp 1713338890
transform 1 0 -8110 0 1 -46423
box -3272 -302 3272 302
use M3_M2_CDNS_69033583165468  M3_M2_CDNS_69033583165468_0
timestamp 1713338890
transform 1 0 -16423 0 1 -46423
box -1292 -302 1292 302
use M3_M2_CDNS_69033583165471  M3_M2_CDNS_69033583165471_0
timestamp 1713338890
transform 1 0 -10487 0 1 -38325
box -434 -1292 434 1292
use M3_M2_CDNS_69033583165472  M3_M2_CDNS_69033583165472_0
timestamp 1713338890
transform 1 0 -9174 0 1 -53792
box -5252 -764 5252 764
use M3_M2_CDNS_69033583165477  M3_M2_CDNS_69033583165477_0
timestamp 1713338890
transform 1 0 -10498 0 1 -33018
box -368 -566 368 566
use M3_M2_CDNS_69033583165478  M3_M2_CDNS_69033583165478_0
timestamp 1713338890
transform 1 0 -5590 0 1 -37452
box -368 -1160 368 1160
use M3_M2_CDNS_69033583165478  M3_M2_CDNS_69033583165478_1
timestamp 1713338890
transform 1 0 -10498 0 1 -29849
box -368 -1160 368 1160
use M3_M2_CDNS_69033583165478  M3_M2_CDNS_69033583165478_2
timestamp 1713338890
transform 1 0 -5590 0 1 -29849
box -368 -1160 368 1160
<< end >>
