* NGSPICE file created from TG_flat_flat.ext - technology: gf180mcuC

.subckt pex_TG VDD SEL VSS OUT IN 
X0 IN a_n2409_n525.t12 OUT.t21 VDD.t44 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 IN SEL.t0 OUT.t73 VSS.t49 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X2 IN a_n2409_n525.t13 OUT.t20 VDD.t43 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X3 OUT a_n2409_n525.t14 IN.t39 VDD.t42 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X4 OUT SEL.t1 IN.t62 VSS.t48 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X5 OUT a_n2409_n525.t15 IN.t38 VDD.t41 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X6 OUT a_n2409_n525.t16 IN.t37 VDD.t40 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X7 VSS SEL.t2 a_n2409_n525.t7 VSS.t45 nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.28u
X8 IN SEL.t3 OUT.t53 VSS.t44 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X9 IN SEL.t4 OUT.t67 VSS.t43 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X10 IN a_n2409_n525.t17 OUT.t19 VDD.t39 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X11 IN SEL.t5 OUT.t68 VSS.t42 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X12 IN SEL.t6 OUT.t54 VSS.t41 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X13 VDD SEL.t7 a_n2409_n525.t3 VDD.t45 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X14 OUT a_n2409_n525.t18 IN.t35 VDD.t38 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X15 OUT SEL.t8 IN.t74 VSS.t40 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X16 OUT SEL.t9 IN.t75 VSS.t39 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X17 OUT a_n2409_n525.t19 IN.t34 VDD.t37 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X18 IN SEL.t11 OUT.t57 VSS.t38 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X19 IN a_n2409_n525.t20 OUT.t18 VDD.t36 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X20 OUT SEL.t12 IN.t64 VSS.t37 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X21 IN a_n2409_n525.t21 OUT.t17 VDD.t35 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X22 VSS SEL.t13 a_n2409_n525.t9 VSS.t34 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X23 OUT a_n2409_n525.t22 IN.t31 VDD.t34 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X24 IN a_n2409_n525.t23 OUT.t16 VDD.t33 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X25 IN a_n2409_n525.t24 OUT.t15 VDD.t32 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X26 IN a_n2409_n525.t25 OUT.t14 VDD.t31 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X27 IN a_n2409_n525.t26 OUT.t13 VDD.t30 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X28 IN SEL.t14 OUT.t44 VSS.t33 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X29 IN SEL.t15 OUT.t45 VSS.t32 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X30 OUT a_n2409_n525.t27 IN.t26 VDD.t29 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X31 OUT SEL.t16 IN.t60 VSS.t31 nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.28u
X32 IN SEL.t17 OUT.t61 VSS.t30 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X33 OUT SEL.t18 IN.t46 VSS.t29 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X34 OUT a_n2409_n525.t28 IN.t25 VDD.t28 pfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.28u
X35 OUT a_n2409_n525.t29 IN.t24 VDD.t27 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X36 OUT SEL.t19 IN.t47 VSS.t28 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X37 IN a_n2409_n525.t30 OUT.t12 VDD.t26 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X38 IN a_n2409_n525.t31 OUT.t11 VDD.t25 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X39 VDD SEL.t20 a_n2409_n525.t1 VDD.t2 pfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.28u
X40 OUT SEL.t21 IN.t1 VSS.t27 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X41 OUT a_n2409_n525.t32 IN.t21 VDD.t24 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X42 OUT SEL.t22 IN.t69 VSS.t26 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X43 OUT SEL.t23 IN.t70 VSS.t25 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X44 OUT a_n2409_n525.t33 IN.t20 VDD.t23 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X45 IN SEL.t25 OUT.t59 VSS.t24 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X46 OUT SEL.t26 IN.t63 VSS.t23 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X47 VDD SEL.t27 a_n2409_n525.t8 VDD.t52 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X48 IN a_n2409_n525.t34 OUT.t10 VDD.t22 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X49 IN a_n2409_n525.t35 OUT.t9 VDD.t21 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X50 IN SEL.t28 OUT.t65 VSS.t22 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X51 IN SEL.t29 OUT.t66 VSS.t21 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X52 IN a_n2409_n525.t36 OUT.t8 VDD.t20 pfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.28u
X53 IN SEL.t30 OUT.t51 VSS.t20 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X54 OUT SEL.t31 IN.t52 VSS.t19 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X55 OUT a_n2409_n525.t37 IN.t16 VDD.t19 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X56 OUT a_n2409_n525.t38 IN.t15 VDD.t18 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X57 OUT a_n2409_n525.t39 IN.t14 VDD.t17 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X58 OUT SEL.t32 IN.t71 VSS.t18 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X59 IN SEL.t33 OUT.t72 VSS.t17 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X60 IN a_n2409_n525.t40 OUT.t7 VDD.t16 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X61 IN a_n2409_n525.t41 OUT.t6 VDD.t15 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X62 OUT a_n2409_n525.t42 IN.t11 VDD.t14 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X63 IN SEL.t34 OUT.t77 VSS.t16 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X64 OUT a_n2409_n525.t43 IN.t10 VDD.t13 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X65 IN a_n2409_n525.t44 OUT.t5 VDD.t12 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X66 OUT SEL.t35 IN.t78 VSS.t15 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X67 IN a_n2409_n525.t45 OUT.t4 VDD.t11 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X68 IN SEL.t36 OUT.t55 VSS.t14 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X69 OUT SEL.t37 IN.t56 VSS.t13 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X70 VDD SEL.t38 a_n2409_n525.t10 VDD.t55 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X71 IN SEL.t39 OUT.t76 VSS.t12 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X72 IN SEL.t40 OUT.t0 VSS.t11 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X73 OUT a_n2409_n525.t46 IN.t7 VDD.t10 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X74 OUT SEL.t43 IN.t58 VSS.t8 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X75 IN a_n2409_n525.t47 OUT.t3 VDD.t9 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X76 IN a_n2409_n525.t48 OUT.t2 VDD.t8 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X77 OUT SEL.t45 IN.t79 VSS.t7 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X78 OUT a_n2409_n525.t49 IN.t4 VDD.t7 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X79 OUT a_n2409_n525.t50 IN.t3 VDD.t6 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X80 IN SEL.t46 OUT.t42 VSS.t6 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X81 OUT SEL.t47 IN.t43 VSS.t5 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X82 IN SEL.t48 OUT.t48 VSS.t4 nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.28u
X83 OUT a_n2409_n525.t51 IN.t2 VDD.t5 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X84 OUT SEL.t50 IN.t49 VSS.t1 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X85 OUT SEL.t51 IN.t50 VSS.t0 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
R0 a_n2409_n525.n42 a_n2409_n525.t28 103.075
R1 a_n2409_n525.n4 a_n2409_n525.t36 49.5689
R2 a_n2409_n525.t28 a_n2409_n525.n41 49.5689
R3 a_n2409_n525.n4 a_n2409_n525.t39 26.0719
R4 a_n2409_n525.n5 a_n2409_n525.t35 26.0719
R5 a_n2409_n525.n6 a_n2409_n525.t38 26.0719
R6 a_n2409_n525.n7 a_n2409_n525.t48 26.0719
R7 a_n2409_n525.n8 a_n2409_n525.t19 26.0719
R8 a_n2409_n525.n9 a_n2409_n525.t20 26.0719
R9 a_n2409_n525.n10 a_n2409_n525.t33 26.0719
R10 a_n2409_n525.n11 a_n2409_n525.t34 26.0719
R11 a_n2409_n525.n12 a_n2409_n525.t32 26.0719
R12 a_n2409_n525.n13 a_n2409_n525.t45 26.0719
R13 a_n2409_n525.n14 a_n2409_n525.t46 26.0719
R14 a_n2409_n525.n15 a_n2409_n525.t17 26.0719
R15 a_n2409_n525.n16 a_n2409_n525.t18 26.0719
R16 a_n2409_n525.n17 a_n2409_n525.t31 26.0719
R17 a_n2409_n525.n18 a_n2409_n525.t29 26.0719
R18 a_n2409_n525.n19 a_n2409_n525.t30 26.0719
R19 a_n2409_n525.n20 a_n2409_n525.t42 26.0719
R20 a_n2409_n525.n21 a_n2409_n525.t44 26.0719
R21 a_n2409_n525.n22 a_n2409_n525.t16 26.0719
R22 a_n2409_n525.n23 a_n2409_n525.t26 26.0719
R23 a_n2409_n525.n24 a_n2409_n525.t14 26.0719
R24 a_n2409_n525.n25 a_n2409_n525.t25 26.0719
R25 a_n2409_n525.n26 a_n2409_n525.t27 26.0719
R26 a_n2409_n525.n27 a_n2409_n525.t40 26.0719
R27 a_n2409_n525.n28 a_n2409_n525.t50 26.0719
R28 a_n2409_n525.n29 a_n2409_n525.t12 26.0719
R29 a_n2409_n525.n30 a_n2409_n525.t22 26.0719
R30 a_n2409_n525.n31 a_n2409_n525.t24 26.0719
R31 a_n2409_n525.n32 a_n2409_n525.t37 26.0719
R32 a_n2409_n525.n33 a_n2409_n525.t47 26.0719
R33 a_n2409_n525.n34 a_n2409_n525.t51 26.0719
R34 a_n2409_n525.n35 a_n2409_n525.t21 26.0719
R35 a_n2409_n525.n36 a_n2409_n525.t49 26.0719
R36 a_n2409_n525.n37 a_n2409_n525.t23 26.0719
R37 a_n2409_n525.n38 a_n2409_n525.t15 26.0719
R38 a_n2409_n525.n39 a_n2409_n525.t13 26.0719
R39 a_n2409_n525.n40 a_n2409_n525.t43 26.0719
R40 a_n2409_n525.n41 a_n2409_n525.t41 26.0719
R41 a_n2409_n525.n5 a_n2409_n525.n4 19.6341
R42 a_n2409_n525.n6 a_n2409_n525.n5 19.6341
R43 a_n2409_n525.n7 a_n2409_n525.n6 19.6341
R44 a_n2409_n525.n8 a_n2409_n525.n7 19.6341
R45 a_n2409_n525.n9 a_n2409_n525.n8 19.6341
R46 a_n2409_n525.n10 a_n2409_n525.n9 19.6341
R47 a_n2409_n525.n11 a_n2409_n525.n10 19.6341
R48 a_n2409_n525.n12 a_n2409_n525.n11 19.6341
R49 a_n2409_n525.n13 a_n2409_n525.n12 19.6341
R50 a_n2409_n525.n14 a_n2409_n525.n13 19.6341
R51 a_n2409_n525.n15 a_n2409_n525.n14 19.6341
R52 a_n2409_n525.n16 a_n2409_n525.n15 19.6341
R53 a_n2409_n525.n17 a_n2409_n525.n16 19.6341
R54 a_n2409_n525.n18 a_n2409_n525.n17 19.6341
R55 a_n2409_n525.n19 a_n2409_n525.n18 19.6341
R56 a_n2409_n525.n20 a_n2409_n525.n19 19.6341
R57 a_n2409_n525.n21 a_n2409_n525.n20 19.6341
R58 a_n2409_n525.n22 a_n2409_n525.n21 19.6341
R59 a_n2409_n525.n23 a_n2409_n525.n22 19.6341
R60 a_n2409_n525.n24 a_n2409_n525.n23 19.6341
R61 a_n2409_n525.n25 a_n2409_n525.n24 19.6341
R62 a_n2409_n525.n26 a_n2409_n525.n25 19.6341
R63 a_n2409_n525.n27 a_n2409_n525.n26 19.6341
R64 a_n2409_n525.n28 a_n2409_n525.n27 19.6341
R65 a_n2409_n525.n29 a_n2409_n525.n28 19.6341
R66 a_n2409_n525.n30 a_n2409_n525.n29 19.6341
R67 a_n2409_n525.n31 a_n2409_n525.n30 19.6341
R68 a_n2409_n525.n32 a_n2409_n525.n31 19.6341
R69 a_n2409_n525.n33 a_n2409_n525.n32 19.6341
R70 a_n2409_n525.n34 a_n2409_n525.n33 19.6341
R71 a_n2409_n525.n35 a_n2409_n525.n34 19.6341
R72 a_n2409_n525.n36 a_n2409_n525.n35 19.6341
R73 a_n2409_n525.n37 a_n2409_n525.n36 19.6341
R74 a_n2409_n525.n38 a_n2409_n525.n37 19.6341
R75 a_n2409_n525.n39 a_n2409_n525.n38 19.6341
R76 a_n2409_n525.n40 a_n2409_n525.n39 19.6341
R77 a_n2409_n525.n41 a_n2409_n525.n40 19.6341
R78 a_n2409_n525.n50 a_n2409_n525.n1 3.7805
R79 a_n2409_n525.n49 a_n2409_n525.n46 3.7805
R80 a_n2409_n525.n49 a_n2409_n525.n48 3.7255
R81 a_n2409_n525.n42 a_n2409_n525.n3 3.13775
R82 a_n2409_n525.n49 a_n2409_n525.n44 3.09941
R83 a_n2409_n525.n51 a_n2409_n525.n50 3.09941
R84 a_n2409_n525.n3 a_n2409_n525.t1 0.9105
R85 a_n2409_n525.n3 a_n2409_n525.n2 0.9105
R86 a_n2409_n525.n44 a_n2409_n525.t10 0.9105
R87 a_n2409_n525.n44 a_n2409_n525.n43 0.9105
R88 a_n2409_n525.n48 a_n2409_n525.t8 0.9105
R89 a_n2409_n525.n48 a_n2409_n525.n47 0.9105
R90 a_n2409_n525.n51 a_n2409_n525.t3 0.9105
R91 a_n2409_n525.n52 a_n2409_n525.n51 0.9105
R92 a_n2409_n525.n1 a_n2409_n525.t7 0.8195
R93 a_n2409_n525.n1 a_n2409_n525.n0 0.8195
R94 a_n2409_n525.n46 a_n2409_n525.t9 0.8195
R95 a_n2409_n525.n46 a_n2409_n525.n45 0.8195
R96 a_n2409_n525.n50 a_n2409_n525.n49 0.626587
R97 a_n2409_n525.n50 a_n2409_n525.n42 0.565935
R98 OUT.n4 OUT.n1 3.81941
R99 OUT.n9 OUT.n6 3.81941
R100 OUT.n14 OUT.n11 3.81941
R101 OUT.n19 OUT.n16 3.81941
R102 OUT.n24 OUT.n21 3.81941
R103 OUT.n29 OUT.n26 3.81941
R104 OUT.n34 OUT.n31 3.81941
R105 OUT.n39 OUT.n36 3.81941
R106 OUT.n44 OUT.n41 3.81941
R107 OUT.n49 OUT.n46 3.81941
R108 OUT.n54 OUT.n51 3.81941
R109 OUT.n59 OUT.n56 3.81941
R110 OUT.n64 OUT.n61 3.81941
R111 OUT.n69 OUT.n66 3.81941
R112 OUT.n74 OUT.n71 3.81941
R113 OUT.n79 OUT.n76 3.81941
R114 OUT.n84 OUT.n81 3.81941
R115 OUT.n89 OUT.n86 3.81941
R116 OUT.n94 OUT.n91 3.81941
R117 OUT.n99 OUT.n96 3.81941
R118 OUT.n4 OUT.n3 3.1505
R119 OUT.n9 OUT.n8 3.1505
R120 OUT.n14 OUT.n13 3.1505
R121 OUT.n19 OUT.n18 3.1505
R122 OUT.n24 OUT.n23 3.1505
R123 OUT.n29 OUT.n28 3.1505
R124 OUT.n34 OUT.n33 3.1505
R125 OUT.n39 OUT.n38 3.1505
R126 OUT.n44 OUT.n43 3.1505
R127 OUT.n49 OUT.n48 3.1505
R128 OUT.n54 OUT.n53 3.1505
R129 OUT.n59 OUT.n58 3.1505
R130 OUT.n64 OUT.n63 3.1505
R131 OUT.n69 OUT.n68 3.1505
R132 OUT.n74 OUT.n73 3.1505
R133 OUT.n79 OUT.n78 3.1505
R134 OUT.n84 OUT.n83 3.1505
R135 OUT.n89 OUT.n88 3.1505
R136 OUT.n94 OUT.n93 3.1505
R137 OUT.n99 OUT.n98 3.1505
R138 OUT.n1 OUT.t8 0.9105
R139 OUT.n1 OUT.n0 0.9105
R140 OUT.n6 OUT.t9 0.9105
R141 OUT.n6 OUT.n5 0.9105
R142 OUT.n11 OUT.t2 0.9105
R143 OUT.n11 OUT.n10 0.9105
R144 OUT.n16 OUT.t18 0.9105
R145 OUT.n16 OUT.n15 0.9105
R146 OUT.n21 OUT.t10 0.9105
R147 OUT.n21 OUT.n20 0.9105
R148 OUT.n26 OUT.t4 0.9105
R149 OUT.n26 OUT.n25 0.9105
R150 OUT.n31 OUT.t19 0.9105
R151 OUT.n31 OUT.n30 0.9105
R152 OUT.n36 OUT.t11 0.9105
R153 OUT.n36 OUT.n35 0.9105
R154 OUT.n41 OUT.t12 0.9105
R155 OUT.n41 OUT.n40 0.9105
R156 OUT.n46 OUT.t5 0.9105
R157 OUT.n46 OUT.n45 0.9105
R158 OUT.n51 OUT.t13 0.9105
R159 OUT.n51 OUT.n50 0.9105
R160 OUT.n56 OUT.t14 0.9105
R161 OUT.n56 OUT.n55 0.9105
R162 OUT.n61 OUT.t7 0.9105
R163 OUT.n61 OUT.n60 0.9105
R164 OUT.n66 OUT.t21 0.9105
R165 OUT.n66 OUT.n65 0.9105
R166 OUT.n71 OUT.t15 0.9105
R167 OUT.n71 OUT.n70 0.9105
R168 OUT.n76 OUT.t3 0.9105
R169 OUT.n76 OUT.n75 0.9105
R170 OUT.n81 OUT.t17 0.9105
R171 OUT.n81 OUT.n80 0.9105
R172 OUT.n86 OUT.t16 0.9105
R173 OUT.n86 OUT.n85 0.9105
R174 OUT.n91 OUT.t20 0.9105
R175 OUT.n91 OUT.n90 0.9105
R176 OUT.n96 OUT.t6 0.9105
R177 OUT.n96 OUT.n95 0.9105
R178 OUT.n3 OUT.t48 0.8195
R179 OUT.n3 OUT.n2 0.8195
R180 OUT.n8 OUT.t0 0.8195
R181 OUT.n8 OUT.n7 0.8195
R182 OUT.n13 OUT.t66 0.8195
R183 OUT.n13 OUT.n12 0.8195
R184 OUT.n18 OUT.t45 0.8195
R185 OUT.n18 OUT.n17 0.8195
R186 OUT.n23 OUT.t67 0.8195
R187 OUT.n23 OUT.n22 0.8195
R188 OUT.n28 OUT.t72 0.8195
R189 OUT.n28 OUT.n27 0.8195
R190 OUT.n33 OUT.t61 0.8195
R191 OUT.n33 OUT.n32 0.8195
R192 OUT.n38 OUT.t54 0.8195
R193 OUT.n38 OUT.n37 0.8195
R194 OUT.n43 OUT.t73 0.8195
R195 OUT.n43 OUT.n42 0.8195
R196 OUT.n48 OUT.t55 0.8195
R197 OUT.n48 OUT.n47 0.8195
R198 OUT.n53 OUT.t57 0.8195
R199 OUT.n53 OUT.n52 0.8195
R200 OUT.n58 OUT.t53 0.8195
R201 OUT.n58 OUT.n57 0.8195
R202 OUT.n63 OUT.t76 0.8195
R203 OUT.n63 OUT.n62 0.8195
R204 OUT.n68 OUT.t65 0.8195
R205 OUT.n68 OUT.n67 0.8195
R206 OUT.n73 OUT.t59 0.8195
R207 OUT.n73 OUT.n72 0.8195
R208 OUT.n78 OUT.t42 0.8195
R209 OUT.n78 OUT.n77 0.8195
R210 OUT.n83 OUT.t77 0.8195
R211 OUT.n83 OUT.n82 0.8195
R212 OUT.n88 OUT.t68 0.8195
R213 OUT.n88 OUT.n87 0.8195
R214 OUT.n93 OUT.t44 0.8195
R215 OUT.n93 OUT.n92 0.8195
R216 OUT.n98 OUT.t51 0.8195
R217 OUT.n98 OUT.n97 0.8195
R218 OUT.n100 OUT.n99 0.730098
R219 OUT.n118 OUT.n4 0.503326
R220 OUT.n117 OUT.n9 0.503326
R221 OUT.n116 OUT.n14 0.503326
R222 OUT.n115 OUT.n19 0.503326
R223 OUT.n114 OUT.n24 0.503326
R224 OUT.n113 OUT.n29 0.503326
R225 OUT.n112 OUT.n34 0.503326
R226 OUT.n111 OUT.n39 0.503326
R227 OUT.n110 OUT.n44 0.503326
R228 OUT.n109 OUT.n49 0.503326
R229 OUT.n108 OUT.n54 0.503326
R230 OUT.n107 OUT.n59 0.503326
R231 OUT.n106 OUT.n64 0.503326
R232 OUT.n105 OUT.n69 0.503326
R233 OUT.n104 OUT.n74 0.503326
R234 OUT.n103 OUT.n79 0.503326
R235 OUT.n102 OUT.n84 0.503326
R236 OUT.n101 OUT.n89 0.503326
R237 OUT.n100 OUT.n94 0.503326
R238 OUT OUT.n118 0.267665
R239 OUT.n118 OUT.n117 0.227272
R240 OUT.n117 OUT.n116 0.227272
R241 OUT.n116 OUT.n115 0.227272
R242 OUT.n115 OUT.n114 0.227272
R243 OUT.n114 OUT.n113 0.227272
R244 OUT.n113 OUT.n112 0.227272
R245 OUT.n112 OUT.n111 0.227272
R246 OUT.n111 OUT.n110 0.227272
R247 OUT.n110 OUT.n109 0.227272
R248 OUT.n109 OUT.n108 0.227272
R249 OUT.n108 OUT.n107 0.227272
R250 OUT.n107 OUT.n106 0.227272
R251 OUT.n106 OUT.n105 0.227272
R252 OUT.n105 OUT.n104 0.227272
R253 OUT.n104 OUT.n103 0.227272
R254 OUT.n103 OUT.n102 0.227272
R255 OUT.n102 OUT.n101 0.227272
R256 OUT.n101 OUT.n100 0.227272
R257 IN.n97 IN.n96 5.18841
R258 IN.n4 IN.n3 4.36941
R259 IN.n9 IN.n8 4.36941
R260 IN.n14 IN.n13 4.36941
R261 IN.n19 IN.n18 4.36941
R262 IN.n24 IN.n23 4.36941
R263 IN.n29 IN.n28 4.36941
R264 IN.n34 IN.n33 4.36941
R265 IN.n39 IN.n38 4.36941
R266 IN.n44 IN.n43 4.36941
R267 IN.n49 IN.n48 4.36941
R268 IN.n54 IN.n53 4.36941
R269 IN.n59 IN.n58 4.36941
R270 IN.n64 IN.n63 4.36941
R271 IN.n69 IN.n68 4.36941
R272 IN.n74 IN.n73 4.36941
R273 IN.n79 IN.n78 4.36941
R274 IN.n84 IN.n83 4.36941
R275 IN.n89 IN.n88 4.36941
R276 IN.n94 IN.n93 4.36941
R277 IN.n118 IN.t60 4.08655
R278 IN.n117 IN.t25 3.5105
R279 IN.n97 IN.n95 3.5105
R280 IN.n120 IN.n118 3.22511
R281 IN.n4 IN.n1 2.6005
R282 IN.n9 IN.n6 2.6005
R283 IN.n14 IN.n11 2.6005
R284 IN.n19 IN.n16 2.6005
R285 IN.n24 IN.n21 2.6005
R286 IN.n29 IN.n26 2.6005
R287 IN.n34 IN.n31 2.6005
R288 IN.n39 IN.n36 2.6005
R289 IN.n44 IN.n41 2.6005
R290 IN.n49 IN.n46 2.6005
R291 IN.n54 IN.n51 2.6005
R292 IN.n59 IN.n56 2.6005
R293 IN.n64 IN.n61 2.6005
R294 IN.n69 IN.n66 2.6005
R295 IN.n74 IN.n71 2.6005
R296 IN.n79 IN.n76 2.6005
R297 IN.n84 IN.n81 2.6005
R298 IN.n89 IN.n86 2.6005
R299 IN.n94 IN.n91 2.6005
R300 IN.n120 IN.n119 2.25773
R301 IN.n1 IN.t10 0.9105
R302 IN.n1 IN.n0 0.9105
R303 IN.n6 IN.t38 0.9105
R304 IN.n6 IN.n5 0.9105
R305 IN.n11 IN.t4 0.9105
R306 IN.n11 IN.n10 0.9105
R307 IN.n16 IN.t2 0.9105
R308 IN.n16 IN.n15 0.9105
R309 IN.n21 IN.t16 0.9105
R310 IN.n21 IN.n20 0.9105
R311 IN.n26 IN.t31 0.9105
R312 IN.n26 IN.n25 0.9105
R313 IN.n31 IN.t3 0.9105
R314 IN.n31 IN.n30 0.9105
R315 IN.n36 IN.t26 0.9105
R316 IN.n36 IN.n35 0.9105
R317 IN.n41 IN.t39 0.9105
R318 IN.n41 IN.n40 0.9105
R319 IN.n46 IN.t37 0.9105
R320 IN.n46 IN.n45 0.9105
R321 IN.n51 IN.t11 0.9105
R322 IN.n51 IN.n50 0.9105
R323 IN.n56 IN.t24 0.9105
R324 IN.n56 IN.n55 0.9105
R325 IN.n61 IN.t35 0.9105
R326 IN.n61 IN.n60 0.9105
R327 IN.n66 IN.t7 0.9105
R328 IN.n66 IN.n65 0.9105
R329 IN.n71 IN.t21 0.9105
R330 IN.n71 IN.n70 0.9105
R331 IN.n76 IN.t20 0.9105
R332 IN.n76 IN.n75 0.9105
R333 IN.n81 IN.t34 0.9105
R334 IN.n81 IN.n80 0.9105
R335 IN.n86 IN.t15 0.9105
R336 IN.n86 IN.n85 0.9105
R337 IN.n91 IN.t14 0.9105
R338 IN.n91 IN.n90 0.9105
R339 IN.n3 IN.t74 0.8195
R340 IN.n3 IN.n2 0.8195
R341 IN.n8 IN.t79 0.8195
R342 IN.n8 IN.n7 0.8195
R343 IN.n13 IN.t71 0.8195
R344 IN.n13 IN.n12 0.8195
R345 IN.n18 IN.t69 0.8195
R346 IN.n18 IN.n17 0.8195
R347 IN.n23 IN.t78 0.8195
R348 IN.n23 IN.n22 0.8195
R349 IN.n28 IN.t49 0.8195
R350 IN.n28 IN.n27 0.8195
R351 IN.n33 IN.t62 0.8195
R352 IN.n33 IN.n32 0.8195
R353 IN.n38 IN.t52 0.8195
R354 IN.n38 IN.n37 0.8195
R355 IN.n43 IN.t58 0.8195
R356 IN.n43 IN.n42 0.8195
R357 IN.n48 IN.t50 0.8195
R358 IN.n48 IN.n47 0.8195
R359 IN.n53 IN.t64 0.8195
R360 IN.n53 IN.n52 0.8195
R361 IN.n58 IN.t1 0.8195
R362 IN.n58 IN.n57 0.8195
R363 IN.n63 IN.t43 0.8195
R364 IN.n63 IN.n62 0.8195
R365 IN.n68 IN.t75 0.8195
R366 IN.n68 IN.n67 0.8195
R367 IN.n73 IN.t47 0.8195
R368 IN.n73 IN.n72 0.8195
R369 IN.n78 IN.t63 0.8195
R370 IN.n78 IN.n77 0.8195
R371 IN.n83 IN.t56 0.8195
R372 IN.n83 IN.n82 0.8195
R373 IN.n88 IN.t46 0.8195
R374 IN.n88 IN.n87 0.8195
R375 IN.n93 IN.t70 0.8195
R376 IN.n93 IN.n92 0.8195
R377 IN.n98 IN.n97 0.688999
R378 IN.n116 IN.n4 0.481804
R379 IN.n115 IN.n9 0.481804
R380 IN.n114 IN.n14 0.481804
R381 IN.n113 IN.n19 0.481804
R382 IN.n112 IN.n24 0.481804
R383 IN.n111 IN.n29 0.481804
R384 IN.n110 IN.n34 0.481804
R385 IN.n109 IN.n39 0.481804
R386 IN.n108 IN.n44 0.481804
R387 IN.n107 IN.n49 0.481804
R388 IN.n106 IN.n54 0.481804
R389 IN.n105 IN.n59 0.481804
R390 IN.n104 IN.n64 0.481804
R391 IN.n103 IN.n69 0.481804
R392 IN.n102 IN.n74 0.481804
R393 IN.n101 IN.n79 0.481804
R394 IN.n100 IN.n84 0.481804
R395 IN.n99 IN.n89 0.481804
R396 IN.n98 IN.n94 0.481804
R397 IN.n117 IN.n116 0.437976
R398 IN.n118 IN.n117 0.434305
R399 IN.n99 IN.n98 0.207694
R400 IN.n100 IN.n99 0.207694
R401 IN.n101 IN.n100 0.207694
R402 IN.n102 IN.n101 0.207694
R403 IN.n103 IN.n102 0.207694
R404 IN.n104 IN.n103 0.207694
R405 IN.n105 IN.n104 0.207694
R406 IN.n106 IN.n105 0.207694
R407 IN.n107 IN.n106 0.207694
R408 IN.n108 IN.n107 0.207694
R409 IN.n109 IN.n108 0.207694
R410 IN.n110 IN.n109 0.207694
R411 IN.n111 IN.n110 0.207694
R412 IN.n112 IN.n111 0.207694
R413 IN.n113 IN.n112 0.207694
R414 IN.n114 IN.n113 0.207694
R415 IN.n115 IN.n114 0.207694
R416 IN.n116 IN.n115 0.207694
R417 IN IN.n120 0.00772628
R418 VDD.n106 VDD.t45 131.47
R419 VDD.n121 VDD.t50 131.47
R420 VDD.n83 VDD.t41 106.912
R421 VDD.n17 VDD.t23 101.513
R422 VDD.n29 VDD.t39 101.513
R423 VDD.n41 VDD.t26 98.2726
R424 VDD.n53 VDD.t42 98.2726
R425 VDD.n106 VDD.t48 92.3082
R426 VDD.n121 VDD.t52 92.3082
R427 VDD.n62 VDD.t44 90.7132
R428 VDD.n74 VDD.t5 90.7132
R429 VDD.n8 VDD.t21 87.4735
R430 VDD.n8 VDD.t18 85.3137
R431 VDD.n62 VDD.t6 82.0739
R432 VDD.n74 VDD.t9 82.0739
R433 VDD.n110 VDD.t0 75.525
R434 VDD.n41 VDD.t14 74.5145
R435 VDD.n53 VDD.t31 74.5145
R436 VDD.n17 VDD.t36 71.2748
R437 VDD.n29 VDD.t10 71.2748
R438 VDD.n83 VDD.t33 65.8752
R439 VDD.n95 VDD.t28 65.8752
R440 VDD.n86 VDD.t43 63.7154
R441 VDD.n20 VDD.t22 58.3158
R442 VDD.n32 VDD.t38 58.3158
R443 VDD.n38 VDD.t27 55.0761
R444 VDD.n50 VDD.t30 55.0761
R445 VDD.n65 VDD.t34 47.5167
R446 VDD.n77 VDD.t35 47.5167
R447 VDD.n4 VDD.t17 44.277
R448 VDD.n11 VDD.t8 42.1171
R449 VDD.n59 VDD.t16 38.8774
R450 VDD.n71 VDD.t19 38.8774
R451 VDD.n103 VDD.t2 36.3641
R452 VDD.n125 VDD.t58 36.3641
R453 VDD.n44 VDD.t12 31.318
R454 VDD.n56 VDD.t29 31.318
R455 VDD.n26 VDD.t11 28.0783
R456 VDD.n80 VDD.t7 22.6787
R457 VDD.n92 VDD.t15 22.6787
R458 VDD.n89 VDD.t13 20.5189
R459 VDD.n114 VDD.t55 19.5809
R460 VDD.n23 VDD.t24 15.1193
R461 VDD.n35 VDD.t25 15.1193
R462 VDD.n47 VDD.t40 11.8796
R463 VDD.n7 VDD.n6 5.41383
R464 VDD.n68 VDD.t32 4.32015
R465 VDD.n102 VDD.n101 4.00449
R466 VDD.n120 VDD.t51 3.98789
R467 VDD.n120 VDD.n119 3.1671
R468 VDD.n5 VDD.n4 3.1505
R469 VDD.n10 VDD.n9 3.1505
R470 VDD.n9 VDD.n8 3.1505
R471 VDD.n13 VDD.n12 3.1505
R472 VDD.n12 VDD.n11 3.1505
R473 VDD.n16 VDD.n15 3.1505
R474 VDD.n15 VDD.n14 3.1505
R475 VDD.n19 VDD.n18 3.1505
R476 VDD.n18 VDD.n17 3.1505
R477 VDD.n22 VDD.n21 3.1505
R478 VDD.n21 VDD.n20 3.1505
R479 VDD.n25 VDD.n24 3.1505
R480 VDD.n24 VDD.n23 3.1505
R481 VDD.n28 VDD.n27 3.1505
R482 VDD.n27 VDD.n26 3.1505
R483 VDD.n31 VDD.n30 3.1505
R484 VDD.n30 VDD.n29 3.1505
R485 VDD.n34 VDD.n33 3.1505
R486 VDD.n33 VDD.n32 3.1505
R487 VDD.n37 VDD.n36 3.1505
R488 VDD.n36 VDD.n35 3.1505
R489 VDD.n40 VDD.n39 3.1505
R490 VDD.n39 VDD.n38 3.1505
R491 VDD.n43 VDD.n42 3.1505
R492 VDD.n42 VDD.n41 3.1505
R493 VDD.n46 VDD.n45 3.1505
R494 VDD.n45 VDD.n44 3.1505
R495 VDD.n49 VDD.n48 3.1505
R496 VDD.n48 VDD.n47 3.1505
R497 VDD.n52 VDD.n51 3.1505
R498 VDD.n51 VDD.n50 3.1505
R499 VDD.n55 VDD.n54 3.1505
R500 VDD.n54 VDD.n53 3.1505
R501 VDD.n58 VDD.n57 3.1505
R502 VDD.n57 VDD.n56 3.1505
R503 VDD.n61 VDD.n60 3.1505
R504 VDD.n60 VDD.n59 3.1505
R505 VDD.n64 VDD.n63 3.1505
R506 VDD.n63 VDD.n62 3.1505
R507 VDD.n67 VDD.n66 3.1505
R508 VDD.n66 VDD.n65 3.1505
R509 VDD.n70 VDD.n69 3.1505
R510 VDD.n69 VDD.n68 3.1505
R511 VDD.n73 VDD.n72 3.1505
R512 VDD.n72 VDD.n71 3.1505
R513 VDD.n76 VDD.n75 3.1505
R514 VDD.n75 VDD.n74 3.1505
R515 VDD.n79 VDD.n78 3.1505
R516 VDD.n78 VDD.n77 3.1505
R517 VDD.n82 VDD.n81 3.1505
R518 VDD.n81 VDD.n80 3.1505
R519 VDD.n85 VDD.n84 3.1505
R520 VDD.n84 VDD.n83 3.1505
R521 VDD.n88 VDD.n87 3.1505
R522 VDD.n87 VDD.n86 3.1505
R523 VDD.n91 VDD.n90 3.1505
R524 VDD.n90 VDD.n89 3.1505
R525 VDD.n94 VDD.n93 3.1505
R526 VDD.n93 VDD.n92 3.1505
R527 VDD.n97 VDD.n96 3.1505
R528 VDD.n96 VDD.n95 3.1505
R529 VDD.n100 VDD.n99 3.1505
R530 VDD.n99 VDD.n98 3.1505
R531 VDD.n108 VDD.n107 3.1505
R532 VDD.n107 VDD.n106 3.1505
R533 VDD.n112 VDD.n111 3.1505
R534 VDD.n111 VDD.n110 3.1505
R535 VDD.n116 VDD.n115 3.1505
R536 VDD.n115 VDD.n114 3.1505
R537 VDD.n127 VDD.n126 3.1505
R538 VDD.n126 VDD.n125 3.1505
R539 VDD.n123 VDD.n122 3.1505
R540 VDD.n122 VDD.n121 3.1505
R541 VDD.n105 VDD.n104 3.1505
R542 VDD.n104 VDD.n103 3.1505
R543 VDD.n124 VDD.n118 3.07789
R544 VDD.n113 VDD.n1 3.07789
R545 VDD.n109 VDD.n3 3.07789
R546 VDD.n7 VDD.n5 2.17513
R547 VDD.n6 VDD.t20 1.08041
R548 VDD.n14 VDD.t37 1.08041
R549 VDD.n118 VDD.t59 0.9105
R550 VDD.n118 VDD.n117 0.9105
R551 VDD.n1 VDD.t1 0.9105
R552 VDD.n1 VDD.n0 0.9105
R553 VDD.n3 VDD.t49 0.9105
R554 VDD.n3 VDD.n2 0.9105
R555 VDD.n10 VDD.n7 0.626574
R556 VDD.n19 VDD.n16 0.144117
R557 VDD.n40 VDD.n37 0.144117
R558 VDD.n61 VDD.n58 0.144117
R559 VDD.n82 VDD.n79 0.144117
R560 VDD.n13 VDD.n10 0.12816
R561 VDD.n16 VDD.n13 0.12816
R562 VDD.n22 VDD.n19 0.12816
R563 VDD.n25 VDD.n22 0.12816
R564 VDD.n28 VDD.n25 0.12816
R565 VDD.n31 VDD.n28 0.12816
R566 VDD.n34 VDD.n31 0.12816
R567 VDD.n37 VDD.n34 0.12816
R568 VDD.n43 VDD.n40 0.12816
R569 VDD.n46 VDD.n43 0.12816
R570 VDD.n49 VDD.n46 0.12816
R571 VDD.n52 VDD.n49 0.12816
R572 VDD.n55 VDD.n52 0.12816
R573 VDD.n58 VDD.n55 0.12816
R574 VDD.n64 VDD.n61 0.12816
R575 VDD.n67 VDD.n64 0.12816
R576 VDD.n70 VDD.n67 0.12816
R577 VDD.n73 VDD.n70 0.12816
R578 VDD.n76 VDD.n73 0.12816
R579 VDD.n79 VDD.n76 0.12816
R580 VDD.n85 VDD.n82 0.12816
R581 VDD.n88 VDD.n85 0.12816
R582 VDD.n91 VDD.n88 0.12816
R583 VDD.n94 VDD.n91 0.12816
R584 VDD.n97 VDD.n94 0.12816
R585 VDD.n100 VDD.n97 0.12816
R586 VDD.n108 VDD.n105 0.12816
R587 VDD.n102 VDD.n100 0.122257
R588 VDD.n112 VDD.n109 0.119223
R589 VDD.n123 VDD.n120 0.111564
R590 VDD.n124 VDD.n123 0.0936915
R591 VDD.n113 VDD.n112 0.0860319
R592 VDD VDD.n116 0.0687979
R593 VDD VDD.n127 0.0598617
R594 VDD.n105 VDD.n102 0.0515638
R595 VDD.n116 VDD.n113 0.0426277
R596 VDD.n127 VDD.n124 0.0349681
R597 VDD.n109 VDD.n108 0.00943617
R598 SEL.n48 SEL.n38 57.8439
R599 SEL.n39 SEL.t20 51.4916
R600 SEL.n0 SEL.t48 48.0881
R601 SEL.n40 SEL.t2 43.2791
R602 SEL.n41 SEL.t42 43.2791
R603 SEL.n42 SEL.t13 43.2791
R604 SEL.n43 SEL.t49 43.2791
R605 SEL.n0 SEL.t23 34.2844
R606 SEL.n1 SEL.t40 34.2844
R607 SEL.n2 SEL.t18 34.2844
R608 SEL.n3 SEL.t29 34.2844
R609 SEL.n4 SEL.t37 34.2844
R610 SEL.n5 SEL.t15 34.2844
R611 SEL.n6 SEL.t26 34.2844
R612 SEL.n7 SEL.t4 34.2844
R613 SEL.n8 SEL.t19 34.2844
R614 SEL.n9 SEL.t33 34.2844
R615 SEL.n10 SEL.t9 34.2844
R616 SEL.n11 SEL.t17 34.2844
R617 SEL.n12 SEL.t47 34.2844
R618 SEL.n13 SEL.t6 34.2844
R619 SEL.n14 SEL.t21 34.2844
R620 SEL.n15 SEL.t0 34.2844
R621 SEL.n16 SEL.t12 34.2844
R622 SEL.n17 SEL.t36 34.2844
R623 SEL.n18 SEL.t51 34.2844
R624 SEL.n19 SEL.t11 34.2844
R625 SEL.n20 SEL.t43 34.2844
R626 SEL.n21 SEL.t3 34.2844
R627 SEL.n22 SEL.t31 34.2844
R628 SEL.n23 SEL.t39 34.2844
R629 SEL.n24 SEL.t1 34.2844
R630 SEL.n25 SEL.t28 34.2844
R631 SEL.n26 SEL.t50 34.2844
R632 SEL.n27 SEL.t25 34.2844
R633 SEL.n28 SEL.t35 34.2844
R634 SEL.n29 SEL.t46 34.2844
R635 SEL.n30 SEL.t22 34.2844
R636 SEL.n31 SEL.t34 34.2844
R637 SEL.n32 SEL.t32 34.2844
R638 SEL.n33 SEL.t5 34.2844
R639 SEL.n34 SEL.t45 34.2844
R640 SEL.n35 SEL.t14 34.2844
R641 SEL.n36 SEL.t8 34.2844
R642 SEL.n37 SEL.t30 34.2844
R643 SEL.n45 SEL.t24 30.6344
R644 SEL.n39 SEL.t10 30.6344
R645 SEL.n40 SEL.t7 30.6344
R646 SEL.n41 SEL.t41 30.6344
R647 SEL.n42 SEL.t38 30.6344
R648 SEL.n43 SEL.t44 30.6344
R649 SEL.n44 SEL.t27 30.6344
R650 SEL.n38 SEL.t16 30.5041
R651 SEL.n40 SEL.n39 20.8576
R652 SEL.n41 SEL.n40 20.8576
R653 SEL.n42 SEL.n41 20.8576
R654 SEL.n43 SEL.n42 20.8576
R655 SEL.n44 SEL.n43 20.8576
R656 SEL.n45 SEL.n44 20.8576
R657 SEL.n47 SEL.n45 19.6891
R658 SEL.n38 SEL.n37 17.4541
R659 SEL.n1 SEL.n0 13.8041
R660 SEL.n2 SEL.n1 13.8041
R661 SEL.n3 SEL.n2 13.8041
R662 SEL.n4 SEL.n3 13.8041
R663 SEL.n5 SEL.n4 13.8041
R664 SEL.n6 SEL.n5 13.8041
R665 SEL.n7 SEL.n6 13.8041
R666 SEL.n8 SEL.n7 13.8041
R667 SEL.n9 SEL.n8 13.8041
R668 SEL.n10 SEL.n9 13.8041
R669 SEL.n11 SEL.n10 13.8041
R670 SEL.n12 SEL.n11 13.8041
R671 SEL.n13 SEL.n12 13.8041
R672 SEL.n14 SEL.n13 13.8041
R673 SEL.n15 SEL.n14 13.8041
R674 SEL.n16 SEL.n15 13.8041
R675 SEL.n17 SEL.n16 13.8041
R676 SEL.n18 SEL.n17 13.8041
R677 SEL.n19 SEL.n18 13.8041
R678 SEL.n20 SEL.n19 13.8041
R679 SEL.n21 SEL.n20 13.8041
R680 SEL.n22 SEL.n21 13.8041
R681 SEL.n23 SEL.n22 13.8041
R682 SEL.n24 SEL.n23 13.8041
R683 SEL.n25 SEL.n24 13.8041
R684 SEL.n26 SEL.n25 13.8041
R685 SEL.n27 SEL.n26 13.8041
R686 SEL.n28 SEL.n27 13.8041
R687 SEL.n29 SEL.n28 13.8041
R688 SEL.n30 SEL.n29 13.8041
R689 SEL.n31 SEL.n30 13.8041
R690 SEL.n32 SEL.n31 13.8041
R691 SEL.n33 SEL.n32 13.8041
R692 SEL.n34 SEL.n33 13.8041
R693 SEL.n35 SEL.n34 13.8041
R694 SEL.n36 SEL.n35 13.8041
R695 SEL.n37 SEL.n36 13.8041
R696 SEL.n48 SEL.n47 4.0005
R697 SEL.n47 SEL.n46 0.440259
R698 SEL SEL.n48 0.00592169
R699 VSS.n51 VSS.t16 388.923
R700 VSS.n45 VSS.t1 381.221
R701 VSS.n7 VSS.t21 369.668
R702 VSS.n74 VSS.t9 361.967
R703 VSS.n15 VSS.t43 342.714
R704 VSS.n23 VSS.t5 342.714
R705 VSS.n29 VSS.t14 331.161
R706 VSS.n37 VSS.t19 331.161
R707 VSS.n59 VSS.t33 323.461
R708 VSS.n59 VSS.t40 292.654
R709 VSS.n29 VSS.t37 284.954
R710 VSS.n37 VSS.t44 284.954
R711 VSS.n15 VSS.t28 273.401
R712 VSS.n23 VSS.t41 273.401
R713 VSS.n74 VSS.t34 254.148
R714 VSS.n7 VSS.t29 246.446
R715 VSS.n45 VSS.t24 234.893
R716 VSS.n43 VSS.t22 227.192
R717 VSS.n51 VSS.t26 227.192
R718 VSS.n9 VSS.t13 215.641
R719 VSS.n71 VSS.t45 207.939
R720 VSS.n13 VSS.t23 188.685
R721 VSS.n21 VSS.t30 188.685
R722 VSS.n31 VSS.t0 177.133
R723 VSS.n57 VSS.t7 169.431
R724 VSS.n4 VSS.t4 156.946
R725 VSS.n53 VSS.t18 138.626
R726 VSS.n61 VSS.t20 138.626
R727 VSS.n27 VSS.t49 130.924
R728 VSS.n35 VSS.t8 130.924
R729 VSS.n17 VSS.t17 119.373
R730 VSS.n76 VSS.t2 100.118
R731 VSS.n5 VSS.t11 92.4176
R732 VSS.n39 VSS.t12 80.8654
R733 VSS.n47 VSS.t15 80.8654
R734 VSS.n41 VSS.t48 73.164
R735 VSS.n49 VSS.t6 73.164
R736 VSS.n4 VSS.t25 65.306
R737 VSS.n11 VSS.t32 34.6569
R738 VSS.n19 VSS.t39 34.6569
R739 VSS.n25 VSS.t27 23.1048
R740 VSS.n33 VSS.t38 23.1048
R741 VSS.n55 VSS.t42 15.4033
R742 VSS.n63 VSS.t31 15.4033
R743 VSS.n66 VSS.n65 5.2005
R744 VSS.n64 VSS.n63 5.2005
R745 VSS.n62 VSS.n61 5.2005
R746 VSS.n60 VSS.n59 5.2005
R747 VSS.n58 VSS.n57 5.2005
R748 VSS.n56 VSS.n55 5.2005
R749 VSS.n54 VSS.n53 5.2005
R750 VSS.n52 VSS.n51 5.2005
R751 VSS.n50 VSS.n49 5.2005
R752 VSS.n48 VSS.n47 5.2005
R753 VSS.n46 VSS.n45 5.2005
R754 VSS.n44 VSS.n43 5.2005
R755 VSS.n42 VSS.n41 5.2005
R756 VSS.n40 VSS.n39 5.2005
R757 VSS.n38 VSS.n37 5.2005
R758 VSS.n36 VSS.n35 5.2005
R759 VSS.n34 VSS.n33 5.2005
R760 VSS.n32 VSS.n31 5.2005
R761 VSS.n30 VSS.n29 5.2005
R762 VSS.n28 VSS.n27 5.2005
R763 VSS.n26 VSS.n25 5.2005
R764 VSS.n24 VSS.n23 5.2005
R765 VSS.n22 VSS.n21 5.2005
R766 VSS.n20 VSS.n19 5.2005
R767 VSS.n18 VSS.n17 5.2005
R768 VSS.n16 VSS.n15 5.2005
R769 VSS.n14 VSS.n13 5.2005
R770 VSS.n12 VSS.n11 5.2005
R771 VSS.n10 VSS.n9 5.2005
R772 VSS.n8 VSS.n7 5.2005
R773 VSS.n6 VSS.n5 5.2005
R774 VSS.n67 VSS.n3 5.2005
R775 VSS.n78 VSS.n76 5.2005
R776 VSS.n75 VSS.n74 5.2005
R777 VSS.n72 VSS.n71 5.2005
R778 VSS.n69 VSS.n68 5.2005
R779 VSS.n70 VSS.n2 4.48602
R780 VSS.n77 VSS.t3 4.48602
R781 VSS.n73 VSS.n1 3.66702
R782 VSS.n6 VSS.n4 1.62155
R783 VSS.n1 VSS.t10 0.8195
R784 VSS.n1 VSS.n0 0.8195
R785 VSS.n12 VSS.n10 0.167855
R786 VSS.n26 VSS.n24 0.167855
R787 VSS.n40 VSS.n38 0.167855
R788 VSS.n54 VSS.n52 0.167855
R789 VSS.n67 VSS.n66 0.149347
R790 VSS.n8 VSS.n6 0.14926
R791 VSS.n10 VSS.n8 0.14926
R792 VSS.n14 VSS.n12 0.14926
R793 VSS.n16 VSS.n14 0.14926
R794 VSS.n18 VSS.n16 0.14926
R795 VSS.n20 VSS.n18 0.14926
R796 VSS.n22 VSS.n20 0.14926
R797 VSS.n24 VSS.n22 0.14926
R798 VSS.n28 VSS.n26 0.14926
R799 VSS.n30 VSS.n28 0.14926
R800 VSS.n32 VSS.n30 0.14926
R801 VSS.n34 VSS.n32 0.14926
R802 VSS.n36 VSS.n34 0.14926
R803 VSS.n38 VSS.n36 0.14926
R804 VSS.n42 VSS.n40 0.14926
R805 VSS.n44 VSS.n42 0.14926
R806 VSS.n46 VSS.n44 0.14926
R807 VSS.n48 VSS.n46 0.14926
R808 VSS.n50 VSS.n48 0.14926
R809 VSS.n52 VSS.n50 0.14926
R810 VSS.n56 VSS.n54 0.14926
R811 VSS.n58 VSS.n56 0.14926
R812 VSS.n60 VSS.n58 0.14926
R813 VSS.n62 VSS.n60 0.14926
R814 VSS.n64 VSS.n62 0.14926
R815 VSS.n66 VSS.n64 0.14926
R816 VSS.n73 VSS.n72 0.132311
R817 VSS.n69 VSS.n67 0.116167
R818 VSS.n72 VSS.n70 0.0954606
R819 VSS.n78 VSS.n77 0.0756181
R820 VSS VSS.n75 0.0742008
R821 VSS VSS.n78 0.0685315
R822 VSS.n70 VSS.n69 0.0472717
R823 VSS.n75 VSS.n73 0.0104213
C0 VDD SEL 1.36f
C1 IN VDD 5.83f
C2 OUT SEL 1.33f
C3 IN OUT 18.1f
C4 OUT VDD 0.321f
C5 IN SEL 0.933f
.ends

