magic
tech gf180mcuC
magscale 1 10
timestamp 1690971400
<< error_p >>
rect -34 781 -23 827
rect 23 781 34 792
rect -80 550 -57 561
rect 57 550 80 561
rect -34 469 -23 515
rect -34 349 -23 395
rect 23 349 34 360
rect -80 118 -57 129
rect 57 118 80 129
rect -34 37 -23 83
rect -34 -83 -23 -37
rect 23 -83 34 -72
rect -80 -314 -57 -303
rect 57 -314 80 -303
rect -34 -395 -23 -349
rect -34 -515 -23 -469
rect 23 -515 34 -504
rect -80 -746 -57 -735
rect 57 -746 80 -735
rect -34 -827 -23 -781
<< nwell >>
rect -278 -956 278 956
<< pmos >>
rect -28 548 28 748
rect -28 116 28 316
rect -28 -316 28 -116
rect -28 -748 28 -548
<< pdiff >>
rect -116 735 -28 748
rect -116 561 -103 735
rect -57 561 -28 735
rect -116 548 -28 561
rect 28 735 116 748
rect 28 561 57 735
rect 103 561 116 735
rect 28 548 116 561
rect -116 303 -28 316
rect -116 129 -103 303
rect -57 129 -28 303
rect -116 116 -28 129
rect 28 303 116 316
rect 28 129 57 303
rect 103 129 116 303
rect 28 116 116 129
rect -116 -129 -28 -116
rect -116 -303 -103 -129
rect -57 -303 -28 -129
rect -116 -316 -28 -303
rect 28 -129 116 -116
rect 28 -303 57 -129
rect 103 -303 116 -129
rect 28 -316 116 -303
rect -116 -561 -28 -548
rect -116 -735 -103 -561
rect -57 -735 -28 -561
rect -116 -748 -28 -735
rect 28 -561 116 -548
rect 28 -735 57 -561
rect 103 -735 116 -561
rect 28 -748 116 -735
<< pdiffc >>
rect -103 561 -57 735
rect 57 561 103 735
rect -103 129 -57 303
rect 57 129 103 303
rect -103 -303 -57 -129
rect 57 -303 103 -129
rect -103 -735 -57 -561
rect 57 -735 103 -561
<< nsubdiff >>
rect -254 860 254 932
rect -254 816 -182 860
rect -254 -816 -241 816
rect -195 -816 -182 816
rect 182 816 254 860
rect -254 -860 -182 -816
rect 182 -816 195 816
rect 241 -816 254 816
rect 182 -860 254 -816
rect -254 -932 254 -860
<< nsubdiffcont >>
rect -241 -816 -195 816
rect 195 -816 241 816
<< polysilicon >>
rect -36 827 36 840
rect -36 781 -23 827
rect 23 781 36 827
rect -36 768 36 781
rect -28 748 28 768
rect -28 528 28 548
rect -36 515 36 528
rect -36 469 -23 515
rect 23 469 36 515
rect -36 456 36 469
rect -36 395 36 408
rect -36 349 -23 395
rect 23 349 36 395
rect -36 336 36 349
rect -28 316 28 336
rect -28 96 28 116
rect -36 83 36 96
rect -36 37 -23 83
rect 23 37 36 83
rect -36 24 36 37
rect -36 -37 36 -24
rect -36 -83 -23 -37
rect 23 -83 36 -37
rect -36 -96 36 -83
rect -28 -116 28 -96
rect -28 -336 28 -316
rect -36 -349 36 -336
rect -36 -395 -23 -349
rect 23 -395 36 -349
rect -36 -408 36 -395
rect -36 -469 36 -456
rect -36 -515 -23 -469
rect 23 -515 36 -469
rect -36 -528 36 -515
rect -28 -548 28 -528
rect -28 -768 28 -748
rect -36 -781 36 -768
rect -36 -827 -23 -781
rect 23 -827 36 -781
rect -36 -840 36 -827
<< polycontact >>
rect -23 781 23 827
rect -23 469 23 515
rect -23 349 23 395
rect -23 37 23 83
rect -23 -83 23 -37
rect -23 -395 23 -349
rect -23 -515 23 -469
rect -23 -827 23 -781
<< metal1 >>
rect -241 873 241 919
rect -241 816 -195 873
rect -34 781 -23 827
rect 23 781 34 827
rect 195 816 241 873
rect -103 735 -57 746
rect -103 550 -57 561
rect 57 735 103 746
rect 57 550 103 561
rect -34 469 -23 515
rect 23 469 34 515
rect -34 349 -23 395
rect 23 349 34 395
rect -103 303 -57 314
rect -103 118 -57 129
rect 57 303 103 314
rect 57 118 103 129
rect -34 37 -23 83
rect 23 37 34 83
rect -34 -83 -23 -37
rect 23 -83 34 -37
rect -103 -129 -57 -118
rect -103 -314 -57 -303
rect 57 -129 103 -118
rect 57 -314 103 -303
rect -34 -395 -23 -349
rect 23 -395 34 -349
rect -34 -515 -23 -469
rect 23 -515 34 -469
rect -103 -561 -57 -550
rect -103 -746 -57 -735
rect 57 -561 103 -550
rect 57 -746 103 -735
rect -241 -873 -195 -816
rect -34 -827 -23 -781
rect 23 -827 34 -781
rect 195 -873 241 -816
rect -241 -919 241 -873
<< properties >>
string FIXED_BBOX -218 -896 218 896
string gencell pmos_3p3
string library gf180mcu
string parameters w 1 l 0.280 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 1 compatible {pmos_3p3 pmos_6p0}
<< end >>
