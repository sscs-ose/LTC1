magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2088 -2044 2960 2644
<< mvnmos >>
rect 0 0 140 600
rect 244 0 384 600
rect 488 0 628 600
rect 732 0 872 600
<< mvndiff >>
rect -88 587 0 600
rect -88 541 -75 587
rect -29 541 0 587
rect -88 482 0 541
rect -88 436 -75 482
rect -29 436 0 482
rect -88 377 0 436
rect -88 331 -75 377
rect -29 331 0 377
rect -88 271 0 331
rect -88 225 -75 271
rect -29 225 0 271
rect -88 165 0 225
rect -88 119 -75 165
rect -29 119 0 165
rect -88 59 0 119
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 140 587 244 600
rect 140 541 169 587
rect 215 541 244 587
rect 140 482 244 541
rect 140 436 169 482
rect 215 436 244 482
rect 140 377 244 436
rect 140 331 169 377
rect 215 331 244 377
rect 140 271 244 331
rect 140 225 169 271
rect 215 225 244 271
rect 140 165 244 225
rect 140 119 169 165
rect 215 119 244 165
rect 140 59 244 119
rect 140 13 169 59
rect 215 13 244 59
rect 140 0 244 13
rect 384 587 488 600
rect 384 541 413 587
rect 459 541 488 587
rect 384 482 488 541
rect 384 436 413 482
rect 459 436 488 482
rect 384 377 488 436
rect 384 331 413 377
rect 459 331 488 377
rect 384 271 488 331
rect 384 225 413 271
rect 459 225 488 271
rect 384 165 488 225
rect 384 119 413 165
rect 459 119 488 165
rect 384 59 488 119
rect 384 13 413 59
rect 459 13 488 59
rect 384 0 488 13
rect 628 587 732 600
rect 628 541 657 587
rect 703 541 732 587
rect 628 482 732 541
rect 628 436 657 482
rect 703 436 732 482
rect 628 377 732 436
rect 628 331 657 377
rect 703 331 732 377
rect 628 271 732 331
rect 628 225 657 271
rect 703 225 732 271
rect 628 165 732 225
rect 628 119 657 165
rect 703 119 732 165
rect 628 59 732 119
rect 628 13 657 59
rect 703 13 732 59
rect 628 0 732 13
rect 872 587 960 600
rect 872 541 901 587
rect 947 541 960 587
rect 872 482 960 541
rect 872 436 901 482
rect 947 436 960 482
rect 872 377 960 436
rect 872 331 901 377
rect 947 331 960 377
rect 872 271 960 331
rect 872 225 901 271
rect 947 225 960 271
rect 872 165 960 225
rect 872 119 901 165
rect 947 119 960 165
rect 872 59 960 119
rect 872 13 901 59
rect 947 13 960 59
rect 872 0 960 13
<< mvndiffc >>
rect -75 541 -29 587
rect -75 436 -29 482
rect -75 331 -29 377
rect -75 225 -29 271
rect -75 119 -29 165
rect -75 13 -29 59
rect 169 541 215 587
rect 169 436 215 482
rect 169 331 215 377
rect 169 225 215 271
rect 169 119 215 165
rect 169 13 215 59
rect 413 541 459 587
rect 413 436 459 482
rect 413 331 459 377
rect 413 225 459 271
rect 413 119 459 165
rect 413 13 459 59
rect 657 541 703 587
rect 657 436 703 482
rect 657 331 703 377
rect 657 225 703 271
rect 657 119 703 165
rect 657 13 703 59
rect 901 541 947 587
rect 901 436 947 482
rect 901 331 947 377
rect 901 225 947 271
rect 901 119 947 165
rect 901 13 947 59
<< polysilicon >>
rect 0 600 140 644
rect 244 600 384 644
rect 488 600 628 644
rect 732 600 872 644
rect 0 -44 140 0
rect 244 -44 384 0
rect 488 -44 628 0
rect 732 -44 872 0
<< metal1 >>
rect -75 587 -29 600
rect -75 482 -29 541
rect -75 377 -29 436
rect -75 271 -29 331
rect -75 165 -29 225
rect -75 59 -29 119
rect -75 0 -29 13
rect 169 587 215 600
rect 169 482 215 541
rect 169 377 215 436
rect 169 271 215 331
rect 169 165 215 225
rect 169 59 215 119
rect 169 0 215 13
rect 413 587 459 600
rect 413 482 459 541
rect 413 377 459 436
rect 413 271 459 331
rect 413 165 459 225
rect 413 59 459 119
rect 413 0 459 13
rect 657 587 703 600
rect 657 482 703 541
rect 657 377 703 436
rect 657 271 703 331
rect 657 165 703 225
rect 657 59 703 119
rect 657 0 703 13
rect 901 587 947 600
rect 901 482 947 541
rect 901 377 947 436
rect 901 271 947 331
rect 901 165 947 225
rect 901 59 947 119
rect 901 0 947 13
<< labels >>
rlabel metal1 680 300 680 300 4 S
rlabel metal1 436 300 436 300 4 D
rlabel metal1 192 300 192 300 4 S
rlabel metal1 924 300 924 300 4 D
rlabel metal1 -52 300 -52 300 4 D
<< end >>
