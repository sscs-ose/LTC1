magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1071 -1695 1071 1695
<< metal1 >>
rect -71 689 71 695
rect -71 -689 -65 689
rect 65 -689 71 689
rect -71 -695 71 -689
<< via1 >>
rect -65 -689 65 689
<< metal2 >>
rect -71 689 71 695
rect -71 -689 -65 689
rect 65 -689 71 689
rect -71 -695 71 -689
<< end >>
