magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -4395 -2045 4395 2045
<< ndiff >>
rect -2395 23 2395 45
rect -2395 -23 -2373 23
rect 2373 -23 2395 23
rect -2395 -45 2395 -23
<< ndiffc >>
rect -2373 -23 2373 23
<< metal1 >>
rect -2384 23 2384 34
rect -2384 -23 -2373 23
rect 2373 -23 2384 23
rect -2384 -34 2384 -23
<< end >>
