magic
tech gf180mcuC
magscale 1 10
timestamp 1695109904
<< nwell >>
rect 1912 890 2133 892
rect 3801 890 3944 891
rect 1912 888 3944 890
rect 928 835 1020 842
rect 928 773 1021 835
rect 1912 830 3945 888
rect 1764 805 1855 809
rect 1764 773 1856 805
rect 928 771 1856 773
rect 929 720 1856 771
rect 952 715 1856 720
rect 380 654 744 670
rect 531 609 616 654
rect 489 606 616 609
rect 531 600 616 606
rect 380 574 743 600
rect 952 578 1001 715
rect 1912 658 1973 830
rect 2267 828 3945 830
rect 3776 775 3945 828
rect 2036 774 2127 775
rect 2035 771 2127 774
rect 2035 715 2258 771
rect 2035 685 2127 715
rect 2035 684 2126 685
rect 1442 607 1613 657
rect 531 563 616 574
rect 952 553 1000 578
rect 1417 575 1613 607
rect 1835 600 1973 658
rect 2466 625 2539 637
rect 2320 622 3358 625
rect 2466 612 2539 622
rect 2421 607 2539 612
rect 1417 564 1582 575
rect 2466 566 2539 607
rect 3245 608 3359 616
rect 3416 608 3510 632
rect 3841 613 3900 775
rect 3245 599 3510 608
rect 3245 589 3359 599
rect 3416 589 3510 599
rect 3245 566 3510 589
rect -384 517 -254 520
rect 952 519 953 553
rect 1417 551 1505 564
rect 3245 556 3462 566
rect 3245 542 3359 556
<< pwell >>
rect 3822 482 3852 490
rect 3822 433 3837 482
rect 4091 395 4190 409
rect 4074 394 4190 395
rect 836 330 888 382
rect 4072 374 4190 394
rect 4071 331 4190 374
rect 4071 316 4189 331
<< ndiff >>
rect 836 330 888 382
<< pdiff >>
rect 1781 727 1837 785
rect 2051 700 2107 759
<< psubdiff >>
rect 3851 163 3892 242
<< nsubdiff >>
rect 3848 949 3895 1021
<< metal1 >>
rect 1870 920 2080 1020
rect 928 835 1020 842
rect 3835 835 3912 842
rect 928 834 1021 835
rect 928 779 950 834
rect 1003 779 1021 834
rect 928 771 1021 779
rect 3835 783 3847 835
rect 3899 783 3912 835
rect 3835 775 3912 783
rect 531 647 616 670
rect 531 609 550 647
rect 489 606 550 609
rect 531 593 550 606
rect 603 593 616 647
rect 531 563 616 593
rect -389 516 -254 542
rect -389 464 -361 516
rect -304 464 -254 516
rect 132 512 213 522
rect -389 452 -254 464
rect -134 508 213 512
rect -134 456 146 508
rect 132 453 146 456
rect 200 453 213 508
rect 132 442 213 453
rect 952 510 1001 771
rect 2204 650 2261 749
rect 1492 638 1582 649
rect 1492 624 1511 638
rect 1476 607 1511 624
rect 1417 585 1511 607
rect 1564 585 1582 638
rect 1417 564 1582 585
rect 2203 647 2261 650
rect 1417 551 1505 564
rect 2054 510 2146 521
rect 952 452 1167 510
rect 2054 458 2083 510
rect 2135 458 2146 510
rect 2054 452 2146 458
rect 2203 448 2260 647
rect 2466 628 2539 637
rect 2466 612 2479 628
rect 2421 607 2479 612
rect 2466 576 2479 607
rect 2531 576 2539 628
rect 3416 627 3510 632
rect 3416 608 3439 627
rect 2466 566 2539 576
rect 3313 574 3439 608
rect 3492 574 3510 627
rect 3313 566 3510 574
rect 3313 551 3436 566
rect 3841 539 3900 775
rect 3829 535 3900 539
rect 3829 505 3958 535
rect 3826 482 3958 505
rect 3826 430 3838 482
rect 3891 456 3958 482
rect 4013 529 4080 544
rect 4013 468 4024 529
rect 4076 468 4080 529
rect 3891 430 3903 456
rect 4013 454 4080 468
rect 3829 425 3902 430
rect 3829 424 3888 425
rect 810 382 922 396
rect 4091 395 4190 409
rect 4074 394 4190 395
rect 810 330 836 382
rect 888 330 922 382
rect 810 315 922 330
rect 1770 380 1886 392
rect 1770 327 1798 380
rect 1852 327 1886 380
rect 1770 312 1886 327
rect 2737 375 2856 389
rect 2737 322 2766 375
rect 2820 322 2856 375
rect 2737 310 2856 322
rect 3666 383 3773 394
rect 3666 328 3688 383
rect 3743 328 3773 383
rect 4072 380 4190 394
rect 4072 374 4094 380
rect 3666 314 3773 328
rect 4071 328 4094 374
rect 4146 331 4190 380
rect 4146 328 4189 331
rect 4071 316 4189 328
rect -377 75 -286 88
rect -377 8 -362 75
rect -299 8 -286 75
rect -377 -5 -286 8
rect -29 0 22 261
rect 788 76 900 89
rect 788 23 817 76
rect 871 23 900 76
rect 788 10 900 23
rect 948 0 998 260
rect 1732 79 1849 91
rect 1732 26 1759 79
rect 1813 26 1849 79
rect 1732 10 1849 26
rect 1918 4 1968 264
rect 2351 17 2535 101
rect 2704 80 2823 96
rect 2704 27 2734 80
rect 2788 27 2823 80
rect 2704 17 2823 27
rect 2882 2 2932 262
rect 3851 163 3892 242
rect 3674 82 3793 95
rect 3674 29 3704 82
rect 3758 29 3793 82
rect 3674 16 3793 29
rect 4010 80 4087 89
rect 4010 20 4020 80
rect 4078 20 4087 80
rect 4010 10 4087 20
<< via1 >>
rect 950 779 1003 834
rect 3847 783 3899 835
rect 550 593 603 647
rect -361 464 -304 516
rect 146 453 200 508
rect 1511 585 1564 638
rect 2083 458 2135 510
rect 2479 576 2531 628
rect 3439 574 3492 627
rect 3048 457 3101 509
rect 3838 430 3891 482
rect 4024 468 4076 529
rect 836 330 888 382
rect 1798 327 1852 380
rect 2766 322 2820 375
rect 3688 328 3743 383
rect 4094 328 4146 380
rect -362 8 -299 75
rect 817 23 871 76
rect 1759 26 1813 79
rect 2734 27 2788 80
rect 3704 29 3758 82
rect 4020 20 4078 80
<< metal2 >>
rect -222 837 1020 895
rect -376 519 -292 520
rect -222 519 -166 837
rect 928 835 1020 837
rect 1912 890 2133 892
rect 3801 890 3944 891
rect 1912 888 3944 890
rect 1912 835 3945 888
rect 928 834 1021 835
rect 928 779 950 834
rect 1003 779 1021 834
rect 1912 830 3847 835
rect 928 773 1021 779
rect 1765 785 1856 805
rect 1765 773 1781 785
rect 928 771 1781 773
rect 929 727 1781 771
rect 1837 727 1856 785
rect 929 720 1856 727
rect 986 715 1856 720
rect 380 657 744 670
rect 1912 658 1973 830
rect 2267 828 3847 830
rect 3776 783 3847 828
rect 3899 783 3945 835
rect 3776 775 3945 783
rect 2035 771 2126 774
rect 2035 759 2258 771
rect 2035 700 2051 759
rect 2107 749 2258 759
rect 2107 715 2261 749
rect 2107 700 2126 715
rect 2035 684 2126 700
rect 1835 657 1973 658
rect 380 647 1973 657
rect 2204 650 2261 715
rect 380 593 550 647
rect 603 638 1973 647
rect 603 600 1511 638
rect 603 593 743 600
rect 380 574 743 593
rect 1442 585 1511 600
rect 1564 600 1973 638
rect 2203 647 2261 650
rect 1564 585 1613 600
rect 1442 575 1613 585
rect 1472 574 1582 575
rect -376 516 -166 519
rect -376 464 -361 516
rect -304 464 -166 516
rect -376 453 -166 464
rect -369 88 -298 453
rect -222 452 -166 453
rect 132 518 213 522
rect 2049 518 2146 523
rect 132 517 1881 518
rect 2005 517 2146 518
rect 132 510 2146 517
rect 132 508 2083 510
rect 132 453 146 508
rect 200 458 2083 508
rect 2135 458 2146 510
rect 200 453 2146 458
rect 132 452 2146 453
rect 132 442 213 452
rect 2049 443 2146 452
rect 2203 508 2260 647
rect 2466 628 2539 637
rect 2466 625 2479 628
rect 2320 576 2479 625
rect 2531 625 2539 628
rect 3416 627 3510 632
rect 2531 616 3358 625
rect 2531 603 3359 616
rect 3416 603 3439 627
rect 2531 576 3439 603
rect 2320 574 3439 576
rect 3492 603 3510 627
rect 3492 574 4100 603
rect 2320 568 4100 574
rect 2320 566 2490 568
rect 3245 546 4100 568
rect 3245 542 3359 546
rect 4012 544 4100 546
rect 4012 529 4101 544
rect 3031 509 3138 511
rect 3031 508 3048 509
rect 2203 457 3048 508
rect 3101 457 3138 509
rect 2203 449 3138 457
rect 2203 448 2260 449
rect 3031 443 3138 449
rect 3822 482 3948 490
rect 3822 430 3838 482
rect 3891 433 3948 482
rect 4012 468 4024 529
rect 4076 518 4101 529
rect 4216 518 4274 519
rect 4076 468 4274 518
rect 4012 454 4274 468
rect 3891 430 3900 433
rect 3822 424 3900 430
rect 809 382 922 396
rect 809 330 836 382
rect 888 330 922 382
rect 809 315 922 330
rect 1770 380 1886 392
rect 1770 327 1798 380
rect 1852 327 1886 380
rect 828 89 888 315
rect 1770 312 1886 327
rect 2737 375 2856 389
rect 2737 322 2766 375
rect 2820 322 2856 375
rect 1792 91 1849 312
rect 2737 310 2856 322
rect 3666 383 3773 394
rect 3666 328 3688 383
rect 3743 328 3773 383
rect 3666 314 3773 328
rect 3829 374 3900 424
rect 4072 380 4158 398
rect 4072 374 4094 380
rect 3829 328 4094 374
rect 4146 328 4158 380
rect 3829 315 4158 328
rect 2750 96 2807 310
rect -377 75 -286 88
rect -377 8 -362 75
rect -299 8 -286 75
rect 788 76 900 89
rect 788 23 817 76
rect 871 23 900 76
rect 788 10 900 23
rect 1732 79 1849 91
rect 1732 26 1759 79
rect 1813 26 1849 79
rect 1732 10 1849 26
rect 2704 80 2823 96
rect 3703 95 3760 314
rect 2704 27 2734 80
rect 2788 27 2823 80
rect 2704 16 2823 27
rect 3674 82 3793 95
rect 3674 29 3704 82
rect 3758 29 3793 82
rect 3674 16 3793 29
rect 4010 81 4087 89
rect 4216 81 4274 454
rect 4010 80 4274 81
rect 4010 20 4020 80
rect 4078 20 4274 80
rect 4010 17 4274 20
rect 4010 10 4087 17
rect -377 -5 -286 8
<< via2 >>
rect 1781 727 1837 785
rect 2051 700 2107 759
<< metal3 >>
rect 1764 785 1855 809
rect 1764 727 1781 785
rect 1837 773 1855 785
rect 2036 773 2127 775
rect 1837 759 2127 773
rect 1837 727 2051 759
rect 1764 719 2051 727
rect 1784 716 2051 719
rect 2036 700 2051 716
rect 2107 700 2127 759
rect 2036 685 2127 700
use and_2_ibr  and_2_ibr_0
timestamp 1695109904
transform 1 0 -257 0 1 -996
box 257 996 1231 2047
use and_2_ibr  and_2_ibr_1
timestamp 1695109904
transform 1 0 709 0 1 -995
box 257 996 1231 2047
use and_2_ibr  and_2_ibr_2
timestamp 1695109904
transform 1 0 1675 0 1 -995
box 257 996 1231 2047
use and_2_ibr  and_2_ibr_3
timestamp 1695109904
transform 1 0 2641 0 1 -995
box 257 996 1231 2047
use nand2  nand2_0 ~/GF180Projects/Top_test/top/magic
timestamp 1694691991
transform 1 0 70 0 1 188
box -70 -188 502 863
use nand2  nand2_1
timestamp 1694691991
transform 1 0 1036 0 1 189
box -70 -188 502 863
use nand2  nand2_2
timestamp 1694691991
transform 1 0 2002 0 1 189
box -70 -188 502 863
use nand2  nand2_3
timestamp 1694691991
transform 1 0 2968 0 1 189
box -70 -188 502 863
use nverterlayout_ibr  nverterlayout_ibr_0 ~/GF180Projects/Top_test/top/magic
timestamp 1695109904
transform 1 0 -308 0 1 -79
box -88 220 316 1130
use nverterlayout_ibr  nverterlayout_ibr_1
timestamp 1695109904
transform 1 0 3959 0 1 -78
box -88 220 316 1130
<< labels >>
flabel via1 -331 38 -331 38 0 FreeSans 480 0 0 0 IN1
port 1 nsew
flabel via1 4046 46 4046 46 0 FreeSans 480 0 0 0 IN2
port 2 nsew
flabel via1 845 50 845 50 0 FreeSans 480 0 0 0 D0
port 3 nsew
flabel via1 1786 42 1786 42 0 FreeSans 480 0 0 0 D1
port 4 nsew
flabel via1 2761 50 2761 50 0 FreeSans 480 0 0 0 D2
port 5 nsew
flabel via1 3729 50 3729 50 0 FreeSans 480 0 0 0 D3
port 6 nsew
flabel metal1 2436 63 2436 63 0 FreeSans 480 0 0 0 VSS
port 7 nsew
flabel metal1 1978 970 1978 970 0 FreeSans 480 0 0 0 VDD
port 8 nsew
<< end >>
