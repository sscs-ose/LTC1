* NGSPICE file created from CLK_div_110_mag_flat.ext - technology: gf180mcuC

.subckt CLK_div_110_mag_flat RST CLK Vdiv110 VSS VDD
X0 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN VSS.t282 VSS.t167 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X1 Vdiv110 CLK_div_10_mag_0.Q3 a_12478_n2129# VDD.t162 pfet_03v3 ad=1.06p pd=5.68u as=0.624p ps=2.92u w=2.4u l=0.28u
X2 VDD CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.Q0 VDD.t467 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q2 a_n1595_3762# VSS.t266 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X4 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_DIV_11_mag_new_0.Q3 a_9506_4996# VDD.t415 pfet_03v3 ad=1.06p pd=5.68u as=0.624p ps=2.92u w=2.4u l=0.28u
X5 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.Q2 a_9414_759# VSS.t40 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X6 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_2874_2775# VSS.t236 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X7 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t164 VDD.t163 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X8 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t148 VSS.t147 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X9 a_11143_759# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t146 VSS.t145 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X10 VDD CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VDD.t152 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X11 VDD CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.QB VDD.t182 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X12 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD.t268 VDD.t270 VDD.t269 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X13 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_2310_2775# VSS.t245 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X14 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 a_n358_4884# VDD.t243 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X15 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_10_mag_0.Q3 VDD.t161 VDD.t160 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X16 a_2874_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t241 VSS.t240 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X17 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q0 VDD.t26 VDD.t25 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X18 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t491 VDD.t490 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X19 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_0.and2_mag_1.OUT VSS.t284 VSS.t283 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X20 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t483 VDD.t482 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X21 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_10_mag_0.Q0 a_1528_759# VSS.t15 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X22 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD.t156 VDD.t155 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X23 a_5904_4934# CLK_DIV_11_mag_new_0.Q0 a_5744_4934# VSS.t88 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X24 VDD RST.t0 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t387 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X25 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK.t0 VDD.t41 VDD.t40 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X26 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.K VDD.t283 VDD.t282 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X27 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_5833_759# VSS.t275 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X28 VDD CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t142 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X29 a_3380_759# CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t30 VSS.t29 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X30 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t475 VDD.t474 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X31 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t132 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X32 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q2 VDD.t431 VDD.t430 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X33 a_9123_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS.t46 VSS.t45 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X34 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t487 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X35 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t343 VDD.t342 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X36 a_12436_1674# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS.t110 VSS.t109 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X37 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_8713_1678# VSS.t135 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X38 a_5035_1632# RST.t1 a_4875_1632# VSS.t237 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X39 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK.t1 a_5904_4934# VSS.t26 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X40 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN VSS.t312 VSS.t311 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X41 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 VSS.t286 VSS.t285 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X42 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q3 a_n1762_4447# VSS.t253 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X43 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t479 VDD.t478 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X44 a_1016_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_0.K VSS.t162 VSS.t66 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X45 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_3.QB a_7568_n338# VSS.t126 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X46 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK.t2 VSS.t28 VSS.t27 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X47 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VDD.t126 VDD.t125 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X48 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_5269_759# VSS.t59 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X49 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q2 a_4311_1632# VSS.t265 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X50 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t99 VDD.t98 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X51 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t464 VDD.t463 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X52 a_4875_1632# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t205 VSS.t204 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X53 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS.t203 VSS.t202 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X54 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_8696_n338# VSS.t63 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X55 a_10419_759# VDD.t492 VSS.t92 VSS.t91 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X56 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_0.and2_mag_1.OUT VDD.t455 VDD.t454 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X57 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.Q0 VSS.t14 VSS.t13 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X58 a_7568_n338# CLK_div_10_mag_0.Q1 a_7408_n338# VSS.t117 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X59 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 a_5035_1632# VSS.t304 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X60 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.JK_FF_mag_2.K.t3 a_12277_n338# VSS.t19 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X61 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD.t49 VDD.t48 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X62 a_11149_n338# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t190 VSS.t19 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X63 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK.t3 VDD.t43 VDD.t42 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X64 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_8132_n338# VSS.t33 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X65 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.K VDD.t281 VDD.t280 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X66 VDD CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD.t22 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X67 CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VSS.t306 VSS.t305 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X68 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_3.QB VDD.t209 VDD.t208 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X69 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.Q3 a_12431_759# VSS.t106 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X70 a_11718_2771# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS.t232 VSS.t231 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X71 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VSS.t75 VSS.t74 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X72 a_8286_759# RST.t2 a_8126_759# VSS.t238 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X73 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t39 VDD.t38 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X74 a_12277_n338# CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t20 VSS.t19 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X75 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT VDD.t84 VDD.t83 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X76 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_4317_2729# VSS.t220 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X77 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_12282_2771# VSS.t187 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X78 a_3226_n338# CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t199 VSS.t198 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X79 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t307 VDD.t306 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X80 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD.t109 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X81 a_11154_2771# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VSS.t22 VSS.t21 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X82 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT VDD.t89 VDD.t88 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X83 a_1022_2731# CLK_DIV_11_mag_new_0.JK_FF_mag_0.K VSS.t161 VSS.t160 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X84 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.QB a_4551_n338# VSS.t175 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X85 VDD CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD.t179 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X86 VDD CLK.t4 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT VDD.t194 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X87 VDD CLK_div_10_mag_0.JK_FF_mag_2.K.t4 CLK_div_10_mag_0.Q3 VDD.t185 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X88 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t323 VDD.t322 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X89 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t46 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X90 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD.t265 VDD.t267 VDD.t266 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X91 a_12282_2771# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS.t197 VSS.t196 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X92 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.Q0 a_3380_759# VSS.t12 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X93 a_7989_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT VSS.t48 VSS.t47 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X94 VDD RST.t3 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD.t390 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X95 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 a_8149_1634# VSS.t180 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X96 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q1 a_9282_n1435# VSS.t37 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X97 a_1746_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t301 VSS.t300 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X98 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_5599_1676# VSS.t78 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X99 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t33 VDD.t32 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X100 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.K VDD.t473 VDD.t472 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X101 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t341 VDD.t340 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X102 CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD.t303 VDD.t302 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X103 a_7425_1634# CLK.t5 a_7265_1634# VSS.t123 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X104 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.Q0 VDD.t21 VDD.t20 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X105 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t337 VDD.t336 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X106 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_5115_n338# VSS.t157 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X107 VDD CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.QB VDD.t70 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X108 a_9506_4996# CLK_DIV_11_mag_new_0.and2_mag_3.OUT a_9346_4996# VDD.t422 pfet_03v3 ad=0.624p pd=2.92u as=0.624p ps=2.92u w=2.4u l=0.28u
X109 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK.t6 VDD.t198 VDD.t197 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X110 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.QB VDD.t301 VDD.t300 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X111 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t240 VDD.t239 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X112 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q2 a_8314_n1435# VSS.t37 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X113 Vdiv110 CLK_div_10_mag_0.nor_3_mag_0.IN3 VSS.t201 VSS.t200 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X114 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t3 VDD.t128 VDD.t127 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X115 CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS.t177 VSS.t176 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X116 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_8850_759# VSS.t62 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X117 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT VDD.t421 VDD.t420 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X118 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.and2_mag_3.IN1 VDD.t348 VDD.t347 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X119 a_6397_759# CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS.t137 VSS.t136 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X120 a_7265_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_2.K VSS.t299 VSS.t298 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X121 a_n1755_2260# CLK_DIV_11_mag_new_0.Q1 VSS.t218 VSS.t217 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X122 a_2310_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t56 VSS.t55 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X123 CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS.t247 VSS.t246 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X124 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_10_mag_0.Q1 a_4545_759# VSS.t116 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X125 a_2092_759# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t243 VSS.t242 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X126 VDD CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VDD.t344 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X127 VDD CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t176 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X128 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD.t93 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X129 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_1.QB a_1534_n338# VSS.t295 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X130 a_11867_759# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t80 VSS.t79 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X131 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q0 VDD.t151 VDD.t150 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X132 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t275 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X133 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_10_mag_0.Q0 VDD.t19 VDD.t18 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X134 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t4 a_7431_2731# VSS.t76 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X135 a_5744_4934# CLK_DIV_11_mag_new_0.and2_mag_3.IN1 VSS.t208 VSS.t207 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X136 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t379 VDD.t378 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X137 VDD CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t67 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X138 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_8286_759# VSS.t256 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X139 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD.t443 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X140 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VDD.t296 VDD.t295 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X141 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN VDD.t453 VDD.t452 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X142 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t45 VDD.t44 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X143 VDD CLK.t7 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT VDD.t199 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X144 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t234 VDD.t233 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X145 a_7562_759# CLK_div_10_mag_0.Q1 a_7402_759# VSS.t115 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X146 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q0 a_10584_1630# VSS.t87 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X147 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.Q2 VDD.t429 VDD.t428 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X148 VDD CLK.t8 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t202 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X149 a_2816_759# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t18 VSS.t17 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X150 a_8713_1678# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT VSS.t51 VSS.t50 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X151 VDD CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB VDD.t425 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X152 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_1.QB VDD.t466 VDD.t465 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X153 CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS.t133 VSS.t132 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X154 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB VDD.t319 VDD.t318 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X155 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q1 VDD.t363 VDD.t351 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X156 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 a_11308_1630# VSS.t230 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X157 a_n1755_3762# CLK_DIV_11_mag_new_0.Q1 VSS.t216 VSS.t215 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X158 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.Q2 VSS.t264 VSS.t263 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X159 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t273 VSS.t272 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X160 a_10584_1630# CLK.t9 a_10424_1630# VSS.t124 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X161 CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD.t404 VDD.t403 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X162 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t103 VDD.t102 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X163 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK.t10 VSS.t70 VSS.t69 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X164 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t230 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X165 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD.t90 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X166 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t222 VSS.t221 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X167 a_4311_1632# CLK.t11 a_4151_1632# VSS.t71 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X168 a_11303_759# RST.t4 a_11143_759# VSS.t239 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X169 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t285 VDD.t284 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X170 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK.t12 VDD.t121 VDD.t120 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X171 VDD RST.t5 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t51 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X172 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT VSS.t168 VSS.t167 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X173 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t262 VDD.t264 VDD.t263 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X174 VDD CLK.t13 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VDD.t122 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X175 a_8696_n338# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS.t255 VSS.t254 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X176 VSS CLK_div_10_mag_0.and2_mag_0.OUT Vdiv110.t3 VSS.t289 nfet_03v3 ad=86.8f pd=0.92u as=86.8f ps=0.92u w=0.22u l=0.28u
X177 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_10590_2727# VSS.t186 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X178 a_7408_n338# VDD.t493 VSS.t94 VSS.t93 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X179 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t400 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X180 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t292 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X181 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.QB a_9260_n338# VSS.t125 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X182 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB VDD.t368 VDD.t367 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X183 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t314 VDD.t313 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X184 a_8132_n338# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VSS.t154 VSS.t153 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X185 a_1368_759# VDD.t494 VSS.t96 VSS.t95 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X186 VDD CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.JK_FF_mag_2.K.t1 VDD.t157 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X187 a_7995_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT VSS.t258 VSS.t257 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X188 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t129 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X189 a_1900_1634# RST.t6 a_1740_1634# VSS.t34 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X190 a_10590_2727# CLK.t14 a_10430_2727# VSS.t72 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X191 VDD RST.t7 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD.t54 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X192 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t97 VDD.t96 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X193 a_2252_759# RST.t8 a_2092_759# VSS.t35 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X194 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q0 VDD.t149 VDD.t148 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X195 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t312 VDD.t311 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X196 a_9260_n338# CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS.t227 VSS.t226 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X197 VDD CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t1 VDD.t360 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X198 a_4317_2729# CLK.t15 a_4157_2729# VSS.t73 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X199 Vdiv110 CLK_div_10_mag_0.Q3 VSS.t105 VSS.t104 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X200 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.and2_mag_3.IN1 a_6609_4975# VSS.t206 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X201 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_11867_759# VSS.t195 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X202 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_11872_1674# VSS.t53 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X203 VDD RST.t9 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT VDD.t57 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X204 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_5679_n338# VSS.t274 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X205 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t419 VDD.t418 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X206 a_8314_n1435# CLK_div_10_mag_0.Q1 VSS.t114 VSS.t37 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X207 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD.t259 VDD.t261 VDD.t260 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X208 a_4551_n338# CLK_div_10_mag_0.Q0 a_4391_n338# VSS.t11 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X209 CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t219 VDD.t218 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X210 VDD CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.Q2 VDD.t205 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X211 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD.t272 VDD.t271 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X212 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 a_1900_1634# VSS.t54 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X213 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD.t447 VDD.t446 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X214 VDD CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.QB VDD.t15 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X215 a_4157_2729# CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t2 VSS.t229 VSS.t228 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X216 a_12478_n2129# CLK_div_10_mag_0.and2_mag_0.OUT a_12318_n2129# VDD.t460 pfet_03v3 ad=0.624p pd=2.92u as=0.624p ps=2.92u w=2.4u l=0.28u
X217 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK.t16 VSS.t128 VSS.t127 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X218 a_11872_1674# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VSS.t173 VSS.t172 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X219 a_5679_n338# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS.t58 VSS.t57 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X220 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_10_mag_0.Q2 a_7562_759# VSS.t39 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X221 a_5109_759# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VSS.t270 VSS.t269 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X222 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VDD.t449 VDD.t448 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X223 a_8149_1634# RST.t10 a_7989_1634# VSS.t36 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X224 a_n350_4053# CLK_DIV_11_mag_new_0.Q0 VSS.t86 VSS.t85 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X225 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t370 VDD.t369 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X226 a_4391_n338# CLK_div_10_mag_0.JK_FF_mag_2.K.t5 VSS.t119 VSS.t118 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X227 a_5599_1676# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t140 VSS.t139 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X228 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.QB a_6243_n338# VSS.t174 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X229 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD.t373 VDD.t372 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X230 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t5 a_1114_4881# VDD.t190 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X231 a_5115_n338# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VSS.t192 VSS.t191 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X232 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.K.t6 a_10585_n338# VSS.t9 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X233 a_9414_759# CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS.t194 VSS.t193 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X234 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.Q2 a_6163_1676# VSS.t262 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X235 a_9346_4996# CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 VDD.t457 VDD.t456 pfet_03v3 ad=0.624p pd=2.92u as=1.06p ps=5.68u w=2.4u l=0.28u
X236 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD.t440 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X237 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q1 VDD.t175 VDD.t174 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X238 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK.t17 VDD.t211 VDD.t210 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X239 a_10579_759# CLK_div_10_mag_0.Q0 a_10419_759# VSS.t10 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X240 VDD CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD.t12 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X241 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD.t225 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X242 VDD CLK.t18 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT VDD.t212 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X243 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD.t106 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X244 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD.t229 VDD.t228 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X245 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q1 VDD.t359 VDD.t358 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X246 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_11713_n338# VSS.t19 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X247 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_4881_2773# VSS.t138 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X248 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q3 a_n1755_2260# VSS.t252 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X249 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t85 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X250 a_10585_n338# CLK_div_10_mag_0.Q0 a_10425_n338# VSS.t9 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X251 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_2662_n338# VSS.t310 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X252 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_10_mag_0.Q1 VDD.t173 VDD.t172 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X253 a_6163_1676# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t164 VSS.t163 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X254 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t101 VDD.t100 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X255 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t396 VDD.t395 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X256 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q1 VDD.t357 VDD.t356 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X257 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.K.t7 VDD.t189 VDD.t188 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X258 a_1534_n338# CLK_div_10_mag_0.CLK a_1374_n338# VSS.t44 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X259 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t305 VDD.t304 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X260 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t139 VDD.t138 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X261 VDD CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.Q1 VDD.t297 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X262 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.CLK VSS.t43 VSS.t42 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X263 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_2464_1678# VSS.t244 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X264 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.K VDD.t471 VDD.t470 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X265 a_1528_759# CLK_div_10_mag_0.CLK a_1368_759# VSS.t41 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X266 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT VDD.t451 VDD.t450 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X267 a_7431_2731# CLK.t19 a_7271_2731# VSS.t129 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X268 VDD CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t6 CLK_DIV_11_mag_new_0.Q1 VDD.t191 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X269 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD.t325 VDD.t324 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X270 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.K.t8 VDD.t221 VDD.t220 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X271 a_4881_2773# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t185 VSS.t184 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X272 VDD CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB VDD.t145 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X273 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q0 VSS.t84 VSS.t83 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X274 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_2098_n338# VSS.t16 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X275 a_2662_n338# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t25 VSS.t24 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X276 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t417 VDD.t416 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X277 VDD RST.t11 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VDD.t244 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X278 a_5833_759# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VSS.t156 VSS.t155 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X279 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_5445_2773# VSS.t77 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X280 a_1374_n338# VDD.t495 VSS.t98 VSS.t97 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X281 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.K VDD.t3 VDD.t2 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X282 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t331 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X283 a_2464_1678# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t183 VSS.t182 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X284 VDD CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD.t169 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X285 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q1 a_9277_1678# VSS.t214 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X286 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VDD.t291 VDD.t290 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X287 a_7271_2731# CLK_DIV_11_mag_new_0.JK_FF_mag_2.K VSS.t297 VSS.t296 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X288 VDD CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t9 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X289 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t484 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X290 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t31 VDD.t30 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X291 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t3 VDD.t375 VDD.t374 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X292 a_n796_2646# CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 VDD.t433 VDD.t432 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X293 VSS CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t7 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VSS.t120 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X294 VDD CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t78 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X295 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.Q0 VSS.t8 VSS.t7 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X296 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK.t20 VSS.t131 VSS.t130 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X297 VDD CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT VDD.t142 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X298 a_11308_1630# RST.t12 a_11148_1630# VSS.t151 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X299 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_DIV_11_mag_new_0.Q3 VSS.t251 VSS.t250 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X300 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VDD.t242 VDD.t241 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X301 a_n1595_3762# CLK_DIV_11_mag_new_0.Q0 a_n1755_3762# VSS.t82 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X302 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t27 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X303 a_10424_1630# CLK_DIV_11_mag_new_0.JK_FF_mag_3.K VSS.t3 VSS.t2 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X304 a_9277_1678# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS.t277 VSS.t276 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X305 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t37 VDD.t36 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X306 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t113 VDD.t112 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X307 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t377 VDD.t376 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X308 VSS CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VSS.t83 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X309 VDD RST.t13 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t247 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X310 a_4151_1632# CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t4 VSS.t144 VSS.t143 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X311 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t256 VDD.t258 VDD.t257 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X312 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q3 VDD.t412 VDD.t411 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X313 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t236 VDD.t235 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X314 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.K VDD.t1 VDD.t0 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X315 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.Q1 a_6397_759# VSS.t113 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X316 a_4385_759# VDD.t496 VSS.t100 VSS.t99 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X317 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.Q0 VDD.t315 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X318 a_n358_4884# CLK_DIV_11_mag_new_0.Q0 VDD.t141 VDD.t140 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X319 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_10_mag_0.Q3 a_10579_759# VSS.t103 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X320 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VDD.t35 VDD.t34 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X321 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t287 VDD.t286 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X322 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.CLK VDD.t77 VDD.t76 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X323 a_12318_n2129# CLK_div_10_mag_0.nor_3_mag_0.IN3 VDD.t339 VDD.t338 pfet_03v3 ad=0.624p pd=2.92u as=1.06p ps=5.68u w=2.4u l=0.28u
X324 VDD CLK.t21 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t215 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X325 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t253 VDD.t255 VDD.t254 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X326 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_8559_2775# VSS.t134 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X327 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VSS.t235 VSS.t234 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X328 VDD CLK.t22 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t114 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X329 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q2 a_10250_n1435# VSS.t4 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X330 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q3 a_1176_1634# VSS.t249 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X331 a_12431_759# CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t308 VSS.t307 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X332 VDD CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VDD.t408 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X333 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t477 VDD.t476 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X334 a_8126_759# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VSS.t90 VSS.t89 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X335 a_1740_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t142 VSS.t141 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X336 a_10430_2727# CLK_DIV_11_mag_new_0.JK_FF_mag_3.K VSS.t1 VSS.t0 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X337 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD.t335 VDD.t334 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X338 VSS CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT VSS.t259 nfet_03v3 ad=86.8f pd=0.92u as=86.8f ps=0.92u w=0.22u l=0.28u
X339 VDD RST.t14 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t250 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X340 VDD CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t353 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X341 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_7995_2775# VSS.t49 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X342 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t5 VDD.t238 VDD.t237 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X343 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t328 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X344 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q1 VDD.t352 VDD.t351 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X345 a_6609_4975# CLK_DIV_11_mag_new_0.Q1 VSS.t213 VSS.t212 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X346 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.Q1 VSS.t112 VSS.t111 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X347 a_8559_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS.t179 VSS.t178 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X348 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.Q2 VDD.t364 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X349 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t308 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X350 a_1176_1634# CLK.t23 a_1016_1634# VSS.t66 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X351 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.Q0 VDD.t8 VDD.t7 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X352 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t8 a_9123_2775# VSS.t68 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X353 a_9282_n1435# CLK_div_10_mag_0.Q2 VSS.t38 VSS.t37 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X354 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_2816_759# VSS.t309 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X355 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.Q0 a_12436_1674# VSS.t81 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X356 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t439 VDD.t438 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X357 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT VDD.t289 VDD.t288 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X358 VDD CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.Q3 VDD.t384 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X359 a_n1762_4447# CLK_DIV_11_mag_new_0.Q1 VSS.t211 VSS.t210 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X360 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VDD.t383 VDD.t382 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X361 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VDD.t459 VDD.t458 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X362 VDD CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t64 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X363 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_10_mag_0.Q2 VDD.t63 VDD.t62 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X364 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD.t435 VDD.t434 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X365 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q1 a_n350_4053# VSS.t85 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X366 a_6243_n338# CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS.t189 VSS.t188 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X367 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VSS.t279 VSS.t278 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X368 a_1114_4881# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VDD.t381 VDD.t380 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X369 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t397 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X370 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD.t327 VDD.t326 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X371 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_11303_759# VSS.t293 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X372 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t394 VDD.t393 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X373 VDD CLK.t24 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t117 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X374 VDD CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t4 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X375 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_1182_2731# VSS.t233 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X376 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT VDD.t279 VDD.t278 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X377 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q2 VDD.t61 VDD.t60 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X378 a_8850_759# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VSS.t32 VSS.t31 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X379 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 VSS.t268 VSS.t267 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X380 CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t481 VDD.t480 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X381 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_11149_n338# VSS.t19 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X382 VDD CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t405 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X383 a_11713_n338# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t292 VSS.t19 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X384 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VSS.t288 VSS.t287 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X385 a_3028_1678# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t65 VSS.t64 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X386 a_4545_759# CLK_div_10_mag_0.Q0 a_4385_759# VSS.t6 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X387 a_10425_n338# CLK_div_10_mag_0.JK_FF_mag_0.K VSS.t271 VSS.t9 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X388 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_11718_2771# VSS.t52 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X389 a_1182_2731# CLK.t25 a_1022_2731# VSS.t67 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X390 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.Q1 VDD.t168 VDD.t167 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X391 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_2252_759# VSS.t23 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X392 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD.t321 VDD.t320 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X393 VDD CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t73 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X394 a_6009_2773# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t166 VSS.t165 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X395 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.QB a_3226_n338# VSS.t294 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X396 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD.t82 VDD.t81 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X397 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_11154_2771# VSS.t171 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X398 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD.t222 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X399 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD.t166 VDD.t165 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X400 a_2098_n338# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t108 VSS.t107 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X401 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT VSS.t159 VSS.t158 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X402 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT VSS.t281 VSS.t280 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X403 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT VDD.t105 VDD.t104 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X404 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q1 VDD.t350 VDD.t349 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X405 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD.t274 VDD.t273 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X406 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.Q3 a_3028_1678# VSS.t248 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X407 a_5445_2773# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t303 VSS.t302 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X408 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t135 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X409 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t462 VDD.t461 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X410 a_7402_759# VDD.t497 VSS.t102 VSS.t101 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X411 VSS CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t223 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X412 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.K VDD.t437 VDD.t436 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X413 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 a_n796_2646# VDD.t371 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X414 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_6009_2773# VSS.t219 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X415 a_5269_759# RST.t15 a_5109_759# VSS.t152 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X416 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VSS.t170 VSS.t169 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X417 a_10250_n1435# CLK_div_10_mag_0.Q0 VSS.t5 VSS.t4 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X418 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_1746_2775# VSS.t181 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X419 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q2 VDD.t424 VDD.t423 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X420 a_11148_1630# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT VSS.t61 VSS.t60 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X421 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.Q1 a_7425_1634# VSS.t209 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
R0 VSS.n12 VSS.n11 19658.7
R1 VSS.n228 VSS.n115 18801.2
R2 VSS.n309 VSS.n308 18801.2
R3 VSS.t127 VSS.n70 17230
R4 VSS.n14 VSS.n12 16362.9
R5 VSS.n392 VSS.n391 14314
R6 VSS.n68 VSS.n14 12989.3
R7 VSS.n371 VSS.t259 10467.5
R8 VSS.n211 VSS.n210 9589.42
R9 VSS.n132 VSS.n131 9415.54
R10 VSS.n67 VSS.n15 8023.75
R11 VSS.n135 VSS.n133 7478.84
R12 VSS.n8 VSS.n7 7059.24
R13 VSS.n130 VSS.t250 7006.49
R14 VSS.n164 VSS.n163 6991.69
R15 VSS.n14 VSS.n13 6944.83
R16 VSS.n416 VSS.n415 6785.63
R17 VSS.n52 VSS.n29 6418.54
R18 VSS.n181 VSS.n180 5437.96
R19 VSS.n135 VSS.n134 4690.81
R20 VSS.n52 VSS.n28 4416.33
R21 VSS.n227 VSS.n120 3893.61
R22 VSS.n282 VSS.n281 3472.05
R23 VSS.n152 VSS.n151 3262.63
R24 VSS.n191 VSS.t200 3112.87
R25 VSS.n159 VSS.n152 3004.05
R26 VSS.n371 VSS.n370 2588.5
R27 VSS.n285 VSS.n284 2416.67
R28 VSS.t77 VSS.t165 2307.56
R29 VSS.t302 VSS.t138 2307.56
R30 VSS.t220 VSS.t184 2307.56
R31 VSS.t134 VSS.t45 2307.56
R32 VSS.t178 VSS.t49 2307.56
R33 VSS.t76 VSS.t257 2307.56
R34 VSS.t52 VSS.t196 2307.56
R35 VSS.t21 VSS.t186 2307.56
R36 VSS.t245 VSS.t240 2307.56
R37 VSS.t55 VSS.t181 2307.56
R38 VSS.t233 VSS.t300 2307.56
R39 VSS.t198 VSS.t310 2307.56
R40 VSS.t24 VSS.t16 2307.56
R41 VSS.t107 VSS.t295 2307.56
R42 VSS.t254 VSS.t33 2307.56
R43 VSS.t126 VSS.t153 2307.56
R44 VSS.t93 VSS.t111 2307.56
R45 VSS.t274 VSS.t188 2307.56
R46 VSS.t175 VSS.t191 2307.56
R47 VSS.n311 VSS.n285 2213.34
R48 VSS.n370 VSS.t285 2166.67
R49 VSS.t66 VSS.n8 1984.24
R50 VSS.n67 VSS.t287 1957.66
R51 VSS.t283 VSS.n126 1878.69
R52 VSS.t118 VSS.n314 1862.04
R53 VSS.n132 VSS.t68 1731.96
R54 VSS.t236 VSS.n392 1719.63
R55 VSS.n309 VSS.t294 1713.53
R56 VSS.t125 VSS.n211 1713.53
R57 VSS.t174 VSS.n228 1713.53
R58 VSS.n376 VSS.t169 1635.55
R59 VSS.n228 VSS.n227 1565.03
R60 VSS.n52 VSS.t234 1564.96
R61 VSS.n302 VSS.t42 1439.29
R62 VSS.t210 VSS.n40 1390.8
R63 VSS.n149 VSS.t27 1272.1
R64 VSS.n151 VSS.n132 1249.34
R65 VSS.n261 VSS.t296 1199.47
R66 VSS.n150 VSS.t0 1199.47
R67 VSS.t160 VSS.n416 1199.47
R68 VSS.t97 VSS.n303 1199.47
R69 VSS.t219 VSS.n262 1153.78
R70 VSS.t187 VSS.n135 1153.78
R71 VSS.t289 VSS.n181 1150.77
R72 VSS.n390 VSS.t176 1143.48
R73 VSS.n373 VSS.n372 1139.06
R74 VSS.n34 VSS.t158 1134.57
R75 VSS.n278 VSS.n10 1119.51
R76 VSS.n391 VSS.t263 1104.59
R77 VSS.n134 VSS.t81 1093.68
R78 VSS.n163 VSS.n162 1062.21
R79 VSS.t26 VSS.t212 1058.09
R80 VSS.n52 VSS.n51 988.177
R81 VSS.t307 VSS.t53 952.793
R82 VSS.t87 VSS.t145 952.793
R83 VSS.n391 VSS.n68 949.904
R84 VSS.n74 VSS.t280 927.716
R85 VSS.t73 VSS.t220 913.885
R86 VSS.t129 VSS.t76 913.885
R87 VSS.t186 VSS.t72 913.885
R88 VSS.t67 VSS.t233 913.885
R89 VSS.t295 VSS.t44 913.885
R90 VSS.t117 VSS.t126 913.885
R91 VSS.t11 VSS.t175 913.885
R92 VSS.n310 VSS.n309 902.461
R93 VSS.n311 VSS.n310 839.713
R94 VSS.n128 VSS.t132 838.187
R95 VSS.n314 VSS.n311 756.466
R96 VSS.n260 VSS.t127 730.073
R97 VSS.n120 VSS.t298 680.952
R98 VSS.n190 VSS.t289 671.942
R99 VSS.n50 VSS.t266 663.793
R100 VSS.n281 VSS.n280 650.433
R101 VSS.t62 VSS.t276 635.715
R102 VSS.t39 VSS.t47 635.715
R103 VSS.n403 VSS.t69 598.279
R104 VSS.n51 VSS.t305 596.024
R105 VSS.n372 VSS.t206 578.554
R106 VSS.n119 VSS.t113 564.287
R107 VSS.n265 VSS.t219 548.331
R108 VSS.n266 VSS.t77 548.331
R109 VSS.n272 VSS.t138 548.331
R110 VSS.n273 VSS.t73 548.331
R111 VSS.n248 VSS.t134 548.331
R112 VSS.n254 VSS.t49 548.331
R113 VSS.n255 VSS.t129 548.331
R114 VSS.n138 VSS.t187 548.331
R115 VSS.n139 VSS.t52 548.331
R116 VSS.n142 VSS.t171 548.331
R117 VSS.n147 VSS.t72 548.331
R118 VSS.n395 VSS.t236 548.331
R119 VSS.n396 VSS.t245 548.331
R120 VSS.n401 VSS.t181 548.331
R121 VSS.n417 VSS.t67 548.331
R122 VSS.t294 VSS.n307 548.331
R123 VSS.t310 VSS.n306 548.331
R124 VSS.t16 VSS.n305 548.331
R125 VSS.t44 VSS.n304 548.331
R126 VSS.n212 VSS.t125 548.331
R127 VSS.n215 VSS.t63 548.331
R128 VSS.n220 VSS.t33 548.331
R129 VSS.n221 VSS.t117 548.331
R130 VSS.n231 VSS.t174 548.331
R131 VSS.n232 VSS.t274 548.331
R132 VSS.n237 VSS.t157 548.331
R133 VSS.n315 VSS.t11 548.331
R134 VSS.n280 VSS.n279 545.501
R135 VSS.t200 VSS.n190 479.959
R136 VSS.t91 VSS.n164 470.426
R137 VSS.t29 VSS.t248 457.144
R138 VSS.n211 VSS.n125 451.231
R139 VSS.n314 VSS.t13 445.519
R140 VSS.n120 VSS.n119 440.476
R141 VSS.n151 VSS.n150 426.769
R142 VSS.n18 VSS.t83 426.396
R143 VSS.t275 VSS.t163 405.356
R144 VSS.t139 VSS.t59 405.356
R145 VSS.t116 VSS.t204 405.356
R146 VSS.t4 VSS.t202 398.623
R147 VSS.t207 VSS.n382 396.058
R148 VSS.n162 VSS.n129 383.952
R149 VSS.t6 VSS.t116 381.512
R150 VSS.t41 VSS.t15 380.952
R151 VSS.t249 VSS.t66 380.952
R152 VSS.n159 VSS.t40 373.81
R153 VSS.t151 VSS.t293 370.132
R154 VSS.t124 VSS.t103 370.132
R155 VSS.t165 VSS.n265 365.555
R156 VSS.n266 VSS.t302 365.555
R157 VSS.t184 VSS.n272 365.555
R158 VSS.n273 VSS.t228 365.555
R159 VSS.t45 VSS.n247 365.555
R160 VSS.n248 VSS.t178 365.555
R161 VSS.t257 VSS.n254 365.555
R162 VSS.n255 VSS.t296 365.555
R163 VSS.t196 VSS.n138 365.555
R164 VSS.n139 VSS.t231 365.555
R165 VSS.n142 VSS.t21 365.555
R166 VSS.t0 VSS.n147 365.555
R167 VSS.t240 VSS.n395 365.555
R168 VSS.n396 VSS.t55 365.555
R169 VSS.t300 VSS.n401 365.555
R170 VSS.n417 VSS.t160 365.555
R171 VSS.n307 VSS.t198 365.555
R172 VSS.n306 VSS.t24 365.555
R173 VSS.n305 VSS.t107 365.555
R174 VSS.n304 VSS.t97 365.555
R175 VSS.n212 VSS.t226 365.555
R176 VSS.n215 VSS.t254 365.555
R177 VSS.t153 VSS.n220 365.555
R178 VSS.n221 VSS.t93 365.555
R179 VSS.t188 VSS.n231 365.555
R180 VSS.n232 VSS.t57 365.555
R181 VSS.t191 VSS.n237 365.555
R182 VSS.n315 VSS.t118 365.555
R183 VSS.n372 VSS.n371 345.394
R184 VSS.n392 VSS.n10 329.483
R185 VSS.t85 VSS.t311 329.029
R186 VSS.t180 VSS.t256 326.19
R187 VSS.t209 VSS.t39 326.19
R188 VSS.n131 VSS.n130 297.363
R189 VSS.n284 VSS.n283 287.072
R190 VSS.n71 VSS.t278 281.091
R191 VSS.n17 VSS.t120 269.688
R192 VSS.t272 VSS.t267 259.553
R193 VSS.n37 VSS.t253 255.748
R194 VSS.n127 VSS.t4 231.852
R195 VSS.n103 VSS.t262 228.907
R196 VSS.n106 VSS.t275 228.907
R197 VSS.n105 VSS.t78 228.907
R198 VSS.n110 VSS.t237 228.907
R199 VSS.n238 VSS.t71 228.907
R200 VSS.t113 VSS.n118 228.796
R201 VSS.t40 VSS.n158 228.571
R202 VSS.n153 VSS.t62 228.571
R203 VSS.n96 VSS.t238 228.571
R204 VSS.n121 VSS.t115 228.571
R205 VSS.t248 VSS.n3 228.571
R206 VSS.n239 VSS.t309 228.571
R207 VSS.n4 VSS.t244 228.571
R208 VSS.n294 VSS.t35 228.571
R209 VSS.n6 VSS.t34 228.571
R210 VSS.n297 VSS.t41 228.571
R211 VSS.t106 VSS.n77 217.304
R212 VSS.t195 VSS.n79 217.304
R213 VSS.n84 VSS.t239 217.304
R214 VSS.n89 VSS.t10 217.304
R215 VSS.t37 VSS.t221 211.208
R216 VSS.n180 VSS.n129 206.661
R217 VSS.n284 VSS.t143 202.679
R218 VSS.n210 VSS.n126 195.244
R219 VSS.t234 VSS.n17 192.633
R220 VSS.n19 VSS.t85 191.375
R221 VSS.n383 VSS.t88 186.381
R222 VSS.n381 VSS.t26 176.673
R223 VSS.t304 VSS.t152 176.45
R224 VSS.t265 VSS.t6 176.45
R225 VSS.t193 VSS.n92 173.81
R226 VSS.t12 VSS.n282 166.667
R227 VSS.n160 VSS.n159 164.286
R228 VSS.n41 VSS.t215 163.793
R229 VSS.n118 VSS.t136 152.606
R230 VSS.t163 VSS.n103 152.606
R231 VSS.n106 VSS.t155 152.606
R232 VSS.n105 VSS.t139 152.606
R233 VSS.n111 VSS.t269 152.606
R234 VSS.t204 VSS.n110 152.606
R235 VSS.n114 VSS.t99 152.606
R236 VSS.t143 VSS.n238 152.606
R237 VSS.t276 VSS.n92 152.381
R238 VSS.n93 VSS.t50 152.381
R239 VSS.t47 VSS.n95 152.381
R240 VSS.t298 VSS.n100 152.381
R241 VSS.n244 VSS.t29 152.381
R242 VSS.t64 VSS.n3 152.381
R243 VSS.n239 VSS.t17 152.381
R244 VSS.n4 VSS.t182 152.381
R245 VSS.n294 VSS.t242 152.381
R246 VSS.t141 VSS.n6 152.381
R247 VSS.n297 VSS.t95 152.381
R248 VSS.n191 VSS.t246 150.845
R249 VSS.n194 VSS.t283 150.845
R250 VSS.n180 VSS.n125 142.794
R251 VSS.n184 VSS.t109 140.889
R252 VSS.n80 VSS.t172 140.889
R253 VSS.t60 VSS.n88 140.889
R254 VSS.n165 VSS.t2 140.889
R255 VSS.t88 VSS.n381 133.962
R256 VSS.n415 VSS.t147 132.734
R257 VSS.t212 VSS.n380 124.254
R258 VSS.n383 VSS.t207 124.254
R259 VSS.t309 VSS.t64 123.811
R260 VSS.t182 VSS.t23 123.811
R261 VSS.t15 VSS.t141 123.811
R262 VSS.n209 VSS.t37 122.846
R263 VSS.n227 VSS.n226 119.948
R264 VSS.t19 VSS.t7 113.144
R265 VSS.t206 VSS.n70 99.0148
R266 VSS.n158 VSS.t214 97.6195
R267 VSS.n153 VSS.t135 97.6195
R268 VSS.n96 VSS.t36 97.6195
R269 VSS.n121 VSS.t123 97.6195
R270 VSS.t83 VSS.t74 94.0088
R271 VSS.n380 VSS.n70 87.3661
R272 VSS.n53 VSS.n52 77.2216
R273 VSS.t242 VSS.t54 76.191
R274 VSS.t95 VSS.t249 76.191
R275 VSS.n405 VSS.t223 64.396
R276 VSS.n42 VSS.t252 63.0818
R277 VSS.n282 VSS.n244 61.9053
R278 VSS.n161 VSS.n160 57.1434
R279 VSS.t214 VSS.t193 54.7624
R280 VSS.t135 VSS.t31 54.7624
R281 VSS.t238 VSS.t180 54.7624
R282 VSS.t36 VSS.t89 54.7624
R283 VSS.t115 VSS.t209 54.7624
R284 VSS.t123 VSS.t101 54.7624
R285 VSS.n251 VSS.n102 54.1355
R286 VSS.n111 VSS.t304 52.4583
R287 VSS.n114 VSS.t265 52.4583
R288 VSS.n386 VSS.t176 47.8266
R289 VSS.t263 VSS.n390 47.8266
R290 VSS.t267 VSS.n405 45.9973
R291 VSS.n42 VSS.t217 42.0547
R292 VSS.n150 VSS.n149 41.0359
R293 VSS.n179 VSS.t9 40.409
R294 VSS.n303 VSS.n302 37.1434
R295 VSS.n226 VSS.t111 34.2711
R296 VSS.t13 VSS.n313 34.2711
R297 VSS.n423 VSS.n8 30.9563
R298 VSS.n269 VSS.n2 27.068
R299 VSS.n283 VSS.t12 25.9531
R300 VSS.t9 VSS.t19 25.4001
R301 VSS.n261 VSS.n260 23.5512
R302 VSS.n279 VSS.t130 22.8476
R303 VSS.n210 VSS.n128 21.6311
R304 VSS.n68 VSS.n67 21.1044
R305 VSS.t253 VSS.t82 20.1154
R306 VSS.t215 VSS.t210 20.1154
R307 VSS.n416 VSS.n403 19.2998
R308 VSS.t305 VSS.n50 17.2419
R309 VSS.t287 VSS.n66 16.5119
R310 VSS.n164 VSS.n161 16.3322
R311 VSS.n210 VSS.n127 16.2708
R312 VSS.n421 VSS.n9 13.2511
R313 VSS.t81 VSS.t106 11.9402
R314 VSS.t109 VSS.t307 11.9402
R315 VSS.t53 VSS.t195 11.9402
R316 VSS.t172 VSS.t79 11.9402
R317 VSS.t293 VSS.t230 11.9402
R318 VSS.t239 VSS.t151 11.9402
R319 VSS.t145 VSS.t60 11.9402
R320 VSS.t103 VSS.t87 11.9402
R321 VSS.t10 VSS.t124 11.9402
R322 VSS.t2 VSS.t91 11.9402
R323 VSS.n279 VSS.n278 11.424
R324 VSS.n407 VSS.t273 10.2623
R325 VSS.n262 VSS.n261 9.42079
R326 VSS.n389 VSS.t264 9.40866
R327 VSS.n188 VSS.t201 9.37686
R328 VSS.n225 VSS.t112 9.3736
R329 VSS.n312 VSS.t14 9.3736
R330 VSS.n301 VSS.t43 9.3736
R331 VSS.n277 VSS.t131 9.3736
R332 VSS.n178 VSS.t8 9.3736
R333 VSS.n148 VSS.t28 9.3736
R334 VSS.n259 VSS.t128 9.3736
R335 VSS.n402 VSS.t70 9.3736
R336 VSS.n59 VSS.t75 9.3645
R337 VSS.n63 VSS.n16 9.3221
R338 VSS.n61 VSS.t235 9.3221
R339 VSS.n57 VSS.n22 9.3221
R340 VSS.n31 VSS.t84 9.3221
R341 VSS.n378 VSS.t170 9.30652
R342 VSS.n360 VSS.t168 9.30652
R343 VSS.n76 VSS.t281 9.30652
R344 VSS.n64 VSS.t288 9.30652
R345 VSS.n21 VSS.t312 9.30652
R346 VSS.n48 VSS.t306 9.30652
R347 VSS.n36 VSS.t159 9.30652
R348 VSS.n207 VSS.t222 9.30652
R349 VSS.n202 VSS.t133 9.30652
R350 VSS.n198 VSS.t203 9.30652
R351 VSS.n375 VSS.t279 9.30518
R352 VSS.n362 VSS.t282 9.30518
R353 VSS.n193 VSS.t247 9.30518
R354 VSS.n368 VSS.t286 9.30323
R355 VSS.n412 VSS.t148 9.30204
R356 VSS.n388 VSS.t177 9.29981
R357 VSS.n410 VSS.n404 9.29009
R358 VSS.n408 VSS.t268 9.29009
R359 VSS.n196 VSS.t284 9.25414
R360 VSS.n210 VSS.n209 8.62119
R361 VSS.n32 VSS.n27 7.39136
R362 VSS VSS.t114 7.30633
R363 VSS.n240 VSS.t18 7.19156
R364 VSS.n242 VSS.t30 7.19156
R365 VSS.n108 VSS.t156 7.19156
R366 VSS.n116 VSS.t137 7.19156
R367 VSS.n154 VSS.t32 7.19156
R368 VSS.n156 VSS.t194 7.19156
R369 VSS.n82 VSS.t80 7.19156
R370 VSS.n185 VSS.t308 7.19156
R371 VSS.n218 VSS.t154 7.19156
R372 VSS.n217 VSS.t255 7.19156
R373 VSS.n214 VSS.t227 7.19156
R374 VSS.n235 VSS.t192 7.19156
R375 VSS.n234 VSS.t58 7.19156
R376 VSS.n229 VSS.t189 7.19156
R377 VSS.n291 VSS.t108 7.19156
R378 VSS.n289 VSS.t25 7.19156
R379 VSS.n287 VSS.t199 7.19156
R380 VSS.n174 VSS.t190 7.19156
R381 VSS.n172 VSS.t292 7.19156
R382 VSS.n170 VSS.t20 7.19156
R383 VSS.n30 VSS.t86 7.19156
R384 VSS.n342 VSS.t277 7.17323
R385 VSS.n340 VSS.t51 7.17323
R386 VSS.n429 VSS.t65 7.17323
R387 VSS.n426 VSS.t183 7.17323
R388 VSS.n69 VSS.t213 7.17156
R389 VSS.n329 VSS.t164 7.16989
R390 VSS.n327 VSS.t140 7.16989
R391 VSS.n355 VSS.t110 7.16656
R392 VSS.n352 VSS.t173 7.16656
R393 VSS.n45 VSS.t211 7.16085
R394 VSS.n44 VSS.t218 7.15156
R395 VSS.n245 VSS.t46 7.13489
R396 VSS.n250 VSS.t179 7.13489
R397 VSS.n252 VSS.t258 7.13489
R398 VSS.n393 VSS.t241 7.13323
R399 VSS.n398 VSS.t56 7.13323
R400 VSS.n399 VSS.t301 7.13323
R401 VSS.n263 VSS.t166 7.13156
R402 VSS.n268 VSS.t303 7.13156
R403 VSS.n270 VSS.t185 7.13156
R404 VSS.n367 VSS.n366 7.1285
R405 VSS.n136 VSS.t197 7.12823
R406 VSS.n141 VSS.t232 7.12823
R407 VSS.n144 VSS.t22 7.12823
R408 VSS.n200 VSS.t5 6.88656
R409 VSS.n203 VSS.t38 6.88656
R410 VSS.n45 VSS.n44 6.41993
R411 VSS VSS.t216 6.02876
R412 VSS.n73 VSS.n72 6.01414
R413 VSS.n73 VSS.t251 6.01414
R414 VSS.n183 VSS.n182 6.01414
R415 VSS.n183 VSS.t105 6.01414
R416 VSS.n299 VSS.t96 5.91399
R417 VSS.n296 VSS.t243 5.91399
R418 VSS.n320 VSS.t100 5.91399
R419 VSS.n113 VSS.t270 5.91399
R420 VSS.n123 VSS.t102 5.91399
R421 VSS.n98 VSS.t90 5.91399
R422 VSS.n167 VSS.t92 5.91399
R423 VSS.n86 VSS.t146 5.91399
R424 VSS.n223 VSS.t94 5.91399
R425 VSS.n317 VSS.t119 5.91399
R426 VSS.n293 VSS.t98 5.91399
R427 VSS.n176 VSS.t271 5.91399
R428 VSS.n385 VSS.t208 5.89898
R429 VSS.n337 VSS.t48 5.89565
R430 VSS.n334 VSS.t299 5.89565
R431 VSS.n424 VSS.t142 5.89565
R432 VSS.n422 VSS.t162 5.89565
R433 VSS.n324 VSS.t205 5.89232
R434 VSS.n433 VSS.t144 5.89232
R435 VSS.n349 VSS.t61 5.88898
R436 VSS.n346 VSS.t3 5.88898
R437 VSS.n257 VSS.t297 5.85732
R438 VSS.n419 VSS.t161 5.85565
R439 VSS.n275 VSS.t229 5.85398
R440 VSS.n145 VSS.t1 5.85065
R441 VSS VSS.n406 5.20234
R442 VSS.n278 VSS 5.20137
R443 VSS.n265 VSS.n264 5.2005
R444 VSS.n267 VSS.n266 5.2005
R445 VSS.n272 VSS.n271 5.2005
R446 VSS.n274 VSS.n273 5.2005
R447 VSS.n377 VSS.n376 5.2005
R448 VSS.n374 VSS.n373 5.2005
R449 VSS.n361 VSS.n71 5.2005
R450 VSS.n365 VSS.n364 5.2005
R451 VSS.n370 VSS.n369 5.2005
R452 VSS.n247 VSS.n246 5.2005
R453 VSS.n249 VSS.n248 5.2005
R454 VSS.n254 VSS.n253 5.2005
R455 VSS.n256 VSS.n255 5.2005
R456 VSS.n75 VSS.n74 5.2005
R457 VSS.n138 VSS.n137 5.2005
R458 VSS.n140 VSS.n139 5.2005
R459 VSS.n143 VSS.n142 5.2005
R460 VSS.n147 VSS.n146 5.2005
R461 VSS.n149 VSS.n148 5.2005
R462 VSS.n175 VSS.n129 5.2005
R463 VSS.n173 VSS.n129 5.2005
R464 VSS.n171 VSS.n129 5.2005
R465 VSS.n169 VSS.n129 5.2005
R466 VSS.n179 VSS.n178 5.2005
R467 VSS.n260 VSS.n259 5.2005
R468 VSS.n384 VSS.n383 5.2005
R469 VSS.n380 VSS.n379 5.2005
R470 VSS.n390 VSS.n389 5.2005
R471 VSS.n387 VSS.n386 5.2005
R472 VSS.n395 VSS.n394 5.2005
R473 VSS.n397 VSS.n396 5.2005
R474 VSS.n401 VSS.n400 5.2005
R475 VSS.n418 VSS.n417 5.2005
R476 VSS.n66 VSS.n65 5.2005
R477 VSS.n62 VSS.n17 5.2005
R478 VSS.n25 VSS.n24 5.2005
R479 VSS.n20 VSS.n19 5.2005
R480 VSS.n60 VSS.n18 5.2005
R481 VSS.n35 VSS.n34 5.2005
R482 VSS.n50 VSS.n49 5.2005
R483 VSS.n38 VSS.n37 5.2005
R484 VSS.n46 VSS.n41 5.2005
R485 VSS.n43 VSS.n42 5.2005
R486 VSS.n409 VSS.n405 5.2005
R487 VSS.n414 VSS.n413 5.2005
R488 VSS.n403 VSS.n402 5.2005
R489 VSS.n302 VSS.n301 5.2005
R490 VSS.n425 VSS.n6 5.2005
R491 VSS.n304 VSS.n292 5.2005
R492 VSS.n305 VSS.n290 5.2005
R493 VSS.n306 VSS.n288 5.2005
R494 VSS.n307 VSS.n286 5.2005
R495 VSS.n316 VSS.n315 5.2005
R496 VSS.n237 VSS.n236 5.2005
R497 VSS.n233 VSS.n232 5.2005
R498 VSS.n231 VSS.n230 5.2005
R499 VSS.n313 VSS.n312 5.2005
R500 VSS.n222 VSS.n221 5.2005
R501 VSS.n220 VSS.n219 5.2005
R502 VSS.n216 VSS.n215 5.2005
R503 VSS.n213 VSS.n212 5.2005
R504 VSS.n226 VSS.n225 5.2005
R505 VSS.n206 VSS.n205 5.2005
R506 VSS.n209 VSS.n208 5.2005
R507 VSS.n205 VSS.n204 5.2005
R508 VSS.n197 VSS.n127 5.2005
R509 VSS.n195 VSS.n194 5.2005
R510 VSS.n192 VSS.n191 5.2005
R511 VSS.n190 VSS.n189 5.2005
R512 VSS.n298 VSS.n297 5.2005
R513 VSS.n295 VSS.n294 5.2005
R514 VSS.n241 VSS.n239 5.2005
R515 VSS.n244 VSS.n243 5.2005
R516 VSS.n321 VSS.n114 5.2005
R517 VSS.n112 VSS.n111 5.2005
R518 VSS.n107 VSS.n106 5.2005
R519 VSS.n118 VSS.n117 5.2005
R520 VSS.n122 VSS.n121 5.2005
R521 VSS.n97 VSS.n96 5.2005
R522 VSS.n155 VSS.n153 5.2005
R523 VSS.n158 VSS.n157 5.2005
R524 VSS.n166 VSS.n165 5.2005
R525 VSS.n88 VSS.n87 5.2005
R526 VSS.n81 VSS.n80 5.2005
R527 VSS.n186 VSS.n184 5.2005
R528 VSS.n428 VSS.n4 5.2005
R529 VSS.n430 VSS.n3 5.2005
R530 VSS.n335 VSS.n100 5.2005
R531 VSS.n338 VSS.n95 5.2005
R532 VSS.n341 VSS.n93 5.2005
R533 VSS.n343 VSS.n92 5.2005
R534 VSS.n347 VSS.n89 5.2005
R535 VSS.n350 VSS.n84 5.2005
R536 VSS.n353 VSS.n79 5.2005
R537 VSS.n356 VSS.n77 5.2005
R538 VSS.n331 VSS.n103 5.2005
R539 VSS.n328 VSS.n105 5.2005
R540 VSS.n325 VSS.n110 5.2005
R541 VSS.n238 VSS.n0 5.2005
R542 VSS.n180 VSS.n179 4.61862
R543 VSS.n33 VSS.n32 4.5005
R544 VSS VSS.n33 4.12455
R545 VSS.t147 VSS.n414 3.94308
R546 VSS.n406 VSS.t272 3.94308
R547 VSS.t278 VSS.t167 3.67489
R548 VSS.n373 VSS.n71 3.67489
R549 VSS.n187 VSS.n183 3.36323
R550 VSS.n358 VSS.n73 3.28959
R551 VSS.n366 VSS.n365 3.03722
R552 VSS.n55 VSS.n54 2.6005
R553 VSS.n54 VSS.n53 2.6005
R554 VSS.n187 VSS 2.40845
R555 VSS.n368 VSS.n367 2.13777
R556 VSS.n357 VSS 2.03762
R557 VSS.n61 VSS 1.09141
R558 VSS.n300 VSS.n299 1.03389
R559 VSS.n366 VSS.n71 1.00481
R560 VSS.n181 VSS.t104 0.878786
R561 VSS.n224 VSS.n124 0.846463
R562 VSS.n319 VSS.n318 0.846463
R563 VSS.n177 VSS.n168 0.846463
R564 VSS.n345 VSS.n90 0.843955
R565 VSS.n43 VSS.n9 0.734346
R566 VSS.n332 VSS.n102 0.70444
R567 VSS VSS.n375 0.676801
R568 VSS.n421 VSS.n420 0.623774
R569 VSS.n357 VSS.n76 0.616742
R570 VSS.n431 VSS.n2 0.574895
R571 VSS.n365 VSS.n359 0.486611
R572 VSS.n298 VSS.n296 0.480225
R573 VSS.n384 VSS.n69 0.439554
R574 VSS VSS.n101 0.43894
R575 VSS.n207 VSS.n206 0.395692
R576 VSS.n204 VSS.n202 0.395692
R577 VSS.n199 VSS.n198 0.395692
R578 VSS.n188 VSS 0.378121
R579 VSS.n27 VSS.n26 0.365463
R580 VSS.n168 VSS.n91 0.35472
R581 VSS.n166 VSS.n85 0.348115
R582 VSS VSS.n214 0.343161
R583 VSS VSS.n217 0.343161
R584 VSS.n229 VSS 0.343161
R585 VSS VSS.n234 0.343161
R586 VSS VSS.n287 0.343161
R587 VSS VSS.n289 0.343161
R588 VSS VSS.n170 0.343161
R589 VSS VSS.n172 0.343161
R590 VSS.n156 VSS 0.343161
R591 VSS.n242 VSS 0.343161
R592 VSS.n39 VSS.n36 0.338437
R593 VSS.n87 VSS.n83 0.325821
R594 VSS.n379 VSS.n378 0.316175
R595 VSS.n97 VSS.n94 0.313436
R596 VSS VSS.n385 0.311851
R597 VSS VSS.n193 0.310668
R598 VSS.n295 VSS.n5 0.294445
R599 VSS.n222 VSS 0.289491
R600 VSS.n316 VSS 0.289491
R601 VSS.n292 VSS 0.289491
R602 VSS.n175 VSS 0.289491
R603 VSS.n426 VSS.n425 0.286539
R604 VSS.n408 VSS.n407 0.284276
R605 VSS.n203 VSS 0.27984
R606 VSS VSS.n200 0.27984
R607 VSS.n47 VSS.n46 0.277931
R608 VSS.n39 VSS.n38 0.272151
R609 VSS.n122 VSS.n99 0.268849
R610 VSS.n263 VSS 0.265394
R611 VSS.n245 VSS 0.265394
R612 VSS.n393 VSS 0.259875
R613 VSS VSS.n398 0.259875
R614 VSS.n136 VSS 0.254582
R615 VSS VSS.n141 0.254582
R616 VSS.n322 VSS.n321 0.252335
R617 VSS.n109 VSS.n108 0.250683
R618 VSS VSS.n196 0.250123
R619 VSS.n196 VSS.n195 0.247195
R620 VSS VSS.n203 0.243604
R621 VSS.n200 VSS 0.243604
R622 VSS.n422 VSS.n421 0.241304
R623 VSS VSS.n78 0.240775
R624 VSS VSS.n104 0.23417
R625 VSS.n112 VSS.n109 0.230041
R626 VSS.n322 VSS.n113 0.22839
R627 VSS.n274 VSS 0.223904
R628 VSS.n256 VSS 0.223904
R629 VSS VSS.n388 0.223676
R630 VSS.n418 VSS 0.21925
R631 VSS.n146 VSS 0.214786
R632 VSS.n99 VSS.n98 0.211876
R633 VSS.n319 VSS.n1 0.201142
R634 VSS.n332 VSS 0.192251
R635 VSS.n412 VSS.n411 0.19152
R636 VSS.n218 VSS 0.191234
R637 VSS.n235 VSS 0.191234
R638 VSS VSS.n291 0.191234
R639 VSS VSS.n174 0.191234
R640 VSS.n168 VSS.n167 0.187931
R641 VSS.n124 VSS.n123 0.187931
R642 VSS.n320 VSS.n319 0.187931
R643 VSS.n58 VSS.n21 0.187704
R644 VSS.n240 VSS.n5 0.18628
R645 VSS.n64 VSS.n63 0.184546
R646 VSS.n362 VSS 0.182492
R647 VSS.n358 VSS.n357 0.180913
R648 VSS.n154 VSS.n94 0.167289
R649 VSS.n410 VSS.n409 0.165806
R650 VSS VSS.n91 0.165638
R651 VSS VSS.n45 0.158206
R652 VSS.n424 VSS.n423 0.156125
R653 VSS.n83 VSS.n82 0.154904
R654 VSS.n193 VSS.n192 0.152211
R655 VSS.n270 VSS 0.147947
R656 VSS.n252 VSS 0.147947
R657 VSS.n399 VSS 0.144875
R658 VSS.n323 VSS.n0 0.144447
R659 VSS VSS.n144 0.141929
R660 VSS VSS.n408 0.140092
R661 VSS.n189 VSS.n187 0.138903
R662 VSS.n339 VSS.n338 0.138304
R663 VSS.n326 VSS.n325 0.137236
R664 VSS VSS.n224 0.137136
R665 VSS.n318 VSS 0.137136
R666 VSS VSS.n300 0.137136
R667 VSS VSS.n177 0.137136
R668 VSS.n63 VSS.n62 0.136634
R669 VSS.n269 VSS.n268 0.133266
R670 VSS.n251 VSS.n250 0.133266
R671 VSS VSS.n269 0.132628
R672 VSS VSS.n251 0.132628
R673 VSS.n86 VSS.n85 0.13261
R674 VSS.n420 VSS 0.127807
R675 VSS VSS.n90 0.127258
R676 VSS.n48 VSS.n47 0.12579
R677 VSS.n336 VSS.n335 0.123883
R678 VSS.n214 VSS.n213 0.118573
R679 VSS.n217 VSS.n216 0.118573
R680 VSS.n219 VSS.n218 0.118573
R681 VSS.n230 VSS.n229 0.118573
R682 VSS.n234 VSS.n233 0.118573
R683 VSS.n236 VSS.n235 0.118573
R684 VSS.n287 VSS.n286 0.118573
R685 VSS.n289 VSS.n288 0.118573
R686 VSS.n291 VSS.n290 0.118573
R687 VSS.n170 VSS.n169 0.118573
R688 VSS.n172 VSS.n171 0.118573
R689 VSS.n174 VSS.n173 0.118573
R690 VSS.n186 VSS.n185 0.118573
R691 VSS.n82 VSS.n81 0.118573
R692 VSS.n157 VSS.n156 0.118573
R693 VSS.n155 VSS.n154 0.118573
R694 VSS.n117 VSS.n116 0.118573
R695 VSS.n108 VSS.n107 0.118573
R696 VSS.n243 VSS.n242 0.118573
R697 VSS.n241 VSS.n240 0.118573
R698 VSS.n345 VSS.n344 0.116405
R699 VSS VSS.n61 0.115458
R700 VSS.n223 VSS 0.115271
R701 VSS.n317 VSS 0.115271
R702 VSS.n293 VSS 0.115271
R703 VSS.n176 VSS 0.115271
R704 VSS VSS.n86 0.115271
R705 VSS.n167 VSS 0.115271
R706 VSS.n98 VSS 0.115271
R707 VSS.n123 VSS 0.115271
R708 VSS.n113 VSS 0.115271
R709 VSS VSS.n320 0.115271
R710 VSS.n296 VSS 0.115271
R711 VSS.n299 VSS 0.115271
R712 VSS VSS.n188 0.113945
R713 VSS.n348 VSS.n347 0.111598
R714 VSS.n342 VSS 0.111331
R715 VSS.n329 VSS 0.111331
R716 VSS.n360 VSS 0.109909
R717 VSS.n116 VSS.n104 0.109491
R718 VSS.n388 VSS.n387 0.109351
R719 VSS VSS.n258 0.106075
R720 VSS.n351 VSS.n350 0.104387
R721 VSS.n185 VSS.n78 0.102885
R722 VSS.n224 VSS.n223 0.10206
R723 VSS.n318 VSS.n317 0.10206
R724 VSS.n300 VSS.n293 0.10206
R725 VSS.n177 VSS.n176 0.10206
R726 VSS.n264 VSS.n263 0.0917766
R727 VSS.n268 VSS.n267 0.0917766
R728 VSS.n271 VSS.n270 0.0917766
R729 VSS.n246 VSS.n245 0.0917766
R730 VSS.n250 VSS.n249 0.0917766
R731 VSS.n253 VSS.n252 0.0917766
R732 VSS.n344 VSS 0.0905
R733 VSS.n394 VSS.n393 0.089875
R734 VSS.n398 VSS.n397 0.089875
R735 VSS.n400 VSS.n399 0.089875
R736 VSS.n361 VSS.n360 0.0895055
R737 VSS.n275 VSS 0.0892234
R738 VSS.n257 VSS 0.0892234
R739 VSS.n137 VSS.n136 0.088051
R740 VSS.n141 VSS.n140 0.088051
R741 VSS.n144 VSS.n143 0.088051
R742 VSS.n44 VSS 0.0879825
R743 VSS.n419 VSS 0.087375
R744 VSS.n363 VSS.n362 0.0869264
R745 VSS VSS.n145 0.085602
R746 VSS VSS.n69 0.085027
R747 VSS.n385 VSS 0.085027
R748 VSS.n351 VSS.n83 0.0847202
R749 VSS.n348 VSS.n85 0.0847202
R750 VSS.n344 VSS.n91 0.0847202
R751 VSS.n339 VSS.n94 0.0847202
R752 VSS.n336 VSS.n99 0.0847202
R753 VSS.n333 VSS.n101 0.0847202
R754 VSS.n330 VSS.n104 0.0847202
R755 VSS.n326 VSS.n109 0.0847202
R756 VSS.n323 VSS.n322 0.0847202
R757 VSS.n432 VSS.n1 0.0847202
R758 VSS.n427 VSS.n5 0.0847202
R759 VSS.n354 VSS.n78 0.0847202
R760 VSS.n124 VSS.n101 0.0814174
R761 VSS.n276 VSS.n275 0.0790106
R762 VSS.n258 VSS.n257 0.0790106
R763 VSS.n47 VSS.n39 0.0777727
R764 VSS.n420 VSS.n419 0.077375
R765 VSS.n354 VSS 0.0768798
R766 VSS.n431 VSS 0.0760786
R767 VSS.n369 VSS.n358 0.0760505
R768 VSS.n145 VSS.n90 0.0758061
R769 VSS.n413 VSS.n412 0.073051
R770 VSS.n277 VSS.n276 0.0718942
R771 VSS.n54 VSS.n27 0.071566
R772 VSS.n57 VSS.n56 0.0706762
R773 VSS.n367 VSS 0.0691188
R774 VSS.n378 VSS.n377 0.0675755
R775 VSS.n76 VSS.n75 0.0675755
R776 VSS.n65 VSS.n64 0.0675755
R777 VSS.n21 VSS.n20 0.0675755
R778 VSS.n49 VSS.n48 0.0675755
R779 VSS.n36 VSS.n35 0.0675755
R780 VSS.n208 VSS.n207 0.0675755
R781 VSS.n202 VSS.n201 0.0675755
R782 VSS.n198 VSS.n197 0.0675755
R783 VSS VSS.n424 0.0666607
R784 VSS.n433 VSS.n432 0.0635267
R785 VSS VSS.n368 0.0624266
R786 VSS.n346 VSS.n345 0.0611231
R787 VSS.n30 VSS 0.0548172
R788 VSS.n352 VSS.n351 0.051776
R789 VSS.n334 VSS.n333 0.0507077
R790 VSS.n58 VSS.n57 0.0449053
R791 VSS.n349 VSS.n348 0.0445653
R792 VSS.n375 VSS.n374 0.04
R793 VSS.n356 VSS.n355 0.0386899
R794 VSS.n353 VSS.n352 0.0386899
R795 VSS.n343 VSS.n342 0.0386899
R796 VSS.n341 VSS.n340 0.0386899
R797 VSS.n328 VSS.n327 0.0386899
R798 VSS.n430 VSS.n429 0.0386899
R799 VSS VSS.n422 0.0377321
R800 VSS VSS.n349 0.0376217
R801 VSS VSS.n346 0.0376217
R802 VSS VSS.n337 0.0376217
R803 VSS VSS.n334 0.0376217
R804 VSS VSS.n324 0.0376217
R805 VSS VSS.n433 0.0376217
R806 VSS.n54 VSS.n25 0.036033
R807 VSS.n258 VSS.n102 0.036
R808 VSS.n355 VSS.n354 0.034951
R809 VSS.n427 VSS.n426 0.0344169
R810 VSS.n337 VSS.n336 0.0322804
R811 VSS.n276 VSS.n2 0.0316538
R812 VSS.n330 VSS.n329 0.0277404
R813 VSS.n60 VSS.n59 0.0263107
R814 VSS.n33 VSS.n31 0.0211167
R815 VSS.n411 VSS.n410 0.0197857
R816 VSS.n327 VSS.n326 0.0189273
R817 VSS.n340 VSS.n339 0.017859
R818 VSS VSS.n1 0.0161881
R819 VSS.n429 VSS 0.0154555
R820 VSS.n333 VSS.n332 0.0130519
R821 VSS.n324 VSS.n323 0.0117166
R822 VSS.n331 VSS.n330 0.0114496
R823 VSS.n59 VSS.n58 0.00961702
R824 VSS.n31 VSS.n30 0.00644714
R825 VSS.n213 VSS 0.00545413
R826 VSS.n216 VSS 0.00545413
R827 VSS.n219 VSS 0.00545413
R828 VSS.n230 VSS 0.00545413
R829 VSS.n233 VSS 0.00545413
R830 VSS.n236 VSS 0.00545413
R831 VSS.n286 VSS 0.00545413
R832 VSS.n288 VSS 0.00545413
R833 VSS.n290 VSS 0.00545413
R834 VSS.n169 VSS 0.00545413
R835 VSS.n171 VSS 0.00545413
R836 VSS.n173 VSS 0.00545413
R837 VSS VSS.n186 0.00545413
R838 VSS.n81 VSS 0.00545413
R839 VSS.n157 VSS 0.00545413
R840 VSS VSS.n155 0.00545413
R841 VSS.n117 VSS 0.00545413
R842 VSS.n107 VSS 0.00545413
R843 VSS.n243 VSS 0.00545413
R844 VSS VSS.n241 0.00545413
R845 VSS.n428 VSS.n427 0.004773
R846 VSS.n264 VSS 0.00432979
R847 VSS.n267 VSS 0.00432979
R848 VSS.n271 VSS 0.00432979
R849 VSS.n246 VSS 0.00432979
R850 VSS.n249 VSS 0.00432979
R851 VSS.n253 VSS 0.00432979
R852 VSS.n394 VSS 0.00425
R853 VSS.n397 VSS 0.00425
R854 VSS.n400 VSS 0.00425
R855 VSS.n137 VSS 0.00417347
R856 VSS.n140 VSS 0.00417347
R857 VSS.n143 VSS 0.00417347
R858 VSS.n409 VSS 0.00417347
R859 VSS.n407 VSS 0.00417347
R860 VSS.n432 VSS.n431 0.00397181
R861 VSS VSS.n222 0.00380275
R862 VSS VSS.n316 0.00380275
R863 VSS VSS.n292 0.00380275
R864 VSS VSS.n175 0.00380275
R865 VSS.n38 VSS 0.00380275
R866 VSS.n46 VSS 0.00380275
R867 VSS.n206 VSS 0.00380275
R868 VSS.n204 VSS 0.00380275
R869 VSS VSS.n199 0.00380275
R870 VSS.n87 VSS 0.00380275
R871 VSS VSS.n166 0.00380275
R872 VSS VSS.n97 0.00380275
R873 VSS VSS.n122 0.00380275
R874 VSS VSS.n112 0.00380275
R875 VSS.n321 VSS 0.00380275
R876 VSS VSS.n295 0.00380275
R877 VSS VSS.n298 0.00380275
R878 VSS.n62 VSS 0.00352521
R879 VSS.n189 VSS 0.00352521
R880 VSS.n425 VSS 0.0035
R881 VSS.n411 VSS.n9 0.00324928
R882 VSS VSS.n274 0.00305319
R883 VSS VSS.n256 0.00305319
R884 VSS VSS.n43 0.00301748
R885 VSS VSS.n418 0.003
R886 VSS.n364 VSS.n363 0.00298619
R887 VSS.n146 VSS 0.00294898
R888 VSS.n379 VSS 0.00293243
R889 VSS VSS.n384 0.00293243
R890 VSS.n413 VSS 0.00233673
R891 VSS.n225 VSS 0.00219811
R892 VSS.n312 VSS 0.00219811
R893 VSS.n301 VSS 0.00219811
R894 VSS.n178 VSS 0.00219811
R895 VSS.n148 VSS 0.00219811
R896 VSS.n377 VSS 0.00219811
R897 VSS.n75 VSS 0.00219811
R898 VSS.n259 VSS 0.00219811
R899 VSS.n402 VSS 0.00219811
R900 VSS.n65 VSS 0.00219811
R901 VSS.n20 VSS 0.00219811
R902 VSS.n49 VSS 0.00219811
R903 VSS.n35 VSS 0.00219811
R904 VSS.n208 VSS 0.00219811
R905 VSS.n201 VSS 0.00219811
R906 VSS.n197 VSS 0.00219811
R907 VSS.n195 VSS 0.00219811
R908 VSS.n192 VSS 0.00219811
R909 VSS.n369 VSS 0.00215138
R910 VSS VSS.n356 0.00210237
R911 VSS VSS.n353 0.00210237
R912 VSS VSS.n343 0.00210237
R913 VSS VSS.n341 0.00210237
R914 VSS VSS.n331 0.00210237
R915 VSS VSS.n328 0.00210237
R916 VSS VSS.n430 0.00210237
R917 VSS VSS.n428 0.00210237
R918 VSS.n387 VSS 0.00171622
R919 VSS.n389 VSS 0.00171622
R920 VSS.n423 VSS 0.00157143
R921 VSS.n350 VSS 0.00156825
R922 VSS.n347 VSS 0.00156825
R923 VSS.n338 VSS 0.00156825
R924 VSS.n335 VSS 0.00156825
R925 VSS.n325 VSS 0.00156825
R926 VSS VSS.n0 0.00156825
R927 VSS.n374 VSS 0.0015
R928 VSS VSS.n361 0.00149448
R929 VSS.n364 VSS 0.00149448
R930 VSS VSS.n277 0.00136539
R931 VSS VSS.n60 0.0013
R932 VSS.n55 VSS.n23 0.00129295
R933 VSS VSS.n23 0.00129295
R934 VSS.n56 VSS.n55 0.000896476
R935 Vdiv110.n3 Vdiv110.n2 9.28805
R936 Vdiv110.n1 Vdiv110.n0 6.01414
R937 Vdiv110.n1 Vdiv110.t3 6.01414
R938 Vdiv110.n5 Vdiv110.n4 3.87405
R939 Vdiv110.n3 Vdiv110.n1 3.74829
R940 Vdiv110.n5 Vdiv110.n3 0.0422391
R941 Vdiv110 Vdiv110.n5 0.003
R942 VDD.t266 VDD.n150 57397.6
R943 VDD.t254 VDD.n207 57397.6
R944 VDD.n404 VDD.t456 2529.02
R945 VDD.n429 VDD 2301.38
R946 VDD.n411 VDD 2301.38
R947 VDD.n430 VDD.n429 1842.37
R948 VDD.n412 VDD.n411 1842.37
R949 VDD.n415 VDD.t152 1403.56
R950 VDD.n417 VDD.t302 1242.86
R951 VDD.n407 VDD.t452 1105.93
R952 VDD.n43 VDD.t403 1105.93
R953 VDD.n400 VDD.t415 1011.51
R954 VDD.t106 VDD.t326 961.905
R955 VDD.t62 VDD.t155 961.905
R956 VDD.t443 VDD.t228 961.905
R957 VDD.t172 VDD.t434 961.905
R958 VDD.t487 VDD.t44 961.905
R959 VDD.t18 VDD.t395 961.905
R960 VDD.n150 VDD.t48 864.287
R961 VDD.n12 VDD.t273 864.287
R962 VDD.n207 VDD.t30 864.287
R963 VDD.t243 VDD.n424 857.144
R964 VDD.t190 VDD.n421 857.144
R965 VDD.n429 VDD.t480 812.681
R966 VDD.n411 VDD.t290 812.681
R967 VDD.t393 VDD.t397 765.152
R968 VDD.t308 VDD.t98 765.152
R969 VDD.t474 VDD.t382 765.152
R970 VDD.t286 VDD.t129 765.152
R971 VDD.t230 VDD.t476 765.152
R972 VDD.t313 VDD.t367 765.152
R973 VDD.t81 VDD.t225 765.152
R974 VDD.t85 VDD.t304 765.152
R975 VDD.t420 VDD.t127 765.152
R976 VDD.t334 VDD.t90 765.152
R977 VDD.t292 VDD.t376 765.152
R978 VDD.t34 VDD.t318 765.152
R979 VDD.t93 VDD.t165 765.152
R980 VDD.t378 VDD.t295 765.152
R981 VDD.t150 VDD.t104 765.152
R982 VDD.t222 VDD.t446 765.152
R983 VDD.t306 VDD.t88 765.152
R984 VDD.t349 VDD.t83 765.152
R985 VDD.t132 VDD.t284 765.152
R986 VDD.t478 VDD.t233 765.152
R987 VDD.t430 VDD.t342 765.152
R988 VDD.t400 VDD.t112 765.152
R989 VDD.t96 VDD.t311 765.152
R990 VDD.t411 VDD.t235 765.152
R991 VDD.t484 VDD.t336 765.152
R992 VDD.t27 VDD.t36 765.152
R993 VDD.t465 VDD.t163 765.152
R994 VDD.t320 VDD.t440 765.152
R995 VDD.t275 VDD.t100 765.152
R996 VDD.t324 VDD.t300 765.152
R997 VDD.t372 VDD.t109 765.152
R998 VDD.t46 VDD.t418 765.152
R999 VDD.t271 VDD.t208 765.152
R1000 VDD.t32 VDD.t331 765.152
R1001 VDD.t135 VDD.t461 765.152
R1002 VDD.t322 VDD.t220 765.152
R1003 VDD.t328 VDD.t482 765.152
R1004 VDD.t463 VDD.t138 765.152
R1005 VDD.t160 VDD.t239 765.152
R1006 VDD.n40 VDD.t338 747.159
R1007 VDD.t340 VDD.t454 642.843
R1008 VDD.n408 VDD.t288 581.375
R1009 VDD VDD.n408 572.967
R1010 VDD.n468 VDD.t278 480.199
R1011 VDD.t405 VDD.t358 461.096
R1012 VDD.t152 VDD.t40 461.096
R1013 VDD.t152 VDD.t347 461.096
R1014 VDD.t344 VDD.t356 461.096
R1015 VDD VDD.n361 429.187
R1016 VDD VDD.n378 429.187
R1017 VDD VDD.n442 429.187
R1018 VDD VDD.n229 426.699
R1019 VDD VDD.n197 426.699
R1020 VDD VDD.n179 426.699
R1021 VDD VDD.n139 426.699
R1022 VDD.n55 VDD 424.618
R1023 VDD VDD.n49 424.618
R1024 VDD VDD.n44 422.557
R1025 VDD.n479 VDD.n478 421.611
R1026 VDD.n400 VDD.t450 420.793
R1027 VDD.n460 VDD.t280 386.365
R1028 VDD.n442 VDD.t237 386.365
R1029 VDD.n378 VDD.t470 386.365
R1030 VDD.n361 VDD.t0 386.365
R1031 VDD.n229 VDD.t257 386.365
R1032 VDD.n197 VDD.t188 386.365
R1033 VDD.n179 VDD.t260 386.365
R1034 VDD.n139 VDD.t436 386.365
R1035 VDD.n55 VDD.t60 386.365
R1036 VDD.n49 VDD.t25 386.365
R1037 VDD.t416 VDD.t54 380.952
R1038 VDD.t169 VDD.t62 380.952
R1039 VDD.t390 VDD.t102 380.952
R1040 VDD.t22 VDD.t172 380.952
R1041 VDD.t38 VDD.t250 380.952
R1042 VDD.t73 VDD.t18 380.952
R1043 VDD.t67 VDD.n55 378.788
R1044 VDD.n49 VDD.t176 378.788
R1045 VDD.n44 VDD.t64 378.788
R1046 VDD.t353 VDD.n463 375
R1047 VDD.n461 VDD.n460 368.159
R1048 VDD.n429 VDD.t405 351.586
R1049 VDD.n411 VDD.t344 351.586
R1050 VDD.n463 VDD.n462 343.137
R1051 VDD.t371 VDD.n479 306.118
R1052 VDD.t382 VDD.t117 303.031
R1053 VDD.t367 VDD.t215 303.031
R1054 VDD.t127 VDD.t212 303.031
R1055 VDD.t318 VDD.t122 303.031
R1056 VDD.t244 VDD.t378 303.031
R1057 VDD.t199 VDD.t150 303.031
R1058 VDD.t57 VDD.t306 303.031
R1059 VDD.t194 VDD.t349 303.031
R1060 VDD.t387 VDD.t478 303.031
R1061 VDD.t202 VDD.t430 303.031
R1062 VDD.t51 VDD.t96 303.031
R1063 VDD.t114 VDD.t411 303.031
R1064 VDD.t78 VDD.t465 303.031
R1065 VDD.t300 VDD.t12 303.031
R1066 VDD.t208 VDD.t179 303.031
R1067 VDD.t220 VDD.t9 303.031
R1068 VDD.t247 VDD.t463 303.031
R1069 VDD.t4 VDD.t160 303.031
R1070 VDD.n483 VDD.n467 298.536
R1071 VDD.n468 VDD.n467 288
R1072 VDD.n142 VDD.t70 242.857
R1073 VDD.n144 VDD.t106 242.857
R1074 VDD.t54 VDD.n147 242.857
R1075 VDD.n151 VDD.t169 242.857
R1076 VDD.n7 VDD.t182 242.857
R1077 VDD.n9 VDD.t443 242.857
R1078 VDD.n13 VDD.t390 242.857
R1079 VDD.n16 VDD.t22 242.857
R1080 VDD.n199 VDD.t15 242.857
R1081 VDD.n201 VDD.t487 242.857
R1082 VDD.t250 VDD.n204 242.857
R1083 VDD.n208 VDD.t73 242.857
R1084 VDD.n433 VDD.n425 199.562
R1085 VDD.n436 VDD.n422 199.562
R1086 VDD.n464 VDD.t353 193.183
R1087 VDD.n446 VDD.t384 193.183
R1088 VDD.n452 VDD.t397 193.183
R1089 VDD.n453 VDD.t308 193.183
R1090 VDD.n459 VDD.t117 193.183
R1091 VDD.n382 VDD.t364 193.183
R1092 VDD.n388 VDD.t129 193.183
R1093 VDD.n389 VDD.t230 193.183
R1094 VDD.n441 VDD.t215 193.183
R1095 VDD.n365 VDD.t191 193.183
R1096 VDD.n371 VDD.t225 193.183
R1097 VDD.n372 VDD.t85 193.183
R1098 VDD.n377 VDD.t212 193.183
R1099 VDD.n348 VDD.t315 193.183
R1100 VDD.n354 VDD.t90 193.183
R1101 VDD.n355 VDD.t292 193.183
R1102 VDD.n360 VDD.t122 193.183
R1103 VDD.n327 VDD.t145 193.183
R1104 VDD.n329 VDD.t93 193.183
R1105 VDD.n332 VDD.t244 193.183
R1106 VDD.n335 VDD.t199 193.183
R1107 VDD.n299 VDD.t360 193.183
R1108 VDD.n301 VDD.t222 193.183
R1109 VDD.n304 VDD.t57 193.183
R1110 VDD.n307 VDD.t194 193.183
R1111 VDD.n271 VDD.t425 193.183
R1112 VDD.n273 VDD.t132 193.183
R1113 VDD.n276 VDD.t387 193.183
R1114 VDD.n279 VDD.t202 193.183
R1115 VDD.n243 VDD.t408 193.183
R1116 VDD.n245 VDD.t400 193.183
R1117 VDD.n248 VDD.t51 193.183
R1118 VDD.n251 VDD.t114 193.183
R1119 VDD.n221 VDD.t467 193.183
R1120 VDD.n223 VDD.t484 193.183
R1121 VDD.n225 VDD.t27 193.183
R1122 VDD.n228 VDD.t78 193.183
R1123 VDD.n183 VDD.t297 193.183
R1124 VDD.n189 VDD.t440 193.183
R1125 VDD.n190 VDD.t275 193.183
R1126 VDD.n196 VDD.t12 193.183
R1127 VDD.n165 VDD.t205 193.183
R1128 VDD.n171 VDD.t109 193.183
R1129 VDD.n172 VDD.t46 193.183
R1130 VDD.n178 VDD.t179 193.183
R1131 VDD.n126 VDD.t185 193.183
R1132 VDD.n132 VDD.t331 193.183
R1133 VDD.n133 VDD.t135 193.183
R1134 VDD.n138 VDD.t9 193.183
R1135 VDD.n71 VDD.t157 193.183
R1136 VDD.n73 VDD.t328 193.183
R1137 VDD.n76 VDD.t247 193.183
R1138 VDD.n79 VDD.t4 193.183
R1139 VDD.n56 VDD.t67 193.183
R1140 VDD.n54 VDD.t176 193.183
R1141 VDD.n48 VDD.t64 193.183
R1142 VDD.n482 VDD.t423 191.288
R1143 VDD.t415 VDD.t422 175.631
R1144 VDD.t460 VDD.t162 175.631
R1145 VDD.n425 VDD.t243 170.577
R1146 VDD.n425 VDD.t140 170.577
R1147 VDD.n422 VDD.t190 170.577
R1148 VDD.n422 VDD.t380 170.577
R1149 VDD.t456 VDD.n403 153.678
R1150 VDD.t338 VDD.n39 153.678
R1151 VDD.t423 VDD.t142 151.516
R1152 VDD.t326 VDD.n142 138.095
R1153 VDD.t48 VDD.n144 138.095
R1154 VDD.t155 VDD.n147 138.095
R1155 VDD.n151 VDD.t266 138.095
R1156 VDD.t228 VDD.n7 138.095
R1157 VDD.t273 VDD.n9 138.095
R1158 VDD.t434 VDD.n13 138.095
R1159 VDD.n16 VDD.t269 138.095
R1160 VDD.t44 VDD.n199 138.095
R1161 VDD.t30 VDD.n201 138.095
R1162 VDD.t395 VDD.n204 138.095
R1163 VDD.n208 VDD.t254 138.095
R1164 VDD.n463 VDD.t490 132.353
R1165 VDD.n480 VDD.t438 124.511
R1166 VDD.n483 VDD.n482 117.216
R1167 VDD.n462 VDD.n461 112.746
R1168 VDD.n464 VDD.t148 109.849
R1169 VDD.n446 VDD.t393 109.849
R1170 VDD.t98 VDD.n452 109.849
R1171 VDD.n453 VDD.t474 109.849
R1172 VDD.t280 VDD.n459 109.849
R1173 VDD.n382 VDD.t286 109.849
R1174 VDD.t476 VDD.n388 109.849
R1175 VDD.n389 VDD.t313 109.849
R1176 VDD.t237 VDD.n441 109.849
R1177 VDD.n365 VDD.t81 109.849
R1178 VDD.t304 VDD.n371 109.849
R1179 VDD.n372 VDD.t420 109.849
R1180 VDD.t470 VDD.n377 109.849
R1181 VDD.n348 VDD.t334 109.849
R1182 VDD.t376 VDD.n354 109.849
R1183 VDD.n355 VDD.t34 109.849
R1184 VDD.t0 VDD.n360 109.849
R1185 VDD.t165 VDD.n327 109.849
R1186 VDD.t295 VDD.n329 109.849
R1187 VDD.t104 VDD.n332 109.849
R1188 VDD.n335 VDD.t2 109.849
R1189 VDD.t446 VDD.n299 109.849
R1190 VDD.t88 VDD.n301 109.849
R1191 VDD.t83 VDD.n304 109.849
R1192 VDD.n307 VDD.t472 109.849
R1193 VDD.t284 VDD.n271 109.849
R1194 VDD.t233 VDD.n273 109.849
R1195 VDD.t342 VDD.n276 109.849
R1196 VDD.n279 VDD.t374 109.849
R1197 VDD.t112 VDD.n243 109.849
R1198 VDD.t311 VDD.n245 109.849
R1199 VDD.t235 VDD.n248 109.849
R1200 VDD.n251 VDD.t282 109.849
R1201 VDD.t336 VDD.n221 109.849
R1202 VDD.t36 VDD.n223 109.849
R1203 VDD.t163 VDD.n225 109.849
R1204 VDD.t257 VDD.n228 109.849
R1205 VDD.n183 VDD.t320 109.849
R1206 VDD.t100 VDD.n189 109.849
R1207 VDD.n190 VDD.t324 109.849
R1208 VDD.t188 VDD.n196 109.849
R1209 VDD.n165 VDD.t372 109.849
R1210 VDD.t418 VDD.n171 109.849
R1211 VDD.n172 VDD.t271 109.849
R1212 VDD.t260 VDD.n178 109.849
R1213 VDD.n126 VDD.t32 109.849
R1214 VDD.t461 VDD.n132 109.849
R1215 VDD.n133 VDD.t322 109.849
R1216 VDD.t436 VDD.n138 109.849
R1217 VDD.t482 VDD.n71 109.849
R1218 VDD.t138 VDD.n73 109.849
R1219 VDD.t239 VDD.n76 109.849
R1220 VDD.n79 VDD.t263 109.849
R1221 VDD.n56 VDD.t174 109.849
R1222 VDD.t60 VDD.n54 109.849
R1223 VDD.t25 VDD.n48 109.849
R1224 VDD.n150 VDD.t416 97.6195
R1225 VDD.t102 VDD.n12 97.6195
R1226 VDD.n207 VDD.t38 97.6195
R1227 VDD.t142 VDD.n475 96.5914
R1228 VDD.n481 VDD.n480 90.2261
R1229 VDD.n408 VDD.t448 80.0005
R1230 VDD.n481 VDD.t371 76.2337
R1231 VDD.t302 VDD 68.2053
R1232 VDD VDD.n400 65.7064
R1233 VDD.n229 VDD.t76 62.1896
R1234 VDD.n197 VDD.t20 62.1896
R1235 VDD.n179 VDD.t167 62.1896
R1236 VDD.n139 VDD.t7 62.1896
R1237 VDD.n417 VDD.t428 61.9053
R1238 VDD.n55 VDD.t369 61.8817
R1239 VDD.n49 VDD.t218 61.8817
R1240 VDD.n44 VDD.t340 61.5769
R1241 VDD.n461 VDD 61.0269
R1242 VDD.n460 VDD.t42 59.702
R1243 VDD.n442 VDD.t120 59.702
R1244 VDD.n378 VDD.t197 59.702
R1245 VDD.n361 VDD.t210 59.702
R1246 VDD.n479 VDD.t241 59.4064
R1247 VDD.n404 VDD.t452 55.0852
R1248 VDD.t288 VDD.n407 55.0852
R1249 VDD.n40 VDD.t403 55.0852
R1250 VDD.t454 VDD.n43 55.0852
R1251 VDD.n475 VDD.t351 54.9247
R1252 VDD.n109 VDD.t262 30.9379
R1253 VDD.n81 VDD.t268 30.9379
R1254 VDD.n100 VDD.t259 30.7203
R1255 VDD.n87 VDD.t256 30.7203
R1256 VDD.n105 VDD.t265 30.2877
R1257 VDD.n93 VDD.t253 29.1661
R1258 VDD.n105 VDD.t497 24.9141
R1259 VDD.n109 VDD.t492 24.5101
R1260 VDD.n95 VDD.t494 24.5101
R1261 VDD.n81 VDD.t496 24.5101
R1262 VDD.n87 VDD.t495 24.4814
R1263 VDD.n100 VDD.t493 24.4814
R1264 VDD.n403 VDD.t422 21.9544
R1265 VDD.n39 VDD.t460 21.9544
R1266 VDD.n482 VDD.n481 20.147
R1267 VDD.n405 VDD.t453 12.3869
R1268 VDD.n393 VDD.t303 12.3869
R1269 VDD.n41 VDD.t404 12.3869
R1270 VDD.n485 VDD.n484 9.64171
R1271 VDD.n95 VDD.n94 8.0005
R1272 VDD.n93 VDD.n92 8.0005
R1273 VDD.n478 VDD.n477 7.01389
R1274 VDD.n486 VDD.n485 6.69176
R1275 VDD.n110 VDD.n108 6.39748
R1276 VDD.n39 VDD 6.30126
R1277 VDD VDD.n483 6.3005
R1278 VDD VDD.n468 6.3005
R1279 VDD.n488 VDD.n467 6.3005
R1280 VDD.n424 VDD 6.3005
R1281 VDD.n421 VDD 6.3005
R1282 VDD.n403 VDD.n402 6.3005
R1283 VDD VDD.n404 6.3005
R1284 VDD.n407 VDD.n406 6.3005
R1285 VDD.n418 VDD.n417 6.3005
R1286 VDD.n336 VDD.n335 6.3005
R1287 VDD.n339 VDD.n332 6.3005
R1288 VDD.n342 VDD.n329 6.3005
R1289 VDD.n345 VDD.n327 6.3005
R1290 VDD.n349 VDD.n348 6.3005
R1291 VDD.n354 VDD.n353 6.3005
R1292 VDD.n356 VDD.n355 6.3005
R1293 VDD.n360 VDD.n359 6.3005
R1294 VDD.n308 VDD.n307 6.3005
R1295 VDD.n311 VDD.n304 6.3005
R1296 VDD.n314 VDD.n301 6.3005
R1297 VDD.n317 VDD.n299 6.3005
R1298 VDD.n366 VDD.n365 6.3005
R1299 VDD.n371 VDD.n370 6.3005
R1300 VDD.n373 VDD.n372 6.3005
R1301 VDD.n377 VDD.n376 6.3005
R1302 VDD.n280 VDD.n279 6.3005
R1303 VDD.n283 VDD.n276 6.3005
R1304 VDD.n286 VDD.n273 6.3005
R1305 VDD.n289 VDD.n271 6.3005
R1306 VDD.n383 VDD.n382 6.3005
R1307 VDD.n388 VDD.n387 6.3005
R1308 VDD.n390 VDD.n389 6.3005
R1309 VDD.n441 VDD.n440 6.3005
R1310 VDD.n252 VDD.n251 6.3005
R1311 VDD.n255 VDD.n248 6.3005
R1312 VDD.n258 VDD.n245 6.3005
R1313 VDD.n261 VDD.n243 6.3005
R1314 VDD.n447 VDD.n446 6.3005
R1315 VDD.n452 VDD.n451 6.3005
R1316 VDD.n454 VDD.n453 6.3005
R1317 VDD.n459 VDD.n458 6.3005
R1318 VDD.n462 VDD 6.3005
R1319 VDD.n465 VDD.n464 6.3005
R1320 VDD.n504 VDD.n221 6.3005
R1321 VDD.n501 VDD.n223 6.3005
R1322 VDD.n498 VDD.n225 6.3005
R1323 VDD.n495 VDD.n228 6.3005
R1324 VDD.n123 VDD.n71 6.3005
R1325 VDD.n120 VDD.n73 6.3005
R1326 VDD.n117 VDD.n76 6.3005
R1327 VDD.n114 VDD.n79 6.3005
R1328 VDD.n127 VDD.n126 6.3005
R1329 VDD.n132 VDD.n131 6.3005
R1330 VDD.n134 VDD.n133 6.3005
R1331 VDD.n138 VDD.n137 6.3005
R1332 VDD.n161 VDD.n142 6.3005
R1333 VDD.n158 VDD.n144 6.3005
R1334 VDD.n155 VDD.n147 6.3005
R1335 VDD.n152 VDD.n151 6.3005
R1336 VDD.n166 VDD.n165 6.3005
R1337 VDD.n171 VDD.n170 6.3005
R1338 VDD.n173 VDD.n172 6.3005
R1339 VDD VDD.n40 6.3005
R1340 VDD.n43 VDD.n42 6.3005
R1341 VDD.n48 VDD.n47 6.3005
R1342 VDD.n54 VDD.n53 6.3005
R1343 VDD.n57 VDD.n56 6.3005
R1344 VDD.n178 VDD.n177 6.3005
R1345 VDD.n26 VDD.n7 6.3005
R1346 VDD.n23 VDD.n9 6.3005
R1347 VDD.n20 VDD.n13 6.3005
R1348 VDD.n17 VDD.n16 6.3005
R1349 VDD.n184 VDD.n183 6.3005
R1350 VDD.n189 VDD.n188 6.3005
R1351 VDD.n191 VDD.n190 6.3005
R1352 VDD.n196 VDD.n195 6.3005
R1353 VDD.n218 VDD.n199 6.3005
R1354 VDD.n215 VDD.n201 6.3005
R1355 VDD.n212 VDD.n204 6.3005
R1356 VDD.n209 VDD.n208 6.3005
R1357 VDD.n439 VDD.n438 5.69603
R1358 VDD.n98 VDD.n97 5.30733
R1359 VDD.n336 VDD.t3 5.213
R1360 VDD.n308 VDD.t473 5.213
R1361 VDD.n280 VDD.t375 5.213
R1362 VDD.n252 VDD.t283 5.213
R1363 VDD.n152 VDD.t267 5.213
R1364 VDD.n17 VDD.t270 5.213
R1365 VDD.n209 VDD.t255 5.213
R1366 VDD.n174 VDD.t272 5.16792
R1367 VDD.n466 VDD.t149 5.15377
R1368 VDD.n472 VDD.n471 5.13287
R1369 VDD.n473 VDD.t363 5.13287
R1370 VDD.n473 VDD.t352 5.13287
R1371 VDD.n431 VDD.t359 5.13287
R1372 VDD.n427 VDD.n426 5.13287
R1373 VDD.n413 VDD.t357 5.13287
R1374 VDD.n397 VDD.n396 5.13287
R1375 VDD.n416 VDD.t348 5.13287
R1376 VDD.n319 VDD.t1 5.13287
R1377 VDD.n357 VDD.t35 5.13287
R1378 VDD.n323 VDD.n322 5.13287
R1379 VDD.n352 VDD.t377 5.13287
R1380 VDD.n351 VDD.n324 5.13287
R1381 VDD.n350 VDD.t335 5.13287
R1382 VDD.n347 VDD.n325 5.13287
R1383 VDD.n338 VDD.t105 5.13287
R1384 VDD.n341 VDD.t296 5.13287
R1385 VDD.n343 VDD.n328 5.13287
R1386 VDD.n344 VDD.t166 5.13287
R1387 VDD.n346 VDD.n326 5.13287
R1388 VDD.n310 VDD.t84 5.13287
R1389 VDD.n313 VDD.t89 5.13287
R1390 VDD.n315 VDD.n300 5.13287
R1391 VDD.n316 VDD.t447 5.13287
R1392 VDD.n318 VDD.n298 5.13287
R1393 VDD.n291 VDD.t471 5.13287
R1394 VDD.n374 VDD.t421 5.13287
R1395 VDD.n295 VDD.n294 5.13287
R1396 VDD.n369 VDD.t305 5.13287
R1397 VDD.n368 VDD.n296 5.13287
R1398 VDD.n367 VDD.t82 5.13287
R1399 VDD.n364 VDD.n297 5.13287
R1400 VDD.n263 VDD.t238 5.13287
R1401 VDD.n391 VDD.t314 5.13287
R1402 VDD.n267 VDD.n266 5.13287
R1403 VDD.n386 VDD.t477 5.13287
R1404 VDD.n385 VDD.n268 5.13287
R1405 VDD.n384 VDD.t287 5.13287
R1406 VDD.n381 VDD.n269 5.13287
R1407 VDD.n282 VDD.t343 5.13287
R1408 VDD.n285 VDD.t234 5.13287
R1409 VDD.n287 VDD.n272 5.13287
R1410 VDD.n288 VDD.t285 5.13287
R1411 VDD.n290 VDD.n270 5.13287
R1412 VDD.n457 VDD.t281 5.13287
R1413 VDD.n455 VDD.t475 5.13287
R1414 VDD.n239 VDD.n238 5.13287
R1415 VDD.n450 VDD.t99 5.13287
R1416 VDD.n449 VDD.n240 5.13287
R1417 VDD.n448 VDD.t394 5.13287
R1418 VDD.n445 VDD.n241 5.13287
R1419 VDD.n254 VDD.t236 5.13287
R1420 VDD.n257 VDD.t312 5.13287
R1421 VDD.n259 VDD.n244 5.13287
R1422 VDD.n260 VDD.t113 5.13287
R1423 VDD.n262 VDD.n242 5.13287
R1424 VDD.n233 VDD.n232 5.13287
R1425 VDD.n505 VDD.n220 5.13287
R1426 VDD.n503 VDD.t337 5.13287
R1427 VDD.n502 VDD.n222 5.13287
R1428 VDD.n500 VDD.t37 5.13287
R1429 VDD.n499 VDD.n224 5.13287
R1430 VDD.n497 VDD.t164 5.13287
R1431 VDD.n494 VDD.t258 5.13287
R1432 VDD.n124 VDD.n70 5.13287
R1433 VDD.n122 VDD.t483 5.13287
R1434 VDD.n121 VDD.n72 5.13287
R1435 VDD.n119 VDD.t139 5.13287
R1436 VDD.n116 VDD.t240 5.13287
R1437 VDD.n125 VDD.n69 5.13287
R1438 VDD.n128 VDD.t33 5.13287
R1439 VDD.n129 VDD.n68 5.13287
R1440 VDD.n130 VDD.t462 5.13287
R1441 VDD.n67 VDD.n66 5.13287
R1442 VDD.n135 VDD.t323 5.13287
R1443 VDD.n63 VDD.t437 5.13287
R1444 VDD.n162 VDD.n141 5.13287
R1445 VDD.n160 VDD.t327 5.13287
R1446 VDD.n159 VDD.n143 5.13287
R1447 VDD.n157 VDD.t49 5.13287
R1448 VDD.n154 VDD.t156 5.13287
R1449 VDD.n164 VDD.n62 5.13287
R1450 VDD.n167 VDD.t373 5.13287
R1451 VDD.n168 VDD.n61 5.13287
R1452 VDD.n169 VDD.t419 5.13287
R1453 VDD.n60 VDD.n59 5.13287
R1454 VDD.n28 VDD.t261 5.13287
R1455 VDD.n46 VDD.n36 5.13287
R1456 VDD.n35 VDD.t26 5.13287
R1457 VDD.n51 VDD.n34 5.13287
R1458 VDD.n52 VDD.t61 5.13287
R1459 VDD.n32 VDD.n31 5.13287
R1460 VDD.n58 VDD.t175 5.13287
R1461 VDD.n27 VDD.n6 5.13287
R1462 VDD.n25 VDD.t229 5.13287
R1463 VDD.n24 VDD.n8 5.13287
R1464 VDD.n22 VDD.t274 5.13287
R1465 VDD.n19 VDD.t435 5.13287
R1466 VDD.n182 VDD.n5 5.13287
R1467 VDD.n185 VDD.t321 5.13287
R1468 VDD.n186 VDD.n4 5.13287
R1469 VDD.n187 VDD.t101 5.13287
R1470 VDD.n3 VDD.n2 5.13287
R1471 VDD.n192 VDD.t325 5.13287
R1472 VDD.n194 VDD.t189 5.13287
R1473 VDD.n219 VDD.n198 5.13287
R1474 VDD.n217 VDD.t45 5.13287
R1475 VDD.n216 VDD.n200 5.13287
R1476 VDD.n214 VDD.t31 5.13287
R1477 VDD.n211 VDD.t396 5.13287
R1478 VDD.n37 VDD.t455 5.09836
R1479 VDD.n398 VDD.t289 5.0955
R1480 VDD.n484 VDD.t439 5.09407
R1481 VDD.n486 VDD.t279 5.09407
R1482 VDD.n428 VDD.t481 5.09407
R1483 VDD.n423 VDD.t126 5.09407
R1484 VDD.n420 VDD.t459 5.09407
R1485 VDD.n401 VDD.t451 5.09407
R1486 VDD.n409 VDD.t449 5.09407
R1487 VDD.n410 VDD.t291 5.09407
R1488 VDD.n362 VDD.t211 5.09407
R1489 VDD.n379 VDD.t198 5.09407
R1490 VDD.n443 VDD.t121 5.09407
R1491 VDD.n235 VDD.t43 5.09407
R1492 VDD.n234 VDD.t491 5.09407
R1493 VDD.n476 VDD.t242 5.09407
R1494 VDD.n493 VDD.t77 5.09407
R1495 VDD.n140 VDD.t8 5.09407
R1496 VDD.n45 VDD.t341 5.09407
R1497 VDD.n50 VDD.t219 5.09407
R1498 VDD.n33 VDD.t370 5.09407
R1499 VDD.n180 VDD.t168 5.09407
R1500 VDD.n507 VDD.t21 5.09407
R1501 VDD.n493 VDD.n492 4.97776
R1502 VDD.n419 VDD.t429 4.9655
R1503 VDD.n478 VDD 4.91677
R1504 VDD.n113 VDD.t264 4.8755
R1505 VDD.n108 VDD.n98 4.84121
R1506 VDD.n490 VDD.n230 4.5005
R1507 VDD.n492 VDD.n491 4.5005
R1508 VDD.n88 VDD.n86 4.5005
R1509 VDD.n89 VDD.n86 4.5005
R1510 VDD.n82 VDD.n80 4.5005
R1511 VDD.n83 VDD.n80 4.5005
R1512 VDD.n101 VDD.n99 4.5005
R1513 VDD.n102 VDD.n99 4.5005
R1514 VDD.n424 VDD.t125 4.26489
R1515 VDD.n421 VDD.t458 4.26489
R1516 VDD.n432 VDD.t141 4.12326
R1517 VDD.n435 VDD.t381 4.12326
R1518 VDD.n487 VDD.t433 4.11379
R1519 VDD.n38 VDD.t339 3.94862
R1520 VDD.n399 VDD.t457 3.94479
R1521 VDD.n363 VDD.n318 3.90405
R1522 VDD.n475 VDD.n474 3.15287
R1523 VDD.n110 VDD.n109 2.88182
R1524 VDD.n96 VDD.n95 2.88074
R1525 VDD.n472 VDD.n470 2.85787
R1526 VDD.n414 VDD.n395 2.85787
R1527 VDD.n358 VDD.n321 2.85787
R1528 VDD.n337 VDD.n334 2.85787
R1529 VDD.n340 VDD.n331 2.85787
R1530 VDD.n309 VDD.n306 2.85787
R1531 VDD.n312 VDD.n303 2.85787
R1532 VDD.n375 VDD.n293 2.85787
R1533 VDD.n392 VDD.n265 2.85787
R1534 VDD.n281 VDD.n278 2.85787
R1535 VDD.n284 VDD.n275 2.85787
R1536 VDD.n456 VDD.n237 2.85787
R1537 VDD.n253 VDD.n250 2.85787
R1538 VDD.n256 VDD.n247 2.85787
R1539 VDD.n496 VDD.n227 2.85787
R1540 VDD.n118 VDD.n75 2.85787
R1541 VDD.n115 VDD.n78 2.85787
R1542 VDD.n136 VDD.n65 2.85787
R1543 VDD.n156 VDD.n146 2.85787
R1544 VDD.n153 VDD.n149 2.85787
R1545 VDD.n176 VDD.n30 2.85787
R1546 VDD.n21 VDD.n11 2.85787
R1547 VDD.n18 VDD.n15 2.85787
R1548 VDD.n193 VDD.n1 2.85787
R1549 VDD.n213 VDD.n203 2.85787
R1550 VDD.n210 VDD.n206 2.85787
R1551 VDD.n470 VDD.t424 2.2755
R1552 VDD.n470 VDD.n469 2.2755
R1553 VDD.n395 VDD.t41 2.2755
R1554 VDD.n395 VDD.n394 2.2755
R1555 VDD.n321 VDD.t319 2.2755
R1556 VDD.n321 VDD.n320 2.2755
R1557 VDD.n334 VDD.t151 2.2755
R1558 VDD.n334 VDD.n333 2.2755
R1559 VDD.n331 VDD.t379 2.2755
R1560 VDD.n331 VDD.n330 2.2755
R1561 VDD.n306 VDD.t350 2.2755
R1562 VDD.n306 VDD.n305 2.2755
R1563 VDD.n303 VDD.t307 2.2755
R1564 VDD.n303 VDD.n302 2.2755
R1565 VDD.n293 VDD.t128 2.2755
R1566 VDD.n293 VDD.n292 2.2755
R1567 VDD.n265 VDD.t368 2.2755
R1568 VDD.n265 VDD.n264 2.2755
R1569 VDD.n278 VDD.t431 2.2755
R1570 VDD.n278 VDD.n277 2.2755
R1571 VDD.n275 VDD.t479 2.2755
R1572 VDD.n275 VDD.n274 2.2755
R1573 VDD.n237 VDD.t383 2.2755
R1574 VDD.n237 VDD.n236 2.2755
R1575 VDD.n250 VDD.t412 2.2755
R1576 VDD.n250 VDD.n249 2.2755
R1577 VDD.n247 VDD.t97 2.2755
R1578 VDD.n247 VDD.n246 2.2755
R1579 VDD.n227 VDD.t466 2.2755
R1580 VDD.n227 VDD.n226 2.2755
R1581 VDD.n75 VDD.t464 2.2755
R1582 VDD.n75 VDD.n74 2.2755
R1583 VDD.n78 VDD.t161 2.2755
R1584 VDD.n78 VDD.n77 2.2755
R1585 VDD.n65 VDD.t221 2.2755
R1586 VDD.n65 VDD.n64 2.2755
R1587 VDD.n146 VDD.t417 2.2755
R1588 VDD.n146 VDD.n145 2.2755
R1589 VDD.n149 VDD.t63 2.2755
R1590 VDD.n149 VDD.n148 2.2755
R1591 VDD.n30 VDD.t209 2.2755
R1592 VDD.n30 VDD.n29 2.2755
R1593 VDD.n11 VDD.t103 2.2755
R1594 VDD.n11 VDD.n10 2.2755
R1595 VDD.n15 VDD.t173 2.2755
R1596 VDD.n15 VDD.n14 2.2755
R1597 VDD.n1 VDD.t301 2.2755
R1598 VDD.n1 VDD.n0 2.2755
R1599 VDD.n203 VDD.t39 2.2755
R1600 VDD.n203 VDD.n202 2.2755
R1601 VDD.n206 VDD.t19 2.2755
R1602 VDD.n206 VDD.n205 2.2755
R1603 VDD.n457 VDD 2.25904
R1604 VDD.n91 VDD.n90 2.2439
R1605 VDD.n104 VDD.n103 2.2439
R1606 VDD.n85 VDD.n84 2.24362
R1607 VDD.n82 VDD.n81 2.12277
R1608 VDD.n402 VDD.n401 1.96666
R1609 VDD.n106 VDD.n105 1.82213
R1610 VDD VDD.n63 1.81785
R1611 VDD.n95 VDD.n93 1.77234
R1612 VDD.n97 VDD.n91 1.6239
R1613 VDD.n107 VDD.n104 1.6239
R1614 VDD.n231 VDD.n230 1.50339
R1615 VDD VDD.n38 1.44207
R1616 VDD.n101 VDD.n100 1.39846
R1617 VDD.n88 VDD.n87 1.39728
R1618 VDD.n125 VDD.n124 1.16167
R1619 VDD.n97 VDD.n96 1.12314
R1620 VDD.n107 VDD.n106 1.12224
R1621 VDD.n163 VDD.n162 1.07428
R1622 VDD.n380 VDD.n290 1.02928
R1623 VDD.n444 VDD.n262 1.02928
R1624 VDD.n181 VDD.n27 1.01882
R1625 VDD.n506 VDD.n219 1.01882
R1626 VDD VDD.n416 0.973239
R1627 VDD.n347 VDD.n346 0.881662
R1628 VDD.n480 VDD.t432 0.783764
R1629 VDD.n108 VDD.n107 0.52356
R1630 VDD.n98 VDD.n85 0.497812
R1631 VDD.n438 VDD.n437 0.493148
R1632 VDD.n432 VDD.n431 0.38985
R1633 VDD.n114 VDD.n113 0.337997
R1634 VDD.n175 VDD.n58 0.334229
R1635 VDD.n113 VDD.n112 0.333658
R1636 VDD.n341 VDD.n340 0.233919
R1637 VDD.n338 VDD.n337 0.233919
R1638 VDD.n313 VDD.n312 0.233919
R1639 VDD.n310 VDD.n309 0.233919
R1640 VDD.n285 VDD.n284 0.233919
R1641 VDD.n282 VDD.n281 0.233919
R1642 VDD.n257 VDD.n256 0.233919
R1643 VDD.n254 VDD.n253 0.233919
R1644 VDD.n119 VDD.n118 0.233919
R1645 VDD.n116 VDD.n115 0.233919
R1646 VDD.n157 VDD.n156 0.233919
R1647 VDD.n154 VDD.n153 0.233919
R1648 VDD.n22 VDD.n21 0.233919
R1649 VDD.n19 VDD.n18 0.233919
R1650 VDD.n214 VDD.n213 0.233919
R1651 VDD.n211 VDD.n210 0.233919
R1652 VDD.n489 VDD.n488 0.224447
R1653 VDD.n235 VDD 0.205357
R1654 VDD.n489 VDD.n466 0.202146
R1655 VDD VDD.n409 0.200279
R1656 VDD.n414 VDD.n413 0.199441
R1657 VDD VDD.n399 0.177304
R1658 VDD.n435 VDD.n434 0.173131
R1659 VDD.n428 VDD.n427 0.170231
R1660 VDD.n444 VDD.n443 0.167533
R1661 VDD VDD.n38 0.16613
R1662 VDD VDD.n291 0.160716
R1663 VDD VDD.n263 0.158984
R1664 VDD VDD.n319 0.157289
R1665 VDD.n380 VDD.n379 0.155496
R1666 VDD.n363 VDD.n362 0.154581
R1667 VDD.n164 VDD.n163 0.144547
R1668 VDD.n344 VDD.n343 0.141016
R1669 VDD.n316 VDD.n315 0.141016
R1670 VDD.n288 VDD.n287 0.141016
R1671 VDD.n260 VDD.n259 0.141016
R1672 VDD.n122 VDD.n121 0.141016
R1673 VDD.n129 VDD.n128 0.141016
R1674 VDD.n130 VDD.n67 0.141016
R1675 VDD.n160 VDD.n159 0.141016
R1676 VDD.n168 VDD.n167 0.141016
R1677 VDD.n169 VDD.n60 0.141016
R1678 VDD.n25 VDD.n24 0.141016
R1679 VDD.n217 VDD.n216 0.141016
R1680 VDD.n163 VDD.n140 0.138896
R1681 VDD.n434 VDD.n423 0.13637
R1682 VDD.n437 VDD.n420 0.13637
R1683 VDD.n364 VDD.n363 0.131861
R1684 VDD.n234 VDD.n233 0.130567
R1685 VDD.n368 VDD.n367 0.123551
R1686 VDD.n369 VDD.n295 0.123551
R1687 VDD.n449 VDD.n448 0.123551
R1688 VDD.n450 VDD.n239 0.123551
R1689 VDD VDD.n135 0.122435
R1690 VDD.n385 VDD.n384 0.122176
R1691 VDD.n386 VDD.n267 0.122176
R1692 VDD.n351 VDD.n350 0.120831
R1693 VDD.n352 VDD.n323 0.120831
R1694 VDD.n445 VDD.n444 0.116432
R1695 VDD.n381 VDD.n380 0.115137
R1696 VDD.n136 VDD 0.111984
R1697 VDD.n106 VDD 0.110941
R1698 VDD.n406 VDD.n405 0.107626
R1699 VDD.n430 VDD.n427 0.107339
R1700 VDD.n346 VDD.n345 0.107339
R1701 VDD.n343 VDD.n342 0.107339
R1702 VDD.n318 VDD.n317 0.107339
R1703 VDD.n315 VDD.n314 0.107339
R1704 VDD.n290 VDD.n289 0.107339
R1705 VDD.n287 VDD.n286 0.107339
R1706 VDD.n262 VDD.n261 0.107339
R1707 VDD.n259 VDD.n258 0.107339
R1708 VDD.n465 VDD.n233 0.107339
R1709 VDD.n124 VDD.n123 0.107339
R1710 VDD.n121 VDD.n120 0.107339
R1711 VDD.n127 VDD.n125 0.107339
R1712 VDD.n131 VDD.n129 0.107339
R1713 VDD.n134 VDD.n67 0.107339
R1714 VDD.n162 VDD.n161 0.107339
R1715 VDD.n159 VDD.n158 0.107339
R1716 VDD.n166 VDD.n164 0.107339
R1717 VDD.n170 VDD.n168 0.107339
R1718 VDD.n173 VDD.n60 0.107339
R1719 VDD.n27 VDD.n26 0.107339
R1720 VDD.n24 VDD.n23 0.107339
R1721 VDD.n219 VDD.n218 0.107339
R1722 VDD.n216 VDD.n215 0.107339
R1723 VDD VDD.n374 0.10728
R1724 VDD VDD.n455 0.10728
R1725 VDD.n340 VDD 0.106177
R1726 VDD.n337 VDD 0.106177
R1727 VDD.n312 VDD 0.106177
R1728 VDD.n309 VDD 0.106177
R1729 VDD.n284 VDD 0.106177
R1730 VDD.n281 VDD 0.106177
R1731 VDD.n256 VDD 0.106177
R1732 VDD.n253 VDD 0.106177
R1733 VDD.n118 VDD 0.106177
R1734 VDD.n115 VDD 0.106177
R1735 VDD VDD.n136 0.106177
R1736 VDD.n156 VDD 0.106177
R1737 VDD.n153 VDD 0.106177
R1738 VDD.n21 VDD 0.106177
R1739 VDD.n18 VDD 0.106177
R1740 VDD.n213 VDD 0.106177
R1741 VDD.n210 VDD 0.106177
R1742 VDD VDD.n391 0.106087
R1743 VDD VDD.n357 0.10492
R1744 VDD.n375 VDD 0.0981271
R1745 VDD.n456 VDD 0.0981271
R1746 VDD.n392 VDD 0.0970363
R1747 VDD.n358 VDD 0.0959696
R1748 VDD.n366 VDD.n364 0.0940593
R1749 VDD.n370 VDD.n368 0.0940593
R1750 VDD.n373 VDD.n295 0.0940593
R1751 VDD.n447 VDD.n445 0.0940593
R1752 VDD.n451 VDD.n449 0.0940593
R1753 VDD.n454 VDD.n239 0.0940593
R1754 VDD.n405 VDD 0.0930506
R1755 VDD VDD.n375 0.0930424
R1756 VDD VDD.n456 0.0930424
R1757 VDD.n383 VDD.n381 0.093014
R1758 VDD.n387 VDD.n385 0.093014
R1759 VDD.n390 VDD.n267 0.093014
R1760 VDD.n349 VDD.n347 0.0919917
R1761 VDD.n353 VDD.n351 0.0919917
R1762 VDD.n356 VDD.n323 0.0919917
R1763 VDD VDD.n358 0.0909972
R1764 VDD VDD.n35 0.0862422
R1765 VDD.n52 VDD 0.0862422
R1766 VDD VDD.n37 0.085945
R1767 VDD.n494 VDD 0.0854968
R1768 VDD VDD.n28 0.0854968
R1769 VDD.n94 VDD 0.0839415
R1770 VDD VDD.n398 0.0825482
R1771 VDD.n490 VDD.n489 0.0819374
R1772 VDD.n89 VDD 0.0816915
R1773 VDD.n339 VDD.n338 0.080629
R1774 VDD.n311 VDD.n310 0.080629
R1775 VDD.n283 VDD.n282 0.080629
R1776 VDD.n255 VDD.n254 0.080629
R1777 VDD.n117 VDD.n116 0.080629
R1778 VDD.n137 VDD.n63 0.080629
R1779 VDD.n155 VDD.n154 0.080629
R1780 VDD.n20 VDD.n19 0.080629
R1781 VDD.n212 VDD.n211 0.080629
R1782 VDD.n102 VDD 0.0805665
R1783 VDD VDD.n344 0.0794677
R1784 VDD VDD.n341 0.0794677
R1785 VDD VDD.n316 0.0794677
R1786 VDD VDD.n313 0.0794677
R1787 VDD VDD.n288 0.0794677
R1788 VDD VDD.n285 0.0794677
R1789 VDD VDD.n260 0.0794677
R1790 VDD VDD.n257 0.0794677
R1791 VDD VDD.n122 0.0794677
R1792 VDD VDD.n119 0.0794677
R1793 VDD.n128 VDD 0.0794677
R1794 VDD VDD.n130 0.0794677
R1795 VDD.n135 VDD 0.0794677
R1796 VDD VDD.n160 0.0794677
R1797 VDD VDD.n157 0.0794677
R1798 VDD.n167 VDD 0.0794677
R1799 VDD VDD.n169 0.0794677
R1800 VDD VDD.n25 0.0794677
R1801 VDD VDD.n22 0.0794677
R1802 VDD VDD.n217 0.0794677
R1803 VDD VDD.n214 0.0794677
R1804 VDD.n174 VDD 0.0765085
R1805 VDD.n431 VDD 0.0759839
R1806 VDD.n83 VDD 0.0738165
R1807 VDD.n112 VDD.n110 0.0725
R1808 VDD.n484 VDD 0.0709717
R1809 VDD VDD.n428 0.0709717
R1810 VDD VDD.n423 0.0709717
R1811 VDD VDD.n420 0.0709717
R1812 VDD VDD.n235 0.0709717
R1813 VDD.n476 VDD 0.0709717
R1814 VDD.n140 VDD 0.0709717
R1815 VDD.n376 VDD.n291 0.0706695
R1816 VDD.n458 VDD.n457 0.0706695
R1817 VDD.n440 VDD.n263 0.0698855
R1818 VDD.n410 VDD.n397 0.0697857
R1819 VDD.n367 VDD 0.0696525
R1820 VDD VDD.n369 0.0696525
R1821 VDD.n374 VDD 0.0696525
R1822 VDD.n448 VDD 0.0696525
R1823 VDD VDD.n450 0.0696525
R1824 VDD.n455 VDD 0.0696525
R1825 VDD.n359 VDD.n319 0.0691188
R1826 VDD.n384 VDD 0.0688799
R1827 VDD VDD.n386 0.0688799
R1828 VDD.n391 VDD 0.0688799
R1829 VDD.n350 VDD 0.0681243
R1830 VDD VDD.n352 0.0681243
R1831 VDD.n357 VDD 0.0681243
R1832 VDD.n111 VDD 0.0659545
R1833 VDD.n503 VDD.n502 0.0647478
R1834 VDD.n500 VDD.n499 0.0647478
R1835 VDD.n186 VDD.n185 0.0647478
R1836 VDD.n187 VDD.n3 0.0647478
R1837 VDD.n418 VDD.n393 0.064413
R1838 VDD.n46 VDD.n45 0.0630764
R1839 VDD.n51 VDD.n50 0.0630764
R1840 VDD.n33 VDD.n32 0.0630764
R1841 VDD VDD.n398 0.062714
R1842 VDD.n42 VDD.n41 0.060911
R1843 VDD.n506 VDD.n505 0.0607039
R1844 VDD.n182 VDD.n181 0.0607039
R1845 VDD.n497 VDD 0.0562522
R1846 VDD VDD.n192 0.0562522
R1847 VDD VDD.n393 0.0557174
R1848 VDD VDD.n487 0.0555633
R1849 VDD.n412 VDD.n397 0.0551535
R1850 VDD VDD.n414 0.0551
R1851 VDD.n466 VDD 0.0550806
R1852 VDD.n434 VDD.n433 0.0545
R1853 VDD.n181 VDD.n180 0.0536232
R1854 VDD VDD.n472 0.0533387
R1855 VDD.n439 VDD.n392 0.0532933
R1856 VDD VDD.n399 0.0529202
R1857 VDD.n41 VDD 0.0526918
R1858 VDD VDD.n496 0.0514734
R1859 VDD.n176 VDD 0.0514734
R1860 VDD.n193 VDD 0.0514734
R1861 VDD.n47 VDD.n46 0.0497857
R1862 VDD.n53 VDD.n51 0.0497857
R1863 VDD.n57 VDD.n32 0.0497857
R1864 VDD.n505 VDD.n504 0.0493496
R1865 VDD.n502 VDD.n501 0.0493496
R1866 VDD.n499 VDD.n498 0.0493496
R1867 VDD.n184 VDD.n182 0.0493496
R1868 VDD.n188 VDD.n186 0.0493496
R1869 VDD.n191 VDD.n3 0.0493496
R1870 VDD.n496 VDD 0.0488186
R1871 VDD VDD.n176 0.0488186
R1872 VDD VDD.n193 0.0488186
R1873 VDD.n112 VDD.n111 0.0455
R1874 VDD VDD.n234 0.043431
R1875 VDD.n416 VDD.n415 0.0419
R1876 VDD.n379 VDD 0.0404465
R1877 VDD.n443 VDD 0.0400238
R1878 VDD.n362 VDD 0.0396099
R1879 VDD VDD.n439 0.0392151
R1880 VDD.n507 VDD 0.039182
R1881 VDD.n413 VDD 0.0391139
R1882 VDD VDD.n473 0.0382419
R1883 VDD.n194 VDD 0.0377891
R1884 VDD.n175 VDD.n174 0.0371957
R1885 VDD.n495 VDD.n494 0.0371372
R1886 VDD.n177 VDD.n28 0.0371372
R1887 VDD.n195 VDD.n194 0.0371372
R1888 VDD VDD.n503 0.0366062
R1889 VDD VDD.n500 0.0366062
R1890 VDD VDD.n497 0.0366062
R1891 VDD.n185 VDD 0.0366062
R1892 VDD VDD.n187 0.0366062
R1893 VDD.n192 VDD 0.0366062
R1894 VDD.n419 VDD 0.0363979
R1895 VDD VDD.n37 0.035637
R1896 VDD VDD.n35 0.0353214
R1897 VDD VDD.n52 0.0353214
R1898 VDD.n58 VDD 0.0353214
R1899 VDD.n485 VDD.n472 0.0344677
R1900 VDD.n477 VDD.n476 0.0327642
R1901 VDD VDD.n436 0.0325968
R1902 VDD VDD.n486 0.032019
R1903 VDD.n409 VDD 0.0305
R1904 VDD.n401 VDD 0.030261
R1905 VDD.n90 VDD.n89 0.0275
R1906 VDD.n94 VDD.n92 0.0275
R1907 VDD.n103 VDD.n102 0.026375
R1908 VDD.n91 VDD.n86 0.025705
R1909 VDD.n104 VDD.n99 0.025705
R1910 VDD.n438 VDD.n419 0.024997
R1911 VDD VDD.n410 0.0243658
R1912 VDD VDD.n432 0.0240135
R1913 VDD VDD.n435 0.0238871
R1914 VDD.n491 VDD.n490 0.0225755
R1915 VDD.n437 VDD 0.0221129
R1916 VDD.n45 VDD 0.0220896
R1917 VDD.n50 VDD 0.0220896
R1918 VDD VDD.n33 0.0220896
R1919 VDD VDD.n493 0.021904
R1920 VDD.n180 VDD 0.021904
R1921 VDD VDD.n507 0.021904
R1922 VDD VDD.n175 0.0214735
R1923 VDD.n84 VDD.n83 0.02075
R1924 VDD.n492 VDD.n230 0.0193811
R1925 VDD.n85 VDD.n80 0.0169383
R1926 VDD VDD.n506 0.0149413
R1927 VDD.n84 VDD.n82 0.0095
R1928 VDD.n111 VDD 0.00868182
R1929 VDD.n487 VDD 0.00543671
R1930 VDD VDD.n430 0.00514516
R1931 VDD VDD.n465 0.00514516
R1932 VDD.n103 VDD.n101 0.003875
R1933 VDD.n488 VDD 0.00315823
R1934 VDD VDD.n412 0.00287624
R1935 VDD.n474 VDD 0.00282258
R1936 VDD.n90 VDD.n88 0.00275
R1937 VDD.n47 VDD 0.00264286
R1938 VDD.n53 VDD 0.00264286
R1939 VDD VDD.n57 0.00264286
R1940 VDD.n96 VDD.n92 0.00171994
R1941 VDD.n345 VDD 0.00166129
R1942 VDD.n342 VDD 0.00166129
R1943 VDD VDD.n339 0.00166129
R1944 VDD VDD.n336 0.00166129
R1945 VDD.n317 VDD 0.00166129
R1946 VDD.n314 VDD 0.00166129
R1947 VDD VDD.n311 0.00166129
R1948 VDD VDD.n308 0.00166129
R1949 VDD.n289 VDD 0.00166129
R1950 VDD.n286 VDD 0.00166129
R1951 VDD VDD.n283 0.00166129
R1952 VDD VDD.n280 0.00166129
R1953 VDD.n261 VDD 0.00166129
R1954 VDD.n258 VDD 0.00166129
R1955 VDD VDD.n255 0.00166129
R1956 VDD VDD.n252 0.00166129
R1957 VDD.n123 VDD 0.00166129
R1958 VDD.n120 VDD 0.00166129
R1959 VDD VDD.n117 0.00166129
R1960 VDD VDD.n114 0.00166129
R1961 VDD VDD.n127 0.00166129
R1962 VDD.n131 VDD 0.00166129
R1963 VDD VDD.n134 0.00166129
R1964 VDD.n137 VDD 0.00166129
R1965 VDD.n161 VDD 0.00166129
R1966 VDD.n158 VDD 0.00166129
R1967 VDD VDD.n155 0.00166129
R1968 VDD VDD.n152 0.00166129
R1969 VDD VDD.n166 0.00166129
R1970 VDD.n170 VDD 0.00166129
R1971 VDD VDD.n173 0.00166129
R1972 VDD.n26 VDD 0.00166129
R1973 VDD.n23 VDD 0.00166129
R1974 VDD VDD.n20 0.00166129
R1975 VDD VDD.n17 0.00166129
R1976 VDD.n218 VDD 0.00166129
R1977 VDD.n215 VDD 0.00166129
R1978 VDD VDD.n212 0.00166129
R1979 VDD VDD.n209 0.00166129
R1980 VDD.n433 VDD 0.00163514
R1981 VDD.n436 VDD 0.00162903
R1982 VDD.n477 VDD.n231 0.00156548
R1983 VDD VDD.n366 0.00151695
R1984 VDD.n370 VDD 0.00151695
R1985 VDD VDD.n373 0.00151695
R1986 VDD.n376 VDD 0.00151695
R1987 VDD VDD.n447 0.00151695
R1988 VDD.n451 VDD 0.00151695
R1989 VDD VDD.n454 0.00151695
R1990 VDD.n458 VDD 0.00151695
R1991 VDD VDD.n383 0.00150559
R1992 VDD.n387 VDD 0.00150559
R1993 VDD VDD.n390 0.00150559
R1994 VDD.n440 VDD 0.00150559
R1995 VDD VDD.n349 0.00149448
R1996 VDD.n353 VDD 0.00149448
R1997 VDD VDD.n356 0.00149448
R1998 VDD.n359 VDD 0.00149448
R1999 VDD.n491 VDD.n231 0.00128347
R2000 VDD.n406 VDD 0.00122874
R2001 VDD.n415 VDD 0.0011
R2002 VDD.n474 VDD 0.00108064
R2003 VDD.n504 VDD 0.00103097
R2004 VDD.n501 VDD 0.00103097
R2005 VDD.n498 VDD 0.00103097
R2006 VDD VDD.n495 0.00103097
R2007 VDD.n177 VDD 0.00103097
R2008 VDD VDD.n184 0.00103097
R2009 VDD.n188 VDD 0.00103097
R2010 VDD VDD.n191 0.00103097
R2011 VDD.n195 VDD 0.00103097
R2012 VDD VDD.n418 0.000934783
R2013 VDD.n42 VDD 0.000910959
R2014 VDD.n402 VDD 0.000739362
R2015 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t3 30.9379
R2016 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n0 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t5 30.664
R2017 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n0 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t2 24.5385
R2018 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t4 24.5101
R2019 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n2 7.46763
R2020 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n3 5.28703
R2021 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n1 4.09208
R2022 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 3.12156
R2023 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 1.86016
R2024 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n0 1.4252
R2025 CLK_div_10_mag_0.JK_FF_mag_2.K.n2 CLK_div_10_mag_0.JK_FF_mag_2.K.t6 37.1981
R2026 CLK_div_10_mag_0.JK_FF_mag_2.K.n4 CLK_div_10_mag_0.JK_FF_mag_2.K.t3 31.528
R2027 CLK_div_10_mag_0.JK_FF_mag_2.K.n1 CLK_div_10_mag_0.JK_FF_mag_2.K.t7 30.5752
R2028 CLK_div_10_mag_0.JK_FF_mag_2.K.n1 CLK_div_10_mag_0.JK_FF_mag_2.K.t5 24.6493
R2029 CLK_div_10_mag_0.JK_FF_mag_2.K.n2 CLK_div_10_mag_0.JK_FF_mag_2.K.t8 17.6611
R2030 CLK_div_10_mag_0.JK_FF_mag_2.K.n3 CLK_div_10_mag_0.JK_FF_mag_2.K 17.0533
R2031 CLK_div_10_mag_0.JK_FF_mag_2.K.n4 CLK_div_10_mag_0.JK_FF_mag_2.K.t4 15.3826
R2032 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_2.K.n4 7.62758
R2033 CLK_div_10_mag_0.JK_FF_mag_2.K.n5 CLK_div_10_mag_0.JK_FF_mag_2.K.n3 3.28711
R2034 CLK_div_10_mag_0.JK_FF_mag_2.K.n0 CLK_div_10_mag_0.JK_FF_mag_2.K.n7 2.99416
R2035 CLK_div_10_mag_0.JK_FF_mag_2.K.n3 CLK_div_10_mag_0.JK_FF_mag_2.K 2.81128
R2036 CLK_div_10_mag_0.JK_FF_mag_2.K.n5 CLK_div_10_mag_0.JK_FF_mag_2.K 2.66613
R2037 CLK_div_10_mag_0.JK_FF_mag_2.K.n7 CLK_div_10_mag_0.JK_FF_mag_2.K.t1 2.2755
R2038 CLK_div_10_mag_0.JK_FF_mag_2.K.n7 CLK_div_10_mag_0.JK_FF_mag_2.K.n6 2.2755
R2039 CLK_div_10_mag_0.JK_FF_mag_2.K.n0 CLK_div_10_mag_0.JK_FF_mag_2.K.n5 2.2505
R2040 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_2.K.n1 1.80834
R2041 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_2.K.n2 1.43706
R2042 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_2.K.n0 0.281955
R2043 RST.n54 RST.t4 36.935
R2044 RST.n52 RST.t2 36.935
R2045 RST.n48 RST.t15 36.935
R2046 RST.n58 RST.t8 36.935
R2047 RST.n7 RST.t12 36.935
R2048 RST.n0 RST.t10 36.935
R2049 RST.n20 RST.t1 36.935
R2050 RST.n34 RST.t6 36.935
R2051 RST.n54 RST.t13 18.1962
R2052 RST.n52 RST.t7 18.1962
R2053 RST.n58 RST.t14 18.1962
R2054 RST.n7 RST.t11 18.1962
R2055 RST.n0 RST.t9 18.1962
R2056 RST.n20 RST.t0 18.1962
R2057 RST.n34 RST.t5 18.1962
R2058 RST.n49 RST.t3 16.3712
R2059 RST.n50 RST.n49 8.0005
R2060 RST.n56 RST.n55 5.39866
R2061 RST.n27 RST.n26 4.51211
R2062 RST.n44 RST.n43 4.5005
R2063 RST.n51 RST.n45 4.5005
R2064 RST.n51 RST.n50 4.5005
R2065 RST.n22 RST.n19 4.5005
R2066 RST.n22 RST.n21 4.5005
R2067 RST.n25 RST.n23 4.5005
R2068 RST.n25 RST.n24 4.5005
R2069 RST.n57 RST.n56 3.52872
R2070 RST RST.n57 3.47469
R2071 RST.n63 RST.n62 2.25544
R2072 RST.n10 RST.n9 2.2505
R2073 RST.n28 RST.n27 2.24707
R2074 RST.n55 RST.n54 2.13714
R2075 RST.n53 RST.n52 2.13714
R2076 RST.n59 RST.n58 2.1359
R2077 RST.n1 RST.n0 2.12318
R2078 RST.n21 RST.n20 2.12318
R2079 RST.n35 RST.n34 2.1224
R2080 RST.n8 RST.n7 2.12188
R2081 RST.n48 RST.n47 2.12075
R2082 RST.n15 RST.n14 1.90023
R2083 RST.n17 RST.n16 1.88263
R2084 RST.n56 RST.n53 1.8704
R2085 RST.n30 RST.n29 1.86678
R2086 RST.n63 RST.n61 1.83032
R2087 RST.n49 RST.n48 1.8255
R2088 RST.n60 RST.n59 1.76243
R2089 RST.n46 RST.n43 1.51223
R2090 RST.n37 RST.n36 1.5005
R2091 RST.n39 RST.n38 1.5005
R2092 RST.n13 RST.n12 1.5005
R2093 RST.n16 RST.n4 1.13307
R2094 RST.n57 RST.n51 1.1235
R2095 RST.n3 RST.n2 0.898107
R2096 RST.n61 RST.n42 0.839477
R2097 RST.n42 RST.n41 0.627203
R2098 RST.n61 RST.n60 0.388998
R2099 RST.n59 RST 0.0687763
R2100 RST.n53 RST 0.0675415
R2101 RST.n55 RST 0.0675409
R2102 RST.n60 RST 0.0544779
R2103 RST.n2 RST 0.0518307
R2104 RST.n44 RST 0.0394837
R2105 RST.n46 RST.n45 0.0367013
R2106 RST.n33 RST 0.0363802
R2107 RST.n9 RST.n6 0.0361897
R2108 RST.n36 RST.n33 0.0346379
R2109 RST.n6 RST 0.031725
R2110 RST.n2 RST.n1 0.0249551
R2111 RST.n23 RST 0.0239664
R2112 RST.n22 RST.n18 0.0236959
R2113 RST.n14 RST.n13 0.0205676
R2114 RST.n39 RST.n30 0.0193514
R2115 RST.n38 RST.n31 0.0181289
R2116 RST.n29 RST.n28 0.0144865
R2117 RST.n27 RST.n25 0.0130264
R2118 RST.n9 RST.n8 0.0129138
R2119 RST.n16 RST.n15 0.0117735
R2120 RST.n10 RST.n5 0.0116103
R2121 RST.n36 RST.n35 0.00825862
R2122 RST.n28 RST.n17 0.0077973
R2123 RST RST.n63 0.00543902
R2124 RST.n47 RST.n46 0.00540913
R2125 RST.n12 RST.n11 0.00513918
R2126 RST.n37 RST.n32 0.00513918
R2127 RST.n51 RST.n43 0.003875
R2128 RST.n12 RST.n10 0.00328351
R2129 RST.n4 RST.n3 0.00328351
R2130 RST.n38 RST.n37 0.00328351
R2131 RST.n40 RST.n39 0.00232432
R2132 RST.n41 RST.n40 0.00232432
R2133 RST.n45 RST.n44 0.00205172
R2134 RST.n50 RST.n47 0.00173095
R2135 RST.n25 RST.n22 0.00142783
R2136 RST.n42 RST 0.00104041
R2137 CLK.n9 CLK.t25 36.935
R2138 CLK.n3 CLK.t23 36.935
R2139 CLK.n67 CLK.t19 36.935
R2140 CLK.n61 CLK.t5 36.935
R2141 CLK.n54 CLK.t1 36.935
R2142 CLK.n43 CLK.t14 36.935
R2143 CLK.n37 CLK.t9 36.935
R2144 CLK.n25 CLK.t15 36.935
R2145 CLK.n19 CLK.t11 36.935
R2146 CLK.n14 CLK.t3 25.5364
R2147 CLK.n48 CLK.t17 25.5364
R2148 CLK.n30 CLK.t12 25.5364
R2149 CLK.n72 CLK.t6 25.5361
R2150 CLK.n9 CLK.t24 18.1962
R2151 CLK.n3 CLK.t22 18.1962
R2152 CLK.n67 CLK.t18 18.1962
R2153 CLK.n61 CLK.t4 18.1962
R2154 CLK.n54 CLK.t0 18.1962
R2155 CLK.n43 CLK.t13 18.1962
R2156 CLK.n37 CLK.t7 18.1962
R2157 CLK.n25 CLK.t21 18.1962
R2158 CLK.n19 CLK.t8 18.1962
R2159 CLK.n48 CLK.t2 14.0749
R2160 CLK.n30 CLK.t20 14.0749
R2161 CLK.n14 CLK.t10 14.0749
R2162 CLK.n72 CLK.t16 14.0734
R2163 CLK.n77 CLK 5.77906
R2164 CLK.n79 CLK.n78 5.11659
R2165 CLK.n5 CLK.n2 4.5005
R2166 CLK.n5 CLK.n4 4.5005
R2167 CLK.n8 CLK.n7 4.5005
R2168 CLK.n10 CLK.n7 4.5005
R2169 CLK.n63 CLK.n60 4.5005
R2170 CLK.n63 CLK.n62 4.5005
R2171 CLK.n66 CLK.n65 4.5005
R2172 CLK.n68 CLK.n65 4.5005
R2173 CLK.n75 CLK.n74 4.5005
R2174 CLK.n74 CLK.n73 4.5005
R2175 CLK.n55 CLK.n52 4.5005
R2176 CLK.n39 CLK.n36 4.5005
R2177 CLK.n39 CLK.n38 4.5005
R2178 CLK.n42 CLK.n41 4.5005
R2179 CLK.n44 CLK.n41 4.5005
R2180 CLK.n51 CLK.n50 4.5005
R2181 CLK.n50 CLK.n49 4.5005
R2182 CLK.n21 CLK.n18 4.5005
R2183 CLK.n21 CLK.n20 4.5005
R2184 CLK.n24 CLK.n23 4.5005
R2185 CLK.n26 CLK.n23 4.5005
R2186 CLK.n33 CLK.n32 4.5005
R2187 CLK.n32 CLK.n31 4.5005
R2188 CLK.n79 CLK.n15 4.5005
R2189 CLK.n80 CLK.n79 4.5005
R2190 CLK.n78 CLK 4.43149
R2191 CLK.n81 CLK 4.16645
R2192 CLK.n76 CLK.n57 4.05348
R2193 CLK.n77 CLK.n76 3.5258
R2194 CLK.n76 CLK 2.3355
R2195 CLK.n81 CLK 2.27103
R2196 CLK.n12 CLK.n11 2.25107
R2197 CLK.n70 CLK.n69 2.25107
R2198 CLK.n46 CLK.n45 2.25107
R2199 CLK.n28 CLK.n27 2.25107
R2200 CLK.n53 CLK.n52 2.24763
R2201 CLK.n57 CLK.n56 2.2455
R2202 CLK.n71 CLK.n58 2.24235
R2203 CLK.n47 CLK.n34 2.24235
R2204 CLK.n29 CLK.n16 2.24235
R2205 CLK.n13 CLK.n0 2.24235
R2206 CLK.n55 CLK.n54 2.12246
R2207 CLK.n4 CLK.n3 2.12175
R2208 CLK.n62 CLK.n61 2.12175
R2209 CLK.n38 CLK.n37 2.12175
R2210 CLK.n20 CLK.n19 2.12175
R2211 CLK.n10 CLK.n9 2.12075
R2212 CLK.n68 CLK.n67 2.12075
R2213 CLK.n44 CLK.n43 2.12075
R2214 CLK.n26 CLK.n25 2.12075
R2215 CLK.n7 CLK.n6 1.74297
R2216 CLK.n65 CLK.n64 1.74297
R2217 CLK.n41 CLK.n40 1.74297
R2218 CLK.n23 CLK.n22 1.74297
R2219 CLK.n78 CLK.n77 1.62556
R2220 CLK.n6 CLK.n1 1.49778
R2221 CLK.n64 CLK.n59 1.49778
R2222 CLK.n40 CLK.n35 1.49778
R2223 CLK.n22 CLK.n17 1.49778
R2224 CLK.n73 CLK.n72 1.42775
R2225 CLK.n49 CLK.n48 1.42706
R2226 CLK.n31 CLK.n30 1.42706
R2227 CLK.n15 CLK.n14 1.42706
R2228 CLK.n13 CLK.n12 0.97145
R2229 CLK.n71 CLK.n70 0.97145
R2230 CLK.n47 CLK.n46 0.97145
R2231 CLK.n29 CLK.n28 0.97145
R2232 CLK CLK.n75 0.1605
R2233 CLK CLK.n51 0.1605
R2234 CLK CLK.n33 0.1605
R2235 CLK CLK.n80 0.1605
R2236 CLK.n53 CLK 0.052998
R2237 CLK.n8 CLK 0.0473512
R2238 CLK.n2 CLK 0.0473512
R2239 CLK.n66 CLK 0.0473512
R2240 CLK.n60 CLK 0.0473512
R2241 CLK.n42 CLK 0.0473512
R2242 CLK.n36 CLK 0.0473512
R2243 CLK.n24 CLK 0.0473512
R2244 CLK.n18 CLK 0.0473512
R2245 CLK.n11 CLK.n8 0.0361897
R2246 CLK.n2 CLK.n1 0.0361897
R2247 CLK.n69 CLK.n66 0.0361897
R2248 CLK.n60 CLK.n59 0.0361897
R2249 CLK.n45 CLK.n42 0.0361897
R2250 CLK.n36 CLK.n35 0.0361897
R2251 CLK.n27 CLK.n24 0.0361897
R2252 CLK.n18 CLK.n17 0.0361897
R2253 CLK.n75 CLK.n58 0.03175
R2254 CLK.n51 CLK.n34 0.03175
R2255 CLK.n33 CLK.n16 0.03175
R2256 CLK.n80 CLK.n0 0.03175
R2257 CLK.n74 CLK.n71 0.0246174
R2258 CLK.n50 CLK.n47 0.0246174
R2259 CLK.n32 CLK.n29 0.0246174
R2260 CLK.n79 CLK.n13 0.0246174
R2261 CLK.n56 CLK.n55 0.0210263
R2262 CLK.n56 CLK.n53 0.0183424
R2263 CLK.n6 CLK.n5 0.0131772
R2264 CLK.n64 CLK.n63 0.0131772
R2265 CLK.n40 CLK.n39 0.0131772
R2266 CLK.n22 CLK.n21 0.0131772
R2267 CLK.n57 CLK.n52 0.0128848
R2268 CLK.n12 CLK.n7 0.0122182
R2269 CLK.n70 CLK.n65 0.0122182
R2270 CLK.n46 CLK.n41 0.0122182
R2271 CLK.n28 CLK.n23 0.0122182
R2272 CLK CLK.n81 0.00567241
R2273 CLK.n11 CLK.n10 0.00515517
R2274 CLK.n4 CLK.n1 0.00515517
R2275 CLK.n69 CLK.n68 0.00515517
R2276 CLK.n62 CLK.n59 0.00515517
R2277 CLK.n45 CLK.n44 0.00515517
R2278 CLK.n38 CLK.n35 0.00515517
R2279 CLK.n27 CLK.n26 0.00515517
R2280 CLK.n20 CLK.n17 0.00515517
R2281 CLK.n73 CLK.n58 0.00175
R2282 CLK.n49 CLK.n34 0.00175
R2283 CLK.n31 CLK.n16 0.00175
R2284 CLK.n15 CLK.n0 0.00175
R2285 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n2 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t4 37.1986
R2286 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t8 31.528
R2287 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n0 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t5 30.6344
R2288 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n0 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t7 27.3855
R2289 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n2 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t3 17.6614
R2290 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t6 15.3826
R2291 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n1 7.62751
R2292 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n3 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 6.09789
R2293 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n0 2.8877
R2294 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n3 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 2.67866
R2295 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n3 2.2505
R2296 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n2 1.43709
R2297 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.4325
C0 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 2.92f
C1 a_8126_759# a_8286_759# 0.0504f
C2 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q2 0.109f
C3 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0622f
C4 a_7562_759# CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.46e-19
C5 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK 0.00104f
C6 a_4875_1632# CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.00695f
C7 CLK_div_10_mag_0.nor_3_mag_0.IN3 VDD 0.396f
C8 CLK CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 6.86e-20
C9 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 3.97e-19
C10 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 4.69e-20
C11 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 2.19f
C12 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 5.73e-20
C13 CLK CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 1.52e-20
C14 CLK_div_10_mag_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 2.44e-20
C15 a_8149_1634# CLK_DIV_11_mag_new_0.Q1 0.0101f
C16 a_3226_n338# VDD 3.56e-19
C17 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 2.04e-19
C18 RST CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0316f
C19 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.QB 0.25f
C20 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 7.55e-19
C21 a_1176_1634# CLK_DIV_11_mag_new_0.Q3 0.0152f
C22 a_1016_1634# a_1176_1634# 0.0504f
C23 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C24 CLK_div_10_mag_0.and2_mag_0.OUT a_12318_n2129# 0.0294f
C25 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C26 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.Q1 8.51e-22
C27 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 2.6e-20
C28 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.161f
C29 a_7562_759# CLK_div_10_mag_0.Q1 0.00166f
C30 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK 0.779f
C31 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_12277_n338# 0.00118f
C32 CLK_div_10_mag_0.JK_FF_mag_2.K a_12277_n338# 0.0114f
C33 RST a_1368_759# 0.00334f
C34 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C35 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.012f
C36 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.013f
C37 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_12282_2771# 0.00118f
C38 a_5035_1632# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0733f
C39 a_6243_n338# CLK_div_10_mag_0.Q1 0.069f
C40 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0833f
C41 CLK_DIV_11_mag_new_0.Q3 CLK 0.48f
C42 CLK_DIV_11_mag_new_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 1.93e-20
C43 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 1.1e-19
C44 VDD a_12282_2771# 3.56e-19
C45 a_4385_759# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 1.17e-20
C46 CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.111f
C47 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00975f
C48 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN VDD 0.512f
C49 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_6243_n338# 0.00118f
C50 a_1016_1634# CLK 0.00224f
C51 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 VDD 9.71f
C52 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.321f
C53 CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK 0.0765f
C54 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 0.647f
C55 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.Q1 3.09e-19
C56 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD 0.391f
C57 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 6.32e-22
C58 a_8132_n338# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0697f
C59 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q1 2.57f
C60 a_8286_759# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 3.66e-20
C61 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 0.00101f
C62 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00183f
C63 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 8.26e-20
C64 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q0 0.00525f
C65 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 7.08e-20
C66 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.198f
C67 a_2252_759# CLK_div_10_mag_0.JK_FF_mag_1.QB 0.00696f
C68 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.0116f
C69 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.109f
C70 a_7989_1634# VDD 2.21e-19
C71 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.Q3 0.133f
C72 a_1016_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 8.64e-19
C73 a_7425_1634# CLK_DIV_11_mag_new_0.Q2 4.66e-19
C74 a_2662_n338# VDD 3.14e-19
C75 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN a_n796_2646# 1.14e-19
C76 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 1.88e-19
C77 a_7989_1634# CLK_DIV_11_mag_new_0.Q1 0.0102f
C78 a_1016_1634# CLK_DIV_11_mag_new_0.Q3 0.0124f
C79 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.119f
C80 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT RST 0.268f
C81 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.529f
C82 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.K 0.783f
C83 CLK_div_10_mag_0.JK_FF_mag_2.K a_11713_n338# 2.96e-19
C84 CLK_div_10_mag_0.Q0 a_11149_n338# 6.43e-21
C85 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.Q3 3.89e-20
C86 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_11718_2771# 0.011f
C87 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_11713_n338# 0.011f
C88 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 8.76e-20
C89 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 1.32e-19
C90 a_5679_n338# CLK_div_10_mag_0.Q1 6.06e-21
C91 a_4875_1632# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0203f
C92 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00393f
C93 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_5679_n338# 0.011f
C94 VDD CLK_div_10_mag_0.Q3 1.18f
C95 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN Vdiv110 1.82e-19
C96 VDD a_11718_2771# 3.14e-19
C97 Vdiv110 a_12478_n2129# 0.198f
C98 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.Q2 0.888f
C99 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_1.QB 0.198f
C100 a_8126_759# VDD 0.00123f
C101 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.01f
C102 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00158f
C103 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 1.89e-20
C104 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.36f
C105 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_1.QB 0.307f
C106 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.Q0 0.0709f
C107 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 0.342f
C108 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q0 8.33e-20
C109 a_2464_1678# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0036f
C110 RST CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.192f
C111 a_9123_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00372f
C112 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK 1.48e-20
C113 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT RST 0.268f
C114 CLK a_1368_759# 4.62e-19
C115 CLK_div_10_mag_0.JK_FF_mag_0.K VDD 0.496f
C116 CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00264f
C117 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 6.82e-19
C118 a_7265_1634# CLK_DIV_11_mag_new_0.Q2 6.02e-19
C119 a_7425_1634# CLK_DIV_11_mag_new_0.Q1 0.00789f
C120 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.343f
C121 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C122 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 5.45e-20
C123 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 8.16e-20
C124 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q0 0.0399f
C125 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.K 0.283f
C126 CLK_DIV_11_mag_new_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 2.15e-20
C127 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.768f
C128 a_1528_759# VDD 0.00892f
C129 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C130 CLK_DIV_11_mag_new_0.Q0 VDD 3.77f
C131 CLK_div_10_mag_0.JK_FF_mag_2.K a_11149_n338# 3.25e-19
C132 a_4311_1632# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 1.5e-20
C133 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_11154_2771# 1.43e-19
C134 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_11149_n338# 1.43e-19
C135 a_2092_759# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 9.1e-19
C136 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 6.04e-21
C137 a_4317_2729# CLK_div_10_mag_0.CLK 1.88e-19
C138 CLK_div_10_mag_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 1.37e-20
C139 VDD a_11154_2771# 3.14e-19
C140 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_5115_n338# 1.43e-19
C141 Vdiv110 a_12318_n2129# 0.0132f
C142 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.Q1 3.23f
C143 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 2.54e-20
C144 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.and2_mag_0.OUT 0.125f
C145 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.651f
C146 a_9282_n1435# CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.069f
C147 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K RST 0.0872f
C148 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 3.61e-20
C149 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 6.82e-19
C150 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 RST 0.0717f
C151 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 9.94e-21
C152 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00403f
C153 a_9123_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 4.52e-20
C154 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 2.81e-20
C155 CLK CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 3.15e-20
C156 a_7265_1634# VDD 2.76e-19
C157 a_8559_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.069f
C158 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 2.03e-20
C159 a_7265_1634# CLK_DIV_11_mag_new_0.Q1 0.00335f
C160 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 2.33e-19
C161 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_2.K 0.00586f
C162 a_6163_1676# CLK_DIV_11_mag_new_0.Q2 0.0157f
C163 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_8696_n338# 4.52e-20
C164 CLK_div_10_mag_0.JK_FF_mag_3.QB a_7568_n338# 0.00392f
C165 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00157f
C166 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_2662_n338# 4.52e-20
C167 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.00253f
C168 a_12431_759# CLK_div_10_mag_0.JK_FF_mag_2.K 0.0811f
C169 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00183f
C170 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 1.08f
C171 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.36f
C172 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_10590_2727# 0.00119f
C173 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 5.53e-20
C174 a_4151_1632# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 1.17e-20
C175 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 5.52e-20
C176 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C177 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 4.67e-22
C178 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 2.47e-20
C179 a_4157_2729# CLK_div_10_mag_0.CLK 2.69e-19
C180 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD 0.442f
C181 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.769f
C182 RST CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0697f
C183 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK 3.86e-20
C184 a_9282_n1435# CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 1.29e-22
C185 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_2.K 0.00586f
C186 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0377f
C187 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 6.57e-19
C188 a_5109_759# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0203f
C189 CLK_div_10_mag_0.JK_FF_mag_2.QB a_7568_n338# 1.41e-20
C190 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 1.77e-19
C191 a_4881_2773# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00378f
C192 a_7402_759# CLK_div_10_mag_0.Q2 0.00335f
C193 a_6163_1676# VDD 3.14e-19
C194 CLK_div_10_mag_0.CLK a_2098_n338# 6.43e-21
C195 CLK_DIV_11_mag_new_0.Q3 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 2.61e-20
C196 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.122f
C197 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.00252f
C198 a_5599_1676# CLK_DIV_11_mag_new_0.Q2 0.00859f
C199 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 9.58e-19
C200 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_8132_n338# 0.0202f
C201 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK 0.579f
C202 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_12478_n2129# 5.39e-20
C203 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 1.5e-20
C204 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_2.K 2.02e-20
C205 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C206 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q3 0.329f
C207 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD 0.994f
C208 a_11867_759# CLK_div_10_mag_0.JK_FF_mag_2.K 0.00964f
C209 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_11867_759# 0.0036f
C210 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.28f
C211 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.289f
C212 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 1.94e-20
C213 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB VDD 0.904f
C214 a_10250_n1435# VDD 3.14e-19
C215 VDD a_10430_2727# 2.21e-19
C216 a_2092_759# a_2252_759# 0.0504f
C217 a_1528_759# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1.5e-20
C218 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.Q1 1.76e-21
C219 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 4.36e-19
C220 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0106f
C221 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT RST 3.84e-20
C222 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 2.48e-19
C223 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.00388f
C224 a_2816_759# RST 0.0015f
C225 CLK_DIV_11_mag_new_0.Q2 CLK_div_10_mag_0.Q1 9.64e-20
C226 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 2.12e-19
C227 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.Q3 0.076f
C228 CLK_DIV_11_mag_new_0.Q2 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 7.49e-20
C229 CLK_div_10_mag_0.JK_FF_mag_2.QB a_7408_n338# 1.86e-20
C230 a_1176_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 8.66e-20
C231 a_5445_2773# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0059f
C232 CLK_DIV_11_mag_new_0.Q3 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 3.07e-20
C233 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 0.209f
C234 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 1.36e-19
C235 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.00243f
C236 a_4317_2729# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0732f
C237 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 VDD 1.08f
C238 a_5599_1676# VDD 3.14e-19
C239 a_5035_1632# CLK_DIV_11_mag_new_0.Q2 0.0101f
C240 CLK_DIV_11_mag_new_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 9e-20
C241 a_12318_n2129# a_12478_n2129# 0.186f
C242 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_12318_n2129# 9.16e-20
C243 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.519f
C244 a_7431_2731# CLK 0.0105f
C245 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.338f
C246 a_2874_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00372f
C247 a_11303_759# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 8.64e-19
C248 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 VDD 0.514f
C249 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.0432f
C250 a_10584_1630# CLK_div_10_mag_0.Q0 7.56e-21
C251 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 1.29e-19
C252 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00156f
C253 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 6.18e-19
C254 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_DIV_11_mag_new_0.Q1 4.07e-19
C255 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.768f
C256 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK 1.48e-19
C257 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 2.92e-20
C258 a_11308_1630# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 2.88e-20
C259 VDD a_9123_2775# 3.56e-19
C260 CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_10_mag_0.Q2 3.87e-19
C261 VDD CLK_div_10_mag_0.Q1 4.14f
C262 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 VDD 1.03f
C263 a_n358_4884# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 2.69e-22
C264 RST CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.295f
C265 CLK_DIV_11_mag_new_0.Q1 a_9123_2775# 0.069f
C266 CLK_DIV_11_mag_new_0.Q1 CLK_div_10_mag_0.Q1 9.86e-19
C267 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0502f
C268 a_2252_759# VDD 0.00101f
C269 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.122f
C270 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.Q2 0.253f
C271 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0281f
C272 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C273 a_4881_2773# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0697f
C274 CLK_div_10_mag_0.JK_FF_mag_2.QB a_6243_n338# 0.0114f
C275 a_4157_2729# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0203f
C276 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.0275f
C277 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.00117f
C278 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.16f
C279 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 1.4e-20
C280 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VDD 0.994f
C281 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 2.11e-20
C282 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK 5.45e-20
C283 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_2.QB 2.59e-21
C284 a_4875_1632# CLK_DIV_11_mag_new_0.Q2 0.0102f
C285 a_11308_1630# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 8.64e-19
C286 a_7271_2731# CLK 0.0114f
C287 a_2310_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.069f
C288 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.and2_mag_1.OUT 0.0693f
C289 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 a_6243_n338# 0.00372f
C290 a_11143_759# VDD 2.21e-19
C291 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_10_mag_0.Q2 1.23e-19
C292 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_1114_4881# 8.64e-19
C293 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD 0.395f
C294 CLK_div_10_mag_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 2.84e-20
C295 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 2.25e-21
C296 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.298f
C297 a_11148_1630# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 9.1e-19
C298 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 6.62e-20
C299 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.CLK 1.86e-19
C300 VDD a_8559_2775# 3.14e-19
C301 CLK_div_10_mag_0.CLK VDD 4f
C302 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 7e-19
C303 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.161f
C304 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0998f
C305 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 1.48e-19
C306 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 1.34e-19
C307 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 3.43e-19
C308 CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 9.8e-19
C309 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.Q1 0.25f
C310 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00115f
C311 CLK_div_10_mag_0.JK_FF_mag_2.QB a_5679_n338# 2.96e-19
C312 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.321f
C313 a_8850_759# VDD 0.00152f
C314 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 7.24e-19
C315 a_4875_1632# VDD 2.21e-19
C316 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C317 a_1114_4881# CLK 1.64e-20
C318 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.221f
C319 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 6.35e-19
C320 a_4311_1632# CLK_DIV_11_mag_new_0.Q2 0.00789f
C321 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_10_mag_0.Q1 7.89e-20
C322 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.484f
C323 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT VDD 0.569f
C324 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.Q3 9.83e-19
C325 a_6009_2773# CLK 9.33e-19
C326 RST CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.286f
C327 a_10579_759# VDD 0.00299f
C328 a_8126_759# CLK_div_10_mag_0.Q2 0.0102f
C329 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 a_5679_n338# 0.069f
C330 a_11148_1630# a_11308_1630# 0.0504f
C331 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.397f
C332 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_DIV_11_mag_new_0.Q1 3.09e-19
C333 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 1.32e-19
C334 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.1f
C335 CLK_div_10_mag_0.Q0 a_4551_n338# 0.00939f
C336 VDD a_7995_2775# 3.14e-19
C337 a_10584_1630# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0731f
C338 CLK_div_10_mag_0.and2_mag_1.OUT RST 4.25e-20
C339 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_8132_n338# 0.00378f
C340 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 6.91e-20
C341 a_5035_1632# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 2.88e-20
C342 a_7562_759# RST 0.00247f
C343 a_5833_759# VDD 0.00152f
C344 a_9506_4996# VDD 0.0418f
C345 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00178f
C346 CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_10_mag_0.Q2 0.289f
C347 a_8713_1678# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0036f
C348 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_DIV_11_mag_new_0.Q2 0.127f
C349 a_4881_2773# RST 3.08e-20
C350 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.233f
C351 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 9.05e-22
C352 CLK_div_10_mag_0.JK_FF_mag_2.QB a_5115_n338# 3.25e-19
C353 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 3.22e-20
C354 CLK_div_10_mag_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00115f
C355 a_2252_759# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0733f
C356 CLK_div_10_mag_0.Q0 a_1534_n338# 2.79e-20
C357 a_4311_1632# VDD 1.04e-19
C358 CLK_div_10_mag_0.JK_FF_mag_1.QB RST 0.253f
C359 CLK_div_10_mag_0.Q0 a_3380_759# 0.0157f
C360 CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_DIV_11_mag_new_0.Q3 0.0145f
C361 a_4151_1632# CLK_DIV_11_mag_new_0.Q2 0.00335f
C362 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 a_n796_2646# 0.0178f
C363 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 9.75e-19
C364 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00262f
C365 a_5445_2773# CLK 9.25e-19
C366 CLK_div_10_mag_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 2.89e-20
C367 CLK_div_10_mag_0.nor_3_mag_0.IN3 a_12277_n338# 2.1e-20
C368 a_10419_759# VDD 0.00727f
C369 a_4151_1632# CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 8.64e-19
C370 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0951f
C371 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 5.7e-20
C372 a_8286_759# CLK_div_10_mag_0.JK_FF_mag_3.QB 0.00696f
C373 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.Q0 1.76f
C374 CLK_div_10_mag_0.JK_FF_mag_2.K a_4551_n338# 9.32e-19
C375 CLK_div_10_mag_0.Q0 a_4391_n338# 0.0101f
C376 a_10424_1630# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0202f
C377 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 VDD 0.69f
C378 a_4875_1632# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 9.1e-19
C379 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C380 a_9346_4996# VDD 0.235f
C381 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00154f
C382 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_DIV_11_mag_new_0.Q1 0.00103f
C383 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 2.98e-19
C384 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 9.12e-19
C385 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0834f
C386 a_4151_1632# VDD 2.21e-19
C387 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0129f
C388 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 0.648f
C389 a_7265_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 8.64e-19
C390 a_9277_1678# CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 4.81e-20
C391 a_6609_4975# CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 0.069f
C392 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 1.17e-19
C393 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0622f
C394 RST CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 1.36e-19
C395 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 7.32e-20
C396 a_4881_2773# CLK 3.81e-19
C397 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q2 0.305f
C398 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.338f
C399 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.306f
C400 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00118f
C401 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0899f
C402 a_3028_1678# CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 1.44e-21
C403 CLK_div_10_mag_0.Q0 a_3226_n338# 0.069f
C404 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 0.342f
C405 a_4317_2729# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 1.24e-20
C406 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00544f
C407 CLK_div_10_mag_0.JK_FF_mag_2.K a_4391_n338# 0.00876f
C408 CLK CLK_div_10_mag_0.JK_FF_mag_1.QB 1.61e-19
C409 a_6609_4975# VDD 3.14e-19
C410 a_4311_1632# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0731f
C411 a_5035_1632# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 1.04e-19
C412 a_5115_n338# RST 1.23e-20
C413 a_6397_759# CLK_div_10_mag_0.Q1 0.0157f
C414 a_6609_4975# CLK_DIV_11_mag_new_0.Q1 0.015f
C415 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 1.84e-21
C416 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 7.07e-19
C417 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q0 0.305f
C418 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0151f
C419 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q2 0.00675f
C420 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.Q2 2.45e-22
C421 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0432f
C422 a_12277_n338# CLK_div_10_mag_0.Q3 0.069f
C423 a_3028_1678# VDD 3.14e-19
C424 a_5904_4934# CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 4.43e-21
C425 CLK_DIV_11_mag_new_0.Q2 CLK_div_10_mag_0.JK_FF_mag_2.QB 3.98e-20
C426 CLK_DIV_11_mag_new_0.Q3 CLK_div_10_mag_0.JK_FF_mag_1.QB 7.16e-20
C427 RST CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0298f
C428 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00391f
C429 a_2098_n338# RST 2.66e-19
C430 a_10250_n1435# CLK_div_10_mag_0.Q2 0.0096f
C431 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 0.275f
C432 a_4317_2729# CLK 0.0105f
C433 CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 4.39e-19
C434 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 2.59e-19
C435 CLK_div_10_mag_0.JK_FF_mag_3.QB VDD 0.913f
C436 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 2.56e-19
C437 a_2464_1678# CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 4.96e-22
C438 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.132f
C439 CLK_DIV_11_mag_new_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.QB 2.31e-19
C440 CLK_DIV_11_mag_new_0.Q2 a_4385_759# 1.04e-19
C441 CLK_div_10_mag_0.Q0 a_2662_n338# 6.06e-21
C442 a_4157_2729# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 1.59e-20
C443 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C444 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_2816_759# 0.0036f
C445 a_4151_1632# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0202f
C446 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00183f
C447 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 3.83e-19
C448 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C449 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD 0.648f
C450 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK 5.92e-19
C451 a_7425_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 1.46e-19
C452 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.Q2 0.0209f
C453 a_5269_759# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 8.64e-19
C454 a_5904_4934# CLK_DIV_11_mag_new_0.Q1 5.19e-20
C455 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0934f
C456 a_n1595_3762# CLK_DIV_11_mag_new_0.Q0 0.0177f
C457 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VDD 0.497f
C458 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00637f
C459 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 1.35e-20
C460 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00107f
C461 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 2.67e-20
C462 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.Q3 0.149f
C463 a_8286_759# RST 0.00211f
C464 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q1 7.47e-19
C465 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 RST 2.96e-19
C466 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 4.01e-20
C467 CLK_div_10_mag_0.JK_FF_mag_2.QB VDD 0.914f
C468 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.651f
C469 a_2464_1678# VDD 3.14e-19
C470 a_5744_4934# CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 3.44e-21
C471 a_n1762_4447# CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 0.069f
C472 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 a_12436_1674# 0.00372f
C473 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_2.K 4.2e-20
C474 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 7.04e-20
C475 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 1.17e-19
C476 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0143f
C477 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.359f
C478 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 3.41e-19
C479 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.11f
C480 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.Q2 0.98f
C481 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_DIV_11_mag_new_0.Q3 0.00935f
C482 a_4157_2729# CLK 0.0114f
C483 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 1.76e-20
C484 a_4385_759# VDD 0.0123f
C485 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00975f
C486 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.233f
C487 a_10424_1630# a_10584_1630# 0.0504f
C488 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 2.03e-20
C489 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 7.97e-19
C490 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD 0.398f
C491 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.K 0.487f
C492 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 3.18e-19
C493 a_2874_2775# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.0114f
C494 CLK_div_10_mag_0.and2_mag_0.OUT VDD 1.03f
C495 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 6.69e-19
C496 a_7271_2731# a_7431_2731# 0.0504f
C497 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 4.26e-19
C498 a_5744_4934# VDD 5.08e-19
C499 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.01f
C500 a_2092_759# RST 0.00283f
C501 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 1.74e-19
C502 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN a_1182_2731# 1.03e-20
C503 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_10_mag_0.Q1 5.37e-19
C504 a_5744_4934# CLK_DIV_11_mag_new_0.Q1 3.35e-20
C505 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.642f
C506 a_n1755_3762# CLK_DIV_11_mag_new_0.Q0 0.00765f
C507 CLK_div_10_mag_0.Q0 a_1528_759# 0.00789f
C508 a_n796_2646# VDD 0.173f
C509 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD 0.398f
C510 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.Q3 2f
C511 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.338f
C512 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.Q3 0.0263f
C513 Vdiv110 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 3.1e-22
C514 a_8286_759# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 8.64e-19
C515 a_11143_759# CLK_div_10_mag_0.Q2 3.6e-22
C516 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 0.00296f
C517 a_n358_4884# CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 0.132f
C518 CLK_DIV_11_mag_new_0.Q2 RST 0.166f
C519 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_0.K 0.125f
C520 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 1.2e-19
C521 a_7562_759# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 1.5e-20
C522 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 a_11872_1674# 0.069f
C523 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 1.47e-20
C524 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.122f
C525 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K RST 0.0775f
C526 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.Q2 3.3e-19
C527 a_2874_2775# CLK 9.34e-19
C528 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_0.K 0.0156f
C529 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_0.K 0.0836f
C530 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 3.79e-19
C531 a_2310_2775# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 2.96e-19
C532 a_7431_2731# CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 1.16e-20
C533 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 1.19e-19
C534 a_n1762_4447# VDD 3.14e-19
C535 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00156f
C536 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q0 0.00123f
C537 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 4.42e-19
C538 a_10425_n338# VDD 2.21e-19
C539 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.0262f
C540 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN a_1114_4881# 2.4e-20
C541 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN a_1022_2731# 1.29e-20
C542 a_8850_759# CLK_div_10_mag_0.Q2 0.00859f
C543 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 RST 0.00535f
C544 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.Q2 0.0661f
C545 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 3.21e-20
C546 a_n1762_4447# CLK_DIV_11_mag_new_0.Q1 0.00544f
C547 RST CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.152f
C548 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT a_11154_2771# 0.00378f
C549 a_12436_1674# CLK_DIV_11_mag_new_0.Q0 0.0157f
C550 CLK_DIV_11_mag_new_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.K 8.75e-20
C551 VDD RST 2.38f
C552 CLK_DIV_11_mag_new_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 3.71e-20
C553 a_2874_2775# CLK_DIV_11_mag_new_0.Q3 0.069f
C554 a_12431_759# CLK_div_10_mag_0.Q3 0.0157f
C555 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0979f
C556 CLK_DIV_11_mag_new_0.Q1 RST 0.163f
C557 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.412f
C558 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C559 a_1740_1634# VDD 2.21e-19
C560 a_10579_759# CLK_div_10_mag_0.Q2 1.86e-20
C561 a_8314_n1435# CLK_div_10_mag_0.Q1 0.0105f
C562 CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 0.205f
C563 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0384f
C564 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 9.58e-20
C565 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_10_mag_0.Q3 4.22e-20
C566 a_1114_4881# CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.132f
C567 a_2310_2775# CLK 9.23e-19
C568 a_4545_759# CLK_div_10_mag_0.Q1 0.00789f
C569 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 2.01e-19
C570 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 0.299f
C571 a_1746_2775# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 3.33e-19
C572 a_4545_759# CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.46e-19
C573 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.101f
C574 CLK CLK_DIV_11_mag_new_0.Q2 1.48f
C575 a_7271_2731# CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 1.49e-20
C576 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 2.86e-19
C577 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VDD 1.32f
C578 a_7568_n338# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0732f
C579 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K a_7995_2775# 1.39e-19
C580 a_4551_n338# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0732f
C581 a_9260_n338# VDD 3.56e-19
C582 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 9.9e-19
C583 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.129f
C584 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.Q1 0.0161f
C585 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 9.45e-20
C586 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 1.05e-20
C587 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_0.Q3 1.89e-20
C588 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 a_11718_2771# 0.00605f
C589 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_11713_n338# 4.52e-20
C590 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK 0.631f
C591 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK 5.73e-19
C592 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT a_10590_2727# 0.0732f
C593 a_9414_759# CLK_div_10_mag_0.JK_FF_mag_3.QB 0.0811f
C594 a_11872_1674# CLK_DIV_11_mag_new_0.Q0 0.00859f
C595 Vdiv110 VDD 0.0768f
C596 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_5679_n338# 4.52e-20
C597 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_DIV_11_mag_new_0.Q0 6.99e-20
C598 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.653f
C599 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_1.QB 0.28f
C600 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_2.K 9.73e-19
C601 a_11867_759# CLK_div_10_mag_0.Q3 0.00859f
C602 CLK_div_10_mag_0.Q0 a_10250_n1435# 0.01f
C603 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00213f
C604 a_n350_4053# CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.069f
C605 a_10419_759# CLK_div_10_mag_0.Q2 2.55e-20
C606 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.338f
C607 CLK_DIV_11_mag_new_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 1.84e-20
C608 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.Q2 0.0579f
C609 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C610 CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 a_n358_4884# 0.0202f
C611 a_2874_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C612 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C613 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.Q2 1.19f
C614 CLK_DIV_11_mag_new_0.and2_mag_3.OUT VDD 0.303f
C615 CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q2 0.00392f
C616 a_1746_2775# CLK 3.8e-19
C617 a_9123_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00118f
C618 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 3.43e-19
C619 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK 0.416f
C620 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD 0.52f
C621 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.Q1 0.209f
C622 CLK VDD 5.66f
C623 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.Q3 0.0703f
C624 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 9.5e-19
C625 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.857f
C626 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.126f
C627 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 4.78e-20
C628 RST CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0915f
C629 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.Q1 7.38e-19
C630 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00157f
C631 CLK CLK_DIV_11_mag_new_0.Q1 0.554f
C632 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.294f
C633 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.792f
C634 a_1182_2731# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.00392f
C635 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 8.64e-20
C636 a_6009_2773# CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.0114f
C637 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_10250_n1435# 5.1e-20
C638 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.321f
C639 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 1.06e-19
C640 a_7408_n338# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0203f
C641 a_4391_n338# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0203f
C642 a_1534_n338# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0732f
C643 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.Q0 0.00425f
C644 a_5109_759# VDD 0.00123f
C645 a_8696_n338# VDD 3.14e-19
C646 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.K 0.251f
C647 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.103f
C648 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 0.342f
C649 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C650 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 a_11154_2771# 0.0697f
C651 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_11149_n338# 0.0202f
C652 a_11308_1630# CLK_DIV_11_mag_new_0.Q0 0.0101f
C653 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT a_10430_2727# 0.0203f
C654 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_5115_n338# 0.0202f
C655 a_12436_1674# CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 0.0811f
C656 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K VDD 0.623f
C657 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 7.16e-20
C658 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.46e-20
C659 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.995f
C660 CLK_DIV_11_mag_new_0.Q3 VDD 4.33f
C661 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.Q1 1.16f
C662 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.Q1 9.69e-19
C663 a_1016_1634# VDD 2.21e-19
C664 a_4385_759# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0202f
C665 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.3f
C666 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 1.83e-19
C667 CLK_DIV_11_mag_new_0.and2_mag_3.IN1 VDD 0.795f
C668 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 2e-19
C669 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT RST 0.288f
C670 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0346f
C671 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.Q1 1.83f
C672 CLK_div_10_mag_0.Q0 a_2252_759# 0.0101f
C673 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.122f
C674 a_6397_759# CLK_div_10_mag_0.JK_FF_mag_2.QB 0.0811f
C675 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 7.36e-21
C676 a_1900_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 8.64e-19
C677 CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q1 0.106f
C678 a_8559_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.011f
C679 a_1182_2731# CLK 0.0105f
C680 a_2098_n338# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0697f
C681 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 1.85e-19
C682 a_5904_4934# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 4.33e-21
C683 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.K 0.0501f
C684 a_8286_759# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0733f
C685 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 2.39e-21
C686 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C687 a_7408_n338# a_7568_n338# 0.0504f
C688 a_5445_2773# CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 2.96e-19
C689 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q1 0.303f
C690 a_8132_n338# VDD 3.14e-19
C691 a_1374_n338# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0203f
C692 a_4391_n338# a_4551_n338# 0.0504f
C693 a_11303_759# CLK_div_10_mag_0.JK_FF_mag_2.K 0.00696f
C694 a_6609_4975# CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 2.5e-19
C695 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C696 a_8850_759# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 5.02e-20
C697 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0635f
C698 a_11148_1630# CLK_DIV_11_mag_new_0.Q0 0.0102f
C699 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 6.91e-20
C700 a_1182_2731# CLK_DIV_11_mag_new_0.Q3 3.43e-19
C701 a_2816_759# CLK_div_10_mag_0.JK_FF_mag_1.QB 0.00964f
C702 a_11872_1674# CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 0.00964f
C703 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 1.32e-21
C704 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.CLK 0.158f
C705 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.Q1 0.0871f
C706 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.26f
C707 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.Q2 1.96f
C708 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 0.139f
C709 RST CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.188f
C710 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.K 0.0905f
C711 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.103f
C712 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_2098_n338# 1.43e-19
C713 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C714 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.25f
C715 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 7.17e-19
C716 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.321f
C717 a_1022_2731# CLK 0.0114f
C718 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.Q0 0.242f
C719 a_7402_759# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0202f
C720 a_9414_759# RST 0.00122f
C721 a_7995_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 1.43e-19
C722 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.36f
C723 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.Q2 8.27e-19
C724 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.00126f
C725 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 2.76e-19
C726 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0622f
C727 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD 0.397f
C728 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0591f
C729 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 1.29e-19
C730 VDD a_1368_759# 0.0132f
C731 a_12478_n2129# VDD 0.0407f
C732 RST CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0792f
C733 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD 0.517f
C734 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 3.57e-20
C735 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.K 2.44e-20
C736 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 3.6e-21
C737 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.43e-20
C738 a_4881_2773# CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 3.12e-19
C739 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 3.26e-20
C740 CLK CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 9.92e-20
C741 a_1374_n338# a_1534_n338# 0.0504f
C742 a_9282_n1435# CLK_div_10_mag_0.Q1 0.0084f
C743 CLK_div_10_mag_0.Q0 a_10579_759# 0.00164f
C744 a_5269_759# CLK_div_10_mag_0.Q1 0.0101f
C745 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0404f
C746 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_11867_759# 0.00378f
C747 a_11143_759# CLK_div_10_mag_0.JK_FF_mag_2.K 0.00695f
C748 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 0.0121f
C749 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_2.K 1.54e-19
C750 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0379f
C751 a_10584_1630# CLK_DIV_11_mag_new_0.Q0 0.00789f
C752 a_1022_2731# CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 0.00472f
C753 a_1022_2731# CLK_DIV_11_mag_new_0.Q3 4.47e-19
C754 a_11308_1630# CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 0.00696f
C755 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_0.CLK 2.18e-21
C756 a_6397_759# RST 0.00122f
C757 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_2.K 0.002f
C758 a_9277_1678# CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.0811f
C759 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00254f
C760 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 2.57e-19
C761 CLK_DIV_11_mag_new_0.Q2 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 5.98e-20
C762 a_5445_2773# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 4.52e-20
C763 CLK_DIV_11_mag_new_0.Q3 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 8.64e-20
C764 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.Q2 0.179f
C765 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD 1f
C766 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q2 0.0609f
C767 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_10_mag_0.Q1 0.0635f
C768 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_10_mag_0.Q2 4.88e-19
C769 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.321f
C770 a_11872_1674# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.00378f
C771 a_12318_n2129# VDD 0.234f
C772 CLK_DIV_11_mag_new_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 4.93e-20
C773 a_4317_2729# CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.00392f
C774 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0844f
C775 a_2874_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C776 RST CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 1.38e-19
C777 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0231f
C778 CLK_div_10_mag_0.Q0 a_10419_759# 0.00117f
C779 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.121f
C780 a_10579_759# CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.46e-19
C781 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 2.48e-19
C782 a_10424_1630# CLK_DIV_11_mag_new_0.Q0 0.00335f
C783 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.105f
C784 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.Q2 4.54f
C785 a_11148_1630# CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 0.00695f
C786 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.653f
C787 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD 1f
C788 a_8713_1678# CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.00964f
C789 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_div_10_mag_0.CLK 0.123f
C790 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.00238f
C791 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 4.11e-19
C792 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q0 0.107f
C793 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_8850_759# 0.069f
C794 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VDD 0.434f
C795 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00397f
C796 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00265f
C797 a_4881_2773# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0195f
C798 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q1 0.116f
C799 a_10425_n338# CLK_div_10_mag_0.Q2 6.36e-19
C800 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 1.65e-21
C801 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 5.2e-20
C802 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 6.36e-20
C803 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.777f
C804 a_5109_759# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 9.1e-19
C805 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 2.48e-19
C806 a_11308_1630# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0733f
C807 RST CLK_div_10_mag_0.Q2 0.11f
C808 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 3.8e-20
C809 a_2310_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.011f
C810 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.0715f
C811 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K VDD 0.829f
C812 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_1368_759# 1.17e-20
C813 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VDD 1.24f
C814 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.Q1 3.7f
C815 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00952f
C816 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_0.CLK 6.94e-19
C817 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K RST 0.0789f
C818 a_7989_1634# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 5.49e-20
C819 a_8149_1634# CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.00696f
C820 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 RST 9.24e-20
C821 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 3.54e-20
C822 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT a_9506_4996# 0.198f
C823 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0135f
C824 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q2 0.0766f
C825 a_n350_4053# CLK_DIV_11_mag_new_0.Q0 0.00379f
C826 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 3.32e-20
C827 a_4385_759# a_4545_759# 0.0504f
C828 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00639f
C829 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 1.03e-19
C830 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN a_n358_4884# 2.7e-20
C831 a_9260_n338# CLK_div_10_mag_0.Q2 0.069f
C832 a_7989_1634# a_8149_1634# 0.0504f
C833 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_5833_759# 0.069f
C834 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0187f
C835 a_11148_1630# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0203f
C836 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00545f
C837 a_1746_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 1.43e-19
C838 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 1.2e-19
C839 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C840 a_8126_759# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 9.1e-19
C841 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 1.93f
C842 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 0.343f
C843 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 1.15f
C844 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 a_12282_2771# 4.52e-20
C845 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q2 0.0515f
C846 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_3.QB 0.0615f
C847 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00367f
C848 CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_10_mag_0.Q3 0.00442f
C849 a_7431_2731# CLK_DIV_11_mag_new_0.Q1 2.79e-20
C850 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_9260_n338# 0.00372f
C851 a_6163_1676# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.00372f
C852 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VDD 0.408f
C853 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD 0.457f
C854 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 2.04e-19
C855 CLK_div_10_mag_0.and2_mag_0.OUT a_12277_n338# 1.54e-19
C856 a_7989_1634# CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.00695f
C857 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.109f
C858 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.27f
C859 CLK CLK_div_10_mag_0.Q2 8.66e-20
C860 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT a_9346_4996# 0.0135f
C861 a_n358_4884# CLK_DIV_11_mag_new_0.Q2 0.00186f
C862 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q1 0.0365f
C863 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.768f
C864 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.98e-19
C865 CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 0.124f
C866 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.QB 0.348f
C867 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 4.04e-19
C868 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_3.QB 1e-19
C869 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK 0.925f
C870 a_10584_1630# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 1.5e-20
C871 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 9.96e-20
C872 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00118f
C873 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VDD 0.409f
C874 a_1182_2731# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00119f
C875 a_4545_759# RST 0.00247f
C876 CLK_div_10_mag_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 8.64e-20
C877 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD 0.741f
C878 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_10_mag_0.Q3 2.27e-20
C879 a_7271_2731# VDD 2.21e-19
C880 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q1 0.0248f
C881 a_1114_4881# CLK_DIV_11_mag_new_0.Q2 0.0115f
C882 a_2816_759# VDD 0.00152f
C883 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_2.K 0.0835f
C884 CLK_div_10_mag_0.Q0 a_4385_759# 0.001f
C885 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 7.08e-20
C886 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0205f
C887 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 1.97f
C888 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_8696_n338# 0.069f
C889 a_6009_2773# CLK_DIV_11_mag_new_0.Q2 0.069f
C890 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 2.21e-19
C891 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.and2_mag_0.OUT 0.026f
C892 a_n358_4884# VDD 0.165f
C893 a_5599_1676# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.069f
C894 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.16f
C895 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.0683f
C896 a_10584_1630# CLK_div_10_mag_0.CLK 0.00194f
C897 a_8149_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 8.64e-19
C898 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.00188f
C899 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 7.07e-19
C900 a_n358_4884# CLK_DIV_11_mag_new_0.Q1 0.0186f
C901 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.346f
C902 CLK_div_10_mag_0.Q0 a_10585_n338# 0.00939f
C903 CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_DIV_11_mag_new_0.Q2 0.026f
C904 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_0.Q1 7.24e-19
C905 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.00441f
C906 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_11149_n338# 0.00378f
C907 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 0.131f
C908 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0894f
C909 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0854f
C910 a_8314_n1435# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 2.36e-22
C911 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.108f
C912 a_9282_n1435# CLK_div_10_mag_0.JK_FF_mag_3.QB 1.45e-20
C913 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.K 0.0838f
C914 CLK_div_10_mag_0.JK_FF_mag_1.QB a_2098_n338# 3.33e-19
C915 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.Q0 1.61e-19
C916 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 5.55e-21
C917 CLK_DIV_11_mag_new_0.Q0 a_12282_2771# 0.069f
C918 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q0 4.75f
C919 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_3.QB 0.198f
C920 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 3.4e-19
C921 a_10424_1630# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 1.17e-20
C922 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_10_mag_0.Q1 8.56e-20
C923 RST CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0698f
C924 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 8.58e-20
C925 a_1114_4881# VDD 0.165f
C926 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.Q0 0.0635f
C927 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_0.and2_mag_0.OUT 0.0758f
C928 a_4157_2729# a_4317_2729# 0.0504f
C929 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.904f
C930 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0385f
C931 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.122f
C932 a_1114_4881# CLK_DIV_11_mag_new_0.Q1 0.015f
C933 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.121f
C934 a_6009_2773# VDD 3.56e-19
C935 a_7568_n338# VDD 2.66e-19
C936 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK 1.69e-19
C937 a_4385_759# CLK_div_10_mag_0.JK_FF_mag_2.K 2.81e-19
C938 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 6.01e-19
C939 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00488f
C940 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 8.28e-20
C941 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.nor_3_mag_0.IN3 4.85e-20
C942 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 7.33e-20
C943 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.K 0.00656f
C944 CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 VDD 0.338f
C945 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.065f
C946 a_10424_1630# CLK_div_10_mag_0.CLK 0.00194f
C947 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_10585_n338# 0.00119f
C948 a_5599_1676# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0036f
C949 CLK_div_10_mag_0.JK_FF_mag_2.K a_10585_n338# 0.00486f
C950 CLK_div_10_mag_0.Q0 a_10425_n338# 0.0101f
C951 CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_DIV_11_mag_new_0.Q1 0.203f
C952 a_5269_759# CLK_div_10_mag_0.JK_FF_mag_2.QB 0.00696f
C953 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 1.19e-19
C954 a_4551_n338# CLK_div_10_mag_0.Q1 2.79e-20
C955 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 2.71e-21
C956 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 3.88e-20
C957 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_4551_n338# 0.00119f
C958 CLK_div_10_mag_0.Q0 RST 0.237f
C959 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_0.Q2 0.00311f
C960 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q3 0.00154f
C961 a_7402_759# CLK_div_10_mag_0.Q1 0.00119f
C962 CLK_DIV_11_mag_new_0.Q0 CLK_div_10_mag_0.Q3 0.00274f
C963 a_9346_4996# CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 8.09e-22
C964 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0345f
C965 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 8.16e-20
C966 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 6.03e-20
C967 a_9282_n1435# CLK_div_10_mag_0.and2_mag_0.OUT 0.00138f
C968 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_10590_2727# 1.19e-20
C969 CLK_div_10_mag_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 1.7e-20
C970 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.267f
C971 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 2.51e-19
C972 a_7408_n338# VDD 0.00746f
C973 a_5445_2773# VDD 3.14e-19
C974 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_2.QB 0.198f
C975 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C976 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C977 a_2092_759# CLK_div_10_mag_0.JK_FF_mag_1.QB 0.00695f
C978 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_2816_759# 0.00378f
C979 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00359f
C980 CLK_div_10_mag_0.Q0 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 3.61e-20
C981 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00118f
C982 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 1.54e-21
C983 CLK_div_10_mag_0.Q0 a_9260_n338# 9.45e-19
C984 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.Q2 0.0352f
C985 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C986 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT RST 0.00543f
C987 CLK_div_10_mag_0.JK_FF_mag_2.K a_10425_n338# 0.00111f
C988 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.527f
C989 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 8.16e-20
C990 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0126f
C991 CLK_div_10_mag_0.JK_FF_mag_2.K RST 3.04f
C992 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.103f
C993 a_11149_n338# RST 2.78e-19
C994 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 RST 0.00237f
C995 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.995f
C996 a_n1595_3762# CLK_DIV_11_mag_new_0.Q3 6.63e-20
C997 a_7265_1634# a_7425_1634# 0.0504f
C998 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 8.26e-20
C999 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 3.56e-19
C1000 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 1.36e-19
C1001 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_12282_2771# 0.0114f
C1002 CLK_div_10_mag_0.and2_mag_1.OUT VDD 0.582f
C1003 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 4.42e-19
C1004 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00975f
C1005 a_6609_4975# CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 2.05e-19
C1006 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_3380_759# 0.00372f
C1007 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.235f
C1008 a_7562_759# VDD 0.00891f
C1009 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00335f
C1010 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_10430_2727# 1.52e-20
C1011 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 8.24e-19
C1012 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 0.198f
C1013 CLK_div_10_mag_0.CLK a_1534_n338# 0.00939f
C1014 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.16f
C1015 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.231f
C1016 a_6243_n338# VDD 3.56e-19
C1017 a_4881_2773# VDD 3.14e-19
C1018 CLK_DIV_11_mag_new_0.Q1 a_7562_759# 3.66e-20
C1019 CLK_div_10_mag_0.Q0 CLK 0.00187f
C1020 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 1.85e-19
C1021 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 8.93e-19
C1022 a_4317_2729# CLK_DIV_11_mag_new_0.Q2 2.79e-20
C1023 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.235f
C1024 a_5269_759# RST 0.00211f
C1025 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 RST 0.0189f
C1026 CLK_div_10_mag_0.JK_FF_mag_1.QB VDD 0.92f
C1027 CLK_div_10_mag_0.Q0 a_5109_759# 3.6e-22
C1028 CLK_div_10_mag_0.Q0 a_8696_n338# 6.06e-21
C1029 CLK_div_10_mag_0.JK_FF_mag_2.K a_9260_n338# 7.4e-19
C1030 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_0.K 0.0275f
C1031 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 3.43e-19
C1032 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 7.22e-20
C1033 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0432f
C1034 Vdiv110 CLK_div_10_mag_0.JK_FF_mag_2.K 4.19e-19
C1035 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_DIV_11_mag_new_0.Q2 0.0599f
C1036 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 0.00574f
C1037 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.Q3 0.0345f
C1038 a_n1755_3762# CLK_DIV_11_mag_new_0.Q3 4.15e-19
C1039 CLK_div_10_mag_0.Q0 CLK_DIV_11_mag_new_0.Q3 1.12e-19
C1040 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 0.104f
C1041 CLK_DIV_11_mag_new_0.Q0 a_10590_2727# 2.79e-20
C1042 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 6.71e-19
C1043 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_10_mag_0.Q3 7.16e-20
C1044 RST CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.097f
C1045 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_11718_2771# 2.96e-19
C1046 a_1528_759# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0731f
C1047 a_5904_4934# CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 0.0731f
C1048 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_9123_2775# 0.0114f
C1049 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 3.21e-20
C1050 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 RST 0.0189f
C1051 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 2.59e-19
C1052 a_1746_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00378f
C1053 CLK_div_10_mag_0.CLK a_1374_n338# 0.0101f
C1054 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK 0.267f
C1055 a_5679_n338# VDD 3.14e-19
C1056 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 0.647f
C1057 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.195f
C1058 CLK CLK_div_10_mag_0.JK_FF_mag_2.K 8.07e-21
C1059 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.K 0.00174f
C1060 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_9260_n338# 4.52e-20
C1061 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_8314_n1435# 3.38e-20
C1062 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.11f
C1063 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.121f
C1064 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00118f
C1065 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.109f
C1066 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_3226_n338# 4.52e-20
C1067 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD 0.398f
C1068 a_10250_n1435# CLK_div_10_mag_0.JK_FF_mag_0.K 0.0027f
C1069 CLK_div_10_mag_0.JK_FF_mag_2.K a_8696_n338# 7.4e-19
C1070 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 RST 0.16f
C1071 a_4311_1632# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 1.46e-19
C1072 a_4157_2729# CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.00472f
C1073 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 VDD 0.434f
C1074 CLK_DIV_11_mag_new_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 1.93e-20
C1075 a_11308_1630# RST 0.0017f
C1076 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.122f
C1077 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.397f
C1078 a_11303_759# CLK_div_10_mag_0.Q3 0.0101f
C1079 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_DIV_11_mag_new_0.Q1 3.8e-20
C1080 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 4.44e-20
C1081 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 3.77e-20
C1082 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.Q0 1.99f
C1083 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.11f
C1084 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_11154_2771# 3.33e-19
C1085 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_0.K 1.41e-20
C1086 a_5744_4934# CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 0.0202f
C1087 CLK_div_10_mag_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 4.8e-20
C1088 CLK CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 3.39e-20
C1089 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 9.87e-20
C1090 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q2 0.322f
C1091 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_8559_2775# 2.96e-19
C1092 a_1182_2731# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0732f
C1093 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 1.71e-21
C1094 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.163f
C1095 a_8126_759# CLK_div_10_mag_0.Q1 3.6e-22
C1096 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.0159f
C1097 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00808f
C1098 a_4157_2729# VDD 2.21e-19
C1099 a_5115_n338# VDD 3.14e-19
C1100 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 2.17e-21
C1101 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_10_mag_0.CLK 1.79e-19
C1102 a_7431_2731# CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 8.21e-19
C1103 a_5109_759# a_5269_759# 0.0504f
C1104 a_4545_759# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 1.5e-20
C1105 CLK_div_10_mag_0.Q0 a_1368_759# 0.00335f
C1106 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.237f
C1107 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.133f
C1108 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_11713_n338# 5.94e-20
C1109 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0894f
C1110 CLK_div_10_mag_0.JK_FF_mag_2.K a_8132_n338# 3.12e-19
C1111 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.Q3 2.27e-20
C1112 CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_10_mag_0.Q1 0.0685f
C1113 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 5.18e-19
C1114 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_11718_2771# 4.52e-20
C1115 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.392f
C1116 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00136f
C1117 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 6.88e-21
C1118 a_2098_n338# VDD 3.14e-19
C1119 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_DIV_11_mag_new_0.Q0 1.32e-19
C1120 a_11148_1630# RST 0.00199f
C1121 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.QB 0.25f
C1122 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 0.116f
C1123 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0635f
C1124 a_11143_759# CLK_div_10_mag_0.Q3 0.0102f
C1125 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 1.2e-19
C1126 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_0.Q2 0.00125f
C1127 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_DIV_11_mag_new_0.Q3 0.257f
C1128 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 6.23e-19
C1129 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q2 9.25e-19
C1130 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C1131 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_10590_2727# 0.00392f
C1132 a_2464_1678# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00378f
C1133 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.343f
C1134 a_6009_2773# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00372f
C1135 a_10430_2727# a_10590_2727# 0.0504f
C1136 a_10250_n1435# CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.069f
C1137 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 1.84e-19
C1138 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 a_n1755_2260# 4.44e-20
C1139 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.Q3 0.313f
C1140 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK 9.85e-20
C1141 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_7995_2775# 3.08e-19
C1142 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.00584f
C1143 a_1022_2731# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0203f
C1144 a_9506_4996# CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 2.31e-19
C1145 a_7995_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 0.00378f
C1146 a_9506_4996# CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 1.9e-19
C1147 a_2874_2775# VDD 3.56e-19
C1148 a_7271_2731# CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.00598f
C1149 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.00395f
C1150 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 8.65e-20
C1151 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 6.24e-20
C1152 a_8286_759# VDD 0.00101f
C1153 a_12478_n2129# CLK_div_10_mag_0.JK_FF_mag_2.K 3.02e-19
C1154 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD 0.391f
C1155 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.Q0 0.0349f
C1156 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00943f
C1157 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 3.79e-20
C1158 a_7425_1634# CLK_div_10_mag_0.CLK 0.00192f
C1159 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 5.63e-21
C1160 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_11154_2771# 0.0195f
C1161 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_0.K 6.37e-19
C1162 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 2.85e-20
C1163 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 2.54e-20
C1164 a_10584_1630# RST 0.00256f
C1165 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VDD 0.423f
C1166 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00356f
C1167 a_10579_759# CLK_div_10_mag_0.Q3 0.00789f
C1168 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_8314_n1435# 0.069f
C1169 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.00481f
C1170 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.Q2 0.0398f
C1171 a_7568_n338# CLK_div_10_mag_0.Q2 2.79e-20
C1172 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0129f
C1173 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q1 0.146f
C1174 CLK_div_10_mag_0.CLK a_1528_759# 0.00164f
C1175 a_5445_2773# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.069f
C1176 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.Q0 0.937f
C1177 CLK_div_10_mag_0.JK_FF_mag_2.QB a_4551_n338# 0.00392f
C1178 a_1900_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0733f
C1179 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN a_n350_4053# 3.01e-20
C1180 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q1 1.17e-19
C1181 a_8559_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0059f
C1182 a_9346_4996# CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 3.59e-19
C1183 a_2092_759# VDD 0.00123f
C1184 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.00916f
C1185 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 5.6e-19
C1186 a_2310_2775# VDD 3.14e-19
C1187 a_6009_2773# CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 8.11e-19
C1188 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.K 0.0334f
C1189 a_2252_759# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 2.88e-20
C1190 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C1191 a_12318_n2129# CLK_div_10_mag_0.JK_FF_mag_2.K 9.21e-20
C1192 CLK_DIV_11_mag_new_0.Q2 VDD 2.82f
C1193 a_11303_759# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0733f
C1194 CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 2.75e-19
C1195 a_7265_1634# CLK_div_10_mag_0.CLK 0.00192f
C1196 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 6.18e-19
C1197 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_DIV_11_mag_new_0.Q0 1.61e-19
C1198 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0228f
C1199 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.233f
C1200 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C1201 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 3.98e-20
C1202 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 0.109f
C1203 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.Q1 2.34f
C1204 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 2.13e-20
C1205 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K VDD 0.881f
C1206 a_10424_1630# RST 0.00256f
C1207 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 2.25e-19
C1208 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK 0.32f
C1209 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VDD 0.423f
C1210 a_10419_759# CLK_div_10_mag_0.Q3 0.00335f
C1211 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.103f
C1212 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.Q1 0.00825f
C1213 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT RST 3.84e-20
C1214 RST CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.28f
C1215 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.K 0.0334f
C1216 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_2098_n338# 0.0202f
C1217 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q1 0.111f
C1218 a_7431_2731# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00119f
C1219 a_1740_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0203f
C1220 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.122f
C1221 CLK_div_10_mag_0.CLK a_10590_2727# 1.88e-19
C1222 a_7995_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0697f
C1223 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.236f
C1224 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.109f
C1225 a_1746_2775# VDD 3.14e-19
C1226 a_5445_2773# CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 3.47e-19
C1227 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 VDD 1.16f
C1228 a_10584_1630# CLK 0.00164f
C1229 RST CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0298f
C1230 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 0.299f
C1231 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.652f
C1232 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00125f
C1233 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT RST 0.00539f
C1234 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.0951f
C1235 CLK_DIV_11_mag_new_0.Q1 VDD 3.43f
C1236 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.407f
C1237 a_1900_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 2.88e-20
C1238 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0378f
C1239 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.249f
C1240 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_10_mag_0.JK_FF_mag_2.K 2.11e-21
C1241 a_11143_759# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0203f
C1242 CLK_div_10_mag_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 8.71e-20
C1243 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.Q1 0.447f
C1244 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.K 1.48e-19
C1245 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.25f
C1246 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00233f
C1247 a_5269_759# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0733f
C1248 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.Q2 0.0163f
C1249 a_9277_1678# RST 0.0013f
C1250 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 4.36e-20
C1251 a_7562_759# CLK_div_10_mag_0.Q2 0.00789f
C1252 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 2.63e-19
C1253 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 1.74e-19
C1254 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 3.72e-19
C1255 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.109f
C1256 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_DIV_11_mag_new_0.Q0 0.0444f
C1257 a_1176_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 1.5e-20
C1258 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_10_mag_0.CLK 0.0312f
C1259 CLK_div_10_mag_0.CLK a_10430_2727# 2.7e-19
C1260 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C1261 a_7402_759# RST 0.00247f
C1262 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.Q1 0.018f
C1263 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT RST 0.0596f
C1264 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 5.79e-20
C1265 a_10424_1630# CLK 0.00117f
C1266 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.122f
C1267 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.105f
C1268 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 3.38e-19
C1269 a_1534_n338# RST 7.81e-19
C1270 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.nor_3_mag_0.IN3 0.144f
C1271 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0854f
C1272 RST CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0705f
C1273 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 2.86e-19
C1274 a_2092_759# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0203f
C1275 a_3380_759# RST 0.00138f
C1276 a_1740_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 9.1e-19
C1277 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 6.51e-19
C1278 CLK_div_10_mag_0.Q0 a_2816_759# 0.00859f
C1279 a_10579_759# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 1.5e-20
C1280 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0285f
C1281 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 2.57e-19
C1282 a_11143_759# a_11303_759# 0.0504f
C1283 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 0.00134f
C1284 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK 0.00323f
C1285 a_8149_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 2.88e-20
C1286 a_8713_1678# RST 0.00129f
C1287 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.105f
C1288 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.00995f
C1289 a_8126_759# CLK_div_10_mag_0.JK_FF_mag_3.QB 0.00695f
C1290 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 5.48e-20
C1291 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.642f
C1292 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_3226_n338# 0.00372f
C1293 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0346f
C1294 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_8850_759# 0.0036f
C1295 a_1016_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 1.17e-20
C1296 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.103f
C1297 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 4.68e-20
C1298 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.Q3 8.98e-19
C1299 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.Q1 5.55e-19
C1300 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 5.42e-20
C1301 a_1022_2731# VDD 2.21e-19
C1302 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 2.57e-19
C1303 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 2.01e-19
C1304 RST CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0784f
C1305 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_0.K 5.7e-19
C1306 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.103f
C1307 RST CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.178f
C1308 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 2.51e-19
C1309 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 0.00183f
C1310 a_1374_n338# RST 9.37e-19
C1311 a_2310_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0059f
C1312 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_9282_n1435# 5.1e-20
C1313 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 1.5e-20
C1314 a_1176_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0731f
C1315 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD 1f
C1316 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00602f
C1317 a_10419_759# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 1.17e-20
C1318 CLK a_7402_759# 3.76e-20
C1319 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 1.12e-19
C1320 CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.106f
C1321 a_7989_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 9.1e-19
C1322 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.CLK 1.9e-19
C1323 a_8149_1634# RST 0.00216f
C1324 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.271f
C1325 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 3.27e-20
C1326 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 a_9506_4996# 2.84e-20
C1327 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 3.6e-19
C1328 a_3226_n338# RST 6.14e-19
C1329 a_4875_1632# a_5035_1632# 0.0504f
C1330 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_2662_n338# 0.069f
C1331 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 2.48e-19
C1332 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.519f
C1333 a_5904_4934# CLK_DIV_11_mag_new_0.Q0 0.0121f
C1334 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.Q3 0.124f
C1335 a_10585_n338# CLK_div_10_mag_0.Q3 2.79e-20
C1336 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.122f
C1337 a_1022_2731# a_1182_2731# 0.0504f
C1338 a_5833_759# CLK_div_10_mag_0.Q1 0.00859f
C1339 CLK_DIV_11_mag_new_0.Q2 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 1.87e-19
C1340 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q0 0.00127f
C1341 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_5833_759# 0.0036f
C1342 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_10_mag_0.Q2 8.64e-20
C1343 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 3.53e-19
C1344 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00157f
C1345 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 RST 0.378f
C1346 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.105f
C1347 RST CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 5.36e-20
C1348 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.349f
C1349 a_1746_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0697f
C1350 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 RST 0.00146f
C1351 a_1016_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0202f
C1352 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.651f
C1353 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.K 0.0659f
C1354 CLK_div_10_mag_0.JK_FF_mag_2.K a_7568_n338# 9.32e-19
C1355 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 1.86e-19
C1356 a_7425_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0731f
C1357 CLK_div_10_mag_0.nor_3_mag_0.IN3 Vdiv110 0.0263f
C1358 a_7989_1634# RST 0.00199f
C1359 a_9414_759# VDD 0.00152f
C1360 CLK_div_10_mag_0.CLK a_10579_759# 0.0024f
C1361 CLK CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 8.88e-20
C1362 a_8713_1678# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.00378f
C1363 a_2662_n338# RST 6.14e-19
C1364 CLK CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 7.37e-20
C1365 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 2.03e-20
C1366 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 a_9346_4996# 9.09e-19
C1367 CLK_DIV_11_mag_new_0.Q1 a_9414_759# 5.02e-20
C1368 a_5744_4934# CLK_DIV_11_mag_new_0.Q0 0.00747f
C1369 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 0.00452f
C1370 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.748f
C1371 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 0.00125f
C1372 a_8286_759# CLK_div_10_mag_0.Q2 0.0101f
C1373 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.211f
C1374 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 1.98e-19
C1375 a_n796_2646# CLK_DIV_11_mag_new_0.Q0 3.17e-19
C1376 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C1377 RST CLK_div_10_mag_0.Q3 0.0409f
C1378 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00158f
C1379 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 2.21e-20
C1380 a_6397_759# VDD 0.00152f
C1381 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.and2_mag_1.OUT 1.59e-20
C1382 CLK_DIV_11_mag_new_0.Q3 a_n1755_2260# 0.0111f
C1383 a_8126_759# RST 0.00198f
C1384 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 1.18e-19
C1385 a_4311_1632# CLK_div_10_mag_0.CLK 0.00193f
C1386 CLK_div_10_mag_0.JK_FF_mag_2.K a_7408_n338# 0.00111f
C1387 CLK_div_10_mag_0.Q0 a_6243_n338# 9.26e-19
C1388 CLK_div_10_mag_0.JK_FF_mag_0.K a_10425_n338# 8.64e-19
C1389 a_7265_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0202f
C1390 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 0.0022f
C1391 a_7425_1634# RST 0.00257f
C1392 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.00165f
C1393 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 1.64e-20
C1394 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 1.39e-19
C1395 CLK_div_10_mag_0.JK_FF_mag_0.K RST 1.55e-19
C1396 a_8149_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0733f
C1397 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00109f
C1398 CLK_div_10_mag_0.CLK a_10419_759# 0.0024f
C1399 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 1.74e-19
C1400 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.QB 1.96f
C1401 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0622f
C1402 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK 0.748f
C1403 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 1.72e-19
C1404 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_12277_n338# 0.00372f
C1405 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 0.276f
C1406 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0622f
C1407 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0496f
C1408 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.397f
C1409 CLK_DIV_11_mag_new_0.Q0 RST 0.0676f
C1410 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 9.61e-21
C1411 a_1528_759# RST 0.0037f
C1412 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 1.17e-19
C1413 a_11154_2771# RST 2.67e-19
C1414 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.QB 0.28f
C1415 Vdiv110 CLK_div_10_mag_0.Q3 0.246f
C1416 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 1.7e-19
C1417 RST CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.186f
C1418 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 0.029f
C1419 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C1420 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00718f
C1421 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.25f
C1422 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.0631f
C1423 CLK_div_10_mag_0.and2_mag_1.OUT a_11149_n338# 5.94e-20
C1424 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.36f
C1425 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0622f
C1426 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.Q2 0.291f
C1427 a_7402_759# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 1.17e-20
C1428 a_10424_1630# CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 8.64e-19
C1429 a_4151_1632# CLK_div_10_mag_0.CLK 0.00193f
C1430 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_DIV_11_mag_new_0.and2_mag_3.IN1 2.29e-19
C1431 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 2.18e-21
C1432 a_10419_759# a_10579_759# 0.0504f
C1433 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 4e-19
C1434 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.and2_mag_3.IN1 2.11e-19
C1435 CLK_div_10_mag_0.JK_FF_mag_2.K a_6243_n338# 7.4e-19
C1436 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 5.2e-20
C1437 a_7265_1634# RST 0.00257f
C1438 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 1.57f
C1439 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 3.38e-19
C1440 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.00118f
C1441 a_7989_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0203f
C1442 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.Q1 0.311f
C1443 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 5.08e-20
C1444 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_2.K 9.14e-19
C1445 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_11713_n338# 0.069f
C1446 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.Q0 0.0485f
C1447 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 3.49e-19
C1448 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C1449 VDD CLK_div_10_mag_0.Q2 2.86f
C1450 CLK_div_10_mag_0.and2_mag_0.OUT a_10250_n1435# 0.00138f
C1451 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 1.01e-19
C1452 CLK_DIV_11_mag_new_0.Q1 CLK_div_10_mag_0.Q2 9.88e-20
C1453 a_9346_4996# a_9506_4996# 0.186f
C1454 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0894f
C1455 a_8713_1678# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 4.81e-20
C1456 a_7425_1634# CLK 0.00164f
C1457 CLK_div_10_mag_0.nor_3_mag_0.IN3 a_12478_n2129# 2.44e-20
C1458 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.321f
C1459 a_10590_2727# RST 7.84e-19
C1460 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K VDD 0.866f
C1461 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 2.11e-19
C1462 RST CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0979f
C1463 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_0.nor_3_mag_0.IN3 0.11f
C1464 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.Q1 1.93f
C1465 CLK_div_10_mag_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 2.52e-20
C1466 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD 0.397f
C1467 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 6.22e-20
C1468 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.Q1 1.96f
C1469 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.Q0 0.00187f
C1470 a_9277_1678# CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 2.75e-21
C1471 CLK_div_10_mag_0.Q0 a_5115_n338# 6.43e-21
C1472 CLK_div_10_mag_0.JK_FF_mag_2.K a_5679_n338# 7.4e-19
C1473 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.QB 0.28f
C1474 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.001f
C1475 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00776f
C1476 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 3.61e-21
C1477 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C1478 CLK a_1528_759# 4.62e-19
C1479 CLK_DIV_11_mag_new_0.Q0 CLK 0.538f
C1480 a_6163_1676# RST 0.00129f
C1481 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 2.22e-20
C1482 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.121f
C1483 CLK_DIV_11_mag_new_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 5.36e-20
C1484 CLK a_11154_2771# 6.43e-21
C1485 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_12277_n338# 4.52e-20
C1486 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_3.QB 2.71e-21
C1487 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q2 0.306f
C1488 a_7425_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 1.5e-20
C1489 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0592f
C1490 a_4385_759# CLK_div_10_mag_0.Q1 0.00335f
C1491 a_5035_1632# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 8.64e-19
C1492 a_4151_1632# a_4311_1632# 0.0504f
C1493 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C1494 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_10_mag_0.Q1 0.108f
C1495 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 a_12282_2771# 0.00372f
C1496 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0846f
C1497 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.359f
C1498 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_6243_n338# 4.52e-20
C1499 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 9.75e-21
C1500 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 8.16e-20
C1501 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT RST 0.256f
C1502 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.Q1 0.0529f
C1503 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 7.98e-20
C1504 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 0.00165f
C1505 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 3.44e-20
C1506 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00301f
C1507 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB RST 0.141f
C1508 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_1534_n338# 0.00119f
C1509 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 3.14e-20
C1510 a_7265_1634# CLK 0.00117f
C1511 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 3.94e-19
C1512 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.Q0 0.128f
C1513 a_8850_759# CLK_div_10_mag_0.JK_FF_mag_3.QB 0.00964f
C1514 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_10_mag_0.Q1 1.83e-20
C1515 a_10430_2727# RST 9.41e-19
C1516 CLK_div_10_mag_0.nor_3_mag_0.IN3 a_12318_n2129# 9.02e-19
C1517 CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_DIV_11_mag_new_0.Q0 0.104f
C1518 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.768f
C1519 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.768f
C1520 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_2.QB 2.71e-21
C1521 a_8713_1678# CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 5.58e-22
C1522 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 5.62e-19
C1523 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN a_n1755_2260# 0.069f
C1524 CLK_div_10_mag_0.JK_FF_mag_2.K a_5115_n338# 3.12e-19
C1525 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT VDD 0.664f
C1526 a_5599_1676# RST 0.00129f
C1527 a_8314_n1435# VDD 6e-19
C1528 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 RST 0.0555f
C1529 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.Q1 0.117f
C1530 CLK a_10590_2727# 0.00939f
C1531 a_7265_1634# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 1.17e-20
C1532 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 3.31e-20
C1533 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 a_11718_2771# 0.069f
C1534 a_n1595_3762# CLK_DIV_11_mag_new_0.Q2 8.95e-19
C1535 CLK CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 8.16e-19
C1536 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_0.Q3 0.00357f
C1537 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 1.36e-20
C1538 a_12478_n2129# CLK_div_10_mag_0.Q3 0.019f
C1539 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 3.77e-20
C1540 a_11303_759# RST 0.00146f
C1541 a_4545_759# VDD 0.00863f
C1542 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C1543 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 8.16e-20
C1544 CLK_div_10_mag_0.CLK a_10585_n338# 2.06e-19
C1545 RST CLK_div_10_mag_0.Q1 0.138f
C1546 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00262f
C1547 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 RST 0.0573f
C1548 CLK_DIV_11_mag_new_0.Q3 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 4.08e-20
C1549 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 4.69e-20
C1550 a_2252_759# RST 0.00283f
C1551 a_5833_759# CLK_div_10_mag_0.JK_FF_mag_2.QB 0.00964f
C1552 CLK_div_10_mag_0.Q0 a_2092_759# 0.0102f
C1553 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_9260_n338# 0.00118f
C1554 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 5.51e-20
C1555 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_3226_n338# 0.00118f
C1556 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C1557 a_5035_1632# RST 0.00216f
C1558 a_12277_n338# VDD 3.56e-19
C1559 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_DIV_11_mag_new_0.Q0 0.11f
C1560 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_2.K 0.199f
C1561 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK 0.307f
C1562 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.231f
C1563 a_1528_759# a_1368_759# 0.0504f
C1564 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C1565 a_n1595_3762# CLK_DIV_11_mag_new_0.Q1 1.75e-19
C1566 CLK a_10430_2727# 0.0101f
C1567 CLK_div_10_mag_0.Q0 CLK_DIV_11_mag_new_0.Q2 2.6e-19
C1568 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT RST 0.265f
C1569 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 2.57e-20
C1570 a_8126_759# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0203f
C1571 a_2662_n338# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0059f
C1572 CLK_div_10_mag_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 3.08e-21
C1573 a_11143_759# RST 0.00195f
C1574 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 1.17f
C1575 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.198f
C1576 a_6009_2773# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C1577 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 1.89e-19
C1578 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 RST 0.0225f
C1579 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 2.39e-20
C1580 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.507f
C1581 CLK_div_10_mag_0.CLK a_10425_n338# 2.94e-19
C1582 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 1.83e-19
C1583 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0309f
C1584 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 0.0497f
C1585 CLK CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 7.51e-20
C1586 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00152f
C1587 CLK_div_10_mag_0.CLK RST 0.533f
C1588 a_9414_759# CLK_div_10_mag_0.Q2 0.0157f
C1589 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.191f
C1590 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 2.01e-19
C1591 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_8696_n338# 0.011f
C1592 CLK_div_10_mag_0.Q0 VDD 5.17f
C1593 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 5.11e-19
C1594 a_n1755_3762# VDD 2.21e-19
C1595 a_11303_759# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 2.88e-20
C1596 a_11713_n338# VDD 3.14e-19
C1597 a_11713_n338# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0059f
C1598 a_8850_759# RST 0.00119f
C1599 a_4875_1632# RST 0.00199f
C1600 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_2662_n338# 0.011f
C1601 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_12431_759# 0.00372f
C1602 CLK a_9123_2775# 9.36e-19
C1603 a_n1755_3762# CLK_DIV_11_mag_new_0.Q1 0.00369f
C1604 CLK_DIV_11_mag_new_0.Q2 CLK_div_10_mag_0.JK_FF_mag_2.K 6.12e-21
C1605 CLK CLK_div_10_mag_0.Q1 1.96e-19
C1606 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 2.25e-19
C1607 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C1608 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 2.49e-20
C1609 CLK CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 7.06e-20
C1610 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 3.38e-19
C1611 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_1368_759# 0.0202f
C1612 a_10579_759# RST 0.00247f
C1613 RST CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 1.36e-19
C1614 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.00774f
C1615 a_n350_4053# CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 1.78e-20
C1616 a_5109_759# CLK_div_10_mag_0.Q1 0.0102f
C1617 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00183f
C1618 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0306f
C1619 a_7431_2731# CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.00392f
C1620 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_DIV_11_mag_new_0.Q3 0.0224f
C1621 a_7431_2731# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0732f
C1622 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.28f
C1623 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD 0.432f
C1624 a_n796_2646# CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 0.0177f
C1625 a_7995_2775# RST 3.68e-20
C1626 a_6009_2773# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C1627 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK 9.66e-19
C1628 a_5833_759# RST 0.00119f
C1629 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 2.61e-19
C1630 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q0 0.00115f
C1631 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 9.22e-20
C1632 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0894f
C1633 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VDD 0.647f
C1634 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0013f
C1635 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.K 1.23e-20
C1636 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_8132_n338# 1.43e-19
C1637 CLK CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 3.99e-20
C1638 a_12436_1674# VDD 3.14e-19
C1639 CLK_div_10_mag_0.JK_FF_mag_2.K VDD 1.66f
C1640 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.038f
C1641 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VDD 1.14f
C1642 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.233f
C1643 a_4311_1632# RST 0.00257f
C1644 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.122f
C1645 a_11149_n338# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0697f
C1646 a_11143_759# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.1e-19
C1647 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 4.25e-20
C1648 a_11149_n338# VDD 3.14e-19
C1649 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_11867_759# 0.069f
C1650 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0592f
C1651 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0593f
C1652 CLK a_8559_2775# 9.24e-19
C1653 CLK_DIV_11_mag_new_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.K 7.1e-22
C1654 CLK_div_10_mag_0.CLK CLK 0.0585f
C1655 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C1656 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_12318_n2129# 2.85e-20
C1657 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.Q0 2.42f
C1658 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 3.38e-20
C1659 a_1528_759# CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.46e-19
C1660 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0032f
C1661 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 2.81e-20
C1662 a_10419_759# RST 0.00247f
C1663 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.211f
C1664 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 6.46e-20
C1665 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0052f
C1666 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 1.83e-19
C1667 a_8132_n338# CLK_div_10_mag_0.Q1 1.25e-20
C1668 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_3.QB 2.59e-21
C1669 CLK_DIV_11_mag_new_0.Q2 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.00111f
C1670 CLK_DIV_11_mag_new_0.Q3 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 7.43e-20
C1671 a_7271_2731# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0203f
C1672 a_5445_2773# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.011f
C1673 CLK_div_10_mag_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 2.87e-19
C1674 a_9282_n1435# VDD 3.14e-19
C1675 CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 0.00982f
C1676 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00164f
C1677 a_8559_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 4.52e-20
C1678 a_5269_759# VDD 0.00101f
C1679 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD 0.395f
C1680 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 5.85e-19
C1681 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C1682 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 1.87e-19
C1683 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.Q3 0.341f
C1684 CLK a_10579_759# 1.84e-20
C1685 a_11872_1674# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0036f
C1686 CLK_DIV_11_mag_new_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 5.49e-19
C1687 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C1688 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00637f
C1689 a_11872_1674# VDD 3.14e-19
C1690 a_12431_759# VDD 3.14e-19
C1691 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT VDD 0.343f
C1692 a_10579_759# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0731f
C1693 a_4151_1632# RST 0.00257f
C1694 RST CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 5.45e-20
C1695 a_9506_4996# CLK_DIV_11_mag_new_0.and2_mag_3.OUT 8.64e-19
C1696 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_3.QB 1.33e-20
C1697 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00118f
C1698 a_4545_759# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0731f
C1699 CLK a_7995_2775# 3.8e-19
C1700 a_7402_759# a_7562_759# 0.0504f
C1701 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.16f
C1702 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 4.31e-20
C1703 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0343f
C1704 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.642f
C1705 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_DIV_11_mag_new_0.Q1 3.11e-19
C1706 CLK_div_10_mag_0.JK_FF_mag_3.QB a_10585_n338# 1.41e-20
C1707 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 7.24e-20
C1708 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 3.39e-20
C1709 CLK_div_10_mag_0.JK_FF_mag_1.QB a_4551_n338# 1.41e-20
C1710 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD 0.395f
C1711 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_1114_4881# 0.0131f
C1712 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 0.0238f
C1713 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 8.94e-19
C1714 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_10_mag_0.Q2 0.113f
C1715 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.00147f
C1716 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.00209f
C1717 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 2.46e-20
C1718 a_5744_4934# a_5904_4934# 0.0504f
C1719 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q0 0.0582f
C1720 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C1721 a_10585_n338# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0732f
C1722 CLK_DIV_11_mag_new_0.Q3 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.11f
C1723 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0591f
C1724 a_4311_1632# CLK 0.00164f
C1725 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 3.37e-21
C1726 a_4881_2773# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 1.43e-19
C1727 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.159f
C1728 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 1.03e-19
C1729 a_7995_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0195f
C1730 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00975f
C1731 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.24f
C1732 CLK_div_10_mag_0.JK_FF_mag_1.QB a_1534_n338# 0.00392f
C1733 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00122f
C1734 a_9506_4996# CLK_DIV_11_mag_new_0.Q3 0.0504f
C1735 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 2.62e-20
C1736 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD 0.66f
C1737 a_n796_2646# CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.132f
C1738 a_3380_759# CLK_div_10_mag_0.JK_FF_mag_1.QB 0.0811f
C1739 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 1.77e-19
C1740 a_10419_759# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0202f
C1741 a_11867_759# VDD 3.14e-19
C1742 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_5115_n338# 0.00378f
C1743 a_9346_4996# CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.0105f
C1744 a_3028_1678# RST 0.00154f
C1745 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 5.25e-20
C1746 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.Q1 0.00335f
C1747 CLK_div_10_mag_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 2.97e-20
C1748 a_4311_1632# CLK_DIV_11_mag_new_0.Q3 4.52e-19
C1749 CLK_div_10_mag_0.JK_FF_mag_3.QB a_10425_n338# 1.86e-20
C1750 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.K 4.24e-20
C1751 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q0 0.0072f
C1752 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK 6.61e-20
C1753 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_10_mag_0.CLK 9.82e-21
C1754 CLK_div_10_mag_0.JK_FF_mag_1.QB a_4391_n338# 1.86e-20
C1755 CLK_div_10_mag_0.CLK a_1368_759# 0.00117f
C1756 a_7562_759# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0731f
C1757 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 6.93e-19
C1758 CLK_div_10_mag_0.JK_FF_mag_3.QB RST 0.182f
C1759 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K a_10430_2727# 0.00472f
C1760 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C1761 a_10425_n338# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0203f
C1762 a_n358_4884# CLK_DIV_11_mag_new_0.Q0 0.00718f
C1763 a_4151_1632# CLK 0.00117f
C1764 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 0.275f
C1765 a_4317_2729# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00119f
C1766 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT RST 0.00229f
C1767 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C1768 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.233f
C1769 a_8314_n1435# CLK_div_10_mag_0.Q2 0.00929f
C1770 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_DIV_11_mag_new_0.Q3 8.02e-19
C1771 a_9346_4996# CLK_DIV_11_mag_new_0.Q3 0.0186f
C1772 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.Q1 0.0343f
C1773 a_3028_1678# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.0811f
C1774 a_2252_759# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 8.64e-19
C1775 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.159f
C1776 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 0.048f
C1777 a_11148_1630# VDD 2.21e-19
C1778 RST CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.187f
C1779 CLK_div_10_mag_0.JK_FF_mag_2.QB RST 0.182f
C1780 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_2098_n338# 0.00378f
C1781 a_2464_1678# RST 0.00184f
C1782 a_6609_4975# CLK_DIV_11_mag_new_0.and2_mag_3.OUT 6.43e-19
C1783 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 7.11e-19
C1784 a_1114_4881# CLK_DIV_11_mag_new_0.Q0 0.00589f
C1785 a_6609_4975# CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 3.04e-20
C1786 a_4151_1632# CLK_DIV_11_mag_new_0.Q3 5.83e-19
C1787 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 2.48e-19
C1788 CLK_div_10_mag_0.JK_FF_mag_3.QB a_9260_n338# 0.0114f
C1789 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 1.82e-19
C1790 a_9277_1678# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.00372f
C1791 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.00121f
C1792 CLK_div_10_mag_0.JK_FF_mag_1.QB a_3226_n338# 0.0114f
C1793 a_4385_759# RST 0.00247f
C1794 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0378f
C1795 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 RST 9.24e-20
C1796 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VDD 1.19f
C1797 a_5679_n338# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0059f
C1798 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_8850_759# 0.00378f
C1799 CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_DIV_11_mag_new_0.Q0 0.205f
C1800 a_10425_n338# a_10585_n338# 0.0504f
C1801 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.Q1 0.0409f
C1802 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0286f
C1803 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 3.25e-19
C1804 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 2.48e-19
C1805 a_2464_1678# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.00964f
C1806 RST CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0914f
C1807 a_6609_4975# CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.00476f
C1808 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 RST 0.00434f
C1809 a_10584_1630# CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 1.46e-19
C1810 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 2.47e-19
C1811 a_2310_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C1812 CLK_div_10_mag_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 5.24e-20
C1813 a_1900_1634# RST 0.00349f
C1814 CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 7.14e-19
C1815 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00137f
C1816 a_10584_1630# CLK_DIV_11_mag_new_0.Q1 4.28e-19
C1817 a_5904_4934# CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 8.5e-20
C1818 a_3028_1678# CLK_DIV_11_mag_new_0.Q3 0.0157f
C1819 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_9414_759# 0.00372f
C1820 a_5904_4934# CLK 0.00487f
C1821 a_1740_1634# a_1900_1634# 0.0504f
C1822 CLK_div_10_mag_0.JK_FF_mag_3.QB a_8696_n338# 2.96e-19
C1823 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.Q3 0.00132f
C1824 a_8713_1678# CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.069f
C1825 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 1.05e-19
C1826 CLK_div_10_mag_0.JK_FF_mag_1.QB a_2662_n338# 2.96e-19
C1827 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.321f
C1828 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C1829 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK 0.0011f
C1830 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0707f
C1831 a_5269_759# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 2.88e-20
C1832 a_5115_n338# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0697f
C1833 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q2 0.0549f
C1834 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 3.98e-19
C1835 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 6.91e-20
C1836 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_10_mag_0.CLK 0.0212f
C1837 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 6.36e-19
C1838 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.415f
C1839 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0843f
C1840 CLK_div_10_mag_0.and2_mag_0.OUT Vdiv110 0.119f
C1841 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.Q2 0.622f
C1842 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q1 0.0995f
C1843 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0635f
C1844 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.121f
C1845 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.K 2.08e-20
C1846 a_1900_1634# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.00696f
C1847 a_5109_759# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 1.04e-19
C1848 a_5109_759# CLK_div_10_mag_0.JK_FF_mag_2.QB 0.00695f
C1849 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_5833_759# 0.00378f
C1850 a_6163_1676# CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.0811f
C1851 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 0.129f
C1852 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 3.92e-19
C1853 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0854f
C1854 a_5904_4934# CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.00107f
C1855 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_DIV_11_mag_new_0.Q3 1.51e-19
C1856 a_10424_1630# VDD 2.21e-19
C1857 a_1746_2775# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0195f
C1858 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0598f
C1859 a_1740_1634# RST 0.00207f
C1860 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 1.89e-19
C1861 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.994f
C1862 a_10424_1630# CLK_DIV_11_mag_new_0.Q1 5.5e-19
C1863 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD 0.648f
C1864 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0215f
C1865 a_5744_4934# CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 1.32e-19
C1866 a_2464_1678# CLK_DIV_11_mag_new_0.Q3 0.00859f
C1867 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 8.28e-20
C1868 CLK_div_10_mag_0.JK_FF_mag_3.QB a_8132_n338# 3.25e-19
C1869 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN VDD 0.424f
C1870 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q2 0.103f
C1871 a_3028_1678# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.00372f
C1872 CLK CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.26f
C1873 a_n1595_3762# CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 0.0732f
C1874 a_n796_2646# CLK 2.02e-20
C1875 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.Q1 0.316f
C1876 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_6397_759# 0.00372f
C1877 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.392f
C1878 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 1.82e-19
C1879 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_0.Q1 0.273f
C1880 a_7431_2731# CLK_div_10_mag_0.CLK 1.87e-19
C1881 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 4.27e-20
C1882 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD 0.742f
C1883 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 RST 0.301f
C1884 a_8286_759# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 2.88e-20
C1885 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.Q2 0.0626f
C1886 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.Q2 0.0569f
C1887 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_10_mag_0.Q3 0.11f
C1888 a_5599_1676# CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.00964f
C1889 a_1740_1634# CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.00695f
C1890 CLK_DIV_11_mag_new_0.Q2 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0274f
C1891 RST CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.178f
C1892 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.121f
C1893 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_7568_n338# 0.00119f
C1894 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.198f
C1895 a_5744_4934# CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.00271f
C1896 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 0.0108f
C1897 a_9277_1678# VDD 3.14e-19
C1898 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_2.K 3.88e-20
C1899 a_1176_1634# RST 9.47e-19
C1900 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0702f
C1901 a_9277_1678# CLK_DIV_11_mag_new_0.Q1 0.0157f
C1902 a_4551_n338# VDD 2.66e-19
C1903 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00488f
C1904 a_1900_1634# CLK_DIV_11_mag_new_0.Q3 0.0101f
C1905 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C1906 CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 8.2e-19
C1907 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.and2_mag_1.OUT 0.124f
C1908 a_9282_n1435# CLK_div_10_mag_0.Q2 0.0112f
C1909 a_n350_4053# VDD 3.85e-19
C1910 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_2816_759# 0.069f
C1911 a_7402_759# VDD 0.0132f
C1912 a_2464_1678# CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.069f
C1913 a_n1755_3762# CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 0.0202f
C1914 CLK_div_10_mag_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 7.34e-20
C1915 CLK RST 3.52f
C1916 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_10_mag_0.Q2 0.0635f
C1917 a_7568_n338# CLK_div_10_mag_0.Q1 0.00939f
C1918 a_n350_4053# CLK_DIV_11_mag_new_0.Q1 0.0205f
C1919 a_7271_2731# CLK_div_10_mag_0.CLK 2.69e-19
C1920 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 6.87e-20
C1921 RST CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0779f
C1922 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 2.71e-21
C1923 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.642f
C1924 a_1740_1634# CLK 6.8e-19
C1925 a_1534_n338# VDD 2.66e-19
C1926 VDD CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 1.18f
C1927 a_5109_759# RST 0.00195f
C1928 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_DIV_11_mag_new_0.Q0 0.0128f
C1929 a_3380_759# VDD 0.00152f
C1930 CLK_DIV_11_mag_new_0.Q2 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 7.94e-20
C1931 a_n1762_4447# CLK_DIV_11_mag_new_0.Q3 0.00572f
C1932 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C1933 CLK_div_10_mag_0.Q0 a_4545_759# 0.00166f
C1934 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 3.4e-19
C1935 CLK_DIV_11_mag_new_0.Q1 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00917f
C1936 a_5035_1632# CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.00696f
C1937 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 8.26e-20
C1938 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.00125f
C1939 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 8.16e-20
C1940 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.QB 0.25f
C1941 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K RST 0.00458f
C1942 RST CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.285f
C1943 CLK_DIV_11_mag_new_0.Q3 RST 0.151f
C1944 a_8713_1678# VDD 3.14e-19
C1945 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00243f
C1946 a_1016_1634# RST 8.14e-19
C1947 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.109f
C1948 a_8713_1678# CLK_DIV_11_mag_new_0.Q1 0.00859f
C1949 a_4391_n338# VDD 3.78e-19
C1950 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK 0.64f
C1951 a_1740_1634# CLK_DIV_11_mag_new_0.Q3 0.0102f
C1952 CLK_div_10_mag_0.and2_mag_0.OUT a_12478_n2129# 0.00894f
C1953 a_10250_n1435# CLK_div_10_mag_0.and2_mag_1.OUT 2.94e-20
C1954 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 9.06e-20
C1955 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.0654f
C1956 a_n1755_3762# a_n1595_3762# 0.0504f
C1957 CLK CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 2.51e-20
C1958 a_5599_1676# CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.00378f
C1959 a_7408_n338# CLK_div_10_mag_0.Q1 0.0101f
C1960 CLK_div_10_mag_0.CLK CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.00119f
C1961 VDD a_n1755_2260# 3.14e-19
C1962 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.768f
C1963 a_1176_1634# CLK 0.00253f
C1964 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.653f
C1965 a_1374_n338# VDD 0.00752f
C1966 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 2.8e-19
C1967 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_10_mag_0.Q3 0.0635f
C1968 a_8132_n338# RST 1.23e-20
C1969 CLK_DIV_11_mag_new_0.Q0 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 1.71e-21
C1970 CLK_DIV_11_mag_new_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 5.5e-20
C1971 a_8696_n338# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0059f
C1972 CLK_DIV_11_mag_new_0.Q1 a_n1755_2260# 0.00347f
C1973 a_12478_n2129# VSS 0.0371f
C1974 a_12318_n2129# VSS 0.038f
C1975 Vdiv110 VSS 0.525f
C1976 CLK_div_10_mag_0.nor_3_mag_0.IN3 VSS 0.337f
C1977 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS 0.669f
C1978 CLK_div_10_mag_0.and2_mag_1.OUT VSS 0.706f
C1979 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS 0.435f
C1980 a_10250_n1435# VSS 0.0679f
C1981 CLK_div_10_mag_0.and2_mag_0.OUT VSS 0.823f
C1982 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS 0.438f
C1983 a_9282_n1435# VSS 0.0679f
C1984 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.436f
C1985 a_8314_n1435# VSS 0.0676f
C1986 a_12277_n338# VSS 0.0676f
C1987 a_11713_n338# VSS 0.0676f
C1988 a_11149_n338# VSS 0.0676f
C1989 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.414f
C1990 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C1991 a_10585_n338# VSS 0.0343f
C1992 a_10425_n338# VSS 0.0881f
C1993 a_9260_n338# VSS 0.0676f
C1994 a_8696_n338# VSS 0.0676f
C1995 a_8132_n338# VSS 0.0676f
C1996 CLK_div_10_mag_0.JK_FF_mag_0.K VSS 0.633f
C1997 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS 0.414f
C1998 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VSS 0.509f
C1999 a_7568_n338# VSS 0.0343f
C2000 a_7408_n338# VSS 0.0881f
C2001 a_6243_n338# VSS 0.0676f
C2002 a_5679_n338# VSS 0.0676f
C2003 a_5115_n338# VSS 0.0676f
C2004 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS 0.415f
C2005 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VSS 0.509f
C2006 a_4551_n338# VSS 0.0343f
C2007 a_4391_n338# VSS 0.0881f
C2008 a_3226_n338# VSS 0.0676f
C2009 a_2662_n338# VSS 0.0676f
C2010 a_2098_n338# VSS 0.0676f
C2011 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C2012 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.509f
C2013 a_1534_n338# VSS 0.0343f
C2014 a_1374_n338# VSS 0.0881f
C2015 CLK_div_10_mag_0.JK_FF_mag_2.K VSS 3.1f
C2016 a_12431_759# VSS 0.0675f
C2017 a_11867_759# VSS 0.0676f
C2018 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.415f
C2019 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.753f
C2020 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.807f
C2021 a_11303_759# VSS 0.0343f
C2022 a_11143_759# VSS 0.0881f
C2023 a_10579_759# VSS 0.0343f
C2024 a_10419_759# VSS 0.0881f
C2025 CLK_div_10_mag_0.JK_FF_mag_3.QB VSS 0.877f
C2026 a_9414_759# VSS 0.0675f
C2027 a_8850_759# VSS 0.0676f
C2028 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS 0.416f
C2029 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 VSS 0.693f
C2030 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VSS 0.808f
C2031 a_8286_759# VSS 0.0343f
C2032 a_8126_759# VSS 0.0881f
C2033 a_7562_759# VSS 0.0343f
C2034 a_7402_759# VSS 0.0881f
C2035 CLK_div_10_mag_0.JK_FF_mag_2.QB VSS 0.879f
C2036 a_6397_759# VSS 0.0675f
C2037 a_5833_759# VSS 0.0676f
C2038 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS 0.415f
C2039 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 VSS 0.696f
C2040 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VSS 0.809f
C2041 a_5269_759# VSS 0.0343f
C2042 a_5109_759# VSS 0.0881f
C2043 a_4545_759# VSS 0.0343f
C2044 a_4385_759# VSS 0.0881f
C2045 CLK_div_10_mag_0.JK_FF_mag_1.QB VSS 0.9f
C2046 a_3380_759# VSS 0.0675f
C2047 a_2816_759# VSS 0.0676f
C2048 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.416f
C2049 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.902f
C2050 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.81f
C2051 a_2252_759# VSS 0.0343f
C2052 a_2092_759# VSS 0.0881f
C2053 a_1528_759# VSS 0.0343f
C2054 a_1368_759# VSS 0.0881f
C2055 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.724f
C2056 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.519f
C2057 CLK_div_10_mag_0.Q3 VSS 1.67f
C2058 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS 0.725f
C2059 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VSS 0.54f
C2060 CLK_div_10_mag_0.Q2 VSS 2.23f
C2061 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS 0.726f
C2062 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VSS 0.539f
C2063 CLK_div_10_mag_0.Q1 VSS 2.6f
C2064 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.724f
C2065 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.539f
C2066 CLK_div_10_mag_0.Q0 VSS 3.5f
C2067 a_12436_1674# VSS 0.0696f
C2068 a_11872_1674# VSS 0.0698f
C2069 a_11308_1630# VSS 0.0378f
C2070 a_11148_1630# VSS 0.0916f
C2071 a_10584_1630# VSS 0.0378f
C2072 a_10424_1630# VSS 0.0917f
C2073 a_9277_1678# VSS 0.069f
C2074 a_8713_1678# VSS 0.0691f
C2075 a_8149_1634# VSS 0.0367f
C2076 a_7989_1634# VSS 0.0905f
C2077 a_7425_1634# VSS 0.0368f
C2078 a_7265_1634# VSS 0.0906f
C2079 a_6163_1676# VSS 0.0693f
C2080 a_5599_1676# VSS 0.0694f
C2081 a_5035_1632# VSS 0.0372f
C2082 a_4875_1632# VSS 0.0911f
C2083 a_4311_1632# VSS 0.0373f
C2084 a_4151_1632# VSS 0.0911f
C2085 a_3028_1678# VSS 0.069f
C2086 a_2464_1678# VSS 0.0691f
C2087 a_1900_1634# VSS 0.0367f
C2088 a_1740_1634# VSS 0.0905f
C2089 a_1176_1634# VSS 0.0368f
C2090 a_1016_1634# VSS 0.0906f
C2091 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS 0.419f
C2092 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT VSS 0.551f
C2093 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS 0.419f
C2094 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT VSS 0.549f
C2095 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.42f
C2096 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.551f
C2097 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.418f
C2098 RST VSS 4.92f
C2099 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.547f
C2100 a_n1755_2260# VSS 0.0716f
C2101 a_12282_2771# VSS 0.0744f
C2102 a_11718_2771# VSS 0.0745f
C2103 a_11154_2771# VSS 0.0744f
C2104 a_10590_2727# VSS 0.047f
C2105 a_10430_2727# VSS 0.101f
C2106 a_9123_2775# VSS 0.0734f
C2107 a_8559_2775# VSS 0.0735f
C2108 a_7995_2775# VSS 0.0735f
C2109 a_7431_2731# VSS 0.0449f
C2110 a_7271_2731# VSS 0.0987f
C2111 a_6009_2773# VSS 0.0739f
C2112 a_5445_2773# VSS 0.074f
C2113 a_4881_2773# VSS 0.0739f
C2114 a_4317_2729# VSS 0.0459f
C2115 a_4157_2729# VSS 0.0997f
C2116 a_2874_2775# VSS 0.0737f
C2117 a_2310_2775# VSS 0.0737f
C2118 a_1746_2775# VSS 0.0737f
C2119 a_1182_2731# VSS 0.0454f
C2120 a_1022_2731# VSS 0.0992f
C2121 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS 0.425f
C2122 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 VSS 0.906f
C2123 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS 0.754f
C2124 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VSS 0.83f
C2125 CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VSS 0.549f
C2126 CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB VSS 0.954f
C2127 CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.612f
C2128 a_n796_2646# VSS 0.0247f
C2129 CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.45f
C2130 CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 VSS 0.504f
C2131 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS 0.424f
C2132 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 VSS 0.86f
C2133 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS 0.742f
C2134 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT VSS 0.827f
C2135 CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT VSS 0.543f
C2136 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.424f
C2137 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.831f
C2138 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.743f
C2139 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.829f
C2140 CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.546f
C2141 CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB VSS 0.912f
C2142 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.424f
C2143 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.844f
C2144 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.741f
C2145 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.826f
C2146 CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.544f
C2147 CLK_DIV_11_mag_new_0.JK_FF_mag_0.K VSS 1.92f
C2148 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K VSS 3.1f
C2149 CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 VSS 0.401f
C2150 CLK_DIV_11_mag_new_0.nand3_mag_0.OUT VSS 0.585f
C2151 a_n1595_3762# VSS 0.0343f
C2152 a_n1755_3762# VSS 0.0881f
C2153 CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN VSS 0.464f
C2154 a_n350_4053# VSS 0.0676f
C2155 CLK_div_10_mag_0.CLK VSS 11.8f
C2156 a_9506_4996# VSS 0.0376f
C2157 a_9346_4996# VSS 0.0391f
C2158 a_6609_4975# VSS 0.0693f
C2159 a_5904_4934# VSS 0.0362f
C2160 a_5744_4934# VSS 0.0901f
C2161 a_n1762_4447# VSS 0.0678f
C2162 CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT VSS 1.03f
C2163 CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 VSS 0.555f
C2164 CLK_DIV_11_mag_new_0.JK_FF_mag_3.K VSS 2.89f
C2165 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN VSS 0.676f
C2166 CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT VSS 0.678f
C2167 CLK_DIV_11_mag_new_0.and2_mag_3.OUT VSS 1.93f
C2168 CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VSS 0.597f
C2169 a_1114_4881# VSS 0.0247f
C2170 CLK_DIV_11_mag_new_0.JK_FF_mag_2.K VSS 2.86f
C2171 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 VSS 18.6f
C2172 CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VSS 2.52f
C2173 CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VSS 0.589f
C2174 a_n358_4884# VSS 0.0247f
C2175 CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VSS 0.453f
C2176 CLK_DIV_11_mag_new_0.Q3 VSS 7.03f
C2177 CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 VSS 0.532f
C2178 CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VSS 0.457f
C2179 CLK_DIV_11_mag_new_0.Q1 VSS 6.68f
C2180 CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS 0.701f
C2181 CLK_DIV_11_mag_new_0.Q2 VSS 6.59f
C2182 CLK VSS 7.58f
C2183 CLK_DIV_11_mag_new_0.Q0 VSS 6.01f
C2184 CLK_DIV_11_mag_new_0.and2_mag_3.IN1 VSS 0.834f
C2185 CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VSS 0.741f
C2186 VDD VSS 0.149p
C2187 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t5 VSS 0.154f
C2188 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t7 VSS 0.0457f
C2189 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n0 VSS 0.158f
C2190 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t6 VSS 0.0621f
C2191 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t8 VSS 0.0779f
C2192 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n1 VSS 0.184f
C2193 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t4 VSS 0.109f
C2194 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t3 VSS 0.0696f
C2195 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n2 VSS 0.193f
C2196 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n3 VSS 1.79f
C2197 CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t1 VSS 0.589f
C2198 CLK.n0 VSS 0.00273f
C2199 CLK.n1 VSS 0.00224f
C2200 CLK.n2 VSS 0.00449f
C2201 CLK.t22 VSS 0.0178f
C2202 CLK.t23 VSS 0.027f
C2203 CLK.n3 VSS 0.0478f
C2204 CLK.n4 VSS 0.00616f
C2205 CLK.n5 VSS 0.00873f
C2206 CLK.n6 VSS 0.0884f
C2207 CLK.n7 VSS 0.0897f
C2208 CLK.n8 VSS 0.00449f
C2209 CLK.t24 VSS 0.0178f
C2210 CLK.t25 VSS 0.027f
C2211 CLK.n9 VSS 0.0478f
C2212 CLK.n10 VSS 0.00616f
C2213 CLK.n11 VSS 0.00222f
C2214 CLK.n12 VSS 0.0566f
C2215 CLK.n13 VSS 0.0561f
C2216 CLK.t3 VSS 0.0224f
C2217 CLK.t10 VSS 0.00571f
C2218 CLK.n14 VSS 0.037f
C2219 CLK.n15 VSS 0.00785f
C2220 CLK.n16 VSS 0.00273f
C2221 CLK.n17 VSS 0.00224f
C2222 CLK.n18 VSS 0.00449f
C2223 CLK.t8 VSS 0.0178f
C2224 CLK.t11 VSS 0.027f
C2225 CLK.n19 VSS 0.0478f
C2226 CLK.n20 VSS 0.00616f
C2227 CLK.n21 VSS 0.00873f
C2228 CLK.n22 VSS 0.0884f
C2229 CLK.n23 VSS 0.0897f
C2230 CLK.n24 VSS 0.00449f
C2231 CLK.t21 VSS 0.0178f
C2232 CLK.t15 VSS 0.027f
C2233 CLK.n25 VSS 0.0478f
C2234 CLK.n26 VSS 0.00616f
C2235 CLK.n27 VSS 0.00222f
C2236 CLK.n28 VSS 0.0566f
C2237 CLK.n29 VSS 0.0561f
C2238 CLK.t12 VSS 0.0224f
C2239 CLK.t20 VSS 0.00571f
C2240 CLK.n30 VSS 0.037f
C2241 CLK.n31 VSS 0.00785f
C2242 CLK.n32 VSS 0.00775f
C2243 CLK.n33 VSS 0.0161f
C2244 CLK.n34 VSS 0.00273f
C2245 CLK.n35 VSS 0.00224f
C2246 CLK.n36 VSS 0.00449f
C2247 CLK.t7 VSS 0.0178f
C2248 CLK.t9 VSS 0.027f
C2249 CLK.n37 VSS 0.0478f
C2250 CLK.n38 VSS 0.00616f
C2251 CLK.n39 VSS 0.00873f
C2252 CLK.n40 VSS 0.0884f
C2253 CLK.n41 VSS 0.0897f
C2254 CLK.n42 VSS 0.00449f
C2255 CLK.t13 VSS 0.0178f
C2256 CLK.t14 VSS 0.027f
C2257 CLK.n43 VSS 0.0478f
C2258 CLK.n44 VSS 0.00616f
C2259 CLK.n45 VSS 0.00222f
C2260 CLK.n46 VSS 0.0566f
C2261 CLK.n47 VSS 0.0561f
C2262 CLK.t17 VSS 0.0224f
C2263 CLK.t2 VSS 0.00571f
C2264 CLK.n48 VSS 0.037f
C2265 CLK.n49 VSS 0.00785f
C2266 CLK.n50 VSS 0.00775f
C2267 CLK.n51 VSS 0.0161f
C2268 CLK.n52 VSS 0.0144f
C2269 CLK.n53 VSS 0.00242f
C2270 CLK.t0 VSS 0.0178f
C2271 CLK.t1 VSS 0.027f
C2272 CLK.n54 VSS 0.048f
C2273 CLK.n55 VSS 0.00721f
C2274 CLK.n56 VSS 0.00294f
C2275 CLK.n57 VSS 0.241f
C2276 CLK.n58 VSS 0.00273f
C2277 CLK.n59 VSS 0.00224f
C2278 CLK.n60 VSS 0.00449f
C2279 CLK.t4 VSS 0.0178f
C2280 CLK.t5 VSS 0.027f
C2281 CLK.n61 VSS 0.0478f
C2282 CLK.n62 VSS 0.00616f
C2283 CLK.n63 VSS 0.00873f
C2284 CLK.n64 VSS 0.0884f
C2285 CLK.n65 VSS 0.0897f
C2286 CLK.n66 VSS 0.00449f
C2287 CLK.t18 VSS 0.0178f
C2288 CLK.t19 VSS 0.027f
C2289 CLK.n67 VSS 0.0478f
C2290 CLK.n68 VSS 0.00616f
C2291 CLK.n69 VSS 0.00222f
C2292 CLK.n70 VSS 0.0566f
C2293 CLK.n71 VSS 0.0561f
C2294 CLK.t16 VSS 0.00571f
C2295 CLK.t6 VSS 0.0224f
C2296 CLK.n72 VSS 0.037f
C2297 CLK.n73 VSS 0.00785f
C2298 CLK.n74 VSS 0.00775f
C2299 CLK.n75 VSS 0.0161f
C2300 CLK.n76 VSS 0.377f
C2301 CLK.n77 VSS 2.22f
C2302 CLK.n78 VSS 2.13f
C2303 CLK.n79 VSS 0.37f
C2304 CLK.n80 VSS 0.0161f
C2305 CLK.n81 VSS 0.331f
C2306 RST.t9 VSS 0.019f
C2307 RST.t10 VSS 0.0288f
C2308 RST.n0 VSS 0.051f
C2309 RST.n1 VSS 0.00933f
C2310 RST.n2 VSS 0.00315f
C2311 RST.n3 VSS 0.0115f
C2312 RST.n4 VSS 0.0175f
C2313 RST.n5 VSS 0.0105f
C2314 RST.n6 VSS 0.00391f
C2315 RST.t11 VSS 0.019f
C2316 RST.t12 VSS 0.0288f
C2317 RST.n7 VSS 0.051f
C2318 RST.n8 VSS 0.0072f
C2319 RST.n9 VSS 0.0028f
C2320 RST.n10 VSS 0.00392f
C2321 RST.n11 VSS 0.0137f
C2322 RST.n12 VSS 0.0012f
C2323 RST.n13 VSS 0.0361f
C2324 RST.n14 VSS 0.727f
C2325 RST.n15 VSS 0.725f
C2326 RST.n16 VSS 0.715f
C2327 RST.n17 VSS 0.716f
C2328 RST.n18 VSS 0.011f
C2329 RST.n19 VSS 0.00208f
C2330 RST.t0 VSS 0.019f
C2331 RST.t1 VSS 0.0288f
C2332 RST.n20 VSS 0.051f
C2333 RST.n21 VSS 0.00764f
C2334 RST.n22 VSS 0.00392f
C2335 RST.n23 VSS 0.0018f
C2336 RST.n24 VSS 8.12e-19
C2337 RST.n25 VSS 0.00379f
C2338 RST.n26 VSS 0.00201f
C2339 RST.n27 VSS 0.0111f
C2340 RST.n28 VSS 0.00808f
C2341 RST.n29 VSS 0.712f
C2342 RST.n30 VSS 0.714f
C2343 RST.n31 VSS 0.0107f
C2344 RST.n32 VSS 0.0122f
C2345 RST.n33 VSS 0.00406f
C2346 RST.t5 VSS 0.019f
C2347 RST.t6 VSS 0.0288f
C2348 RST.n34 VSS 0.051f
C2349 RST.n35 VSS 0.0071f
C2350 RST.n36 VSS 0.00244f
C2351 RST.n37 VSS 0.0012f
C2352 RST.n38 VSS 0.00332f
C2353 RST.n39 VSS 0.00783f
C2354 RST.n40 VSS 0.00138f
C2355 RST.n41 VSS 0.0923f
C2356 RST.n42 VSS 0.215f
C2357 RST.n43 VSS 0.0149f
C2358 RST.n44 VSS 0.00235f
C2359 RST.n45 VSS 0.00221f
C2360 RST.n46 VSS 0.00236f
C2361 RST.n47 VSS 2.64e-19
C2362 RST.t15 VSS 0.0288f
C2363 RST.n48 VSS 0.0357f
C2364 RST.t3 VSS 0.0173f
C2365 RST.n49 VSS 0.017f
C2366 RST.n50 VSS 0.00639f
C2367 RST.n51 VSS 0.0115f
C2368 RST.t2 VSS 0.0288f
C2369 RST.t7 VSS 0.019f
C2370 RST.n52 VSS 0.051f
C2371 RST.n53 VSS 0.0275f
C2372 RST.t4 VSS 0.0288f
C2373 RST.t13 VSS 0.019f
C2374 RST.n54 VSS 0.051f
C2375 RST.n55 VSS 0.278f
C2376 RST.n56 VSS 0.866f
C2377 RST.n57 VSS 0.717f
C2378 RST.t8 VSS 0.0288f
C2379 RST.t14 VSS 0.019f
C2380 RST.n58 VSS 0.051f
C2381 RST.n59 VSS 0.026f
C2382 RST.n60 VSS 0.053f
C2383 RST.n61 VSS 0.345f
C2384 RST.n62 VSS 0.209f
C2385 RST.n63 VSS 0.252f
C2386 CLK_div_10_mag_0.JK_FF_mag_2.K.n0 VSS 0.0639f
C2387 CLK_div_10_mag_0.JK_FF_mag_2.K.t7 VSS 0.0298f
C2388 CLK_div_10_mag_0.JK_FF_mag_2.K.t5 VSS 0.023f
C2389 CLK_div_10_mag_0.JK_FF_mag_2.K.n1 VSS 0.059f
C2390 CLK_div_10_mag_0.JK_FF_mag_2.K.t8 VSS 0.0207f
C2391 CLK_div_10_mag_0.JK_FF_mag_2.K.t6 VSS 0.0324f
C2392 CLK_div_10_mag_0.JK_FF_mag_2.K.n2 VSS 0.0574f
C2393 CLK_div_10_mag_0.JK_FF_mag_2.K.n3 VSS 1.11f
C2394 CLK_div_10_mag_0.JK_FF_mag_2.K.t4 VSS 0.0185f
C2395 CLK_div_10_mag_0.JK_FF_mag_2.K.t3 VSS 0.0231f
C2396 CLK_div_10_mag_0.JK_FF_mag_2.K.n4 VSS 0.0547f
C2397 CLK_div_10_mag_0.JK_FF_mag_2.K.n5 VSS 0.368f
C2398 CLK_div_10_mag_0.JK_FF_mag_2.K.t1 VSS 0.0144f
C2399 CLK_div_10_mag_0.JK_FF_mag_2.K.n6 VSS 0.0144f
C2400 CLK_div_10_mag_0.JK_FF_mag_2.K.n7 VSS 0.0308f
C2401 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t2 VSS 0.0207f
C2402 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t5 VSS 0.0271f
C2403 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n0 VSS 0.0537f
C2404 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t3 VSS 0.0273f
C2405 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t4 VSS 0.0207f
C2406 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n1 VSS 0.0537f
C2407 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n2 VSS 0.675f
C2408 CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n3 VSS 0.0327f
C2409 VDD.t20 VSS 0.0721f
C2410 VDD.t12 VSS 0.0558f
C2411 VDD.t301 VSS 0.00335f
C2412 VDD.n0 VSS 0.00335f
C2413 VDD.n1 VSS 0.00732f
C2414 VDD.t325 VSS 0.00816f
C2415 VDD.n2 VSS 0.00815f
C2416 VDD.n3 VSS 0.072f
C2417 VDD.t440 VSS 0.108f
C2418 VDD.n4 VSS 0.00815f
C2419 VDD.t321 VSS 0.00816f
C2420 VDD.n5 VSS 0.00815f
C2421 VDD.n6 VSS 0.00815f
C2422 VDD.t182 VSS 0.0857f
C2423 VDD.n7 VSS 0.0436f
C2424 VDD.t229 VSS 0.00816f
C2425 VDD.n8 VSS 0.00815f
C2426 VDD.t228 VSS 0.0782f
C2427 VDD.t443 VSS 0.0857f
C2428 VDD.n9 VSS 0.0436f
C2429 VDD.t274 VSS 0.00816f
C2430 VDD.t103 VSS 0.00335f
C2431 VDD.n10 VSS 0.00335f
C2432 VDD.n11 VSS 0.00732f
C2433 VDD.t273 VSS 0.0713f
C2434 VDD.n12 VSS 0.281f
C2435 VDD.t102 VSS 0.034f
C2436 VDD.t390 VSS 0.0444f
C2437 VDD.n13 VSS 0.0436f
C2438 VDD.t435 VSS 0.00816f
C2439 VDD.t173 VSS 0.00335f
C2440 VDD.n14 VSS 0.00335f
C2441 VDD.n15 VSS 0.00732f
C2442 VDD.t434 VSS 0.0782f
C2443 VDD.t172 VSS 0.0955f
C2444 VDD.t22 VSS 0.0444f
C2445 VDD.t269 VSS 0.0897f
C2446 VDD.n16 VSS 0.0436f
C2447 VDD.t270 VSS 0.00874f
C2448 VDD.n17 VSS 0.0628f
C2449 VDD.n18 VSS 0.0464f
C2450 VDD.n19 VSS 0.0477f
C2451 VDD.n20 VSS 0.0253f
C2452 VDD.n21 VSS 0.0464f
C2453 VDD.n22 VSS 0.0475f
C2454 VDD.n23 VSS 0.0282f
C2455 VDD.n24 VSS 0.0404f
C2456 VDD.n25 VSS 0.0376f
C2457 VDD.n26 VSS 0.0282f
C2458 VDD.n27 VSS 0.0704f
C2459 VDD.t168 VSS 0.00812f
C2460 VDD.t261 VSS 0.00816f
C2461 VDD.n28 VSS 0.0775f
C2462 VDD.t167 VSS 0.0721f
C2463 VDD.t179 VSS 0.0558f
C2464 VDD.t209 VSS 0.00335f
C2465 VDD.n29 VSS 0.00335f
C2466 VDD.n30 VSS 0.00732f
C2467 VDD.t175 VSS 0.00816f
C2468 VDD.n31 VSS 0.00815f
C2469 VDD.n32 VSS 0.0708f
C2470 VDD.t369 VSS 0.0725f
C2471 VDD.t370 VSS 0.00812f
C2472 VDD.n33 VSS 0.0597f
C2473 VDD.t176 VSS 0.0643f
C2474 VDD.n34 VSS 0.00815f
C2475 VDD.t219 VSS 0.00812f
C2476 VDD.t26 VSS 0.00816f
C2477 VDD.n35 VSS 0.0759f
C2478 VDD.t218 VSS 0.0725f
C2479 VDD.t64 VSS 0.0643f
C2480 VDD.n36 VSS 0.00815f
C2481 VDD.t341 VSS 0.00812f
C2482 VDD.t455 VSS 0.00812f
C2483 VDD.n37 VSS 0.095f
C2484 VDD.t403 VSS 0.104f
C2485 VDD.t404 VSS 0.017f
C2486 VDD.t339 VSS 0.0317f
C2487 VDD.n38 VSS 0.0509f
C2488 VDD.t162 VSS 0.207f
C2489 VDD.t460 VSS 0.0661f
C2490 VDD.n39 VSS 0.0766f
C2491 VDD.t338 VSS 0.211f
C2492 VDD.n40 VSS 0.0988f
C2493 VDD.n41 VSS 0.103f
C2494 VDD.n42 VSS 0.0629f
C2495 VDD.n43 VSS 0.115f
C2496 VDD.t454 VSS 0.0675f
C2497 VDD.t340 VSS 0.116f
C2498 VDD.n44 VSS 0.0752f
C2499 VDD.n45 VSS 0.0597f
C2500 VDD.n46 VSS 0.0708f
C2501 VDD.n47 VSS 0.0426f
C2502 VDD.n48 VSS 0.0506f
C2503 VDD.t25 VSS 0.0558f
C2504 VDD.n49 VSS 0.118f
C2505 VDD.n50 VSS 0.0597f
C2506 VDD.n51 VSS 0.0708f
C2507 VDD.t61 VSS 0.00816f
C2508 VDD.n52 VSS 0.0759f
C2509 VDD.n53 VSS 0.0426f
C2510 VDD.n54 VSS 0.0506f
C2511 VDD.t60 VSS 0.0558f
C2512 VDD.n55 VSS 0.118f
C2513 VDD.t67 VSS 0.0643f
C2514 VDD.t174 VSS 0.098f
C2515 VDD.n56 VSS 0.0506f
C2516 VDD.n57 VSS 0.0426f
C2517 VDD.n58 VSS 0.196f
C2518 VDD.t272 VSS 0.00819f
C2519 VDD.n59 VSS 0.00815f
C2520 VDD.n60 VSS 0.0404f
C2521 VDD.t109 VSS 0.108f
C2522 VDD.n61 VSS 0.00815f
C2523 VDD.t373 VSS 0.00816f
C2524 VDD.n62 VSS 0.00815f
C2525 VDD.t8 VSS 0.00812f
C2526 VDD.t437 VSS 0.00816f
C2527 VDD.n63 VSS 0.0385f
C2528 VDD.t7 VSS 0.0721f
C2529 VDD.t9 VSS 0.0558f
C2530 VDD.t221 VSS 0.00335f
C2531 VDD.n64 VSS 0.00335f
C2532 VDD.n65 VSS 0.00732f
C2533 VDD.t323 VSS 0.00816f
C2534 VDD.n66 VSS 0.00815f
C2535 VDD.n67 VSS 0.0404f
C2536 VDD.t331 VSS 0.108f
C2537 VDD.n68 VSS 0.00815f
C2538 VDD.t33 VSS 0.00816f
C2539 VDD.n69 VSS 0.00815f
C2540 VDD.n70 VSS 0.00815f
C2541 VDD.t157 VSS 0.106f
C2542 VDD.n71 VSS 0.0506f
C2543 VDD.t483 VSS 0.00816f
C2544 VDD.n72 VSS 0.00815f
C2545 VDD.t482 VSS 0.0983f
C2546 VDD.t328 VSS 0.108f
C2547 VDD.n73 VSS 0.0506f
C2548 VDD.t139 VSS 0.00816f
C2549 VDD.t464 VSS 0.00335f
C2550 VDD.n74 VSS 0.00335f
C2551 VDD.n75 VSS 0.00732f
C2552 VDD.t138 VSS 0.0983f
C2553 VDD.t463 VSS 0.12f
C2554 VDD.t247 VSS 0.0558f
C2555 VDD.n76 VSS 0.0506f
C2556 VDD.t240 VSS 0.00816f
C2557 VDD.t161 VSS 0.00335f
C2558 VDD.n77 VSS 0.00335f
C2559 VDD.n78 VSS 0.00732f
C2560 VDD.t239 VSS 0.0983f
C2561 VDD.t160 VSS 0.12f
C2562 VDD.t4 VSS 0.0558f
C2563 VDD.t263 VSS 0.098f
C2564 VDD.n79 VSS 0.0506f
C2565 VDD.n80 VSS 0.00242f
C2566 VDD.t496 VSS 0.0053f
C2567 VDD.t268 VSS 0.007f
C2568 VDD.n81 VSS 0.0137f
C2569 VDD.n82 VSS 0.00321f
C2570 VDD.n83 VSS 0.00166f
C2571 VDD.n84 VSS 8.38e-19
C2572 VDD.n85 VSS 0.00747f
C2573 VDD.n86 VSS 0.00204f
C2574 VDD.t256 VSS 0.00696f
C2575 VDD.t495 VSS 0.00531f
C2576 VDD.n87 VSS 0.0137f
C2577 VDD.n88 VSS 0.00257f
C2578 VDD.n89 VSS 0.00218f
C2579 VDD.n90 VSS 8.38e-19
C2580 VDD.n91 VSS 0.0264f
C2581 VDD.n92 VSS 8.06e-19
C2582 VDD.t494 VSS 0.0053f
C2583 VDD.t253 VSS 0.00661f
C2584 VDD.n93 VSS 0.00677f
C2585 VDD.n94 VSS 0.00227f
C2586 VDD.n95 VSS 0.00728f
C2587 VDD.n96 VSS 0.00247f
C2588 VDD.n97 VSS 0.102f
C2589 VDD.n98 VSS 0.15f
C2590 VDD.n99 VSS 0.00204f
C2591 VDD.t259 VSS 0.00696f
C2592 VDD.t493 VSS 0.00531f
C2593 VDD.n100 VSS 0.0137f
C2594 VDD.n101 VSS 0.00267f
C2595 VDD.n102 VSS 0.0021f
C2596 VDD.n103 VSS 8.38e-19
C2597 VDD.n104 VSS 0.0264f
C2598 VDD.t497 VSS 0.00542f
C2599 VDD.t265 VSS 0.00686f
C2600 VDD.n105 VSS 0.0137f
C2601 VDD.n106 VSS 0.00499f
C2602 VDD.n107 VSS 0.0346f
C2603 VDD.n108 VSS 0.166f
C2604 VDD.t492 VSS 0.0053f
C2605 VDD.t262 VSS 0.007f
C2606 VDD.n109 VSS 0.0137f
C2607 VDD.n110 VSS 0.0698f
C2608 VDD.n111 VSS 7.92e-19
C2609 VDD.n112 VSS 0.00655f
C2610 VDD.t264 VSS 0.00762f
C2611 VDD.n113 VSS 0.0189f
C2612 VDD.n114 VSS 0.0465f
C2613 VDD.n115 VSS 0.0464f
C2614 VDD.n116 VSS 0.0477f
C2615 VDD.n117 VSS 0.0253f
C2616 VDD.n118 VSS 0.0464f
C2617 VDD.n119 VSS 0.0475f
C2618 VDD.n120 VSS 0.0282f
C2619 VDD.n121 VSS 0.0404f
C2620 VDD.n122 VSS 0.0376f
C2621 VDD.n123 VSS 0.0282f
C2622 VDD.n124 VSS 0.0769f
C2623 VDD.n125 VSS 0.0874f
C2624 VDD.t185 VSS 0.106f
C2625 VDD.t32 VSS 0.0983f
C2626 VDD.n126 VSS 0.0506f
C2627 VDD.n127 VSS 0.0282f
C2628 VDD.n128 VSS 0.0376f
C2629 VDD.n129 VSS 0.0404f
C2630 VDD.t462 VSS 0.00816f
C2631 VDD.n130 VSS 0.0376f
C2632 VDD.n131 VSS 0.0282f
C2633 VDD.n132 VSS 0.0506f
C2634 VDD.t461 VSS 0.0983f
C2635 VDD.t135 VSS 0.108f
C2636 VDD.t220 VSS 0.12f
C2637 VDD.t322 VSS 0.0983f
C2638 VDD.n133 VSS 0.0506f
C2639 VDD.n134 VSS 0.0282f
C2640 VDD.n135 VSS 0.0356f
C2641 VDD.n136 VSS 0.0333f
C2642 VDD.n137 VSS 0.0253f
C2643 VDD.n138 VSS 0.0506f
C2644 VDD.t436 VSS 0.0558f
C2645 VDD.n139 VSS 0.0757f
C2646 VDD.n140 VSS 0.0256f
C2647 VDD.n141 VSS 0.00815f
C2648 VDD.t70 VSS 0.0857f
C2649 VDD.n142 VSS 0.0436f
C2650 VDD.t327 VSS 0.00816f
C2651 VDD.n143 VSS 0.00815f
C2652 VDD.t326 VSS 0.0782f
C2653 VDD.t106 VSS 0.0857f
C2654 VDD.n144 VSS 0.0436f
C2655 VDD.t49 VSS 0.00816f
C2656 VDD.t417 VSS 0.00335f
C2657 VDD.n145 VSS 0.00335f
C2658 VDD.n146 VSS 0.00732f
C2659 VDD.n147 VSS 0.0436f
C2660 VDD.t156 VSS 0.00816f
C2661 VDD.t63 VSS 0.00335f
C2662 VDD.n148 VSS 0.00335f
C2663 VDD.n149 VSS 0.00732f
C2664 VDD.t155 VSS 0.0782f
C2665 VDD.t62 VSS 0.0955f
C2666 VDD.t169 VSS 0.0444f
C2667 VDD.t48 VSS 0.0713f
C2668 VDD.t54 VSS 0.0444f
C2669 VDD.t416 VSS 0.034f
C2670 VDD.n150 VSS 0.281f
C2671 VDD.t266 VSS 0.0897f
C2672 VDD.n151 VSS 0.0436f
C2673 VDD.t267 VSS 0.00874f
C2674 VDD.n152 VSS 0.0628f
C2675 VDD.n153 VSS 0.0464f
C2676 VDD.n154 VSS 0.0477f
C2677 VDD.n155 VSS 0.0253f
C2678 VDD.n156 VSS 0.0464f
C2679 VDD.n157 VSS 0.0475f
C2680 VDD.n158 VSS 0.0282f
C2681 VDD.n159 VSS 0.0404f
C2682 VDD.n160 VSS 0.0376f
C2683 VDD.n161 VSS 0.0282f
C2684 VDD.n162 VSS 0.0722f
C2685 VDD.n163 VSS 0.0576f
C2686 VDD.n164 VSS 0.0414f
C2687 VDD.t205 VSS 0.106f
C2688 VDD.t372 VSS 0.0983f
C2689 VDD.n165 VSS 0.0506f
C2690 VDD.n166 VSS 0.0282f
C2691 VDD.n167 VSS 0.0376f
C2692 VDD.n168 VSS 0.0404f
C2693 VDD.t419 VSS 0.00816f
C2694 VDD.n169 VSS 0.0376f
C2695 VDD.n170 VSS 0.0282f
C2696 VDD.n171 VSS 0.0506f
C2697 VDD.t418 VSS 0.0983f
C2698 VDD.t46 VSS 0.108f
C2699 VDD.t208 VSS 0.12f
C2700 VDD.t271 VSS 0.0983f
C2701 VDD.n172 VSS 0.0506f
C2702 VDD.n173 VSS 0.0282f
C2703 VDD.n174 VSS 0.0402f
C2704 VDD.n175 VSS 0.154f
C2705 VDD.n176 VSS 0.0611f
C2706 VDD.n177 VSS 0.0357f
C2707 VDD.n178 VSS 0.0506f
C2708 VDD.t260 VSS 0.0558f
C2709 VDD.n179 VSS 0.0757f
C2710 VDD.n180 VSS 0.0557f
C2711 VDD.n181 VSS 0.0947f
C2712 VDD.n182 VSS 0.07f
C2713 VDD.t297 VSS 0.106f
C2714 VDD.t320 VSS 0.0983f
C2715 VDD.n183 VSS 0.0506f
C2716 VDD.n184 VSS 0.042f
C2717 VDD.n185 VSS 0.0656f
C2718 VDD.n186 VSS 0.072f
C2719 VDD.t101 VSS 0.00816f
C2720 VDD.n187 VSS 0.0656f
C2721 VDD.n188 VSS 0.042f
C2722 VDD.n189 VSS 0.0506f
C2723 VDD.t100 VSS 0.0983f
C2724 VDD.t275 VSS 0.108f
C2725 VDD.t300 VSS 0.12f
C2726 VDD.t324 VSS 0.0983f
C2727 VDD.n190 VSS 0.0506f
C2728 VDD.n191 VSS 0.042f
C2729 VDD.n192 VSS 0.0612f
C2730 VDD.n193 VSS 0.0611f
C2731 VDD.t189 VSS 0.00816f
C2732 VDD.n194 VSS 0.052f
C2733 VDD.n195 VSS 0.0357f
C2734 VDD.n196 VSS 0.0506f
C2735 VDD.t188 VSS 0.0558f
C2736 VDD.n197 VSS 0.0757f
C2737 VDD.t21 VSS 0.00812f
C2738 VDD.n198 VSS 0.00815f
C2739 VDD.t15 VSS 0.0857f
C2740 VDD.n199 VSS 0.0436f
C2741 VDD.t45 VSS 0.00816f
C2742 VDD.n200 VSS 0.00815f
C2743 VDD.t44 VSS 0.0782f
C2744 VDD.t487 VSS 0.0857f
C2745 VDD.n201 VSS 0.0436f
C2746 VDD.t31 VSS 0.00816f
C2747 VDD.t39 VSS 0.00335f
C2748 VDD.n202 VSS 0.00335f
C2749 VDD.n203 VSS 0.00732f
C2750 VDD.n204 VSS 0.0436f
C2751 VDD.t396 VSS 0.00816f
C2752 VDD.t19 VSS 0.00335f
C2753 VDD.n205 VSS 0.00335f
C2754 VDD.n206 VSS 0.00732f
C2755 VDD.t395 VSS 0.0782f
C2756 VDD.t18 VSS 0.0955f
C2757 VDD.t73 VSS 0.0444f
C2758 VDD.t30 VSS 0.0713f
C2759 VDD.t250 VSS 0.0444f
C2760 VDD.t38 VSS 0.034f
C2761 VDD.n207 VSS 0.281f
C2762 VDD.t254 VSS 0.0897f
C2763 VDD.n208 VSS 0.0436f
C2764 VDD.t255 VSS 0.00874f
C2765 VDD.n209 VSS 0.0628f
C2766 VDD.n210 VSS 0.0464f
C2767 VDD.n211 VSS 0.0477f
C2768 VDD.n212 VSS 0.0253f
C2769 VDD.n213 VSS 0.0464f
C2770 VDD.n214 VSS 0.0475f
C2771 VDD.n215 VSS 0.0282f
C2772 VDD.n216 VSS 0.0404f
C2773 VDD.n217 VSS 0.0376f
C2774 VDD.n218 VSS 0.0282f
C2775 VDD.n219 VSS 0.0704f
C2776 VDD.n220 VSS 0.00815f
C2777 VDD.t467 VSS 0.106f
C2778 VDD.n221 VSS 0.0506f
C2779 VDD.t337 VSS 0.00816f
C2780 VDD.n222 VSS 0.00815f
C2781 VDD.t336 VSS 0.0983f
C2782 VDD.t484 VSS 0.108f
C2783 VDD.n223 VSS 0.0506f
C2784 VDD.t37 VSS 0.00816f
C2785 VDD.n224 VSS 0.00815f
C2786 VDD.t36 VSS 0.0983f
C2787 VDD.t27 VSS 0.108f
C2788 VDD.n225 VSS 0.0506f
C2789 VDD.t164 VSS 0.00816f
C2790 VDD.t466 VSS 0.00335f
C2791 VDD.n226 VSS 0.00335f
C2792 VDD.n227 VSS 0.00732f
C2793 VDD.t163 VSS 0.0983f
C2794 VDD.t465 VSS 0.12f
C2795 VDD.t78 VSS 0.0558f
C2796 VDD.n228 VSS 0.0506f
C2797 VDD.t258 VSS 0.00816f
C2798 VDD.t257 VSS 0.0558f
C2799 VDD.t76 VSS 0.0721f
C2800 VDD.n229 VSS 0.0757f
C2801 VDD.t77 VSS 0.00812f
C2802 VDD.n230 VSS 0.00828f
C2803 VDD.n232 VSS 0.00815f
C2804 VDD.n233 VSS 0.0401f
C2805 VDD.t490 VSS 0.078f
C2806 VDD.t491 VSS 0.00812f
C2807 VDD.n234 VSS 0.0375f
C2808 VDD.t43 VSS 0.00812f
C2809 VDD.n235 VSS 0.0336f
C2810 VDD.t42 VSS 0.0719f
C2811 VDD.t117 VSS 0.0558f
C2812 VDD.t383 VSS 0.00335f
C2813 VDD.n236 VSS 0.00335f
C2814 VDD.n237 VSS 0.00732f
C2815 VDD.t475 VSS 0.00816f
C2816 VDD.n238 VSS 0.00815f
C2817 VDD.n239 VSS 0.0442f
C2818 VDD.t397 VSS 0.108f
C2819 VDD.n240 VSS 0.00815f
C2820 VDD.t394 VSS 0.00816f
C2821 VDD.n241 VSS 0.00815f
C2822 VDD.n242 VSS 0.00815f
C2823 VDD.t408 VSS 0.106f
C2824 VDD.n243 VSS 0.0506f
C2825 VDD.t113 VSS 0.00816f
C2826 VDD.n244 VSS 0.00815f
C2827 VDD.t112 VSS 0.0983f
C2828 VDD.t400 VSS 0.108f
C2829 VDD.n245 VSS 0.0506f
C2830 VDD.t312 VSS 0.00816f
C2831 VDD.t97 VSS 0.00335f
C2832 VDD.n246 VSS 0.00335f
C2833 VDD.n247 VSS 0.00732f
C2834 VDD.t311 VSS 0.0983f
C2835 VDD.t96 VSS 0.12f
C2836 VDD.t51 VSS 0.0558f
C2837 VDD.n248 VSS 0.0506f
C2838 VDD.t236 VSS 0.00816f
C2839 VDD.t412 VSS 0.00335f
C2840 VDD.n249 VSS 0.00335f
C2841 VDD.n250 VSS 0.00732f
C2842 VDD.t235 VSS 0.0983f
C2843 VDD.t411 VSS 0.12f
C2844 VDD.t114 VSS 0.0558f
C2845 VDD.t282 VSS 0.098f
C2846 VDD.n251 VSS 0.0506f
C2847 VDD.t283 VSS 0.00874f
C2848 VDD.n252 VSS 0.0628f
C2849 VDD.n253 VSS 0.0464f
C2850 VDD.n254 VSS 0.0477f
C2851 VDD.n255 VSS 0.0253f
C2852 VDD.n256 VSS 0.0464f
C2853 VDD.n257 VSS 0.0475f
C2854 VDD.n258 VSS 0.0282f
C2855 VDD.n259 VSS 0.0404f
C2856 VDD.n260 VSS 0.0376f
C2857 VDD.n261 VSS 0.0282f
C2858 VDD.n262 VSS 0.0707f
C2859 VDD.t121 VSS 0.00812f
C2860 VDD.t238 VSS 0.00816f
C2861 VDD.n263 VSS 0.0476f
C2862 VDD.t120 VSS 0.0719f
C2863 VDD.t215 VSS 0.0558f
C2864 VDD.t368 VSS 0.00335f
C2865 VDD.n264 VSS 0.00335f
C2866 VDD.n265 VSS 0.00732f
C2867 VDD.t314 VSS 0.00816f
C2868 VDD.n266 VSS 0.00815f
C2869 VDD.n267 VSS 0.0445f
C2870 VDD.t129 VSS 0.108f
C2871 VDD.n268 VSS 0.00815f
C2872 VDD.t287 VSS 0.00816f
C2873 VDD.n269 VSS 0.00815f
C2874 VDD.n270 VSS 0.00815f
C2875 VDD.t425 VSS 0.106f
C2876 VDD.n271 VSS 0.0506f
C2877 VDD.t285 VSS 0.00816f
C2878 VDD.n272 VSS 0.00815f
C2879 VDD.t284 VSS 0.0983f
C2880 VDD.t132 VSS 0.108f
C2881 VDD.n273 VSS 0.0506f
C2882 VDD.t234 VSS 0.00816f
C2883 VDD.t479 VSS 0.00335f
C2884 VDD.n274 VSS 0.00335f
C2885 VDD.n275 VSS 0.00732f
C2886 VDD.t233 VSS 0.0983f
C2887 VDD.t478 VSS 0.12f
C2888 VDD.t387 VSS 0.0558f
C2889 VDD.n276 VSS 0.0506f
C2890 VDD.t343 VSS 0.00816f
C2891 VDD.t431 VSS 0.00335f
C2892 VDD.n277 VSS 0.00335f
C2893 VDD.n278 VSS 0.00732f
C2894 VDD.t342 VSS 0.0983f
C2895 VDD.t430 VSS 0.12f
C2896 VDD.t202 VSS 0.0558f
C2897 VDD.t374 VSS 0.098f
C2898 VDD.n279 VSS 0.0506f
C2899 VDD.t375 VSS 0.00874f
C2900 VDD.n280 VSS 0.0628f
C2901 VDD.n281 VSS 0.0464f
C2902 VDD.n282 VSS 0.0477f
C2903 VDD.n283 VSS 0.0253f
C2904 VDD.n284 VSS 0.0464f
C2905 VDD.n285 VSS 0.0475f
C2906 VDD.n286 VSS 0.0282f
C2907 VDD.n287 VSS 0.0404f
C2908 VDD.n288 VSS 0.0376f
C2909 VDD.n289 VSS 0.0282f
C2910 VDD.n290 VSS 0.0707f
C2911 VDD.t198 VSS 0.00812f
C2912 VDD.t471 VSS 0.00816f
C2913 VDD.n291 VSS 0.0472f
C2914 VDD.t197 VSS 0.0719f
C2915 VDD.t212 VSS 0.0558f
C2916 VDD.t128 VSS 0.00335f
C2917 VDD.n292 VSS 0.00335f
C2918 VDD.n293 VSS 0.00732f
C2919 VDD.t421 VSS 0.00816f
C2920 VDD.n294 VSS 0.00815f
C2921 VDD.n295 VSS 0.0442f
C2922 VDD.t225 VSS 0.108f
C2923 VDD.n296 VSS 0.00815f
C2924 VDD.t82 VSS 0.00816f
C2925 VDD.n297 VSS 0.00815f
C2926 VDD.n298 VSS 0.00815f
C2927 VDD.t360 VSS 0.106f
C2928 VDD.n299 VSS 0.0506f
C2929 VDD.t447 VSS 0.00816f
C2930 VDD.n300 VSS 0.00815f
C2931 VDD.t446 VSS 0.0983f
C2932 VDD.t222 VSS 0.108f
C2933 VDD.n301 VSS 0.0506f
C2934 VDD.t89 VSS 0.00816f
C2935 VDD.t307 VSS 0.00335f
C2936 VDD.n302 VSS 0.00335f
C2937 VDD.n303 VSS 0.00732f
C2938 VDD.t88 VSS 0.0983f
C2939 VDD.t306 VSS 0.12f
C2940 VDD.t57 VSS 0.0558f
C2941 VDD.n304 VSS 0.0506f
C2942 VDD.t84 VSS 0.00816f
C2943 VDD.t350 VSS 0.00335f
C2944 VDD.n305 VSS 0.00335f
C2945 VDD.n306 VSS 0.00732f
C2946 VDD.t83 VSS 0.0983f
C2947 VDD.t349 VSS 0.12f
C2948 VDD.t194 VSS 0.0558f
C2949 VDD.t472 VSS 0.098f
C2950 VDD.n307 VSS 0.0506f
C2951 VDD.t473 VSS 0.00874f
C2952 VDD.n308 VSS 0.0628f
C2953 VDD.n309 VSS 0.0464f
C2954 VDD.n310 VSS 0.0477f
C2955 VDD.n311 VSS 0.0253f
C2956 VDD.n312 VSS 0.0464f
C2957 VDD.n313 VSS 0.0475f
C2958 VDD.n314 VSS 0.0282f
C2959 VDD.n315 VSS 0.0404f
C2960 VDD.n316 VSS 0.0376f
C2961 VDD.n317 VSS 0.0282f
C2962 VDD.n318 VSS 0.0959f
C2963 VDD.t211 VSS 0.00812f
C2964 VDD.t1 VSS 0.00816f
C2965 VDD.n319 VSS 0.048f
C2966 VDD.t210 VSS 0.0719f
C2967 VDD.t122 VSS 0.0558f
C2968 VDD.t319 VSS 0.00335f
C2969 VDD.n320 VSS 0.00335f
C2970 VDD.n321 VSS 0.00732f
C2971 VDD.t35 VSS 0.00816f
C2972 VDD.n322 VSS 0.00815f
C2973 VDD.n323 VSS 0.0449f
C2974 VDD.t90 VSS 0.108f
C2975 VDD.n324 VSS 0.00815f
C2976 VDD.t335 VSS 0.00816f
C2977 VDD.n325 VSS 0.00815f
C2978 VDD.n326 VSS 0.00815f
C2979 VDD.t145 VSS 0.106f
C2980 VDD.n327 VSS 0.0506f
C2981 VDD.t166 VSS 0.00816f
C2982 VDD.n328 VSS 0.00815f
C2983 VDD.t165 VSS 0.0983f
C2984 VDD.t93 VSS 0.108f
C2985 VDD.n329 VSS 0.0506f
C2986 VDD.t296 VSS 0.00816f
C2987 VDD.t379 VSS 0.00335f
C2988 VDD.n330 VSS 0.00335f
C2989 VDD.n331 VSS 0.00732f
C2990 VDD.t295 VSS 0.0983f
C2991 VDD.t378 VSS 0.12f
C2992 VDD.t244 VSS 0.0558f
C2993 VDD.n332 VSS 0.0506f
C2994 VDD.t105 VSS 0.00816f
C2995 VDD.t151 VSS 0.00335f
C2996 VDD.n333 VSS 0.00335f
C2997 VDD.n334 VSS 0.00732f
C2998 VDD.t104 VSS 0.0983f
C2999 VDD.t150 VSS 0.12f
C3000 VDD.t199 VSS 0.0558f
C3001 VDD.t2 VSS 0.098f
C3002 VDD.n335 VSS 0.0506f
C3003 VDD.t3 VSS 0.00874f
C3004 VDD.n336 VSS 0.0628f
C3005 VDD.n337 VSS 0.0464f
C3006 VDD.n338 VSS 0.0477f
C3007 VDD.n339 VSS 0.0253f
C3008 VDD.n340 VSS 0.0464f
C3009 VDD.n341 VSS 0.0475f
C3010 VDD.n342 VSS 0.0282f
C3011 VDD.n343 VSS 0.0404f
C3012 VDD.n344 VSS 0.0376f
C3013 VDD.n345 VSS 0.0282f
C3014 VDD.n346 VSS 0.0962f
C3015 VDD.n347 VSS 0.111f
C3016 VDD.t315 VSS 0.106f
C3017 VDD.t334 VSS 0.0983f
C3018 VDD.n348 VSS 0.0506f
C3019 VDD.n349 VSS 0.0301f
C3020 VDD.n350 VSS 0.0415f
C3021 VDD.n351 VSS 0.0449f
C3022 VDD.t377 VSS 0.00816f
C3023 VDD.n352 VSS 0.0415f
C3024 VDD.n353 VSS 0.0301f
C3025 VDD.n354 VSS 0.0506f
C3026 VDD.t376 VSS 0.0983f
C3027 VDD.t292 VSS 0.108f
C3028 VDD.t318 VSS 0.12f
C3029 VDD.t34 VSS 0.0983f
C3030 VDD.n355 VSS 0.0506f
C3031 VDD.n356 VSS 0.0301f
C3032 VDD.n357 VSS 0.0392f
C3033 VDD.n358 VSS 0.0372f
C3034 VDD.n359 VSS 0.0268f
C3035 VDD.n360 VSS 0.0506f
C3036 VDD.t0 VSS 0.0558f
C3037 VDD.n361 VSS 0.0757f
C3038 VDD.n362 VSS 0.0456f
C3039 VDD.n363 VSS 0.0508f
C3040 VDD.n364 VSS 0.0454f
C3041 VDD.t191 VSS 0.106f
C3042 VDD.t81 VSS 0.0983f
C3043 VDD.n365 VSS 0.0506f
C3044 VDD.n366 VSS 0.0298f
C3045 VDD.n367 VSS 0.0409f
C3046 VDD.n368 VSS 0.0442f
C3047 VDD.t305 VSS 0.00816f
C3048 VDD.n369 VSS 0.0409f
C3049 VDD.n370 VSS 0.0298f
C3050 VDD.n371 VSS 0.0506f
C3051 VDD.t304 VSS 0.0983f
C3052 VDD.t85 VSS 0.108f
C3053 VDD.t127 VSS 0.12f
C3054 VDD.t420 VSS 0.0983f
C3055 VDD.n372 VSS 0.0506f
C3056 VDD.n373 VSS 0.0298f
C3057 VDD.n374 VSS 0.0386f
C3058 VDD.n375 VSS 0.0366f
C3059 VDD.n376 VSS 0.0265f
C3060 VDD.n377 VSS 0.0506f
C3061 VDD.t470 VSS 0.0558f
C3062 VDD.n378 VSS 0.0757f
C3063 VDD.n379 VSS 0.0437f
C3064 VDD.n380 VSS 0.0716f
C3065 VDD.n381 VSS 0.0435f
C3066 VDD.t364 VSS 0.106f
C3067 VDD.t286 VSS 0.0983f
C3068 VDD.n382 VSS 0.0506f
C3069 VDD.n383 VSS 0.03f
C3070 VDD.n384 VSS 0.0412f
C3071 VDD.n385 VSS 0.0445f
C3072 VDD.t477 VSS 0.00816f
C3073 VDD.n386 VSS 0.0412f
C3074 VDD.n387 VSS 0.03f
C3075 VDD.n388 VSS 0.0506f
C3076 VDD.t476 VSS 0.0983f
C3077 VDD.t230 VSS 0.108f
C3078 VDD.t367 VSS 0.12f
C3079 VDD.t313 VSS 0.0983f
C3080 VDD.n389 VSS 0.0506f
C3081 VDD.n390 VSS 0.03f
C3082 VDD.n391 VSS 0.0389f
C3083 VDD.n392 VSS 0.0314f
C3084 VDD.t429 VSS 0.00779f
C3085 VDD.t303 VSS 0.017f
C3086 VDD.n393 VSS 0.0978f
C3087 VDD.t348 VSS 0.00816f
C3088 VDD.t41 VSS 0.00335f
C3089 VDD.n394 VSS 0.00335f
C3090 VDD.n395 VSS 0.00732f
C3091 VDD.t357 VSS 0.00816f
C3092 VDD.n396 VSS 0.00815f
C3093 VDD.n397 VSS 0.0652f
C3094 VDD.t290 VSS 0.0959f
C3095 VDD.t356 VSS 0.0789f
C3096 VDD.t344 VSS 0.0394f
C3097 VDD.t449 VSS 0.00812f
C3098 VDD.t289 VSS 0.00812f
C3099 VDD.n398 VSS 0.0548f
C3100 VDD.t448 VSS 0.0537f
C3101 VDD.t452 VSS 0.104f
C3102 VDD.t453 VSS 0.017f
C3103 VDD.t457 VSS 0.0316f
C3104 VDD.n399 VSS 0.115f
C3105 VDD.t422 VSS 0.0661f
C3106 VDD.t451 VSS 0.00812f
C3107 VDD.t415 VSS 0.199f
C3108 VDD.t450 VSS 0.0961f
C3109 VDD.n400 VSS 0.0633f
C3110 VDD.n401 VSS 0.101f
C3111 VDD.n402 VSS 0.0959f
C3112 VDD.n403 VSS 0.0766f
C3113 VDD.t456 VSS 0.21f
C3114 VDD.n404 VSS 0.119f
C3115 VDD.n405 VSS 0.0609f
C3116 VDD.n406 VSS 0.0401f
C3117 VDD.n407 VSS 0.115f
C3118 VDD.t288 VSS 0.0571f
C3119 VDD.n408 VSS 0.0759f
C3120 VDD.n409 VSS 0.0739f
C3121 VDD.t291 VSS 0.00812f
C3122 VDD.n410 VSS 0.0554f
C3123 VDD.n411 VSS 0.0791f
C3124 VDD.n412 VSS 0.0688f
C3125 VDD.n413 VSS 0.0856f
C3126 VDD.n414 VSS 0.0868f
C3127 VDD.t40 VSS 0.0789f
C3128 VDD.t347 VSS 0.0789f
C3129 VDD.t152 VSS 0.0594f
C3130 VDD.n415 VSS 0.029f
C3131 VDD.n416 VSS 0.104f
C3132 VDD.t302 VSS 0.0809f
C3133 VDD.t428 VSS 0.0972f
C3134 VDD.n417 VSS 0.0844f
C3135 VDD.n418 VSS 0.0601f
C3136 VDD.n419 VSS 0.0704f
C3137 VDD.t459 VSS 0.00812f
C3138 VDD.n420 VSS 0.0265f
C3139 VDD.t458 VSS 0.0768f
C3140 VDD.n421 VSS 0.087f
C3141 VDD.t190 VSS 0.0911f
C3142 VDD.t380 VSS 0.0915f
C3143 VDD.n422 VSS 0.0574f
C3144 VDD.t381 VSS 0.0195f
C3145 VDD.t126 VSS 0.00812f
C3146 VDD.n423 VSS 0.0265f
C3147 VDD.t125 VSS 0.0768f
C3148 VDD.n424 VSS 0.087f
C3149 VDD.t243 VSS 0.0911f
C3150 VDD.t140 VSS 0.0915f
C3151 VDD.n425 VSS 0.0574f
C3152 VDD.t141 VSS 0.0195f
C3153 VDD.t359 VSS 0.00816f
C3154 VDD.n426 VSS 0.00815f
C3155 VDD.n427 VSS 0.0401f
C3156 VDD.t480 VSS 0.0959f
C3157 VDD.t358 VSS 0.0789f
C3158 VDD.t405 VSS 0.0394f
C3159 VDD.t481 VSS 0.00812f
C3160 VDD.n428 VSS 0.0287f
C3161 VDD.n429 VSS 0.0791f
C3162 VDD.n430 VSS 0.0574f
C3163 VDD.n431 VSS 0.254f
C3164 VDD.n432 VSS 0.47f
C3165 VDD.n433 VSS 0.168f
C3166 VDD.n434 VSS 0.283f
C3167 VDD.n435 VSS 0.262f
C3168 VDD.n436 VSS 0.139f
C3169 VDD.n437 VSS 0.607f
C3170 VDD.n438 VSS 0.707f
C3171 VDD.n439 VSS 0.125f
C3172 VDD.n440 VSS 0.0267f
C3173 VDD.n441 VSS 0.0506f
C3174 VDD.t237 VSS 0.0558f
C3175 VDD.n442 VSS 0.0757f
C3176 VDD.n443 VSS 0.0453f
C3177 VDD.n444 VSS 0.0725f
C3178 VDD.n445 VSS 0.0432f
C3179 VDD.t384 VSS 0.106f
C3180 VDD.t393 VSS 0.0983f
C3181 VDD.n446 VSS 0.0506f
C3182 VDD.n447 VSS 0.0298f
C3183 VDD.n448 VSS 0.0409f
C3184 VDD.n449 VSS 0.0442f
C3185 VDD.t99 VSS 0.00816f
C3186 VDD.n450 VSS 0.0409f
C3187 VDD.n451 VSS 0.0298f
C3188 VDD.n452 VSS 0.0506f
C3189 VDD.t98 VSS 0.0983f
C3190 VDD.t308 VSS 0.108f
C3191 VDD.t382 VSS 0.12f
C3192 VDD.t474 VSS 0.0983f
C3193 VDD.n453 VSS 0.0506f
C3194 VDD.n454 VSS 0.0298f
C3195 VDD.n455 VSS 0.0386f
C3196 VDD.n456 VSS 0.0366f
C3197 VDD.t281 VSS 0.00816f
C3198 VDD.n457 VSS 0.0418f
C3199 VDD.n458 VSS 0.0265f
C3200 VDD.n459 VSS 0.0506f
C3201 VDD.t280 VSS 0.0558f
C3202 VDD.n460 VSS 0.0713f
C3203 VDD.n461 VSS 0.0674f
C3204 VDD.n462 VSS 0.0413f
C3205 VDD.n463 VSS 0.074f
C3206 VDD.t353 VSS 0.0638f
C3207 VDD.t148 VSS 0.098f
C3208 VDD.n464 VSS 0.0506f
C3209 VDD.n465 VSS 0.0285f
C3210 VDD.t149 VSS 0.00829f
C3211 VDD.n466 VSS 0.0453f
C3212 VDD.n467 VSS 0.0872f
C3213 VDD.t433 VSS 0.0194f
C3214 VDD.t278 VSS 0.1f
C3215 VDD.n468 VSS 0.0694f
C3216 VDD.t279 VSS 0.00812f
C3217 VDD.t424 VSS 0.00335f
C3218 VDD.n469 VSS 0.00335f
C3219 VDD.n470 VSS 0.00732f
C3220 VDD.n471 VSS 0.00815f
C3221 VDD.n472 VSS 0.0611f
C3222 VDD.t439 VSS 0.00812f
C3223 VDD.t363 VSS 0.00816f
C3224 VDD.t352 VSS 0.00816f
C3225 VDD.n473 VSS 0.0751f
C3226 VDD.n474 VSS 0.0344f
C3227 VDD.t351 VSS 0.196f
C3228 VDD.n475 VSS 0.101f
C3229 VDD.t142 VSS 0.112f
C3230 VDD.t423 VSS 0.154f
C3231 VDD.t242 VSS 0.00812f
C3232 VDD.n476 VSS 0.0202f
C3233 VDD.n477 VSS 0.00414f
C3234 VDD.n478 VSS 0.0622f
C3235 VDD.t241 VSS 0.0723f
C3236 VDD.n479 VSS 0.0848f
C3237 VDD.t371 VSS 0.0681f
C3238 VDD.t432 VSS 0.0262f
C3239 VDD.t438 VSS 0.108f
C3240 VDD.n481 VSS 0.0291f
C3241 VDD.n482 VSS 0.102f
C3242 VDD.n483 VSS 0.0606f
C3243 VDD.n484 VSS 0.0288f
C3244 VDD.n485 VSS 0.0156f
C3245 VDD.n486 VSS 0.0848f
C3246 VDD.n487 VSS 0.0366f
C3247 VDD.n488 VSS 0.0406f
C3248 VDD.n489 VSS 0.0278f
C3249 VDD.n490 VSS 0.00706f
C3250 VDD.n491 VSS 0.00118f
C3251 VDD.n492 VSS 0.354f
C3252 VDD.n493 VSS 0.483f
C3253 VDD.n494 VSS 0.0775f
C3254 VDD.n495 VSS 0.0357f
C3255 VDD.n496 VSS 0.0611f
C3256 VDD.n497 VSS 0.0612f
C3257 VDD.n498 VSS 0.042f
C3258 VDD.n499 VSS 0.072f
C3259 VDD.n500 VSS 0.0656f
C3260 VDD.n501 VSS 0.042f
C3261 VDD.n502 VSS 0.072f
C3262 VDD.n503 VSS 0.0656f
C3263 VDD.n504 VSS 0.042f
C3264 VDD.n505 VSS 0.07f
C3265 VDD.n506 VSS 0.0736f
C3266 VDD.n507 VSS 0.0478f
.ends

