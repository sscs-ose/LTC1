magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2961 -2038 2961 2038
<< metal2 >>
rect -961 28 961 38
rect -961 -28 -951 28
rect -895 -28 -809 28
rect -753 -28 -667 28
rect -611 -28 -525 28
rect -469 -28 -383 28
rect -327 -28 -241 28
rect -185 -28 -99 28
rect -43 -28 43 28
rect 99 -28 185 28
rect 241 -28 327 28
rect 383 -28 469 28
rect 525 -28 611 28
rect 667 -28 753 28
rect 809 -28 895 28
rect 951 -28 961 28
rect -961 -38 961 -28
<< via2 >>
rect -951 -28 -895 28
rect -809 -28 -753 28
rect -667 -28 -611 28
rect -525 -28 -469 28
rect -383 -28 -327 28
rect -241 -28 -185 28
rect -99 -28 -43 28
rect 43 -28 99 28
rect 185 -28 241 28
rect 327 -28 383 28
rect 469 -28 525 28
rect 611 -28 667 28
rect 753 -28 809 28
rect 895 -28 951 28
<< metal3 >>
rect -961 28 961 38
rect -961 -28 -951 28
rect -895 -28 -809 28
rect -753 -28 -667 28
rect -611 -28 -525 28
rect -469 -28 -383 28
rect -327 -28 -241 28
rect -185 -28 -99 28
rect -43 -28 43 28
rect 99 -28 185 28
rect 241 -28 327 28
rect 383 -28 469 28
rect 525 -28 611 28
rect 667 -28 753 28
rect 809 -28 895 28
rect 951 -28 961 28
rect -961 -38 961 -28
<< end >>
