* NGSPICE file created from Current_Mirror_Top_flat.ext - technology: gf180mcuC

.subckt Current_Mirror_Top_flat VDD G_source_up G_source_dn VSS G_sink_up G_sink_dn
+ SD0_1 G1_2 G1_1 SD1_1 G2_1 SD2_1 ITAIL
X0 VSS G2_1.t24 G2_1.t25 VSS.t16 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X1 G2_1 ITAIL.t38 ITAIL.t39 VSS.t45 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X2 VDD G1_2.t26 G1_2.t27 VDD.t5 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X3 G2_1 ITAIL.t36 ITAIL.t37 VSS.t6 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X4 G1_2 G1_2.t42 VDD.t86 VDD.t85 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X5 SD0_1 G_sink_dn.t24 VSS.t96 VSS.t95 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X6 ITAIL ITAIL.t34 G2_1.t57 VSS.t31 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X7 SD2_1 G2_1.t60 VSS.t77 VSS.t53 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X8 G_sink_dn G_sink_dn.t21 VSS.t89 VSS.t88 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X9 G1_1 G1_1.t38 G1_2.t51 VDD.t72 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X10 G1_2 G1_2.t44 VDD.t84 VDD.t83 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X11 VDD G1_2.t24 G1_2.t25 VDD.t80 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X12 ITAIL ITAIL.t32 G2_1.t56 VSS.t13 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X13 G1_2 G1_1.t36 G1_1.t37 VDD.t59 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X14 G_sink_dn G_sink_up.t24 G_sink_up.t25 VSS.t93 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X15 VSS G2_1.t61 SD2_1.t18 VSS.t21 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X16 VSS G_sink_dn.t26 SD0_1.t14 VSS.t99 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X17 G_sink_up G1_1.t61 SD1_1.t9 VDD.t7 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X18 VSS G2_1.t62 SD2_1.t17 VSS.t48 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X19 VSS G2_1.t22 G2_1.t23 VSS.t62 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X20 SD2_1 G2_1.t63 VSS.t70 VSS.t24 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X21 VSS G2_1.t20 G2_1.t21 VSS.t26 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X22 G_source_dn G_source_dn.t18 G_source_up.t23 VDD.t91 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X23 G_sink_up G1_1.t62 SD1_1.t8 VDD.t8 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X24 VSS G2_1.t64 SD2_1.t15 VSS.t2 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X25 G_sink_up G_sink_up.t22 G_sink_dn.t3 VSS.t100 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X26 G2_1 ITAIL.t30 ITAIL.t31 VSS.t24 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X27 G1_1 G1_1.t34 G1_2.t57 VDD.t38 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X28 VSS G_sink_dn.t19 G_sink_dn.t20 VSS.t85 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X29 VSS G_sink_dn.t27 SD0_1.t13 VSS.t103 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X30 SD1_1 G1_2.t62 VDD.t36 VDD.t35 pfet_03v3 ad=0.104p pd=0.92u as=0.176p ps=1.68u w=0.4u l=0.5u
X31 G1_1 ITAIL.t42 SD2_1.t35 VSS.t42 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X32 SD2_1 G2_1.t65 VSS.t64 VSS.t57 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X33 G1_1 G1_1.t32 G1_2.t56 VDD.t7 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X34 VSS G2_1.t66 SD2_1.t13 VSS.t62 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X35 SD2_1 ITAIL.t43 G1_1.t58 VSS.t6 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X36 G2_1 ITAIL.t28 ITAIL.t29 VSS.t29 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X37 G2_1 G2_1.t38 VSS.t61 VSS.t11 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X38 G_source_up G_source_up.t14 VDD.t25 VDD.t24 pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X39 G_source_up G_source_up.t12 VDD.t31 VDD.t30 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X40 G_sink_dn G_sink_up.t20 G_sink_up.t21 VSS.t111 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X41 SD1_1 G1_2.t63 VDD.t34 VDD.t33 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X42 G1_1 G1_1.t30 G1_2.t55 VDD.t8 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X43 VSS G2_1.t18 G2_1.t19 VSS.t37 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X44 SD0_1 G_sink_up.t27 G_source_dn.t7 VSS.t97 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X45 G1_2 G1_2.t40 VDD.t79 VDD.t35 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X46 G2_1 G2_1.t30 VSS.t58 VSS.t57 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X47 G1_1 ITAIL.t44 SD2_1.t34 VSS.t13 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X48 G1_2 G1_1.t28 G1_1.t29 VDD.t45 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X49 VSS G2_1.t16 G2_1.t17 VSS.t42 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X50 G_source_up G_source_dn.t16 G_source_dn.t17 VDD.t90 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X51 G2_1 ITAIL.t26 ITAIL.t27 VSS.t8 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X52 VSS G_sink_dn.t28 SD0_1.t12 VSS.t80 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X53 G_sink_dn G_sink_up.t18 G_sink_up.t19 VSS.t109 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X54 G1_2 G1_2.t32 VDD.t77 VDD.t33 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X55 G1_1 ITAIL.t45 SD2_1.t33 VSS.t31 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X56 ITAIL ITAIL.t24 G2_1.t52 VSS.t21 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X57 G1_1 G1_1.t26 G1_2.t58 VDD.t41 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X58 G_sink_up G1_1.t67 SD1_1.t7 VDD.t4 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X59 G1_1 G1_1.t24 G1_2.t5 VDD.t6 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X60 G_sink_up G_sink_up.t16 G_sink_dn.t6 VSS.t106 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X61 G2_1 G2_1.t32 VSS.t54 VSS.t53 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X62 G1_1 ITAIL.t47 SD2_1.t32 VSS.t26 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X63 G_source_dn G_sink_up.t29 SD0_1.t3 VSS.t98 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X64 VDD G1_2.t66 SD1_1.t17 VDD.t69 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X65 SD0_1 G_sink_up.t30 G_source_dn.t5 VSS.t112 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X66 SD2_1 G2_1.t70 VSS.t52 VSS.t45 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X67 SD2_1 ITAIL.t48 G1_1.t54 VSS.t53 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X68 G1_1 G1_1.t22 G1_2.t4 VDD.t5 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X69 SD1_1 G1_2.t67 VDD.t75 VDD.t67 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X70 G2_1 G2_1.t0 VSS.t51 VSS.t0 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X71 VDD G_source_up.t10 G_source_up.t11 VDD.t15 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X72 VSS G2_1.t14 G2_1.t15 VSS.t48 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X73 VDD G1_2.t22 G1_2.t23 VDD.t72 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X74 SD1_1 G1_1.t70 G_sink_up.t4 VDD.t0 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X75 G1_1 G1_1.t20 G1_2.t3 VDD.t4 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X76 G_sink_dn G_sink_up.t14 G_sink_up.t15 VSS.t88 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X77 SD2_1 G2_1.t72 VSS.t47 VSS.t29 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X78 SD1_1 G1_1.t72 G_sink_up.t3 VDD.t2 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X79 VDD G1_2.t20 G1_2.t21 VDD.t69 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X80 G1_1 ITAIL.t49 SD2_1.t31 VSS.t21 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X81 SD0_1 G_sink_dn.t29 VSS.t84 VSS.t83 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X82 G2_1 ITAIL.t22 ITAIL.t23 VSS.t4 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X83 G1_1 ITAIL.t50 SD2_1.t30 VSS.t48 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X84 G_source_up G_source_dn.t14 G_source_dn.t15 VDD.t89 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X85 G2_1 G2_1.t34 VSS.t46 VSS.t45 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X86 G_source_up G_source_dn.t12 G_source_dn.t13 VDD.t27 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X87 G_sink_dn G_sink_dn.t17 VSS.t94 VSS.t93 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X88 SD1_1 G1_1.t73 G_sink_up.t2 VDD.t1 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X89 G1_2 G1_2.t30 VDD.t68 VDD.t67 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X90 ITAIL ITAIL.t20 G2_1.t47 VSS.t16 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X91 G1_2 G1_1.t18 G1_1.t19 VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X92 G2_1 G2_1.t2 VSS.t7 VSS.t6 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X93 G1_1 ITAIL.t52 SD2_1.t29 VSS.t2 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X94 G1_2 G1_1.t16 G1_1.t17 VDD.t2 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X95 ITAIL ITAIL.t18 G2_1.t46 VSS.t2 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X96 VSS G2_1.t75 SD2_1.t10 VSS.t42 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X97 G1_1 ITAIL.t54 SD2_1.t28 VSS.t16 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X98 G_source_dn G_source_dn.t22 G_source_up.t19 VDD.t3 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X99 G_source_dn G_sink_up.t31 SD0_1.t7 VSS.t103 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X100 G1_2 G1_1.t14 G1_1.t15 VDD.t1 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X101 VSS G2_1.t12 G2_1.t13 VSS.t13 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X102 VDD G1_2.t18 G1_2.t19 VDD.t7 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X103 VSS G2_1.t76 SD2_1.t9 VSS.t37 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X104 VSS G_sink_dn.t15 G_sink_dn.t16 VSS.t90 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X105 ITAIL ITAIL.t16 G2_1.t45 VSS.t62 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X106 VDD G1_2.t16 G1_2.t17 VDD.t8 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X107 G1_2 G1_1.t12 G1_1.t13 VDD.t35 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X108 ITAIL ITAIL.t14 G2_1.t44 VSS.t26 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X109 VSS G2_1.t10 G2_1.t11 VSS.t31 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X110 SD2_1 G2_1.t77 VSS.t34 VSS.t4 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X111 SD0_1 G_sink_dn.t31 VSS.t117 VSS.t97 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X112 SD1_1 G1_1.t74 G_sink_up.t1 VDD.t85 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X113 SD2_1 ITAIL.t57 G1_1.t49 VSS.t11 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X114 SD2_1 ITAIL.t58 G1_1.t48 VSS.t8 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X115 VSS G2_1.t78 SD2_1.t7 VSS.t31 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X116 G_source_up G_source_dn.t10 G_source_dn.t11 VDD.t9 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X117 SD1_1 G1_1.t75 G_sink_up.t0 VDD.t83 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X118 G2_1 G2_1.t36 VSS.t30 VSS.t29 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X119 G2_1 ITAIL.t12 ITAIL.t13 VSS.t11 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X120 G1_2 G1_1.t10 G1_1.t11 VDD.t33 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X121 G_sink_dn G_sink_dn.t13 VSS.t110 VSS.t109 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X122 G_sink_up G1_1.t76 SD1_1.t1 VDD.t80 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X123 SD1_1 G1_2.t69 VDD.t62 VDD.t59 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X124 SD2_1 ITAIL.t59 G1_1.t47 VSS.t0 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X125 G_source_up G_source_up.t8 VDD.t14 VDD.t13 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X126 SD0_1 G_sink_up.t32 G_source_dn.t3 VSS.t95 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X127 G1_2 G1_1.t8 G1_1.t9 VDD.t85 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X128 VSS G2_1.t80 SD2_1.t6 VSS.t26 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X129 G_source_dn G_source_dn.t20 G_source_up.t17 VDD.t92 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X130 SD2_1 ITAIL.t60 G1_1.t46 VSS.t45 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X131 G_source_up G_source_up.t6 VDD.t29 VDD.t28 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X132 G2_1 ITAIL.t10 ITAIL.t11 VSS.t57 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X133 G2_1 G2_1.t4 VSS.t25 VSS.t24 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X134 VSS G_sink_dn.t11 G_sink_dn.t12 VSS.t106 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X135 G1_2 G1_1.t6 G1_1.t7 VDD.t83 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X136 ITAIL ITAIL.t8 G2_1.t41 VSS.t42 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X137 VDD G1_2.t70 SD1_1.t14 VDD.t38 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X138 G1_1 G1_1.t4 G1_2.t48 VDD.t80 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X139 G1_2 G1_2.t6 VDD.t60 VDD.t59 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X140 G_source_dn G_sink_up.t33 SD0_1.t5 VSS.t99 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X141 SD2_1 ITAIL.t62 G1_1.t45 VSS.t29 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X142 VSS G2_1.t8 G2_1.t9 VSS.t21 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X143 VDD G1_2.t14 G1_2.t15 VDD.t4 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X144 VDD G_source_up.t4 G_source_up.t5 VDD.t10 pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X145 G1_1 G1_1.t2 G1_2.t54 VDD.t69 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X146 ITAIL ITAIL.t6 G2_1.t40 VSS.t37 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X147 VSS G_sink_dn.t9 G_sink_dn.t10 VSS.t100 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X148 G_sink_up G_sink_up.t12 G_sink_dn.t0 VSS.t85 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X149 SD2_1 ITAIL.t64 G1_1.t44 VSS.t24 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X150 SD0_1 G_sink_up.t35 G_source_dn.t1 VSS.t83 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X151 VDD G1_2.t12 G1_2.t13 VDD.t38 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X152 G1_2 G1_1.t0 G1_1.t1 VDD.t67 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X153 G1_2 G1_2.t34 VDD.t54 VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X154 SD1_1 G1_2.t73 VDD.t53 VDD.t45 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X155 G2_1 ITAIL.t4 ITAIL.t5 VSS.t0 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X156 G2_1 G2_1.t28 VSS.t18 VSS.t8 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X157 SD2_1 ITAIL.t65 G1_1.t43 VSS.t57 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X158 G1_2 G1_2.t28 VDD.t52 VDD.t2 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X159 G_sink_dn G_sink_dn.t7 VSS.t113 VSS.t111 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X160 G1_1 ITAIL.t66 SD2_1.t27 VSS.t62 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X161 SD2_1 G2_1.t83 VSS.t20 VSS.t6 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X162 VSS G2_1.t84 SD2_1.t4 VSS.t16 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X163 G2_1 G2_1.t26 VSS.t5 VSS.t4 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X164 G1_1 ITAIL.t67 SD2_1.t26 VSS.t37 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X165 G1_2 G1_2.t36 VDD.t51 VDD.t1 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X166 VDD G1_2.t76 SD1_1.t12 VDD.t41 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X167 G2_1 ITAIL.t2 ITAIL.t3 VSS.t53 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X168 VDD G1_2.t77 SD1_1.t11 VDD.t6 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X169 VDD G_source_up.t2 G_source_up.t3 VDD.t21 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X170 G1_2 G1_2.t38 VDD.t46 VDD.t45 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X171 SD2_1 ITAIL.t68 G1_1.t40 VSS.t4 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X172 G_source_dn G_sink_up.t36 SD0_1.t1 VSS.t80 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X173 G_sink_up G_sink_up.t10 G_sink_dn.t23 VSS.t90 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X174 VSS G2_1.t86 SD2_1.t3 VSS.t13 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X175 SD2_1 G2_1.t87 VSS.t12 VSS.t11 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X176 VSS G2_1.t6 G2_1.t7 VSS.t2 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X177 SD2_1 G2_1.t88 VSS.t9 VSS.t8 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X178 VDD G_source_up.t0 G_source_up.t1 VDD.t18 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X179 VDD G1_2.t79 SD1_1.t10 VDD.t5 pfet_03v3 ad=0.176p pd=1.68u as=0.104p ps=0.92u w=0.4u l=0.5u
X180 ITAIL ITAIL.t0 G2_1.t49 VSS.t48 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X181 G_source_dn G_source_dn.t8 G_source_up.t16 VDD.t26 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X182 G_sink_up G1_1.t79 SD1_1.t0 VDD.t72 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X183 VDD G1_2.t10 G1_2.t11 VDD.t41 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X184 VSS G_sink_dn.t34 SD0_1.t9 VSS.t98 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X185 VDD G1_2.t8 G1_2.t9 VDD.t6 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X186 SD0_1 G_sink_dn.t35 VSS.t116 VSS.t112 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X187 SD2_1 G2_1.t89 VSS.t1 VSS.t0 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
R0 G2_1.n133 G2_1.n132 74.2622
R1 G2_1.n26 G2_1.n23 71.202
R2 G2_1.n28 G2_1.t6 37.4414
R3 G2_1.n116 G2_1.t34 37.4414
R4 G2_1.n132 G2_1.n131 21.0894
R5 G2_1.n131 G2_1.n130 21.0894
R6 G2_1.n130 G2_1.n129 21.0894
R7 G2_1.n129 G2_1.n128 21.0894
R8 G2_1.n128 G2_1.n127 21.0894
R9 G2_1.n127 G2_1.n126 21.0894
R10 G2_1.n126 G2_1.n125 21.0894
R11 G2_1.n125 G2_1.n124 21.0894
R12 G2_1.n124 G2_1.n123 21.0894
R13 G2_1.n15 G2_1.n14 21.0894
R14 G2_1.n16 G2_1.n15 21.0894
R15 G2_1.n17 G2_1.n16 21.0894
R16 G2_1.n18 G2_1.n17 21.0894
R17 G2_1.n19 G2_1.n18 21.0894
R18 G2_1.n20 G2_1.n19 21.0894
R19 G2_1.n21 G2_1.n20 21.0894
R20 G2_1.n22 G2_1.n21 21.0894
R21 G2_1.n23 G2_1.n22 21.0894
R22 G2_1.n131 G2_1.t66 16.5715
R23 G2_1.n130 G2_1.t87 16.5715
R24 G2_1.n127 G2_1.t78 16.5715
R25 G2_1.n126 G2_1.t63 16.5715
R26 G2_1.n123 G2_1.t84 16.5715
R27 G2_1.n14 G2_1.t88 16.5715
R28 G2_1.n17 G2_1.t80 16.5715
R29 G2_1.n18 G2_1.t65 16.5715
R30 G2_1.n21 G2_1.t75 16.5715
R31 G2_1.n22 G2_1.t89 16.5715
R32 G2_1.n132 G2_1.t70 16.3525
R33 G2_1.n129 G2_1.t61 16.3525
R34 G2_1.n128 G2_1.t77 16.3525
R35 G2_1.n125 G2_1.t76 16.3525
R36 G2_1.n124 G2_1.t60 16.3525
R37 G2_1.n15 G2_1.t62 16.3525
R38 G2_1.n16 G2_1.t83 16.3525
R39 G2_1.n19 G2_1.t86 16.3525
R40 G2_1.n20 G2_1.t72 16.3525
R41 G2_1.n23 G2_1.t64 16.3525
R42 G2_1.n104 G2_1.t8 14.0165
R43 G2_1.n101 G2_1.t26 14.0165
R44 G2_1.n92 G2_1.t10 14.0165
R45 G2_1.n89 G2_1.t4 14.0165
R46 G2_1.n82 G2_1.t18 14.0165
R47 G2_1.n79 G2_1.t32 14.0165
R48 G2_1.n70 G2_1.t24 14.0165
R49 G2_1.n67 G2_1.t28 14.0165
R50 G2_1.n62 G2_1.t14 14.0165
R51 G2_1.n59 G2_1.t2 14.0165
R52 G2_1.n52 G2_1.t20 14.0165
R53 G2_1.n49 G2_1.t30 14.0165
R54 G2_1.n44 G2_1.t12 14.0165
R55 G2_1.n41 G2_1.t36 14.0165
R56 G2_1.n32 G2_1.t16 14.0165
R57 G2_1.n29 G2_1.t0 14.0165
R58 G2_1.n113 G2_1.t38 14.0165
R59 G2_1.n115 G2_1.t22 13.7245
R60 G2_1.n30 G2_1.n29 4.0005
R61 G2_1.n33 G2_1.n32 4.0005
R62 G2_1.n42 G2_1.n41 4.0005
R63 G2_1.n45 G2_1.n44 4.0005
R64 G2_1.n50 G2_1.n49 4.0005
R65 G2_1.n53 G2_1.n52 4.0005
R66 G2_1.n60 G2_1.n59 4.0005
R67 G2_1.n63 G2_1.n62 4.0005
R68 G2_1.n68 G2_1.n67 4.0005
R69 G2_1.n71 G2_1.n70 4.0005
R70 G2_1.n80 G2_1.n79 4.0005
R71 G2_1.n83 G2_1.n82 4.0005
R72 G2_1.n90 G2_1.n89 4.0005
R73 G2_1.n93 G2_1.n92 4.0005
R74 G2_1.n102 G2_1.n101 4.0005
R75 G2_1.n105 G2_1.n104 4.0005
R76 G2_1.n114 G2_1.n113 4.0005
R77 G2_1.n118 G2_1.n117 4.0005
R78 G2_1.n26 G2_1.n25 3.58493
R79 G2_1.n108 G2_1.n107 3.57898
R80 G2_1.n86 G2_1.n85 3.57507
R81 G2_1.n133 G2_1.n122 3.5665
R82 G2_1.n46 G2_1.n11 3.53988
R83 G2_1.n99 G2_1.n98 3.53861
R84 G2_1.n77 G2_1.n76 3.53721
R85 G2_1.n74 G2_1.n73 3.53202
R86 G2_1.n96 G2_1.n95 3.53202
R87 G2_1.n87 G2_1.n1 3.52224
R88 G2_1.n65 G2_1.n3 3.51637
R89 G2_1.n47 G2_1.n9 3.51246
R90 G2_1.n57 G2_1.n56 3.51057
R91 G2_1.n36 G2_1.n35 3.50854
R92 G2_1.n111 G2_1.n110 3.50645
R93 G2_1.n39 G2_1.n38 3.49699
R94 G2_1.n64 G2_1.n5 3.49116
R95 G2_1.n54 G2_1.n7 3.4806
R96 G2_1.n134 G2_1.n120 3.46399
R97 G2_1.n27 G2_1.n13 3.45496
R98 G2_1.n104 G2_1.n103 2.3365
R99 G2_1.n101 G2_1.n100 2.3365
R100 G2_1.n92 G2_1.n91 2.3365
R101 G2_1.n89 G2_1.n88 2.3365
R102 G2_1.n82 G2_1.n81 2.3365
R103 G2_1.n79 G2_1.n78 2.3365
R104 G2_1.n70 G2_1.n69 2.3365
R105 G2_1.n67 G2_1.n66 2.3365
R106 G2_1.n62 G2_1.n61 2.3365
R107 G2_1.n59 G2_1.n58 2.3365
R108 G2_1.n52 G2_1.n51 2.3365
R109 G2_1.n49 G2_1.n48 2.3365
R110 G2_1.n44 G2_1.n43 2.3365
R111 G2_1.n41 G2_1.n40 2.3365
R112 G2_1.n32 G2_1.n31 2.3365
R113 G2_1.n29 G2_1.n28 2.3365
R114 G2_1.n113 G2_1.n112 2.3365
R115 G2_1.n117 G2_1.n116 2.3365
R116 G2_1.n107 G2_1.t9 1.6385
R117 G2_1.n107 G2_1.n106 1.6385
R118 G2_1.n110 G2_1.t52 1.6385
R119 G2_1.n110 G2_1.n109 1.6385
R120 G2_1.n95 G2_1.t11 1.6385
R121 G2_1.n95 G2_1.n94 1.6385
R122 G2_1.n98 G2_1.t57 1.6385
R123 G2_1.n98 G2_1.n97 1.6385
R124 G2_1.n85 G2_1.t19 1.6385
R125 G2_1.n85 G2_1.n84 1.6385
R126 G2_1.n1 G2_1.t40 1.6385
R127 G2_1.n1 G2_1.n0 1.6385
R128 G2_1.n73 G2_1.t25 1.6385
R129 G2_1.n73 G2_1.n72 1.6385
R130 G2_1.n76 G2_1.t47 1.6385
R131 G2_1.n76 G2_1.n75 1.6385
R132 G2_1.n5 G2_1.t15 1.6385
R133 G2_1.n5 G2_1.n4 1.6385
R134 G2_1.n3 G2_1.t49 1.6385
R135 G2_1.n3 G2_1.n2 1.6385
R136 G2_1.n7 G2_1.t21 1.6385
R137 G2_1.n7 G2_1.n6 1.6385
R138 G2_1.n56 G2_1.t44 1.6385
R139 G2_1.n56 G2_1.n55 1.6385
R140 G2_1.n11 G2_1.t13 1.6385
R141 G2_1.n11 G2_1.n10 1.6385
R142 G2_1.n9 G2_1.t56 1.6385
R143 G2_1.n9 G2_1.n8 1.6385
R144 G2_1.n35 G2_1.t17 1.6385
R145 G2_1.n35 G2_1.n34 1.6385
R146 G2_1.n38 G2_1.t41 1.6385
R147 G2_1.n38 G2_1.n37 1.6385
R148 G2_1.n120 G2_1.t23 1.6385
R149 G2_1.n120 G2_1.n119 1.6385
R150 G2_1.n122 G2_1.t45 1.6385
R151 G2_1.n122 G2_1.n121 1.6385
R152 G2_1.n13 G2_1.t46 1.6385
R153 G2_1.n13 G2_1.n12 1.6385
R154 G2_1.n25 G2_1.t7 1.6385
R155 G2_1.n25 G2_1.n24 1.6385
R156 G2_1 G2_1.n134 0.362318
R157 G2_1.n117 G2_1.n115 0.2925
R158 G2_1.n83 G2_1.n80 0.253351
R159 G2_1.n118 G2_1.n114 0.197599
R160 G2_1.n33 G2_1.n30 0.197599
R161 G2_1.n53 G2_1.n50 0.197599
R162 G2_1.n71 G2_1.n68 0.197599
R163 G2_1.n93 G2_1.n90 0.197599
R164 G2_1.n45 G2_1.n42 0.172031
R165 G2_1.n63 G2_1.n60 0.172031
R166 G2_1.n105 G2_1.n102 0.172031
R167 G2_1.n39 G2_1.n36 0.100499
R168 G2_1.n47 G2_1.n46 0.093148
R169 G2_1.n65 G2_1.n64 0.0926899
R170 G2_1.n57 G2_1.n54 0.0817532
R171 G2_1.n87 G2_1.n86 0.0807174
R172 G2_1.n77 G2_1.n74 0.0742956
R173 G2_1.n99 G2_1.n96 0.0727632
R174 G2_1.n74 G2_1.n71 0.0708476
R175 G2_1.n96 G2_1.n93 0.0705535
R176 G2_1.n111 G2_1.n108 0.0688207
R177 G2_1.n114 G2_1.n111 0.0665096
R178 G2_1.n90 G2_1.n87 0.0655603
R179 G2_1.n68 G2_1.n65 0.0636092
R180 G2_1.n54 G2_1.n53 0.061636
R181 G2_1.n50 G2_1.n47 0.0606109
R182 G2_1.n36 G2_1.n33 0.0579026
R183 G2_1.n108 G2_1.n105 0.049875
R184 G2_1.n86 G2_1.n83 0.0488673
R185 G2_1.n102 G2_1.n99 0.0443624
R186 G2_1.n46 G2_1.n45 0.0432184
R187 G2_1.n80 G2_1.n77 0.0423084
R188 G2_1.n60 G2_1.n57 0.0409019
R189 G2_1.n64 G2_1.n63 0.0397098
R190 G2_1.n42 G2_1.n39 0.0396398
R191 G2_1.n30 G2_1.n27 0.0223182
R192 G2_1.n134 G2_1.n133 0.00742308
R193 G2_1 G2_1.n118 0.00504545
R194 G2_1.n27 G2_1.n26 0.00495545
R195 VSS.n105 VSS.t106 223.469
R196 VSS.n102 VSS.t93 208.894
R197 VSS.n100 VSS.t90 194.321
R198 VSS.n98 VSS.t88 179.746
R199 VSS.n96 VSS.t85 165.173
R200 VSS.n93 VSS.t109 150.599
R201 VSS.n116 VSS.t111 150.599
R202 VSS.n73 VSS.t97 138.453
R203 VSS.n91 VSS.t100 136.024
R204 VSS.n76 VSS.t99 123.879
R205 VSS.n167 VSS.t62 114.472
R206 VSS.n78 VSS.t112 109.305
R207 VSS.n164 VSS.t11 107.007
R208 VSS.n162 VSS.t21 99.5411
R209 VSS.n80 VSS.t103 94.7314
R210 VSS.n160 VSS.t4 92.0755
R211 VSS.n158 VSS.t31 84.61
R212 VSS.n82 VSS.t95 80.1575
R213 VSS.n155 VSS.t24 77.1445
R214 VSS.n177 VSS.t45 77.1445
R215 VSS.n153 VSS.t37 69.6789
R216 VSS.n85 VSS.t80 65.5835
R217 VSS.n151 VSS.t53 62.2134
R218 VSS.n69 VSS.t98 58.2965
R219 VSS.n149 VSS.t16 54.7478
R220 VSS.n87 VSS.t83 51.0095
R221 VSS.n146 VSS.t8 47.2823
R222 VSS.n144 VSS.t48 39.8167
R223 VSS.n142 VSS.t6 32.3512
R224 VSS.n140 VSS.t26 24.8856
R225 VSS.n137 VSS.t57 17.4201
R226 VSS.n30 VSS.t2 13.6873
R227 VSS.n128 VSS.t0 12.4431
R228 VSS.n135 VSS.t13 9.95456
R229 VSS.n17 VSS.n16 6.40927
R230 VSS.n283 VSS.t113 6.40764
R231 VSS.n270 VSS.t84 6.4068
R232 VSS.n272 VSS.n259 6.4068
R233 VSS.n255 VSS.n201 6.35296
R234 VSS.n57 VSS.n56 5.4245
R235 VSS.n35 VSS.n34 5.41019
R236 VSS.n253 VSS.t52 5.3939
R237 VSS.n200 VSS.t46 5.3802
R238 VSS.n173 VSS.n170 5.2005
R239 VSS.n180 VSS.n178 5.2005
R240 VSS.n31 VSS.n29 5.2005
R241 VSS.n31 VSS.n27 5.2005
R242 VSS.n129 VSS.n128 5.2005
R243 VSS.n132 VSS.n131 5.2005
R244 VSS.n134 VSS.n133 5.2005
R245 VSS.n136 VSS.n135 5.2005
R246 VSS.n138 VSS.n137 5.2005
R247 VSS.n141 VSS.n140 5.2005
R248 VSS.n143 VSS.n142 5.2005
R249 VSS.n145 VSS.n144 5.2005
R250 VSS.n147 VSS.n146 5.2005
R251 VSS.n150 VSS.n149 5.2005
R252 VSS.n152 VSS.n151 5.2005
R253 VSS.n154 VSS.n153 5.2005
R254 VSS.n156 VSS.n155 5.2005
R255 VSS.n159 VSS.n158 5.2005
R256 VSS.n161 VSS.n160 5.2005
R257 VSS.n163 VSS.n162 5.2005
R258 VSS.n165 VSS.n164 5.2005
R259 VSS.n168 VSS.n167 5.2005
R260 VSS.n180 VSS.n177 5.2005
R261 VSS.n111 VSS.n110 5.2005
R262 VSS.n12 VSS.n11 5.2005
R263 VSS.n117 VSS.n116 5.2005
R264 VSS.n117 VSS.n114 5.2005
R265 VSS.n71 VSS.n69 5.2005
R266 VSS.n71 VSS.n68 5.2005
R267 VSS.n74 VSS.n73 5.2005
R268 VSS.n77 VSS.n76 5.2005
R269 VSS.n79 VSS.n78 5.2005
R270 VSS.n81 VSS.n80 5.2005
R271 VSS.n83 VSS.n82 5.2005
R272 VSS.n86 VSS.n85 5.2005
R273 VSS.n88 VSS.n87 5.2005
R274 VSS.n90 VSS.n89 5.2005
R275 VSS.n92 VSS.n91 5.2005
R276 VSS.n94 VSS.n93 5.2005
R277 VSS.n97 VSS.n96 5.2005
R278 VSS.n99 VSS.n98 5.2005
R279 VSS.n101 VSS.n100 5.2005
R280 VSS.n103 VSS.n102 5.2005
R281 VSS.n106 VSS.n105 5.2005
R282 VSS.n131 VSS.t42 4.97753
R283 VSS.n31 VSS.n30 4.5005
R284 VSS.n180 VSS.n179 4.5005
R285 VSS.n117 VSS.n115 4.5005
R286 VSS.n71 VSS.n70 4.5005
R287 VSS.n64 VSS.n55 4.1554
R288 VSS.n66 VSS.n65 3.92314
R289 VSS.n286 VSS.n285 3.87094
R290 VSS.n67 VSS.n66 3.84637
R291 VSS.n166 VSS.n119 3.75507
R292 VSS.n157 VSS.n121 3.75507
R293 VSS.n148 VSS.n123 3.75507
R294 VSS.n139 VSS.n125 3.75507
R295 VSS.n130 VSS.n127 3.75507
R296 VSS.n224 VSS.n217 3.75507
R297 VSS.n230 VSS.n213 3.75507
R298 VSS.n236 VSS.n209 3.75507
R299 VSS.n242 VSS.n205 3.75507
R300 VSS.n245 VSS.n203 3.75507
R301 VSS.n239 VSS.n207 3.75507
R302 VSS.n233 VSS.n211 3.75507
R303 VSS.n227 VSS.n215 3.75507
R304 VSS.n221 VSS.n219 3.75507
R305 VSS.n50 VSS.n41 3.74137
R306 VSS.n45 VSS.n43 3.74137
R307 VSS.n189 VSS.n185 3.74137
R308 VSS.n194 VSS.n183 3.74137
R309 VSS.n265 VSS.n261 3.6768
R310 VSS.n277 VSS.n258 3.6768
R311 VSS.n104 VSS.n1 3.64159
R312 VSS.n95 VSS.n3 3.64159
R313 VSS.n84 VSS.n5 3.64159
R314 VSS.n75 VSS.n7 3.64159
R315 VSS.n285 VSS.n256 3.51026
R316 VSS.n261 VSS.t116 2.7305
R317 VSS.n261 VSS.n260 2.7305
R318 VSS.n258 VSS.t89 2.7305
R319 VSS.n258 VSS.n257 2.7305
R320 VSS.n1 VSS.t94 2.7305
R321 VSS.n1 VSS.n0 2.7305
R322 VSS.n3 VSS.t110 2.7305
R323 VSS.n3 VSS.n2 2.7305
R324 VSS.n5 VSS.t96 2.7305
R325 VSS.n5 VSS.n4 2.7305
R326 VSS.n7 VSS.t117 2.7305
R327 VSS.n7 VSS.n6 2.7305
R328 VSS.n37 VSS.n36 2.60175
R329 VSS.n174 VSS.n173 2.60175
R330 VSS.n59 VSS.n58 2.60175
R331 VSS.n249 VSS.n248 2.60175
R332 VSS.n25 VSS.n23 2.60175
R333 VSS.n112 VSS.n111 2.60175
R334 VSS.n15 VSS.n13 2.60175
R335 VSS.n13 VSS.n12 2.601
R336 VSS.n12 VSS.n10 2.601
R337 VSS.n111 VSS.n109 2.601
R338 VSS.n23 VSS.n22 2.601
R339 VSS.n173 VSS.n172 2.601
R340 VSS.n175 VSS.n174 2.601
R341 VSS.n287 VSS.n112 2.601
R342 VSS.n22 VSS.n21 2.48901
R343 VSS.n29 VSS.n28 2.48901
R344 VSS.n133 VSS.t29 2.48901
R345 VSS.n286 VSS.n117 2.41864
R346 VSS.n253 VSS.n252 2.41785
R347 VSS.n181 VSS.n180 2.41764
R348 VSS.n62 VSS.n61 2.40802
R349 VSS.n32 VSS.n31 2.40802
R350 VSS.n72 VSS.n71 2.40802
R351 VSS.n54 VSS.n39 2.40786
R352 VSS.n65 VSS.n33 2.25997
R353 VSS.n256 VSS.n181 2.25167
R354 VSS.n285 VSS.n284 2.2505
R355 VSS.n66 VSS.n20 2.2505
R356 VSS.n64 VSS.n63 2.2505
R357 VSS.n255 VSS.n254 2.2505
R358 VSS.n15 VSS.n14 2.17323
R359 VSS.n25 VSS.n24 2.16377
R360 VSS.n61 VSS.n60 2.13331
R361 VSS.n39 VSS.n38 2.13331
R362 VSS.n180 VSS.n176 2.02394
R363 VSS.n252 VSS.n250 2.02394
R364 VSS.n117 VSS.n113 2.02394
R365 VSS.n65 VSS.n64 1.87545
R366 VSS.n256 VSS.n255 1.87428
R367 VSS.n119 VSS.t12 1.6385
R368 VSS.n119 VSS.n118 1.6385
R369 VSS.n121 VSS.t70 1.6385
R370 VSS.n121 VSS.n120 1.6385
R371 VSS.n123 VSS.t9 1.6385
R372 VSS.n123 VSS.n122 1.6385
R373 VSS.n125 VSS.t64 1.6385
R374 VSS.n125 VSS.n124 1.6385
R375 VSS.n127 VSS.t1 1.6385
R376 VSS.n127 VSS.n126 1.6385
R377 VSS.n217 VSS.t47 1.6385
R378 VSS.n217 VSS.n216 1.6385
R379 VSS.n213 VSS.t20 1.6385
R380 VSS.n213 VSS.n212 1.6385
R381 VSS.n209 VSS.t77 1.6385
R382 VSS.n209 VSS.n208 1.6385
R383 VSS.n205 VSS.t34 1.6385
R384 VSS.n205 VSS.n204 1.6385
R385 VSS.n203 VSS.t61 1.6385
R386 VSS.n203 VSS.n202 1.6385
R387 VSS.n207 VSS.t25 1.6385
R388 VSS.n207 VSS.n206 1.6385
R389 VSS.n211 VSS.t18 1.6385
R390 VSS.n211 VSS.n210 1.6385
R391 VSS.n215 VSS.t58 1.6385
R392 VSS.n215 VSS.n214 1.6385
R393 VSS.n219 VSS.t51 1.6385
R394 VSS.n219 VSS.n218 1.6385
R395 VSS.n41 VSS.t30 1.6385
R396 VSS.n41 VSS.n40 1.6385
R397 VSS.n43 VSS.t7 1.6385
R398 VSS.n43 VSS.n42 1.6385
R399 VSS.n185 VSS.t54 1.6385
R400 VSS.n185 VSS.n184 1.6385
R401 VSS.n183 VSS.t5 1.6385
R402 VSS.n183 VSS.n182 1.6385
R403 VSS.n27 VSS.n26 1.24476
R404 VSS.n10 VSS.n9 0.556908
R405 VSS.n109 VSS.n108 0.447533
R406 VSS.n172 VSS.n171 0.447533
R407 VSS.n252 VSS.n251 0.430411
R408 VSS.n9 VSS.n8 0.248057
R409 VSS.n108 VSS.n107 0.24188
R410 VSS.n134 VSS.n132 0.129952
R411 VSS.n136 VSS.n134 0.129952
R412 VSS.n138 VSS.n136 0.129952
R413 VSS.n143 VSS.n141 0.129952
R414 VSS.n145 VSS.n143 0.129952
R415 VSS.n147 VSS.n145 0.129952
R416 VSS.n152 VSS.n150 0.129952
R417 VSS.n154 VSS.n152 0.129952
R418 VSS.n156 VSS.n154 0.129952
R419 VSS.n161 VSS.n159 0.129952
R420 VSS.n163 VSS.n161 0.129952
R421 VSS.n165 VSS.n163 0.129952
R422 VSS.n263 VSS.n262 0.129952
R423 VSS.n264 VSS.n263 0.129952
R424 VSS.n267 VSS.n266 0.129952
R425 VSS.n268 VSS.n267 0.129952
R426 VSS.n269 VSS.n268 0.129952
R427 VSS.n274 VSS.n273 0.129952
R428 VSS.n275 VSS.n274 0.129952
R429 VSS.n276 VSS.n275 0.129952
R430 VSS.n279 VSS.n278 0.129952
R431 VSS.n280 VSS.n279 0.129952
R432 VSS.n223 VSS.n222 0.129952
R433 VSS.n226 VSS.n225 0.129952
R434 VSS.n229 VSS.n228 0.129952
R435 VSS.n232 VSS.n231 0.129952
R436 VSS.n235 VSS.n234 0.129952
R437 VSS.n238 VSS.n237 0.129952
R438 VSS.n241 VSS.n240 0.129952
R439 VSS.n244 VSS.n243 0.129952
R440 VSS.n53 VSS.n52 0.129952
R441 VSS.n52 VSS.n51 0.129952
R442 VSS.n49 VSS.n48 0.129952
R443 VSS.n48 VSS.n47 0.129952
R444 VSS.n47 VSS.n46 0.129952
R445 VSS.n187 VSS.n186 0.129952
R446 VSS.n188 VSS.n187 0.129952
R447 VSS.n191 VSS.n190 0.129952
R448 VSS.n192 VSS.n191 0.129952
R449 VSS.n193 VSS.n192 0.129952
R450 VSS.n196 VSS.n195 0.129952
R451 VSS.n197 VSS.n196 0.129952
R452 VSS.n79 VSS.n77 0.129952
R453 VSS.n81 VSS.n79 0.129952
R454 VSS.n83 VSS.n81 0.129952
R455 VSS.n88 VSS.n86 0.129952
R456 VSS.n90 VSS.n88 0.129952
R457 VSS.n92 VSS.n90 0.129952
R458 VSS.n94 VSS.n92 0.129952
R459 VSS.n99 VSS.n97 0.129952
R460 VSS.n101 VSS.n99 0.129952
R461 VSS.n103 VSS.n101 0.129952
R462 VSS.n168 VSS.n166 0.120089
R463 VSS.n246 VSS.n245 0.120089
R464 VSS.n106 VSS.n104 0.120089
R465 VSS.n54 VSS.n53 0.118897
R466 VSS.n74 VSS.n72 0.117951
R467 VSS.n278 VSS.n277 0.112692
R468 VSS.n243 VSS.n242 0.112692
R469 VSS.n195 VSS.n194 0.112692
R470 VSS.n169 VSS.n168 0.10776
R471 VSS.n281 VSS.n280 0.10776
R472 VSS.n247 VSS.n246 0.10776
R473 VSS.n198 VSS.n197 0.10776
R474 VSS.n159 VSS.n157 0.105295
R475 VSS.n240 VSS.n239 0.105295
R476 VSS.n97 VSS.n95 0.105295
R477 VSS.n75 VSS.n74 0.0985137
R478 VSS.n273 VSS.n272 0.0978973
R479 VSS.n237 VSS.n236 0.0978973
R480 VSS.n190 VSS.n189 0.0978973
R481 VSS.n265 VSS.n264 0.0911164
R482 VSS.n150 VSS.n148 0.0905
R483 VSS.n234 VSS.n233 0.0905
R484 VSS.n84 VSS.n83 0.0837192
R485 VSS.n231 VSS.n230 0.0831027
R486 VSS.n45 VSS.n44 0.0831027
R487 VSS.n270 VSS.n269 0.0763219
R488 VSS.n141 VSS.n139 0.0757055
R489 VSS.n228 VSS.n227 0.0757055
R490 VSS VSS.n106 0.075089
R491 VSS.n130 VSS.n129 0.0695411
R492 VSS.n221 VSS.n220 0.0695411
R493 VSS.n225 VSS.n224 0.0683082
R494 VSS.n50 VSS.n49 0.0683082
R495 VSS.n224 VSS.n223 0.0621438
R496 VSS.n51 VSS.n50 0.0621438
R497 VSS.n132 VSS.n130 0.060911
R498 VSS.n222 VSS.n221 0.060911
R499 VSS.n139 VSS.n138 0.0547466
R500 VSS.n227 VSS.n226 0.0547466
R501 VSS.n271 VSS.n270 0.0541301
R502 VSS.n230 VSS.n229 0.0473493
R503 VSS.n46 VSS.n45 0.0473493
R504 VSS.n86 VSS.n84 0.0467329
R505 VSS.n148 VSS.n147 0.0399521
R506 VSS.n233 VSS.n232 0.0399521
R507 VSS.n266 VSS.n265 0.0393356
R508 VSS VSS.n288 0.0331712
R509 VSS.n272 VSS.n271 0.0325548
R510 VSS.n236 VSS.n235 0.0325548
R511 VSS.n189 VSS.n188 0.0325548
R512 VSS.n77 VSS.n75 0.0319384
R513 VSS.n157 VSS.n156 0.0251575
R514 VSS.n239 VSS.n238 0.0251575
R515 VSS.n95 VSS.n94 0.0251575
R516 VSS.n175 VSS.n169 0.0226918
R517 VSS.n282 VSS.n281 0.0226918
R518 VSS.n249 VSS.n247 0.0226918
R519 VSS.n37 VSS.n35 0.0226918
R520 VSS.n199 VSS.n198 0.0226918
R521 VSS.n288 VSS.n287 0.0226918
R522 VSS.n18 VSS.n17 0.0220753
R523 VSS.n59 VSS.n57 0.0220753
R524 VSS.n277 VSS.n276 0.0177603
R525 VSS.n242 VSS.n241 0.0177603
R526 VSS.n194 VSS.n193 0.0177603
R527 VSS.n55 VSS.n54 0.0112717
R528 VSS.n63 VSS.n62 0.010987
R529 VSS.n33 VSS.n32 0.010987
R530 VSS.n20 VSS.n19 0.010987
R531 VSS.n72 VSS.n67 0.010987
R532 VSS.n166 VSS.n165 0.010363
R533 VSS.n245 VSS.n244 0.010363
R534 VSS.n104 VSS.n103 0.010363
R535 VSS.n33 VSS.n25 0.00358219
R536 VSS.n63 VSS.n59 0.00358219
R537 VSS.n20 VSS.n18 0.00296575
R538 VSS.n67 VSS.n15 0.00296575
R539 VSS.n181 VSS.n175 0.00234932
R540 VSS.n284 VSS.n282 0.00234932
R541 VSS.n254 VSS.n249 0.00234932
R542 VSS.n201 VSS.n199 0.00234932
R543 VSS.n287 VSS.n286 0.00234932
R544 VSS.n55 VSS.n37 0.00173288
R545 VSS.n254 VSS.n253 0.00128532
R546 VSS.n201 VSS.n200 0.00128532
R547 VSS.n284 VSS.n283 0.00128532
R548 ITAIL.n22 ITAIL.t52 120.174
R549 ITAIL.n75 ITAIL.t60 120.174
R550 ITAIL.n49 ITAIL.n48 106.159
R551 ITAIL.n130 ITAIL.n129 103.823
R552 ITAIL.n24 ITAIL.n23 103.823
R553 ITAIL.n77 ITAIL.n76 103.823
R554 ITAIL.n68 ITAIL.n67 103.823
R555 ITAIL.n12 ITAIL.n11 103.823
R556 ITAIL.n93 ITAIL.n92 103.823
R557 ITAIL.n54 ITAIL.n53 103.823
R558 ITAIL.n140 ITAIL.n139 103.823
R559 ITAIL.n145 ITAIL.n144 103.823
R560 ITAIL.n67 ITAIL.t66 37.2224
R561 ITAIL.n11 ITAIL.t59 37.2224
R562 ITAIL.n23 ITAIL.n22 21.0894
R563 ITAIL.n25 ITAIL.n24 21.0894
R564 ITAIL.n76 ITAIL.n75 21.0894
R565 ITAIL.n78 ITAIL.n77 21.0894
R566 ITAIL.n13 ITAIL.n12 21.0894
R567 ITAIL.n34 ITAIL.n33 21.0894
R568 ITAIL.n69 ITAIL.n68 21.0894
R569 ITAIL.n22 ITAIL.t62 16.3525
R570 ITAIL.n23 ITAIL.t44 16.3525
R571 ITAIL.n24 ITAIL.t43 16.3525
R572 ITAIL.n75 ITAIL.t49 16.3525
R573 ITAIL.n76 ITAIL.t68 16.3525
R574 ITAIL.n77 ITAIL.t67 16.3525
R575 ITAIL.n67 ITAIL.t57 16.1335
R576 ITAIL.n68 ITAIL.t45 16.1335
R577 ITAIL.n11 ITAIL.t42 16.1335
R578 ITAIL.n12 ITAIL.t65 16.1335
R579 ITAIL.n33 ITAIL.t54 16.1335
R580 ITAIL.n48 ITAIL.t18 14.0165
R581 ITAIL.n50 ITAIL.t28 14.0165
R582 ITAIL.n52 ITAIL.t32 14.0165
R583 ITAIL.n55 ITAIL.t36 14.0165
R584 ITAIL.n7 ITAIL.t2 14.0165
R585 ITAIL.n141 ITAIL.t22 14.0165
R586 ITAIL.n143 ITAIL.t24 13.9435
R587 ITAIL.n89 ITAIL.t4 13.7975
R588 ITAIL.n91 ITAIL.t8 13.7975
R589 ITAIL.n126 ITAIL.t16 13.7975
R590 ITAIL.n128 ITAIL.t12 13.7975
R591 ITAIL.n119 ITAIL.t30 13.7975
R592 ITAIL.n111 ITAIL.t26 13.7975
R593 ITAIL.n94 ITAIL.t10 13.7975
R594 ITAIL.n79 ITAIL.t48 13.3985
R595 ITAIL.n26 ITAIL.t50 13.3702
R596 ITAIL.n147 ITAIL.t38 12.7902
R597 ITAIL.n59 ITAIL.t0 12.7453
R598 ITAIL.n122 ITAIL.t34 12.5263
R599 ITAIL.n71 ITAIL.t64 12.5263
R600 ITAIL.n15 ITAIL.t47 12.4812
R601 ITAIL.n36 ITAIL.t58 12.4812
R602 ITAIL.n105 ITAIL.t20 12.4795
R603 ITAIL.n97 ITAIL.t14 12.4359
R604 ITAIL.n2 ITAIL.t6 11.6805
R605 ITAIL.n48 ITAIL.n47 9.23263
R606 ITAIL.n148 ITAIL.t39 5.20163
R607 ITAIL.n90 ITAIL.n89 4.15465
R608 ITAIL.n91 ITAIL.n90 4.15465
R609 ITAIL.n127 ITAIL.n126 4.15465
R610 ITAIL.n128 ITAIL.n127 4.15465
R611 ITAIL.n120 ITAIL.n119 4.15465
R612 ITAIL.n112 ITAIL.n111 4.15465
R613 ITAIL.n95 ITAIL.n94 4.15465
R614 ITAIL.n51 ITAIL.n50 4.15465
R615 ITAIL.n52 ITAIL.n51 4.15465
R616 ITAIL.n56 ITAIL.n55 4.15465
R617 ITAIL.n8 ITAIL.n7 4.15465
R618 ITAIL.n142 ITAIL.n141 4.15465
R619 ITAIL.n143 ITAIL.n142 4.15465
R620 ITAIL.n80 ITAIL.n79 3.75668
R621 ITAIL.n27 ITAIL.n26 3.75431
R622 ITAIL.n16 ITAIL.n14 3.549
R623 ITAIL.n149 ITAIL.n147 3.51942
R624 ITAIL.n72 ITAIL.n70 3.51322
R625 ITAIL.n106 ITAIL.n104 3.50928
R626 ITAIL.n123 ITAIL.n122 3.50535
R627 ITAIL.n72 ITAIL.n71 3.50535
R628 ITAIL.n138 ITAIL.n137 3.50535
R629 ITAIL.n37 ITAIL.n35 3.49926
R630 ITAIL.n106 ITAIL.n105 3.49877
R631 ITAIL.n16 ITAIL.n15 3.4914
R632 ITAIL.n37 ITAIL.n36 3.4914
R633 ITAIL.n98 ITAIL.n97 3.47756
R634 ITAIL.n152 ITAIL.n150 3.46513
R635 ITAIL.n51 ITAIL.n46 3.43811
R636 ITAIL.n56 ITAIL.n44 3.43811
R637 ITAIL.n8 ITAIL.n5 3.43811
R638 ITAIL.n142 ITAIL.n1 3.43615
R639 ITAIL.n90 ITAIL.n88 3.43224
R640 ITAIL.n127 ITAIL.n125 3.43224
R641 ITAIL.n120 ITAIL.n117 3.43224
R642 ITAIL.n112 ITAIL.n109 3.43224
R643 ITAIL.n95 ITAIL.n86 3.43224
R644 ITAIL.n102 ITAIL.n101 2.90675
R645 ITAIL.n74 ITAIL.n73 2.88464
R646 ITAIL.n18 ITAIL.n17 2.88464
R647 ITAIL.n39 ITAIL.n38 2.88464
R648 ITAIL.n101 ITAIL.n100 2.88464
R649 ITAIL.n150 ITAIL.n146 2.88451
R650 ITAIL.n132 ITAIL.n131 2.88438
R651 ITAIL.n133 ITAIL.n132 2.87461
R652 ITAIL.n113 ITAIL.n107 2.8741
R653 ITAIL.n144 ITAIL.n143 2.4095
R654 ITAIL.n92 ITAIL.n91 2.3365
R655 ITAIL.n129 ITAIL.n128 2.3365
R656 ITAIL.n119 ITAIL.n118 2.3365
R657 ITAIL.n111 ITAIL.n110 2.3365
R658 ITAIL.n100 ITAIL.n99 2.3365
R659 ITAIL.n94 ITAIL.n93 2.3365
R660 ITAIL.n50 ITAIL.n49 2.3365
R661 ITAIL.n53 ITAIL.n52 2.3365
R662 ITAIL.n55 ITAIL.n54 2.3365
R663 ITAIL.n7 ITAIL.n6 2.3365
R664 ITAIL.n141 ITAIL.n140 2.3365
R665 ITAIL.n131 ITAIL.n130 2.2635
R666 ITAIL.n3 ITAIL.n2 2.2635
R667 ITAIL.n152 ITAIL.n151 2.2565
R668 ITAIL.n83 ITAIL.n74 2.2505
R669 ITAIL.n20 ITAIL.n18 2.2505
R670 ITAIL.n40 ITAIL.n39 2.2505
R671 ITAIL.n115 ITAIL.n114 2.2505
R672 ITAIL.n63 ITAIL.n62 2.2505
R673 ITAIL.n136 ITAIL.n135 2.2505
R674 ITAIL.n60 ITAIL.n58 2.1905
R675 ITAIL.n146 ITAIL.n145 2.1175
R676 ITAIL.n61 ITAIL.n60 2.11497
R677 ITAIL.n26 ITAIL.n25 1.92893
R678 ITAIL.n79 ITAIL.n78 1.9031
R679 ITAIL.n88 ITAIL.t5 1.6385
R680 ITAIL.n88 ITAIL.n87 1.6385
R681 ITAIL.n125 ITAIL.t13 1.6385
R682 ITAIL.n125 ITAIL.n124 1.6385
R683 ITAIL.n117 ITAIL.t31 1.6385
R684 ITAIL.n117 ITAIL.n116 1.6385
R685 ITAIL.n109 ITAIL.t27 1.6385
R686 ITAIL.n109 ITAIL.n108 1.6385
R687 ITAIL.n86 ITAIL.t11 1.6385
R688 ITAIL.n86 ITAIL.n85 1.6385
R689 ITAIL.n46 ITAIL.t29 1.6385
R690 ITAIL.n46 ITAIL.n45 1.6385
R691 ITAIL.n44 ITAIL.t37 1.6385
R692 ITAIL.n44 ITAIL.n43 1.6385
R693 ITAIL.n5 ITAIL.t3 1.6385
R694 ITAIL.n5 ITAIL.n4 1.6385
R695 ITAIL.n1 ITAIL.t23 1.6385
R696 ITAIL.n1 ITAIL.n0 1.6385
R697 ITAIL.n134 ITAIL.n133 1.22514
R698 ITAIL.n28 ITAIL.n27 1.16042
R699 ITAIL.n21 ITAIL.n10 1.12967
R700 ITAIL.n40 ITAIL.n31 1.12556
R701 ITAIL.n81 ITAIL.n80 1.12469
R702 ITAIL.n60 ITAIL.n59 1.06529
R703 ITAIL.n139 ITAIL.n138 1.06529
R704 ITAIL.n138 ITAIL.n3 1.06529
R705 ITAIL.n104 ITAIL.n103 1.02542
R706 ITAIL.n35 ITAIL.n34 1.01842
R707 ITAIL.n135 ITAIL.n65 1.01782
R708 ITAIL.n14 ITAIL.n13 1.00064
R709 ITAIL.n70 ITAIL.n69 0.99056
R710 ITAIL.n83 ITAIL.n82 0.933875
R711 ITAIL.n42 ITAIL.n21 0.850862
R712 ITAIL.n134 ITAIL.n84 0.785857
R713 ITAIL.n133 ITAIL.n115 0.652981
R714 ITAIL.n115 ITAIL.n102 0.604805
R715 ITAIL.n82 ITAIL.n81 0.558332
R716 ITAIL.n65 ITAIL.n42 0.503536
R717 ITAIL.n29 ITAIL.n28 0.249615
R718 ITAIL.n65 ITAIL.n64 0.245589
R719 ITAIL.n61 ITAIL.n56 0.147502
R720 ITAIL.n113 ITAIL.n112 0.141303
R721 ITAIL.n121 ITAIL.n120 0.124649
R722 ITAIL.n9 ITAIL.n8 0.123649
R723 ITAIL.n96 ITAIL.n95 0.122649
R724 ITAIL.n58 ITAIL.n57 0.0735
R725 ITAIL.n41 ITAIL.n40 0.0374863
R726 ITAIL.n40 ITAIL.n32 0.0362534
R727 ITAIL.n98 ITAIL.n96 0.0325
R728 ITAIL.n20 ITAIL.n19 0.0315
R729 ITAIL.n137 ITAIL.n9 0.0315
R730 ITAIL.n149 ITAIL.n148 0.0315
R731 ITAIL.n123 ITAIL.n121 0.0305
R732 ITAIL.n31 ITAIL.n29 0.0305
R733 ITAIL.n31 ITAIL.n30 0.0295
R734 ITAIL.n64 ITAIL.n63 0.0215938
R735 ITAIL.n84 ITAIL.n66 0.0205
R736 ITAIL.n114 ITAIL.n113 0.0117741
R737 ITAIL.n84 ITAIL.n83 0.0105
R738 ITAIL.n62 ITAIL.n61 0.00955805
R739 ITAIL.n135 ITAIL.n134 0.00692857
R740 ITAIL ITAIL.n152 0.0065
R741 ITAIL.n42 ITAIL.n41 0.00543151
R742 ITAIL.n114 ITAIL.n106 0.0035
R743 ITAIL.n132 ITAIL.n123 0.0025
R744 ITAIL.n18 ITAIL.n16 0.0025
R745 ITAIL.n137 ITAIL.n136 0.0025
R746 ITAIL.n21 ITAIL.n20 0.00187264
R747 ITAIL.n39 ITAIL.n37 0.0015
R748 ITAIL.n74 ITAIL.n72 0.0015
R749 ITAIL.n101 ITAIL.n98 0.0015
R750 ITAIL.n150 ITAIL.n149 0.0015
R751 G1_2.n130 G1_2.n129 103.823
R752 G1_2.n128 G1_2.n127 103.823
R753 G1_2.n126 G1_2.n125 103.823
R754 G1_2.n124 G1_2.n123 103.823
R755 G1_2.n108 G1_2.n105 90.2366
R756 G1_2.n54 G1_2.n51 90.0338
R757 G1_2.n21 G1_2.n18 89.6266
R758 G1_2.n113 G1_2.n112 89.2199
R759 G1_2.n86 G1_2.n85 86.0167
R760 G1_2.n46 G1_2.n43 85.9783
R761 G1_2.n48 G1_2.n47 25.6154
R762 G1_2.n102 G1_2.n101 25.6154
R763 G1_2.n112 G1_2.n109 25.6154
R764 G1_2.n59 G1_2.n55 25.5424
R765 G1_2.n91 G1_2.n90 25.3234
R766 G1_2.n84 G1_2.n83 25.3234
R767 G1_2.n70 G1_2.n69 25.3234
R768 G1_2.n25 G1_2.n22 25.3234
R769 G1_2.n15 G1_2.n14 25.1774
R770 G1_2.n129 G1_2.n128 21.0894
R771 G1_2.n127 G1_2.n126 21.0894
R772 G1_2.n125 G1_2.n124 21.0894
R773 G1_2.n123 G1_2.n122 21.0894
R774 G1_2.n15 G1_2.t22 14.1625
R775 G1_2.n47 G1_2.t32 14.0895
R776 G1_2.n48 G1_2.t12 14.0895
R777 G1_2.n55 G1_2.t6 14.0895
R778 G1_2.n58 G1_2.t8 14.0895
R779 G1_2.n101 G1_2.t38 14.0895
R780 G1_2.n102 G1_2.t20 14.0895
R781 G1_2.n109 G1_2.t30 14.0895
R782 G1_2.n112 G1_2.t10 14.0895
R783 G1_2.n41 G1_2.t26 14.0535
R784 G1_2.n90 G1_2.t42 14.0165
R785 G1_2.n83 G1_2.t24 14.0165
R786 G1_2.n84 G1_2.t34 14.0165
R787 G1_2.n70 G1_2.t14 14.0165
R788 G1_2.n69 G1_2.t28 14.0165
R789 G1_2.n14 G1_2.t36 14.0165
R790 G1_2.n22 G1_2.t44 14.0165
R791 G1_2.n118 G1_2.t40 14.0165
R792 G1_2.n92 G1_2.t18 13.8688
R793 G1_2.n26 G1_2.t16 13.6515
R794 G1_2.n129 G1_2.t76 13.4325
R795 G1_2.n128 G1_2.t67 13.4325
R796 G1_2.n127 G1_2.t66 13.4325
R797 G1_2.n126 G1_2.t73 13.4325
R798 G1_2.n125 G1_2.t77 13.4325
R799 G1_2.n124 G1_2.t69 13.4325
R800 G1_2.n123 G1_2.t70 13.4325
R801 G1_2.n122 G1_2.t63 13.4325
R802 G1_2.n33 G1_2.t79 9.73306
R803 G1_2.n133 G1_2.t62 8.6145
R804 G1_2.n94 G1_2.n86 8.02477
R805 G1_2.n130 G1_2.n0 8.0005
R806 G1_2.n83 G1_2.n82 7.31048
R807 G1_2.n14 G1_2.n13 7.28939
R808 G1_2.n112 G1_2.n111 6.99488
R809 G1_2.n18 G1_2.n17 6.98985
R810 G1_2.n89 G1_2.n88 6.98577
R811 G1_2.n105 G1_2.n104 6.9857
R812 G1_2.n46 G1_2.n45 6.98386
R813 G1_2.n54 G1_2.n53 6.98202
R814 G1_2.n51 G1_2.n50 6.98202
R815 G1_2.n68 G1_2.n67 6.92657
R816 G1_2.n85 G1_2.n80 6.92657
R817 G1_2.n21 G1_2.n20 6.92657
R818 G1_2.n108 G1_2.n107 6.92646
R819 G1_2.n38 G1_2.n37 5.62918
R820 G1_2.n135 G1_2.n121 5.6219
R821 G1_2.n96 G1_2.n95 4.5005
R822 G1_2.n121 G1_2.n120 4.5005
R823 G1_2.n57 G1_2.n56 4.3805
R824 G1_2.n43 G1_2.n42 4.11505
R825 G1_2.n93 G1_2.n92 3.94099
R826 G1_2.n35 G1_2.n34 3.4914
R827 G1_2.n35 G1_2.n33 3.48541
R828 G1_2.n117 G1_2.n113 3.152
R829 G1_2.n74 G1_2.n73 2.96161
R830 G1_2.n39 G1_2.n31 2.95451
R831 G1_2.n116 G1_2.n115 2.94775
R832 G1_2.n97 G1_2.n78 2.94616
R833 G1_2.n62 G1_2.n61 2.93059
R834 G1_2.n4 G1_2.n3 2.92692
R835 G1_2.n9 G1_2.n8 2.9268
R836 G1_2.n29 G1_2.n28 2.91729
R837 G1_2.n64 G1_2.n59 2.88761
R838 G1_2.n101 G1_2.n100 2.88761
R839 G1_2.n135 G1_2.n134 2.88564
R840 G1_2.n37 G1_2.n36 2.88464
R841 G1_2.n27 G1_2.n26 2.86878
R842 G1_2.n40 G1_2.n39 2.86794
R843 G1_2.n98 G1_2.n97 2.62905
R844 G1_2.n134 G1_2.n133 2.3365
R845 G1_2.n76 G1_2.n75 2.2505
R846 G1_2.n65 G1_2.n64 2.2505
R847 G1_2.n100 G1_2.n99 2.2505
R848 G1_2.n24 G1_2.n23 2.22892
R849 G1_2.n131 G1_2.n130 2.1175
R850 G1_2.n111 G1_2.t11 1.8205
R851 G1_2.n111 G1_2.n110 1.8205
R852 G1_2.n107 G1_2.t56 1.8205
R853 G1_2.n107 G1_2.n106 1.8205
R854 G1_2.n104 G1_2.t21 1.8205
R855 G1_2.n104 G1_2.n103 1.8205
R856 G1_2.n8 G1_2.t17 1.8205
R857 G1_2.n8 G1_2.n7 1.8205
R858 G1_2.n67 G1_2.t5 1.8205
R859 G1_2.n67 G1_2.n66 1.8205
R860 G1_2.n88 G1_2.t54 1.8205
R861 G1_2.n88 G1_2.n87 1.8205
R862 G1_2.n78 G1_2.t19 1.8205
R863 G1_2.n78 G1_2.n77 1.8205
R864 G1_2.n80 G1_2.t58 1.8205
R865 G1_2.n80 G1_2.n79 1.8205
R866 G1_2.n82 G1_2.t25 1.8205
R867 G1_2.n82 G1_2.n81 1.8205
R868 G1_2.n73 G1_2.t15 1.8205
R869 G1_2.n73 G1_2.n72 1.8205
R870 G1_2.n20 G1_2.t57 1.8205
R871 G1_2.n20 G1_2.n19 1.8205
R872 G1_2.n17 G1_2.t23 1.8205
R873 G1_2.n17 G1_2.n16 1.8205
R874 G1_2.n13 G1_2.t4 1.8205
R875 G1_2.n13 G1_2.n12 1.8205
R876 G1_2.n53 G1_2.t55 1.8205
R877 G1_2.n53 G1_2.n52 1.8205
R878 G1_2.n50 G1_2.t13 1.8205
R879 G1_2.n50 G1_2.n49 1.8205
R880 G1_2.n45 G1_2.t51 1.8205
R881 G1_2.n45 G1_2.n44 1.8205
R882 G1_2.n31 G1_2.t27 1.8205
R883 G1_2.n31 G1_2.n30 1.8205
R884 G1_2.n61 G1_2.t9 1.8205
R885 G1_2.n61 G1_2.n60 1.8205
R886 G1_2.n3 G1_2.t3 1.8205
R887 G1_2.n3 G1_2.n2 1.8205
R888 G1_2.n115 G1_2.t48 1.8205
R889 G1_2.n115 G1_2.n114 1.8205
R890 G1_2.n75 G1_2.n71 1.61816
R891 G1_2.n65 G1_2.n29 1.41264
R892 G1_2.n99 G1_2.n98 1.38535
R893 G1_2.n101 G1_2.n1 1.20181
R894 G1_2.n71 G1_2.n70 0.853387
R895 G1_2.n99 G1_2.n65 0.696503
R896 G1_2.n18 G1_2.n15 0.642258
R897 G1_2.n85 G1_2.n84 0.384711
R898 G1_2.n69 G1_2.n68 0.384711
R899 G1_2.n22 G1_2.n21 0.384711
R900 G1_2.n26 G1_2.n25 0.3655
R901 G1_2.n109 G1_2.n108 0.298459
R902 G1_2.n132 G1_2.n131 0.292201
R903 G1_2.n25 G1_2.n24 0.231026
R904 G1_2.n51 G1_2.n48 0.223969
R905 G1_2.n55 G1_2.n54 0.223969
R906 G1_2.n90 G1_2.n89 0.154184
R907 G1_2.n47 G1_2.n46 0.14948
R908 G1_2.n58 G1_2.n57 0.1465
R909 G1_2.n92 G1_2.n91 0.143972
R910 G1_2.n120 G1_2.n119 0.140885
R911 G1_2.n42 G1_2.n40 0.133227
R912 G1_2.n98 G1_2.n76 0.120105
R913 G1_2.n105 G1_2.n102 0.0749898
R914 G1_2.n59 G1_2.n58 0.0735
R915 G1_2.n119 G1_2.n118 0.0735
R916 G1_2.n134 G1_2.n132 0.0734811
R917 G1_2.n63 G1_2.n62 0.055602
R918 G1_2.n5 G1_2.n4 0.0537653
R919 G1_2.n10 G1_2.n9 0.0519286
R920 G1_2.n42 G1_2.n41 0.037206
R921 G1_2.n117 G1_2.n116 0.0356143
R922 G1_2.n39 G1_2.n38 0.021405
R923 G1_2.n28 G1_2.n27 0.0200941
R924 G1_2.n75 G1_2.n74 0.019821
R925 G1_2.n97 G1_2.n96 0.019259
R926 G1_2.n96 G1_2.n94 0.01175
R927 G1_2.n28 G1_2.n11 0.0060102
R928 G1_2.n100 G1_2.n5 0.0060102
R929 G1_2.n94 G1_2.n93 0.00425
R930 G1_2.n64 G1_2.n63 0.00417347
R931 G1_2.n121 G1_2.n117 0.00417347
R932 G1_2.n10 G1_2.n6 0.00293243
R933 G1_2 G1_2.n0 0.0025
R934 G1_2.n11 G1_2.n10 0.00233673
R935 G1_2.n38 G1_2.n32 0.00233673
R936 G1_2.n37 G1_2.n35 0.0015
R937 G1_2 G1_2.n135 0.0015
R938 VDD.n151 VDD.t30 151.695
R939 VDD.n151 VDD.t15 148.749
R940 VDD.n136 VDD.t10 122.648
R941 VDD.n167 VDD.t24 122.444
R942 VDD.n148 VDD.t26 113.403
R943 VDD.n153 VDD.t9 110.457
R944 VDD.n164 VDD.t92 81.002
R945 VDD.n137 VDD.t90 78.0565
R946 VDD.n146 VDD.t27 75.111
R947 VDD.n155 VDD.t91 72.1654
R948 VDD.n76 VDD.t4 56.5849
R949 VDD.n60 VDD.t1 54.5272
R950 VDD.n60 VDD.t72 50.412
R951 VDD.n76 VDD.t45 48.3544
R952 VDD.n91 VDD.t80 45.268
R953 VDD.n75 VDD.t2 43.2104
R954 VDD.n162 VDD.t89 42.7104
R955 VDD.n59 VDD.t5 41.1528
R956 VDD.n139 VDD.t3 39.7649
R957 VDD.n61 VDD.t33 37.0375
R958 VDD.n144 VDD.t18 36.8194
R959 VDD.n81 VDD.t69 34.9799
R960 VDD.n157 VDD.t13 33.8738
R961 VDD.n93 VDD.t35 32.4079
R962 VDD.n90 VDD.t0 31.8935
R963 VDD.n74 VDD.t6 29.8359
R964 VDD.n66 VDD.t38 23.663
R965 VDD.n82 VDD.t85 21.6054
R966 VDD.n89 VDD.t41 18.519
R967 VDD.n69 VDD.t59 16.4614
R968 VDD.n67 VDD.t83 10.2886
R969 VDD.n83 VDD.t7 8.23095
R970 VDD.n108 VDD.t36 7.62593
R971 VDD.n134 VDD.n7 7.1505
R972 VDD.n57 VDD.n56 6.54575
R973 VDD.n102 VDD.n101 6.50606
R974 VDD.n110 VDD.n91 6.3005
R975 VDD.n111 VDD.n90 6.3005
R976 VDD.n112 VDD.n89 6.3005
R977 VDD.n114 VDD.n84 6.3005
R978 VDD.n115 VDD.n83 6.3005
R979 VDD.n116 VDD.n82 6.3005
R980 VDD.n117 VDD.n81 6.3005
R981 VDD.n119 VDD.n76 6.3005
R982 VDD.n120 VDD.n75 6.3005
R983 VDD.n121 VDD.n74 6.3005
R984 VDD.n123 VDD.n69 6.3005
R985 VDD.n124 VDD.n68 6.3005
R986 VDD.n125 VDD.n67 6.3005
R987 VDD.n126 VDD.n66 6.3005
R988 VDD.n128 VDD.n61 6.3005
R989 VDD.n129 VDD.n60 6.3005
R990 VDD.n130 VDD.n59 6.3005
R991 VDD.n12 VDD.n10 6.3005
R992 VDD.n96 VDD.n94 6.3005
R993 VDD.n12 VDD.n9 6.3005
R994 VDD.n138 VDD.n137 6.3005
R995 VDD.n140 VDD.n139 6.3005
R996 VDD.n142 VDD.n141 6.3005
R997 VDD.n145 VDD.n144 6.3005
R998 VDD.n147 VDD.n146 6.3005
R999 VDD.n149 VDD.n148 6.3005
R1000 VDD.n152 VDD.n151 6.3005
R1001 VDD.n154 VDD.n153 6.3005
R1002 VDD.n156 VDD.n155 6.3005
R1003 VDD.n158 VDD.n157 6.3005
R1004 VDD.n161 VDD.n160 6.3005
R1005 VDD.n163 VDD.n162 6.3005
R1006 VDD.n165 VDD.n164 6.3005
R1007 VDD.n168 VDD.t25 6.22476
R1008 VDD.n135 VDD.n6 6.21492
R1009 VDD.n84 VDD.t67 5.14453
R1010 VDD.n94 VDD.n93 5.14453
R1011 VDD.n108 VDD.t79 5.00941
R1012 VDD.n132 VDD.n58 5.00941
R1013 VDD.n63 VDD.t34 4.5505
R1014 VDD.n63 VDD.n62 4.5505
R1015 VDD.n71 VDD.t62 4.5505
R1016 VDD.n71 VDD.n70 4.5505
R1017 VDD.n78 VDD.t53 4.5505
R1018 VDD.n78 VDD.n77 4.5505
R1019 VDD.n86 VDD.t75 4.5505
R1020 VDD.n86 VDD.n85 4.5505
R1021 VDD.n12 VDD.n11 4.5005
R1022 VDD.n160 VDD.t21 4.41876
R1023 VDD.n16 VDD.n15 3.60132
R1024 VDD.n53 VDD.n23 3.18941
R1025 VDD.n48 VDD.n25 3.18941
R1026 VDD.n43 VDD.n27 3.18941
R1027 VDD.n39 VDD.n29 3.18941
R1028 VDD.n34 VDD.n31 3.18941
R1029 VDD.n127 VDD.n65 3.18941
R1030 VDD.n122 VDD.n73 3.18941
R1031 VDD.n118 VDD.n80 3.18941
R1032 VDD.n113 VDD.n88 3.18941
R1033 VDD.n159 VDD.n1 3.18159
R1034 VDD.n150 VDD.n3 3.18159
R1035 VDD.n143 VDD.n5 3.18159
R1036 VDD.n107 VDD.n106 3.15175
R1037 VDD.n18 VDD.n17 3.15175
R1038 VDD.n17 VDD.n16 3.151
R1039 VDD.n106 VDD.n105 3.151
R1040 VDD.n16 VDD.n14 3.151
R1041 VDD.n105 VDD.n104 3.151
R1042 VDD.n168 VDD.n167 3.1505
R1043 VDD.n68 VDD.t8 3.08692
R1044 VDD.n127 VDD.n63 3.07593
R1045 VDD.n122 VDD.n71 3.07593
R1046 VDD.n118 VDD.n78 3.07593
R1047 VDD.n113 VDD.n86 3.07593
R1048 VDD.n1 VDD.t14 3.03383
R1049 VDD.n1 VDD.n0 3.03383
R1050 VDD.n3 VDD.t31 3.03383
R1051 VDD.n3 VDD.n2 3.03383
R1052 VDD.n5 VDD.t29 3.03383
R1053 VDD.n5 VDD.n4 3.03383
R1054 VDD.n18 VDD.n13 2.76626
R1055 VDD.n20 VDD.n19 2.75233
R1056 VDD.n102 VDD.n96 2.62983
R1057 VDD.n100 VDD.n98 2.62936
R1058 VDD.n55 VDD.n21 2.62088
R1059 VDD.n135 VDD.n134 2.24061
R1060 VDD.n105 VDD.n103 2.05811
R1061 VDD.n23 VDD.t51 1.8205
R1062 VDD.n23 VDD.n22 1.8205
R1063 VDD.n25 VDD.t84 1.8205
R1064 VDD.n25 VDD.n24 1.8205
R1065 VDD.n27 VDD.t52 1.8205
R1066 VDD.n27 VDD.n26 1.8205
R1067 VDD.n29 VDD.t86 1.8205
R1068 VDD.n29 VDD.n28 1.8205
R1069 VDD.n31 VDD.t54 1.8205
R1070 VDD.n31 VDD.n30 1.8205
R1071 VDD.n65 VDD.t77 1.8205
R1072 VDD.n65 VDD.n64 1.8205
R1073 VDD.n73 VDD.t60 1.8205
R1074 VDD.n73 VDD.n72 1.8205
R1075 VDD.n80 VDD.t46 1.8205
R1076 VDD.n80 VDD.n79 1.8205
R1077 VDD.n88 VDD.t68 1.8205
R1078 VDD.n88 VDD.n87 1.8205
R1079 VDD.n96 VDD.n92 1.77932
R1080 VDD.n96 VDD.n95 1.61584
R1081 VDD.n98 VDD.n97 1.48285
R1082 VDD.n141 VDD.t28 1.47325
R1083 VDD.n9 VDD.n8 1.02931
R1084 VDD.n13 VDD.n12 0.78178
R1085 VDD.n134 VDD.n133 0.19404
R1086 VDD.n167 VDD.n166 0.111676
R1087 VDD.n52 VDD.n51 0.108313
R1088 VDD.n51 VDD.n50 0.108313
R1089 VDD.n50 VDD.n49 0.108313
R1090 VDD.n47 VDD.n46 0.108313
R1091 VDD.n46 VDD.n45 0.108313
R1092 VDD.n45 VDD.n44 0.108313
R1093 VDD.n42 VDD.n41 0.108313
R1094 VDD.n41 VDD.n40 0.108313
R1095 VDD.n38 VDD.n37 0.108313
R1096 VDD.n37 VDD.n36 0.108313
R1097 VDD.n36 VDD.n35 0.108313
R1098 VDD.n130 VDD.n129 0.108313
R1099 VDD.n129 VDD.n128 0.108313
R1100 VDD.n126 VDD.n125 0.108313
R1101 VDD.n125 VDD.n124 0.108313
R1102 VDD.n124 VDD.n123 0.108313
R1103 VDD.n121 VDD.n120 0.108313
R1104 VDD.n120 VDD.n119 0.108313
R1105 VDD.n117 VDD.n116 0.108313
R1106 VDD.n116 VDD.n115 0.108313
R1107 VDD.n115 VDD.n114 0.108313
R1108 VDD.n112 VDD.n111 0.108313
R1109 VDD.n111 VDD.n110 0.108313
R1110 VDD.n138 VDD.n136 0.108313
R1111 VDD.n140 VDD.n138 0.108313
R1112 VDD.n142 VDD.n140 0.108313
R1113 VDD.n147 VDD.n145 0.108313
R1114 VDD.n149 VDD.n147 0.108313
R1115 VDD.n154 VDD.n152 0.108313
R1116 VDD.n156 VDD.n154 0.108313
R1117 VDD.n158 VDD.n156 0.108313
R1118 VDD.n163 VDD.n161 0.108313
R1119 VDD.n165 VDD.n163 0.108313
R1120 VDD.n150 VDD.n149 0.107844
R1121 VDD VDD.n165 0.107375
R1122 VDD.n54 VDD.n53 0.106438
R1123 VDD.n43 VDD.n42 0.099875
R1124 VDD.n55 VDD.n54 0.0967182
R1125 VDD.n119 VDD.n118 0.092375
R1126 VDD.n34 VDD.n33 0.0895625
R1127 VDD.n110 VDD.n109 0.0890938
R1128 VDD.n33 VDD.n32 0.0844062
R1129 VDD.n131 VDD.n130 0.083
R1130 VDD.n128 VDD.n127 0.0820625
R1131 VDD.n122 VDD.n121 0.0755
R1132 VDD.n40 VDD.n39 0.068
R1133 VDD.n113 VDD.n112 0.0651875
R1134 VDD.n145 VDD.n143 0.0600312
R1135 VDD.n159 VDD.n158 0.0590938
R1136 VDD.n49 VDD.n48 0.0576875
R1137 VDD.n48 VDD.n47 0.051125
R1138 VDD.n161 VDD.n159 0.0497188
R1139 VDD.n143 VDD.n142 0.0487812
R1140 VDD.n114 VDD.n113 0.043625
R1141 VDD.n39 VDD.n38 0.0408125
R1142 VDD.n123 VDD.n122 0.0333125
R1143 VDD.n127 VDD.n126 0.02675
R1144 VDD.n35 VDD.n34 0.01925
R1145 VDD.n118 VDD.n117 0.0164375
R1146 VDD.n133 VDD.n132 0.0159688
R1147 VDD.n109 VDD.n108 0.0140938
R1148 VDD.n136 VDD.n135 0.0112812
R1149 VDD.n56 VDD.n55 0.00977193
R1150 VDD.n44 VDD.n43 0.0089375
R1151 VDD.n107 VDD.n102 0.008
R1152 VDD.n108 VDD.n107 0.006125
R1153 VDD.n57 VDD.n18 0.00565625
R1154 VDD.n56 VDD.n20 0.00378125
R1155 VDD.n132 VDD.n131 0.0033125
R1156 VDD.n53 VDD.n52 0.002375
R1157 VDD.n133 VDD.n57 0.002375
R1158 VDD.n100 VDD.n99 0.00209515
R1159 VDD.n101 VDD.n100 0.00177952
R1160 VDD VDD.n168 0.0014375
R1161 VDD.n152 VDD.n150 0.00096875
R1162 G_sink_dn.n11 G_sink_dn.n10 49.2755
R1163 G_sink_dn.n4 G_sink_dn.t34 33.7914
R1164 G_sink_dn.n35 G_sink_dn.t7 33.7914
R1165 G_sink_dn.n5 G_sink_dn.n4 21.0894
R1166 G_sink_dn.n6 G_sink_dn.n5 21.0894
R1167 G_sink_dn.n7 G_sink_dn.n6 21.0894
R1168 G_sink_dn.n8 G_sink_dn.n7 21.0894
R1169 G_sink_dn.n9 G_sink_dn.n8 21.0894
R1170 G_sink_dn.n10 G_sink_dn.n9 21.0894
R1171 G_sink_dn.n18 G_sink_dn.n11 21.0894
R1172 G_sink_dn.n25 G_sink_dn.n18 21.0894
R1173 G_sink_dn.n26 G_sink_dn.n25 21.0894
R1174 G_sink_dn.n27 G_sink_dn.n26 21.0894
R1175 G_sink_dn.n34 G_sink_dn.n27 21.0894
R1176 G_sink_dn.n35 G_sink_dn.n34 21.0894
R1177 G_sink_dn.n4 G_sink_dn.t31 13.0675
R1178 G_sink_dn.n5 G_sink_dn.t26 13.0675
R1179 G_sink_dn.n8 G_sink_dn.t24 13.0675
R1180 G_sink_dn.n9 G_sink_dn.t28 13.0675
R1181 G_sink_dn.n6 G_sink_dn.t35 12.7025
R1182 G_sink_dn.n7 G_sink_dn.t27 12.7025
R1183 G_sink_dn.n10 G_sink_dn.t29 12.7025
R1184 G_sink_dn.n11 G_sink_dn.t9 12.7025
R1185 G_sink_dn.n26 G_sink_dn.t21 12.7025
R1186 G_sink_dn.n27 G_sink_dn.t15 12.7025
R1187 G_sink_dn.n17 G_sink_dn.t13 10.7315
R1188 G_sink_dn.n24 G_sink_dn.t19 10.7315
R1189 G_sink_dn.n33 G_sink_dn.t17 10.7315
R1190 G_sink_dn.n36 G_sink_dn.t11 10.7315
R1191 G_sink_dn.n17 G_sink_dn.n16 4.1025
R1192 G_sink_dn.n24 G_sink_dn.n23 4.1025
R1193 G_sink_dn.n33 G_sink_dn.n32 4.1025
R1194 G_sink_dn.n37 G_sink_dn.n36 4.1025
R1195 G_sink_dn.n16 G_sink_dn.n15 3.4655
R1196 G_sink_dn.n23 G_sink_dn.n22 3.4655
R1197 G_sink_dn.n32 G_sink_dn.n31 3.4655
R1198 G_sink_dn.n37 G_sink_dn.n3 3.4655
R1199 G_sink_dn.n16 G_sink_dn.n13 3.35007
R1200 G_sink_dn.n23 G_sink_dn.n20 3.35007
R1201 G_sink_dn.n32 G_sink_dn.n29 3.35007
R1202 G_sink_dn.n37 G_sink_dn.n1 3.35007
R1203 G_sink_dn.n15 G_sink_dn.t10 2.7305
R1204 G_sink_dn.n15 G_sink_dn.n14 2.7305
R1205 G_sink_dn.n13 G_sink_dn.t3 2.7305
R1206 G_sink_dn.n13 G_sink_dn.n12 2.7305
R1207 G_sink_dn.n22 G_sink_dn.t0 2.7305
R1208 G_sink_dn.n22 G_sink_dn.n21 2.7305
R1209 G_sink_dn.n20 G_sink_dn.t20 2.7305
R1210 G_sink_dn.n20 G_sink_dn.n19 2.7305
R1211 G_sink_dn.n31 G_sink_dn.t16 2.7305
R1212 G_sink_dn.n31 G_sink_dn.n30 2.7305
R1213 G_sink_dn.n29 G_sink_dn.t23 2.7305
R1214 G_sink_dn.n29 G_sink_dn.n28 2.7305
R1215 G_sink_dn.n3 G_sink_dn.t6 2.7305
R1216 G_sink_dn.n3 G_sink_dn.n2 2.7305
R1217 G_sink_dn.n1 G_sink_dn.t12 2.7305
R1218 G_sink_dn.n1 G_sink_dn.n0 2.7305
R1219 G_sink_dn.n18 G_sink_dn.n17 2.3365
R1220 G_sink_dn.n25 G_sink_dn.n24 2.3365
R1221 G_sink_dn.n34 G_sink_dn.n33 2.3365
R1222 G_sink_dn.n36 G_sink_dn.n35 2.3365
R1223 G_sink_dn G_sink_dn.n37 0.496
R1224 SD0_1.n18 SD0_1.n3 3.41579
R1225 SD0_1.n13 SD0_1.n10 3.00682
R1226 SD0_1.n24 SD0_1.n1 3.0043
R1227 SD0_1.n15 SD0_1.n5 3.00256
R1228 SD0_1.n27 SD0_1.t12 2.7305
R1229 SD0_1.n27 SD0_1.n26 2.7305
R1230 SD0_1.n3 SD0_1.t13 2.7305
R1231 SD0_1.n3 SD0_1.n2 2.7305
R1232 SD0_1.n20 SD0_1.t7 2.7305
R1233 SD0_1.n20 SD0_1.n19 2.7305
R1234 SD0_1.n7 SD0_1.t14 2.7305
R1235 SD0_1.n7 SD0_1.n6 2.7305
R1236 SD0_1.n12 SD0_1.t3 2.7305
R1237 SD0_1.n12 SD0_1.n11 2.7305
R1238 SD0_1.n10 SD0_1.t9 2.7305
R1239 SD0_1.n10 SD0_1.n9 2.7305
R1240 SD0_1.n5 SD0_1.t5 2.7305
R1241 SD0_1.n5 SD0_1.n4 2.7305
R1242 SD0_1.n1 SD0_1.t1 2.7305
R1243 SD0_1.n1 SD0_1.n0 2.7305
R1244 SD0_1.n13 SD0_1.n12 2.56463
R1245 SD0_1.n22 SD0_1.n21 2.24419
R1246 SD0_1 SD0_1.n29 1.50504
R1247 SD0_1.n14 SD0_1.n8 1.4943
R1248 SD0_1.n8 SD0_1.n7 1.43801
R1249 SD0_1.n28 SD0_1.n27 1.43776
R1250 SD0_1.n21 SD0_1.n20 1.43749
R1251 SD0_1.n14 SD0_1.n13 0.603471
R1252 SD0_1.n23 SD0_1.n22 0.57715
R1253 SD0_1.n17 SD0_1.n16 0.576682
R1254 SD0_1.n16 SD0_1.n15 0.0255633
R1255 SD0_1.n24 SD0_1.n23 0.0244241
R1256 SD0_1.n18 SD0_1.n17 0.0180472
R1257 SD0_1.n22 SD0_1.n18 0.0146295
R1258 SD0_1.n15 SD0_1.n14 0.0145334
R1259 SD0_1 SD0_1.n24 0.00391772
R1260 SD0_1.n28 SD0_1.n25 0.00358243
R1261 SD0_1.n29 SD0_1.n28 0.00181665
R1262 SD2_1.n68 SD2_1.n1 3.5764
R1263 SD2_1.n26 SD2_1.n25 3.18472
R1264 SD2_1.n30 SD2_1.n17 3.17597
R1265 SD2_1.n39 SD2_1.n15 3.17588
R1266 SD2_1.n41 SD2_1.n13 3.17454
R1267 SD2_1.n44 SD2_1.n9 3.17453
R1268 SD2_1.n56 SD2_1.n5 3.1741
R1269 SD2_1.n27 SD2_1.n21 3.17375
R1270 SD2_1.n72 SD2_1.n69 3.17335
R1271 SD2_1.n50 SD2_1.n7 3.17318
R1272 SD2_1.n65 SD2_1.n3 3.17219
R1273 SD2_1.n74 SD2_1.n73 3.01386
R1274 SD2_1.n42 SD2_1.n11 2.93559
R1275 SD2_1.n26 SD2_1.n23 2.56337
R1276 SD2_1.n28 SD2_1.n19 2.56302
R1277 SD2_1.n75 SD2_1.n74 2.25469
R1278 SD2_1.n64 SD2_1.n63 2.24989
R1279 SD2_1.n38 SD2_1.n37 2.24988
R1280 SD2_1.n34 SD2_1.n33 2.24511
R1281 SD2_1.n48 SD2_1.n47 2.24483
R1282 SD2_1.n60 SD2_1.n59 2.24483
R1283 SD2_1.n54 SD2_1.n53 2.24455
R1284 SD2_1.n62 SD2_1.n61 1.74882
R1285 SD2_1.n58 SD2_1.n57 1.74881
R1286 SD2_1.n46 SD2_1.n45 1.74881
R1287 SD2_1.n36 SD2_1.n35 1.74881
R1288 SD2_1.n19 SD2_1.n18 1.74881
R1289 SD2_1.n32 SD2_1.n31 1.73459
R1290 SD2_1.n52 SD2_1.t26 1.6385
R1291 SD2_1.n52 SD2_1.n51 1.6385
R1292 SD2_1.n11 SD2_1.t30 1.6385
R1293 SD2_1.n11 SD2_1.n10 1.6385
R1294 SD2_1.n23 SD2_1.t29 1.6385
R1295 SD2_1.n23 SD2_1.n22 1.6385
R1296 SD2_1.n25 SD2_1.t15 1.6385
R1297 SD2_1.n25 SD2_1.n24 1.6385
R1298 SD2_1.n21 SD2_1.t35 1.6385
R1299 SD2_1.n21 SD2_1.n20 1.6385
R1300 SD2_1.n17 SD2_1.t3 1.6385
R1301 SD2_1.n17 SD2_1.n16 1.6385
R1302 SD2_1.n15 SD2_1.t32 1.6385
R1303 SD2_1.n15 SD2_1.n14 1.6385
R1304 SD2_1.n13 SD2_1.t17 1.6385
R1305 SD2_1.n13 SD2_1.n12 1.6385
R1306 SD2_1.n9 SD2_1.t28 1.6385
R1307 SD2_1.n9 SD2_1.n8 1.6385
R1308 SD2_1.n7 SD2_1.t9 1.6385
R1309 SD2_1.n7 SD2_1.n6 1.6385
R1310 SD2_1.n5 SD2_1.t33 1.6385
R1311 SD2_1.n5 SD2_1.n4 1.6385
R1312 SD2_1.n3 SD2_1.t18 1.6385
R1313 SD2_1.n3 SD2_1.n2 1.6385
R1314 SD2_1.n1 SD2_1.t27 1.6385
R1315 SD2_1.n1 SD2_1.n0 1.6385
R1316 SD2_1.n71 SD2_1.n70 1.5755
R1317 SD2_1.n32 SD2_1.t34 1.48949
R1318 SD2_1.n58 SD2_1.t7 1.47237
R1319 SD2_1.n46 SD2_1.t4 1.47237
R1320 SD2_1.n36 SD2_1.t6 1.47237
R1321 SD2_1.n19 SD2_1.t10 1.47237
R1322 SD2_1.n62 SD2_1.t31 1.47236
R1323 SD2_1.n53 SD2_1.n52 1.44171
R1324 SD2_1.n73 SD2_1.t13 1.28985
R1325 SD2_1.n63 SD2_1.n62 1.07211
R1326 SD2_1.n37 SD2_1.n36 1.07199
R1327 SD2_1.n47 SD2_1.n46 1.07199
R1328 SD2_1.n59 SD2_1.n58 1.07199
R1329 SD2_1.n33 SD2_1.n32 1.07053
R1330 SD2_1.n29 SD2_1.n28 0.626751
R1331 SD2_1.n27 SD2_1.n26 0.622777
R1332 SD2_1.n43 SD2_1.n42 0.612573
R1333 SD2_1.n55 SD2_1.n54 0.606132
R1334 SD2_1.n64 SD2_1.n60 0.605265
R1335 SD2_1.n38 SD2_1.n34 0.603102
R1336 SD2_1.n49 SD2_1.n48 0.601395
R1337 SD2_1.n67 SD2_1.n66 0.593475
R1338 SD2_1.n41 SD2_1.n40 0.584536
R1339 SD2_1.n73 SD2_1.n72 0.31735
R1340 SD2_1.n72 SD2_1.n71 0.0635
R1341 SD2_1.n28 SD2_1.n27 0.0264198
R1342 SD2_1.n66 SD2_1.n65 0.0249444
R1343 SD2_1.n40 SD2_1.n39 0.024125
R1344 SD2_1.n42 SD2_1.n41 0.0174125
R1345 SD2_1.n34 SD2_1.n30 0.0172816
R1346 SD2_1.n48 SD2_1.n44 0.0167161
R1347 SD2_1.n54 SD2_1.n50 0.0161504
R1348 SD2_1.n60 SD2_1.n56 0.0144661
R1349 SD2_1.n68 SD2_1.n67 0.0061962
R1350 SD2_1.n39 SD2_1.n38 0.00549888
R1351 SD2_1.n74 SD2_1.n69 0.00543151
R1352 SD2_1.n56 SD2_1.n55 0.005
R1353 SD2_1.n75 SD2_1.n68 0.00441168
R1354 SD2_1.n65 SD2_1.n64 0.00433224
R1355 SD2_1 SD2_1.n75 0.00328222
R1356 SD2_1.n30 SD2_1.n29 0.00275
R1357 SD2_1.n44 SD2_1.n43 0.00275
R1358 SD2_1.n50 SD2_1.n49 0.00275
R1359 G1_1.n5 G1_1.n2 103.823
R1360 G1_1.n54 G1_1.n53 103.823
R1361 G1_1.n4 G1_1.n3 103.823
R1362 G1_1.n55 G1_1.n52 103.823
R1363 G1_1.n2 G1_1.t76 32.8424
R1364 G1_1.n53 G1_1.t73 32.8424
R1365 G1_1.n117 G1_1.t12 31.6661
R1366 G1_1.n33 G1_1.t22 31.5165
R1367 G1_1.n5 G1_1.n4 21.0894
R1368 G1_1.n55 G1_1.n54 21.0894
R1369 G1_1.n116 G1_1.t18 15.4035
R1370 G1_1.n117 G1_1.t4 15.4035
R1371 G1_1.n69 G1_1.t16 15.1845
R1372 G1_1.n70 G1_1.t20 15.1845
R1373 G1_1.n33 G1_1.t14 15.0385
R1374 G1_1.n34 G1_1.t38 15.0385
R1375 G1_1.n79 G1_1.t8 15.0385
R1376 G1_1.n81 G1_1.t32 15.0385
R1377 G1_1.n45 G1_1.t6 14.8925
R1378 G1_1.n47 G1_1.t30 14.8925
R1379 G1_1.n65 G1_1.t24 12.0455
R1380 G1_1.n64 G1_1.t36 12.0455
R1381 G1_1.n89 G1_1.t26 11.9725
R1382 G1_1.n88 G1_1.t0 11.9725
R1383 G1_1.n39 G1_1.t34 11.8995
R1384 G1_1.n38 G1_1.t10 11.8995
R1385 G1_1.n2 G1_1.t70 11.7535
R1386 G1_1.n53 G1_1.t79 11.7535
R1387 G1_1.n54 G1_1.t75 11.7535
R1388 G1_1.n4 G1_1.t74 11.7535
R1389 G1_1.n3 G1_1.t67 11.7535
R1390 G1_1.n52 G1_1.t72 11.7535
R1391 G1_1.n74 G1_1.t2 11.6805
R1392 G1_1.n73 G1_1.t28 11.6805
R1393 G1_1.n57 G1_1.t62 8.14629
R1394 G1_1.n0 G1_1.t61 8.14629
R1395 G1_1.n5 G1_1.n1 8.0005
R1396 G1_1.n118 G1_1.n116 7.97643
R1397 G1_1.n66 G1_1.n64 7.49604
R1398 G1_1.n35 G1_1.n34 7.2359
R1399 G1_1.n90 G1_1.n88 6.91289
R1400 G1_1.n71 G1_1.n69 6.84014
R1401 G1_1.n75 G1_1.n74 6.80135
R1402 G1_1.n40 G1_1.n39 6.66015
R1403 G1_1.n71 G1_1.n70 6.57708
R1404 G1_1.n40 G1_1.n38 6.40401
R1405 G1_1.n90 G1_1.n89 6.26687
R1406 G1_1.n35 G1_1.n33 5.94386
R1407 G1_1.n75 G1_1.n73 5.92785
R1408 G1_1.n61 G1_1.n60 5.92398
R1409 G1_1.n125 G1_1.n124 5.90903
R1410 G1_1.n118 G1_1.n117 5.81346
R1411 G1_1.n66 G1_1.n65 5.80139
R1412 G1_1.n30 G1_1.n23 5.1485
R1413 G1_1.n114 G1_1.t46 5.1485
R1414 G1_1.n32 G1_1.n31 4.4205
R1415 G1_1.n115 G1_1.t13 4.4205
R1416 G1_1.n46 G1_1.n45 4.19007
R1417 G1_1.n80 G1_1.n79 4.07041
R1418 G1_1.n82 G1_1.n81 4.07041
R1419 G1_1.n121 G1_1.n90 4.0005
R1420 G1_1.n119 G1_1.n118 4.0005
R1421 G1_1.n36 G1_1.n35 4.0005
R1422 G1_1.n41 G1_1.n40 4.0005
R1423 G1_1.n67 G1_1.n66 4.0005
R1424 G1_1.n72 G1_1.n71 4.0005
R1425 G1_1.n76 G1_1.n75 4.0005
R1426 G1_1.n48 G1_1.n47 3.8092
R1427 G1_1.n113 G1_1.n94 3.54572
R1428 G1_1.n111 G1_1.n98 3.54572
R1429 G1_1.n109 G1_1.n102 3.54572
R1430 G1_1.n107 G1_1.n106 3.54572
R1431 G1_1.n29 G1_1.n25 3.54572
R1432 G1_1.n58 G1_1.n56 3.53093
R1433 G1_1.n28 G1_1.n27 3.5105
R1434 G1_1.n108 G1_1.n104 3.5105
R1435 G1_1.n110 G1_1.n100 3.5105
R1436 G1_1.n112 G1_1.n96 3.5105
R1437 G1_1.n58 G1_1.n57 3.50535
R1438 G1_1.n1 G1_1.n0 3.50535
R1439 G1_1.n120 G1_1.n92 3.02311
R1440 G1_1.n68 G1_1.n14 3.01724
R1441 G1_1.n124 G1_1.n10 3.01333
R1442 G1_1.n37 G1_1.n22 3.01333
R1443 G1_1.n44 G1_1.n18 3.00941
R1444 G1_1.n63 G1_1.n16 2.93311
R1445 G1_1.n122 G1_1.n87 2.93115
R1446 G1_1.n42 G1_1.n20 2.9292
R1447 G1_1.n77 G1_1.n12 2.92333
R1448 G1_1.n8 G1_1.n7 2.88455
R1449 G1_1.n60 G1_1.n59 2.88451
R1450 G1_1.n51 G1_1.n50 2.66717
R1451 G1_1.n85 G1_1.n84 2.66717
R1452 G1_1.n83 G1_1.n82 2.51997
R1453 G1_1.n84 G1_1.n80 2.45537
R1454 G1_1.n32 G1_1.n30 2.44296
R1455 G1_1.n50 G1_1.n46 2.41267
R1456 G1_1.n49 G1_1.n48 2.41267
R1457 G1_1.n115 G1_1.n114 2.14942
R1458 G1_1.n6 G1_1.n5 1.9715
R1459 G1_1.n10 G1_1.t9 1.8205
R1460 G1_1.n10 G1_1.n9 1.8205
R1461 G1_1.n87 G1_1.t1 1.8205
R1462 G1_1.n87 G1_1.n86 1.8205
R1463 G1_1.n92 G1_1.t19 1.8205
R1464 G1_1.n92 G1_1.n91 1.8205
R1465 G1_1.n22 G1_1.t15 1.8205
R1466 G1_1.n22 G1_1.n21 1.8205
R1467 G1_1.n20 G1_1.t11 1.8205
R1468 G1_1.n20 G1_1.n19 1.8205
R1469 G1_1.n18 G1_1.t7 1.8205
R1470 G1_1.n18 G1_1.n17 1.8205
R1471 G1_1.n16 G1_1.t37 1.8205
R1472 G1_1.n16 G1_1.n15 1.8205
R1473 G1_1.n14 G1_1.t17 1.8205
R1474 G1_1.n14 G1_1.n13 1.8205
R1475 G1_1.n12 G1_1.t29 1.8205
R1476 G1_1.n12 G1_1.n11 1.8205
R1477 G1_1.n27 G1_1.t45 1.6385
R1478 G1_1.n27 G1_1.n26 1.6385
R1479 G1_1.n104 G1_1.t58 1.6385
R1480 G1_1.n104 G1_1.n103 1.6385
R1481 G1_1.n100 G1_1.t54 1.6385
R1482 G1_1.n100 G1_1.n99 1.6385
R1483 G1_1.n96 G1_1.t40 1.6385
R1484 G1_1.n96 G1_1.n95 1.6385
R1485 G1_1.n94 G1_1.t49 1.6385
R1486 G1_1.n94 G1_1.n93 1.6385
R1487 G1_1.n98 G1_1.t44 1.6385
R1488 G1_1.n98 G1_1.n97 1.6385
R1489 G1_1.n102 G1_1.t48 1.6385
R1490 G1_1.n102 G1_1.n101 1.6385
R1491 G1_1.n106 G1_1.t43 1.6385
R1492 G1_1.n106 G1_1.n105 1.6385
R1493 G1_1.n25 G1_1.t47 1.6385
R1494 G1_1.n25 G1_1.n24 1.6385
R1495 G1_1.n119 G1_1.n115 1.14702
R1496 G1_1.n36 G1_1.n32 1.14051
R1497 G1_1.n56 G1_1.n55 0.995675
R1498 G1_1.n121 G1_1.n120 0.692144
R1499 G1_1.n41 G1_1.n37 0.686551
R1500 G1_1.n68 G1_1.n67 0.660185
R1501 G1_1.n76 G1_1.n72 0.659391
R1502 G1_1.n63 G1_1.n62 0.656587
R1503 G1_1.n123 G1_1.n122 0.651709
R1504 G1_1.n43 G1_1.n42 0.651372
R1505 G1_1.n78 G1_1.n77 0.648302
R1506 G1_1.n30 G1_1.n29 0.565423
R1507 G1_1.n29 G1_1.n28 0.565423
R1508 G1_1.n108 G1_1.n107 0.565423
R1509 G1_1.n109 G1_1.n108 0.565423
R1510 G1_1.n110 G1_1.n109 0.565423
R1511 G1_1.n111 G1_1.n110 0.565423
R1512 G1_1.n112 G1_1.n111 0.565423
R1513 G1_1.n113 G1_1.n112 0.565423
R1514 G1_1.n114 G1_1.n113 0.565423
R1515 G1_1.n7 G1_1.n6 0.3655
R1516 G1_1.n50 G1_1.n49 0.127457
R1517 G1_1.n84 G1_1.n83 0.0651018
R1518 G1_1.n124 G1_1.n123 0.0345777
R1519 G1_1.n85 G1_1.n78 0.0337039
R1520 G1_1.n62 G1_1.n61 0.0330714
R1521 G1_1.n44 G1_1.n43 0.0313571
R1522 G1_1.n120 G1_1.n119 0.0151939
R1523 G1_1.n67 G1_1.n63 0.0106739
R1524 G1_1.n37 G1_1.n36 0.00923786
R1525 G1_1.n77 G1_1.n76 0.00575
R1526 G1_1 G1_1.n125 0.0055
R1527 G1_1.n122 G1_1.n121 0.00437931
R1528 G1_1.n60 G1_1.n58 0.0025
R1529 G1_1.n72 G1_1.n68 0.00228218
R1530 G1_1.n8 G1_1.n1 0.00228158
R1531 G1_1.n51 G1_1.n44 0.00221429
R1532 G1_1.n61 G1_1.n51 0.00221429
R1533 G1_1.n42 G1_1.n41 0.00203846
R1534 G1_1.n125 G1_1.n8 0.0017181
R1535 G1_1.n124 G1_1.n85 0.00137379
R1536 G_sink_up.n22 G_sink_up.n18 132.008
R1537 G_sink_up.n0 G_sink_up.t29 116.525
R1538 G_sink_up.n48 G_sink_up.n47 106.159
R1539 G_sink_up.n2 G_sink_up.n1 103.823
R1540 G_sink_up.n6 G_sink_up.n5 103.823
R1541 G_sink_up.n17 G_sink_up.n16 103.823
R1542 G_sink_up.n24 G_sink_up.n23 103.823
R1543 G_sink_up.n5 G_sink_up.n2 49.2755
R1544 G_sink_up.n16 G_sink_up.t27 33.7914
R1545 G_sink_up.n27 G_sink_up.n24 22.4014
R1546 G_sink_up.n1 G_sink_up.n0 21.0894
R1547 G_sink_up.n47 G_sink_up.n6 21.0894
R1548 G_sink_up.n18 G_sink_up.n17 21.0894
R1549 G_sink_up.n23 G_sink_up.n22 21.0894
R1550 G_sink_up.n0 G_sink_up.t30 12.7025
R1551 G_sink_up.n1 G_sink_up.t31 12.7025
R1552 G_sink_up.n2 G_sink_up.t35 12.7025
R1553 G_sink_up.n6 G_sink_up.t14 12.7025
R1554 G_sink_up.n16 G_sink_up.t33 12.7025
R1555 G_sink_up.n17 G_sink_up.t32 12.7025
R1556 G_sink_up.n18 G_sink_up.t36 12.7025
R1557 G_sink_up.n23 G_sink_up.t12 12.7025
R1558 G_sink_up.n24 G_sink_up.t24 12.7025
R1559 G_sink_up.n4 G_sink_up.t22 10.3665
R1560 G_sink_up.n21 G_sink_up.t18 10.3665
R1561 G_sink_up.n48 G_sink_up.t20 10.3665
R1562 G_sink_up.n4 G_sink_up.n3 10.2268
R1563 G_sink_up.n25 G_sink_up.t16 9.14366
R1564 G_sink_up.n7 G_sink_up.t10 7.9575
R1565 G_sink_up.n21 G_sink_up.n20 7.48719
R1566 G_sink_up.n49 G_sink_up.t21 6.05659
R1567 G_sink_up.n30 G_sink_up.t1 4.5505
R1568 G_sink_up.n30 G_sink_up.n29 4.5505
R1569 G_sink_up.n32 G_sink_up.t3 4.5505
R1570 G_sink_up.n32 G_sink_up.n31 4.5505
R1571 G_sink_up.n34 G_sink_up.t0 4.5505
R1572 G_sink_up.n34 G_sink_up.n33 4.5505
R1573 G_sink_up.n36 G_sink_up.t2 4.5505
R1574 G_sink_up.n36 G_sink_up.n35 4.5505
R1575 G_sink_up.n41 G_sink_up.t4 4.5505
R1576 G_sink_up.n41 G_sink_up.n40 4.5505
R1577 G_sink_up.n49 G_sink_up.n48 4.15442
R1578 G_sink_up.n37 G_sink_up.n36 3.98849
R1579 G_sink_up.n44 G_sink_up.n43 3.83414
R1580 G_sink_up.n46 G_sink_up.n45 3.50535
R1581 G_sink_up.n14 G_sink_up.n13 3.46045
R1582 G_sink_up.n11 G_sink_up.n10 3.45688
R1583 G_sink_up.n43 G_sink_up.n42 3.13411
R1584 G_sink_up.n39 G_sink_up.n30 2.80398
R1585 G_sink_up.n38 G_sink_up.n32 2.80398
R1586 G_sink_up.n37 G_sink_up.n34 2.80398
R1587 G_sink_up.n42 G_sink_up.n41 2.78907
R1588 G_sink_up.n13 G_sink_up.t25 2.7305
R1589 G_sink_up.n13 G_sink_up.n12 2.7305
R1590 G_sink_up.n20 G_sink_up.t19 2.7305
R1591 G_sink_up.n20 G_sink_up.n19 2.7305
R1592 G_sink_up.n10 G_sink_up.t15 2.7305
R1593 G_sink_up.n10 G_sink_up.n9 2.7305
R1594 G_sink_up.n5 G_sink_up.n4 2.3365
R1595 G_sink_up.n22 G_sink_up.n21 2.3365
R1596 G_sink_up.n8 G_sink_up.n7 2.2635
R1597 G_sink_up.n43 G_sink_up.n28 2.2505
R1598 G_sink_up.n28 G_sink_up.n27 1.78431
R1599 G_sink_up.n38 G_sink_up.n37 1.18502
R1600 G_sink_up.n39 G_sink_up.n38 1.18502
R1601 G_sink_up.n26 G_sink_up.n25 1.18043
R1602 G_sink_up.n42 G_sink_up.n39 1.1582
R1603 G_sink_up.n46 G_sink_up.n8 1.13829
R1604 G_sink_up.n47 G_sink_up.n46 1.06529
R1605 G_sink_up.n27 G_sink_up.n26 0.465838
R1606 G_sink_up G_sink_up.n49 0.207891
R1607 G_sink_up.n45 G_sink_up.n11 0.0315
R1608 G_sink_up.n15 G_sink_up.n14 0.0227581
R1609 G_sink_up.n28 G_sink_up.n15 0.00569231
R1610 G_sink_up.n45 G_sink_up.n44 0.0035
R1611 SD1_1.n28 SD1_1.t1 4.5505
R1612 SD1_1.n28 SD1_1.n27 4.5505
R1613 SD1_1.n1 SD1_1.t12 4.5505
R1614 SD1_1.n1 SD1_1.n0 4.5505
R1615 SD1_1.n3 SD1_1.t9 4.5505
R1616 SD1_1.n3 SD1_1.n2 4.5505
R1617 SD1_1.n5 SD1_1.t17 4.5505
R1618 SD1_1.n5 SD1_1.n4 4.5505
R1619 SD1_1.n7 SD1_1.t7 4.5505
R1620 SD1_1.n7 SD1_1.n6 4.5505
R1621 SD1_1.n9 SD1_1.t11 4.5505
R1622 SD1_1.n9 SD1_1.n8 4.5505
R1623 SD1_1.n11 SD1_1.t8 4.5505
R1624 SD1_1.n11 SD1_1.n10 4.5505
R1625 SD1_1.n13 SD1_1.t14 4.5505
R1626 SD1_1.n13 SD1_1.n12 4.5505
R1627 SD1_1.n15 SD1_1.t0 4.5505
R1628 SD1_1.n15 SD1_1.n14 4.5505
R1629 SD1_1.n17 SD1_1.t10 4.5505
R1630 SD1_1.n17 SD1_1.n16 4.5505
R1631 SD1_1.n18 SD1_1.n17 3.17149
R1632 SD1_1.n19 SD1_1.n13 2.77857
R1633 SD1_1.n25 SD1_1.n1 2.54881
R1634 SD1_1.n18 SD1_1.n15 2.54881
R1635 SD1_1.n24 SD1_1.n3 2.54872
R1636 SD1_1.n23 SD1_1.n5 2.54872
R1637 SD1_1.n22 SD1_1.n7 2.54872
R1638 SD1_1.n20 SD1_1.n11 2.54872
R1639 SD1_1.n21 SD1_1.n9 2.54854
R1640 SD1_1.n31 SD1_1.n30 2.25795
R1641 SD1_1.n29 SD1_1.n26 2.2439
R1642 SD1_1.n29 SD1_1.n28 1.65397
R1643 SD1_1.n19 SD1_1.n18 0.635915
R1644 SD1_1.n24 SD1_1.n23 0.627793
R1645 SD1_1.n21 SD1_1.n20 0.626983
R1646 SD1_1.n25 SD1_1.n24 0.623305
R1647 SD1_1.n22 SD1_1.n21 0.622387
R1648 SD1_1.n23 SD1_1.n22 0.621579
R1649 SD1_1.n20 SD1_1.n19 0.614074
R1650 SD1_1.n26 SD1_1.n25 0.609182
R1651 SD1_1.n31 SD1_1.n26 0.0151956
R1652 SD1_1.n30 SD1_1.n29 0.010363
R1653 SD1_1 SD1_1.n31 0.00163924
R1654 G_source_dn.n47 G_source_dn.t20 34.3024
R1655 G_source_dn.n48 G_source_dn.t14 10.8775
R1656 G_source_dn.n45 G_source_dn.t18 10.8775
R1657 G_source_dn.n18 G_source_dn.t12 10.8775
R1658 G_source_dn.n15 G_source_dn.t22 10.8775
R1659 G_source_dn.n12 G_source_dn.t16 10.8775
R1660 G_source_dn.n27 G_source_dn.t10 9.65117
R1661 G_source_dn.n23 G_source_dn.t8 9.65117
R1662 G_source_dn.n36 G_source_dn.n35 6.96833
R1663 G_source_dn.n39 G_source_dn.t1 6.17107
R1664 G_source_dn.n13 G_source_dn.n12 4.15702
R1665 G_source_dn.n16 G_source_dn.n15 4.0005
R1666 G_source_dn.n19 G_source_dn.n18 4.0005
R1667 G_source_dn.n46 G_source_dn.n45 4.0005
R1668 G_source_dn.n49 G_source_dn.n48 4.0005
R1669 G_source_dn.n24 G_source_dn.n23 3.51942
R1670 G_source_dn.n28 G_source_dn.n27 3.51942
R1671 G_source_dn.n38 G_source_dn.n30 3.46159
R1672 G_source_dn.n36 G_source_dn.n34 3.46159
R1673 G_source_dn.n37 G_source_dn.n32 3.44007
R1674 G_source_dn.n40 G_source_dn.n39 3.34436
R1675 G_source_dn.n1 G_source_dn.t15 3.03383
R1676 G_source_dn.n1 G_source_dn.n0 3.03383
R1677 G_source_dn.n11 G_source_dn.t17 3.03383
R1678 G_source_dn.n11 G_source_dn.n10 3.03383
R1679 G_source_dn.n9 G_source_dn.t13 3.03383
R1680 G_source_dn.n9 G_source_dn.n8 3.03383
R1681 G_source_dn.n3 G_source_dn.t11 3.03383
R1682 G_source_dn.n3 G_source_dn.n2 3.03383
R1683 G_source_dn.n21 G_source_dn.n7 2.8741
R1684 G_source_dn.n42 G_source_dn.n5 2.8741
R1685 G_source_dn.n41 G_source_dn.n40 2.84271
R1686 G_source_dn.n50 G_source_dn.n1 2.80398
R1687 G_source_dn.n13 G_source_dn.n11 2.80398
R1688 G_source_dn.n20 G_source_dn.n9 2.80398
R1689 G_source_dn.n43 G_source_dn.n3 2.80398
R1690 G_source_dn.n32 G_source_dn.t5 2.7305
R1691 G_source_dn.n32 G_source_dn.n31 2.7305
R1692 G_source_dn.n30 G_source_dn.t3 2.7305
R1693 G_source_dn.n30 G_source_dn.n29 2.7305
R1694 G_source_dn.n34 G_source_dn.t7 2.7305
R1695 G_source_dn.n34 G_source_dn.n33 2.7305
R1696 G_source_dn.n48 G_source_dn.n47 2.3365
R1697 G_source_dn.n45 G_source_dn.n44 2.3365
R1698 G_source_dn.n18 G_source_dn.n17 2.3365
R1699 G_source_dn.n15 G_source_dn.n14 2.3365
R1700 G_source_dn.n5 G_source_dn.n4 2.1175
R1701 G_source_dn.n7 G_source_dn.n6 2.1175
R1702 G_source_dn G_source_dn.n50 1.15876
R1703 G_source_dn.n19 G_source_dn.n16 1.1118
R1704 G_source_dn.n49 G_source_dn.n46 1.1118
R1705 G_source_dn.n26 G_source_dn.n25 1.0508
R1706 G_source_dn.n37 G_source_dn.n36 0.798761
R1707 G_source_dn.n38 G_source_dn.n37 0.798761
R1708 G_source_dn.n39 G_source_dn.n38 0.710717
R1709 G_source_dn.n16 G_source_dn.n13 0.157022
R1710 G_source_dn.n20 G_source_dn.n19 0.157022
R1711 G_source_dn.n46 G_source_dn.n43 0.157022
R1712 G_source_dn.n21 G_source_dn.n20 0.143676
R1713 G_source_dn.n43 G_source_dn.n42 0.142676
R1714 G_source_dn.n50 G_source_dn.n49 0.1025
R1715 G_source_dn.n25 G_source_dn.n24 0.0315
R1716 G_source_dn.n28 G_source_dn.n26 0.0305
R1717 G_source_dn.n22 G_source_dn.n21 0.0117741
R1718 G_source_dn.n42 G_source_dn.n41 0.0117741
R1719 G_source_dn.n41 G_source_dn.n28 0.0045
R1720 G_source_dn.n24 G_source_dn.n22 0.0035
R1721 G_source_up.n13 G_source_up.n12 27.2758
R1722 G_source_up.n21 G_source_up.n20 27.2758
R1723 G_source_up.n29 G_source_up.n28 27.2758
R1724 G_source_up.n6 G_source_up.t4 10.4831
R1725 G_source_up.n34 G_source_up.t14 10.1908
R1726 G_source_up.n12 G_source_up.t6 7.5925
R1727 G_source_up.n13 G_source_up.t0 7.5925
R1728 G_source_up.n20 G_source_up.t12 7.5925
R1729 G_source_up.n21 G_source_up.t10 7.5925
R1730 G_source_up.n28 G_source_up.t8 7.5925
R1731 G_source_up.n29 G_source_up.t2 7.5925
R1732 G_source_up.n7 G_source_up.n6 4.0005
R1733 G_source_up.n11 G_source_up.n10 4.0005
R1734 G_source_up.n15 G_source_up.n14 4.0005
R1735 G_source_up.n19 G_source_up.n18 4.0005
R1736 G_source_up.n23 G_source_up.n22 4.0005
R1737 G_source_up.n27 G_source_up.n26 4.0005
R1738 G_source_up.n33 G_source_up.n30 4.0005
R1739 G_source_up.n35 G_source_up.n34 4.0005
R1740 G_source_up.n37 G_source_up.t17 3.03383
R1741 G_source_up.n37 G_source_up.n36 3.03383
R1742 G_source_up.n25 G_source_up.t23 3.03383
R1743 G_source_up.n25 G_source_up.n24 3.03383
R1744 G_source_up.n1 G_source_up.t11 3.03383
R1745 G_source_up.n1 G_source_up.n0 3.03383
R1746 G_source_up.n17 G_source_up.t16 3.03383
R1747 G_source_up.n17 G_source_up.n16 3.03383
R1748 G_source_up.n3 G_source_up.t1 3.03383
R1749 G_source_up.n3 G_source_up.n2 3.03383
R1750 G_source_up.n9 G_source_up.t19 3.03383
R1751 G_source_up.n9 G_source_up.n8 3.03383
R1752 G_source_up.n5 G_source_up.t5 3.03383
R1753 G_source_up.n5 G_source_up.n4 3.03383
R1754 G_source_up.n32 G_source_up.t3 3.03383
R1755 G_source_up.n32 G_source_up.n31 3.03383
R1756 G_source_up.n26 G_source_up.n25 2.84924
R1757 G_source_up.n23 G_source_up.n1 2.84924
R1758 G_source_up.n18 G_source_up.n17 2.84924
R1759 G_source_up.n15 G_source_up.n3 2.84924
R1760 G_source_up.n10 G_source_up.n9 2.84924
R1761 G_source_up.n33 G_source_up.n32 2.84924
R1762 G_source_up.n7 G_source_up.n5 2.84872
R1763 G_source_up.n38 G_source_up.n37 2.6005
R1764 G_source_up.n12 G_source_up.n11 2.59881
R1765 G_source_up.n14 G_source_up.n13 2.59881
R1766 G_source_up.n20 G_source_up.n19 2.59881
R1767 G_source_up.n22 G_source_up.n21 2.59881
R1768 G_source_up.n28 G_source_up.n27 2.59881
R1769 G_source_up.n30 G_source_up.n29 2.59881
R1770 G_source_up G_source_up.n38 0.959196
R1771 G_source_up.n35 G_source_up.n33 0.732411
R1772 G_source_up.n10 G_source_up.n7 0.728327
R1773 G_source_up.n26 G_source_up.n23 0.724527
R1774 G_source_up.n18 G_source_up.n15 0.720586
R1775 G_source_up.n38 G_source_up.n35 0.249235
C0 G1_2 SD1_1 0.376f
C1 SD0_1 VDD 0.0216f
C2 G1_1 VDD 9.89f
C3 G1_1 ITAIL 0.618f
C4 G1_2 G2_1 0.00451f
C5 G_source_up G_source_dn 2.18f
C6 G1_1 SD2_1 2.49f
C7 ITAIL VDD 0.207f
C8 G_source_dn G_sink_up 0.408f
C9 SD2_1 VDD 0.0868f
C10 ITAIL SD2_1 1.02f
C11 G_sink_up G_sink_dn 1.71f
C12 G_source_dn SD0_1 0.852f
C13 G_source_up G1_2 4.84e-20
C14 G_sink_dn SD0_1 0.16f
C15 G_sink_up G1_2 0.556f
C16 G_source_up SD1_1 9.69e-20
C17 G_source_dn G1_1 4.33e-19
C18 G_sink_up SD1_1 1.28f
C19 G_sink_dn G1_1 4.2e-19
C20 SD0_1 G1_2 0.00621f
C21 G_source_dn VDD 1.83f
C22 G1_2 G1_1 4.36f
C23 SD0_1 SD1_1 0.0712f
C24 G_sink_dn VDD 0.00582f
C25 G1_2 ITAIL 0.127f
C26 G1_1 SD1_1 0.351f
C27 G1_2 VDD 13.9f
C28 G1_1 G2_1 0.874f
C29 G1_2 SD2_1 0.118f
C30 SD1_1 VDD 0.848f
C31 G_source_up G_sink_up 0.0161f
C32 G2_1 VDD 0.00603f
C33 ITAIL G2_1 5.61f
C34 G_source_up SD0_1 0.0116f
C35 G_source_dn G_sink_dn 0.302f
C36 G2_1 SD2_1 0.473f
C37 G_sink_up SD0_1 0.164f
C38 G_source_dn G1_2 0.00127f
C39 G_sink_up G1_1 0.246f
C40 G_sink_dn G1_2 0.0111f
C41 G_source_dn SD1_1 0.0263f
C42 G_source_up VDD 5.28f
C43 G_sink_dn SD1_1 0.0316f
C44 SD0_1 G1_1 0.00104f
C45 G_sink_up VDD 0.781f
.ends

