magic
tech gf180mcuC
magscale 1 10
timestamp 1694680735
<< nwell >>
rect -1809 6092 86 7070
rect -1809 6078 -1527 6092
rect -1450 6088 86 6092
rect -1450 6078 -302 6088
rect -1809 6075 -302 6078
rect -225 6075 86 6088
rect -1809 6032 86 6075
rect -1809 5947 -197 6032
rect -193 5947 86 6032
rect -1809 5664 86 5947
rect 360 6065 3868 6364
rect 360 5929 3861 6065
rect 360 5685 740 5929
rect -62 4310 4299 4347
rect -62 4136 298 4310
rect 4262 4136 4299 4310
rect -62 3627 4299 4136
rect -62 3565 1081 3627
rect 1086 3565 4299 3627
rect -62 3490 661 3565
rect 4261 3490 4299 3565
rect -62 2767 4299 3490
rect 159 2695 619 2767
rect 4262 2695 4299 2767
rect -62 2403 4299 2695
<< pwell >>
rect 480 5270 560 5350
rect 676 5063 757 5067
rect 773 5063 776 5067
rect 1956 5040 2387 5296
rect 1975 4687 2387 4943
<< psubdiff >>
rect -1778 5546 -1650 5562
rect -1778 5435 -1761 5546
rect -1667 5435 -1650 5546
rect -1778 5416 -1650 5435
rect -1511 5546 -1383 5562
rect -1511 5435 -1494 5546
rect -1400 5435 -1383 5546
rect -1511 5416 -1383 5435
rect -1301 5546 -1173 5562
rect -1301 5435 -1284 5546
rect -1190 5435 -1173 5546
rect -1301 5416 -1173 5435
rect -1091 5546 -963 5562
rect -1091 5435 -1074 5546
rect -980 5435 -963 5546
rect -1091 5416 -963 5435
rect -881 5546 -753 5562
rect -881 5435 -864 5546
rect -770 5435 -753 5546
rect -881 5416 -753 5435
rect -671 5546 -543 5562
rect -671 5435 -654 5546
rect -560 5435 -543 5546
rect -671 5416 -543 5435
rect -461 5546 -333 5562
rect -461 5435 -444 5546
rect -350 5435 -333 5546
rect -461 5416 -333 5435
rect -251 5546 -123 5562
rect -251 5435 -234 5546
rect -140 5435 -123 5546
rect -251 5416 -123 5435
rect 360 5549 488 5565
rect 360 5438 377 5549
rect 471 5438 488 5549
rect 360 5419 488 5438
rect 570 5549 698 5565
rect 570 5438 587 5549
rect 681 5438 698 5549
rect 570 5419 698 5438
rect 780 5549 908 5565
rect 780 5438 797 5549
rect 891 5438 908 5549
rect 780 5419 908 5438
rect 990 5549 1118 5565
rect 990 5438 1007 5549
rect 1101 5438 1118 5549
rect 990 5419 1118 5438
rect 1200 5549 1328 5565
rect 1200 5438 1217 5549
rect 1311 5438 1328 5549
rect 1200 5419 1328 5438
rect 1410 5549 1538 5565
rect 1410 5438 1427 5549
rect 1521 5438 1538 5549
rect 1410 5419 1538 5438
rect 1620 5549 1748 5565
rect 1620 5438 1637 5549
rect 1731 5438 1748 5549
rect 1620 5419 1748 5438
rect 1830 5549 1958 5565
rect 1830 5438 1847 5549
rect 1941 5438 1958 5549
rect 1830 5419 1958 5438
rect 2040 5549 2168 5565
rect 2040 5438 2057 5549
rect 2151 5438 2168 5549
rect 2040 5419 2168 5438
rect 2250 5549 2378 5565
rect 2250 5438 2267 5549
rect 2361 5438 2378 5549
rect 2250 5419 2378 5438
rect 2460 5549 2588 5565
rect 2460 5438 2477 5549
rect 2571 5438 2588 5549
rect 2460 5419 2588 5438
rect 2670 5549 2798 5565
rect 2670 5438 2687 5549
rect 2781 5438 2798 5549
rect 2670 5419 2798 5438
rect 2880 5549 3008 5565
rect 2880 5438 2897 5549
rect 2991 5438 3008 5549
rect 2880 5419 3008 5438
rect 3090 5549 3218 5565
rect 3090 5438 3107 5549
rect 3201 5438 3218 5549
rect 3090 5419 3218 5438
rect 3300 5549 3428 5565
rect 3300 5438 3317 5549
rect 3411 5438 3428 5549
rect 3300 5419 3428 5438
rect 3510 5549 3638 5565
rect 3510 5438 3527 5549
rect 3621 5438 3638 5549
rect 3510 5419 3638 5438
rect 3720 5549 3848 5565
rect 3720 5438 3737 5549
rect 3831 5438 3848 5549
rect 3720 5419 3848 5438
rect -1637 4545 -1509 4561
rect -1637 4434 -1620 4545
rect -1526 4434 -1509 4545
rect -1637 4415 -1509 4434
rect -1427 4545 -1299 4561
rect -1427 4434 -1410 4545
rect -1316 4434 -1299 4545
rect -1427 4415 -1299 4434
rect -1217 4545 -1089 4561
rect -1217 4434 -1200 4545
rect -1106 4434 -1089 4545
rect -1217 4415 -1089 4434
rect -1007 4545 -879 4561
rect -1007 4434 -990 4545
rect -896 4434 -879 4545
rect -1007 4415 -879 4434
rect -797 4545 -669 4561
rect -797 4434 -780 4545
rect -686 4434 -669 4545
rect -797 4415 -669 4434
rect -587 4545 -459 4561
rect -587 4434 -570 4545
rect -476 4434 -459 4545
rect -587 4415 -459 4434
rect -377 4545 -249 4561
rect -377 4434 -360 4545
rect -266 4434 -249 4545
rect -377 4415 -249 4434
rect -167 4545 -39 4561
rect -167 4434 -150 4545
rect -56 4434 -39 4545
rect -167 4415 -39 4434
rect 360 4530 488 4546
rect 360 4419 377 4530
rect 471 4419 488 4530
rect 360 4400 488 4419
rect 570 4530 698 4546
rect 570 4419 587 4530
rect 681 4419 698 4530
rect 570 4400 698 4419
rect 780 4530 908 4546
rect 780 4419 797 4530
rect 891 4419 908 4530
rect 780 4400 908 4419
rect 990 4530 1118 4546
rect 990 4419 1007 4530
rect 1101 4419 1118 4530
rect 990 4400 1118 4419
rect 1200 4530 1328 4546
rect 1200 4419 1217 4530
rect 1311 4419 1328 4530
rect 1200 4400 1328 4419
rect 1410 4530 1538 4546
rect 1410 4419 1427 4530
rect 1521 4419 1538 4530
rect 1410 4400 1538 4419
rect 1620 4530 1748 4546
rect 1620 4419 1637 4530
rect 1731 4419 1748 4530
rect 1620 4400 1748 4419
rect 1830 4530 1958 4546
rect 1830 4419 1847 4530
rect 1941 4419 1958 4530
rect 1830 4400 1958 4419
rect 2040 4530 2168 4546
rect 2040 4419 2057 4530
rect 2151 4419 2168 4530
rect 2040 4400 2168 4419
rect 2250 4530 2378 4546
rect 2250 4419 2267 4530
rect 2361 4419 2378 4530
rect 2250 4400 2378 4419
rect 2460 4530 2588 4546
rect 2460 4419 2477 4530
rect 2571 4419 2588 4530
rect 2460 4400 2588 4419
rect 2670 4530 2798 4546
rect 2670 4419 2687 4530
rect 2781 4419 2798 4530
rect 2670 4400 2798 4419
rect 2880 4530 3008 4546
rect 2880 4419 2897 4530
rect 2991 4419 3008 4530
rect 2880 4400 3008 4419
rect 3090 4530 3218 4546
rect 3090 4419 3107 4530
rect 3201 4419 3218 4530
rect 3090 4400 3218 4419
rect 3300 4530 3428 4546
rect 3300 4419 3317 4530
rect 3411 4419 3428 4530
rect 3300 4400 3428 4419
rect 3510 4530 3638 4546
rect 3510 4419 3527 4530
rect 3621 4419 3638 4530
rect 3510 4400 3638 4419
rect 3720 4530 3848 4546
rect 3720 4419 3737 4530
rect 3831 4419 3848 4530
rect 3720 4400 3848 4419
rect 0 2341 128 2357
rect 0 2230 17 2341
rect 111 2230 128 2341
rect 0 2211 128 2230
rect 210 2341 338 2357
rect 210 2230 227 2341
rect 321 2230 338 2341
rect 210 2211 338 2230
rect 420 2341 548 2357
rect 420 2230 437 2341
rect 531 2230 548 2341
rect 420 2211 548 2230
rect 630 2341 758 2357
rect 630 2230 647 2341
rect 741 2230 758 2341
rect 630 2211 758 2230
rect 840 2341 968 2357
rect 840 2230 857 2341
rect 951 2230 968 2341
rect 840 2211 968 2230
rect 1050 2341 1178 2357
rect 1050 2230 1067 2341
rect 1161 2230 1178 2341
rect 1050 2211 1178 2230
rect 1260 2341 1388 2357
rect 1260 2230 1277 2341
rect 1371 2230 1388 2341
rect 1260 2211 1388 2230
rect 1470 2341 1598 2357
rect 1470 2230 1487 2341
rect 1581 2230 1598 2341
rect 1470 2211 1598 2230
rect 1680 2341 1808 2357
rect 1680 2230 1697 2341
rect 1791 2230 1808 2341
rect 1680 2211 1808 2230
rect 1890 2341 2018 2357
rect 1890 2230 1907 2341
rect 2001 2230 2018 2341
rect 1890 2211 2018 2230
rect 2100 2341 2228 2357
rect 2100 2230 2117 2341
rect 2211 2230 2228 2341
rect 2100 2211 2228 2230
rect 2310 2341 2438 2357
rect 2310 2230 2327 2341
rect 2421 2230 2438 2341
rect 2310 2211 2438 2230
rect 2520 2341 2648 2357
rect 2520 2230 2537 2341
rect 2631 2230 2648 2341
rect 2520 2211 2648 2230
rect 2730 2341 2858 2357
rect 2730 2230 2747 2341
rect 2841 2230 2858 2341
rect 2730 2211 2858 2230
rect 2940 2341 3068 2357
rect 2940 2230 2957 2341
rect 3051 2230 3068 2341
rect 2940 2211 3068 2230
rect 3150 2341 3278 2357
rect 3150 2230 3167 2341
rect 3261 2230 3278 2341
rect 3150 2211 3278 2230
rect 3360 2341 3488 2357
rect 3360 2230 3377 2341
rect 3471 2230 3488 2341
rect 3360 2211 3488 2230
rect 3570 2341 3698 2357
rect 3570 2230 3587 2341
rect 3681 2230 3698 2341
rect 3570 2211 3698 2230
rect 3780 2341 3908 2357
rect 3780 2230 3797 2341
rect 3891 2230 3908 2341
rect 3780 2211 3908 2230
rect 3990 2341 4118 2357
rect 3990 2230 4007 2341
rect 4101 2230 4118 2341
rect 3990 2211 4118 2230
rect 0 1126 128 1142
rect 0 1015 17 1126
rect 111 1015 128 1126
rect 0 996 128 1015
rect 210 1126 338 1142
rect 210 1015 227 1126
rect 321 1015 338 1126
rect 210 996 338 1015
rect 420 1126 548 1142
rect 420 1015 437 1126
rect 531 1015 548 1126
rect 420 996 548 1015
rect 630 1126 758 1142
rect 630 1015 647 1126
rect 741 1015 758 1126
rect 630 996 758 1015
rect 840 1126 968 1142
rect 840 1015 857 1126
rect 951 1015 968 1126
rect 840 996 968 1015
rect 1050 1126 1178 1142
rect 1050 1015 1067 1126
rect 1161 1015 1178 1126
rect 1050 996 1178 1015
rect 1260 1126 1388 1142
rect 1260 1015 1277 1126
rect 1371 1015 1388 1126
rect 1260 996 1388 1015
rect 1470 1126 1598 1142
rect 1470 1015 1487 1126
rect 1581 1015 1598 1126
rect 1470 996 1598 1015
rect 1680 1126 1808 1142
rect 1680 1015 1697 1126
rect 1791 1015 1808 1126
rect 1680 996 1808 1015
rect 1890 1126 2018 1142
rect 1890 1015 1907 1126
rect 2001 1015 2018 1126
rect 1890 996 2018 1015
rect 2100 1126 2228 1142
rect 2100 1015 2117 1126
rect 2211 1015 2228 1126
rect 2100 996 2228 1015
rect 2310 1126 2438 1142
rect 2310 1015 2327 1126
rect 2421 1015 2438 1126
rect 2310 996 2438 1015
rect 2520 1126 2648 1142
rect 2520 1015 2537 1126
rect 2631 1015 2648 1126
rect 2520 996 2648 1015
rect 2730 1126 2858 1142
rect 2730 1015 2747 1126
rect 2841 1015 2858 1126
rect 2730 996 2858 1015
rect 2940 1126 3068 1142
rect 2940 1015 2957 1126
rect 3051 1015 3068 1126
rect 2940 996 3068 1015
rect 3150 1126 3278 1142
rect 3150 1015 3167 1126
rect 3261 1015 3278 1126
rect 3150 996 3278 1015
rect 3360 1126 3488 1142
rect 3360 1015 3377 1126
rect 3471 1015 3488 1126
rect 3360 996 3488 1015
rect 3570 1126 3698 1142
rect 3570 1015 3587 1126
rect 3681 1015 3698 1126
rect 3570 996 3698 1015
rect 3780 1126 3908 1142
rect 3780 1015 3797 1126
rect 3891 1015 3908 1126
rect 3780 996 3908 1015
rect 3990 1126 4118 1142
rect 3990 1015 4007 1126
rect 4101 1015 4118 1126
rect 3990 996 4118 1015
rect 0 -79 128 -63
rect 0 -190 17 -79
rect 111 -190 128 -79
rect 0 -209 128 -190
rect 210 -79 338 -63
rect 210 -190 227 -79
rect 321 -190 338 -79
rect 210 -209 338 -190
rect 420 -79 548 -63
rect 420 -190 437 -79
rect 531 -190 548 -79
rect 420 -209 548 -190
rect 630 -79 758 -63
rect 630 -190 647 -79
rect 741 -190 758 -79
rect 630 -209 758 -190
rect 840 -79 968 -63
rect 840 -190 857 -79
rect 951 -190 968 -79
rect 840 -209 968 -190
rect 1050 -79 1178 -63
rect 1050 -190 1067 -79
rect 1161 -190 1178 -79
rect 1050 -209 1178 -190
rect 1260 -79 1388 -63
rect 1260 -190 1277 -79
rect 1371 -190 1388 -79
rect 1260 -209 1388 -190
rect 1470 -79 1598 -63
rect 1470 -190 1487 -79
rect 1581 -190 1598 -79
rect 1470 -209 1598 -190
rect 1680 -79 1808 -63
rect 1680 -190 1697 -79
rect 1791 -190 1808 -79
rect 1680 -209 1808 -190
rect 1890 -79 2018 -63
rect 1890 -190 1907 -79
rect 2001 -190 2018 -79
rect 1890 -209 2018 -190
rect 2100 -79 2228 -63
rect 2100 -190 2117 -79
rect 2211 -190 2228 -79
rect 2100 -209 2228 -190
rect 2310 -79 2438 -63
rect 2310 -190 2327 -79
rect 2421 -190 2438 -79
rect 2310 -209 2438 -190
rect 2520 -79 2648 -63
rect 2520 -190 2537 -79
rect 2631 -190 2648 -79
rect 2520 -209 2648 -190
rect 2730 -79 2858 -63
rect 2730 -190 2747 -79
rect 2841 -190 2858 -79
rect 2730 -209 2858 -190
rect 2940 -79 3068 -63
rect 2940 -190 2957 -79
rect 3051 -190 3068 -79
rect 2940 -209 3068 -190
rect 3150 -79 3278 -63
rect 3150 -190 3167 -79
rect 3261 -190 3278 -79
rect 3150 -209 3278 -190
rect 3360 -79 3488 -63
rect 3360 -190 3377 -79
rect 3471 -190 3488 -79
rect 3360 -209 3488 -190
rect 3570 -79 3698 -63
rect 3570 -190 3587 -79
rect 3681 -190 3698 -79
rect 3570 -209 3698 -190
rect 3780 -79 3908 -63
rect 3780 -190 3797 -79
rect 3891 -190 3908 -79
rect 3780 -209 3908 -190
rect 3990 -79 4118 -63
rect 3990 -190 4007 -79
rect 4101 -190 4118 -79
rect 3990 -209 4118 -190
<< nsubdiff >>
rect -1758 7033 -1588 7046
rect -1758 6891 -1745 7033
rect -1604 6891 -1588 7033
rect -1758 6878 -1588 6891
rect -1528 7033 -1358 7046
rect -1528 6891 -1515 7033
rect -1374 6891 -1358 7033
rect -1528 6878 -1358 6891
rect -1298 7033 -1128 7046
rect -1298 6891 -1285 7033
rect -1144 6891 -1128 7033
rect -1298 6878 -1128 6891
rect -1068 7033 -898 7046
rect -1068 6891 -1055 7033
rect -914 6891 -898 7033
rect -1068 6878 -898 6891
rect -838 7033 -668 7046
rect -838 6891 -825 7033
rect -684 6891 -668 7033
rect -838 6878 -668 6891
rect -608 7033 -438 7046
rect -608 6891 -595 7033
rect -454 6891 -438 7033
rect -608 6878 -438 6891
rect -378 7033 -208 7046
rect -378 6891 -365 7033
rect -224 6891 -208 7033
rect -378 6878 -208 6891
rect -133 7033 37 7046
rect -133 6891 -120 7033
rect 21 6891 37 7033
rect -133 6878 37 6891
rect 420 6327 590 6340
rect 420 6185 433 6327
rect 574 6185 590 6327
rect 420 6172 590 6185
rect 650 6327 820 6340
rect 650 6185 663 6327
rect 804 6185 820 6327
rect 650 6172 820 6185
rect 880 6327 1050 6340
rect 880 6185 893 6327
rect 1034 6185 1050 6327
rect 880 6172 1050 6185
rect 1110 6327 1280 6340
rect 1110 6185 1123 6327
rect 1264 6185 1280 6327
rect 1110 6172 1280 6185
rect 1340 6327 1510 6340
rect 1340 6185 1353 6327
rect 1494 6185 1510 6327
rect 1340 6172 1510 6185
rect 1570 6327 1740 6340
rect 1570 6185 1583 6327
rect 1724 6185 1740 6327
rect 1570 6172 1740 6185
rect 1800 6327 1970 6340
rect 1800 6185 1813 6327
rect 1954 6185 1970 6327
rect 1800 6172 1970 6185
rect 2030 6327 2200 6340
rect 2030 6185 2043 6327
rect 2184 6185 2200 6327
rect 2030 6172 2200 6185
rect 2260 6327 2430 6340
rect 2260 6185 2273 6327
rect 2414 6185 2430 6327
rect 2260 6172 2430 6185
rect 2490 6327 2660 6340
rect 2490 6185 2503 6327
rect 2644 6185 2660 6327
rect 2490 6172 2660 6185
rect 2720 6327 2890 6340
rect 2720 6185 2733 6327
rect 2874 6185 2890 6327
rect 2720 6172 2890 6185
rect 2950 6327 3120 6340
rect 2950 6185 2963 6327
rect 3104 6185 3120 6327
rect 2950 6172 3120 6185
rect 3180 6327 3350 6340
rect 3180 6185 3193 6327
rect 3334 6185 3350 6327
rect 3180 6172 3350 6185
rect 3410 6327 3580 6340
rect 3410 6185 3423 6327
rect 3564 6185 3580 6327
rect 3410 6172 3580 6185
rect 3640 6327 3810 6340
rect 3640 6185 3653 6327
rect 3794 6185 3810 6327
rect 3640 6172 3810 6185
rect -1758 5843 -1588 5856
rect -1758 5701 -1745 5843
rect -1604 5701 -1588 5843
rect -1758 5688 -1588 5701
rect -1528 5843 -1358 5856
rect -1528 5701 -1515 5843
rect -1374 5701 -1358 5843
rect -1528 5688 -1358 5701
rect -1298 5843 -1128 5856
rect -1298 5701 -1285 5843
rect -1144 5701 -1128 5843
rect -1298 5688 -1128 5701
rect -1068 5843 -898 5856
rect -1068 5701 -1055 5843
rect -914 5701 -898 5843
rect -1068 5688 -898 5701
rect -838 5843 -668 5856
rect -838 5701 -825 5843
rect -684 5701 -668 5843
rect -838 5688 -668 5701
rect -608 5843 -438 5856
rect -608 5701 -595 5843
rect -454 5701 -438 5843
rect -608 5688 -438 5701
rect -378 5843 -208 5856
rect -378 5701 -365 5843
rect -224 5701 -208 5843
rect -378 5688 -208 5701
rect -133 5843 37 5856
rect -133 5701 -120 5843
rect 21 5701 37 5843
rect -133 5688 37 5701
rect -35 3877 135 3890
rect -35 3735 -22 3877
rect 119 3735 135 3877
rect -35 3722 135 3735
rect 195 3877 365 3890
rect 195 3735 208 3877
rect 349 3735 365 3877
rect 195 3722 365 3735
rect 425 3877 595 3890
rect 425 3735 438 3877
rect 579 3735 595 3877
rect 425 3722 595 3735
rect 655 3877 825 3890
rect 655 3735 668 3877
rect 809 3735 825 3877
rect 655 3722 825 3735
rect 885 3877 1055 3890
rect 885 3735 898 3877
rect 1039 3735 1055 3877
rect 885 3722 1055 3735
rect 1115 3877 1285 3890
rect 1115 3735 1128 3877
rect 1269 3735 1285 3877
rect 1115 3722 1285 3735
rect 1345 3877 1515 3890
rect 1345 3735 1358 3877
rect 1499 3735 1515 3877
rect 1345 3722 1515 3735
rect 1575 3877 1745 3890
rect 1575 3735 1588 3877
rect 1729 3735 1745 3877
rect 1575 3722 1745 3735
rect 1805 3877 1975 3890
rect 1805 3735 1818 3877
rect 1959 3735 1975 3877
rect 1805 3722 1975 3735
rect 2035 3877 2205 3890
rect 2035 3735 2048 3877
rect 2189 3735 2205 3877
rect 2035 3722 2205 3735
rect 2265 3877 2435 3890
rect 2265 3735 2278 3877
rect 2419 3735 2435 3877
rect 2265 3722 2435 3735
rect 2495 3877 2665 3890
rect 2495 3735 2508 3877
rect 2649 3735 2665 3877
rect 2495 3722 2665 3735
rect 2725 3877 2895 3890
rect 2725 3735 2738 3877
rect 2879 3735 2895 3877
rect 2725 3722 2895 3735
rect 2955 3877 3125 3890
rect 2955 3735 2968 3877
rect 3109 3735 3125 3877
rect 2955 3722 3125 3735
rect 3185 3877 3355 3890
rect 3185 3735 3198 3877
rect 3339 3735 3355 3877
rect 3185 3722 3355 3735
rect 3415 3877 3585 3890
rect 3415 3735 3428 3877
rect 3569 3735 3585 3877
rect 3415 3722 3585 3735
rect 3645 3877 3815 3890
rect 3645 3735 3658 3877
rect 3799 3735 3815 3877
rect 3645 3722 3815 3735
rect 3875 3877 4045 3890
rect 3875 3735 3888 3877
rect 4029 3735 4045 3877
rect 3875 3722 4045 3735
rect 4105 3877 4275 3890
rect 4105 3735 4118 3877
rect 4259 3735 4275 3877
rect 4105 3722 4275 3735
rect -35 2582 135 2595
rect -35 2440 -22 2582
rect 119 2440 135 2582
rect -35 2427 135 2440
rect 195 2582 365 2595
rect 195 2440 208 2582
rect 349 2440 365 2582
rect 195 2427 365 2440
rect 425 2582 595 2595
rect 425 2440 438 2582
rect 579 2440 595 2582
rect 425 2427 595 2440
rect 655 2582 825 2595
rect 655 2440 668 2582
rect 809 2440 825 2582
rect 655 2427 825 2440
rect 885 2582 1055 2595
rect 885 2440 898 2582
rect 1039 2440 1055 2582
rect 885 2427 1055 2440
rect 1115 2582 1285 2595
rect 1115 2440 1128 2582
rect 1269 2440 1285 2582
rect 1115 2427 1285 2440
rect 1345 2582 1515 2595
rect 1345 2440 1358 2582
rect 1499 2440 1515 2582
rect 1345 2427 1515 2440
rect 1575 2582 1745 2595
rect 1575 2440 1588 2582
rect 1729 2440 1745 2582
rect 1575 2427 1745 2440
rect 1805 2582 1975 2595
rect 1805 2440 1818 2582
rect 1959 2440 1975 2582
rect 1805 2427 1975 2440
rect 2035 2582 2205 2595
rect 2035 2440 2048 2582
rect 2189 2440 2205 2582
rect 2035 2427 2205 2440
rect 2265 2582 2435 2595
rect 2265 2440 2278 2582
rect 2419 2440 2435 2582
rect 2265 2427 2435 2440
rect 2495 2582 2665 2595
rect 2495 2440 2508 2582
rect 2649 2440 2665 2582
rect 2495 2427 2665 2440
rect 2725 2582 2895 2595
rect 2725 2440 2738 2582
rect 2879 2440 2895 2582
rect 2725 2427 2895 2440
rect 2955 2582 3125 2595
rect 2955 2440 2968 2582
rect 3109 2440 3125 2582
rect 2955 2427 3125 2440
rect 3185 2582 3355 2595
rect 3185 2440 3198 2582
rect 3339 2440 3355 2582
rect 3185 2427 3355 2440
rect 3415 2582 3585 2595
rect 3415 2440 3428 2582
rect 3569 2440 3585 2582
rect 3415 2427 3585 2440
rect 3645 2582 3815 2595
rect 3645 2440 3658 2582
rect 3799 2440 3815 2582
rect 3645 2427 3815 2440
rect 3875 2582 4045 2595
rect 3875 2440 3888 2582
rect 4029 2440 4045 2582
rect 3875 2427 4045 2440
rect 4105 2582 4275 2595
rect 4105 2440 4118 2582
rect 4259 2440 4275 2582
rect 4105 2427 4275 2440
<< psubdiffcont >>
rect -1761 5435 -1667 5546
rect -1494 5435 -1400 5546
rect -1284 5435 -1190 5546
rect -1074 5435 -980 5546
rect -864 5435 -770 5546
rect -654 5435 -560 5546
rect -444 5435 -350 5546
rect -234 5435 -140 5546
rect 377 5438 471 5549
rect 587 5438 681 5549
rect 797 5438 891 5549
rect 1007 5438 1101 5549
rect 1217 5438 1311 5549
rect 1427 5438 1521 5549
rect 1637 5438 1731 5549
rect 1847 5438 1941 5549
rect 2057 5438 2151 5549
rect 2267 5438 2361 5549
rect 2477 5438 2571 5549
rect 2687 5438 2781 5549
rect 2897 5438 2991 5549
rect 3107 5438 3201 5549
rect 3317 5438 3411 5549
rect 3527 5438 3621 5549
rect 3737 5438 3831 5549
rect -1620 4434 -1526 4545
rect -1410 4434 -1316 4545
rect -1200 4434 -1106 4545
rect -990 4434 -896 4545
rect -780 4434 -686 4545
rect -570 4434 -476 4545
rect -360 4434 -266 4545
rect -150 4434 -56 4545
rect 377 4419 471 4530
rect 587 4419 681 4530
rect 797 4419 891 4530
rect 1007 4419 1101 4530
rect 1217 4419 1311 4530
rect 1427 4419 1521 4530
rect 1637 4419 1731 4530
rect 1847 4419 1941 4530
rect 2057 4419 2151 4530
rect 2267 4419 2361 4530
rect 2477 4419 2571 4530
rect 2687 4419 2781 4530
rect 2897 4419 2991 4530
rect 3107 4419 3201 4530
rect 3317 4419 3411 4530
rect 3527 4419 3621 4530
rect 3737 4419 3831 4530
rect 17 2230 111 2341
rect 227 2230 321 2341
rect 437 2230 531 2341
rect 647 2230 741 2341
rect 857 2230 951 2341
rect 1067 2230 1161 2341
rect 1277 2230 1371 2341
rect 1487 2230 1581 2341
rect 1697 2230 1791 2341
rect 1907 2230 2001 2341
rect 2117 2230 2211 2341
rect 2327 2230 2421 2341
rect 2537 2230 2631 2341
rect 2747 2230 2841 2341
rect 2957 2230 3051 2341
rect 3167 2230 3261 2341
rect 3377 2230 3471 2341
rect 3587 2230 3681 2341
rect 3797 2230 3891 2341
rect 4007 2230 4101 2341
rect 17 1015 111 1126
rect 227 1015 321 1126
rect 437 1015 531 1126
rect 647 1015 741 1126
rect 857 1015 951 1126
rect 1067 1015 1161 1126
rect 1277 1015 1371 1126
rect 1487 1015 1581 1126
rect 1697 1015 1791 1126
rect 1907 1015 2001 1126
rect 2117 1015 2211 1126
rect 2327 1015 2421 1126
rect 2537 1015 2631 1126
rect 2747 1015 2841 1126
rect 2957 1015 3051 1126
rect 3167 1015 3261 1126
rect 3377 1015 3471 1126
rect 3587 1015 3681 1126
rect 3797 1015 3891 1126
rect 4007 1015 4101 1126
rect 17 -190 111 -79
rect 227 -190 321 -79
rect 437 -190 531 -79
rect 647 -190 741 -79
rect 857 -190 951 -79
rect 1067 -190 1161 -79
rect 1277 -190 1371 -79
rect 1487 -190 1581 -79
rect 1697 -190 1791 -79
rect 1907 -190 2001 -79
rect 2117 -190 2211 -79
rect 2327 -190 2421 -79
rect 2537 -190 2631 -79
rect 2747 -190 2841 -79
rect 2957 -190 3051 -79
rect 3167 -190 3261 -79
rect 3377 -190 3471 -79
rect 3587 -190 3681 -79
rect 3797 -190 3891 -79
rect 4007 -190 4101 -79
<< nsubdiffcont >>
rect -1745 6891 -1604 7033
rect -1515 6891 -1374 7033
rect -1285 6891 -1144 7033
rect -1055 6891 -914 7033
rect -825 6891 -684 7033
rect -595 6891 -454 7033
rect -365 6891 -224 7033
rect -120 6891 21 7033
rect 433 6185 574 6327
rect 663 6185 804 6327
rect 893 6185 1034 6327
rect 1123 6185 1264 6327
rect 1353 6185 1494 6327
rect 1583 6185 1724 6327
rect 1813 6185 1954 6327
rect 2043 6185 2184 6327
rect 2273 6185 2414 6327
rect 2503 6185 2644 6327
rect 2733 6185 2874 6327
rect 2963 6185 3104 6327
rect 3193 6185 3334 6327
rect 3423 6185 3564 6327
rect 3653 6185 3794 6327
rect -1745 5701 -1604 5843
rect -1515 5701 -1374 5843
rect -1285 5701 -1144 5843
rect -1055 5701 -914 5843
rect -825 5701 -684 5843
rect -595 5701 -454 5843
rect -365 5701 -224 5843
rect -120 5701 21 5843
rect -22 3735 119 3877
rect 208 3735 349 3877
rect 438 3735 579 3877
rect 668 3735 809 3877
rect 898 3735 1039 3877
rect 1128 3735 1269 3877
rect 1358 3735 1499 3877
rect 1588 3735 1729 3877
rect 1818 3735 1959 3877
rect 2048 3735 2189 3877
rect 2278 3735 2419 3877
rect 2508 3735 2649 3877
rect 2738 3735 2879 3877
rect 2968 3735 3109 3877
rect 3198 3735 3339 3877
rect 3428 3735 3569 3877
rect 3658 3735 3799 3877
rect 3888 3735 4029 3877
rect 4118 3735 4259 3877
rect -22 2440 119 2582
rect 208 2440 349 2582
rect 438 2440 579 2582
rect 668 2440 809 2582
rect 898 2440 1039 2582
rect 1128 2440 1269 2582
rect 1358 2440 1499 2582
rect 1588 2440 1729 2582
rect 1818 2440 1959 2582
rect 2048 2440 2189 2582
rect 2278 2440 2419 2582
rect 2508 2440 2649 2582
rect 2738 2440 2879 2582
rect 2968 2440 3109 2582
rect 3198 2440 3339 2582
rect 3428 2440 3569 2582
rect 3658 2440 3799 2582
rect 3888 2440 4029 2582
rect 4118 2440 4259 2582
<< polysilicon >>
rect -1635 6797 -107 6815
rect -1635 6762 -224 6797
rect -1635 6701 -1536 6762
rect -1635 6657 -1535 6701
rect -1023 6657 -923 6762
rect -819 6657 -719 6762
rect -240 6744 -224 6762
rect -172 6744 -107 6797
rect -240 6726 -107 6744
rect -207 6657 -107 6726
rect -1431 6310 -1331 6518
rect -1227 6310 -1127 6499
rect -615 6310 -515 6511
rect -411 6310 -311 6514
rect -1635 6270 -107 6310
rect -1635 6221 -1536 6270
rect -1635 6177 -1535 6221
rect -1023 6177 -923 6270
rect -819 6177 -719 6270
rect -1431 6007 -1331 6059
rect -1456 5987 -1331 6007
rect -1456 5931 -1428 5987
rect -1382 5958 -1331 5987
rect -1227 5958 -1127 6059
rect -615 5958 -515 6059
rect -411 5958 -311 6059
rect -1382 5931 -311 5958
rect -207 6020 -107 6270
rect -207 5959 -183 6020
rect -130 5959 -107 6020
rect -207 5940 -107 5959
rect 534 6083 3694 6097
rect 534 5993 581 6083
rect 671 6061 1109 6083
rect 671 5993 685 6061
rect 534 5979 685 5993
rect 1095 5993 1109 6061
rect 1199 6061 1397 6083
rect 1199 5993 1246 6061
rect 1095 5979 1246 5993
rect 534 5935 634 5979
rect 1146 5935 1246 5979
rect 1350 5993 1397 6061
rect 1487 6061 1925 6083
rect 1487 5993 1501 6061
rect 1350 5979 1501 5993
rect 1911 5993 1925 6061
rect 2015 6061 2213 6083
rect 2015 5993 2062 6061
rect 1911 5979 2062 5993
rect 1350 5935 1450 5979
rect 1962 5935 2062 5979
rect 2166 5993 2213 6061
rect 2303 6061 2741 6083
rect 2303 5993 2317 6061
rect 2166 5979 2317 5993
rect 2727 5993 2741 6061
rect 2831 6061 3029 6083
rect 2831 5993 2878 6061
rect 2727 5979 2878 5993
rect 2166 5935 2266 5979
rect 2778 5935 2878 5979
rect 2982 5993 3029 6061
rect 3119 6061 3559 6083
rect 3119 5993 3133 6061
rect 2982 5979 3133 5993
rect 3545 5993 3559 6061
rect 3649 5993 3694 6083
rect 3545 5979 3694 5993
rect 2982 5935 3082 5979
rect 3594 5935 3694 5979
rect -1456 5919 -311 5931
rect -1456 5918 -1374 5919
rect 738 5712 838 5815
rect 942 5762 1042 5815
rect 942 5712 956 5762
rect 738 5690 956 5712
rect 1028 5712 1042 5762
rect 1554 5762 1654 5815
rect 1554 5712 1568 5762
rect 1028 5690 1568 5712
rect 1640 5712 1654 5762
rect 1758 5762 1858 5815
rect 1758 5712 1772 5762
rect 1640 5690 1772 5712
rect 1844 5712 1858 5762
rect 2370 5762 2470 5815
rect 2370 5712 2384 5762
rect 1844 5690 2384 5712
rect 2456 5712 2470 5762
rect 2574 5762 2674 5815
rect 2574 5712 2588 5762
rect 2456 5690 2588 5712
rect 2660 5712 2674 5762
rect 3186 5762 3286 5815
rect 3186 5712 3200 5762
rect 2660 5690 3200 5712
rect 3272 5712 3286 5762
rect 3390 5762 3490 5815
rect 3390 5712 3404 5762
rect 3272 5690 3404 5712
rect 3476 5690 3490 5762
rect 738 5676 3490 5690
rect -1678 5360 508 5363
rect -1678 5346 3771 5360
rect -1678 5340 1098 5346
rect -1678 5310 490 5340
rect -1678 5249 -1579 5310
rect -1066 5249 -966 5310
rect -862 5249 -762 5310
rect -250 5249 -150 5310
rect 472 5290 490 5310
rect 540 5324 1098 5340
rect 540 5290 572 5324
rect 472 5260 572 5290
rect 1084 5274 1098 5324
rect 1170 5324 1914 5346
rect 1170 5274 1184 5324
rect 1084 5260 1184 5274
rect 1288 5272 1388 5324
rect 1900 5274 1914 5324
rect 1986 5324 3771 5346
rect 1986 5274 2000 5324
rect 1900 5260 2000 5274
rect 2243 5228 2343 5324
rect 2855 5228 2955 5324
rect 3059 5228 3159 5324
rect 3671 5228 3771 5324
rect 676 5043 776 5071
rect -1474 4992 -1374 5041
rect -1270 4992 -1170 5042
rect -658 4992 -558 5043
rect -454 4992 -354 5043
rect 676 5007 694 5043
rect 472 4993 694 5007
rect 744 5007 776 5043
rect 880 5068 980 5071
rect 880 5064 894 5068
rect 880 5043 980 5064
rect 880 5007 906 5043
rect 744 4993 906 5007
rect 956 5007 980 5043
rect 1492 5057 1592 5071
rect 1492 5007 1506 5057
rect 956 4993 1506 5007
rect 472 4992 1506 4993
rect -1678 4985 1506 4992
rect 1578 5007 1592 5057
rect 1696 5057 1796 5071
rect 1696 5007 1710 5057
rect 1578 4985 1710 5007
rect 1782 5007 1796 5057
rect 2447 5007 2547 5108
rect 2651 5007 2751 5108
rect 3263 5007 3363 5108
rect 3467 5007 3567 5108
rect 1782 4985 3771 5007
rect -1678 4971 3771 4985
rect -1678 4952 572 4971
rect -1678 4903 -1579 4952
rect -1678 4859 -1578 4903
rect -1066 4859 -966 4952
rect -862 4859 -762 4952
rect -250 4911 572 4952
rect -250 4859 -150 4911
rect 472 4875 572 4911
rect 1084 4875 1184 4971
rect 1288 4875 1388 4971
rect 1900 4875 2000 4971
rect 2243 4875 2343 4971
rect 2855 4875 2955 4971
rect 3059 4875 3159 4971
rect 3671 4875 3771 4971
rect 676 4721 776 4723
rect 676 4714 771 4721
rect 676 4709 776 4714
rect -1474 4638 -1374 4695
rect -1270 4638 -1170 4695
rect -658 4638 -558 4695
rect -454 4638 -354 4695
rect 676 4659 690 4709
rect -75 4638 690 4659
rect -1474 4637 690 4638
rect 762 4659 776 4709
rect 880 4659 980 4711
rect 1492 4659 1592 4711
rect 1696 4709 1796 4723
rect 1696 4659 1710 4709
rect 762 4637 1710 4659
rect 1782 4659 1796 4709
rect 2447 4659 2547 4755
rect 2651 4659 2751 4755
rect 3263 4659 3363 4755
rect 3467 4659 3567 4755
rect 1782 4637 3567 4659
rect -1474 4623 3567 4637
rect -1474 4599 784 4623
rect 112 4345 4088 4359
rect 112 4273 126 4345
rect 198 4323 4002 4345
rect 198 4273 212 4323
rect 112 4217 212 4273
rect 724 4217 824 4323
rect 928 4217 1028 4323
rect 1540 4217 1640 4323
rect 1744 4217 1844 4323
rect 2356 4217 2456 4323
rect 2560 4217 2660 4323
rect 3172 4217 3272 4323
rect 3376 4217 3476 4323
rect 3988 4273 4002 4323
rect 4074 4273 4088 4345
rect 3988 4217 4088 4273
rect 316 4014 416 4117
rect 520 4014 620 4117
rect 1132 4064 1232 4117
rect 1132 4014 1146 4064
rect 316 3992 1146 4014
rect 1218 4014 1232 4064
rect 1336 4014 1436 4117
rect 1948 4014 2048 4117
rect 2152 4014 2252 4117
rect 2764 4064 2864 4117
rect 2764 4014 2778 4064
rect 1218 3992 2778 4014
rect 2850 4014 2864 4064
rect 2968 4014 3068 4117
rect 3580 4014 3680 4117
rect 3784 4014 3884 4117
rect 2850 3992 3884 4014
rect 316 3978 3884 3992
rect 112 3649 4088 3663
rect 112 3579 180 3649
rect 250 3627 693 3649
rect 250 3579 264 3627
rect 112 3565 264 3579
rect 679 3579 693 3627
rect 763 3627 997 3649
rect 763 3579 824 3627
rect 679 3565 824 3579
rect 112 3521 212 3565
rect 724 3521 824 3565
rect 928 3579 997 3627
rect 1067 3627 1504 3649
rect 1067 3579 1081 3627
rect 928 3565 1081 3579
rect 1490 3579 1504 3627
rect 1574 3627 1813 3649
rect 1574 3579 1640 3627
rect 1490 3565 1640 3579
rect 928 3521 1028 3565
rect 1540 3521 1640 3565
rect 1744 3579 1813 3627
rect 1883 3627 2320 3649
rect 1883 3579 1897 3627
rect 1744 3565 1897 3579
rect 2306 3579 2320 3627
rect 2390 3627 2628 3649
rect 2390 3579 2456 3627
rect 2306 3565 2456 3579
rect 1744 3521 1844 3565
rect 2356 3521 2456 3565
rect 2560 3579 2628 3627
rect 2698 3627 3134 3649
rect 2698 3579 2712 3627
rect 2560 3565 2712 3579
rect 3120 3579 3134 3627
rect 3204 3627 3443 3649
rect 3204 3579 3272 3627
rect 3120 3565 3272 3579
rect 2560 3521 2660 3565
rect 3172 3521 3272 3565
rect 3376 3579 3443 3627
rect 3513 3627 3947 3649
rect 3513 3579 3527 3627
rect 3376 3565 3527 3579
rect 3933 3579 3947 3627
rect 4017 3579 4088 3649
rect 3933 3565 4088 3579
rect 3376 3521 3476 3565
rect 3988 3521 4088 3565
rect 316 3210 416 3321
rect 520 3210 620 3321
rect 316 3196 620 3210
rect 316 3173 412 3196
rect 112 3116 412 3173
rect 492 3173 620 3196
rect 1132 3215 1232 3321
rect 1336 3215 1436 3321
rect 1132 3201 1436 3215
rect 1132 3173 1241 3201
rect 492 3159 1241 3173
rect 492 3116 827 3159
rect 112 3102 827 3116
rect 112 2996 212 3102
rect 724 3074 827 3102
rect 915 3116 1241 3159
rect 1329 3173 1436 3201
rect 1948 3213 2048 3321
rect 2152 3213 2252 3321
rect 1948 3199 2252 3213
rect 1948 3173 2055 3199
rect 1329 3159 2055 3173
rect 1329 3116 1653 3159
rect 915 3102 1653 3116
rect 915 3074 1028 3102
rect 724 3060 1028 3074
rect 724 2996 824 3060
rect 928 2996 1028 3060
rect 1540 3070 1653 3102
rect 1745 3116 2055 3159
rect 2141 3173 2252 3199
rect 2764 3217 2864 3321
rect 2968 3217 3068 3321
rect 2764 3203 3068 3217
rect 2764 3173 2869 3203
rect 2141 3159 2869 3173
rect 2141 3116 2453 3159
rect 1745 3102 2453 3116
rect 1745 3070 1844 3102
rect 1540 3056 1844 3070
rect 1540 2996 1640 3056
rect 1744 2996 1844 3056
rect 2356 3075 2453 3102
rect 2537 3116 2869 3159
rect 2959 3173 3068 3203
rect 3580 3215 3680 3321
rect 3784 3215 3884 3321
rect 3580 3201 3884 3215
rect 3580 3173 3698 3201
rect 2959 3159 3698 3173
rect 2959 3116 3283 3159
rect 2537 3102 3283 3116
rect 2537 3075 2660 3102
rect 2356 3061 2660 3075
rect 2356 2996 2456 3061
rect 2560 2996 2660 3061
rect 3172 3073 3283 3102
rect 3369 3116 3698 3159
rect 3786 3173 3884 3201
rect 3786 3116 4088 3173
rect 3369 3102 4088 3116
rect 3369 3073 3476 3102
rect 3172 3059 3476 3073
rect 3172 2996 3272 3059
rect 3376 2996 3476 3059
rect 3988 2996 4088 3102
rect 316 2752 416 2796
rect 264 2738 416 2752
rect 264 2671 278 2738
rect 345 2693 416 2738
rect 520 2752 620 2796
rect 1132 2752 1232 2796
rect 520 2738 673 2752
rect 520 2693 592 2738
rect 345 2671 592 2693
rect 659 2693 673 2738
rect 1079 2738 1232 2752
rect 1079 2693 1093 2738
rect 659 2671 1093 2693
rect 1160 2693 1232 2738
rect 1336 2752 1436 2796
rect 1948 2752 2048 2796
rect 1336 2738 1486 2752
rect 1336 2693 1405 2738
rect 1160 2671 1405 2693
rect 1472 2693 1486 2738
rect 1900 2738 2048 2752
rect 1900 2693 1914 2738
rect 1472 2671 1914 2693
rect 1981 2693 2048 2738
rect 2152 2752 2252 2796
rect 2764 2752 2864 2796
rect 2152 2738 2305 2752
rect 2152 2693 2224 2738
rect 1981 2671 2224 2693
rect 2291 2693 2305 2738
rect 2714 2738 2864 2752
rect 2714 2693 2728 2738
rect 2291 2671 2728 2693
rect 2795 2693 2864 2738
rect 2968 2752 3068 2796
rect 2968 2738 3121 2752
rect 3580 2748 3680 2796
rect 2968 2693 3040 2738
rect 2795 2671 3040 2693
rect 3107 2693 3121 2738
rect 3527 2734 3680 2748
rect 3527 2693 3541 2734
rect 3107 2671 3541 2693
rect 3604 2693 3680 2734
rect 3784 2752 3884 2796
rect 3784 2738 3936 2752
rect 3784 2693 3855 2738
rect 3604 2671 3855 2693
rect 3922 2671 3936 2738
rect 264 2657 3936 2671
rect 112 2130 4088 2144
rect 112 2108 1758 2130
rect 112 2046 212 2108
rect 724 2046 824 2108
rect 928 2046 1028 2108
rect 1540 2046 1640 2108
rect 1744 2058 1758 2108
rect 1830 2128 4088 2130
rect 1830 2108 2370 2128
rect 1830 2058 1844 2108
rect 1744 2044 1844 2058
rect 2356 2056 2370 2108
rect 2442 2108 4088 2128
rect 2442 2056 2456 2108
rect 2356 2042 2456 2056
rect 2560 2046 2660 2108
rect 3172 2046 3272 2108
rect 3376 2046 3476 2108
rect 3988 2046 4088 2108
rect 316 1693 416 1758
rect 520 1693 620 1758
rect 1132 1693 1232 1758
rect 1336 1693 1436 1758
rect 1948 1693 2048 1758
rect 2152 1693 2252 1758
rect 2764 1693 2864 1758
rect 2968 1693 3068 1758
rect 3580 1693 3680 1758
rect 3784 1693 3884 1758
rect -151 1657 4354 1693
rect -151 1579 -115 1657
rect -181 1564 -92 1579
rect -181 1513 -165 1564
rect -111 1513 -92 1564
rect 112 1551 212 1657
rect 724 1551 824 1657
rect 928 1551 1028 1657
rect 1540 1551 1640 1657
rect 1744 1551 1844 1657
rect 2356 1551 2456 1657
rect 2560 1551 2660 1657
rect 3172 1551 3272 1657
rect 3376 1551 3476 1657
rect 3988 1551 4088 1657
rect 4318 1598 4354 1657
rect 4296 1582 4385 1598
rect 4296 1528 4312 1582
rect 4368 1528 4385 1582
rect 4296 1515 4385 1528
rect -181 1498 -92 1513
rect 316 1248 416 1307
rect 520 1248 620 1307
rect 1132 1248 1232 1307
rect 1336 1298 1436 1312
rect 1336 1248 1350 1298
rect 316 1226 1350 1248
rect 1422 1248 1436 1298
rect 1948 1248 2048 1307
rect 2152 1298 2252 1312
rect 2152 1248 2166 1298
rect 1422 1226 2166 1248
rect 2238 1248 2252 1298
rect 2764 1298 2864 1312
rect 2764 1248 2778 1298
rect 2238 1226 2778 1248
rect 2850 1248 2864 1298
rect 2968 1248 3068 1307
rect 3580 1248 3680 1307
rect 3784 1248 3884 1307
rect 2850 1226 3884 1248
rect 316 1212 3884 1226
rect 112 915 4088 929
rect 112 843 126 915
rect 198 914 942 915
rect 198 893 738 914
rect 198 843 212 893
rect 112 829 212 843
rect 724 842 738 893
rect 810 893 942 914
rect 810 842 824 893
rect 724 828 824 842
rect 928 843 942 893
rect 1014 893 1554 915
rect 1014 843 1028 893
rect 928 829 1028 843
rect 1540 843 1554 893
rect 1626 893 1758 915
rect 1626 843 1640 893
rect 1540 829 1640 843
rect 1744 843 1758 893
rect 1830 893 2370 915
rect 1830 843 1844 893
rect 1744 829 1844 843
rect 2356 843 2370 893
rect 2442 893 2574 915
rect 2442 843 2456 893
rect 2356 829 2456 843
rect 2560 843 2574 893
rect 2646 893 3186 915
rect 2646 843 2660 893
rect 2560 829 2660 843
rect 3172 843 3186 893
rect 3258 893 3390 915
rect 3258 843 3272 893
rect 3172 829 3272 843
rect 3376 843 3390 893
rect 3462 893 4002 915
rect 3462 843 3476 893
rect 3376 829 3476 843
rect 3988 843 4002 893
rect 4074 843 4088 915
rect 3988 829 4088 843
rect 316 531 416 545
rect 316 481 330 531
rect 112 459 330 481
rect 402 481 416 531
rect 520 531 620 545
rect 520 481 534 531
rect 402 459 534 481
rect 606 481 620 531
rect 1132 531 1232 545
rect 1132 481 1146 531
rect 606 467 1146 481
rect 606 459 738 467
rect 112 445 738 459
rect 112 339 212 445
rect 724 395 738 445
rect 810 445 942 467
rect 810 395 824 445
rect 724 339 824 395
rect 928 395 942 445
rect 1014 459 1146 467
rect 1218 481 1232 531
rect 1336 531 1436 545
rect 1336 481 1350 531
rect 1218 459 1350 481
rect 1422 481 1436 531
rect 1948 531 2048 545
rect 1948 481 1962 531
rect 1422 467 1962 481
rect 1422 459 1554 467
rect 1014 445 1554 459
rect 1014 395 1028 445
rect 928 339 1028 395
rect 1540 395 1554 445
rect 1626 445 1758 467
rect 1626 395 1640 445
rect 1540 339 1640 395
rect 1744 395 1758 445
rect 1830 459 1962 467
rect 2034 481 2048 531
rect 2152 531 2252 545
rect 2152 481 2166 531
rect 2034 459 2166 481
rect 2238 481 2252 531
rect 2764 531 2864 545
rect 2764 481 2778 531
rect 2238 467 2778 481
rect 2238 459 2370 467
rect 1830 445 2370 459
rect 1830 395 1844 445
rect 1744 339 1844 395
rect 2356 395 2370 445
rect 2442 445 2574 467
rect 2442 395 2456 445
rect 2356 339 2456 395
rect 2560 395 2574 445
rect 2646 459 2778 467
rect 2850 481 2864 531
rect 2968 531 3068 545
rect 2968 481 2982 531
rect 2850 459 2982 481
rect 3054 481 3068 531
rect 3580 531 3680 545
rect 3580 481 3594 531
rect 3054 467 3594 481
rect 3054 459 3186 467
rect 2646 445 3186 459
rect 2646 395 2660 445
rect 2560 339 2660 395
rect 3172 395 3186 445
rect 3258 445 3390 467
rect 3258 395 3272 445
rect 3172 339 3272 395
rect 3376 395 3390 445
rect 3462 459 3594 467
rect 3666 481 3680 531
rect 3784 531 3884 545
rect 3784 481 3798 531
rect 3666 459 3798 481
rect 3870 481 3884 531
rect 3870 459 4088 481
rect 3462 445 4088 459
rect 3462 395 3476 445
rect 3376 339 3476 395
rect 3988 339 4088 445
rect 316 86 416 100
rect 316 14 330 86
rect 402 36 416 86
rect 520 86 620 100
rect 520 36 534 86
rect 402 14 534 36
rect 606 36 620 86
rect 1132 86 1232 100
rect 1132 36 1146 86
rect 606 14 1146 36
rect 1218 36 1232 86
rect 1336 86 1436 100
rect 1336 36 1350 86
rect 1218 14 1350 36
rect 1422 36 1436 86
rect 1948 86 2048 100
rect 1948 36 1962 86
rect 1422 14 1962 36
rect 2034 36 2048 86
rect 2152 86 2252 100
rect 2152 36 2166 86
rect 2034 14 2166 36
rect 2238 36 2252 86
rect 2764 86 2864 100
rect 2764 36 2778 86
rect 2238 14 2778 36
rect 2850 36 2864 86
rect 2968 86 3068 100
rect 2968 36 2982 86
rect 2850 14 2982 36
rect 3054 36 3068 86
rect 3580 86 3680 100
rect 3580 36 3594 86
rect 3054 14 3594 36
rect 3666 36 3680 86
rect 3784 86 3884 100
rect 3784 36 3798 86
rect 3666 14 3798 36
rect 3870 14 3884 86
rect 316 0 3884 14
<< polycontact >>
rect -224 6744 -172 6797
rect -1428 5931 -1382 5987
rect -183 5959 -130 6020
rect 581 5993 671 6083
rect 1109 5993 1199 6083
rect 1397 5993 1487 6083
rect 1925 5993 2015 6083
rect 2213 5993 2303 6083
rect 2741 5993 2831 6083
rect 3029 5993 3119 6083
rect 3559 5993 3649 6083
rect 956 5690 1028 5762
rect 1568 5690 1640 5762
rect 1772 5690 1844 5762
rect 2384 5690 2456 5762
rect 2588 5690 2660 5762
rect 3200 5690 3272 5762
rect 3404 5690 3476 5762
rect 490 5290 540 5340
rect 1098 5274 1170 5346
rect 1914 5274 1986 5346
rect 694 4993 744 5043
rect 906 4993 956 5043
rect 1506 4985 1578 5057
rect 1710 4985 1782 5057
rect 690 4637 762 4709
rect 1710 4637 1782 4709
rect 126 4273 198 4345
rect 4002 4273 4074 4345
rect 1146 3992 1218 4064
rect 2778 3992 2850 4064
rect 180 3579 250 3649
rect 693 3579 763 3649
rect 997 3579 1067 3649
rect 1504 3579 1574 3649
rect 1813 3579 1883 3649
rect 2320 3579 2390 3649
rect 2628 3579 2698 3649
rect 3134 3579 3204 3649
rect 3443 3579 3513 3649
rect 3947 3579 4017 3649
rect 412 3116 492 3196
rect 827 3074 915 3159
rect 1241 3116 1329 3201
rect 1653 3070 1745 3159
rect 2055 3116 2141 3199
rect 2453 3075 2537 3159
rect 2869 3116 2959 3203
rect 3283 3073 3369 3159
rect 3698 3116 3786 3201
rect 278 2671 345 2738
rect 592 2671 659 2738
rect 1093 2671 1160 2738
rect 1405 2671 1472 2738
rect 1914 2671 1981 2738
rect 2224 2671 2291 2738
rect 2728 2671 2795 2738
rect 3040 2671 3107 2738
rect 3541 2671 3604 2734
rect 3855 2671 3922 2738
rect 1758 2058 1830 2130
rect 2370 2056 2442 2128
rect -165 1513 -111 1564
rect 4312 1528 4368 1582
rect 1350 1226 1422 1298
rect 2166 1226 2238 1298
rect 2778 1226 2850 1298
rect 126 843 198 915
rect 738 842 810 914
rect 942 843 1014 915
rect 1554 843 1626 915
rect 1758 843 1830 915
rect 2370 843 2442 915
rect 2574 843 2646 915
rect 3186 843 3258 915
rect 3390 843 3462 915
rect 4002 843 4074 915
rect 330 459 402 531
rect 534 459 606 531
rect 738 395 810 467
rect 942 395 1014 467
rect 1146 459 1218 531
rect 1350 459 1422 531
rect 1554 395 1626 467
rect 1758 395 1830 467
rect 1962 459 2034 531
rect 2166 459 2238 531
rect 2370 395 2442 467
rect 2574 395 2646 467
rect 2778 459 2850 531
rect 2982 459 3054 531
rect 3186 395 3258 467
rect 3390 395 3462 467
rect 3594 459 3666 531
rect 3798 459 3870 531
rect 330 14 402 86
rect 534 14 606 86
rect 1146 14 1218 86
rect 1350 14 1422 86
rect 1962 14 2034 86
rect 2166 14 2238 86
rect 2778 14 2850 86
rect 2982 14 3054 86
rect 3594 14 3666 86
rect 3798 14 3870 86
<< metal1 >>
rect -1809 7033 314 7070
rect -1809 6891 -1745 7033
rect -1604 6891 -1515 7033
rect -1374 6891 -1285 7033
rect -1144 6891 -1055 7033
rect -914 6891 -825 7033
rect -684 6891 -595 7033
rect -454 6891 -365 7033
rect -224 6891 -120 7033
rect 21 6891 314 7033
rect -1809 6878 314 6891
rect -1710 6655 -1664 6878
rect -894 6655 -848 6878
rect -238 6797 -164 6811
rect -238 6744 -224 6797
rect -172 6744 -164 6797
rect -238 6729 -164 6744
rect -78 6655 -32 6878
rect -1527 6626 -1450 6637
rect -1527 6574 -1513 6626
rect -1461 6574 -1450 6626
rect -1527 6560 -1450 6574
rect -1116 6625 -1039 6636
rect -1116 6573 -1102 6625
rect -1050 6573 -1039 6625
rect -1116 6559 -1039 6573
rect -708 6625 -631 6636
rect -708 6573 -694 6625
rect -642 6573 -631 6625
rect -708 6559 -631 6573
rect -302 6625 -225 6636
rect -302 6573 -288 6625
rect -236 6573 -225 6625
rect -302 6559 -225 6573
rect -1302 6413 -1256 6539
rect -487 6413 -441 6557
rect -1992 6316 -32 6413
rect -1710 6175 -1664 6316
rect -894 6175 -848 6316
rect -78 6175 -32 6316
rect 166 6364 314 6878
rect 166 6327 3868 6364
rect 166 6185 433 6327
rect 574 6185 663 6327
rect 804 6185 893 6327
rect 1034 6185 1123 6327
rect 1264 6185 1353 6327
rect 1494 6185 1583 6327
rect 1724 6185 1813 6327
rect 1954 6185 2043 6327
rect 2184 6185 2273 6327
rect 2414 6185 2503 6327
rect 2644 6185 2733 6327
rect 2874 6185 2963 6327
rect 3104 6185 3193 6327
rect 3334 6185 3423 6327
rect 3564 6185 3653 6327
rect 3794 6324 3868 6327
rect 3794 6226 4230 6324
rect 3794 6185 3868 6226
rect 166 6172 3868 6185
rect -1527 6158 -1450 6169
rect -1527 6106 -1513 6158
rect -1461 6106 -1450 6158
rect -1527 6092 -1450 6106
rect -1116 6144 -1039 6155
rect -1116 6092 -1102 6144
rect -1050 6092 -1039 6144
rect -1116 6078 -1039 6092
rect -711 6144 -634 6155
rect -711 6092 -697 6144
rect -645 6092 -634 6144
rect -711 6078 -634 6092
rect -302 6154 -225 6165
rect -302 6102 -288 6154
rect -236 6102 -225 6154
rect -302 6088 -225 6102
rect -1441 5988 -1368 6004
rect -1441 5931 -1428 5988
rect -1376 5931 -1368 5988
rect -1441 5914 -1368 5931
rect -1302 5856 -1256 6078
rect -486 5856 -440 6075
rect -193 6021 -116 6032
rect -193 6020 -177 6021
rect -193 5959 -183 6020
rect -125 5962 -116 6021
rect -130 5959 -116 5962
rect -193 5947 -116 5959
rect 166 5856 314 6172
rect 459 5933 505 6172
rect 572 6083 680 6092
rect 572 5993 581 6083
rect 671 6079 680 6083
rect 1100 6083 1208 6092
rect 1100 6079 1109 6083
rect 671 6033 1109 6079
rect 671 5993 709 6033
rect 572 5984 709 5993
rect -1809 5843 314 5856
rect -1809 5701 -1745 5843
rect -1604 5701 -1515 5843
rect -1374 5701 -1285 5843
rect -1144 5701 -1055 5843
rect -914 5701 -825 5843
rect -684 5701 -595 5843
rect -454 5701 -365 5843
rect -224 5701 -120 5843
rect 21 5708 314 5843
rect 663 5812 709 5984
rect 1071 5993 1109 6033
rect 1199 5993 1208 6083
rect 1071 5984 1208 5993
rect 1071 5933 1117 5984
rect 1275 5933 1321 6172
rect 1388 6083 1496 6092
rect 1388 5993 1397 6083
rect 1487 6073 1496 6083
rect 1916 6083 2024 6092
rect 1916 6073 1925 6083
rect 1487 6027 1925 6073
rect 1487 5993 1525 6027
rect 1388 5984 1525 5993
rect 1479 5933 1525 5984
rect 1887 5993 1925 6027
rect 2015 5993 2024 6083
rect 1887 5984 2024 5993
rect 1887 5933 1933 5984
rect 2091 5933 2137 6172
rect 2204 6083 2312 6092
rect 2204 5993 2213 6083
rect 2303 6070 2312 6083
rect 2732 6083 2840 6092
rect 2732 6070 2741 6083
rect 2303 6024 2741 6070
rect 2303 5993 2341 6024
rect 2204 5984 2341 5993
rect 2295 5933 2341 5984
rect 2703 5993 2741 6024
rect 2831 5993 2840 6083
rect 2703 5984 2840 5993
rect 2703 5933 2749 5984
rect 2907 5933 2953 6172
rect 3020 6083 3128 6092
rect 3020 5993 3029 6083
rect 3119 6076 3128 6083
rect 3550 6083 3658 6092
rect 3550 6076 3559 6083
rect 3119 6030 3559 6076
rect 3119 5993 3157 6030
rect 3020 5984 3157 5993
rect 3111 5933 3157 5984
rect 3519 5993 3559 6030
rect 3649 5993 3658 6083
rect 3519 5984 3658 5993
rect 3519 5933 3565 5984
rect 3723 5933 3769 6172
rect 636 5724 709 5812
rect 867 5771 913 5817
rect 1683 5771 1729 5817
rect 2499 5771 2545 5817
rect 3315 5771 3361 5817
rect 867 5762 3485 5771
rect 867 5716 956 5762
rect 21 5701 86 5708
rect -1809 5664 86 5701
rect 835 5690 956 5716
rect 1028 5725 1568 5762
rect 1028 5690 1037 5725
rect 835 5681 1037 5690
rect 1559 5690 1568 5725
rect 1640 5725 1772 5762
rect 1640 5690 1649 5725
rect 1559 5681 1649 5690
rect 1763 5690 1772 5725
rect 1844 5725 2384 5762
rect 1844 5690 1853 5725
rect 1763 5681 1853 5690
rect 2375 5690 2384 5725
rect 2456 5725 2588 5762
rect 2456 5690 2465 5725
rect 2375 5681 2465 5690
rect 2579 5690 2588 5725
rect 2660 5725 3200 5762
rect 2660 5690 2669 5725
rect 2579 5681 2669 5690
rect 3191 5690 3200 5725
rect 3272 5725 3404 5762
rect 3272 5690 3281 5725
rect 3191 5681 3281 5690
rect 3395 5690 3404 5725
rect 3476 5690 3485 5762
rect 3395 5681 3485 5690
rect 835 5632 913 5681
rect 360 5562 3883 5565
rect -1793 5549 3883 5562
rect -1793 5546 377 5549
rect -1793 5435 -1761 5546
rect -1667 5435 -1494 5546
rect -1400 5435 -1284 5546
rect -1190 5435 -1074 5546
rect -980 5435 -864 5546
rect -770 5435 -654 5546
rect -560 5435 -444 5546
rect -350 5435 -234 5546
rect -140 5438 377 5546
rect 471 5438 587 5549
rect 681 5438 797 5549
rect 891 5438 1007 5549
rect 1101 5438 1217 5549
rect 1311 5438 1427 5549
rect 1521 5438 1637 5549
rect 1731 5438 1847 5549
rect 1941 5438 2057 5549
rect 2151 5438 2267 5549
rect 2361 5438 2477 5549
rect 2571 5438 2687 5549
rect 2781 5438 2897 5549
rect 2991 5438 3107 5549
rect 3201 5438 3317 5549
rect 3411 5438 3527 5549
rect 3621 5438 3737 5549
rect 3831 5438 3883 5549
rect -140 5435 3883 5438
rect -1793 5419 3883 5435
rect -1793 5416 448 5419
rect -1345 5203 -1299 5416
rect -529 5203 -483 5416
rect 477 5340 567 5355
rect 477 5311 490 5340
rect 291 5290 490 5311
rect 540 5290 567 5340
rect 291 5265 567 5290
rect 291 5258 513 5265
rect 397 5226 443 5258
rect 805 5226 851 5419
rect 1089 5346 1179 5355
rect 1089 5274 1098 5346
rect 1170 5315 1179 5346
rect 1170 5274 1259 5315
rect 1089 5265 1259 5274
rect 1213 5226 1259 5265
rect 1621 5226 1667 5419
rect 1905 5346 1995 5355
rect 1905 5274 1914 5346
rect 1986 5311 1995 5346
rect 1986 5274 2075 5311
rect 1905 5265 2075 5274
rect 2029 5226 2075 5265
rect 2576 5226 2622 5419
rect 3392 5226 3438 5419
rect 2355 5200 2430 5210
rect -1565 5176 -1488 5187
rect -1565 5124 -1551 5176
rect -1499 5124 -1488 5176
rect -1565 5110 -1488 5124
rect -1158 5175 -1081 5186
rect -1158 5123 -1144 5175
rect -1092 5123 -1081 5175
rect -1158 5109 -1081 5123
rect -751 5175 -674 5186
rect -751 5123 -737 5175
rect -685 5123 -674 5175
rect -751 5109 -674 5123
rect -343 5175 -266 5186
rect -343 5123 -329 5175
rect -277 5123 -266 5175
rect 2355 5142 2365 5200
rect 2420 5142 2430 5200
rect -343 5109 -266 5123
rect -1753 5016 -1707 5087
rect -937 5016 -891 5087
rect -121 5016 -75 5087
rect 601 5067 647 5132
rect 601 5046 757 5067
rect 1009 5064 1055 5117
rect -1905 4948 -75 5016
rect 289 5043 757 5046
rect 289 4993 694 5043
rect 744 4993 757 5043
rect 289 4990 757 4993
rect 601 4976 757 4990
rect 890 5043 1055 5064
rect 890 4993 906 5043
rect 956 4993 1055 5043
rect -1345 4857 -1299 4948
rect -529 4857 -483 4948
rect 601 4873 647 4976
rect 890 4971 1055 4993
rect 1009 4873 1055 4971
rect 1417 5066 1463 5121
rect 1825 5066 1871 5116
rect 1417 5057 1587 5066
rect 1417 4985 1506 5057
rect 1578 4985 1587 5057
rect 1417 4976 1587 4985
rect 1701 5057 1871 5066
rect 1701 4985 1710 5057
rect 1782 4985 1871 5057
rect 2168 5043 2214 5135
rect 2355 5131 2430 5142
rect 2763 5196 2838 5206
rect 2763 5138 2773 5196
rect 2828 5138 2838 5196
rect 2763 5127 2838 5138
rect 3170 5197 3245 5207
rect 3170 5139 3180 5197
rect 3235 5139 3245 5197
rect 1701 4976 1871 4985
rect 1417 4873 1463 4976
rect 1825 4873 1871 4976
rect 2146 5024 2236 5043
rect 2146 4970 2164 5024
rect 2218 5020 2236 5024
rect 2984 5020 3030 5137
rect 3170 5128 3245 5139
rect 3580 5197 3655 5207
rect 3580 5139 3590 5197
rect 3645 5139 3655 5197
rect 3580 5128 3655 5139
rect 3800 5020 3846 5143
rect 2218 4974 3846 5020
rect 2218 4970 2236 4974
rect 2146 4953 2236 4970
rect 2576 4873 2622 4974
rect 3392 4873 3438 4974
rect 2356 4851 2431 4861
rect -1566 4830 -1489 4841
rect -1566 4778 -1552 4830
rect -1500 4778 -1489 4830
rect -1566 4764 -1489 4778
rect -1158 4830 -1081 4841
rect -1158 4778 -1144 4830
rect -1092 4778 -1081 4830
rect -1158 4764 -1081 4778
rect -751 4830 -674 4841
rect -751 4778 -737 4830
rect -685 4778 -674 4830
rect -751 4764 -674 4778
rect -343 4830 -266 4841
rect -343 4778 -329 4830
rect -277 4778 -266 4830
rect -343 4764 -266 4778
rect -1753 4561 -1707 4741
rect -937 4561 -891 4742
rect -121 4561 -75 4743
rect -1753 4545 -39 4561
rect 397 4546 443 4757
rect 805 4714 851 4764
rect 678 4709 851 4714
rect 678 4637 690 4709
rect 762 4668 851 4709
rect 762 4637 771 4668
rect 678 4626 771 4637
rect 687 4625 771 4626
rect 1213 4546 1259 4760
rect 1621 4722 1667 4757
rect 1621 4718 1743 4722
rect 1621 4709 1791 4718
rect 1621 4676 1710 4709
rect 1701 4637 1710 4676
rect 1782 4637 1791 4709
rect 1701 4628 1791 4637
rect 2029 4546 2075 4757
rect 2168 4546 2214 4826
rect 2356 4793 2366 4851
rect 2421 4793 2431 4851
rect 2356 4782 2431 4793
rect 2761 4849 2836 4859
rect 2761 4791 2771 4849
rect 2826 4791 2836 4849
rect 2761 4780 2836 4791
rect 2984 4546 3030 4861
rect 3171 4849 3246 4859
rect 3171 4791 3181 4849
rect 3236 4791 3246 4849
rect 3171 4780 3246 4791
rect 3580 4851 3655 4861
rect 3580 4793 3590 4851
rect 3645 4793 3655 4851
rect 3580 4782 3655 4793
rect 3800 4546 3846 4852
rect -1753 4434 -1620 4545
rect -1526 4434 -1410 4545
rect -1316 4434 -1200 4545
rect -1106 4434 -990 4545
rect -896 4434 -780 4545
rect -686 4434 -570 4545
rect -476 4434 -360 4545
rect -266 4434 -150 4545
rect -56 4434 -39 4545
rect -1753 4415 -39 4434
rect 360 4530 3883 4546
rect 360 4419 377 4530
rect 471 4419 587 4530
rect 681 4419 797 4530
rect 891 4419 1007 4530
rect 1101 4419 1217 4530
rect 1311 4419 1427 4530
rect 1521 4419 1637 4530
rect 1731 4419 1847 4530
rect 1941 4419 2057 4530
rect 2151 4419 2267 4530
rect 2361 4419 2477 4530
rect 2571 4419 2687 4530
rect 2781 4419 2897 4530
rect 2991 4419 3107 4530
rect 3201 4419 3317 4530
rect 3411 4419 3527 4530
rect 3621 4419 3737 4530
rect 3831 4419 3883 4530
rect 360 4400 3883 4419
rect 117 4345 207 4354
rect 117 4273 126 4345
rect 198 4273 207 4345
rect 3993 4345 4083 4354
rect 117 4264 207 4273
rect 431 4323 516 4333
rect 431 4322 3755 4323
rect 431 4262 446 4322
rect 506 4262 3755 4322
rect 3993 4273 4002 4345
rect 4074 4273 4083 4345
rect 3993 4264 4083 4273
rect 431 4261 3755 4262
rect 431 4249 516 4261
rect 228 4199 301 4209
rect 228 4141 237 4199
rect 291 4141 301 4199
rect 445 4163 491 4249
rect 636 4199 709 4209
rect 228 4130 301 4141
rect 636 4141 645 4199
rect 699 4141 709 4199
rect 636 4130 709 4141
rect 1043 4199 1116 4209
rect 1043 4141 1052 4199
rect 1106 4141 1116 4199
rect 1261 4173 1307 4261
rect 1453 4199 1526 4209
rect 1043 4130 1116 4141
rect 1453 4141 1462 4199
rect 1516 4141 1526 4199
rect 1453 4130 1526 4141
rect 1859 4199 1932 4209
rect 1859 4141 1868 4199
rect 1922 4141 1932 4199
rect 2077 4161 2123 4261
rect 2265 4199 2338 4209
rect 1859 4130 1932 4141
rect 2265 4141 2274 4199
rect 2328 4141 2338 4199
rect 2265 4130 2338 4141
rect 2675 4199 2748 4209
rect 2675 4141 2684 4199
rect 2738 4141 2748 4199
rect 2893 4169 2939 4261
rect 3080 4199 3153 4209
rect 2675 4130 2748 4141
rect 3080 4141 3089 4199
rect 3143 4141 3153 4199
rect 3080 4130 3153 4141
rect 3492 4199 3565 4209
rect 3492 4141 3501 4199
rect 3555 4141 3565 4199
rect 3709 4172 3755 4261
rect 3899 4199 3972 4209
rect 3492 4130 3565 4141
rect 3899 4141 3908 4199
rect 3962 4141 3972 4199
rect 3899 4130 3972 4141
rect 4132 4119 4230 6226
rect 37 3914 83 4119
rect 853 3914 899 4119
rect 1137 4064 1227 4073
rect 1137 3992 1146 4064
rect 1218 3992 1227 4064
rect 1137 3983 1227 3992
rect 1669 3914 1715 4119
rect 2485 3914 2531 4119
rect 2769 4064 2859 4073
rect 2769 3992 2778 4064
rect 2850 3992 2859 4064
rect 2769 3983 2859 3992
rect 3301 3914 3347 4119
rect 4117 3914 4230 4119
rect -62 3877 4299 3914
rect -62 3735 -22 3877
rect 119 3735 208 3877
rect 349 3735 438 3877
rect 579 3735 668 3877
rect 809 3735 898 3877
rect 1039 3735 1128 3877
rect 1269 3735 1358 3877
rect 1499 3735 1588 3877
rect 1729 3735 1818 3877
rect 1959 3735 2048 3877
rect 2189 3735 2278 3877
rect 2419 3735 2508 3877
rect 2649 3735 2738 3877
rect 2879 3735 2968 3877
rect 3109 3735 3198 3877
rect 3339 3735 3428 3877
rect 3569 3735 3658 3877
rect 3799 3735 3888 3877
rect 4029 3735 4118 3877
rect 4259 3735 4299 3877
rect -62 3722 4299 3735
rect 37 3519 83 3722
rect 171 3649 259 3658
rect 171 3579 180 3649
rect 250 3619 259 3649
rect 684 3649 772 3658
rect 684 3619 693 3649
rect 250 3579 287 3619
rect 171 3570 287 3579
rect 241 3519 287 3570
rect 649 3579 693 3619
rect 763 3579 772 3649
rect 649 3570 772 3579
rect 649 3519 695 3570
rect 853 3519 899 3722
rect 988 3649 1076 3658
rect 988 3579 997 3649
rect 1067 3619 1076 3649
rect 1495 3649 1583 3658
rect 1495 3619 1504 3649
rect 1067 3579 1103 3619
rect 988 3570 1103 3579
rect 1057 3519 1103 3570
rect 1465 3579 1504 3619
rect 1574 3579 1583 3649
rect 1465 3570 1583 3579
rect 1465 3519 1511 3570
rect 1669 3519 1715 3722
rect 1804 3649 1892 3658
rect 1804 3579 1813 3649
rect 1883 3619 1892 3649
rect 2311 3649 2399 3658
rect 2311 3619 2320 3649
rect 1883 3579 1919 3619
rect 1804 3570 1919 3579
rect 1873 3519 1919 3570
rect 2281 3579 2320 3619
rect 2390 3579 2399 3649
rect 2281 3570 2399 3579
rect 2281 3519 2327 3570
rect 2485 3519 2531 3722
rect 2619 3649 2707 3658
rect 2619 3579 2628 3649
rect 2698 3619 2707 3649
rect 3125 3649 3213 3658
rect 3125 3619 3134 3649
rect 2698 3579 2735 3619
rect 2619 3570 2735 3579
rect 2689 3519 2735 3570
rect 3097 3579 3134 3619
rect 3204 3579 3213 3649
rect 3097 3570 3213 3579
rect 3097 3519 3143 3570
rect 3301 3519 3347 3722
rect 3434 3649 3522 3658
rect 3434 3579 3443 3649
rect 3513 3619 3522 3649
rect 3938 3649 4026 3658
rect 3938 3619 3947 3649
rect 3513 3579 3551 3619
rect 3434 3570 3551 3579
rect 3505 3519 3551 3570
rect 3913 3579 3947 3619
rect 4017 3579 4026 3649
rect 3913 3570 4026 3579
rect 3913 3519 3959 3570
rect 4117 3519 4163 3722
rect 445 3205 491 3323
rect 1261 3210 1307 3323
rect 403 3196 501 3205
rect 403 3181 412 3196
rect 37 3135 412 3181
rect 37 2994 83 3135
rect 403 3116 412 3135
rect 492 3181 501 3196
rect 1232 3201 1338 3210
rect 2077 3208 2123 3323
rect 2893 3212 2939 3323
rect 1232 3181 1241 3201
rect 492 3159 1241 3181
rect 492 3135 827 3159
rect 492 3116 501 3135
rect 403 3107 501 3116
rect 818 3074 827 3135
rect 915 3135 1241 3159
rect 915 3074 924 3135
rect 1232 3116 1241 3135
rect 1329 3181 1338 3201
rect 2046 3199 2150 3208
rect 2046 3181 2055 3199
rect 1329 3159 2055 3181
rect 1329 3135 1653 3159
rect 1329 3116 1338 3135
rect 1232 3107 1338 3116
rect 818 3065 924 3074
rect 1644 3070 1653 3135
rect 1745 3135 2055 3159
rect 1745 3070 1754 3135
rect 2046 3116 2055 3135
rect 2141 3181 2150 3199
rect 2860 3203 2968 3212
rect 3709 3210 3755 3323
rect 2860 3181 2869 3203
rect 2141 3159 2869 3181
rect 2141 3135 2453 3159
rect 2141 3116 2150 3135
rect 2046 3107 2150 3116
rect 853 2994 899 3065
rect 1644 3061 1754 3070
rect 2444 3075 2453 3135
rect 2537 3135 2869 3159
rect 2537 3075 2546 3135
rect 2860 3116 2869 3135
rect 2959 3181 2968 3203
rect 3689 3201 3795 3210
rect 3689 3181 3698 3201
rect 2959 3159 3698 3181
rect 2959 3135 3283 3159
rect 2959 3116 2968 3135
rect 2860 3107 2968 3116
rect 2444 3066 2546 3075
rect 3274 3073 3283 3135
rect 3369 3135 3698 3159
rect 3369 3073 3378 3135
rect 3689 3116 3698 3135
rect 3786 3181 3795 3201
rect 3786 3135 4163 3181
rect 3786 3116 3795 3135
rect 3689 3107 3795 3116
rect 1669 2994 1715 3061
rect 2485 2994 2531 3066
rect 3274 3064 3378 3073
rect 3301 2994 3347 3064
rect 4117 2994 4163 3135
rect -182 2850 60 2915
rect 4131 2856 4486 2921
rect -182 1718 -117 2850
rect 241 2747 287 2798
rect 241 2738 354 2747
rect 241 2699 278 2738
rect 269 2671 278 2699
rect 345 2671 354 2738
rect 269 2662 354 2671
rect 445 2595 491 2798
rect 649 2747 695 2798
rect 583 2738 695 2747
rect 583 2671 592 2738
rect 659 2699 695 2738
rect 1057 2747 1103 2798
rect 1057 2738 1169 2747
rect 1057 2737 1093 2738
rect 1057 2699 1089 2737
rect 659 2671 668 2699
rect 583 2662 668 2671
rect 1080 2679 1089 2699
rect 1080 2671 1093 2679
rect 1160 2671 1169 2738
rect 1080 2668 1169 2671
rect 1084 2662 1169 2668
rect 1261 2595 1307 2798
rect 1465 2747 1511 2798
rect 1396 2738 1511 2747
rect 1396 2671 1405 2738
rect 1472 2699 1511 2738
rect 1873 2747 1919 2798
rect 1873 2738 1990 2747
rect 1873 2699 1914 2738
rect 1472 2671 1481 2699
rect 1396 2662 1481 2671
rect 1905 2671 1914 2699
rect 1981 2671 1990 2738
rect 1905 2662 1990 2671
rect 2077 2595 2123 2798
rect 2281 2747 2327 2798
rect 2215 2738 2327 2747
rect 2215 2671 2224 2738
rect 2291 2699 2327 2738
rect 2689 2748 2735 2798
rect 2689 2747 2801 2748
rect 2689 2738 2804 2747
rect 2689 2699 2728 2738
rect 2291 2671 2300 2699
rect 2215 2662 2300 2671
rect 2719 2671 2728 2699
rect 2795 2671 2804 2738
rect 2719 2662 2804 2671
rect 2893 2595 2939 2798
rect 3097 2747 3143 2798
rect 3031 2738 3143 2747
rect 3031 2671 3040 2738
rect 3107 2699 3143 2738
rect 3505 2743 3551 2798
rect 3505 2734 3613 2743
rect 3505 2699 3541 2734
rect 3107 2671 3116 2699
rect 3031 2662 3116 2671
rect 3532 2671 3541 2699
rect 3604 2671 3613 2734
rect 3532 2662 3613 2671
rect 3709 2595 3755 2798
rect 3913 2747 3959 2798
rect 3846 2738 3959 2747
rect 3846 2671 3855 2738
rect 3922 2699 3959 2738
rect 3922 2671 3931 2699
rect 3846 2662 3931 2671
rect -62 2582 4299 2595
rect -62 2440 -22 2582
rect 119 2440 208 2582
rect 349 2440 438 2582
rect 579 2440 668 2582
rect 809 2440 898 2582
rect 1039 2440 1128 2582
rect 1269 2440 1358 2582
rect 1499 2440 1588 2582
rect 1729 2440 1818 2582
rect 1959 2440 2048 2582
rect 2189 2440 2278 2582
rect 2419 2440 2508 2582
rect 2649 2440 2738 2582
rect 2879 2440 2968 2582
rect 3109 2440 3198 2582
rect 3339 2440 3428 2582
rect 3569 2440 3658 2582
rect 3799 2440 3888 2582
rect 4029 2440 4118 2582
rect 4259 2440 4299 2582
rect -62 2403 4299 2440
rect 0 2341 4200 2357
rect 0 2230 17 2341
rect 111 2230 227 2341
rect 321 2230 437 2341
rect 531 2230 647 2341
rect 741 2230 857 2341
rect 951 2230 1067 2341
rect 1161 2230 1277 2341
rect 1371 2230 1487 2341
rect 1581 2230 1697 2341
rect 1791 2230 1907 2341
rect 2001 2230 2117 2341
rect 2211 2230 2327 2341
rect 2421 2230 2537 2341
rect 2631 2230 2747 2341
rect 2841 2230 2957 2341
rect 3051 2230 3167 2341
rect 3261 2230 3377 2341
rect 3471 2230 3587 2341
rect 3681 2230 3797 2341
rect 3891 2230 4007 2341
rect 4101 2230 4200 2341
rect 0 2211 4200 2230
rect 445 2000 491 2211
rect 1261 2000 1307 2211
rect 1749 2130 1839 2139
rect 1749 2058 1758 2130
rect 1830 2058 1839 2130
rect 1749 2049 1839 2058
rect 2077 2000 2123 2211
rect 2361 2128 2451 2137
rect 2361 2056 2370 2128
rect 2442 2056 2451 2128
rect 2361 2047 2451 2056
rect 2893 2000 2939 2211
rect 3709 2000 3755 2211
rect 220 1926 293 1936
rect 220 1868 229 1926
rect 283 1868 293 1926
rect 220 1857 293 1868
rect 631 1934 704 1944
rect 631 1876 640 1934
rect 694 1876 704 1934
rect 631 1865 704 1876
rect 1038 1933 1111 1943
rect 1038 1875 1047 1933
rect 1101 1875 1111 1933
rect 1038 1864 1111 1875
rect 1448 1933 1521 1943
rect 1448 1875 1457 1933
rect 1511 1875 1521 1933
rect 1448 1864 1521 1875
rect 1854 1933 1927 1943
rect 1854 1875 1863 1933
rect 1917 1875 1927 1933
rect 1854 1864 1927 1875
rect 2264 1933 2337 1943
rect 2264 1875 2273 1933
rect 2327 1875 2337 1933
rect 2264 1864 2337 1875
rect 2671 1933 2744 1943
rect 2671 1875 2680 1933
rect 2734 1875 2744 1933
rect 2671 1864 2744 1875
rect 3076 1933 3149 1943
rect 3076 1875 3085 1933
rect 3139 1875 3149 1933
rect 3076 1864 3149 1875
rect 3486 1933 3559 1943
rect 3486 1875 3495 1933
rect 3549 1875 3559 1933
rect 3486 1864 3559 1875
rect 3897 1937 3970 1947
rect 3897 1879 3906 1937
rect 3960 1879 3970 1937
rect 3897 1868 3970 1879
rect 37 1718 83 1804
rect 853 1718 899 1809
rect 1669 1718 1715 1808
rect 2485 1718 2531 1811
rect 3301 1718 3347 1810
rect 4117 1718 4163 1807
rect 4421 1718 4486 2856
rect -182 1653 4486 1718
rect -181 1564 -92 1579
rect -181 1513 -165 1564
rect -111 1513 -92 1564
rect 445 1549 491 1653
rect 1261 1549 1307 1653
rect 2077 1549 2123 1653
rect 2893 1549 2939 1653
rect 3709 1549 3755 1653
rect 4296 1582 4385 1598
rect -181 530 -92 1513
rect 4296 1528 4312 1582
rect 4368 1528 4385 1582
rect 224 1482 297 1492
rect 224 1424 233 1482
rect 287 1424 297 1482
rect 224 1413 297 1424
rect 634 1481 707 1491
rect 634 1423 643 1481
rect 697 1423 707 1481
rect 634 1412 707 1423
rect 1043 1480 1116 1490
rect 1043 1422 1052 1480
rect 1106 1422 1116 1480
rect 1043 1411 1116 1422
rect 1452 1479 1525 1489
rect 1452 1421 1461 1479
rect 1515 1421 1525 1479
rect 1452 1410 1525 1421
rect 1861 1479 1934 1489
rect 1861 1421 1870 1479
rect 1924 1421 1934 1479
rect 1861 1410 1934 1421
rect 2267 1479 2340 1489
rect 2267 1421 2276 1479
rect 2330 1421 2340 1479
rect 2267 1410 2340 1421
rect 2674 1479 2747 1489
rect 2674 1421 2683 1479
rect 2737 1421 2747 1479
rect 2674 1410 2747 1421
rect 3082 1478 3155 1488
rect 3082 1420 3091 1478
rect 3145 1420 3155 1478
rect 3082 1409 3155 1420
rect 3490 1480 3563 1490
rect 3490 1422 3499 1480
rect 3553 1422 3563 1480
rect 3490 1411 3563 1422
rect 3898 1479 3971 1489
rect 3898 1421 3907 1479
rect 3961 1421 3971 1479
rect 3898 1410 3971 1421
rect 37 1142 83 1353
rect 853 1142 899 1353
rect 1341 1298 1431 1307
rect 1341 1226 1350 1298
rect 1422 1226 1431 1298
rect 1341 1217 1431 1226
rect 1669 1142 1715 1353
rect 2157 1298 2247 1307
rect 2157 1226 2166 1298
rect 2238 1226 2247 1298
rect 2157 1217 2247 1226
rect 2485 1142 2531 1353
rect 2769 1298 2859 1307
rect 2769 1226 2778 1298
rect 2850 1226 2859 1298
rect 2769 1217 2859 1226
rect 3301 1142 3347 1353
rect 4117 1142 4163 1353
rect 0 1126 4200 1142
rect 0 1015 17 1126
rect 111 1015 227 1126
rect 321 1015 437 1126
rect 531 1015 647 1126
rect 741 1015 857 1126
rect 951 1015 1067 1126
rect 1161 1015 1277 1126
rect 1371 1015 1487 1126
rect 1581 1015 1697 1126
rect 1791 1015 1907 1126
rect 2001 1015 2117 1126
rect 2211 1015 2327 1126
rect 2421 1015 2537 1126
rect 2631 1015 2747 1126
rect 2841 1015 2957 1126
rect 3051 1015 3167 1126
rect 3261 1015 3377 1126
rect 3471 1015 3587 1126
rect 3681 1015 3797 1126
rect 3891 1015 4007 1126
rect 4101 1015 4200 1126
rect 0 996 4200 1015
rect 117 915 207 924
rect 117 880 126 915
rect 37 843 126 880
rect 198 843 207 915
rect 37 834 207 843
rect 37 785 83 834
rect 445 785 491 996
rect 729 914 819 923
rect 729 842 738 914
rect 810 880 819 914
rect 933 915 1023 924
rect 933 880 942 915
rect 810 843 942 880
rect 1014 843 1023 915
rect 810 842 1023 843
rect 729 834 1023 842
rect 729 833 933 834
rect 853 785 899 833
rect 1261 785 1307 996
rect 1545 915 1635 924
rect 1545 843 1554 915
rect 1626 881 1635 915
rect 1749 915 1839 924
rect 1749 881 1758 915
rect 1626 843 1758 881
rect 1830 843 1839 915
rect 1545 834 1839 843
rect 1669 785 1715 834
rect 2077 785 2123 996
rect 2361 915 2451 924
rect 2361 843 2370 915
rect 2442 881 2451 915
rect 2565 915 2655 924
rect 2565 881 2574 915
rect 2442 843 2574 881
rect 2646 843 2655 915
rect 2361 834 2655 843
rect 2485 785 2531 834
rect 2893 785 2939 996
rect 3177 915 3267 924
rect 3177 843 3186 915
rect 3258 881 3267 915
rect 3381 915 3471 924
rect 3381 881 3390 915
rect 3258 843 3390 881
rect 3462 843 3471 915
rect 3177 834 3471 843
rect 3301 785 3347 834
rect 3709 785 3755 996
rect 3993 915 4083 924
rect 3993 843 4002 915
rect 4074 880 4083 915
rect 4074 843 4163 880
rect 3993 834 4163 843
rect 4117 785 4163 834
rect 241 548 287 589
rect 241 540 359 548
rect 649 547 695 589
rect 601 540 695 547
rect 241 531 411 540
rect 241 530 330 531
rect -181 459 330 530
rect 402 530 411 531
rect 525 531 695 540
rect 525 530 534 531
rect 402 459 534 530
rect 606 530 695 531
rect 1057 543 1103 594
rect 1465 554 1511 597
rect 1057 540 1169 543
rect 1405 540 1511 554
rect 1057 531 1227 540
rect 1057 530 1146 531
rect 606 467 1146 530
rect 606 459 738 467
rect -181 441 738 459
rect 241 430 358 441
rect 241 337 287 430
rect 649 395 738 441
rect 810 441 942 467
rect 810 395 819 441
rect 649 386 819 395
rect 933 395 942 441
rect 1014 459 1146 467
rect 1218 530 1227 531
rect 1341 531 1511 540
rect 1341 530 1350 531
rect 1218 459 1350 530
rect 1422 530 1511 531
rect 1873 543 1919 599
rect 2281 560 2327 596
rect 1873 540 1974 543
rect 2224 540 2327 560
rect 1873 531 2043 540
rect 1873 530 1962 531
rect 1422 467 1962 530
rect 1422 459 1554 467
rect 1014 441 1554 459
rect 1014 395 1103 441
rect 933 386 1103 395
rect 649 337 695 386
rect 987 379 1103 386
rect 1057 337 1103 379
rect 1465 395 1554 441
rect 1626 441 1758 467
rect 1626 395 1635 441
rect 1465 386 1635 395
rect 1749 395 1758 441
rect 1830 459 1962 467
rect 2034 530 2043 531
rect 2157 531 2327 540
rect 2157 530 2166 531
rect 2034 459 2166 530
rect 2238 530 2327 531
rect 2689 556 2735 598
rect 3097 564 3143 596
rect 2689 540 2785 556
rect 3031 540 3143 564
rect 2689 531 2859 540
rect 2689 530 2778 531
rect 2238 467 2778 530
rect 2238 459 2370 467
rect 1830 441 2370 459
rect 1830 395 1919 441
rect 1749 386 1919 395
rect 1465 383 1610 386
rect 1465 337 1511 383
rect 1781 377 1919 386
rect 1873 337 1919 377
rect 2281 395 2370 441
rect 2442 441 2574 467
rect 2442 395 2451 441
rect 2281 386 2451 395
rect 2565 395 2574 441
rect 2646 459 2778 467
rect 2850 530 2859 531
rect 2973 531 3143 540
rect 2973 530 2982 531
rect 2850 459 2982 530
rect 3054 530 3143 531
rect 3505 567 3551 600
rect 3505 540 3625 567
rect 3913 566 3959 600
rect 3858 540 3959 566
rect 3505 531 3675 540
rect 3505 530 3594 531
rect 3054 467 3594 530
rect 3054 459 3186 467
rect 2646 441 3186 459
rect 2646 395 2735 441
rect 2565 386 2735 395
rect 2281 367 2389 386
rect 2622 372 2735 386
rect 2281 337 2327 367
rect 2689 337 2735 372
rect 3097 395 3186 441
rect 3258 441 3390 467
rect 3258 395 3267 441
rect 3097 386 3267 395
rect 3381 395 3390 441
rect 3462 459 3594 467
rect 3666 530 3675 531
rect 3789 531 3959 540
rect 3789 530 3798 531
rect 3666 459 3798 530
rect 3870 530 3959 531
rect 4296 530 4385 1528
rect 3870 459 4385 530
rect 3462 441 4385 459
rect 3462 395 3551 441
rect 3381 386 3551 395
rect 3097 378 3229 386
rect 3097 337 3143 378
rect 3439 368 3551 386
rect 3505 337 3551 368
rect 3913 337 3959 441
rect -186 176 -87 196
rect -186 103 -171 176
rect -98 103 -87 176
rect -186 76 -87 103
rect 37 -63 83 141
rect 445 95 491 141
rect 321 86 615 95
rect 321 14 330 86
rect 402 48 534 86
rect 402 14 411 48
rect 321 5 411 14
rect 525 14 534 48
rect 606 14 615 86
rect 525 5 615 14
rect 853 -63 899 141
rect 1261 95 1307 141
rect 1137 86 1431 95
rect 1137 14 1146 86
rect 1218 48 1350 86
rect 1218 14 1227 48
rect 1137 5 1227 14
rect 1341 14 1350 48
rect 1422 14 1431 86
rect 1341 5 1431 14
rect 1669 -63 1715 141
rect 2077 95 2123 141
rect 1953 86 2247 95
rect 1953 14 1962 86
rect 2034 48 2166 86
rect 2034 14 2043 48
rect 1953 5 2043 14
rect 2157 14 2166 48
rect 2238 14 2247 86
rect 2157 5 2247 14
rect 2485 -63 2531 141
rect 2893 95 2939 141
rect 2769 86 3063 95
rect 2769 14 2778 86
rect 2850 48 2982 86
rect 2850 14 2859 48
rect 2769 5 2859 14
rect 2973 14 2982 48
rect 3054 14 3063 86
rect 2973 5 3063 14
rect 3301 -63 3347 141
rect 3709 95 3755 141
rect 3585 86 3879 95
rect 3585 14 3594 86
rect 3666 48 3798 86
rect 3666 14 3675 48
rect 3585 5 3675 14
rect 3789 14 3798 48
rect 3870 14 3879 86
rect 3789 5 3879 14
rect 4117 -63 4163 141
rect 0 -79 4200 -63
rect 0 -190 17 -79
rect 111 -190 227 -79
rect 321 -190 437 -79
rect 531 -190 647 -79
rect 741 -190 857 -79
rect 951 -190 1067 -79
rect 1161 -190 1277 -79
rect 1371 -190 1487 -79
rect 1581 -190 1697 -79
rect 1791 -190 1907 -79
rect 2001 -190 2117 -79
rect 2211 -190 2327 -79
rect 2421 -190 2537 -79
rect 2631 -190 2747 -79
rect 2841 -190 2957 -79
rect 3051 -190 3167 -79
rect 3261 -190 3377 -79
rect 3471 -190 3587 -79
rect 3681 -190 3797 -79
rect 3891 -190 4007 -79
rect 4101 -190 4200 -79
rect 0 -209 4200 -190
<< via1 >>
rect -224 6744 -172 6797
rect -1513 6574 -1461 6626
rect -1102 6573 -1050 6625
rect -694 6573 -642 6625
rect -288 6573 -236 6625
rect -1513 6106 -1461 6158
rect -1102 6092 -1050 6144
rect -697 6092 -645 6144
rect -288 6102 -236 6154
rect -1428 5987 -1376 5988
rect -1428 5931 -1382 5987
rect -1382 5931 -1376 5987
rect -177 6020 -125 6021
rect -177 5962 -130 6020
rect -130 5962 -125 6020
rect 596 6008 655 6068
rect 1776 5695 1832 5751
rect 2395 5695 2451 5751
rect 394 5476 449 5529
rect 3753 5455 3808 5513
rect 1103 5280 1160 5336
rect -1551 5124 -1499 5176
rect -1144 5123 -1092 5175
rect -737 5123 -685 5175
rect -329 5123 -277 5175
rect 2365 5142 2420 5200
rect 2773 5138 2828 5196
rect 3180 5139 3235 5197
rect 2164 4970 2218 5024
rect 3590 5139 3645 5197
rect -1552 4778 -1500 4830
rect -1144 4778 -1092 4830
rect -737 4778 -685 4830
rect -329 4778 -277 4830
rect 696 4643 751 4697
rect 2366 4793 2421 4851
rect 2771 4791 2826 4849
rect 3181 4791 3236 4849
rect 3590 4793 3645 4851
rect -128 4462 -73 4515
rect 394 4447 449 4500
rect 3753 4442 3808 4500
rect 129 4277 189 4337
rect 446 4262 506 4322
rect 4008 4280 4066 4338
rect 237 4141 291 4199
rect 645 4141 699 4199
rect 1052 4141 1106 4199
rect 1462 4141 1516 4199
rect 1868 4141 1922 4199
rect 2274 4141 2328 4199
rect 2684 4141 2738 4199
rect 3089 4141 3143 4199
rect 3501 4141 3555 4199
rect 3908 4141 3962 4199
rect 1152 4001 1209 4055
rect 2784 3999 2841 4055
rect 5 3772 59 3830
rect 4150 3772 4204 3830
rect 184 3584 243 3642
rect 1818 3585 1872 3643
rect 2330 3586 2384 3644
rect 3953 3585 4009 3642
rect 1250 3125 1318 3190
rect 2880 3127 2945 3190
rect 1089 2679 1093 2737
rect 1093 2679 1143 2737
rect 1916 2675 1970 2733
rect 2737 2680 2791 2738
rect 25 2502 79 2560
rect 4154 2481 4208 2539
rect 34 2268 89 2321
rect 4022 2256 4077 2309
rect 1764 2064 1819 2120
rect 2379 2065 2434 2121
rect 229 1868 283 1926
rect 640 1876 694 1934
rect 1047 1875 1101 1933
rect 1457 1875 1511 1933
rect 1863 1875 1917 1933
rect 2273 1875 2327 1933
rect 2680 1875 2734 1933
rect 3085 1875 3139 1933
rect 3495 1875 3549 1933
rect 3906 1879 3960 1937
rect 233 1424 287 1482
rect 643 1423 697 1481
rect 1052 1422 1106 1480
rect 1461 1421 1515 1479
rect 1870 1421 1924 1479
rect 2276 1421 2330 1479
rect 2683 1421 2737 1479
rect 3091 1420 3145 1478
rect 3499 1422 3553 1480
rect 3907 1421 3961 1479
rect 1357 1234 1414 1289
rect 2173 1235 2230 1290
rect 2782 1231 2842 1291
rect 34 1053 89 1106
rect 4022 1041 4077 1094
rect 136 855 190 909
rect 1561 851 1616 906
rect 2380 854 2432 906
rect -171 103 -98 176
rect 1154 21 1207 77
rect 1974 21 2029 79
rect 2785 21 2842 80
rect 34 -162 89 -109
rect 4025 -165 4080 -112
<< metal2 >>
rect -1705 6797 657 6815
rect -1705 6748 -224 6797
rect -1705 5978 -1638 6748
rect -235 6744 -224 6748
rect -172 6748 657 6797
rect -172 6744 -167 6748
rect -235 6732 -167 6744
rect -1527 6626 -1450 6637
rect -1527 6574 -1513 6626
rect -1461 6616 -1450 6626
rect -1116 6625 -1039 6636
rect -1116 6616 -1102 6625
rect -1461 6574 -1102 6616
rect -1527 6573 -1102 6574
rect -1050 6616 -1039 6625
rect -708 6625 -631 6636
rect -708 6616 -694 6625
rect -1050 6573 -694 6616
rect -642 6616 -631 6625
rect -302 6625 -225 6636
rect -302 6616 -288 6625
rect -642 6573 -288 6616
rect -236 6573 -225 6625
rect -1527 6560 -225 6573
rect -1516 6559 -225 6560
rect -1516 6205 -1459 6559
rect -1099 6205 -1042 6559
rect -694 6205 -637 6559
rect -287 6205 -230 6559
rect -1516 6169 -230 6205
rect -1527 6165 -230 6169
rect -1527 6158 -225 6165
rect -1527 6106 -1513 6158
rect -1461 6154 -225 6158
rect -1461 6148 -288 6154
rect -1461 6106 -1450 6148
rect -1527 6092 -1450 6106
rect -1116 6144 -1039 6148
rect -1116 6092 -1102 6144
rect -1050 6092 -1039 6144
rect -1116 6078 -1039 6092
rect -711 6144 -634 6148
rect -711 6092 -697 6144
rect -645 6092 -634 6144
rect -711 6078 -634 6092
rect -302 6102 -288 6148
rect -236 6102 -225 6154
rect -302 6088 -225 6102
rect 590 6085 657 6748
rect 579 6068 674 6085
rect -130 6033 -74 6034
rect -188 6021 -74 6033
rect -1441 5988 -1368 6004
rect -1441 5978 -1428 5988
rect -1705 5931 -1428 5978
rect -1376 5931 -1368 5988
rect -188 5962 -177 6021
rect -125 5962 -74 6021
rect 579 6008 596 6068
rect 655 6008 674 6068
rect 579 5992 674 6008
rect -188 5938 -74 5962
rect -1705 5914 -1368 5931
rect -1705 5911 -1394 5914
rect -130 5751 -74 5938
rect 1763 5751 1853 5771
rect 2375 5751 2465 5771
rect -130 5695 1776 5751
rect 1832 5695 2395 5751
rect 2451 5695 2465 5751
rect 1763 5681 1853 5695
rect 384 5529 461 5540
rect 384 5476 394 5529
rect 449 5476 461 5529
rect 384 5464 461 5476
rect -1565 5178 -1488 5187
rect -1158 5178 -1081 5186
rect -751 5178 -674 5186
rect -343 5178 -266 5186
rect -1565 5176 -266 5178
rect -1565 5124 -1551 5176
rect -1499 5175 -266 5176
rect -1499 5124 -1144 5175
rect -1565 5123 -1144 5124
rect -1092 5123 -737 5175
rect -685 5123 -329 5175
rect -277 5123 -266 5175
rect -1565 5120 -266 5123
rect -1565 5110 -1488 5120
rect -1555 4841 -1497 5110
rect -1158 5109 -1081 5120
rect -751 5109 -674 5120
rect -343 5109 -266 5120
rect -1146 4841 -1088 5109
rect -736 4841 -678 5109
rect -333 4841 -275 5109
rect -1566 4830 -1489 4841
rect -1566 4778 -1552 4830
rect -1500 4825 -1489 4830
rect -1158 4830 -1081 4841
rect -1158 4825 -1144 4830
rect -1500 4778 -1144 4825
rect -1092 4825 -1081 4830
rect -751 4830 -674 4841
rect -751 4825 -737 4830
rect -1092 4778 -737 4825
rect -685 4825 -674 4830
rect -343 4830 -266 4841
rect -343 4825 -329 4830
rect -685 4778 -329 4825
rect -277 4778 -266 4830
rect -1566 4767 -266 4778
rect -1566 4764 -1489 4767
rect -1158 4764 -1081 4767
rect -751 4764 -674 4767
rect -343 4764 -266 4767
rect -128 4526 -72 4561
rect -140 4521 -63 4526
rect -140 4515 -39 4521
rect -140 4499 -128 4515
rect -182 4462 -128 4499
rect -73 4499 -39 4515
rect 393 4511 449 5464
rect 1089 5336 1179 5355
rect 1089 5332 1103 5336
rect 690 5280 1103 5332
rect 1160 5280 1179 5336
rect 690 5276 1179 5280
rect 690 4723 746 5276
rect 1089 5265 1179 5276
rect 2163 5043 2219 5695
rect 2375 5681 2465 5695
rect 3743 5513 3818 5523
rect 3743 5455 3753 5513
rect 3808 5455 3818 5513
rect 3743 5444 3818 5455
rect 2355 5200 2430 5210
rect 2355 5142 2365 5200
rect 2420 5198 2430 5200
rect 2763 5198 2838 5206
rect 3170 5198 3245 5207
rect 3580 5198 3655 5207
rect 2420 5197 3655 5198
rect 2420 5196 3180 5197
rect 2420 5142 2773 5196
rect 2355 5131 2430 5142
rect 2763 5138 2773 5142
rect 2828 5142 3180 5196
rect 2828 5138 2838 5142
rect 2146 5024 2236 5043
rect 2146 4970 2164 5024
rect 2218 4970 2236 5024
rect 2146 4953 2236 4970
rect 2370 4861 2426 5131
rect 2763 5127 2838 5138
rect 3170 5139 3180 5142
rect 3235 5142 3590 5197
rect 3235 5139 3245 5142
rect 3170 5128 3245 5139
rect 3580 5139 3590 5142
rect 3645 5139 3655 5197
rect 3580 5128 3655 5139
rect 2356 4851 2431 4861
rect 2772 4859 2828 5127
rect 3178 4859 3234 5128
rect 3585 4861 3641 5128
rect 2356 4793 2366 4851
rect 2421 4793 2431 4851
rect 2356 4782 2431 4793
rect 2761 4849 2836 4859
rect 2761 4791 2771 4849
rect 2826 4791 2836 4849
rect 2761 4780 2836 4791
rect 3171 4849 3246 4859
rect 3171 4791 3181 4849
rect 3236 4791 3246 4849
rect 3171 4780 3246 4791
rect 3580 4851 3655 4861
rect 3580 4793 3590 4851
rect 3645 4793 3655 4851
rect 3580 4782 3655 4793
rect 678 4722 746 4723
rect 678 4697 771 4722
rect 678 4643 696 4697
rect 751 4643 771 4697
rect 678 4626 771 4643
rect 687 4625 771 4626
rect 384 4506 461 4511
rect 256 4500 461 4506
rect 256 4499 394 4500
rect -73 4462 394 4499
rect -182 4447 394 4462
rect 449 4447 461 4500
rect -182 4435 461 4447
rect -182 4434 446 4435
rect -182 4427 418 4434
rect -182 2329 -110 4427
rect 117 4348 206 4355
rect 92 4337 206 4348
rect 92 4277 129 4337
rect 189 4277 206 4337
rect 690 4333 746 4625
rect 3757 4510 3813 5444
rect 3743 4502 3818 4510
rect 3743 4500 4484 4502
rect 3743 4442 3753 4500
rect 3808 4442 4484 4500
rect 3743 4431 4484 4442
rect 3766 4430 4484 4431
rect 92 4264 206 4277
rect 431 4322 746 4333
rect 92 4021 148 4264
rect 431 4262 446 4322
rect 506 4277 746 4322
rect 3993 4346 4083 4354
rect 3993 4338 4115 4346
rect 3993 4280 4008 4338
rect 4066 4280 4115 4338
rect 506 4262 516 4277
rect 3993 4264 4115 4280
rect 431 4249 516 4262
rect 228 4199 301 4209
rect 228 4141 237 4199
rect 291 4193 301 4199
rect 636 4199 709 4209
rect 636 4193 645 4199
rect 291 4141 645 4193
rect 699 4193 709 4199
rect 1043 4199 1116 4209
rect 1043 4193 1052 4199
rect 699 4141 1052 4193
rect 1106 4193 1116 4199
rect 1453 4199 1526 4209
rect 1453 4193 1462 4199
rect 1106 4141 1462 4193
rect 1516 4193 1526 4199
rect 1859 4199 1932 4209
rect 1859 4193 1868 4199
rect 1516 4141 1868 4193
rect 1922 4193 1932 4199
rect 2265 4199 2338 4209
rect 2265 4193 2274 4199
rect 1922 4141 2274 4193
rect 2328 4193 2338 4199
rect 2675 4199 2748 4209
rect 2675 4193 2684 4199
rect 2328 4141 2684 4193
rect 2738 4193 2748 4199
rect 3080 4199 3153 4209
rect 3080 4193 3089 4199
rect 2738 4141 3089 4193
rect 3143 4193 3153 4199
rect 3492 4199 3565 4209
rect 3492 4193 3501 4199
rect 3143 4141 3501 4193
rect 3555 4193 3565 4199
rect 3899 4199 3972 4209
rect 3899 4193 3908 4199
rect 3555 4141 3908 4193
rect 3962 4141 3972 4199
rect 228 4137 3972 4141
rect 228 4130 301 4137
rect 636 4130 709 4137
rect 1043 4130 1116 4137
rect 1453 4130 1526 4137
rect 1859 4130 1932 4137
rect 2265 4130 2338 4137
rect 2675 4130 2748 4137
rect 3080 4130 3153 4137
rect 3492 4130 3565 4137
rect 3899 4130 3972 4137
rect 1137 4055 1227 4073
rect 92 3965 246 4021
rect 1137 4001 1152 4055
rect 1209 4033 1227 4055
rect 2769 4055 2859 4073
rect 1209 4001 1309 4033
rect 1137 3983 1309 4001
rect 2769 3999 2784 4055
rect 2841 4035 2859 4055
rect 2841 3999 2946 4035
rect 4059 4021 4115 4264
rect 2769 3983 2946 3999
rect 1153 3977 1309 3983
rect 2810 3979 2946 3983
rect -4 3832 69 3840
rect -4 3830 79 3832
rect -4 3772 5 3830
rect 59 3772 79 3830
rect -4 3761 79 3772
rect 23 2570 79 3761
rect 190 3658 246 3965
rect 171 3642 259 3658
rect 171 3584 184 3642
rect 243 3584 259 3642
rect 171 3570 259 3584
rect 1253 3210 1309 3977
rect 1809 3646 1882 3653
rect 2321 3646 2394 3654
rect 1809 3644 2394 3646
rect 1809 3643 2330 3644
rect 1809 3585 1818 3643
rect 1872 3590 2330 3643
rect 1872 3585 1882 3590
rect 1809 3574 1882 3585
rect 2310 3586 2330 3590
rect 2384 3586 2394 3644
rect 2310 3575 2394 3586
rect 1231 3190 1337 3210
rect 1231 3125 1250 3190
rect 1318 3125 1337 3190
rect 1231 3108 1337 3125
rect 1080 2737 1153 2747
rect 1080 2679 1089 2737
rect 1143 2723 1153 2737
rect 1814 2743 1870 3574
rect 1814 2733 1980 2743
rect 1814 2723 1916 2733
rect 1143 2679 1916 2723
rect 1080 2675 1916 2679
rect 1970 2723 1980 2733
rect 2310 2723 2366 3575
rect 2890 3208 2946 3979
rect 3956 3965 4115 4021
rect 3956 3658 4012 3965
rect 4141 3830 4214 3840
rect 4141 3772 4150 3830
rect 4204 3772 4214 3830
rect 4141 3761 4214 3772
rect 3938 3642 4026 3658
rect 3938 3585 3953 3642
rect 4009 3585 4026 3642
rect 3938 3570 4026 3585
rect 2863 3190 2964 3208
rect 2863 3127 2880 3190
rect 2945 3127 2964 3190
rect 2863 3111 2964 3127
rect 2728 2738 2801 2748
rect 2728 2723 2737 2738
rect 1970 2680 2737 2723
rect 2791 2680 2801 2738
rect 1970 2675 2801 2680
rect 1080 2669 2801 2675
rect 1080 2668 2772 2669
rect 1123 2667 2772 2668
rect 1907 2664 1980 2667
rect 16 2560 89 2570
rect 16 2502 25 2560
rect 79 2502 89 2560
rect 4151 2549 4207 3761
rect 16 2491 89 2502
rect 4145 2539 4218 2549
rect 4145 2481 4154 2539
rect 4208 2481 4218 2539
rect 4145 2470 4218 2481
rect 24 2329 101 2332
rect -182 2321 101 2329
rect -182 2268 34 2321
rect 89 2268 101 2321
rect -182 2257 101 2268
rect 24 2256 101 2257
rect 4012 2316 4089 2320
rect 4412 2316 4484 4430
rect 4012 2309 4484 2316
rect 4012 2256 4022 2309
rect 4077 2256 4484 2309
rect 33 1117 89 2256
rect 4012 2244 4484 2256
rect 1749 2126 1839 2139
rect 1749 2063 1762 2126
rect 1826 2063 1839 2126
rect 1749 2049 1839 2063
rect 2361 2123 2451 2137
rect 2361 2061 2375 2123
rect 2437 2061 2451 2123
rect 2361 2047 2451 2061
rect 220 1926 293 1936
rect 220 1868 229 1926
rect 283 1919 293 1926
rect 631 1934 704 1944
rect 631 1919 640 1934
rect 283 1876 640 1919
rect 694 1919 704 1934
rect 1038 1933 1111 1943
rect 1038 1919 1047 1933
rect 694 1876 1047 1919
rect 283 1875 1047 1876
rect 1101 1919 1111 1933
rect 1448 1933 1521 1943
rect 1448 1919 1457 1933
rect 1101 1875 1457 1919
rect 1511 1919 1521 1933
rect 1854 1933 1927 1943
rect 1854 1919 1863 1933
rect 1511 1875 1863 1919
rect 1917 1919 1927 1933
rect 2264 1933 2337 1943
rect 2264 1919 2273 1933
rect 1917 1875 2273 1919
rect 2327 1919 2337 1933
rect 2671 1933 2744 1943
rect 2671 1919 2680 1933
rect 2327 1875 2680 1919
rect 2734 1919 2744 1933
rect 3076 1933 3149 1943
rect 3076 1919 3085 1933
rect 2734 1875 3085 1919
rect 3139 1919 3149 1933
rect 3486 1933 3559 1943
rect 3486 1919 3495 1933
rect 3139 1875 3495 1919
rect 3549 1919 3559 1933
rect 3897 1937 3970 1947
rect 3897 1919 3906 1937
rect 3549 1879 3906 1919
rect 3960 1879 3970 1937
rect 3549 1875 3970 1879
rect 283 1868 3970 1875
rect 220 1863 3966 1868
rect 220 1857 293 1863
rect 229 1492 285 1857
rect 224 1482 297 1492
rect 638 1491 694 1863
rect 224 1424 233 1482
rect 287 1424 297 1482
rect 224 1413 297 1424
rect 634 1481 707 1491
rect 1047 1490 1103 1863
rect 634 1423 643 1481
rect 697 1423 707 1481
rect 634 1412 707 1423
rect 1043 1480 1116 1490
rect 1458 1489 1514 1863
rect 1865 1489 1921 1863
rect 2280 1489 2336 1863
rect 2677 1489 2733 1863
rect 1043 1422 1052 1480
rect 1106 1422 1116 1480
rect 1043 1411 1116 1422
rect 1452 1479 1525 1489
rect 1452 1421 1461 1479
rect 1515 1421 1525 1479
rect 1452 1410 1525 1421
rect 1861 1479 1934 1489
rect 1861 1421 1870 1479
rect 1924 1421 1934 1479
rect 1861 1410 1934 1421
rect 2267 1479 2340 1489
rect 2267 1421 2276 1479
rect 2330 1421 2340 1479
rect 2267 1410 2340 1421
rect 2674 1479 2747 1489
rect 3088 1488 3144 1863
rect 3504 1490 3560 1863
rect 2674 1421 2683 1479
rect 2737 1421 2747 1479
rect 2674 1410 2747 1421
rect 3082 1478 3155 1488
rect 3082 1420 3091 1478
rect 3145 1420 3155 1478
rect 3082 1409 3155 1420
rect 3490 1480 3563 1490
rect 3910 1489 3966 1863
rect 3490 1422 3499 1480
rect 3553 1422 3563 1480
rect 3490 1411 3563 1422
rect 3898 1479 3971 1489
rect 3898 1421 3907 1479
rect 3961 1421 3971 1479
rect 3898 1410 3971 1421
rect 1341 1293 1431 1307
rect 1341 1230 1353 1293
rect 1417 1290 1431 1293
rect 2157 1293 2246 1307
rect 2157 1290 2171 1293
rect 2232 1290 2246 1293
rect 2769 1292 2859 1307
rect 2769 1290 2782 1292
rect 1417 1234 2171 1290
rect 1417 1230 1431 1234
rect 1341 1217 1431 1230
rect 2157 1231 2171 1234
rect 2232 1234 2782 1290
rect 2232 1231 2263 1234
rect 2157 1217 2263 1231
rect 2769 1230 2782 1234
rect 2843 1230 2859 1292
rect 2769 1217 2859 1230
rect 24 1106 101 1117
rect 24 1053 34 1106
rect 89 1084 101 1106
rect 89 1053 808 1084
rect 24 1041 808 1053
rect 27 1028 808 1041
rect 127 909 200 919
rect 127 855 136 909
rect 190 855 200 909
rect -186 176 -87 196
rect 127 176 200 855
rect -186 103 -171 176
rect -98 103 200 176
rect -186 76 -87 103
rect 24 -109 101 -98
rect 24 -162 34 -109
rect 89 -112 101 -109
rect 752 -112 808 1028
rect 1367 904 1423 1217
rect 1548 906 1630 921
rect 1548 904 1561 906
rect 1367 851 1561 904
rect 1616 904 1630 906
rect 2207 904 2263 1217
rect 2366 906 2447 920
rect 2366 904 2380 906
rect 1616 854 2380 904
rect 2432 904 2447 906
rect 2799 904 2855 1217
rect 4029 1105 4085 2244
rect 4012 1094 4089 1105
rect 4012 1041 4022 1094
rect 4077 1041 4089 1094
rect 4012 1029 4089 1041
rect 2432 854 2855 904
rect 1616 851 2855 854
rect 1367 848 2855 851
rect 1548 837 1630 848
rect 2363 840 2447 848
rect 1139 77 1222 91
rect 1139 21 1154 77
rect 1207 75 1222 77
rect 1554 75 1610 837
rect 1961 79 2044 91
rect 1961 75 1974 79
rect 1207 21 1974 75
rect 2029 75 2044 79
rect 2363 75 2419 840
rect 2772 80 2855 92
rect 2772 75 2785 80
rect 2029 21 2785 75
rect 2842 21 2855 80
rect 1139 19 2855 21
rect 1139 8 1222 19
rect 1961 8 2044 19
rect 2772 8 2855 19
rect 4029 -101 4085 1029
rect 89 -162 808 -112
rect 24 -168 808 -162
rect 4015 -112 4092 -101
rect 4015 -165 4025 -112
rect 4080 -165 4092 -112
rect 24 -174 101 -168
rect 4015 -177 4092 -165
<< via2 >>
rect 1762 2120 1826 2126
rect 1762 2064 1764 2120
rect 1764 2064 1819 2120
rect 1819 2064 1826 2120
rect 1762 2063 1826 2064
rect 2375 2121 2437 2123
rect 2375 2065 2379 2121
rect 2379 2065 2434 2121
rect 2434 2065 2437 2121
rect 2375 2061 2437 2065
rect 1353 1289 1417 1293
rect 2171 1290 2232 1293
rect 2782 1291 2843 1292
rect 1353 1234 1357 1289
rect 1357 1234 1414 1289
rect 1414 1234 1417 1289
rect 2171 1235 2173 1290
rect 2173 1235 2230 1290
rect 2230 1235 2232 1290
rect 1353 1230 1417 1234
rect 2171 1231 2232 1235
rect 2782 1231 2842 1291
rect 2842 1231 2843 1291
rect 2782 1230 2843 1231
<< metal3 >>
rect 1749 2128 1839 2139
rect 2361 2128 2451 2137
rect 1749 2126 2451 2128
rect 1749 2063 1762 2126
rect 1826 2123 2451 2126
rect 1826 2067 2375 2123
rect 1826 2063 1839 2067
rect 1749 2049 1839 2063
rect 2361 2061 2375 2067
rect 2437 2061 2451 2123
rect 1341 1293 1431 1307
rect 1341 1230 1353 1293
rect 1417 1291 1431 1293
rect 1417 1290 1478 1291
rect 1769 1290 1830 2049
rect 2361 2047 2451 2061
rect 2157 1293 2247 1307
rect 2157 1290 2171 1293
rect 1417 1231 2171 1290
rect 2232 1290 2247 1293
rect 2375 1290 2436 2047
rect 2769 1292 2859 1307
rect 2769 1290 2782 1292
rect 2232 1231 2782 1290
rect 1417 1230 2782 1231
rect 2843 1230 2859 1292
rect 1341 1229 2859 1230
rect 1341 1217 1431 1229
rect 2157 1217 2247 1229
rect 2769 1217 2859 1229
use nmos_3p3_AJEA3B  nmos_3p3_AJEA3B_0
timestamp 1694665332
transform 1 0 1236 0 1 5168
box -876 -128 876 128
use nmos_3p3_AJEA3B  nmos_3p3_AJEA3B_1
timestamp 1694665332
transform 1 0 3007 0 1 4815
box -876 -128 876 128
use nmos_3p3_AJEA3B  nmos_3p3_AJEA3B_2
timestamp 1694665332
transform 1 0 -914 0 1 5145
box -876 -128 876 128
use nmos_3p3_AJEA3B  nmos_3p3_AJEA3B_3
timestamp 1694665332
transform 1 0 3007 0 1 5168
box -876 -128 876 128
use nmos_3p3_AJEA3B  nmos_3p3_AJEA3B_4
timestamp 1694665332
transform 1 0 1236 0 1 4815
box -876 -128 876 128
use nmos_3p3_AJEA3B  nmos_3p3_AJEA3B_5
timestamp 1694665332
transform 1 0 -914 0 1 4799
box -876 -128 876 128
use nmos_3p3_Z2JHD6  nmos_3p3_Z2JHD6_0
timestamp 1693483456
transform 1 0 2100 0 1 1902
box -2100 -168 2100 168
use nmos_3p3_Z2JHD6  nmos_3p3_Z2JHD6_1
timestamp 1693483456
transform 1 0 2100 0 1 239
box -2100 -168 2100 168
use nmos_3p3_Z2JHD6  nmos_3p3_Z2JHD6_2
timestamp 1693483456
transform 1 0 2100 0 1 687
box -2100 -168 2100 168
use nmos_3p3_Z2JHD6  nmos_3p3_Z2JHD6_3
timestamp 1693483456
transform 1 0 2100 0 1 1451
box -2100 -168 2100 168
use pfet_03v3_TTE2U8  pfet_03v3_TTE2U8_0
timestamp 1694679271
transform 1 0 -871 0 1 6117
box -938 -190 938 190
use pfet_03v3_TTE2U8  pfet_03v3_TTE2U8_1
timestamp 1694679271
transform 1 0 -871 0 1 6597
box -938 -190 938 190
use pmos_3p3_5QR9E7  pmos_3p3_5QR9E7_0
timestamp 1693564975
transform 1 0 2100 0 1 4157
box -2162 -170 2162 170
use pmos_3p3_DVJ9E7  pmos_3p3_DVJ9E7_0
timestamp 1693295468
transform 1 0 2114 0 1 5875
box -1754 -190 1754 190
use pmos_3p3_ZBCND7  pmos_3p3_ZBCND7_0
timestamp 1693543231
transform 1 0 2100 0 1 3421
box -2162 -230 2162 230
use pmos_3p3_ZBCND7  pmos_3p3_ZBCND7_1
timestamp 1693543231
transform 1 0 2100 0 1 2896
box -2162 -230 2162 230
<< labels >>
flabel nsubdiffcont 505 6259 505 6259 0 FreeSans 480 0 0 0 VDD
port 0 nsew
flabel metal1 513 5478 513 5478 0 FreeSans 480 0 0 0 VSS
port 3 nsew
flabel metal1 314 5279 314 5279 0 FreeSans 480 0 0 0 G_sink_up
port 4 nsew
flabel metal1 307 5018 307 5018 0 FreeSans 480 0 0 0 G_sink_dn
port 5 nsew
flabel via1 2395 5173 2395 5173 0 FreeSans 480 0 0 0 SD0_1
port 6 nsew
flabel polycontact 160 4312 160 4312 0 FreeSans 480 0 0 0 G1_2
port 7 nsew
flabel via1 263 4170 263 4170 0 FreeSans 480 0 0 0 SD1_1
port 9 nsew
flabel polycontact 1175 4023 1175 4023 0 FreeSans 480 0 0 0 G1_1
port 8 nsew
flabel polycontact 361 499 361 499 0 FreeSans 480 0 0 0 G2_1
port 10 nsew
flabel via1 252 1901 252 1901 0 FreeSans 480 0 0 0 SD2_1
port 11 nsew
flabel via1 -143 136 -143 141 0 FreeSans 480 0 0 0 ITAIL
port 12 nsew
flabel metal1 651 5747 651 5747 0 FreeSans 480 0 0 0 G_source_up
port 1 nsew
flabel metal1 851 5654 851 5654 0 FreeSans 480 0 0 0 G_source_dn
port 2 nsew
flabel metal1 -1875 4982 -1875 4982 0 FreeSans 1600 0 0 0 ITAIL_SINK
port 13 nsew
flabel metal1 -1963 6357 -1963 6357 0 FreeSans 1600 0 0 0 ITAIL_SRC
port 14 nsew
flabel via1 -260 6600 -260 6600 0 FreeSans 1600 0 0 0 A1
port 15 nsew
flabel via1 -303 5146 -303 5146 0 FreeSans 1600 0 0 0 A2
port 16 nsew
<< end >>
