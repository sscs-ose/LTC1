magic
tech gf180mcuC
magscale 1 10
timestamp 1692985371
<< nwell >>
rect 0 428 1060 569
rect 815 342 870 380
rect 397 -180 398 -151
rect 145 -341 916 -337
<< pwell >>
rect 205 -475 206 -466
rect 217 -480 269 -434
rect 609 -1130 620 -442
<< pmos >>
rect 662 -180 663 -151
<< psubdiff >>
rect 58 -1160 187 -1141
rect 58 -1210 73 -1160
rect 168 -1210 187 -1160
rect 58 -1223 187 -1210
rect 258 -1160 387 -1141
rect 258 -1210 273 -1160
rect 368 -1210 387 -1160
rect 258 -1223 387 -1210
rect 458 -1160 587 -1141
rect 458 -1210 473 -1160
rect 568 -1210 587 -1160
rect 458 -1223 587 -1210
rect 658 -1160 787 -1141
rect 658 -1210 673 -1160
rect 768 -1210 787 -1160
rect 658 -1223 787 -1210
<< nsubdiff >>
rect 58 529 176 545
rect 58 483 78 529
rect 147 483 176 529
rect 58 469 176 483
rect 258 529 376 545
rect 258 483 278 529
rect 347 483 376 529
rect 258 469 376 483
rect 478 529 596 545
rect 478 483 498 529
rect 567 483 596 529
rect 478 469 596 483
rect 698 529 816 545
rect 698 483 718 529
rect 787 483 816 529
rect 698 469 816 483
rect 898 529 1016 545
rect 898 483 918 529
rect 987 483 1016 529
rect 898 469 1016 483
<< psubdiffcont >>
rect 73 -1210 168 -1160
rect 273 -1210 368 -1160
rect 473 -1210 568 -1160
rect 673 -1210 768 -1160
<< nsubdiffcont >>
rect 78 483 147 529
rect 278 483 347 529
rect 498 483 567 529
rect 718 483 787 529
rect 918 483 987 529
<< polysilicon >>
rect 174 342 886 394
rect 113 89 174 97
rect 113 84 274 89
rect 113 37 126 84
rect 174 37 274 84
rect 113 21 274 37
rect 786 -25 886 4
rect 786 -28 807 -25
rect 174 -72 807 -28
rect 862 -72 886 -25
rect 174 -81 886 -72
rect 192 -431 498 -418
rect 192 -466 217 -431
rect 205 -477 217 -466
rect 269 -466 498 -431
rect 269 -477 478 -466
rect 204 -490 478 -477
rect 490 -490 498 -466
rect 732 -770 832 -722
rect 192 -1063 212 -1025
rect 264 -1063 832 -1025
rect 192 -1081 832 -1063
<< polycontact >>
rect 126 37 174 84
rect 807 -72 862 -25
rect 217 -477 269 -431
rect 212 -1063 264 -1016
<< metal1 >>
rect 0 529 1060 569
rect 0 483 78 529
rect 147 483 278 529
rect 347 483 498 529
rect 567 483 718 529
rect 787 483 918 529
rect 987 483 1060 529
rect 0 455 1060 483
rect 885 405 961 455
rect 99 355 961 405
rect 99 285 145 355
rect 507 285 553 355
rect 915 285 961 355
rect 270 249 369 265
rect 270 191 284 249
rect 358 191 369 249
rect 270 178 369 191
rect -52 84 185 85
rect -52 37 126 84
rect 174 37 185 84
rect -52 30 185 37
rect 303 84 349 132
rect 711 86 757 132
rect 711 84 886 86
rect 303 36 886 84
rect -52 -722 3 30
rect 786 -25 886 36
rect 302 -75 648 -26
rect 302 -288 351 -75
rect 599 -127 648 -75
rect 786 -72 807 -25
rect 862 -72 886 -25
rect 786 -80 886 -72
rect 599 -172 771 -127
rect 599 -226 695 -172
rect 663 -240 695 -226
rect 759 -195 771 -172
rect 1011 -170 1187 -155
rect 759 -240 770 -195
rect 663 -263 770 -240
rect 1011 -238 1024 -170
rect 1088 -238 1187 -170
rect 1011 -252 1187 -238
rect 99 -336 145 -290
rect 507 -336 553 -290
rect 915 -336 961 -290
rect 99 -382 961 -336
rect 205 -431 280 -429
rect 205 -477 217 -431
rect 269 -477 280 -431
rect 205 -490 280 -477
rect 81 -570 154 -558
rect 81 -623 95 -570
rect 153 -623 154 -570
rect 81 -635 154 -623
rect 211 -722 269 -490
rect 657 -540 703 -509
rect 329 -555 409 -542
rect 329 -617 331 -555
rect 398 -617 409 -555
rect 329 -629 409 -617
rect 494 -561 567 -549
rect 494 -614 507 -561
rect 565 -614 567 -561
rect 494 -626 567 -614
rect 657 -551 743 -540
rect 657 -608 671 -551
rect 731 -608 743 -551
rect 657 -620 743 -608
rect -52 -762 269 -722
rect -53 -770 269 -762
rect -53 -1026 -6 -770
rect 106 -853 212 -833
rect 657 -834 703 -620
rect 859 -665 906 -382
rect 859 -667 907 -665
rect 106 -919 118 -853
rect 189 -919 212 -853
rect 106 -932 212 -919
rect 510 -856 703 -834
rect 510 -922 526 -856
rect 597 -922 703 -856
rect 510 -927 703 -922
rect 205 -1016 273 -1003
rect 205 -1026 212 -1016
rect -53 -1063 212 -1026
rect 264 -1063 273 -1016
rect -53 -1073 273 -1063
rect 321 -1027 368 -953
rect 657 -977 703 -927
rect 860 -717 907 -667
rect 860 -763 1001 -717
rect 860 -953 906 -763
rect 861 -1027 908 -954
rect 321 -1067 908 -1027
rect 321 -1072 907 -1067
rect 321 -1075 906 -1072
rect 38 -1133 957 -1121
rect 38 -1160 743 -1133
rect 38 -1210 73 -1160
rect 168 -1210 273 -1160
rect 368 -1210 473 -1160
rect 568 -1210 673 -1160
rect 38 -1214 743 -1210
rect 850 -1214 957 -1133
rect 38 -1233 957 -1214
<< via1 >>
rect 284 191 358 249
rect 695 -240 759 -172
rect 1024 -238 1088 -170
rect 95 -623 153 -570
rect 331 -617 398 -555
rect 507 -614 565 -561
rect 671 -608 731 -551
rect 118 -919 189 -853
rect 526 -922 597 -856
rect 743 -1160 850 -1133
rect 743 -1210 768 -1160
rect 768 -1210 850 -1160
rect 743 -1214 850 -1210
<< metal2 >>
rect 270 265 375 270
rect 270 249 376 265
rect 270 191 284 249
rect 358 191 376 249
rect 270 -298 375 191
rect 663 -170 1111 -151
rect 663 -172 1024 -170
rect 663 -240 695 -172
rect 759 -238 1024 -172
rect 1088 -238 1111 -170
rect 759 -240 1111 -238
rect 663 -264 1111 -240
rect 80 -404 583 -298
rect 80 -550 190 -404
rect 373 -405 583 -404
rect 81 -570 190 -550
rect 81 -623 95 -570
rect 153 -623 190 -570
rect 81 -635 190 -623
rect 327 -542 408 -535
rect 327 -555 409 -542
rect 327 -617 331 -555
rect 398 -617 409 -555
rect 327 -629 409 -617
rect 490 -561 583 -405
rect 490 -614 507 -561
rect 565 -614 583 -561
rect 327 -682 408 -629
rect 490 -635 583 -614
rect 666 -551 757 -264
rect 1015 -265 1111 -264
rect 666 -608 671 -551
rect 731 -608 757 -551
rect 666 -620 757 -608
rect 325 -707 408 -682
rect 325 -708 807 -707
rect 325 -763 828 -708
rect 106 -853 703 -834
rect 106 -919 118 -853
rect 189 -856 703 -853
rect 189 -919 526 -856
rect 106 -922 526 -919
rect 597 -922 703 -856
rect 106 -932 703 -922
rect 772 -1126 828 -763
rect 731 -1133 867 -1126
rect 731 -1214 743 -1133
rect 850 -1214 867 -1133
rect 731 -1223 867 -1214
use nmos_3p3_UKFAHE  nmos_3p3_UKFAHE_0
timestamp 1691656227
transform 1 0 243 0 1 -898
box -162 -152 162 152
use nmos_3p3_UKFAHE  nmos_3p3_UKFAHE_1
timestamp 1691656227
transform 1 0 447 0 1 -898
box -162 -152 162 152
use nmos_3p3_UKFAHE  nmos_3p3_UKFAHE_2
timestamp 1691656227
transform 1 0 782 0 1 -594
box -162 -152 162 152
use nmos_3p3_UKFAHE  nmos_3p3_UKFAHE_3
timestamp 1691656227
transform 1 0 782 0 1 -898
box -162 -152 162 152
use nmos_3p3_UKFAHE  nmos_3p3_UKFAHE_4
timestamp 1691656227
transform 1 0 447 0 1 -594
box -162 -152 162 152
use nmos_3p3_UKFAHE  nmos_3p3_UKFAHE_5
timestamp 1691656227
transform 1 0 243 0 1 -594
box -162 -152 162 152
use pmos_3p3_YMKZL5  pmos_3p3_YMKZL5_0
timestamp 1691652503
transform 1 0 428 0 1 -208
box -224 -214 224 214
use pmos_3p3_YMKZL5  pmos_3p3_YMKZL5_1
timestamp 1691652503
transform 1 0 632 0 1 -208
box -224 -214 224 214
use pmos_3p3_YMKZL5  pmos_3p3_YMKZL5_2
timestamp 1691652503
transform 1 0 836 0 1 -208
box -224 -214 224 214
use pmos_3p3_YMKZL5  pmos_3p3_YMKZL5_3
timestamp 1691652503
transform 1 0 224 0 1 -208
box -224 -214 224 214
use pmos_3p3_YMKZL5  pmos_3p3_YMKZL5_4
timestamp 1691652503
transform 1 0 836 0 1 214
box -224 -214 224 214
use pmos_3p3_YMKZL5  pmos_3p3_YMKZL5_5
timestamp 1691652503
transform 1 0 632 0 1 214
box -224 -214 224 214
use pmos_3p3_YMKZL5  pmos_3p3_YMKZL5_6
timestamp 1691652503
transform 1 0 428 0 1 214
box -224 -214 224 214
use pmos_3p3_YMKZL5  pmos_3p3_YMKZL5_7
timestamp 1691652503
transform 1 0 224 0 1 214
box -224 -214 224 214
<< labels >>
flabel psubdiffcont 514 -1187 514 -1187 0 FreeSans 480 0 0 0 VSS
port 0 nsew
flabel metal1 1133 -218 1133 -218 0 FreeSans 480 0 0 0 OUT
port 1 nsew
flabel metal1 966 -741 966 -741 0 FreeSans 480 0 0 0 IN
port 2 nsew
flabel metal1 -37 -344 -37 -344 0 FreeSans 480 0 0 0 CLK
port 3 nsew
flabel nsubdiffcont 533 506 533 506 0 FreeSans 640 0 0 0 VDD
port 5 nsew
<< end >>
