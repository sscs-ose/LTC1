* NGSPICE file created from MSB_Unit_Cell_flat.ext - technology: gf180mcuC

.subckt MSB_Unit_Cell_flat IM VSS Ri Ci Ri-1 VDD QB Q OUT OUT+ OUT- SD IM_T
X0 OUT- QB.t3 OUT.t55 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 OUT IM_T.t0 SD.t48 VSS.t102 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X2 OUT+ Q.t3 OUT.t120 VSS.t33 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X3 VSS IM.t0 SD.t3 VSS.t43 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X4 Local_Enc_0.NAND_5.A Local_Enc_0.NAND_6.B VDD.t10 VDD.t9 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X5 OUT- QB.t4 OUT.t54 VSS.t21 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X6 OUT+ Q.t4 OUT.t121 VSS.t31 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X7 OUT Q.t5 OUT+.t61 VSS.t8 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X8 OUT- QB.t5 OUT.t53 VSS.t33 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X9 OUT+ Q.t6 OUT.t138 VSS.t10 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X10 OUT+ Q.t7 OUT.t15 VSS.t21 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X11 SD IM_T.t1 OUT.t10 VSS.t14 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X12 OUT+ Q.t8 OUT.t16 VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X13 SD IM_T.t2 OUT.t116 VSS.t63 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X14 OUT- QB.t6 OUT.t52 VSS.t19 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X15 OUT QB.t7 OUT-.t59 VSS.t32 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X16 OUT- QB.t8 OUT.t51 VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X17 OUT QB.t9 OUT-.t57 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X18 OUT Q.t9 OUT+.t57 VSS.t30 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X19 SD IM_T.t3 OUT.t92 VSS.t36 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X20 OUT Q.t10 OUT+.t56 VSS.t32 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X21 OUT Q.t11 OUT+.t55 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X22 OUT Q.t12 OUT+.t54 VSS.t9 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X23 OUT+ Q.t13 OUT.t104 VSS.t19 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X24 OUT+ Q.t14 OUT.t105 VSS.t28 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X25 OUT Q.t15 OUT+.t51 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X26 OUT QB.t10 OUT-.t56 VSS.t30 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X27 OUT QB.t11 OUT-.t55 VSS.t9 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X28 OUT- QB.t12 OUT.t50 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X29 OUT IM_T.t4 SD.t44 VSS.t105 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X30 OUT Q.t16 OUT+.t50 VSS.t29 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X31 OUT IM_T.t5 SD.t43 VSS.t78 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X32 OUT+ Q.t17 OUT.t123 VSS.t31 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X33 OUT Q.t18 OUT+.t48 VSS.t8 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X34 VSS IM.t1 SD.t58 VSS.t53 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X35 SD IM_T.t6 OUT.t126 VSS.t90 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X36 OUT+ Q.t19 OUT.t6 VSS.t10 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X37 OUT QB.t13 OUT-.t53 VSS.t29 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X38 Q Local_Enc_0.NAND_8.A Local_Enc_0.NAND_8.SD VSS.t49 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X39 OUT Q.t20 OUT+.t46 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X40 SD IM_T.t7 OUT.t131 VSS.t111 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X41 OUT IM_T.t8 SD.t40 VSS.t68 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X42 OUT+ Q.t21 OUT.t143 VSS.t28 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X43 Local_Enc_0.NAND_8.SD QB.t14 VSS.t35 VSS.t34 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X44 OUT+ Q.t22 OUT.t144 VSS.t33 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X45 OUT QB.t15 OUT-.t52 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X46 SD IM_T.t9 OUT.t127 VSS.t91 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X47 SD IM_T.t10 OUT.t133 VSS.t81 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X48 VSS IM.t2 SD.t2 VSS.t40 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X49 Local_Enc_0.NAND_8.A Local_Enc_0.NAND_5.B VDD.t26 VDD.t25 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X50 OUT- QB.t16 OUT.t49 VSS.t21 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X51 Local_Enc_0.NAND_6.SD Local_Enc_0.NAND_6.B VSS.t39 VSS.t38 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X52 OUT+ Q.t23 OUT.t149 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X53 SD IM.t3 VSS.t85 VSS.t12 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X54 OUT+ Q.t24 OUT.t150 VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X55 OUT+ Q.t25 OUT.t88 VSS.t21 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X56 OUT QB.t17 OUT-.t50 VSS.t32 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X57 OUT- QB.t18 OUT.t48 VSS.t31 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X58 OUT- QB.t19 OUT.t47 VSS.t19 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X59 SD IM.t4 VSS.t75 VSS.t74 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X60 OUT QB.t20 OUT-.t47 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X61 OUT- QB.t21 OUT.t46 VSS.t10 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X62 SD IM.t5 VSS.t118 VSS.t23 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X63 OUT Q.t26 OUT+.t40 VSS.t30 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X64 VDD Local_Enc_0.NAND_6.A Local_Enc_0.NAND_5.A VDD.t42 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X65 Local_Enc_0.NAND_6.B Ci.t0 VDD.t36 VDD.t35 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X66 VSS IM.t6 SD.t50 VSS.t24 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X67 OUT Q.t27 OUT+.t39 VSS.t9 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X68 OUT Q.t28 OUT+.t38 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X69 OUT IM_T.t11 SD.t37 VSS.t92 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X70 SD IM.t7 VSS.t112 VSS.t37 nfet_03v3 ad=0.312p pd=1.72u as=0.528p ps=3.28u w=1.2u l=0.5u
X71 OUT Q.t29 OUT+.t37 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X72 OUT QB.t22 OUT-.t45 VSS.t30 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X73 OUT QB.t23 OUT-.t44 VSS.t8 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X74 OUT+ Q.t30 OUT.t113 VSS.t33 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X75 OUT QB.t24 OUT-.t43 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X76 OUT QB.t25 OUT-.t42 VSS.t9 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X77 VDD Ci.t1 Local_Enc_0.NAND_6.B VDD.t32 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X78 OUT Q.t31 OUT+.t35 VSS.t29 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X79 OUT Q.t32 OUT+.t34 VSS.t8 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X80 VSS IM.t8 SD.t14 VSS.t56 nfet_03v3 ad=0.528p pd=3.28u as=0.312p ps=1.72u w=1.2u l=0.5u
X81 OUT+ Q.t33 OUT.t102 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X82 VSS IM.t9 SD.t0 VSS.t0 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X83 OUT+ Q.t34 OUT.t103 VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X84 OUT IM_T.t12 SD.t36 VSS.t108 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X85 SD IM_T.t13 OUT.t132 VSS.t97 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X86 OUT QB.t26 OUT-.t41 VSS.t32 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X87 OUT- QB.t27 OUT.t45 VSS.t31 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X88 OUT- QB.t28 OUT.t44 VSS.t19 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X89 OUT- QB.t29 OUT.t43 VSS.t28 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X90 VSS IM.t10 SD.t54 VSS.t102 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X91 OUT- QB.t30 OUT.t42 VSS.t10 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X92 OUT IM_T.t14 SD.t34 VSS.t43 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X93 OUT+ Q.t35 OUT.t122 VSS.t28 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X94 VDD Q.t36 QB.t1 VDD.t27 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X95 QB Q.t37 Local_Enc_0.NAND_4.SD VSS.t114 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X96 Local_Enc_0.NAND_6.A Ri.t0 VDD.t41 VDD.t40 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X97 Local_Enc_0.NAND_4.SD Local_Enc_0.NAND_4.B VSS.t27 VSS.t26 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X98 SD IM.t11 VSS.t84 VSS.t14 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X99 QB Local_Enc_0.NAND_4.B VDD.t6 VDD.t5 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X100 OUT- QB.t31 OUT.t41 VSS.t21 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X101 SD IM.t12 VSS.t117 VSS.t63 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X102 Local_Enc_0.NAND_5.SD Local_Enc_0.NAND_5.B VSS.t55 VSS.t54 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X103 OUT- QB.t32 OUT.t40 VSS.t33 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X104 VDD Ri.t1 Local_Enc_0.NAND_6.A VDD.t37 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X105 OUT Q.t38 OUT+.t30 VSS.t29 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X106 SD IM.t13 VSS.t88 VSS.t36 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X107 SD IM_T.t15 OUT.t129 VSS.t99 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X108 VSS IM.t14 SD.t63 VSS.t71 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X109 OUT- QB.t33 OUT.t39 VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X110 OUT QB.t34 OUT-.t33 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X111 OUT Q.t39 OUT+.t29 VSS.t30 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X112 SD IM_T.t16 OUT.t134 VSS.t72 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X113 OUT QB.t35 OUT-.t32 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X114 VDD Local_Enc_0.NAND_5.A Local_Enc_0.NAND_8.A VDD.t22 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X115 OUT Q.t40 OUT+.t28 VSS.t32 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X116 SD IM.t15 VSS.t89 VSS.t13 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X117 OUT Q.t41 OUT+.t27 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X118 OUT Q.t42 OUT+.t26 VSS.t9 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X119 OUT+ Q.t43 OUT.t158 VSS.t19 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X120 VSS IM.t16 SD.t55 VSS.t105 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X121 OUT Q.t44 OUT+.t24 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X122 OUT Q.t45 OUT+.t23 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X123 Local_Enc_0.NAND_5.A Local_Enc_0.NAND_6.A Local_Enc_0.NAND_6.SD VSS.t113 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X124 Local_Enc_0.NAND_2.SD Ci.t2 VSS.t52 VSS.t51 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X125 OUT IM_T.t17 SD.t31 VSS.t62 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X126 OUT QB.t36 OUT-.t31 VSS.t8 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X127 OUT QB.t37 OUT-.t30 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X128 SD IM_T.t18 OUT.t11 VSS.t18 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X129 OUT- QB.t38 OUT.t38 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X130 OUT IM_T.t19 SD.t29 VSS.t3 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X131 OUT- QB.t39 OUT.t37 VSS.t21 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X132 OUT+ Q.t46 OUT.t87 VSS.t31 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X133 OUT Q.t47 OUT+.t21 VSS.t8 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X134 Local_Enc_0.NAND_6.B Ci.t3 Local_Enc_0.NAND_2.SD VSS.t83 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X135 VSS IM.t17 SD.t5 VSS.t25 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X136 OUT+ Q.t48 OUT.t3 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X137 OUT- QB.t40 OUT.t36 VSS.t33 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X138 OUT+ Q.t49 OUT.t141 VSS.t10 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X139 OUT QB.t41 OUT-.t26 VSS.t29 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X140 OUT- QB.t42 OUT.t35 VSS.t31 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X141 OUT- QB.t43 OUT.t34 VSS.t28 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X142 OUT- QB.t44 OUT.t33 VSS.t10 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X143 OUT- QB.t45 OUT.t32 VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X144 SD IM.t18 VSS.t82 VSS.t81 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X145 OUT Q.t50 OUT+.t18 VSS.t30 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X146 OUT Q.t51 OUT+.t17 VSS.t32 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X147 OUT Q.t52 OUT+.t16 VSS.t9 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X148 OUT+ Q.t53 OUT.t156 VSS.t19 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X149 OUT+ Q.t54 OUT.t157 VSS.t28 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X150 SD IM_T.t20 OUT.t8 VSS.t12 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X151 Local_Enc_0.NAND_3.SD Ri.t2 VSS.t67 VSS.t66 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X152 Local_Enc_0.NAND_1.SD Local_Enc_0.NAND_1.B VSS.t17 VSS.t16 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X153 Local_Enc_0.NAND_5.B Local_Enc_0.NAND_1.B VDD.t4 VDD.t3 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X154 SD IM_T.t21 OUT.t17 VSS.t23 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X155 Local_Enc_0.NAND_6.A Ri.t3 Local_Enc_0.NAND_3.SD VSS.t59 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X156 OUT+ Q.t55 OUT.t99 VSS.t21 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X157 OUT IM_T.t22 SD.t26 VSS.t24 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X158 VSS IM.t19 SD.t49 VSS.t92 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X159 SD IM_T.t23 OUT.t93 VSS.t37 nfet_03v3 ad=0.312p pd=1.72u as=0.528p ps=3.28u w=1.2u l=0.5u
X160 OUT QB.t46 OUT-.t21 VSS.t29 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X161 OUT QB.t47 OUT-.t20 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X162 OUT QB.t48 OUT-.t19 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X163 VSS IM.t20 SD.t10 VSS.t78 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X164 OUT IM_T.t24 SD.t24 VSS.t53 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X165 VDD Local_Enc_0.NAND_8.A Local_Enc_0.NAND_4.B VDD.t19 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X166 Local_Enc_0.NAND_8.A Local_Enc_0.NAND_5.A Local_Enc_0.NAND_5.SD VSS.t50 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X167 SD IM.t21 VSS.t120 VSS.t90 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X168 OUT Q.t56 OUT+.t12 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X169 OUT Q.t57 OUT+.t11 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X170 OUT QB.t49 OUT-.t18 VSS.t30 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X171 Local_Enc_0.NAND_4.B Local_Enc_0.NAND_8.A VDD.t18 VDD.t17 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X172 Local_Enc_0.NAND_1.B Ri-1.t0 VDD.t31 VDD.t30 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X173 Local_Enc_0.NAND_0.SD Ri-1.t1 VSS.t65 VSS.t64 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X174 OUT QB.t50 OUT-.t17 VSS.t8 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X175 OUT IM_T.t25 SD.t23 VSS.t56 nfet_03v3 ad=0.528p pd=3.28u as=0.312p ps=1.72u w=1.2u l=0.5u
X176 OUT+ Q.t58 OUT.t96 VSS.t33 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X177 OUT QB.t51 OUT-.t16 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X178 OUT QB.t52 OUT-.t15 VSS.t9 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X179 OUT- QB.t53 OUT.t31 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X180 SD IM.t22 VSS.t119 VSS.t111 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X181 OUT- QB.t54 OUT.t30 VSS.t33 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X182 VDD Ri-1.t2 Local_Enc_0.NAND_1.B VDD.t11 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X183 Local_Enc_0.NAND_1.B Ri-1.t3 Local_Enc_0.NAND_0.SD VSS.t57 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X184 VSS IM.t23 SD.t6 VSS.t68 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X185 OUT+ Q.t59 OUT.t85 VSS.t31 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X186 OUT+ Q.t60 OUT.t1 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X187 SD IM.t24 VSS.t101 VSS.t91 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X188 OUT+ Q.t61 OUT.t155 VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X189 OUT IM_T.t26 SD.t22 VSS.t40 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X190 OUT+ Q.t62 OUT.t98 VSS.t10 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X191 OUT+ Q.t63 OUT.t94 VSS.t21 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X192 OUT QB.t55 OUT-.t12 VSS.t32 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X193 OUT- QB.t56 OUT.t29 VSS.t31 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X194 OUT- QB.t57 OUT.t28 VSS.t19 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X195 OUT- QB.t58 OUT.t27 VSS.t28 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X196 OUT- QB.t59 OUT.t26 VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X197 OUT- QB.t60 OUT.t25 VSS.t10 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X198 OUT QB.t61 OUT-.t6 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X199 OUT Q.t64 OUT+.t4 VSS.t32 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X200 OUT+ Q.t65 OUT.t12 VSS.t19 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X201 SD IM_T.t27 OUT.t125 VSS.t74 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X202 OUT QB.t62 OUT-.t5 VSS.t30 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X203 OUT QB.t63 OUT-.t4 VSS.t8 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X204 SD IM.t25 VSS.t100 VSS.t99 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X205 OUT QB.t64 OUT-.t3 VSS.t9 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X206 OUT Q.t66 OUT+.t2 VSS.t29 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X207 OUT IM_T.t28 SD.t20 VSS.t71 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X208 SD IM.t26 VSS.t73 VSS.t72 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X209 SD IM_T.t29 OUT.t9 VSS.t13 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X210 OUT QB.t65 OUT-.t2 VSS.t29 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X211 OUT QB.t66 OUT-.t1 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X212 VSS IM.t27 SD.t9 VSS.t62 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X213 OUT- QB.t67 OUT.t24 VSS.t28 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X214 VDD Local_Enc_0.NAND_8.A Q.t1 VDD.t14 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X215 OUT Q.t67 OUT+.t1 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X216 VSS IM.t28 SD.t1 VSS.t3 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X217 SD IM.t29 VSS.t58 VSS.t18 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X218 OUT Q.t68 OUT+.t0 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X219 OUT IM_T.t30 SD.t18 VSS.t0 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X220 Local_Enc_0.NAND_5.B Local_Enc_0.NAND_1.B Local_Enc_0.NAND_1.SD VSS.t15 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X221 Q QB.t68 VDD.t8 VDD.t7 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X222 OUT IM_T.t31 SD.t17 VSS.t25 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X223 Local_Enc_0.NAND_4.B Local_Enc_0.NAND_8.A Local_Enc_0.NAND_7.SD VSS.t48 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X224 VDD Local_Enc_0.NAND_1.B Local_Enc_0.NAND_5.B VDD.t0 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X225 VSS IM.t30 SD.t56 VSS.t108 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X226 SD IM.t31 VSS.t98 VSS.t97 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X227 Local_Enc_0.NAND_7.SD Local_Enc_0.NAND_8.A VSS.t47 VSS.t46 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
R0 QB.n4 QB.t14 26.9784
R1 QB.n20 QB.t29 24.9712
R2 QB.n35 QB.t58 24.9712
R3 QB.n50 QB.t43 24.9712
R4 QB.n5 QB.t67 24.9712
R5 QB.n65 QB.n64 21.4076
R6 QB.n67 QB.n19 21.1997
R7 QB.n66 QB.n34 20.1581
R8 QB.n65 QB.n49 20.1567
R9 QB.n22 QB.t23 15.1115
R10 QB.n23 QB.t57 15.1115
R11 QB.n26 QB.t34 15.1115
R12 QB.n27 QB.t4 15.1115
R13 QB.n30 QB.t20 15.1115
R14 QB.n31 QB.t38 15.1115
R15 QB.n37 QB.t50 15.1115
R16 QB.n38 QB.t19 15.1115
R17 QB.n41 QB.t66 15.1115
R18 QB.n42 QB.t31 15.1115
R19 QB.n45 QB.t47 15.1115
R20 QB.n46 QB.t3 15.1115
R21 QB.n52 QB.t36 15.1115
R22 QB.n53 QB.t6 15.1115
R23 QB.n56 QB.t48 15.1115
R24 QB.n57 QB.t16 15.1115
R25 QB.n60 QB.t35 15.1115
R26 QB.n61 QB.t53 15.1115
R27 QB.n7 QB.t63 15.1115
R28 QB.n8 QB.t28 15.1115
R29 QB.n11 QB.t9 15.1115
R30 QB.n12 QB.t39 15.1115
R31 QB.n15 QB.t61 15.1115
R32 QB.n16 QB.t12 15.1115
R33 QB.n4 QB.t68 14.7248
R34 QB.n20 QB.t46 14.4545
R35 QB.n21 QB.t45 14.4545
R36 QB.n24 QB.t64 14.4545
R37 QB.n25 QB.t30 14.4545
R38 QB.n28 QB.t24 14.4545
R39 QB.n29 QB.t40 14.4545
R40 QB.n32 QB.t62 14.4545
R41 QB.n33 QB.t27 14.4545
R42 QB.n35 QB.t13 14.4545
R43 QB.n36 QB.t8 14.4545
R44 QB.n39 QB.t25 14.4545
R45 QB.n40 QB.t60 14.4545
R46 QB.n43 QB.t51 14.4545
R47 QB.n44 QB.t5 14.4545
R48 QB.n47 QB.t22 14.4545
R49 QB.n48 QB.t56 14.4545
R50 QB.n50 QB.t41 14.4545
R51 QB.n51 QB.t33 14.4545
R52 QB.n54 QB.t52 14.4545
R53 QB.n55 QB.t21 14.4545
R54 QB.n58 QB.t15 14.4545
R55 QB.n59 QB.t32 14.4545
R56 QB.n62 QB.t49 14.4545
R57 QB.n63 QB.t18 14.4545
R58 QB.n5 QB.t65 14.4545
R59 QB.n6 QB.t59 14.4545
R60 QB.n9 QB.t11 14.4545
R61 QB.n10 QB.t44 14.4545
R62 QB.n13 QB.t37 14.4545
R63 QB.n14 QB.t54 14.4545
R64 QB.n17 QB.t10 14.4545
R65 QB.n18 QB.t42 14.4545
R66 QB.n34 QB.n33 12.7802
R67 QB.n49 QB.n48 12.7802
R68 QB.n64 QB.n63 12.7802
R69 QB.n19 QB.n18 12.7802
R70 QB.n34 QB.t55 12.1915
R71 QB.n49 QB.t17 12.1915
R72 QB.n64 QB.t7 12.1915
R73 QB.n19 QB.t26 12.1915
R74 QB.n21 QB.n20 9.86024
R75 QB.n22 QB.n21 9.86024
R76 QB.n23 QB.n22 9.86024
R77 QB.n24 QB.n23 9.86024
R78 QB.n25 QB.n24 9.86024
R79 QB.n26 QB.n25 9.86024
R80 QB.n27 QB.n26 9.86024
R81 QB.n28 QB.n27 9.86024
R82 QB.n29 QB.n28 9.86024
R83 QB.n30 QB.n29 9.86024
R84 QB.n31 QB.n30 9.86024
R85 QB.n32 QB.n31 9.86024
R86 QB.n33 QB.n32 9.86024
R87 QB.n36 QB.n35 9.86024
R88 QB.n37 QB.n36 9.86024
R89 QB.n38 QB.n37 9.86024
R90 QB.n39 QB.n38 9.86024
R91 QB.n40 QB.n39 9.86024
R92 QB.n41 QB.n40 9.86024
R93 QB.n42 QB.n41 9.86024
R94 QB.n43 QB.n42 9.86024
R95 QB.n44 QB.n43 9.86024
R96 QB.n45 QB.n44 9.86024
R97 QB.n46 QB.n45 9.86024
R98 QB.n47 QB.n46 9.86024
R99 QB.n48 QB.n47 9.86024
R100 QB.n51 QB.n50 9.86024
R101 QB.n52 QB.n51 9.86024
R102 QB.n53 QB.n52 9.86024
R103 QB.n54 QB.n53 9.86024
R104 QB.n55 QB.n54 9.86024
R105 QB.n56 QB.n55 9.86024
R106 QB.n57 QB.n56 9.86024
R107 QB.n58 QB.n57 9.86024
R108 QB.n59 QB.n58 9.86024
R109 QB.n60 QB.n59 9.86024
R110 QB.n61 QB.n60 9.86024
R111 QB.n62 QB.n61 9.86024
R112 QB.n63 QB.n62 9.86024
R113 QB.n6 QB.n5 9.86024
R114 QB.n7 QB.n6 9.86024
R115 QB.n8 QB.n7 9.86024
R116 QB.n9 QB.n8 9.86024
R117 QB.n10 QB.n9 9.86024
R118 QB.n11 QB.n10 9.86024
R119 QB.n12 QB.n11 9.86024
R120 QB.n13 QB.n12 9.86024
R121 QB.n14 QB.n13 9.86024
R122 QB.n15 QB.n14 9.86024
R123 QB.n16 QB.n15 9.86024
R124 QB.n17 QB.n16 9.86024
R125 QB.n18 QB.n17 9.86024
R126 QB.n68 QB 8.0222
R127 QB.n3 QB.n0 6.8765
R128 QB QB.n4 4.18544
R129 QB.n2 QB.t1 3.6405
R130 QB.n2 QB.n1 3.6405
R131 QB.n3 QB.n2 3.08447
R132 QB.n69 QB.n68 2.2505
R133 QB.n66 QB.n65 1.23881
R134 QB QB.n67 0.749429
R135 QB.n69 QB 0.241152
R136 QB.n67 QB.n66 0.182313
R137 QB QB.n3 0.17463
R138 QB QB.n69 0.112881
R139 QB.n68 QB 0.10226
R140 OUT.n228 OUT.t93 5.37963
R141 OUT.n243 OUT.n197 4.86963
R142 OUT OUT.n196 4.78467
R143 OUT.n70 OUT.n69 3.9342
R144 OUT.n65 OUT.n64 3.9339
R145 OUT.n190 OUT.n189 3.78102
R146 OUT.n228 OUT.n227 3.61615
R147 OUT.n230 OUT.n223 3.61615
R148 OUT.n232 OUT.n219 3.61615
R149 OUT.n234 OUT.n215 3.61615
R150 OUT.n236 OUT.n211 3.61615
R151 OUT.n238 OUT.n207 3.61615
R152 OUT.n240 OUT.n203 3.61615
R153 OUT.n242 OUT.n199 3.61615
R154 OUT.n126 OUT.n125 3.50723
R155 OUT.n105 OUT.n104 3.50723
R156 OUT.n84 OUT.n83 3.50723
R157 OUT.n70 OUT.n67 3.50518
R158 OUT.n127 OUT.n121 3.50518
R159 OUT.n106 OUT.n100 3.50518
R160 OUT.n85 OUT.n79 3.50518
R161 OUT.n241 OUT.n201 3.50463
R162 OUT.n239 OUT.n205 3.50463
R163 OUT.n237 OUT.n209 3.50463
R164 OUT.n235 OUT.n213 3.50463
R165 OUT.n233 OUT.n217 3.50463
R166 OUT.n231 OUT.n221 3.50463
R167 OUT.n229 OUT.n225 3.50463
R168 OUT.n22 OUT.n16 3.5031
R169 OUT.n21 OUT.n20 3.5031
R170 OUT.n36 OUT.n30 3.5031
R171 OUT.n35 OUT.n34 3.5031
R172 OUT.n53 OUT.n47 3.5031
R173 OUT.n52 OUT.n51 3.5031
R174 OUT.n65 OUT.n62 3.5031
R175 OUT.n22 OUT.n14 3.41897
R176 OUT.n21 OUT.n18 3.41897
R177 OUT.n36 OUT.n28 3.41897
R178 OUT.n35 OUT.n32 3.41897
R179 OUT.n53 OUT.n45 3.41897
R180 OUT.n52 OUT.n49 3.41897
R181 OUT.n126 OUT.n123 3.41897
R182 OUT.n127 OUT.n119 3.41897
R183 OUT.n105 OUT.n102 3.41897
R184 OUT.n106 OUT.n98 3.41897
R185 OUT.n84 OUT.n81 3.41897
R186 OUT.n85 OUT.n77 3.41897
R187 OUT.n196 OUT.n1 3.37397
R188 OUT.n195 OUT.n3 3.37397
R189 OUT.n190 OUT.n187 3.37397
R190 OUT.n88 OUT.n87 3.1505
R191 OUT.n91 OUT.n90 3.1505
R192 OUT.n109 OUT.n108 3.1505
R193 OUT.n112 OUT.n111 3.1505
R194 OUT.n130 OUT.n129 3.1505
R195 OUT.n133 OUT.n132 3.1505
R196 OUT.n136 OUT.n135 3.1505
R197 OUT.n6 OUT.n5 3.1505
R198 OUT.n148 OUT.n75 3.1505
R199 OUT.n149 OUT.n73 3.1505
R200 OUT.n145 OUT.n96 3.1505
R201 OUT.n146 OUT.n94 3.1505
R202 OUT.n142 OUT.n117 3.1505
R203 OUT.n143 OUT.n115 3.1505
R204 OUT.n9 OUT.n8 3.1505
R205 OUT.n140 OUT.n139 3.1505
R206 OUT.n155 OUT.n154 3.1505
R207 OUT.n156 OUT.n152 3.1505
R208 OUT.n58 OUT.n57 3.1505
R209 OUT.n59 OUT.n55 3.1505
R210 OUT.n41 OUT.n40 3.1505
R211 OUT.n42 OUT.n38 3.1505
R212 OUT.n12 OUT.n11 3.1505
R213 OUT.n25 OUT.n24 3.1505
R214 OUT.n164 OUT.n163 3.1505
R215 OUT.n161 OUT.n160 3.1505
R216 OUT.n171 OUT.n170 3.1505
R217 OUT.n168 OUT.n167 3.1505
R218 OUT.n178 OUT.n177 3.1505
R219 OUT.n175 OUT.n174 3.1505
R220 OUT.n185 OUT.n184 3.1505
R221 OUT.n182 OUT.n181 3.1505
R222 OUT.n1 OUT.t34 2.7305
R223 OUT.n1 OUT.n0 2.7305
R224 OUT.n3 OUT.t16 2.7305
R225 OUT.n3 OUT.n2 2.7305
R226 OUT.n181 OUT.t40 2.7305
R227 OUT.n181 OUT.n180 2.7305
R228 OUT.n184 OUT.t120 2.7305
R229 OUT.n184 OUT.n183 2.7305
R230 OUT.n174 OUT.t53 2.7305
R231 OUT.n174 OUT.n173 2.7305
R232 OUT.n177 OUT.t144 2.7305
R233 OUT.n177 OUT.n176 2.7305
R234 OUT.n167 OUT.t36 2.7305
R235 OUT.n167 OUT.n166 2.7305
R236 OUT.n170 OUT.t96 2.7305
R237 OUT.n170 OUT.n169 2.7305
R238 OUT.n160 OUT.t30 2.7305
R239 OUT.n160 OUT.n159 2.7305
R240 OUT.n163 OUT.t113 2.7305
R241 OUT.n163 OUT.n162 2.7305
R242 OUT.n16 OUT.t149 2.7305
R243 OUT.n16 OUT.n15 2.7305
R244 OUT.n14 OUT.t55 2.7305
R245 OUT.n14 OUT.n13 2.7305
R246 OUT.n20 OUT.t48 2.7305
R247 OUT.n20 OUT.n19 2.7305
R248 OUT.n18 OUT.t121 2.7305
R249 OUT.n18 OUT.n17 2.7305
R250 OUT.n30 OUT.t1 2.7305
R251 OUT.n30 OUT.n29 2.7305
R252 OUT.n28 OUT.t38 2.7305
R253 OUT.n28 OUT.n27 2.7305
R254 OUT.n34 OUT.t29 2.7305
R255 OUT.n34 OUT.n33 2.7305
R256 OUT.n32 OUT.t87 2.7305
R257 OUT.n32 OUT.n31 2.7305
R258 OUT.n47 OUT.t102 2.7305
R259 OUT.n47 OUT.n46 2.7305
R260 OUT.n45 OUT.t50 2.7305
R261 OUT.n45 OUT.n44 2.7305
R262 OUT.n51 OUT.t45 2.7305
R263 OUT.n51 OUT.n50 2.7305
R264 OUT.n49 OUT.t123 2.7305
R265 OUT.n49 OUT.n48 2.7305
R266 OUT.n24 OUT.t99 2.7305
R267 OUT.n24 OUT.n23 2.7305
R268 OUT.n11 OUT.t49 2.7305
R269 OUT.n11 OUT.n10 2.7305
R270 OUT.n38 OUT.t88 2.7305
R271 OUT.n38 OUT.n37 2.7305
R272 OUT.n40 OUT.t41 2.7305
R273 OUT.n40 OUT.n39 2.7305
R274 OUT.n55 OUT.t94 2.7305
R275 OUT.n55 OUT.n54 2.7305
R276 OUT.n57 OUT.t54 2.7305
R277 OUT.n57 OUT.n56 2.7305
R278 OUT.n152 OUT.t15 2.7305
R279 OUT.n152 OUT.n151 2.7305
R280 OUT.n154 OUT.t37 2.7305
R281 OUT.n154 OUT.n153 2.7305
R282 OUT.n139 OUT.t46 2.7305
R283 OUT.n139 OUT.n138 2.7305
R284 OUT.n8 OUT.t98 2.7305
R285 OUT.n8 OUT.n7 2.7305
R286 OUT.n115 OUT.t25 2.7305
R287 OUT.n115 OUT.n114 2.7305
R288 OUT.n117 OUT.t138 2.7305
R289 OUT.n117 OUT.n116 2.7305
R290 OUT.n94 OUT.t42 2.7305
R291 OUT.n94 OUT.n93 2.7305
R292 OUT.n96 OUT.t141 2.7305
R293 OUT.n96 OUT.n95 2.7305
R294 OUT.n73 OUT.t33 2.7305
R295 OUT.n73 OUT.n72 2.7305
R296 OUT.n75 OUT.t6 2.7305
R297 OUT.n75 OUT.n74 2.7305
R298 OUT.n67 OUT.t26 2.7305
R299 OUT.n67 OUT.n66 2.7305
R300 OUT.n69 OUT.t122 2.7305
R301 OUT.n69 OUT.n68 2.7305
R302 OUT.n5 OUT.t52 2.7305
R303 OUT.n5 OUT.n4 2.7305
R304 OUT.n135 OUT.t158 2.7305
R305 OUT.n135 OUT.n134 2.7305
R306 OUT.n132 OUT.t47 2.7305
R307 OUT.n132 OUT.n131 2.7305
R308 OUT.n129 OUT.t104 2.7305
R309 OUT.n129 OUT.n128 2.7305
R310 OUT.n111 OUT.t28 2.7305
R311 OUT.n111 OUT.n110 2.7305
R312 OUT.n108 OUT.t156 2.7305
R313 OUT.n108 OUT.n107 2.7305
R314 OUT.n90 OUT.t44 2.7305
R315 OUT.n90 OUT.n89 2.7305
R316 OUT.n87 OUT.t12 2.7305
R317 OUT.n87 OUT.n86 2.7305
R318 OUT.n125 OUT.t105 2.7305
R319 OUT.n125 OUT.n124 2.7305
R320 OUT.n123 OUT.t27 2.7305
R321 OUT.n123 OUT.n122 2.7305
R322 OUT.n121 OUT.t39 2.7305
R323 OUT.n121 OUT.n120 2.7305
R324 OUT.n119 OUT.t150 2.7305
R325 OUT.n119 OUT.n118 2.7305
R326 OUT.n104 OUT.t157 2.7305
R327 OUT.n104 OUT.n103 2.7305
R328 OUT.n102 OUT.t43 2.7305
R329 OUT.n102 OUT.n101 2.7305
R330 OUT.n100 OUT.t51 2.7305
R331 OUT.n100 OUT.n99 2.7305
R332 OUT.n98 OUT.t155 2.7305
R333 OUT.n98 OUT.n97 2.7305
R334 OUT.n83 OUT.t143 2.7305
R335 OUT.n83 OUT.n82 2.7305
R336 OUT.n81 OUT.t24 2.7305
R337 OUT.n81 OUT.n80 2.7305
R338 OUT.n79 OUT.t32 2.7305
R339 OUT.n79 OUT.n78 2.7305
R340 OUT.n77 OUT.t103 2.7305
R341 OUT.n77 OUT.n76 2.7305
R342 OUT.n64 OUT.t35 2.7305
R343 OUT.n64 OUT.n63 2.7305
R344 OUT.n62 OUT.t3 2.7305
R345 OUT.n62 OUT.n61 2.7305
R346 OUT.n187 OUT.t31 2.7305
R347 OUT.n187 OUT.n186 2.7305
R348 OUT.n189 OUT.t85 2.7305
R349 OUT.n189 OUT.n188 2.7305
R350 OUT.n201 OUT.t17 1.3655
R351 OUT.n201 OUT.n200 1.3655
R352 OUT.n205 OUT.t127 1.3655
R353 OUT.n205 OUT.n204 1.3655
R354 OUT.n209 OUT.t8 1.3655
R355 OUT.n209 OUT.n208 1.3655
R356 OUT.n213 OUT.t131 1.3655
R357 OUT.n213 OUT.n212 1.3655
R358 OUT.n217 OUT.t132 1.3655
R359 OUT.n217 OUT.n216 1.3655
R360 OUT.n221 OUT.t9 1.3655
R361 OUT.n221 OUT.n220 1.3655
R362 OUT.n225 OUT.t126 1.3655
R363 OUT.n225 OUT.n224 1.3655
R364 OUT.n227 OUT.t92 1.3655
R365 OUT.n227 OUT.n226 1.3655
R366 OUT.n223 OUT.t134 1.3655
R367 OUT.n223 OUT.n222 1.3655
R368 OUT.n219 OUT.t133 1.3655
R369 OUT.n219 OUT.n218 1.3655
R370 OUT.n215 OUT.t11 1.3655
R371 OUT.n215 OUT.n214 1.3655
R372 OUT.n211 OUT.t10 1.3655
R373 OUT.n211 OUT.n210 1.3655
R374 OUT.n207 OUT.t129 1.3655
R375 OUT.n207 OUT.n206 1.3655
R376 OUT.n203 OUT.t116 1.3655
R377 OUT.n203 OUT.n202 1.3655
R378 OUT.n199 OUT.t125 1.3655
R379 OUT.n199 OUT.n198 1.3655
R380 OUT.n22 OUT.n21 0.583357
R381 OUT.n36 OUT.n35 0.583357
R382 OUT.n53 OUT.n52 0.583357
R383 OUT.n127 OUT.n126 0.583357
R384 OUT.n106 OUT.n105 0.583357
R385 OUT.n85 OUT.n84 0.583357
R386 OUT.n137 OUT.n127 0.521929
R387 OUT.n113 OUT.n106 0.521929
R388 OUT.n92 OUT.n85 0.521929
R389 OUT.n179 OUT.n22 0.5105
R390 OUT.n172 OUT.n36 0.5105
R391 OUT.n165 OUT.n53 0.5105
R392 OUT.n243 OUT.n242 0.5105
R393 OUT.n242 OUT.n241 0.5105
R394 OUT.n241 OUT.n240 0.5105
R395 OUT.n240 OUT.n239 0.5105
R396 OUT.n239 OUT.n238 0.5105
R397 OUT.n238 OUT.n237 0.5105
R398 OUT.n237 OUT.n236 0.5105
R399 OUT.n236 OUT.n235 0.5105
R400 OUT.n235 OUT.n234 0.5105
R401 OUT.n234 OUT.n233 0.5105
R402 OUT.n233 OUT.n232 0.5105
R403 OUT.n232 OUT.n231 0.5105
R404 OUT.n231 OUT.n230 0.5105
R405 OUT.n230 OUT.n229 0.5105
R406 OUT.n229 OUT.n228 0.5105
R407 OUT.n141 OUT.n26 0.463357
R408 OUT.n144 OUT.n43 0.463357
R409 OUT.n147 OUT.n60 0.463357
R410 OUT.n179 OUT.n26 0.454786
R411 OUT.n172 OUT.n43 0.454786
R412 OUT.n165 OUT.n60 0.454786
R413 OUT.n141 OUT.n137 0.446214
R414 OUT.n144 OUT.n113 0.446214
R415 OUT.n147 OUT.n92 0.446214
R416 OUT.n193 OUT.n192 0.41094
R417 OUT.n195 OUT.n194 0.406984
R418 OUT.n192 OUT.n191 0.405005
R419 OUT.n196 OUT.n195 0.404016
R420 OUT.n91 OUT.n88 0.401049
R421 OUT.n112 OUT.n109 0.401049
R422 OUT.n133 OUT.n130 0.401049
R423 OUT.n136 OUT.n6 0.401049
R424 OUT.n149 OUT.n148 0.401049
R425 OUT.n146 OUT.n145 0.401049
R426 OUT.n143 OUT.n142 0.401049
R427 OUT.n140 OUT.n9 0.401049
R428 OUT.n156 OUT.n155 0.401049
R429 OUT.n59 OUT.n58 0.401049
R430 OUT.n42 OUT.n41 0.401049
R431 OUT.n25 OUT.n12 0.401049
R432 OUT.n164 OUT.n161 0.401049
R433 OUT.n171 OUT.n168 0.401049
R434 OUT.n178 OUT.n175 0.401049
R435 OUT.n185 OUT.n182 0.401049
R436 OUT.n194 OUT.n193 0.399071
R437 OUT.n191 OUT.n190 0.398082
R438 OUT.n71 OUT.n70 0.382477
R439 OUT.n158 OUT.n65 0.374105
R440 OUT.n157 OUT.n150 0.33957
R441 OUT OUT.n243 0.33675
R442 OUT.n158 OUT.n157 0.333291
R443 OUT.n150 OUT.n71 0.327012
R444 OUT.n88 OUT.n71 0.226984
R445 OUT.n150 OUT.n149 0.226984
R446 OUT.n157 OUT.n156 0.226984
R447 OUT.n161 OUT.n158 0.226984
R448 OUT.n109 OUT.n92 0.215115
R449 OUT.n130 OUT.n113 0.215115
R450 OUT.n137 OUT.n136 0.215115
R451 OUT.n147 OUT.n146 0.215115
R452 OUT.n144 OUT.n143 0.215115
R453 OUT.n141 OUT.n140 0.215115
R454 OUT.n60 OUT.n59 0.215115
R455 OUT.n43 OUT.n42 0.215115
R456 OUT.n26 OUT.n25 0.215115
R457 OUT.n168 OUT.n165 0.215115
R458 OUT.n175 OUT.n172 0.215115
R459 OUT.n182 OUT.n179 0.215115
R460 OUT.n92 OUT.n91 0.173577
R461 OUT.n113 OUT.n112 0.173577
R462 OUT.n137 OUT.n133 0.173577
R463 OUT.n148 OUT.n147 0.173577
R464 OUT.n145 OUT.n144 0.173577
R465 OUT.n142 OUT.n141 0.173577
R466 OUT.n155 OUT.n60 0.173577
R467 OUT.n58 OUT.n43 0.173577
R468 OUT.n41 OUT.n26 0.173577
R469 OUT.n165 OUT.n164 0.173577
R470 OUT.n172 OUT.n171 0.173577
R471 OUT.n179 OUT.n178 0.173577
R472 OUT.n194 OUT.n6 0.119181
R473 OUT.n193 OUT.n9 0.119181
R474 OUT.n192 OUT.n12 0.119181
R475 OUT.n191 OUT.n185 0.119181
R476 OUT-.n87 OUT-.t59 9.52957
R477 OUT-.n64 OUT-.t50 9.52957
R478 OUT-.n41 OUT-.t12 9.52957
R479 OUT-.n18 OUT-.t41 9.52957
R480 OUT-.n91 OUT-.n69 8.25388
R481 OUT-.n68 OUT-.n46 8.25388
R482 OUT-.n45 OUT-.n23 8.25388
R483 OUT-.n22 OUT-.n0 8.25388
R484 OUT-.n76 OUT-.n75 6.83298
R485 OUT-.n53 OUT-.n52 6.83298
R486 OUT-.n30 OUT-.n29 6.83298
R487 OUT-.n7 OUT-.n6 6.83298
R488 OUT-.n80 OUT-.n79 5.5481
R489 OUT-.n77 OUT-.n71 5.5481
R490 OUT-.n76 OUT-.n73 5.5481
R491 OUT-.n57 OUT-.n56 5.5481
R492 OUT-.n54 OUT-.n48 5.5481
R493 OUT-.n53 OUT-.n50 5.5481
R494 OUT-.n34 OUT-.n33 5.5481
R495 OUT-.n31 OUT-.n25 5.5481
R496 OUT-.n30 OUT-.n27 5.5481
R497 OUT-.n11 OUT-.n10 5.5481
R498 OUT-.n8 OUT-.n2 5.5481
R499 OUT-.n7 OUT-.n4 5.5481
R500 OUT-.n87 OUT-.n86 5.53001
R501 OUT-.n64 OUT-.n63 5.53001
R502 OUT-.n41 OUT-.n40 5.53001
R503 OUT-.n18 OUT-.n17 5.53001
R504 OUT-.n88 OUT-.n84 5.52516
R505 OUT-.n65 OUT-.n61 5.52516
R506 OUT-.n42 OUT-.n38 5.52516
R507 OUT-.n19 OUT-.n15 5.52516
R508 OUT-.n89 OUT-.n82 5.51961
R509 OUT-.n66 OUT-.n59 5.51961
R510 OUT-.n43 OUT-.n36 5.51961
R511 OUT-.n20 OUT-.n13 5.51961
R512 OUT-.n82 OUT-.t31 2.7305
R513 OUT-.n82 OUT-.n81 2.7305
R514 OUT-.n84 OUT-.t19 2.7305
R515 OUT-.n84 OUT-.n83 2.7305
R516 OUT-.n86 OUT-.t32 2.7305
R517 OUT-.n86 OUT-.n85 2.7305
R518 OUT-.n79 OUT-.t26 2.7305
R519 OUT-.n79 OUT-.n78 2.7305
R520 OUT-.n71 OUT-.t15 2.7305
R521 OUT-.n71 OUT-.n70 2.7305
R522 OUT-.n73 OUT-.t52 2.7305
R523 OUT-.n73 OUT-.n72 2.7305
R524 OUT-.n75 OUT-.t18 2.7305
R525 OUT-.n75 OUT-.n74 2.7305
R526 OUT-.n59 OUT-.t17 2.7305
R527 OUT-.n59 OUT-.n58 2.7305
R528 OUT-.n61 OUT-.t1 2.7305
R529 OUT-.n61 OUT-.n60 2.7305
R530 OUT-.n63 OUT-.t20 2.7305
R531 OUT-.n63 OUT-.n62 2.7305
R532 OUT-.n56 OUT-.t53 2.7305
R533 OUT-.n56 OUT-.n55 2.7305
R534 OUT-.n48 OUT-.t42 2.7305
R535 OUT-.n48 OUT-.n47 2.7305
R536 OUT-.n50 OUT-.t16 2.7305
R537 OUT-.n50 OUT-.n49 2.7305
R538 OUT-.n52 OUT-.t45 2.7305
R539 OUT-.n52 OUT-.n51 2.7305
R540 OUT-.n36 OUT-.t44 2.7305
R541 OUT-.n36 OUT-.n35 2.7305
R542 OUT-.n38 OUT-.t33 2.7305
R543 OUT-.n38 OUT-.n37 2.7305
R544 OUT-.n40 OUT-.t47 2.7305
R545 OUT-.n40 OUT-.n39 2.7305
R546 OUT-.n33 OUT-.t21 2.7305
R547 OUT-.n33 OUT-.n32 2.7305
R548 OUT-.n25 OUT-.t3 2.7305
R549 OUT-.n25 OUT-.n24 2.7305
R550 OUT-.n27 OUT-.t43 2.7305
R551 OUT-.n27 OUT-.n26 2.7305
R552 OUT-.n29 OUT-.t5 2.7305
R553 OUT-.n29 OUT-.n28 2.7305
R554 OUT-.n13 OUT-.t4 2.7305
R555 OUT-.n13 OUT-.n12 2.7305
R556 OUT-.n15 OUT-.t57 2.7305
R557 OUT-.n15 OUT-.n14 2.7305
R558 OUT-.n17 OUT-.t6 2.7305
R559 OUT-.n17 OUT-.n16 2.7305
R560 OUT-.n10 OUT-.t2 2.7305
R561 OUT-.n10 OUT-.n9 2.7305
R562 OUT-.n2 OUT-.t55 2.7305
R563 OUT-.n2 OUT-.n1 2.7305
R564 OUT-.n4 OUT-.t30 2.7305
R565 OUT-.n4 OUT-.n3 2.7305
R566 OUT-.n6 OUT-.t56 2.7305
R567 OUT-.n6 OUT-.n5 2.7305
R568 OUT-.n96 OUT-.n95 2.25828
R569 OUT-.n89 OUT-.n88 1.28037
R570 OUT-.n66 OUT-.n65 1.28037
R571 OUT-.n43 OUT-.n42 1.28037
R572 OUT-.n20 OUT-.n19 1.28037
R573 OUT-.n77 OUT-.n76 1.27854
R574 OUT-.n54 OUT-.n53 1.27854
R575 OUT-.n31 OUT-.n30 1.27854
R576 OUT-.n8 OUT-.n7 1.27854
R577 OUT-.n80 OUT-.n77 1.27492
R578 OUT-.n57 OUT-.n54 1.27492
R579 OUT-.n34 OUT-.n31 1.27492
R580 OUT-.n11 OUT-.n8 1.27492
R581 OUT-.n88 OUT-.n87 1.26834
R582 OUT-.n65 OUT-.n64 1.26834
R583 OUT-.n42 OUT-.n41 1.26834
R584 OUT-.n19 OUT-.n18 1.26834
R585 OUT-.n96 OUT-.n94 0.915071
R586 OUT-.n92 OUT-.n91 0.832625
R587 OUT-.n94 OUT-.n93 0.687929
R588 OUT-.n93 OUT-.n92 0.686214
R589 OUT-.n91 OUT-.n90 0.637571
R590 OUT-.n68 OUT-.n67 0.637571
R591 OUT-.n45 OUT-.n44 0.637571
R592 OUT-.n22 OUT-.n21 0.637571
R593 OUT-.n90 OUT-.n89 0.636636
R594 OUT-.n67 OUT-.n66 0.636636
R595 OUT-.n44 OUT-.n43 0.636636
R596 OUT-.n21 OUT-.n20 0.636636
R597 OUT-.n90 OUT-.n80 0.550143
R598 OUT-.n67 OUT-.n57 0.550143
R599 OUT-.n44 OUT-.n34 0.550143
R600 OUT-.n21 OUT-.n11 0.550143
R601 OUT-.n92 OUT-.n68 0.146911
R602 OUT-.n93 OUT-.n45 0.146911
R603 OUT-.n94 OUT-.n22 0.146911
R604 OUT- OUT-.n96 0.00392857
R605 VSS.n430 VSS.n427 4305.43
R606 VSS.t26 VSS.n20 2298.26
R607 VSS.t34 VSS.n413 2273.61
R608 VSS.n12 VSS.t16 2129.07
R609 VSS.t57 VSS.n12 2122.02
R610 VSS.n420 VSS.t54 2106.22
R611 VSS.t83 VSS.n420 2102.28
R612 VSS.n10 VSS.n9 2074.41
R613 VSS.n412 VSS.n10 1813.46
R614 VSS.n412 VSS.t114 1424.08
R615 VSS.t64 VSS.n13 1424.08
R616 VSS.t51 VSS.n421 1411.83
R617 VSS.t49 VSS.n412 1408.8
R618 VSS.t114 VSS.n21 599.241
R619 VSS.n11 VSS.t15 599.241
R620 VSS.n14 VSS.t57 599.241
R621 VSS.n422 VSS.t83 594.087
R622 VSS.n414 VSS.t49 592.812
R623 VSS.n419 VSS.t50 592.812
R624 VSS.n21 VSS.t26 528.742
R625 VSS.t16 VSS.n11 528.742
R626 VSS.n14 VSS.t64 528.742
R627 VSS.n422 VSS.t51 524.194
R628 VSS.n414 VSS.t34 523.069
R629 VSS.t54 VSS.n419 523.069
R630 VSS.n4 VSS.t36 239.559
R631 VSS.n377 VSS.t113 135.75
R632 VSS.n7 VSS.t66 119.779
R633 VSS.n30 VSS.t72 105.406
R634 VSS.t72 VSS.n29 102.212
R635 VSS.t48 VSS.t0 99.0177
R636 VSS.n369 VSS.t13 91.0324
R637 VSS.t113 VSS.t102 91.0324
R638 VSS.n388 VSS.t25 86.2413
R639 VSS.n431 VSS.t37 67.0767
R640 VSS.n395 VSS.t90 60.6885
R641 VSS.n3 VSS.n0 55.8973
R642 VSS.n202 VSS.t32 48.8215
R643 VSS.n93 VSS.t78 43.1446
R644 VSS.n401 VSS.t43 41.5238
R645 VSS.n358 VSS.t97 40.8739
R646 VSS.n350 VSS.t18 36.3324
R647 VSS.n412 VSS.t81 36.3324
R648 VSS.n346 VSS.t24 34.0616
R649 VSS.n337 VSS.t62 29.5201
R650 VSS.t13 VSS.t46 28.7474
R651 VSS.n331 VSS.t14 27.2494
R652 VSS.n405 VSS.t48 25.5533
R653 VSS.n0 VSS.t40 23.9563
R654 VSS.n322 VSS.t12 22.7079
R655 VSS.t90 VSS.t38 20.7622
R656 VSS.n317 VSS.t53 20.4372
R657 VSS.n307 VSS.t108 15.8957
R658 VSS.n238 VSS.t9 14.7603
R659 VSS.n301 VSS.t91 13.625
R660 VSS.n295 VSS.t3 11.3542
R661 VSS.n373 VSS.n31 11.2304
R662 VSS.n393 VSS.n31 11.2304
R663 VSS.t74 VSS.t28 9.08347
R664 VSS.t105 VSS.t29 9.08347
R665 VSS.t23 VSS.t22 9.08347
R666 VSS.t68 VSS.t8 9.08347
R667 VSS.n290 VSS.t63 9.08347
R668 VSS.t63 VSS.t19 9.08347
R669 VSS.t91 VSS.t10 9.08347
R670 VSS.t108 VSS.t11 9.08347
R671 VSS.t21 VSS.t99 9.08347
R672 VSS.t53 VSS.t20 9.08347
R673 VSS.t12 VSS.t33 9.08347
R674 VSS.t6 VSS.t71 9.08347
R675 VSS.t14 VSS.t7 9.08347
R676 VSS.t62 VSS.t30 9.08347
R677 VSS.n229 VSS.t21 7.9481
R678 VSS.t81 VSS.n411 7.9481
R679 VSS.n284 VSS.t68 6.81273
R680 VSS.n18 VSS.t27 6.65541
R681 VSS.n16 VSS.t17 6.65541
R682 VSS.n8 VSS.t65 6.65541
R683 VSS.n416 VSS.t35 6.65541
R684 VSS.n417 VSS.t55 6.65541
R685 VSS.n424 VSS.t52 6.65541
R686 VSS.n371 VSS.t47 6.65541
R687 VSS.n391 VSS.t39 6.65541
R688 VSS.n434 VSS.t67 6.65541
R689 VSS.n406 VSS.n405 6.38871
R690 VSS.n395 VSS.n394 6.38871
R691 VSS.n388 VSS.n387 6.38871
R692 VSS.n4 VSS.n3 6.38871
R693 VSS.t40 VSS.t59 6.38871
R694 VSS.n431 VSS.n430 6.38871
R695 VSS.n260 VSS.n259 6.21452
R696 VSS.n423 VSS.n422 5.2005
R697 VSS.n415 VSS.n414 5.2005
R698 VSS.n419 VSS.n418 5.2005
R699 VSS.n21 VSS.n19 5.2005
R700 VSS.n17 VSS.n11 5.2005
R701 VSS.n15 VSS.n14 5.2005
R702 VSS.n370 VSS.n369 5.2005
R703 VSS.n378 VSS.n377 5.2005
R704 VSS.n435 VSS.n7 5.2005
R705 VSS.n428 VSS.t112 5.13332
R706 VSS.n259 VSS.n182 5.10637
R707 VSS.n278 VSS.t23 4.54198
R708 VSS.n425 VSS.n8 3.81335
R709 VSS.n353 VSS.n98 3.78833
R710 VSS.n334 VSS.n100 3.78833
R711 VSS.n315 VSS.n102 3.78833
R712 VSS.n293 VSS.n104 3.78833
R713 VSS.n270 VSS.n106 3.78833
R714 VSS.n366 VSS.n35 3.78833
R715 VSS.n376 VSS.n33 3.78833
R716 VSS.n381 VSS.n380 3.78833
R717 VSS.n246 VSS.n184 3.74137
R718 VSS.n237 VSS.n186 3.74137
R719 VSS.n222 VSS.n188 3.74137
R720 VSS.n206 VSS.n190 3.74137
R721 VSS.n26 VSS.n25 3.74137
R722 VSS.n404 VSS.n28 3.74137
R723 VSS.n384 VSS.n383 3.74137
R724 VSS.n426 VSS.n425 3.52971
R725 VSS.n208 VSS.t111 3.40661
R726 VSS.n209 VSS.t31 3.40661
R727 VSS.n150 VSS.n149 2.64635
R728 VSS.n153 VSS.n152 2.64635
R729 VSS.n156 VSS.n155 2.64635
R730 VSS.n181 VSS.n109 2.60322
R731 VSS.n408 VSS.n407 2.6005
R732 VSS.n407 VSS.n406 2.6005
R733 VSS.n403 VSS.n402 2.6005
R734 VSS.n402 VSS.n401 2.6005
R735 VSS.n400 VSS.n399 2.6005
R736 VSS.n399 VSS.n398 2.6005
R737 VSS.n397 VSS.n396 2.6005
R738 VSS.n396 VSS.n395 2.6005
R739 VSS.n386 VSS.n385 2.6005
R740 VSS.n387 VSS.n386 2.6005
R741 VSS.n2 VSS.n1 2.6005
R742 VSS.n3 VSS.n2 2.6005
R743 VSS.n429 VSS.n428 2.6005
R744 VSS.n430 VSS.n429 2.6005
R745 VSS.n258 VSS.n257 2.6005
R746 VSS.n257 VSS.n256 2.6005
R747 VSS.n254 VSS.n253 2.6005
R748 VSS.n253 VSS.n252 2.6005
R749 VSS.n250 VSS.n249 2.6005
R750 VSS.n249 VSS.n248 2.6005
R751 VSS.n245 VSS.n244 2.6005
R752 VSS.n244 VSS.n243 2.6005
R753 VSS.n241 VSS.n240 2.6005
R754 VSS.n240 VSS.n239 2.6005
R755 VSS.n236 VSS.n235 2.6005
R756 VSS.n235 VSS.n234 2.6005
R757 VSS.n232 VSS.n231 2.6005
R758 VSS.n231 VSS.n230 2.6005
R759 VSS.n227 VSS.n226 2.6005
R760 VSS.n226 VSS.n225 2.6005
R761 VSS.n221 VSS.n220 2.6005
R762 VSS.n220 VSS.n219 2.6005
R763 VSS.n216 VSS.n215 2.6005
R764 VSS.n215 VSS.n214 2.6005
R765 VSS.n211 VSS.n210 2.6005
R766 VSS.n210 VSS.n209 2.6005
R767 VSS.n205 VSS.n204 2.6005
R768 VSS.n204 VSS.n203 2.6005
R769 VSS.n200 VSS.n199 2.6005
R770 VSS.n199 VSS.n198 2.6005
R771 VSS.n195 VSS.n194 2.6005
R772 VSS.n194 VSS.n193 2.6005
R773 VSS.n410 VSS.n409 2.6005
R774 VSS.n411 VSS.n410 2.6005
R775 VSS.n96 VSS.n95 2.6005
R776 VSS.n56 VSS.n55 2.6005
R777 VSS.n58 VSS.n57 2.6005
R778 VSS.n60 VSS.n59 2.6005
R779 VSS.n62 VSS.n61 2.6005
R780 VSS.n64 VSS.n63 2.6005
R781 VSS.n66 VSS.n65 2.6005
R782 VSS.n68 VSS.n67 2.6005
R783 VSS.n70 VSS.n69 2.6005
R784 VSS.n72 VSS.n71 2.6005
R785 VSS.n74 VSS.n73 2.6005
R786 VSS.n76 VSS.n75 2.6005
R787 VSS.n78 VSS.n77 2.6005
R788 VSS.n80 VSS.n79 2.6005
R789 VSS.n83 VSS.n82 2.6005
R790 VSS.n85 VSS.n84 2.6005
R791 VSS.n54 VSS.n53 2.6005
R792 VSS.n52 VSS.n51 2.6005
R793 VSS.n120 VSS.n119 2.6005
R794 VSS.n108 VSS.n107 2.6005
R795 VSS.n262 VSS.n261 2.6005
R796 VSS.t74 VSS.n267 2.6005
R797 VSS.n274 VSS.n273 2.6005
R798 VSS.n278 VSS.n277 2.6005
R799 VSS.n284 VSS.n283 2.6005
R800 VSS.n290 VSS.n289 2.6005
R801 VSS.n295 VSS.n294 2.6005
R802 VSS.n301 VSS.n300 2.6005
R803 VSS.n307 VSS.n306 2.6005
R804 VSS.n311 VSS.n310 2.6005
R805 VSS.n317 VSS.n316 2.6005
R806 VSS.n322 VSS.n321 2.6005
R807 VSS.n326 VSS.n325 2.6005
R808 VSS.n331 VSS.n330 2.6005
R809 VSS.n337 VSS.n336 2.6005
R810 VSS.n341 VSS.n340 2.6005
R811 VSS.n346 VSS.n345 2.6005
R812 VSS.n46 VSS.n45 2.6005
R813 VSS.n48 VSS.n47 2.6005
R814 VSS.n50 VSS.n49 2.6005
R815 VSS.n124 VSS.n123 2.6005
R816 VSS.n174 VSS.n173 2.6005
R817 VSS.n157 VSS.n156 2.6005
R818 VSS.n154 VSS.n153 2.6005
R819 VSS.n151 VSS.n150 2.6005
R820 VSS.n148 VSS.n147 2.6005
R821 VSS.n146 VSS.n145 2.6005
R822 VSS.n144 VSS.n143 2.6005
R823 VSS.n142 VSS.n141 2.6005
R824 VSS.n140 VSS.n139 2.6005
R825 VSS.n138 VSS.n137 2.6005
R826 VSS.n136 VSS.n135 2.6005
R827 VSS.n134 VSS.n133 2.6005
R828 VSS.n132 VSS.n131 2.6005
R829 VSS.n130 VSS.n129 2.6005
R830 VSS.n128 VSS.n127 2.6005
R831 VSS.n126 VSS.n125 2.6005
R832 VSS.n122 VSS.n121 2.6005
R833 VSS.n177 VSS.n176 2.6005
R834 VSS.n180 VSS.n179 2.6005
R835 VSS.n179 VSS.n178 2.6005
R836 VSS.n364 VSS.n363 2.6005
R837 VSS.n360 VSS.n359 2.6005
R838 VSS.n359 VSS.n358 2.6005
R839 VSS.n356 VSS.n355 2.6005
R840 VSS.n355 VSS.n354 2.6005
R841 VSS.n352 VSS.n351 2.6005
R842 VSS.n351 VSS.n350 2.6005
R843 VSS.n348 VSS.n347 2.6005
R844 VSS.n347 VSS.n346 2.6005
R845 VSS.n343 VSS.n342 2.6005
R846 VSS.n342 VSS.n341 2.6005
R847 VSS.n339 VSS.n338 2.6005
R848 VSS.n338 VSS.n337 2.6005
R849 VSS.n333 VSS.n332 2.6005
R850 VSS.n332 VSS.n331 2.6005
R851 VSS.n328 VSS.n327 2.6005
R852 VSS.n327 VSS.n326 2.6005
R853 VSS.n324 VSS.n323 2.6005
R854 VSS.n323 VSS.n322 2.6005
R855 VSS.n319 VSS.n318 2.6005
R856 VSS.n318 VSS.n317 2.6005
R857 VSS.n313 VSS.n312 2.6005
R858 VSS.n312 VSS.n311 2.6005
R859 VSS.n309 VSS.n308 2.6005
R860 VSS.n308 VSS.n307 2.6005
R861 VSS.n303 VSS.n302 2.6005
R862 VSS.n302 VSS.n301 2.6005
R863 VSS.n297 VSS.n296 2.6005
R864 VSS.n296 VSS.n295 2.6005
R865 VSS.n292 VSS.n291 2.6005
R866 VSS.n291 VSS.n290 2.6005
R867 VSS.n286 VSS.n285 2.6005
R868 VSS.n285 VSS.n284 2.6005
R869 VSS.n280 VSS.n279 2.6005
R870 VSS.n279 VSS.n278 2.6005
R871 VSS.n276 VSS.n275 2.6005
R872 VSS.n275 VSS.n274 2.6005
R873 VSS.n269 VSS.n268 2.6005
R874 VSS.n268 VSS.t74 2.6005
R875 VSS.n264 VSS.n263 2.6005
R876 VSS.n263 VSS.n262 2.6005
R877 VSS.n109 VSS.n108 2.6005
R878 VSS.n192 VSS.n191 2.6005
R879 VSS.n272 VSS.n271 2.6005
R880 VSS.n282 VSS.n281 2.6005
R881 VSS.n288 VSS.n287 2.6005
R882 VSS.n299 VSS.n298 2.6005
R883 VSS.n305 VSS.n304 2.6005
R884 VSS.n229 VSS.n228 2.6005
R885 VSS.n224 VSS.n223 2.6005
R886 VSS.n218 VSS.n217 2.6005
R887 VSS.n213 VSS.n212 2.6005
R888 VSS.n208 VSS.n207 2.6005
R889 VSS.n202 VSS.n201 2.6005
R890 VSS.n197 VSS.n196 2.6005
R891 VSS.n266 VSS.n265 2.6005
R892 VSS.n23 VSS.n22 2.6005
R893 VSS.n368 VSS.n367 2.6005
R894 VSS.n374 VSS.n373 2.6005
R895 VSS.n373 VSS.n372 2.6005
R896 VSS.n375 VSS.n31 2.6005
R897 VSS.n31 VSS.n30 2.6005
R898 VSS.n393 VSS.n392 2.6005
R899 VSS.n394 VSS.n393 2.6005
R900 VSS.n390 VSS.n389 2.6005
R901 VSS.n389 VSS.n388 2.6005
R902 VSS.n6 VSS.n5 2.6005
R903 VSS.n5 VSS.n4 2.6005
R904 VSS.n433 VSS.n432 2.6005
R905 VSS.n432 VSS.n431 2.6005
R906 VSS.n425 VSS.n424 2.53474
R907 VSS.n262 VSS.t56 2.27124
R908 VSS.n256 VSS.n255 2.27124
R909 VSS.n252 VSS.n251 2.27124
R910 VSS.n274 VSS.t105 2.27124
R911 VSS.n248 VSS.n247 2.27124
R912 VSS.n243 VSS.n242 2.27124
R913 VSS.n239 VSS.n238 2.27124
R914 VSS.n234 VSS.n233 2.27124
R915 VSS.n230 VSS.n229 2.27124
R916 VSS.n225 VSS.n224 2.27124
R917 VSS.n219 VSS.n218 2.27124
R918 VSS.n214 VSS.n213 2.27124
R919 VSS.n209 VSS.n208 2.27124
R920 VSS.n203 VSS.n202 2.27124
R921 VSS.n198 VSS.n197 2.27124
R922 VSS.n193 VSS.n192 2.27124
R923 VSS.n411 VSS.n23 2.27124
R924 VSS.n95 VSS.n94 1.75437
R925 VSS.n82 VSS.n81 1.75437
R926 VSS.n173 VSS.n172 1.50887
R927 VSS.n184 VSS.t118 1.3655
R928 VSS.n184 VSS.n183 1.3655
R929 VSS.n186 VSS.t101 1.3655
R930 VSS.n186 VSS.n185 1.3655
R931 VSS.n188 VSS.t85 1.3655
R932 VSS.n188 VSS.n187 1.3655
R933 VSS.n190 VSS.t119 1.3655
R934 VSS.n190 VSS.n189 1.3655
R935 VSS.n25 VSS.t98 1.3655
R936 VSS.n25 VSS.n24 1.3655
R937 VSS.n28 VSS.t89 1.3655
R938 VSS.n28 VSS.n27 1.3655
R939 VSS.n383 VSS.t120 1.3655
R940 VSS.n383 VSS.n382 1.3655
R941 VSS.n98 VSS.t58 1.3655
R942 VSS.n98 VSS.n97 1.3655
R943 VSS.n100 VSS.t84 1.3655
R944 VSS.n100 VSS.n99 1.3655
R945 VSS.n102 VSS.t100 1.3655
R946 VSS.n102 VSS.n101 1.3655
R947 VSS.n104 VSS.t117 1.3655
R948 VSS.n104 VSS.n103 1.3655
R949 VSS.n106 VSS.t75 1.3655
R950 VSS.n106 VSS.n105 1.3655
R951 VSS.n35 VSS.t82 1.3655
R952 VSS.n35 VSS.n34 1.3655
R953 VSS.n33 VSS.t73 1.3655
R954 VSS.n33 VSS.n32 1.3655
R955 VSS.n380 VSS.t88 1.3655
R956 VSS.n380 VSS.n379 1.3655
R957 VSS.n171 VSS.n158 1.27833
R958 VSS.n171 VSS.n159 1.27833
R959 VSS.n171 VSS.n160 1.27833
R960 VSS.n171 VSS.n161 1.27833
R961 VSS.n171 VSS.n162 1.27833
R962 VSS.n171 VSS.n163 1.27833
R963 VSS.n171 VSS.n164 1.27833
R964 VSS.n171 VSS.n165 1.27833
R965 VSS.n171 VSS.n166 1.27833
R966 VSS.n171 VSS.n167 1.27833
R967 VSS.n171 VSS.n168 1.27833
R968 VSS.n171 VSS.n169 1.27833
R969 VSS.n181 VSS.n180 1.2289
R970 VSS.n218 VSS.t6 1.13587
R971 VSS.n198 VSS.t92 1.13587
R972 VSS.n171 VSS.n170 0.729291
R973 VSS.n172 VSS.n171 0.729086
R974 VSS.n18 VSS 0.684889
R975 VSS VSS.n416 0.684889
R976 VSS.n16 VSS 0.620412
R977 VSS.n417 VSS 0.620412
R978 VSS.n94 VSS.n93 0.424314
R979 VSS.n93 VSS.n92 0.424314
R980 VSS.n93 VSS.n91 0.424314
R981 VSS.n93 VSS.n90 0.424314
R982 VSS.n93 VSS.n89 0.424314
R983 VSS.n93 VSS.n88 0.424314
R984 VSS.n93 VSS.n87 0.424314
R985 VSS.n93 VSS.n86 0.424314
R986 VSS.n426 VSS 0.341269
R987 VSS.n174 VSS.n157 0.240099
R988 VSS.n157 VSS.n154 0.240099
R989 VSS.n154 VSS.n151 0.240099
R990 VSS.n151 VSS.n148 0.240099
R991 VSS.n148 VSS.n146 0.240099
R992 VSS.n146 VSS.n144 0.240099
R993 VSS.n144 VSS.n142 0.240099
R994 VSS.n142 VSS.n140 0.240099
R995 VSS.n140 VSS.n138 0.240099
R996 VSS.n138 VSS.n136 0.240099
R997 VSS.n136 VSS.n134 0.240099
R998 VSS.n134 VSS.n132 0.240099
R999 VSS.n132 VSS.n130 0.240099
R1000 VSS.n130 VSS.n128 0.240099
R1001 VSS.n128 VSS.n126 0.240099
R1002 VSS.n126 VSS.n124 0.240099
R1003 VSS.n56 VSS.n54 0.240099
R1004 VSS.n58 VSS.n56 0.240099
R1005 VSS.n60 VSS.n58 0.240099
R1006 VSS.n62 VSS.n60 0.240099
R1007 VSS.n64 VSS.n62 0.240099
R1008 VSS.n66 VSS.n64 0.240099
R1009 VSS.n68 VSS.n66 0.240099
R1010 VSS.n70 VSS.n68 0.240099
R1011 VSS.n72 VSS.n70 0.240099
R1012 VSS.n74 VSS.n72 0.240099
R1013 VSS.n76 VSS.n74 0.240099
R1014 VSS.n78 VSS.n76 0.240099
R1015 VSS.n80 VSS.n78 0.240099
R1016 VSS.n83 VSS.n80 0.240099
R1017 VSS.n85 VSS.n83 0.240099
R1018 VSS.n96 VSS.n85 0.240099
R1019 VSS.n122 VSS.n120 0.234957
R1020 VSS.n120 VSS.n118 0.234957
R1021 VSS.n118 VSS.n117 0.234957
R1022 VSS.n117 VSS.n116 0.234957
R1023 VSS.n116 VSS.n115 0.234957
R1024 VSS.n115 VSS.n114 0.234957
R1025 VSS.n114 VSS.n113 0.234957
R1026 VSS.n113 VSS.n112 0.234957
R1027 VSS.n112 VSS.n111 0.234957
R1028 VSS.n111 VSS.n110 0.234957
R1029 VSS.n37 VSS.n36 0.234957
R1030 VSS.n38 VSS.n37 0.234957
R1031 VSS.n39 VSS.n38 0.234957
R1032 VSS.n40 VSS.n39 0.234957
R1033 VSS.n41 VSS.n40 0.234957
R1034 VSS.n42 VSS.n41 0.234957
R1035 VSS.n43 VSS.n42 0.234957
R1036 VSS.n44 VSS.n43 0.234957
R1037 VSS.n46 VSS.n44 0.234957
R1038 VSS.n48 VSS.n46 0.234957
R1039 VSS.n50 VSS.n48 0.234957
R1040 VSS.n52 VSS.n50 0.234957
R1041 VSS.n180 VSS.n177 0.234957
R1042 VSS.n364 VSS.n96 0.220714
R1043 VSS.n54 VSS.n52 0.209695
R1044 VSS.n124 VSS.n122 0.199945
R1045 VSS.n177 VSS.n174 0.197176
R1046 VSS.n433 VSS.n426 0.159446
R1047 VSS.n258 VSS.n254 0.144885
R1048 VSS.n254 VSS.n250 0.144885
R1049 VSS.n245 VSS.n241 0.144885
R1050 VSS.n236 VSS.n232 0.144885
R1051 VSS.n232 VSS.n227 0.144885
R1052 VSS.n221 VSS.n216 0.144885
R1053 VSS.n216 VSS.n211 0.144885
R1054 VSS.n205 VSS.n200 0.144885
R1055 VSS.n200 VSS.n195 0.144885
R1056 VSS.n409 VSS.n408 0.144885
R1057 VSS.n403 VSS.n400 0.144885
R1058 VSS.n400 VSS.n397 0.144885
R1059 VSS.n19 VSS.n18 0.142847
R1060 VSS.n15 VSS.n8 0.142847
R1061 VSS.n416 VSS.n415 0.142847
R1062 VSS.n418 VSS.n417 0.142847
R1063 VSS.n424 VSS.n423 0.142847
R1064 VSS.n409 VSS.n26 0.141035
R1065 VSS VSS.n16 0.130908
R1066 VSS.n241 VSS.n237 0.125634
R1067 VSS.n246 VSS.n245 0.123709
R1068 VSS.n408 VSS.n404 0.108307
R1069 VSS.n363 VSS.n362 0.108192
R1070 VSS.n176 VSS.n175 0.108192
R1071 VSS.n206 VSS.n205 0.100607
R1072 VSS.n227 VSS.n222 0.0852059
R1073 VSS.n259 VSS.n258 0.0832807
R1074 VSS.n385 VSS.n384 0.0775053
R1075 VSS.n222 VSS.n221 0.0601791
R1076 VSS.n365 VSS.n364 0.055041
R1077 VSS.n390 VSS.n381 0.0549122
R1078 VSS VSS.n376 0.0523246
R1079 VSS.n211 VSS.n206 0.0447781
R1080 VSS.n280 VSS.n276 0.0390439
R1081 VSS.n313 VSS.n309 0.0390439
R1082 VSS.n328 VSS.n324 0.0390439
R1083 VSS.n343 VSS.n339 0.0390439
R1084 VSS.n368 VSS.n366 0.0388886
R1085 VSS.n404 VSS.n403 0.0370775
R1086 VSS.n391 VSS.n390 0.035798
R1087 VSS.n375 VSS 0.0353367
R1088 VSS.n371 VSS.n370 0.0335569
R1089 VSS.n435 VSS.n434 0.0334787
R1090 VSS.n353 VSS.n352 0.0324914
R1091 VSS.n288 VSS.n286 0.0317206
R1092 VSS.n305 VSS.n303 0.0317206
R1093 VSS.n320 VSS.n319 0.0317206
R1094 VSS.n349 VSS.n348 0.0317206
R1095 VSS.n361 VSS.n360 0.0317206
R1096 VSS VSS.n374 0.0307574
R1097 VSS VSS.n6 0.0307128
R1098 VSS.n334 VSS.n333 0.0294079
R1099 VSS.n392 VSS.n391 0.0292915
R1100 VSS.n269 VSS.n266 0.0270953
R1101 VSS.n286 VSS.n282 0.0270953
R1102 VSS.n303 VSS.n299 0.0270953
R1103 VSS.n333 VSS.n329 0.0270953
R1104 VSS.n348 VSS.n344 0.0270953
R1105 VSS.n360 VSS.n357 0.0270953
R1106 VSS.n366 VSS.n365 0.0260924
R1107 VSS.n264 VSS.n260 0.0253608
R1108 VSS.n293 VSS.n292 0.0232409
R1109 VSS.n250 VSS.n246 0.0216765
R1110 VSS.n270 VSS.n269 0.0201574
R1111 VSS.n237 VSS.n236 0.0197513
R1112 VSS.n374 VSS.n371 0.0167085
R1113 VSS.n297 VSS.n293 0.016303
R1114 VSS VSS.n368 0.0150024
R1115 VSS.n315 VSS.n314 0.0143758
R1116 VSS.n319 VSS.n315 0.0132195
R1117 VSS.n260 VSS.n181 0.0124649
R1118 VSS.n266 VSS.n264 0.0124486
R1119 VSS.n282 VSS.n280 0.0124486
R1120 VSS.n299 VSS.n297 0.0124486
R1121 VSS.n314 VSS.n313 0.0124486
R1122 VSS.n329 VSS.n328 0.0124486
R1123 VSS.n344 VSS.n343 0.0124486
R1124 VSS.n357 VSS.n356 0.0124486
R1125 VSS.n17 VSS 0.0124388
R1126 VSS.n272 VSS.n270 0.0120632
R1127 VSS.n381 VSS.n6 0.0107128
R1128 VSS.n376 VSS.n375 0.00817773
R1129 VSS.n276 VSS.n272 0.00782334
R1130 VSS.n292 VSS.n288 0.00782334
R1131 VSS.n309 VSS.n305 0.00782334
R1132 VSS.n324 VSS.n320 0.00782334
R1133 VSS.n339 VSS.n335 0.00782334
R1134 VSS.n352 VSS.n349 0.00782334
R1135 VSS.n364 VSS.n361 0.00782334
R1136 VSS.n356 VSS.n353 0.00705246
R1137 VSS.n392 VSS.n378 0.0047654
R1138 VSS.n195 VSS.n26 0.00435027
R1139 VSS.n335 VSS.n334 0.00281263
R1140 VSS.n19 VSS 0.00141837
R1141 VSS VSS.n17 0.00141837
R1142 VSS VSS.n15 0.00141837
R1143 VSS.n415 VSS 0.00141837
R1144 VSS.n418 VSS 0.00141837
R1145 VSS.n423 VSS 0.00141837
R1146 VSS.n434 VSS.n433 0.000925532
R1147 VSS.n370 VSS 0.00071327
R1148 VSS.n378 VSS 0.00071327
R1149 VSS VSS.n435 0.000712766
R1150 IM_T.n18 IM_T.t25 84.5899
R1151 IM_T.n20 IM_T.n19 64.4419
R1152 IM_T.n22 IM_T.n21 64.4419
R1153 IM_T.n24 IM_T.n23 64.4419
R1154 IM_T.n26 IM_T.n25 64.4419
R1155 IM_T.n28 IM_T.n27 64.4419
R1156 IM_T.n30 IM_T.n29 64.4419
R1157 IM_T.n32 IM_T.n31 64.4419
R1158 IM_T.n3 IM_T.n2 63.3497
R1159 IM_T.n5 IM_T.n4 63.3497
R1160 IM_T.n7 IM_T.n6 63.3497
R1161 IM_T.n9 IM_T.n8 63.3497
R1162 IM_T.n11 IM_T.n10 63.3497
R1163 IM_T.n13 IM_T.n12 63.3497
R1164 IM_T.n15 IM_T.n14 63.3497
R1165 IM_T.n17 IM_T.n16 57.704
R1166 IM_T.n2 IM_T.t27 31.3373
R1167 IM_T.n33 IM_T.n32 31.1676
R1168 IM_T.n18 IM_T.t21 20.1485
R1169 IM_T.n19 IM_T.t8 20.1485
R1170 IM_T.n20 IM_T.t9 20.1485
R1171 IM_T.n21 IM_T.t12 20.1485
R1172 IM_T.n22 IM_T.t20 20.1485
R1173 IM_T.n23 IM_T.t28 20.1485
R1174 IM_T.n24 IM_T.t7 20.1485
R1175 IM_T.n25 IM_T.t22 20.1485
R1176 IM_T.n26 IM_T.t13 20.1485
R1177 IM_T.n27 IM_T.t5 20.1485
R1178 IM_T.n28 IM_T.t29 20.1485
R1179 IM_T.n29 IM_T.t14 20.1485
R1180 IM_T.n30 IM_T.t6 20.1485
R1181 IM_T.n31 IM_T.t31 20.1485
R1182 IM_T.n32 IM_T.t23 20.1485
R1183 IM_T.n2 IM_T.t4 18.4695
R1184 IM_T.n3 IM_T.t2 18.4695
R1185 IM_T.n4 IM_T.t19 18.4695
R1186 IM_T.n5 IM_T.t15 18.4695
R1187 IM_T.n6 IM_T.t24 18.4695
R1188 IM_T.n7 IM_T.t1 18.4695
R1189 IM_T.n8 IM_T.t17 18.4695
R1190 IM_T.n9 IM_T.t18 18.4695
R1191 IM_T.n10 IM_T.t11 18.4695
R1192 IM_T.n11 IM_T.t10 18.4695
R1193 IM_T.n12 IM_T.t30 18.4695
R1194 IM_T.n13 IM_T.t16 18.4695
R1195 IM_T.n14 IM_T.t0 18.4695
R1196 IM_T.n15 IM_T.t3 18.4695
R1197 IM_T.n16 IM_T.t26 18.4695
R1198 IM_T.n19 IM_T.n18 13.0902
R1199 IM_T.n21 IM_T.n20 13.0902
R1200 IM_T.n23 IM_T.n22 13.0902
R1201 IM_T.n25 IM_T.n24 13.0902
R1202 IM_T.n27 IM_T.n26 13.0902
R1203 IM_T.n29 IM_T.n28 13.0902
R1204 IM_T.n31 IM_T.n30 13.0902
R1205 IM_T.n4 IM_T.n3 12.8683
R1206 IM_T.n6 IM_T.n5 12.8683
R1207 IM_T.n8 IM_T.n7 12.8683
R1208 IM_T.n10 IM_T.n9 12.8683
R1209 IM_T.n12 IM_T.n11 12.8683
R1210 IM_T.n14 IM_T.n13 12.8683
R1211 IM_T.n16 IM_T.n15 12.8683
R1212 IM_T.n34 IM_T.n33 2.25726
R1213 IM_T.n34 IM_T.n1 2.24397
R1214 IM_T.n1 IM_T 0.530288
R1215 IM_T.n34 IM_T.n17 0.0277093
R1216 IM_T.n1 IM_T.n0 0.0150524
R1217 IM_T IM_T.n34 0.00154651
R1218 SD.n81 SD.n78 4.5005
R1219 SD.n82 SD.n81 4.5005
R1220 SD.n68 SD.n13 3.63741
R1221 SD.n42 SD.n41 3.28149
R1222 SD.n53 SD.n27 3.28101
R1223 SD.n65 SD.n18 3.27542
R1224 SD.n2 SD.n1 3.26817
R1225 SD.n106 SD.n88 3.258
R1226 SD.n44 SD.n34 3.25644
R1227 SD.n77 SD.n4 3.24511
R1228 SD.n95 SD.n92 3.23798
R1229 SD.n97 SD.n90 3.23061
R1230 SD.n74 SD.n11 3.2111
R1231 SD.n59 SD.n20 3.20644
R1232 SD.n56 SD.n22 3.20496
R1233 SD.n50 SD.n32 3.204
R1234 SD.n108 SD.n86 3.19428
R1235 SD.n113 SD.n84 3.16815
R1236 SD.n111 SD.n110 2.58749
R1237 SD.n76 SD.n6 2.5852
R1238 SD.n42 SD.n39 2.57457
R1239 SD.n95 SD.n94 2.56564
R1240 SD.n49 SD.n48 2.24976
R1241 SD.n63 SD.n62 2.24638
R1242 SD.n101 SD.n100 2.24631
R1243 SD.n72 SD.n71 2.24557
R1244 SD.n117 SD.n116 2.24508
R1245 SD.n55 SD.n25 1.49577
R1246 SD.n105 SD.n104 1.49553
R1247 SD.n75 SD.n9 1.49548
R1248 SD.n43 SD.n37 1.49542
R1249 SD.n66 SD.n16 1.49542
R1250 SD.n52 SD.n30 1.49542
R1251 SD.n110 SD.t3 1.47093
R1252 SD.n27 SD.t1 1.47081
R1253 SD.n1 SD.t43 1.4708
R1254 SD.n18 SD.t20 1.46022
R1255 SD.n6 SD.t37 1.4602
R1256 SD.n88 SD.t54 1.46017
R1257 SD.n34 SD.t55 1.46008
R1258 SD.n70 SD.n69 1.45967
R1259 SD.n47 SD.n46 1.45927
R1260 SD.n4 SD.n3 1.45919
R1261 SD.n61 SD.n60 1.45916
R1262 SD.n116 SD.n115 1.4476
R1263 SD.n80 SD.n79 1.44746
R1264 SD.n104 SD.n103 1.44722
R1265 SD.n16 SD.n15 1.44631
R1266 SD.n37 SD.n36 1.4456
R1267 SD.n30 SD.n29 1.44501
R1268 SD.n9 SD.n8 1.44371
R1269 SD.n25 SD.n24 1.44299
R1270 SD.n99 SD.t5 1.42418
R1271 SD.n41 SD.n40 1.41105
R1272 SD.n115 SD.t18 1.3655
R1273 SD.n115 SD.n114 1.3655
R1274 SD.n103 SD.t48 1.3655
R1275 SD.n103 SD.n102 1.3655
R1276 SD.n94 SD.t22 1.3655
R1277 SD.n94 SD.n93 1.3655
R1278 SD.n92 SD.t2 1.3655
R1279 SD.n92 SD.n91 1.3655
R1280 SD.n90 SD.t17 1.3655
R1281 SD.n90 SD.n89 1.3655
R1282 SD.n86 SD.t34 1.3655
R1283 SD.n86 SD.n85 1.3655
R1284 SD.n84 SD.t0 1.3655
R1285 SD.n84 SD.n83 1.3655
R1286 SD.n8 SD.t50 1.3655
R1287 SD.n8 SD.n7 1.3655
R1288 SD.n15 SD.t63 1.3655
R1289 SD.n15 SD.n14 1.3655
R1290 SD.n24 SD.t56 1.3655
R1291 SD.n24 SD.n23 1.3655
R1292 SD.n29 SD.t29 1.3655
R1293 SD.n29 SD.n28 1.3655
R1294 SD.n36 SD.t44 1.3655
R1295 SD.n36 SD.n35 1.3655
R1296 SD.n39 SD.t14 1.3655
R1297 SD.n39 SD.n38 1.3655
R1298 SD.n32 SD.t40 1.3655
R1299 SD.n32 SD.n31 1.3655
R1300 SD.n22 SD.t36 1.3655
R1301 SD.n22 SD.n21 1.3655
R1302 SD.n20 SD.t58 1.3655
R1303 SD.n20 SD.n19 1.3655
R1304 SD.n13 SD.t9 1.3655
R1305 SD.n13 SD.n12 1.3655
R1306 SD.n11 SD.t26 1.3655
R1307 SD.n11 SD.n10 1.3655
R1308 SD.n41 SD.t23 1.28824
R1309 SD.n99 SD.n98 1.2738
R1310 SD.n80 SD.t10 1.24719
R1311 SD.n61 SD.t24 1.23341
R1312 SD.n4 SD.t49 1.23339
R1313 SD.n47 SD.t6 1.23331
R1314 SD.n70 SD.t31 1.23295
R1315 SD.n34 SD.n33 1.23247
R1316 SD.n88 SD.n87 1.23239
R1317 SD.n6 SD.n5 1.23236
R1318 SD.n18 SD.n17 1.23234
R1319 SD.n1 SD.n0 1.21851
R1320 SD.n27 SD.n26 1.21849
R1321 SD.n110 SD.n109 1.21839
R1322 SD.n71 SD.n70 1.09468
R1323 SD.n48 SD.n47 1.09004
R1324 SD.n81 SD.n80 1.08925
R1325 SD.n62 SD.n61 1.08871
R1326 SD.n100 SD.n99 1.08617
R1327 SD.n78 SD.n77 0.605393
R1328 SD.n96 SD.n95 0.603024
R1329 SD.n67 SD.n66 0.590381
R1330 SD.n49 SD.n45 0.57793
R1331 SD.n108 SD.n107 0.571801
R1332 SD.n43 SD.n42 0.571708
R1333 SD.n58 SD.n57 0.570677
R1334 SD.n76 SD.n75 0.57026
R1335 SD.n112 SD.n111 0.56537
R1336 SD.n55 SD.n54 0.560195
R1337 SD.n105 SD.n101 0.558901
R1338 SD.n52 SD.n51 0.553694
R1339 SD.n118 SD.n117 0.551536
R1340 SD.n73 SD.n72 0.54879
R1341 SD.n64 SD.n63 0.545974
R1342 SD.n74 SD.n73 0.0239783
R1343 SD.n65 SD.n64 0.0232473
R1344 SD.n54 SD.n53 0.0202802
R1345 SD.n107 SD.n106 0.0192912
R1346 SD.n45 SD.n44 0.0192912
R1347 SD.n57 SD.n56 0.0181289
R1348 SD.n44 SD.n43 0.0164699
R1349 SD.n101 SD.n97 0.0163101
R1350 SD SD.n118 0.0153352
R1351 SD.n106 SD.n105 0.0151457
R1352 SD.n56 SD.n55 0.0149378
R1353 SD.n53 SD.n52 0.0148219
R1354 SD.n113 SD.n112 0.0148149
R1355 SD.n51 SD.n50 0.0143462
R1356 SD.n72 SD.n68 0.0138309
R1357 SD.n77 SD.n76 0.0138281
R1358 SD.n117 SD.n113 0.0138259
R1359 SD.n111 SD.n108 0.0134986
R1360 SD.n63 SD.n59 0.0119156
R1361 SD.n66 SD.n65 0.0115197
R1362 SD.n50 SD.n49 0.0113833
R1363 SD.n75 SD.n74 0.011083
R1364 SD SD.n82 0.00643407
R1365 SD.n68 SD.n67 0.00445604
R1366 SD.n59 SD.n58 0.00386449
R1367 SD.n78 SD 0.00346703
R1368 SD.n97 SD.n96 0.00247802
R1369 SD.n82 SD.n2 0.00247802
R1370 SD SD.n2 0.00148901
R1371 Q.n56 Q.n55 74.7525
R1372 Q.n58 Q.n57 74.7525
R1373 Q.n60 Q.n59 74.7525
R1374 Q.n16 Q.t35 63.1408
R1375 Q.n62 Q.n61 60.196
R1376 Q.n22 Q.n21 50.8038
R1377 Q.n18 Q.n17 48.5408
R1378 Q.n20 Q.n19 48.5408
R1379 Q.n66 Q.t36 28.2228
R1380 Q.n55 Q.t16 28.1785
R1381 Q.n1 Q.t14 24.4602
R1382 Q.n39 Q.t54 24.4602
R1383 Q.n23 Q.t21 24.4602
R1384 Q.n57 Q.n56 15.1845
R1385 Q.n59 Q.n58 15.1845
R1386 Q.n61 Q.n60 15.1845
R1387 Q.n3 Q.t5 14.6005
R1388 Q.n4 Q.t43 14.6005
R1389 Q.n7 Q.t20 14.6005
R1390 Q.n8 Q.t55 14.6005
R1391 Q.n11 Q.t68 14.6005
R1392 Q.n12 Q.t23 14.6005
R1393 Q.n41 Q.t47 14.6005
R1394 Q.n42 Q.t13 14.6005
R1395 Q.n45 Q.t57 14.6005
R1396 Q.n46 Q.t25 14.6005
R1397 Q.n49 Q.t45 14.6005
R1398 Q.n50 Q.t60 14.6005
R1399 Q.n25 Q.t18 14.6005
R1400 Q.n26 Q.t53 14.6005
R1401 Q.n29 Q.t29 14.6005
R1402 Q.n30 Q.t63 14.6005
R1403 Q.n33 Q.t15 14.6005
R1404 Q.n34 Q.t33 14.6005
R1405 Q.n16 Q.t32 14.6005
R1406 Q.n17 Q.t65 14.6005
R1407 Q.n18 Q.t44 14.6005
R1408 Q.n19 Q.t7 14.6005
R1409 Q.n20 Q.t28 14.6005
R1410 Q.n21 Q.t48 14.6005
R1411 Q.n66 Q.t37 14.4701
R1412 Q.n1 Q.t31 14.0165
R1413 Q.n2 Q.t24 14.0165
R1414 Q.n5 Q.t42 14.0165
R1415 Q.n6 Q.t6 14.0165
R1416 Q.n9 Q.t67 14.0165
R1417 Q.n10 Q.t22 14.0165
R1418 Q.n13 Q.t39 14.0165
R1419 Q.n14 Q.t4 14.0165
R1420 Q.n39 Q.t66 14.0165
R1421 Q.n40 Q.t61 14.0165
R1422 Q.n43 Q.t12 14.0165
R1423 Q.n44 Q.t49 14.0165
R1424 Q.n47 Q.t41 14.0165
R1425 Q.n48 Q.t58 14.0165
R1426 Q.n51 Q.t9 14.0165
R1427 Q.n52 Q.t46 14.0165
R1428 Q.n23 Q.t38 14.0165
R1429 Q.n24 Q.t34 14.0165
R1430 Q.n27 Q.t52 14.0165
R1431 Q.n28 Q.t19 14.0165
R1432 Q.n31 Q.t11 14.0165
R1433 Q.n32 Q.t30 14.0165
R1434 Q.n35 Q.t50 14.0165
R1435 Q.n36 Q.t17 14.0165
R1436 Q.n55 Q.t8 12.9945
R1437 Q.n56 Q.t27 12.9945
R1438 Q.n57 Q.t62 12.9945
R1439 Q.n58 Q.t56 12.9945
R1440 Q.n59 Q.t3 12.9945
R1441 Q.n60 Q.t26 12.9945
R1442 Q.n61 Q.t59 12.9945
R1443 Q.n15 Q.t40 12.3375
R1444 Q.n53 Q.t10 12.3375
R1445 Q.n37 Q.t51 12.3375
R1446 Q.n22 Q.t64 12.3375
R1447 Q.n15 Q.n14 12.1232
R1448 Q.n53 Q.n52 12.1232
R1449 Q.n37 Q.n36 12.1232
R1450 Q.n2 Q.n1 9.86024
R1451 Q.n3 Q.n2 9.86024
R1452 Q.n4 Q.n3 9.86024
R1453 Q.n5 Q.n4 9.86024
R1454 Q.n6 Q.n5 9.86024
R1455 Q.n7 Q.n6 9.86024
R1456 Q.n8 Q.n7 9.86024
R1457 Q.n9 Q.n8 9.86024
R1458 Q.n10 Q.n9 9.86024
R1459 Q.n11 Q.n10 9.86024
R1460 Q.n12 Q.n11 9.86024
R1461 Q.n13 Q.n12 9.86024
R1462 Q.n14 Q.n13 9.86024
R1463 Q.n40 Q.n39 9.86024
R1464 Q.n41 Q.n40 9.86024
R1465 Q.n42 Q.n41 9.86024
R1466 Q.n43 Q.n42 9.86024
R1467 Q.n44 Q.n43 9.86024
R1468 Q.n45 Q.n44 9.86024
R1469 Q.n46 Q.n45 9.86024
R1470 Q.n47 Q.n46 9.86024
R1471 Q.n48 Q.n47 9.86024
R1472 Q.n49 Q.n48 9.86024
R1473 Q.n50 Q.n49 9.86024
R1474 Q.n51 Q.n50 9.86024
R1475 Q.n52 Q.n51 9.86024
R1476 Q.n24 Q.n23 9.86024
R1477 Q.n25 Q.n24 9.86024
R1478 Q.n26 Q.n25 9.86024
R1479 Q.n27 Q.n26 9.86024
R1480 Q.n28 Q.n27 9.86024
R1481 Q.n29 Q.n28 9.86024
R1482 Q.n30 Q.n29 9.86024
R1483 Q.n31 Q.n30 9.86024
R1484 Q.n32 Q.n31 9.86024
R1485 Q.n33 Q.n32 9.86024
R1486 Q.n34 Q.n33 9.86024
R1487 Q.n35 Q.n34 9.86024
R1488 Q.n36 Q.n35 9.86024
R1489 Q.n17 Q.n16 9.86024
R1490 Q.n19 Q.n18 9.86024
R1491 Q.n21 Q.n20 9.86024
R1492 Q.n38 Q.n22 9.72687
R1493 Q.n54 Q.n53 8.44029
R1494 Q.n38 Q.n37 8.44029
R1495 Q.n70 Q.n65 6.8765
R1496 Q.n63 Q.n15 6.14729
R1497 Q.n69 Q 6.04981
R1498 Q Q.n66 4.53357
R1499 Q.n68 Q.t1 3.6405
R1500 Q.n68 Q.n67 3.6405
R1501 Q Q.n63 3.63115
R1502 Q.n69 Q.n68 2.6005
R1503 Q.n64 Q 2.26759
R1504 Q.n63 Q.n62 2.2505
R1505 Q.n54 Q.n38 1.24534
R1506 Q.n62 Q.n54 1.24509
R1507 Q.n70 Q.n69 0.484465
R1508 Q Q.n70 0.17463
R1509 Q Q.n64 0.00252247
R1510 Q.n64 Q.n0 0.00151124
R1511 OUT+.n15 OUT+.t4 9.53443
R1512 OUT+.n84 OUT+.t28 9.53443
R1513 OUT+.n61 OUT+.t56 9.53443
R1514 OUT+.n38 OUT+.t17 9.53443
R1515 OUT+.n92 OUT+.n70 6.13289
R1516 OUT+.n46 OUT+.n24 6.13289
R1517 OUT+.n23 OUT+.n1 6.08789
R1518 OUT+.n69 OUT+.n47 6.08789
R1519 OUT+.n20 OUT+.n19 5.91472
R1520 OUT+.n89 OUT+.n88 5.91472
R1521 OUT+.n66 OUT+.n65 5.91472
R1522 OUT+.n43 OUT+.n42 5.91472
R1523 OUT+.n16 OUT+.n9 5.84965
R1524 OUT+.n85 OUT+.n78 5.84965
R1525 OUT+.n62 OUT+.n55 5.84965
R1526 OUT+.n39 OUT+.n32 5.84965
R1527 OUT+.n17 OUT+.n7 5.54055
R1528 OUT+.n86 OUT+.n76 5.54055
R1529 OUT+.n63 OUT+.n53 5.54055
R1530 OUT+.n40 OUT+.n30 5.54055
R1531 OUT+.n14 OUT+.n13 4.38877
R1532 OUT+.n83 OUT+.n82 4.38877
R1533 OUT+.n60 OUT+.n59 4.38877
R1534 OUT+.n37 OUT+.n36 4.38877
R1535 OUT+.n22 OUT+.n3 3.64354
R1536 OUT+.n91 OUT+.n72 3.64354
R1537 OUT+.n68 OUT+.n49 3.64354
R1538 OUT+.n45 OUT+.n26 3.64354
R1539 OUT+.n93 OUT+.n92 3.49643
R1540 OUT+.n21 OUT+.n5 3.29178
R1541 OUT+.n90 OUT+.n74 3.29178
R1542 OUT+.n67 OUT+.n51 3.29178
R1543 OUT+.n44 OUT+.n28 3.29178
R1544 OUT+.n14 OUT+.n11 3.29055
R1545 OUT+.n83 OUT+.n80 3.29055
R1546 OUT+.n60 OUT+.n57 3.29055
R1547 OUT+.n37 OUT+.n34 3.29055
R1548 OUT+.n21 OUT+.n20 3.08985
R1549 OUT+.n90 OUT+.n89 3.08985
R1550 OUT+.n67 OUT+.n66 3.08985
R1551 OUT+.n44 OUT+.n43 3.08985
R1552 OUT+.n95 OUT+.n23 2.87408
R1553 OUT+.n93 OUT+.n69 2.87254
R1554 OUT+.n94 OUT+.n46 2.83004
R1555 OUT+.n19 OUT+.t16 2.7305
R1556 OUT+.n19 OUT+.n18 2.7305
R1557 OUT+.n7 OUT+.t24 2.7305
R1558 OUT+.n7 OUT+.n6 2.7305
R1559 OUT+.n9 OUT+.t55 2.7305
R1560 OUT+.n9 OUT+.n8 2.7305
R1561 OUT+.n11 OUT+.t38 2.7305
R1562 OUT+.n11 OUT+.n10 2.7305
R1563 OUT+.n13 OUT+.t18 2.7305
R1564 OUT+.n13 OUT+.n12 2.7305
R1565 OUT+.n5 OUT+.t34 2.7305
R1566 OUT+.n5 OUT+.n4 2.7305
R1567 OUT+.n3 OUT+.t30 2.7305
R1568 OUT+.n3 OUT+.n2 2.7305
R1569 OUT+.n88 OUT+.t39 2.7305
R1570 OUT+.n88 OUT+.n87 2.7305
R1571 OUT+.n76 OUT+.t46 2.7305
R1572 OUT+.n76 OUT+.n75 2.7305
R1573 OUT+.n78 OUT+.t12 2.7305
R1574 OUT+.n78 OUT+.n77 2.7305
R1575 OUT+.n80 OUT+.t0 2.7305
R1576 OUT+.n80 OUT+.n79 2.7305
R1577 OUT+.n82 OUT+.t40 2.7305
R1578 OUT+.n82 OUT+.n81 2.7305
R1579 OUT+.n74 OUT+.t61 2.7305
R1580 OUT+.n74 OUT+.n73 2.7305
R1581 OUT+.n72 OUT+.t50 2.7305
R1582 OUT+.n72 OUT+.n71 2.7305
R1583 OUT+.n65 OUT+.t26 2.7305
R1584 OUT+.n65 OUT+.n64 2.7305
R1585 OUT+.n53 OUT+.t11 2.7305
R1586 OUT+.n53 OUT+.n52 2.7305
R1587 OUT+.n55 OUT+.t1 2.7305
R1588 OUT+.n55 OUT+.n54 2.7305
R1589 OUT+.n57 OUT+.t23 2.7305
R1590 OUT+.n57 OUT+.n56 2.7305
R1591 OUT+.n59 OUT+.t29 2.7305
R1592 OUT+.n59 OUT+.n58 2.7305
R1593 OUT+.n51 OUT+.t21 2.7305
R1594 OUT+.n51 OUT+.n50 2.7305
R1595 OUT+.n49 OUT+.t35 2.7305
R1596 OUT+.n49 OUT+.n48 2.7305
R1597 OUT+.n42 OUT+.t54 2.7305
R1598 OUT+.n42 OUT+.n41 2.7305
R1599 OUT+.n30 OUT+.t37 2.7305
R1600 OUT+.n30 OUT+.n29 2.7305
R1601 OUT+.n32 OUT+.t27 2.7305
R1602 OUT+.n32 OUT+.n31 2.7305
R1603 OUT+.n34 OUT+.t51 2.7305
R1604 OUT+.n34 OUT+.n33 2.7305
R1605 OUT+.n36 OUT+.t57 2.7305
R1606 OUT+.n36 OUT+.n35 2.7305
R1607 OUT+.n28 OUT+.t48 2.7305
R1608 OUT+.n28 OUT+.n27 2.7305
R1609 OUT+.n26 OUT+.t2 2.7305
R1610 OUT+.n26 OUT+.n25 2.7305
R1611 OUT+ OUT+.n0 2.25494
R1612 OUT+.n15 OUT+.n14 2.2505
R1613 OUT+.n84 OUT+.n83 2.2505
R1614 OUT+.n61 OUT+.n60 2.2505
R1615 OUT+.n38 OUT+.n37 2.2505
R1616 OUT+.n69 OUT+.n68 0.797345
R1617 OUT+.n23 OUT+.n22 0.797304
R1618 OUT+.n22 OUT+.n21 0.76828
R1619 OUT+.n91 OUT+.n90 0.76828
R1620 OUT+.n68 OUT+.n67 0.76828
R1621 OUT+.n45 OUT+.n44 0.76828
R1622 OUT+.n92 OUT+.n91 0.755717
R1623 OUT+.n46 OUT+.n45 0.755717
R1624 OUT+.n95 OUT+.n94 0.666333
R1625 OUT+.n94 OUT+.n93 0.6655
R1626 OUT+ OUT+.n95 0.618
R1627 OUT+.n16 OUT+.n15 0.60021
R1628 OUT+.n85 OUT+.n84 0.60021
R1629 OUT+.n62 OUT+.n61 0.60021
R1630 OUT+.n39 OUT+.n38 0.60021
R1631 OUT+.n17 OUT+.n16 0.59455
R1632 OUT+.n86 OUT+.n85 0.59455
R1633 OUT+.n63 OUT+.n62 0.59455
R1634 OUT+.n40 OUT+.n39 0.59455
R1635 OUT+.n20 OUT+.n17 0.58347
R1636 OUT+.n89 OUT+.n86 0.58347
R1637 OUT+.n66 OUT+.n63 0.58347
R1638 OUT+.n43 OUT+.n40 0.58347
R1639 IM IM.n30 32.4335
R1640 IM.n0 IM.t8 30.5343
R1641 IM.n0 IM.t4 18.1775
R1642 IM.n1 IM.t16 18.1775
R1643 IM.n4 IM.t12 18.1775
R1644 IM.n5 IM.t28 18.1775
R1645 IM.n8 IM.t25 18.1775
R1646 IM.n9 IM.t1 18.1775
R1647 IM.n12 IM.t11 18.1775
R1648 IM.n13 IM.t27 18.1775
R1649 IM.n16 IM.t29 18.1775
R1650 IM.n17 IM.t19 18.1775
R1651 IM.n20 IM.t18 18.1775
R1652 IM.n21 IM.t9 18.1775
R1653 IM.n24 IM.t26 18.1775
R1654 IM.n25 IM.t10 18.1775
R1655 IM.n28 IM.t13 18.1775
R1656 IM.n29 IM.t2 18.1775
R1657 IM.n2 IM.t5 17.6665
R1658 IM.n3 IM.t23 17.6665
R1659 IM.n6 IM.t24 17.6665
R1660 IM.n7 IM.t30 17.6665
R1661 IM.n10 IM.t3 17.6665
R1662 IM.n11 IM.t14 17.6665
R1663 IM.n14 IM.t22 17.6665
R1664 IM.n15 IM.t6 17.6665
R1665 IM.n18 IM.t31 17.6665
R1666 IM.n19 IM.t20 17.6665
R1667 IM.n22 IM.t15 17.6665
R1668 IM.n23 IM.t0 17.6665
R1669 IM.n26 IM.t21 17.6665
R1670 IM.n27 IM.t17 17.6665
R1671 IM.n30 IM.t7 17.6665
R1672 IM.n1 IM.n0 12.8683
R1673 IM.n2 IM.n1 12.8683
R1674 IM.n3 IM.n2 12.8683
R1675 IM.n4 IM.n3 12.8683
R1676 IM.n5 IM.n4 12.8683
R1677 IM.n6 IM.n5 12.8683
R1678 IM.n7 IM.n6 12.8683
R1679 IM.n8 IM.n7 12.8683
R1680 IM.n9 IM.n8 12.8683
R1681 IM.n10 IM.n9 12.8683
R1682 IM.n11 IM.n10 12.8683
R1683 IM.n12 IM.n11 12.8683
R1684 IM.n13 IM.n12 12.8683
R1685 IM.n14 IM.n13 12.8683
R1686 IM.n15 IM.n14 12.8683
R1687 IM.n16 IM.n15 12.8683
R1688 IM.n17 IM.n16 12.8683
R1689 IM.n18 IM.n17 12.8683
R1690 IM.n19 IM.n18 12.8683
R1691 IM.n20 IM.n19 12.8683
R1692 IM.n21 IM.n20 12.8683
R1693 IM.n22 IM.n21 12.8683
R1694 IM.n23 IM.n22 12.8683
R1695 IM.n24 IM.n23 12.8683
R1696 IM.n25 IM.n24 12.8683
R1697 IM.n26 IM.n25 12.8683
R1698 IM.n27 IM.n26 12.8683
R1699 IM.n28 IM.n27 12.8683
R1700 IM.n29 IM.n28 12.8683
R1701 IM.n30 IM.n29 12.8683
R1702 VDD.n11 VDD.t11 178.431
R1703 VDD.n24 VDD.t32 178.431
R1704 VDD.n20 VDD.t22 178.431
R1705 VDD.n16 VDD.t14 178.431
R1706 VDD.n38 VDD.t37 178.431
R1707 VDD.n34 VDD.t42 178.431
R1708 VDD.n30 VDD.t19 178.431
R1709 VDD.n7 VDD.t0 178.431
R1710 VDD.n3 VDD.t27 178.431
R1711 VDD.n11 VDD.t30 135.294
R1712 VDD.n24 VDD.t35 135.294
R1713 VDD.n20 VDD.t25 135.294
R1714 VDD.n16 VDD.t7 135.294
R1715 VDD.n38 VDD.t40 135.294
R1716 VDD.n34 VDD.t9 135.294
R1717 VDD.n30 VDD.t17 135.294
R1718 VDD.n7 VDD.t3 135.294
R1719 VDD.n3 VDD.t5 135.294
R1720 VDD.n17 VDD.n15 6.69527
R1721 VDD.n31 VDD.n29 6.69527
R1722 VDD.n4 VDD.n2 6.69527
R1723 VDD.n19 VDD.n14 6.59267
R1724 VDD.n23 VDD.n13 6.59267
R1725 VDD.n33 VDD.n28 6.59267
R1726 VDD.n37 VDD.n27 6.59267
R1727 VDD.n6 VDD.n1 6.59267
R1728 VDD.n10 VDD.n0 6.59267
R1729 VDD.n18 VDD.t8 6.55815
R1730 VDD.n22 VDD.t26 6.55815
R1731 VDD.n26 VDD.t36 6.55815
R1732 VDD.n32 VDD.t18 6.55815
R1733 VDD.n36 VDD.t10 6.55815
R1734 VDD.n40 VDD.t41 6.55815
R1735 VDD.n5 VDD.t6 6.55815
R1736 VDD.n9 VDD.t4 6.55815
R1737 VDD.n43 VDD.t31 6.55815
R1738 VDD.n17 VDD.n16 6.3005
R1739 VDD.n21 VDD.n20 6.3005
R1740 VDD.n25 VDD.n24 6.3005
R1741 VDD.n31 VDD.n30 6.3005
R1742 VDD.n35 VDD.n34 6.3005
R1743 VDD.n39 VDD.n38 6.3005
R1744 VDD.n4 VDD.n3 6.3005
R1745 VDD.n8 VDD.n7 6.3005
R1746 VDD.n12 VDD.n11 6.3005
R1747 VDD.n41 VDD.n40 3.87957
R1748 VDD.n42 VDD.n41 3.48326
R1749 VDD.n41 VDD.n26 2.58214
R1750 VDD.n19 VDD.n18 0.339604
R1751 VDD.n33 VDD.n32 0.339604
R1752 VDD.n6 VDD.n5 0.339604
R1753 VDD.n23 VDD.n22 0.302039
R1754 VDD.n37 VDD.n36 0.302039
R1755 VDD.n10 VDD.n9 0.302039
R1756 VDD.n43 VDD.n42 0.2717
R1757 VDD.n42 VDD 0.1883
R1758 VDD.n21 VDD.n19 0.1031
R1759 VDD.n25 VDD.n23 0.1031
R1760 VDD.n35 VDD.n33 0.1031
R1761 VDD.n39 VDD.n37 0.1031
R1762 VDD.n8 VDD.n6 0.1031
R1763 VDD.n12 VDD.n10 0.1031
R1764 VDD.n18 VDD 0.0893
R1765 VDD.n22 VDD 0.0893
R1766 VDD.n26 VDD 0.0893
R1767 VDD.n32 VDD 0.0893
R1768 VDD.n36 VDD 0.0893
R1769 VDD.n40 VDD 0.0893
R1770 VDD.n5 VDD 0.0893
R1771 VDD VDD.n43 0.0893
R1772 VDD.n9 VDD 0.0839
R1773 VDD VDD.n17 0.0017
R1774 VDD VDD.n21 0.0017
R1775 VDD VDD.n25 0.0017
R1776 VDD VDD.n31 0.0017
R1777 VDD VDD.n35 0.0017
R1778 VDD VDD.n39 0.0017
R1779 VDD VDD.n4 0.0017
R1780 VDD VDD.n8 0.0017
R1781 VDD VDD.n12 0.0017
R1782 Ci.n3 Ci.t1 28.2228
R1783 Ci.n0 Ci.t2 26.9784
R1784 Ci.n0 Ci.t0 14.7248
R1785 Ci.n3 Ci.t3 14.4701
R1786 Ci.n4 Ci.n3 4.5003
R1787 Ci.n1 Ci.n0 4.14631
R1788 Ci.n2 Ci 0.70023
R1789 Ci Ci.n4 0.0779
R1790 Ci.n2 Ci.n1 0.0635
R1791 Ci Ci.n2 0.0293
R1792 Ci.n4 Ci 0.0059
R1793 Ci.n1 Ci 0.0023
R1794 Ri.n3 Ri.t1 28.2228
R1795 Ri.n0 Ri.t2 26.9784
R1796 Ri.n0 Ri.t0 14.7248
R1797 Ri.n3 Ri.t3 14.4701
R1798 Ri.n4 Ri.n3 4.50813
R1799 Ri.n1 Ri.n0 4.15413
R1800 Ri.n2 Ri 0.4205
R1801 Ri.n2 Ri.n1 0.0924565
R1802 Ri Ri.n4 0.0885435
R1803 Ri.n4 Ri 0.00636957
R1804 Ri Ri.n2 0.00441304
R1805 Ri.n1 Ri 0.00245652
R1806 Ri-1.n2 Ri-1.t2 28.2228
R1807 Ri-1.n0 Ri-1.t1 26.9784
R1808 Ri-1.n0 Ri-1.t0 14.7248
R1809 Ri-1.n2 Ri-1.t3 14.4701
R1810 Ri-1.n3 Ri-1.n2 4.50813
R1811 Ri-1.n1 Ri-1.n0 4.15413
R1812 Ri-1.n4 Ri-1 0.768793
R1813 Ri-1 Ri-1.n1 0.086587
R1814 Ri-1.n4 Ri-1.n3 0.0787609
R1815 Ri-1 Ri-1.n4 0.0200652
R1816 Ri-1.n3 Ri-1 0.00636957
R1817 Ri-1.n1 Ri-1 0.00245652
C0 SD Ri 9.7e-19
C1 SD QB 0.00262f
C2 Local_Enc_0.NAND_7.SD Q 1.23e-19
C3 Local_Enc_0.NAND_5.A Local_Enc_0.NAND_6.A 0.216f
C4 IM_T Local_Enc_0.NAND_6.A 0.00339f
C5 Local_Enc_0.NAND_5.A OUT 0.00106f
C6 OUT- OUT 8.42f
C7 IM_T OUT 0.762f
C8 VDD Q 0.588f
C9 VDD Local_Enc_0.NAND_6.B 0.618f
C10 Local_Enc_0.NAND_6.SD Local_Enc_0.NAND_6.B 0.00403f
C11 IM Local_Enc_0.NAND_4.B 1.99e-19
C12 VDD Local_Enc_0.NAND_0.SD 8.42e-19
C13 OUT+ OUT- 8.48f
C14 VDD Local_Enc_0.NAND_6.A 0.358f
C15 OUT+ IM_T 0.00188f
C16 Local_Enc_0.NAND_6.SD Local_Enc_0.NAND_6.A 0.0812f
C17 QB Local_Enc_0.NAND_5.B 0.00682f
C18 Local_Enc_0.NAND_8.A Local_Enc_0.NAND_4.B 0.345f
C19 Ci Local_Enc_0.NAND_5.A 0.00328f
C20 IM Q 7.41e-19
C21 IM Local_Enc_0.NAND_6.B 0.00136f
C22 Local_Enc_0.NAND_2.SD Ri 5.71e-20
C23 Q Local_Enc_0.NAND_8.A 0.208f
C24 IM OUT 1.33f
C25 Local_Enc_0.NAND_1.B Local_Enc_0.NAND_5.B 0.344f
C26 Local_Enc_0.NAND_8.A Local_Enc_0.NAND_6.B 0.00405f
C27 Ci VDD 0.478f
C28 Local_Enc_0.NAND_1.SD Local_Enc_0.NAND_5.A 5.76e-20
C29 Ri Local_Enc_0.NAND_3.SD 0.0852f
C30 SD Local_Enc_0.NAND_4.B 0.00299f
C31 Local_Enc_0.NAND_8.A Local_Enc_0.NAND_6.A 0.0124f
C32 OUT Local_Enc_0.NAND_8.A 1.41e-19
C33 OUT+ IM 8.52e-21
C34 VDD Ri-1 0.546f
C35 SD Q 0.00613f
C36 OUT+ Local_Enc_0.NAND_8.A 7.56e-20
C37 SD Local_Enc_0.NAND_6.B 0.00526f
C38 Local_Enc_0.NAND_4.B Local_Enc_0.NAND_5.B 0.026f
C39 SD Local_Enc_0.NAND_6.A 0.00198f
C40 Ci Local_Enc_0.NAND_8.A 9.39e-19
C41 SD OUT 4.67f
C42 Local_Enc_0.NAND_4.SD Local_Enc_0.NAND_8.A 5.76e-20
C43 Q Local_Enc_0.NAND_5.B 0.0478f
C44 OUT+ SD 0.00427f
C45 Local_Enc_0.NAND_6.B Local_Enc_0.NAND_5.B 0.0342f
C46 Local_Enc_0.NAND_6.B Local_Enc_0.NAND_5.SD 2.79e-20
C47 Local_Enc_0.NAND_5.B Local_Enc_0.NAND_0.SD 0.00175f
C48 IM_T Local_Enc_0.NAND_5.A 0.00438f
C49 OUT- IM_T 0.0213f
C50 Local_Enc_0.NAND_5.SD Local_Enc_0.NAND_6.A 5.69e-20
C51 Local_Enc_0.NAND_6.B Local_Enc_0.NAND_2.SD 0.0444f
C52 Local_Enc_0.NAND_7.SD Local_Enc_0.NAND_5.A 1.88e-20
C53 Local_Enc_0.NAND_7.SD IM_T 2.11e-19
C54 Local_Enc_0.NAND_5.A VDD 0.503f
C55 IM_T VDD 0.00972f
C56 Local_Enc_0.NAND_6.SD Local_Enc_0.NAND_5.A 0.0451f
C57 Local_Enc_0.NAND_6.A Local_Enc_0.NAND_3.SD 0.0419f
C58 Ci Local_Enc_0.NAND_5.B 0.0105f
C59 Local_Enc_0.NAND_6.SD IM_T 2.11e-19
C60 Local_Enc_0.NAND_4.SD Local_Enc_0.NAND_5.B 6.99e-20
C61 Ri-1 Local_Enc_0.NAND_5.B 0.0106f
C62 Ci Local_Enc_0.NAND_2.SD 0.0852f
C63 IM Local_Enc_0.NAND_5.A 0.00213f
C64 OUT- IM 0.0126f
C65 IM_T IM 2.05f
C66 Local_Enc_0.NAND_1.SD Local_Enc_0.NAND_5.B 0.0469f
C67 Local_Enc_0.NAND_5.A Local_Enc_0.NAND_8.A 0.333f
C68 OUT- Local_Enc_0.NAND_8.A 1.62e-19
C69 IM_T Local_Enc_0.NAND_8.A 0.0073f
C70 Local_Enc_0.NAND_7.SD Local_Enc_0.NAND_8.A 0.0852f
C71 VDD Local_Enc_0.NAND_8.A 0.864f
C72 SD Local_Enc_0.NAND_5.A 0.0153f
C73 OUT- SD 0.0307f
C74 IM_T SD 1f
C75 QB Local_Enc_0.NAND_8.SD 0.0055f
C76 Local_Enc_0.NAND_7.SD SD 3.62e-19
C77 IM Local_Enc_0.NAND_8.A 3.24e-19
C78 QB Local_Enc_0.NAND_1.B 1.31e-19
C79 SD VDD 0.00235f
C80 Local_Enc_0.NAND_6.SD SD 3.72e-19
C81 Local_Enc_0.NAND_5.A Local_Enc_0.NAND_5.B 0.316f
C82 Local_Enc_0.NAND_5.A Local_Enc_0.NAND_5.SD 0.0874f
C83 IM_T Local_Enc_0.NAND_5.SD 1.47e-20
C84 IM SD 0.916f
C85 VDD Local_Enc_0.NAND_5.B 0.864f
C86 Local_Enc_0.NAND_5.A Local_Enc_0.NAND_2.SD 2.15e-19
C87 IM_T Local_Enc_0.NAND_2.SD 1.47e-20
C88 Ri Local_Enc_0.NAND_4.B 2.34e-22
C89 QB Local_Enc_0.NAND_4.B 0.495f
C90 SD Local_Enc_0.NAND_8.A 0.00473f
C91 IM_T Local_Enc_0.NAND_3.SD 2.11e-19
C92 Local_Enc_0.NAND_8.SD Local_Enc_0.NAND_4.B 0.00331f
C93 Q QB 5.71f
C94 Local_Enc_0.NAND_6.B Ri 0.0132f
C95 QB Local_Enc_0.NAND_6.B 4.6e-19
C96 Local_Enc_0.NAND_1.B Local_Enc_0.NAND_4.B 0.00819f
C97 Q Local_Enc_0.NAND_8.SD 0.043f
C98 Ri Local_Enc_0.NAND_6.A 0.233f
C99 QB OUT 2.71f
C100 Local_Enc_0.NAND_8.A Local_Enc_0.NAND_5.B 0.0646f
C101 Q Local_Enc_0.NAND_1.B 0.004f
C102 Local_Enc_0.NAND_8.A Local_Enc_0.NAND_5.SD 0.045f
C103 Local_Enc_0.NAND_6.B Local_Enc_0.NAND_1.B 1.35e-19
C104 OUT+ QB 1.83f
C105 Local_Enc_0.NAND_1.B Local_Enc_0.NAND_0.SD 0.0419f
C106 Ci Ri 0.0212f
C107 Ci QB 5.92e-19
C108 Local_Enc_0.NAND_4.SD QB 0.0423f
C109 Q Local_Enc_0.NAND_4.B 0.686f
C110 Local_Enc_0.NAND_6.B Local_Enc_0.NAND_4.B 2.09e-20
C111 SD Local_Enc_0.NAND_3.SD 4.2e-19
C112 Local_Enc_0.NAND_6.A Local_Enc_0.NAND_4.B 1.31e-19
C113 OUT Local_Enc_0.NAND_4.B 2.29e-19
C114 Ri-1 Local_Enc_0.NAND_1.B 0.24f
C115 Local_Enc_0.NAND_5.SD Local_Enc_0.NAND_5.B 0.0043f
C116 Local_Enc_0.NAND_1.SD Local_Enc_0.NAND_1.B 0.0852f
C117 Q OUT 4.21f
C118 Local_Enc_0.NAND_6.B Local_Enc_0.NAND_6.A 0.429f
C119 OUT Local_Enc_0.NAND_6.B 1.93e-19
C120 OUT+ Q 1.2f
C121 Local_Enc_0.NAND_4.SD Local_Enc_0.NAND_4.B 0.00495f
C122 Ri-1 Local_Enc_0.NAND_4.B 1.08e-19
C123 Ci Local_Enc_0.NAND_6.B 0.235f
C124 OUT+ OUT 7.38f
C125 Local_Enc_0.NAND_4.SD Q 0.0961f
C126 Ci Local_Enc_0.NAND_0.SD 5.76e-20
C127 Local_Enc_0.NAND_5.A Ri 9.5e-19
C128 Ci Local_Enc_0.NAND_6.A 1.17e-19
C129 IM_T Ri 0.00546f
C130 OUT- QB 1.7f
C131 Local_Enc_0.NAND_5.A QB 0.00927f
C132 IM_T QB 0.00321f
C133 Ri-1 Local_Enc_0.NAND_6.B 1.18e-19
C134 Local_Enc_0.NAND_1.SD Q 6.06e-19
C135 Local_Enc_0.NAND_7.SD Ri 3.42e-22
C136 IM_T Local_Enc_0.NAND_8.SD 1.47e-20
C137 Local_Enc_0.NAND_7.SD QB 3.34e-19
C138 Ri-1 Local_Enc_0.NAND_0.SD 0.0852f
C139 VDD Ri 0.406f
C140 VDD QB 0.639f
C141 Local_Enc_0.NAND_6.SD Ri 1.61e-21
C142 Local_Enc_0.NAND_5.A Local_Enc_0.NAND_1.B 0.00251f
C143 VDD Local_Enc_0.NAND_1.B 0.628f
C144 Ci Ri-1 0.0236f
C145 IM Ri 1.66e-21
C146 IM QB 7.5e-19
C147 Local_Enc_0.NAND_8.A Ri 5.57e-19
C148 QB Local_Enc_0.NAND_8.A 0.43f
C149 Local_Enc_0.NAND_5.A Local_Enc_0.NAND_4.B 0.00496f
C150 IM_T Local_Enc_0.NAND_4.B 0.00103f
C151 Local_Enc_0.NAND_8.A Local_Enc_0.NAND_8.SD 0.0821f
C152 Local_Enc_0.NAND_7.SD Local_Enc_0.NAND_4.B 0.0419f
C153 Local_Enc_0.NAND_5.A Q 2.28e-19
C154 OUT- Q 1.19f
C155 Local_Enc_0.NAND_8.A Local_Enc_0.NAND_1.B 1.18e-19
C156 IM_T Q 0.0573f
C157 VDD Local_Enc_0.NAND_4.B 0.673f
C158 Local_Enc_0.NAND_5.A Local_Enc_0.NAND_6.B 0.232f
C159 IM_T Local_Enc_0.NAND_6.B 0.00448f
C160 OUT- VSS 3.05f
C161 OUT+ VSS 3.87f
C162 SD VSS 5.44f
C163 IM VSS 8.4f
C164 IM_T VSS 15.2f
C165 Local_Enc_0.NAND_7.SD VSS 0.0983f
C166 Local_Enc_0.NAND_6.SD VSS 0.0986f
C167 Local_Enc_0.NAND_3.SD VSS 0.0998f
C168 Local_Enc_0.NAND_6.A VSS 0.56f
C169 Ri VSS 0.977f
C170 Local_Enc_0.NAND_8.SD VSS 0.0983f
C171 Local_Enc_0.NAND_5.SD VSS 0.0983f
C172 Local_Enc_0.NAND_2.SD VSS 0.0997f
C173 Local_Enc_0.NAND_6.B VSS 0.669f
C174 Local_Enc_0.NAND_8.A VSS 1.42f
C175 Local_Enc_0.NAND_5.A VSS 0.674f
C176 Ci VSS 0.927f
C177 Local_Enc_0.NAND_4.SD VSS 0.0983f
C178 Local_Enc_0.NAND_1.SD VSS 0.0983f
C179 Local_Enc_0.NAND_0.SD VSS 0.0983f
C180 Local_Enc_0.NAND_5.B VSS 0.695f
C181 Local_Enc_0.NAND_4.B VSS 0.67f
C182 Local_Enc_0.NAND_1.B VSS 0.754f
C183 Ri-1 VSS 0.848f
C184 OUT VSS 9.62f
C185 QB VSS 18.2f
C186 Q VSS 20f
C187 VDD VSS 14f
C188 IM.t8 VSS 0.0417f
C189 IM.t4 VSS 0.0306f
C190 IM.n0 VSS 0.0488f
C191 IM.t16 VSS 0.0306f
C192 IM.n1 VSS 0.0328f
C193 IM.t5 VSS 0.03f
C194 IM.n2 VSS 0.0324f
C195 IM.t23 VSS 0.03f
C196 IM.n3 VSS 0.0324f
C197 IM.t12 VSS 0.0306f
C198 IM.n4 VSS 0.0328f
C199 IM.t28 VSS 0.0306f
C200 IM.n5 VSS 0.0328f
C201 IM.t24 VSS 0.03f
C202 IM.n6 VSS 0.0324f
C203 IM.t30 VSS 0.03f
C204 IM.n7 VSS 0.0324f
C205 IM.t25 VSS 0.0306f
C206 IM.n8 VSS 0.0328f
C207 IM.t1 VSS 0.0306f
C208 IM.n9 VSS 0.0328f
C209 IM.t3 VSS 0.03f
C210 IM.n10 VSS 0.0324f
C211 IM.t14 VSS 0.03f
C212 IM.n11 VSS 0.0324f
C213 IM.t11 VSS 0.0306f
C214 IM.n12 VSS 0.0328f
C215 IM.t27 VSS 0.0306f
C216 IM.n13 VSS 0.0328f
C217 IM.t22 VSS 0.03f
C218 IM.n14 VSS 0.0324f
C219 IM.t6 VSS 0.03f
C220 IM.n15 VSS 0.0324f
C221 IM.t29 VSS 0.0306f
C222 IM.n16 VSS 0.0328f
C223 IM.t19 VSS 0.0306f
C224 IM.n17 VSS 0.0328f
C225 IM.t31 VSS 0.03f
C226 IM.n18 VSS 0.0324f
C227 IM.t20 VSS 0.03f
C228 IM.n19 VSS 0.0324f
C229 IM.t18 VSS 0.0306f
C230 IM.n20 VSS 0.0328f
C231 IM.t9 VSS 0.0306f
C232 IM.n21 VSS 0.0328f
C233 IM.t15 VSS 0.03f
C234 IM.n22 VSS 0.0324f
C235 IM.t0 VSS 0.03f
C236 IM.n23 VSS 0.0324f
C237 IM.t26 VSS 0.0306f
C238 IM.n24 VSS 0.0328f
C239 IM.t10 VSS 0.0306f
C240 IM.n25 VSS 0.0328f
C241 IM.t21 VSS 0.03f
C242 IM.n26 VSS 0.0324f
C243 IM.t17 VSS 0.03f
C244 IM.n27 VSS 0.0324f
C245 IM.t13 VSS 0.0306f
C246 IM.n28 VSS 0.0328f
C247 IM.t2 VSS 0.0306f
C248 IM.n29 VSS 0.0328f
C249 IM.t7 VSS 0.03f
C250 IM.n30 VSS 0.0405f
C251 OUT+.n0 VSS 0.0484f
C252 OUT+.n1 VSS 0.0527f
C253 OUT+.t30 VSS 0.0222f
C254 OUT+.n2 VSS 0.0222f
C255 OUT+.n3 VSS 0.0526f
C256 OUT+.t34 VSS 0.0222f
C257 OUT+.n4 VSS 0.0222f
C258 OUT+.n5 VSS 0.0459f
C259 OUT+.t24 VSS 0.0222f
C260 OUT+.n6 VSS 0.0222f
C261 OUT+.n7 VSS 0.077f
C262 OUT+.t55 VSS 0.0222f
C263 OUT+.n8 VSS 0.0222f
C264 OUT+.n9 VSS 0.101f
C265 OUT+.t38 VSS 0.0222f
C266 OUT+.n10 VSS 0.0222f
C267 OUT+.n11 VSS 0.0459f
C268 OUT+.t18 VSS 0.0222f
C269 OUT+.n12 VSS 0.0222f
C270 OUT+.n13 VSS 0.081f
C271 OUT+.n14 VSS 0.285f
C272 OUT+.t4 VSS 0.115f
C273 OUT+.n15 VSS 0.479f
C274 OUT+.n16 VSS 0.295f
C275 OUT+.n17 VSS 0.21f
C276 OUT+.t16 VSS 0.0222f
C277 OUT+.n18 VSS 0.0222f
C278 OUT+.n19 VSS 0.1f
C279 OUT+.n20 VSS 0.37f
C280 OUT+.n21 VSS 0.177f
C281 OUT+.n22 VSS 0.226f
C282 OUT+.n23 VSS 0.266f
C283 OUT+.n24 VSS 0.0533f
C284 OUT+.t2 VSS 0.0222f
C285 OUT+.n25 VSS 0.0222f
C286 OUT+.n26 VSS 0.0526f
C287 OUT+.t48 VSS 0.0222f
C288 OUT+.n27 VSS 0.0222f
C289 OUT+.n28 VSS 0.0459f
C290 OUT+.t37 VSS 0.0222f
C291 OUT+.n29 VSS 0.0222f
C292 OUT+.n30 VSS 0.077f
C293 OUT+.t27 VSS 0.0222f
C294 OUT+.n31 VSS 0.0222f
C295 OUT+.n32 VSS 0.101f
C296 OUT+.t51 VSS 0.0222f
C297 OUT+.n33 VSS 0.0222f
C298 OUT+.n34 VSS 0.0459f
C299 OUT+.t57 VSS 0.0222f
C300 OUT+.n35 VSS 0.0222f
C301 OUT+.n36 VSS 0.081f
C302 OUT+.n37 VSS 0.285f
C303 OUT+.t17 VSS 0.115f
C304 OUT+.n38 VSS 0.479f
C305 OUT+.n39 VSS 0.295f
C306 OUT+.n40 VSS 0.21f
C307 OUT+.t54 VSS 0.0222f
C308 OUT+.n41 VSS 0.0222f
C309 OUT+.n42 VSS 0.1f
C310 OUT+.n43 VSS 0.37f
C311 OUT+.n44 VSS 0.177f
C312 OUT+.n45 VSS 0.222f
C313 OUT+.n46 VSS 0.27f
C314 OUT+.n47 VSS 0.0527f
C315 OUT+.t35 VSS 0.0222f
C316 OUT+.n48 VSS 0.0222f
C317 OUT+.n49 VSS 0.0526f
C318 OUT+.t21 VSS 0.0222f
C319 OUT+.n50 VSS 0.0222f
C320 OUT+.n51 VSS 0.0459f
C321 OUT+.t11 VSS 0.0222f
C322 OUT+.n52 VSS 0.0222f
C323 OUT+.n53 VSS 0.077f
C324 OUT+.t1 VSS 0.0222f
C325 OUT+.n54 VSS 0.0222f
C326 OUT+.n55 VSS 0.101f
C327 OUT+.t23 VSS 0.0222f
C328 OUT+.n56 VSS 0.0222f
C329 OUT+.n57 VSS 0.0459f
C330 OUT+.t29 VSS 0.0222f
C331 OUT+.n58 VSS 0.0222f
C332 OUT+.n59 VSS 0.081f
C333 OUT+.n60 VSS 0.285f
C334 OUT+.t56 VSS 0.115f
C335 OUT+.n61 VSS 0.479f
C336 OUT+.n62 VSS 0.295f
C337 OUT+.n63 VSS 0.21f
C338 OUT+.t26 VSS 0.0222f
C339 OUT+.n64 VSS 0.0222f
C340 OUT+.n65 VSS 0.1f
C341 OUT+.n66 VSS 0.37f
C342 OUT+.n67 VSS 0.177f
C343 OUT+.n68 VSS 0.226f
C344 OUT+.n69 VSS 0.265f
C345 OUT+.n70 VSS 0.0533f
C346 OUT+.t50 VSS 0.0222f
C347 OUT+.n71 VSS 0.0222f
C348 OUT+.n72 VSS 0.0526f
C349 OUT+.t61 VSS 0.0222f
C350 OUT+.n73 VSS 0.0222f
C351 OUT+.n74 VSS 0.0459f
C352 OUT+.t46 VSS 0.0222f
C353 OUT+.n75 VSS 0.0222f
C354 OUT+.n76 VSS 0.077f
C355 OUT+.t12 VSS 0.0222f
C356 OUT+.n77 VSS 0.0222f
C357 OUT+.n78 VSS 0.101f
C358 OUT+.t0 VSS 0.0222f
C359 OUT+.n79 VSS 0.0222f
C360 OUT+.n80 VSS 0.0459f
C361 OUT+.t40 VSS 0.0222f
C362 OUT+.n81 VSS 0.0222f
C363 OUT+.n82 VSS 0.081f
C364 OUT+.n83 VSS 0.285f
C365 OUT+.t28 VSS 0.115f
C366 OUT+.n84 VSS 0.479f
C367 OUT+.n85 VSS 0.295f
C368 OUT+.n86 VSS 0.21f
C369 OUT+.t39 VSS 0.0222f
C370 OUT+.n87 VSS 0.0222f
C371 OUT+.n88 VSS 0.1f
C372 OUT+.n89 VSS 0.37f
C373 OUT+.n90 VSS 0.177f
C374 OUT+.n91 VSS 0.222f
C375 OUT+.n92 VSS 0.338f
C376 OUT+.n93 VSS 0.912f
C377 OUT+.n94 VSS 0.625f
C378 OUT+.n95 VSS 0.605f
C379 Q.n0 VSS 0.0122f
C380 Q.t14 VSS 0.0669f
C381 Q.t31 VSS 0.0398f
C382 Q.n1 VSS 0.114f
C383 Q.t24 VSS 0.0398f
C384 Q.n2 VSS 0.0761f
C385 Q.t5 VSS 0.0412f
C386 Q.n3 VSS 0.0779f
C387 Q.t43 VSS 0.0412f
C388 Q.n4 VSS 0.0779f
C389 Q.t42 VSS 0.0398f
C390 Q.n5 VSS 0.0761f
C391 Q.t6 VSS 0.0398f
C392 Q.n6 VSS 0.0761f
C393 Q.t20 VSS 0.0412f
C394 Q.n7 VSS 0.0779f
C395 Q.t55 VSS 0.0412f
C396 Q.n8 VSS 0.0779f
C397 Q.t67 VSS 0.0398f
C398 Q.n9 VSS 0.0761f
C399 Q.t22 VSS 0.0398f
C400 Q.n10 VSS 0.0761f
C401 Q.t68 VSS 0.0412f
C402 Q.n11 VSS 0.0779f
C403 Q.t23 VSS 0.0412f
C404 Q.n12 VSS 0.0779f
C405 Q.t39 VSS 0.0398f
C406 Q.n13 VSS 0.0761f
C407 Q.t4 VSS 0.0398f
C408 Q.n14 VSS 0.0824f
C409 Q.t40 VSS 0.0357f
C410 Q.n15 VSS 0.0765f
C411 Q.t35 VSS 0.133f
C412 Q.t32 VSS 0.0412f
C413 Q.n16 VSS 0.161f
C414 Q.t65 VSS 0.0412f
C415 Q.n17 VSS 0.134f
C416 Q.t44 VSS 0.0412f
C417 Q.n18 VSS 0.134f
C418 Q.t7 VSS 0.0412f
C419 Q.n19 VSS 0.134f
C420 Q.t28 VSS 0.0412f
C421 Q.n20 VSS 0.134f
C422 Q.t48 VSS 0.0412f
C423 Q.n21 VSS 0.138f
C424 Q.t64 VSS 0.0357f
C425 Q.n22 VSS 0.169f
C426 Q.t21 VSS 0.0669f
C427 Q.t38 VSS 0.0398f
C428 Q.n23 VSS 0.114f
C429 Q.t34 VSS 0.0398f
C430 Q.n24 VSS 0.0761f
C431 Q.t18 VSS 0.0412f
C432 Q.n25 VSS 0.0779f
C433 Q.t53 VSS 0.0412f
C434 Q.n26 VSS 0.0779f
C435 Q.t52 VSS 0.0398f
C436 Q.n27 VSS 0.0761f
C437 Q.t19 VSS 0.0398f
C438 Q.n28 VSS 0.0761f
C439 Q.t29 VSS 0.0412f
C440 Q.n29 VSS 0.0779f
C441 Q.t63 VSS 0.0412f
C442 Q.n30 VSS 0.0779f
C443 Q.t11 VSS 0.0398f
C444 Q.n31 VSS 0.0761f
C445 Q.t30 VSS 0.0398f
C446 Q.n32 VSS 0.0761f
C447 Q.t15 VSS 0.0412f
C448 Q.n33 VSS 0.0779f
C449 Q.t33 VSS 0.0412f
C450 Q.n34 VSS 0.0779f
C451 Q.t50 VSS 0.0398f
C452 Q.n35 VSS 0.0761f
C453 Q.t17 VSS 0.0398f
C454 Q.n36 VSS 0.0824f
C455 Q.t51 VSS 0.0357f
C456 Q.n37 VSS 0.0942f
C457 Q.n38 VSS 0.333f
C458 Q.t54 VSS 0.0669f
C459 Q.t66 VSS 0.0398f
C460 Q.n39 VSS 0.114f
C461 Q.t61 VSS 0.0398f
C462 Q.n40 VSS 0.0761f
C463 Q.t47 VSS 0.0412f
C464 Q.n41 VSS 0.0779f
C465 Q.t13 VSS 0.0412f
C466 Q.n42 VSS 0.0779f
C467 Q.t12 VSS 0.0398f
C468 Q.n43 VSS 0.0761f
C469 Q.t49 VSS 0.0398f
C470 Q.n44 VSS 0.0761f
C471 Q.t57 VSS 0.0412f
C472 Q.n45 VSS 0.0779f
C473 Q.t25 VSS 0.0412f
C474 Q.n46 VSS 0.0779f
C475 Q.t41 VSS 0.0398f
C476 Q.n47 VSS 0.0761f
C477 Q.t58 VSS 0.0398f
C478 Q.n48 VSS 0.0761f
C479 Q.t45 VSS 0.0412f
C480 Q.n49 VSS 0.0779f
C481 Q.t60 VSS 0.0412f
C482 Q.n50 VSS 0.0779f
C483 Q.t9 VSS 0.0398f
C484 Q.n51 VSS 0.0761f
C485 Q.t46 VSS 0.0398f
C486 Q.n52 VSS 0.0824f
C487 Q.t10 VSS 0.0357f
C488 Q.n53 VSS 0.0942f
C489 Q.n54 VSS 0.212f
C490 Q.t16 VSS 0.0641f
C491 Q.t8 VSS 0.0373f
C492 Q.n55 VSS 0.118f
C493 Q.t27 VSS 0.0373f
C494 Q.n56 VSS 0.0952f
C495 Q.t62 VSS 0.0373f
C496 Q.n57 VSS 0.0952f
C497 Q.t56 VSS 0.0373f
C498 Q.n58 VSS 0.0952f
C499 Q.t3 VSS 0.0373f
C500 Q.n59 VSS 0.0952f
C501 Q.t26 VSS 0.0373f
C502 Q.n60 VSS 0.0952f
C503 Q.t59 VSS 0.0373f
C504 Q.n61 VSS 0.0913f
C505 Q.n62 VSS 0.336f
C506 Q.n63 VSS 0.163f
C507 Q.n64 VSS 5.71e-19
C508 Q.n65 VSS 0.0225f
C509 Q.t36 VSS 0.0234f
C510 Q.t37 VSS 0.0134f
C511 Q.n66 VSS 0.0611f
C512 Q.t1 VSS 0.00924f
C513 Q.n67 VSS 0.00924f
C514 Q.n68 VSS 0.0185f
C515 Q.n69 VSS 0.158f
C516 Q.n70 VSS 0.0836f
C517 SD.n0 VSS 0.0127f
C518 SD.t43 VSS 0.0151f
C519 SD.n1 VSS 0.0561f
C520 SD.n2 VSS 0.0689f
C521 SD.t49 VSS 0.0128f
C522 SD.n3 VSS 0.0149f
C523 SD.n4 VSS 0.0557f
C524 SD.t37 VSS 0.015f
C525 SD.n5 VSS 0.0128f
C526 SD.n6 VSS 0.0452f
C527 SD.t50 VSS 0.0136f
C528 SD.n7 VSS 0.0136f
C529 SD.n8 VSS 0.0276f
C530 SD.n9 VSS 0.0312f
C531 SD.t26 VSS 0.0136f
C532 SD.n10 VSS 0.0136f
C533 SD.n11 VSS 0.0532f
C534 SD.t9 VSS 0.0136f
C535 SD.n12 VSS 0.0136f
C536 SD.n13 VSS 0.0541f
C537 SD.t63 VSS 0.0136f
C538 SD.n14 VSS 0.0136f
C539 SD.n15 VSS 0.0276f
C540 SD.n16 VSS 0.0312f
C541 SD.t20 VSS 0.015f
C542 SD.n17 VSS 0.0128f
C543 SD.n18 VSS 0.0563f
C544 SD.t58 VSS 0.0136f
C545 SD.n19 VSS 0.0136f
C546 SD.n20 VSS 0.053f
C547 SD.t36 VSS 0.0136f
C548 SD.n21 VSS 0.0136f
C549 SD.n22 VSS 0.053f
C550 SD.t56 VSS 0.0136f
C551 SD.n23 VSS 0.0136f
C552 SD.n24 VSS 0.0276f
C553 SD.n25 VSS 0.0312f
C554 SD.n26 VSS 0.0127f
C555 SD.t1 VSS 0.0151f
C556 SD.n27 VSS 0.0563f
C557 SD.t29 VSS 0.0136f
C558 SD.n28 VSS 0.0136f
C559 SD.n29 VSS 0.0276f
C560 SD.n30 VSS 0.0312f
C561 SD.t40 VSS 0.0136f
C562 SD.n31 VSS 0.0136f
C563 SD.n32 VSS 0.0529f
C564 SD.t55 VSS 0.0149f
C565 SD.n33 VSS 0.0128f
C566 SD.n34 VSS 0.0559f
C567 SD.t44 VSS 0.0136f
C568 SD.n35 VSS 0.0136f
C569 SD.n36 VSS 0.0276f
C570 SD.n37 VSS 0.0312f
C571 SD.t14 VSS 0.0136f
C572 SD.n38 VSS 0.0136f
C573 SD.n39 VSS 0.0413f
C574 SD.t23 VSS 0.0133f
C575 SD.n40 VSS 0.0144f
C576 SD.n41 VSS 0.0567f
C577 SD.n42 VSS 0.125f
C578 SD.n43 VSS 0.0272f
C579 SD.n44 VSS 0.0724f
C580 SD.n45 VSS 0.0268f
C581 SD.t6 VSS 0.0128f
C582 SD.n46 VSS 0.0149f
C583 SD.n47 VSS 0.0271f
C584 SD.n48 VSS 0.0312f
C585 SD.n49 VSS 0.0284f
C586 SD.n50 VSS 0.0746f
C587 SD.n51 VSS 0.0258f
C588 SD.n52 VSS 0.0263f
C589 SD.n53 VSS 0.0737f
C590 SD.n54 VSS 0.0262f
C591 SD.n55 VSS 0.0273f
C592 SD.n56 VSS 0.077f
C593 SD.n57 VSS 0.0269f
C594 SD.n58 VSS 0.029f
C595 SD.n59 VSS 0.0756f
C596 SD.n60 VSS 0.0149f
C597 SD.t24 VSS 0.0128f
C598 SD.n61 VSS 0.0271f
C599 SD.n62 VSS 0.0312f
C600 SD.n63 VSS 0.027f
C601 SD.n64 VSS 0.026f
C602 SD.n65 VSS 0.0738f
C603 SD.n66 VSS 0.027f
C604 SD.n67 VSS 0.0282f
C605 SD.n68 VSS 0.075f
C606 SD.t31 VSS 0.0128f
C607 SD.n69 VSS 0.015f
C608 SD.n70 VSS 0.0273f
C609 SD.n71 VSS 0.0312f
C610 SD.n72 VSS 0.0256f
C611 SD.n73 VSS 0.0263f
C612 SD.n74 VSS 0.0778f
C613 SD.n75 VSS 0.0262f
C614 SD.n76 VSS 0.0402f
C615 SD.n77 VSS 0.0979f
C616 SD.n78 VSS 0.0286f
C617 SD.t10 VSS 0.0129f
C618 SD.n79 VSS 0.0148f
C619 SD.n80 VSS 0.0272f
C620 SD.n81 VSS 0.0312f
C621 SD.n82 VSS 7.96e-19
C622 SD.t0 VSS 0.0136f
C623 SD.n83 VSS 0.0136f
C624 SD.n84 VSS 0.0522f
C625 SD.t34 VSS 0.0136f
C626 SD.n85 VSS 0.0136f
C627 SD.n86 VSS 0.0527f
C628 SD.t54 VSS 0.015f
C629 SD.n87 VSS 0.0128f
C630 SD.n88 VSS 0.0558f
C631 SD.t17 VSS 0.0136f
C632 SD.n89 VSS 0.0136f
C633 SD.n90 VSS 0.0535f
C634 SD.t2 VSS 0.0136f
C635 SD.n91 VSS 0.0136f
C636 SD.n92 VSS 0.0538f
C637 SD.t22 VSS 0.0136f
C638 SD.n93 VSS 0.0136f
C639 SD.n94 VSS 0.0412f
C640 SD.n95 VSS 0.129f
C641 SD.n96 VSS 0.0282f
C642 SD.n97 VSS 0.0761f
C643 SD.t5 VSS 0.0146f
C644 SD.n98 VSS 0.0132f
C645 SD.n99 VSS 0.0272f
C646 SD.n100 VSS 0.0312f
C647 SD.n101 VSS 0.027f
C648 SD.t48 VSS 0.0136f
C649 SD.n102 VSS 0.0136f
C650 SD.n103 VSS 0.0277f
C651 SD.n104 VSS 0.0311f
C652 SD.n105 VSS 0.0265f
C653 SD.n106 VSS 0.0723f
C654 SD.n107 VSS 0.0267f
C655 SD.n108 VSS 0.101f
C656 SD.n109 VSS 0.0127f
C657 SD.t3 VSS 0.0151f
C658 SD.n110 VSS 0.0451f
C659 SD.n111 VSS 0.0398f
C660 SD.n112 VSS 0.0263f
C661 SD.n113 VSS 0.0752f
C662 SD.t18 VSS 0.0136f
C663 SD.n114 VSS 0.0136f
C664 SD.n115 VSS 0.0277f
C665 SD.n116 VSS 0.0311f
C666 SD.n117 VSS 0.0252f
C667 SD.n118 VSS 0.0258f
C668 IM_T.n0 VSS 0.00126f
C669 IM_T.n1 VSS 0.0159f
C670 IM_T.t27 VSS 0.0309f
C671 IM_T.t4 VSS 0.0225f
C672 IM_T.n2 VSS 0.0496f
C673 IM_T.t2 VSS 0.0225f
C674 IM_T.n3 VSS 0.0374f
C675 IM_T.t19 VSS 0.0225f
C676 IM_T.n4 VSS 0.0374f
C677 IM_T.t15 VSS 0.0225f
C678 IM_T.n5 VSS 0.0374f
C679 IM_T.t24 VSS 0.0225f
C680 IM_T.n6 VSS 0.0374f
C681 IM_T.t1 VSS 0.0225f
C682 IM_T.n7 VSS 0.0374f
C683 IM_T.t17 VSS 0.0225f
C684 IM_T.n8 VSS 0.0374f
C685 IM_T.t18 VSS 0.0225f
C686 IM_T.n9 VSS 0.0374f
C687 IM_T.t11 VSS 0.0225f
C688 IM_T.n10 VSS 0.0374f
C689 IM_T.t10 VSS 0.0225f
C690 IM_T.n11 VSS 0.0374f
C691 IM_T.t30 VSS 0.0225f
C692 IM_T.n12 VSS 0.0374f
C693 IM_T.t16 VSS 0.0225f
C694 IM_T.n13 VSS 0.0374f
C695 IM_T.t0 VSS 0.0225f
C696 IM_T.n14 VSS 0.0374f
C697 IM_T.t3 VSS 0.0225f
C698 IM_T.n15 VSS 0.0374f
C699 IM_T.t26 VSS 0.0225f
C700 IM_T.n16 VSS 0.0378f
C701 IM_T.n17 VSS 0.0979f
C702 IM_T.t25 VSS 0.0504f
C703 IM_T.t21 VSS 0.0237f
C704 IM_T.n18 VSS 0.0467f
C705 IM_T.t8 VSS 0.0237f
C706 IM_T.n19 VSS 0.0383f
C707 IM_T.t9 VSS 0.0237f
C708 IM_T.n20 VSS 0.0383f
C709 IM_T.t12 VSS 0.0237f
C710 IM_T.n21 VSS 0.0383f
C711 IM_T.t20 VSS 0.0237f
C712 IM_T.n22 VSS 0.0383f
C713 IM_T.t28 VSS 0.0237f
C714 IM_T.n23 VSS 0.0383f
C715 IM_T.t7 VSS 0.0237f
C716 IM_T.n24 VSS 0.0383f
C717 IM_T.t22 VSS 0.0237f
C718 IM_T.n25 VSS 0.0383f
C719 IM_T.t13 VSS 0.0237f
C720 IM_T.n26 VSS 0.0383f
C721 IM_T.t5 VSS 0.0237f
C722 IM_T.n27 VSS 0.0383f
C723 IM_T.t29 VSS 0.0237f
C724 IM_T.n28 VSS 0.0383f
C725 IM_T.t14 VSS 0.0237f
C726 IM_T.n29 VSS 0.0383f
C727 IM_T.t6 VSS 0.0237f
C728 IM_T.n30 VSS 0.0383f
C729 IM_T.t31 VSS 0.0237f
C730 IM_T.n31 VSS 0.0383f
C731 IM_T.t23 VSS 0.0237f
C732 IM_T.n32 VSS 0.0436f
C733 IM_T.n33 VSS 0.0159f
C734 IM_T.n34 VSS 0.00131f
C735 OUT-.n0 VSS 0.0699f
C736 OUT-.t55 VSS 0.0197f
C737 OUT-.n1 VSS 0.0197f
C738 OUT-.n2 VSS 0.0689f
C739 OUT-.t30 VSS 0.0197f
C740 OUT-.n3 VSS 0.0197f
C741 OUT-.n4 VSS 0.0689f
C742 OUT-.t56 VSS 0.0197f
C743 OUT-.n5 VSS 0.0197f
C744 OUT-.n6 VSS 0.108f
C745 OUT-.n7 VSS 0.51f
C746 OUT-.n8 VSS 0.339f
C747 OUT-.t2 VSS 0.0197f
C748 OUT-.n9 VSS 0.0197f
C749 OUT-.n10 VSS 0.0689f
C750 OUT-.n11 VSS 0.27f
C751 OUT-.t4 VSS 0.0197f
C752 OUT-.n12 VSS 0.0197f
C753 OUT-.n13 VSS 0.0676f
C754 OUT-.t57 VSS 0.0197f
C755 OUT-.n14 VSS 0.0197f
C756 OUT-.n15 VSS 0.0686f
C757 OUT-.t6 VSS 0.0197f
C758 OUT-.n16 VSS 0.0197f
C759 OUT-.n17 VSS 0.0674f
C760 OUT-.t41 VSS 0.119f
C761 OUT-.n18 VSS 0.52f
C762 OUT-.n19 VSS 0.34f
C763 OUT-.n20 VSS 0.268f
C764 OUT-.n21 VSS 0.201f
C765 OUT-.n22 VSS 0.17f
C766 OUT-.n23 VSS 0.0699f
C767 OUT-.t3 VSS 0.0197f
C768 OUT-.n24 VSS 0.0197f
C769 OUT-.n25 VSS 0.0689f
C770 OUT-.t43 VSS 0.0197f
C771 OUT-.n26 VSS 0.0197f
C772 OUT-.n27 VSS 0.0689f
C773 OUT-.t5 VSS 0.0197f
C774 OUT-.n28 VSS 0.0197f
C775 OUT-.n29 VSS 0.108f
C776 OUT-.n30 VSS 0.51f
C777 OUT-.n31 VSS 0.339f
C778 OUT-.t21 VSS 0.0197f
C779 OUT-.n32 VSS 0.0197f
C780 OUT-.n33 VSS 0.0689f
C781 OUT-.n34 VSS 0.27f
C782 OUT-.t44 VSS 0.0197f
C783 OUT-.n35 VSS 0.0197f
C784 OUT-.n36 VSS 0.0676f
C785 OUT-.t33 VSS 0.0197f
C786 OUT-.n37 VSS 0.0197f
C787 OUT-.n38 VSS 0.0686f
C788 OUT-.t47 VSS 0.0197f
C789 OUT-.n39 VSS 0.0197f
C790 OUT-.n40 VSS 0.0674f
C791 OUT-.t12 VSS 0.119f
C792 OUT-.n41 VSS 0.52f
C793 OUT-.n42 VSS 0.34f
C794 OUT-.n43 VSS 0.268f
C795 OUT-.n44 VSS 0.201f
C796 OUT-.n45 VSS 0.17f
C797 OUT-.n46 VSS 0.0699f
C798 OUT-.t42 VSS 0.0197f
C799 OUT-.n47 VSS 0.0197f
C800 OUT-.n48 VSS 0.0689f
C801 OUT-.t16 VSS 0.0197f
C802 OUT-.n49 VSS 0.0197f
C803 OUT-.n50 VSS 0.0689f
C804 OUT-.t45 VSS 0.0197f
C805 OUT-.n51 VSS 0.0197f
C806 OUT-.n52 VSS 0.108f
C807 OUT-.n53 VSS 0.51f
C808 OUT-.n54 VSS 0.339f
C809 OUT-.t53 VSS 0.0197f
C810 OUT-.n55 VSS 0.0197f
C811 OUT-.n56 VSS 0.0689f
C812 OUT-.n57 VSS 0.27f
C813 OUT-.t17 VSS 0.0197f
C814 OUT-.n58 VSS 0.0197f
C815 OUT-.n59 VSS 0.0676f
C816 OUT-.t1 VSS 0.0197f
C817 OUT-.n60 VSS 0.0197f
C818 OUT-.n61 VSS 0.0686f
C819 OUT-.t20 VSS 0.0197f
C820 OUT-.n62 VSS 0.0197f
C821 OUT-.n63 VSS 0.0674f
C822 OUT-.t50 VSS 0.119f
C823 OUT-.n64 VSS 0.52f
C824 OUT-.n65 VSS 0.34f
C825 OUT-.n66 VSS 0.268f
C826 OUT-.n67 VSS 0.201f
C827 OUT-.n68 VSS 0.17f
C828 OUT-.n69 VSS 0.0699f
C829 OUT-.t15 VSS 0.0197f
C830 OUT-.n70 VSS 0.0197f
C831 OUT-.n71 VSS 0.0689f
C832 OUT-.t52 VSS 0.0197f
C833 OUT-.n72 VSS 0.0197f
C834 OUT-.n73 VSS 0.0689f
C835 OUT-.t18 VSS 0.0197f
C836 OUT-.n74 VSS 0.0197f
C837 OUT-.n75 VSS 0.108f
C838 OUT-.n76 VSS 0.51f
C839 OUT-.n77 VSS 0.339f
C840 OUT-.t26 VSS 0.0197f
C841 OUT-.n78 VSS 0.0197f
C842 OUT-.n79 VSS 0.0689f
C843 OUT-.n80 VSS 0.27f
C844 OUT-.t31 VSS 0.0197f
C845 OUT-.n81 VSS 0.0197f
C846 OUT-.n82 VSS 0.0676f
C847 OUT-.t19 VSS 0.0197f
C848 OUT-.n83 VSS 0.0197f
C849 OUT-.n84 VSS 0.0686f
C850 OUT-.t32 VSS 0.0197f
C851 OUT-.n85 VSS 0.0197f
C852 OUT-.n86 VSS 0.0674f
C853 OUT-.t59 VSS 0.119f
C854 OUT-.n87 VSS 0.52f
C855 OUT-.n88 VSS 0.34f
C856 OUT-.n89 VSS 0.268f
C857 OUT-.n90 VSS 0.201f
C858 OUT-.n91 VSS 0.418f
C859 OUT-.n92 VSS 0.6f
C860 OUT-.n93 VSS 0.548f
C861 OUT-.n94 VSS 0.642f
C862 OUT-.n95 VSS 0.0428f
C863 OUT-.n96 VSS 0.392f
C864 OUT.t34 VSS 0.0182f
C865 OUT.n0 VSS 0.0182f
C866 OUT.n1 VSS 0.0387f
C867 OUT.t16 VSS 0.0182f
C868 OUT.n2 VSS 0.0182f
C869 OUT.n3 VSS 0.0387f
C870 OUT.t52 VSS 0.0182f
C871 OUT.n4 VSS 0.0182f
C872 OUT.n5 VSS 0.0363f
C873 OUT.n6 VSS 0.139f
C874 OUT.t98 VSS 0.0182f
C875 OUT.n7 VSS 0.0182f
C876 OUT.n8 VSS 0.0363f
C877 OUT.n9 VSS 0.139f
C878 OUT.t49 VSS 0.0182f
C879 OUT.n10 VSS 0.0182f
C880 OUT.n11 VSS 0.0363f
C881 OUT.n12 VSS 0.139f
C882 OUT.t55 VSS 0.0182f
C883 OUT.n13 VSS 0.0182f
C884 OUT.n14 VSS 0.0394f
C885 OUT.t149 VSS 0.0182f
C886 OUT.n15 VSS 0.0182f
C887 OUT.n16 VSS 0.0408f
C888 OUT.t121 VSS 0.0182f
C889 OUT.n17 VSS 0.0182f
C890 OUT.n18 VSS 0.0394f
C891 OUT.t48 VSS 0.0182f
C892 OUT.n19 VSS 0.0182f
C893 OUT.n20 VSS 0.0408f
C894 OUT.n21 VSS 0.202f
C895 OUT.n22 VSS 0.259f
C896 OUT.t99 VSS 0.0182f
C897 OUT.n23 VSS 0.0182f
C898 OUT.n24 VSS 0.0363f
C899 OUT.n25 VSS 0.165f
C900 OUT.n26 VSS 0.222f
C901 OUT.t38 VSS 0.0182f
C902 OUT.n27 VSS 0.0182f
C903 OUT.n28 VSS 0.0394f
C904 OUT.t1 VSS 0.0182f
C905 OUT.n29 VSS 0.0182f
C906 OUT.n30 VSS 0.0408f
C907 OUT.t87 VSS 0.0182f
C908 OUT.n31 VSS 0.0182f
C909 OUT.n32 VSS 0.0394f
C910 OUT.t29 VSS 0.0182f
C911 OUT.n33 VSS 0.0182f
C912 OUT.n34 VSS 0.0408f
C913 OUT.n35 VSS 0.202f
C914 OUT.n36 VSS 0.259f
C915 OUT.t88 VSS 0.0182f
C916 OUT.n37 VSS 0.0182f
C917 OUT.n38 VSS 0.0363f
C918 OUT.t41 VSS 0.0182f
C919 OUT.n39 VSS 0.0182f
C920 OUT.n40 VSS 0.0363f
C921 OUT.n41 VSS 0.154f
C922 OUT.n42 VSS 0.165f
C923 OUT.n43 VSS 0.222f
C924 OUT.t50 VSS 0.0182f
C925 OUT.n44 VSS 0.0182f
C926 OUT.n45 VSS 0.0394f
C927 OUT.t102 VSS 0.0182f
C928 OUT.n46 VSS 0.0182f
C929 OUT.n47 VSS 0.0408f
C930 OUT.t123 VSS 0.0182f
C931 OUT.n48 VSS 0.0182f
C932 OUT.n49 VSS 0.0394f
C933 OUT.t45 VSS 0.0182f
C934 OUT.n50 VSS 0.0182f
C935 OUT.n51 VSS 0.0408f
C936 OUT.n52 VSS 0.202f
C937 OUT.n53 VSS 0.259f
C938 OUT.t94 VSS 0.0182f
C939 OUT.n54 VSS 0.0182f
C940 OUT.n55 VSS 0.0363f
C941 OUT.t54 VSS 0.0182f
C942 OUT.n56 VSS 0.0182f
C943 OUT.n57 VSS 0.0363f
C944 OUT.n58 VSS 0.154f
C945 OUT.n59 VSS 0.165f
C946 OUT.n60 VSS 0.222f
C947 OUT.t3 VSS 0.0182f
C948 OUT.n61 VSS 0.0182f
C949 OUT.n62 VSS 0.0408f
C950 OUT.t35 VSS 0.0182f
C951 OUT.n63 VSS 0.0182f
C952 OUT.n64 VSS 0.06f
C953 OUT.n65 VSS 0.413f
C954 OUT.t26 VSS 0.0182f
C955 OUT.n66 VSS 0.0182f
C956 OUT.n67 VSS 0.0408f
C957 OUT.t122 VSS 0.0182f
C958 OUT.n68 VSS 0.0182f
C959 OUT.n69 VSS 0.0597f
C960 OUT.n70 VSS 0.414f
C961 OUT.n71 VSS 0.253f
C962 OUT.t33 VSS 0.0182f
C963 OUT.n72 VSS 0.0182f
C964 OUT.n73 VSS 0.0363f
C965 OUT.t6 VSS 0.0182f
C966 OUT.n74 VSS 0.0182f
C967 OUT.n75 VSS 0.0363f
C968 OUT.t103 VSS 0.0182f
C969 OUT.n76 VSS 0.0182f
C970 OUT.n77 VSS 0.0394f
C971 OUT.t32 VSS 0.0182f
C972 OUT.n78 VSS 0.0182f
C973 OUT.n79 VSS 0.0408f
C974 OUT.t24 VSS 0.0182f
C975 OUT.n80 VSS 0.0182f
C976 OUT.n81 VSS 0.0394f
C977 OUT.t143 VSS 0.0182f
C978 OUT.n82 VSS 0.0182f
C979 OUT.n83 VSS 0.0407f
C980 OUT.n84 VSS 0.203f
C981 OUT.n85 VSS 0.26f
C982 OUT.t12 VSS 0.0182f
C983 OUT.n86 VSS 0.0182f
C984 OUT.n87 VSS 0.0363f
C985 OUT.n88 VSS 0.168f
C986 OUT.t44 VSS 0.0182f
C987 OUT.n89 VSS 0.0182f
C988 OUT.n90 VSS 0.0363f
C989 OUT.n91 VSS 0.154f
C990 OUT.n92 VSS 0.228f
C991 OUT.t42 VSS 0.0182f
C992 OUT.n93 VSS 0.0182f
C993 OUT.n94 VSS 0.0363f
C994 OUT.t141 VSS 0.0182f
C995 OUT.n95 VSS 0.0182f
C996 OUT.n96 VSS 0.0363f
C997 OUT.t155 VSS 0.0182f
C998 OUT.n97 VSS 0.0182f
C999 OUT.n98 VSS 0.0394f
C1000 OUT.t51 VSS 0.0182f
C1001 OUT.n99 VSS 0.0182f
C1002 OUT.n100 VSS 0.0408f
C1003 OUT.t43 VSS 0.0182f
C1004 OUT.n101 VSS 0.0182f
C1005 OUT.n102 VSS 0.0394f
C1006 OUT.t157 VSS 0.0182f
C1007 OUT.n103 VSS 0.0182f
C1008 OUT.n104 VSS 0.0407f
C1009 OUT.n105 VSS 0.203f
C1010 OUT.n106 VSS 0.26f
C1011 OUT.t156 VSS 0.0182f
C1012 OUT.n107 VSS 0.0182f
C1013 OUT.n108 VSS 0.0363f
C1014 OUT.n109 VSS 0.165f
C1015 OUT.t28 VSS 0.0182f
C1016 OUT.n110 VSS 0.0182f
C1017 OUT.n111 VSS 0.0363f
C1018 OUT.n112 VSS 0.154f
C1019 OUT.n113 VSS 0.228f
C1020 OUT.t25 VSS 0.0182f
C1021 OUT.n114 VSS 0.0182f
C1022 OUT.n115 VSS 0.0363f
C1023 OUT.t138 VSS 0.0182f
C1024 OUT.n116 VSS 0.0182f
C1025 OUT.n117 VSS 0.0363f
C1026 OUT.t150 VSS 0.0182f
C1027 OUT.n118 VSS 0.0182f
C1028 OUT.n119 VSS 0.0394f
C1029 OUT.t39 VSS 0.0182f
C1030 OUT.n120 VSS 0.0182f
C1031 OUT.n121 VSS 0.0408f
C1032 OUT.t27 VSS 0.0182f
C1033 OUT.n122 VSS 0.0182f
C1034 OUT.n123 VSS 0.0394f
C1035 OUT.t105 VSS 0.0182f
C1036 OUT.n124 VSS 0.0182f
C1037 OUT.n125 VSS 0.0407f
C1038 OUT.n126 VSS 0.203f
C1039 OUT.n127 VSS 0.26f
C1040 OUT.t104 VSS 0.0182f
C1041 OUT.n128 VSS 0.0182f
C1042 OUT.n129 VSS 0.0363f
C1043 OUT.n130 VSS 0.165f
C1044 OUT.t47 VSS 0.0182f
C1045 OUT.n131 VSS 0.0182f
C1046 OUT.n132 VSS 0.0363f
C1047 OUT.n133 VSS 0.154f
C1048 OUT.t158 VSS 0.0182f
C1049 OUT.n134 VSS 0.0182f
C1050 OUT.n135 VSS 0.0363f
C1051 OUT.n136 VSS 0.165f
C1052 OUT.n137 VSS 0.228f
C1053 OUT.t46 VSS 0.0182f
C1054 OUT.n138 VSS 0.0182f
C1055 OUT.n139 VSS 0.0363f
C1056 OUT.n140 VSS 0.165f
C1057 OUT.n141 VSS 0.221f
C1058 OUT.n142 VSS 0.154f
C1059 OUT.n143 VSS 0.165f
C1060 OUT.n144 VSS 0.221f
C1061 OUT.n145 VSS 0.154f
C1062 OUT.n146 VSS 0.165f
C1063 OUT.n147 VSS 0.221f
C1064 OUT.n148 VSS 0.154f
C1065 OUT.n149 VSS 0.168f
C1066 OUT.n150 VSS 0.243f
C1067 OUT.t15 VSS 0.0182f
C1068 OUT.n151 VSS 0.0182f
C1069 OUT.n152 VSS 0.0363f
C1070 OUT.t37 VSS 0.0182f
C1071 OUT.n153 VSS 0.0182f
C1072 OUT.n154 VSS 0.0363f
C1073 OUT.n155 VSS 0.154f
C1074 OUT.n156 VSS 0.168f
C1075 OUT.n157 VSS 0.244f
C1076 OUT.n158 VSS 0.253f
C1077 OUT.t30 VSS 0.0182f
C1078 OUT.n159 VSS 0.0182f
C1079 OUT.n160 VSS 0.0363f
C1080 OUT.n161 VSS 0.168f
C1081 OUT.t113 VSS 0.0182f
C1082 OUT.n162 VSS 0.0182f
C1083 OUT.n163 VSS 0.0363f
C1084 OUT.n164 VSS 0.154f
C1085 OUT.n165 VSS 0.228f
C1086 OUT.t36 VSS 0.0182f
C1087 OUT.n166 VSS 0.0182f
C1088 OUT.n167 VSS 0.0363f
C1089 OUT.n168 VSS 0.165f
C1090 OUT.t96 VSS 0.0182f
C1091 OUT.n169 VSS 0.0182f
C1092 OUT.n170 VSS 0.0363f
C1093 OUT.n171 VSS 0.154f
C1094 OUT.n172 VSS 0.228f
C1095 OUT.t53 VSS 0.0182f
C1096 OUT.n173 VSS 0.0182f
C1097 OUT.n174 VSS 0.0363f
C1098 OUT.n175 VSS 0.165f
C1099 OUT.t144 VSS 0.0182f
C1100 OUT.n176 VSS 0.0182f
C1101 OUT.n177 VSS 0.0363f
C1102 OUT.n178 VSS 0.154f
C1103 OUT.n179 VSS 0.228f
C1104 OUT.t40 VSS 0.0182f
C1105 OUT.n180 VSS 0.0182f
C1106 OUT.n181 VSS 0.0363f
C1107 OUT.n182 VSS 0.165f
C1108 OUT.t120 VSS 0.0182f
C1109 OUT.n183 VSS 0.0182f
C1110 OUT.n184 VSS 0.0363f
C1111 OUT.n185 VSS 0.139f
C1112 OUT.t31 VSS 0.0182f
C1113 OUT.n186 VSS 0.0182f
C1114 OUT.n187 VSS 0.0387f
C1115 OUT.t85 VSS 0.0182f
C1116 OUT.n188 VSS 0.0182f
C1117 OUT.n189 VSS 0.0567f
C1118 OUT.n190 VSS 0.414f
C1119 OUT.n191 VSS 0.247f
C1120 OUT.n192 VSS 0.25f
C1121 OUT.n193 VSS 0.249f
C1122 OUT.n194 VSS 0.248f
C1123 OUT.n195 VSS 0.266f
C1124 OUT.n196 VSS 1.22f
C1125 OUT.n197 VSS 0.103f
C1126 OUT.t125 VSS 0.0363f
C1127 OUT.n198 VSS 0.0363f
C1128 OUT.n199 VSS 0.0809f
C1129 OUT.t17 VSS 0.0363f
C1130 OUT.n200 VSS 0.0363f
C1131 OUT.n201 VSS 0.0783f
C1132 OUT.t116 VSS 0.0363f
C1133 OUT.n202 VSS 0.0363f
C1134 OUT.n203 VSS 0.0809f
C1135 OUT.t127 VSS 0.0363f
C1136 OUT.n204 VSS 0.0363f
C1137 OUT.n205 VSS 0.0783f
C1138 OUT.t129 VSS 0.0363f
C1139 OUT.n206 VSS 0.0363f
C1140 OUT.n207 VSS 0.0809f
C1141 OUT.t8 VSS 0.0363f
C1142 OUT.n208 VSS 0.0363f
C1143 OUT.n209 VSS 0.0783f
C1144 OUT.t10 VSS 0.0363f
C1145 OUT.n210 VSS 0.0363f
C1146 OUT.n211 VSS 0.0809f
C1147 OUT.t131 VSS 0.0363f
C1148 OUT.n212 VSS 0.0363f
C1149 OUT.n213 VSS 0.0783f
C1150 OUT.t11 VSS 0.0363f
C1151 OUT.n214 VSS 0.0363f
C1152 OUT.n215 VSS 0.0809f
C1153 OUT.t132 VSS 0.0363f
C1154 OUT.n216 VSS 0.0363f
C1155 OUT.n217 VSS 0.0783f
C1156 OUT.t133 VSS 0.0363f
C1157 OUT.n218 VSS 0.0363f
C1158 OUT.n219 VSS 0.0809f
C1159 OUT.t9 VSS 0.0363f
C1160 OUT.n220 VSS 0.0363f
C1161 OUT.n221 VSS 0.0783f
C1162 OUT.t134 VSS 0.0363f
C1163 OUT.n222 VSS 0.0363f
C1164 OUT.n223 VSS 0.0809f
C1165 OUT.t126 VSS 0.0363f
C1166 OUT.n224 VSS 0.0363f
C1167 OUT.n225 VSS 0.0783f
C1168 OUT.t92 VSS 0.0363f
C1169 OUT.n226 VSS 0.0363f
C1170 OUT.n227 VSS 0.0809f
C1171 OUT.t93 VSS 0.121f
C1172 OUT.n228 VSS 0.435f
C1173 OUT.n229 VSS 0.246f
C1174 OUT.n230 VSS 0.258f
C1175 OUT.n231 VSS 0.246f
C1176 OUT.n232 VSS 0.258f
C1177 OUT.n233 VSS 0.246f
C1178 OUT.n234 VSS 0.258f
C1179 OUT.n235 VSS 0.246f
C1180 OUT.n236 VSS 0.258f
C1181 OUT.n237 VSS 0.246f
C1182 OUT.n238 VSS 0.258f
C1183 OUT.n239 VSS 0.246f
C1184 OUT.n240 VSS 0.258f
C1185 OUT.n241 VSS 0.246f
C1186 OUT.n242 VSS 0.258f
C1187 OUT.n243 VSS 0.242f
C1188 QB.n0 VSS 0.02f
C1189 QB.t1 VSS 0.00819f
C1190 QB.n1 VSS 0.00819f
C1191 QB.n2 VSS 0.0207f
C1192 QB.n3 VSS 0.0971f
C1193 QB.t68 VSS 0.0123f
C1194 QB.t14 VSS 0.02f
C1195 QB.n4 VSS 0.0569f
C1196 QB.t67 VSS 0.0603f
C1197 QB.t65 VSS 0.0362f
C1198 QB.n5 VSS 0.103f
C1199 QB.t59 VSS 0.0362f
C1200 QB.n6 VSS 0.0684f
C1201 QB.t63 VSS 0.0376f
C1202 QB.n7 VSS 0.0701f
C1203 QB.t28 VSS 0.0376f
C1204 QB.n8 VSS 0.0701f
C1205 QB.t11 VSS 0.0362f
C1206 QB.n9 VSS 0.0684f
C1207 QB.t44 VSS 0.0362f
C1208 QB.n10 VSS 0.0684f
C1209 QB.t9 VSS 0.0376f
C1210 QB.n11 VSS 0.0701f
C1211 QB.t39 VSS 0.0376f
C1212 QB.n12 VSS 0.0701f
C1213 QB.t37 VSS 0.0362f
C1214 QB.n13 VSS 0.0684f
C1215 QB.t54 VSS 0.0362f
C1216 QB.n14 VSS 0.0684f
C1217 QB.t61 VSS 0.0376f
C1218 QB.n15 VSS 0.0701f
C1219 QB.t12 VSS 0.0376f
C1220 QB.n16 VSS 0.0701f
C1221 QB.t10 VSS 0.0362f
C1222 QB.n17 VSS 0.0684f
C1223 QB.t42 VSS 0.0362f
C1224 QB.n18 VSS 0.0755f
C1225 QB.t26 VSS 0.0313f
C1226 QB.n19 VSS 0.0976f
C1227 QB.t29 VSS 0.0603f
C1228 QB.t46 VSS 0.0362f
C1229 QB.n20 VSS 0.103f
C1230 QB.t45 VSS 0.0362f
C1231 QB.n21 VSS 0.0684f
C1232 QB.t23 VSS 0.0376f
C1233 QB.n22 VSS 0.0701f
C1234 QB.t57 VSS 0.0376f
C1235 QB.n23 VSS 0.0701f
C1236 QB.t64 VSS 0.0362f
C1237 QB.n24 VSS 0.0684f
C1238 QB.t30 VSS 0.0362f
C1239 QB.n25 VSS 0.0684f
C1240 QB.t34 VSS 0.0376f
C1241 QB.n26 VSS 0.0701f
C1242 QB.t4 VSS 0.0376f
C1243 QB.n27 VSS 0.0701f
C1244 QB.t24 VSS 0.0362f
C1245 QB.n28 VSS 0.0684f
C1246 QB.t40 VSS 0.0362f
C1247 QB.n29 VSS 0.0684f
C1248 QB.t20 VSS 0.0376f
C1249 QB.n30 VSS 0.0701f
C1250 QB.t38 VSS 0.0376f
C1251 QB.n31 VSS 0.0701f
C1252 QB.t62 VSS 0.0362f
C1253 QB.n32 VSS 0.0684f
C1254 QB.t27 VSS 0.0362f
C1255 QB.n33 VSS 0.0755f
C1256 QB.t55 VSS 0.0313f
C1257 QB.n34 VSS 0.0917f
C1258 QB.t58 VSS 0.0603f
C1259 QB.t13 VSS 0.0362f
C1260 QB.n35 VSS 0.103f
C1261 QB.t8 VSS 0.0362f
C1262 QB.n36 VSS 0.0684f
C1263 QB.t50 VSS 0.0376f
C1264 QB.n37 VSS 0.0701f
C1265 QB.t19 VSS 0.0376f
C1266 QB.n38 VSS 0.0701f
C1267 QB.t25 VSS 0.0362f
C1268 QB.n39 VSS 0.0684f
C1269 QB.t60 VSS 0.0362f
C1270 QB.n40 VSS 0.0684f
C1271 QB.t66 VSS 0.0376f
C1272 QB.n41 VSS 0.0701f
C1273 QB.t31 VSS 0.0376f
C1274 QB.n42 VSS 0.0701f
C1275 QB.t51 VSS 0.0362f
C1276 QB.n43 VSS 0.0684f
C1277 QB.t5 VSS 0.0362f
C1278 QB.n44 VSS 0.0684f
C1279 QB.t47 VSS 0.0376f
C1280 QB.n45 VSS 0.0701f
C1281 QB.t3 VSS 0.0376f
C1282 QB.n46 VSS 0.0701f
C1283 QB.t22 VSS 0.0362f
C1284 QB.n47 VSS 0.0684f
C1285 QB.t56 VSS 0.0362f
C1286 QB.n48 VSS 0.0755f
C1287 QB.t17 VSS 0.0313f
C1288 QB.n49 VSS 0.0917f
C1289 QB.t43 VSS 0.0603f
C1290 QB.t41 VSS 0.0362f
C1291 QB.n50 VSS 0.103f
C1292 QB.t33 VSS 0.0362f
C1293 QB.n51 VSS 0.0684f
C1294 QB.t36 VSS 0.0376f
C1295 QB.n52 VSS 0.0701f
C1296 QB.t6 VSS 0.0376f
C1297 QB.n53 VSS 0.0701f
C1298 QB.t52 VSS 0.0362f
C1299 QB.n54 VSS 0.0684f
C1300 QB.t21 VSS 0.0362f
C1301 QB.n55 VSS 0.0684f
C1302 QB.t48 VSS 0.0376f
C1303 QB.n56 VSS 0.0701f
C1304 QB.t16 VSS 0.0376f
C1305 QB.n57 VSS 0.0701f
C1306 QB.t15 VSS 0.0362f
C1307 QB.n58 VSS 0.0684f
C1308 QB.t32 VSS 0.0362f
C1309 QB.n59 VSS 0.0684f
C1310 QB.t35 VSS 0.0376f
C1311 QB.n60 VSS 0.0701f
C1312 QB.t53 VSS 0.0376f
C1313 QB.n61 VSS 0.0701f
C1314 QB.t49 VSS 0.0362f
C1315 QB.n62 VSS 0.0684f
C1316 QB.t18 VSS 0.0362f
C1317 QB.n63 VSS 0.0755f
C1318 QB.t7 VSS 0.0313f
C1319 QB.n64 VSS 0.101f
C1320 QB.n65 VSS 0.37f
C1321 QB.n66 VSS 0.16f
C1322 QB.n67 VSS 0.242f
C1323 QB.n68 VSS 0.247f
C1324 QB.n69 VSS 0.0254f
.ends

