magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2051 -2857 14313 58440
<< isosubstrate >>
rect -51 -51 12313 14512
<< nwell >>
rect 601 591 11661 6463
<< psubdiff >>
rect 684 13543 11578 13787
rect 684 12537 928 13543
rect 11334 12537 11578 13543
rect 684 12139 11578 12537
rect 684 11133 928 12139
rect 11334 11133 11578 12139
rect 684 10735 11578 11133
rect 684 9729 928 10735
rect 11334 9729 11578 10735
rect 684 9331 11578 9729
rect 684 8325 928 9331
rect 11334 8325 11578 9331
rect 684 8081 11578 8325
<< nsubdiff >>
rect 684 6136 11578 6380
rect 684 5130 928 6136
rect 11334 5130 11578 6136
rect 684 4732 11578 5130
rect 684 3726 928 4732
rect 11334 3726 11578 4732
rect 684 3328 11578 3726
rect 684 2322 928 3328
rect 11334 2322 11578 3328
rect 684 1924 11578 2322
rect 684 918 928 1924
rect 11334 918 11578 1924
rect 684 674 11578 918
<< metal1 >>
rect 511 13950 597 14418
rect 11665 13950 11751 14418
rect 695 13554 11567 13776
rect 695 12526 917 13554
rect 11345 12526 11567 13554
rect 695 12150 11567 12526
rect 695 11122 917 12150
rect 11345 11122 11567 12150
rect 695 10746 11567 11122
rect 695 9718 917 10746
rect 11345 9718 11567 10746
rect 695 9342 11567 9718
rect 695 8314 917 9342
rect 11345 8314 11567 9342
rect 695 8092 11567 8314
rect 511 7450 597 7918
rect 11665 7450 11751 7918
rect 511 6543 597 7011
rect 11665 6543 11751 7011
rect 695 6147 11567 6369
rect 695 5119 917 6147
rect 11345 5119 11567 6147
rect 695 4743 11567 5119
rect 695 3715 917 4743
rect 11345 3715 11567 4743
rect 695 3339 11567 3715
rect 695 2311 917 3339
rect 11345 2311 11567 3339
rect 695 1935 11567 2311
rect 695 907 917 1935
rect 11345 907 11567 1935
rect 695 685 11567 907
rect 511 43 597 511
rect 11665 43 11751 511
<< metal2 >>
rect -5 43 503 14905
rect 563 43 1071 14905
rect 1131 43 1639 14905
rect 1699 -857 2207 56440
rect 2267 43 2775 14905
rect 2835 -857 3343 56440
rect 3403 43 3911 14905
rect 3971 -857 4479 56440
rect 4539 43 5047 14905
rect 5107 -857 5615 56440
rect 5675 43 6101 14905
rect 6161 43 6587 14905
rect 6647 -857 7155 56440
rect 7215 43 7723 14905
rect 7783 -857 8291 56440
rect 8351 43 8859 14905
rect 8919 -857 9427 56440
rect 9487 43 9995 14905
rect 10055 -857 10563 56440
rect 10623 43 11131 14905
rect 11191 43 11699 14905
rect 11759 43 12267 14905
use M1_NWELL_CDNS_40661953145217  M1_NWELL_CDNS_40661953145217_0
timestamp 1713338890
transform 1 0 883 0 1 1421
box -128 -645 128 645
use M1_NWELL_CDNS_40661953145217  M1_NWELL_CDNS_40661953145217_1
timestamp 1713338890
transform 1 0 11379 0 1 1421
box -128 -645 128 645
use M1_NWELL_CDNS_40661953145217  M1_NWELL_CDNS_40661953145217_2
timestamp 1713338890
transform 1 0 883 0 1 2825
box -128 -645 128 645
use M1_NWELL_CDNS_40661953145217  M1_NWELL_CDNS_40661953145217_3
timestamp 1713338890
transform 1 0 11379 0 1 2825
box -128 -645 128 645
use M1_NWELL_CDNS_40661953145217  M1_NWELL_CDNS_40661953145217_4
timestamp 1713338890
transform 1 0 883 0 1 4229
box -128 -645 128 645
use M1_NWELL_CDNS_40661953145217  M1_NWELL_CDNS_40661953145217_5
timestamp 1713338890
transform 1 0 11379 0 1 4229
box -128 -645 128 645
use M1_NWELL_CDNS_40661953145217  M1_NWELL_CDNS_40661953145217_6
timestamp 1713338890
transform 1 0 883 0 1 5633
box -128 -645 128 645
use M1_NWELL_CDNS_40661953145217  M1_NWELL_CDNS_40661953145217_7
timestamp 1713338890
transform 1 0 11379 0 1 5633
box -128 -645 128 645
use M1_NWELL_CDNS_40661953145397  M1_NWELL_CDNS_40661953145397_0
timestamp 1713338890
transform 1 0 6131 0 1 2123
box -5345 -128 5345 128
use M1_NWELL_CDNS_40661953145397  M1_NWELL_CDNS_40661953145397_1
timestamp 1713338890
transform 1 0 6131 0 1 3527
box -5345 -128 5345 128
use M1_NWELL_CDNS_40661953145397  M1_NWELL_CDNS_40661953145397_2
timestamp 1713338890
transform 1 0 6131 0 1 4931
box -5345 -128 5345 128
use M1_NWELL_CDNS_40661953145398  M1_NWELL_CDNS_40661953145398_0
timestamp 1713338890
transform 1 0 6131 0 1 719
box -5486 -128 5486 128
use M1_NWELL_CDNS_40661953145398  M1_NWELL_CDNS_40661953145398_1
timestamp 1713338890
transform 1 0 6131 0 1 6335
box -5486 -128 5486 128
use M1_NWELL_CDNS_40661953145399  M1_NWELL_CDNS_40661953145399_0
timestamp 1713338890
transform 1 0 6131 0 1 873
box -5204 -128 5204 128
use M1_NWELL_CDNS_40661953145399  M1_NWELL_CDNS_40661953145399_1
timestamp 1713338890
transform 1 0 6131 0 1 1969
box -5204 -128 5204 128
use M1_NWELL_CDNS_40661953145399  M1_NWELL_CDNS_40661953145399_2
timestamp 1713338890
transform 1 0 6131 0 1 2277
box -5204 -128 5204 128
use M1_NWELL_CDNS_40661953145399  M1_NWELL_CDNS_40661953145399_3
timestamp 1713338890
transform 1 0 6131 0 1 3681
box -5204 -128 5204 128
use M1_NWELL_CDNS_40661953145399  M1_NWELL_CDNS_40661953145399_4
timestamp 1713338890
transform 1 0 6131 0 1 3373
box -5204 -128 5204 128
use M1_NWELL_CDNS_40661953145399  M1_NWELL_CDNS_40661953145399_5
timestamp 1713338890
transform 1 0 6131 0 1 4777
box -5204 -128 5204 128
use M1_NWELL_CDNS_40661953145399  M1_NWELL_CDNS_40661953145399_6
timestamp 1713338890
transform 1 0 6131 0 1 5085
box -5204 -128 5204 128
use M1_NWELL_CDNS_40661953145399  M1_NWELL_CDNS_40661953145399_7
timestamp 1713338890
transform 1 0 6131 0 1 6181
box -5204 -128 5204 128
use M1_NWELL_CDNS_40661953145400  M1_NWELL_CDNS_40661953145400_0
timestamp 1713338890
transform 1 0 729 0 1 3527
box -128 -2760 128 2760
use M1_NWELL_CDNS_40661953145400  M1_NWELL_CDNS_40661953145400_1
timestamp 1713338890
transform 1 0 11533 0 1 3527
box -128 -2760 128 2760
use M1_NWELL_CDNS_40661953145407  M1_NWELL_CDNS_40661953145407_0
timestamp 1713338890
transform 1 0 6131 0 1 7684
box -5628 -328 5628 328
use M1_NWELL_CDNS_40661953145407  M1_NWELL_CDNS_40661953145407_1
timestamp 1713338890
transform 1 0 6131 0 1 14184
box -5628 -328 5628 328
use M1_NWELL_CDNS_40661953145412  M1_NWELL_CDNS_40661953145412_0
timestamp 1713338890
transform 1 0 11985 0 1 10934
box -328 -3578 328 3578
use M1_NWELL_CDNS_40661953145412  M1_NWELL_CDNS_40661953145412_1
timestamp 1713338890
transform 1 0 277 0 1 10934
box -328 -3578 328 3578
use M1_PSUB_CDNS_6903358316550  M1_PSUB_CDNS_6903358316550_0
timestamp 1713338890
transform 1 0 6131 0 1 277
box -5545 -245 5545 245
use M1_PSUB_CDNS_6903358316550  M1_PSUB_CDNS_6903358316550_1
timestamp 1713338890
transform 1 0 6131 0 1 6777
box -5545 -245 5545 245
use M1_PSUB_CDNS_6903358316551  M1_PSUB_CDNS_6903358316551_0
timestamp 1713338890
transform 1 0 6131 0 1 9530
box -5262 -45 5262 45
use M1_PSUB_CDNS_6903358316551  M1_PSUB_CDNS_6903358316551_1
timestamp 1713338890
transform 1 0 6131 0 1 10934
box -5262 -45 5262 45
use M1_PSUB_CDNS_6903358316551  M1_PSUB_CDNS_6903358316551_2
timestamp 1713338890
transform 1 0 6131 0 1 12338
box -5262 -45 5262 45
use M1_PSUB_CDNS_6903358316552  M1_PSUB_CDNS_6903358316552_0
timestamp 1713338890
transform 1 0 6131 0 1 8280
box -5121 -45 5121 45
use M1_PSUB_CDNS_6903358316552  M1_PSUB_CDNS_6903358316552_1
timestamp 1713338890
transform 1 0 6131 0 1 9376
box -5121 -45 5121 45
use M1_PSUB_CDNS_6903358316552  M1_PSUB_CDNS_6903358316552_2
timestamp 1713338890
transform 1 0 6131 0 1 9684
box -5121 -45 5121 45
use M1_PSUB_CDNS_6903358316552  M1_PSUB_CDNS_6903358316552_3
timestamp 1713338890
transform 1 0 6131 0 1 10780
box -5121 -45 5121 45
use M1_PSUB_CDNS_6903358316552  M1_PSUB_CDNS_6903358316552_4
timestamp 1713338890
transform 1 0 6131 0 1 11088
box -5121 -45 5121 45
use M1_PSUB_CDNS_6903358316552  M1_PSUB_CDNS_6903358316552_5
timestamp 1713338890
transform 1 0 6131 0 1 12492
box -5121 -45 5121 45
use M1_PSUB_CDNS_6903358316552  M1_PSUB_CDNS_6903358316552_6
timestamp 1713338890
transform 1 0 6131 0 1 12184
box -5121 -45 5121 45
use M1_PSUB_CDNS_6903358316552  M1_PSUB_CDNS_6903358316552_7
timestamp 1713338890
transform 1 0 6131 0 1 13588
box -5121 -45 5121 45
use M1_PSUB_CDNS_6903358316553  M1_PSUB_CDNS_6903358316553_0
timestamp 1713338890
transform 1 0 6131 0 1 8126
box -5403 -45 5403 45
use M1_PSUB_CDNS_6903358316553  M1_PSUB_CDNS_6903358316553_1
timestamp 1713338890
transform 1 0 6131 0 1 13742
box -5403 -45 5403 45
use M1_PSUB_CDNS_6903358316555  M1_PSUB_CDNS_6903358316555_0
timestamp 1713338890
transform 1 0 11379 0 1 8828
box -45 -562 45 562
use M1_PSUB_CDNS_6903358316555  M1_PSUB_CDNS_6903358316555_1
timestamp 1713338890
transform 1 0 883 0 1 8828
box -45 -562 45 562
use M1_PSUB_CDNS_6903358316555  M1_PSUB_CDNS_6903358316555_2
timestamp 1713338890
transform 1 0 883 0 1 10232
box -45 -562 45 562
use M1_PSUB_CDNS_6903358316555  M1_PSUB_CDNS_6903358316555_3
timestamp 1713338890
transform 1 0 11379 0 1 10232
box -45 -562 45 562
use M1_PSUB_CDNS_6903358316555  M1_PSUB_CDNS_6903358316555_4
timestamp 1713338890
transform 1 0 883 0 1 11636
box -45 -562 45 562
use M1_PSUB_CDNS_6903358316555  M1_PSUB_CDNS_6903358316555_5
timestamp 1713338890
transform 1 0 11379 0 1 11636
box -45 -562 45 562
use M1_PSUB_CDNS_6903358316555  M1_PSUB_CDNS_6903358316555_6
timestamp 1713338890
transform 1 0 883 0 1 13040
box -45 -562 45 562
use M1_PSUB_CDNS_6903358316555  M1_PSUB_CDNS_6903358316555_7
timestamp 1713338890
transform 1 0 11379 0 1 13040
box -45 -562 45 562
use M1_PSUB_CDNS_6903358316556  M1_PSUB_CDNS_6903358316556_0
timestamp 1713338890
transform 1 0 11533 0 1 10934
box -45 -2677 45 2677
use M1_PSUB_CDNS_6903358316556  M1_PSUB_CDNS_6903358316556_1
timestamp 1713338890
transform 1 0 729 0 1 10934
box -45 -2677 45 2677
use M1_PSUB_CDNS_6903358316558  M1_PSUB_CDNS_6903358316558_0
timestamp 1713338890
transform 1 0 277 0 1 3527
box -245 -3495 245 3495
use M1_PSUB_CDNS_6903358316558  M1_PSUB_CDNS_6903358316558_1
timestamp 1713338890
transform 1 0 11985 0 1 3527
box -245 -3495 245 3495
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_0
timestamp 1713338890
transform 1 0 2521 0 1 2123
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_1
timestamp 1713338890
transform 1 0 4793 0 1 2123
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_2
timestamp 1713338890
transform -1 0 7469 0 1 2123
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_3
timestamp 1713338890
transform -1 0 9741 0 1 2123
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_4
timestamp 1713338890
transform 1 0 2521 0 1 3527
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_5
timestamp 1713338890
transform 1 0 4793 0 1 3527
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_6
timestamp 1713338890
transform -1 0 9741 0 1 3527
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_7
timestamp 1713338890
transform -1 0 7469 0 1 3527
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_8
timestamp 1713338890
transform 1 0 2521 0 1 4931
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_9
timestamp 1713338890
transform 1 0 4793 0 1 4931
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_10
timestamp 1713338890
transform -1 0 7469 0 1 4931
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_11
timestamp 1713338890
transform -1 0 9741 0 1 4931
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_12
timestamp 1713338890
transform 1 0 3657 0 1 9530
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_13
timestamp 1713338890
transform 1 0 1385 0 1 9530
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_14
timestamp 1713338890
transform -1 0 10877 0 1 9530
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_15
timestamp 1713338890
transform -1 0 8605 0 1 9530
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_16
timestamp 1713338890
transform 1 0 1385 0 1 10934
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_17
timestamp 1713338890
transform 1 0 3657 0 1 10934
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_18
timestamp 1713338890
transform -1 0 8605 0 1 10934
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_19
timestamp 1713338890
transform -1 0 10877 0 1 10934
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_20
timestamp 1713338890
transform 1 0 3657 0 1 12338
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_21
timestamp 1713338890
transform 1 0 1385 0 1 12338
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_22
timestamp 1713338890
transform -1 0 10877 0 1 12338
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_23
timestamp 1713338890
transform -1 0 8605 0 1 12338
box -254 -146 254 146
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_0
timestamp 1713338890
transform 1 0 1953 0 1 1421
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_1
timestamp 1713338890
transform 1 0 5361 0 1 1421
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_2
timestamp 1713338890
transform 1 0 3089 0 1 1421
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_3
timestamp 1713338890
transform 1 0 4225 0 1 1421
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_4
timestamp 1713338890
transform 1 0 10309 0 1 1421
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_5
timestamp 1713338890
transform 1 0 8037 0 1 1421
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_6
timestamp 1713338890
transform 1 0 9173 0 1 1421
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_7
timestamp 1713338890
transform 1 0 6901 0 1 1421
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_8
timestamp 1713338890
transform 1 0 4225 0 1 2825
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_9
timestamp 1713338890
transform 1 0 3089 0 1 2825
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_10
timestamp 1713338890
transform 1 0 5361 0 1 2825
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_11
timestamp 1713338890
transform 1 0 1953 0 1 2825
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_12
timestamp 1713338890
transform 1 0 9173 0 1 2825
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_13
timestamp 1713338890
transform 1 0 8037 0 1 2825
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_14
timestamp 1713338890
transform 1 0 10309 0 1 2825
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_15
timestamp 1713338890
transform 1 0 6901 0 1 2825
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_16
timestamp 1713338890
transform 1 0 3089 0 1 4229
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_17
timestamp 1713338890
transform 1 0 1953 0 1 4229
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_18
timestamp 1713338890
transform 1 0 5361 0 1 4229
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_19
timestamp 1713338890
transform 1 0 4225 0 1 4229
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_20
timestamp 1713338890
transform 1 0 6901 0 1 4229
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_21
timestamp 1713338890
transform 1 0 9173 0 1 4229
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_22
timestamp 1713338890
transform 1 0 8037 0 1 4229
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_23
timestamp 1713338890
transform 1 0 10309 0 1 4229
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_24
timestamp 1713338890
transform 1 0 4225 0 1 5633
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_25
timestamp 1713338890
transform 1 0 1953 0 1 5633
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_26
timestamp 1713338890
transform 1 0 5361 0 1 5633
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_27
timestamp 1713338890
transform 1 0 3089 0 1 5633
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_28
timestamp 1713338890
transform 1 0 6901 0 1 5633
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_29
timestamp 1713338890
transform 1 0 10309 0 1 5633
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_30
timestamp 1713338890
transform 1 0 8037 0 1 5633
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_31
timestamp 1713338890
transform 1 0 9173 0 1 5633
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_32
timestamp 1713338890
transform 1 0 3089 0 1 8828
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_33
timestamp 1713338890
transform 1 0 5361 0 1 8828
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_34
timestamp 1713338890
transform 1 0 1953 0 1 8828
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_35
timestamp 1713338890
transform 1 0 4225 0 1 8828
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_36
timestamp 1713338890
transform 1 0 6901 0 1 8828
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_37
timestamp 1713338890
transform 1 0 10309 0 1 8828
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_38
timestamp 1713338890
transform 1 0 8037 0 1 8828
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_39
timestamp 1713338890
transform 1 0 9173 0 1 8828
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_40
timestamp 1713338890
transform 1 0 4225 0 1 10232
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_41
timestamp 1713338890
transform 1 0 3089 0 1 10232
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_42
timestamp 1713338890
transform 1 0 5361 0 1 10232
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_43
timestamp 1713338890
transform 1 0 1953 0 1 10232
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_44
timestamp 1713338890
transform 1 0 9173 0 1 10232
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_45
timestamp 1713338890
transform 1 0 8037 0 1 10232
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_46
timestamp 1713338890
transform 1 0 10309 0 1 10232
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_47
timestamp 1713338890
transform 1 0 6901 0 1 10232
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_48
timestamp 1713338890
transform 1 0 4225 0 1 11636
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_49
timestamp 1713338890
transform 1 0 3089 0 1 11636
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_50
timestamp 1713338890
transform 1 0 5361 0 1 11636
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_51
timestamp 1713338890
transform 1 0 1953 0 1 11636
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_52
timestamp 1713338890
transform 1 0 9173 0 1 11636
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_53
timestamp 1713338890
transform 1 0 8037 0 1 11636
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_54
timestamp 1713338890
transform 1 0 10309 0 1 11636
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_55
timestamp 1713338890
transform 1 0 6901 0 1 11636
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_56
timestamp 1713338890
transform 1 0 4225 0 1 13040
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_57
timestamp 1713338890
transform 1 0 3089 0 1 13040
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_58
timestamp 1713338890
transform 1 0 5361 0 1 13040
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_59
timestamp 1713338890
transform 1 0 1953 0 1 13040
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_60
timestamp 1713338890
transform 1 0 9173 0 1 13040
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_61
timestamp 1713338890
transform 1 0 10309 0 1 13040
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_62
timestamp 1713338890
transform 1 0 6901 0 1 13040
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_63
timestamp 1713338890
transform 1 0 8037 0 1 13040
box -224 -286 224 286
use M2_M1_CDNS_6903358316540  M2_M1_CDNS_6903358316540_0
timestamp 1713338890
transform 1 0 5888 0 1 9530
box -200 -146 200 146
use M2_M1_CDNS_6903358316540  M2_M1_CDNS_6903358316540_1
timestamp 1713338890
transform -1 0 6374 0 1 9530
box -200 -146 200 146
use M2_M1_CDNS_6903358316540  M2_M1_CDNS_6903358316540_2
timestamp 1713338890
transform 1 0 5888 0 1 10934
box -200 -146 200 146
use M2_M1_CDNS_6903358316540  M2_M1_CDNS_6903358316540_3
timestamp 1713338890
transform -1 0 6374 0 1 10934
box -200 -146 200 146
use M2_M1_CDNS_6903358316540  M2_M1_CDNS_6903358316540_4
timestamp 1713338890
transform 1 0 5888 0 1 12338
box -200 -146 200 146
use M2_M1_CDNS_6903358316540  M2_M1_CDNS_6903358316540_5
timestamp 1713338890
transform -1 0 6374 0 1 12338
box -200 -146 200 146
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_0
timestamp 1713338890
transform 1 0 2521 0 1 796
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_1
timestamp 1713338890
transform 1 0 4793 0 1 796
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_2
timestamp 1713338890
transform -1 0 7469 0 1 796
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_3
timestamp 1713338890
transform -1 0 9741 0 1 796
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_4
timestamp 1713338890
transform 1 0 4793 0 1 6258
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_5
timestamp 1713338890
transform 1 0 2521 0 1 6258
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_6
timestamp 1713338890
transform -1 0 9741 0 1 6258
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_7
timestamp 1713338890
transform -1 0 7469 0 1 6258
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_8
timestamp 1713338890
transform -1 0 8605 0 1 8203
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_9
timestamp 1713338890
transform -1 0 10877 0 1 8203
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_10
timestamp 1713338890
transform 1 0 3657 0 1 8203
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_11
timestamp 1713338890
transform 1 0 1385 0 1 8203
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_12
timestamp 1713338890
transform -1 0 10877 0 1 13665
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_13
timestamp 1713338890
transform -1 0 8605 0 1 13665
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_14
timestamp 1713338890
transform 1 0 3657 0 1 13665
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_15
timestamp 1713338890
transform 1 0 1385 0 1 13665
box -254 -92 254 92
use M2_M1_CDNS_6903358316547  M2_M1_CDNS_6903358316547_0
timestamp 1713338890
transform -1 0 6374 0 1 8203
box -200 -92 200 92
use M2_M1_CDNS_6903358316547  M2_M1_CDNS_6903358316547_1
timestamp 1713338890
transform 1 0 5888 0 1 8203
box -200 -92 200 92
use M2_M1_CDNS_6903358316547  M2_M1_CDNS_6903358316547_2
timestamp 1713338890
transform -1 0 6374 0 1 13665
box -200 -92 200 92
use M2_M1_CDNS_6903358316547  M2_M1_CDNS_6903358316547_3
timestamp 1713338890
transform 1 0 5888 0 1 13665
box -200 -92 200 92
use M2_M1_CDNS_6903358316554  M2_M1_CDNS_6903358316554_0
timestamp 1713338890
transform 1 0 1385 0 1 277
box -224 -224 224 224
use M2_M1_CDNS_6903358316554  M2_M1_CDNS_6903358316554_1
timestamp 1713338890
transform 1 0 3657 0 1 277
box -224 -224 224 224
use M2_M1_CDNS_6903358316554  M2_M1_CDNS_6903358316554_2
timestamp 1713338890
transform -1 0 10877 0 1 277
box -224 -224 224 224
use M2_M1_CDNS_6903358316554  M2_M1_CDNS_6903358316554_3
timestamp 1713338890
transform -1 0 8605 0 1 277
box -224 -224 224 224
use M2_M1_CDNS_6903358316554  M2_M1_CDNS_6903358316554_4
timestamp 1713338890
transform 1 0 1385 0 1 6777
box -224 -224 224 224
use M2_M1_CDNS_6903358316554  M2_M1_CDNS_6903358316554_5
timestamp 1713338890
transform 1 0 3657 0 1 6777
box -224 -224 224 224
use M2_M1_CDNS_6903358316554  M2_M1_CDNS_6903358316554_6
timestamp 1713338890
transform -1 0 10877 0 1 6777
box -224 -224 224 224
use M2_M1_CDNS_6903358316554  M2_M1_CDNS_6903358316554_7
timestamp 1713338890
transform -1 0 8605 0 1 6777
box -224 -224 224 224
use M2_M1_CDNS_6903358316554  M2_M1_CDNS_6903358316554_8
timestamp 1713338890
transform -1 0 11445 0 1 7684
box -224 -224 224 224
use M2_M1_CDNS_6903358316554  M2_M1_CDNS_6903358316554_9
timestamp 1713338890
transform -1 0 9741 0 1 7684
box -224 -224 224 224
use M2_M1_CDNS_6903358316554  M2_M1_CDNS_6903358316554_10
timestamp 1713338890
transform -1 0 7469 0 1 7684
box -224 -224 224 224
use M2_M1_CDNS_6903358316554  M2_M1_CDNS_6903358316554_11
timestamp 1713338890
transform 1 0 4793 0 1 7684
box -224 -224 224 224
use M2_M1_CDNS_6903358316554  M2_M1_CDNS_6903358316554_12
timestamp 1713338890
transform 1 0 2521 0 1 7684
box -224 -224 224 224
use M2_M1_CDNS_6903358316554  M2_M1_CDNS_6903358316554_13
timestamp 1713338890
transform 1 0 817 0 1 7684
box -224 -224 224 224
use M2_M1_CDNS_6903358316554  M2_M1_CDNS_6903358316554_14
timestamp 1713338890
transform -1 0 9741 0 1 14184
box -224 -224 224 224
use M2_M1_CDNS_6903358316554  M2_M1_CDNS_6903358316554_15
timestamp 1713338890
transform -1 0 11445 0 1 14184
box -224 -224 224 224
use M2_M1_CDNS_6903358316554  M2_M1_CDNS_6903358316554_16
timestamp 1713338890
transform -1 0 7469 0 1 14184
box -224 -224 224 224
use M2_M1_CDNS_6903358316554  M2_M1_CDNS_6903358316554_17
timestamp 1713338890
transform 1 0 4793 0 1 14184
box -224 -224 224 224
use M2_M1_CDNS_6903358316554  M2_M1_CDNS_6903358316554_18
timestamp 1713338890
transform 1 0 2521 0 1 14184
box -224 -224 224 224
use M2_M1_CDNS_6903358316554  M2_M1_CDNS_6903358316554_19
timestamp 1713338890
transform 1 0 817 0 1 14184
box -224 -224 224 224
use M2_M1_CDNS_6903358316557  M2_M1_CDNS_6903358316557_0
timestamp 1713338890
transform 1 0 5888 0 1 277
box -162 -224 162 224
use M2_M1_CDNS_6903358316557  M2_M1_CDNS_6903358316557_1
timestamp 1713338890
transform -1 0 6374 0 1 277
box -162 -224 162 224
use M2_M1_CDNS_6903358316557  M2_M1_CDNS_6903358316557_2
timestamp 1713338890
transform 1 0 5888 0 1 6777
box -162 -224 162 224
use M2_M1_CDNS_6903358316557  M2_M1_CDNS_6903358316557_3
timestamp 1713338890
transform -1 0 6374 0 1 6777
box -162 -224 162 224
use M2_M1_CDNS_6903358316559  M2_M1_CDNS_6903358316559_0
timestamp 1713338890
transform 1 0 323 0 1 3527
box -146 -3440 146 3440
use M2_M1_CDNS_6903358316559  M2_M1_CDNS_6903358316559_1
timestamp 1713338890
transform -1 0 11939 0 1 3527
box -146 -3440 146 3440
use M2_M1_CDNS_6903358316560  M2_M1_CDNS_6903358316560_0
timestamp 1713338890
transform 1 0 817 0 1 3527
box -92 -2792 92 2792
use M2_M1_CDNS_6903358316560  M2_M1_CDNS_6903358316560_1
timestamp 1713338890
transform -1 0 11445 0 1 3527
box -92 -2792 92 2792
use M2_M1_CDNS_6903358316561  M2_M1_CDNS_6903358316561_0
timestamp 1713338890
transform 1 0 11939 0 1 3527
box -146 -3332 146 3332
use np_6p0_CDNS_4066195314553  np_6p0_CDNS_4066195314553_0
timestamp 1713338890
transform 0 -1 11131 1 0 8528
box 0 0 600 10000
use np_6p0_CDNS_4066195314553  np_6p0_CDNS_4066195314553_1
timestamp 1713338890
transform 0 -1 11131 1 0 9932
box 0 0 600 10000
use np_6p0_CDNS_4066195314553  np_6p0_CDNS_4066195314553_2
timestamp 1713338890
transform 0 -1 11131 1 0 11336
box 0 0 600 10000
use np_6p0_CDNS_4066195314553  np_6p0_CDNS_4066195314553_3
timestamp 1713338890
transform 0 -1 11131 1 0 12740
box 0 0 600 10000
use pn_6p0_CDNS_4066195314552  pn_6p0_CDNS_4066195314552_0
timestamp 1713338890
transform 0 -1 11131 1 0 1121
box -120 -120 720 10120
use pn_6p0_CDNS_4066195314552  pn_6p0_CDNS_4066195314552_1
timestamp 1713338890
transform 0 -1 11131 1 0 2525
box -120 -120 720 10120
use pn_6p0_CDNS_4066195314552  pn_6p0_CDNS_4066195314552_2
timestamp 1713338890
transform 0 -1 11131 1 0 3929
box -120 -120 720 10120
use pn_6p0_CDNS_4066195314552  pn_6p0_CDNS_4066195314552_3
timestamp 1713338890
transform 0 -1 11131 1 0 5333
box -120 -120 720 10120
<< end >>
