magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1000 -994 2040 5126
use pmos_6p0_esd_40  pmos_6p0_esd_40_0
timestamp 1713338890
transform 1 0 0 0 1 0
box 0 6 598 4126
use pmos_6p0_esd_40  pmos_6p0_esd_40_1
timestamp 1713338890
transform -1 0 1040 0 1 0
box 0 6 598 4126
<< end >>
