magic
tech gf180mcuC
magscale 1 10
timestamp 1694939250
<< pwell >>
rect -820 -536 820 536
<< nmos >>
rect -708 68 -508 468
rect -404 68 -204 468
rect -100 68 100 468
rect 204 68 404 468
rect 508 68 708 468
rect -708 -468 -508 -68
rect -404 -468 -204 -68
rect -100 -468 100 -68
rect 204 -468 404 -68
rect 508 -468 708 -68
<< ndiff >>
rect -796 455 -708 468
rect -796 81 -783 455
rect -737 81 -708 455
rect -796 68 -708 81
rect -508 455 -404 468
rect -508 81 -479 455
rect -433 81 -404 455
rect -508 68 -404 81
rect -204 455 -100 468
rect -204 81 -175 455
rect -129 81 -100 455
rect -204 68 -100 81
rect 100 455 204 468
rect 100 81 129 455
rect 175 81 204 455
rect 100 68 204 81
rect 404 455 508 468
rect 404 81 433 455
rect 479 81 508 455
rect 404 68 508 81
rect 708 455 796 468
rect 708 81 737 455
rect 783 81 796 455
rect 708 68 796 81
rect -796 -81 -708 -68
rect -796 -455 -783 -81
rect -737 -455 -708 -81
rect -796 -468 -708 -455
rect -508 -81 -404 -68
rect -508 -455 -479 -81
rect -433 -455 -404 -81
rect -508 -468 -404 -455
rect -204 -81 -100 -68
rect -204 -455 -175 -81
rect -129 -455 -100 -81
rect -204 -468 -100 -455
rect 100 -81 204 -68
rect 100 -455 129 -81
rect 175 -455 204 -81
rect 100 -468 204 -455
rect 404 -81 508 -68
rect 404 -455 433 -81
rect 479 -455 508 -81
rect 404 -468 508 -455
rect 708 -81 796 -68
rect 708 -455 737 -81
rect 783 -455 796 -81
rect 708 -468 796 -455
<< ndiffc >>
rect -783 81 -737 455
rect -479 81 -433 455
rect -175 81 -129 455
rect 129 81 175 455
rect 433 81 479 455
rect 737 81 783 455
rect -783 -455 -737 -81
rect -479 -455 -433 -81
rect -175 -455 -129 -81
rect 129 -455 175 -81
rect 433 -455 479 -81
rect 737 -455 783 -81
<< polysilicon >>
rect -708 468 -508 512
rect -404 468 -204 512
rect -100 468 100 512
rect 204 468 404 512
rect 508 468 708 512
rect -708 24 -508 68
rect -404 24 -204 68
rect -100 24 100 68
rect 204 24 404 68
rect 508 24 708 68
rect -708 -68 -508 -24
rect -404 -68 -204 -24
rect -100 -68 100 -24
rect 204 -68 404 -24
rect 508 -68 708 -24
rect -708 -512 -508 -468
rect -404 -512 -204 -468
rect -100 -512 100 -468
rect 204 -512 404 -468
rect 508 -512 708 -468
<< metal1 >>
rect -783 455 -737 466
rect -783 70 -737 81
rect -479 455 -433 466
rect -479 70 -433 81
rect -175 455 -129 466
rect -175 70 -129 81
rect 129 455 175 466
rect 129 70 175 81
rect 433 455 479 466
rect 433 70 479 81
rect 737 455 783 466
rect 737 70 783 81
rect -783 -81 -737 -70
rect -783 -466 -737 -455
rect -479 -81 -433 -70
rect -479 -466 -433 -455
rect -175 -81 -129 -70
rect -175 -466 -129 -455
rect 129 -81 175 -70
rect 129 -466 175 -455
rect 433 -81 479 -70
rect 433 -466 479 -455
rect 737 -81 783 -70
rect 737 -466 783 -455
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 2 l 1 m 2 nf 5 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
