magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1298 -1019 1298 1019
<< metal2 >>
rect -298 14 298 19
rect -298 -14 -293 14
rect -265 -14 -231 14
rect -203 -14 -169 14
rect -141 -14 -107 14
rect -79 -14 -45 14
rect -17 -14 17 14
rect 45 -14 79 14
rect 107 -14 141 14
rect 169 -14 203 14
rect 231 -14 265 14
rect 293 -14 298 14
rect -298 -19 298 -14
<< via2 >>
rect -293 -14 -265 14
rect -231 -14 -203 14
rect -169 -14 -141 14
rect -107 -14 -79 14
rect -45 -14 -17 14
rect 17 -14 45 14
rect 79 -14 107 14
rect 141 -14 169 14
rect 203 -14 231 14
rect 265 -14 293 14
<< metal3 >>
rect -298 14 298 19
rect -298 -14 -293 14
rect -265 -14 -231 14
rect -203 -14 -169 14
rect -141 -14 -107 14
rect -79 -14 -45 14
rect -17 -14 17 14
rect 45 -14 79 14
rect 107 -14 141 14
rect 169 -14 203 14
rect 231 -14 265 14
rect 293 -14 298 14
rect -298 -19 298 -14
<< end >>
