magic
tech gf180mcuC
magscale 1 10
timestamp 1692959041
<< error_s >>
rect -3685 -2473 -3529 -2459
rect -3685 -2505 -3668 -2473
rect -3639 -2551 -3622 -2505
rect -3639 -2569 -3575 -2551
rect -3546 -2569 -3529 -2473
rect -3681 -2707 -3525 -2693
rect -3681 -2739 -3664 -2707
rect -3635 -2785 -3618 -2739
rect -3635 -2803 -3571 -2785
rect -3542 -2803 -3525 -2707
rect -1768 -2723 -1620 -2698
rect -1768 -2743 -1666 -2723
rect -1754 -2744 -1666 -2743
rect -1754 -2747 -1722 -2744
rect -1708 -2747 -1697 -2744
rect -1719 -2753 -1676 -2747
rect -1722 -2754 -1676 -2753
rect -1722 -2800 -1666 -2754
rect -1642 -2800 -1620 -2723
rect -2649 -2953 -2481 -2911
rect -2008 -2952 -1840 -2911
rect -2649 -2967 -2607 -2953
rect -2524 -2965 -2481 -2953
rect -2524 -2967 -2491 -2965
rect -1998 -2967 -1965 -2952
rect -1882 -2967 -1840 -2952
rect -2593 -2969 -2547 -2967
rect -2537 -2969 -2491 -2967
rect -2593 -3023 -2491 -2969
rect -1952 -2980 -1906 -2967
rect -1896 -2980 -1840 -2967
rect -1952 -3023 -1840 -2980
rect -2808 -3105 -2640 -3063
rect -2808 -3116 -2766 -3105
rect -2798 -3119 -2766 -3116
rect -2683 -3116 -2640 -3105
rect -2489 -3104 -2321 -3062
rect -2489 -3116 -2447 -3104
rect -2683 -3119 -2650 -3116
rect -2479 -3118 -2447 -3116
rect -2364 -3116 -2321 -3104
rect -2167 -3104 -1999 -3062
rect -2167 -3116 -2125 -3104
rect -2364 -3118 -2331 -3116
rect -2157 -3118 -2125 -3116
rect -2042 -3116 -1999 -3104
rect -1852 -3104 -1684 -3062
rect -1852 -3116 -1810 -3104
rect -2042 -3118 -2009 -3116
rect -1842 -3118 -1810 -3116
rect -1727 -3118 -1684 -3104
rect -2752 -3121 -2706 -3119
rect -2696 -3121 -2650 -3119
rect -2752 -3175 -2650 -3121
rect -2433 -3121 -2387 -3118
rect -2377 -3121 -2331 -3118
rect -2433 -3174 -2331 -3121
rect -2111 -3121 -2065 -3118
rect -2055 -3121 -2009 -3118
rect -2111 -3174 -2009 -3121
rect -1796 -3130 -1750 -3118
rect -1740 -3130 -1684 -3118
rect -1796 -3174 -1684 -3130
rect -3130 -3259 -2801 -3218
rect -3130 -3260 -2927 -3259
rect -3130 -3274 -3088 -3260
rect -3004 -3272 -2927 -3260
rect -3004 -3274 -2972 -3272
rect -2959 -3274 -2927 -3272
rect -2843 -3272 -2801 -3259
rect -2330 -3260 -2160 -3218
rect -2330 -3272 -2288 -3260
rect -2843 -3274 -2811 -3272
rect -2320 -3274 -2288 -3272
rect -2202 -3272 -2160 -3260
rect -1689 -3259 -1361 -3218
rect -1689 -3272 -1647 -3259
rect -2202 -3274 -2170 -3272
rect -1679 -3274 -1647 -3272
rect -1563 -3260 -1361 -3259
rect -1563 -3272 -1487 -3260
rect -1563 -3274 -1531 -3272
rect -1519 -3274 -1487 -3272
rect -1403 -3274 -1361 -3260
rect -3074 -3276 -3028 -3274
rect -3018 -3276 -2972 -3274
rect -3074 -3330 -2972 -3276
rect -2913 -3276 -2867 -3274
rect -2857 -3276 -2811 -3274
rect -2913 -3330 -2811 -3276
rect -2274 -3276 -2228 -3274
rect -2216 -3276 -2170 -3274
rect -2274 -3330 -2170 -3276
rect -1633 -3276 -1587 -3274
rect -1577 -3276 -1531 -3274
rect -1633 -3330 -1531 -3276
rect -1473 -3288 -1427 -3274
rect -1417 -3288 -1361 -3274
rect -1473 -3330 -1361 -3288
rect -2877 -3561 -2729 -3515
rect -2852 -3580 -2806 -3561
rect -2775 -3563 -2729 -3561
rect -2794 -3573 -2783 -3569
rect -2775 -3573 -2737 -3563
rect -2797 -3580 -2737 -3573
rect -2831 -3617 -2785 -3580
rect -2783 -3617 -2737 -3580
rect -2649 -3806 -2481 -3766
rect -2649 -3808 -2491 -3806
rect -2649 -3822 -2607 -3808
rect -2524 -3822 -2491 -3808
rect -2008 -3809 -1840 -3766
rect -2008 -3820 -1965 -3809
rect -1998 -3822 -1965 -3820
rect -1882 -3822 -1840 -3809
rect -2593 -3834 -2547 -3822
rect -2537 -3834 -2491 -3822
rect -2593 -3878 -2491 -3834
rect -1952 -3835 -1906 -3822
rect -1896 -3835 -1840 -3822
rect -1952 -3878 -1840 -3835
rect -2809 -3961 -2641 -3919
rect -2809 -3973 -2767 -3961
rect -2799 -3975 -2767 -3973
rect -2684 -3973 -2641 -3961
rect -2491 -3960 -2317 -3915
rect -2491 -3971 -2446 -3960
rect -2363 -3971 -2317 -3960
rect -2684 -3975 -2651 -3973
rect -2753 -3978 -2707 -3975
rect -2697 -3978 -2651 -3975
rect -2753 -4031 -2651 -3978
rect -2435 -3978 -2389 -3971
rect -2373 -3973 -2317 -3971
rect -2168 -3960 -2000 -3918
rect -2168 -3973 -2126 -3960
rect -2373 -3978 -2327 -3973
rect -2158 -3974 -2126 -3973
rect -2043 -3973 -2000 -3960
rect -1848 -3961 -1680 -3919
rect -1848 -3973 -1806 -3961
rect -2043 -3974 -2010 -3973
rect -2435 -4033 -2327 -3978
rect -2112 -3978 -2066 -3974
rect -2056 -3978 -2010 -3974
rect -1838 -3975 -1806 -3973
rect -1723 -3975 -1680 -3961
rect -2112 -4030 -2010 -3978
rect -1792 -3987 -1746 -3975
rect -1736 -3987 -1680 -3975
rect -1792 -4031 -1680 -3987
rect -3130 -4119 -2801 -4078
rect -3130 -4120 -2927 -4119
rect -3130 -4134 -3088 -4120
rect -3004 -4132 -2927 -4120
rect -3004 -4134 -2972 -4132
rect -2959 -4134 -2927 -4132
rect -2843 -4132 -2801 -4119
rect -2330 -4120 -2160 -4078
rect -2330 -4132 -2288 -4120
rect -2843 -4134 -2811 -4132
rect -2320 -4134 -2288 -4132
rect -2202 -4132 -2160 -4120
rect -1689 -4119 -1361 -4078
rect -1689 -4132 -1647 -4119
rect -2202 -4134 -2170 -4132
rect -1679 -4134 -1647 -4132
rect -1563 -4120 -1361 -4119
rect -1563 -4132 -1487 -4120
rect -1563 -4134 -1531 -4132
rect -1519 -4134 -1487 -4132
rect -1403 -4134 -1361 -4120
rect -3074 -4136 -3028 -4134
rect -3018 -4136 -2972 -4134
rect -3074 -4190 -2972 -4136
rect -2913 -4136 -2867 -4134
rect -2857 -4136 -2811 -4134
rect -2913 -4190 -2811 -4136
rect -2274 -4136 -2228 -4134
rect -2216 -4136 -2170 -4134
rect -2274 -4190 -2170 -4136
rect -1633 -4136 -1587 -4134
rect -1577 -4136 -1531 -4134
rect -1633 -4190 -1531 -4136
rect -1473 -4148 -1427 -4134
rect -1417 -4148 -1361 -4134
rect -1473 -4190 -1361 -4148
rect -1772 -4386 -1618 -4358
rect -1772 -4404 -1745 -4386
rect -1726 -4415 -1699 -4404
rect -1726 -4437 -1699 -4425
rect -1726 -4465 -1664 -4437
rect -1644 -4465 -1618 -4386
rect -2649 -4666 -2481 -4626
rect -2649 -4668 -2491 -4666
rect -2649 -4682 -2607 -4668
rect -2524 -4682 -2491 -4668
rect -2008 -4669 -1840 -4626
rect -2008 -4680 -1965 -4669
rect -1998 -4682 -1965 -4680
rect -1882 -4682 -1840 -4669
rect -2593 -4694 -2547 -4682
rect -2537 -4694 -2491 -4682
rect -2593 -4738 -2491 -4694
rect -1952 -4695 -1906 -4682
rect -1896 -4695 -1840 -4682
rect -1952 -4738 -1840 -4695
rect -2809 -4825 -2641 -4783
rect -2809 -4837 -2767 -4825
rect -2799 -4839 -2767 -4837
rect -2684 -4837 -2641 -4825
rect -2489 -4826 -2321 -4784
rect -2489 -4837 -2447 -4826
rect -2684 -4839 -2651 -4837
rect -2753 -4842 -2707 -4839
rect -2697 -4842 -2651 -4839
rect -2479 -4840 -2447 -4837
rect -2364 -4837 -2321 -4826
rect -2169 -4824 -2001 -4782
rect -2169 -4837 -2127 -4824
rect -2364 -4840 -2331 -4837
rect -2159 -4838 -2127 -4837
rect -2044 -4837 -2001 -4824
rect -1849 -4825 -1681 -4783
rect -1849 -4837 -1807 -4825
rect -2044 -4838 -2011 -4837
rect -2753 -4895 -2651 -4842
rect -2433 -4842 -2387 -4840
rect -2377 -4842 -2331 -4840
rect -2433 -4896 -2331 -4842
rect -2113 -4842 -2067 -4838
rect -2057 -4842 -2011 -4838
rect -1839 -4839 -1807 -4837
rect -1724 -4839 -1681 -4825
rect -2113 -4894 -2011 -4842
rect -1793 -4851 -1747 -4839
rect -1737 -4851 -1681 -4839
rect -1793 -4895 -1681 -4851
rect -2972 -4930 -2798 -4929
rect -3133 -4974 -2798 -4930
rect -3133 -4975 -2927 -4974
rect -3133 -4986 -3088 -4975
rect -3004 -4985 -2927 -4975
rect -2843 -4985 -2798 -4974
rect -3004 -4986 -2959 -4985
rect -3077 -4991 -3031 -4986
rect -3015 -4987 -2959 -4986
rect -3015 -4991 -2969 -4987
rect -3077 -5047 -2969 -4991
rect -2916 -4991 -2870 -4985
rect -2854 -4987 -2798 -4985
rect -2332 -4975 -2158 -4930
rect -2332 -4986 -2288 -4975
rect -2202 -4986 -2158 -4975
rect -1692 -4974 -1358 -4930
rect -1692 -4986 -1647 -4974
rect -1563 -4975 -1358 -4974
rect -1563 -4986 -1487 -4975
rect -1403 -4986 -1358 -4975
rect -2854 -4991 -2808 -4987
rect -2916 -5047 -2808 -4991
rect -2276 -4991 -2230 -4986
rect -2214 -4987 -2158 -4986
rect -2214 -4991 -2168 -4987
rect -2276 -5047 -2168 -4991
rect -1636 -4991 -1590 -4986
rect -1574 -4987 -1518 -4986
rect -1574 -4991 -1528 -4987
rect -1636 -5047 -1528 -4991
rect -1476 -5003 -1430 -4986
rect -1414 -5003 -1358 -4986
rect -3077 -5048 -2959 -5047
rect -2276 -5048 -2158 -5047
rect -1636 -5048 -1518 -5047
rect -1476 -5048 -1358 -5003
rect -2876 -5245 -2728 -5220
rect -2876 -5266 -2851 -5245
rect -2750 -5266 -2728 -5245
rect -2830 -5276 -2784 -5266
rect -2774 -5267 -2728 -5266
rect -2830 -5277 -2783 -5276
rect -2774 -5277 -2737 -5267
rect -2830 -5306 -2737 -5277
rect -2830 -5322 -2774 -5306
rect -2649 -5528 -2481 -5486
rect -2008 -5527 -1840 -5486
rect -2649 -5542 -2607 -5528
rect -2524 -5540 -2481 -5528
rect -2524 -5542 -2491 -5540
rect -1998 -5542 -1965 -5527
rect -1882 -5542 -1840 -5527
rect -2593 -5544 -2547 -5542
rect -2537 -5544 -2491 -5542
rect -2593 -5598 -2491 -5544
rect -1952 -5555 -1906 -5542
rect -1896 -5555 -1840 -5542
rect -1952 -5598 -1840 -5555
rect -2811 -5680 -2643 -5638
rect -2811 -5691 -2769 -5680
rect -2801 -5694 -2769 -5691
rect -2686 -5691 -2643 -5680
rect -2489 -5679 -2321 -5637
rect -2489 -5691 -2447 -5679
rect -2686 -5694 -2653 -5691
rect -2479 -5693 -2447 -5691
rect -2364 -5691 -2321 -5679
rect -2171 -5679 -2003 -5637
rect -2171 -5691 -2129 -5679
rect -2364 -5693 -2331 -5691
rect -2161 -5693 -2129 -5691
rect -2046 -5691 -2003 -5679
rect -1848 -5679 -1680 -5637
rect -1848 -5691 -1806 -5679
rect -2046 -5693 -2013 -5691
rect -1838 -5693 -1806 -5691
rect -1723 -5693 -1680 -5679
rect -2755 -5696 -2709 -5694
rect -2699 -5696 -2653 -5694
rect -2755 -5750 -2653 -5696
rect -2433 -5696 -2387 -5693
rect -2377 -5696 -2331 -5693
rect -2433 -5749 -2331 -5696
rect -2115 -5696 -2069 -5693
rect -2059 -5696 -2013 -5693
rect -2115 -5749 -2013 -5696
rect -1792 -5705 -1746 -5693
rect -1736 -5705 -1680 -5693
rect -1792 -5749 -1680 -5705
rect -3130 -5834 -2801 -5793
rect -3130 -5835 -2927 -5834
rect -3130 -5849 -3088 -5835
rect -3004 -5847 -2927 -5835
rect -3004 -5849 -2972 -5847
rect -2959 -5849 -2927 -5847
rect -2843 -5847 -2801 -5834
rect -2330 -5835 -2160 -5793
rect -2330 -5847 -2288 -5835
rect -2843 -5849 -2811 -5847
rect -2320 -5849 -2288 -5847
rect -2202 -5847 -2160 -5835
rect -1689 -5834 -1361 -5793
rect -1689 -5847 -1647 -5834
rect -2202 -5849 -2170 -5847
rect -1679 -5849 -1647 -5847
rect -1563 -5835 -1361 -5834
rect -1563 -5847 -1487 -5835
rect -1563 -5849 -1531 -5847
rect -1519 -5849 -1487 -5847
rect -1403 -5849 -1361 -5835
rect -3074 -5851 -3028 -5849
rect -3018 -5851 -2972 -5849
rect -3074 -5905 -2972 -5851
rect -2913 -5851 -2867 -5849
rect -2857 -5851 -2811 -5849
rect -2913 -5905 -2811 -5851
rect -2274 -5851 -2228 -5849
rect -2216 -5851 -2170 -5849
rect -2274 -5905 -2170 -5851
rect -1633 -5851 -1587 -5849
rect -1577 -5851 -1531 -5849
rect -1633 -5905 -1531 -5851
rect -1473 -5863 -1427 -5849
rect -1417 -5863 -1361 -5849
rect -1473 -5905 -1361 -5863
rect -1767 -6066 -1619 -6041
rect -1767 -6087 -1665 -6066
rect -1754 -6093 -1721 -6087
rect -1708 -6093 -1697 -6087
rect -1719 -6097 -1675 -6093
rect -1721 -6143 -1665 -6097
rect -1641 -6143 -1619 -6066
<< nwell >>
rect -3356 -2050 -1223 1494
rect -3327 -6363 -1192 -2523
rect -801 -3402 1273 1072
rect -515 -6334 1318 -4010
rect 2632 -6145 5214 -5425
rect 2632 -6339 4327 -6145
rect 4440 -6339 5214 -6145
rect 2632 -6568 5214 -6339
rect 2632 -6704 3180 -6568
rect 3236 -6704 5214 -6568
rect 2632 -7048 5214 -6704
<< pwell >>
rect -3356 -10473 -1146 -6788
rect -610 -10718 1318 -6466
rect 2853 -8434 4966 -7343
<< pdiff >>
rect -2435 -4033 -2373 -3971
<< psubdiff >>
rect -564 -6512 1276 -6497
rect -564 -6558 -549 -6512
rect -503 -6558 -451 -6512
rect -405 -6558 -353 -6512
rect -307 -6558 -255 -6512
rect -209 -6558 -157 -6512
rect -111 -6558 -59 -6512
rect -13 -6558 39 -6512
rect 85 -6558 137 -6512
rect 183 -6558 235 -6512
rect 281 -6558 333 -6512
rect 379 -6558 431 -6512
rect 477 -6558 529 -6512
rect 575 -6558 627 -6512
rect 673 -6558 725 -6512
rect 771 -6558 823 -6512
rect 869 -6558 921 -6512
rect 967 -6558 1019 -6512
rect 1065 -6558 1117 -6512
rect 1163 -6558 1215 -6512
rect 1261 -6558 1276 -6512
rect -564 -6573 1276 -6558
rect -564 -6610 -488 -6573
rect -564 -6656 -549 -6610
rect -503 -6656 -488 -6610
rect -564 -6708 -488 -6656
rect -564 -6754 -549 -6708
rect -503 -6754 -488 -6708
rect -564 -6806 -488 -6754
rect -3310 -6842 -1176 -6827
rect -3310 -6888 -3295 -6842
rect -3249 -6888 -3197 -6842
rect -3151 -6888 -3099 -6842
rect -3053 -6888 -3001 -6842
rect -2955 -6888 -2903 -6842
rect -2857 -6888 -2805 -6842
rect -2759 -6888 -2707 -6842
rect -2661 -6888 -2609 -6842
rect -2563 -6888 -2511 -6842
rect -2465 -6888 -2413 -6842
rect -2367 -6888 -2315 -6842
rect -2269 -6888 -2217 -6842
rect -2171 -6888 -2119 -6842
rect -2073 -6888 -2021 -6842
rect -1975 -6888 -1923 -6842
rect -1877 -6888 -1825 -6842
rect -1779 -6888 -1727 -6842
rect -1681 -6888 -1629 -6842
rect -1583 -6888 -1531 -6842
rect -1485 -6888 -1433 -6842
rect -1387 -6888 -1335 -6842
rect -1289 -6888 -1237 -6842
rect -1191 -6888 -1176 -6842
rect -3310 -6903 -1176 -6888
rect -3310 -6940 -3234 -6903
rect -3310 -6986 -3295 -6940
rect -3249 -6986 -3234 -6940
rect -3310 -7038 -3234 -6986
rect -3310 -7084 -3295 -7038
rect -3249 -7084 -3234 -7038
rect -1252 -6940 -1176 -6903
rect -1252 -6986 -1237 -6940
rect -1191 -6986 -1176 -6940
rect -1252 -7038 -1176 -6986
rect -3310 -7136 -3234 -7084
rect -3310 -7182 -3295 -7136
rect -3249 -7182 -3234 -7136
rect -1252 -7084 -1237 -7038
rect -1191 -7084 -1176 -7038
rect -1252 -7136 -1176 -7084
rect -3310 -7234 -3234 -7182
rect -3310 -7280 -3295 -7234
rect -3249 -7280 -3234 -7234
rect -3310 -7332 -3234 -7280
rect -3310 -7378 -3295 -7332
rect -3249 -7378 -3234 -7332
rect -3310 -7430 -3234 -7378
rect -3310 -7476 -3295 -7430
rect -3249 -7476 -3234 -7430
rect -3310 -7528 -3234 -7476
rect -3310 -7574 -3295 -7528
rect -3249 -7574 -3234 -7528
rect -3310 -7626 -3234 -7574
rect -3310 -7672 -3295 -7626
rect -3249 -7672 -3234 -7626
rect -3310 -7724 -3234 -7672
rect -3310 -7770 -3295 -7724
rect -3249 -7770 -3234 -7724
rect -1252 -7182 -1237 -7136
rect -1191 -7182 -1176 -7136
rect -1252 -7234 -1176 -7182
rect -1252 -7280 -1237 -7234
rect -1191 -7280 -1176 -7234
rect -1252 -7332 -1176 -7280
rect -1252 -7378 -1237 -7332
rect -1191 -7378 -1176 -7332
rect -1252 -7430 -1176 -7378
rect -1252 -7476 -1237 -7430
rect -1191 -7476 -1176 -7430
rect -1252 -7528 -1176 -7476
rect -1252 -7574 -1237 -7528
rect -1191 -7574 -1176 -7528
rect -1252 -7626 -1176 -7574
rect -1252 -7672 -1237 -7626
rect -1191 -7672 -1176 -7626
rect -1252 -7724 -1176 -7672
rect -3310 -7822 -3234 -7770
rect -3310 -7868 -3295 -7822
rect -3249 -7868 -3234 -7822
rect -1252 -7770 -1237 -7724
rect -1191 -7770 -1176 -7724
rect -3310 -7920 -3234 -7868
rect -1252 -7822 -1176 -7770
rect -3310 -7966 -3295 -7920
rect -3249 -7966 -3234 -7920
rect -1252 -7868 -1237 -7822
rect -1191 -7868 -1176 -7822
rect -1252 -7920 -1176 -7868
rect -3310 -8018 -3234 -7966
rect -3310 -8064 -3295 -8018
rect -3249 -8064 -3234 -8018
rect -3310 -8116 -3234 -8064
rect -3310 -8162 -3295 -8116
rect -3249 -8162 -3234 -8116
rect -3310 -8214 -3234 -8162
rect -3310 -8260 -3295 -8214
rect -3249 -8260 -3234 -8214
rect -3310 -8312 -3234 -8260
rect -3310 -8358 -3295 -8312
rect -3249 -8358 -3234 -8312
rect -3310 -8410 -3234 -8358
rect -3310 -8456 -3295 -8410
rect -3249 -8456 -3234 -8410
rect -3310 -8508 -3234 -8456
rect -3310 -8554 -3295 -8508
rect -3249 -8554 -3234 -8508
rect -1252 -7966 -1237 -7920
rect -1191 -7966 -1176 -7920
rect -1252 -8018 -1176 -7966
rect -1252 -8064 -1237 -8018
rect -1191 -8064 -1176 -8018
rect -1252 -8116 -1176 -8064
rect -1252 -8162 -1237 -8116
rect -1191 -8162 -1176 -8116
rect -1252 -8214 -1176 -8162
rect -1252 -8260 -1237 -8214
rect -1191 -8260 -1176 -8214
rect -1252 -8312 -1176 -8260
rect -1252 -8358 -1237 -8312
rect -1191 -8358 -1176 -8312
rect -1252 -8410 -1176 -8358
rect -1252 -8456 -1237 -8410
rect -1191 -8456 -1176 -8410
rect -1252 -8508 -1176 -8456
rect -3310 -8606 -3234 -8554
rect -3310 -8652 -3295 -8606
rect -3249 -8652 -3234 -8606
rect -1252 -8554 -1237 -8508
rect -1191 -8554 -1176 -8508
rect -3310 -8704 -3234 -8652
rect -3310 -8750 -3295 -8704
rect -3249 -8750 -3234 -8704
rect -1252 -8606 -1176 -8554
rect -1252 -8652 -1237 -8606
rect -1191 -8652 -1176 -8606
rect -1252 -8704 -1176 -8652
rect -3310 -8802 -3234 -8750
rect -3310 -8848 -3295 -8802
rect -3249 -8848 -3234 -8802
rect -3310 -8900 -3234 -8848
rect -3310 -8946 -3295 -8900
rect -3249 -8946 -3234 -8900
rect -3310 -8998 -3234 -8946
rect -3310 -9044 -3295 -8998
rect -3249 -9044 -3234 -8998
rect -3310 -9096 -3234 -9044
rect -3310 -9142 -3295 -9096
rect -3249 -9142 -3234 -9096
rect -3310 -9194 -3234 -9142
rect -3310 -9240 -3295 -9194
rect -3249 -9240 -3234 -9194
rect -3310 -9292 -3234 -9240
rect -3310 -9338 -3295 -9292
rect -3249 -9338 -3234 -9292
rect -1252 -8750 -1237 -8704
rect -1191 -8750 -1176 -8704
rect -1252 -8802 -1176 -8750
rect -1252 -8848 -1237 -8802
rect -1191 -8848 -1176 -8802
rect -1252 -8900 -1176 -8848
rect -1252 -8946 -1237 -8900
rect -1191 -8946 -1176 -8900
rect -1252 -8998 -1176 -8946
rect -1252 -9044 -1237 -8998
rect -1191 -9044 -1176 -8998
rect -1252 -9096 -1176 -9044
rect -1252 -9142 -1237 -9096
rect -1191 -9142 -1176 -9096
rect -1252 -9194 -1176 -9142
rect -1252 -9240 -1237 -9194
rect -1191 -9240 -1176 -9194
rect -1252 -9292 -1176 -9240
rect -3310 -9390 -3234 -9338
rect -3310 -9436 -3295 -9390
rect -3249 -9436 -3234 -9390
rect -3310 -9488 -3234 -9436
rect -1252 -9338 -1237 -9292
rect -1191 -9338 -1176 -9292
rect -3310 -9534 -3295 -9488
rect -3249 -9534 -3234 -9488
rect -3310 -9586 -3234 -9534
rect -1252 -9390 -1176 -9338
rect -1252 -9436 -1237 -9390
rect -1191 -9436 -1176 -9390
rect -1252 -9488 -1176 -9436
rect -1252 -9534 -1237 -9488
rect -1191 -9534 -1176 -9488
rect -3310 -9632 -3295 -9586
rect -3249 -9632 -3234 -9586
rect -3310 -9684 -3234 -9632
rect -3310 -9730 -3295 -9684
rect -3249 -9730 -3234 -9684
rect -3310 -9782 -3234 -9730
rect -3310 -9828 -3295 -9782
rect -3249 -9828 -3234 -9782
rect -3310 -9880 -3234 -9828
rect -3310 -9926 -3295 -9880
rect -3249 -9926 -3234 -9880
rect -3310 -9978 -3234 -9926
rect -3310 -10024 -3295 -9978
rect -3249 -10024 -3234 -9978
rect -3310 -10076 -3234 -10024
rect -3310 -10122 -3295 -10076
rect -3249 -10122 -3234 -10076
rect -3310 -10174 -3234 -10122
rect -1252 -9586 -1176 -9534
rect -1252 -9632 -1237 -9586
rect -1191 -9632 -1176 -9586
rect -1252 -9684 -1176 -9632
rect -1252 -9730 -1237 -9684
rect -1191 -9730 -1176 -9684
rect -1252 -9782 -1176 -9730
rect -1252 -9828 -1237 -9782
rect -1191 -9828 -1176 -9782
rect -1252 -9880 -1176 -9828
rect -1252 -9926 -1237 -9880
rect -1191 -9926 -1176 -9880
rect -1252 -9978 -1176 -9926
rect -1252 -10024 -1237 -9978
rect -1191 -10024 -1176 -9978
rect -1252 -10076 -1176 -10024
rect -1252 -10122 -1237 -10076
rect -1191 -10122 -1176 -10076
rect -3310 -10220 -3295 -10174
rect -3249 -10220 -3234 -10174
rect -1252 -10174 -1176 -10122
rect -3310 -10272 -3234 -10220
rect -3310 -10318 -3295 -10272
rect -3249 -10318 -3234 -10272
rect -3310 -10355 -3234 -10318
rect -1252 -10220 -1237 -10174
rect -1191 -10220 -1176 -10174
rect -1252 -10272 -1176 -10220
rect -1252 -10318 -1237 -10272
rect -1191 -10318 -1176 -10272
rect -1252 -10355 -1176 -10318
rect -3310 -10370 -1176 -10355
rect -3310 -10416 -3295 -10370
rect -3249 -10416 -3197 -10370
rect -3151 -10416 -3099 -10370
rect -3053 -10416 -3001 -10370
rect -2955 -10416 -2903 -10370
rect -2857 -10416 -2805 -10370
rect -2759 -10416 -2707 -10370
rect -2661 -10416 -2609 -10370
rect -2563 -10416 -2511 -10370
rect -2465 -10416 -2413 -10370
rect -2367 -10416 -2315 -10370
rect -2269 -10416 -2217 -10370
rect -2171 -10416 -2119 -10370
rect -2073 -10416 -2021 -10370
rect -1975 -10416 -1923 -10370
rect -1877 -10416 -1825 -10370
rect -1779 -10416 -1727 -10370
rect -1681 -10416 -1629 -10370
rect -1583 -10416 -1531 -10370
rect -1485 -10416 -1433 -10370
rect -1387 -10416 -1335 -10370
rect -1289 -10416 -1237 -10370
rect -1191 -10416 -1176 -10370
rect -3310 -10431 -1176 -10416
rect -564 -6852 -549 -6806
rect -503 -6852 -488 -6806
rect 1200 -6610 1276 -6573
rect 1200 -6656 1215 -6610
rect 1261 -6656 1276 -6610
rect 1200 -6708 1276 -6656
rect 1200 -6754 1215 -6708
rect 1261 -6754 1276 -6708
rect 1200 -6806 1276 -6754
rect -564 -6904 -488 -6852
rect -564 -6950 -549 -6904
rect -503 -6950 -488 -6904
rect 1200 -6852 1215 -6806
rect 1261 -6852 1276 -6806
rect 1200 -6904 1276 -6852
rect -564 -7002 -488 -6950
rect -564 -7048 -549 -7002
rect -503 -7048 -488 -7002
rect -564 -7100 -488 -7048
rect -564 -7146 -549 -7100
rect -503 -7146 -488 -7100
rect -564 -7198 -488 -7146
rect -564 -7244 -549 -7198
rect -503 -7244 -488 -7198
rect -564 -7296 -488 -7244
rect -564 -7342 -549 -7296
rect -503 -7342 -488 -7296
rect -564 -7394 -488 -7342
rect -564 -7440 -549 -7394
rect -503 -7440 -488 -7394
rect -564 -7492 -488 -7440
rect -564 -7538 -549 -7492
rect -503 -7538 -488 -7492
rect -564 -7590 -488 -7538
rect -564 -7636 -549 -7590
rect -503 -7636 -488 -7590
rect 1200 -6950 1215 -6904
rect 1261 -6950 1276 -6904
rect 1200 -7002 1276 -6950
rect 1200 -7048 1215 -7002
rect 1261 -7048 1276 -7002
rect 1200 -7100 1276 -7048
rect 1200 -7146 1215 -7100
rect 1261 -7146 1276 -7100
rect 1200 -7198 1276 -7146
rect 1200 -7244 1215 -7198
rect 1261 -7244 1276 -7198
rect 1200 -7296 1276 -7244
rect 1200 -7342 1215 -7296
rect 1261 -7342 1276 -7296
rect 1200 -7394 1276 -7342
rect 1200 -7440 1215 -7394
rect 1261 -7440 1276 -7394
rect 1200 -7492 1276 -7440
rect 1200 -7538 1215 -7492
rect 1261 -7538 1276 -7492
rect 1200 -7590 1276 -7538
rect -564 -7688 -488 -7636
rect -564 -7734 -549 -7688
rect -503 -7734 -488 -7688
rect -564 -7786 -488 -7734
rect -564 -7832 -549 -7786
rect -503 -7832 -488 -7786
rect 1200 -7636 1215 -7590
rect 1261 -7636 1276 -7590
rect 1200 -7688 1276 -7636
rect 1200 -7734 1215 -7688
rect 1261 -7734 1276 -7688
rect 1200 -7786 1276 -7734
rect -564 -7884 -488 -7832
rect -564 -7930 -549 -7884
rect -503 -7930 -488 -7884
rect -564 -7982 -488 -7930
rect -564 -8028 -549 -7982
rect -503 -8028 -488 -7982
rect -564 -8080 -488 -8028
rect -564 -8126 -549 -8080
rect -503 -8126 -488 -8080
rect -564 -8178 -488 -8126
rect -564 -8224 -549 -8178
rect -503 -8224 -488 -8178
rect -564 -8276 -488 -8224
rect -564 -8322 -549 -8276
rect -503 -8322 -488 -8276
rect -564 -8374 -488 -8322
rect -564 -8420 -549 -8374
rect -503 -8420 -488 -8374
rect -564 -8472 -488 -8420
rect -564 -8518 -549 -8472
rect -503 -8518 -488 -8472
rect 1200 -7832 1215 -7786
rect 1261 -7832 1276 -7786
rect 1200 -7884 1276 -7832
rect 1200 -7930 1215 -7884
rect 1261 -7930 1276 -7884
rect 1200 -7982 1276 -7930
rect 1200 -8028 1215 -7982
rect 1261 -8028 1276 -7982
rect 1200 -8080 1276 -8028
rect 1200 -8126 1215 -8080
rect 1261 -8126 1276 -8080
rect 1200 -8178 1276 -8126
rect 1200 -8224 1215 -8178
rect 1261 -8224 1276 -8178
rect 1200 -8276 1276 -8224
rect 1200 -8322 1215 -8276
rect 1261 -8322 1276 -8276
rect 1200 -8374 1276 -8322
rect 3046 -8156 4681 -8126
rect 3046 -8294 3076 -8156
rect 4649 -8294 4681 -8156
rect 3046 -8326 4681 -8294
rect 1200 -8420 1215 -8374
rect 1261 -8420 1276 -8374
rect 1200 -8472 1276 -8420
rect -564 -8570 -488 -8518
rect -564 -8616 -549 -8570
rect -503 -8616 -488 -8570
rect -564 -8668 -488 -8616
rect -564 -8714 -549 -8668
rect -503 -8714 -488 -8668
rect -564 -8766 -488 -8714
rect -564 -8812 -549 -8766
rect -503 -8812 -488 -8766
rect 1200 -8518 1215 -8472
rect 1261 -8518 1276 -8472
rect 1200 -8570 1276 -8518
rect 1200 -8616 1215 -8570
rect 1261 -8616 1276 -8570
rect 1200 -8668 1276 -8616
rect 1200 -8714 1215 -8668
rect 1261 -8714 1276 -8668
rect 1200 -8766 1276 -8714
rect -564 -8864 -488 -8812
rect -564 -8910 -549 -8864
rect -503 -8910 -488 -8864
rect -564 -8962 -488 -8910
rect -564 -9008 -549 -8962
rect -503 -9008 -488 -8962
rect -564 -9060 -488 -9008
rect -564 -9106 -549 -9060
rect -503 -9106 -488 -9060
rect -564 -9158 -488 -9106
rect -564 -9204 -549 -9158
rect -503 -9204 -488 -9158
rect -564 -9256 -488 -9204
rect -564 -9302 -549 -9256
rect -503 -9302 -488 -9256
rect -564 -9354 -488 -9302
rect -564 -9400 -549 -9354
rect -503 -9400 -488 -9354
rect -564 -9452 -488 -9400
rect -564 -9498 -549 -9452
rect -503 -9498 -488 -9452
rect 1200 -8812 1215 -8766
rect 1261 -8812 1276 -8766
rect 1200 -8864 1276 -8812
rect 1200 -8910 1215 -8864
rect 1261 -8910 1276 -8864
rect 1200 -8962 1276 -8910
rect 1200 -9008 1215 -8962
rect 1261 -9008 1276 -8962
rect 1200 -9060 1276 -9008
rect 1200 -9106 1215 -9060
rect 1261 -9106 1276 -9060
rect 1200 -9158 1276 -9106
rect 1200 -9204 1215 -9158
rect 1261 -9204 1276 -9158
rect 1200 -9256 1276 -9204
rect 1200 -9302 1215 -9256
rect 1261 -9302 1276 -9256
rect 1200 -9354 1276 -9302
rect 1200 -9400 1215 -9354
rect 1261 -9400 1276 -9354
rect 1200 -9452 1276 -9400
rect -564 -9550 -488 -9498
rect -564 -9596 -549 -9550
rect -503 -9596 -488 -9550
rect -564 -9648 -488 -9596
rect 1200 -9498 1215 -9452
rect 1261 -9498 1276 -9452
rect 1200 -9550 1276 -9498
rect 1200 -9596 1215 -9550
rect 1261 -9596 1276 -9550
rect -564 -9694 -549 -9648
rect -503 -9694 -488 -9648
rect -564 -9746 -488 -9694
rect -564 -9792 -549 -9746
rect -503 -9792 -488 -9746
rect -564 -9844 -488 -9792
rect -564 -9890 -549 -9844
rect -503 -9890 -488 -9844
rect -564 -9942 -488 -9890
rect -564 -9988 -549 -9942
rect -503 -9988 -488 -9942
rect -564 -10040 -488 -9988
rect -564 -10086 -549 -10040
rect -503 -10086 -488 -10040
rect -564 -10138 -488 -10086
rect -564 -10184 -549 -10138
rect -503 -10184 -488 -10138
rect -564 -10236 -488 -10184
rect -564 -10282 -549 -10236
rect -503 -10282 -488 -10236
rect -564 -10334 -488 -10282
rect 1200 -9648 1276 -9596
rect 1200 -9694 1215 -9648
rect 1261 -9694 1276 -9648
rect 1200 -9746 1276 -9694
rect 1200 -9792 1215 -9746
rect 1261 -9792 1276 -9746
rect 1200 -9844 1276 -9792
rect 1200 -9890 1215 -9844
rect 1261 -9890 1276 -9844
rect 1200 -9942 1276 -9890
rect 1200 -9988 1215 -9942
rect 1261 -9988 1276 -9942
rect 1200 -10040 1276 -9988
rect 1200 -10086 1215 -10040
rect 1261 -10086 1276 -10040
rect 1200 -10138 1276 -10086
rect 1200 -10184 1215 -10138
rect 1261 -10184 1276 -10138
rect 1200 -10236 1276 -10184
rect 1200 -10282 1215 -10236
rect 1261 -10282 1276 -10236
rect -564 -10380 -549 -10334
rect -503 -10380 -488 -10334
rect -564 -10432 -488 -10380
rect 1200 -10334 1276 -10282
rect 1200 -10380 1215 -10334
rect 1261 -10380 1276 -10334
rect -564 -10478 -549 -10432
rect -503 -10478 -488 -10432
rect -564 -10530 -488 -10478
rect -564 -10576 -549 -10530
rect -503 -10576 -488 -10530
rect -564 -10613 -488 -10576
rect 1200 -10432 1276 -10380
rect 1200 -10478 1215 -10432
rect 1261 -10478 1276 -10432
rect 1200 -10530 1276 -10478
rect 1200 -10576 1215 -10530
rect 1261 -10576 1276 -10530
rect 1200 -10613 1276 -10576
rect -564 -10628 1276 -10613
rect -564 -10674 -549 -10628
rect -503 -10674 -451 -10628
rect -405 -10674 -353 -10628
rect -307 -10674 -255 -10628
rect -209 -10674 -157 -10628
rect -111 -10674 -59 -10628
rect -13 -10674 39 -10628
rect 85 -10674 137 -10628
rect 183 -10674 235 -10628
rect 281 -10674 333 -10628
rect 379 -10674 431 -10628
rect 477 -10674 529 -10628
rect 575 -10674 627 -10628
rect 673 -10674 725 -10628
rect 771 -10674 823 -10628
rect 869 -10674 921 -10628
rect 967 -10674 1019 -10628
rect 1065 -10674 1117 -10628
rect 1163 -10674 1215 -10628
rect 1261 -10674 1276 -10628
rect -564 -10689 1276 -10674
<< nsubdiff >>
rect -3309 1441 -1257 1456
rect -3309 1394 -3294 1441
rect -3247 1395 -3199 1441
rect -3153 1395 -3105 1441
rect -3059 1395 -3011 1441
rect -2965 1395 -2917 1441
rect -2871 1395 -2823 1441
rect -2777 1395 -2729 1441
rect -2683 1395 -2635 1441
rect -2589 1395 -2541 1441
rect -2495 1395 -2447 1441
rect -2401 1395 -2353 1441
rect -2307 1395 -2259 1441
rect -2213 1395 -2165 1441
rect -2119 1395 -2071 1441
rect -2025 1395 -1977 1441
rect -1931 1395 -1883 1441
rect -1837 1395 -1789 1441
rect -1743 1395 -1695 1441
rect -1649 1395 -1601 1441
rect -1555 1395 -1507 1441
rect -1461 1395 -1413 1441
rect -1367 1395 -1319 1441
rect -3247 1394 -1319 1395
rect -1272 1394 -1257 1441
rect -3309 1380 -1257 1394
rect -3309 1346 -3233 1380
rect -3309 1300 -3294 1346
rect -3248 1300 -3233 1346
rect -3309 1252 -3233 1300
rect -1333 1346 -1257 1380
rect -1333 1300 -1318 1346
rect -1272 1300 -1257 1346
rect -3309 1206 -3294 1252
rect -3248 1206 -3233 1252
rect -3309 1158 -3233 1206
rect -1333 1252 -1257 1300
rect -1333 1206 -1318 1252
rect -1272 1206 -1257 1252
rect -3309 1112 -3294 1158
rect -3248 1112 -3233 1158
rect -3309 1064 -3233 1112
rect -3309 1018 -3294 1064
rect -3248 1018 -3233 1064
rect -3309 970 -3233 1018
rect -3309 924 -3294 970
rect -3248 924 -3233 970
rect -3309 876 -3233 924
rect -3309 830 -3294 876
rect -3248 830 -3233 876
rect -3309 782 -3233 830
rect -3309 736 -3294 782
rect -3248 736 -3233 782
rect -3309 688 -3233 736
rect -3309 642 -3294 688
rect -3248 642 -3233 688
rect -3309 594 -3233 642
rect -3309 548 -3294 594
rect -3248 548 -3233 594
rect -3309 500 -3233 548
rect -1333 1158 -1257 1206
rect -1333 1112 -1318 1158
rect -1272 1112 -1257 1158
rect -1333 1064 -1257 1112
rect -1333 1018 -1318 1064
rect -1272 1018 -1257 1064
rect -1333 970 -1257 1018
rect -1333 924 -1318 970
rect -1272 924 -1257 970
rect -1333 876 -1257 924
rect -1333 830 -1318 876
rect -1272 830 -1257 876
rect -1333 782 -1257 830
rect -1333 736 -1318 782
rect -1272 736 -1257 782
rect -1333 688 -1257 736
rect -1333 642 -1318 688
rect -1272 642 -1257 688
rect -1333 594 -1257 642
rect -1333 548 -1318 594
rect -1272 548 -1257 594
rect -3309 454 -3294 500
rect -3248 454 -3233 500
rect -1333 500 -1257 548
rect -3309 406 -3233 454
rect -1333 454 -1318 500
rect -1272 454 -1257 500
rect -3309 360 -3294 406
rect -3248 360 -3233 406
rect -3309 312 -3233 360
rect -3309 266 -3294 312
rect -3248 266 -3233 312
rect -3309 218 -3233 266
rect -3309 172 -3294 218
rect -3248 172 -3233 218
rect -3309 124 -3233 172
rect -3309 78 -3294 124
rect -3248 78 -3233 124
rect -3309 30 -3233 78
rect -3309 -16 -3294 30
rect -3248 -16 -3233 30
rect -3309 -64 -3233 -16
rect -3309 -110 -3294 -64
rect -3248 -110 -3233 -64
rect -3309 -158 -3233 -110
rect -3309 -204 -3294 -158
rect -3248 -204 -3233 -158
rect -3309 -252 -3233 -204
rect -1333 406 -1257 454
rect -1333 360 -1318 406
rect -1272 360 -1257 406
rect -1333 312 -1257 360
rect -1333 266 -1318 312
rect -1272 266 -1257 312
rect -1333 218 -1257 266
rect -1333 172 -1318 218
rect -1272 172 -1257 218
rect -1333 124 -1257 172
rect -1333 78 -1318 124
rect -1272 78 -1257 124
rect -1333 30 -1257 78
rect -1333 -16 -1318 30
rect -1272 -16 -1257 30
rect -1333 -64 -1257 -16
rect -1333 -110 -1318 -64
rect -1272 -110 -1257 -64
rect -1333 -158 -1257 -110
rect -1333 -204 -1318 -158
rect -1272 -204 -1257 -158
rect -3309 -298 -3294 -252
rect -3248 -298 -3233 -252
rect -1333 -252 -1257 -204
rect -3309 -346 -3233 -298
rect -3309 -392 -3294 -346
rect -3248 -392 -3233 -346
rect -3309 -440 -3233 -392
rect -3309 -486 -3294 -440
rect -3248 -486 -3233 -440
rect -3309 -534 -3233 -486
rect -3309 -580 -3294 -534
rect -3248 -580 -3233 -534
rect -3309 -628 -3233 -580
rect -3309 -674 -3294 -628
rect -3248 -674 -3233 -628
rect -3309 -722 -3233 -674
rect -3309 -768 -3294 -722
rect -3248 -768 -3233 -722
rect -3309 -816 -3233 -768
rect -3309 -862 -3294 -816
rect -3248 -862 -3233 -816
rect -3309 -910 -3233 -862
rect -3309 -956 -3294 -910
rect -3248 -956 -3233 -910
rect -1333 -298 -1318 -252
rect -1272 -298 -1257 -252
rect -1333 -346 -1257 -298
rect -1333 -392 -1318 -346
rect -1272 -392 -1257 -346
rect -1333 -440 -1257 -392
rect -1333 -486 -1318 -440
rect -1272 -486 -1257 -440
rect -1333 -534 -1257 -486
rect -1333 -580 -1318 -534
rect -1272 -580 -1257 -534
rect -1333 -628 -1257 -580
rect -1333 -674 -1318 -628
rect -1272 -674 -1257 -628
rect -1333 -722 -1257 -674
rect -1333 -768 -1318 -722
rect -1272 -768 -1257 -722
rect -1333 -816 -1257 -768
rect -1333 -862 -1318 -816
rect -1272 -862 -1257 -816
rect -1333 -910 -1257 -862
rect -3309 -1004 -3233 -956
rect -3309 -1050 -3294 -1004
rect -3248 -1050 -3233 -1004
rect -1333 -956 -1318 -910
rect -1272 -956 -1257 -910
rect -1333 -1004 -1257 -956
rect -3309 -1098 -3233 -1050
rect -3309 -1144 -3294 -1098
rect -3248 -1144 -3233 -1098
rect -3309 -1192 -3233 -1144
rect -3309 -1238 -3294 -1192
rect -3248 -1238 -3233 -1192
rect -3309 -1286 -3233 -1238
rect -3309 -1332 -3294 -1286
rect -3248 -1332 -3233 -1286
rect -3309 -1380 -3233 -1332
rect -3309 -1426 -3294 -1380
rect -3248 -1426 -3233 -1380
rect -3309 -1474 -3233 -1426
rect -3309 -1520 -3294 -1474
rect -3248 -1520 -3233 -1474
rect -3309 -1568 -3233 -1520
rect -3309 -1614 -3294 -1568
rect -3248 -1614 -3233 -1568
rect -3309 -1662 -3233 -1614
rect -3309 -1708 -3294 -1662
rect -3248 -1708 -3233 -1662
rect -3309 -1756 -3233 -1708
rect -3309 -1802 -3294 -1756
rect -3248 -1802 -3233 -1756
rect -3309 -1850 -3233 -1802
rect -3309 -1896 -3294 -1850
rect -3248 -1896 -3233 -1850
rect -3309 -1929 -3233 -1896
rect -1333 -1050 -1318 -1004
rect -1272 -1050 -1257 -1004
rect -1333 -1098 -1257 -1050
rect -1333 -1144 -1318 -1098
rect -1272 -1144 -1257 -1098
rect -1333 -1192 -1257 -1144
rect -1333 -1238 -1318 -1192
rect -1272 -1238 -1257 -1192
rect -1333 -1286 -1257 -1238
rect -1333 -1332 -1318 -1286
rect -1272 -1332 -1257 -1286
rect -1333 -1380 -1257 -1332
rect -1333 -1426 -1318 -1380
rect -1272 -1426 -1257 -1380
rect -1333 -1474 -1257 -1426
rect -1333 -1520 -1318 -1474
rect -1272 -1520 -1257 -1474
rect -1333 -1568 -1257 -1520
rect -1333 -1614 -1318 -1568
rect -1272 -1614 -1257 -1568
rect -1333 -1662 -1257 -1614
rect -1333 -1708 -1318 -1662
rect -1272 -1708 -1257 -1662
rect -1333 -1756 -1257 -1708
rect -1333 -1802 -1318 -1756
rect -1272 -1802 -1257 -1756
rect -1333 -1850 -1257 -1802
rect -1333 -1896 -1318 -1850
rect -1272 -1896 -1257 -1850
rect -1333 -1929 -1257 -1896
rect -3309 -1944 -1257 -1929
rect -3309 -1990 -3293 -1944
rect -3247 -1990 -3199 -1944
rect -3153 -1990 -3105 -1944
rect -3059 -1990 -3011 -1944
rect -2965 -1990 -2917 -1944
rect -2871 -1990 -2823 -1944
rect -2777 -1990 -2729 -1944
rect -2683 -1990 -2635 -1944
rect -2589 -1990 -2541 -1944
rect -2495 -1990 -2447 -1944
rect -2401 -1990 -2353 -1944
rect -2307 -1990 -2259 -1944
rect -2213 -1990 -2165 -1944
rect -2119 -1990 -2071 -1944
rect -2025 -1990 -1977 -1944
rect -1931 -1990 -1883 -1944
rect -1837 -1990 -1789 -1944
rect -1743 -1990 -1695 -1944
rect -1649 -1990 -1601 -1944
rect -1555 -1990 -1507 -1944
rect -1461 -1990 -1413 -1944
rect -1367 -1990 -1319 -1944
rect -1273 -1990 -1257 -1944
rect -3309 -2005 -1257 -1990
rect -762 1013 1233 1028
rect -762 967 -747 1013
rect -701 967 -653 1013
rect -607 967 -552 1013
rect -506 967 -458 1013
rect -412 967 -362 1013
rect -316 967 -268 1013
rect -222 967 -167 1013
rect -121 967 -73 1013
rect -27 967 21 1013
rect 67 967 115 1013
rect 161 967 216 1013
rect 262 967 310 1013
rect 356 967 406 1013
rect 452 967 500 1013
rect 546 967 601 1013
rect 647 967 695 1013
rect 741 967 789 1013
rect 835 967 883 1013
rect 929 967 984 1013
rect 1030 967 1078 1013
rect 1124 967 1172 1013
rect 1218 967 1233 1013
rect -762 952 1233 967
rect -762 917 -686 952
rect -762 871 -747 917
rect -701 871 -686 917
rect -762 823 -686 871
rect 1157 917 1233 952
rect 1157 871 1172 917
rect 1218 871 1233 917
rect -762 777 -747 823
rect -701 777 -686 823
rect -762 727 -686 777
rect 1157 816 1233 871
rect 1157 770 1172 816
rect 1218 770 1233 816
rect -762 681 -747 727
rect -701 681 -686 727
rect -762 633 -686 681
rect -762 587 -747 633
rect -701 587 -686 633
rect -762 539 -686 587
rect -762 493 -747 539
rect -701 493 -686 539
rect -762 438 -686 493
rect -762 392 -747 438
rect -701 392 -686 438
rect -762 344 -686 392
rect -762 298 -747 344
rect -701 298 -686 344
rect -762 248 -686 298
rect -762 202 -747 248
rect -701 202 -686 248
rect -762 154 -686 202
rect -762 108 -747 154
rect -701 108 -686 154
rect -762 53 -686 108
rect 1157 722 1233 770
rect 1157 676 1172 722
rect 1218 676 1233 722
rect 1157 628 1233 676
rect 1157 582 1172 628
rect 1218 582 1233 628
rect 1157 534 1233 582
rect 1157 488 1172 534
rect 1218 488 1233 534
rect 1157 433 1233 488
rect 1157 387 1172 433
rect 1218 387 1233 433
rect 1157 339 1233 387
rect 1157 293 1172 339
rect 1218 293 1233 339
rect 1157 243 1233 293
rect 1157 197 1172 243
rect 1218 197 1233 243
rect 1157 149 1233 197
rect 1157 103 1172 149
rect 1218 103 1233 149
rect -762 7 -747 53
rect -701 7 -686 53
rect -762 -41 -686 7
rect -762 -87 -747 -41
rect -701 -87 -686 -41
rect -762 -135 -686 -87
rect -762 -181 -747 -135
rect -701 -181 -686 -135
rect -762 -229 -686 -181
rect -762 -275 -747 -229
rect -701 -275 -686 -229
rect -762 -330 -686 -275
rect 1157 48 1233 103
rect 1157 2 1172 48
rect 1218 2 1233 48
rect 1157 -46 1233 2
rect 1157 -92 1172 -46
rect 1218 -92 1233 -46
rect 1157 -140 1233 -92
rect 1157 -186 1172 -140
rect 1218 -186 1233 -140
rect 1157 -234 1233 -186
rect 1157 -280 1172 -234
rect 1218 -280 1233 -234
rect -762 -376 -747 -330
rect -701 -376 -686 -330
rect -762 -424 -686 -376
rect -762 -470 -747 -424
rect -701 -470 -686 -424
rect -762 -520 -686 -470
rect -762 -566 -747 -520
rect -701 -566 -686 -520
rect -762 -614 -686 -566
rect -762 -660 -747 -614
rect -701 -660 -686 -614
rect -762 -715 -686 -660
rect -762 -761 -747 -715
rect -701 -761 -686 -715
rect -762 -809 -686 -761
rect -762 -855 -747 -809
rect -701 -855 -686 -809
rect -762 -903 -686 -855
rect -762 -949 -747 -903
rect -701 -949 -686 -903
rect -762 -997 -686 -949
rect 1157 -335 1233 -280
rect 1157 -381 1172 -335
rect 1218 -381 1233 -335
rect 1157 -429 1233 -381
rect 1157 -475 1172 -429
rect 1218 -475 1233 -429
rect 1157 -525 1233 -475
rect 1157 -571 1172 -525
rect 1218 -571 1233 -525
rect 1157 -619 1233 -571
rect 1157 -665 1172 -619
rect 1218 -665 1233 -619
rect 1157 -720 1233 -665
rect 1157 -766 1172 -720
rect 1218 -766 1233 -720
rect 1157 -814 1233 -766
rect 1157 -860 1172 -814
rect 1218 -860 1233 -814
rect 1157 -908 1233 -860
rect 1157 -954 1172 -908
rect 1218 -954 1233 -908
rect -762 -1043 -747 -997
rect -701 -1043 -686 -997
rect -762 -1098 -686 -1043
rect -762 -1144 -747 -1098
rect -701 -1144 -686 -1098
rect -762 -1192 -686 -1144
rect -762 -1238 -747 -1192
rect -701 -1238 -686 -1192
rect -762 -1288 -686 -1238
rect -762 -1334 -747 -1288
rect -701 -1334 -686 -1288
rect 1157 -1004 1233 -954
rect 1157 -1050 1172 -1004
rect 1218 -1050 1233 -1004
rect 1157 -1098 1233 -1050
rect 1157 -1144 1172 -1098
rect 1218 -1144 1233 -1098
rect 1157 -1199 1233 -1144
rect 1157 -1245 1172 -1199
rect 1218 -1245 1233 -1199
rect 1157 -1293 1233 -1245
rect -762 -1382 -686 -1334
rect -762 -1428 -747 -1382
rect -701 -1428 -686 -1382
rect -762 -1476 -686 -1428
rect -762 -1522 -747 -1476
rect -701 -1522 -686 -1476
rect -762 -1577 -686 -1522
rect -762 -1623 -747 -1577
rect -701 -1623 -686 -1577
rect -762 -1671 -686 -1623
rect -762 -1717 -747 -1671
rect -701 -1717 -686 -1671
rect -762 -1767 -686 -1717
rect -762 -1813 -747 -1767
rect -701 -1813 -686 -1767
rect -762 -1861 -686 -1813
rect -762 -1907 -747 -1861
rect -701 -1907 -686 -1861
rect -762 -1962 -686 -1907
rect -762 -2008 -747 -1962
rect -701 -2008 -686 -1962
rect 1157 -1339 1172 -1293
rect 1218 -1339 1233 -1293
rect 1157 -1387 1233 -1339
rect 1157 -1433 1172 -1387
rect 1218 -1433 1233 -1387
rect 1157 -1481 1233 -1433
rect 1157 -1527 1172 -1481
rect 1218 -1527 1233 -1481
rect 1157 -1582 1233 -1527
rect 1157 -1628 1172 -1582
rect 1218 -1628 1233 -1582
rect 1157 -1676 1233 -1628
rect 1157 -1722 1172 -1676
rect 1218 -1722 1233 -1676
rect 1157 -1772 1233 -1722
rect 1157 -1818 1172 -1772
rect 1218 -1818 1233 -1772
rect 1157 -1866 1233 -1818
rect 1157 -1912 1172 -1866
rect 1218 -1912 1233 -1866
rect 1157 -1967 1233 -1912
rect -762 -2056 -686 -2008
rect -762 -2102 -747 -2056
rect -701 -2102 -686 -2056
rect -762 -2150 -686 -2102
rect -762 -2196 -747 -2150
rect -701 -2196 -686 -2150
rect -762 -2244 -686 -2196
rect -762 -2290 -747 -2244
rect -701 -2290 -686 -2244
rect -762 -2345 -686 -2290
rect -762 -2391 -747 -2345
rect -701 -2391 -686 -2345
rect 1157 -2013 1172 -1967
rect 1218 -2013 1233 -1967
rect 1157 -2061 1233 -2013
rect 1157 -2107 1172 -2061
rect 1218 -2107 1233 -2061
rect 1157 -2155 1233 -2107
rect 1157 -2201 1172 -2155
rect 1218 -2201 1233 -2155
rect 1157 -2249 1233 -2201
rect 1157 -2295 1172 -2249
rect 1218 -2295 1233 -2249
rect 1157 -2350 1233 -2295
rect -762 -2439 -686 -2391
rect -762 -2485 -747 -2439
rect -701 -2485 -686 -2439
rect -762 -2535 -686 -2485
rect -3282 -2593 -1230 -2578
rect -3282 -2640 -3267 -2593
rect -3220 -2639 -3172 -2593
rect -3126 -2639 -3078 -2593
rect -3032 -2639 -2984 -2593
rect -2938 -2639 -2890 -2593
rect -2844 -2639 -2796 -2593
rect -2750 -2639 -2702 -2593
rect -2656 -2639 -2608 -2593
rect -2562 -2639 -2514 -2593
rect -2468 -2639 -2420 -2593
rect -2374 -2639 -2326 -2593
rect -2280 -2639 -2232 -2593
rect -2186 -2639 -2138 -2593
rect -2092 -2639 -2044 -2593
rect -1998 -2639 -1950 -2593
rect -1904 -2639 -1856 -2593
rect -1810 -2639 -1762 -2593
rect -1716 -2639 -1668 -2593
rect -1622 -2639 -1574 -2593
rect -1528 -2639 -1480 -2593
rect -1434 -2639 -1386 -2593
rect -1340 -2639 -1292 -2593
rect -3220 -2640 -1292 -2639
rect -1245 -2640 -1230 -2593
rect -3282 -2654 -1230 -2640
rect -3282 -2688 -3206 -2654
rect -3282 -2734 -3267 -2688
rect -3221 -2734 -3206 -2688
rect -1306 -2688 -1230 -2654
rect -3282 -2782 -3206 -2734
rect -3282 -2828 -3267 -2782
rect -3221 -2828 -3206 -2782
rect -3282 -2876 -3206 -2828
rect -1306 -2734 -1291 -2688
rect -1245 -2734 -1230 -2688
rect -1306 -2782 -1230 -2734
rect -1306 -2828 -1291 -2782
rect -1245 -2828 -1230 -2782
rect -3282 -2922 -3267 -2876
rect -3221 -2922 -3206 -2876
rect -3282 -2970 -3206 -2922
rect -3282 -3016 -3267 -2970
rect -3221 -3016 -3206 -2970
rect -3282 -3064 -3206 -3016
rect -3282 -3110 -3267 -3064
rect -3221 -3110 -3206 -3064
rect -3282 -3158 -3206 -3110
rect -3282 -3204 -3267 -3158
rect -3221 -3204 -3206 -3158
rect -3282 -3252 -3206 -3204
rect -3282 -3298 -3267 -3252
rect -3221 -3298 -3206 -3252
rect -3282 -3346 -3206 -3298
rect -3282 -3392 -3267 -3346
rect -3221 -3392 -3206 -3346
rect -3282 -3440 -3206 -3392
rect -3282 -3486 -3267 -3440
rect -3221 -3486 -3206 -3440
rect -3282 -3534 -3206 -3486
rect -1306 -2876 -1230 -2828
rect -1306 -2922 -1291 -2876
rect -1245 -2922 -1230 -2876
rect -1306 -2970 -1230 -2922
rect -1306 -3016 -1291 -2970
rect -1245 -3016 -1230 -2970
rect -1306 -3064 -1230 -3016
rect -1306 -3110 -1291 -3064
rect -1245 -3110 -1230 -3064
rect -1306 -3158 -1230 -3110
rect -1306 -3204 -1291 -3158
rect -1245 -3204 -1230 -3158
rect -1306 -3252 -1230 -3204
rect -1306 -3298 -1291 -3252
rect -1245 -3298 -1230 -3252
rect -1306 -3346 -1230 -3298
rect -1306 -3392 -1291 -3346
rect -1245 -3392 -1230 -3346
rect -762 -2581 -747 -2535
rect -701 -2581 -686 -2535
rect -762 -2629 -686 -2581
rect -762 -2675 -747 -2629
rect -701 -2675 -686 -2629
rect -762 -2730 -686 -2675
rect -762 -2776 -747 -2730
rect -701 -2776 -686 -2730
rect -762 -2824 -686 -2776
rect -762 -2870 -747 -2824
rect -701 -2870 -686 -2824
rect -762 -2918 -686 -2870
rect -762 -2964 -747 -2918
rect -701 -2964 -686 -2918
rect -762 -3012 -686 -2964
rect -762 -3058 -747 -3012
rect -701 -3058 -686 -3012
rect 1157 -2396 1172 -2350
rect 1218 -2396 1233 -2350
rect 1157 -2444 1233 -2396
rect 1157 -2490 1172 -2444
rect 1218 -2490 1233 -2444
rect 1157 -2540 1233 -2490
rect 1157 -2586 1172 -2540
rect 1218 -2586 1233 -2540
rect 1157 -2634 1233 -2586
rect 1157 -2680 1172 -2634
rect 1218 -2680 1233 -2634
rect 1157 -2735 1233 -2680
rect 1157 -2781 1172 -2735
rect 1218 -2781 1233 -2735
rect 1157 -2829 1233 -2781
rect 1157 -2875 1172 -2829
rect 1218 -2875 1233 -2829
rect 1157 -2923 1233 -2875
rect 1157 -2969 1172 -2923
rect 1218 -2969 1233 -2923
rect 1157 -3019 1233 -2969
rect -762 -3113 -686 -3058
rect -762 -3159 -747 -3113
rect -701 -3159 -686 -3113
rect -762 -3207 -686 -3159
rect 1157 -3065 1172 -3019
rect 1218 -3065 1233 -3019
rect 1157 -3113 1233 -3065
rect 1157 -3159 1172 -3113
rect 1218 -3159 1233 -3113
rect -762 -3253 -747 -3207
rect -701 -3253 -686 -3207
rect -762 -3288 -686 -3253
rect 1157 -3207 1233 -3159
rect 1157 -3253 1172 -3207
rect 1218 -3253 1233 -3207
rect 1157 -3288 1233 -3253
rect -762 -3303 1233 -3288
rect -762 -3349 -747 -3303
rect -701 -3349 -653 -3303
rect -607 -3349 -552 -3303
rect -506 -3349 -458 -3303
rect -412 -3349 -362 -3303
rect -316 -3349 -268 -3303
rect -222 -3349 -167 -3303
rect -121 -3349 -73 -3303
rect -27 -3349 21 -3303
rect 67 -3349 115 -3303
rect 161 -3349 216 -3303
rect 262 -3349 310 -3303
rect 356 -3349 406 -3303
rect 452 -3349 500 -3303
rect 546 -3349 601 -3303
rect 647 -3349 695 -3303
rect 741 -3349 789 -3303
rect 835 -3349 883 -3303
rect 929 -3349 984 -3303
rect 1030 -3349 1078 -3303
rect 1124 -3349 1172 -3303
rect 1218 -3349 1233 -3303
rect -762 -3364 1233 -3349
rect -1306 -3440 -1230 -3392
rect -1306 -3486 -1291 -3440
rect -1245 -3486 -1230 -3440
rect -3282 -3580 -3267 -3534
rect -3221 -3580 -3206 -3534
rect -3282 -3628 -3206 -3580
rect -3282 -3674 -3267 -3628
rect -3221 -3674 -3206 -3628
rect -1306 -3534 -1230 -3486
rect -1306 -3580 -1291 -3534
rect -1245 -3580 -1230 -3534
rect -1306 -3628 -1230 -3580
rect -3282 -3722 -3206 -3674
rect -1306 -3674 -1291 -3628
rect -1245 -3674 -1230 -3628
rect -3282 -3768 -3267 -3722
rect -3221 -3768 -3206 -3722
rect -3282 -3816 -3206 -3768
rect -3282 -3862 -3267 -3816
rect -3221 -3862 -3206 -3816
rect -3282 -3910 -3206 -3862
rect -3282 -3956 -3267 -3910
rect -3221 -3956 -3206 -3910
rect -3282 -4004 -3206 -3956
rect -1306 -3722 -1230 -3674
rect -1306 -3768 -1291 -3722
rect -1245 -3768 -1230 -3722
rect -1306 -3816 -1230 -3768
rect -1306 -3862 -1291 -3816
rect -1245 -3862 -1230 -3816
rect -1306 -3910 -1230 -3862
rect -1306 -3956 -1291 -3910
rect -1245 -3956 -1230 -3910
rect -3282 -4050 -3267 -4004
rect -3221 -4050 -3206 -4004
rect -1306 -4004 -1230 -3956
rect -3282 -4098 -3206 -4050
rect -3282 -4144 -3267 -4098
rect -3221 -4144 -3206 -4098
rect -3282 -4192 -3206 -4144
rect -3282 -4238 -3267 -4192
rect -3221 -4238 -3206 -4192
rect -3282 -4286 -3206 -4238
rect -3282 -4332 -3267 -4286
rect -3221 -4332 -3206 -4286
rect -3282 -4380 -3206 -4332
rect -1306 -4050 -1291 -4004
rect -1245 -4050 -1230 -4004
rect -1306 -4098 -1230 -4050
rect -1306 -4144 -1291 -4098
rect -1245 -4144 -1230 -4098
rect -1306 -4192 -1230 -4144
rect -1306 -4238 -1291 -4192
rect -1245 -4238 -1230 -4192
rect -1306 -4286 -1230 -4238
rect -1306 -4332 -1291 -4286
rect -1245 -4332 -1230 -4286
rect -3282 -4426 -3267 -4380
rect -3221 -4426 -3206 -4380
rect -3282 -4474 -3206 -4426
rect -3282 -4520 -3267 -4474
rect -3221 -4520 -3206 -4474
rect -1306 -4380 -1230 -4332
rect -1306 -4426 -1291 -4380
rect -1245 -4426 -1230 -4380
rect -3282 -4568 -3206 -4520
rect -3282 -4614 -3267 -4568
rect -3221 -4614 -3206 -4568
rect -1306 -4474 -1230 -4426
rect -1306 -4520 -1291 -4474
rect -1245 -4520 -1230 -4474
rect -1306 -4568 -1230 -4520
rect -3282 -4662 -3206 -4614
rect -3282 -4708 -3267 -4662
rect -3221 -4708 -3206 -4662
rect -3282 -4756 -3206 -4708
rect -3282 -4802 -3267 -4756
rect -3221 -4802 -3206 -4756
rect -3282 -4850 -3206 -4802
rect -3282 -4896 -3267 -4850
rect -3221 -4896 -3206 -4850
rect -3282 -4944 -3206 -4896
rect -3282 -4990 -3267 -4944
rect -3221 -4990 -3206 -4944
rect -3282 -5038 -3206 -4990
rect -3282 -5084 -3267 -5038
rect -3221 -5084 -3206 -5038
rect -3282 -5132 -3206 -5084
rect -3282 -5178 -3267 -5132
rect -3221 -5178 -3206 -5132
rect -1306 -4614 -1291 -4568
rect -1245 -4614 -1230 -4568
rect -1306 -4662 -1230 -4614
rect -1306 -4708 -1291 -4662
rect -1245 -4708 -1230 -4662
rect -1306 -4756 -1230 -4708
rect -1306 -4802 -1291 -4756
rect -1245 -4802 -1230 -4756
rect -1306 -4850 -1230 -4802
rect -1306 -4896 -1291 -4850
rect -1245 -4896 -1230 -4850
rect -1306 -4944 -1230 -4896
rect -1306 -4990 -1291 -4944
rect -1245 -4990 -1230 -4944
rect -1306 -5038 -1230 -4990
rect -1306 -5084 -1291 -5038
rect -1245 -5084 -1230 -5038
rect -1306 -5132 -1230 -5084
rect -3282 -5226 -3206 -5178
rect -3282 -5272 -3267 -5226
rect -3221 -5272 -3206 -5226
rect -3282 -5320 -3206 -5272
rect -1306 -5178 -1291 -5132
rect -1245 -5178 -1230 -5132
rect -3282 -5366 -3267 -5320
rect -3221 -5366 -3206 -5320
rect -1306 -5226 -1230 -5178
rect -1306 -5272 -1291 -5226
rect -1245 -5272 -1230 -5226
rect -1306 -5320 -1230 -5272
rect -3282 -5414 -3206 -5366
rect -3282 -5460 -3267 -5414
rect -3221 -5460 -3206 -5414
rect -1306 -5366 -1291 -5320
rect -1245 -5366 -1230 -5320
rect -1306 -5414 -1230 -5366
rect -3282 -5508 -3206 -5460
rect -3282 -5554 -3267 -5508
rect -3221 -5554 -3206 -5508
rect -3282 -5602 -3206 -5554
rect -3282 -5648 -3267 -5602
rect -3221 -5648 -3206 -5602
rect -3282 -5696 -3206 -5648
rect -3282 -5742 -3267 -5696
rect -3221 -5742 -3206 -5696
rect -3282 -5790 -3206 -5742
rect -3282 -5836 -3267 -5790
rect -3221 -5836 -3206 -5790
rect -3282 -5884 -3206 -5836
rect -3282 -5930 -3267 -5884
rect -3221 -5930 -3206 -5884
rect -3282 -5978 -3206 -5930
rect -3282 -6024 -3267 -5978
rect -3221 -6024 -3206 -5978
rect -1306 -5460 -1291 -5414
rect -1245 -5460 -1230 -5414
rect -1306 -5508 -1230 -5460
rect -1306 -5554 -1291 -5508
rect -1245 -5554 -1230 -5508
rect -1306 -5602 -1230 -5554
rect -1306 -5648 -1291 -5602
rect -1245 -5648 -1230 -5602
rect -1306 -5696 -1230 -5648
rect -1306 -5742 -1291 -5696
rect -1245 -5742 -1230 -5696
rect -1306 -5790 -1230 -5742
rect -1306 -5836 -1291 -5790
rect -1245 -5836 -1230 -5790
rect -1306 -5884 -1230 -5836
rect -1306 -5930 -1291 -5884
rect -1245 -5930 -1230 -5884
rect -1306 -5978 -1230 -5930
rect -3282 -6072 -3206 -6024
rect -3282 -6118 -3267 -6072
rect -3221 -6118 -3206 -6072
rect -3282 -6166 -3206 -6118
rect -1306 -6024 -1291 -5978
rect -1245 -6024 -1230 -5978
rect -1306 -6072 -1230 -6024
rect -1306 -6118 -1291 -6072
rect -1245 -6118 -1230 -6072
rect -3282 -6212 -3267 -6166
rect -3221 -6212 -3206 -6166
rect -3282 -6245 -3206 -6212
rect -1306 -6166 -1230 -6118
rect -1306 -6212 -1291 -6166
rect -1245 -6212 -1230 -6166
rect -1306 -6245 -1230 -6212
rect -3282 -6260 -1230 -6245
rect -3282 -6306 -3266 -6260
rect -3220 -6306 -3172 -6260
rect -3126 -6306 -3078 -6260
rect -3032 -6306 -2984 -6260
rect -2938 -6306 -2890 -6260
rect -2844 -6306 -2796 -6260
rect -2750 -6306 -2702 -6260
rect -2656 -6306 -2608 -6260
rect -2562 -6306 -2514 -6260
rect -2468 -6306 -2420 -6260
rect -2374 -6306 -2326 -6260
rect -2280 -6306 -2232 -6260
rect -2186 -6306 -2138 -6260
rect -2092 -6306 -2044 -6260
rect -1998 -6306 -1950 -6260
rect -1904 -6306 -1856 -6260
rect -1810 -6306 -1762 -6260
rect -1716 -6306 -1668 -6260
rect -1622 -6306 -1574 -6260
rect -1528 -6306 -1480 -6260
rect -1434 -6306 -1386 -6260
rect -1340 -6306 -1292 -6260
rect -1246 -6306 -1230 -6260
rect -477 -4068 1293 -4053
rect -477 -4115 -462 -4068
rect -415 -4114 -367 -4068
rect -321 -4114 -273 -4068
rect -227 -4114 -179 -4068
rect -133 -4114 -85 -4068
rect -39 -4114 9 -4068
rect 55 -4114 103 -4068
rect 149 -4114 197 -4068
rect 243 -4114 291 -4068
rect 337 -4114 385 -4068
rect 431 -4114 479 -4068
rect 525 -4114 573 -4068
rect 619 -4114 667 -4068
rect 713 -4114 761 -4068
rect 807 -4114 855 -4068
rect 901 -4114 949 -4068
rect 995 -4114 1043 -4068
rect 1089 -4114 1137 -4068
rect 1183 -4114 1231 -4068
rect -415 -4115 1231 -4114
rect 1278 -4115 1293 -4068
rect -477 -4129 1293 -4115
rect -477 -4163 -401 -4129
rect -477 -4213 -462 -4163
rect -416 -4213 -401 -4163
rect -477 -4261 -401 -4213
rect 1217 -4163 1293 -4129
rect 1217 -4213 1232 -4163
rect 1278 -4213 1293 -4163
rect -477 -4307 -462 -4261
rect -416 -4307 -401 -4261
rect -477 -4355 -401 -4307
rect -477 -4401 -462 -4355
rect -416 -4401 -401 -4355
rect -477 -4449 -401 -4401
rect 1217 -4261 1293 -4213
rect 1217 -4307 1232 -4261
rect 1278 -4307 1293 -4261
rect 1217 -4355 1293 -4307
rect 1217 -4401 1232 -4355
rect 1278 -4401 1293 -4355
rect -477 -4495 -462 -4449
rect -416 -4495 -401 -4449
rect -477 -4543 -401 -4495
rect -477 -4589 -462 -4543
rect -416 -4589 -401 -4543
rect -477 -4637 -401 -4589
rect -477 -4683 -462 -4637
rect -416 -4683 -401 -4637
rect -477 -4731 -401 -4683
rect -477 -4777 -462 -4731
rect -416 -4777 -401 -4731
rect -477 -4825 -401 -4777
rect -477 -4871 -462 -4825
rect -416 -4871 -401 -4825
rect -477 -4919 -401 -4871
rect -477 -4965 -462 -4919
rect -416 -4965 -401 -4919
rect -477 -5013 -401 -4965
rect -477 -5059 -462 -5013
rect -416 -5059 -401 -5013
rect -477 -5107 -401 -5059
rect -477 -5153 -462 -5107
rect -416 -5153 -401 -5107
rect 1217 -4449 1293 -4401
rect 1217 -4495 1232 -4449
rect 1278 -4495 1293 -4449
rect 1217 -4543 1293 -4495
rect 1217 -4589 1232 -4543
rect 1278 -4589 1293 -4543
rect 1217 -4637 1293 -4589
rect 1217 -4683 1232 -4637
rect 1278 -4683 1293 -4637
rect 1217 -4731 1293 -4683
rect 1217 -4777 1232 -4731
rect 1278 -4777 1293 -4731
rect 1217 -4825 1293 -4777
rect 1217 -4871 1232 -4825
rect 1278 -4871 1293 -4825
rect 1217 -4919 1293 -4871
rect 1217 -4965 1232 -4919
rect 1278 -4965 1293 -4919
rect 1217 -5013 1293 -4965
rect 1217 -5059 1232 -5013
rect 1278 -5059 1293 -5013
rect 1217 -5107 1293 -5059
rect -477 -5201 -401 -5153
rect -477 -5247 -462 -5201
rect -416 -5247 -401 -5201
rect 1217 -5153 1232 -5107
rect 1278 -5153 1293 -5107
rect 1217 -5201 1293 -5153
rect -477 -5295 -401 -5247
rect -477 -5341 -462 -5295
rect -416 -5341 -401 -5295
rect -477 -5389 -401 -5341
rect -477 -5435 -462 -5389
rect -416 -5435 -401 -5389
rect -477 -5483 -401 -5435
rect -477 -5529 -462 -5483
rect -416 -5529 -401 -5483
rect -477 -5577 -401 -5529
rect -477 -5623 -462 -5577
rect -416 -5623 -401 -5577
rect -477 -5671 -401 -5623
rect -477 -5717 -462 -5671
rect -416 -5717 -401 -5671
rect -477 -5765 -401 -5717
rect -477 -5811 -462 -5765
rect -416 -5811 -401 -5765
rect -477 -5859 -401 -5811
rect -477 -5905 -462 -5859
rect -416 -5905 -401 -5859
rect -477 -5953 -401 -5905
rect -477 -5999 -462 -5953
rect -416 -5999 -401 -5953
rect -477 -6047 -401 -5999
rect -477 -6093 -462 -6047
rect -416 -6093 -401 -6047
rect -477 -6141 -401 -6093
rect -477 -6187 -462 -6141
rect -416 -6187 -401 -6141
rect -477 -6221 -401 -6187
rect 1217 -5247 1232 -5201
rect 1278 -5247 1293 -5201
rect 1217 -5295 1293 -5247
rect 1217 -5341 1232 -5295
rect 1278 -5341 1293 -5295
rect 1217 -5389 1293 -5341
rect 1217 -5435 1232 -5389
rect 1278 -5435 1293 -5389
rect 1217 -5483 1293 -5435
rect 1217 -5529 1232 -5483
rect 1278 -5529 1293 -5483
rect 1217 -5577 1293 -5529
rect 1217 -5623 1232 -5577
rect 1278 -5623 1293 -5577
rect 1217 -5671 1293 -5623
rect 1217 -5717 1232 -5671
rect 1278 -5717 1293 -5671
rect 1217 -5765 1293 -5717
rect 2977 -5557 4766 -5524
rect 2977 -5693 3066 -5557
rect 4667 -5693 4766 -5557
rect 2977 -5722 4766 -5693
rect 1217 -5811 1232 -5765
rect 1278 -5811 1293 -5765
rect 1217 -5859 1293 -5811
rect 1217 -5905 1232 -5859
rect 1278 -5905 1293 -5859
rect 1217 -5953 1293 -5905
rect 1217 -5999 1232 -5953
rect 1278 -5999 1293 -5953
rect 1217 -6047 1293 -5999
rect 1217 -6093 1232 -6047
rect 1278 -6093 1293 -6047
rect 1217 -6141 1293 -6093
rect 1217 -6187 1232 -6141
rect 1278 -6187 1293 -6141
rect 1217 -6221 1293 -6187
rect -477 -6235 1293 -6221
rect -477 -6282 -462 -6235
rect -415 -6236 1231 -6235
rect -415 -6282 -367 -6236
rect -321 -6282 -273 -6236
rect -227 -6282 -179 -6236
rect -133 -6282 -85 -6236
rect -39 -6282 9 -6236
rect 55 -6282 103 -6236
rect 149 -6282 197 -6236
rect 243 -6282 291 -6236
rect 337 -6282 385 -6236
rect 431 -6282 479 -6236
rect 525 -6282 573 -6236
rect 619 -6282 667 -6236
rect 713 -6282 761 -6236
rect 807 -6282 855 -6236
rect 901 -6282 949 -6236
rect 995 -6282 1043 -6236
rect 1089 -6282 1137 -6236
rect 1183 -6282 1231 -6236
rect 1278 -6282 1293 -6235
rect -477 -6297 1293 -6282
rect -3282 -6321 -1230 -6306
<< psubdiffcont >>
rect -549 -6558 -503 -6512
rect -451 -6558 -405 -6512
rect -353 -6558 -307 -6512
rect -255 -6558 -209 -6512
rect -157 -6558 -111 -6512
rect -59 -6558 -13 -6512
rect 39 -6558 85 -6512
rect 137 -6558 183 -6512
rect 235 -6558 281 -6512
rect 333 -6558 379 -6512
rect 431 -6558 477 -6512
rect 529 -6558 575 -6512
rect 627 -6558 673 -6512
rect 725 -6558 771 -6512
rect 823 -6558 869 -6512
rect 921 -6558 967 -6512
rect 1019 -6558 1065 -6512
rect 1117 -6558 1163 -6512
rect 1215 -6558 1261 -6512
rect -549 -6656 -503 -6610
rect -549 -6754 -503 -6708
rect -3295 -6888 -3249 -6842
rect -3197 -6888 -3151 -6842
rect -3099 -6888 -3053 -6842
rect -3001 -6888 -2955 -6842
rect -2903 -6888 -2857 -6842
rect -2805 -6888 -2759 -6842
rect -2707 -6888 -2661 -6842
rect -2609 -6888 -2563 -6842
rect -2511 -6888 -2465 -6842
rect -2413 -6888 -2367 -6842
rect -2315 -6888 -2269 -6842
rect -2217 -6888 -2171 -6842
rect -2119 -6888 -2073 -6842
rect -2021 -6888 -1975 -6842
rect -1923 -6888 -1877 -6842
rect -1825 -6888 -1779 -6842
rect -1727 -6888 -1681 -6842
rect -1629 -6888 -1583 -6842
rect -1531 -6888 -1485 -6842
rect -1433 -6888 -1387 -6842
rect -1335 -6888 -1289 -6842
rect -1237 -6888 -1191 -6842
rect -3295 -6986 -3249 -6940
rect -3295 -7084 -3249 -7038
rect -1237 -6986 -1191 -6940
rect -3295 -7182 -3249 -7136
rect -1237 -7084 -1191 -7038
rect -3295 -7280 -3249 -7234
rect -3295 -7378 -3249 -7332
rect -3295 -7476 -3249 -7430
rect -3295 -7574 -3249 -7528
rect -3295 -7672 -3249 -7626
rect -3295 -7770 -3249 -7724
rect -1237 -7182 -1191 -7136
rect -1237 -7280 -1191 -7234
rect -1237 -7378 -1191 -7332
rect -1237 -7476 -1191 -7430
rect -1237 -7574 -1191 -7528
rect -1237 -7672 -1191 -7626
rect -3295 -7868 -3249 -7822
rect -1237 -7770 -1191 -7724
rect -3295 -7966 -3249 -7920
rect -1237 -7868 -1191 -7822
rect -3295 -8064 -3249 -8018
rect -3295 -8162 -3249 -8116
rect -3295 -8260 -3249 -8214
rect -3295 -8358 -3249 -8312
rect -3295 -8456 -3249 -8410
rect -3295 -8554 -3249 -8508
rect -1237 -7966 -1191 -7920
rect -1237 -8064 -1191 -8018
rect -1237 -8162 -1191 -8116
rect -1237 -8260 -1191 -8214
rect -1237 -8358 -1191 -8312
rect -1237 -8456 -1191 -8410
rect -3295 -8652 -3249 -8606
rect -1237 -8554 -1191 -8508
rect -3295 -8750 -3249 -8704
rect -1237 -8652 -1191 -8606
rect -3295 -8848 -3249 -8802
rect -3295 -8946 -3249 -8900
rect -3295 -9044 -3249 -8998
rect -3295 -9142 -3249 -9096
rect -3295 -9240 -3249 -9194
rect -3295 -9338 -3249 -9292
rect -1237 -8750 -1191 -8704
rect -1237 -8848 -1191 -8802
rect -1237 -8946 -1191 -8900
rect -1237 -9044 -1191 -8998
rect -1237 -9142 -1191 -9096
rect -1237 -9240 -1191 -9194
rect -3295 -9436 -3249 -9390
rect -1237 -9338 -1191 -9292
rect -3295 -9534 -3249 -9488
rect -1237 -9436 -1191 -9390
rect -1237 -9534 -1191 -9488
rect -3295 -9632 -3249 -9586
rect -3295 -9730 -3249 -9684
rect -3295 -9828 -3249 -9782
rect -3295 -9926 -3249 -9880
rect -3295 -10024 -3249 -9978
rect -3295 -10122 -3249 -10076
rect -1237 -9632 -1191 -9586
rect -1237 -9730 -1191 -9684
rect -1237 -9828 -1191 -9782
rect -1237 -9926 -1191 -9880
rect -1237 -10024 -1191 -9978
rect -1237 -10122 -1191 -10076
rect -3295 -10220 -3249 -10174
rect -3295 -10318 -3249 -10272
rect -1237 -10220 -1191 -10174
rect -1237 -10318 -1191 -10272
rect -3295 -10416 -3249 -10370
rect -3197 -10416 -3151 -10370
rect -3099 -10416 -3053 -10370
rect -3001 -10416 -2955 -10370
rect -2903 -10416 -2857 -10370
rect -2805 -10416 -2759 -10370
rect -2707 -10416 -2661 -10370
rect -2609 -10416 -2563 -10370
rect -2511 -10416 -2465 -10370
rect -2413 -10416 -2367 -10370
rect -2315 -10416 -2269 -10370
rect -2217 -10416 -2171 -10370
rect -2119 -10416 -2073 -10370
rect -2021 -10416 -1975 -10370
rect -1923 -10416 -1877 -10370
rect -1825 -10416 -1779 -10370
rect -1727 -10416 -1681 -10370
rect -1629 -10416 -1583 -10370
rect -1531 -10416 -1485 -10370
rect -1433 -10416 -1387 -10370
rect -1335 -10416 -1289 -10370
rect -1237 -10416 -1191 -10370
rect -549 -6852 -503 -6806
rect 1215 -6656 1261 -6610
rect 1215 -6754 1261 -6708
rect -549 -6950 -503 -6904
rect 1215 -6852 1261 -6806
rect -549 -7048 -503 -7002
rect -549 -7146 -503 -7100
rect -549 -7244 -503 -7198
rect -549 -7342 -503 -7296
rect -549 -7440 -503 -7394
rect -549 -7538 -503 -7492
rect -549 -7636 -503 -7590
rect 1215 -6950 1261 -6904
rect 1215 -7048 1261 -7002
rect 1215 -7146 1261 -7100
rect 1215 -7244 1261 -7198
rect 1215 -7342 1261 -7296
rect 1215 -7440 1261 -7394
rect 1215 -7538 1261 -7492
rect -549 -7734 -503 -7688
rect -549 -7832 -503 -7786
rect 1215 -7636 1261 -7590
rect 1215 -7734 1261 -7688
rect -549 -7930 -503 -7884
rect -549 -8028 -503 -7982
rect -549 -8126 -503 -8080
rect -549 -8224 -503 -8178
rect -549 -8322 -503 -8276
rect -549 -8420 -503 -8374
rect -549 -8518 -503 -8472
rect 1215 -7832 1261 -7786
rect 1215 -7930 1261 -7884
rect 1215 -8028 1261 -7982
rect 1215 -8126 1261 -8080
rect 1215 -8224 1261 -8178
rect 1215 -8322 1261 -8276
rect 3076 -8294 4649 -8156
rect 1215 -8420 1261 -8374
rect -549 -8616 -503 -8570
rect -549 -8714 -503 -8668
rect -549 -8812 -503 -8766
rect 1215 -8518 1261 -8472
rect 1215 -8616 1261 -8570
rect 1215 -8714 1261 -8668
rect -549 -8910 -503 -8864
rect -549 -9008 -503 -8962
rect -549 -9106 -503 -9060
rect -549 -9204 -503 -9158
rect -549 -9302 -503 -9256
rect -549 -9400 -503 -9354
rect -549 -9498 -503 -9452
rect 1215 -8812 1261 -8766
rect 1215 -8910 1261 -8864
rect 1215 -9008 1261 -8962
rect 1215 -9106 1261 -9060
rect 1215 -9204 1261 -9158
rect 1215 -9302 1261 -9256
rect 1215 -9400 1261 -9354
rect -549 -9596 -503 -9550
rect 1215 -9498 1261 -9452
rect 1215 -9596 1261 -9550
rect -549 -9694 -503 -9648
rect -549 -9792 -503 -9746
rect -549 -9890 -503 -9844
rect -549 -9988 -503 -9942
rect -549 -10086 -503 -10040
rect -549 -10184 -503 -10138
rect -549 -10282 -503 -10236
rect 1215 -9694 1261 -9648
rect 1215 -9792 1261 -9746
rect 1215 -9890 1261 -9844
rect 1215 -9988 1261 -9942
rect 1215 -10086 1261 -10040
rect 1215 -10184 1261 -10138
rect 1215 -10282 1261 -10236
rect -549 -10380 -503 -10334
rect 1215 -10380 1261 -10334
rect -549 -10478 -503 -10432
rect -549 -10576 -503 -10530
rect 1215 -10478 1261 -10432
rect 1215 -10576 1261 -10530
rect -549 -10674 -503 -10628
rect -451 -10674 -405 -10628
rect -353 -10674 -307 -10628
rect -255 -10674 -209 -10628
rect -157 -10674 -111 -10628
rect -59 -10674 -13 -10628
rect 39 -10674 85 -10628
rect 137 -10674 183 -10628
rect 235 -10674 281 -10628
rect 333 -10674 379 -10628
rect 431 -10674 477 -10628
rect 529 -10674 575 -10628
rect 627 -10674 673 -10628
rect 725 -10674 771 -10628
rect 823 -10674 869 -10628
rect 921 -10674 967 -10628
rect 1019 -10674 1065 -10628
rect 1117 -10674 1163 -10628
rect 1215 -10674 1261 -10628
<< nsubdiffcont >>
rect -3294 1394 -3247 1441
rect -3199 1395 -3153 1441
rect -3105 1395 -3059 1441
rect -3011 1395 -2965 1441
rect -2917 1395 -2871 1441
rect -2823 1395 -2777 1441
rect -2729 1395 -2683 1441
rect -2635 1395 -2589 1441
rect -2541 1395 -2495 1441
rect -2447 1395 -2401 1441
rect -2353 1395 -2307 1441
rect -2259 1395 -2213 1441
rect -2165 1395 -2119 1441
rect -2071 1395 -2025 1441
rect -1977 1395 -1931 1441
rect -1883 1395 -1837 1441
rect -1789 1395 -1743 1441
rect -1695 1395 -1649 1441
rect -1601 1395 -1555 1441
rect -1507 1395 -1461 1441
rect -1413 1395 -1367 1441
rect -1319 1394 -1272 1441
rect -3294 1300 -3248 1346
rect -1318 1300 -1272 1346
rect -3294 1206 -3248 1252
rect -1318 1206 -1272 1252
rect -3294 1112 -3248 1158
rect -3294 1018 -3248 1064
rect -3294 924 -3248 970
rect -3294 830 -3248 876
rect -3294 736 -3248 782
rect -3294 642 -3248 688
rect -3294 548 -3248 594
rect -1318 1112 -1272 1158
rect -1318 1018 -1272 1064
rect -1318 924 -1272 970
rect -1318 830 -1272 876
rect -1318 736 -1272 782
rect -1318 642 -1272 688
rect -1318 548 -1272 594
rect -3294 454 -3248 500
rect -1318 454 -1272 500
rect -3294 360 -3248 406
rect -3294 266 -3248 312
rect -3294 172 -3248 218
rect -3294 78 -3248 124
rect -3294 -16 -3248 30
rect -3294 -110 -3248 -64
rect -3294 -204 -3248 -158
rect -1318 360 -1272 406
rect -1318 266 -1272 312
rect -1318 172 -1272 218
rect -1318 78 -1272 124
rect -1318 -16 -1272 30
rect -1318 -110 -1272 -64
rect -1318 -204 -1272 -158
rect -3294 -298 -3248 -252
rect -3294 -392 -3248 -346
rect -3294 -486 -3248 -440
rect -3294 -580 -3248 -534
rect -3294 -674 -3248 -628
rect -3294 -768 -3248 -722
rect -3294 -862 -3248 -816
rect -3294 -956 -3248 -910
rect -1318 -298 -1272 -252
rect -1318 -392 -1272 -346
rect -1318 -486 -1272 -440
rect -1318 -580 -1272 -534
rect -1318 -674 -1272 -628
rect -1318 -768 -1272 -722
rect -1318 -862 -1272 -816
rect -3294 -1050 -3248 -1004
rect -1318 -956 -1272 -910
rect -3294 -1144 -3248 -1098
rect -3294 -1238 -3248 -1192
rect -3294 -1332 -3248 -1286
rect -3294 -1426 -3248 -1380
rect -3294 -1520 -3248 -1474
rect -3294 -1614 -3248 -1568
rect -3294 -1708 -3248 -1662
rect -3294 -1802 -3248 -1756
rect -3294 -1896 -3248 -1850
rect -1318 -1050 -1272 -1004
rect -1318 -1144 -1272 -1098
rect -1318 -1238 -1272 -1192
rect -1318 -1332 -1272 -1286
rect -1318 -1426 -1272 -1380
rect -1318 -1520 -1272 -1474
rect -1318 -1614 -1272 -1568
rect -1318 -1708 -1272 -1662
rect -1318 -1802 -1272 -1756
rect -1318 -1896 -1272 -1850
rect -3293 -1990 -3247 -1944
rect -3199 -1990 -3153 -1944
rect -3105 -1990 -3059 -1944
rect -3011 -1990 -2965 -1944
rect -2917 -1990 -2871 -1944
rect -2823 -1990 -2777 -1944
rect -2729 -1990 -2683 -1944
rect -2635 -1990 -2589 -1944
rect -2541 -1990 -2495 -1944
rect -2447 -1990 -2401 -1944
rect -2353 -1990 -2307 -1944
rect -2259 -1990 -2213 -1944
rect -2165 -1990 -2119 -1944
rect -2071 -1990 -2025 -1944
rect -1977 -1990 -1931 -1944
rect -1883 -1990 -1837 -1944
rect -1789 -1990 -1743 -1944
rect -1695 -1990 -1649 -1944
rect -1601 -1990 -1555 -1944
rect -1507 -1990 -1461 -1944
rect -1413 -1990 -1367 -1944
rect -1319 -1990 -1273 -1944
rect -747 967 -701 1013
rect -653 967 -607 1013
rect -552 967 -506 1013
rect -458 967 -412 1013
rect -362 967 -316 1013
rect -268 967 -222 1013
rect -167 967 -121 1013
rect -73 967 -27 1013
rect 21 967 67 1013
rect 115 967 161 1013
rect 216 967 262 1013
rect 310 967 356 1013
rect 406 967 452 1013
rect 500 967 546 1013
rect 601 967 647 1013
rect 695 967 741 1013
rect 789 967 835 1013
rect 883 967 929 1013
rect 984 967 1030 1013
rect 1078 967 1124 1013
rect 1172 967 1218 1013
rect -747 871 -701 917
rect 1172 871 1218 917
rect -747 777 -701 823
rect 1172 770 1218 816
rect -747 681 -701 727
rect -747 587 -701 633
rect -747 493 -701 539
rect -747 392 -701 438
rect -747 298 -701 344
rect -747 202 -701 248
rect -747 108 -701 154
rect 1172 676 1218 722
rect 1172 582 1218 628
rect 1172 488 1218 534
rect 1172 387 1218 433
rect 1172 293 1218 339
rect 1172 197 1218 243
rect 1172 103 1218 149
rect -747 7 -701 53
rect -747 -87 -701 -41
rect -747 -181 -701 -135
rect -747 -275 -701 -229
rect 1172 2 1218 48
rect 1172 -92 1218 -46
rect 1172 -186 1218 -140
rect 1172 -280 1218 -234
rect -747 -376 -701 -330
rect -747 -470 -701 -424
rect -747 -566 -701 -520
rect -747 -660 -701 -614
rect -747 -761 -701 -715
rect -747 -855 -701 -809
rect -747 -949 -701 -903
rect 1172 -381 1218 -335
rect 1172 -475 1218 -429
rect 1172 -571 1218 -525
rect 1172 -665 1218 -619
rect 1172 -766 1218 -720
rect 1172 -860 1218 -814
rect 1172 -954 1218 -908
rect -747 -1043 -701 -997
rect -747 -1144 -701 -1098
rect -747 -1238 -701 -1192
rect -747 -1334 -701 -1288
rect 1172 -1050 1218 -1004
rect 1172 -1144 1218 -1098
rect 1172 -1245 1218 -1199
rect -747 -1428 -701 -1382
rect -747 -1522 -701 -1476
rect -747 -1623 -701 -1577
rect -747 -1717 -701 -1671
rect -747 -1813 -701 -1767
rect -747 -1907 -701 -1861
rect -747 -2008 -701 -1962
rect 1172 -1339 1218 -1293
rect 1172 -1433 1218 -1387
rect 1172 -1527 1218 -1481
rect 1172 -1628 1218 -1582
rect 1172 -1722 1218 -1676
rect 1172 -1818 1218 -1772
rect 1172 -1912 1218 -1866
rect -747 -2102 -701 -2056
rect -747 -2196 -701 -2150
rect -747 -2290 -701 -2244
rect -747 -2391 -701 -2345
rect 1172 -2013 1218 -1967
rect 1172 -2107 1218 -2061
rect 1172 -2201 1218 -2155
rect 1172 -2295 1218 -2249
rect -747 -2485 -701 -2439
rect -3267 -2640 -3220 -2593
rect -3172 -2639 -3126 -2593
rect -3078 -2639 -3032 -2593
rect -2984 -2639 -2938 -2593
rect -2890 -2639 -2844 -2593
rect -2796 -2639 -2750 -2593
rect -2702 -2639 -2656 -2593
rect -2608 -2639 -2562 -2593
rect -2514 -2639 -2468 -2593
rect -2420 -2639 -2374 -2593
rect -2326 -2639 -2280 -2593
rect -2232 -2639 -2186 -2593
rect -2138 -2639 -2092 -2593
rect -2044 -2639 -1998 -2593
rect -1950 -2639 -1904 -2593
rect -1856 -2639 -1810 -2593
rect -1762 -2639 -1716 -2593
rect -1668 -2639 -1622 -2593
rect -1574 -2639 -1528 -2593
rect -1480 -2639 -1434 -2593
rect -1386 -2639 -1340 -2593
rect -1292 -2640 -1245 -2593
rect -3267 -2734 -3221 -2688
rect -3267 -2828 -3221 -2782
rect -1291 -2734 -1245 -2688
rect -1291 -2828 -1245 -2782
rect -3267 -2922 -3221 -2876
rect -3267 -3016 -3221 -2970
rect -3267 -3110 -3221 -3064
rect -3267 -3204 -3221 -3158
rect -3267 -3298 -3221 -3252
rect -3267 -3392 -3221 -3346
rect -3267 -3486 -3221 -3440
rect -1291 -2922 -1245 -2876
rect -1291 -3016 -1245 -2970
rect -1291 -3110 -1245 -3064
rect -1291 -3204 -1245 -3158
rect -1291 -3298 -1245 -3252
rect -1291 -3392 -1245 -3346
rect -747 -2581 -701 -2535
rect -747 -2675 -701 -2629
rect -747 -2776 -701 -2730
rect -747 -2870 -701 -2824
rect -747 -2964 -701 -2918
rect -747 -3058 -701 -3012
rect 1172 -2396 1218 -2350
rect 1172 -2490 1218 -2444
rect 1172 -2586 1218 -2540
rect 1172 -2680 1218 -2634
rect 1172 -2781 1218 -2735
rect 1172 -2875 1218 -2829
rect 1172 -2969 1218 -2923
rect -747 -3159 -701 -3113
rect 1172 -3065 1218 -3019
rect 1172 -3159 1218 -3113
rect -747 -3253 -701 -3207
rect 1172 -3253 1218 -3207
rect -747 -3349 -701 -3303
rect -653 -3349 -607 -3303
rect -552 -3349 -506 -3303
rect -458 -3349 -412 -3303
rect -362 -3349 -316 -3303
rect -268 -3349 -222 -3303
rect -167 -3349 -121 -3303
rect -73 -3349 -27 -3303
rect 21 -3349 67 -3303
rect 115 -3349 161 -3303
rect 216 -3349 262 -3303
rect 310 -3349 356 -3303
rect 406 -3349 452 -3303
rect 500 -3349 546 -3303
rect 601 -3349 647 -3303
rect 695 -3349 741 -3303
rect 789 -3349 835 -3303
rect 883 -3349 929 -3303
rect 984 -3349 1030 -3303
rect 1078 -3349 1124 -3303
rect 1172 -3349 1218 -3303
rect -1291 -3486 -1245 -3440
rect -3267 -3580 -3221 -3534
rect -3267 -3674 -3221 -3628
rect -1291 -3580 -1245 -3534
rect -1291 -3674 -1245 -3628
rect -3267 -3768 -3221 -3722
rect -3267 -3862 -3221 -3816
rect -3267 -3956 -3221 -3910
rect -1291 -3768 -1245 -3722
rect -1291 -3862 -1245 -3816
rect -1291 -3956 -1245 -3910
rect -3267 -4050 -3221 -4004
rect -3267 -4144 -3221 -4098
rect -3267 -4238 -3221 -4192
rect -3267 -4332 -3221 -4286
rect -1291 -4050 -1245 -4004
rect -1291 -4144 -1245 -4098
rect -1291 -4238 -1245 -4192
rect -1291 -4332 -1245 -4286
rect -3267 -4426 -3221 -4380
rect -3267 -4520 -3221 -4474
rect -1291 -4426 -1245 -4380
rect -3267 -4614 -3221 -4568
rect -1291 -4520 -1245 -4474
rect -3267 -4708 -3221 -4662
rect -3267 -4802 -3221 -4756
rect -3267 -4896 -3221 -4850
rect -3267 -4990 -3221 -4944
rect -3267 -5084 -3221 -5038
rect -3267 -5178 -3221 -5132
rect -1291 -4614 -1245 -4568
rect -1291 -4708 -1245 -4662
rect -1291 -4802 -1245 -4756
rect -1291 -4896 -1245 -4850
rect -1291 -4990 -1245 -4944
rect -1291 -5084 -1245 -5038
rect -3267 -5272 -3221 -5226
rect -1291 -5178 -1245 -5132
rect -3267 -5366 -3221 -5320
rect -1291 -5272 -1245 -5226
rect -3267 -5460 -3221 -5414
rect -1291 -5366 -1245 -5320
rect -3267 -5554 -3221 -5508
rect -3267 -5648 -3221 -5602
rect -3267 -5742 -3221 -5696
rect -3267 -5836 -3221 -5790
rect -3267 -5930 -3221 -5884
rect -3267 -6024 -3221 -5978
rect -1291 -5460 -1245 -5414
rect -1291 -5554 -1245 -5508
rect -1291 -5648 -1245 -5602
rect -1291 -5742 -1245 -5696
rect -1291 -5836 -1245 -5790
rect -1291 -5930 -1245 -5884
rect -3267 -6118 -3221 -6072
rect -1291 -6024 -1245 -5978
rect -1291 -6118 -1245 -6072
rect -3267 -6212 -3221 -6166
rect -1291 -6212 -1245 -6166
rect -3266 -6306 -3220 -6260
rect -3172 -6306 -3126 -6260
rect -3078 -6306 -3032 -6260
rect -2984 -6306 -2938 -6260
rect -2890 -6306 -2844 -6260
rect -2796 -6306 -2750 -6260
rect -2702 -6306 -2656 -6260
rect -2608 -6306 -2562 -6260
rect -2514 -6306 -2468 -6260
rect -2420 -6306 -2374 -6260
rect -2326 -6306 -2280 -6260
rect -2232 -6306 -2186 -6260
rect -2138 -6306 -2092 -6260
rect -2044 -6306 -1998 -6260
rect -1950 -6306 -1904 -6260
rect -1856 -6306 -1810 -6260
rect -1762 -6306 -1716 -6260
rect -1668 -6306 -1622 -6260
rect -1574 -6306 -1528 -6260
rect -1480 -6306 -1434 -6260
rect -1386 -6306 -1340 -6260
rect -1292 -6306 -1246 -6260
rect -462 -4115 -415 -4068
rect -367 -4114 -321 -4068
rect -273 -4114 -227 -4068
rect -179 -4114 -133 -4068
rect -85 -4114 -39 -4068
rect 9 -4114 55 -4068
rect 103 -4114 149 -4068
rect 197 -4114 243 -4068
rect 291 -4114 337 -4068
rect 385 -4114 431 -4068
rect 479 -4114 525 -4068
rect 573 -4114 619 -4068
rect 667 -4114 713 -4068
rect 761 -4114 807 -4068
rect 855 -4114 901 -4068
rect 949 -4114 995 -4068
rect 1043 -4114 1089 -4068
rect 1137 -4114 1183 -4068
rect 1231 -4115 1278 -4068
rect -462 -4213 -416 -4163
rect 1232 -4213 1278 -4163
rect -462 -4307 -416 -4261
rect -462 -4401 -416 -4355
rect 1232 -4307 1278 -4261
rect 1232 -4401 1278 -4355
rect -462 -4495 -416 -4449
rect -462 -4589 -416 -4543
rect -462 -4683 -416 -4637
rect -462 -4777 -416 -4731
rect -462 -4871 -416 -4825
rect -462 -4965 -416 -4919
rect -462 -5059 -416 -5013
rect -462 -5153 -416 -5107
rect 1232 -4495 1278 -4449
rect 1232 -4589 1278 -4543
rect 1232 -4683 1278 -4637
rect 1232 -4777 1278 -4731
rect 1232 -4871 1278 -4825
rect 1232 -4965 1278 -4919
rect 1232 -5059 1278 -5013
rect -462 -5247 -416 -5201
rect 1232 -5153 1278 -5107
rect -462 -5341 -416 -5295
rect -462 -5435 -416 -5389
rect -462 -5529 -416 -5483
rect -462 -5623 -416 -5577
rect -462 -5717 -416 -5671
rect -462 -5811 -416 -5765
rect -462 -5905 -416 -5859
rect -462 -5999 -416 -5953
rect -462 -6093 -416 -6047
rect -462 -6187 -416 -6141
rect 1232 -5247 1278 -5201
rect 1232 -5341 1278 -5295
rect 1232 -5435 1278 -5389
rect 1232 -5529 1278 -5483
rect 1232 -5623 1278 -5577
rect 1232 -5717 1278 -5671
rect 3066 -5693 4667 -5557
rect 1232 -5811 1278 -5765
rect 1232 -5905 1278 -5859
rect 1232 -5999 1278 -5953
rect 1232 -6093 1278 -6047
rect 1232 -6187 1278 -6141
rect -462 -6282 -415 -6235
rect -367 -6282 -321 -6236
rect -273 -6282 -227 -6236
rect -179 -6282 -133 -6236
rect -85 -6282 -39 -6236
rect 9 -6282 55 -6236
rect 103 -6282 149 -6236
rect 197 -6282 243 -6236
rect 291 -6282 337 -6236
rect 385 -6282 431 -6236
rect 479 -6282 525 -6236
rect 573 -6282 619 -6236
rect 667 -6282 713 -6236
rect 761 -6282 807 -6236
rect 855 -6282 901 -6236
rect 949 -6282 995 -6236
rect 1043 -6282 1089 -6236
rect 1137 -6282 1183 -6236
rect 1231 -6282 1278 -6235
<< polysilicon >>
rect -2679 1260 -1919 1276
rect -2679 1214 -2323 1260
rect -2277 1214 -1919 1260
rect -2679 1192 -1919 1214
rect -2679 507 -1919 517
rect -2895 504 -2783 505
rect -2895 458 -2864 504
rect -2818 458 -2783 504
rect -2895 457 -2783 458
rect -2679 461 -2428 507
rect -2382 504 -1919 507
rect -2382 461 -2215 504
rect -2679 457 -2215 461
rect -2167 457 -1919 504
rect -1815 504 -1703 505
rect -1815 458 -1782 504
rect -1736 458 -1703 504
rect -1815 457 -1703 458
rect -2679 444 -1919 457
rect -2895 -232 -2783 -231
rect -2895 -278 -2864 -232
rect -2818 -278 -2783 -232
rect -2895 -279 -2783 -278
rect -2679 -232 -1919 -219
rect -2679 -278 -2428 -232
rect -2382 -278 -2215 -232
rect -2679 -279 -2215 -278
rect -2167 -279 -1919 -232
rect -1815 -232 -1703 -231
rect -1815 -278 -1781 -232
rect -1735 -278 -1703 -232
rect -1815 -279 -1703 -278
rect -2679 -292 -1919 -279
rect -2895 -968 -2783 -967
rect -2895 -1014 -2863 -968
rect -2817 -1014 -2783 -968
rect -2895 -1015 -2783 -1014
rect -2679 -970 -1919 -955
rect -2679 -971 -2215 -970
rect -2679 -1017 -2428 -971
rect -2382 -1017 -2215 -971
rect -2167 -1017 -1919 -970
rect -1815 -968 -1703 -967
rect -1815 -1014 -1781 -968
rect -1735 -1014 -1703 -968
rect -1815 -1015 -1703 -1014
rect -2679 -1028 -1919 -1017
rect -365 842 -253 863
rect -365 796 -336 842
rect -290 796 -253 842
rect -365 758 -253 796
rect 715 844 827 864
rect 715 798 750 844
rect 796 798 827 844
rect 715 758 827 798
rect -149 -7 -37 70
rect 67 -7 179 70
rect 283 -7 395 70
rect 499 -7 611 70
rect -149 -60 611 -7
rect -149 -106 99 -60
rect 145 -106 611 -60
rect -149 -153 611 -106
rect -149 -280 -37 -153
rect 67 -280 179 -153
rect 283 -280 395 -153
rect 499 -280 611 -153
rect -365 -1122 -253 -968
rect -365 -1170 -330 -1122
rect -283 -1170 -253 -1122
rect -365 -1320 -253 -1170
rect -149 -1080 -37 -968
rect 67 -1080 179 -968
rect 283 -1080 395 -968
rect 499 -1080 611 -968
rect -149 -1135 611 -1080
rect -149 -1181 99 -1135
rect 145 -1181 611 -1135
rect -149 -1226 611 -1181
rect -149 -1320 -37 -1226
rect 67 -1320 179 -1226
rect 283 -1320 395 -1226
rect 499 -1320 611 -1226
rect 715 -1123 827 -968
rect 715 -1169 752 -1123
rect 798 -1169 827 -1123
rect 715 -1320 827 -1169
rect -149 -2117 -37 -2008
rect 67 -2117 179 -2008
rect 283 -2117 395 -2008
rect 499 -2117 611 -2008
rect -149 -2171 611 -2117
rect -149 -2217 130 -2171
rect 176 -2217 611 -2171
rect -149 -2263 611 -2217
rect -149 -2358 -37 -2263
rect 67 -2358 179 -2263
rect 283 -2358 395 -2263
rect 499 -2358 611 -2263
rect -2849 -2747 -2762 -2733
rect -2849 -2793 -2828 -2747
rect -2782 -2793 -2762 -2747
rect -2849 -2813 -2762 -2793
rect -2370 -2747 -2283 -2731
rect -2370 -2793 -2348 -2747
rect -2302 -2793 -2283 -2747
rect -2370 -2811 -2283 -2793
rect -2207 -2747 -2120 -2731
rect -2207 -2793 -2188 -2747
rect -2142 -2793 -2120 -2747
rect -2207 -2811 -2120 -2793
rect -1728 -2747 -1642 -2733
rect -1728 -2793 -1708 -2747
rect -1662 -2793 -1642 -2747
rect -2833 -2865 -2777 -2813
rect -2353 -2821 -2297 -2811
rect -2193 -2821 -2137 -2811
rect -1728 -2813 -1642 -2793
rect -1713 -2865 -1657 -2813
rect -365 -3132 -253 -3045
rect -365 -3184 -333 -3132
rect -276 -3184 -253 -3132
rect -365 -3206 -253 -3184
rect 715 -3128 827 -3046
rect 715 -3182 738 -3128
rect 796 -3182 827 -3128
rect 715 -3202 827 -3182
rect -3077 -3534 -2937 -3509
rect -3077 -3580 -3061 -3534
rect -3015 -3580 -2937 -3534
rect -2673 -3542 -2617 -3497
rect -2513 -3542 -2457 -3497
rect -2033 -3542 -1977 -3497
rect -1873 -3542 -1817 -3497
rect -1553 -3525 -1403 -3509
rect -2684 -3559 -2606 -3542
rect -3077 -3595 -2937 -3580
rect -2845 -3580 -2767 -3563
rect -2845 -3626 -2829 -3580
rect -2783 -3626 -2767 -3580
rect -2684 -3605 -2668 -3559
rect -2622 -3605 -2606 -3559
rect -2684 -3619 -2606 -3605
rect -2524 -3558 -2446 -3542
rect -2524 -3604 -2508 -3558
rect -2462 -3604 -2446 -3558
rect -2044 -3558 -1966 -3542
rect -2524 -3619 -2446 -3604
rect -2363 -3577 -2285 -3563
rect -2845 -3640 -2767 -3626
rect -2363 -3623 -2348 -3577
rect -2302 -3623 -2285 -3577
rect -2363 -3640 -2285 -3623
rect -2205 -3577 -2127 -3563
rect -2205 -3623 -2188 -3577
rect -2142 -3623 -2127 -3577
rect -2044 -3604 -2028 -3558
rect -1982 -3604 -1966 -3558
rect -2044 -3619 -1966 -3604
rect -1884 -3559 -1806 -3542
rect -1884 -3605 -1868 -3559
rect -1822 -3605 -1806 -3559
rect -1884 -3619 -1806 -3605
rect -1723 -3580 -1645 -3563
rect -2205 -3640 -2127 -3623
rect -1723 -3626 -1707 -3580
rect -1661 -3626 -1645 -3580
rect -1553 -3571 -1468 -3525
rect -1422 -3571 -1403 -3525
rect -1553 -3596 -1403 -3571
rect -1723 -3640 -1645 -3626
rect -2833 -3685 -2777 -3640
rect -2353 -3685 -2297 -3640
rect -2193 -3685 -2137 -3640
rect -1713 -3685 -1657 -3640
rect -3086 -4380 -2937 -4361
rect -3086 -4426 -3068 -4380
rect -3022 -4426 -2937 -4380
rect -2673 -4402 -2617 -4361
rect -3086 -4453 -2937 -4426
rect -2688 -4420 -2601 -4402
rect -2513 -4403 -2457 -4361
rect -2033 -4403 -1977 -4361
rect -1873 -4402 -1817 -4361
rect -1553 -4381 -1396 -4361
rect -2688 -4466 -2667 -4420
rect -2621 -4466 -2601 -4420
rect -2688 -4484 -2601 -4466
rect -2529 -4420 -2442 -4403
rect -2529 -4466 -2507 -4420
rect -2461 -4466 -2442 -4420
rect -2529 -4483 -2442 -4466
rect -2048 -4420 -1961 -4403
rect -2048 -4466 -2029 -4420
rect -1983 -4466 -1961 -4420
rect -2048 -4483 -1961 -4466
rect -1889 -4420 -1802 -4402
rect -1889 -4466 -1869 -4420
rect -1823 -4466 -1802 -4420
rect -1553 -4427 -1468 -4381
rect -1422 -4427 -1396 -4381
rect -1553 -4448 -1396 -4427
rect -2993 -4569 -2937 -4525
rect -2833 -4569 -2777 -4525
rect -2673 -4569 -2617 -4484
rect -2513 -4569 -2457 -4483
rect -2353 -4569 -2297 -4525
rect -2193 -4569 -2137 -4525
rect -2033 -4569 -1977 -4483
rect -1889 -4484 -1802 -4466
rect -1873 -4569 -1817 -4484
rect -1713 -4569 -1657 -4525
rect -1553 -4569 -1497 -4525
rect -2993 -5213 -2937 -5169
rect -3083 -5231 -2937 -5213
rect -3083 -5277 -3068 -5231
rect -3022 -5277 -2937 -5231
rect -2833 -5246 -2777 -5169
rect -2673 -5213 -2617 -5169
rect -2513 -5213 -2457 -5169
rect -2353 -5246 -2297 -5169
rect -2193 -5246 -2137 -5169
rect -2033 -5213 -1977 -5169
rect -1873 -5213 -1817 -5169
rect -1713 -5246 -1657 -5169
rect -1553 -5213 -1497 -5169
rect -1553 -5232 -1403 -5213
rect -3083 -5296 -2937 -5277
rect -2845 -5260 -2767 -5246
rect -2845 -5306 -2829 -5260
rect -2783 -5306 -2767 -5260
rect -2363 -5263 -2285 -5246
rect -2845 -5323 -2767 -5306
rect -2684 -5281 -2606 -5267
rect -2684 -5327 -2668 -5281
rect -2622 -5327 -2606 -5281
rect -2684 -5344 -2606 -5327
rect -2524 -5282 -2446 -5267
rect -2524 -5328 -2508 -5282
rect -2462 -5328 -2446 -5282
rect -2363 -5309 -2348 -5263
rect -2302 -5309 -2285 -5263
rect -2363 -5323 -2285 -5309
rect -2205 -5263 -2127 -5246
rect -2205 -5309 -2188 -5263
rect -2142 -5309 -2127 -5263
rect -1723 -5260 -1645 -5246
rect -2205 -5323 -2127 -5309
rect -2044 -5282 -1966 -5267
rect -2524 -5344 -2446 -5328
rect -2044 -5328 -2028 -5282
rect -1982 -5328 -1966 -5282
rect -2044 -5344 -1966 -5328
rect -1884 -5281 -1806 -5267
rect -1884 -5327 -1868 -5281
rect -1822 -5327 -1806 -5281
rect -1723 -5306 -1707 -5260
rect -1661 -5306 -1645 -5260
rect -1553 -5278 -1468 -5232
rect -1422 -5278 -1403 -5232
rect -1553 -5305 -1403 -5278
rect -1723 -5323 -1645 -5306
rect -1884 -5344 -1806 -5327
rect -2993 -5421 -2937 -5377
rect -2833 -5421 -2777 -5377
rect -2673 -5421 -2617 -5344
rect -2513 -5421 -2457 -5344
rect -2353 -5421 -2297 -5377
rect -2193 -5421 -2137 -5377
rect -2033 -5421 -1977 -5344
rect -1873 -5421 -1817 -5344
rect -1713 -5421 -1657 -5377
rect -1553 -5421 -1497 -5377
rect -2993 -6065 -2937 -6021
rect -3086 -6081 -2937 -6065
rect -2833 -6073 -2777 -6021
rect -2673 -6065 -2617 -6021
rect -2513 -6065 -2457 -6021
rect -3086 -6127 -3068 -6081
rect -3022 -6127 -2937 -6081
rect -3086 -6147 -2937 -6127
rect -2849 -6093 -2762 -6073
rect -2353 -6075 -2297 -6021
rect -2193 -6075 -2137 -6021
rect -2033 -6065 -1977 -6021
rect -1873 -6065 -1817 -6021
rect -1713 -6073 -1657 -6021
rect -1553 -6065 -1497 -6021
rect -2849 -6139 -2828 -6093
rect -2782 -6139 -2762 -6093
rect -2849 -6153 -2762 -6139
rect -2370 -6093 -2283 -6075
rect -2370 -6139 -2348 -6093
rect -2302 -6139 -2283 -6093
rect -2370 -6155 -2283 -6139
rect -2207 -6093 -2120 -6075
rect -2207 -6139 -2188 -6093
rect -2142 -6139 -2120 -6093
rect -2207 -6155 -2120 -6139
rect -1728 -6093 -1641 -6073
rect -1728 -6139 -1708 -6093
rect -1662 -6139 -1641 -6093
rect -1728 -6153 -1641 -6139
rect -1553 -6085 -1403 -6065
rect -1553 -6131 -1468 -6085
rect -1422 -6131 -1403 -6085
rect -1553 -6152 -1403 -6131
rect -168 -4248 80 -4235
rect -168 -4303 -154 -4248
rect -90 -4303 80 -4248
rect -168 -4318 80 -4303
rect -1 -4361 80 -4318
rect -1 -4444 791 -4361
rect -173 -5148 -90 -5132
rect -173 -5194 -156 -5148
rect -110 -5194 -90 -5148
rect -173 -5211 -90 -5194
rect -161 -5224 -105 -5211
rect -1 -5224 791 -5132
rect 895 -5135 951 -5132
rect 884 -5152 967 -5135
rect 884 -5198 901 -5152
rect 947 -5198 967 -5152
rect 884 -5214 967 -5198
rect 895 -5224 951 -5214
rect -3063 -7053 -2918 -7040
rect -3063 -7099 -3049 -7053
rect -3003 -7099 -2918 -7053
rect -1534 -7053 -1389 -7040
rect -3063 -7112 -2918 -7099
rect -2974 -7139 -2918 -7112
rect -2174 -7139 -2118 -7095
rect -2014 -7139 -1958 -7095
rect -1854 -7139 -1798 -7095
rect -1694 -7139 -1638 -7095
rect -1534 -7099 -1449 -7053
rect -1403 -7099 -1389 -7053
rect -1534 -7112 -1389 -7099
rect -1534 -7139 -1478 -7112
rect -2814 -7789 -2758 -7783
rect -2654 -7789 -2598 -7783
rect -2494 -7789 -2438 -7783
rect -2334 -7789 -2278 -7783
rect -2174 -7789 -2118 -7739
rect -2014 -7789 -1958 -7739
rect -1854 -7789 -1798 -7739
rect -1694 -7789 -1638 -7739
rect -1534 -7783 -1478 -7739
rect -2814 -7815 -1638 -7789
rect -3063 -7853 -2918 -7840
rect -3063 -7899 -3049 -7853
rect -3003 -7899 -2918 -7853
rect -2814 -7864 -2251 -7815
rect -2202 -7864 -1638 -7815
rect -2814 -7887 -1638 -7864
rect -2814 -7895 -2758 -7887
rect -2654 -7895 -2598 -7887
rect -2494 -7895 -2438 -7887
rect -2334 -7895 -2278 -7887
rect -3063 -7912 -2918 -7899
rect -2974 -7939 -2918 -7912
rect -2174 -7939 -2118 -7887
rect -2014 -7939 -1958 -7887
rect -1854 -7939 -1798 -7887
rect -1694 -7939 -1638 -7887
rect -1534 -7853 -1389 -7840
rect -1534 -7899 -1449 -7853
rect -1403 -7899 -1389 -7853
rect -1534 -7912 -1389 -7899
rect -1534 -7939 -1478 -7912
rect -2814 -8589 -2758 -8583
rect -2654 -8589 -2598 -8583
rect -2494 -8589 -2438 -8583
rect -2334 -8589 -2278 -8583
rect -2174 -8589 -2118 -8539
rect -2014 -8589 -1958 -8539
rect -1854 -8589 -1798 -8539
rect -1694 -8589 -1638 -8539
rect -1534 -8583 -1478 -8539
rect -2814 -8616 -1638 -8589
rect -3063 -8651 -2918 -8638
rect -3063 -8697 -3049 -8651
rect -3003 -8697 -2918 -8651
rect -3063 -8710 -2918 -8697
rect -2974 -8737 -2918 -8710
rect -2814 -8665 -2251 -8616
rect -2202 -8665 -1638 -8616
rect -2814 -8687 -1638 -8665
rect -2814 -8737 -2758 -8687
rect -2654 -8737 -2598 -8687
rect -2494 -8737 -2438 -8687
rect -2334 -8737 -2278 -8687
rect -2174 -8737 -2118 -8687
rect -2014 -8737 -1958 -8687
rect -1854 -8737 -1798 -8687
rect -1694 -8737 -1638 -8687
rect -1534 -8651 -1389 -8638
rect -1534 -8697 -1449 -8651
rect -1403 -8697 -1389 -8651
rect -1534 -8710 -1389 -8697
rect -1534 -8737 -1478 -8710
rect -2974 -9381 -2918 -9337
rect -2814 -9389 -2758 -9337
rect -2654 -9389 -2598 -9337
rect -2494 -9389 -2438 -9337
rect -2334 -9389 -2278 -9337
rect -2174 -9389 -2118 -9337
rect -2014 -9389 -1958 -9337
rect -1854 -9389 -1798 -9337
rect -1694 -9389 -1638 -9337
rect -1534 -9381 -1478 -9337
rect -2814 -9416 -1638 -9389
rect -3063 -9451 -2918 -9438
rect -3063 -9497 -3049 -9451
rect -3003 -9497 -2918 -9451
rect -3063 -9510 -2918 -9497
rect -2974 -9537 -2918 -9510
rect -2814 -9465 -2252 -9416
rect -2203 -9465 -1638 -9416
rect -2814 -9487 -1638 -9465
rect -2814 -9537 -2758 -9487
rect -2654 -9537 -2598 -9487
rect -2494 -9537 -2438 -9487
rect -2334 -9537 -2278 -9487
rect -2174 -9537 -2118 -9487
rect -2014 -9537 -1958 -9487
rect -1854 -9537 -1798 -9487
rect -1694 -9537 -1638 -9487
rect -1534 -9451 -1389 -9438
rect -1534 -9497 -1449 -9451
rect -1403 -9497 -1389 -9451
rect -1534 -9510 -1389 -9497
rect -1534 -9537 -1478 -9510
rect -2974 -10181 -2918 -10137
rect -2814 -10181 -2758 -10137
rect -2654 -10181 -2598 -10137
rect -2494 -10181 -2438 -10137
rect -2334 -10181 -2278 -10137
rect -2174 -10181 -2118 -10137
rect -2014 -10181 -1958 -10137
rect -1854 -10181 -1798 -10137
rect -1694 -10181 -1638 -10137
rect -1534 -10181 -1478 -10137
rect -262 -6863 -183 -6842
rect -262 -6909 -245 -6863
rect -199 -6909 -183 -6863
rect -262 -6938 -183 -6909
rect 863 -6885 940 -6871
rect 863 -6931 878 -6885
rect 924 -6931 940 -6885
rect 863 -6946 940 -6931
rect 2869 -6927 3083 -6885
rect 3561 -6920 3673 -6886
rect 4225 -6920 4337 -6887
rect 2869 -6979 2893 -6927
rect 2945 -6939 3083 -6927
rect 3515 -6939 3722 -6920
rect 4164 -6939 4337 -6920
rect 2945 -6979 4337 -6939
rect 2869 -7002 4337 -6979
rect 4890 -6912 5105 -6885
rect 4890 -6960 5026 -6912
rect 5082 -6960 5105 -6912
rect 4890 -6997 5105 -6960
rect 2869 -7061 3012 -7002
rect 3086 -7008 4224 -7002
rect 3086 -7061 3582 -7008
rect 2869 -7067 3582 -7061
rect 3656 -7061 4224 -7008
rect 4298 -7061 4337 -7002
rect 3656 -7067 4337 -7061
rect 2869 -7085 4337 -7067
rect 3293 -7410 3500 -7380
rect 3293 -7470 3310 -7410
rect 3363 -7470 3500 -7410
rect 3293 -7492 3500 -7470
rect 3734 -7390 3944 -7377
rect 3734 -7412 4373 -7390
rect 3734 -7471 3754 -7412
rect 3806 -7471 4373 -7412
rect 3734 -7480 4373 -7471
rect 3734 -7493 3944 -7480
rect 4261 -7491 4373 -7480
rect -89 -7645 -33 -7626
rect 232 -7645 288 -7626
rect 392 -7645 448 -7626
rect 713 -7645 769 -7626
rect -89 -7682 769 -7645
rect -260 -7725 -180 -7705
rect -260 -7771 -243 -7725
rect -197 -7771 -180 -7725
rect -260 -7788 -180 -7771
rect -89 -7740 313 -7682
rect 371 -7740 769 -7682
rect -89 -7769 769 -7740
rect -89 -7788 -33 -7769
rect 232 -7788 288 -7769
rect 392 -7788 448 -7769
rect 713 -7788 769 -7769
rect 862 -7743 939 -7729
rect 862 -7789 877 -7743
rect 923 -7789 939 -7743
rect 862 -7803 939 -7789
rect -89 -8562 -33 -8476
rect 232 -8562 288 -8476
rect 392 -8562 448 -8476
rect 713 -8562 769 -8476
rect -89 -8593 984 -8562
rect -89 -8651 908 -8593
rect 966 -8651 984 -8593
rect -89 -8686 984 -8651
rect -89 -8768 -33 -8686
rect 232 -8768 288 -8686
rect 392 -8768 448 -8686
rect 713 -8768 769 -8686
rect -264 -9468 -175 -9453
rect -264 -9514 -243 -9468
rect -197 -9514 -175 -9468
rect -264 -9531 -175 -9514
rect -89 -9475 -33 -9456
rect 232 -9475 288 -9456
rect 392 -9475 448 -9456
rect 713 -9475 769 -9456
rect -89 -9511 769 -9475
rect -89 -9569 304 -9511
rect 362 -9569 769 -9511
rect 858 -9474 948 -9456
rect 858 -9520 880 -9474
rect 926 -9520 948 -9474
rect 858 -9534 948 -9520
rect -89 -9599 769 -9569
rect -89 -9618 -33 -9599
rect 232 -9618 288 -9599
rect 392 -9618 448 -9599
rect 713 -9618 769 -9599
rect -261 -10321 -185 -10306
rect -261 -10367 -246 -10321
rect -200 -10367 -185 -10321
rect -261 -10381 -185 -10367
rect 873 -10329 1019 -10306
rect 873 -10375 957 -10329
rect 1003 -10375 1019 -10329
rect 873 -10396 1019 -10375
<< polycontact >>
rect -2323 1214 -2277 1260
rect -2864 458 -2818 504
rect -2428 461 -2382 507
rect -2215 457 -2167 504
rect -1782 458 -1736 504
rect -2864 -278 -2818 -232
rect -2428 -278 -2382 -232
rect -2215 -279 -2167 -232
rect -1781 -278 -1735 -232
rect -2863 -1014 -2817 -968
rect -2428 -1017 -2382 -971
rect -2215 -1017 -2167 -970
rect -1781 -1014 -1735 -968
rect -336 796 -290 842
rect 750 798 796 844
rect 99 -106 145 -60
rect -330 -1170 -283 -1122
rect 99 -1181 145 -1135
rect 752 -1169 798 -1123
rect 130 -2217 176 -2171
rect -2828 -2793 -2782 -2747
rect -2348 -2793 -2302 -2747
rect -2188 -2793 -2142 -2747
rect -1708 -2793 -1662 -2747
rect -333 -3184 -276 -3132
rect 738 -3182 796 -3128
rect -3061 -3580 -3015 -3534
rect -2829 -3626 -2783 -3580
rect -2668 -3605 -2622 -3559
rect -2508 -3604 -2462 -3558
rect -2348 -3623 -2302 -3577
rect -2188 -3623 -2142 -3577
rect -2028 -3604 -1982 -3558
rect -1868 -3605 -1822 -3559
rect -1707 -3626 -1661 -3580
rect -1468 -3571 -1422 -3525
rect -3068 -4426 -3022 -4380
rect -2667 -4466 -2621 -4420
rect -2507 -4466 -2461 -4420
rect -2029 -4466 -1983 -4420
rect -1869 -4466 -1823 -4420
rect -1468 -4427 -1422 -4381
rect -3068 -5277 -3022 -5231
rect -2829 -5306 -2783 -5260
rect -2668 -5327 -2622 -5281
rect -2508 -5328 -2462 -5282
rect -2348 -5309 -2302 -5263
rect -2188 -5309 -2142 -5263
rect -2028 -5328 -1982 -5282
rect -1868 -5327 -1822 -5281
rect -1707 -5306 -1661 -5260
rect -1468 -5278 -1422 -5232
rect -3068 -6127 -3022 -6081
rect -2828 -6139 -2782 -6093
rect -2348 -6139 -2302 -6093
rect -2188 -6139 -2142 -6093
rect -1708 -6139 -1662 -6093
rect -1468 -6131 -1422 -6085
rect -154 -4303 -90 -4248
rect -156 -5194 -110 -5148
rect 901 -5198 947 -5152
rect -3049 -7099 -3003 -7053
rect -1449 -7099 -1403 -7053
rect -3049 -7899 -3003 -7853
rect -2251 -7864 -2202 -7815
rect -1449 -7899 -1403 -7853
rect -3049 -8697 -3003 -8651
rect -2251 -8665 -2202 -8616
rect -1449 -8697 -1403 -8651
rect -3049 -9497 -3003 -9451
rect -2252 -9465 -2203 -9416
rect -1449 -9497 -1403 -9451
rect -245 -6909 -199 -6863
rect 878 -6931 924 -6885
rect 2893 -6979 2945 -6927
rect 5026 -6960 5082 -6912
rect 3012 -7061 3086 -7002
rect 3582 -7067 3656 -7008
rect 4224 -7061 4298 -7002
rect 3310 -7470 3363 -7410
rect 3754 -7471 3806 -7412
rect -243 -7771 -197 -7725
rect 313 -7740 371 -7682
rect 877 -7789 923 -7743
rect 908 -8651 966 -8593
rect -243 -9514 -197 -9468
rect 304 -9569 362 -9511
rect 880 -9520 926 -9474
rect -246 -10367 -200 -10321
rect 957 -10375 1003 -10329
<< metal1 >>
rect 435 1736 564 2004
rect 406 1708 587 1736
rect 406 1601 432 1708
rect 561 1601 587 1708
rect 406 1576 587 1601
rect -3320 1441 -1246 1467
rect 1556 1465 1694 1480
rect 1556 1464 1571 1465
rect -3320 1394 -3294 1441
rect -3247 1395 -3199 1441
rect -3153 1395 -3105 1441
rect -3059 1395 -3011 1441
rect -2965 1395 -2917 1441
rect -2871 1395 -2823 1441
rect -2777 1395 -2729 1441
rect -2683 1395 -2635 1441
rect -2589 1395 -2541 1441
rect -2495 1395 -2447 1441
rect -2401 1395 -2353 1441
rect -2307 1395 -2259 1441
rect -2213 1395 -2165 1441
rect -2119 1395 -2071 1441
rect -2025 1395 -1977 1441
rect -1931 1395 -1883 1441
rect -1837 1395 -1789 1441
rect -1743 1395 -1695 1441
rect -1649 1395 -1601 1441
rect -1555 1395 -1507 1441
rect -1461 1395 -1413 1441
rect -1367 1395 -1319 1441
rect -3247 1394 -1319 1395
rect -1272 1394 -1246 1441
rect -3320 1369 -1246 1394
rect -3320 1346 -3222 1369
rect -3320 1300 -3294 1346
rect -3248 1300 -3222 1346
rect -3320 1252 -3222 1300
rect -3320 1206 -3294 1252
rect -3248 1206 -3222 1252
rect -3320 1158 -3222 1206
rect -3320 1112 -3294 1158
rect -3248 1112 -3222 1158
rect -3320 1064 -3222 1112
rect -3320 1018 -3294 1064
rect -3248 1018 -3222 1064
rect -3320 970 -3222 1018
rect -3320 924 -3294 970
rect -3248 924 -3222 970
rect -3320 876 -3222 924
rect -3320 830 -3294 876
rect -3248 830 -3222 876
rect -3320 782 -3222 830
rect -3320 736 -3294 782
rect -3248 736 -3222 782
rect -3320 688 -3222 736
rect -3320 642 -3294 688
rect -3248 642 -3222 688
rect -3320 594 -3222 642
rect -3320 548 -3294 594
rect -3248 548 -3222 594
rect -3320 500 -3222 548
rect -3320 454 -3294 500
rect -3248 454 -3222 500
rect -3320 406 -3222 454
rect -3320 360 -3294 406
rect -3248 360 -3222 406
rect -3320 312 -3222 360
rect -3320 266 -3294 312
rect -3248 266 -3222 312
rect -3320 218 -3222 266
rect -3320 172 -3294 218
rect -3248 172 -3222 218
rect -3320 124 -3222 172
rect -3320 78 -3294 124
rect -3248 78 -3222 124
rect -3320 30 -3222 78
rect -3320 -16 -3294 30
rect -3248 -16 -3222 30
rect -3320 -64 -3222 -16
rect -3320 -110 -3294 -64
rect -3248 -110 -3222 -64
rect -3320 -158 -3222 -110
rect -3320 -204 -3294 -158
rect -3248 -204 -3222 -158
rect -3320 -252 -3222 -204
rect -3320 -298 -3294 -252
rect -3248 -298 -3222 -252
rect -3320 -346 -3222 -298
rect -3320 -392 -3294 -346
rect -3248 -392 -3222 -346
rect -3320 -440 -3222 -392
rect -3320 -486 -3294 -440
rect -3248 -486 -3222 -440
rect -3320 -534 -3222 -486
rect -3320 -580 -3294 -534
rect -3248 -580 -3222 -534
rect -3320 -628 -3222 -580
rect -3320 -674 -3294 -628
rect -3248 -674 -3222 -628
rect -3320 -722 -3222 -674
rect -3320 -768 -3294 -722
rect -3248 -768 -3222 -722
rect -3320 -816 -3222 -768
rect -3320 -862 -3294 -816
rect -3248 -862 -3222 -816
rect -3320 -910 -3222 -862
rect -3320 -956 -3294 -910
rect -3248 -956 -3222 -910
rect -3320 -1004 -3222 -956
rect -3320 -1050 -3294 -1004
rect -3248 -1050 -3222 -1004
rect -3320 -1098 -3222 -1050
rect -3320 -1144 -3294 -1098
rect -3248 -1144 -3222 -1098
rect -3320 -1192 -3222 -1144
rect -3320 -1238 -3294 -1192
rect -3248 -1238 -3222 -1192
rect -3320 -1286 -3222 -1238
rect -3320 -1332 -3294 -1286
rect -3248 -1332 -3222 -1286
rect -3320 -1380 -3222 -1332
rect -3320 -1426 -3294 -1380
rect -3248 -1426 -3222 -1380
rect -3320 -1474 -3222 -1426
rect -3320 -1520 -3294 -1474
rect -3248 -1520 -3222 -1474
rect -3320 -1568 -3222 -1520
rect -3320 -1614 -3294 -1568
rect -3248 -1614 -3222 -1568
rect -3320 -1662 -3222 -1614
rect -2973 508 -2921 1149
rect -2757 508 -2705 1150
rect -2973 504 -2705 508
rect -2973 458 -2864 504
rect -2818 458 -2705 504
rect -2973 454 -2705 458
rect -2973 -228 -2921 454
rect -2757 -228 -2705 454
rect -2973 -232 -2705 -228
rect -2973 -278 -2864 -232
rect -2818 -278 -2705 -232
rect -2973 -282 -2705 -278
rect -2973 -964 -2921 -282
rect -2757 -964 -2705 -282
rect -2973 -968 -2705 -964
rect -2973 -1014 -2863 -968
rect -2817 -1014 -2705 -968
rect -2973 -1018 -2705 -1014
rect -2973 -1660 -2921 -1018
rect -3320 -1708 -3294 -1662
rect -3248 -1708 -3222 -1662
rect -3320 -1756 -3222 -1708
rect -3320 -1802 -3294 -1756
rect -3248 -1802 -3222 -1756
rect -2757 -1764 -2705 -1018
rect -3320 -1850 -3222 -1802
rect -2773 -1774 -2689 -1764
rect -2773 -1828 -2758 -1774
rect -2704 -1828 -2689 -1774
rect -2773 -1842 -2689 -1828
rect -3320 -1896 -3294 -1850
rect -3248 -1896 -3222 -1850
rect -3320 -1918 -3222 -1896
rect -2541 -1918 -2489 1369
rect -2431 1289 -2312 1320
rect -2431 1229 -2402 1289
rect -2342 1281 -2312 1289
rect -2342 1260 -2165 1281
rect -2342 1229 -2323 1260
rect -2431 1214 -2323 1229
rect -2277 1214 -2165 1260
rect -2431 1201 -2165 1214
rect -2431 507 -2379 1201
rect -2431 461 -2428 507
rect -2382 461 -2379 507
rect -2431 -232 -2379 461
rect -2431 -278 -2428 -232
rect -2382 -278 -2379 -232
rect -2431 -971 -2379 -278
rect -2431 -1017 -2428 -971
rect -2382 -1017 -2379 -971
rect -2431 -1032 -2379 -1017
rect -2325 -1764 -2273 1150
rect -2217 504 -2165 1201
rect -2217 457 -2215 504
rect -2167 457 -2165 504
rect -2217 -232 -2165 457
rect -2217 -279 -2215 -232
rect -2167 -279 -2165 -232
rect -2217 -970 -2165 -279
rect -2217 -1017 -2215 -970
rect -2167 -1017 -2165 -970
rect -2217 -1032 -2165 -1017
rect -2343 -1774 -2259 -1764
rect -2343 -1828 -2326 -1774
rect -2272 -1828 -2259 -1774
rect -2343 -1842 -2259 -1828
rect -2109 -1918 -2057 1369
rect -1344 1346 -1246 1369
rect -524 1441 1571 1464
rect -524 1383 196 1441
rect 258 1383 1571 1441
rect -524 1362 1571 1383
rect -1344 1300 -1318 1346
rect -1272 1300 -1246 1346
rect 1556 1360 1571 1362
rect 1681 1360 1694 1465
rect 1556 1345 1694 1360
rect -1344 1252 -1246 1300
rect 1353 1257 1487 1272
rect -1344 1206 -1318 1252
rect -1272 1206 -1246 1252
rect -1344 1158 -1246 1206
rect -1893 507 -1841 1150
rect -1677 507 -1625 1150
rect -1893 504 -1625 507
rect -1893 458 -1782 504
rect -1736 458 -1625 504
rect -1893 453 -1625 458
rect -1893 -228 -1841 453
rect -1677 -228 -1625 453
rect -1893 -232 -1625 -228
rect -1893 -278 -1781 -232
rect -1735 -278 -1625 -232
rect -1893 -282 -1625 -278
rect -1893 -964 -1841 -282
rect -1677 -964 -1625 -282
rect -1893 -968 -1625 -964
rect -1893 -1014 -1781 -968
rect -1735 -1014 -1625 -968
rect -1893 -1018 -1625 -1014
rect -1893 -1766 -1841 -1018
rect -1677 -1659 -1625 -1018
rect -1344 1112 -1318 1158
rect -1272 1112 -1246 1158
rect -523 1231 1365 1257
rect -523 1175 -229 1231
rect -171 1229 1365 1231
rect -171 1175 631 1229
rect -523 1172 631 1175
rect 691 1172 1365 1229
rect -523 1153 1365 1172
rect 1474 1153 1487 1257
rect 1353 1137 1487 1153
rect -1344 1064 -1246 1112
rect -1344 1018 -1318 1064
rect -1272 1018 -1246 1064
rect -1344 970 -1246 1018
rect -1344 924 -1318 970
rect -1272 924 -1246 970
rect -1344 876 -1246 924
rect -1344 830 -1318 876
rect -1272 845 -1246 876
rect -773 1013 1244 1039
rect -773 967 -747 1013
rect -701 967 -653 1013
rect -607 967 -552 1013
rect -506 967 -458 1013
rect -412 967 -362 1013
rect -316 967 -268 1013
rect -222 967 -167 1013
rect -121 967 -73 1013
rect -27 967 21 1013
rect 67 967 115 1013
rect 161 967 216 1013
rect 262 967 310 1013
rect 356 967 406 1013
rect 452 967 500 1013
rect 546 967 601 1013
rect 647 967 695 1013
rect 741 967 789 1013
rect 835 967 883 1013
rect 929 967 984 1013
rect 1030 967 1078 1013
rect 1124 967 1172 1013
rect 1218 967 1244 1013
rect -773 941 1244 967
rect -773 917 -675 941
rect -773 871 -747 917
rect -701 871 -675 917
rect -773 845 -675 871
rect -1272 830 -675 845
rect -1344 823 -675 830
rect -1344 782 -747 823
rect -1344 736 -1318 782
rect -1272 777 -747 782
rect -701 777 -675 823
rect -1272 736 -675 777
rect -1344 727 -675 736
rect -1344 708 -747 727
rect -1344 688 -1246 708
rect -1344 642 -1318 688
rect -1272 642 -1246 688
rect -1344 594 -1246 642
rect -1344 548 -1318 594
rect -1272 548 -1246 594
rect -1344 500 -1246 548
rect -1344 454 -1318 500
rect -1272 454 -1246 500
rect -1344 406 -1246 454
rect -1344 360 -1318 406
rect -1272 360 -1246 406
rect -1344 312 -1246 360
rect -1344 266 -1318 312
rect -1272 266 -1246 312
rect -1344 218 -1246 266
rect -1344 172 -1318 218
rect -1272 172 -1246 218
rect -1344 124 -1246 172
rect -1344 78 -1318 124
rect -1272 78 -1246 124
rect -1344 58 -1246 78
rect -773 681 -747 708
rect -701 681 -675 727
rect -440 848 -160 860
rect -440 842 -230 848
rect -440 796 -336 842
rect -290 796 -230 842
rect -440 792 -230 796
rect -172 792 -160 848
rect -440 780 -160 792
rect -440 712 -394 780
rect -224 712 -178 780
rect -8 689 38 941
rect 183 847 273 860
rect 183 789 199 847
rect 259 789 273 847
rect 183 775 273 789
rect 208 712 254 775
rect 424 712 470 941
rect 1146 917 1244 941
rect 1146 871 1172 917
rect 1218 871 1244 917
rect 619 851 902 864
rect 619 794 632 851
rect 692 844 902 851
rect 692 798 750 844
rect 796 798 902 844
rect 692 794 902 798
rect 619 782 902 794
rect 640 712 686 782
rect 856 712 902 782
rect 1146 816 1244 871
rect 1146 770 1172 816
rect 1218 770 1244 816
rect 1146 722 1244 770
rect -773 633 -675 681
rect -773 587 -747 633
rect -701 587 -675 633
rect -773 539 -675 587
rect -773 493 -747 539
rect -701 493 -675 539
rect -773 438 -675 493
rect -773 392 -747 438
rect -701 392 -675 438
rect -773 344 -675 392
rect -773 298 -747 344
rect -701 298 -675 344
rect -773 248 -675 298
rect -773 202 -747 248
rect -701 202 -675 248
rect -773 154 -675 202
rect -773 108 -747 154
rect -701 108 -675 154
rect 1146 676 1172 722
rect 1218 676 1244 722
rect 1146 628 1244 676
rect 1146 582 1172 628
rect 1218 582 1244 628
rect 1146 534 1244 582
rect 1146 488 1172 534
rect 1218 488 1244 534
rect 1146 433 1244 488
rect 1146 387 1172 433
rect 1218 387 1244 433
rect 1146 339 1244 387
rect 1146 293 1172 339
rect 1218 293 1244 339
rect 1146 243 1244 293
rect 1146 197 1172 243
rect 1218 197 1244 243
rect 1146 149 1244 197
rect -773 58 -675 108
rect -1344 53 -675 58
rect -1344 30 -747 53
rect -1344 -16 -1318 30
rect -1272 7 -747 30
rect -701 7 -675 53
rect -1272 -16 -675 7
rect -1344 -41 -675 -16
rect -1344 -64 -747 -41
rect -1344 -110 -1318 -64
rect -1272 -79 -747 -64
rect -1272 -110 -1246 -79
rect -1344 -158 -1246 -110
rect -1344 -204 -1318 -158
rect -1272 -204 -1246 -158
rect -1344 -252 -1246 -204
rect -1344 -298 -1318 -252
rect -1272 -298 -1246 -252
rect -1344 -346 -1246 -298
rect -1344 -392 -1318 -346
rect -1272 -392 -1246 -346
rect -1344 -440 -1246 -392
rect -1344 -486 -1318 -440
rect -1272 -486 -1246 -440
rect -1344 -534 -1246 -486
rect -1344 -580 -1318 -534
rect -1272 -580 -1246 -534
rect -1344 -614 -1246 -580
rect -773 -87 -747 -79
rect -701 -87 -675 -41
rect -773 -135 -675 -87
rect -773 -181 -747 -135
rect -701 -181 -675 -135
rect -260 -66 -144 -44
rect -260 -145 -242 -66
rect -160 -145 -144 -66
rect -260 -160 -144 -145
rect -773 -229 -675 -181
rect -773 -275 -747 -229
rect -701 -275 -675 -229
rect -773 -330 -675 -275
rect -224 -326 -178 -160
rect -8 -326 38 116
rect 96 -60 148 -36
rect 96 -106 99 -60
rect 145 -106 148 -60
rect -773 -376 -747 -330
rect -701 -376 -675 -330
rect -773 -424 -675 -376
rect -773 -470 -747 -424
rect -701 -470 -675 -424
rect -773 -520 -675 -470
rect -773 -566 -747 -520
rect -701 -566 -675 -520
rect -773 -614 -675 -566
rect -1344 -628 -747 -614
rect -1344 -674 -1318 -628
rect -1272 -660 -747 -628
rect -701 -660 -675 -614
rect -1272 -674 -675 -660
rect -1344 -715 -675 -674
rect -1344 -722 -747 -715
rect -1344 -768 -1318 -722
rect -1272 -751 -747 -722
rect -1272 -768 -1246 -751
rect -1344 -816 -1246 -768
rect -1344 -862 -1318 -816
rect -1272 -862 -1246 -816
rect -1344 -910 -1246 -862
rect -1344 -956 -1318 -910
rect -1272 -956 -1246 -910
rect -1344 -1004 -1246 -956
rect -1344 -1050 -1318 -1004
rect -1272 -1050 -1246 -1004
rect -1344 -1098 -1246 -1050
rect -1344 -1144 -1318 -1098
rect -1272 -1144 -1246 -1098
rect -1344 -1192 -1246 -1144
rect -1344 -1238 -1318 -1192
rect -1272 -1238 -1246 -1192
rect -773 -761 -747 -751
rect -701 -761 -675 -715
rect -773 -809 -675 -761
rect -773 -855 -747 -809
rect -701 -855 -675 -809
rect -773 -903 -675 -855
rect -773 -949 -747 -903
rect -701 -949 -675 -903
rect -773 -997 -675 -949
rect -773 -1043 -747 -997
rect -701 -1043 -675 -997
rect -773 -1098 -675 -1043
rect -773 -1144 -747 -1098
rect -701 -1144 -675 -1098
rect -773 -1192 -675 -1144
rect -773 -1238 -747 -1192
rect -701 -1238 -675 -1192
rect -1344 -1286 -675 -1238
rect -1344 -1332 -1318 -1286
rect -1272 -1288 -675 -1286
rect -1272 -1332 -747 -1288
rect -1344 -1334 -747 -1332
rect -701 -1334 -675 -1288
rect -1344 -1375 -675 -1334
rect -440 -1121 -394 -922
rect -224 -1121 -178 -922
rect -440 -1122 -178 -1121
rect -440 -1170 -330 -1122
rect -283 -1170 -178 -1122
rect -440 -1172 -178 -1170
rect -440 -1366 -394 -1172
rect -224 -1366 -178 -1172
rect -8 -1366 38 -922
rect 96 -1135 148 -106
rect 424 -326 470 116
rect 1146 103 1172 149
rect 1218 103 1244 149
rect 1146 48 1244 103
rect 1146 2 1172 48
rect 1218 2 1244 48
rect 1146 -46 1244 2
rect 605 -71 721 -51
rect 605 -150 621 -71
rect 703 -150 721 -71
rect 605 -167 721 -150
rect 1146 -92 1172 -46
rect 1218 -92 1244 -46
rect 1146 -140 1244 -92
rect 640 -326 686 -167
rect 1146 -186 1172 -140
rect 1218 -186 1244 -140
rect 1146 -234 1244 -186
rect 1146 -280 1172 -234
rect 1218 -280 1244 -234
rect 1146 -335 1244 -280
rect 1146 -381 1172 -335
rect 1218 -381 1244 -335
rect 1146 -429 1244 -381
rect 1146 -475 1172 -429
rect 1218 -475 1244 -429
rect 1146 -525 1244 -475
rect 1146 -571 1172 -525
rect 1218 -571 1244 -525
rect 1146 -619 1244 -571
rect 1146 -665 1172 -619
rect 1218 -665 1244 -619
rect 1146 -720 1244 -665
rect 1146 -766 1172 -720
rect 1218 -766 1244 -720
rect 1146 -814 1244 -766
rect 1146 -860 1172 -814
rect 1218 -860 1244 -814
rect 1146 -908 1244 -860
rect 96 -1181 99 -1135
rect 145 -1181 148 -1135
rect -1344 -1380 -1246 -1375
rect -1344 -1426 -1318 -1380
rect -1272 -1426 -1246 -1380
rect -1344 -1474 -1246 -1426
rect -1344 -1520 -1318 -1474
rect -1272 -1520 -1246 -1474
rect -1344 -1568 -1246 -1520
rect -1344 -1614 -1318 -1568
rect -1272 -1614 -1246 -1568
rect -1344 -1662 -1246 -1614
rect -1344 -1708 -1318 -1662
rect -1272 -1708 -1246 -1662
rect -1344 -1756 -1246 -1708
rect -1909 -1777 -1825 -1766
rect -1909 -1831 -1894 -1777
rect -1840 -1831 -1825 -1777
rect -1909 -1844 -1825 -1831
rect -1344 -1802 -1318 -1756
rect -1272 -1802 -1246 -1756
rect -1344 -1813 -1246 -1802
rect -773 -1382 -675 -1375
rect -773 -1428 -747 -1382
rect -701 -1428 -675 -1382
rect -773 -1476 -675 -1428
rect -773 -1522 -747 -1476
rect -701 -1522 -675 -1476
rect -773 -1577 -675 -1522
rect -773 -1623 -747 -1577
rect -701 -1623 -675 -1577
rect -773 -1671 -675 -1623
rect -773 -1717 -747 -1671
rect -701 -1717 -675 -1671
rect -773 -1767 -675 -1717
rect -773 -1813 -747 -1767
rect -701 -1813 -675 -1767
rect -1344 -1850 -675 -1813
rect -1344 -1896 -1318 -1850
rect -1272 -1861 -675 -1850
rect -1272 -1896 -747 -1861
rect -1344 -1907 -747 -1896
rect -701 -1907 -675 -1861
rect -1344 -1918 -675 -1907
rect -3320 -1944 -675 -1918
rect -3320 -1990 -3293 -1944
rect -3247 -1990 -3199 -1944
rect -3153 -1990 -3105 -1944
rect -3059 -1990 -3011 -1944
rect -2965 -1990 -2917 -1944
rect -2871 -1990 -2823 -1944
rect -2777 -1990 -2729 -1944
rect -2683 -1990 -2635 -1944
rect -2589 -1990 -2541 -1944
rect -2495 -1990 -2447 -1944
rect -2401 -1990 -2353 -1944
rect -2307 -1990 -2259 -1944
rect -2213 -1990 -2165 -1944
rect -2119 -1990 -2071 -1944
rect -2025 -1990 -1977 -1944
rect -1931 -1990 -1883 -1944
rect -1837 -1990 -1789 -1944
rect -1743 -1990 -1695 -1944
rect -1649 -1990 -1601 -1944
rect -1555 -1990 -1507 -1944
rect -1461 -1990 -1413 -1944
rect -1367 -1990 -1319 -1944
rect -1273 -1950 -675 -1944
rect -1273 -1990 -1246 -1950
rect -3320 -2016 -1246 -1990
rect -773 -1962 -675 -1950
rect -773 -2008 -747 -1962
rect -701 -2008 -675 -1962
rect -3472 -2206 -1779 -2187
rect -3472 -2262 -3452 -2206
rect -3396 -2262 -3341 -2206
rect -3285 -2208 -1779 -2206
rect -3285 -2212 -2327 -2208
rect -3285 -2262 -2759 -2212
rect -3472 -2268 -2759 -2262
rect -2703 -2264 -2327 -2212
rect -2271 -2216 -1779 -2208
rect -2271 -2264 -1895 -2216
rect -2703 -2268 -1895 -2264
rect -3472 -2272 -1895 -2268
rect -1839 -2272 -1779 -2216
rect -3472 -2309 -1779 -2272
rect -3472 -2316 -3250 -2309
rect -3472 -2372 -3453 -2316
rect -3397 -2372 -3342 -2316
rect -3286 -2372 -3250 -2316
rect -3472 -2404 -3250 -2372
rect -3668 -2505 -3546 -2473
rect -3668 -2569 -3639 -2505
rect -3575 -2569 -3546 -2505
rect -1536 -2567 -1372 -2016
rect -773 -2056 -675 -2008
rect -773 -2102 -747 -2056
rect -701 -2102 -675 -2056
rect -773 -2150 -675 -2102
rect -773 -2196 -747 -2150
rect -701 -2196 -675 -2150
rect -773 -2244 -675 -2196
rect -328 -2169 -135 -2154
rect -328 -2170 -205 -2169
rect -328 -2223 -313 -2170
rect -260 -2221 -205 -2170
rect -153 -2221 -135 -2169
rect -260 -2223 -135 -2221
rect -328 -2236 -135 -2223
rect -773 -2290 -747 -2244
rect -701 -2290 -675 -2244
rect -773 -2345 -675 -2290
rect -773 -2391 -747 -2345
rect -701 -2391 -675 -2345
rect -773 -2439 -675 -2391
rect -8 -2404 38 -1962
rect 96 -2154 148 -1181
rect 208 -1103 254 -922
rect 208 -1117 353 -1103
rect 208 -1181 283 -1117
rect 341 -1181 353 -1117
rect 208 -1194 353 -1181
rect 208 -1366 254 -1194
rect 424 -1366 470 -922
rect 640 -1121 686 -922
rect 856 -1121 902 -922
rect 640 -1123 902 -1121
rect 640 -1169 752 -1123
rect 798 -1169 902 -1123
rect 640 -1172 902 -1169
rect 640 -1366 686 -1172
rect 856 -1366 902 -1172
rect 1146 -954 1172 -908
rect 1218 -954 1244 -908
rect 1146 -1004 1244 -954
rect 1146 -1050 1172 -1004
rect 1218 -1050 1244 -1004
rect 1146 -1098 1244 -1050
rect 1146 -1144 1172 -1098
rect 1218 -1144 1244 -1098
rect 1146 -1199 1244 -1144
rect 1146 -1245 1172 -1199
rect 1218 -1245 1244 -1199
rect 1146 -1293 1244 -1245
rect 1146 -1339 1172 -1293
rect 1218 -1339 1244 -1293
rect 1146 -1387 1244 -1339
rect 1146 -1433 1172 -1387
rect 1218 -1433 1244 -1387
rect 1146 -1481 1244 -1433
rect 1146 -1527 1172 -1481
rect 1218 -1527 1244 -1481
rect 1146 -1582 1244 -1527
rect 1146 -1628 1172 -1582
rect 1218 -1628 1244 -1582
rect 1146 -1676 1244 -1628
rect 1146 -1722 1172 -1676
rect 1218 -1722 1244 -1676
rect 1146 -1772 1244 -1722
rect 1146 -1818 1172 -1772
rect 1218 -1818 1244 -1772
rect 1146 -1866 1244 -1818
rect 1146 -1912 1172 -1866
rect 1218 -1912 1244 -1866
rect 96 -2167 259 -2154
rect 96 -2171 195 -2167
rect 96 -2217 130 -2171
rect 176 -2217 195 -2171
rect 96 -2219 195 -2217
rect 247 -2219 259 -2167
rect 96 -2237 259 -2219
rect 424 -2404 470 -1962
rect 1146 -1967 1244 -1912
rect 1146 -2013 1172 -1967
rect 1218 -2013 1244 -1967
rect 1146 -2061 1244 -2013
rect 1146 -2107 1172 -2061
rect 1218 -2107 1244 -2061
rect 1146 -2155 1244 -2107
rect 1146 -2201 1172 -2155
rect 1218 -2201 1244 -2155
rect 1146 -2249 1244 -2201
rect 1146 -2295 1172 -2249
rect 1218 -2295 1244 -2249
rect 1146 -2350 1244 -2295
rect 1146 -2396 1172 -2350
rect 1218 -2396 1244 -2350
rect -773 -2485 -747 -2439
rect -701 -2485 -675 -2439
rect -773 -2535 -675 -2485
rect -3668 -2597 -3546 -2569
rect -3293 -2593 -1219 -2567
rect -3293 -2640 -3267 -2593
rect -3220 -2639 -3172 -2593
rect -3126 -2639 -3078 -2593
rect -3032 -2639 -2984 -2593
rect -2938 -2639 -2890 -2593
rect -2844 -2639 -2796 -2593
rect -2750 -2639 -2702 -2593
rect -2656 -2639 -2608 -2593
rect -2562 -2639 -2514 -2593
rect -2468 -2639 -2420 -2593
rect -2374 -2639 -2326 -2593
rect -2280 -2639 -2232 -2593
rect -2186 -2639 -2138 -2593
rect -2092 -2639 -2044 -2593
rect -1998 -2639 -1950 -2593
rect -1904 -2639 -1856 -2593
rect -1810 -2639 -1762 -2593
rect -1716 -2639 -1668 -2593
rect -1622 -2639 -1574 -2593
rect -1528 -2639 -1480 -2593
rect -1434 -2639 -1386 -2593
rect -1340 -2639 -1292 -2593
rect -3220 -2640 -1292 -2639
rect -1245 -2640 -1219 -2593
rect -3293 -2654 -1219 -2640
rect -773 -2581 -747 -2535
rect -701 -2581 -675 -2535
rect -773 -2629 -675 -2581
rect -773 -2654 -747 -2629
rect -3293 -2665 -747 -2654
rect -3293 -2688 -3195 -2665
rect -3664 -2739 -3542 -2707
rect -3664 -2803 -3635 -2739
rect -3571 -2803 -3542 -2739
rect -3664 -2831 -3542 -2803
rect -3293 -2734 -3267 -2688
rect -3221 -2734 -3195 -2688
rect -1317 -2675 -747 -2665
rect -701 -2675 -675 -2629
rect -1317 -2688 -675 -2675
rect -3293 -2782 -3195 -2734
rect -1743 -2743 -1642 -2723
rect -3293 -2828 -3267 -2782
rect -3221 -2828 -3195 -2782
rect -2849 -2744 -1642 -2743
rect -2849 -2747 -1722 -2744
rect -1666 -2747 -1642 -2744
rect -2849 -2793 -2828 -2747
rect -2782 -2793 -2348 -2747
rect -2302 -2793 -2188 -2747
rect -2142 -2793 -1722 -2747
rect -1662 -2793 -1642 -2747
rect -2849 -2799 -1722 -2793
rect -1743 -2800 -1722 -2799
rect -1666 -2800 -1642 -2793
rect -1743 -2820 -1642 -2800
rect -1317 -2734 -1291 -2688
rect -1245 -2730 -675 -2688
rect -1245 -2734 -747 -2730
rect -1317 -2776 -747 -2734
rect -701 -2776 -675 -2730
rect -1317 -2782 -675 -2776
rect -3293 -2876 -3195 -2828
rect -3293 -2922 -3267 -2876
rect -3221 -2922 -3195 -2876
rect -3293 -2970 -3195 -2922
rect -1317 -2828 -1291 -2782
rect -1245 -2793 -675 -2782
rect -1245 -2828 -1219 -2793
rect -1317 -2876 -1219 -2828
rect -1317 -2922 -1291 -2876
rect -1245 -2922 -1219 -2876
rect -3293 -3016 -3267 -2970
rect -3221 -3016 -3195 -2970
rect -3293 -3064 -3195 -3016
rect -2607 -2967 -2524 -2953
rect -2607 -3023 -2593 -2967
rect -2537 -3023 -2524 -2967
rect -2607 -3035 -2524 -3023
rect -1965 -2967 -1882 -2952
rect -1965 -3023 -1952 -2967
rect -1896 -3023 -1882 -2967
rect -1965 -3036 -1882 -3023
rect -1317 -2970 -1219 -2922
rect -1317 -3016 -1291 -2970
rect -1245 -3016 -1219 -2970
rect -3293 -3110 -3267 -3064
rect -3221 -3110 -3195 -3064
rect -1317 -3064 -1219 -3016
rect -3293 -3158 -3195 -3110
rect -3293 -3204 -3267 -3158
rect -3221 -3204 -3195 -3158
rect -2766 -3119 -2683 -3105
rect -2766 -3175 -2752 -3119
rect -2696 -3175 -2683 -3119
rect -2766 -3187 -2683 -3175
rect -2447 -3118 -2364 -3104
rect -2447 -3174 -2433 -3118
rect -2377 -3174 -2364 -3118
rect -2447 -3186 -2364 -3174
rect -2125 -3118 -2042 -3104
rect -2125 -3174 -2111 -3118
rect -2055 -3174 -2042 -3118
rect -2125 -3186 -2042 -3174
rect -1810 -3118 -1727 -3104
rect -1810 -3174 -1796 -3118
rect -1740 -3174 -1727 -3118
rect -1810 -3186 -1727 -3174
rect -1317 -3110 -1291 -3064
rect -1245 -3110 -1219 -3064
rect -1317 -3158 -1219 -3110
rect -3293 -3252 -3195 -3204
rect -3293 -3298 -3267 -3252
rect -3221 -3298 -3195 -3252
rect -1317 -3204 -1291 -3158
rect -1245 -3189 -1219 -3158
rect -773 -2824 -675 -2793
rect -773 -2870 -747 -2824
rect -701 -2870 -675 -2824
rect -773 -2918 -675 -2870
rect -773 -2964 -747 -2918
rect -701 -2964 -675 -2918
rect -773 -3012 -675 -2964
rect 1146 -2444 1244 -2396
rect 1146 -2490 1172 -2444
rect 1218 -2490 1244 -2444
rect 1146 -2540 1244 -2490
rect 1146 -2586 1172 -2540
rect 1218 -2586 1244 -2540
rect 1146 -2634 1244 -2586
rect 1146 -2680 1172 -2634
rect 1218 -2680 1244 -2634
rect 1146 -2735 1244 -2680
rect 1146 -2781 1172 -2735
rect 1218 -2781 1244 -2735
rect 1146 -2829 1244 -2781
rect 1146 -2875 1172 -2829
rect 1218 -2875 1244 -2829
rect 1146 -2923 1244 -2875
rect 1146 -2969 1172 -2923
rect 1218 -2969 1244 -2923
rect -773 -3058 -747 -3012
rect -701 -3058 -675 -3012
rect -773 -3113 -675 -3058
rect -773 -3159 -747 -3113
rect -701 -3159 -675 -3113
rect -773 -3189 -675 -3159
rect -1245 -3204 -675 -3189
rect -440 -3114 -394 -3000
rect -224 -3114 -178 -3000
rect -440 -3126 -160 -3114
rect -440 -3132 -233 -3126
rect -440 -3184 -333 -3132
rect -276 -3184 -233 -3132
rect -440 -3185 -233 -3184
rect -172 -3185 -160 -3126
rect -440 -3198 -160 -3185
rect -1317 -3207 -675 -3204
rect -1317 -3252 -747 -3207
rect -3293 -3346 -3195 -3298
rect -3088 -3274 -3004 -3260
rect -3088 -3330 -3074 -3274
rect -3018 -3330 -3004 -3274
rect -3088 -3344 -3004 -3330
rect -2927 -3274 -2843 -3259
rect -2927 -3330 -2913 -3274
rect -2857 -3330 -2843 -3274
rect -2927 -3343 -2843 -3330
rect -2288 -3274 -2202 -3260
rect -2288 -3330 -2274 -3274
rect -2216 -3330 -2202 -3274
rect -2288 -3344 -2202 -3330
rect -1647 -3274 -1563 -3259
rect -1647 -3330 -1633 -3274
rect -1577 -3330 -1563 -3274
rect -1647 -3343 -1563 -3330
rect -1487 -3274 -1403 -3260
rect -1487 -3330 -1473 -3274
rect -1417 -3330 -1403 -3274
rect -1487 -3344 -1403 -3330
rect -1317 -3298 -1291 -3252
rect -1245 -3253 -747 -3252
rect -701 -3253 -675 -3207
rect -1245 -3277 -675 -3253
rect -8 -3277 38 -2999
rect 208 -3116 254 -3000
rect 208 -3117 255 -3116
rect 188 -3129 273 -3117
rect 188 -3188 200 -3129
rect 261 -3188 273 -3129
rect 188 -3201 273 -3188
rect 424 -3277 470 -2999
rect 640 -3112 686 -3000
rect 856 -3112 902 -3000
rect 620 -3126 902 -3112
rect 620 -3185 632 -3126
rect 693 -3128 902 -3126
rect 693 -3182 738 -3128
rect 796 -3182 902 -3128
rect 693 -3185 902 -3182
rect 620 -3198 902 -3185
rect 1146 -3019 1244 -2969
rect 1146 -3065 1172 -3019
rect 1218 -3065 1244 -3019
rect 1146 -3113 1244 -3065
rect 1146 -3159 1172 -3113
rect 1218 -3159 1244 -3113
rect 1146 -3207 1244 -3159
rect 1146 -3253 1172 -3207
rect 1218 -3253 1244 -3207
rect 1146 -3277 1244 -3253
rect -1245 -3298 1244 -3277
rect -1317 -3303 1244 -3298
rect -1317 -3328 -747 -3303
rect -3293 -3392 -3267 -3346
rect -3221 -3392 -3195 -3346
rect -3293 -3440 -3195 -3392
rect -3293 -3486 -3267 -3440
rect -3221 -3486 -3195 -3440
rect -1317 -3346 -1219 -3328
rect -1317 -3392 -1291 -3346
rect -1245 -3392 -1219 -3346
rect -1317 -3440 -1219 -3392
rect -3293 -3534 -3195 -3486
rect -3068 -3509 -3022 -3461
rect -3293 -3580 -3267 -3534
rect -3221 -3580 -3195 -3534
rect -3293 -3628 -3195 -3580
rect -3077 -3534 -3003 -3509
rect -1468 -3515 -1422 -3463
rect -1317 -3486 -1291 -3440
rect -1245 -3486 -1219 -3440
rect -3077 -3580 -3061 -3534
rect -3015 -3580 -3003 -3534
rect -1480 -3525 -1410 -3515
rect -3077 -3595 -3003 -3580
rect -2852 -3561 -2751 -3540
rect -3293 -3674 -3267 -3628
rect -3221 -3674 -3195 -3628
rect -2852 -3617 -2831 -3561
rect -2775 -3563 -2751 -3561
rect -2684 -3559 -2606 -3542
rect -2684 -3563 -2668 -3559
rect -2852 -3626 -2829 -3617
rect -2775 -3605 -2668 -3563
rect -2622 -3563 -2606 -3559
rect -2524 -3558 -2446 -3542
rect -2524 -3563 -2508 -3558
rect -2622 -3604 -2508 -3563
rect -2462 -3563 -2446 -3558
rect -2044 -3558 -1966 -3542
rect -2044 -3563 -2028 -3558
rect -2462 -3577 -2028 -3563
rect -2462 -3604 -2348 -3577
rect -2622 -3605 -2348 -3604
rect -2775 -3617 -2348 -3605
rect -2783 -3619 -2348 -3617
rect -2783 -3626 -2751 -3619
rect -2852 -3637 -2751 -3626
rect -2363 -3623 -2348 -3619
rect -2302 -3619 -2188 -3577
rect -2302 -3623 -2285 -3619
rect -2845 -3640 -2767 -3637
rect -2363 -3640 -2285 -3623
rect -2205 -3623 -2188 -3619
rect -2142 -3604 -2028 -3577
rect -1982 -3563 -1966 -3558
rect -1884 -3559 -1806 -3542
rect -1884 -3563 -1868 -3559
rect -1982 -3604 -1868 -3563
rect -2142 -3605 -1868 -3604
rect -1822 -3563 -1806 -3559
rect -1822 -3580 -1645 -3563
rect -1822 -3605 -1707 -3580
rect -2142 -3619 -1707 -3605
rect -2142 -3623 -2127 -3619
rect -2205 -3640 -2127 -3623
rect -1723 -3626 -1707 -3619
rect -1661 -3626 -1645 -3580
rect -1480 -3571 -1468 -3525
rect -1422 -3571 -1410 -3525
rect -1480 -3583 -1410 -3571
rect -1317 -3534 -1219 -3486
rect -1317 -3580 -1291 -3534
rect -1245 -3580 -1219 -3534
rect -1723 -3640 -1645 -3626
rect -1317 -3628 -1219 -3580
rect -3293 -3722 -3195 -3674
rect -3293 -3768 -3267 -3722
rect -3221 -3768 -3195 -3722
rect -3293 -3816 -3195 -3768
rect -1317 -3674 -1291 -3628
rect -1245 -3674 -1219 -3628
rect -1317 -3722 -1219 -3674
rect -1317 -3768 -1291 -3722
rect -1245 -3768 -1219 -3722
rect -3293 -3862 -3267 -3816
rect -3221 -3862 -3195 -3816
rect -3293 -3910 -3195 -3862
rect -2607 -3822 -2524 -3808
rect -2607 -3878 -2593 -3822
rect -2537 -3878 -2524 -3822
rect -2607 -3890 -2524 -3878
rect -1965 -3822 -1882 -3809
rect -1965 -3878 -1952 -3822
rect -1896 -3878 -1882 -3822
rect -1965 -3891 -1882 -3878
rect -1317 -3816 -1219 -3768
rect -1317 -3862 -1291 -3816
rect -1245 -3862 -1219 -3816
rect -3293 -3956 -3267 -3910
rect -3221 -3956 -3195 -3910
rect -3293 -4004 -3195 -3956
rect -1317 -3910 -1219 -3862
rect -1317 -3956 -1291 -3910
rect -1245 -3956 -1219 -3910
rect -3293 -4050 -3267 -4004
rect -3221 -4050 -3195 -4004
rect -2767 -3975 -2684 -3961
rect -2767 -4031 -2753 -3975
rect -2697 -4031 -2684 -3975
rect -2767 -4043 -2684 -4031
rect -2446 -3971 -2363 -3960
rect -2446 -4033 -2435 -3971
rect -2373 -4033 -2363 -3971
rect -2446 -4042 -2363 -4033
rect -2126 -3974 -2043 -3960
rect -2126 -4030 -2112 -3974
rect -2056 -4030 -2043 -3974
rect -2126 -4042 -2043 -4030
rect -1806 -3975 -1723 -3961
rect -1806 -4031 -1792 -3975
rect -1736 -4031 -1723 -3975
rect -1806 -4043 -1723 -4031
rect -1317 -4004 -1219 -3956
rect -3293 -4098 -3195 -4050
rect -3293 -4144 -3267 -4098
rect -3221 -4144 -3195 -4098
rect -1317 -4050 -1291 -4004
rect -1245 -4050 -1219 -4004
rect -1317 -4098 -1219 -4050
rect -3293 -4192 -3195 -4144
rect -3293 -4238 -3267 -4192
rect -3221 -4238 -3195 -4192
rect -3088 -4134 -3004 -4120
rect -3088 -4190 -3074 -4134
rect -3018 -4190 -3004 -4134
rect -3088 -4204 -3004 -4190
rect -2927 -4134 -2843 -4119
rect -2927 -4190 -2913 -4134
rect -2857 -4190 -2843 -4134
rect -2927 -4203 -2843 -4190
rect -2288 -4134 -2202 -4120
rect -2288 -4190 -2274 -4134
rect -2216 -4190 -2202 -4134
rect -2288 -4204 -2202 -4190
rect -1647 -4134 -1563 -4119
rect -1647 -4190 -1633 -4134
rect -1577 -4190 -1563 -4134
rect -1647 -4203 -1563 -4190
rect -1487 -4134 -1403 -4120
rect -1487 -4190 -1473 -4134
rect -1417 -4190 -1403 -4134
rect -1487 -4204 -1403 -4190
rect -1317 -4144 -1291 -4098
rect -1245 -4121 -1219 -4098
rect -1071 -4121 -912 -3328
rect -773 -3349 -747 -3328
rect -701 -3349 -653 -3303
rect -607 -3349 -552 -3303
rect -506 -3349 -458 -3303
rect -412 -3349 -362 -3303
rect -316 -3349 -268 -3303
rect -222 -3349 -167 -3303
rect -121 -3349 -73 -3303
rect -27 -3349 21 -3303
rect 67 -3349 115 -3303
rect 161 -3349 216 -3303
rect 262 -3349 310 -3303
rect 356 -3349 406 -3303
rect 452 -3349 500 -3303
rect 546 -3349 601 -3303
rect 647 -3349 695 -3303
rect 741 -3349 789 -3303
rect 835 -3349 883 -3303
rect 929 -3349 984 -3303
rect 1030 -3349 1078 -3303
rect 1124 -3349 1172 -3303
rect 1218 -3349 1244 -3303
rect -773 -3375 1244 -3349
rect 1352 -3497 1486 -3482
rect -308 -3513 1364 -3497
rect -308 -3573 -233 -3513
rect -171 -3516 1364 -3513
rect -171 -3573 634 -3516
rect -308 -3577 634 -3573
rect 695 -3577 1364 -3516
rect -308 -3601 1364 -3577
rect 1473 -3601 1486 -3497
rect 1352 -3617 1486 -3601
rect 1550 -3693 1688 -3678
rect 1550 -3694 1565 -3693
rect -308 -3710 1565 -3694
rect -308 -3773 198 -3710
rect 260 -3773 1565 -3710
rect -308 -3796 1565 -3773
rect 1550 -3798 1565 -3796
rect 1675 -3798 1688 -3693
rect 1550 -3813 1688 -3798
rect -488 -4068 1304 -4042
rect -488 -4115 -462 -4068
rect -415 -4114 -367 -4068
rect -321 -4114 -273 -4068
rect -227 -4114 -179 -4068
rect -133 -4114 -85 -4068
rect -39 -4114 9 -4068
rect 55 -4114 103 -4068
rect 149 -4114 197 -4068
rect 243 -4114 291 -4068
rect 337 -4114 385 -4068
rect 431 -4114 479 -4068
rect 525 -4114 573 -4068
rect 619 -4114 667 -4068
rect 713 -4114 761 -4068
rect 807 -4114 855 -4068
rect 901 -4114 949 -4068
rect 995 -4114 1043 -4068
rect 1089 -4114 1137 -4068
rect 1183 -4114 1231 -4068
rect -415 -4115 1231 -4114
rect 1278 -4115 1304 -4068
rect -488 -4121 1304 -4115
rect -1245 -4140 1304 -4121
rect -1245 -4144 -390 -4140
rect -1317 -4163 -390 -4144
rect -1317 -4192 -462 -4163
rect -3293 -4286 -3195 -4238
rect -3293 -4332 -3267 -4286
rect -3221 -4332 -3195 -4286
rect -1317 -4238 -1291 -4192
rect -1245 -4213 -462 -4192
rect -416 -4213 -390 -4163
rect -1245 -4238 -390 -4213
rect 1206 -4163 1304 -4140
rect 1206 -4213 1232 -4163
rect 1278 -4213 1304 -4163
rect -1317 -4261 -390 -4238
rect -1317 -4268 -462 -4261
rect -1317 -4286 -1219 -4268
rect -3293 -4380 -3195 -4332
rect -3068 -4373 -3022 -4315
rect -1468 -4369 -1422 -4315
rect -1317 -4332 -1291 -4286
rect -1245 -4332 -1219 -4286
rect -3293 -4426 -3267 -4380
rect -3221 -4426 -3195 -4380
rect -3293 -4474 -3195 -4426
rect -3080 -4380 -3010 -4373
rect -3080 -4426 -3068 -4380
rect -3022 -4426 -3010 -4380
rect -1480 -4381 -1410 -4369
rect -1745 -4404 -1644 -4386
rect -1745 -4415 -1726 -4404
rect -3080 -4439 -3010 -4426
rect -2688 -4420 -1726 -4415
rect -2688 -4466 -2667 -4420
rect -2621 -4466 -2507 -4420
rect -2461 -4466 -2029 -4420
rect -1983 -4466 -1869 -4420
rect -1823 -4465 -1726 -4420
rect -1664 -4465 -1644 -4404
rect -1480 -4427 -1468 -4381
rect -1422 -4427 -1410 -4381
rect -1480 -4439 -1410 -4427
rect -1317 -4380 -1219 -4332
rect -1317 -4426 -1291 -4380
rect -1245 -4426 -1219 -4380
rect -1823 -4466 -1644 -4465
rect -2688 -4471 -1644 -4466
rect -3293 -4520 -3267 -4474
rect -3221 -4520 -3195 -4474
rect -1745 -4483 -1644 -4471
rect -1317 -4474 -1219 -4426
rect -3293 -4568 -3195 -4520
rect -3293 -4614 -3267 -4568
rect -3221 -4614 -3195 -4568
rect -1317 -4520 -1291 -4474
rect -1245 -4520 -1219 -4474
rect -1317 -4568 -1219 -4520
rect -3068 -4582 -3022 -4571
rect -2908 -4582 -2862 -4571
rect -2748 -4582 -2702 -4571
rect -2588 -4582 -2542 -4571
rect -2428 -4582 -2382 -4571
rect -2268 -4582 -2222 -4571
rect -2108 -4582 -2062 -4571
rect -1948 -4582 -1902 -4571
rect -1788 -4582 -1742 -4571
rect -1628 -4582 -1582 -4571
rect -1468 -4582 -1422 -4571
rect -3293 -4662 -3195 -4614
rect -3293 -4708 -3267 -4662
rect -3221 -4708 -3195 -4662
rect -1317 -4614 -1291 -4568
rect -1245 -4614 -1219 -4568
rect -1317 -4619 -1219 -4614
rect -488 -4307 -462 -4268
rect -416 -4307 -390 -4261
rect -488 -4355 -390 -4307
rect -176 -4238 -66 -4223
rect 187 -4229 267 -4215
rect 187 -4232 200 -4229
rect -176 -4310 -164 -4238
rect -83 -4310 -66 -4238
rect -176 -4325 -66 -4310
rect 82 -4282 200 -4232
rect -488 -4401 -462 -4355
rect -416 -4401 -390 -4355
rect -488 -4449 -390 -4401
rect -488 -4495 -462 -4449
rect -416 -4495 -390 -4449
rect -488 -4543 -390 -4495
rect -488 -4589 -462 -4543
rect -416 -4589 -390 -4543
rect -488 -4619 -390 -4589
rect -1317 -4637 -390 -4619
rect -1317 -4662 -462 -4637
rect -3293 -4756 -3195 -4708
rect -2607 -4682 -2524 -4668
rect -2607 -4738 -2593 -4682
rect -2537 -4738 -2524 -4682
rect -2607 -4750 -2524 -4738
rect -1965 -4682 -1882 -4669
rect -1965 -4738 -1952 -4682
rect -1896 -4738 -1882 -4682
rect -1965 -4751 -1882 -4738
rect -1317 -4708 -1291 -4662
rect -1245 -4683 -462 -4662
rect -416 -4683 -390 -4637
rect -1245 -4708 -390 -4683
rect -1317 -4731 -390 -4708
rect -3293 -4802 -3267 -4756
rect -3221 -4802 -3195 -4756
rect -3293 -4850 -3195 -4802
rect -1317 -4756 -462 -4731
rect -1317 -4802 -1291 -4756
rect -1245 -4766 -462 -4756
rect -1245 -4802 -1219 -4766
rect -3293 -4896 -3267 -4850
rect -3221 -4896 -3195 -4850
rect -3293 -4944 -3195 -4896
rect -2767 -4839 -2684 -4825
rect -2767 -4895 -2753 -4839
rect -2697 -4895 -2684 -4839
rect -2767 -4907 -2684 -4895
rect -2447 -4840 -2364 -4826
rect -2447 -4896 -2433 -4840
rect -2377 -4896 -2364 -4840
rect -2447 -4908 -2364 -4896
rect -2127 -4838 -2044 -4824
rect -2127 -4894 -2113 -4838
rect -2057 -4894 -2044 -4838
rect -2127 -4906 -2044 -4894
rect -1807 -4839 -1724 -4825
rect -1807 -4895 -1793 -4839
rect -1737 -4895 -1724 -4839
rect -1807 -4907 -1724 -4895
rect -1317 -4850 -1219 -4802
rect -1317 -4896 -1291 -4850
rect -1245 -4896 -1219 -4850
rect -3293 -4990 -3267 -4944
rect -3221 -4990 -3195 -4944
rect -1317 -4944 -1219 -4896
rect -3293 -5038 -3195 -4990
rect -3293 -5084 -3267 -5038
rect -3221 -5084 -3195 -5038
rect -3088 -4986 -3004 -4975
rect -3088 -5048 -3077 -4986
rect -3015 -5048 -3004 -4986
rect -3088 -5059 -3004 -5048
rect -2927 -4985 -2843 -4974
rect -2927 -5047 -2916 -4985
rect -2854 -5047 -2843 -4985
rect -2927 -5058 -2843 -5047
rect -2288 -4986 -2202 -4975
rect -2288 -5048 -2276 -4986
rect -2214 -5048 -2202 -4986
rect -2288 -5059 -2202 -5048
rect -1647 -4986 -1563 -4974
rect -1647 -5048 -1636 -4986
rect -1574 -5048 -1563 -4986
rect -1647 -5058 -1563 -5048
rect -1487 -4986 -1403 -4975
rect -1487 -5048 -1476 -4986
rect -1414 -5048 -1403 -4986
rect -1487 -5059 -1403 -5048
rect -1317 -4990 -1291 -4944
rect -1245 -4990 -1219 -4944
rect -1317 -5038 -1219 -4990
rect -3293 -5132 -3195 -5084
rect -3293 -5178 -3267 -5132
rect -3221 -5178 -3195 -5132
rect -1317 -5084 -1291 -5038
rect -1245 -5084 -1219 -5038
rect -1317 -5132 -1219 -5084
rect -3293 -5226 -3195 -5178
rect -3068 -5219 -3022 -5156
rect -2908 -5167 -2862 -5156
rect -2748 -5167 -2702 -5156
rect -2588 -5167 -2542 -5156
rect -2428 -5167 -2382 -5156
rect -2268 -5167 -2222 -5156
rect -2108 -5167 -2062 -5156
rect -1948 -5167 -1902 -5156
rect -1788 -5167 -1742 -5156
rect -1628 -5167 -1582 -5156
rect -3293 -5272 -3267 -5226
rect -3221 -5272 -3195 -5226
rect -3293 -5320 -3195 -5272
rect -3081 -5231 -3009 -5219
rect -1468 -5223 -1422 -5156
rect -1317 -5178 -1291 -5132
rect -1245 -5178 -1219 -5132
rect -3081 -5277 -3068 -5231
rect -3022 -5277 -3009 -5231
rect -1480 -5232 -1410 -5223
rect -3081 -5289 -3009 -5277
rect -2851 -5260 -2750 -5245
rect -2851 -5266 -2829 -5260
rect -3293 -5366 -3267 -5320
rect -3221 -5366 -3195 -5320
rect -2851 -5322 -2830 -5266
rect -2783 -5266 -2750 -5260
rect -2774 -5267 -2750 -5266
rect -2363 -5263 -2285 -5246
rect -2363 -5267 -2348 -5263
rect -2774 -5281 -2348 -5267
rect -2774 -5322 -2668 -5281
rect -2851 -5323 -2668 -5322
rect -2851 -5342 -2750 -5323
rect -2684 -5327 -2668 -5323
rect -2622 -5282 -2348 -5281
rect -2622 -5323 -2508 -5282
rect -2622 -5327 -2606 -5323
rect -2684 -5344 -2606 -5327
rect -2524 -5328 -2508 -5323
rect -2462 -5309 -2348 -5282
rect -2302 -5267 -2285 -5263
rect -2205 -5263 -2127 -5246
rect -2205 -5267 -2188 -5263
rect -2302 -5309 -2188 -5267
rect -2142 -5267 -2127 -5263
rect -1723 -5260 -1645 -5246
rect -1723 -5267 -1707 -5260
rect -2142 -5281 -1707 -5267
rect -2142 -5282 -1868 -5281
rect -2142 -5309 -2028 -5282
rect -2462 -5323 -2028 -5309
rect -2462 -5328 -2446 -5323
rect -2524 -5344 -2446 -5328
rect -2044 -5328 -2028 -5323
rect -1982 -5323 -1868 -5282
rect -1982 -5328 -1966 -5323
rect -2044 -5344 -1966 -5328
rect -1884 -5327 -1868 -5323
rect -1822 -5306 -1707 -5281
rect -1661 -5306 -1645 -5260
rect -1480 -5278 -1468 -5232
rect -1422 -5278 -1410 -5232
rect -1480 -5291 -1410 -5278
rect -1317 -5226 -1219 -5178
rect -1317 -5272 -1291 -5226
rect -1245 -5272 -1219 -5226
rect -1822 -5323 -1645 -5306
rect -1317 -5320 -1219 -5272
rect -1822 -5327 -1806 -5323
rect -1884 -5344 -1806 -5327
rect -3293 -5414 -3195 -5366
rect -3293 -5460 -3267 -5414
rect -3221 -5460 -3195 -5414
rect -1317 -5366 -1291 -5320
rect -1245 -5366 -1219 -5320
rect -1317 -5414 -1219 -5366
rect -3068 -5434 -3022 -5423
rect -2908 -5434 -2862 -5423
rect -2748 -5434 -2702 -5423
rect -2588 -5434 -2542 -5423
rect -2428 -5434 -2382 -5423
rect -2268 -5434 -2222 -5423
rect -2108 -5434 -2062 -5423
rect -1948 -5434 -1902 -5423
rect -1788 -5434 -1742 -5423
rect -1628 -5434 -1582 -5423
rect -1468 -5434 -1422 -5423
rect -3293 -5508 -3195 -5460
rect -3293 -5554 -3267 -5508
rect -3221 -5554 -3195 -5508
rect -1317 -5460 -1291 -5414
rect -1245 -5460 -1219 -5414
rect -1317 -5469 -1219 -5460
rect -488 -4777 -462 -4766
rect -416 -4777 -390 -4731
rect -488 -4825 -390 -4777
rect -488 -4871 -462 -4825
rect -416 -4871 -390 -4825
rect -488 -4919 -390 -4871
rect -488 -4965 -462 -4919
rect -416 -4965 -390 -4919
rect -488 -5013 -390 -4965
rect -488 -5059 -462 -5013
rect -416 -5059 -390 -5013
rect -488 -5107 -390 -5059
rect -488 -5153 -462 -5107
rect -416 -5153 -390 -5107
rect -488 -5201 -390 -5153
rect -488 -5247 -462 -5201
rect -416 -5247 -390 -5201
rect -488 -5295 -390 -5247
rect -488 -5341 -462 -5295
rect -416 -5341 -390 -5295
rect -488 -5389 -390 -5341
rect -488 -5435 -462 -5389
rect -416 -5435 -390 -5389
rect -488 -5469 -390 -5435
rect -1317 -5483 -390 -5469
rect -1317 -5508 -462 -5483
rect -3293 -5602 -3195 -5554
rect -3293 -5648 -3267 -5602
rect -3221 -5648 -3195 -5602
rect -2607 -5542 -2524 -5528
rect -2607 -5598 -2593 -5542
rect -2537 -5598 -2524 -5542
rect -2607 -5610 -2524 -5598
rect -1965 -5542 -1882 -5527
rect -1965 -5598 -1952 -5542
rect -1896 -5598 -1882 -5542
rect -1965 -5611 -1882 -5598
rect -1317 -5554 -1291 -5508
rect -1245 -5529 -462 -5508
rect -416 -5529 -390 -5483
rect -1245 -5554 -390 -5529
rect -1317 -5577 -390 -5554
rect -1317 -5602 -462 -5577
rect -3293 -5696 -3195 -5648
rect -1317 -5648 -1291 -5602
rect -1245 -5616 -462 -5602
rect -1245 -5648 -1219 -5616
rect -3293 -5742 -3267 -5696
rect -3221 -5742 -3195 -5696
rect -3293 -5790 -3195 -5742
rect -2769 -5694 -2686 -5680
rect -2769 -5750 -2755 -5694
rect -2699 -5750 -2686 -5694
rect -2769 -5762 -2686 -5750
rect -2447 -5693 -2364 -5679
rect -2447 -5749 -2433 -5693
rect -2377 -5749 -2364 -5693
rect -2447 -5761 -2364 -5749
rect -2129 -5693 -2046 -5679
rect -2129 -5749 -2115 -5693
rect -2059 -5749 -2046 -5693
rect -2129 -5761 -2046 -5749
rect -1806 -5693 -1723 -5679
rect -1806 -5749 -1792 -5693
rect -1736 -5749 -1723 -5693
rect -1806 -5761 -1723 -5749
rect -1317 -5696 -1219 -5648
rect -1317 -5742 -1291 -5696
rect -1245 -5742 -1219 -5696
rect -3293 -5836 -3267 -5790
rect -3221 -5836 -3195 -5790
rect -1317 -5790 -1219 -5742
rect -3293 -5884 -3195 -5836
rect -3293 -5930 -3267 -5884
rect -3221 -5930 -3195 -5884
rect -3088 -5849 -3004 -5835
rect -3088 -5905 -3074 -5849
rect -3018 -5905 -3004 -5849
rect -3088 -5919 -3004 -5905
rect -2927 -5849 -2843 -5834
rect -2927 -5905 -2913 -5849
rect -2857 -5905 -2843 -5849
rect -2927 -5918 -2843 -5905
rect -2288 -5849 -2202 -5835
rect -2288 -5905 -2274 -5849
rect -2216 -5905 -2202 -5849
rect -2288 -5919 -2202 -5905
rect -1647 -5849 -1563 -5834
rect -1647 -5905 -1633 -5849
rect -1577 -5905 -1563 -5849
rect -1647 -5918 -1563 -5905
rect -1487 -5849 -1403 -5835
rect -1487 -5905 -1473 -5849
rect -1417 -5905 -1403 -5849
rect -1487 -5919 -1403 -5905
rect -1317 -5836 -1291 -5790
rect -1245 -5836 -1219 -5790
rect -1317 -5884 -1219 -5836
rect -3293 -5978 -3195 -5930
rect -3293 -6024 -3267 -5978
rect -3221 -6024 -3195 -5978
rect -1317 -5930 -1291 -5884
rect -1245 -5930 -1219 -5884
rect -1317 -5978 -1219 -5930
rect -3293 -6072 -3195 -6024
rect -3068 -6069 -3022 -6008
rect -2908 -6019 -2862 -6008
rect -2748 -6019 -2702 -6008
rect -2588 -6019 -2542 -6008
rect -2428 -6019 -2382 -6008
rect -2268 -6019 -2222 -6008
rect -2108 -6019 -2062 -6008
rect -1948 -6019 -1902 -6008
rect -1788 -6019 -1742 -6008
rect -1628 -6019 -1582 -6008
rect -3293 -6118 -3267 -6072
rect -3221 -6118 -3195 -6072
rect -3293 -6166 -3195 -6118
rect -3080 -6081 -3011 -6069
rect -3080 -6127 -3068 -6081
rect -3022 -6127 -3011 -6081
rect -1742 -6087 -1641 -6066
rect -1468 -6074 -1422 -6008
rect -1317 -6024 -1291 -5978
rect -1245 -6011 -1219 -5978
rect -488 -5623 -462 -5616
rect -416 -5623 -390 -5577
rect -488 -5671 -390 -5623
rect -488 -5717 -462 -5671
rect -416 -5717 -390 -5671
rect -488 -5765 -390 -5717
rect -488 -5811 -462 -5765
rect -416 -5811 -390 -5765
rect -488 -5859 -390 -5811
rect -488 -5905 -462 -5859
rect -416 -5905 -390 -5859
rect -238 -5142 -188 -4488
rect -78 -5142 -28 -4488
rect -238 -5148 -28 -5142
rect -238 -5194 -156 -5148
rect -110 -5194 -28 -5148
rect -238 -5201 -28 -5194
rect -238 -5868 -188 -5201
rect -488 -5953 -390 -5905
rect -488 -5999 -462 -5953
rect -416 -5999 -390 -5953
rect -488 -6011 -390 -5999
rect -1245 -6024 -390 -6011
rect -1317 -6047 -390 -6024
rect -1317 -6072 -462 -6047
rect -3080 -6139 -3011 -6127
rect -2849 -6093 -1721 -6087
rect -1665 -6093 -1641 -6087
rect -2849 -6139 -2828 -6093
rect -2782 -6139 -2348 -6093
rect -2302 -6139 -2188 -6093
rect -2142 -6139 -1721 -6093
rect -1662 -6139 -1641 -6093
rect -2849 -6143 -1721 -6139
rect -1665 -6143 -1641 -6139
rect -1481 -6085 -1410 -6074
rect -1481 -6131 -1468 -6085
rect -1422 -6131 -1410 -6085
rect -1481 -6143 -1410 -6131
rect -1317 -6118 -1291 -6072
rect -1245 -6093 -462 -6072
rect -416 -6093 -390 -6047
rect -1245 -6118 -390 -6093
rect -78 -6064 -28 -5201
rect 82 -5868 132 -4282
rect 187 -4284 200 -4282
rect 255 -4232 267 -4229
rect 255 -4282 708 -4232
rect 255 -4284 267 -4282
rect 187 -4299 267 -4284
rect 356 -4350 433 -4337
rect 356 -4404 368 -4350
rect 422 -4404 433 -4350
rect 356 -4414 433 -4404
rect 210 -5950 260 -4488
rect 370 -5868 420 -4414
rect 357 -5948 434 -5939
rect 357 -5950 367 -5948
rect 210 -6000 367 -5950
rect 357 -6004 367 -6000
rect 423 -5950 434 -5948
rect 530 -5950 580 -4488
rect 658 -5868 708 -4282
rect 1206 -4261 1304 -4213
rect 1206 -4307 1232 -4261
rect 1278 -4307 1304 -4261
rect 1206 -4355 1304 -4307
rect 1206 -4401 1232 -4355
rect 1278 -4401 1304 -4355
rect 1206 -4449 1304 -4401
rect 818 -5146 868 -4488
rect 978 -5146 1028 -4488
rect 818 -5152 1028 -5146
rect 818 -5198 901 -5152
rect 947 -5198 1028 -5152
rect 818 -5205 1028 -5198
rect 423 -6000 580 -5950
rect 423 -6004 434 -6000
rect 357 -6014 434 -6004
rect 49 -6061 133 -6046
rect 49 -6064 63 -6061
rect -78 -6114 63 -6064
rect -1317 -6141 -390 -6118
rect 49 -6117 63 -6114
rect 119 -6064 133 -6061
rect 818 -6064 868 -5205
rect 978 -5868 1028 -5205
rect 1206 -4495 1232 -4449
rect 1278 -4495 1304 -4449
rect 1206 -4543 1304 -4495
rect 1206 -4589 1232 -4543
rect 1278 -4589 1304 -4543
rect 1206 -4637 1304 -4589
rect 1206 -4683 1232 -4637
rect 1278 -4683 1304 -4637
rect 1206 -4731 1304 -4683
rect 1206 -4777 1232 -4731
rect 1278 -4777 1304 -4731
rect 1206 -4825 1304 -4777
rect 1206 -4871 1232 -4825
rect 1278 -4871 1304 -4825
rect 1206 -4919 1304 -4871
rect 1206 -4965 1232 -4919
rect 1278 -4965 1304 -4919
rect 1206 -5013 1304 -4965
rect 1206 -5059 1232 -5013
rect 1278 -5059 1304 -5013
rect 1206 -5107 1304 -5059
rect 1206 -5153 1232 -5107
rect 1278 -5153 1304 -5107
rect 1206 -5201 1304 -5153
rect 1206 -5247 1232 -5201
rect 1278 -5247 1304 -5201
rect 1206 -5295 1304 -5247
rect 1206 -5341 1232 -5295
rect 1278 -5341 1304 -5295
rect 1206 -5389 1304 -5341
rect 1206 -5435 1232 -5389
rect 1278 -5435 1304 -5389
rect 1206 -5483 1304 -5435
rect 1206 -5529 1232 -5483
rect 1278 -5529 1304 -5483
rect 1206 -5577 1304 -5529
rect 1206 -5623 1232 -5577
rect 1278 -5579 1304 -5577
rect 2934 -5557 4809 -5488
rect 2934 -5579 3066 -5557
rect 1278 -5623 3066 -5579
rect 1206 -5671 3066 -5623
rect 1206 -5717 1232 -5671
rect 1278 -5693 3066 -5671
rect 4667 -5693 4809 -5557
rect 1278 -5711 4809 -5693
rect 1278 -5717 1304 -5711
rect 1206 -5765 1304 -5717
rect 2934 -5749 4809 -5711
rect 1206 -5811 1232 -5765
rect 1278 -5811 1304 -5765
rect 1206 -5859 1304 -5811
rect 119 -6114 868 -6064
rect 1206 -5905 1232 -5859
rect 1278 -5905 1304 -5859
rect 1206 -5953 1304 -5905
rect 1206 -5999 1232 -5953
rect 1278 -5999 1304 -5953
rect 1206 -6047 1304 -5999
rect 3112 -6044 3158 -5749
rect 3486 -6044 3532 -5749
rect 4150 -6045 4196 -5749
rect 4656 -6025 4714 -5749
rect 1206 -6093 1232 -6047
rect 1278 -6093 1304 -6047
rect 4656 -6083 4868 -6025
rect 119 -6117 133 -6114
rect 49 -6131 133 -6117
rect -1742 -6163 -1641 -6143
rect -1317 -6158 -462 -6141
rect -3293 -6212 -3267 -6166
rect -3221 -6212 -3195 -6166
rect -3293 -6234 -3195 -6212
rect -1317 -6166 -1219 -6158
rect -1317 -6212 -1291 -6166
rect -1245 -6212 -1219 -6166
rect -1317 -6234 -1219 -6212
rect -3293 -6260 -1219 -6234
rect -3293 -6306 -3266 -6260
rect -3220 -6306 -3172 -6260
rect -3126 -6306 -3078 -6260
rect -3032 -6306 -2984 -6260
rect -2938 -6306 -2890 -6260
rect -2844 -6306 -2796 -6260
rect -2750 -6306 -2702 -6260
rect -2656 -6306 -2608 -6260
rect -2562 -6306 -2514 -6260
rect -2468 -6306 -2420 -6260
rect -2374 -6306 -2326 -6260
rect -2280 -6306 -2232 -6260
rect -2186 -6306 -2138 -6260
rect -2092 -6306 -2044 -6260
rect -1998 -6306 -1950 -6260
rect -1904 -6306 -1856 -6260
rect -1810 -6306 -1762 -6260
rect -1716 -6306 -1668 -6260
rect -1622 -6306 -1574 -6260
rect -1528 -6306 -1480 -6260
rect -1434 -6306 -1386 -6260
rect -1340 -6306 -1292 -6260
rect -1246 -6306 -1219 -6260
rect -3293 -6332 -1219 -6306
rect -488 -6187 -462 -6158
rect -416 -6187 -390 -6141
rect -488 -6210 -390 -6187
rect 1206 -6141 1304 -6093
rect 1206 -6187 1232 -6141
rect 1278 -6187 1304 -6141
rect 1206 -6210 1304 -6187
rect -488 -6235 1304 -6210
rect -488 -6282 -462 -6235
rect -415 -6236 1231 -6235
rect -415 -6282 -367 -6236
rect -321 -6282 -273 -6236
rect -227 -6282 -179 -6236
rect -133 -6282 -85 -6236
rect -39 -6282 9 -6236
rect 55 -6282 103 -6236
rect 149 -6282 197 -6236
rect 243 -6282 291 -6236
rect 337 -6282 385 -6236
rect 431 -6282 479 -6236
rect 525 -6282 573 -6236
rect 619 -6282 667 -6236
rect 713 -6282 761 -6236
rect 807 -6282 855 -6236
rect 901 -6282 949 -6236
rect 995 -6282 1043 -6236
rect 1089 -6282 1137 -6236
rect 1183 -6282 1231 -6236
rect 1278 -6282 1304 -6235
rect -488 -6308 1304 -6282
rect 4350 -6215 4447 -6200
rect 4350 -6282 4363 -6215
rect 4434 -6282 4447 -6215
rect 4350 -6295 4447 -6282
rect -574 -6512 1287 -6487
rect -574 -6558 -549 -6512
rect -503 -6558 -451 -6512
rect -405 -6558 -353 -6512
rect -307 -6558 -255 -6512
rect -209 -6558 -157 -6512
rect -111 -6558 -59 -6512
rect -13 -6558 39 -6512
rect 85 -6558 137 -6512
rect 183 -6558 235 -6512
rect 281 -6558 333 -6512
rect 379 -6558 431 -6512
rect 477 -6558 529 -6512
rect 575 -6558 627 -6512
rect 673 -6558 725 -6512
rect 771 -6558 823 -6512
rect 869 -6558 921 -6512
rect 967 -6558 1019 -6512
rect 1065 -6558 1117 -6512
rect 1163 -6558 1215 -6512
rect 1261 -6558 1287 -6512
rect -574 -6584 1287 -6558
rect -574 -6610 -477 -6584
rect -574 -6656 -549 -6610
rect -503 -6656 -477 -6610
rect -574 -6708 -477 -6656
rect -574 -6754 -549 -6708
rect -503 -6754 -477 -6708
rect 1190 -6610 1287 -6584
rect 1190 -6656 1215 -6610
rect 1261 -6656 1287 -6610
rect 1190 -6708 1287 -6656
rect -574 -6806 -477 -6754
rect -3320 -6842 -1166 -6817
rect -3320 -6888 -3295 -6842
rect -3249 -6888 -3197 -6842
rect -3151 -6888 -3099 -6842
rect -3053 -6888 -3001 -6842
rect -2955 -6888 -2903 -6842
rect -2857 -6888 -2805 -6842
rect -2759 -6888 -2707 -6842
rect -2661 -6888 -2609 -6842
rect -2563 -6888 -2511 -6842
rect -2465 -6888 -2413 -6842
rect -2367 -6888 -2315 -6842
rect -2269 -6888 -2217 -6842
rect -2171 -6888 -2119 -6842
rect -2073 -6888 -2021 -6842
rect -1975 -6888 -1923 -6842
rect -1877 -6888 -1825 -6842
rect -1779 -6888 -1727 -6842
rect -1681 -6888 -1629 -6842
rect -1583 -6888 -1531 -6842
rect -1485 -6888 -1433 -6842
rect -1387 -6888 -1335 -6842
rect -1289 -6888 -1237 -6842
rect -1191 -6888 -1166 -6842
rect -3320 -6914 -1166 -6888
rect -3320 -6940 -3223 -6914
rect -3320 -6986 -3295 -6940
rect -3249 -6986 -3223 -6940
rect -3320 -7038 -3223 -6986
rect -3320 -7084 -3295 -7038
rect -3249 -7084 -3223 -7038
rect -3320 -7136 -3223 -7084
rect -3060 -7053 -2992 -7040
rect -3060 -7099 -3049 -7053
rect -3003 -7099 -2992 -7053
rect -3060 -7107 -2992 -7099
rect -3320 -7182 -3295 -7136
rect -3249 -7182 -3223 -7136
rect -3049 -7141 -3003 -7107
rect -3320 -7234 -3223 -7182
rect -3320 -7280 -3295 -7234
rect -3249 -7280 -3223 -7234
rect -3320 -7332 -3223 -7280
rect -3067 -7227 -2984 -7214
rect -3067 -7283 -3053 -7227
rect -2997 -7283 -2984 -7227
rect -3067 -7296 -2984 -7283
rect -2907 -7229 -2824 -7216
rect -2907 -7285 -2893 -7229
rect -2837 -7285 -2824 -7229
rect -2907 -7298 -2824 -7285
rect -3320 -7378 -3295 -7332
rect -3249 -7378 -3223 -7332
rect -3320 -7430 -3223 -7378
rect -3320 -7476 -3295 -7430
rect -3249 -7476 -3223 -7430
rect -3320 -7528 -3223 -7476
rect -3320 -7574 -3295 -7528
rect -3249 -7574 -3223 -7528
rect -3320 -7626 -3223 -7574
rect -3320 -7672 -3295 -7626
rect -3249 -7672 -3223 -7626
rect -3320 -7724 -3223 -7672
rect -3320 -7770 -3295 -7724
rect -3249 -7770 -3223 -7724
rect -3320 -7822 -3223 -7770
rect -3320 -7868 -3295 -7822
rect -3249 -7868 -3223 -7822
rect -3320 -7920 -3223 -7868
rect -3060 -7853 -2992 -7840
rect -3060 -7899 -3049 -7853
rect -3003 -7899 -2992 -7853
rect -3060 -7907 -2992 -7899
rect -3320 -7966 -3295 -7920
rect -3249 -7966 -3223 -7920
rect -3049 -7941 -3003 -7907
rect -3320 -8018 -3223 -7966
rect -3320 -8064 -3295 -8018
rect -3249 -8064 -3223 -8018
rect -3320 -8116 -3223 -8064
rect -3066 -8029 -2983 -8016
rect -3066 -8085 -3052 -8029
rect -2996 -8085 -2983 -8029
rect -3066 -8098 -2983 -8085
rect -2907 -8030 -2824 -8017
rect -2907 -8086 -2893 -8030
rect -2837 -8086 -2824 -8030
rect -2907 -8099 -2824 -8086
rect -3320 -8162 -3295 -8116
rect -3249 -8162 -3223 -8116
rect -3320 -8214 -3223 -8162
rect -3320 -8260 -3295 -8214
rect -3249 -8260 -3223 -8214
rect -3320 -8312 -3223 -8260
rect -3320 -8358 -3295 -8312
rect -3249 -8358 -3223 -8312
rect -3320 -8410 -3223 -8358
rect -3320 -8456 -3295 -8410
rect -3249 -8456 -3223 -8410
rect -3320 -8508 -3223 -8456
rect -3320 -8554 -3295 -8508
rect -3249 -8554 -3223 -8508
rect -3320 -8606 -3223 -8554
rect -3320 -8652 -3295 -8606
rect -3249 -8652 -3223 -8606
rect -3320 -8704 -3223 -8652
rect -3320 -8750 -3295 -8704
rect -3249 -8750 -3223 -8704
rect -3060 -8651 -2992 -8638
rect -3060 -8697 -3049 -8651
rect -3003 -8697 -2992 -8651
rect -3060 -8705 -2992 -8697
rect -3049 -8750 -3003 -8705
rect -2889 -8750 -2843 -8739
rect -3320 -8802 -3223 -8750
rect -3320 -8848 -3295 -8802
rect -3249 -8848 -3223 -8802
rect -3320 -8900 -3223 -8848
rect -3069 -8831 -2986 -8818
rect -3069 -8887 -3055 -8831
rect -2999 -8887 -2986 -8831
rect -3069 -8900 -2986 -8887
rect -2907 -8831 -2824 -8818
rect -2907 -8887 -2893 -8831
rect -2837 -8887 -2824 -8831
rect -2907 -8900 -2824 -8887
rect -3320 -8946 -3295 -8900
rect -3249 -8946 -3223 -8900
rect -3320 -8998 -3223 -8946
rect -3320 -9044 -3295 -8998
rect -3249 -9044 -3223 -8998
rect -3320 -9096 -3223 -9044
rect -3320 -9142 -3295 -9096
rect -3249 -9142 -3223 -9096
rect -3320 -9194 -3223 -9142
rect -3320 -9240 -3295 -9194
rect -3249 -9240 -3223 -9194
rect -3320 -9292 -3223 -9240
rect -3320 -9338 -3295 -9292
rect -3249 -9338 -3223 -9292
rect -3049 -9335 -3003 -9324
rect -2889 -9335 -2843 -9324
rect -3320 -9390 -3223 -9338
rect -3320 -9436 -3295 -9390
rect -3249 -9436 -3223 -9390
rect -3320 -9488 -3223 -9436
rect -3320 -9534 -3295 -9488
rect -3249 -9534 -3223 -9488
rect -3060 -9451 -2992 -9438
rect -3060 -9497 -3049 -9451
rect -3003 -9497 -2992 -9451
rect -3060 -9505 -2992 -9497
rect -3320 -9586 -3223 -9534
rect -3049 -9550 -3003 -9505
rect -2889 -9550 -2843 -9539
rect -3320 -9632 -3295 -9586
rect -3249 -9632 -3223 -9586
rect -3320 -9684 -3223 -9632
rect -3320 -9730 -3295 -9684
rect -3249 -9730 -3223 -9684
rect -3069 -9630 -2986 -9617
rect -3069 -9686 -3055 -9630
rect -2999 -9686 -2986 -9630
rect -3069 -9699 -2986 -9686
rect -2907 -9632 -2824 -9619
rect -2907 -9688 -2893 -9632
rect -2837 -9688 -2824 -9632
rect -2907 -9701 -2824 -9688
rect -3320 -9782 -3223 -9730
rect -3320 -9828 -3295 -9782
rect -3249 -9828 -3223 -9782
rect -3320 -9880 -3223 -9828
rect -3320 -9926 -3295 -9880
rect -3249 -9926 -3223 -9880
rect -3320 -9978 -3223 -9926
rect -3320 -10024 -3295 -9978
rect -3249 -10024 -3223 -9978
rect -3320 -10076 -3223 -10024
rect -3320 -10122 -3295 -10076
rect -3249 -10122 -3223 -10076
rect -3320 -10174 -3223 -10122
rect -3049 -10135 -3003 -10124
rect -2889 -10135 -2843 -10124
rect -3320 -10220 -3295 -10174
rect -3249 -10220 -3223 -10174
rect -3320 -10272 -3223 -10220
rect -3320 -10318 -3295 -10272
rect -3249 -10318 -3223 -10272
rect -3320 -10344 -3223 -10318
rect -2731 -10344 -2681 -6914
rect -2587 -7542 -2504 -7529
rect -2587 -7598 -2573 -7542
rect -2517 -7598 -2504 -7542
rect -2587 -7611 -2504 -7598
rect -2587 -8343 -2504 -8330
rect -2587 -8399 -2573 -8343
rect -2517 -8399 -2504 -8343
rect -2587 -8412 -2504 -8399
rect -2569 -8750 -2523 -8739
rect -2587 -9144 -2504 -9131
rect -2587 -9200 -2573 -9144
rect -2517 -9200 -2504 -9144
rect -2587 -9213 -2504 -9200
rect -2569 -9335 -2523 -9324
rect -2569 -9550 -2523 -9539
rect -2587 -9945 -2504 -9932
rect -2587 -10001 -2573 -9945
rect -2517 -10001 -2504 -9945
rect -2587 -10014 -2504 -10001
rect -2569 -10135 -2523 -10124
rect -2411 -10344 -2361 -6914
rect -2249 -7152 -2203 -7141
rect -2268 -7229 -2185 -7216
rect -2268 -7285 -2254 -7229
rect -2198 -7285 -2185 -7229
rect -2268 -7298 -2185 -7285
rect -2249 -7737 -2203 -7726
rect -2268 -7809 -2184 -7797
rect -2268 -7869 -2256 -7809
rect -2196 -7869 -2184 -7809
rect -2268 -7881 -2184 -7869
rect -2249 -7952 -2203 -7941
rect -2268 -8030 -2185 -8017
rect -2268 -8086 -2254 -8030
rect -2198 -8086 -2185 -8030
rect -2268 -8099 -2185 -8086
rect -2249 -8537 -2203 -8526
rect -2268 -8610 -2184 -8598
rect -2268 -8670 -2256 -8610
rect -2196 -8670 -2184 -8610
rect -2268 -8682 -2184 -8670
rect -2249 -8750 -2203 -8739
rect -2268 -8831 -2185 -8818
rect -2268 -8887 -2254 -8831
rect -2198 -8887 -2185 -8831
rect -2268 -8900 -2185 -8887
rect -2249 -9335 -2203 -9324
rect -2269 -9410 -2185 -9398
rect -2269 -9470 -2257 -9410
rect -2197 -9470 -2185 -9410
rect -2269 -9482 -2185 -9470
rect -2249 -9550 -2203 -9539
rect -2268 -9632 -2185 -9619
rect -2268 -9688 -2254 -9632
rect -2198 -9688 -2185 -9632
rect -2268 -9701 -2185 -9688
rect -2249 -10135 -2203 -10124
rect -2091 -10344 -2041 -6914
rect -1929 -7152 -1883 -7141
rect -1949 -7543 -1866 -7530
rect -1949 -7599 -1935 -7543
rect -1879 -7599 -1866 -7543
rect -1949 -7612 -1866 -7599
rect -1929 -7737 -1883 -7726
rect -1929 -7952 -1883 -7941
rect -1949 -8344 -1866 -8331
rect -1949 -8400 -1935 -8344
rect -1879 -8400 -1866 -8344
rect -1949 -8413 -1866 -8400
rect -1929 -8537 -1883 -8526
rect -1929 -8750 -1883 -8739
rect -1949 -9145 -1866 -9132
rect -1949 -9201 -1935 -9145
rect -1879 -9201 -1866 -9145
rect -1949 -9214 -1866 -9201
rect -1929 -9335 -1883 -9324
rect -1929 -9550 -1883 -9539
rect -1949 -9946 -1866 -9933
rect -1949 -10002 -1935 -9946
rect -1879 -10002 -1866 -9946
rect -1949 -10015 -1866 -10002
rect -1929 -10135 -1883 -10124
rect -1771 -10344 -1721 -6914
rect -1263 -6940 -1166 -6914
rect -1263 -6986 -1237 -6940
rect -1191 -6982 -1166 -6940
rect -574 -6852 -549 -6806
rect -503 -6852 -477 -6806
rect -574 -6904 -477 -6852
rect -164 -6760 844 -6714
rect -164 -6863 -118 -6760
rect 127 -6824 229 -6811
rect 127 -6829 143 -6824
rect -574 -6950 -549 -6904
rect -503 -6950 -477 -6904
rect -574 -6982 -477 -6950
rect -1191 -6986 -477 -6982
rect -1263 -7002 -477 -6986
rect -324 -6909 -245 -6863
rect -199 -6909 -118 -6863
rect -324 -6990 -278 -6909
rect -323 -7001 -278 -6990
rect -164 -6992 -118 -6909
rect -4 -6875 143 -6829
rect -4 -6984 42 -6875
rect 127 -6880 143 -6875
rect 215 -6829 229 -6824
rect 215 -6875 684 -6829
rect 215 -6880 229 -6875
rect 127 -6894 229 -6880
rect 638 -6984 684 -6875
rect 798 -6885 844 -6760
rect 1190 -6754 1215 -6708
rect 1261 -6754 1287 -6708
rect 3675 -6551 3777 -6530
rect 3675 -6709 3691 -6551
rect 3759 -6709 3777 -6551
rect 3675 -6724 3777 -6709
rect 1190 -6806 1287 -6754
rect 1190 -6852 1215 -6806
rect 1261 -6852 1287 -6806
rect 798 -6931 878 -6885
rect 924 -6931 1004 -6885
rect 798 -6992 844 -6931
rect 958 -6988 1004 -6931
rect 960 -6997 1004 -6988
rect 1190 -6904 1287 -6852
rect 1190 -6950 1215 -6904
rect 1261 -6950 1287 -6904
rect -1263 -7038 -549 -7002
rect -1460 -7053 -1392 -7040
rect -1460 -7099 -1449 -7053
rect -1403 -7099 -1392 -7053
rect -1460 -7107 -1392 -7099
rect -1263 -7084 -1237 -7038
rect -1191 -7048 -549 -7038
rect -503 -7048 -477 -7002
rect 1190 -7002 1287 -6950
rect -1191 -7084 -477 -7048
rect -1263 -7100 -477 -7084
rect -1263 -7104 -549 -7100
rect -1609 -7152 -1563 -7141
rect -1449 -7152 -1403 -7107
rect -1263 -7136 -1166 -7104
rect -1263 -7182 -1237 -7136
rect -1191 -7182 -1166 -7136
rect -1629 -7228 -1546 -7215
rect -1629 -7284 -1615 -7228
rect -1559 -7284 -1546 -7228
rect -1629 -7297 -1546 -7284
rect -1471 -7230 -1388 -7217
rect -1471 -7286 -1457 -7230
rect -1401 -7286 -1388 -7230
rect -1471 -7299 -1388 -7286
rect -1263 -7234 -1166 -7182
rect -1263 -7280 -1237 -7234
rect -1191 -7280 -1166 -7234
rect -1263 -7332 -1166 -7280
rect -1263 -7378 -1237 -7332
rect -1191 -7378 -1166 -7332
rect -1263 -7430 -1166 -7378
rect -1263 -7476 -1237 -7430
rect -1191 -7476 -1166 -7430
rect -1263 -7528 -1166 -7476
rect -1263 -7574 -1237 -7528
rect -1191 -7574 -1166 -7528
rect -1263 -7626 -1166 -7574
rect -1263 -7672 -1237 -7626
rect -1191 -7672 -1166 -7626
rect -1263 -7687 -1166 -7672
rect -574 -7146 -549 -7104
rect -503 -7146 -477 -7100
rect -184 -7047 -99 -7032
rect -184 -7129 -169 -7047
rect -113 -7129 -99 -7047
rect -184 -7142 -99 -7129
rect 1190 -7048 1215 -7002
rect 1261 -7048 1287 -7002
rect 1190 -7100 1287 -7048
rect -574 -7198 -477 -7146
rect -574 -7244 -549 -7198
rect -503 -7244 -477 -7198
rect 1190 -7146 1215 -7100
rect 1261 -7146 1287 -7100
rect 2301 -6913 2561 -6869
rect 2896 -6913 2942 -6840
rect 4810 -6845 4868 -6083
rect 5031 -6899 5077 -6840
rect 5014 -6912 5094 -6899
rect 2301 -6920 2958 -6913
rect 2301 -7089 2349 -6920
rect 2506 -6927 2958 -6920
rect 2506 -6979 2893 -6927
rect 2945 -6959 2958 -6927
rect 2945 -6979 4337 -6959
rect 5014 -6960 5026 -6912
rect 5082 -6960 5094 -6912
rect 5014 -6972 5094 -6960
rect 2506 -7002 4337 -6979
rect 2506 -7061 3012 -7002
rect 3086 -7008 4224 -7002
rect 3086 -7061 3582 -7008
rect 2506 -7067 3582 -7061
rect 3656 -7061 4224 -7008
rect 4298 -7061 4337 -7002
rect 3656 -7067 4337 -7061
rect 2506 -7068 4337 -7067
rect 2506 -7082 4325 -7068
rect 2506 -7089 2561 -7082
rect 2301 -7126 2561 -7089
rect 1190 -7198 1287 -7146
rect 3914 -7197 4022 -7182
rect -574 -7296 -477 -7244
rect -574 -7342 -549 -7296
rect -503 -7342 -477 -7296
rect 298 -7215 381 -7199
rect 298 -7287 312 -7215
rect 368 -7287 381 -7215
rect 298 -7301 381 -7287
rect 1190 -7244 1215 -7198
rect 1261 -7244 1287 -7198
rect 3262 -7218 3366 -7198
rect 3914 -7209 3934 -7197
rect 3262 -7223 3274 -7218
rect 1190 -7296 1287 -7244
rect -574 -7394 -477 -7342
rect -574 -7440 -549 -7394
rect -503 -7440 -477 -7394
rect -574 -7492 -477 -7440
rect -574 -7538 -549 -7492
rect -503 -7538 -477 -7492
rect -574 -7590 -477 -7538
rect 1190 -7342 1215 -7296
rect 1261 -7342 1287 -7296
rect 1190 -7394 1287 -7342
rect 1190 -7440 1215 -7394
rect 1261 -7440 1287 -7394
rect 1190 -7492 1287 -7440
rect 1190 -7538 1215 -7492
rect 1261 -7538 1287 -7492
rect -574 -7636 -549 -7590
rect -503 -7636 -477 -7590
rect -574 -7687 -477 -7636
rect -1263 -7688 -477 -7687
rect -1263 -7724 -549 -7688
rect -1609 -7737 -1563 -7726
rect -1449 -7737 -1403 -7726
rect -1263 -7770 -1237 -7724
rect -1191 -7734 -549 -7724
rect -503 -7734 -477 -7688
rect 157 -7693 203 -7579
rect -1191 -7770 -477 -7734
rect -1263 -7786 -477 -7770
rect -1263 -7809 -549 -7786
rect -1263 -7822 -1166 -7809
rect -1460 -7853 -1392 -7840
rect -1460 -7899 -1449 -7853
rect -1403 -7899 -1392 -7853
rect -1460 -7907 -1392 -7899
rect -1263 -7868 -1237 -7822
rect -1191 -7868 -1166 -7822
rect -1609 -7952 -1563 -7941
rect -1449 -7952 -1403 -7907
rect -1263 -7920 -1166 -7868
rect -1263 -7966 -1237 -7920
rect -1191 -7966 -1166 -7920
rect -1629 -8029 -1546 -8016
rect -1629 -8085 -1615 -8029
rect -1559 -8085 -1546 -8029
rect -1629 -8098 -1546 -8085
rect -1470 -8030 -1387 -8017
rect -1470 -8086 -1456 -8030
rect -1400 -8086 -1387 -8030
rect -1470 -8099 -1387 -8086
rect -1263 -8018 -1166 -7966
rect -1263 -8064 -1237 -8018
rect -1191 -8064 -1166 -8018
rect -1263 -8116 -1166 -8064
rect -1263 -8162 -1237 -8116
rect -1191 -8162 -1166 -8116
rect -1263 -8191 -1166 -8162
rect -574 -7832 -549 -7809
rect -503 -7832 -477 -7786
rect -574 -7884 -477 -7832
rect -324 -7771 -243 -7725
rect -197 -7771 -118 -7725
rect -324 -7835 -278 -7771
rect -574 -7930 -549 -7884
rect -503 -7930 -477 -7884
rect -574 -7982 -477 -7930
rect -574 -8028 -549 -7982
rect -503 -8028 -477 -7982
rect -574 -8080 -477 -8028
rect -574 -8126 -549 -8080
rect -503 -8126 -477 -8080
rect -574 -8178 -477 -8126
rect -574 -8191 -549 -8178
rect -1263 -8214 -549 -8191
rect -1263 -8260 -1237 -8214
rect -1191 -8224 -549 -8214
rect -503 -8224 -477 -8178
rect -1191 -8260 -477 -8224
rect -1263 -8276 -477 -8260
rect -1263 -8312 -549 -8276
rect -1263 -8358 -1237 -8312
rect -1191 -8313 -549 -8312
rect -1191 -8358 -1166 -8313
rect -1263 -8410 -1166 -8358
rect -1263 -8456 -1237 -8410
rect -1191 -8456 -1166 -8410
rect -1263 -8508 -1166 -8456
rect -1609 -8537 -1563 -8526
rect -1449 -8537 -1403 -8526
rect -1263 -8554 -1237 -8508
rect -1191 -8554 -1166 -8508
rect -1263 -8606 -1166 -8554
rect -1460 -8651 -1392 -8638
rect -1460 -8697 -1449 -8651
rect -1403 -8697 -1392 -8651
rect -1460 -8705 -1392 -8697
rect -1263 -8652 -1237 -8606
rect -1191 -8652 -1166 -8606
rect -1263 -8704 -1166 -8652
rect -1609 -8750 -1563 -8739
rect -1449 -8750 -1403 -8705
rect -1263 -8750 -1237 -8704
rect -1191 -8750 -1166 -8704
rect -1263 -8787 -1166 -8750
rect -574 -8322 -549 -8313
rect -503 -8322 -477 -8276
rect -164 -8279 -118 -7771
rect -4 -7739 203 -7693
rect 297 -7677 387 -7665
rect -574 -8374 -477 -8322
rect -574 -8420 -549 -8374
rect -503 -8420 -477 -8374
rect -183 -8295 -100 -8279
rect -183 -8367 -169 -8295
rect -113 -8367 -100 -8295
rect -183 -8381 -100 -8367
rect -574 -8472 -477 -8420
rect -574 -8518 -549 -8472
rect -503 -8518 -477 -8472
rect -574 -8570 -477 -8518
rect -574 -8616 -549 -8570
rect -503 -8616 -477 -8570
rect -574 -8668 -477 -8616
rect -574 -8714 -549 -8668
rect -503 -8714 -477 -8668
rect -574 -8766 -477 -8714
rect -574 -8787 -549 -8766
rect -1263 -8802 -549 -8787
rect -1629 -8830 -1546 -8817
rect -1629 -8886 -1615 -8830
rect -1559 -8886 -1546 -8830
rect -1629 -8899 -1546 -8886
rect -1468 -8830 -1385 -8817
rect -1468 -8886 -1454 -8830
rect -1398 -8886 -1385 -8830
rect -1468 -8899 -1385 -8886
rect -1263 -8848 -1237 -8802
rect -1191 -8812 -549 -8802
rect -503 -8812 -477 -8766
rect -1191 -8848 -477 -8812
rect -1263 -8864 -477 -8848
rect -1263 -8900 -549 -8864
rect -1263 -8946 -1237 -8900
rect -1191 -8909 -549 -8900
rect -1191 -8946 -1166 -8909
rect -1263 -8998 -1166 -8946
rect -1263 -9044 -1237 -8998
rect -1191 -9044 -1166 -8998
rect -1263 -9096 -1166 -9044
rect -1263 -9142 -1237 -9096
rect -1191 -9142 -1166 -9096
rect -1263 -9194 -1166 -9142
rect -1263 -9240 -1237 -9194
rect -1191 -9240 -1166 -9194
rect -1263 -9270 -1166 -9240
rect -574 -8910 -549 -8909
rect -503 -8910 -477 -8864
rect -574 -8962 -477 -8910
rect -574 -9008 -549 -8962
rect -503 -9008 -477 -8962
rect -574 -9060 -477 -9008
rect -574 -9106 -549 -9060
rect -503 -9106 -477 -9060
rect -574 -9158 -477 -9106
rect -574 -9204 -549 -9158
rect -503 -9204 -477 -9158
rect -574 -9256 -477 -9204
rect -574 -9270 -549 -9256
rect -1263 -9292 -549 -9270
rect -1609 -9335 -1563 -9324
rect -1449 -9335 -1403 -9324
rect -1263 -9338 -1237 -9292
rect -1191 -9302 -549 -9292
rect -503 -9302 -477 -9256
rect -1191 -9338 -477 -9302
rect -1263 -9354 -477 -9338
rect -1263 -9390 -549 -9354
rect -1263 -9436 -1237 -9390
rect -1191 -9392 -549 -9390
rect -1191 -9436 -1166 -9392
rect -1460 -9451 -1392 -9438
rect -1460 -9497 -1449 -9451
rect -1403 -9497 -1392 -9451
rect -1460 -9505 -1392 -9497
rect -1263 -9488 -1166 -9436
rect -1609 -9550 -1563 -9539
rect -1449 -9550 -1403 -9505
rect -1263 -9534 -1237 -9488
rect -1191 -9534 -1166 -9488
rect -1263 -9586 -1166 -9534
rect -1629 -9631 -1546 -9618
rect -1629 -9687 -1615 -9631
rect -1559 -9687 -1546 -9631
rect -1629 -9700 -1546 -9687
rect -1469 -9630 -1386 -9617
rect -1469 -9686 -1455 -9630
rect -1399 -9686 -1386 -9630
rect -1469 -9699 -1386 -9686
rect -1263 -9632 -1237 -9586
rect -1191 -9632 -1166 -9586
rect -1263 -9684 -1166 -9632
rect -1263 -9730 -1237 -9684
rect -1191 -9730 -1166 -9684
rect -1263 -9744 -1166 -9730
rect -574 -9400 -549 -9392
rect -503 -9400 -477 -9354
rect -574 -9452 -477 -9400
rect -574 -9498 -549 -9452
rect -503 -9498 -477 -9452
rect -574 -9550 -477 -9498
rect -324 -9468 -278 -9410
rect -164 -9468 -118 -8381
rect -4 -8645 42 -7739
rect 297 -7743 309 -7677
rect 375 -7743 387 -7677
rect 477 -7693 523 -7569
rect 1190 -7590 1287 -7538
rect 1190 -7636 1215 -7590
rect 1261 -7636 1287 -7590
rect 3016 -7296 3274 -7223
rect 3352 -7296 3366 -7218
rect 3016 -7301 3366 -7296
rect 3016 -7398 3094 -7301
rect 3262 -7310 3366 -7301
rect 3749 -7265 3934 -7209
rect 4001 -7265 4022 -7197
rect 5029 -7225 5075 -6972
rect 3749 -7270 4022 -7265
rect 3016 -7410 3376 -7398
rect 3749 -7399 3810 -7270
rect 3914 -7280 4022 -7270
rect 4979 -7250 5111 -7225
rect 4979 -7274 5000 -7250
rect 4186 -7320 5000 -7274
rect 3016 -7470 3310 -7410
rect 3363 -7470 3376 -7410
rect 3016 -7476 3376 -7470
rect 1190 -7688 1287 -7636
rect 477 -7739 684 -7693
rect 297 -7755 387 -7743
rect 157 -7897 203 -7834
rect 139 -7913 222 -7897
rect 139 -7985 153 -7913
rect 209 -7985 222 -7913
rect 139 -7999 222 -7985
rect 157 -8489 203 -7999
rect 317 -8067 363 -7834
rect 289 -8080 391 -8067
rect 289 -8136 305 -8080
rect 377 -8136 391 -8080
rect 289 -8150 391 -8136
rect 317 -8410 363 -8150
rect 477 -8488 523 -7834
rect 134 -8505 217 -8489
rect 134 -8577 148 -8505
rect 204 -8577 217 -8505
rect 134 -8591 217 -8577
rect 460 -8504 543 -8488
rect 460 -8576 474 -8504
rect 530 -8576 543 -8504
rect 460 -8590 543 -8576
rect -23 -8661 60 -8645
rect -23 -8733 -9 -8661
rect 47 -8733 60 -8661
rect -23 -8747 60 -8733
rect -324 -9514 -243 -9468
rect -197 -9514 -118 -9468
rect -4 -9509 42 -8747
rect 157 -9410 203 -8591
rect 317 -9085 363 -8824
rect 288 -9098 390 -9085
rect 288 -9154 304 -9098
rect 376 -9154 390 -9098
rect 288 -9168 390 -9154
rect 317 -9410 363 -9168
rect 477 -9212 523 -8590
rect 638 -8645 684 -7739
rect 1190 -7734 1215 -7688
rect 1261 -7734 1287 -7688
rect 1372 -7622 1494 -7595
rect 3016 -7598 3094 -7476
rect 3298 -7482 3376 -7476
rect 3742 -7412 3818 -7399
rect 3742 -7471 3754 -7412
rect 3806 -7471 3818 -7412
rect 3313 -7542 3359 -7482
rect 3742 -7483 3818 -7471
rect 3757 -7538 3803 -7483
rect 4186 -7537 4232 -7320
rect 4979 -7333 5000 -7320
rect 5089 -7333 5111 -7250
rect 4979 -7354 5111 -7333
rect 1372 -7696 1396 -7622
rect 1469 -7696 1494 -7622
rect 1372 -7719 1494 -7696
rect 3001 -7618 3109 -7598
rect 3001 -7696 3016 -7618
rect 3095 -7696 3109 -7618
rect 3001 -7712 3109 -7696
rect 798 -7789 877 -7743
rect 923 -7789 1004 -7743
rect 798 -8284 844 -7789
rect 958 -7843 1004 -7789
rect 1190 -7786 1287 -7734
rect 1190 -7832 1215 -7786
rect 1261 -7832 1287 -7786
rect 1190 -7884 1287 -7832
rect 1190 -7930 1215 -7884
rect 1261 -7930 1287 -7884
rect 1190 -7982 1287 -7930
rect 1190 -8028 1215 -7982
rect 1261 -8028 1287 -7982
rect 1190 -8080 1287 -8028
rect 1190 -8126 1215 -8080
rect 1261 -8126 1287 -8080
rect 3529 -8109 3575 -7932
rect 3973 -8109 4019 -7933
rect 4402 -8109 4448 -7933
rect 1190 -8160 1287 -8126
rect 2973 -8156 4757 -8109
rect 2973 -8160 3076 -8156
rect 1190 -8178 3076 -8160
rect 1190 -8224 1215 -8178
rect 1261 -8224 3076 -8178
rect 1190 -8263 3076 -8224
rect 1190 -8276 1287 -8263
rect 779 -8300 862 -8284
rect 779 -8372 793 -8300
rect 849 -8372 862 -8300
rect 779 -8386 862 -8372
rect 1190 -8322 1215 -8276
rect 1261 -8322 1287 -8276
rect 1190 -8374 1287 -8322
rect 2973 -8294 3076 -8263
rect 4649 -8294 4757 -8156
rect 2973 -8344 4757 -8294
rect 620 -8661 703 -8645
rect 620 -8733 634 -8661
rect 690 -8733 703 -8661
rect 620 -8747 703 -8733
rect 457 -9228 540 -9212
rect 457 -9300 471 -9228
rect 527 -9300 540 -9228
rect 457 -9314 540 -9300
rect 477 -9410 523 -9314
rect 288 -9506 378 -9494
rect -574 -9596 -549 -9550
rect -503 -9596 -477 -9550
rect -4 -9555 203 -9509
rect -574 -9648 -477 -9596
rect -574 -9694 -549 -9648
rect -503 -9694 -477 -9648
rect 157 -9681 203 -9555
rect 288 -9572 300 -9506
rect 366 -9572 378 -9506
rect 638 -9509 684 -8747
rect 288 -9584 378 -9572
rect 477 -9555 684 -9509
rect 798 -9473 844 -8386
rect 1190 -8420 1215 -8374
rect 1261 -8420 1287 -8374
rect 1190 -8472 1287 -8420
rect 1190 -8518 1215 -8472
rect 1261 -8518 1287 -8472
rect 1190 -8570 1287 -8518
rect 892 -8588 982 -8576
rect 892 -8654 904 -8588
rect 970 -8654 982 -8588
rect 892 -8666 982 -8654
rect 1190 -8616 1215 -8570
rect 1261 -8616 1287 -8570
rect 1190 -8668 1287 -8616
rect 1190 -8714 1215 -8668
rect 1261 -8714 1287 -8668
rect 1190 -8766 1287 -8714
rect 1190 -8812 1215 -8766
rect 1261 -8812 1287 -8766
rect 1190 -8864 1287 -8812
rect 1190 -8910 1215 -8864
rect 1261 -8910 1287 -8864
rect 1190 -8962 1287 -8910
rect 1190 -9008 1215 -8962
rect 1261 -9008 1287 -8962
rect 1190 -9060 1287 -9008
rect 1190 -9106 1215 -9060
rect 1261 -9106 1287 -9060
rect 1190 -9158 1287 -9106
rect 1190 -9204 1215 -9158
rect 1261 -9204 1287 -9158
rect 1190 -9256 1287 -9204
rect 1190 -9302 1215 -9256
rect 1261 -9302 1287 -9256
rect 1190 -9354 1287 -9302
rect 1190 -9400 1215 -9354
rect 1261 -9400 1287 -9354
rect 958 -9473 1004 -9410
rect 798 -9474 1004 -9473
rect 798 -9520 880 -9474
rect 926 -9520 1004 -9474
rect 1190 -9452 1287 -9400
rect 1190 -9498 1215 -9452
rect 1261 -9498 1287 -9452
rect 1190 -9550 1287 -9498
rect 477 -9681 523 -9555
rect 1190 -9596 1215 -9550
rect 1261 -9596 1287 -9550
rect 1190 -9648 1287 -9596
rect -574 -9744 -477 -9694
rect -1263 -9746 -477 -9744
rect -1263 -9782 -549 -9746
rect -1263 -9828 -1237 -9782
rect -1191 -9792 -549 -9782
rect -503 -9792 -477 -9746
rect -1191 -9828 -477 -9792
rect 1190 -9694 1215 -9648
rect 1261 -9694 1287 -9648
rect 1190 -9746 1287 -9694
rect 1190 -9792 1215 -9746
rect 1261 -9792 1287 -9746
rect -1263 -9844 -477 -9828
rect -1263 -9866 -549 -9844
rect -1263 -9880 -1166 -9866
rect -1263 -9926 -1237 -9880
rect -1191 -9926 -1166 -9880
rect -1263 -9978 -1166 -9926
rect -1263 -10024 -1237 -9978
rect -1191 -10024 -1166 -9978
rect -1263 -10076 -1166 -10024
rect -1263 -10122 -1237 -10076
rect -1191 -10122 -1166 -10076
rect -1609 -10135 -1563 -10124
rect -1449 -10135 -1403 -10124
rect -1263 -10174 -1166 -10122
rect -1263 -10220 -1237 -10174
rect -1191 -10191 -1166 -10174
rect -574 -9890 -549 -9866
rect -503 -9890 -477 -9844
rect -574 -9942 -477 -9890
rect 299 -9835 382 -9819
rect 299 -9907 313 -9835
rect 369 -9907 382 -9835
rect 299 -9921 382 -9907
rect 1190 -9844 1287 -9792
rect 1190 -9890 1215 -9844
rect 1261 -9890 1287 -9844
rect -574 -9988 -549 -9942
rect -503 -9988 -477 -9942
rect -574 -10040 -477 -9988
rect 1190 -9942 1287 -9890
rect 1190 -9988 1215 -9942
rect 1261 -9988 1287 -9942
rect -574 -10086 -549 -10040
rect -503 -10086 -477 -10040
rect -574 -10138 -477 -10086
rect -184 -10036 -99 -10021
rect -184 -10118 -169 -10036
rect -113 -10118 -99 -10036
rect -184 -10131 -99 -10118
rect 1190 -10040 1287 -9988
rect 1190 -10086 1215 -10040
rect 1261 -10086 1287 -10040
rect -574 -10184 -549 -10138
rect -503 -10184 -477 -10138
rect -574 -10191 -477 -10184
rect -1191 -10220 -477 -10191
rect -1263 -10236 -477 -10220
rect -1263 -10272 -549 -10236
rect -1263 -10318 -1237 -10272
rect -1191 -10282 -549 -10272
rect -503 -10282 -477 -10236
rect 1190 -10138 1287 -10086
rect 1190 -10184 1215 -10138
rect 1261 -10184 1287 -10138
rect 1190 -10236 1287 -10184
rect -1191 -10313 -477 -10282
rect -1191 -10318 -1166 -10313
rect -1263 -10344 -1166 -10318
rect -3320 -10370 -1166 -10344
rect -3320 -10416 -3295 -10370
rect -3249 -10416 -3197 -10370
rect -3151 -10416 -3099 -10370
rect -3053 -10416 -3001 -10370
rect -2955 -10416 -2903 -10370
rect -2857 -10416 -2805 -10370
rect -2759 -10416 -2707 -10370
rect -2661 -10416 -2609 -10370
rect -2563 -10416 -2511 -10370
rect -2465 -10416 -2413 -10370
rect -2367 -10416 -2315 -10370
rect -2269 -10416 -2217 -10370
rect -2171 -10416 -2119 -10370
rect -2073 -10416 -2021 -10370
rect -1975 -10416 -1923 -10370
rect -1877 -10416 -1825 -10370
rect -1779 -10416 -1727 -10370
rect -1681 -10416 -1629 -10370
rect -1583 -10416 -1531 -10370
rect -1485 -10416 -1433 -10370
rect -1387 -10416 -1335 -10370
rect -1289 -10416 -1237 -10370
rect -1191 -10416 -1166 -10370
rect -3320 -10441 -1166 -10416
rect -574 -10334 -477 -10313
rect -574 -10380 -549 -10334
rect -503 -10380 -477 -10334
rect -324 -10321 -278 -10237
rect -164 -10321 -118 -10254
rect -324 -10367 -246 -10321
rect -200 -10367 -118 -10321
rect -574 -10432 -477 -10380
rect -574 -10478 -549 -10432
rect -503 -10478 -477 -10432
rect -574 -10530 -477 -10478
rect -164 -10481 -118 -10367
rect -4 -10369 42 -10260
rect 444 -10364 546 -10351
rect 444 -10369 460 -10364
rect -4 -10415 460 -10369
rect 444 -10420 460 -10415
rect 532 -10369 546 -10364
rect 638 -10369 684 -10260
rect 532 -10415 684 -10369
rect 798 -10328 844 -10260
rect 958 -10318 1004 -10259
rect 1190 -10282 1215 -10236
rect 1261 -10282 1287 -10236
rect 944 -10328 1011 -10318
rect 798 -10329 1011 -10328
rect 798 -10375 957 -10329
rect 1003 -10375 1011 -10329
rect 798 -10376 1011 -10375
rect 532 -10420 546 -10415
rect 444 -10434 546 -10420
rect 798 -10481 844 -10376
rect 944 -10388 1011 -10376
rect 1190 -10334 1287 -10282
rect 1190 -10380 1215 -10334
rect 1261 -10380 1287 -10334
rect -164 -10527 844 -10481
rect 1190 -10432 1287 -10380
rect 1190 -10478 1215 -10432
rect 1261 -10478 1287 -10432
rect -574 -10576 -549 -10530
rect -503 -10576 -477 -10530
rect -574 -10602 -477 -10576
rect 1190 -10530 1287 -10478
rect 1190 -10576 1215 -10530
rect 1261 -10576 1287 -10530
rect 1190 -10602 1287 -10576
rect -574 -10628 1287 -10602
rect -574 -10674 -549 -10628
rect -503 -10674 -451 -10628
rect -405 -10674 -353 -10628
rect -307 -10674 -255 -10628
rect -209 -10674 -157 -10628
rect -111 -10674 -59 -10628
rect -13 -10674 39 -10628
rect 85 -10674 137 -10628
rect 183 -10674 235 -10628
rect 281 -10674 333 -10628
rect 379 -10674 431 -10628
rect 477 -10674 529 -10628
rect 575 -10674 627 -10628
rect 673 -10674 725 -10628
rect 771 -10674 823 -10628
rect 869 -10674 921 -10628
rect 967 -10674 1019 -10628
rect 1065 -10674 1117 -10628
rect 1163 -10674 1215 -10628
rect 1261 -10674 1287 -10628
rect -574 -10699 1287 -10674
<< via1 >>
rect 432 1601 561 1708
rect -2758 -1828 -2704 -1774
rect -2402 1229 -2342 1289
rect -2326 -1828 -2272 -1774
rect 196 1383 258 1441
rect 1571 1360 1681 1465
rect -229 1175 -171 1231
rect 631 1172 691 1229
rect 1365 1153 1474 1257
rect -230 792 -172 848
rect 199 789 259 847
rect 632 794 692 851
rect -242 -145 -160 -66
rect 621 -150 703 -71
rect -1894 -1831 -1840 -1777
rect -3452 -2262 -3396 -2206
rect -3341 -2262 -3285 -2206
rect -2759 -2268 -2703 -2212
rect -2327 -2264 -2271 -2208
rect -1895 -2272 -1839 -2216
rect -3453 -2372 -3397 -2316
rect -3342 -2372 -3286 -2316
rect -313 -2223 -260 -2170
rect -205 -2221 -153 -2169
rect 283 -1181 341 -1117
rect 195 -2219 247 -2167
rect -233 -3185 -172 -3126
rect 200 -3188 261 -3129
rect 632 -3185 693 -3126
rect -233 -3573 -171 -3513
rect 634 -3577 695 -3516
rect 1364 -3601 1473 -3497
rect 198 -3773 260 -3710
rect 1565 -3798 1675 -3693
rect -164 -4248 -83 -4238
rect -164 -4303 -154 -4248
rect -154 -4303 -90 -4248
rect -90 -4303 -83 -4248
rect -164 -4310 -83 -4303
rect 200 -4284 255 -4229
rect 368 -4404 422 -4350
rect 367 -6004 423 -5948
rect 63 -6117 119 -6061
rect 4363 -6282 4434 -6215
rect -3053 -7283 -2997 -7227
rect -2893 -7285 -2837 -7229
rect -3052 -8085 -2996 -8029
rect -2893 -8086 -2837 -8030
rect -3055 -8887 -2999 -8831
rect -2893 -8887 -2837 -8831
rect -3055 -9686 -2999 -9630
rect -2893 -9688 -2837 -9632
rect -2573 -7598 -2517 -7542
rect -2573 -8399 -2517 -8343
rect -2573 -9200 -2517 -9144
rect -2573 -10001 -2517 -9945
rect -2254 -7285 -2198 -7229
rect -2256 -7815 -2196 -7809
rect -2256 -7864 -2251 -7815
rect -2251 -7864 -2202 -7815
rect -2202 -7864 -2196 -7815
rect -2256 -7869 -2196 -7864
rect -2254 -8086 -2198 -8030
rect -2256 -8616 -2196 -8610
rect -2256 -8665 -2251 -8616
rect -2251 -8665 -2202 -8616
rect -2202 -8665 -2196 -8616
rect -2256 -8670 -2196 -8665
rect -2254 -8887 -2198 -8831
rect -2257 -9416 -2197 -9410
rect -2257 -9465 -2252 -9416
rect -2252 -9465 -2203 -9416
rect -2203 -9465 -2197 -9416
rect -2257 -9470 -2197 -9465
rect -2254 -9688 -2198 -9632
rect -1935 -7599 -1879 -7543
rect -1935 -8400 -1879 -8344
rect -1935 -9201 -1879 -9145
rect -1935 -10002 -1879 -9946
rect 143 -6880 215 -6824
rect 3691 -6709 3759 -6551
rect -1615 -7284 -1559 -7228
rect -1457 -7286 -1401 -7230
rect -169 -7129 -113 -7047
rect 2349 -7089 2506 -6920
rect 312 -7287 368 -7215
rect -1615 -8085 -1559 -8029
rect -1456 -8086 -1400 -8030
rect -169 -8367 -113 -8295
rect -1615 -8886 -1559 -8830
rect -1454 -8886 -1398 -8830
rect -1615 -9687 -1559 -9631
rect -1455 -9686 -1399 -9630
rect 309 -7682 375 -7677
rect 309 -7740 313 -7682
rect 313 -7740 371 -7682
rect 371 -7740 375 -7682
rect 309 -7743 375 -7740
rect 3274 -7296 3352 -7218
rect 3934 -7265 4001 -7197
rect 153 -7985 209 -7913
rect 305 -8136 377 -8080
rect 148 -8577 204 -8505
rect 474 -8576 530 -8504
rect -9 -8733 47 -8661
rect 304 -9154 376 -9098
rect 5000 -7333 5089 -7250
rect 1396 -7696 1469 -7622
rect 3016 -7696 3095 -7618
rect 793 -8372 849 -8300
rect 634 -8733 690 -8661
rect 471 -9300 527 -9228
rect 300 -9511 366 -9506
rect 300 -9569 304 -9511
rect 304 -9569 362 -9511
rect 362 -9569 366 -9511
rect 300 -9572 366 -9569
rect 904 -8593 970 -8588
rect 904 -8651 908 -8593
rect 908 -8651 966 -8593
rect 966 -8651 970 -8593
rect 904 -8654 970 -8651
rect 313 -9907 369 -9835
rect -169 -10118 -113 -10036
rect 460 -10420 532 -10364
<< metal2 >>
rect 406 1708 587 1736
rect 406 1692 432 1708
rect -986 1610 432 1692
rect -986 1442 -904 1610
rect 406 1601 432 1610
rect 561 1692 587 1708
rect 2339 1692 2460 1712
rect 561 1610 2460 1692
rect 561 1601 587 1610
rect 406 1576 587 1601
rect 1558 1465 1693 1479
rect -2407 1360 -576 1442
rect 184 1441 266 1451
rect 184 1383 196 1441
rect 258 1383 266 1441
rect 184 1372 266 1383
rect -2407 1320 -2312 1360
rect -2431 1289 -2312 1320
rect -2431 1229 -2402 1289
rect -2342 1229 -2312 1289
rect -2431 1201 -2312 1229
rect -2773 -1774 -2689 -1764
rect -2773 -1828 -2758 -1774
rect -2704 -1828 -2689 -1774
rect -2773 -1842 -2689 -1828
rect -2343 -1774 -2259 -1764
rect -2343 -1828 -2326 -1774
rect -2272 -1828 -2259 -1774
rect -2343 -1842 -2259 -1828
rect -1909 -1777 -1825 -1766
rect -1909 -1831 -1894 -1777
rect -1840 -1831 -1825 -1777
rect -3472 -2206 -3250 -2187
rect -3472 -2262 -3452 -2206
rect -3396 -2262 -3341 -2206
rect -3285 -2262 -3250 -2206
rect -2759 -2207 -2703 -1842
rect -2327 -2201 -2271 -1842
rect -1909 -1844 -1825 -1831
rect -3472 -2316 -3250 -2262
rect -2773 -2212 -2689 -2207
rect -2773 -2268 -2759 -2212
rect -2703 -2268 -2689 -2212
rect -2773 -2285 -2689 -2268
rect -2341 -2208 -2257 -2201
rect -1895 -2208 -1839 -1844
rect -658 -2154 -576 1360
rect -240 1231 -158 1244
rect -240 1175 -229 1231
rect -171 1175 -158 1231
rect -240 1164 -158 1175
rect -229 860 -172 1164
rect 199 860 256 1372
rect 1558 1360 1571 1465
rect 1681 1360 1693 1465
rect 1558 1344 1693 1360
rect 1352 1257 1487 1272
rect 618 1229 702 1245
rect 618 1172 631 1229
rect 691 1172 702 1229
rect 618 1161 702 1172
rect 632 866 690 1161
rect 1352 1153 1365 1257
rect 1474 1153 1487 1257
rect 1352 1137 1487 1153
rect -242 848 -160 860
rect -242 792 -230 848
rect -172 792 -160 848
rect -242 780 -160 792
rect 184 847 272 860
rect 184 789 199 847
rect 259 789 272 847
rect 184 776 272 789
rect 618 851 702 866
rect 618 794 632 851
rect 692 794 702 851
rect 618 782 702 794
rect -260 -66 -144 -44
rect -260 -145 -242 -66
rect -160 -145 -144 -66
rect -260 -160 -144 -145
rect 605 -71 721 -51
rect 605 -150 621 -71
rect 703 -150 721 -71
rect 605 -167 721 -150
rect 1363 -1108 1474 1137
rect 272 -1117 351 -1108
rect 272 -1181 283 -1117
rect 341 -1181 351 -1117
rect 272 -1191 351 -1181
rect 1363 -1186 1377 -1108
rect 1461 -1186 1474 -1108
rect -658 -2167 259 -2154
rect -658 -2169 195 -2167
rect -658 -2170 -205 -2169
rect -2341 -2264 -2327 -2208
rect -2271 -2264 -2257 -2208
rect -2341 -2279 -2257 -2264
rect -1909 -2216 -1825 -2208
rect -1909 -2272 -1895 -2216
rect -1839 -2272 -1825 -2216
rect -658 -2223 -313 -2170
rect -260 -2221 -205 -2170
rect -153 -2219 195 -2169
rect 247 -2219 259 -2167
rect -153 -2221 259 -2219
rect -260 -2223 259 -2221
rect -658 -2236 259 -2223
rect -1909 -2286 -1825 -2272
rect -3472 -2372 -3453 -2316
rect -3397 -2372 -3342 -2316
rect -3286 -2372 -3250 -2316
rect -3472 -2404 -3250 -2372
rect -3668 -2505 -3546 -2473
rect -3668 -2569 -3639 -2505
rect -3575 -2569 -3546 -2505
rect -3668 -2597 -3546 -2569
rect -3664 -2739 -3542 -2707
rect -3664 -2803 -3635 -2739
rect -3571 -2803 -3542 -2739
rect -3664 -2831 -3542 -2803
rect -3472 -3116 -3352 -2404
rect -1743 -2744 -1642 -2723
rect -1743 -2800 -1722 -2744
rect -1666 -2800 -1642 -2744
rect -1743 -2820 -1642 -2800
rect -2607 -2965 -2524 -2953
rect -2156 -2965 -1882 -2952
rect -2607 -2967 -2142 -2965
rect -2607 -3023 -2593 -2967
rect -2537 -3021 -2142 -2967
rect -2086 -3021 -2032 -2965
rect -1976 -2967 -1882 -2965
rect -1976 -3021 -1952 -2967
rect -2537 -3023 -1952 -3021
rect -1896 -3023 -1882 -2967
rect -2607 -3025 -1882 -3023
rect -2607 -3035 -2524 -3025
rect -2156 -3036 -1882 -3025
rect -2766 -3116 -2683 -3105
rect -2447 -3116 -2364 -3104
rect -2125 -3116 -2042 -3104
rect -1810 -3116 -1727 -3104
rect -3472 -3118 -1727 -3116
rect -3472 -3119 -2433 -3118
rect -3472 -3175 -2752 -3119
rect -2696 -3174 -2433 -3119
rect -2377 -3174 -2111 -3118
rect -2055 -3174 -1796 -3118
rect -1740 -3174 -1727 -3118
rect -2696 -3175 -1727 -3174
rect -3472 -3177 -1727 -3175
rect -3472 -3973 -3352 -3177
rect -2766 -3187 -2683 -3177
rect -2447 -3186 -2364 -3177
rect -2125 -3186 -2042 -3177
rect -1810 -3186 -1727 -3177
rect -245 -3126 -160 -3114
rect -245 -3185 -233 -3126
rect -172 -3185 -160 -3126
rect -245 -3198 -160 -3185
rect 188 -3129 273 -3117
rect 188 -3188 200 -3129
rect 261 -3188 273 -3129
rect -3088 -3272 -3004 -3260
rect -2927 -3272 -2843 -3259
rect -2547 -3272 -2355 -3260
rect -2288 -3272 -2202 -3260
rect -1647 -3272 -1563 -3259
rect -1487 -3272 -1403 -3260
rect -3088 -3273 -1403 -3272
rect -3088 -3274 -2533 -3273
rect -3088 -3330 -3074 -3274
rect -3018 -3330 -2913 -3274
rect -2857 -3329 -2533 -3274
rect -2477 -3329 -2423 -3273
rect -2367 -3274 -1403 -3273
rect -2367 -3329 -2274 -3274
rect -2857 -3330 -2274 -3329
rect -2216 -3330 -1633 -3274
rect -1577 -3330 -1473 -3274
rect -1417 -3330 -1403 -3274
rect -3088 -3332 -1403 -3330
rect -3088 -3344 -3004 -3332
rect -2927 -3343 -2843 -3332
rect -2547 -3344 -2355 -3332
rect -2288 -3344 -2202 -3332
rect -1647 -3343 -1563 -3332
rect -1487 -3344 -1403 -3332
rect -238 -3507 -168 -3198
rect 188 -3201 273 -3188
rect 620 -3126 705 -3112
rect 620 -3185 632 -3126
rect 693 -3185 705 -3126
rect 620 -3198 705 -3185
rect 194 -3202 265 -3201
rect -244 -3513 -162 -3507
rect -2852 -3561 -2751 -3540
rect -2852 -3617 -2831 -3561
rect -2775 -3617 -2751 -3561
rect -244 -3573 -233 -3513
rect -171 -3573 -162 -3513
rect -244 -3582 -162 -3573
rect -2852 -3637 -2751 -3617
rect 194 -3699 264 -3202
rect 634 -3453 693 -3198
rect 633 -3504 694 -3453
rect 1363 -3482 1474 -1186
rect 1567 -71 1681 1344
rect 1567 -149 1583 -71
rect 1666 -149 1681 -71
rect 1352 -3497 1486 -3482
rect 620 -3516 707 -3504
rect 620 -3577 634 -3516
rect 695 -3577 707 -3516
rect 620 -3590 707 -3577
rect 185 -3710 274 -3699
rect 185 -3773 198 -3710
rect 260 -3773 274 -3710
rect 185 -3788 274 -3773
rect -2524 -3808 -2332 -3806
rect -2607 -3819 -2332 -3808
rect -2607 -3822 -2510 -3819
rect -2607 -3878 -2593 -3822
rect -2537 -3875 -2510 -3822
rect -2454 -3875 -2400 -3819
rect -2344 -3820 -2332 -3819
rect -1965 -3820 -1882 -3809
rect -2344 -3822 -1882 -3820
rect -2344 -3875 -1952 -3822
rect -2537 -3878 -1952 -3875
rect -1896 -3878 -1882 -3822
rect -2607 -3880 -1882 -3878
rect -2607 -3890 -2332 -3880
rect -1965 -3891 -1882 -3880
rect -2767 -3973 -2684 -3961
rect -2446 -3971 -2363 -3960
rect -2446 -3973 -2435 -3971
rect -3472 -3975 -2435 -3973
rect -3472 -4031 -2753 -3975
rect -2697 -4031 -2435 -3975
rect -3472 -4033 -2435 -4031
rect -2373 -3973 -2363 -3971
rect -2126 -3973 -2043 -3960
rect -1806 -3973 -1723 -3961
rect -2373 -3974 -1723 -3973
rect -2373 -4030 -2112 -3974
rect -2056 -3975 -1723 -3974
rect -2056 -4030 -1792 -3975
rect -2373 -4031 -1792 -4030
rect -1736 -4031 -1723 -3975
rect -2373 -4033 -1723 -4031
rect -3472 -4034 -1723 -4033
rect -3472 -4837 -3352 -4034
rect -2767 -4043 -2684 -4034
rect -2446 -4042 -2363 -4034
rect -2126 -4042 -2043 -4034
rect -1806 -4043 -1723 -4034
rect -3088 -4132 -3004 -4120
rect -2927 -4132 -2843 -4119
rect -2288 -4132 -2202 -4120
rect -2121 -4131 -1929 -4118
rect -2121 -4132 -2107 -4131
rect -3088 -4134 -2107 -4132
rect -3088 -4190 -3074 -4134
rect -3018 -4190 -2913 -4134
rect -2857 -4190 -2274 -4134
rect -2216 -4187 -2107 -4134
rect -2051 -4187 -1997 -4131
rect -1941 -4132 -1929 -4131
rect -1647 -4132 -1563 -4119
rect -1487 -4132 -1403 -4120
rect -1941 -4134 -1403 -4132
rect -1941 -4187 -1633 -4134
rect -2216 -4190 -1633 -4187
rect -1577 -4190 -1473 -4134
rect -1417 -4190 -1403 -4134
rect -3088 -4192 -1403 -4190
rect -3088 -4204 -3004 -4192
rect -2927 -4203 -2843 -4192
rect -2288 -4204 -2202 -4192
rect -2121 -4202 -1929 -4192
rect -1647 -4203 -1563 -4192
rect -1487 -4204 -1403 -4192
rect 194 -4215 264 -3788
rect -176 -4238 -66 -4223
rect -176 -4310 -164 -4238
rect -83 -4310 -66 -4238
rect 187 -4229 267 -4215
rect 187 -4284 200 -4229
rect 255 -4284 267 -4229
rect 187 -4299 267 -4284
rect -176 -4325 -66 -4310
rect -1745 -4404 -1644 -4386
rect -1745 -4465 -1726 -4404
rect -1664 -4465 -1644 -4404
rect -1745 -4483 -1644 -4465
rect -2524 -4668 -2332 -4666
rect -2607 -4679 -2332 -4668
rect -2607 -4682 -2510 -4679
rect -2607 -4738 -2593 -4682
rect -2537 -4735 -2510 -4682
rect -2454 -4735 -2400 -4679
rect -2344 -4680 -2332 -4679
rect -1965 -4680 -1882 -4669
rect -2344 -4682 -1882 -4680
rect -2344 -4735 -1952 -4682
rect -2537 -4738 -1952 -4735
rect -1896 -4738 -1882 -4682
rect -2607 -4740 -1882 -4738
rect -2607 -4750 -2332 -4740
rect -1965 -4751 -1882 -4740
rect -158 -4696 -82 -4325
rect 633 -4337 694 -3590
rect 1352 -3601 1364 -3497
rect 1473 -3601 1486 -3497
rect 1352 -3616 1486 -3601
rect 1567 -3679 1681 -149
rect 1552 -3693 1687 -3679
rect 1552 -3798 1565 -3693
rect 1675 -3798 1687 -3693
rect 1552 -3814 1687 -3798
rect 356 -4350 694 -4337
rect 356 -4404 368 -4350
rect 422 -4398 694 -4350
rect 422 -4404 433 -4398
rect 356 -4414 433 -4404
rect -158 -4772 1952 -4696
rect -2767 -4837 -2684 -4825
rect -2447 -4837 -2364 -4826
rect -2127 -4837 -2044 -4824
rect -1807 -4837 -1724 -4825
rect -3472 -4838 -1724 -4837
rect -3472 -4839 -2113 -4838
rect -3472 -4895 -2753 -4839
rect -2697 -4840 -2113 -4839
rect -2697 -4895 -2433 -4840
rect -3472 -4896 -2433 -4895
rect -2377 -4894 -2113 -4840
rect -2057 -4839 -1724 -4838
rect -2057 -4894 -1793 -4839
rect -2377 -4895 -1793 -4894
rect -1737 -4895 -1724 -4839
rect -2377 -4896 -1724 -4895
rect -3472 -4898 -1724 -4896
rect -3472 -5691 -3352 -4898
rect -2767 -4907 -2684 -4898
rect -2447 -4908 -2364 -4898
rect -2127 -4906 -2044 -4898
rect -1807 -4907 -1724 -4898
rect -3088 -4986 -3004 -4975
rect -3088 -5048 -3077 -4986
rect -3015 -4987 -3004 -4986
rect -2927 -4985 -2843 -4974
rect -2927 -4987 -2916 -4985
rect -3015 -5047 -2916 -4987
rect -2854 -4987 -2843 -4985
rect -2288 -4986 -2202 -4975
rect -2288 -4987 -2276 -4986
rect -2854 -5047 -2276 -4987
rect -3015 -5048 -3004 -5047
rect -3088 -5059 -3004 -5048
rect -2927 -5058 -2843 -5047
rect -2288 -5048 -2276 -5047
rect -2214 -4987 -2202 -4986
rect -2120 -4987 -1928 -4976
rect -1647 -4986 -1563 -4974
rect -1647 -4987 -1636 -4986
rect -2214 -4989 -1636 -4987
rect -2214 -5045 -2106 -4989
rect -2050 -5045 -1996 -4989
rect -1940 -5045 -1636 -4989
rect -2214 -5047 -1636 -5045
rect -2214 -5048 -2202 -5047
rect -2288 -5059 -2202 -5048
rect -2120 -5060 -1928 -5047
rect -1647 -5048 -1636 -5047
rect -1574 -4987 -1563 -4986
rect -1487 -4986 -1403 -4975
rect -1487 -4987 -1476 -4986
rect -1574 -5047 -1476 -4987
rect -1574 -5048 -1563 -5047
rect -1647 -5058 -1563 -5048
rect -1487 -5048 -1476 -5047
rect -1414 -5048 -1403 -4986
rect -1487 -5059 -1403 -5048
rect -2851 -5266 -2750 -5245
rect -2851 -5322 -2830 -5266
rect -2774 -5322 -2750 -5266
rect -2851 -5342 -2750 -5322
rect -2607 -5540 -2524 -5528
rect -2155 -5540 -1882 -5527
rect -2607 -5542 -2141 -5540
rect -2607 -5598 -2593 -5542
rect -2537 -5596 -2141 -5542
rect -2085 -5596 -2031 -5540
rect -1975 -5542 -1882 -5540
rect -1975 -5596 -1952 -5542
rect -2537 -5598 -1952 -5596
rect -1896 -5598 -1882 -5542
rect -2607 -5600 -1882 -5598
rect -2607 -5610 -2524 -5600
rect -2155 -5611 -1882 -5600
rect -2769 -5691 -2686 -5680
rect -2447 -5691 -2364 -5679
rect -2129 -5691 -2046 -5679
rect -1806 -5691 -1723 -5679
rect -3472 -5693 -1723 -5691
rect -3472 -5694 -2433 -5693
rect -3472 -5750 -2755 -5694
rect -2699 -5749 -2433 -5694
rect -2377 -5749 -2115 -5693
rect -2059 -5749 -1792 -5693
rect -1736 -5749 -1723 -5693
rect -2699 -5750 -1723 -5749
rect -3472 -5752 -1723 -5750
rect -3472 -5826 -3352 -5752
rect -2769 -5762 -2686 -5752
rect -2447 -5761 -2364 -5752
rect -2129 -5761 -2046 -5752
rect -1806 -5761 -1723 -5752
rect -3088 -5847 -3004 -5835
rect -2927 -5847 -2843 -5834
rect -2540 -5847 -2348 -5835
rect -2288 -5847 -2202 -5835
rect -1647 -5847 -1563 -5834
rect -1487 -5847 -1403 -5835
rect -3088 -5848 -1403 -5847
rect -3088 -5849 -2526 -5848
rect -3088 -5905 -3074 -5849
rect -3018 -5905 -2913 -5849
rect -2857 -5904 -2526 -5849
rect -2470 -5904 -2416 -5848
rect -2360 -5849 -1403 -5848
rect -2360 -5904 -2274 -5849
rect -2857 -5905 -2274 -5904
rect -2216 -5905 -1633 -5849
rect -1577 -5905 -1473 -5849
rect -1417 -5905 -1403 -5849
rect -3088 -5907 -1403 -5905
rect -3088 -5919 -3004 -5907
rect -2927 -5918 -2843 -5907
rect -2540 -5919 -2348 -5907
rect -2288 -5919 -2202 -5907
rect -1647 -5918 -1563 -5907
rect -1487 -5919 -1403 -5907
rect 342 -5942 446 -5928
rect 342 -6014 356 -5942
rect 428 -6014 446 -5942
rect 342 -6027 446 -6014
rect 38 -6054 142 -6041
rect -1742 -6087 -1641 -6066
rect -1742 -6143 -1721 -6087
rect -1665 -6143 -1641 -6087
rect 38 -6126 55 -6054
rect 127 -6126 142 -6054
rect 38 -6140 142 -6126
rect -1742 -6163 -1641 -6143
rect -2286 -6657 -2167 -6644
rect -2286 -6738 -2267 -6657
rect -2186 -6670 -2167 -6657
rect -424 -6663 -329 -6651
rect -424 -6670 -411 -6663
rect -2186 -6733 -411 -6670
rect -341 -6670 -329 -6663
rect -341 -6733 372 -6670
rect -2186 -6734 372 -6733
rect -2186 -6738 -2167 -6734
rect -2286 -6749 -2167 -6738
rect -424 -6745 -329 -6734
rect 127 -6824 229 -6811
rect 127 -6880 143 -6824
rect 215 -6880 229 -6824
rect 127 -6894 229 -6880
rect -184 -7047 -99 -7032
rect -184 -7129 -169 -7047
rect -113 -7129 -99 -7047
rect -184 -7142 -99 -7129
rect -3067 -7225 -2984 -7214
rect -2907 -7225 -2824 -7216
rect -2590 -7223 -2505 -7210
rect -2590 -7225 -2577 -7223
rect -3067 -7227 -2577 -7225
rect -3067 -7283 -3053 -7227
rect -2997 -7229 -2577 -7227
rect -2997 -7283 -2893 -7229
rect -3067 -7285 -2893 -7283
rect -2837 -7285 -2577 -7229
rect -3067 -7289 -2577 -7285
rect -3067 -7296 -2984 -7289
rect -2907 -7298 -2824 -7289
rect -2590 -7290 -2577 -7289
rect -2516 -7225 -2505 -7223
rect -2268 -7225 -2185 -7216
rect -1629 -7225 -1546 -7215
rect -1471 -7225 -1388 -7217
rect -2516 -7228 -1388 -7225
rect -2516 -7229 -1615 -7228
rect -2516 -7285 -2254 -7229
rect -2198 -7284 -1615 -7229
rect -1559 -7230 -1388 -7228
rect -1559 -7284 -1457 -7230
rect -2198 -7285 -1457 -7284
rect -2516 -7286 -1457 -7285
rect -1401 -7286 -1388 -7230
rect -2516 -7289 -1388 -7286
rect -2516 -7290 -2505 -7289
rect -2590 -7301 -2505 -7290
rect -2268 -7298 -2185 -7289
rect -1629 -7297 -1546 -7289
rect -1471 -7299 -1388 -7289
rect -2587 -7538 -2504 -7529
rect -1953 -7538 -1863 -7523
rect -2587 -7539 -732 -7538
rect -2587 -7542 -1939 -7539
rect -2587 -7598 -2573 -7542
rect -2517 -7598 -1939 -7542
rect -2587 -7602 -1939 -7598
rect -2587 -7611 -2504 -7602
rect -1953 -7608 -1939 -7602
rect -1875 -7602 -732 -7539
rect -1875 -7608 -1863 -7602
rect -1953 -7615 -1863 -7608
rect -2268 -7809 -2184 -7797
rect -2268 -7869 -2256 -7809
rect -2196 -7869 -2184 -7809
rect -2268 -7881 -2184 -7869
rect -3066 -8026 -2983 -8016
rect -2907 -8026 -2824 -8017
rect -2268 -8026 -2185 -8017
rect -1954 -8024 -1864 -8012
rect -1954 -8026 -1940 -8024
rect -3066 -8029 -1940 -8026
rect -3066 -8085 -3052 -8029
rect -2996 -8030 -1940 -8029
rect -2996 -8085 -2893 -8030
rect -3066 -8086 -2893 -8085
rect -2837 -8086 -2254 -8030
rect -2198 -8086 -1940 -8030
rect -3066 -8090 -1940 -8086
rect -3066 -8098 -2983 -8090
rect -2907 -8099 -2824 -8090
rect -2268 -8099 -2185 -8090
rect -1954 -8093 -1940 -8090
rect -1876 -8026 -1864 -8024
rect -1629 -8026 -1546 -8016
rect -1470 -8026 -1387 -8017
rect -1876 -8029 -1387 -8026
rect -1876 -8085 -1615 -8029
rect -1559 -8030 -1387 -8029
rect -1559 -8085 -1456 -8030
rect -1876 -8086 -1456 -8085
rect -1400 -8086 -1387 -8030
rect -1876 -8090 -1387 -8086
rect -1876 -8093 -1864 -8090
rect -1954 -8104 -1864 -8093
rect -1629 -8098 -1546 -8090
rect -1470 -8099 -1387 -8090
rect -2589 -8337 -2504 -8325
rect -2589 -8405 -2576 -8337
rect -2515 -8339 -2504 -8337
rect -1949 -8339 -1866 -8331
rect -2515 -8344 -962 -8339
rect -2515 -8400 -1935 -8344
rect -1879 -8400 -962 -8344
rect -2515 -8402 -962 -8400
rect -2515 -8403 -1866 -8402
rect -2515 -8405 -2504 -8403
rect -2589 -8416 -2504 -8405
rect -1949 -8413 -1866 -8403
rect -2268 -8610 -2184 -8598
rect -2268 -8670 -2256 -8610
rect -2196 -8670 -2184 -8610
rect -2268 -8682 -2184 -8670
rect -1025 -8664 -962 -8402
rect -796 -8506 -732 -7602
rect 148 -7897 211 -6894
rect 308 -7199 372 -6734
rect 298 -7215 381 -7199
rect 298 -7287 312 -7215
rect 368 -7287 381 -7215
rect 298 -7301 381 -7287
rect 1876 -7407 1952 -4772
rect 2339 -6869 2460 1610
rect 4326 -6196 4456 -6187
rect 3924 -6215 4456 -6196
rect 3924 -6282 4363 -6215
rect 4434 -6282 4456 -6215
rect 3924 -6295 4456 -6282
rect 3675 -6551 3777 -6530
rect 3675 -6577 3691 -6551
rect 3268 -6680 3691 -6577
rect 2301 -6920 2561 -6869
rect 2301 -7089 2349 -6920
rect 2506 -7089 2561 -6920
rect 2301 -7126 2561 -7089
rect 3268 -7198 3357 -6680
rect 3675 -6709 3691 -6680
rect 3759 -6709 3777 -6551
rect 3675 -6724 3777 -6709
rect 3924 -7182 4011 -6295
rect 4326 -6307 4456 -6295
rect 3914 -7197 4022 -7182
rect 3262 -7218 3366 -7198
rect 3262 -7296 3274 -7218
rect 3352 -7296 3366 -7218
rect 3914 -7265 3934 -7197
rect 4001 -7265 4022 -7197
rect 3914 -7280 4022 -7265
rect 4979 -7250 5123 -7222
rect 3262 -7310 3366 -7296
rect 4979 -7333 5000 -7250
rect 5089 -7333 5123 -7250
rect 4979 -7407 5123 -7333
rect 1876 -7483 5123 -7407
rect 1372 -7606 1494 -7595
rect 3001 -7606 3109 -7598
rect 1372 -7618 3109 -7606
rect 1372 -7622 3016 -7618
rect 297 -7677 387 -7665
rect 297 -7743 309 -7677
rect 375 -7743 387 -7677
rect 1372 -7696 1396 -7622
rect 1469 -7696 3016 -7622
rect 3095 -7696 3109 -7618
rect 1372 -7704 3109 -7696
rect 1372 -7719 1494 -7704
rect 3001 -7712 3109 -7704
rect 297 -7755 387 -7743
rect 139 -7913 222 -7897
rect 139 -7985 153 -7913
rect 209 -7985 222 -7913
rect 139 -7999 222 -7985
rect -188 -8074 -93 -8062
rect -188 -8144 -175 -8074
rect -105 -8079 -93 -8074
rect 289 -8079 391 -8067
rect -105 -8080 391 -8079
rect -105 -8136 305 -8080
rect 377 -8136 391 -8080
rect -105 -8140 391 -8136
rect -105 -8144 -93 -8140
rect -188 -8156 -93 -8144
rect 289 -8150 391 -8140
rect -422 -8293 -327 -8283
rect -183 -8293 -100 -8279
rect -422 -8295 -100 -8293
rect -422 -8365 -409 -8295
rect -339 -8365 -169 -8295
rect -422 -8367 -169 -8365
rect -113 -8299 -100 -8295
rect 779 -8299 862 -8284
rect -113 -8300 862 -8299
rect -113 -8367 793 -8300
rect -422 -8368 793 -8367
rect -422 -8377 -327 -8368
rect -183 -8370 793 -8368
rect -183 -8381 -100 -8370
rect 779 -8372 793 -8370
rect 849 -8372 862 -8300
rect 779 -8386 862 -8372
rect 134 -8505 217 -8489
rect 134 -8506 148 -8505
rect -796 -8572 148 -8506
rect 134 -8577 148 -8572
rect 204 -8506 217 -8505
rect 460 -8504 543 -8488
rect 460 -8506 474 -8504
rect 204 -8572 474 -8506
rect 204 -8577 217 -8572
rect 134 -8591 217 -8577
rect 460 -8576 474 -8572
rect 530 -8576 543 -8504
rect 460 -8590 543 -8576
rect 892 -8588 982 -8576
rect -23 -8661 60 -8645
rect -23 -8664 -9 -8661
rect -1025 -8729 -9 -8664
rect -23 -8733 -9 -8729
rect 47 -8664 60 -8661
rect 620 -8661 703 -8645
rect 620 -8664 634 -8661
rect 47 -8729 634 -8664
rect 47 -8733 60 -8729
rect -23 -8747 60 -8733
rect 620 -8733 634 -8729
rect 690 -8733 703 -8661
rect 892 -8654 904 -8588
rect 970 -8654 982 -8588
rect 892 -8666 982 -8654
rect 620 -8747 703 -8733
rect -3069 -8827 -2986 -8818
rect -2907 -8827 -2824 -8818
rect -2268 -8827 -2185 -8818
rect -1954 -8823 -1864 -8811
rect -1954 -8827 -1940 -8823
rect -3069 -8831 -1940 -8827
rect -3069 -8887 -3055 -8831
rect -2999 -8887 -2893 -8831
rect -2837 -8887 -2254 -8831
rect -2198 -8887 -1940 -8831
rect -3069 -8891 -1940 -8887
rect -3069 -8900 -2986 -8891
rect -2907 -8900 -2824 -8891
rect -2268 -8900 -2185 -8891
rect -1954 -8892 -1940 -8891
rect -1876 -8827 -1864 -8823
rect -1629 -8827 -1546 -8817
rect -1468 -8827 -1385 -8817
rect -1876 -8830 -1385 -8827
rect -1876 -8886 -1615 -8830
rect -1559 -8886 -1454 -8830
rect -1398 -8886 -1385 -8830
rect -1876 -8891 -1385 -8886
rect -1876 -8892 -1864 -8891
rect -1954 -8903 -1864 -8892
rect -1629 -8899 -1546 -8891
rect -1468 -8899 -1385 -8891
rect -186 -9093 -91 -9081
rect -2587 -9139 -2504 -9129
rect -2587 -9207 -2576 -9139
rect -2515 -9140 -2504 -9139
rect -1949 -9140 -1866 -9132
rect -2515 -9145 -1866 -9140
rect -2515 -9201 -1935 -9145
rect -1879 -9201 -1866 -9145
rect -186 -9163 -173 -9093
rect -103 -9096 -91 -9093
rect 288 -9096 390 -9085
rect -103 -9098 390 -9096
rect -103 -9154 304 -9098
rect 376 -9154 390 -9098
rect -103 -9157 390 -9154
rect -103 -9163 -91 -9157
rect -186 -9175 -91 -9163
rect 288 -9168 390 -9157
rect -2515 -9204 -1866 -9201
rect -2515 -9207 -2504 -9204
rect -2587 -9214 -2504 -9207
rect -1949 -9214 -1866 -9204
rect 457 -9228 540 -9212
rect 457 -9300 471 -9228
rect 527 -9300 540 -9228
rect 457 -9314 540 -9300
rect -2269 -9410 -2185 -9398
rect -2269 -9470 -2257 -9410
rect -2197 -9470 -2185 -9410
rect -2269 -9482 -2185 -9470
rect 288 -9506 378 -9494
rect 288 -9572 300 -9506
rect 366 -9572 378 -9506
rect 288 -9584 378 -9572
rect -3069 -9628 -2986 -9617
rect -2907 -9628 -2824 -9619
rect -2590 -9626 -2504 -9615
rect -2590 -9628 -2578 -9626
rect -3069 -9630 -2578 -9628
rect -3069 -9686 -3055 -9630
rect -2999 -9632 -2578 -9630
rect -2999 -9686 -2893 -9632
rect -3069 -9688 -2893 -9686
rect -2837 -9688 -2578 -9632
rect -3069 -9692 -2578 -9688
rect -3069 -9699 -2986 -9692
rect -2907 -9701 -2824 -9692
rect -2590 -9694 -2578 -9692
rect -2516 -9628 -2504 -9626
rect -2268 -9628 -2185 -9619
rect -1629 -9628 -1546 -9618
rect -1469 -9628 -1386 -9617
rect -2516 -9630 -1386 -9628
rect -2516 -9631 -1455 -9630
rect -2516 -9632 -1615 -9631
rect -2516 -9688 -2254 -9632
rect -2198 -9687 -1615 -9632
rect -1559 -9686 -1455 -9631
rect -1399 -9686 -1386 -9630
rect -1559 -9687 -1386 -9686
rect -2198 -9688 -1386 -9687
rect -2516 -9692 -1386 -9688
rect -2516 -9694 -2504 -9692
rect -2590 -9705 -2504 -9694
rect -2268 -9701 -2185 -9692
rect -1629 -9700 -1546 -9692
rect -1469 -9699 -1386 -9692
rect -425 -9834 -330 -9822
rect 299 -9834 382 -9819
rect -425 -9904 -412 -9834
rect -342 -9835 382 -9834
rect -342 -9904 313 -9835
rect -425 -9907 313 -9904
rect 369 -9907 382 -9835
rect -425 -9908 382 -9907
rect -425 -9916 -330 -9908
rect 299 -9921 382 -9908
rect -2587 -9941 -2504 -9932
rect -1955 -9941 -1865 -9927
rect -2587 -9945 -1940 -9941
rect -2587 -10001 -2573 -9945
rect -2517 -10001 -1940 -9945
rect -2587 -10005 -1940 -10001
rect -2587 -10014 -2504 -10005
rect -1955 -10010 -1940 -10005
rect -1876 -10010 -1865 -9941
rect -1955 -10019 -1865 -10010
rect -184 -10036 -99 -10021
rect -184 -10118 -169 -10036
rect -113 -10118 -99 -10036
rect -184 -10131 -99 -10118
rect 469 -10351 529 -9314
rect 444 -10364 546 -10351
rect 444 -10420 460 -10364
rect 532 -10420 546 -10364
rect 444 -10434 546 -10420
<< via2 >>
rect -242 -145 -160 -66
rect 621 -150 703 -71
rect 283 -1181 341 -1117
rect 1377 -1186 1461 -1108
rect -3639 -2569 -3575 -2505
rect -3635 -2803 -3571 -2739
rect -1722 -2800 -1666 -2744
rect -2142 -3021 -2086 -2965
rect -2032 -3021 -1976 -2965
rect -2533 -3329 -2477 -3273
rect -2423 -3329 -2367 -3273
rect -2831 -3617 -2775 -3561
rect 1583 -149 1666 -71
rect -2510 -3875 -2454 -3819
rect -2400 -3875 -2344 -3819
rect -2107 -4187 -2051 -4131
rect -1997 -4187 -1941 -4131
rect -1726 -4465 -1664 -4404
rect -2510 -4735 -2454 -4679
rect -2400 -4735 -2344 -4679
rect -2106 -5045 -2050 -4989
rect -1996 -5045 -1940 -4989
rect -2830 -5322 -2774 -5266
rect -2141 -5596 -2085 -5540
rect -2031 -5596 -1975 -5540
rect -2526 -5904 -2470 -5848
rect -2416 -5904 -2360 -5848
rect 356 -5948 428 -5942
rect 356 -6004 367 -5948
rect 367 -6004 423 -5948
rect 423 -6004 428 -5948
rect 356 -6014 428 -6004
rect -1721 -6143 -1665 -6087
rect 55 -6061 127 -6054
rect 55 -6117 63 -6061
rect 63 -6117 119 -6061
rect 119 -6117 127 -6061
rect 55 -6126 127 -6117
rect -2267 -6738 -2186 -6657
rect -411 -6733 -341 -6663
rect -169 -7129 -113 -7047
rect -2577 -7290 -2516 -7223
rect -1939 -7543 -1875 -7539
rect -1939 -7599 -1935 -7543
rect -1935 -7599 -1879 -7543
rect -1879 -7599 -1875 -7543
rect -1939 -7608 -1875 -7599
rect -2256 -7869 -2196 -7809
rect -1940 -8093 -1876 -8024
rect -2576 -8343 -2515 -8337
rect -2576 -8399 -2573 -8343
rect -2573 -8399 -2517 -8343
rect -2517 -8399 -2515 -8343
rect -2576 -8405 -2515 -8399
rect -2256 -8670 -2196 -8610
rect 309 -7743 375 -7677
rect 1396 -7696 1469 -7622
rect -175 -8144 -105 -8074
rect -409 -8365 -339 -8295
rect 904 -8654 970 -8588
rect -1940 -8892 -1876 -8823
rect -2576 -9144 -2515 -9139
rect -2576 -9200 -2573 -9144
rect -2573 -9200 -2517 -9144
rect -2517 -9200 -2515 -9144
rect -2576 -9207 -2515 -9200
rect -173 -9163 -103 -9093
rect -2257 -9470 -2197 -9410
rect 300 -9572 366 -9506
rect -2578 -9694 -2516 -9626
rect -412 -9904 -342 -9834
rect -1940 -9946 -1876 -9941
rect -1940 -10002 -1935 -9946
rect -1935 -10002 -1879 -9946
rect -1879 -10002 -1876 -9946
rect -1940 -10010 -1876 -10002
rect -169 -10118 -113 -10036
<< metal3 >>
rect -260 -65 -144 -44
rect 605 -65 721 -51
rect 1573 -65 1680 -50
rect -260 -66 1680 -65
rect -260 -145 -242 -66
rect -160 -71 1680 -66
rect -160 -145 621 -71
rect -260 -150 621 -145
rect 703 -149 1583 -71
rect 1666 -149 1680 -71
rect 703 -150 1680 -149
rect -260 -153 1680 -150
rect -260 -160 -144 -153
rect 605 -167 721 -153
rect 1573 -169 1680 -153
rect 1366 -1100 1473 -1090
rect 269 -1108 1473 -1100
rect 269 -1117 1377 -1108
rect 269 -1181 283 -1117
rect 341 -1181 1377 -1117
rect 269 -1186 1377 -1181
rect 1461 -1186 1473 -1108
rect 269 -1196 1473 -1186
rect 1366 -1206 1473 -1196
rect -3668 -2505 -3546 -2473
rect -3668 -2569 -3639 -2505
rect -3575 -2506 -3546 -2505
rect -3575 -2569 -1660 -2506
rect -3668 -2572 -1660 -2569
rect -3668 -2597 -3546 -2572
rect -3664 -2738 -3542 -2707
rect -1726 -2723 -1660 -2572
rect -3664 -2739 -2767 -2738
rect -3664 -2803 -3635 -2739
rect -3571 -2803 -2767 -2739
rect -3664 -2804 -2767 -2803
rect -3664 -2831 -3542 -2804
rect -2833 -3540 -2767 -2804
rect -1743 -2744 -1642 -2723
rect -1743 -2800 -1722 -2744
rect -1666 -2800 -1642 -2744
rect -1743 -2820 -1642 -2800
rect -2156 -2965 -1964 -2952
rect -2156 -3021 -2142 -2965
rect -2086 -3021 -2032 -2965
rect -1976 -3021 -1964 -2965
rect -2156 -3036 -1964 -3021
rect -2547 -3273 -2355 -3260
rect -2547 -3329 -2533 -3273
rect -2477 -3329 -2423 -3273
rect -2367 -3329 -2355 -3273
rect -2547 -3344 -2355 -3329
rect -2852 -3561 -2751 -3540
rect -2852 -3617 -2831 -3561
rect -2775 -3617 -2751 -3561
rect -2852 -3637 -2751 -3617
rect -2833 -5245 -2767 -3637
rect -2458 -3806 -2392 -3344
rect -2524 -3819 -2332 -3806
rect -2524 -3875 -2510 -3819
rect -2454 -3875 -2400 -3819
rect -2344 -3875 -2332 -3819
rect -2524 -3890 -2332 -3875
rect -2458 -4666 -2392 -3890
rect -2097 -4118 -2031 -3036
rect -2121 -4131 -1929 -4118
rect -2121 -4187 -2107 -4131
rect -2051 -4187 -1997 -4131
rect -1941 -4187 -1929 -4131
rect -2121 -4202 -1929 -4187
rect -2524 -4679 -2332 -4666
rect -2524 -4735 -2510 -4679
rect -2454 -4735 -2400 -4679
rect -2344 -4735 -2332 -4679
rect -2524 -4750 -2332 -4735
rect -2851 -5266 -2750 -5245
rect -2851 -5322 -2830 -5266
rect -2774 -5322 -2750 -5266
rect -2851 -5342 -2750 -5322
rect -2833 -6171 -2767 -5342
rect -2458 -5835 -2392 -4750
rect -2097 -4976 -2031 -4202
rect -1726 -4386 -1660 -2820
rect -1745 -4404 -1644 -4386
rect -1745 -4465 -1726 -4404
rect -1664 -4465 -1644 -4404
rect -1745 -4483 -1644 -4465
rect -2120 -4989 -1928 -4976
rect -2120 -5045 -2106 -4989
rect -2050 -5045 -1996 -4989
rect -1940 -5045 -1928 -4989
rect -2120 -5060 -1928 -5045
rect -2097 -5527 -2031 -5060
rect -2155 -5540 -1963 -5527
rect -2155 -5596 -2141 -5540
rect -2085 -5596 -2031 -5540
rect -1975 -5596 -1963 -5540
rect -2155 -5611 -1963 -5596
rect -2540 -5848 -2348 -5835
rect -2540 -5904 -2526 -5848
rect -2470 -5904 -2416 -5848
rect -2360 -5904 -2348 -5848
rect -2540 -5919 -2348 -5904
rect -2493 -6470 -2388 -5919
rect -2596 -6566 -2388 -6470
rect -2120 -6457 -2011 -5611
rect -1726 -6066 -1660 -4483
rect -421 -5906 438 -5816
rect -1742 -6087 -1641 -6066
rect -1742 -6143 -1721 -6087
rect -1665 -6143 -1641 -6087
rect -1742 -6163 -1641 -6143
rect -2120 -6553 -1861 -6457
rect -2596 -7223 -2500 -6566
rect -2286 -6657 -2167 -6644
rect -2286 -6738 -2267 -6657
rect -2186 -6738 -2167 -6657
rect -2286 -6749 -2167 -6738
rect -2596 -7290 -2577 -7223
rect -2516 -7290 -2500 -7223
rect -2596 -7291 -2500 -7290
rect -2590 -8337 -2504 -7291
rect -2590 -8405 -2576 -8337
rect -2515 -8405 -2504 -8337
rect -2590 -9139 -2504 -8405
rect -2590 -9207 -2576 -9139
rect -2515 -9207 -2504 -9139
rect -2590 -9626 -2504 -9207
rect -2273 -7809 -2180 -6749
rect -1957 -7539 -1861 -6553
rect -421 -6651 -331 -5906
rect 342 -5928 438 -5906
rect 342 -5942 446 -5928
rect 342 -6014 356 -5942
rect 428 -6014 446 -5942
rect 342 -6027 446 -6014
rect 38 -6053 142 -6041
rect -180 -6054 142 -6053
rect -180 -6126 55 -6054
rect 127 -6126 142 -6054
rect -180 -6129 142 -6126
rect -424 -6663 -329 -6651
rect -424 -6733 -411 -6663
rect -341 -6733 -329 -6663
rect -424 -6745 -329 -6733
rect -1957 -7608 -1939 -7539
rect -1875 -7608 -1861 -7539
rect -1957 -7611 -1861 -7608
rect -2273 -7869 -2256 -7809
rect -2196 -7869 -2180 -7809
rect -2273 -8610 -2180 -7869
rect -2273 -8670 -2256 -8610
rect -2196 -8670 -2180 -8610
rect -2273 -9410 -2180 -8670
rect -2273 -9470 -2257 -9410
rect -2197 -9470 -2180 -9410
rect -2273 -9490 -2180 -9470
rect -1951 -8024 -1865 -7611
rect -1951 -8093 -1940 -8024
rect -1876 -8093 -1865 -8024
rect -1951 -8823 -1865 -8093
rect -421 -8283 -331 -6745
rect -180 -7032 -104 -6129
rect 38 -6140 142 -6129
rect -184 -7047 -99 -7032
rect -184 -7129 -169 -7047
rect -113 -7129 -99 -7047
rect -184 -7142 -99 -7129
rect -180 -8062 -104 -7142
rect 1020 -7623 1096 -7574
rect 1372 -7622 1494 -7595
rect 1372 -7623 1396 -7622
rect 297 -7669 387 -7665
rect 1020 -7669 1396 -7623
rect 297 -7677 1396 -7669
rect 297 -7743 309 -7677
rect 375 -7696 1396 -7677
rect 1469 -7696 1494 -7622
rect 375 -7697 1494 -7696
rect 375 -7743 1096 -7697
rect 1372 -7719 1494 -7697
rect 297 -7752 1096 -7743
rect 297 -7755 387 -7752
rect -188 -8074 -93 -8062
rect -188 -8144 -175 -8074
rect -105 -8144 -93 -8074
rect -188 -8156 -93 -8144
rect -422 -8295 -327 -8283
rect -422 -8365 -409 -8295
rect -339 -8365 -327 -8295
rect -422 -8377 -327 -8365
rect -1951 -8892 -1940 -8823
rect -1876 -8892 -1865 -8823
rect -2590 -9694 -2578 -9626
rect -2516 -9694 -2504 -9626
rect -2590 -9705 -2504 -9694
rect -1951 -9941 -1865 -8892
rect -421 -9822 -331 -8377
rect -180 -9081 -104 -8156
rect 1020 -8545 1096 -7752
rect 891 -8588 1096 -8545
rect 891 -8654 904 -8588
rect 970 -8654 1096 -8588
rect 891 -8684 1096 -8654
rect -186 -9093 -91 -9081
rect -186 -9163 -173 -9093
rect -103 -9163 -91 -9093
rect -186 -9175 -91 -9163
rect -425 -9834 -330 -9822
rect -425 -9904 -412 -9834
rect -342 -9904 -330 -9834
rect -425 -9916 -330 -9904
rect -1951 -10010 -1940 -9941
rect -1876 -10010 -1865 -9941
rect -1951 -10020 -1865 -10010
rect -180 -10021 -104 -9175
rect 288 -9497 378 -9494
rect 1020 -9497 1096 -8684
rect 288 -9506 1096 -9497
rect 288 -9572 300 -9506
rect 366 -9572 1096 -9506
rect 288 -9580 1096 -9572
rect 288 -9584 378 -9580
rect 1020 -9670 1096 -9580
rect -184 -10036 -99 -10021
rect -184 -10118 -169 -10036
rect -113 -10118 -99 -10036
rect -184 -10131 -99 -10118
use nmos_3p3_77EFTS  nmos_3p3_77EFTS_0
timestamp 1692885173
transform 1 0 4317 0 1 -7735
box -168 -268 168 268
use nmos_3p3_77EFTS  nmos_3p3_77EFTS_1
timestamp 1692885173
transform 1 0 3444 0 1 -7735
box -168 -268 168 268
use nmos_3p3_77EFTS  nmos_3p3_77EFTS_2
timestamp 1692885173
transform 1 0 3888 0 1 -7736
box -168 -268 168 268
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_0
timestamp 1692712407
transform 1 0 -2546 0 -1 -9037
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_1
timestamp 1692712407
transform 1 0 -2546 0 -1 -9837
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_2
timestamp 1692712407
transform -1 0 -1906 0 -1 -9037
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_3
timestamp 1692712407
transform -1 0 -1906 0 -1 -9837
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_4
timestamp 1692712407
transform 1 0 -2546 0 1 -8239
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_5
timestamp 1692712407
transform -1 0 -1906 0 1 -8239
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_6
timestamp 1692712407
transform 1 0 -2546 0 1 -7439
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_7
timestamp 1692712407
transform -1 0 -1906 0 1 -7439
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_8
timestamp 1692712407
transform 1 0 340 0 1 -9962
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_9
timestamp 1692712407
transform 1 0 340 0 1 -9112
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_10
timestamp 1692712407
transform 1 0 340 0 1 -8132
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_11
timestamp 1692712407
transform 1 0 340 0 1 -7282
box -220 -368 220 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_0
timestamp 1692712407
transform 1 0 -2946 0 -1 -9037
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_1
timestamp 1692712407
transform 1 0 -2306 0 -1 -9037
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_2
timestamp 1692712407
transform 1 0 -2786 0 -1 -9037
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_3
timestamp 1692712407
transform 1 0 -2306 0 -1 -9837
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_4
timestamp 1692712407
transform 1 0 -2946 0 -1 -9837
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_5
timestamp 1692712407
transform 1 0 -2786 0 -1 -9837
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_6
timestamp 1692712407
transform -1 0 -2146 0 -1 -9037
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_7
timestamp 1692712407
transform -1 0 -1666 0 -1 -9037
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_8
timestamp 1692712407
transform -1 0 -1506 0 -1 -9037
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_9
timestamp 1692712407
transform -1 0 -2146 0 -1 -9837
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_10
timestamp 1692712407
transform -1 0 -1506 0 -1 -9837
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_11
timestamp 1692712407
transform -1 0 -1666 0 -1 -9837
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_12
timestamp 1692712407
transform 1 0 -2306 0 1 -8239
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_13
timestamp 1692712407
transform 1 0 -2786 0 1 -8239
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_14
timestamp 1692712407
transform 1 0 -2946 0 1 -8239
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_15
timestamp 1692712407
transform -1 0 -1506 0 1 -8239
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_16
timestamp 1692712407
transform -1 0 -1666 0 1 -8239
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_17
timestamp 1692712407
transform -1 0 -2146 0 1 -8239
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_18
timestamp 1692712407
transform 1 0 -2306 0 1 -7439
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_19
timestamp 1692712407
transform 1 0 -2946 0 1 -7439
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_20
timestamp 1692712407
transform 1 0 -2786 0 1 -7439
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_21
timestamp 1692712407
transform -1 0 -2146 0 1 -7439
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_22
timestamp 1692712407
transform -1 0 -1666 0 1 -7439
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_23
timestamp 1692712407
transform -1 0 -1506 0 1 -7439
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_24
timestamp 1692712407
transform -1 0 741 0 1 -9962
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_25
timestamp 1692712407
transform -1 0 901 0 1 -9962
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_26
timestamp 1692712407
transform -1 0 -221 0 1 -9962
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_27
timestamp 1692712407
transform -1 0 -61 0 1 -9962
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_28
timestamp 1692712407
transform -1 0 901 0 1 -9112
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_29
timestamp 1692712407
transform -1 0 741 0 1 -9112
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_30
timestamp 1692712407
transform -1 0 -221 0 1 -9112
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_31
timestamp 1692712407
transform -1 0 -61 0 1 -9112
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_32
timestamp 1692712407
transform -1 0 -61 0 1 -8132
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_33
timestamp 1692712407
transform -1 0 -221 0 1 -8132
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_34
timestamp 1692712407
transform -1 0 901 0 1 -8132
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_35
timestamp 1692712407
transform -1 0 741 0 1 -8132
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_36
timestamp 1692712407
transform -1 0 -221 0 1 -7282
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_37
timestamp 1692712407
transform -1 0 -61 0 1 -7282
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_38
timestamp 1692712407
transform -1 0 901 0 1 -7282
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_39
timestamp 1692712407
transform -1 0 741 0 1 -7282
box -140 -368 140 368
use pmos_3p3_9BLZD7  pmos_3p3_9BLZD7_0
timestamp 1692615943
transform 1 0 -2299 0 1 -255
box -554 -1534 554 1534
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_0
timestamp 1692615943
transform 1 0 771 0 1 -1664
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_1
timestamp 1692615943
transform 1 0 -309 0 1 -2702
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_2
timestamp 1692615943
transform 1 0 -93 0 1 -2702
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_3
timestamp 1692615943
transform 1 0 555 0 1 -1664
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_4
timestamp 1692615943
transform 1 0 771 0 1 -2702
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_5
timestamp 1692615943
transform 1 0 555 0 1 -2702
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_6
timestamp 1692615943
transform 1 0 -309 0 1 -1664
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_7
timestamp 1692615943
transform 1 0 -93 0 1 -1664
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_8
timestamp 1692615943
transform 1 0 771 0 1 -624
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_9
timestamp 1692615943
transform 1 0 555 0 1 -624
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_10
timestamp 1692615943
transform 1 0 555 0 1 414
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_11
timestamp 1692615943
transform 1 0 771 0 1 414
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_12
timestamp 1692615943
transform 1 0 -93 0 1 -624
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_13
timestamp 1692615943
transform 1 0 -309 0 1 -624
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_14
timestamp 1692615943
transform 1 0 -309 0 1 414
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_15
timestamp 1692615943
transform 1 0 -93 0 1 414
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_16
timestamp 1692615943
transform 1 0 -2839 0 1 -1359
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_17
timestamp 1692615943
transform 1 0 -1759 0 1 -1359
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_18
timestamp 1692615943
transform 1 0 -2839 0 1 113
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_19
timestamp 1692615943
transform 1 0 -2839 0 1 -623
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_20
timestamp 1692615943
transform 1 0 -2839 0 1 849
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_21
timestamp 1692615943
transform 1 0 -1759 0 1 849
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_22
timestamp 1692615943
transform 1 0 -1759 0 1 113
box -230 -430 230 430
use pmos_3p3_9K6RD7  pmos_3p3_9K6RD7_23
timestamp 1692615943
transform 1 0 -1759 0 1 -623
box -230 -430 230 430
use pmos_3p3_M6GBWP  pmos_3p3_M6GBWP_0
timestamp 1692885173
transform 1 0 4946 0 1 -6753
box -230 -220 230 220
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_0
timestamp 1692683681
transform 1 0 395 0 1 -5568
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_1
timestamp 1692683681
transform 1 0 395 0 1 -4788
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_2
timestamp 1692683681
transform -1 0 -1925 0 -1 -4869
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_3
timestamp 1692683681
transform -1 0 -1925 0 -1 -5721
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_4
timestamp 1692683681
transform 1 0 -2565 0 -1 -4869
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_5
timestamp 1692683681
transform 1 0 -2565 0 -1 -5721
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_6
timestamp 1692683681
transform 1 0 -2565 0 1 -4017
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_7
timestamp 1692683681
transform -1 0 -1925 0 1 -4017
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_8
timestamp 1692683681
transform 1 0 -2565 0 1 -3165
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_9
timestamp 1692683681
transform -1 0 -1925 0 1 -3165
box -282 -430 282 430
use pmos_3p3_M22VUP  pmos_3p3_M22VUP_0
timestamp 1691491496
transform 1 0 231 0 1 -1664
box -338 -430 338 430
use pmos_3p3_M22VUP  pmos_3p3_M22VUP_1
timestamp 1691491496
transform 1 0 231 0 1 -2702
box -338 -430 338 430
use pmos_3p3_M22VUP  pmos_3p3_M22VUP_2
timestamp 1691491496
transform 1 0 231 0 1 -624
box -338 -430 338 430
use pmos_3p3_M22VUP  pmos_3p3_M22VUP_3
timestamp 1691491496
transform 1 0 231 0 1 414
box -338 -430 338 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_0
timestamp 1692683681
transform 1 0 27 0 1 -5568
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_1
timestamp 1692683681
transform 1 0 -133 0 1 -5568
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_2
timestamp 1692683681
transform 1 0 923 0 1 -5568
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_3
timestamp 1692683681
transform 1 0 763 0 1 -5568
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_4
timestamp 1692683681
transform 1 0 -133 0 1 -4788
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_5
timestamp 1692683681
transform 1 0 27 0 1 -4788
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_6
timestamp 1692683681
transform 1 0 923 0 1 -4788
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_7
timestamp 1692683681
transform 1 0 763 0 1 -4788
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_8
timestamp 1692683681
transform -1 0 -1525 0 -1 -4869
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_9
timestamp 1692683681
transform -1 0 -1685 0 -1 -4869
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_10
timestamp 1692683681
transform -1 0 -2165 0 -1 -4869
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_11
timestamp 1692683681
transform -1 0 -1685 0 -1 -5721
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_12
timestamp 1692683681
transform -1 0 -1525 0 -1 -5721
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_13
timestamp 1692683681
transform -1 0 -2165 0 -1 -5721
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_14
timestamp 1692683681
transform 1 0 -2805 0 1 -4017
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_15
timestamp 1692683681
transform 1 0 -2965 0 1 -4017
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_16
timestamp 1692683681
transform 1 0 -2805 0 -1 -4869
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_17
timestamp 1692683681
transform 1 0 -2965 0 -1 -4869
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_18
timestamp 1692683681
transform 1 0 -2325 0 -1 -4869
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_19
timestamp 1692683681
transform -1 0 -2165 0 1 -4017
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_20
timestamp 1692683681
transform 1 0 -2805 0 -1 -5721
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_21
timestamp 1692683681
transform 1 0 -2965 0 -1 -5721
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_22
timestamp 1692683681
transform 1 0 -2325 0 -1 -5721
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_23
timestamp 1692683681
transform 1 0 -2325 0 1 -4017
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_24
timestamp 1692683681
transform 1 0 -2805 0 1 -3165
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_25
timestamp 1692683681
transform 1 0 -2965 0 1 -3165
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_26
timestamp 1692683681
transform -1 0 -2165 0 1 -3165
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_27
timestamp 1692683681
transform -1 0 -1685 0 1 -4017
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_28
timestamp 1692683681
transform -1 0 -1525 0 1 -4017
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_29
timestamp 1692683681
transform -1 0 -1525 0 1 -3165
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_30
timestamp 1692683681
transform -1 0 -1685 0 1 -3165
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_31
timestamp 1692683681
transform 1 0 -2325 0 1 -3165
box -202 -430 202 430
use pmos_3p3_MYZUUP  pmos_3p3_MYZUUP_0
timestamp 1692885173
transform 1 0 4281 0 1 -6443
box -230 -530 230 530
use pmos_3p3_MYZUUP  pmos_3p3_MYZUUP_1
timestamp 1692885173
transform 1 0 3027 0 1 -6442
box -230 -530 230 530
use pmos_3p3_MYZUUP  pmos_3p3_MYZUUP_2
timestamp 1692885173
transform 1 0 3617 0 1 -6442
box -230 -530 230 530
<< labels >>
flabel metal1 -1062 792 -1062 792 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
flabel metal1 -883 -7043 -883 -7043 0 FreeSans 1600 0 0 0 VSS
port 1 nsew
flabel via2 -3597 -2535 -3597 -2535 0 FreeSans 480 0 0 0 VINN
port 3 nsew
flabel via2 -3593 -2778 -3593 -2778 0 FreeSans 480 0 0 0 VINP
port 2 nsew
flabel metal1 672 -6091 672 -6091 0 FreeSans 640 0 0 0 OUT
port 7 nsew
flabel metal1 511 1917 511 1917 0 FreeSans 640 0 0 0 IBIAS
port 8 nsew
<< end >>
