magic
tech gf180mcuC
magscale 1 10
timestamp 1714491929
<< nwell >>
rect -60 958 881 1080
rect -60 908 -28 958
rect 830 908 881 958
<< psubdiff >>
rect -99 -349 894 -321
rect -99 -412 -83 -349
rect -14 -412 42 -349
rect 111 -412 167 -349
rect 236 -412 292 -349
rect 361 -412 417 -349
rect 486 -412 542 -349
rect 611 -412 667 -349
rect 736 -412 792 -349
rect 861 -412 894 -349
rect -99 -438 894 -412
<< nsubdiff >>
rect -9 1022 823 1036
rect -9 972 11 1022
rect 60 972 112 1022
rect 161 972 213 1022
rect 262 972 314 1022
rect 363 972 415 1022
rect 464 972 516 1022
rect 565 972 617 1022
rect 666 972 718 1022
rect 767 972 823 1022
rect -9 958 823 972
<< psubdiffcont >>
rect -83 -412 -14 -349
rect 42 -412 111 -349
rect 167 -412 236 -349
rect 292 -412 361 -349
rect 417 -412 486 -349
rect 542 -412 611 -349
rect 667 -412 736 -349
rect 792 -412 861 -349
<< nsubdiffcont >>
rect 11 972 60 1022
rect 112 972 161 1022
rect 213 972 262 1022
rect 314 972 363 1022
rect 415 972 464 1022
rect 516 972 565 1022
rect 617 972 666 1022
rect 718 972 767 1022
<< polysilicon >>
rect 114 216 184 247
rect 51 203 184 216
rect 51 148 66 203
rect 123 197 184 203
rect 288 197 358 246
rect 462 197 532 245
rect 636 197 706 241
rect 123 148 706 197
rect 51 144 706 148
rect 51 134 184 144
rect 114 103 184 134
rect 288 102 358 144
rect 462 101 532 144
rect 636 97 706 144
<< polycontact >>
rect 66 148 123 203
<< metal1 >>
rect -208 1119 1036 1236
rect -208 -320 -121 1119
rect -9 1022 823 1036
rect -9 972 11 1022
rect 60 972 112 1022
rect 161 972 213 1022
rect 262 972 314 1022
rect 363 972 415 1022
rect 464 972 516 1022
rect 565 972 617 1022
rect 666 972 718 1022
rect 767 972 823 1022
rect -9 958 823 972
rect 39 825 85 958
rect 387 829 433 958
rect 735 827 781 958
rect 51 203 134 216
rect 51 198 66 203
rect 7 152 66 198
rect 51 148 66 152
rect 123 148 134 203
rect 51 134 134 148
rect 213 190 259 302
rect 561 190 607 293
rect 213 144 766 190
rect 213 45 259 144
rect 561 36 607 144
rect -208 -321 -99 -320
rect 39 -321 85 -194
rect 387 -321 433 -188
rect 735 -321 781 -194
rect 927 -321 1036 1119
rect -208 -349 1036 -321
rect -208 -412 -83 -349
rect -14 -412 42 -349
rect 111 -412 167 -349
rect 236 -412 292 -349
rect 361 -412 417 -349
rect 486 -412 542 -349
rect 611 -412 667 -349
rect 736 -412 792 -349
rect 861 -412 1036 -349
rect -208 -438 1036 -412
use nmos_3p3_S7UZWU  nmos_3p3_S7UZWU_0
timestamp 1714126980
transform 1 0 410 0 1 -78
box -408 -208 408 208
use pmos_3p3_MD4UPK  pmos_3p3_MD4UPK_0
timestamp 1714126980
transform 1 0 410 0 1 562
box -470 -410 470 410
<< labels >>
flabel metal1 30 173 30 173 0 FreeSans 320 0 0 0 IN
port 1 nsew
flabel metal1 736 167 736 167 0 FreeSans 320 0 0 0 OUT
port 2 nsew
flabel metal1 403 -309 403 -309 0 FreeSans 320 0 0 0 VSS
port 4 nsew
flabel metal1 277 987 277 987 0 FreeSans 320 0 0 0 VDD
port 0 nsew
<< end >>
