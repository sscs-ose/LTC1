magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2421 -2045 2421 2045
<< psubdiff >>
rect -421 23 421 45
rect -421 -23 -399 23
rect 399 -23 421 23
rect -421 -45 421 -23
<< psubdiffcont >>
rect -399 -23 399 23
<< metal1 >>
rect -410 23 410 34
rect -410 -23 -399 23
rect 399 -23 410 23
rect -410 -34 410 -23
<< end >>
