magic
tech gf180mcuC
magscale 1 10
timestamp 1714558667
<< nwell >>
rect -70 1700 860 2228
<< nsubdiff >>
rect -32 2099 477 2193
<< metal1 >>
rect -70 2063 2901 2241
rect -206 1666 76 1738
rect 389 1675 500 1690
rect 389 1623 402 1675
rect 456 1623 500 1675
rect 389 1610 500 1623
rect 2952 1612 3133 1625
rect 2952 1502 3032 1612
rect 3116 1502 3133 1612
rect 2952 1496 3133 1502
rect -31 689 84 720
rect -31 629 -9 689
rect 51 629 84 689
rect -31 595 84 629
rect 1403 684 1502 686
rect 1403 632 1416 684
rect 1471 632 1502 684
rect 1403 629 1502 632
rect 1403 628 1483 629
rect 363 593 453 602
rect 363 532 377 593
rect 440 532 453 593
rect 363 522 453 532
rect 170 12 2895 189
<< via1 >>
rect 402 1623 456 1675
rect 3032 1502 3116 1612
rect 370 1016 427 1091
rect -9 629 51 689
rect 1416 632 1471 684
rect 377 532 440 593
<< metal2 >>
rect 361 1675 500 1688
rect 361 1623 402 1675
rect 456 1623 500 1675
rect 361 1615 500 1623
rect 364 1610 500 1615
rect 3020 1612 3133 1625
rect 364 1091 434 1610
rect 3020 1578 3032 1612
rect 2674 1522 3032 1578
rect 3020 1502 3032 1522
rect 3116 1502 3133 1612
rect 3020 1496 3133 1502
rect 364 1016 370 1091
rect 427 1016 434 1091
rect -31 689 84 720
rect -31 629 -9 689
rect 51 629 84 689
rect -31 595 84 629
rect 364 602 434 1016
rect 1384 692 1484 697
rect 1384 626 1394 692
rect 1473 626 1484 692
rect 1384 621 1484 626
rect 363 593 453 602
rect 363 532 377 593
rect 440 532 453 593
rect 363 522 453 532
<< via2 >>
rect -9 629 51 689
rect 1394 684 1473 692
rect 1394 632 1416 684
rect 1416 632 1471 684
rect 1471 632 1473 684
rect 1394 626 1473 632
<< metal3 >>
rect -31 696 84 720
rect -31 692 1502 696
rect -31 689 1394 692
rect -31 629 -9 689
rect 51 629 1394 689
rect -31 626 1394 629
rect 1473 626 1502 692
rect -31 620 1502 626
rect -31 595 84 620
use JK_FF_mag  JK_FF_mag_0
timestamp 1714558667
transform 1 0 320 0 1 80
box -430 0 2603 2148
<< labels >>
flabel metal1 925 105 925 105 0 FreeSans 640 0 0 0 VSS
port 0 nsew
flabel metal1 1080 2189 1080 2189 0 FreeSans 640 0 0 0 VDD
port 1 nsew
flabel metal2 2961 1553 2961 1553 0 FreeSans 640 0 0 0 Vdiv2
port 2 nsew
flabel metal1 -171 1702 -171 1702 0 FreeSans 640 0 0 0 CLK
port 3 nsew
flabel via2 20 657 20 657 0 FreeSans 640 0 0 0 RST
port 4 nsew
<< end >>
