magic
tech gf180mcuC
magscale 1 10
timestamp 1694765517
<< mimcap >>
rect -22269 21180 -17269 21260
rect -22269 16340 -22189 21180
rect -17349 16340 -17269 21180
rect -22269 16260 -17269 16340
rect -16655 21180 -11655 21260
rect -16655 16340 -16575 21180
rect -11735 16340 -11655 21180
rect -16655 16260 -11655 16340
rect -11041 21180 -6041 21260
rect -11041 16340 -10961 21180
rect -6121 16340 -6041 21180
rect -11041 16260 -6041 16340
rect -5427 21180 -427 21260
rect -5427 16340 -5347 21180
rect -507 16340 -427 21180
rect -5427 16260 -427 16340
rect 187 21180 5187 21260
rect 187 16340 267 21180
rect 5107 16340 5187 21180
rect 187 16260 5187 16340
rect 5801 21180 10801 21260
rect 5801 16340 5881 21180
rect 10721 16340 10801 21180
rect 5801 16260 10801 16340
rect 11415 21180 16415 21260
rect 11415 16340 11495 21180
rect 16335 16340 16415 21180
rect 11415 16260 16415 16340
rect 17029 21180 22029 21260
rect 17029 16340 17109 21180
rect 21949 16340 22029 21180
rect 17029 16260 22029 16340
rect -22269 15820 -17269 15900
rect -22269 10980 -22189 15820
rect -17349 10980 -17269 15820
rect -22269 10900 -17269 10980
rect -16655 15820 -11655 15900
rect -16655 10980 -16575 15820
rect -11735 10980 -11655 15820
rect -16655 10900 -11655 10980
rect -11041 15820 -6041 15900
rect -11041 10980 -10961 15820
rect -6121 10980 -6041 15820
rect -11041 10900 -6041 10980
rect -5427 15820 -427 15900
rect -5427 10980 -5347 15820
rect -507 10980 -427 15820
rect -5427 10900 -427 10980
rect 187 15820 5187 15900
rect 187 10980 267 15820
rect 5107 10980 5187 15820
rect 187 10900 5187 10980
rect 5801 15820 10801 15900
rect 5801 10980 5881 15820
rect 10721 10980 10801 15820
rect 5801 10900 10801 10980
rect 11415 15820 16415 15900
rect 11415 10980 11495 15820
rect 16335 10980 16415 15820
rect 11415 10900 16415 10980
rect 17029 15820 22029 15900
rect 17029 10980 17109 15820
rect 21949 10980 22029 15820
rect 17029 10900 22029 10980
rect -22269 10460 -17269 10540
rect -22269 5620 -22189 10460
rect -17349 5620 -17269 10460
rect -22269 5540 -17269 5620
rect -16655 10460 -11655 10540
rect -16655 5620 -16575 10460
rect -11735 5620 -11655 10460
rect -16655 5540 -11655 5620
rect -11041 10460 -6041 10540
rect -11041 5620 -10961 10460
rect -6121 5620 -6041 10460
rect -11041 5540 -6041 5620
rect -5427 10460 -427 10540
rect -5427 5620 -5347 10460
rect -507 5620 -427 10460
rect -5427 5540 -427 5620
rect 187 10460 5187 10540
rect 187 5620 267 10460
rect 5107 5620 5187 10460
rect 187 5540 5187 5620
rect 5801 10460 10801 10540
rect 5801 5620 5881 10460
rect 10721 5620 10801 10460
rect 5801 5540 10801 5620
rect 11415 10460 16415 10540
rect 11415 5620 11495 10460
rect 16335 5620 16415 10460
rect 11415 5540 16415 5620
rect 17029 10460 22029 10540
rect 17029 5620 17109 10460
rect 21949 5620 22029 10460
rect 17029 5540 22029 5620
rect -22269 5100 -17269 5180
rect -22269 260 -22189 5100
rect -17349 260 -17269 5100
rect -22269 180 -17269 260
rect -16655 5100 -11655 5180
rect -16655 260 -16575 5100
rect -11735 260 -11655 5100
rect -16655 180 -11655 260
rect -11041 5100 -6041 5180
rect -11041 260 -10961 5100
rect -6121 260 -6041 5100
rect -11041 180 -6041 260
rect -5427 5100 -427 5180
rect -5427 260 -5347 5100
rect -507 260 -427 5100
rect -5427 180 -427 260
rect 187 5100 5187 5180
rect 187 260 267 5100
rect 5107 260 5187 5100
rect 187 180 5187 260
rect 5801 5100 10801 5180
rect 5801 260 5881 5100
rect 10721 260 10801 5100
rect 5801 180 10801 260
rect 11415 5100 16415 5180
rect 11415 260 11495 5100
rect 16335 260 16415 5100
rect 11415 180 16415 260
rect 17029 5100 22029 5180
rect 17029 260 17109 5100
rect 21949 260 22029 5100
rect 17029 180 22029 260
rect -22269 -260 -17269 -180
rect -22269 -5100 -22189 -260
rect -17349 -5100 -17269 -260
rect -22269 -5180 -17269 -5100
rect -16655 -260 -11655 -180
rect -16655 -5100 -16575 -260
rect -11735 -5100 -11655 -260
rect -16655 -5180 -11655 -5100
rect -11041 -260 -6041 -180
rect -11041 -5100 -10961 -260
rect -6121 -5100 -6041 -260
rect -11041 -5180 -6041 -5100
rect -5427 -260 -427 -180
rect -5427 -5100 -5347 -260
rect -507 -5100 -427 -260
rect -5427 -5180 -427 -5100
rect 187 -260 5187 -180
rect 187 -5100 267 -260
rect 5107 -5100 5187 -260
rect 187 -5180 5187 -5100
rect 5801 -260 10801 -180
rect 5801 -5100 5881 -260
rect 10721 -5100 10801 -260
rect 5801 -5180 10801 -5100
rect 11415 -260 16415 -180
rect 11415 -5100 11495 -260
rect 16335 -5100 16415 -260
rect 11415 -5180 16415 -5100
rect 17029 -260 22029 -180
rect 17029 -5100 17109 -260
rect 21949 -5100 22029 -260
rect 17029 -5180 22029 -5100
rect -22269 -5620 -17269 -5540
rect -22269 -10460 -22189 -5620
rect -17349 -10460 -17269 -5620
rect -22269 -10540 -17269 -10460
rect -16655 -5620 -11655 -5540
rect -16655 -10460 -16575 -5620
rect -11735 -10460 -11655 -5620
rect -16655 -10540 -11655 -10460
rect -11041 -5620 -6041 -5540
rect -11041 -10460 -10961 -5620
rect -6121 -10460 -6041 -5620
rect -11041 -10540 -6041 -10460
rect -5427 -5620 -427 -5540
rect -5427 -10460 -5347 -5620
rect -507 -10460 -427 -5620
rect -5427 -10540 -427 -10460
rect 187 -5620 5187 -5540
rect 187 -10460 267 -5620
rect 5107 -10460 5187 -5620
rect 187 -10540 5187 -10460
rect 5801 -5620 10801 -5540
rect 5801 -10460 5881 -5620
rect 10721 -10460 10801 -5620
rect 5801 -10540 10801 -10460
rect 11415 -5620 16415 -5540
rect 11415 -10460 11495 -5620
rect 16335 -10460 16415 -5620
rect 11415 -10540 16415 -10460
rect 17029 -5620 22029 -5540
rect 17029 -10460 17109 -5620
rect 21949 -10460 22029 -5620
rect 17029 -10540 22029 -10460
rect -22269 -10980 -17269 -10900
rect -22269 -15820 -22189 -10980
rect -17349 -15820 -17269 -10980
rect -22269 -15900 -17269 -15820
rect -16655 -10980 -11655 -10900
rect -16655 -15820 -16575 -10980
rect -11735 -15820 -11655 -10980
rect -16655 -15900 -11655 -15820
rect -11041 -10980 -6041 -10900
rect -11041 -15820 -10961 -10980
rect -6121 -15820 -6041 -10980
rect -11041 -15900 -6041 -15820
rect -5427 -10980 -427 -10900
rect -5427 -15820 -5347 -10980
rect -507 -15820 -427 -10980
rect -5427 -15900 -427 -15820
rect 187 -10980 5187 -10900
rect 187 -15820 267 -10980
rect 5107 -15820 5187 -10980
rect 187 -15900 5187 -15820
rect 5801 -10980 10801 -10900
rect 5801 -15820 5881 -10980
rect 10721 -15820 10801 -10980
rect 5801 -15900 10801 -15820
rect 11415 -10980 16415 -10900
rect 11415 -15820 11495 -10980
rect 16335 -15820 16415 -10980
rect 11415 -15900 16415 -15820
rect 17029 -10980 22029 -10900
rect 17029 -15820 17109 -10980
rect 21949 -15820 22029 -10980
rect 17029 -15900 22029 -15820
rect -22269 -16340 -17269 -16260
rect -22269 -21180 -22189 -16340
rect -17349 -21180 -17269 -16340
rect -22269 -21260 -17269 -21180
rect -16655 -16340 -11655 -16260
rect -16655 -21180 -16575 -16340
rect -11735 -21180 -11655 -16340
rect -16655 -21260 -11655 -21180
rect -11041 -16340 -6041 -16260
rect -11041 -21180 -10961 -16340
rect -6121 -21180 -6041 -16340
rect -11041 -21260 -6041 -21180
rect -5427 -16340 -427 -16260
rect -5427 -21180 -5347 -16340
rect -507 -21180 -427 -16340
rect -5427 -21260 -427 -21180
rect 187 -16340 5187 -16260
rect 187 -21180 267 -16340
rect 5107 -21180 5187 -16340
rect 187 -21260 5187 -21180
rect 5801 -16340 10801 -16260
rect 5801 -21180 5881 -16340
rect 10721 -21180 10801 -16340
rect 5801 -21260 10801 -21180
rect 11415 -16340 16415 -16260
rect 11415 -21180 11495 -16340
rect 16335 -21180 16415 -16340
rect 11415 -21260 16415 -21180
rect 17029 -16340 22029 -16260
rect 17029 -21180 17109 -16340
rect 21949 -21180 22029 -16340
rect 17029 -21260 22029 -21180
<< mimcapcontact >>
rect -22189 16340 -17349 21180
rect -16575 16340 -11735 21180
rect -10961 16340 -6121 21180
rect -5347 16340 -507 21180
rect 267 16340 5107 21180
rect 5881 16340 10721 21180
rect 11495 16340 16335 21180
rect 17109 16340 21949 21180
rect -22189 10980 -17349 15820
rect -16575 10980 -11735 15820
rect -10961 10980 -6121 15820
rect -5347 10980 -507 15820
rect 267 10980 5107 15820
rect 5881 10980 10721 15820
rect 11495 10980 16335 15820
rect 17109 10980 21949 15820
rect -22189 5620 -17349 10460
rect -16575 5620 -11735 10460
rect -10961 5620 -6121 10460
rect -5347 5620 -507 10460
rect 267 5620 5107 10460
rect 5881 5620 10721 10460
rect 11495 5620 16335 10460
rect 17109 5620 21949 10460
rect -22189 260 -17349 5100
rect -16575 260 -11735 5100
rect -10961 260 -6121 5100
rect -5347 260 -507 5100
rect 267 260 5107 5100
rect 5881 260 10721 5100
rect 11495 260 16335 5100
rect 17109 260 21949 5100
rect -22189 -5100 -17349 -260
rect -16575 -5100 -11735 -260
rect -10961 -5100 -6121 -260
rect -5347 -5100 -507 -260
rect 267 -5100 5107 -260
rect 5881 -5100 10721 -260
rect 11495 -5100 16335 -260
rect 17109 -5100 21949 -260
rect -22189 -10460 -17349 -5620
rect -16575 -10460 -11735 -5620
rect -10961 -10460 -6121 -5620
rect -5347 -10460 -507 -5620
rect 267 -10460 5107 -5620
rect 5881 -10460 10721 -5620
rect 11495 -10460 16335 -5620
rect 17109 -10460 21949 -5620
rect -22189 -15820 -17349 -10980
rect -16575 -15820 -11735 -10980
rect -10961 -15820 -6121 -10980
rect -5347 -15820 -507 -10980
rect 267 -15820 5107 -10980
rect 5881 -15820 10721 -10980
rect 11495 -15820 16335 -10980
rect 17109 -15820 21949 -10980
rect -22189 -21180 -17349 -16340
rect -16575 -21180 -11735 -16340
rect -10961 -21180 -6121 -16340
rect -5347 -21180 -507 -16340
rect 267 -21180 5107 -16340
rect 5881 -21180 10721 -16340
rect 11495 -21180 16335 -16340
rect 17109 -21180 21949 -16340
<< metal4 >>
rect -22389 21313 -16909 21380
rect -22389 21260 -17059 21313
rect -22389 16260 -22269 21260
rect -17269 16260 -17059 21260
rect -22389 16207 -17059 16260
rect -16971 16207 -16909 21313
rect -22389 16140 -16909 16207
rect -16775 21313 -11295 21380
rect -16775 21260 -11445 21313
rect -16775 16260 -16655 21260
rect -11655 16260 -11445 21260
rect -16775 16207 -11445 16260
rect -11357 16207 -11295 21313
rect -16775 16140 -11295 16207
rect -11161 21313 -5681 21380
rect -11161 21260 -5831 21313
rect -11161 16260 -11041 21260
rect -6041 16260 -5831 21260
rect -11161 16207 -5831 16260
rect -5743 16207 -5681 21313
rect -11161 16140 -5681 16207
rect -5547 21313 -67 21380
rect -5547 21260 -217 21313
rect -5547 16260 -5427 21260
rect -427 16260 -217 21260
rect -5547 16207 -217 16260
rect -129 16207 -67 21313
rect -5547 16140 -67 16207
rect 67 21313 5547 21380
rect 67 21260 5397 21313
rect 67 16260 187 21260
rect 5187 16260 5397 21260
rect 67 16207 5397 16260
rect 5485 16207 5547 21313
rect 67 16140 5547 16207
rect 5681 21313 11161 21380
rect 5681 21260 11011 21313
rect 5681 16260 5801 21260
rect 10801 16260 11011 21260
rect 5681 16207 11011 16260
rect 11099 16207 11161 21313
rect 5681 16140 11161 16207
rect 11295 21313 16775 21380
rect 11295 21260 16625 21313
rect 11295 16260 11415 21260
rect 16415 16260 16625 21260
rect 11295 16207 16625 16260
rect 16713 16207 16775 21313
rect 11295 16140 16775 16207
rect 16909 21313 22389 21380
rect 16909 21260 22239 21313
rect 16909 16260 17029 21260
rect 22029 16260 22239 21260
rect 16909 16207 22239 16260
rect 22327 16207 22389 21313
rect 16909 16140 22389 16207
rect -22389 15953 -16909 16020
rect -22389 15900 -17059 15953
rect -22389 10900 -22269 15900
rect -17269 10900 -17059 15900
rect -22389 10847 -17059 10900
rect -16971 10847 -16909 15953
rect -22389 10780 -16909 10847
rect -16775 15953 -11295 16020
rect -16775 15900 -11445 15953
rect -16775 10900 -16655 15900
rect -11655 10900 -11445 15900
rect -16775 10847 -11445 10900
rect -11357 10847 -11295 15953
rect -16775 10780 -11295 10847
rect -11161 15953 -5681 16020
rect -11161 15900 -5831 15953
rect -11161 10900 -11041 15900
rect -6041 10900 -5831 15900
rect -11161 10847 -5831 10900
rect -5743 10847 -5681 15953
rect -11161 10780 -5681 10847
rect -5547 15953 -67 16020
rect -5547 15900 -217 15953
rect -5547 10900 -5427 15900
rect -427 10900 -217 15900
rect -5547 10847 -217 10900
rect -129 10847 -67 15953
rect -5547 10780 -67 10847
rect 67 15953 5547 16020
rect 67 15900 5397 15953
rect 67 10900 187 15900
rect 5187 10900 5397 15900
rect 67 10847 5397 10900
rect 5485 10847 5547 15953
rect 67 10780 5547 10847
rect 5681 15953 11161 16020
rect 5681 15900 11011 15953
rect 5681 10900 5801 15900
rect 10801 10900 11011 15900
rect 5681 10847 11011 10900
rect 11099 10847 11161 15953
rect 5681 10780 11161 10847
rect 11295 15953 16775 16020
rect 11295 15900 16625 15953
rect 11295 10900 11415 15900
rect 16415 10900 16625 15900
rect 11295 10847 16625 10900
rect 16713 10847 16775 15953
rect 11295 10780 16775 10847
rect 16909 15953 22389 16020
rect 16909 15900 22239 15953
rect 16909 10900 17029 15900
rect 22029 10900 22239 15900
rect 16909 10847 22239 10900
rect 22327 10847 22389 15953
rect 16909 10780 22389 10847
rect -22389 10593 -16909 10660
rect -22389 10540 -17059 10593
rect -22389 5540 -22269 10540
rect -17269 5540 -17059 10540
rect -22389 5487 -17059 5540
rect -16971 5487 -16909 10593
rect -22389 5420 -16909 5487
rect -16775 10593 -11295 10660
rect -16775 10540 -11445 10593
rect -16775 5540 -16655 10540
rect -11655 5540 -11445 10540
rect -16775 5487 -11445 5540
rect -11357 5487 -11295 10593
rect -16775 5420 -11295 5487
rect -11161 10593 -5681 10660
rect -11161 10540 -5831 10593
rect -11161 5540 -11041 10540
rect -6041 5540 -5831 10540
rect -11161 5487 -5831 5540
rect -5743 5487 -5681 10593
rect -11161 5420 -5681 5487
rect -5547 10593 -67 10660
rect -5547 10540 -217 10593
rect -5547 5540 -5427 10540
rect -427 5540 -217 10540
rect -5547 5487 -217 5540
rect -129 5487 -67 10593
rect -5547 5420 -67 5487
rect 67 10593 5547 10660
rect 67 10540 5397 10593
rect 67 5540 187 10540
rect 5187 5540 5397 10540
rect 67 5487 5397 5540
rect 5485 5487 5547 10593
rect 67 5420 5547 5487
rect 5681 10593 11161 10660
rect 5681 10540 11011 10593
rect 5681 5540 5801 10540
rect 10801 5540 11011 10540
rect 5681 5487 11011 5540
rect 11099 5487 11161 10593
rect 5681 5420 11161 5487
rect 11295 10593 16775 10660
rect 11295 10540 16625 10593
rect 11295 5540 11415 10540
rect 16415 5540 16625 10540
rect 11295 5487 16625 5540
rect 16713 5487 16775 10593
rect 11295 5420 16775 5487
rect 16909 10593 22389 10660
rect 16909 10540 22239 10593
rect 16909 5540 17029 10540
rect 22029 5540 22239 10540
rect 16909 5487 22239 5540
rect 22327 5487 22389 10593
rect 16909 5420 22389 5487
rect -22389 5233 -16909 5300
rect -22389 5180 -17059 5233
rect -22389 180 -22269 5180
rect -17269 180 -17059 5180
rect -22389 127 -17059 180
rect -16971 127 -16909 5233
rect -22389 60 -16909 127
rect -16775 5233 -11295 5300
rect -16775 5180 -11445 5233
rect -16775 180 -16655 5180
rect -11655 180 -11445 5180
rect -16775 127 -11445 180
rect -11357 127 -11295 5233
rect -16775 60 -11295 127
rect -11161 5233 -5681 5300
rect -11161 5180 -5831 5233
rect -11161 180 -11041 5180
rect -6041 180 -5831 5180
rect -11161 127 -5831 180
rect -5743 127 -5681 5233
rect -11161 60 -5681 127
rect -5547 5233 -67 5300
rect -5547 5180 -217 5233
rect -5547 180 -5427 5180
rect -427 180 -217 5180
rect -5547 127 -217 180
rect -129 127 -67 5233
rect -5547 60 -67 127
rect 67 5233 5547 5300
rect 67 5180 5397 5233
rect 67 180 187 5180
rect 5187 180 5397 5180
rect 67 127 5397 180
rect 5485 127 5547 5233
rect 67 60 5547 127
rect 5681 5233 11161 5300
rect 5681 5180 11011 5233
rect 5681 180 5801 5180
rect 10801 180 11011 5180
rect 5681 127 11011 180
rect 11099 127 11161 5233
rect 5681 60 11161 127
rect 11295 5233 16775 5300
rect 11295 5180 16625 5233
rect 11295 180 11415 5180
rect 16415 180 16625 5180
rect 11295 127 16625 180
rect 16713 127 16775 5233
rect 11295 60 16775 127
rect 16909 5233 22389 5300
rect 16909 5180 22239 5233
rect 16909 180 17029 5180
rect 22029 180 22239 5180
rect 16909 127 22239 180
rect 22327 127 22389 5233
rect 16909 60 22389 127
rect -22389 -127 -16909 -60
rect -22389 -180 -17059 -127
rect -22389 -5180 -22269 -180
rect -17269 -5180 -17059 -180
rect -22389 -5233 -17059 -5180
rect -16971 -5233 -16909 -127
rect -22389 -5300 -16909 -5233
rect -16775 -127 -11295 -60
rect -16775 -180 -11445 -127
rect -16775 -5180 -16655 -180
rect -11655 -5180 -11445 -180
rect -16775 -5233 -11445 -5180
rect -11357 -5233 -11295 -127
rect -16775 -5300 -11295 -5233
rect -11161 -127 -5681 -60
rect -11161 -180 -5831 -127
rect -11161 -5180 -11041 -180
rect -6041 -5180 -5831 -180
rect -11161 -5233 -5831 -5180
rect -5743 -5233 -5681 -127
rect -11161 -5300 -5681 -5233
rect -5547 -127 -67 -60
rect -5547 -180 -217 -127
rect -5547 -5180 -5427 -180
rect -427 -5180 -217 -180
rect -5547 -5233 -217 -5180
rect -129 -5233 -67 -127
rect -5547 -5300 -67 -5233
rect 67 -127 5547 -60
rect 67 -180 5397 -127
rect 67 -5180 187 -180
rect 5187 -5180 5397 -180
rect 67 -5233 5397 -5180
rect 5485 -5233 5547 -127
rect 67 -5300 5547 -5233
rect 5681 -127 11161 -60
rect 5681 -180 11011 -127
rect 5681 -5180 5801 -180
rect 10801 -5180 11011 -180
rect 5681 -5233 11011 -5180
rect 11099 -5233 11161 -127
rect 5681 -5300 11161 -5233
rect 11295 -127 16775 -60
rect 11295 -180 16625 -127
rect 11295 -5180 11415 -180
rect 16415 -5180 16625 -180
rect 11295 -5233 16625 -5180
rect 16713 -5233 16775 -127
rect 11295 -5300 16775 -5233
rect 16909 -127 22389 -60
rect 16909 -180 22239 -127
rect 16909 -5180 17029 -180
rect 22029 -5180 22239 -180
rect 16909 -5233 22239 -5180
rect 22327 -5233 22389 -127
rect 16909 -5300 22389 -5233
rect -22389 -5487 -16909 -5420
rect -22389 -5540 -17059 -5487
rect -22389 -10540 -22269 -5540
rect -17269 -10540 -17059 -5540
rect -22389 -10593 -17059 -10540
rect -16971 -10593 -16909 -5487
rect -22389 -10660 -16909 -10593
rect -16775 -5487 -11295 -5420
rect -16775 -5540 -11445 -5487
rect -16775 -10540 -16655 -5540
rect -11655 -10540 -11445 -5540
rect -16775 -10593 -11445 -10540
rect -11357 -10593 -11295 -5487
rect -16775 -10660 -11295 -10593
rect -11161 -5487 -5681 -5420
rect -11161 -5540 -5831 -5487
rect -11161 -10540 -11041 -5540
rect -6041 -10540 -5831 -5540
rect -11161 -10593 -5831 -10540
rect -5743 -10593 -5681 -5487
rect -11161 -10660 -5681 -10593
rect -5547 -5487 -67 -5420
rect -5547 -5540 -217 -5487
rect -5547 -10540 -5427 -5540
rect -427 -10540 -217 -5540
rect -5547 -10593 -217 -10540
rect -129 -10593 -67 -5487
rect -5547 -10660 -67 -10593
rect 67 -5487 5547 -5420
rect 67 -5540 5397 -5487
rect 67 -10540 187 -5540
rect 5187 -10540 5397 -5540
rect 67 -10593 5397 -10540
rect 5485 -10593 5547 -5487
rect 67 -10660 5547 -10593
rect 5681 -5487 11161 -5420
rect 5681 -5540 11011 -5487
rect 5681 -10540 5801 -5540
rect 10801 -10540 11011 -5540
rect 5681 -10593 11011 -10540
rect 11099 -10593 11161 -5487
rect 5681 -10660 11161 -10593
rect 11295 -5487 16775 -5420
rect 11295 -5540 16625 -5487
rect 11295 -10540 11415 -5540
rect 16415 -10540 16625 -5540
rect 11295 -10593 16625 -10540
rect 16713 -10593 16775 -5487
rect 11295 -10660 16775 -10593
rect 16909 -5487 22389 -5420
rect 16909 -5540 22239 -5487
rect 16909 -10540 17029 -5540
rect 22029 -10540 22239 -5540
rect 16909 -10593 22239 -10540
rect 22327 -10593 22389 -5487
rect 16909 -10660 22389 -10593
rect -22389 -10847 -16909 -10780
rect -22389 -10900 -17059 -10847
rect -22389 -15900 -22269 -10900
rect -17269 -15900 -17059 -10900
rect -22389 -15953 -17059 -15900
rect -16971 -15953 -16909 -10847
rect -22389 -16020 -16909 -15953
rect -16775 -10847 -11295 -10780
rect -16775 -10900 -11445 -10847
rect -16775 -15900 -16655 -10900
rect -11655 -15900 -11445 -10900
rect -16775 -15953 -11445 -15900
rect -11357 -15953 -11295 -10847
rect -16775 -16020 -11295 -15953
rect -11161 -10847 -5681 -10780
rect -11161 -10900 -5831 -10847
rect -11161 -15900 -11041 -10900
rect -6041 -15900 -5831 -10900
rect -11161 -15953 -5831 -15900
rect -5743 -15953 -5681 -10847
rect -11161 -16020 -5681 -15953
rect -5547 -10847 -67 -10780
rect -5547 -10900 -217 -10847
rect -5547 -15900 -5427 -10900
rect -427 -15900 -217 -10900
rect -5547 -15953 -217 -15900
rect -129 -15953 -67 -10847
rect -5547 -16020 -67 -15953
rect 67 -10847 5547 -10780
rect 67 -10900 5397 -10847
rect 67 -15900 187 -10900
rect 5187 -15900 5397 -10900
rect 67 -15953 5397 -15900
rect 5485 -15953 5547 -10847
rect 67 -16020 5547 -15953
rect 5681 -10847 11161 -10780
rect 5681 -10900 11011 -10847
rect 5681 -15900 5801 -10900
rect 10801 -15900 11011 -10900
rect 5681 -15953 11011 -15900
rect 11099 -15953 11161 -10847
rect 5681 -16020 11161 -15953
rect 11295 -10847 16775 -10780
rect 11295 -10900 16625 -10847
rect 11295 -15900 11415 -10900
rect 16415 -15900 16625 -10900
rect 11295 -15953 16625 -15900
rect 16713 -15953 16775 -10847
rect 11295 -16020 16775 -15953
rect 16909 -10847 22389 -10780
rect 16909 -10900 22239 -10847
rect 16909 -15900 17029 -10900
rect 22029 -15900 22239 -10900
rect 16909 -15953 22239 -15900
rect 22327 -15953 22389 -10847
rect 16909 -16020 22389 -15953
rect -22389 -16207 -16909 -16140
rect -22389 -16260 -17059 -16207
rect -22389 -21260 -22269 -16260
rect -17269 -21260 -17059 -16260
rect -22389 -21313 -17059 -21260
rect -16971 -21313 -16909 -16207
rect -22389 -21380 -16909 -21313
rect -16775 -16207 -11295 -16140
rect -16775 -16260 -11445 -16207
rect -16775 -21260 -16655 -16260
rect -11655 -21260 -11445 -16260
rect -16775 -21313 -11445 -21260
rect -11357 -21313 -11295 -16207
rect -16775 -21380 -11295 -21313
rect -11161 -16207 -5681 -16140
rect -11161 -16260 -5831 -16207
rect -11161 -21260 -11041 -16260
rect -6041 -21260 -5831 -16260
rect -11161 -21313 -5831 -21260
rect -5743 -21313 -5681 -16207
rect -11161 -21380 -5681 -21313
rect -5547 -16207 -67 -16140
rect -5547 -16260 -217 -16207
rect -5547 -21260 -5427 -16260
rect -427 -21260 -217 -16260
rect -5547 -21313 -217 -21260
rect -129 -21313 -67 -16207
rect -5547 -21380 -67 -21313
rect 67 -16207 5547 -16140
rect 67 -16260 5397 -16207
rect 67 -21260 187 -16260
rect 5187 -21260 5397 -16260
rect 67 -21313 5397 -21260
rect 5485 -21313 5547 -16207
rect 67 -21380 5547 -21313
rect 5681 -16207 11161 -16140
rect 5681 -16260 11011 -16207
rect 5681 -21260 5801 -16260
rect 10801 -21260 11011 -16260
rect 5681 -21313 11011 -21260
rect 11099 -21313 11161 -16207
rect 5681 -21380 11161 -21313
rect 11295 -16207 16775 -16140
rect 11295 -16260 16625 -16207
rect 11295 -21260 11415 -16260
rect 16415 -21260 16625 -16260
rect 11295 -21313 16625 -21260
rect 16713 -21313 16775 -16207
rect 11295 -21380 16775 -21313
rect 16909 -16207 22389 -16140
rect 16909 -16260 22239 -16207
rect 16909 -21260 17029 -16260
rect 22029 -21260 22239 -16260
rect 16909 -21313 22239 -21260
rect 22327 -21313 22389 -16207
rect 16909 -21380 22389 -21313
<< via4 >>
rect -17059 16207 -16971 21313
rect -11445 16207 -11357 21313
rect -5831 16207 -5743 21313
rect -217 16207 -129 21313
rect 5397 16207 5485 21313
rect 11011 16207 11099 21313
rect 16625 16207 16713 21313
rect 22239 16207 22327 21313
rect -17059 10847 -16971 15953
rect -11445 10847 -11357 15953
rect -5831 10847 -5743 15953
rect -217 10847 -129 15953
rect 5397 10847 5485 15953
rect 11011 10847 11099 15953
rect 16625 10847 16713 15953
rect 22239 10847 22327 15953
rect -17059 5487 -16971 10593
rect -11445 5487 -11357 10593
rect -5831 5487 -5743 10593
rect -217 5487 -129 10593
rect 5397 5487 5485 10593
rect 11011 5487 11099 10593
rect 16625 5487 16713 10593
rect 22239 5487 22327 10593
rect -17059 127 -16971 5233
rect -11445 127 -11357 5233
rect -5831 127 -5743 5233
rect -217 127 -129 5233
rect 5397 127 5485 5233
rect 11011 127 11099 5233
rect 16625 127 16713 5233
rect 22239 127 22327 5233
rect -17059 -5233 -16971 -127
rect -11445 -5233 -11357 -127
rect -5831 -5233 -5743 -127
rect -217 -5233 -129 -127
rect 5397 -5233 5485 -127
rect 11011 -5233 11099 -127
rect 16625 -5233 16713 -127
rect 22239 -5233 22327 -127
rect -17059 -10593 -16971 -5487
rect -11445 -10593 -11357 -5487
rect -5831 -10593 -5743 -5487
rect -217 -10593 -129 -5487
rect 5397 -10593 5485 -5487
rect 11011 -10593 11099 -5487
rect 16625 -10593 16713 -5487
rect 22239 -10593 22327 -5487
rect -17059 -15953 -16971 -10847
rect -11445 -15953 -11357 -10847
rect -5831 -15953 -5743 -10847
rect -217 -15953 -129 -10847
rect 5397 -15953 5485 -10847
rect 11011 -15953 11099 -10847
rect 16625 -15953 16713 -10847
rect 22239 -15953 22327 -10847
rect -17059 -21313 -16971 -16207
rect -11445 -21313 -11357 -16207
rect -5831 -21313 -5743 -16207
rect -217 -21313 -129 -16207
rect 5397 -21313 5485 -16207
rect 11011 -21313 11099 -16207
rect 16625 -21313 16713 -16207
rect 22239 -21313 22327 -16207
<< metal5 >>
rect -19875 21180 -19663 21440
rect -17121 21313 -16909 21440
rect -19875 15820 -19663 16340
rect -17121 16207 -17059 21313
rect -16971 16207 -16909 21313
rect -14261 21180 -14049 21440
rect -11507 21313 -11295 21440
rect -17121 15953 -16909 16207
rect -19875 10460 -19663 10980
rect -17121 10847 -17059 15953
rect -16971 10847 -16909 15953
rect -14261 15820 -14049 16340
rect -11507 16207 -11445 21313
rect -11357 16207 -11295 21313
rect -8647 21180 -8435 21440
rect -5893 21313 -5681 21440
rect -11507 15953 -11295 16207
rect -17121 10593 -16909 10847
rect -19875 5100 -19663 5620
rect -17121 5487 -17059 10593
rect -16971 5487 -16909 10593
rect -14261 10460 -14049 10980
rect -11507 10847 -11445 15953
rect -11357 10847 -11295 15953
rect -8647 15820 -8435 16340
rect -5893 16207 -5831 21313
rect -5743 16207 -5681 21313
rect -3033 21180 -2821 21440
rect -279 21313 -67 21440
rect -5893 15953 -5681 16207
rect -11507 10593 -11295 10847
rect -17121 5233 -16909 5487
rect -19875 -260 -19663 260
rect -17121 127 -17059 5233
rect -16971 127 -16909 5233
rect -14261 5100 -14049 5620
rect -11507 5487 -11445 10593
rect -11357 5487 -11295 10593
rect -8647 10460 -8435 10980
rect -5893 10847 -5831 15953
rect -5743 10847 -5681 15953
rect -3033 15820 -2821 16340
rect -279 16207 -217 21313
rect -129 16207 -67 21313
rect 2581 21180 2793 21440
rect 5335 21313 5547 21440
rect -279 15953 -67 16207
rect -5893 10593 -5681 10847
rect -11507 5233 -11295 5487
rect -17121 -127 -16909 127
rect -19875 -5620 -19663 -5100
rect -17121 -5233 -17059 -127
rect -16971 -5233 -16909 -127
rect -14261 -260 -14049 260
rect -11507 127 -11445 5233
rect -11357 127 -11295 5233
rect -8647 5100 -8435 5620
rect -5893 5487 -5831 10593
rect -5743 5487 -5681 10593
rect -3033 10460 -2821 10980
rect -279 10847 -217 15953
rect -129 10847 -67 15953
rect 2581 15820 2793 16340
rect 5335 16207 5397 21313
rect 5485 16207 5547 21313
rect 8195 21180 8407 21440
rect 10949 21313 11161 21440
rect 5335 15953 5547 16207
rect -279 10593 -67 10847
rect -5893 5233 -5681 5487
rect -11507 -127 -11295 127
rect -17121 -5487 -16909 -5233
rect -19875 -10980 -19663 -10460
rect -17121 -10593 -17059 -5487
rect -16971 -10593 -16909 -5487
rect -14261 -5620 -14049 -5100
rect -11507 -5233 -11445 -127
rect -11357 -5233 -11295 -127
rect -8647 -260 -8435 260
rect -5893 127 -5831 5233
rect -5743 127 -5681 5233
rect -3033 5100 -2821 5620
rect -279 5487 -217 10593
rect -129 5487 -67 10593
rect 2581 10460 2793 10980
rect 5335 10847 5397 15953
rect 5485 10847 5547 15953
rect 8195 15820 8407 16340
rect 10949 16207 11011 21313
rect 11099 16207 11161 21313
rect 13809 21180 14021 21440
rect 16563 21313 16775 21440
rect 10949 15953 11161 16207
rect 5335 10593 5547 10847
rect -279 5233 -67 5487
rect -5893 -127 -5681 127
rect -11507 -5487 -11295 -5233
rect -17121 -10847 -16909 -10593
rect -19875 -16340 -19663 -15820
rect -17121 -15953 -17059 -10847
rect -16971 -15953 -16909 -10847
rect -14261 -10980 -14049 -10460
rect -11507 -10593 -11445 -5487
rect -11357 -10593 -11295 -5487
rect -8647 -5620 -8435 -5100
rect -5893 -5233 -5831 -127
rect -5743 -5233 -5681 -127
rect -3033 -260 -2821 260
rect -279 127 -217 5233
rect -129 127 -67 5233
rect 2581 5100 2793 5620
rect 5335 5487 5397 10593
rect 5485 5487 5547 10593
rect 8195 10460 8407 10980
rect 10949 10847 11011 15953
rect 11099 10847 11161 15953
rect 13809 15820 14021 16340
rect 16563 16207 16625 21313
rect 16713 16207 16775 21313
rect 19423 21180 19635 21440
rect 22177 21313 22389 21440
rect 16563 15953 16775 16207
rect 10949 10593 11161 10847
rect 5335 5233 5547 5487
rect -279 -127 -67 127
rect -5893 -5487 -5681 -5233
rect -11507 -10847 -11295 -10593
rect -17121 -16207 -16909 -15953
rect -19875 -21440 -19663 -21180
rect -17121 -21313 -17059 -16207
rect -16971 -21313 -16909 -16207
rect -14261 -16340 -14049 -15820
rect -11507 -15953 -11445 -10847
rect -11357 -15953 -11295 -10847
rect -8647 -10980 -8435 -10460
rect -5893 -10593 -5831 -5487
rect -5743 -10593 -5681 -5487
rect -3033 -5620 -2821 -5100
rect -279 -5233 -217 -127
rect -129 -5233 -67 -127
rect 2581 -260 2793 260
rect 5335 127 5397 5233
rect 5485 127 5547 5233
rect 8195 5100 8407 5620
rect 10949 5487 11011 10593
rect 11099 5487 11161 10593
rect 13809 10460 14021 10980
rect 16563 10847 16625 15953
rect 16713 10847 16775 15953
rect 19423 15820 19635 16340
rect 22177 16207 22239 21313
rect 22327 16207 22389 21313
rect 22177 15953 22389 16207
rect 16563 10593 16775 10847
rect 10949 5233 11161 5487
rect 5335 -127 5547 127
rect -279 -5487 -67 -5233
rect -5893 -10847 -5681 -10593
rect -11507 -16207 -11295 -15953
rect -17121 -21440 -16909 -21313
rect -14261 -21440 -14049 -21180
rect -11507 -21313 -11445 -16207
rect -11357 -21313 -11295 -16207
rect -8647 -16340 -8435 -15820
rect -5893 -15953 -5831 -10847
rect -5743 -15953 -5681 -10847
rect -3033 -10980 -2821 -10460
rect -279 -10593 -217 -5487
rect -129 -10593 -67 -5487
rect 2581 -5620 2793 -5100
rect 5335 -5233 5397 -127
rect 5485 -5233 5547 -127
rect 8195 -260 8407 260
rect 10949 127 11011 5233
rect 11099 127 11161 5233
rect 13809 5100 14021 5620
rect 16563 5487 16625 10593
rect 16713 5487 16775 10593
rect 19423 10460 19635 10980
rect 22177 10847 22239 15953
rect 22327 10847 22389 15953
rect 22177 10593 22389 10847
rect 16563 5233 16775 5487
rect 10949 -127 11161 127
rect 5335 -5487 5547 -5233
rect -279 -10847 -67 -10593
rect -5893 -16207 -5681 -15953
rect -11507 -21440 -11295 -21313
rect -8647 -21440 -8435 -21180
rect -5893 -21313 -5831 -16207
rect -5743 -21313 -5681 -16207
rect -3033 -16340 -2821 -15820
rect -279 -15953 -217 -10847
rect -129 -15953 -67 -10847
rect 2581 -10980 2793 -10460
rect 5335 -10593 5397 -5487
rect 5485 -10593 5547 -5487
rect 8195 -5620 8407 -5100
rect 10949 -5233 11011 -127
rect 11099 -5233 11161 -127
rect 13809 -260 14021 260
rect 16563 127 16625 5233
rect 16713 127 16775 5233
rect 19423 5100 19635 5620
rect 22177 5487 22239 10593
rect 22327 5487 22389 10593
rect 22177 5233 22389 5487
rect 16563 -127 16775 127
rect 10949 -5487 11161 -5233
rect 5335 -10847 5547 -10593
rect -279 -16207 -67 -15953
rect -5893 -21440 -5681 -21313
rect -3033 -21440 -2821 -21180
rect -279 -21313 -217 -16207
rect -129 -21313 -67 -16207
rect 2581 -16340 2793 -15820
rect 5335 -15953 5397 -10847
rect 5485 -15953 5547 -10847
rect 8195 -10980 8407 -10460
rect 10949 -10593 11011 -5487
rect 11099 -10593 11161 -5487
rect 13809 -5620 14021 -5100
rect 16563 -5233 16625 -127
rect 16713 -5233 16775 -127
rect 19423 -260 19635 260
rect 22177 127 22239 5233
rect 22327 127 22389 5233
rect 22177 -127 22389 127
rect 16563 -5487 16775 -5233
rect 10949 -10847 11161 -10593
rect 5335 -16207 5547 -15953
rect -279 -21440 -67 -21313
rect 2581 -21440 2793 -21180
rect 5335 -21313 5397 -16207
rect 5485 -21313 5547 -16207
rect 8195 -16340 8407 -15820
rect 10949 -15953 11011 -10847
rect 11099 -15953 11161 -10847
rect 13809 -10980 14021 -10460
rect 16563 -10593 16625 -5487
rect 16713 -10593 16775 -5487
rect 19423 -5620 19635 -5100
rect 22177 -5233 22239 -127
rect 22327 -5233 22389 -127
rect 22177 -5487 22389 -5233
rect 16563 -10847 16775 -10593
rect 10949 -16207 11161 -15953
rect 5335 -21440 5547 -21313
rect 8195 -21440 8407 -21180
rect 10949 -21313 11011 -16207
rect 11099 -21313 11161 -16207
rect 13809 -16340 14021 -15820
rect 16563 -15953 16625 -10847
rect 16713 -15953 16775 -10847
rect 19423 -10980 19635 -10460
rect 22177 -10593 22239 -5487
rect 22327 -10593 22389 -5487
rect 22177 -10847 22389 -10593
rect 16563 -16207 16775 -15953
rect 10949 -21440 11161 -21313
rect 13809 -21440 14021 -21180
rect 16563 -21313 16625 -16207
rect 16713 -21313 16775 -16207
rect 19423 -16340 19635 -15820
rect 22177 -15953 22239 -10847
rect 22327 -15953 22389 -10847
rect 22177 -16207 22389 -15953
rect 16563 -21440 16775 -21313
rect 19423 -21440 19635 -21180
rect 22177 -21313 22239 -16207
rect 22327 -21313 22389 -16207
rect 22177 -21440 22389 -21313
<< properties >>
string FIXED_BBOX 16909 16140 22149 21380
string gencell mim_2p0fF
string library gf180mcu
string parameters w 25 l 25 val 17.625k carea 25.00 cperi 20.00 nx 8 ny 8 dummy 0 square 0 lmin 5.00 wmin 5.00 lmax 100.0 wmax 100.0 dc 0 bconnect 1 tconnect 1
<< end >>
