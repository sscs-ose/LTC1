magic
tech gf180mcuC
magscale 1 10
timestamp 1714126980
<< error_p >>
rect -431 70 -385 166
rect -227 70 -181 166
rect -23 70 23 166
rect 181 70 227 166
rect 385 70 431 166
rect -431 -166 -385 -70
rect -227 -166 -181 -70
rect -23 -166 23 -70
rect 181 -166 227 -70
rect 385 -166 431 -70
<< nwell >>
rect -530 -298 530 298
<< pmos >>
rect -356 68 -256 168
rect -152 68 -52 168
rect 52 68 152 168
rect 256 68 356 168
rect -356 -168 -256 -68
rect -152 -168 -52 -68
rect 52 -168 152 -68
rect 256 -168 356 -68
<< pdiff >>
rect -444 155 -356 168
rect -444 81 -431 155
rect -385 81 -356 155
rect -444 68 -356 81
rect -256 155 -152 168
rect -256 81 -227 155
rect -181 81 -152 155
rect -256 68 -152 81
rect -52 155 52 168
rect -52 81 -23 155
rect 23 81 52 155
rect -52 68 52 81
rect 152 155 256 168
rect 152 81 181 155
rect 227 81 256 155
rect 152 68 256 81
rect 356 155 444 168
rect 356 81 385 155
rect 431 81 444 155
rect 356 68 444 81
rect -444 -81 -356 -68
rect -444 -155 -431 -81
rect -385 -155 -356 -81
rect -444 -168 -356 -155
rect -256 -81 -152 -68
rect -256 -155 -227 -81
rect -181 -155 -152 -81
rect -256 -168 -152 -155
rect -52 -81 52 -68
rect -52 -155 -23 -81
rect 23 -155 52 -81
rect -52 -168 52 -155
rect 152 -81 256 -68
rect 152 -155 181 -81
rect 227 -155 256 -81
rect 152 -168 256 -155
rect 356 -81 444 -68
rect 356 -155 385 -81
rect 431 -155 444 -81
rect 356 -168 444 -155
<< pdiffc >>
rect -431 81 -385 155
rect -227 81 -181 155
rect -23 81 23 155
rect 181 81 227 155
rect 385 81 431 155
rect -431 -155 -385 -81
rect -227 -155 -181 -81
rect -23 -155 23 -81
rect 181 -155 227 -81
rect 385 -155 431 -81
<< polysilicon >>
rect -356 168 -256 212
rect -152 168 -52 212
rect 52 168 152 212
rect 256 168 356 212
rect -356 24 -256 68
rect -152 24 -52 68
rect 52 24 152 68
rect 256 24 356 68
rect -356 -68 -256 -24
rect -152 -68 -52 -24
rect 52 -68 152 -24
rect 256 -68 356 -24
rect -356 -212 -256 -168
rect -152 -212 -52 -168
rect 52 -212 152 -168
rect 256 -212 356 -168
<< metal1 >>
rect -431 155 -385 166
rect -431 70 -385 81
rect -227 155 -181 166
rect -227 70 -181 81
rect -23 155 23 166
rect -23 70 23 81
rect 181 155 227 166
rect 181 70 227 81
rect 385 155 431 166
rect 385 70 431 81
rect -431 -81 -385 -70
rect -431 -166 -385 -155
rect -227 -81 -181 -70
rect -227 -166 -181 -155
rect -23 -81 23 -70
rect -23 -166 23 -155
rect 181 -81 227 -70
rect 181 -166 227 -155
rect 385 -81 431 -70
rect 385 -166 431 -155
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 0.5 l 0.5 m 2 nf 4 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
