magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2045 -2421 2045 2421
<< psubdiff >>
rect -45 399 45 421
rect -45 -399 -23 399
rect 23 -399 45 399
rect -45 -421 45 -399
<< psubdiffcont >>
rect -23 -399 23 399
<< metal1 >>
rect -34 399 34 410
rect -34 -399 -23 399
rect 23 -399 34 399
rect -34 -410 34 -399
<< end >>
