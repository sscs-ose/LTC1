magic
tech gf180mcuC
magscale 1 10
timestamp 1694513024
<< nwell >>
rect -4304 -386 4304 386
<< nsubdiff >>
rect -4280 290 4280 362
rect -4280 -290 -4208 290
rect 4208 -290 4280 290
rect -4280 -362 4280 -290
<< polysilicon >>
rect -4120 189 -3880 202
rect -4120 143 -4107 189
rect -3893 143 -3880 189
rect -4120 100 -3880 143
rect -4120 -143 -3880 -100
rect -4120 -189 -4107 -143
rect -3893 -189 -3880 -143
rect -4120 -202 -3880 -189
rect -3800 189 -3560 202
rect -3800 143 -3787 189
rect -3573 143 -3560 189
rect -3800 100 -3560 143
rect -3800 -143 -3560 -100
rect -3800 -189 -3787 -143
rect -3573 -189 -3560 -143
rect -3800 -202 -3560 -189
rect -3480 189 -3240 202
rect -3480 143 -3467 189
rect -3253 143 -3240 189
rect -3480 100 -3240 143
rect -3480 -143 -3240 -100
rect -3480 -189 -3467 -143
rect -3253 -189 -3240 -143
rect -3480 -202 -3240 -189
rect -3160 189 -2920 202
rect -3160 143 -3147 189
rect -2933 143 -2920 189
rect -3160 100 -2920 143
rect -3160 -143 -2920 -100
rect -3160 -189 -3147 -143
rect -2933 -189 -2920 -143
rect -3160 -202 -2920 -189
rect -2840 189 -2600 202
rect -2840 143 -2827 189
rect -2613 143 -2600 189
rect -2840 100 -2600 143
rect -2840 -143 -2600 -100
rect -2840 -189 -2827 -143
rect -2613 -189 -2600 -143
rect -2840 -202 -2600 -189
rect -2520 189 -2280 202
rect -2520 143 -2507 189
rect -2293 143 -2280 189
rect -2520 100 -2280 143
rect -2520 -143 -2280 -100
rect -2520 -189 -2507 -143
rect -2293 -189 -2280 -143
rect -2520 -202 -2280 -189
rect -2200 189 -1960 202
rect -2200 143 -2187 189
rect -1973 143 -1960 189
rect -2200 100 -1960 143
rect -2200 -143 -1960 -100
rect -2200 -189 -2187 -143
rect -1973 -189 -1960 -143
rect -2200 -202 -1960 -189
rect -1880 189 -1640 202
rect -1880 143 -1867 189
rect -1653 143 -1640 189
rect -1880 100 -1640 143
rect -1880 -143 -1640 -100
rect -1880 -189 -1867 -143
rect -1653 -189 -1640 -143
rect -1880 -202 -1640 -189
rect -1560 189 -1320 202
rect -1560 143 -1547 189
rect -1333 143 -1320 189
rect -1560 100 -1320 143
rect -1560 -143 -1320 -100
rect -1560 -189 -1547 -143
rect -1333 -189 -1320 -143
rect -1560 -202 -1320 -189
rect -1240 189 -1000 202
rect -1240 143 -1227 189
rect -1013 143 -1000 189
rect -1240 100 -1000 143
rect -1240 -143 -1000 -100
rect -1240 -189 -1227 -143
rect -1013 -189 -1000 -143
rect -1240 -202 -1000 -189
rect -920 189 -680 202
rect -920 143 -907 189
rect -693 143 -680 189
rect -920 100 -680 143
rect -920 -143 -680 -100
rect -920 -189 -907 -143
rect -693 -189 -680 -143
rect -920 -202 -680 -189
rect -600 189 -360 202
rect -600 143 -587 189
rect -373 143 -360 189
rect -600 100 -360 143
rect -600 -143 -360 -100
rect -600 -189 -587 -143
rect -373 -189 -360 -143
rect -600 -202 -360 -189
rect -280 189 -40 202
rect -280 143 -267 189
rect -53 143 -40 189
rect -280 100 -40 143
rect -280 -143 -40 -100
rect -280 -189 -267 -143
rect -53 -189 -40 -143
rect -280 -202 -40 -189
rect 40 189 280 202
rect 40 143 53 189
rect 267 143 280 189
rect 40 100 280 143
rect 40 -143 280 -100
rect 40 -189 53 -143
rect 267 -189 280 -143
rect 40 -202 280 -189
rect 360 189 600 202
rect 360 143 373 189
rect 587 143 600 189
rect 360 100 600 143
rect 360 -143 600 -100
rect 360 -189 373 -143
rect 587 -189 600 -143
rect 360 -202 600 -189
rect 680 189 920 202
rect 680 143 693 189
rect 907 143 920 189
rect 680 100 920 143
rect 680 -143 920 -100
rect 680 -189 693 -143
rect 907 -189 920 -143
rect 680 -202 920 -189
rect 1000 189 1240 202
rect 1000 143 1013 189
rect 1227 143 1240 189
rect 1000 100 1240 143
rect 1000 -143 1240 -100
rect 1000 -189 1013 -143
rect 1227 -189 1240 -143
rect 1000 -202 1240 -189
rect 1320 189 1560 202
rect 1320 143 1333 189
rect 1547 143 1560 189
rect 1320 100 1560 143
rect 1320 -143 1560 -100
rect 1320 -189 1333 -143
rect 1547 -189 1560 -143
rect 1320 -202 1560 -189
rect 1640 189 1880 202
rect 1640 143 1653 189
rect 1867 143 1880 189
rect 1640 100 1880 143
rect 1640 -143 1880 -100
rect 1640 -189 1653 -143
rect 1867 -189 1880 -143
rect 1640 -202 1880 -189
rect 1960 189 2200 202
rect 1960 143 1973 189
rect 2187 143 2200 189
rect 1960 100 2200 143
rect 1960 -143 2200 -100
rect 1960 -189 1973 -143
rect 2187 -189 2200 -143
rect 1960 -202 2200 -189
rect 2280 189 2520 202
rect 2280 143 2293 189
rect 2507 143 2520 189
rect 2280 100 2520 143
rect 2280 -143 2520 -100
rect 2280 -189 2293 -143
rect 2507 -189 2520 -143
rect 2280 -202 2520 -189
rect 2600 189 2840 202
rect 2600 143 2613 189
rect 2827 143 2840 189
rect 2600 100 2840 143
rect 2600 -143 2840 -100
rect 2600 -189 2613 -143
rect 2827 -189 2840 -143
rect 2600 -202 2840 -189
rect 2920 189 3160 202
rect 2920 143 2933 189
rect 3147 143 3160 189
rect 2920 100 3160 143
rect 2920 -143 3160 -100
rect 2920 -189 2933 -143
rect 3147 -189 3160 -143
rect 2920 -202 3160 -189
rect 3240 189 3480 202
rect 3240 143 3253 189
rect 3467 143 3480 189
rect 3240 100 3480 143
rect 3240 -143 3480 -100
rect 3240 -189 3253 -143
rect 3467 -189 3480 -143
rect 3240 -202 3480 -189
rect 3560 189 3800 202
rect 3560 143 3573 189
rect 3787 143 3800 189
rect 3560 100 3800 143
rect 3560 -143 3800 -100
rect 3560 -189 3573 -143
rect 3787 -189 3800 -143
rect 3560 -202 3800 -189
rect 3880 189 4120 202
rect 3880 143 3893 189
rect 4107 143 4120 189
rect 3880 100 4120 143
rect 3880 -143 4120 -100
rect 3880 -189 3893 -143
rect 4107 -189 4120 -143
rect 3880 -202 4120 -189
<< polycontact >>
rect -4107 143 -3893 189
rect -4107 -189 -3893 -143
rect -3787 143 -3573 189
rect -3787 -189 -3573 -143
rect -3467 143 -3253 189
rect -3467 -189 -3253 -143
rect -3147 143 -2933 189
rect -3147 -189 -2933 -143
rect -2827 143 -2613 189
rect -2827 -189 -2613 -143
rect -2507 143 -2293 189
rect -2507 -189 -2293 -143
rect -2187 143 -1973 189
rect -2187 -189 -1973 -143
rect -1867 143 -1653 189
rect -1867 -189 -1653 -143
rect -1547 143 -1333 189
rect -1547 -189 -1333 -143
rect -1227 143 -1013 189
rect -1227 -189 -1013 -143
rect -907 143 -693 189
rect -907 -189 -693 -143
rect -587 143 -373 189
rect -587 -189 -373 -143
rect -267 143 -53 189
rect -267 -189 -53 -143
rect 53 143 267 189
rect 53 -189 267 -143
rect 373 143 587 189
rect 373 -189 587 -143
rect 693 143 907 189
rect 693 -189 907 -143
rect 1013 143 1227 189
rect 1013 -189 1227 -143
rect 1333 143 1547 189
rect 1333 -189 1547 -143
rect 1653 143 1867 189
rect 1653 -189 1867 -143
rect 1973 143 2187 189
rect 1973 -189 2187 -143
rect 2293 143 2507 189
rect 2293 -189 2507 -143
rect 2613 143 2827 189
rect 2613 -189 2827 -143
rect 2933 143 3147 189
rect 2933 -189 3147 -143
rect 3253 143 3467 189
rect 3253 -189 3467 -143
rect 3573 143 3787 189
rect 3573 -189 3787 -143
rect 3893 143 4107 189
rect 3893 -189 4107 -143
<< ppolyres >>
rect -4120 -100 -3880 100
rect -3800 -100 -3560 100
rect -3480 -100 -3240 100
rect -3160 -100 -2920 100
rect -2840 -100 -2600 100
rect -2520 -100 -2280 100
rect -2200 -100 -1960 100
rect -1880 -100 -1640 100
rect -1560 -100 -1320 100
rect -1240 -100 -1000 100
rect -920 -100 -680 100
rect -600 -100 -360 100
rect -280 -100 -40 100
rect 40 -100 280 100
rect 360 -100 600 100
rect 680 -100 920 100
rect 1000 -100 1240 100
rect 1320 -100 1560 100
rect 1640 -100 1880 100
rect 1960 -100 2200 100
rect 2280 -100 2520 100
rect 2600 -100 2840 100
rect 2920 -100 3160 100
rect 3240 -100 3480 100
rect 3560 -100 3800 100
rect 3880 -100 4120 100
<< metal1 >>
rect -4118 143 -4107 189
rect -3893 143 -3882 189
rect -3798 143 -3787 189
rect -3573 143 -3562 189
rect -3478 143 -3467 189
rect -3253 143 -3242 189
rect -3158 143 -3147 189
rect -2933 143 -2922 189
rect -2838 143 -2827 189
rect -2613 143 -2602 189
rect -2518 143 -2507 189
rect -2293 143 -2282 189
rect -2198 143 -2187 189
rect -1973 143 -1962 189
rect -1878 143 -1867 189
rect -1653 143 -1642 189
rect -1558 143 -1547 189
rect -1333 143 -1322 189
rect -1238 143 -1227 189
rect -1013 143 -1002 189
rect -918 143 -907 189
rect -693 143 -682 189
rect -598 143 -587 189
rect -373 143 -362 189
rect -278 143 -267 189
rect -53 143 -42 189
rect 42 143 53 189
rect 267 143 278 189
rect 362 143 373 189
rect 587 143 598 189
rect 682 143 693 189
rect 907 143 918 189
rect 1002 143 1013 189
rect 1227 143 1238 189
rect 1322 143 1333 189
rect 1547 143 1558 189
rect 1642 143 1653 189
rect 1867 143 1878 189
rect 1962 143 1973 189
rect 2187 143 2198 189
rect 2282 143 2293 189
rect 2507 143 2518 189
rect 2602 143 2613 189
rect 2827 143 2838 189
rect 2922 143 2933 189
rect 3147 143 3158 189
rect 3242 143 3253 189
rect 3467 143 3478 189
rect 3562 143 3573 189
rect 3787 143 3798 189
rect 3882 143 3893 189
rect 4107 143 4118 189
rect -4118 -189 -4107 -143
rect -3893 -189 -3882 -143
rect -3798 -189 -3787 -143
rect -3573 -189 -3562 -143
rect -3478 -189 -3467 -143
rect -3253 -189 -3242 -143
rect -3158 -189 -3147 -143
rect -2933 -189 -2922 -143
rect -2838 -189 -2827 -143
rect -2613 -189 -2602 -143
rect -2518 -189 -2507 -143
rect -2293 -189 -2282 -143
rect -2198 -189 -2187 -143
rect -1973 -189 -1962 -143
rect -1878 -189 -1867 -143
rect -1653 -189 -1642 -143
rect -1558 -189 -1547 -143
rect -1333 -189 -1322 -143
rect -1238 -189 -1227 -143
rect -1013 -189 -1002 -143
rect -918 -189 -907 -143
rect -693 -189 -682 -143
rect -598 -189 -587 -143
rect -373 -189 -362 -143
rect -278 -189 -267 -143
rect -53 -189 -42 -143
rect 42 -189 53 -143
rect 267 -189 278 -143
rect 362 -189 373 -143
rect 587 -189 598 -143
rect 682 -189 693 -143
rect 907 -189 918 -143
rect 1002 -189 1013 -143
rect 1227 -189 1238 -143
rect 1322 -189 1333 -143
rect 1547 -189 1558 -143
rect 1642 -189 1653 -143
rect 1867 -189 1878 -143
rect 1962 -189 1973 -143
rect 2187 -189 2198 -143
rect 2282 -189 2293 -143
rect 2507 -189 2518 -143
rect 2602 -189 2613 -143
rect 2827 -189 2838 -143
rect 2922 -189 2933 -143
rect 3147 -189 3158 -143
rect 3242 -189 3253 -143
rect 3467 -189 3478 -143
rect 3562 -189 3573 -143
rect 3787 -189 3798 -143
rect 3882 -189 3893 -143
rect 4107 -189 4118 -143
<< properties >>
string FIXED_BBOX -4244 -326 4244 326
string gencell ppolyf_u
string library gf180mcu
string parameters w 1.2 l 1.0 m 1 nx 26 wmin 0.80 lmin 1.00 rho 315 val 278.761 dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0
<< end >>
