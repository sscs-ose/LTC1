magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -7445 -2095 7445 2095
<< psubdiff >>
rect -5445 70 5445 95
rect -5445 -70 -5381 70
rect 5381 -70 5445 70
rect -5445 -95 5445 -70
<< psubdiffcont >>
rect -5381 -70 5381 70
<< metal1 >>
rect -5434 70 5434 84
rect -5434 -70 -5381 70
rect 5381 -70 5434 70
rect -5434 -84 5434 -70
<< end >>
