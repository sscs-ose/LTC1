magic
tech gf180mcuC
magscale 1 10
timestamp 1693893072
<< nwell >>
rect -110 3244 6662 3581
rect -110 2807 6662 3187
rect -110 2335 6662 2715
rect -110 2084 6663 2335
rect -110 1884 270 2084
rect 937 2012 1044 2084
rect 1761 2006 1868 2084
rect 2577 2008 2684 2084
rect 3396 2006 3503 2084
rect 4207 2006 4314 2084
rect 5030 2006 5137 2084
rect 5829 2012 5936 2084
rect -110 1704 6649 1884
rect -110 1577 6662 1704
rect -110 1504 6649 1577
rect -101 1294 6663 1331
rect -101 1201 270 1294
rect 364 1247 6663 1294
rect 364 1201 1425 1247
rect -101 1199 1348 1201
rect 1464 1199 6663 1247
rect -101 1197 6663 1199
rect -110 946 6663 1197
<< psubdiff >>
rect 0 4796 157 4816
rect 0 4678 18 4796
rect 135 4678 157 4796
rect 0 4660 157 4678
rect 230 4796 387 4816
rect 230 4678 248 4796
rect 365 4678 387 4796
rect 230 4660 387 4678
rect 460 4796 617 4816
rect 460 4678 478 4796
rect 595 4678 617 4796
rect 460 4660 617 4678
rect 690 4796 847 4816
rect 690 4678 708 4796
rect 825 4678 847 4796
rect 690 4660 847 4678
rect 920 4796 1077 4816
rect 920 4678 938 4796
rect 1055 4678 1077 4796
rect 920 4660 1077 4678
rect 1150 4796 1307 4816
rect 1150 4678 1168 4796
rect 1285 4678 1307 4796
rect 1150 4660 1307 4678
rect 1380 4796 1537 4816
rect 1380 4678 1398 4796
rect 1515 4678 1537 4796
rect 1380 4660 1537 4678
rect 1610 4796 1767 4816
rect 1610 4678 1628 4796
rect 1745 4678 1767 4796
rect 1610 4660 1767 4678
rect 1840 4796 1997 4816
rect 1840 4678 1858 4796
rect 1975 4678 1997 4796
rect 1840 4660 1997 4678
rect 2070 4796 2227 4816
rect 2070 4678 2088 4796
rect 2205 4678 2227 4796
rect 2070 4660 2227 4678
rect 2300 4796 2457 4816
rect 2300 4678 2318 4796
rect 2435 4678 2457 4796
rect 2300 4660 2457 4678
rect 2530 4796 2687 4816
rect 2530 4678 2548 4796
rect 2665 4678 2687 4796
rect 2530 4660 2687 4678
rect 2760 4796 2917 4816
rect 2760 4678 2778 4796
rect 2895 4678 2917 4796
rect 2760 4660 2917 4678
rect 2990 4796 3147 4816
rect 2990 4678 3008 4796
rect 3125 4678 3147 4796
rect 2990 4660 3147 4678
rect 3220 4796 3377 4816
rect 3220 4678 3238 4796
rect 3355 4678 3377 4796
rect 3220 4660 3377 4678
rect 3450 4796 3607 4816
rect 3450 4678 3468 4796
rect 3585 4678 3607 4796
rect 3450 4660 3607 4678
rect 3680 4796 3837 4816
rect 3680 4678 3698 4796
rect 3815 4678 3837 4796
rect 3680 4660 3837 4678
rect 3910 4796 4067 4816
rect 3910 4678 3928 4796
rect 4045 4678 4067 4796
rect 3910 4660 4067 4678
rect 4140 4796 4297 4816
rect 4140 4678 4158 4796
rect 4275 4678 4297 4796
rect 4140 4660 4297 4678
rect 4370 4796 4527 4816
rect 4370 4678 4388 4796
rect 4505 4678 4527 4796
rect 4370 4660 4527 4678
rect 4600 4796 4757 4816
rect 4600 4678 4618 4796
rect 4735 4678 4757 4796
rect 4600 4660 4757 4678
rect 4830 4796 4987 4816
rect 4830 4678 4848 4796
rect 4965 4678 4987 4796
rect 4830 4660 4987 4678
rect 5060 4796 5217 4816
rect 5060 4678 5078 4796
rect 5195 4678 5217 4796
rect 5060 4660 5217 4678
rect 5290 4796 5447 4816
rect 5290 4678 5308 4796
rect 5425 4678 5447 4796
rect 5290 4660 5447 4678
rect 5520 4796 5677 4816
rect 5520 4678 5538 4796
rect 5655 4678 5677 4796
rect 5520 4660 5677 4678
rect 5750 4796 5907 4816
rect 5750 4678 5768 4796
rect 5885 4678 5907 4796
rect 5750 4660 5907 4678
rect 5980 4796 6137 4816
rect 5980 4678 5998 4796
rect 6115 4678 6137 4796
rect 5980 4660 6137 4678
rect 6210 4796 6367 4816
rect 6210 4678 6228 4796
rect 6345 4678 6367 4796
rect 6210 4660 6367 4678
rect 6440 4796 6597 4816
rect 6440 4678 6458 4796
rect 6575 4678 6597 4796
rect 6440 4660 6597 4678
rect 0 3775 157 3795
rect 0 3657 18 3775
rect 135 3657 157 3775
rect 0 3639 157 3657
rect 230 3775 387 3795
rect 230 3657 248 3775
rect 365 3657 387 3775
rect 230 3639 387 3657
rect 460 3775 617 3795
rect 460 3657 478 3775
rect 595 3657 617 3775
rect 460 3639 617 3657
rect 690 3775 847 3795
rect 690 3657 708 3775
rect 825 3657 847 3775
rect 690 3639 847 3657
rect 920 3775 1077 3795
rect 920 3657 938 3775
rect 1055 3657 1077 3775
rect 920 3639 1077 3657
rect 1150 3775 1307 3795
rect 1150 3657 1168 3775
rect 1285 3657 1307 3775
rect 1150 3639 1307 3657
rect 1380 3775 1537 3795
rect 1380 3657 1398 3775
rect 1515 3657 1537 3775
rect 1380 3639 1537 3657
rect 1610 3775 1767 3795
rect 1610 3657 1628 3775
rect 1745 3657 1767 3775
rect 1610 3639 1767 3657
rect 1840 3775 1997 3795
rect 1840 3657 1858 3775
rect 1975 3657 1997 3775
rect 1840 3639 1997 3657
rect 2070 3775 2227 3795
rect 2070 3657 2088 3775
rect 2205 3657 2227 3775
rect 2070 3639 2227 3657
rect 2300 3775 2457 3795
rect 2300 3657 2318 3775
rect 2435 3657 2457 3775
rect 2300 3639 2457 3657
rect 2530 3775 2687 3795
rect 2530 3657 2548 3775
rect 2665 3657 2687 3775
rect 2530 3639 2687 3657
rect 2760 3775 2917 3795
rect 2760 3657 2778 3775
rect 2895 3657 2917 3775
rect 2760 3639 2917 3657
rect 2990 3775 3147 3795
rect 2990 3657 3008 3775
rect 3125 3657 3147 3775
rect 2990 3639 3147 3657
rect 3220 3775 3377 3795
rect 3220 3657 3238 3775
rect 3355 3657 3377 3775
rect 3220 3639 3377 3657
rect 3450 3775 3607 3795
rect 3450 3657 3468 3775
rect 3585 3657 3607 3775
rect 3450 3639 3607 3657
rect 3680 3775 3837 3795
rect 3680 3657 3698 3775
rect 3815 3657 3837 3775
rect 3680 3639 3837 3657
rect 3910 3775 4067 3795
rect 3910 3657 3928 3775
rect 4045 3657 4067 3775
rect 3910 3639 4067 3657
rect 4140 3775 4297 3795
rect 4140 3657 4158 3775
rect 4275 3657 4297 3775
rect 4140 3639 4297 3657
rect 4370 3775 4527 3795
rect 4370 3657 4388 3775
rect 4505 3657 4527 3775
rect 4370 3639 4527 3657
rect 4600 3775 4757 3795
rect 4600 3657 4618 3775
rect 4735 3657 4757 3775
rect 4600 3639 4757 3657
rect 4830 3775 4987 3795
rect 4830 3657 4848 3775
rect 4965 3657 4987 3775
rect 4830 3639 4987 3657
rect 5060 3775 5217 3795
rect 5060 3657 5078 3775
rect 5195 3657 5217 3775
rect 5060 3639 5217 3657
rect 5290 3775 5447 3795
rect 5290 3657 5308 3775
rect 5425 3657 5447 3775
rect 5290 3639 5447 3657
rect 5520 3775 5677 3795
rect 5520 3657 5538 3775
rect 5655 3657 5677 3775
rect 5520 3639 5677 3657
rect 5750 3775 5907 3795
rect 5750 3657 5768 3775
rect 5885 3657 5907 3775
rect 5750 3639 5907 3657
rect 5980 3775 6137 3795
rect 5980 3657 5998 3775
rect 6115 3657 6137 3775
rect 5980 3639 6137 3657
rect 6210 3775 6367 3795
rect 6210 3657 6228 3775
rect 6345 3657 6367 3775
rect 6210 3639 6367 3657
rect 6440 3775 6597 3795
rect 6440 3657 6458 3775
rect 6575 3657 6597 3775
rect 6440 3639 6597 3657
rect 0 878 157 898
rect 0 760 18 878
rect 135 760 157 878
rect 0 742 157 760
rect 230 878 387 898
rect 230 760 248 878
rect 365 760 387 878
rect 230 742 387 760
rect 460 878 617 898
rect 460 760 478 878
rect 595 760 617 878
rect 460 742 617 760
rect 690 878 847 898
rect 690 760 708 878
rect 825 760 847 878
rect 690 742 847 760
rect 920 878 1077 898
rect 920 760 938 878
rect 1055 760 1077 878
rect 920 742 1077 760
rect 1150 878 1307 898
rect 1150 760 1168 878
rect 1285 760 1307 878
rect 1150 742 1307 760
rect 1380 878 1537 898
rect 1380 760 1398 878
rect 1515 760 1537 878
rect 1380 742 1537 760
rect 1610 878 1767 898
rect 1610 760 1628 878
rect 1745 760 1767 878
rect 1610 742 1767 760
rect 1840 878 1997 898
rect 1840 760 1858 878
rect 1975 760 1997 878
rect 1840 742 1997 760
rect 2070 878 2227 898
rect 2070 760 2088 878
rect 2205 760 2227 878
rect 2070 742 2227 760
rect 2300 878 2457 898
rect 2300 760 2318 878
rect 2435 760 2457 878
rect 2300 742 2457 760
rect 2530 878 2687 898
rect 2530 760 2548 878
rect 2665 760 2687 878
rect 2530 742 2687 760
rect 2760 878 2917 898
rect 2760 760 2778 878
rect 2895 760 2917 878
rect 2760 742 2917 760
rect 2990 878 3147 898
rect 2990 760 3008 878
rect 3125 760 3147 878
rect 2990 742 3147 760
rect 3220 878 3377 898
rect 3220 760 3238 878
rect 3355 760 3377 878
rect 3220 742 3377 760
rect 3450 878 3607 898
rect 3450 760 3468 878
rect 3585 760 3607 878
rect 3450 742 3607 760
rect 3680 878 3837 898
rect 3680 760 3698 878
rect 3815 760 3837 878
rect 3680 742 3837 760
rect 3910 878 4067 898
rect 3910 760 3928 878
rect 4045 760 4067 878
rect 3910 742 4067 760
rect 4140 878 4297 898
rect 4140 760 4158 878
rect 4275 760 4297 878
rect 4140 742 4297 760
rect 4370 878 4527 898
rect 4370 760 4388 878
rect 4505 760 4527 878
rect 4370 742 4527 760
rect 4600 878 4757 898
rect 4600 760 4618 878
rect 4735 760 4757 878
rect 4600 742 4757 760
rect 4830 878 4987 898
rect 4830 760 4848 878
rect 4965 760 4987 878
rect 4830 742 4987 760
rect 5060 878 5217 898
rect 5060 760 5078 878
rect 5195 760 5217 878
rect 5060 742 5217 760
rect 5290 878 5447 898
rect 5290 760 5308 878
rect 5425 760 5447 878
rect 5290 742 5447 760
rect 5520 878 5677 898
rect 5520 760 5538 878
rect 5655 760 5677 878
rect 5520 742 5677 760
rect 5750 878 5907 898
rect 5750 760 5768 878
rect 5885 760 5907 878
rect 5750 742 5907 760
rect 5980 878 6137 898
rect 5980 760 5998 878
rect 6115 760 6137 878
rect 5980 742 6137 760
rect 6210 878 6367 898
rect 6210 760 6228 878
rect 6345 760 6367 878
rect 6210 742 6367 760
rect 6440 878 6597 898
rect 6440 760 6458 878
rect 6575 760 6597 878
rect 6440 742 6597 760
rect 8 -131 165 -111
rect 8 -249 26 -131
rect 143 -249 165 -131
rect 8 -267 165 -249
rect 238 -131 395 -111
rect 238 -249 256 -131
rect 373 -249 395 -131
rect 238 -267 395 -249
rect 468 -131 625 -111
rect 468 -249 486 -131
rect 603 -249 625 -131
rect 468 -267 625 -249
rect 698 -131 855 -111
rect 698 -249 716 -131
rect 833 -249 855 -131
rect 698 -267 855 -249
rect 928 -131 1085 -111
rect 928 -249 946 -131
rect 1063 -249 1085 -131
rect 928 -267 1085 -249
rect 1158 -131 1315 -111
rect 1158 -249 1176 -131
rect 1293 -249 1315 -131
rect 1158 -267 1315 -249
rect 1388 -131 1545 -111
rect 1388 -249 1406 -131
rect 1523 -249 1545 -131
rect 1388 -267 1545 -249
rect 1618 -131 1775 -111
rect 1618 -249 1636 -131
rect 1753 -249 1775 -131
rect 1618 -267 1775 -249
rect 1848 -131 2005 -111
rect 1848 -249 1866 -131
rect 1983 -249 2005 -131
rect 1848 -267 2005 -249
rect 2078 -131 2235 -111
rect 2078 -249 2096 -131
rect 2213 -249 2235 -131
rect 2078 -267 2235 -249
rect 2308 -131 2465 -111
rect 2308 -249 2326 -131
rect 2443 -249 2465 -131
rect 2308 -267 2465 -249
rect 2538 -131 2695 -111
rect 2538 -249 2556 -131
rect 2673 -249 2695 -131
rect 2538 -267 2695 -249
rect 2768 -131 2925 -111
rect 2768 -249 2786 -131
rect 2903 -249 2925 -131
rect 2768 -267 2925 -249
rect 2998 -131 3155 -111
rect 2998 -249 3016 -131
rect 3133 -249 3155 -131
rect 2998 -267 3155 -249
rect 3228 -131 3385 -111
rect 3228 -249 3246 -131
rect 3363 -249 3385 -131
rect 3228 -267 3385 -249
rect 3458 -131 3615 -111
rect 3458 -249 3476 -131
rect 3593 -249 3615 -131
rect 3458 -267 3615 -249
rect 3688 -131 3845 -111
rect 3688 -249 3706 -131
rect 3823 -249 3845 -131
rect 3688 -267 3845 -249
rect 3918 -131 4075 -111
rect 3918 -249 3936 -131
rect 4053 -249 4075 -131
rect 3918 -267 4075 -249
rect 4148 -131 4305 -111
rect 4148 -249 4166 -131
rect 4283 -249 4305 -131
rect 4148 -267 4305 -249
rect 4378 -131 4535 -111
rect 4378 -249 4396 -131
rect 4513 -249 4535 -131
rect 4378 -267 4535 -249
rect 4608 -131 4765 -111
rect 4608 -249 4626 -131
rect 4743 -249 4765 -131
rect 4608 -267 4765 -249
rect 4838 -131 4995 -111
rect 4838 -249 4856 -131
rect 4973 -249 4995 -131
rect 4838 -267 4995 -249
rect 5068 -131 5225 -111
rect 5068 -249 5086 -131
rect 5203 -249 5225 -131
rect 5068 -267 5225 -249
rect 5298 -131 5455 -111
rect 5298 -249 5316 -131
rect 5433 -249 5455 -131
rect 5298 -267 5455 -249
rect 5528 -131 5685 -111
rect 5528 -249 5546 -131
rect 5663 -249 5685 -131
rect 5528 -267 5685 -249
rect 5758 -131 5915 -111
rect 5758 -249 5776 -131
rect 5893 -249 5915 -131
rect 5758 -267 5915 -249
rect 5988 -131 6145 -111
rect 5988 -249 6006 -131
rect 6123 -249 6145 -131
rect 5988 -267 6145 -249
rect 6218 -131 6375 -111
rect 6218 -249 6236 -131
rect 6353 -249 6375 -131
rect 6218 -267 6375 -249
rect 6448 -131 6605 -111
rect 6448 -249 6466 -131
rect 6583 -249 6605 -131
rect 6448 -267 6605 -249
<< nsubdiff >>
rect -61 3533 107 3554
rect -61 3410 -38 3533
rect 87 3410 107 3533
rect -61 3387 107 3410
rect 169 3533 337 3554
rect 169 3410 192 3533
rect 317 3410 337 3533
rect 169 3387 337 3410
rect 399 3533 567 3554
rect 399 3410 422 3533
rect 547 3410 567 3533
rect 399 3387 567 3410
rect 629 3533 797 3554
rect 629 3410 652 3533
rect 777 3410 797 3533
rect 629 3387 797 3410
rect 859 3533 1027 3554
rect 859 3410 882 3533
rect 1007 3410 1027 3533
rect 859 3387 1027 3410
rect 1089 3533 1257 3554
rect 1089 3410 1112 3533
rect 1237 3410 1257 3533
rect 1089 3387 1257 3410
rect 1319 3533 1487 3554
rect 1319 3410 1342 3533
rect 1467 3410 1487 3533
rect 1319 3387 1487 3410
rect 1549 3533 1717 3554
rect 1549 3410 1572 3533
rect 1697 3410 1717 3533
rect 1549 3387 1717 3410
rect 1779 3533 1947 3554
rect 1779 3410 1802 3533
rect 1927 3410 1947 3533
rect 1779 3387 1947 3410
rect 2009 3533 2177 3554
rect 2009 3410 2032 3533
rect 2157 3410 2177 3533
rect 2009 3387 2177 3410
rect 2239 3533 2407 3554
rect 2239 3410 2262 3533
rect 2387 3410 2407 3533
rect 2239 3387 2407 3410
rect 2469 3533 2637 3554
rect 2469 3410 2492 3533
rect 2617 3410 2637 3533
rect 2469 3387 2637 3410
rect 2699 3533 2867 3554
rect 2699 3410 2722 3533
rect 2847 3410 2867 3533
rect 2699 3387 2867 3410
rect 2929 3533 3097 3554
rect 2929 3410 2952 3533
rect 3077 3410 3097 3533
rect 2929 3387 3097 3410
rect 3159 3533 3327 3554
rect 3159 3410 3182 3533
rect 3307 3410 3327 3533
rect 3159 3387 3327 3410
rect 3389 3533 3557 3554
rect 3389 3410 3412 3533
rect 3537 3410 3557 3533
rect 3389 3387 3557 3410
rect 3619 3533 3787 3554
rect 3619 3410 3642 3533
rect 3767 3410 3787 3533
rect 3619 3387 3787 3410
rect 3849 3533 4017 3554
rect 3849 3410 3872 3533
rect 3997 3410 4017 3533
rect 3849 3387 4017 3410
rect 4079 3533 4247 3554
rect 4079 3410 4102 3533
rect 4227 3410 4247 3533
rect 4079 3387 4247 3410
rect 4309 3533 4477 3554
rect 4309 3410 4332 3533
rect 4457 3410 4477 3533
rect 4309 3387 4477 3410
rect 4539 3533 4707 3554
rect 4539 3410 4562 3533
rect 4687 3410 4707 3533
rect 4539 3387 4707 3410
rect 4769 3533 4937 3554
rect 4769 3410 4792 3533
rect 4917 3410 4937 3533
rect 4769 3387 4937 3410
rect 4999 3533 5167 3554
rect 4999 3410 5022 3533
rect 5147 3410 5167 3533
rect 4999 3387 5167 3410
rect 5229 3533 5397 3554
rect 5229 3410 5252 3533
rect 5377 3410 5397 3533
rect 5229 3387 5397 3410
rect 5459 3533 5627 3554
rect 5459 3410 5482 3533
rect 5607 3410 5627 3533
rect 5459 3387 5627 3410
rect 5689 3533 5857 3554
rect 5689 3410 5712 3533
rect 5837 3410 5857 3533
rect 5689 3387 5857 3410
rect 5919 3533 6087 3554
rect 5919 3410 5942 3533
rect 6067 3410 6087 3533
rect 5919 3387 6087 3410
rect 6149 3533 6317 3554
rect 6149 3410 6172 3533
rect 6297 3410 6317 3533
rect 6149 3387 6317 3410
rect 6379 3533 6547 3554
rect 6379 3410 6402 3533
rect 6527 3410 6547 3533
rect 6379 3387 6547 3410
rect -61 2287 107 2308
rect -61 2164 -38 2287
rect 87 2164 107 2287
rect -61 2141 107 2164
rect 169 2287 337 2308
rect 169 2164 192 2287
rect 317 2164 337 2287
rect 169 2141 337 2164
rect 399 2287 567 2308
rect 399 2164 422 2287
rect 547 2164 567 2287
rect 399 2141 567 2164
rect 629 2287 797 2308
rect 629 2164 652 2287
rect 777 2164 797 2287
rect 629 2141 797 2164
rect 859 2287 1027 2308
rect 859 2164 882 2287
rect 1007 2164 1027 2287
rect 859 2141 1027 2164
rect 1089 2287 1257 2308
rect 1089 2164 1112 2287
rect 1237 2164 1257 2287
rect 1089 2141 1257 2164
rect 1319 2287 1487 2308
rect 1319 2164 1342 2287
rect 1467 2164 1487 2287
rect 1319 2141 1487 2164
rect 1549 2287 1717 2308
rect 1549 2164 1572 2287
rect 1697 2164 1717 2287
rect 1549 2141 1717 2164
rect 1779 2287 1947 2308
rect 1779 2164 1802 2287
rect 1927 2164 1947 2287
rect 1779 2141 1947 2164
rect 2009 2287 2177 2308
rect 2009 2164 2032 2287
rect 2157 2164 2177 2287
rect 2009 2141 2177 2164
rect 2239 2287 2407 2308
rect 2239 2164 2262 2287
rect 2387 2164 2407 2287
rect 2239 2141 2407 2164
rect 2469 2287 2637 2308
rect 2469 2164 2492 2287
rect 2617 2164 2637 2287
rect 2469 2141 2637 2164
rect 2699 2287 2867 2308
rect 2699 2164 2722 2287
rect 2847 2164 2867 2287
rect 2699 2141 2867 2164
rect 2929 2287 3097 2308
rect 2929 2164 2952 2287
rect 3077 2164 3097 2287
rect 2929 2141 3097 2164
rect 3159 2287 3327 2308
rect 3159 2164 3182 2287
rect 3307 2164 3327 2287
rect 3159 2141 3327 2164
rect 3389 2287 3557 2308
rect 3389 2164 3412 2287
rect 3537 2164 3557 2287
rect 3389 2141 3557 2164
rect 3619 2287 3787 2308
rect 3619 2164 3642 2287
rect 3767 2164 3787 2287
rect 3619 2141 3787 2164
rect 3849 2287 4017 2308
rect 3849 2164 3872 2287
rect 3997 2164 4017 2287
rect 3849 2141 4017 2164
rect 4079 2287 4247 2308
rect 4079 2164 4102 2287
rect 4227 2164 4247 2287
rect 4079 2141 4247 2164
rect 4309 2287 4477 2308
rect 4309 2164 4332 2287
rect 4457 2164 4477 2287
rect 4309 2141 4477 2164
rect 4539 2287 4707 2308
rect 4539 2164 4562 2287
rect 4687 2164 4707 2287
rect 4539 2141 4707 2164
rect 4769 2287 4937 2308
rect 4769 2164 4792 2287
rect 4917 2164 4937 2287
rect 4769 2141 4937 2164
rect 4999 2287 5167 2308
rect 4999 2164 5022 2287
rect 5147 2164 5167 2287
rect 4999 2141 5167 2164
rect 5229 2287 5397 2308
rect 5229 2164 5252 2287
rect 5377 2164 5397 2287
rect 5229 2141 5397 2164
rect 5459 2287 5627 2308
rect 5459 2164 5482 2287
rect 5607 2164 5627 2287
rect 5459 2141 5627 2164
rect 5689 2287 5857 2308
rect 5689 2164 5712 2287
rect 5837 2164 5857 2287
rect 5689 2141 5857 2164
rect 5919 2287 6087 2308
rect 5919 2164 5942 2287
rect 6067 2164 6087 2287
rect 5919 2141 6087 2164
rect 6149 2287 6317 2308
rect 6149 2164 6172 2287
rect 6297 2164 6317 2287
rect 6149 2141 6317 2164
rect 6379 2287 6547 2308
rect 6379 2164 6402 2287
rect 6527 2164 6547 2287
rect 6379 2141 6547 2164
rect -61 1134 107 1155
rect -61 1011 -38 1134
rect 87 1011 107 1134
rect -61 988 107 1011
rect 169 1134 337 1155
rect 169 1011 192 1134
rect 317 1011 337 1134
rect 169 988 337 1011
rect 399 1134 567 1155
rect 399 1011 422 1134
rect 547 1011 567 1134
rect 399 988 567 1011
rect 629 1134 797 1155
rect 629 1011 652 1134
rect 777 1011 797 1134
rect 629 988 797 1011
rect 859 1134 1027 1155
rect 859 1011 882 1134
rect 1007 1011 1027 1134
rect 859 988 1027 1011
rect 1089 1134 1257 1155
rect 1089 1011 1112 1134
rect 1237 1011 1257 1134
rect 1089 988 1257 1011
rect 1319 1134 1487 1155
rect 1319 1011 1342 1134
rect 1467 1011 1487 1134
rect 1319 988 1487 1011
rect 1549 1134 1717 1155
rect 1549 1011 1572 1134
rect 1697 1011 1717 1134
rect 1549 988 1717 1011
rect 1779 1134 1947 1155
rect 1779 1011 1802 1134
rect 1927 1011 1947 1134
rect 1779 988 1947 1011
rect 2009 1134 2177 1155
rect 2009 1011 2032 1134
rect 2157 1011 2177 1134
rect 2009 988 2177 1011
rect 2239 1134 2407 1155
rect 2239 1011 2262 1134
rect 2387 1011 2407 1134
rect 2239 988 2407 1011
rect 2469 1134 2637 1155
rect 2469 1011 2492 1134
rect 2617 1011 2637 1134
rect 2469 988 2637 1011
rect 2699 1134 2867 1155
rect 2699 1011 2722 1134
rect 2847 1011 2867 1134
rect 2699 988 2867 1011
rect 2929 1134 3097 1155
rect 2929 1011 2952 1134
rect 3077 1011 3097 1134
rect 2929 988 3097 1011
rect 3159 1134 3327 1155
rect 3159 1011 3182 1134
rect 3307 1011 3327 1134
rect 3159 988 3327 1011
rect 3389 1134 3557 1155
rect 3389 1011 3412 1134
rect 3537 1011 3557 1134
rect 3389 988 3557 1011
rect 3619 1134 3787 1155
rect 3619 1011 3642 1134
rect 3767 1011 3787 1134
rect 3619 988 3787 1011
rect 3849 1134 4017 1155
rect 3849 1011 3872 1134
rect 3997 1011 4017 1134
rect 3849 988 4017 1011
rect 4079 1134 4247 1155
rect 4079 1011 4102 1134
rect 4227 1011 4247 1134
rect 4079 988 4247 1011
rect 4309 1134 4477 1155
rect 4309 1011 4332 1134
rect 4457 1011 4477 1134
rect 4309 988 4477 1011
rect 4539 1134 4707 1155
rect 4539 1011 4562 1134
rect 4687 1011 4707 1134
rect 4539 988 4707 1011
rect 4769 1134 4937 1155
rect 4769 1011 4792 1134
rect 4917 1011 4937 1134
rect 4769 988 4937 1011
rect 4999 1134 5167 1155
rect 4999 1011 5022 1134
rect 5147 1011 5167 1134
rect 4999 988 5167 1011
rect 5229 1134 5397 1155
rect 5229 1011 5252 1134
rect 5377 1011 5397 1134
rect 5229 988 5397 1011
rect 5459 1134 5627 1155
rect 5459 1011 5482 1134
rect 5607 1011 5627 1134
rect 5459 988 5627 1011
rect 5689 1134 5857 1155
rect 5689 1011 5712 1134
rect 5837 1011 5857 1134
rect 5689 988 5857 1011
rect 5919 1134 6087 1155
rect 5919 1011 5942 1134
rect 6067 1011 6087 1134
rect 5919 988 6087 1011
rect 6149 1134 6317 1155
rect 6149 1011 6172 1134
rect 6297 1011 6317 1134
rect 6149 988 6317 1011
rect 6379 1134 6547 1155
rect 6379 1011 6402 1134
rect 6527 1011 6547 1134
rect 6379 988 6547 1011
<< psubdiffcont >>
rect 18 4678 135 4796
rect 248 4678 365 4796
rect 478 4678 595 4796
rect 708 4678 825 4796
rect 938 4678 1055 4796
rect 1168 4678 1285 4796
rect 1398 4678 1515 4796
rect 1628 4678 1745 4796
rect 1858 4678 1975 4796
rect 2088 4678 2205 4796
rect 2318 4678 2435 4796
rect 2548 4678 2665 4796
rect 2778 4678 2895 4796
rect 3008 4678 3125 4796
rect 3238 4678 3355 4796
rect 3468 4678 3585 4796
rect 3698 4678 3815 4796
rect 3928 4678 4045 4796
rect 4158 4678 4275 4796
rect 4388 4678 4505 4796
rect 4618 4678 4735 4796
rect 4848 4678 4965 4796
rect 5078 4678 5195 4796
rect 5308 4678 5425 4796
rect 5538 4678 5655 4796
rect 5768 4678 5885 4796
rect 5998 4678 6115 4796
rect 6228 4678 6345 4796
rect 6458 4678 6575 4796
rect 18 3657 135 3775
rect 248 3657 365 3775
rect 478 3657 595 3775
rect 708 3657 825 3775
rect 938 3657 1055 3775
rect 1168 3657 1285 3775
rect 1398 3657 1515 3775
rect 1628 3657 1745 3775
rect 1858 3657 1975 3775
rect 2088 3657 2205 3775
rect 2318 3657 2435 3775
rect 2548 3657 2665 3775
rect 2778 3657 2895 3775
rect 3008 3657 3125 3775
rect 3238 3657 3355 3775
rect 3468 3657 3585 3775
rect 3698 3657 3815 3775
rect 3928 3657 4045 3775
rect 4158 3657 4275 3775
rect 4388 3657 4505 3775
rect 4618 3657 4735 3775
rect 4848 3657 4965 3775
rect 5078 3657 5195 3775
rect 5308 3657 5425 3775
rect 5538 3657 5655 3775
rect 5768 3657 5885 3775
rect 5998 3657 6115 3775
rect 6228 3657 6345 3775
rect 6458 3657 6575 3775
rect 18 760 135 878
rect 248 760 365 878
rect 478 760 595 878
rect 708 760 825 878
rect 938 760 1055 878
rect 1168 760 1285 878
rect 1398 760 1515 878
rect 1628 760 1745 878
rect 1858 760 1975 878
rect 2088 760 2205 878
rect 2318 760 2435 878
rect 2548 760 2665 878
rect 2778 760 2895 878
rect 3008 760 3125 878
rect 3238 760 3355 878
rect 3468 760 3585 878
rect 3698 760 3815 878
rect 3928 760 4045 878
rect 4158 760 4275 878
rect 4388 760 4505 878
rect 4618 760 4735 878
rect 4848 760 4965 878
rect 5078 760 5195 878
rect 5308 760 5425 878
rect 5538 760 5655 878
rect 5768 760 5885 878
rect 5998 760 6115 878
rect 6228 760 6345 878
rect 6458 760 6575 878
rect 26 -249 143 -131
rect 256 -249 373 -131
rect 486 -249 603 -131
rect 716 -249 833 -131
rect 946 -249 1063 -131
rect 1176 -249 1293 -131
rect 1406 -249 1523 -131
rect 1636 -249 1753 -131
rect 1866 -249 1983 -131
rect 2096 -249 2213 -131
rect 2326 -249 2443 -131
rect 2556 -249 2673 -131
rect 2786 -249 2903 -131
rect 3016 -249 3133 -131
rect 3246 -249 3363 -131
rect 3476 -249 3593 -131
rect 3706 -249 3823 -131
rect 3936 -249 4053 -131
rect 4166 -249 4283 -131
rect 4396 -249 4513 -131
rect 4626 -249 4743 -131
rect 4856 -249 4973 -131
rect 5086 -249 5203 -131
rect 5316 -249 5433 -131
rect 5546 -249 5663 -131
rect 5776 -249 5893 -131
rect 6006 -249 6123 -131
rect 6236 -249 6353 -131
rect 6466 -249 6583 -131
<< nsubdiffcont >>
rect -38 3410 87 3533
rect 192 3410 317 3533
rect 422 3410 547 3533
rect 652 3410 777 3533
rect 882 3410 1007 3533
rect 1112 3410 1237 3533
rect 1342 3410 1467 3533
rect 1572 3410 1697 3533
rect 1802 3410 1927 3533
rect 2032 3410 2157 3533
rect 2262 3410 2387 3533
rect 2492 3410 2617 3533
rect 2722 3410 2847 3533
rect 2952 3410 3077 3533
rect 3182 3410 3307 3533
rect 3412 3410 3537 3533
rect 3642 3410 3767 3533
rect 3872 3410 3997 3533
rect 4102 3410 4227 3533
rect 4332 3410 4457 3533
rect 4562 3410 4687 3533
rect 4792 3410 4917 3533
rect 5022 3410 5147 3533
rect 5252 3410 5377 3533
rect 5482 3410 5607 3533
rect 5712 3410 5837 3533
rect 5942 3410 6067 3533
rect 6172 3410 6297 3533
rect 6402 3410 6527 3533
rect -38 2164 87 2287
rect 192 2164 317 2287
rect 422 2164 547 2287
rect 652 2164 777 2287
rect 882 2164 1007 2287
rect 1112 2164 1237 2287
rect 1342 2164 1467 2287
rect 1572 2164 1697 2287
rect 1802 2164 1927 2287
rect 2032 2164 2157 2287
rect 2262 2164 2387 2287
rect 2492 2164 2617 2287
rect 2722 2164 2847 2287
rect 2952 2164 3077 2287
rect 3182 2164 3307 2287
rect 3412 2164 3537 2287
rect 3642 2164 3767 2287
rect 3872 2164 3997 2287
rect 4102 2164 4227 2287
rect 4332 2164 4457 2287
rect 4562 2164 4687 2287
rect 4792 2164 4917 2287
rect 5022 2164 5147 2287
rect 5252 2164 5377 2287
rect 5482 2164 5607 2287
rect 5712 2164 5837 2287
rect 5942 2164 6067 2287
rect 6172 2164 6297 2287
rect 6402 2164 6527 2287
rect -38 1011 87 1134
rect 192 1011 317 1134
rect 422 1011 547 1134
rect 652 1011 777 1134
rect 882 1011 1007 1134
rect 1112 1011 1237 1134
rect 1342 1011 1467 1134
rect 1572 1011 1697 1134
rect 1802 1011 1927 1134
rect 2032 1011 2157 1134
rect 2262 1011 2387 1134
rect 2492 1011 2617 1134
rect 2722 1011 2847 1134
rect 2952 1011 3077 1134
rect 3182 1011 3307 1134
rect 3412 1011 3537 1134
rect 3642 1011 3767 1134
rect 3872 1011 3997 1134
rect 4102 1011 4227 1134
rect 4332 1011 4457 1134
rect 4562 1011 4687 1134
rect 4792 1011 4917 1134
rect 5022 1011 5147 1134
rect 5252 1011 5377 1134
rect 5482 1011 5607 1134
rect 5712 1011 5837 1134
rect 5942 1011 6067 1134
rect 6172 1011 6297 1134
rect 6402 1011 6527 1134
<< polysilicon >>
rect 112 4597 6536 4625
rect 112 4525 126 4597
rect 198 4589 738 4597
rect 198 4525 212 4589
rect 112 4511 212 4525
rect 724 4525 738 4589
rect 810 4589 1554 4597
rect 810 4525 824 4589
rect 724 4511 824 4525
rect 928 4518 1028 4589
rect 1540 4525 1554 4589
rect 1626 4589 2370 4597
rect 1626 4525 1640 4589
rect 1540 4511 1640 4525
rect 1744 4518 1844 4589
rect 2356 4525 2370 4589
rect 2442 4589 3186 4597
rect 2442 4525 2456 4589
rect 2356 4511 2456 4525
rect 2560 4518 2660 4589
rect 3172 4525 3186 4589
rect 3258 4589 4002 4597
rect 3258 4525 3272 4589
rect 3172 4511 3272 4525
rect 3376 4518 3476 4589
rect 3988 4525 4002 4589
rect 4074 4589 4818 4597
rect 4074 4525 4088 4589
rect 3988 4511 4088 4525
rect 4192 4518 4292 4589
rect 4804 4525 4818 4589
rect 4890 4589 5634 4597
rect 4890 4525 4904 4589
rect 4804 4511 4904 4525
rect 5008 4518 5108 4589
rect 5620 4525 5634 4589
rect 5706 4589 6450 4597
rect 5706 4525 5720 4589
rect 5620 4511 5720 4525
rect 5824 4518 5924 4589
rect 6436 4525 6450 4589
rect 6522 4525 6536 4597
rect 6436 4511 6536 4525
rect 316 4285 416 4310
rect 316 4235 330 4285
rect 112 4213 330 4235
rect 402 4235 416 4285
rect 520 4285 620 4310
rect 520 4235 534 4285
rect 402 4213 534 4235
rect 606 4235 620 4285
rect 1132 4292 1232 4310
rect 1132 4235 1146 4292
rect 606 4221 1146 4235
rect 606 4213 738 4221
rect 112 4199 738 4213
rect 112 4142 212 4199
rect 724 4149 738 4199
rect 810 4199 942 4221
rect 810 4149 824 4199
rect 724 4135 824 4149
rect 928 4149 942 4199
rect 1014 4220 1146 4221
rect 1218 4235 1232 4292
rect 1336 4301 1436 4315
rect 1336 4235 1350 4301
rect 1218 4229 1350 4235
rect 1422 4235 1436 4301
rect 1948 4285 2048 4310
rect 1948 4235 1962 4285
rect 1422 4229 1962 4235
rect 1218 4221 1962 4229
rect 1218 4220 1758 4221
rect 1014 4218 1758 4220
rect 1014 4199 1554 4218
rect 1014 4149 1028 4199
rect 928 4135 1028 4149
rect 1540 4146 1554 4199
rect 1626 4199 1758 4218
rect 1626 4146 1640 4199
rect 1540 4132 1640 4146
rect 1744 4149 1758 4199
rect 1830 4213 1962 4221
rect 2034 4235 2048 4285
rect 2152 4285 2252 4310
rect 2152 4235 2166 4285
rect 2034 4213 2166 4235
rect 2238 4235 2252 4285
rect 2764 4285 2864 4310
rect 2764 4235 2778 4285
rect 2238 4221 2778 4235
rect 2238 4213 2370 4221
rect 1830 4199 2370 4213
rect 1830 4149 1844 4199
rect 1744 4135 1844 4149
rect 2356 4149 2370 4199
rect 2442 4199 2574 4221
rect 2442 4149 2456 4199
rect 2356 4135 2456 4149
rect 2560 4149 2574 4199
rect 2646 4213 2778 4221
rect 2850 4235 2864 4285
rect 2968 4285 3068 4310
rect 2968 4235 2982 4285
rect 2850 4213 2982 4235
rect 3054 4235 3068 4285
rect 3580 4285 3680 4310
rect 3580 4235 3594 4285
rect 3054 4221 3594 4235
rect 3054 4213 3186 4221
rect 2646 4199 3186 4213
rect 2646 4149 2660 4199
rect 2560 4135 2660 4149
rect 3172 4149 3186 4199
rect 3258 4199 3390 4221
rect 3258 4149 3272 4199
rect 3172 4135 3272 4149
rect 3376 4149 3390 4199
rect 3462 4213 3594 4221
rect 3666 4235 3680 4285
rect 3784 4285 3884 4310
rect 3784 4235 3798 4285
rect 3666 4213 3798 4235
rect 3870 4235 3884 4285
rect 4396 4285 4496 4310
rect 4396 4235 4410 4285
rect 3870 4221 4410 4235
rect 3870 4213 4002 4221
rect 3462 4199 4002 4213
rect 3462 4149 3476 4199
rect 3376 4135 3476 4149
rect 3988 4149 4002 4199
rect 4074 4199 4206 4221
rect 4074 4149 4088 4199
rect 3988 4135 4088 4149
rect 4192 4149 4206 4199
rect 4278 4213 4410 4221
rect 4482 4235 4496 4285
rect 4600 4285 4700 4310
rect 4600 4235 4614 4285
rect 4482 4213 4614 4235
rect 4686 4235 4700 4285
rect 5212 4285 5312 4310
rect 5212 4235 5226 4285
rect 4686 4221 5226 4235
rect 4686 4213 4818 4221
rect 4278 4199 4818 4213
rect 4278 4149 4292 4199
rect 4192 4135 4292 4149
rect 4804 4149 4818 4199
rect 4890 4199 5022 4221
rect 4890 4149 4904 4199
rect 4804 4135 4904 4149
rect 5008 4149 5022 4199
rect 5094 4213 5226 4221
rect 5298 4235 5312 4285
rect 5416 4285 5516 4310
rect 5416 4235 5430 4285
rect 5298 4213 5430 4235
rect 5502 4235 5516 4285
rect 6028 4285 6128 4310
rect 6028 4235 6042 4285
rect 5502 4221 6042 4235
rect 5502 4213 5634 4221
rect 5094 4199 5634 4213
rect 5094 4149 5108 4199
rect 5008 4135 5108 4149
rect 5620 4149 5634 4199
rect 5706 4199 5838 4221
rect 5706 4149 5720 4199
rect 5620 4135 5720 4149
rect 5824 4149 5838 4199
rect 5910 4213 6042 4221
rect 6114 4235 6128 4285
rect 6232 4285 6332 4310
rect 6232 4235 6246 4285
rect 6114 4213 6246 4235
rect 6318 4235 6332 4285
rect 6318 4221 6536 4235
rect 6318 4213 6450 4221
rect 5910 4199 6450 4213
rect 5910 4149 5924 4199
rect 5824 4135 5924 4149
rect 6436 4149 6450 4199
rect 6522 4149 6536 4221
rect 6436 4135 6536 4149
rect 316 3932 416 3946
rect 316 3860 330 3932
rect 402 3882 416 3932
rect 520 3882 620 3934
rect 1132 3932 1232 3946
rect 1132 3882 1146 3932
rect 402 3860 1146 3882
rect 1218 3882 1232 3932
rect 1336 3882 1436 3934
rect 1948 3932 2048 3946
rect 1948 3882 1962 3932
rect 1218 3860 1962 3882
rect 2034 3882 2048 3932
rect 2152 3882 2252 3934
rect 2764 3932 2864 3946
rect 2764 3882 2778 3932
rect 2034 3860 2778 3882
rect 2850 3882 2864 3932
rect 2968 3882 3068 3934
rect 3580 3932 3680 3946
rect 3580 3882 3594 3932
rect 2850 3860 3594 3882
rect 3666 3882 3680 3932
rect 3784 3882 3884 3934
rect 4396 3932 4496 3946
rect 4396 3882 4410 3932
rect 3666 3860 4410 3882
rect 4482 3882 4496 3932
rect 4600 3882 4700 3934
rect 5212 3932 5312 3946
rect 5212 3882 5226 3932
rect 4482 3860 5226 3882
rect 5298 3882 5312 3932
rect 5416 3882 5516 3934
rect 6028 3882 6128 3934
rect 6232 3932 6332 3946
rect 6232 3882 6246 3932
rect 5298 3860 6246 3882
rect 6318 3860 6332 3932
rect 316 3846 6332 3860
rect 135 3330 217 3341
rect 64 3322 6488 3330
rect 64 3274 150 3322
rect 198 3292 6488 3322
rect 198 3274 217 3292
rect 64 3256 217 3274
rect 64 3244 164 3256
rect 676 3244 776 3292
rect 880 3244 980 3292
rect 1492 3244 1592 3292
rect 1696 3244 1796 3292
rect 2308 3244 2408 3292
rect 2512 3244 2612 3292
rect 3124 3244 3224 3292
rect 3328 3244 3428 3292
rect 3940 3244 4040 3292
rect 4144 3244 4244 3292
rect 4756 3244 4856 3292
rect 4960 3244 5060 3292
rect 5572 3244 5672 3292
rect 5776 3244 5876 3292
rect 6388 3244 6488 3292
rect -200 2840 -127 2845
rect 268 2840 368 3036
rect 472 2840 572 3036
rect 1084 2840 1184 3036
rect 1288 2840 1388 3036
rect 1900 2840 2000 3036
rect 2104 2840 2204 3036
rect 2716 2840 2816 3036
rect 2920 2840 3020 3036
rect 3532 2840 3632 3036
rect 3736 2840 3836 3036
rect 4348 2840 4448 3036
rect 4552 2840 4652 3036
rect 5164 2840 5264 3036
rect 5368 2840 5468 3036
rect 5980 2840 6080 3036
rect 6184 2840 6284 3036
rect -200 2829 6795 2840
rect -200 2781 -187 2829
rect -140 2827 6795 2829
rect -140 2781 6719 2827
rect -200 2769 6719 2781
rect 6775 2769 6795 2827
rect -200 2765 -127 2769
rect 64 2677 164 2769
rect 676 2677 776 2769
rect 880 2677 980 2769
rect 1492 2677 1592 2769
rect 1696 2677 1796 2769
rect 2308 2677 2408 2769
rect 2512 2677 2612 2769
rect 3124 2677 3224 2769
rect 3328 2677 3428 2769
rect 3940 2677 4040 2769
rect 4144 2677 4244 2769
rect 4756 2677 4856 2769
rect 4960 2677 5060 2769
rect 5572 2677 5672 2769
rect 5776 2677 5876 2769
rect 6388 2677 6488 2769
rect 6705 2755 6795 2769
rect 268 2492 368 2513
rect 212 2477 368 2492
rect 212 2418 226 2477
rect 280 2465 368 2477
rect 472 2465 572 2513
rect 1084 2465 1184 2513
rect 1288 2465 1388 2513
rect 1900 2465 2000 2513
rect 2104 2465 2204 2513
rect 2716 2465 2816 2513
rect 2920 2465 3020 2513
rect 3532 2465 3632 2513
rect 3736 2465 3836 2513
rect 4348 2465 4448 2513
rect 4552 2465 4652 2513
rect 5164 2465 5264 2513
rect 5368 2465 5468 2513
rect 5980 2465 6080 2513
rect 6184 2507 6284 2513
rect 6184 2480 6340 2507
rect 6184 2465 6276 2480
rect 280 2430 6276 2465
rect 6326 2430 6340 2480
rect 280 2427 6340 2430
rect 280 2418 296 2427
rect 212 2404 296 2418
rect 6255 2416 6340 2427
rect 133 2084 212 2095
rect 938 2084 1017 2094
rect 1762 2084 1841 2088
rect 2578 2084 2657 2090
rect 3397 2084 3476 2088
rect 4208 2084 4287 2088
rect 5031 2084 5110 2088
rect 5830 2084 5909 2094
rect 64 2082 6488 2084
rect 64 2027 146 2082
rect 195 2081 6488 2082
rect 195 2046 951 2081
rect 195 2027 212 2046
rect 64 2013 212 2027
rect 64 1984 164 2013
rect 676 1998 776 2046
rect 880 2026 951 2046
rect 1000 2077 5843 2081
rect 1000 2075 2591 2077
rect 1000 2046 1775 2075
rect 1000 2045 1044 2046
rect 1000 2026 1017 2045
rect 880 2012 1017 2026
rect 880 1998 980 2012
rect 1492 1998 1592 2046
rect 1696 2020 1775 2046
rect 1824 2046 2591 2075
rect 1824 2039 1868 2046
rect 1824 2020 1841 2039
rect 1696 2006 1841 2020
rect 1696 1998 1796 2006
rect 2308 1998 2408 2046
rect 2512 2022 2591 2046
rect 2640 2075 5843 2077
rect 2640 2046 3410 2075
rect 2640 2041 2684 2046
rect 2640 2022 2657 2041
rect 2512 2008 2657 2022
rect 2512 1998 2612 2008
rect 3124 1998 3224 2046
rect 3328 2020 3410 2046
rect 3459 2046 4221 2075
rect 3459 2039 3503 2046
rect 3459 2020 3476 2039
rect 3328 2006 3476 2020
rect 3328 1998 3428 2006
rect 3940 1998 4040 2046
rect 4144 2020 4221 2046
rect 4270 2046 5044 2075
rect 4270 2039 4314 2046
rect 4270 2020 4287 2039
rect 4144 2006 4287 2020
rect 4144 1998 4244 2006
rect 4756 1998 4856 2046
rect 4960 2020 5044 2046
rect 5093 2046 5843 2075
rect 5093 2039 5137 2046
rect 5093 2020 5110 2039
rect 4960 2006 5110 2020
rect 4960 1998 5060 2006
rect 5572 1998 5672 2046
rect 5776 2026 5843 2046
rect 5892 2046 6488 2081
rect 5892 2045 5936 2046
rect 5892 2026 5909 2045
rect 5776 2012 5909 2026
rect 5776 1998 5876 2012
rect 6388 1998 6488 2046
rect 268 1615 368 1790
rect 472 1615 572 1790
rect 1084 1615 1184 1790
rect 1288 1615 1388 1790
rect 1900 1615 2000 1790
rect 2104 1615 2204 1790
rect 2716 1615 2816 1790
rect 2920 1615 3020 1790
rect 3532 1615 3632 1790
rect 3736 1615 3836 1790
rect 4348 1615 4448 1790
rect 4552 1615 4652 1790
rect 5164 1615 5264 1790
rect 5368 1615 5468 1790
rect 5980 1615 6080 1790
rect 6184 1615 6284 1790
rect 64 1601 6488 1615
rect 64 1553 806 1601
rect 854 1553 1611 1601
rect 1659 1553 2434 1601
rect 2482 1553 3248 1601
rect 3296 1553 4070 1601
rect 4118 1553 4875 1601
rect 4923 1553 5682 1601
rect 5730 1553 6488 1601
rect 64 1539 6488 1553
rect 64 1447 164 1539
rect 676 1447 776 1539
rect 880 1447 980 1539
rect 1492 1447 1592 1539
rect 1696 1447 1796 1539
rect 2308 1447 2408 1539
rect 2512 1447 2612 1539
rect 3124 1447 3224 1539
rect 3328 1447 3428 1539
rect 3940 1447 4040 1539
rect 4144 1447 4244 1539
rect 4756 1447 4856 1539
rect 4960 1447 5060 1539
rect 5572 1447 5672 1539
rect 5776 1447 5876 1539
rect 6388 1447 6488 1539
rect 268 1235 368 1297
rect 2153 1283 2233 1284
rect 2977 1283 3057 1285
rect 3790 1283 3870 1285
rect 4607 1283 4687 1287
rect 5426 1283 5506 1287
rect 472 1282 572 1283
rect 472 1268 604 1282
rect 472 1235 538 1268
rect 268 1213 538 1235
rect 587 1249 604 1268
rect 587 1235 631 1249
rect 1084 1235 1184 1283
rect 1288 1282 1388 1283
rect 1288 1268 1425 1282
rect 1288 1235 1359 1268
rect 587 1213 1359 1235
rect 1408 1235 1425 1268
rect 1900 1235 2000 1283
rect 2104 1270 2233 1283
rect 2104 1235 2167 1270
rect 1408 1215 2167 1235
rect 2216 1251 2233 1270
rect 2216 1235 2260 1251
rect 2716 1235 2816 1283
rect 2920 1271 3057 1283
rect 2920 1235 2991 1271
rect 2216 1216 2991 1235
rect 3040 1252 3057 1271
rect 3040 1235 3084 1252
rect 3532 1235 3632 1283
rect 3736 1271 3870 1283
rect 3736 1235 3804 1271
rect 3040 1216 3804 1235
rect 3853 1252 3870 1271
rect 3853 1235 3897 1252
rect 4348 1235 4448 1283
rect 4552 1273 4687 1283
rect 4552 1235 4621 1273
rect 3853 1218 4621 1235
rect 4670 1254 4687 1273
rect 4670 1235 4714 1254
rect 5164 1235 5264 1283
rect 5368 1273 5506 1283
rect 5368 1235 5440 1273
rect 4670 1218 5440 1235
rect 5489 1254 5506 1273
rect 5489 1235 5533 1254
rect 5980 1235 6080 1283
rect 6184 1235 6284 1283
rect 5489 1218 6284 1235
rect 3853 1216 6284 1218
rect 2216 1215 6284 1216
rect 1408 1213 6284 1215
rect 268 1197 6284 1213
rect 112 681 6536 695
rect 112 609 126 681
rect 198 659 6536 681
rect 198 609 212 659
rect 112 588 212 609
rect 724 588 824 659
rect 928 588 1028 659
rect 1540 588 1640 659
rect 1744 588 1844 659
rect 2356 588 2456 659
rect 2560 588 2660 659
rect 3172 588 3272 659
rect 3376 588 3476 659
rect 3988 588 4088 659
rect 4192 588 4292 659
rect 4804 588 4904 659
rect 5008 588 5108 659
rect 5620 588 5720 659
rect 5824 588 5924 659
rect 6436 588 6536 659
rect 316 319 416 383
rect 520 319 620 383
rect 1132 319 1232 382
rect 1336 319 1436 382
rect 1948 319 2048 381
rect 2152 319 2252 380
rect 2764 319 2864 382
rect 2968 319 3068 381
rect 3580 319 3680 380
rect 3784 319 3884 381
rect 4396 319 4496 381
rect 4600 319 4700 381
rect 5212 319 5312 381
rect 5416 319 5516 381
rect 6028 319 6128 383
rect 6232 319 6332 381
rect -92 283 6536 319
rect -92 223 -56 283
rect -117 205 -37 223
rect -117 157 -103 205
rect -56 157 -37 205
rect 112 168 212 283
rect 724 168 824 283
rect 928 168 1028 283
rect 1540 168 1640 283
rect 1744 168 1844 283
rect 2356 168 2456 283
rect 2560 168 2660 283
rect 3172 168 3272 283
rect 3376 168 3476 283
rect 3988 168 4088 283
rect 4192 168 4292 283
rect 4804 168 4904 283
rect 5008 168 5108 283
rect 5620 168 5720 283
rect 5824 168 5924 283
rect 6436 168 6536 283
rect -117 140 -37 157
rect 316 22 416 36
rect 316 -50 330 22
rect 402 -28 416 22
rect 520 -28 620 28
rect 1132 -28 1232 28
rect 1336 -28 1436 28
rect 1948 -28 2048 27
rect 2152 -28 2252 28
rect 2764 -28 2864 26
rect 2968 -28 3068 26
rect 3580 -28 3680 24
rect 3784 -28 3884 24
rect 4396 -28 4496 27
rect 4600 -28 4700 27
rect 5212 -28 5312 27
rect 5416 -28 5516 26
rect 6028 -28 6128 27
rect 6232 -28 6332 28
rect 402 -50 6332 -28
rect 316 -64 6332 -50
<< polycontact >>
rect 126 4525 198 4597
rect 738 4525 810 4597
rect 1554 4525 1626 4597
rect 2370 4525 2442 4597
rect 3186 4525 3258 4597
rect 4002 4525 4074 4597
rect 4818 4525 4890 4597
rect 5634 4525 5706 4597
rect 6450 4525 6522 4597
rect 330 4213 402 4285
rect 534 4213 606 4285
rect 738 4149 810 4221
rect 942 4149 1014 4221
rect 1146 4220 1218 4292
rect 1350 4229 1422 4301
rect 1554 4146 1626 4218
rect 1758 4149 1830 4221
rect 1962 4213 2034 4285
rect 2166 4213 2238 4285
rect 2370 4149 2442 4221
rect 2574 4149 2646 4221
rect 2778 4213 2850 4285
rect 2982 4213 3054 4285
rect 3186 4149 3258 4221
rect 3390 4149 3462 4221
rect 3594 4213 3666 4285
rect 3798 4213 3870 4285
rect 4002 4149 4074 4221
rect 4206 4149 4278 4221
rect 4410 4213 4482 4285
rect 4614 4213 4686 4285
rect 4818 4149 4890 4221
rect 5022 4149 5094 4221
rect 5226 4213 5298 4285
rect 5430 4213 5502 4285
rect 5634 4149 5706 4221
rect 5838 4149 5910 4221
rect 6042 4213 6114 4285
rect 6246 4213 6318 4285
rect 6450 4149 6522 4221
rect 330 3860 402 3932
rect 1146 3860 1218 3932
rect 1962 3860 2034 3932
rect 2778 3860 2850 3932
rect 3594 3860 3666 3932
rect 4410 3860 4482 3932
rect 5226 3860 5298 3932
rect 6246 3860 6318 3932
rect 150 3274 198 3322
rect -187 2781 -140 2829
rect 6719 2769 6775 2827
rect 226 2418 280 2477
rect 6276 2430 6326 2480
rect 146 2027 195 2082
rect 951 2026 1000 2081
rect 1775 2020 1824 2075
rect 2591 2022 2640 2077
rect 3410 2020 3459 2075
rect 4221 2020 4270 2075
rect 5044 2020 5093 2075
rect 5843 2026 5892 2081
rect 806 1553 854 1601
rect 1611 1553 1659 1601
rect 2434 1553 2482 1601
rect 3248 1553 3296 1601
rect 4070 1553 4118 1601
rect 4875 1553 4923 1601
rect 5682 1553 5730 1601
rect 538 1213 587 1268
rect 1359 1213 1408 1268
rect 2167 1215 2216 1270
rect 2991 1216 3040 1271
rect 3804 1216 3853 1271
rect 4621 1218 4670 1273
rect 5440 1218 5489 1273
rect 126 609 198 681
rect -103 157 -56 205
rect 330 -50 402 22
<< metal1 >>
rect 0 4796 6655 4816
rect 0 4678 18 4796
rect 135 4678 248 4796
rect 365 4678 478 4796
rect 595 4678 708 4796
rect 825 4678 938 4796
rect 1055 4678 1168 4796
rect 1285 4678 1398 4796
rect 1515 4678 1628 4796
rect 1745 4678 1858 4796
rect 1975 4678 2088 4796
rect 2205 4678 2318 4796
rect 2435 4678 2548 4796
rect 2665 4678 2778 4796
rect 2895 4678 3008 4796
rect 3125 4678 3238 4796
rect 3355 4678 3468 4796
rect 3585 4678 3698 4796
rect 3815 4678 3928 4796
rect 4045 4678 4158 4796
rect 4275 4678 4388 4796
rect 4505 4678 4618 4796
rect 4735 4678 4848 4796
rect 4965 4678 5078 4796
rect 5195 4678 5308 4796
rect 5425 4678 5538 4796
rect 5655 4678 5768 4796
rect 5885 4678 5998 4796
rect 6115 4678 6228 4796
rect 6345 4678 6458 4796
rect 6575 4678 6655 4796
rect 0 4660 6655 4678
rect 117 4597 207 4606
rect 117 4593 126 4597
rect -328 4525 126 4593
rect 198 4525 207 4597
rect -328 4516 207 4525
rect -328 4482 160 4516
rect -328 3015 -217 4482
rect 37 4470 83 4482
rect 445 4472 491 4660
rect 729 4597 819 4606
rect 729 4525 738 4597
rect 810 4562 819 4597
rect 810 4525 899 4562
rect 729 4516 899 4525
rect 853 4470 899 4516
rect 1261 4472 1307 4660
rect 1545 4597 1635 4606
rect 1545 4525 1554 4597
rect 1626 4560 1635 4597
rect 1626 4525 1715 4560
rect 1545 4516 1715 4525
rect 1616 4514 1715 4516
rect 1669 4470 1715 4514
rect 2077 4472 2123 4660
rect 2361 4597 2451 4606
rect 2361 4525 2370 4597
rect 2442 4562 2451 4597
rect 2442 4525 2531 4562
rect 2361 4516 2531 4525
rect 2361 4515 2438 4516
rect 2485 4470 2531 4516
rect 2893 4472 2939 4660
rect 3177 4597 3267 4606
rect 3177 4525 3186 4597
rect 3258 4561 3267 4597
rect 3258 4525 3347 4561
rect 3177 4516 3347 4525
rect 3247 4515 3347 4516
rect 3301 4470 3347 4515
rect 3709 4472 3755 4660
rect 3993 4597 4083 4606
rect 3993 4525 4002 4597
rect 4074 4560 4083 4597
rect 4074 4525 4163 4560
rect 3993 4516 4163 4525
rect 4064 4514 4163 4516
rect 4117 4470 4163 4514
rect 4525 4472 4571 4660
rect 4809 4597 4899 4606
rect 4809 4525 4818 4597
rect 4890 4560 4899 4597
rect 4890 4525 4979 4560
rect 4809 4516 4979 4525
rect 4874 4514 4979 4516
rect 4933 4470 4979 4514
rect 5341 4472 5387 4660
rect 5625 4597 5715 4606
rect 5625 4525 5634 4597
rect 5706 4562 5715 4597
rect 5706 4525 5795 4562
rect 5625 4516 5795 4525
rect 5749 4470 5795 4516
rect 6157 4472 6203 4660
rect 6441 4603 6531 4606
rect 6441 4597 6929 4603
rect 6441 4525 6450 4597
rect 6522 4525 6929 4597
rect 6441 4516 6929 4525
rect 6504 4492 6929 4516
rect 6565 4470 6611 4492
rect 241 4294 287 4365
rect 649 4294 695 4356
rect 241 4285 411 4294
rect 241 4213 330 4285
rect 402 4273 411 4285
rect 525 4285 695 4294
rect 525 4273 534 4285
rect 402 4227 534 4273
rect 402 4213 411 4227
rect 241 4204 411 4213
rect 525 4213 534 4227
rect 606 4273 695 4285
rect 1057 4301 1103 4370
rect 1465 4310 1511 4370
rect 1341 4301 1511 4310
rect 1057 4292 1227 4301
rect 1057 4273 1146 4292
rect 606 4227 1146 4273
rect 606 4221 819 4227
rect 606 4213 738 4221
rect 525 4204 738 4213
rect 241 4096 287 4204
rect 649 4149 738 4204
rect 810 4149 819 4221
rect 649 4140 819 4149
rect 933 4221 1146 4227
rect 933 4149 942 4221
rect 1014 4220 1146 4221
rect 1218 4273 1227 4292
rect 1341 4273 1350 4301
rect 1218 4229 1350 4273
rect 1422 4273 1511 4301
rect 1873 4294 1919 4368
rect 2281 4294 2327 4365
rect 1873 4285 2043 4294
rect 1873 4273 1962 4285
rect 1422 4229 1962 4273
rect 1218 4227 1962 4229
rect 1218 4220 1227 4227
rect 1341 4220 1635 4227
rect 1014 4211 1227 4220
rect 1465 4218 1635 4220
rect 1014 4149 1103 4211
rect 933 4140 1103 4149
rect 649 4096 695 4140
rect 1057 4096 1103 4140
rect 1465 4146 1554 4218
rect 1626 4146 1635 4218
rect 1465 4137 1635 4146
rect 1749 4221 1962 4227
rect 1749 4149 1758 4221
rect 1830 4213 1962 4221
rect 2034 4273 2043 4285
rect 2157 4285 2327 4294
rect 2157 4273 2166 4285
rect 2034 4227 2166 4273
rect 2034 4213 2043 4227
rect 1830 4204 2043 4213
rect 2157 4213 2166 4227
rect 2238 4273 2327 4285
rect 2689 4294 2735 4364
rect 3097 4294 3143 4362
rect 2689 4285 2859 4294
rect 2689 4273 2778 4285
rect 2238 4227 2778 4273
rect 2238 4221 2451 4227
rect 2238 4213 2370 4221
rect 2157 4204 2370 4213
rect 1830 4149 1919 4204
rect 1749 4140 1919 4149
rect 1465 4096 1511 4137
rect 1873 4096 1919 4140
rect 2281 4149 2370 4204
rect 2442 4149 2451 4221
rect 2281 4140 2451 4149
rect 2565 4221 2778 4227
rect 2565 4149 2574 4221
rect 2646 4213 2778 4221
rect 2850 4273 2859 4285
rect 2973 4285 3143 4294
rect 2973 4273 2982 4285
rect 2850 4227 2982 4273
rect 2850 4213 2859 4227
rect 2646 4204 2859 4213
rect 2973 4213 2982 4227
rect 3054 4273 3143 4285
rect 3505 4294 3551 4369
rect 3913 4294 3959 4362
rect 3505 4285 3675 4294
rect 3505 4273 3594 4285
rect 3054 4227 3594 4273
rect 3054 4221 3267 4227
rect 3054 4213 3186 4221
rect 2973 4204 3186 4213
rect 2646 4149 2735 4204
rect 2565 4140 2735 4149
rect 2281 4096 2327 4140
rect 2689 4096 2735 4140
rect 3097 4149 3186 4204
rect 3258 4149 3267 4221
rect 3097 4140 3267 4149
rect 3381 4221 3594 4227
rect 3381 4149 3390 4221
rect 3462 4213 3594 4221
rect 3666 4273 3675 4285
rect 3789 4285 3959 4294
rect 3789 4273 3798 4285
rect 3666 4227 3798 4273
rect 3666 4213 3675 4227
rect 3462 4204 3675 4213
rect 3789 4213 3798 4227
rect 3870 4273 3959 4285
rect 4321 4294 4367 4362
rect 4729 4294 4775 4362
rect 4321 4285 4491 4294
rect 4321 4273 4410 4285
rect 3870 4227 4410 4273
rect 3870 4221 4083 4227
rect 3870 4213 4002 4221
rect 3789 4204 4002 4213
rect 3462 4149 3551 4204
rect 3381 4140 3551 4149
rect 3097 4096 3143 4140
rect 3505 4096 3551 4140
rect 3913 4149 4002 4204
rect 4074 4149 4083 4221
rect 3913 4140 4083 4149
rect 4197 4221 4410 4227
rect 4197 4149 4206 4221
rect 4278 4213 4410 4221
rect 4482 4273 4491 4285
rect 4605 4285 4775 4294
rect 4605 4273 4614 4285
rect 4482 4227 4614 4273
rect 4482 4213 4491 4227
rect 4278 4204 4491 4213
rect 4605 4213 4614 4227
rect 4686 4273 4775 4285
rect 5137 4294 5183 4364
rect 5545 4294 5591 4367
rect 5137 4285 5307 4294
rect 5137 4273 5226 4285
rect 4686 4227 5226 4273
rect 4686 4221 4899 4227
rect 4686 4213 4818 4221
rect 4605 4204 4818 4213
rect 4278 4149 4367 4204
rect 4197 4140 4367 4149
rect 3913 4096 3959 4140
rect 4321 4096 4367 4140
rect 4729 4149 4818 4204
rect 4890 4149 4899 4221
rect 4729 4140 4899 4149
rect 5013 4221 5226 4227
rect 5013 4149 5022 4221
rect 5094 4213 5226 4221
rect 5298 4273 5307 4285
rect 5421 4285 5591 4294
rect 5421 4273 5430 4285
rect 5298 4227 5430 4273
rect 5298 4213 5307 4227
rect 5094 4204 5307 4213
rect 5421 4213 5430 4227
rect 5502 4273 5591 4285
rect 5953 4294 5999 4364
rect 6361 4294 6407 4363
rect 5953 4285 6123 4294
rect 5953 4273 6042 4285
rect 5502 4227 6042 4273
rect 5502 4221 5715 4227
rect 5502 4213 5634 4221
rect 5421 4204 5634 4213
rect 5094 4149 5183 4204
rect 5013 4140 5183 4149
rect 4729 4096 4775 4140
rect 5137 4096 5183 4140
rect 5545 4149 5634 4204
rect 5706 4149 5715 4221
rect 5545 4140 5715 4149
rect 5829 4221 6042 4227
rect 5829 4149 5838 4221
rect 5910 4213 6042 4221
rect 6114 4273 6123 4285
rect 6237 4285 6407 4294
rect 6237 4273 6246 4285
rect 6114 4227 6246 4273
rect 6114 4213 6123 4227
rect 5910 4204 6123 4213
rect 6237 4213 6246 4227
rect 6318 4273 6407 4285
rect 6318 4230 6529 4273
rect 6318 4221 6531 4230
rect 6318 4213 6450 4221
rect 6237 4204 6450 4213
rect 5910 4149 5999 4204
rect 5829 4140 5999 4149
rect 5545 4096 5591 4140
rect 5953 4096 5999 4140
rect 6361 4149 6450 4204
rect 6522 4149 6531 4221
rect 6361 4140 6531 4149
rect 6361 4096 6407 4140
rect 37 3795 83 3990
rect 445 3943 491 3989
rect 367 3941 491 3943
rect 321 3932 491 3941
rect 321 3860 330 3932
rect 402 3897 491 3932
rect 402 3860 411 3897
rect 321 3851 411 3860
rect 853 3795 899 3991
rect 1261 3990 1306 3991
rect 1261 3947 1307 3990
rect 1196 3941 1307 3947
rect 1137 3932 1307 3941
rect 1137 3860 1146 3932
rect 1218 3894 1307 3932
rect 1218 3860 1227 3894
rect 1137 3851 1227 3860
rect 1669 3795 1715 3986
rect 2077 3945 2123 3993
rect 2002 3941 2123 3945
rect 1953 3932 2123 3941
rect 1953 3860 1962 3932
rect 2034 3899 2123 3932
rect 2034 3860 2043 3899
rect 1953 3851 2043 3860
rect 2485 3795 2531 3988
rect 2893 3949 2939 3993
rect 3709 3990 3754 3991
rect 2813 3941 2939 3949
rect 2769 3932 2939 3941
rect 2769 3860 2778 3932
rect 2850 3903 2939 3932
rect 2850 3860 2859 3903
rect 2769 3851 2859 3860
rect 3301 3795 3347 3987
rect 3709 3951 3755 3990
rect 3638 3941 3755 3951
rect 3585 3932 3755 3941
rect 3585 3860 3594 3932
rect 3666 3905 3755 3932
rect 3666 3860 3675 3905
rect 3585 3851 3675 3860
rect 4117 3795 4163 3981
rect 4525 3945 4571 3991
rect 4446 3941 4571 3945
rect 4401 3932 4571 3941
rect 4401 3860 4410 3932
rect 4482 3899 4571 3932
rect 4482 3860 4491 3899
rect 4401 3851 4491 3860
rect 4933 3795 4979 3986
rect 5341 3945 5387 3989
rect 5265 3941 5387 3945
rect 5217 3932 5387 3941
rect 5217 3860 5226 3932
rect 5298 3899 5387 3932
rect 5298 3860 5307 3899
rect 5217 3851 5307 3860
rect 5749 3795 5795 3981
rect 6157 3943 6203 3991
rect 6157 3941 6287 3943
rect 6157 3932 6327 3941
rect 6157 3897 6246 3932
rect 6237 3860 6246 3897
rect 6318 3860 6327 3932
rect 6237 3851 6327 3860
rect 6565 3795 6611 3983
rect 0 3775 6655 3795
rect 0 3657 18 3775
rect 135 3657 248 3775
rect 365 3657 478 3775
rect 595 3657 708 3775
rect 825 3657 938 3775
rect 1055 3657 1168 3775
rect 1285 3657 1398 3775
rect 1515 3657 1628 3775
rect 1745 3657 1858 3775
rect 1975 3657 2088 3775
rect 2205 3657 2318 3775
rect 2435 3657 2548 3775
rect 2665 3657 2778 3775
rect 2895 3657 3008 3775
rect 3125 3657 3238 3775
rect 3355 3657 3468 3775
rect 3585 3657 3698 3775
rect 3815 3657 3928 3775
rect 4045 3657 4158 3775
rect 4275 3657 4388 3775
rect 4505 3657 4618 3775
rect 4735 3657 4848 3775
rect 4965 3657 5078 3775
rect 5195 3657 5308 3775
rect 5425 3657 5538 3775
rect 5655 3657 5768 3775
rect 5885 3657 5998 3775
rect 6115 3657 6228 3775
rect 6345 3657 6458 3775
rect 6575 3657 6655 3775
rect 0 3639 6655 3657
rect -110 3533 6662 3581
rect -110 3410 -38 3533
rect 87 3410 192 3533
rect 317 3410 422 3533
rect 547 3410 652 3533
rect 777 3410 882 3533
rect 1007 3410 1112 3533
rect 1237 3410 1342 3533
rect 1467 3410 1572 3533
rect 1697 3410 1802 3533
rect 1927 3410 2032 3533
rect 2157 3410 2262 3533
rect 2387 3410 2492 3533
rect 2617 3410 2722 3533
rect 2847 3410 2952 3533
rect 3077 3410 3182 3533
rect 3307 3410 3412 3533
rect 3537 3410 3642 3533
rect 3767 3410 3872 3533
rect 3997 3410 4102 3533
rect 4227 3410 4332 3533
rect 4457 3410 4562 3533
rect 4687 3410 4792 3533
rect 4917 3410 5022 3533
rect 5147 3410 5252 3533
rect 5377 3410 5482 3533
rect 5607 3410 5712 3533
rect 5837 3410 5942 3533
rect 6067 3410 6172 3533
rect 6297 3410 6402 3533
rect 6527 3519 6662 3533
rect 6528 3463 6662 3519
rect 6527 3410 6662 3463
rect -110 3387 6662 3410
rect -11 3198 35 3387
rect 135 3328 217 3341
rect 135 3270 147 3328
rect 206 3270 217 3328
rect 135 3256 217 3270
rect 805 3198 851 3387
rect 1621 3198 1667 3387
rect 2437 3198 2483 3387
rect 3253 3198 3299 3387
rect 4069 3198 4115 3387
rect 4885 3198 4931 3387
rect 5701 3198 5747 3387
rect 6517 3198 6563 3387
rect 181 3171 258 3183
rect 181 3116 191 3171
rect 245 3116 258 3171
rect 181 3104 258 3116
rect 588 3171 665 3183
rect 588 3116 598 3171
rect 652 3116 665 3171
rect 588 3104 665 3116
rect 999 3167 1076 3179
rect 999 3112 1009 3167
rect 1063 3112 1076 3167
rect 999 3100 1076 3112
rect 1403 3168 1480 3180
rect 1403 3113 1413 3168
rect 1467 3113 1480 3168
rect 1403 3101 1480 3113
rect 1809 3166 1886 3178
rect 1809 3111 1819 3166
rect 1873 3111 1886 3166
rect 1809 3099 1886 3111
rect 2219 3168 2296 3180
rect 2219 3113 2229 3168
rect 2283 3113 2296 3168
rect 2219 3101 2296 3113
rect 2624 3165 2701 3177
rect 2624 3110 2634 3165
rect 2688 3110 2701 3165
rect 2624 3098 2701 3110
rect 3033 3165 3110 3177
rect 3033 3110 3043 3165
rect 3097 3110 3110 3165
rect 3033 3098 3110 3110
rect 3444 3165 3521 3177
rect 3444 3110 3454 3165
rect 3508 3110 3521 3165
rect 3444 3098 3521 3110
rect 3849 3165 3926 3177
rect 3849 3110 3859 3165
rect 3913 3110 3926 3165
rect 3849 3098 3926 3110
rect 4255 3167 4332 3179
rect 4255 3112 4265 3167
rect 4319 3112 4332 3167
rect 4255 3100 4332 3112
rect 4665 3169 4742 3181
rect 4665 3114 4675 3169
rect 4729 3114 4742 3169
rect 4665 3102 4742 3114
rect 5072 3166 5149 3178
rect 5072 3111 5082 3166
rect 5136 3111 5149 3166
rect 5072 3099 5149 3111
rect 5481 3166 5558 3178
rect 5481 3111 5491 3166
rect 5545 3111 5558 3166
rect 5481 3099 5558 3111
rect 5889 3168 5966 3180
rect 5889 3113 5899 3168
rect 5953 3113 5966 3168
rect 5889 3101 5966 3113
rect 6295 3171 6372 3183
rect 6295 3116 6305 3171
rect 6359 3116 6372 3171
rect 6295 3104 6372 3116
rect -328 2931 100 3015
rect 397 2931 443 3085
rect 1213 2931 1259 3089
rect 2029 2931 2075 3092
rect 2845 2931 2891 3086
rect 3661 2931 3707 3087
rect 4477 2931 4523 3085
rect 5293 2931 5339 3089
rect 6109 2931 6155 3087
rect 6818 3006 6929 4492
rect 6452 2931 6929 3006
rect -328 2904 6929 2931
rect -11 2895 6929 2904
rect -200 2840 -127 2845
rect -305 2829 -127 2840
rect -305 2781 -187 2829
rect -140 2781 -127 2829
rect -305 2765 -127 2781
rect -11 2820 6563 2895
rect -305 1414 -235 2765
rect -11 2675 35 2820
rect 805 2675 851 2820
rect 1621 2675 1667 2820
rect 177 2655 254 2667
rect 177 2600 187 2655
rect 241 2600 254 2655
rect 177 2588 254 2600
rect 588 2657 665 2669
rect 588 2602 598 2657
rect 652 2602 665 2657
rect 588 2590 665 2602
rect 991 2660 1068 2672
rect 991 2605 1001 2660
rect 1055 2605 1068 2660
rect 991 2593 1068 2605
rect 1401 2663 1478 2675
rect 1401 2608 1411 2663
rect 1465 2608 1478 2663
rect 1401 2596 1478 2608
rect 1808 2662 1885 2674
rect 1808 2607 1818 2662
rect 1872 2607 1885 2662
rect 1808 2595 1885 2607
rect 2215 2661 2292 2673
rect 2437 2672 2483 2820
rect 3253 2675 3299 2820
rect 4069 2675 4115 2820
rect 2215 2606 2225 2661
rect 2279 2606 2292 2661
rect 2215 2594 2292 2606
rect 2623 2659 2700 2671
rect 2623 2604 2633 2659
rect 2687 2604 2700 2659
rect 2623 2592 2700 2604
rect 3035 2657 3112 2669
rect 3035 2602 3045 2657
rect 3099 2602 3112 2657
rect 3035 2590 3112 2602
rect 3440 2660 3517 2672
rect 3440 2605 3450 2660
rect 3504 2605 3517 2660
rect 3440 2593 3517 2605
rect 3849 2659 3926 2671
rect 4885 2669 4931 2820
rect 5701 2675 5747 2820
rect 6517 2675 6563 2820
rect 6705 2827 6848 2840
rect 6705 2769 6719 2827
rect 6775 2769 6848 2827
rect 6705 2755 6848 2769
rect 3849 2604 3859 2659
rect 3913 2604 3926 2659
rect 3849 2592 3926 2604
rect 4257 2657 4334 2669
rect 4257 2602 4267 2657
rect 4321 2602 4334 2657
rect 4257 2590 4334 2602
rect 4665 2657 4742 2669
rect 4665 2602 4675 2657
rect 4729 2602 4742 2657
rect 4665 2590 4742 2602
rect 5072 2656 5149 2668
rect 5072 2601 5082 2656
rect 5136 2601 5149 2656
rect 5072 2589 5149 2601
rect 5480 2661 5557 2673
rect 5480 2606 5490 2661
rect 5544 2606 5557 2661
rect 5480 2594 5557 2606
rect 5887 2661 5964 2673
rect 5887 2606 5897 2661
rect 5951 2606 5964 2661
rect 5887 2594 5964 2606
rect 6297 2659 6374 2671
rect 6297 2604 6307 2659
rect 6361 2604 6374 2659
rect 6297 2592 6374 2604
rect 212 2477 296 2492
rect 212 2418 226 2477
rect 280 2418 296 2477
rect 212 2404 296 2418
rect 397 2335 443 2559
rect 1213 2335 1259 2576
rect 2029 2335 2075 2572
rect 2845 2335 2891 2573
rect 3661 2335 3707 2569
rect 4477 2335 4523 2572
rect 5293 2335 5339 2570
rect 6109 2335 6155 2560
rect 6255 2483 6340 2507
rect 6255 2427 6269 2483
rect 6325 2480 6340 2483
rect 6326 2430 6340 2480
rect 6325 2427 6340 2430
rect 6255 2416 6340 2427
rect -110 2287 6663 2335
rect -110 2164 -38 2287
rect 87 2271 192 2287
rect 87 2215 184 2271
rect 87 2164 192 2215
rect 317 2164 422 2287
rect 547 2164 652 2287
rect 777 2164 882 2287
rect 1007 2164 1112 2287
rect 1237 2164 1342 2287
rect 1467 2164 1572 2287
rect 1697 2164 1802 2287
rect 1927 2164 2032 2287
rect 2157 2164 2262 2287
rect 2387 2164 2492 2287
rect 2617 2164 2722 2287
rect 2847 2164 2952 2287
rect 3077 2164 3182 2287
rect 3307 2164 3412 2287
rect 3537 2164 3642 2287
rect 3767 2164 3872 2287
rect 3997 2164 4102 2287
rect 4227 2164 4332 2287
rect 4457 2164 4562 2287
rect 4687 2164 4792 2287
rect 4917 2164 5022 2287
rect 5147 2164 5252 2287
rect 5377 2164 5482 2287
rect 5607 2164 5712 2287
rect 5837 2164 5942 2287
rect 6067 2164 6172 2287
rect 6297 2164 6402 2287
rect 6527 2164 6663 2287
rect -110 2141 6663 2164
rect -11 1952 35 2141
rect 135 2082 239 2094
rect 135 2027 146 2082
rect 195 2027 239 2082
rect 135 2014 239 2027
rect 193 1769 239 2014
rect 805 1952 851 2141
rect 940 2082 1044 2093
rect 940 2025 949 2082
rect 1004 2079 1044 2082
rect 1004 2025 1055 2079
rect 940 2013 1055 2025
rect 998 2012 1055 2013
rect 380 1927 456 1940
rect 380 1871 391 1927
rect 446 1871 456 1927
rect 380 1860 456 1871
rect 601 1769 647 1836
rect 1009 1769 1055 2012
rect 1621 1952 1667 2141
rect 1764 2075 1868 2087
rect 1764 2020 1775 2075
rect 1824 2071 1868 2075
rect 1824 2020 1871 2071
rect 1764 2007 1871 2020
rect 1822 2006 1871 2007
rect 1196 1933 1272 1946
rect 1196 1877 1207 1933
rect 1262 1877 1272 1933
rect 1196 1866 1272 1877
rect 1417 1769 1463 1836
rect 1825 1769 1871 2006
rect 2437 1952 2483 2141
rect 2580 2077 2684 2089
rect 2580 2022 2591 2077
rect 2640 2076 2684 2077
rect 2640 2022 2687 2076
rect 2580 2009 2687 2022
rect 2638 2008 2687 2009
rect 2012 1926 2088 1939
rect 2012 1870 2023 1926
rect 2078 1870 2088 1926
rect 2012 1859 2088 1870
rect 2233 1769 2279 1836
rect 2641 1769 2687 2008
rect 3253 1952 3299 2141
rect 3399 2075 3503 2087
rect 3399 2020 3410 2075
rect 3459 2020 3503 2075
rect 3399 2007 3503 2020
rect 2826 1930 2902 1943
rect 2826 1874 2837 1930
rect 2892 1874 2902 1930
rect 2826 1863 2902 1874
rect 3049 1769 3095 1836
rect 3457 1769 3503 2007
rect 4069 1952 4115 2141
rect 4210 2075 4314 2087
rect 4210 2020 4221 2075
rect 4270 2056 4314 2075
rect 4270 2020 4319 2056
rect 4210 2007 4319 2020
rect 4268 2006 4319 2007
rect 3643 1925 3719 1938
rect 3643 1869 3654 1925
rect 3709 1869 3719 1925
rect 3643 1858 3719 1869
rect 3865 1769 3911 1836
rect 4273 1769 4319 2006
rect 4885 1952 4931 2141
rect 5033 2075 5137 2087
rect 5033 2020 5044 2075
rect 5093 2020 5137 2075
rect 5033 2007 5137 2020
rect 5089 2006 5137 2007
rect 4460 1928 4536 1941
rect 4460 1872 4471 1928
rect 4526 1872 4536 1928
rect 4460 1861 4536 1872
rect 4681 1769 4727 1836
rect 5089 1769 5135 2006
rect 5701 1952 5747 2141
rect 5832 2084 5936 2093
rect 5832 2030 5841 2084
rect 5895 2080 5936 2084
rect 5895 2030 5951 2080
rect 5832 2026 5843 2030
rect 5892 2026 5951 2030
rect 5832 2013 5951 2026
rect 5890 2012 5951 2013
rect 5276 1927 5352 1940
rect 5276 1871 5287 1927
rect 5342 1871 5352 1927
rect 5276 1860 5352 1871
rect 5497 1769 5543 1836
rect 5905 1769 5951 2012
rect 6517 1952 6563 2141
rect 6090 1929 6166 1942
rect 6090 1873 6101 1929
rect 6156 1873 6166 1929
rect 6090 1862 6166 1873
rect 6313 1769 6359 1836
rect 193 1686 6359 1769
rect 193 1439 239 1686
rect -28 1416 48 1429
rect -28 1414 -17 1416
rect -305 1360 -17 1414
rect 38 1360 48 1416
rect -305 1349 48 1360
rect -305 1344 30 1349
rect -305 347 -235 1344
rect 397 1155 443 1329
rect 601 1282 647 1686
rect 781 1614 883 1627
rect 781 1540 793 1614
rect 867 1540 883 1614
rect 781 1530 883 1540
rect 805 1445 851 1530
rect 1009 1442 1055 1686
rect 585 1281 647 1282
rect 527 1268 647 1281
rect 527 1213 538 1268
rect 587 1220 647 1268
rect 587 1213 631 1220
rect 527 1201 631 1213
rect 1213 1155 1259 1329
rect 1417 1282 1463 1686
rect 1585 1630 1691 1631
rect 1585 1614 1692 1630
rect 1585 1540 1598 1614
rect 1672 1540 1692 1614
rect 1585 1533 1692 1540
rect 1585 1531 1691 1533
rect 1621 1445 1667 1531
rect 1825 1425 1871 1686
rect 1406 1281 1463 1282
rect 1348 1268 1463 1281
rect 1348 1213 1359 1268
rect 1408 1217 1463 1268
rect 1408 1213 1425 1217
rect 1348 1201 1425 1213
rect 2029 1155 2075 1329
rect 2233 1284 2279 1686
rect 2407 1614 2509 1630
rect 2407 1540 2421 1614
rect 2495 1540 2509 1614
rect 2407 1533 2509 1540
rect 2437 1445 2483 1533
rect 2641 1412 2687 1686
rect 2214 1283 2279 1284
rect 2156 1270 2279 1283
rect 2156 1215 2167 1270
rect 2216 1217 2279 1270
rect 2216 1215 2260 1217
rect 2156 1203 2260 1215
rect 2845 1155 2891 1329
rect 3049 1285 3095 1686
rect 3226 1614 3328 1628
rect 3226 1540 3235 1614
rect 3309 1540 3328 1614
rect 3226 1531 3328 1540
rect 3253 1445 3299 1531
rect 3457 1417 3503 1686
rect 3038 1284 3095 1285
rect 2980 1271 3095 1284
rect 2980 1216 2991 1271
rect 3040 1225 3095 1271
rect 3040 1216 3084 1225
rect 2980 1204 3084 1216
rect 3661 1155 3707 1329
rect 3865 1285 3911 1686
rect 4044 1614 4146 1632
rect 4044 1540 4057 1614
rect 4131 1540 4146 1614
rect 4044 1535 4146 1540
rect 4069 1445 4115 1535
rect 4273 1429 4319 1686
rect 3851 1284 3911 1285
rect 3793 1271 3911 1284
rect 3793 1216 3804 1271
rect 3853 1225 3911 1271
rect 3853 1216 3897 1225
rect 3793 1204 3897 1216
rect 4477 1155 4523 1329
rect 4681 1287 4727 1686
rect 4850 1614 4952 1630
rect 4850 1540 4862 1614
rect 4936 1540 4952 1614
rect 4850 1533 4952 1540
rect 4885 1445 4931 1533
rect 5089 1427 5135 1686
rect 4668 1286 4727 1287
rect 4610 1273 4727 1286
rect 4610 1218 4621 1273
rect 4670 1226 4727 1273
rect 4670 1218 4714 1226
rect 4610 1206 4714 1218
rect 5293 1155 5339 1329
rect 5497 1287 5543 1686
rect 5658 1629 5760 1630
rect 5655 1614 5760 1629
rect 5655 1540 5669 1614
rect 5743 1540 5760 1614
rect 5655 1533 5760 1540
rect 5655 1528 5759 1533
rect 5701 1445 5747 1528
rect 5905 1435 5951 1686
rect 6313 1412 6359 1686
rect 6500 1422 6576 1430
rect 6778 1422 6848 2755
rect 6500 1417 6848 1422
rect 6500 1361 6511 1417
rect 6566 1361 6848 1417
rect 6500 1352 6848 1361
rect 6500 1350 6576 1352
rect 5487 1286 5543 1287
rect 5429 1273 5543 1286
rect 5429 1218 5440 1273
rect 5489 1226 5543 1273
rect 5489 1218 5533 1226
rect 5429 1206 5533 1218
rect 6109 1155 6155 1329
rect -110 1134 6663 1155
rect -110 1011 -38 1134
rect 87 1076 192 1134
rect 87 1020 172 1076
rect 87 1011 192 1020
rect 317 1011 422 1134
rect 547 1011 652 1134
rect 777 1011 882 1134
rect 1007 1011 1112 1134
rect 1237 1011 1342 1134
rect 1467 1011 1572 1134
rect 1697 1011 1802 1134
rect 1927 1011 2032 1134
rect 2157 1011 2262 1134
rect 2387 1011 2492 1134
rect 2617 1011 2722 1134
rect 2847 1011 2952 1134
rect 3077 1011 3182 1134
rect 3307 1011 3412 1134
rect 3537 1011 3642 1134
rect 3767 1011 3872 1134
rect 3997 1011 4102 1134
rect 4227 1011 4332 1134
rect 4457 1011 4562 1134
rect 4687 1011 4792 1134
rect 4917 1011 5022 1134
rect 5147 1011 5252 1134
rect 5377 1011 5482 1134
rect 5607 1011 5712 1134
rect 5837 1011 5942 1134
rect 6067 1011 6172 1134
rect 6297 1011 6402 1134
rect 6527 1011 6663 1134
rect -110 946 6663 1011
rect 0 878 6655 898
rect 0 760 18 878
rect 135 760 248 878
rect 365 760 478 878
rect 595 760 708 878
rect 825 760 938 878
rect 1055 760 1168 878
rect 1285 760 1398 878
rect 1515 760 1628 878
rect 1745 760 1858 878
rect 1975 760 2088 878
rect 2205 760 2318 878
rect 2435 760 2548 878
rect 2665 760 2778 878
rect 2895 760 3008 878
rect 3125 760 3238 878
rect 3355 760 3468 878
rect 3585 760 3698 878
rect 3815 760 3928 878
rect 4045 760 4158 878
rect 4275 760 4388 878
rect 4505 760 4618 878
rect 4735 760 4848 878
rect 4965 760 5078 878
rect 5195 760 5308 878
rect 5425 760 5538 878
rect 5655 760 5768 878
rect 5885 760 5998 878
rect 6115 760 6228 878
rect 6345 760 6458 878
rect 6575 760 6655 878
rect 0 742 6655 760
rect 117 681 207 690
rect 117 609 126 681
rect 198 609 207 681
rect 117 600 207 609
rect 445 542 491 742
rect 1261 542 1307 742
rect 2077 542 2123 742
rect 2893 542 2939 742
rect 3709 542 3755 742
rect 4525 542 4571 742
rect 5341 542 5387 742
rect 6157 542 6203 742
rect 220 511 300 526
rect 220 454 232 511
rect 285 454 300 511
rect 220 442 300 454
rect 629 514 709 529
rect 629 457 641 514
rect 694 457 709 514
rect 629 445 709 457
rect 1034 513 1114 528
rect 1034 456 1046 513
rect 1099 456 1114 513
rect 1034 444 1114 456
rect 1443 514 1523 529
rect 1443 457 1455 514
rect 1508 457 1523 514
rect 1443 445 1523 457
rect 1850 514 1930 529
rect 1850 457 1862 514
rect 1915 457 1930 514
rect 1850 445 1930 457
rect 2261 514 2341 529
rect 2261 457 2273 514
rect 2326 457 2341 514
rect 2261 445 2341 457
rect 2668 515 2748 530
rect 2668 458 2680 515
rect 2733 458 2748 515
rect 2668 446 2748 458
rect 3077 514 3157 529
rect 3077 457 3089 514
rect 3142 457 3157 514
rect 3077 445 3157 457
rect 3485 516 3565 531
rect 3485 459 3497 516
rect 3550 459 3565 516
rect 3485 447 3565 459
rect 3896 516 3976 531
rect 3896 459 3908 516
rect 3961 459 3976 516
rect 3896 447 3976 459
rect 4302 514 4382 529
rect 4302 457 4314 514
rect 4367 457 4382 514
rect 4302 445 4382 457
rect 4711 514 4791 529
rect 4711 457 4723 514
rect 4776 457 4791 514
rect 4711 445 4791 457
rect 5121 514 5201 529
rect 5121 457 5133 514
rect 5186 457 5201 514
rect 5121 445 5201 457
rect 5522 518 5602 533
rect 5522 461 5534 518
rect 5587 461 5602 518
rect 5522 449 5602 461
rect 5934 514 6014 529
rect 5934 457 5946 514
rect 5999 457 6014 514
rect 5934 445 6014 457
rect 6340 518 6420 533
rect 6340 461 6352 518
rect 6405 461 6420 518
rect 6340 449 6420 461
rect 37 347 83 426
rect 853 347 899 426
rect 1669 347 1715 426
rect 2485 347 2531 426
rect 3301 347 3347 427
rect 4117 347 4163 427
rect 4933 347 4979 426
rect 5749 347 5795 427
rect 6565 347 6611 426
rect 6778 347 6848 1352
rect -305 277 6848 347
rect -117 205 -37 223
rect -117 157 -103 205
rect -56 157 -37 205
rect 445 186 491 277
rect 1261 186 1307 277
rect 2077 186 2123 277
rect 2893 186 2939 277
rect 3709 186 3755 277
rect 4525 186 4571 277
rect 5341 186 5387 277
rect 6157 186 6203 277
rect -117 140 -37 157
rect 220 157 300 172
rect 220 100 232 157
rect 285 100 300 157
rect 220 88 300 100
rect 627 162 707 177
rect 627 105 639 162
rect 692 105 707 162
rect 627 93 707 105
rect 1037 157 1117 172
rect 1037 100 1049 157
rect 1102 100 1117 157
rect 1037 88 1117 100
rect 1444 154 1524 169
rect 1444 97 1456 154
rect 1509 97 1524 154
rect 1444 85 1524 97
rect 1854 154 1934 169
rect 1854 97 1866 154
rect 1919 97 1934 154
rect 1854 85 1934 97
rect 2261 161 2341 176
rect 2261 104 2273 161
rect 2326 104 2341 161
rect 2261 92 2341 104
rect 2667 158 2747 173
rect 2667 101 2679 158
rect 2732 101 2747 158
rect 2667 89 2747 101
rect 3078 157 3158 172
rect 3078 100 3090 157
rect 3143 100 3158 157
rect 3078 88 3158 100
rect 3482 157 3562 172
rect 3482 100 3494 157
rect 3547 100 3562 157
rect 3482 88 3562 100
rect 3893 157 3973 172
rect 3893 100 3905 157
rect 3958 100 3973 157
rect 3893 88 3973 100
rect 4300 157 4380 172
rect 4300 100 4312 157
rect 4365 100 4380 157
rect 4300 88 4380 100
rect 4707 162 4787 177
rect 4707 105 4719 162
rect 4772 105 4787 162
rect 4707 93 4787 105
rect 5117 155 5197 170
rect 5117 98 5129 155
rect 5182 98 5197 155
rect 5117 86 5197 98
rect 5523 155 5603 170
rect 5523 98 5535 155
rect 5588 98 5603 155
rect 5523 86 5603 98
rect 5933 155 6013 170
rect 5933 98 5945 155
rect 5998 98 6013 155
rect 5933 86 6013 98
rect 6340 156 6420 171
rect 6340 99 6352 156
rect 6405 99 6420 156
rect 6340 87 6420 99
rect 37 -111 83 70
rect 321 22 412 31
rect 321 -50 330 22
rect 402 -50 412 22
rect 321 -53 412 -50
rect 321 -59 411 -53
rect 853 -111 899 70
rect 1669 -111 1715 70
rect 2485 -111 2531 70
rect 3301 -111 3347 70
rect 4117 -111 4163 70
rect 4933 -111 4979 70
rect 5749 -111 5795 70
rect 6565 -111 6611 70
rect 8 -131 6663 -111
rect 8 -249 26 -131
rect 143 -249 256 -131
rect 373 -249 486 -131
rect 603 -249 716 -131
rect 833 -249 946 -131
rect 1063 -249 1176 -131
rect 1293 -249 1406 -131
rect 1523 -249 1636 -131
rect 1753 -249 1866 -131
rect 1983 -249 2096 -131
rect 2213 -249 2326 -131
rect 2443 -249 2556 -131
rect 2673 -249 2786 -131
rect 2903 -249 3016 -131
rect 3133 -249 3246 -131
rect 3363 -249 3476 -131
rect 3593 -249 3706 -131
rect 3823 -249 3936 -131
rect 4053 -249 4166 -131
rect 4283 -249 4396 -131
rect 4513 -249 4626 -131
rect 4743 -249 4856 -131
rect 4973 -249 5086 -131
rect 5203 -249 5316 -131
rect 5433 -249 5546 -131
rect 5663 -249 5776 -131
rect 5893 -249 6006 -131
rect 6123 -249 6236 -131
rect 6353 -249 6466 -131
rect 6583 -249 6663 -131
rect 8 -267 6663 -249
<< via1 >>
rect 47 4710 101 4765
rect 6488 4705 6542 4760
rect 1558 4533 1612 4588
rect 2371 4527 2425 4582
rect 1965 3865 2019 3920
rect 2782 3873 2836 3928
rect 62 3686 116 3741
rect 6486 3684 6540 3739
rect 29 3472 85 3528
rect 6472 3463 6527 3519
rect 6527 3463 6528 3519
rect 147 3322 206 3328
rect 147 3274 150 3322
rect 150 3274 198 3322
rect 198 3274 206 3322
rect 147 3270 206 3274
rect 191 3116 245 3171
rect 598 3116 652 3171
rect 1009 3112 1063 3167
rect 1413 3113 1467 3168
rect 1819 3111 1873 3166
rect 2229 3113 2283 3168
rect 2634 3110 2688 3165
rect 3043 3110 3097 3165
rect 3454 3110 3508 3165
rect 3859 3110 3913 3165
rect 4265 3112 4319 3167
rect 4675 3114 4729 3169
rect 5082 3111 5136 3166
rect 5491 3111 5545 3166
rect 5899 3113 5953 3168
rect 6305 3116 6359 3171
rect 187 2600 241 2655
rect 598 2602 652 2657
rect 1001 2605 1055 2660
rect 1411 2608 1465 2663
rect 1818 2607 1872 2662
rect 2225 2606 2279 2661
rect 2633 2604 2687 2659
rect 3045 2602 3099 2657
rect 3450 2605 3504 2660
rect 3859 2604 3913 2659
rect 4267 2602 4321 2657
rect 4675 2602 4729 2657
rect 5082 2601 5136 2656
rect 5490 2606 5544 2661
rect 5897 2606 5951 2661
rect 6307 2604 6361 2659
rect 226 2418 280 2477
rect 6269 2480 6325 2483
rect 6269 2430 6276 2480
rect 6276 2430 6325 2480
rect 6269 2427 6325 2430
rect 184 2215 192 2271
rect 192 2215 236 2271
rect 6475 2210 6527 2266
rect 949 2081 1004 2082
rect 949 2026 951 2081
rect 951 2026 1000 2081
rect 1000 2026 1004 2081
rect 949 2025 1004 2026
rect 391 1871 446 1927
rect 1207 1877 1262 1933
rect 2023 1870 2078 1926
rect 2837 1874 2892 1930
rect 3654 1869 3709 1925
rect 4471 1872 4526 1928
rect 5841 2081 5895 2084
rect 5841 2030 5843 2081
rect 5843 2030 5892 2081
rect 5892 2030 5895 2081
rect 5287 1871 5342 1927
rect 6101 1873 6156 1929
rect -17 1360 38 1416
rect 793 1601 867 1614
rect 793 1553 806 1601
rect 806 1553 854 1601
rect 854 1553 867 1601
rect 793 1540 867 1553
rect 1598 1601 1672 1614
rect 1598 1553 1611 1601
rect 1611 1553 1659 1601
rect 1659 1553 1672 1601
rect 1598 1540 1672 1553
rect 2421 1601 2495 1614
rect 2421 1553 2434 1601
rect 2434 1553 2482 1601
rect 2482 1553 2495 1601
rect 2421 1540 2495 1553
rect 3235 1601 3309 1614
rect 3235 1553 3248 1601
rect 3248 1553 3296 1601
rect 3296 1553 3309 1601
rect 3235 1540 3309 1553
rect 4057 1601 4131 1614
rect 4057 1553 4070 1601
rect 4070 1553 4118 1601
rect 4118 1553 4131 1601
rect 4057 1540 4131 1553
rect 4862 1601 4936 1614
rect 4862 1553 4875 1601
rect 4875 1553 4923 1601
rect 4923 1553 4936 1601
rect 4862 1540 4936 1553
rect 5669 1601 5743 1614
rect 5669 1553 5682 1601
rect 5682 1553 5730 1601
rect 5730 1553 5743 1601
rect 5669 1540 5743 1553
rect 6511 1361 6566 1417
rect 172 1020 192 1076
rect 192 1020 224 1076
rect 6441 1050 6493 1106
rect 37 784 89 840
rect 6492 783 6544 839
rect 132 615 185 672
rect 232 454 285 511
rect 641 457 694 514
rect 1046 456 1099 513
rect 1455 457 1508 514
rect 1862 457 1915 514
rect 2273 457 2326 514
rect 2680 458 2733 515
rect 3089 457 3142 514
rect 3497 459 3550 516
rect 3908 459 3961 516
rect 4314 457 4367 514
rect 4723 457 4776 514
rect 5133 457 5186 514
rect 5534 461 5587 518
rect 5946 457 5999 514
rect 6352 461 6405 518
rect 232 100 285 157
rect 639 105 692 162
rect 1049 100 1102 157
rect 1456 97 1509 154
rect 1866 97 1919 154
rect 2273 104 2326 161
rect 2679 101 2732 158
rect 3090 100 3143 157
rect 3494 100 3547 157
rect 3905 100 3958 157
rect 4312 100 4365 157
rect 4719 105 4772 162
rect 5129 98 5182 155
rect 5535 98 5588 155
rect 5945 98 5998 155
rect 6352 99 6405 156
rect 344 -41 397 16
rect 46 -234 98 -178
rect 6509 -233 6561 -177
<< metal2 >>
rect 37 4765 114 4777
rect 37 4710 47 4765
rect 101 4710 114 4765
rect 37 4698 114 4710
rect 6478 4760 6555 4772
rect 6478 4705 6488 4760
rect 6542 4705 6555 4760
rect 56 3790 112 4698
rect 6478 4693 6555 4705
rect 1548 4588 1625 4600
rect 1548 4533 1558 4588
rect 1612 4578 1625 4588
rect 2361 4586 2438 4594
rect 2361 4582 2845 4586
rect 2361 4578 2371 4582
rect 1612 4533 2371 4578
rect 1548 4527 2371 4533
rect 2425 4530 2845 4582
rect 2425 4527 2438 4530
rect 1548 4522 2438 4527
rect 1548 4521 1625 4522
rect 1961 3932 2017 4522
rect 2361 4515 2438 4522
rect 2789 3940 2845 4530
rect 1955 3925 2032 3932
rect 2772 3928 2849 3940
rect 2772 3925 2782 3928
rect 1955 3920 2782 3925
rect 1955 3865 1965 3920
rect 2019 3873 2782 3920
rect 2836 3873 2849 3928
rect 2019 3869 2849 3873
rect 2019 3865 2032 3869
rect 1955 3853 2032 3865
rect 2772 3861 2849 3869
rect -356 3753 112 3790
rect 6483 3778 6539 4693
rect -356 3741 129 3753
rect 6483 3751 6917 3778
rect -356 3686 62 3741
rect 116 3686 129 3741
rect -356 3674 129 3686
rect 6476 3739 6917 3751
rect 6476 3684 6486 3739
rect 6540 3684 6917 3739
rect 6476 3680 6917 3684
rect -356 3673 98 3674
rect -356 833 -239 3673
rect 6476 3672 6553 3680
rect 21 3528 96 3537
rect 6462 3528 6537 3532
rect -123 3472 29 3528
rect 85 3472 96 3528
rect -123 2273 -67 3472
rect 21 3463 96 3472
rect 6460 3519 6537 3528
rect 6460 3463 6472 3519
rect 6528 3463 6707 3519
rect 6460 3458 6537 3463
rect 6460 3454 6535 3458
rect 135 3330 217 3341
rect 53 3328 217 3330
rect 53 3270 147 3328
rect 206 3270 217 3328
rect 53 3256 217 3270
rect 53 2464 109 3256
rect 181 3171 258 3183
rect 181 3116 191 3171
rect 245 3116 258 3171
rect 181 3104 258 3116
rect 588 3171 665 3183
rect 588 3116 598 3171
rect 652 3116 665 3171
rect 588 3104 665 3116
rect 999 3167 1076 3179
rect 999 3112 1009 3167
rect 1063 3112 1076 3167
rect 189 2667 245 3104
rect 595 2669 651 3104
rect 999 3100 1076 3112
rect 1403 3168 1480 3180
rect 1403 3113 1413 3168
rect 1467 3113 1480 3168
rect 1403 3101 1480 3113
rect 1809 3166 1886 3178
rect 1809 3111 1819 3166
rect 1873 3111 1886 3166
rect 1002 2672 1058 3100
rect 1416 2675 1472 3101
rect 1809 3099 1886 3111
rect 2219 3168 2296 3180
rect 2219 3113 2229 3168
rect 2283 3113 2296 3168
rect 2219 3101 2296 3113
rect 2624 3165 2701 3177
rect 2624 3110 2634 3165
rect 2688 3110 2701 3165
rect 177 2661 254 2667
rect 588 2661 665 2669
rect 991 2661 1068 2672
rect 1401 2663 1478 2675
rect 1822 2674 1878 3099
rect 1401 2661 1411 2663
rect 177 2660 1411 2661
rect 177 2657 1001 2660
rect 177 2655 598 2657
rect 177 2600 187 2655
rect 241 2605 598 2655
rect 241 2600 254 2605
rect 177 2588 254 2600
rect 588 2602 598 2605
rect 652 2605 1001 2657
rect 1055 2608 1411 2660
rect 1465 2661 1478 2663
rect 1808 2662 1885 2674
rect 2229 2673 2285 3101
rect 2624 3098 2701 3110
rect 3033 3165 3110 3177
rect 3033 3110 3043 3165
rect 3097 3110 3110 3165
rect 3033 3098 3110 3110
rect 3444 3165 3521 3177
rect 3444 3110 3454 3165
rect 3508 3110 3521 3165
rect 3444 3098 3521 3110
rect 3849 3165 3926 3177
rect 3849 3110 3859 3165
rect 3913 3110 3926 3165
rect 3849 3098 3926 3110
rect 4255 3167 4332 3179
rect 4255 3112 4265 3167
rect 4319 3112 4332 3167
rect 4255 3100 4332 3112
rect 4665 3169 4742 3181
rect 4665 3114 4675 3169
rect 4729 3114 4742 3169
rect 4665 3102 4742 3114
rect 5072 3166 5149 3178
rect 5072 3111 5082 3166
rect 5136 3111 5149 3166
rect 1808 2661 1818 2662
rect 1465 2608 1818 2661
rect 1055 2607 1818 2608
rect 1872 2661 1885 2662
rect 2215 2661 2292 2673
rect 2638 2671 2694 3098
rect 2623 2661 2700 2671
rect 3048 2669 3104 3098
rect 3456 2672 3512 3098
rect 3035 2661 3112 2669
rect 3440 2661 3517 2672
rect 3865 2671 3921 3098
rect 3849 2661 3926 2671
rect 4268 2669 4324 3100
rect 4674 2669 4730 3102
rect 5072 3099 5149 3111
rect 5481 3166 5558 3178
rect 5481 3111 5491 3166
rect 5545 3111 5558 3166
rect 5481 3099 5558 3111
rect 5889 3168 5966 3180
rect 5889 3113 5899 3168
rect 5953 3113 5966 3168
rect 5889 3101 5966 3113
rect 6295 3171 6372 3183
rect 6295 3116 6305 3171
rect 6359 3116 6372 3171
rect 6295 3104 6372 3116
rect 4257 2661 4334 2669
rect 4665 2661 4742 2669
rect 5086 2668 5142 3099
rect 5497 2673 5553 3099
rect 5902 2673 5958 3101
rect 5072 2661 5149 2668
rect 5480 2661 5557 2673
rect 5887 2661 5964 2673
rect 6310 2671 6366 3104
rect 6297 2661 6374 2671
rect 1872 2607 2225 2661
rect 1055 2606 2225 2607
rect 2279 2660 5490 2661
rect 2279 2659 3450 2660
rect 2279 2606 2633 2659
rect 1055 2605 2633 2606
rect 652 2602 665 2605
rect 588 2590 665 2602
rect 991 2593 1068 2605
rect 1401 2596 1478 2605
rect 1808 2595 1885 2605
rect 2215 2594 2292 2605
rect 2623 2604 2633 2605
rect 2687 2657 3450 2659
rect 2687 2605 3045 2657
rect 2687 2604 2700 2605
rect 2623 2592 2700 2604
rect 3035 2602 3045 2605
rect 3099 2605 3450 2657
rect 3504 2659 5490 2660
rect 3504 2605 3859 2659
rect 3099 2602 3112 2605
rect 3035 2590 3112 2602
rect 3440 2593 3517 2605
rect 3849 2604 3859 2605
rect 3913 2657 5490 2659
rect 3913 2605 4267 2657
rect 3913 2604 3926 2605
rect 3849 2592 3926 2604
rect 4257 2602 4267 2605
rect 4321 2605 4675 2657
rect 4321 2602 4334 2605
rect 4257 2590 4334 2602
rect 4665 2602 4675 2605
rect 4729 2656 5490 2657
rect 4729 2605 5082 2656
rect 4729 2602 4742 2605
rect 4665 2590 4742 2602
rect 5072 2601 5082 2605
rect 5136 2606 5490 2656
rect 5544 2606 5897 2661
rect 5951 2659 6374 2661
rect 5951 2606 6307 2659
rect 5136 2605 6307 2606
rect 5136 2601 5149 2605
rect 5072 2589 5149 2601
rect 5480 2594 5557 2605
rect 5887 2594 5964 2605
rect 6297 2604 6307 2605
rect 6361 2604 6374 2659
rect 6297 2592 6374 2604
rect 212 2477 296 2492
rect 6255 2483 6340 2507
rect 212 2464 226 2477
rect 53 2418 226 2464
rect 280 2464 296 2477
rect 280 2418 1001 2464
rect 53 2408 1001 2418
rect 212 2404 296 2408
rect 170 2273 246 2283
rect -123 2271 246 2273
rect -123 2217 184 2271
rect 170 2215 184 2217
rect 236 2215 246 2271
rect 170 2203 246 2215
rect 179 1768 235 2203
rect 945 2093 1001 2408
rect 5840 2427 6269 2483
rect 6325 2427 6340 2483
rect 5840 2093 5896 2427
rect 6255 2416 6340 2427
rect 6461 2269 6537 2278
rect 6651 2269 6707 3463
rect 6461 2266 6707 2269
rect 6461 2210 6475 2266
rect 6527 2213 6707 2266
rect 6527 2210 6537 2213
rect 6461 2198 6537 2210
rect 940 2082 1017 2093
rect 940 2025 949 2082
rect 1004 2025 1017 2082
rect 940 2013 1017 2025
rect 5829 2084 5910 2093
rect 5829 2030 5841 2084
rect 5895 2030 5910 2084
rect 5829 2013 5910 2030
rect 380 1927 456 1940
rect 380 1871 391 1927
rect 446 1871 456 1927
rect 380 1860 456 1871
rect 1196 1933 1272 1946
rect 1196 1877 1207 1933
rect 1262 1877 1272 1933
rect 1196 1866 1272 1877
rect 2012 1926 2088 1939
rect 2012 1870 2023 1926
rect 2078 1870 2088 1926
rect -149 1712 235 1768
rect -149 1080 -93 1712
rect 384 1615 440 1860
rect 781 1615 883 1627
rect 1200 1615 1256 1866
rect 2012 1859 2088 1870
rect 2826 1930 2902 1943
rect 2826 1874 2837 1930
rect 2892 1874 2902 1930
rect 2826 1863 2902 1874
rect 3643 1925 3719 1938
rect 3643 1869 3654 1925
rect 3709 1869 3719 1925
rect 1585 1630 1691 1631
rect 1585 1615 1692 1630
rect 2022 1615 2078 1859
rect 2407 1615 2509 1630
rect 2831 1615 2887 1863
rect 3643 1858 3719 1869
rect 4460 1928 4536 1941
rect 4460 1872 4471 1928
rect 4526 1872 4536 1928
rect 4460 1861 4536 1872
rect 5276 1927 5352 1940
rect 5276 1871 5287 1927
rect 5342 1871 5352 1927
rect 3226 1615 3328 1628
rect 3651 1615 3707 1858
rect 4044 1615 4146 1632
rect 4467 1615 4523 1861
rect 5276 1860 5352 1871
rect 6090 1929 6166 1942
rect 6090 1873 6101 1929
rect 6156 1873 6166 1929
rect 6090 1862 6166 1873
rect 4850 1615 4952 1630
rect 5281 1615 5337 1860
rect 5658 1629 5760 1630
rect 5655 1615 5760 1629
rect 6099 1615 6155 1862
rect 6472 1821 6528 2198
rect 6472 1765 6742 1821
rect -11 1614 6567 1615
rect -11 1613 793 1614
rect -19 1540 793 1613
rect 867 1540 1598 1614
rect 1672 1540 2421 1614
rect 2495 1540 3235 1614
rect 3309 1540 4057 1614
rect 4131 1540 4862 1614
rect 4936 1540 5669 1614
rect 5743 1613 6567 1614
rect 5743 1540 6571 1613
rect -19 1539 6571 1540
rect -19 1429 37 1539
rect 781 1530 883 1539
rect 1585 1533 1692 1539
rect 2407 1533 2509 1539
rect 1585 1531 1691 1533
rect 3226 1531 3328 1539
rect 4044 1535 4146 1539
rect 4850 1533 4952 1539
rect 5655 1533 5760 1539
rect 5655 1528 5759 1533
rect 6515 1430 6571 1539
rect -28 1416 48 1429
rect -28 1360 -17 1416
rect 38 1360 48 1416
rect -28 1349 48 1360
rect 6500 1417 6576 1430
rect 6500 1361 6511 1417
rect 6566 1361 6576 1417
rect 6500 1350 6576 1361
rect 6427 1106 6503 1118
rect 158 1080 234 1088
rect -149 1076 234 1080
rect -149 1024 172 1076
rect 158 1020 172 1024
rect 224 1020 234 1076
rect 6427 1050 6441 1106
rect 6493 1105 6503 1106
rect 6686 1105 6742 1765
rect 6493 1050 6742 1105
rect 6427 1049 6742 1050
rect 6427 1038 6503 1049
rect 158 1008 234 1020
rect 23 840 99 852
rect 23 833 37 840
rect -356 784 37 833
rect 89 784 99 840
rect -356 777 99 784
rect -356 716 -110 777
rect 23 772 99 777
rect 6478 840 6554 851
rect 6478 839 6556 840
rect 6478 783 6492 839
rect 6544 823 6556 839
rect 6544 822 6642 823
rect 6819 822 6917 3680
rect 6544 783 6917 822
rect 6478 771 6917 783
rect -227 713 -110 716
rect 6500 724 6917 771
rect -227 -183 -171 713
rect 120 673 200 687
rect 74 672 200 673
rect 74 615 132 672
rect 185 615 200 672
rect 74 603 200 615
rect 74 26 130 603
rect 220 516 300 526
rect 629 516 709 529
rect 1034 516 1114 528
rect 1443 516 1523 529
rect 1850 516 1930 529
rect 2261 516 2341 529
rect 2668 516 2748 530
rect 3077 516 3157 529
rect 3485 516 3565 531
rect 3896 516 3976 531
rect 4302 516 4382 529
rect 4711 516 4791 529
rect 5121 516 5201 529
rect 5522 518 5602 533
rect 5522 516 5534 518
rect 220 515 3497 516
rect 220 514 2680 515
rect 220 511 641 514
rect 220 454 232 511
rect 285 460 641 511
rect 285 454 300 460
rect 220 442 300 454
rect 629 457 641 460
rect 694 513 1455 514
rect 694 460 1046 513
rect 694 457 709 460
rect 629 445 709 457
rect 1034 456 1046 460
rect 1099 460 1455 513
rect 1099 456 1114 460
rect 232 172 288 442
rect 641 177 697 445
rect 1034 444 1114 456
rect 1443 457 1455 460
rect 1508 460 1862 514
rect 1508 457 1523 460
rect 1443 445 1523 457
rect 1850 457 1862 460
rect 1915 460 2273 514
rect 1915 457 1930 460
rect 1850 445 1930 457
rect 2261 457 2273 460
rect 2326 460 2680 514
rect 2326 457 2341 460
rect 2261 445 2341 457
rect 2668 458 2680 460
rect 2733 514 3497 515
rect 2733 460 3089 514
rect 2733 458 2748 460
rect 2668 446 2748 458
rect 3077 457 3089 460
rect 3142 460 3497 514
rect 3142 457 3157 460
rect 220 157 300 172
rect 220 100 232 157
rect 285 100 300 157
rect 220 88 300 100
rect 627 162 707 177
rect 1045 172 1101 444
rect 627 105 639 162
rect 692 105 707 162
rect 627 93 707 105
rect 1037 157 1117 172
rect 1454 169 1510 445
rect 1862 169 1918 445
rect 2270 176 2326 445
rect 1037 100 1049 157
rect 1102 100 1117 157
rect 1037 88 1117 100
rect 1444 154 1524 169
rect 1444 97 1456 154
rect 1509 97 1524 154
rect 1444 85 1524 97
rect 1854 154 1934 169
rect 1854 97 1866 154
rect 1919 97 1934 154
rect 1854 85 1934 97
rect 2261 161 2341 176
rect 2677 173 2733 446
rect 3077 445 3157 457
rect 3485 459 3497 460
rect 3550 460 3908 516
rect 3550 459 3565 460
rect 3485 447 3565 459
rect 3896 459 3908 460
rect 3961 514 5534 516
rect 3961 460 4314 514
rect 3961 459 3976 460
rect 3896 447 3976 459
rect 4302 457 4314 460
rect 4367 460 4723 514
rect 4367 457 4382 460
rect 2261 104 2273 161
rect 2326 104 2341 161
rect 2261 92 2341 104
rect 2667 158 2747 173
rect 3096 172 3152 445
rect 3494 172 3550 447
rect 3906 172 3962 447
rect 4302 445 4382 457
rect 4711 457 4723 460
rect 4776 460 5133 514
rect 4776 457 4791 460
rect 4711 445 4791 457
rect 5121 457 5133 460
rect 5186 461 5534 514
rect 5587 516 5602 518
rect 5934 516 6014 529
rect 6340 518 6420 533
rect 6340 516 6352 518
rect 5587 514 6352 516
rect 5587 461 5946 514
rect 5186 460 5946 461
rect 5186 457 5201 460
rect 5121 445 5201 457
rect 5522 449 5602 460
rect 5934 457 5946 460
rect 5999 461 6352 514
rect 6405 461 6420 518
rect 5999 460 6420 461
rect 5999 457 6014 460
rect 4311 172 4367 445
rect 4722 177 4778 445
rect 2667 101 2679 158
rect 2732 101 2747 158
rect 2667 89 2747 101
rect 3078 157 3158 172
rect 3078 100 3090 157
rect 3143 100 3158 157
rect 3078 88 3158 100
rect 3482 157 3562 172
rect 3482 100 3494 157
rect 3547 100 3562 157
rect 3482 88 3562 100
rect 3893 157 3973 172
rect 3893 100 3905 157
rect 3958 100 3973 157
rect 3893 88 3973 100
rect 4300 157 4380 172
rect 4300 100 4312 157
rect 4365 100 4380 157
rect 4300 88 4380 100
rect 4707 162 4787 177
rect 5133 170 5189 445
rect 5534 170 5590 449
rect 5934 445 6014 457
rect 6340 449 6420 460
rect 5950 170 6006 445
rect 6356 171 6412 449
rect 4707 105 4719 162
rect 4772 105 4787 162
rect 4707 93 4787 105
rect 5117 155 5197 170
rect 5117 98 5129 155
rect 5182 98 5197 155
rect 5117 86 5197 98
rect 5523 155 5603 170
rect 5523 98 5535 155
rect 5588 98 5603 155
rect 5523 86 5603 98
rect 5933 155 6013 170
rect 5933 98 5945 155
rect 5998 98 6013 155
rect 5933 86 6013 98
rect 6340 156 6420 171
rect 6340 99 6352 156
rect 6405 99 6420 156
rect 6340 87 6420 99
rect 332 26 412 31
rect 74 16 412 26
rect 74 -30 344 16
rect 332 -41 344 -30
rect 397 -41 412 16
rect 332 -53 412 -41
rect 6500 -165 6556 724
rect 32 -178 108 -166
rect 32 -183 46 -178
rect -227 -234 46 -183
rect 98 -234 108 -178
rect -227 -239 108 -234
rect 32 -246 108 -239
rect 6495 -177 6571 -165
rect 6495 -233 6509 -177
rect 6561 -233 6571 -177
rect 6495 -245 6571 -233
use nmos_3p3_9NPLV7  nmos_3p3_9NPLV7_0
timestamp 1693373438
transform 1 0 3324 0 1 4414
box -3324 -128 3324 128
use nmos_3p3_9NPLV7  nmos_3p3_9NPLV7_1
timestamp 1693373438
transform 1 0 3324 0 1 128
box -3324 -128 3324 128
use nmos_3p3_9NPLV7  nmos_3p3_9NPLV7_2
timestamp 1693373438
transform 1 0 3324 0 1 484
box -3324 -128 3324 128
use nmos_3p3_9NPLV7  nmos_3p3_9NPLV7_3
timestamp 1693373438
transform 1 0 3324 0 1 4038
box -3324 -128 3324 128
use pmos_3p3_DVR9E7  pmos_3p3_DVR9E7_0
timestamp 1693394299
transform 1 0 3276 0 1 1894
box -3386 -190 3386 190
use pmos_3p3_DVR9E7  pmos_3p3_DVR9E7_1
timestamp 1693394299
transform 1 0 3276 0 1 3140
box -3386 -190 3386 190
use pmos_3p3_DVR9E7  pmos_3p3_DVR9E7_2
timestamp 1693394299
transform 1 0 3276 0 1 1387
box -3386 -190 3386 190
use pmos_3p3_DVR9E7  pmos_3p3_DVR9E7_3
timestamp 1693394299
transform 1 0 3276 0 1 2617
box -3386 -190 3386 190
<< labels >>
flabel psubdiffcont 1694 -197 1694 -197 0 FreeSans 480 0 0 0 VSS
port 0 nsew
flabel via1 1071 489 1071 489 0 FreeSans 480 0 0 0 SD0_1
port 1 nsew
flabel via1 356 -14 356 -14 0 FreeSans 480 0 0 0 G0_2
port 2 nsew
flabel polycontact -84 182 -84 182 0 FreeSans 480 0 0 0 G0_1
port 3 nsew
flabel nsubdiffcont 1652 1063 1652 1063 0 FreeSans 480 0 0 0 VDD
port 4 nsew
flabel polycontact 554 1242 554 1242 0 FreeSans 480 0 0 0 G1_2
port 5 nsew
flabel via1 4 1395 4 1395 0 FreeSans 480 0 0 0 G1_1
port 6 nsew
flabel via1 623 2625 623 2625 0 FreeSans 480 0 0 0 SD2_0
port 8 nsew
flabel polycontact 359 3894 359 3894 0 FreeSans 480 0 0 0 G3_2
port 9 nsew
flabel polycontact 365 4250 365 4250 0 FreeSans 480 0 0 0 G3_1
port 10 nsew
<< end >>
