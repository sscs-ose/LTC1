magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1931 -1019 1931 1019
<< metal2 >>
rect -931 14 931 19
rect -931 -14 -926 14
rect -898 -14 -850 14
rect -822 -14 -774 14
rect -746 -14 -698 14
rect -670 -14 -622 14
rect -594 -14 -546 14
rect -518 -14 -470 14
rect -442 -14 -394 14
rect -366 -14 -318 14
rect -290 -14 -242 14
rect -214 -14 -166 14
rect -138 -14 -90 14
rect -62 -14 -14 14
rect 14 -14 62 14
rect 90 -14 138 14
rect 166 -14 214 14
rect 242 -14 290 14
rect 318 -14 366 14
rect 394 -14 442 14
rect 470 -14 518 14
rect 546 -14 594 14
rect 622 -14 670 14
rect 698 -14 746 14
rect 774 -14 822 14
rect 850 -14 898 14
rect 926 -14 931 14
rect -931 -19 931 -14
<< via2 >>
rect -926 -14 -898 14
rect -850 -14 -822 14
rect -774 -14 -746 14
rect -698 -14 -670 14
rect -622 -14 -594 14
rect -546 -14 -518 14
rect -470 -14 -442 14
rect -394 -14 -366 14
rect -318 -14 -290 14
rect -242 -14 -214 14
rect -166 -14 -138 14
rect -90 -14 -62 14
rect -14 -14 14 14
rect 62 -14 90 14
rect 138 -14 166 14
rect 214 -14 242 14
rect 290 -14 318 14
rect 366 -14 394 14
rect 442 -14 470 14
rect 518 -14 546 14
rect 594 -14 622 14
rect 670 -14 698 14
rect 746 -14 774 14
rect 822 -14 850 14
rect 898 -14 926 14
<< metal3 >>
rect -931 14 931 19
rect -931 -14 -926 14
rect -898 -14 -850 14
rect -822 -14 -774 14
rect -746 -14 -698 14
rect -670 -14 -622 14
rect -594 -14 -546 14
rect -518 -14 -470 14
rect -442 -14 -394 14
rect -366 -14 -318 14
rect -290 -14 -242 14
rect -214 -14 -166 14
rect -138 -14 -90 14
rect -62 -14 -14 14
rect 14 -14 62 14
rect 90 -14 138 14
rect 166 -14 214 14
rect 242 -14 290 14
rect 318 -14 366 14
rect 394 -14 442 14
rect 470 -14 518 14
rect 546 -14 594 14
rect 622 -14 670 14
rect 698 -14 746 14
rect 774 -14 822 14
rect 850 -14 898 14
rect 926 -14 931 14
rect -931 -19 931 -14
<< end >>
