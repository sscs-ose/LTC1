magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2727 -2045 2727 2045
<< psubdiff >>
rect -727 23 727 45
rect -727 -23 -705 23
rect -659 -23 -581 23
rect -535 -23 -457 23
rect -411 -23 -333 23
rect -287 -23 -209 23
rect -163 -23 -85 23
rect -39 -23 39 23
rect 85 -23 163 23
rect 209 -23 287 23
rect 333 -23 411 23
rect 457 -23 535 23
rect 581 -23 659 23
rect 705 -23 727 23
rect -727 -45 727 -23
<< psubdiffcont >>
rect -705 -23 -659 23
rect -581 -23 -535 23
rect -457 -23 -411 23
rect -333 -23 -287 23
rect -209 -23 -163 23
rect -85 -23 -39 23
rect 39 -23 85 23
rect 163 -23 209 23
rect 287 -23 333 23
rect 411 -23 457 23
rect 535 -23 581 23
rect 659 -23 705 23
<< metal1 >>
rect -716 23 716 34
rect -716 -23 -705 23
rect -659 -23 -581 23
rect -535 -23 -457 23
rect -411 -23 -333 23
rect -287 -23 -209 23
rect -163 -23 -85 23
rect -39 -23 39 23
rect 85 -23 163 23
rect 209 -23 287 23
rect 333 -23 411 23
rect 457 -23 535 23
rect 581 -23 659 23
rect 705 -23 716 23
rect -716 -34 716 -23
<< end >>
