magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1298 -2972 1298 2972
<< metal1 >>
rect -298 1966 298 1972
rect -298 1940 -292 1966
rect -266 1940 -230 1966
rect -204 1940 -168 1966
rect -142 1940 -106 1966
rect -80 1940 -44 1966
rect -18 1940 18 1966
rect 44 1940 80 1966
rect 106 1940 142 1966
rect 168 1940 204 1966
rect 230 1940 266 1966
rect 292 1940 298 1966
rect -298 1904 298 1940
rect -298 1878 -292 1904
rect -266 1878 -230 1904
rect -204 1878 -168 1904
rect -142 1878 -106 1904
rect -80 1878 -44 1904
rect -18 1878 18 1904
rect 44 1878 80 1904
rect 106 1878 142 1904
rect 168 1878 204 1904
rect 230 1878 266 1904
rect 292 1878 298 1904
rect -298 1842 298 1878
rect -298 1816 -292 1842
rect -266 1816 -230 1842
rect -204 1816 -168 1842
rect -142 1816 -106 1842
rect -80 1816 -44 1842
rect -18 1816 18 1842
rect 44 1816 80 1842
rect 106 1816 142 1842
rect 168 1816 204 1842
rect 230 1816 266 1842
rect 292 1816 298 1842
rect -298 1780 298 1816
rect -298 1754 -292 1780
rect -266 1754 -230 1780
rect -204 1754 -168 1780
rect -142 1754 -106 1780
rect -80 1754 -44 1780
rect -18 1754 18 1780
rect 44 1754 80 1780
rect 106 1754 142 1780
rect 168 1754 204 1780
rect 230 1754 266 1780
rect 292 1754 298 1780
rect -298 1718 298 1754
rect -298 1692 -292 1718
rect -266 1692 -230 1718
rect -204 1692 -168 1718
rect -142 1692 -106 1718
rect -80 1692 -44 1718
rect -18 1692 18 1718
rect 44 1692 80 1718
rect 106 1692 142 1718
rect 168 1692 204 1718
rect 230 1692 266 1718
rect 292 1692 298 1718
rect -298 1656 298 1692
rect -298 1630 -292 1656
rect -266 1630 -230 1656
rect -204 1630 -168 1656
rect -142 1630 -106 1656
rect -80 1630 -44 1656
rect -18 1630 18 1656
rect 44 1630 80 1656
rect 106 1630 142 1656
rect 168 1630 204 1656
rect 230 1630 266 1656
rect 292 1630 298 1656
rect -298 1594 298 1630
rect -298 1568 -292 1594
rect -266 1568 -230 1594
rect -204 1568 -168 1594
rect -142 1568 -106 1594
rect -80 1568 -44 1594
rect -18 1568 18 1594
rect 44 1568 80 1594
rect 106 1568 142 1594
rect 168 1568 204 1594
rect 230 1568 266 1594
rect 292 1568 298 1594
rect -298 1532 298 1568
rect -298 1506 -292 1532
rect -266 1506 -230 1532
rect -204 1506 -168 1532
rect -142 1506 -106 1532
rect -80 1506 -44 1532
rect -18 1506 18 1532
rect 44 1506 80 1532
rect 106 1506 142 1532
rect 168 1506 204 1532
rect 230 1506 266 1532
rect 292 1506 298 1532
rect -298 1470 298 1506
rect -298 1444 -292 1470
rect -266 1444 -230 1470
rect -204 1444 -168 1470
rect -142 1444 -106 1470
rect -80 1444 -44 1470
rect -18 1444 18 1470
rect 44 1444 80 1470
rect 106 1444 142 1470
rect 168 1444 204 1470
rect 230 1444 266 1470
rect 292 1444 298 1470
rect -298 1408 298 1444
rect -298 1382 -292 1408
rect -266 1382 -230 1408
rect -204 1382 -168 1408
rect -142 1382 -106 1408
rect -80 1382 -44 1408
rect -18 1382 18 1408
rect 44 1382 80 1408
rect 106 1382 142 1408
rect 168 1382 204 1408
rect 230 1382 266 1408
rect 292 1382 298 1408
rect -298 1346 298 1382
rect -298 1320 -292 1346
rect -266 1320 -230 1346
rect -204 1320 -168 1346
rect -142 1320 -106 1346
rect -80 1320 -44 1346
rect -18 1320 18 1346
rect 44 1320 80 1346
rect 106 1320 142 1346
rect 168 1320 204 1346
rect 230 1320 266 1346
rect 292 1320 298 1346
rect -298 1284 298 1320
rect -298 1258 -292 1284
rect -266 1258 -230 1284
rect -204 1258 -168 1284
rect -142 1258 -106 1284
rect -80 1258 -44 1284
rect -18 1258 18 1284
rect 44 1258 80 1284
rect 106 1258 142 1284
rect 168 1258 204 1284
rect 230 1258 266 1284
rect 292 1258 298 1284
rect -298 1222 298 1258
rect -298 1196 -292 1222
rect -266 1196 -230 1222
rect -204 1196 -168 1222
rect -142 1196 -106 1222
rect -80 1196 -44 1222
rect -18 1196 18 1222
rect 44 1196 80 1222
rect 106 1196 142 1222
rect 168 1196 204 1222
rect 230 1196 266 1222
rect 292 1196 298 1222
rect -298 1160 298 1196
rect -298 1134 -292 1160
rect -266 1134 -230 1160
rect -204 1134 -168 1160
rect -142 1134 -106 1160
rect -80 1134 -44 1160
rect -18 1134 18 1160
rect 44 1134 80 1160
rect 106 1134 142 1160
rect 168 1134 204 1160
rect 230 1134 266 1160
rect 292 1134 298 1160
rect -298 1098 298 1134
rect -298 1072 -292 1098
rect -266 1072 -230 1098
rect -204 1072 -168 1098
rect -142 1072 -106 1098
rect -80 1072 -44 1098
rect -18 1072 18 1098
rect 44 1072 80 1098
rect 106 1072 142 1098
rect 168 1072 204 1098
rect 230 1072 266 1098
rect 292 1072 298 1098
rect -298 1036 298 1072
rect -298 1010 -292 1036
rect -266 1010 -230 1036
rect -204 1010 -168 1036
rect -142 1010 -106 1036
rect -80 1010 -44 1036
rect -18 1010 18 1036
rect 44 1010 80 1036
rect 106 1010 142 1036
rect 168 1010 204 1036
rect 230 1010 266 1036
rect 292 1010 298 1036
rect -298 974 298 1010
rect -298 948 -292 974
rect -266 948 -230 974
rect -204 948 -168 974
rect -142 948 -106 974
rect -80 948 -44 974
rect -18 948 18 974
rect 44 948 80 974
rect 106 948 142 974
rect 168 948 204 974
rect 230 948 266 974
rect 292 948 298 974
rect -298 912 298 948
rect -298 886 -292 912
rect -266 886 -230 912
rect -204 886 -168 912
rect -142 886 -106 912
rect -80 886 -44 912
rect -18 886 18 912
rect 44 886 80 912
rect 106 886 142 912
rect 168 886 204 912
rect 230 886 266 912
rect 292 886 298 912
rect -298 850 298 886
rect -298 824 -292 850
rect -266 824 -230 850
rect -204 824 -168 850
rect -142 824 -106 850
rect -80 824 -44 850
rect -18 824 18 850
rect 44 824 80 850
rect 106 824 142 850
rect 168 824 204 850
rect 230 824 266 850
rect 292 824 298 850
rect -298 788 298 824
rect -298 762 -292 788
rect -266 762 -230 788
rect -204 762 -168 788
rect -142 762 -106 788
rect -80 762 -44 788
rect -18 762 18 788
rect 44 762 80 788
rect 106 762 142 788
rect 168 762 204 788
rect 230 762 266 788
rect 292 762 298 788
rect -298 726 298 762
rect -298 700 -292 726
rect -266 700 -230 726
rect -204 700 -168 726
rect -142 700 -106 726
rect -80 700 -44 726
rect -18 700 18 726
rect 44 700 80 726
rect 106 700 142 726
rect 168 700 204 726
rect 230 700 266 726
rect 292 700 298 726
rect -298 664 298 700
rect -298 638 -292 664
rect -266 638 -230 664
rect -204 638 -168 664
rect -142 638 -106 664
rect -80 638 -44 664
rect -18 638 18 664
rect 44 638 80 664
rect 106 638 142 664
rect 168 638 204 664
rect 230 638 266 664
rect 292 638 298 664
rect -298 602 298 638
rect -298 576 -292 602
rect -266 576 -230 602
rect -204 576 -168 602
rect -142 576 -106 602
rect -80 576 -44 602
rect -18 576 18 602
rect 44 576 80 602
rect 106 576 142 602
rect 168 576 204 602
rect 230 576 266 602
rect 292 576 298 602
rect -298 540 298 576
rect -298 514 -292 540
rect -266 514 -230 540
rect -204 514 -168 540
rect -142 514 -106 540
rect -80 514 -44 540
rect -18 514 18 540
rect 44 514 80 540
rect 106 514 142 540
rect 168 514 204 540
rect 230 514 266 540
rect 292 514 298 540
rect -298 478 298 514
rect -298 452 -292 478
rect -266 452 -230 478
rect -204 452 -168 478
rect -142 452 -106 478
rect -80 452 -44 478
rect -18 452 18 478
rect 44 452 80 478
rect 106 452 142 478
rect 168 452 204 478
rect 230 452 266 478
rect 292 452 298 478
rect -298 416 298 452
rect -298 390 -292 416
rect -266 390 -230 416
rect -204 390 -168 416
rect -142 390 -106 416
rect -80 390 -44 416
rect -18 390 18 416
rect 44 390 80 416
rect 106 390 142 416
rect 168 390 204 416
rect 230 390 266 416
rect 292 390 298 416
rect -298 354 298 390
rect -298 328 -292 354
rect -266 328 -230 354
rect -204 328 -168 354
rect -142 328 -106 354
rect -80 328 -44 354
rect -18 328 18 354
rect 44 328 80 354
rect 106 328 142 354
rect 168 328 204 354
rect 230 328 266 354
rect 292 328 298 354
rect -298 292 298 328
rect -298 266 -292 292
rect -266 266 -230 292
rect -204 266 -168 292
rect -142 266 -106 292
rect -80 266 -44 292
rect -18 266 18 292
rect 44 266 80 292
rect 106 266 142 292
rect 168 266 204 292
rect 230 266 266 292
rect 292 266 298 292
rect -298 230 298 266
rect -298 204 -292 230
rect -266 204 -230 230
rect -204 204 -168 230
rect -142 204 -106 230
rect -80 204 -44 230
rect -18 204 18 230
rect 44 204 80 230
rect 106 204 142 230
rect 168 204 204 230
rect 230 204 266 230
rect 292 204 298 230
rect -298 168 298 204
rect -298 142 -292 168
rect -266 142 -230 168
rect -204 142 -168 168
rect -142 142 -106 168
rect -80 142 -44 168
rect -18 142 18 168
rect 44 142 80 168
rect 106 142 142 168
rect 168 142 204 168
rect 230 142 266 168
rect 292 142 298 168
rect -298 106 298 142
rect -298 80 -292 106
rect -266 80 -230 106
rect -204 80 -168 106
rect -142 80 -106 106
rect -80 80 -44 106
rect -18 80 18 106
rect 44 80 80 106
rect 106 80 142 106
rect 168 80 204 106
rect 230 80 266 106
rect 292 80 298 106
rect -298 44 298 80
rect -298 18 -292 44
rect -266 18 -230 44
rect -204 18 -168 44
rect -142 18 -106 44
rect -80 18 -44 44
rect -18 18 18 44
rect 44 18 80 44
rect 106 18 142 44
rect 168 18 204 44
rect 230 18 266 44
rect 292 18 298 44
rect -298 -18 298 18
rect -298 -44 -292 -18
rect -266 -44 -230 -18
rect -204 -44 -168 -18
rect -142 -44 -106 -18
rect -80 -44 -44 -18
rect -18 -44 18 -18
rect 44 -44 80 -18
rect 106 -44 142 -18
rect 168 -44 204 -18
rect 230 -44 266 -18
rect 292 -44 298 -18
rect -298 -80 298 -44
rect -298 -106 -292 -80
rect -266 -106 -230 -80
rect -204 -106 -168 -80
rect -142 -106 -106 -80
rect -80 -106 -44 -80
rect -18 -106 18 -80
rect 44 -106 80 -80
rect 106 -106 142 -80
rect 168 -106 204 -80
rect 230 -106 266 -80
rect 292 -106 298 -80
rect -298 -142 298 -106
rect -298 -168 -292 -142
rect -266 -168 -230 -142
rect -204 -168 -168 -142
rect -142 -168 -106 -142
rect -80 -168 -44 -142
rect -18 -168 18 -142
rect 44 -168 80 -142
rect 106 -168 142 -142
rect 168 -168 204 -142
rect 230 -168 266 -142
rect 292 -168 298 -142
rect -298 -204 298 -168
rect -298 -230 -292 -204
rect -266 -230 -230 -204
rect -204 -230 -168 -204
rect -142 -230 -106 -204
rect -80 -230 -44 -204
rect -18 -230 18 -204
rect 44 -230 80 -204
rect 106 -230 142 -204
rect 168 -230 204 -204
rect 230 -230 266 -204
rect 292 -230 298 -204
rect -298 -266 298 -230
rect -298 -292 -292 -266
rect -266 -292 -230 -266
rect -204 -292 -168 -266
rect -142 -292 -106 -266
rect -80 -292 -44 -266
rect -18 -292 18 -266
rect 44 -292 80 -266
rect 106 -292 142 -266
rect 168 -292 204 -266
rect 230 -292 266 -266
rect 292 -292 298 -266
rect -298 -328 298 -292
rect -298 -354 -292 -328
rect -266 -354 -230 -328
rect -204 -354 -168 -328
rect -142 -354 -106 -328
rect -80 -354 -44 -328
rect -18 -354 18 -328
rect 44 -354 80 -328
rect 106 -354 142 -328
rect 168 -354 204 -328
rect 230 -354 266 -328
rect 292 -354 298 -328
rect -298 -390 298 -354
rect -298 -416 -292 -390
rect -266 -416 -230 -390
rect -204 -416 -168 -390
rect -142 -416 -106 -390
rect -80 -416 -44 -390
rect -18 -416 18 -390
rect 44 -416 80 -390
rect 106 -416 142 -390
rect 168 -416 204 -390
rect 230 -416 266 -390
rect 292 -416 298 -390
rect -298 -452 298 -416
rect -298 -478 -292 -452
rect -266 -478 -230 -452
rect -204 -478 -168 -452
rect -142 -478 -106 -452
rect -80 -478 -44 -452
rect -18 -478 18 -452
rect 44 -478 80 -452
rect 106 -478 142 -452
rect 168 -478 204 -452
rect 230 -478 266 -452
rect 292 -478 298 -452
rect -298 -514 298 -478
rect -298 -540 -292 -514
rect -266 -540 -230 -514
rect -204 -540 -168 -514
rect -142 -540 -106 -514
rect -80 -540 -44 -514
rect -18 -540 18 -514
rect 44 -540 80 -514
rect 106 -540 142 -514
rect 168 -540 204 -514
rect 230 -540 266 -514
rect 292 -540 298 -514
rect -298 -576 298 -540
rect -298 -602 -292 -576
rect -266 -602 -230 -576
rect -204 -602 -168 -576
rect -142 -602 -106 -576
rect -80 -602 -44 -576
rect -18 -602 18 -576
rect 44 -602 80 -576
rect 106 -602 142 -576
rect 168 -602 204 -576
rect 230 -602 266 -576
rect 292 -602 298 -576
rect -298 -638 298 -602
rect -298 -664 -292 -638
rect -266 -664 -230 -638
rect -204 -664 -168 -638
rect -142 -664 -106 -638
rect -80 -664 -44 -638
rect -18 -664 18 -638
rect 44 -664 80 -638
rect 106 -664 142 -638
rect 168 -664 204 -638
rect 230 -664 266 -638
rect 292 -664 298 -638
rect -298 -700 298 -664
rect -298 -726 -292 -700
rect -266 -726 -230 -700
rect -204 -726 -168 -700
rect -142 -726 -106 -700
rect -80 -726 -44 -700
rect -18 -726 18 -700
rect 44 -726 80 -700
rect 106 -726 142 -700
rect 168 -726 204 -700
rect 230 -726 266 -700
rect 292 -726 298 -700
rect -298 -762 298 -726
rect -298 -788 -292 -762
rect -266 -788 -230 -762
rect -204 -788 -168 -762
rect -142 -788 -106 -762
rect -80 -788 -44 -762
rect -18 -788 18 -762
rect 44 -788 80 -762
rect 106 -788 142 -762
rect 168 -788 204 -762
rect 230 -788 266 -762
rect 292 -788 298 -762
rect -298 -824 298 -788
rect -298 -850 -292 -824
rect -266 -850 -230 -824
rect -204 -850 -168 -824
rect -142 -850 -106 -824
rect -80 -850 -44 -824
rect -18 -850 18 -824
rect 44 -850 80 -824
rect 106 -850 142 -824
rect 168 -850 204 -824
rect 230 -850 266 -824
rect 292 -850 298 -824
rect -298 -886 298 -850
rect -298 -912 -292 -886
rect -266 -912 -230 -886
rect -204 -912 -168 -886
rect -142 -912 -106 -886
rect -80 -912 -44 -886
rect -18 -912 18 -886
rect 44 -912 80 -886
rect 106 -912 142 -886
rect 168 -912 204 -886
rect 230 -912 266 -886
rect 292 -912 298 -886
rect -298 -948 298 -912
rect -298 -974 -292 -948
rect -266 -974 -230 -948
rect -204 -974 -168 -948
rect -142 -974 -106 -948
rect -80 -974 -44 -948
rect -18 -974 18 -948
rect 44 -974 80 -948
rect 106 -974 142 -948
rect 168 -974 204 -948
rect 230 -974 266 -948
rect 292 -974 298 -948
rect -298 -1010 298 -974
rect -298 -1036 -292 -1010
rect -266 -1036 -230 -1010
rect -204 -1036 -168 -1010
rect -142 -1036 -106 -1010
rect -80 -1036 -44 -1010
rect -18 -1036 18 -1010
rect 44 -1036 80 -1010
rect 106 -1036 142 -1010
rect 168 -1036 204 -1010
rect 230 -1036 266 -1010
rect 292 -1036 298 -1010
rect -298 -1072 298 -1036
rect -298 -1098 -292 -1072
rect -266 -1098 -230 -1072
rect -204 -1098 -168 -1072
rect -142 -1098 -106 -1072
rect -80 -1098 -44 -1072
rect -18 -1098 18 -1072
rect 44 -1098 80 -1072
rect 106 -1098 142 -1072
rect 168 -1098 204 -1072
rect 230 -1098 266 -1072
rect 292 -1098 298 -1072
rect -298 -1134 298 -1098
rect -298 -1160 -292 -1134
rect -266 -1160 -230 -1134
rect -204 -1160 -168 -1134
rect -142 -1160 -106 -1134
rect -80 -1160 -44 -1134
rect -18 -1160 18 -1134
rect 44 -1160 80 -1134
rect 106 -1160 142 -1134
rect 168 -1160 204 -1134
rect 230 -1160 266 -1134
rect 292 -1160 298 -1134
rect -298 -1196 298 -1160
rect -298 -1222 -292 -1196
rect -266 -1222 -230 -1196
rect -204 -1222 -168 -1196
rect -142 -1222 -106 -1196
rect -80 -1222 -44 -1196
rect -18 -1222 18 -1196
rect 44 -1222 80 -1196
rect 106 -1222 142 -1196
rect 168 -1222 204 -1196
rect 230 -1222 266 -1196
rect 292 -1222 298 -1196
rect -298 -1258 298 -1222
rect -298 -1284 -292 -1258
rect -266 -1284 -230 -1258
rect -204 -1284 -168 -1258
rect -142 -1284 -106 -1258
rect -80 -1284 -44 -1258
rect -18 -1284 18 -1258
rect 44 -1284 80 -1258
rect 106 -1284 142 -1258
rect 168 -1284 204 -1258
rect 230 -1284 266 -1258
rect 292 -1284 298 -1258
rect -298 -1320 298 -1284
rect -298 -1346 -292 -1320
rect -266 -1346 -230 -1320
rect -204 -1346 -168 -1320
rect -142 -1346 -106 -1320
rect -80 -1346 -44 -1320
rect -18 -1346 18 -1320
rect 44 -1346 80 -1320
rect 106 -1346 142 -1320
rect 168 -1346 204 -1320
rect 230 -1346 266 -1320
rect 292 -1346 298 -1320
rect -298 -1382 298 -1346
rect -298 -1408 -292 -1382
rect -266 -1408 -230 -1382
rect -204 -1408 -168 -1382
rect -142 -1408 -106 -1382
rect -80 -1408 -44 -1382
rect -18 -1408 18 -1382
rect 44 -1408 80 -1382
rect 106 -1408 142 -1382
rect 168 -1408 204 -1382
rect 230 -1408 266 -1382
rect 292 -1408 298 -1382
rect -298 -1444 298 -1408
rect -298 -1470 -292 -1444
rect -266 -1470 -230 -1444
rect -204 -1470 -168 -1444
rect -142 -1470 -106 -1444
rect -80 -1470 -44 -1444
rect -18 -1470 18 -1444
rect 44 -1470 80 -1444
rect 106 -1470 142 -1444
rect 168 -1470 204 -1444
rect 230 -1470 266 -1444
rect 292 -1470 298 -1444
rect -298 -1506 298 -1470
rect -298 -1532 -292 -1506
rect -266 -1532 -230 -1506
rect -204 -1532 -168 -1506
rect -142 -1532 -106 -1506
rect -80 -1532 -44 -1506
rect -18 -1532 18 -1506
rect 44 -1532 80 -1506
rect 106 -1532 142 -1506
rect 168 -1532 204 -1506
rect 230 -1532 266 -1506
rect 292 -1532 298 -1506
rect -298 -1568 298 -1532
rect -298 -1594 -292 -1568
rect -266 -1594 -230 -1568
rect -204 -1594 -168 -1568
rect -142 -1594 -106 -1568
rect -80 -1594 -44 -1568
rect -18 -1594 18 -1568
rect 44 -1594 80 -1568
rect 106 -1594 142 -1568
rect 168 -1594 204 -1568
rect 230 -1594 266 -1568
rect 292 -1594 298 -1568
rect -298 -1630 298 -1594
rect -298 -1656 -292 -1630
rect -266 -1656 -230 -1630
rect -204 -1656 -168 -1630
rect -142 -1656 -106 -1630
rect -80 -1656 -44 -1630
rect -18 -1656 18 -1630
rect 44 -1656 80 -1630
rect 106 -1656 142 -1630
rect 168 -1656 204 -1630
rect 230 -1656 266 -1630
rect 292 -1656 298 -1630
rect -298 -1692 298 -1656
rect -298 -1718 -292 -1692
rect -266 -1718 -230 -1692
rect -204 -1718 -168 -1692
rect -142 -1718 -106 -1692
rect -80 -1718 -44 -1692
rect -18 -1718 18 -1692
rect 44 -1718 80 -1692
rect 106 -1718 142 -1692
rect 168 -1718 204 -1692
rect 230 -1718 266 -1692
rect 292 -1718 298 -1692
rect -298 -1754 298 -1718
rect -298 -1780 -292 -1754
rect -266 -1780 -230 -1754
rect -204 -1780 -168 -1754
rect -142 -1780 -106 -1754
rect -80 -1780 -44 -1754
rect -18 -1780 18 -1754
rect 44 -1780 80 -1754
rect 106 -1780 142 -1754
rect 168 -1780 204 -1754
rect 230 -1780 266 -1754
rect 292 -1780 298 -1754
rect -298 -1816 298 -1780
rect -298 -1842 -292 -1816
rect -266 -1842 -230 -1816
rect -204 -1842 -168 -1816
rect -142 -1842 -106 -1816
rect -80 -1842 -44 -1816
rect -18 -1842 18 -1816
rect 44 -1842 80 -1816
rect 106 -1842 142 -1816
rect 168 -1842 204 -1816
rect 230 -1842 266 -1816
rect 292 -1842 298 -1816
rect -298 -1878 298 -1842
rect -298 -1904 -292 -1878
rect -266 -1904 -230 -1878
rect -204 -1904 -168 -1878
rect -142 -1904 -106 -1878
rect -80 -1904 -44 -1878
rect -18 -1904 18 -1878
rect 44 -1904 80 -1878
rect 106 -1904 142 -1878
rect 168 -1904 204 -1878
rect 230 -1904 266 -1878
rect 292 -1904 298 -1878
rect -298 -1940 298 -1904
rect -298 -1966 -292 -1940
rect -266 -1966 -230 -1940
rect -204 -1966 -168 -1940
rect -142 -1966 -106 -1940
rect -80 -1966 -44 -1940
rect -18 -1966 18 -1940
rect 44 -1966 80 -1940
rect 106 -1966 142 -1940
rect 168 -1966 204 -1940
rect 230 -1966 266 -1940
rect 292 -1966 298 -1940
rect -298 -1972 298 -1966
<< via1 >>
rect -292 1940 -266 1966
rect -230 1940 -204 1966
rect -168 1940 -142 1966
rect -106 1940 -80 1966
rect -44 1940 -18 1966
rect 18 1940 44 1966
rect 80 1940 106 1966
rect 142 1940 168 1966
rect 204 1940 230 1966
rect 266 1940 292 1966
rect -292 1878 -266 1904
rect -230 1878 -204 1904
rect -168 1878 -142 1904
rect -106 1878 -80 1904
rect -44 1878 -18 1904
rect 18 1878 44 1904
rect 80 1878 106 1904
rect 142 1878 168 1904
rect 204 1878 230 1904
rect 266 1878 292 1904
rect -292 1816 -266 1842
rect -230 1816 -204 1842
rect -168 1816 -142 1842
rect -106 1816 -80 1842
rect -44 1816 -18 1842
rect 18 1816 44 1842
rect 80 1816 106 1842
rect 142 1816 168 1842
rect 204 1816 230 1842
rect 266 1816 292 1842
rect -292 1754 -266 1780
rect -230 1754 -204 1780
rect -168 1754 -142 1780
rect -106 1754 -80 1780
rect -44 1754 -18 1780
rect 18 1754 44 1780
rect 80 1754 106 1780
rect 142 1754 168 1780
rect 204 1754 230 1780
rect 266 1754 292 1780
rect -292 1692 -266 1718
rect -230 1692 -204 1718
rect -168 1692 -142 1718
rect -106 1692 -80 1718
rect -44 1692 -18 1718
rect 18 1692 44 1718
rect 80 1692 106 1718
rect 142 1692 168 1718
rect 204 1692 230 1718
rect 266 1692 292 1718
rect -292 1630 -266 1656
rect -230 1630 -204 1656
rect -168 1630 -142 1656
rect -106 1630 -80 1656
rect -44 1630 -18 1656
rect 18 1630 44 1656
rect 80 1630 106 1656
rect 142 1630 168 1656
rect 204 1630 230 1656
rect 266 1630 292 1656
rect -292 1568 -266 1594
rect -230 1568 -204 1594
rect -168 1568 -142 1594
rect -106 1568 -80 1594
rect -44 1568 -18 1594
rect 18 1568 44 1594
rect 80 1568 106 1594
rect 142 1568 168 1594
rect 204 1568 230 1594
rect 266 1568 292 1594
rect -292 1506 -266 1532
rect -230 1506 -204 1532
rect -168 1506 -142 1532
rect -106 1506 -80 1532
rect -44 1506 -18 1532
rect 18 1506 44 1532
rect 80 1506 106 1532
rect 142 1506 168 1532
rect 204 1506 230 1532
rect 266 1506 292 1532
rect -292 1444 -266 1470
rect -230 1444 -204 1470
rect -168 1444 -142 1470
rect -106 1444 -80 1470
rect -44 1444 -18 1470
rect 18 1444 44 1470
rect 80 1444 106 1470
rect 142 1444 168 1470
rect 204 1444 230 1470
rect 266 1444 292 1470
rect -292 1382 -266 1408
rect -230 1382 -204 1408
rect -168 1382 -142 1408
rect -106 1382 -80 1408
rect -44 1382 -18 1408
rect 18 1382 44 1408
rect 80 1382 106 1408
rect 142 1382 168 1408
rect 204 1382 230 1408
rect 266 1382 292 1408
rect -292 1320 -266 1346
rect -230 1320 -204 1346
rect -168 1320 -142 1346
rect -106 1320 -80 1346
rect -44 1320 -18 1346
rect 18 1320 44 1346
rect 80 1320 106 1346
rect 142 1320 168 1346
rect 204 1320 230 1346
rect 266 1320 292 1346
rect -292 1258 -266 1284
rect -230 1258 -204 1284
rect -168 1258 -142 1284
rect -106 1258 -80 1284
rect -44 1258 -18 1284
rect 18 1258 44 1284
rect 80 1258 106 1284
rect 142 1258 168 1284
rect 204 1258 230 1284
rect 266 1258 292 1284
rect -292 1196 -266 1222
rect -230 1196 -204 1222
rect -168 1196 -142 1222
rect -106 1196 -80 1222
rect -44 1196 -18 1222
rect 18 1196 44 1222
rect 80 1196 106 1222
rect 142 1196 168 1222
rect 204 1196 230 1222
rect 266 1196 292 1222
rect -292 1134 -266 1160
rect -230 1134 -204 1160
rect -168 1134 -142 1160
rect -106 1134 -80 1160
rect -44 1134 -18 1160
rect 18 1134 44 1160
rect 80 1134 106 1160
rect 142 1134 168 1160
rect 204 1134 230 1160
rect 266 1134 292 1160
rect -292 1072 -266 1098
rect -230 1072 -204 1098
rect -168 1072 -142 1098
rect -106 1072 -80 1098
rect -44 1072 -18 1098
rect 18 1072 44 1098
rect 80 1072 106 1098
rect 142 1072 168 1098
rect 204 1072 230 1098
rect 266 1072 292 1098
rect -292 1010 -266 1036
rect -230 1010 -204 1036
rect -168 1010 -142 1036
rect -106 1010 -80 1036
rect -44 1010 -18 1036
rect 18 1010 44 1036
rect 80 1010 106 1036
rect 142 1010 168 1036
rect 204 1010 230 1036
rect 266 1010 292 1036
rect -292 948 -266 974
rect -230 948 -204 974
rect -168 948 -142 974
rect -106 948 -80 974
rect -44 948 -18 974
rect 18 948 44 974
rect 80 948 106 974
rect 142 948 168 974
rect 204 948 230 974
rect 266 948 292 974
rect -292 886 -266 912
rect -230 886 -204 912
rect -168 886 -142 912
rect -106 886 -80 912
rect -44 886 -18 912
rect 18 886 44 912
rect 80 886 106 912
rect 142 886 168 912
rect 204 886 230 912
rect 266 886 292 912
rect -292 824 -266 850
rect -230 824 -204 850
rect -168 824 -142 850
rect -106 824 -80 850
rect -44 824 -18 850
rect 18 824 44 850
rect 80 824 106 850
rect 142 824 168 850
rect 204 824 230 850
rect 266 824 292 850
rect -292 762 -266 788
rect -230 762 -204 788
rect -168 762 -142 788
rect -106 762 -80 788
rect -44 762 -18 788
rect 18 762 44 788
rect 80 762 106 788
rect 142 762 168 788
rect 204 762 230 788
rect 266 762 292 788
rect -292 700 -266 726
rect -230 700 -204 726
rect -168 700 -142 726
rect -106 700 -80 726
rect -44 700 -18 726
rect 18 700 44 726
rect 80 700 106 726
rect 142 700 168 726
rect 204 700 230 726
rect 266 700 292 726
rect -292 638 -266 664
rect -230 638 -204 664
rect -168 638 -142 664
rect -106 638 -80 664
rect -44 638 -18 664
rect 18 638 44 664
rect 80 638 106 664
rect 142 638 168 664
rect 204 638 230 664
rect 266 638 292 664
rect -292 576 -266 602
rect -230 576 -204 602
rect -168 576 -142 602
rect -106 576 -80 602
rect -44 576 -18 602
rect 18 576 44 602
rect 80 576 106 602
rect 142 576 168 602
rect 204 576 230 602
rect 266 576 292 602
rect -292 514 -266 540
rect -230 514 -204 540
rect -168 514 -142 540
rect -106 514 -80 540
rect -44 514 -18 540
rect 18 514 44 540
rect 80 514 106 540
rect 142 514 168 540
rect 204 514 230 540
rect 266 514 292 540
rect -292 452 -266 478
rect -230 452 -204 478
rect -168 452 -142 478
rect -106 452 -80 478
rect -44 452 -18 478
rect 18 452 44 478
rect 80 452 106 478
rect 142 452 168 478
rect 204 452 230 478
rect 266 452 292 478
rect -292 390 -266 416
rect -230 390 -204 416
rect -168 390 -142 416
rect -106 390 -80 416
rect -44 390 -18 416
rect 18 390 44 416
rect 80 390 106 416
rect 142 390 168 416
rect 204 390 230 416
rect 266 390 292 416
rect -292 328 -266 354
rect -230 328 -204 354
rect -168 328 -142 354
rect -106 328 -80 354
rect -44 328 -18 354
rect 18 328 44 354
rect 80 328 106 354
rect 142 328 168 354
rect 204 328 230 354
rect 266 328 292 354
rect -292 266 -266 292
rect -230 266 -204 292
rect -168 266 -142 292
rect -106 266 -80 292
rect -44 266 -18 292
rect 18 266 44 292
rect 80 266 106 292
rect 142 266 168 292
rect 204 266 230 292
rect 266 266 292 292
rect -292 204 -266 230
rect -230 204 -204 230
rect -168 204 -142 230
rect -106 204 -80 230
rect -44 204 -18 230
rect 18 204 44 230
rect 80 204 106 230
rect 142 204 168 230
rect 204 204 230 230
rect 266 204 292 230
rect -292 142 -266 168
rect -230 142 -204 168
rect -168 142 -142 168
rect -106 142 -80 168
rect -44 142 -18 168
rect 18 142 44 168
rect 80 142 106 168
rect 142 142 168 168
rect 204 142 230 168
rect 266 142 292 168
rect -292 80 -266 106
rect -230 80 -204 106
rect -168 80 -142 106
rect -106 80 -80 106
rect -44 80 -18 106
rect 18 80 44 106
rect 80 80 106 106
rect 142 80 168 106
rect 204 80 230 106
rect 266 80 292 106
rect -292 18 -266 44
rect -230 18 -204 44
rect -168 18 -142 44
rect -106 18 -80 44
rect -44 18 -18 44
rect 18 18 44 44
rect 80 18 106 44
rect 142 18 168 44
rect 204 18 230 44
rect 266 18 292 44
rect -292 -44 -266 -18
rect -230 -44 -204 -18
rect -168 -44 -142 -18
rect -106 -44 -80 -18
rect -44 -44 -18 -18
rect 18 -44 44 -18
rect 80 -44 106 -18
rect 142 -44 168 -18
rect 204 -44 230 -18
rect 266 -44 292 -18
rect -292 -106 -266 -80
rect -230 -106 -204 -80
rect -168 -106 -142 -80
rect -106 -106 -80 -80
rect -44 -106 -18 -80
rect 18 -106 44 -80
rect 80 -106 106 -80
rect 142 -106 168 -80
rect 204 -106 230 -80
rect 266 -106 292 -80
rect -292 -168 -266 -142
rect -230 -168 -204 -142
rect -168 -168 -142 -142
rect -106 -168 -80 -142
rect -44 -168 -18 -142
rect 18 -168 44 -142
rect 80 -168 106 -142
rect 142 -168 168 -142
rect 204 -168 230 -142
rect 266 -168 292 -142
rect -292 -230 -266 -204
rect -230 -230 -204 -204
rect -168 -230 -142 -204
rect -106 -230 -80 -204
rect -44 -230 -18 -204
rect 18 -230 44 -204
rect 80 -230 106 -204
rect 142 -230 168 -204
rect 204 -230 230 -204
rect 266 -230 292 -204
rect -292 -292 -266 -266
rect -230 -292 -204 -266
rect -168 -292 -142 -266
rect -106 -292 -80 -266
rect -44 -292 -18 -266
rect 18 -292 44 -266
rect 80 -292 106 -266
rect 142 -292 168 -266
rect 204 -292 230 -266
rect 266 -292 292 -266
rect -292 -354 -266 -328
rect -230 -354 -204 -328
rect -168 -354 -142 -328
rect -106 -354 -80 -328
rect -44 -354 -18 -328
rect 18 -354 44 -328
rect 80 -354 106 -328
rect 142 -354 168 -328
rect 204 -354 230 -328
rect 266 -354 292 -328
rect -292 -416 -266 -390
rect -230 -416 -204 -390
rect -168 -416 -142 -390
rect -106 -416 -80 -390
rect -44 -416 -18 -390
rect 18 -416 44 -390
rect 80 -416 106 -390
rect 142 -416 168 -390
rect 204 -416 230 -390
rect 266 -416 292 -390
rect -292 -478 -266 -452
rect -230 -478 -204 -452
rect -168 -478 -142 -452
rect -106 -478 -80 -452
rect -44 -478 -18 -452
rect 18 -478 44 -452
rect 80 -478 106 -452
rect 142 -478 168 -452
rect 204 -478 230 -452
rect 266 -478 292 -452
rect -292 -540 -266 -514
rect -230 -540 -204 -514
rect -168 -540 -142 -514
rect -106 -540 -80 -514
rect -44 -540 -18 -514
rect 18 -540 44 -514
rect 80 -540 106 -514
rect 142 -540 168 -514
rect 204 -540 230 -514
rect 266 -540 292 -514
rect -292 -602 -266 -576
rect -230 -602 -204 -576
rect -168 -602 -142 -576
rect -106 -602 -80 -576
rect -44 -602 -18 -576
rect 18 -602 44 -576
rect 80 -602 106 -576
rect 142 -602 168 -576
rect 204 -602 230 -576
rect 266 -602 292 -576
rect -292 -664 -266 -638
rect -230 -664 -204 -638
rect -168 -664 -142 -638
rect -106 -664 -80 -638
rect -44 -664 -18 -638
rect 18 -664 44 -638
rect 80 -664 106 -638
rect 142 -664 168 -638
rect 204 -664 230 -638
rect 266 -664 292 -638
rect -292 -726 -266 -700
rect -230 -726 -204 -700
rect -168 -726 -142 -700
rect -106 -726 -80 -700
rect -44 -726 -18 -700
rect 18 -726 44 -700
rect 80 -726 106 -700
rect 142 -726 168 -700
rect 204 -726 230 -700
rect 266 -726 292 -700
rect -292 -788 -266 -762
rect -230 -788 -204 -762
rect -168 -788 -142 -762
rect -106 -788 -80 -762
rect -44 -788 -18 -762
rect 18 -788 44 -762
rect 80 -788 106 -762
rect 142 -788 168 -762
rect 204 -788 230 -762
rect 266 -788 292 -762
rect -292 -850 -266 -824
rect -230 -850 -204 -824
rect -168 -850 -142 -824
rect -106 -850 -80 -824
rect -44 -850 -18 -824
rect 18 -850 44 -824
rect 80 -850 106 -824
rect 142 -850 168 -824
rect 204 -850 230 -824
rect 266 -850 292 -824
rect -292 -912 -266 -886
rect -230 -912 -204 -886
rect -168 -912 -142 -886
rect -106 -912 -80 -886
rect -44 -912 -18 -886
rect 18 -912 44 -886
rect 80 -912 106 -886
rect 142 -912 168 -886
rect 204 -912 230 -886
rect 266 -912 292 -886
rect -292 -974 -266 -948
rect -230 -974 -204 -948
rect -168 -974 -142 -948
rect -106 -974 -80 -948
rect -44 -974 -18 -948
rect 18 -974 44 -948
rect 80 -974 106 -948
rect 142 -974 168 -948
rect 204 -974 230 -948
rect 266 -974 292 -948
rect -292 -1036 -266 -1010
rect -230 -1036 -204 -1010
rect -168 -1036 -142 -1010
rect -106 -1036 -80 -1010
rect -44 -1036 -18 -1010
rect 18 -1036 44 -1010
rect 80 -1036 106 -1010
rect 142 -1036 168 -1010
rect 204 -1036 230 -1010
rect 266 -1036 292 -1010
rect -292 -1098 -266 -1072
rect -230 -1098 -204 -1072
rect -168 -1098 -142 -1072
rect -106 -1098 -80 -1072
rect -44 -1098 -18 -1072
rect 18 -1098 44 -1072
rect 80 -1098 106 -1072
rect 142 -1098 168 -1072
rect 204 -1098 230 -1072
rect 266 -1098 292 -1072
rect -292 -1160 -266 -1134
rect -230 -1160 -204 -1134
rect -168 -1160 -142 -1134
rect -106 -1160 -80 -1134
rect -44 -1160 -18 -1134
rect 18 -1160 44 -1134
rect 80 -1160 106 -1134
rect 142 -1160 168 -1134
rect 204 -1160 230 -1134
rect 266 -1160 292 -1134
rect -292 -1222 -266 -1196
rect -230 -1222 -204 -1196
rect -168 -1222 -142 -1196
rect -106 -1222 -80 -1196
rect -44 -1222 -18 -1196
rect 18 -1222 44 -1196
rect 80 -1222 106 -1196
rect 142 -1222 168 -1196
rect 204 -1222 230 -1196
rect 266 -1222 292 -1196
rect -292 -1284 -266 -1258
rect -230 -1284 -204 -1258
rect -168 -1284 -142 -1258
rect -106 -1284 -80 -1258
rect -44 -1284 -18 -1258
rect 18 -1284 44 -1258
rect 80 -1284 106 -1258
rect 142 -1284 168 -1258
rect 204 -1284 230 -1258
rect 266 -1284 292 -1258
rect -292 -1346 -266 -1320
rect -230 -1346 -204 -1320
rect -168 -1346 -142 -1320
rect -106 -1346 -80 -1320
rect -44 -1346 -18 -1320
rect 18 -1346 44 -1320
rect 80 -1346 106 -1320
rect 142 -1346 168 -1320
rect 204 -1346 230 -1320
rect 266 -1346 292 -1320
rect -292 -1408 -266 -1382
rect -230 -1408 -204 -1382
rect -168 -1408 -142 -1382
rect -106 -1408 -80 -1382
rect -44 -1408 -18 -1382
rect 18 -1408 44 -1382
rect 80 -1408 106 -1382
rect 142 -1408 168 -1382
rect 204 -1408 230 -1382
rect 266 -1408 292 -1382
rect -292 -1470 -266 -1444
rect -230 -1470 -204 -1444
rect -168 -1470 -142 -1444
rect -106 -1470 -80 -1444
rect -44 -1470 -18 -1444
rect 18 -1470 44 -1444
rect 80 -1470 106 -1444
rect 142 -1470 168 -1444
rect 204 -1470 230 -1444
rect 266 -1470 292 -1444
rect -292 -1532 -266 -1506
rect -230 -1532 -204 -1506
rect -168 -1532 -142 -1506
rect -106 -1532 -80 -1506
rect -44 -1532 -18 -1506
rect 18 -1532 44 -1506
rect 80 -1532 106 -1506
rect 142 -1532 168 -1506
rect 204 -1532 230 -1506
rect 266 -1532 292 -1506
rect -292 -1594 -266 -1568
rect -230 -1594 -204 -1568
rect -168 -1594 -142 -1568
rect -106 -1594 -80 -1568
rect -44 -1594 -18 -1568
rect 18 -1594 44 -1568
rect 80 -1594 106 -1568
rect 142 -1594 168 -1568
rect 204 -1594 230 -1568
rect 266 -1594 292 -1568
rect -292 -1656 -266 -1630
rect -230 -1656 -204 -1630
rect -168 -1656 -142 -1630
rect -106 -1656 -80 -1630
rect -44 -1656 -18 -1630
rect 18 -1656 44 -1630
rect 80 -1656 106 -1630
rect 142 -1656 168 -1630
rect 204 -1656 230 -1630
rect 266 -1656 292 -1630
rect -292 -1718 -266 -1692
rect -230 -1718 -204 -1692
rect -168 -1718 -142 -1692
rect -106 -1718 -80 -1692
rect -44 -1718 -18 -1692
rect 18 -1718 44 -1692
rect 80 -1718 106 -1692
rect 142 -1718 168 -1692
rect 204 -1718 230 -1692
rect 266 -1718 292 -1692
rect -292 -1780 -266 -1754
rect -230 -1780 -204 -1754
rect -168 -1780 -142 -1754
rect -106 -1780 -80 -1754
rect -44 -1780 -18 -1754
rect 18 -1780 44 -1754
rect 80 -1780 106 -1754
rect 142 -1780 168 -1754
rect 204 -1780 230 -1754
rect 266 -1780 292 -1754
rect -292 -1842 -266 -1816
rect -230 -1842 -204 -1816
rect -168 -1842 -142 -1816
rect -106 -1842 -80 -1816
rect -44 -1842 -18 -1816
rect 18 -1842 44 -1816
rect 80 -1842 106 -1816
rect 142 -1842 168 -1816
rect 204 -1842 230 -1816
rect 266 -1842 292 -1816
rect -292 -1904 -266 -1878
rect -230 -1904 -204 -1878
rect -168 -1904 -142 -1878
rect -106 -1904 -80 -1878
rect -44 -1904 -18 -1878
rect 18 -1904 44 -1878
rect 80 -1904 106 -1878
rect 142 -1904 168 -1878
rect 204 -1904 230 -1878
rect 266 -1904 292 -1878
rect -292 -1966 -266 -1940
rect -230 -1966 -204 -1940
rect -168 -1966 -142 -1940
rect -106 -1966 -80 -1940
rect -44 -1966 -18 -1940
rect 18 -1966 44 -1940
rect 80 -1966 106 -1940
rect 142 -1966 168 -1940
rect 204 -1966 230 -1940
rect 266 -1966 292 -1940
<< metal2 >>
rect -298 1966 298 1972
rect -298 1940 -292 1966
rect -266 1940 -230 1966
rect -204 1940 -168 1966
rect -142 1940 -106 1966
rect -80 1940 -44 1966
rect -18 1940 18 1966
rect 44 1940 80 1966
rect 106 1940 142 1966
rect 168 1940 204 1966
rect 230 1940 266 1966
rect 292 1940 298 1966
rect -298 1904 298 1940
rect -298 1878 -292 1904
rect -266 1878 -230 1904
rect -204 1878 -168 1904
rect -142 1878 -106 1904
rect -80 1878 -44 1904
rect -18 1878 18 1904
rect 44 1878 80 1904
rect 106 1878 142 1904
rect 168 1878 204 1904
rect 230 1878 266 1904
rect 292 1878 298 1904
rect -298 1842 298 1878
rect -298 1816 -292 1842
rect -266 1816 -230 1842
rect -204 1816 -168 1842
rect -142 1816 -106 1842
rect -80 1816 -44 1842
rect -18 1816 18 1842
rect 44 1816 80 1842
rect 106 1816 142 1842
rect 168 1816 204 1842
rect 230 1816 266 1842
rect 292 1816 298 1842
rect -298 1780 298 1816
rect -298 1754 -292 1780
rect -266 1754 -230 1780
rect -204 1754 -168 1780
rect -142 1754 -106 1780
rect -80 1754 -44 1780
rect -18 1754 18 1780
rect 44 1754 80 1780
rect 106 1754 142 1780
rect 168 1754 204 1780
rect 230 1754 266 1780
rect 292 1754 298 1780
rect -298 1718 298 1754
rect -298 1692 -292 1718
rect -266 1692 -230 1718
rect -204 1692 -168 1718
rect -142 1692 -106 1718
rect -80 1692 -44 1718
rect -18 1692 18 1718
rect 44 1692 80 1718
rect 106 1692 142 1718
rect 168 1692 204 1718
rect 230 1692 266 1718
rect 292 1692 298 1718
rect -298 1656 298 1692
rect -298 1630 -292 1656
rect -266 1630 -230 1656
rect -204 1630 -168 1656
rect -142 1630 -106 1656
rect -80 1630 -44 1656
rect -18 1630 18 1656
rect 44 1630 80 1656
rect 106 1630 142 1656
rect 168 1630 204 1656
rect 230 1630 266 1656
rect 292 1630 298 1656
rect -298 1594 298 1630
rect -298 1568 -292 1594
rect -266 1568 -230 1594
rect -204 1568 -168 1594
rect -142 1568 -106 1594
rect -80 1568 -44 1594
rect -18 1568 18 1594
rect 44 1568 80 1594
rect 106 1568 142 1594
rect 168 1568 204 1594
rect 230 1568 266 1594
rect 292 1568 298 1594
rect -298 1532 298 1568
rect -298 1506 -292 1532
rect -266 1506 -230 1532
rect -204 1506 -168 1532
rect -142 1506 -106 1532
rect -80 1506 -44 1532
rect -18 1506 18 1532
rect 44 1506 80 1532
rect 106 1506 142 1532
rect 168 1506 204 1532
rect 230 1506 266 1532
rect 292 1506 298 1532
rect -298 1470 298 1506
rect -298 1444 -292 1470
rect -266 1444 -230 1470
rect -204 1444 -168 1470
rect -142 1444 -106 1470
rect -80 1444 -44 1470
rect -18 1444 18 1470
rect 44 1444 80 1470
rect 106 1444 142 1470
rect 168 1444 204 1470
rect 230 1444 266 1470
rect 292 1444 298 1470
rect -298 1408 298 1444
rect -298 1382 -292 1408
rect -266 1382 -230 1408
rect -204 1382 -168 1408
rect -142 1382 -106 1408
rect -80 1382 -44 1408
rect -18 1382 18 1408
rect 44 1382 80 1408
rect 106 1382 142 1408
rect 168 1382 204 1408
rect 230 1382 266 1408
rect 292 1382 298 1408
rect -298 1346 298 1382
rect -298 1320 -292 1346
rect -266 1320 -230 1346
rect -204 1320 -168 1346
rect -142 1320 -106 1346
rect -80 1320 -44 1346
rect -18 1320 18 1346
rect 44 1320 80 1346
rect 106 1320 142 1346
rect 168 1320 204 1346
rect 230 1320 266 1346
rect 292 1320 298 1346
rect -298 1284 298 1320
rect -298 1258 -292 1284
rect -266 1258 -230 1284
rect -204 1258 -168 1284
rect -142 1258 -106 1284
rect -80 1258 -44 1284
rect -18 1258 18 1284
rect 44 1258 80 1284
rect 106 1258 142 1284
rect 168 1258 204 1284
rect 230 1258 266 1284
rect 292 1258 298 1284
rect -298 1222 298 1258
rect -298 1196 -292 1222
rect -266 1196 -230 1222
rect -204 1196 -168 1222
rect -142 1196 -106 1222
rect -80 1196 -44 1222
rect -18 1196 18 1222
rect 44 1196 80 1222
rect 106 1196 142 1222
rect 168 1196 204 1222
rect 230 1196 266 1222
rect 292 1196 298 1222
rect -298 1160 298 1196
rect -298 1134 -292 1160
rect -266 1134 -230 1160
rect -204 1134 -168 1160
rect -142 1134 -106 1160
rect -80 1134 -44 1160
rect -18 1134 18 1160
rect 44 1134 80 1160
rect 106 1134 142 1160
rect 168 1134 204 1160
rect 230 1134 266 1160
rect 292 1134 298 1160
rect -298 1098 298 1134
rect -298 1072 -292 1098
rect -266 1072 -230 1098
rect -204 1072 -168 1098
rect -142 1072 -106 1098
rect -80 1072 -44 1098
rect -18 1072 18 1098
rect 44 1072 80 1098
rect 106 1072 142 1098
rect 168 1072 204 1098
rect 230 1072 266 1098
rect 292 1072 298 1098
rect -298 1036 298 1072
rect -298 1010 -292 1036
rect -266 1010 -230 1036
rect -204 1010 -168 1036
rect -142 1010 -106 1036
rect -80 1010 -44 1036
rect -18 1010 18 1036
rect 44 1010 80 1036
rect 106 1010 142 1036
rect 168 1010 204 1036
rect 230 1010 266 1036
rect 292 1010 298 1036
rect -298 974 298 1010
rect -298 948 -292 974
rect -266 948 -230 974
rect -204 948 -168 974
rect -142 948 -106 974
rect -80 948 -44 974
rect -18 948 18 974
rect 44 948 80 974
rect 106 948 142 974
rect 168 948 204 974
rect 230 948 266 974
rect 292 948 298 974
rect -298 912 298 948
rect -298 886 -292 912
rect -266 886 -230 912
rect -204 886 -168 912
rect -142 886 -106 912
rect -80 886 -44 912
rect -18 886 18 912
rect 44 886 80 912
rect 106 886 142 912
rect 168 886 204 912
rect 230 886 266 912
rect 292 886 298 912
rect -298 850 298 886
rect -298 824 -292 850
rect -266 824 -230 850
rect -204 824 -168 850
rect -142 824 -106 850
rect -80 824 -44 850
rect -18 824 18 850
rect 44 824 80 850
rect 106 824 142 850
rect 168 824 204 850
rect 230 824 266 850
rect 292 824 298 850
rect -298 788 298 824
rect -298 762 -292 788
rect -266 762 -230 788
rect -204 762 -168 788
rect -142 762 -106 788
rect -80 762 -44 788
rect -18 762 18 788
rect 44 762 80 788
rect 106 762 142 788
rect 168 762 204 788
rect 230 762 266 788
rect 292 762 298 788
rect -298 726 298 762
rect -298 700 -292 726
rect -266 700 -230 726
rect -204 700 -168 726
rect -142 700 -106 726
rect -80 700 -44 726
rect -18 700 18 726
rect 44 700 80 726
rect 106 700 142 726
rect 168 700 204 726
rect 230 700 266 726
rect 292 700 298 726
rect -298 664 298 700
rect -298 638 -292 664
rect -266 638 -230 664
rect -204 638 -168 664
rect -142 638 -106 664
rect -80 638 -44 664
rect -18 638 18 664
rect 44 638 80 664
rect 106 638 142 664
rect 168 638 204 664
rect 230 638 266 664
rect 292 638 298 664
rect -298 602 298 638
rect -298 576 -292 602
rect -266 576 -230 602
rect -204 576 -168 602
rect -142 576 -106 602
rect -80 576 -44 602
rect -18 576 18 602
rect 44 576 80 602
rect 106 576 142 602
rect 168 576 204 602
rect 230 576 266 602
rect 292 576 298 602
rect -298 540 298 576
rect -298 514 -292 540
rect -266 514 -230 540
rect -204 514 -168 540
rect -142 514 -106 540
rect -80 514 -44 540
rect -18 514 18 540
rect 44 514 80 540
rect 106 514 142 540
rect 168 514 204 540
rect 230 514 266 540
rect 292 514 298 540
rect -298 478 298 514
rect -298 452 -292 478
rect -266 452 -230 478
rect -204 452 -168 478
rect -142 452 -106 478
rect -80 452 -44 478
rect -18 452 18 478
rect 44 452 80 478
rect 106 452 142 478
rect 168 452 204 478
rect 230 452 266 478
rect 292 452 298 478
rect -298 416 298 452
rect -298 390 -292 416
rect -266 390 -230 416
rect -204 390 -168 416
rect -142 390 -106 416
rect -80 390 -44 416
rect -18 390 18 416
rect 44 390 80 416
rect 106 390 142 416
rect 168 390 204 416
rect 230 390 266 416
rect 292 390 298 416
rect -298 354 298 390
rect -298 328 -292 354
rect -266 328 -230 354
rect -204 328 -168 354
rect -142 328 -106 354
rect -80 328 -44 354
rect -18 328 18 354
rect 44 328 80 354
rect 106 328 142 354
rect 168 328 204 354
rect 230 328 266 354
rect 292 328 298 354
rect -298 292 298 328
rect -298 266 -292 292
rect -266 266 -230 292
rect -204 266 -168 292
rect -142 266 -106 292
rect -80 266 -44 292
rect -18 266 18 292
rect 44 266 80 292
rect 106 266 142 292
rect 168 266 204 292
rect 230 266 266 292
rect 292 266 298 292
rect -298 230 298 266
rect -298 204 -292 230
rect -266 204 -230 230
rect -204 204 -168 230
rect -142 204 -106 230
rect -80 204 -44 230
rect -18 204 18 230
rect 44 204 80 230
rect 106 204 142 230
rect 168 204 204 230
rect 230 204 266 230
rect 292 204 298 230
rect -298 168 298 204
rect -298 142 -292 168
rect -266 142 -230 168
rect -204 142 -168 168
rect -142 142 -106 168
rect -80 142 -44 168
rect -18 142 18 168
rect 44 142 80 168
rect 106 142 142 168
rect 168 142 204 168
rect 230 142 266 168
rect 292 142 298 168
rect -298 106 298 142
rect -298 80 -292 106
rect -266 80 -230 106
rect -204 80 -168 106
rect -142 80 -106 106
rect -80 80 -44 106
rect -18 80 18 106
rect 44 80 80 106
rect 106 80 142 106
rect 168 80 204 106
rect 230 80 266 106
rect 292 80 298 106
rect -298 44 298 80
rect -298 18 -292 44
rect -266 18 -230 44
rect -204 18 -168 44
rect -142 18 -106 44
rect -80 18 -44 44
rect -18 18 18 44
rect 44 18 80 44
rect 106 18 142 44
rect 168 18 204 44
rect 230 18 266 44
rect 292 18 298 44
rect -298 -18 298 18
rect -298 -44 -292 -18
rect -266 -44 -230 -18
rect -204 -44 -168 -18
rect -142 -44 -106 -18
rect -80 -44 -44 -18
rect -18 -44 18 -18
rect 44 -44 80 -18
rect 106 -44 142 -18
rect 168 -44 204 -18
rect 230 -44 266 -18
rect 292 -44 298 -18
rect -298 -80 298 -44
rect -298 -106 -292 -80
rect -266 -106 -230 -80
rect -204 -106 -168 -80
rect -142 -106 -106 -80
rect -80 -106 -44 -80
rect -18 -106 18 -80
rect 44 -106 80 -80
rect 106 -106 142 -80
rect 168 -106 204 -80
rect 230 -106 266 -80
rect 292 -106 298 -80
rect -298 -142 298 -106
rect -298 -168 -292 -142
rect -266 -168 -230 -142
rect -204 -168 -168 -142
rect -142 -168 -106 -142
rect -80 -168 -44 -142
rect -18 -168 18 -142
rect 44 -168 80 -142
rect 106 -168 142 -142
rect 168 -168 204 -142
rect 230 -168 266 -142
rect 292 -168 298 -142
rect -298 -204 298 -168
rect -298 -230 -292 -204
rect -266 -230 -230 -204
rect -204 -230 -168 -204
rect -142 -230 -106 -204
rect -80 -230 -44 -204
rect -18 -230 18 -204
rect 44 -230 80 -204
rect 106 -230 142 -204
rect 168 -230 204 -204
rect 230 -230 266 -204
rect 292 -230 298 -204
rect -298 -266 298 -230
rect -298 -292 -292 -266
rect -266 -292 -230 -266
rect -204 -292 -168 -266
rect -142 -292 -106 -266
rect -80 -292 -44 -266
rect -18 -292 18 -266
rect 44 -292 80 -266
rect 106 -292 142 -266
rect 168 -292 204 -266
rect 230 -292 266 -266
rect 292 -292 298 -266
rect -298 -328 298 -292
rect -298 -354 -292 -328
rect -266 -354 -230 -328
rect -204 -354 -168 -328
rect -142 -354 -106 -328
rect -80 -354 -44 -328
rect -18 -354 18 -328
rect 44 -354 80 -328
rect 106 -354 142 -328
rect 168 -354 204 -328
rect 230 -354 266 -328
rect 292 -354 298 -328
rect -298 -390 298 -354
rect -298 -416 -292 -390
rect -266 -416 -230 -390
rect -204 -416 -168 -390
rect -142 -416 -106 -390
rect -80 -416 -44 -390
rect -18 -416 18 -390
rect 44 -416 80 -390
rect 106 -416 142 -390
rect 168 -416 204 -390
rect 230 -416 266 -390
rect 292 -416 298 -390
rect -298 -452 298 -416
rect -298 -478 -292 -452
rect -266 -478 -230 -452
rect -204 -478 -168 -452
rect -142 -478 -106 -452
rect -80 -478 -44 -452
rect -18 -478 18 -452
rect 44 -478 80 -452
rect 106 -478 142 -452
rect 168 -478 204 -452
rect 230 -478 266 -452
rect 292 -478 298 -452
rect -298 -514 298 -478
rect -298 -540 -292 -514
rect -266 -540 -230 -514
rect -204 -540 -168 -514
rect -142 -540 -106 -514
rect -80 -540 -44 -514
rect -18 -540 18 -514
rect 44 -540 80 -514
rect 106 -540 142 -514
rect 168 -540 204 -514
rect 230 -540 266 -514
rect 292 -540 298 -514
rect -298 -576 298 -540
rect -298 -602 -292 -576
rect -266 -602 -230 -576
rect -204 -602 -168 -576
rect -142 -602 -106 -576
rect -80 -602 -44 -576
rect -18 -602 18 -576
rect 44 -602 80 -576
rect 106 -602 142 -576
rect 168 -602 204 -576
rect 230 -602 266 -576
rect 292 -602 298 -576
rect -298 -638 298 -602
rect -298 -664 -292 -638
rect -266 -664 -230 -638
rect -204 -664 -168 -638
rect -142 -664 -106 -638
rect -80 -664 -44 -638
rect -18 -664 18 -638
rect 44 -664 80 -638
rect 106 -664 142 -638
rect 168 -664 204 -638
rect 230 -664 266 -638
rect 292 -664 298 -638
rect -298 -700 298 -664
rect -298 -726 -292 -700
rect -266 -726 -230 -700
rect -204 -726 -168 -700
rect -142 -726 -106 -700
rect -80 -726 -44 -700
rect -18 -726 18 -700
rect 44 -726 80 -700
rect 106 -726 142 -700
rect 168 -726 204 -700
rect 230 -726 266 -700
rect 292 -726 298 -700
rect -298 -762 298 -726
rect -298 -788 -292 -762
rect -266 -788 -230 -762
rect -204 -788 -168 -762
rect -142 -788 -106 -762
rect -80 -788 -44 -762
rect -18 -788 18 -762
rect 44 -788 80 -762
rect 106 -788 142 -762
rect 168 -788 204 -762
rect 230 -788 266 -762
rect 292 -788 298 -762
rect -298 -824 298 -788
rect -298 -850 -292 -824
rect -266 -850 -230 -824
rect -204 -850 -168 -824
rect -142 -850 -106 -824
rect -80 -850 -44 -824
rect -18 -850 18 -824
rect 44 -850 80 -824
rect 106 -850 142 -824
rect 168 -850 204 -824
rect 230 -850 266 -824
rect 292 -850 298 -824
rect -298 -886 298 -850
rect -298 -912 -292 -886
rect -266 -912 -230 -886
rect -204 -912 -168 -886
rect -142 -912 -106 -886
rect -80 -912 -44 -886
rect -18 -912 18 -886
rect 44 -912 80 -886
rect 106 -912 142 -886
rect 168 -912 204 -886
rect 230 -912 266 -886
rect 292 -912 298 -886
rect -298 -948 298 -912
rect -298 -974 -292 -948
rect -266 -974 -230 -948
rect -204 -974 -168 -948
rect -142 -974 -106 -948
rect -80 -974 -44 -948
rect -18 -974 18 -948
rect 44 -974 80 -948
rect 106 -974 142 -948
rect 168 -974 204 -948
rect 230 -974 266 -948
rect 292 -974 298 -948
rect -298 -1010 298 -974
rect -298 -1036 -292 -1010
rect -266 -1036 -230 -1010
rect -204 -1036 -168 -1010
rect -142 -1036 -106 -1010
rect -80 -1036 -44 -1010
rect -18 -1036 18 -1010
rect 44 -1036 80 -1010
rect 106 -1036 142 -1010
rect 168 -1036 204 -1010
rect 230 -1036 266 -1010
rect 292 -1036 298 -1010
rect -298 -1072 298 -1036
rect -298 -1098 -292 -1072
rect -266 -1098 -230 -1072
rect -204 -1098 -168 -1072
rect -142 -1098 -106 -1072
rect -80 -1098 -44 -1072
rect -18 -1098 18 -1072
rect 44 -1098 80 -1072
rect 106 -1098 142 -1072
rect 168 -1098 204 -1072
rect 230 -1098 266 -1072
rect 292 -1098 298 -1072
rect -298 -1134 298 -1098
rect -298 -1160 -292 -1134
rect -266 -1160 -230 -1134
rect -204 -1160 -168 -1134
rect -142 -1160 -106 -1134
rect -80 -1160 -44 -1134
rect -18 -1160 18 -1134
rect 44 -1160 80 -1134
rect 106 -1160 142 -1134
rect 168 -1160 204 -1134
rect 230 -1160 266 -1134
rect 292 -1160 298 -1134
rect -298 -1196 298 -1160
rect -298 -1222 -292 -1196
rect -266 -1222 -230 -1196
rect -204 -1222 -168 -1196
rect -142 -1222 -106 -1196
rect -80 -1222 -44 -1196
rect -18 -1222 18 -1196
rect 44 -1222 80 -1196
rect 106 -1222 142 -1196
rect 168 -1222 204 -1196
rect 230 -1222 266 -1196
rect 292 -1222 298 -1196
rect -298 -1258 298 -1222
rect -298 -1284 -292 -1258
rect -266 -1284 -230 -1258
rect -204 -1284 -168 -1258
rect -142 -1284 -106 -1258
rect -80 -1284 -44 -1258
rect -18 -1284 18 -1258
rect 44 -1284 80 -1258
rect 106 -1284 142 -1258
rect 168 -1284 204 -1258
rect 230 -1284 266 -1258
rect 292 -1284 298 -1258
rect -298 -1320 298 -1284
rect -298 -1346 -292 -1320
rect -266 -1346 -230 -1320
rect -204 -1346 -168 -1320
rect -142 -1346 -106 -1320
rect -80 -1346 -44 -1320
rect -18 -1346 18 -1320
rect 44 -1346 80 -1320
rect 106 -1346 142 -1320
rect 168 -1346 204 -1320
rect 230 -1346 266 -1320
rect 292 -1346 298 -1320
rect -298 -1382 298 -1346
rect -298 -1408 -292 -1382
rect -266 -1408 -230 -1382
rect -204 -1408 -168 -1382
rect -142 -1408 -106 -1382
rect -80 -1408 -44 -1382
rect -18 -1408 18 -1382
rect 44 -1408 80 -1382
rect 106 -1408 142 -1382
rect 168 -1408 204 -1382
rect 230 -1408 266 -1382
rect 292 -1408 298 -1382
rect -298 -1444 298 -1408
rect -298 -1470 -292 -1444
rect -266 -1470 -230 -1444
rect -204 -1470 -168 -1444
rect -142 -1470 -106 -1444
rect -80 -1470 -44 -1444
rect -18 -1470 18 -1444
rect 44 -1470 80 -1444
rect 106 -1470 142 -1444
rect 168 -1470 204 -1444
rect 230 -1470 266 -1444
rect 292 -1470 298 -1444
rect -298 -1506 298 -1470
rect -298 -1532 -292 -1506
rect -266 -1532 -230 -1506
rect -204 -1532 -168 -1506
rect -142 -1532 -106 -1506
rect -80 -1532 -44 -1506
rect -18 -1532 18 -1506
rect 44 -1532 80 -1506
rect 106 -1532 142 -1506
rect 168 -1532 204 -1506
rect 230 -1532 266 -1506
rect 292 -1532 298 -1506
rect -298 -1568 298 -1532
rect -298 -1594 -292 -1568
rect -266 -1594 -230 -1568
rect -204 -1594 -168 -1568
rect -142 -1594 -106 -1568
rect -80 -1594 -44 -1568
rect -18 -1594 18 -1568
rect 44 -1594 80 -1568
rect 106 -1594 142 -1568
rect 168 -1594 204 -1568
rect 230 -1594 266 -1568
rect 292 -1594 298 -1568
rect -298 -1630 298 -1594
rect -298 -1656 -292 -1630
rect -266 -1656 -230 -1630
rect -204 -1656 -168 -1630
rect -142 -1656 -106 -1630
rect -80 -1656 -44 -1630
rect -18 -1656 18 -1630
rect 44 -1656 80 -1630
rect 106 -1656 142 -1630
rect 168 -1656 204 -1630
rect 230 -1656 266 -1630
rect 292 -1656 298 -1630
rect -298 -1692 298 -1656
rect -298 -1718 -292 -1692
rect -266 -1718 -230 -1692
rect -204 -1718 -168 -1692
rect -142 -1718 -106 -1692
rect -80 -1718 -44 -1692
rect -18 -1718 18 -1692
rect 44 -1718 80 -1692
rect 106 -1718 142 -1692
rect 168 -1718 204 -1692
rect 230 -1718 266 -1692
rect 292 -1718 298 -1692
rect -298 -1754 298 -1718
rect -298 -1780 -292 -1754
rect -266 -1780 -230 -1754
rect -204 -1780 -168 -1754
rect -142 -1780 -106 -1754
rect -80 -1780 -44 -1754
rect -18 -1780 18 -1754
rect 44 -1780 80 -1754
rect 106 -1780 142 -1754
rect 168 -1780 204 -1754
rect 230 -1780 266 -1754
rect 292 -1780 298 -1754
rect -298 -1816 298 -1780
rect -298 -1842 -292 -1816
rect -266 -1842 -230 -1816
rect -204 -1842 -168 -1816
rect -142 -1842 -106 -1816
rect -80 -1842 -44 -1816
rect -18 -1842 18 -1816
rect 44 -1842 80 -1816
rect 106 -1842 142 -1816
rect 168 -1842 204 -1816
rect 230 -1842 266 -1816
rect 292 -1842 298 -1816
rect -298 -1878 298 -1842
rect -298 -1904 -292 -1878
rect -266 -1904 -230 -1878
rect -204 -1904 -168 -1878
rect -142 -1904 -106 -1878
rect -80 -1904 -44 -1878
rect -18 -1904 18 -1878
rect 44 -1904 80 -1878
rect 106 -1904 142 -1878
rect 168 -1904 204 -1878
rect 230 -1904 266 -1878
rect 292 -1904 298 -1878
rect -298 -1940 298 -1904
rect -298 -1966 -292 -1940
rect -266 -1966 -230 -1940
rect -204 -1966 -168 -1940
rect -142 -1966 -106 -1940
rect -80 -1966 -44 -1940
rect -18 -1966 18 -1940
rect 44 -1966 80 -1940
rect 106 -1966 142 -1940
rect 168 -1966 204 -1940
rect 230 -1966 266 -1940
rect 292 -1966 298 -1940
rect -298 -1972 298 -1966
<< end >>
