magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2088 -2044 2228 2344
<< mvnmos >>
rect 0 0 140 300
<< mvndiff >>
rect -88 287 0 300
rect -88 241 -75 287
rect -29 241 0 287
rect -88 173 0 241
rect -88 127 -75 173
rect -29 127 0 173
rect -88 59 0 127
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 140 287 228 300
rect 140 241 169 287
rect 215 241 228 287
rect 140 173 228 241
rect 140 127 169 173
rect 215 127 228 173
rect 140 59 228 127
rect 140 13 169 59
rect 215 13 228 59
rect 140 0 228 13
<< mvndiffc >>
rect -75 241 -29 287
rect -75 127 -29 173
rect -75 13 -29 59
rect 169 241 215 287
rect 169 127 215 173
rect 169 13 215 59
<< polysilicon >>
rect 0 300 140 344
rect 0 -44 140 0
<< metal1 >>
rect -75 287 -29 300
rect -75 173 -29 241
rect -75 59 -29 127
rect -75 0 -29 13
rect 169 287 215 300
rect 169 173 215 241
rect 169 59 215 127
rect 169 0 215 13
<< labels >>
rlabel mvndiffc 192 150 192 150 4 D
rlabel mvndiffc -52 150 -52 150 4 S
<< end >>
