magic
tech gf180mcuC
magscale 1 10
timestamp 1699521709
<< metal1 >>
rect 2272 1553 2348 1565
rect 2272 1501 2284 1553
rect 2336 1550 2348 1553
rect 2336 1504 2799 1550
rect 2336 1501 2348 1504
rect 2272 1489 2348 1501
rect 690 1446 766 1458
rect 690 1443 702 1446
rect 377 1397 702 1443
rect 690 1394 702 1397
rect 754 1394 766 1446
rect 690 1382 766 1394
rect 2395 1446 2471 1458
rect 2395 1394 2407 1446
rect 2459 1443 2471 1446
rect 2459 1397 2799 1443
rect 2459 1394 2471 1397
rect 2395 1382 2471 1394
rect 554 1339 630 1351
rect 554 1336 566 1339
rect 377 1290 566 1336
rect 554 1287 566 1290
rect 618 1287 630 1339
rect 554 1275 630 1287
rect 2518 1339 2594 1351
rect 2518 1287 2530 1339
rect 2582 1336 2594 1339
rect 2582 1290 2799 1336
rect 2582 1287 2594 1290
rect 2518 1275 2594 1287
rect 2654 1232 2730 1244
rect 2654 1229 2666 1232
rect 377 1183 2666 1229
rect 2654 1180 2666 1183
rect 2718 1180 2730 1232
rect 2654 1168 2730 1180
rect 69 1092 1249 1122
rect 69 1040 99 1092
rect 151 1040 1249 1092
rect 69 1010 1249 1040
rect 1812 1010 3578 1122
rect 2272 798 2348 810
rect 2272 746 2284 798
rect 2336 746 2348 798
rect 4896 749 5362 795
rect 2272 734 2348 746
rect 2652 703 2733 715
rect 237 678 313 690
rect 237 626 249 678
rect 301 626 313 678
rect 688 647 700 703
rect 756 647 1039 703
rect 2652 647 2664 703
rect 2720 647 3436 703
rect 688 635 768 647
rect 2652 635 2733 647
rect 237 614 313 626
rect 682 558 762 570
rect 682 548 694 558
rect 414 502 694 548
rect 750 502 762 558
rect 682 490 762 502
rect -99 237 205 267
rect 2651 251 2732 263
rect 5056 251 5132 261
rect -99 185 -69 237
rect -17 185 205 237
rect -99 155 205 185
rect 552 222 632 234
rect 1082 222 1158 234
rect 552 166 564 222
rect 620 170 1094 222
rect 1146 170 1324 222
rect 2389 195 2663 251
rect 2719 195 2732 251
rect 4882 249 5132 251
rect 2651 183 2732 195
rect 620 166 1324 170
rect 4882 197 5067 249
rect 5119 197 5132 249
rect 4882 195 5132 197
rect 5056 185 5132 195
rect 552 154 632 166
rect 1082 158 1158 166
rect 2225 0 3326 112
rect 552 -54 632 -42
rect 2914 -54 2990 -46
rect 552 -80 564 -54
rect 414 -110 564 -80
rect 620 -110 1274 -54
rect 2914 -58 3720 -54
rect 2780 -83 2860 -71
rect 414 -122 632 -110
rect 414 -126 582 -122
rect 2475 -139 2792 -83
rect 2848 -139 2860 -83
rect 2914 -110 2926 -58
rect 2978 -110 3720 -58
rect 4755 -84 4835 -72
rect 2914 -122 2990 -110
rect 2780 -151 2860 -139
rect 4755 -140 4767 -84
rect 4823 -140 4835 -84
rect 4755 -152 4835 -140
rect 237 -208 313 -196
rect 237 -260 249 -208
rect 301 -260 313 -208
rect 237 -272 313 -260
rect 688 -535 768 -523
rect 2782 -532 2858 -520
rect 69 -618 181 -588
rect 688 -591 700 -535
rect 756 -591 1051 -535
rect 688 -603 768 -591
rect 2782 -594 2794 -532
rect 2846 -535 2858 -532
rect 2846 -591 3431 -535
rect 2846 -594 2858 -591
rect 2782 -606 2858 -594
rect 69 -670 99 -618
rect 151 -670 181 -618
rect 69 -700 181 -670
rect 2395 -634 2471 -622
rect 2395 -686 2407 -634
rect 2459 -686 2471 -634
rect 4896 -683 5362 -637
rect 2395 -698 2471 -686
rect 1812 -1010 2913 -898
rect 235 -1026 315 -1014
rect 235 -1082 247 -1026
rect 303 -1082 315 -1026
rect 235 -1094 315 -1082
rect 427 -1151 507 -1139
rect 427 -1207 439 -1151
rect 495 -1207 507 -1151
rect 427 -1219 507 -1207
rect 2516 -1220 2596 -1208
rect 2516 -1276 2528 -1220
rect 2584 -1276 2596 -1220
rect 5162 -1276 5362 -1230
rect 2516 -1288 2596 -1276
rect 688 -1317 768 -1305
rect 688 -1373 700 -1317
rect 756 -1373 984 -1317
rect 688 -1385 768 -1373
rect -99 -1471 505 -1441
rect -99 -1523 -69 -1471
rect -17 -1523 505 -1471
rect -99 -1553 505 -1523
rect 393 -1908 505 -1553
rect 2915 -1489 2993 -1478
rect 3954 -1488 4196 -1442
rect 2915 -1490 3066 -1489
rect 2915 -1544 2927 -1490
rect 2979 -1544 3066 -1490
rect 2915 -1545 3066 -1544
rect 2915 -1556 2993 -1545
rect 2652 -1769 2732 -1757
rect 2485 -1825 2664 -1769
rect 2720 -1825 2732 -1769
rect 2652 -1837 2732 -1825
rect 2782 -1804 2858 -1792
rect 2782 -1856 2794 -1804
rect 2846 -1811 2858 -1804
rect 2846 -1856 3039 -1811
rect 2782 -1857 3039 -1856
rect 2782 -1868 2858 -1857
rect 393 -2020 806 -1908
rect 2492 -2020 3135 -1914
rect 3735 -2026 4836 -1914
<< via1 >>
rect 2284 1501 2336 1553
rect 702 1394 754 1446
rect 2407 1394 2459 1446
rect 566 1287 618 1339
rect 2530 1287 2582 1339
rect 2666 1180 2718 1232
rect 99 1040 151 1092
rect 1611 1040 1663 1092
rect 2284 746 2336 798
rect 249 626 301 678
rect 700 647 756 703
rect 2664 647 2720 703
rect 694 502 750 558
rect -69 185 -17 237
rect 564 166 620 222
rect 1094 170 1146 222
rect 2663 195 2719 251
rect 3744 169 3796 221
rect 5067 197 5119 249
rect 2033 30 2085 82
rect 564 -110 620 -54
rect 2792 -139 2848 -83
rect 2926 -110 2978 -58
rect 4767 -140 4823 -84
rect 249 -260 301 -208
rect 700 -591 756 -535
rect 2794 -594 2846 -532
rect 99 -670 151 -618
rect 2407 -686 2459 -634
rect 1611 -980 1663 -928
rect 247 -1082 303 -1026
rect 439 -1207 495 -1151
rect 2528 -1276 2584 -1220
rect 700 -1373 756 -1317
rect -69 -1523 -17 -1471
rect 2927 -1544 2979 -1490
rect 1361 -1851 1413 -1799
rect 2664 -1825 2720 -1769
rect 2794 -1856 2846 -1804
rect 5067 -1846 5119 -1794
rect 2033 -1990 2085 -1938
<< metal2 >>
rect 2272 1553 2348 1565
rect 2272 1501 2284 1553
rect 2336 1501 2348 1553
rect 2272 1489 2348 1501
rect 690 1446 766 1458
rect 690 1394 702 1446
rect 754 1394 766 1446
rect 690 1382 766 1394
rect 554 1339 630 1351
rect 554 1287 566 1339
rect 618 1287 630 1339
rect 554 1275 630 1287
rect 69 1092 181 1122
rect 69 1040 99 1092
rect 151 1040 181 1092
rect -99 237 13 267
rect -99 185 -69 237
rect -17 185 13 237
rect -99 -1471 13 185
rect 69 -618 181 1040
rect 237 680 313 690
rect 237 624 247 680
rect 303 624 313 680
rect 237 614 313 624
rect 564 234 620 1275
rect 700 715 756 1382
rect 1581 1092 1693 1122
rect 1581 1040 1611 1092
rect 1663 1040 1693 1092
rect 688 703 768 715
rect 688 647 700 703
rect 756 647 768 703
rect 688 635 768 647
rect 700 570 756 635
rect 682 558 762 570
rect 682 502 694 558
rect 750 502 762 558
rect 682 490 762 502
rect 552 222 632 234
rect 552 166 564 222
rect 620 166 632 222
rect 552 154 632 166
rect 564 -42 620 154
rect 552 -54 632 -42
rect 552 -110 564 -54
rect 620 -110 632 -54
rect 700 -74 756 490
rect 1082 225 1158 234
rect 1082 169 1092 225
rect 1148 169 1158 225
rect 1082 158 1158 169
rect 552 -122 632 -110
rect 690 -84 766 -74
rect 690 -140 700 -84
rect 756 -140 766 -84
rect 690 -150 766 -140
rect 237 -206 313 -196
rect 237 -262 247 -206
rect 303 -262 313 -206
rect 237 -272 313 -262
rect 700 -523 756 -150
rect 688 -535 768 -523
rect 688 -591 700 -535
rect 756 -591 768 -535
rect 688 -603 768 -591
rect 69 -670 99 -618
rect 151 -670 181 -618
rect 69 -700 181 -670
rect 235 -1026 315 -1014
rect 235 -1082 247 -1026
rect 303 -1082 315 -1026
rect 235 -1094 315 -1082
rect 427 -1151 507 -1139
rect 427 -1207 439 -1151
rect 495 -1207 507 -1151
rect 427 -1219 507 -1207
rect 700 -1305 756 -603
rect 1581 -928 1693 1040
rect 2282 810 2338 1489
rect 2395 1446 2471 1458
rect 2395 1394 2407 1446
rect 2459 1394 2471 1446
rect 2395 1382 2471 1394
rect 2272 798 2348 810
rect 2272 746 2284 798
rect 2336 746 2348 798
rect 2272 734 2348 746
rect 1581 -980 1611 -928
rect 1663 -980 1693 -928
rect 1581 -1010 1693 -980
rect 2003 82 2115 112
rect 2003 30 2033 82
rect 2085 30 2115 82
rect 688 -1317 768 -1305
rect 688 -1373 700 -1317
rect 756 -1373 768 -1317
rect 688 -1385 768 -1373
rect -99 -1523 -69 -1471
rect -17 -1523 13 -1471
rect -99 -1553 13 -1523
rect 1349 -1797 1425 -1787
rect 1349 -1853 1359 -1797
rect 1415 -1853 1425 -1797
rect 1349 -1863 1425 -1853
rect 2003 -1938 2115 30
rect 2405 -622 2461 1382
rect 2518 1339 2594 1351
rect 2518 1287 2530 1339
rect 2582 1287 2594 1339
rect 2518 1275 2594 1287
rect 2395 -634 2471 -622
rect 2395 -686 2407 -634
rect 2459 -686 2471 -634
rect 2395 -698 2471 -686
rect 2528 -1208 2584 1275
rect 2654 1232 2730 1244
rect 2654 1180 2666 1232
rect 2718 1180 2730 1232
rect 2654 1168 2730 1180
rect 2664 715 2720 1168
rect 2652 703 2733 715
rect 2652 647 2664 703
rect 2720 647 2733 703
rect 2652 635 2733 647
rect 5065 680 5121 690
rect 2664 263 2720 635
rect 2651 251 2732 263
rect 2651 195 2663 251
rect 2719 195 2732 251
rect 5065 249 5121 624
rect 2651 183 2732 195
rect 3732 223 3808 233
rect 2664 -1141 2720 183
rect 3732 167 3742 223
rect 3798 167 3808 223
rect 3732 157 3808 167
rect 5065 197 5067 249
rect 5119 197 5121 249
rect 2924 -58 2980 -46
rect 2780 -83 2860 -71
rect 2780 -139 2792 -83
rect 2848 -139 2860 -83
rect 2780 -151 2860 -139
rect 2924 -110 2926 -58
rect 2978 -110 2980 -58
rect 2792 -532 2848 -151
rect 2924 -196 2980 -110
rect 4757 -84 4833 -74
rect 4757 -140 4767 -84
rect 4823 -140 4833 -84
rect 4757 -150 4833 -140
rect 2914 -206 2990 -196
rect 2914 -262 2924 -206
rect 2980 -262 2990 -206
rect 2914 -272 2990 -262
rect 2792 -594 2794 -532
rect 2846 -594 2848 -532
rect 2792 -1016 2848 -594
rect 2782 -1026 2858 -1016
rect 2782 -1082 2792 -1026
rect 2848 -1082 2858 -1026
rect 2782 -1092 2858 -1082
rect 2654 -1151 2730 -1141
rect 2654 -1207 2664 -1151
rect 2720 -1207 2730 -1151
rect 2516 -1220 2596 -1208
rect 2654 -1217 2730 -1207
rect 2516 -1276 2528 -1220
rect 2584 -1276 2596 -1220
rect 2516 -1288 2596 -1276
rect 2664 -1757 2720 -1217
rect 2652 -1769 2732 -1757
rect 2652 -1825 2664 -1769
rect 2720 -1825 2732 -1769
rect 2652 -1837 2732 -1825
rect 2792 -1804 2848 -1092
rect 2924 -1478 2980 -272
rect 2915 -1490 2993 -1478
rect 2915 -1544 2927 -1490
rect 2979 -1544 2993 -1490
rect 2915 -1556 2993 -1544
rect 2924 -1787 2980 -1556
rect 2792 -1856 2794 -1804
rect 2846 -1856 2848 -1804
rect 2792 -1868 2848 -1856
rect 2914 -1797 2990 -1787
rect 2914 -1853 2924 -1797
rect 2980 -1853 2990 -1797
rect 2914 -1863 2990 -1853
rect 5065 -1794 5121 197
rect 5065 -1846 5067 -1794
rect 5119 -1846 5121 -1794
rect 5065 -1858 5121 -1846
rect 2003 -1990 2033 -1938
rect 2085 -1990 2115 -1938
rect 2003 -2020 2115 -1990
<< via2 >>
rect 247 678 303 680
rect 247 626 249 678
rect 249 626 301 678
rect 301 626 303 678
rect 247 624 303 626
rect 1092 222 1148 225
rect 1092 170 1094 222
rect 1094 170 1146 222
rect 1146 170 1148 222
rect 1092 169 1148 170
rect 700 -140 756 -84
rect 247 -208 303 -206
rect 247 -260 249 -208
rect 249 -260 301 -208
rect 301 -260 303 -208
rect 247 -262 303 -260
rect 247 -1082 303 -1026
rect 439 -1207 495 -1151
rect 1359 -1799 1415 -1797
rect 1359 -1851 1361 -1799
rect 1361 -1851 1413 -1799
rect 1413 -1851 1415 -1799
rect 1359 -1853 1415 -1851
rect 5065 624 5121 680
rect 3742 221 3798 223
rect 3742 169 3744 221
rect 3744 169 3796 221
rect 3796 169 3798 221
rect 3742 167 3798 169
rect 4767 -140 4823 -84
rect 2924 -262 2980 -206
rect 2792 -1082 2848 -1026
rect 2664 -1207 2720 -1151
rect 2924 -1853 2980 -1797
<< metal3 >>
rect 237 680 313 690
rect 5055 680 5131 690
rect 237 624 247 680
rect 303 624 5065 680
rect 5121 624 5131 680
rect 237 614 313 624
rect 5055 614 5131 624
rect 1082 225 1158 234
rect 1082 169 1092 225
rect 1148 223 1158 225
rect 2234 223 2389 224
rect 3732 223 3808 233
rect 1148 169 3742 223
rect 1082 167 3742 169
rect 3798 167 3808 223
rect 1082 158 1158 167
rect 3732 157 3808 167
rect 690 -84 766 -74
rect 4757 -84 4833 -74
rect 690 -140 700 -84
rect 756 -140 4767 -84
rect 4823 -140 4833 -84
rect 690 -150 766 -140
rect 4757 -150 4833 -140
rect 237 -206 313 -196
rect 2914 -206 2990 -196
rect 237 -262 247 -206
rect 303 -262 2924 -206
rect 2980 -262 2990 -206
rect 237 -272 313 -262
rect 2914 -272 2990 -262
rect 237 -1026 313 -1016
rect 2782 -1026 2858 -1016
rect 237 -1082 247 -1026
rect 303 -1082 2792 -1026
rect 2848 -1082 2858 -1026
rect 237 -1092 313 -1082
rect 2782 -1092 2858 -1082
rect 427 -1151 507 -1139
rect 2654 -1151 2730 -1141
rect 427 -1207 439 -1151
rect 495 -1207 2664 -1151
rect 2720 -1207 2730 -1151
rect 427 -1219 507 -1207
rect 2654 -1217 2730 -1207
rect 1349 -1797 1425 -1787
rect 2914 -1797 2990 -1781
rect 1349 -1853 1359 -1797
rect 1415 -1853 2924 -1797
rect 2980 -1853 2990 -1797
rect 1349 -1863 1425 -1853
rect 2914 -1863 2990 -1853
use AND_2_In_Layout  AND_2_In_Layout_0 ~/GF180Projects/Tapeout/Magic/Logic_Gates/AND_2_Input
timestamp 1695658812
transform 1 0 4124 0 1 -1718
box 0 -308 1085 833
use AND_3_In_Layout  AND_3_In_Layout_0 ~/GF180Projects/Tapeout/Magic/Logic_Gates/AND_3_Input
timestamp 1699521709
transform 1 0 777 0 1 -1713
box 0 -307 1783 828
use AND_3_In_Layout  AND_3_In_Layout_1
timestamp 1699521709
transform 1 0 3160 0 1 307
box 0 -307 1783 828
use AND_3_In_Layout  AND_3_In_Layout_2
timestamp 1699521709
transform 1 0 3160 0 -1 -195
box 0 -307 1783 828
use AND_3_In_Layout  AND_3_In_Layout_3
timestamp 1699521709
transform 1 0 777 0 1 307
box 0 -307 1783 828
use AND_3_In_Layout  AND_3_In_Layout_4
timestamp 1699521709
transform 1 0 777 0 -1 -195
box 0 -307 1783 828
use Inverter_Layout  Inverter_Layout_0 ~/GF180Projects/Tapeout/Magic/Logic_Gates/Inverter
timestamp 1699521709
transform -1 0 495 0 1 -1431
box -62 -124 342 856
use Inverter_Layout  Inverter_Layout_1
timestamp 1699521709
transform -1 0 495 0 1 279
box -62 -124 342 856
use Inverter_Layout  Inverter_Layout_2
timestamp 1699521709
transform -1 0 495 0 -1 143
box -62 -124 342 856
use OR_2_In_Layout  OR_2_In_Layout_0 ~/GF180Projects/Tapeout/Magic/Logic_Gates/OR_2_Input
timestamp 1695658812
transform 1 0 2913 0 1 -1786
box 0 -240 1172 901
<< labels >>
flabel metal1 400 1313 400 1313 0 FreeSans 320 0 0 0 B
port 1 nsew
flabel metal1 400 1206 400 1206 0 FreeSans 320 0 0 0 C
port 2 nsew
flabel metal1 400 1420 400 1420 0 FreeSans 320 0 0 0 A
port 0 nsew
flabel metal1 5339 -1253 5339 -1253 0 FreeSans 320 0 0 0 S1
port 4 nsew
flabel metal1 5339 -660 5339 -660 0 FreeSans 320 0 0 0 S3
port 5 nsew
flabel metal1 5339 772 5339 772 0 FreeSans 320 0 0 0 S2
port 6 nsew
flabel metal1 2776 1527 2776 1527 0 FreeSans 320 0 0 0 S6
port 7 nsew
flabel metal1 2776 1420 2776 1420 0 FreeSans 320 0 0 0 S5
port 8 nsew
flabel metal1 2776 1313 2776 1313 0 FreeSans 320 0 0 0 S4
port 9 nsew
flabel metal1 3209 1066 3209 1066 0 FreeSans 320 0 0 0 VDD
port 11 nsew
flabel metal1 3014 -1964 3014 -1964 0 FreeSans 320 0 0 0 VSS
port 12 nsew
<< end >>
