* NGSPICE file created from folded_single_check4_flat.ext - technology: gf180mcuC


* Top level circuit folded_single_check4_flat

C0 a_n2688_n4475# m1_n2767_n4043# 0.0515f
C1 a_n2688_n4475# m1_n2607_n3890# 0.0335f
C2 m3_n2833_n4475# a_n1553_n4448# 6.65e-20
C3 a_n3086_n4453# a_n2688_n4475# 0.0105f
C4 w_n3327_n4475# a_n2688_n4475# 0.581f
C5 m3_n2833_n4475# m1_n3088_n4204# 0.0409f
C6 m1_n2607_n3890# a_n1553_n4448# 1.16e-19
C7 m1_n2767_n4043# m1_n3088_n4204# 0.523f
C8 a_n3086_n4453# a_n1553_n4448# 0.00192f
C9 w_n3327_n4475# a_n1553_n4448# 0.197f
C10 m1_n2607_n3890# m1_n3088_n4204# 0.221f
C11 a_n3086_n4453# m1_n3088_n4204# 0.0312f
C12 w_n3327_n4475# m1_n3088_n4204# 0.431f
C13 m3_n2833_n4475# m1_n2767_n4043# 0.0518f
C14 m3_n2833_n4475# m1_n2607_n3890# 0.142f
C15 a_n3086_n4453# m3_n2833_n4475# 0.00338f
C16 w_n3327_n4475# m3_n2833_n4475# 0.0616f
C17 m1_n2607_n3890# m1_n2767_n4043# 0.311f
C18 a_n3086_n4453# m1_n2767_n4043# 0.00356f
C19 w_n3327_n4475# m1_n2767_n4043# 0.454f
C20 a_n2435_n4033# m1_n2767_n4043# 0.00293f
C21 a_n3086_n4453# m1_n2607_n3890# 3.17e-19
C22 w_n3327_n4475# m1_n2607_n3890# 0.19f
C23 w_n3327_n4475# a_n3086_n4453# 0.189f
C24 a_n2688_n4475# a_n1553_n4448# 0.028f
C25 a_n2688_n4475# m1_n3088_n4204# 0.268f
C26 a_n1553_n4448# m1_n3088_n4204# 0.0314f
C27 a_n2688_n4475# m3_n2833_n4475# 0.00415f
C28 m3_n2833_n4475# VSUBS 0.0951f $ **FLOATING
C29 m1_n3088_n4204# VSUBS 0.349f $ **FLOATING
C30 m1_n2767_n4043# VSUBS 0.425f $ **FLOATING
C31 m1_n2607_n3890# VSUBS 0.19f $ **FLOATING
C32 a_n1553_n4448# VSUBS 0.0546f $ **FLOATING
C33 a_n2688_n4475# VSUBS 0.47f $ **FLOATING
C34 a_n3086_n4453# VSUBS 0.0535f $ **FLOATING
C35 w_n3327_n4475# VSUBS 5.43f $ **FLOATING
.end

