magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2208 -2120 3080 2620
<< nwell >>
rect -208 -120 1080 620
<< mvpmos >>
rect 0 0 140 500
rect 244 0 384 500
rect 488 0 628 500
rect 732 0 872 500
<< mvpdiff >>
rect -88 487 0 500
rect -88 441 -75 487
rect -29 441 0 487
rect -88 380 0 441
rect -88 334 -75 380
rect -29 334 0 380
rect -88 273 0 334
rect -88 227 -75 273
rect -29 227 0 273
rect -88 166 0 227
rect -88 120 -75 166
rect -29 120 0 166
rect -88 59 0 120
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 140 487 244 500
rect 140 441 169 487
rect 215 441 244 487
rect 140 380 244 441
rect 140 334 169 380
rect 215 334 244 380
rect 140 273 244 334
rect 140 227 169 273
rect 215 227 244 273
rect 140 166 244 227
rect 140 120 169 166
rect 215 120 244 166
rect 140 59 244 120
rect 140 13 169 59
rect 215 13 244 59
rect 140 0 244 13
rect 384 487 488 500
rect 384 441 413 487
rect 459 441 488 487
rect 384 380 488 441
rect 384 334 413 380
rect 459 334 488 380
rect 384 273 488 334
rect 384 227 413 273
rect 459 227 488 273
rect 384 166 488 227
rect 384 120 413 166
rect 459 120 488 166
rect 384 59 488 120
rect 384 13 413 59
rect 459 13 488 59
rect 384 0 488 13
rect 628 487 732 500
rect 628 441 657 487
rect 703 441 732 487
rect 628 380 732 441
rect 628 334 657 380
rect 703 334 732 380
rect 628 273 732 334
rect 628 227 657 273
rect 703 227 732 273
rect 628 166 732 227
rect 628 120 657 166
rect 703 120 732 166
rect 628 59 732 120
rect 628 13 657 59
rect 703 13 732 59
rect 628 0 732 13
rect 872 487 960 500
rect 872 441 901 487
rect 947 441 960 487
rect 872 380 960 441
rect 872 334 901 380
rect 947 334 960 380
rect 872 273 960 334
rect 872 227 901 273
rect 947 227 960 273
rect 872 166 960 227
rect 872 120 901 166
rect 947 120 960 166
rect 872 59 960 120
rect 872 13 901 59
rect 947 13 960 59
rect 872 0 960 13
<< mvpdiffc >>
rect -75 441 -29 487
rect -75 334 -29 380
rect -75 227 -29 273
rect -75 120 -29 166
rect -75 13 -29 59
rect 169 441 215 487
rect 169 334 215 380
rect 169 227 215 273
rect 169 120 215 166
rect 169 13 215 59
rect 413 441 459 487
rect 413 334 459 380
rect 413 227 459 273
rect 413 120 459 166
rect 413 13 459 59
rect 657 441 703 487
rect 657 334 703 380
rect 657 227 703 273
rect 657 120 703 166
rect 657 13 703 59
rect 901 441 947 487
rect 901 334 947 380
rect 901 227 947 273
rect 901 120 947 166
rect 901 13 947 59
<< polysilicon >>
rect 0 500 140 544
rect 244 500 384 544
rect 488 500 628 544
rect 732 500 872 544
rect 0 -44 140 0
rect 244 -44 384 0
rect 488 -44 628 0
rect 732 -44 872 0
<< metal1 >>
rect -75 487 -29 500
rect -75 380 -29 441
rect -75 273 -29 334
rect -75 166 -29 227
rect -75 59 -29 120
rect -75 0 -29 13
rect 169 487 215 500
rect 169 380 215 441
rect 169 273 215 334
rect 169 166 215 227
rect 169 59 215 120
rect 169 0 215 13
rect 413 487 459 500
rect 413 380 459 441
rect 413 273 459 334
rect 413 166 459 227
rect 413 59 459 120
rect 413 0 459 13
rect 657 487 703 500
rect 657 380 703 441
rect 657 273 703 334
rect 657 166 703 227
rect 657 59 703 120
rect 657 0 703 13
rect 901 487 947 500
rect 901 380 947 441
rect 901 273 947 334
rect 901 166 947 227
rect 901 59 947 120
rect 901 0 947 13
<< labels >>
rlabel mvpdiffc 680 250 680 250 4 D
rlabel mvpdiffc 436 250 436 250 4 S
rlabel mvpdiffc 192 250 192 250 4 D
rlabel mvpdiffc 924 250 924 250 4 S
rlabel mvpdiffc -52 250 -52 250 4 S
<< end >>
