magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2145 -6145 2145 6145
<< psubdiff >>
rect -145 4112 145 4145
rect -145 -4112 -117 4112
rect 117 -4112 145 4112
rect -145 -4145 145 -4112
<< psubdiffcont >>
rect -117 -4112 117 4112
<< metal1 >>
rect -134 4112 134 4134
rect -134 -4112 -117 4112
rect 117 -4112 134 4112
rect -134 -4134 134 -4112
<< end >>
