magic
tech gf180mcuC
magscale 1 10
timestamp 1694400330
<< nwell >>
rect -4262 10 -4167 108
<< ndiff >>
rect 4608 -278 4641 -218
rect 4608 -528 4641 -468
<< psubdiff >>
rect 2665 1988 6316 1990
rect 2665 1986 6334 1988
rect 2665 1974 6353 1986
rect 2665 1920 2690 1974
rect 2763 1920 2834 1974
rect 2907 1920 2978 1974
rect 3051 1920 3122 1974
rect 3195 1920 3266 1974
rect 3339 1920 3410 1974
rect 3483 1920 3554 1974
rect 3627 1920 3698 1974
rect 3771 1920 3842 1974
rect 3915 1920 3986 1974
rect 4059 1920 4130 1974
rect 4203 1920 4274 1974
rect 4347 1920 4418 1974
rect 4491 1920 4562 1974
rect 4635 1920 4706 1974
rect 4779 1920 4850 1974
rect 4923 1920 4994 1974
rect 5067 1920 5138 1974
rect 5211 1920 5282 1974
rect 5355 1920 5426 1974
rect 5499 1920 5570 1974
rect 5643 1920 5714 1974
rect 5787 1920 5858 1974
rect 5931 1920 6002 1974
rect 6075 1920 6146 1974
rect 6219 1920 6353 1974
rect 2665 1892 6353 1920
rect 2665 1826 2764 1892
rect 2665 1772 2678 1826
rect 2751 1772 2764 1826
rect 6231 1854 6353 1892
rect 6231 1800 6254 1854
rect 6327 1800 6353 1854
rect 2665 1706 2764 1772
rect 2665 1652 2678 1706
rect 2751 1652 2764 1706
rect 2665 1586 2764 1652
rect 2665 1532 2678 1586
rect 2751 1532 2764 1586
rect 6231 1734 6353 1800
rect 6231 1680 6254 1734
rect 6327 1680 6353 1734
rect 6231 1614 6353 1680
rect 6231 1560 6254 1614
rect 6327 1560 6353 1614
rect 2665 1466 2764 1532
rect 2665 1412 2678 1466
rect 2751 1412 2764 1466
rect 2665 1346 2764 1412
rect 2665 1292 2678 1346
rect 2751 1292 2764 1346
rect 6231 1494 6353 1560
rect 6231 1440 6254 1494
rect 6327 1440 6353 1494
rect 6231 1374 6353 1440
rect 6231 1320 6254 1374
rect 6327 1320 6353 1374
rect 2665 1226 2764 1292
rect 2665 1172 2678 1226
rect 2751 1172 2764 1226
rect 6231 1254 6353 1320
rect 6231 1200 6254 1254
rect 6327 1200 6353 1254
rect 2665 1106 2764 1172
rect 2665 1052 2678 1106
rect 2751 1052 2764 1106
rect 2665 986 2764 1052
rect 2665 932 2678 986
rect 2751 932 2764 986
rect 6231 1134 6353 1200
rect 6231 1080 6254 1134
rect 6327 1080 6353 1134
rect 6231 1014 6353 1080
rect 6231 960 6254 1014
rect 6327 960 6353 1014
rect 2665 866 2764 932
rect 6231 894 6353 960
rect 2665 812 2678 866
rect 2751 812 2764 866
rect 2665 746 2764 812
rect 2665 692 2678 746
rect 2751 692 2764 746
rect 6231 840 6254 894
rect 6327 840 6353 894
rect 6231 774 6353 840
rect 6231 720 6254 774
rect 6327 720 6353 774
rect 2665 626 2764 692
rect 2665 572 2678 626
rect 2751 572 2764 626
rect 6231 654 6353 720
rect 2665 506 2764 572
rect 6231 600 6254 654
rect 6327 600 6353 654
rect 2665 452 2678 506
rect 2751 452 2764 506
rect 2665 386 2764 452
rect 6231 534 6353 600
rect 2665 332 2678 386
rect 2751 332 2764 386
rect 6231 480 6254 534
rect 6327 480 6353 534
rect 6231 414 6353 480
rect 2665 266 2764 332
rect 2665 212 2678 266
rect 2751 212 2764 266
rect 2665 146 2764 212
rect 6231 360 6254 414
rect 6327 360 6353 414
rect 2665 92 2678 146
rect 2751 92 2764 146
rect 6231 294 6353 360
rect 6231 240 6254 294
rect 6327 240 6353 294
rect 6231 174 6353 240
rect 6231 120 6254 174
rect 6327 120 6353 174
rect 2665 26 2764 92
rect 6231 54 6353 120
rect 2665 -28 2678 26
rect 2751 -28 2764 26
rect 2665 -94 2764 -28
rect 2665 -148 2678 -94
rect 2751 -148 2764 -94
rect 2665 -214 2764 -148
rect 6231 0 6254 54
rect 6327 0 6353 54
rect 6231 -66 6353 0
rect 2665 -268 2678 -214
rect 2751 -268 2764 -214
rect 6231 -120 6254 -66
rect 6327 -120 6353 -66
rect 6231 -186 6353 -120
rect 2665 -334 2764 -268
rect 6231 -240 6254 -186
rect 6327 -240 6353 -186
rect 6231 -306 6353 -240
rect 2665 -388 2678 -334
rect 2751 -388 2764 -334
rect 2665 -454 2764 -388
rect 2665 -508 2678 -454
rect 2751 -508 2764 -454
rect 6231 -360 6254 -306
rect 6327 -360 6353 -306
rect 6231 -426 6353 -360
rect 2665 -574 2764 -508
rect 6231 -480 6254 -426
rect 6327 -480 6353 -426
rect 6231 -546 6353 -480
rect 2665 -628 2678 -574
rect 2751 -628 2764 -574
rect 2665 -694 2764 -628
rect 2665 -748 2678 -694
rect 2751 -748 2764 -694
rect 2665 -814 2764 -748
rect 6231 -600 6254 -546
rect 6327 -600 6353 -546
rect 6231 -666 6353 -600
rect 6231 -720 6254 -666
rect 6327 -720 6353 -666
rect 6231 -786 6353 -720
rect 2665 -868 2678 -814
rect 2751 -868 2764 -814
rect 6231 -840 6254 -786
rect 6327 -840 6353 -786
rect 2665 -934 2764 -868
rect 2665 -988 2678 -934
rect 2751 -988 2764 -934
rect 2665 -1054 2764 -988
rect 2665 -1108 2678 -1054
rect 2751 -1108 2764 -1054
rect 2665 -1174 2764 -1108
rect 2665 -1228 2678 -1174
rect 2751 -1228 2764 -1174
rect 6231 -906 6353 -840
rect 6231 -960 6254 -906
rect 6327 -960 6353 -906
rect 6231 -1026 6353 -960
rect 6231 -1080 6254 -1026
rect 6327 -1080 6353 -1026
rect 2665 -1294 2764 -1228
rect 2665 -1348 2678 -1294
rect 2751 -1348 2764 -1294
rect 2665 -1414 2764 -1348
rect 2665 -1468 2678 -1414
rect 2751 -1468 2764 -1414
rect 6231 -1146 6353 -1080
rect 6231 -1200 6254 -1146
rect 6327 -1200 6353 -1146
rect 6231 -1266 6353 -1200
rect 6231 -1320 6254 -1266
rect 6327 -1320 6353 -1266
rect 6231 -1386 6353 -1320
rect 2665 -1550 2764 -1468
rect 6231 -1440 6254 -1386
rect 6327 -1440 6353 -1386
rect 3241 -1549 3435 -1548
rect 6231 -1549 6353 -1440
rect 3241 -1550 6452 -1549
rect 2665 -1564 6452 -1550
rect 2665 -1578 2681 -1564
rect 2667 -1618 2681 -1578
rect 2754 -1618 2806 -1564
rect 2879 -1618 2931 -1564
rect 3004 -1618 3056 -1564
rect 3129 -1618 3181 -1564
rect 3254 -1565 6452 -1564
rect 3254 -1614 3318 -1565
rect 3381 -1566 6229 -1565
rect 3381 -1614 3439 -1566
rect 3254 -1615 3439 -1614
rect 3502 -1615 3560 -1566
rect 3623 -1615 3681 -1566
rect 3744 -1615 3802 -1566
rect 3865 -1615 3923 -1566
rect 3986 -1615 4044 -1566
rect 4107 -1615 4165 -1566
rect 4228 -1615 4286 -1566
rect 4349 -1615 4407 -1566
rect 4470 -1615 4528 -1566
rect 4591 -1615 4649 -1566
rect 4712 -1615 4770 -1566
rect 4833 -1615 4891 -1566
rect 4954 -1615 5012 -1566
rect 5075 -1615 5133 -1566
rect 5196 -1615 5254 -1566
rect 5317 -1615 5375 -1566
rect 5438 -1615 5496 -1566
rect 5559 -1615 5617 -1566
rect 5680 -1615 5738 -1566
rect 5801 -1615 5859 -1566
rect 5922 -1615 5980 -1566
rect 6043 -1615 6101 -1566
rect 6164 -1614 6229 -1566
rect 6292 -1584 6452 -1565
rect 6292 -1614 6375 -1584
rect 6164 -1615 6375 -1614
rect 3254 -1618 6375 -1615
rect 2667 -1629 6375 -1618
rect 2667 -1635 3333 -1629
rect 3240 -1760 3333 -1635
rect 6360 -1633 6375 -1629
rect 6438 -1633 6452 -1584
rect 3240 -1809 3255 -1760
rect 3318 -1809 3333 -1760
rect 6360 -1691 6452 -1633
rect 6360 -1719 6375 -1691
rect 3240 -1871 3333 -1809
rect 6359 -1740 6375 -1719
rect 6438 -1740 6452 -1691
rect 3240 -1920 3255 -1871
rect 3318 -1920 3333 -1871
rect 6359 -1791 6452 -1740
rect 6359 -1840 6374 -1791
rect 6437 -1840 6452 -1791
rect 3240 -1982 3333 -1920
rect 3240 -2031 3255 -1982
rect 3318 -2031 3333 -1982
rect 3240 -2093 3333 -2031
rect 6359 -1902 6452 -1840
rect 6359 -1951 6374 -1902
rect 6437 -1951 6452 -1902
rect 6359 -2013 6452 -1951
rect 6359 -2062 6374 -2013
rect 6437 -2062 6452 -2013
rect 3240 -2142 3255 -2093
rect 3318 -2142 3333 -2093
rect 3240 -2204 3333 -2142
rect 3240 -2253 3255 -2204
rect 3318 -2253 3333 -2204
rect 6359 -2124 6452 -2062
rect 6359 -2173 6374 -2124
rect 6437 -2173 6452 -2124
rect 6359 -2235 6452 -2173
rect 3240 -2315 3333 -2253
rect 3240 -2364 3255 -2315
rect 3318 -2364 3333 -2315
rect 3240 -2426 3333 -2364
rect 3240 -2475 3255 -2426
rect 3318 -2475 3333 -2426
rect 6359 -2284 6374 -2235
rect 6437 -2284 6452 -2235
rect 6359 -2346 6452 -2284
rect 6359 -2395 6374 -2346
rect 6437 -2395 6452 -2346
rect -274 -2548 2823 -2535
rect -274 -2549 502 -2548
rect -274 -2598 -236 -2549
rect -173 -2550 21 -2549
rect -173 -2598 -108 -2550
rect -274 -2599 -108 -2598
rect -45 -2598 21 -2550
rect 84 -2550 373 -2549
rect 84 -2598 138 -2550
rect -45 -2599 138 -2598
rect 201 -2551 373 -2550
rect 201 -2599 250 -2551
rect -274 -2600 250 -2599
rect 313 -2598 373 -2551
rect 436 -2597 502 -2549
rect 565 -2549 1104 -2548
rect 565 -2597 619 -2549
rect 436 -2598 619 -2597
rect 682 -2550 975 -2549
rect 682 -2598 731 -2550
rect 313 -2599 731 -2598
rect 794 -2599 849 -2550
rect 912 -2598 975 -2550
rect 1038 -2597 1104 -2549
rect 1167 -2549 2823 -2548
rect 1167 -2597 1221 -2549
rect 1038 -2598 1221 -2597
rect 1284 -2550 2823 -2549
rect 1284 -2598 1333 -2550
rect 912 -2599 1333 -2598
rect 1396 -2599 1451 -2550
rect 1514 -2599 1574 -2550
rect 1637 -2599 1691 -2550
rect 1754 -2599 1812 -2550
rect 1875 -2599 1934 -2550
rect 1997 -2551 2516 -2550
rect 1997 -2599 2045 -2551
rect 313 -2600 2045 -2599
rect 2108 -2600 2164 -2551
rect 2227 -2600 2276 -2551
rect 2339 -2600 2397 -2551
rect 2460 -2599 2516 -2551
rect 2579 -2552 2742 -2550
rect 2579 -2599 2631 -2552
rect 2460 -2600 2631 -2599
rect -274 -2601 2631 -2600
rect 2694 -2599 2742 -2552
rect 2805 -2599 2823 -2550
rect 2694 -2601 2823 -2599
rect -274 -2615 2823 -2601
rect -274 -2664 -180 -2615
rect -274 -2711 -250 -2664
rect -196 -2711 -180 -2664
rect 2737 -2650 2823 -2615
rect -274 -2765 -180 -2711
rect -274 -2812 -249 -2765
rect -195 -2812 -180 -2765
rect -274 -2862 -180 -2812
rect -274 -2909 -250 -2862
rect -196 -2909 -180 -2862
rect -274 -2970 -180 -2909
rect -274 -3017 -249 -2970
rect -195 -3017 -180 -2970
rect -274 -3095 -180 -3017
rect -274 -3142 -249 -3095
rect -195 -3142 -180 -3095
rect -274 -3209 -180 -3142
rect 2737 -2697 2753 -2650
rect 2807 -2697 2823 -2650
rect 2737 -2751 2823 -2697
rect 2737 -2798 2754 -2751
rect 2808 -2798 2823 -2751
rect 2737 -2848 2823 -2798
rect 2737 -2895 2753 -2848
rect 2807 -2895 2823 -2848
rect 2737 -2956 2823 -2895
rect 2737 -3003 2754 -2956
rect 2808 -3003 2823 -2956
rect 2737 -3081 2823 -3003
rect 2737 -3128 2754 -3081
rect 2808 -3128 2823 -3081
rect -274 -3256 -248 -3209
rect -194 -3256 -180 -3209
rect -274 -3321 -180 -3256
rect 2737 -3195 2823 -3128
rect 2737 -3242 2755 -3195
rect 2809 -3242 2823 -3195
rect -274 -3368 -247 -3321
rect -193 -3368 -180 -3321
rect -274 -3425 -180 -3368
rect -274 -3472 -249 -3425
rect -195 -3472 -180 -3425
rect -274 -3529 -180 -3472
rect -274 -3576 -249 -3529
rect -195 -3576 -180 -3529
rect 2737 -3307 2823 -3242
rect 2737 -3354 2756 -3307
rect 2810 -3354 2823 -3307
rect 2737 -3411 2823 -3354
rect 2737 -3458 2754 -3411
rect 2808 -3458 2823 -3411
rect 2737 -3515 2823 -3458
rect -274 -3624 -180 -3576
rect -274 -3671 -251 -3624
rect -197 -3671 -180 -3624
rect -274 -3733 -180 -3671
rect 2737 -3562 2754 -3515
rect 2808 -3562 2823 -3515
rect 2737 -3610 2823 -3562
rect 2737 -3657 2752 -3610
rect 2806 -3657 2823 -3610
rect -274 -3780 -250 -3733
rect -196 -3780 -180 -3733
rect -274 -3837 -180 -3780
rect -274 -3884 -250 -3837
rect -196 -3884 -180 -3837
rect 2737 -3719 2823 -3657
rect 2737 -3766 2753 -3719
rect 2807 -3766 2823 -3719
rect 2737 -3823 2823 -3766
rect -274 -3932 -180 -3884
rect -274 -3979 -252 -3932
rect -198 -3979 -180 -3932
rect -274 -4042 -180 -3979
rect -274 -4089 -251 -4042
rect -197 -4089 -180 -4042
rect 2737 -3870 2753 -3823
rect 2807 -3870 2823 -3823
rect 2737 -3918 2823 -3870
rect 2737 -3965 2751 -3918
rect 2805 -3965 2823 -3918
rect 2737 -4028 2823 -3965
rect -274 -4146 -180 -4089
rect -274 -4193 -251 -4146
rect -197 -4193 -180 -4146
rect -274 -4241 -180 -4193
rect -274 -4288 -253 -4241
rect -199 -4288 -180 -4241
rect 2737 -4075 2752 -4028
rect 2806 -4075 2823 -4028
rect 2737 -4132 2823 -4075
rect 2737 -4179 2752 -4132
rect 2806 -4179 2823 -4132
rect 2737 -4227 2823 -4179
rect -274 -4342 -180 -4288
rect -274 -4389 -250 -4342
rect -196 -4389 -180 -4342
rect 2737 -4274 2750 -4227
rect 2804 -4274 2823 -4227
rect 2737 -4328 2823 -4274
rect -274 -4446 -180 -4389
rect -274 -4493 -250 -4446
rect -196 -4493 -180 -4446
rect -274 -4541 -180 -4493
rect -274 -4588 -252 -4541
rect -198 -4588 -180 -4541
rect 2737 -4375 2753 -4328
rect 2807 -4375 2823 -4328
rect 2737 -4432 2823 -4375
rect 2737 -4479 2753 -4432
rect 2807 -4479 2823 -4432
rect 2737 -4527 2823 -4479
rect -274 -4651 -180 -4588
rect 2737 -4574 2751 -4527
rect 2805 -4574 2823 -4527
rect -274 -4698 -251 -4651
rect -197 -4698 -180 -4651
rect -274 -4755 -180 -4698
rect 2737 -4637 2823 -4574
rect 2737 -4684 2752 -4637
rect 2806 -4684 2823 -4637
rect -274 -4802 -251 -4755
rect -197 -4802 -180 -4755
rect -274 -4850 -180 -4802
rect -274 -4897 -253 -4850
rect -199 -4897 -180 -4850
rect -274 -4954 -180 -4897
rect 2737 -4741 2823 -4684
rect 2737 -4788 2752 -4741
rect 2806 -4788 2823 -4741
rect 2737 -4836 2823 -4788
rect 2737 -4883 2750 -4836
rect 2804 -4883 2823 -4836
rect -274 -5001 -249 -4954
rect -195 -5001 -180 -4954
rect -274 -5064 -180 -5001
rect -274 -5111 -248 -5064
rect -194 -5111 -180 -5064
rect 2737 -4940 2823 -4883
rect 2737 -4987 2754 -4940
rect 2808 -4987 2823 -4940
rect 2737 -5050 2823 -4987
rect -274 -5168 -180 -5111
rect -274 -5215 -248 -5168
rect -194 -5215 -180 -5168
rect -274 -5272 -180 -5215
rect 2737 -5097 2755 -5050
rect 2809 -5097 2823 -5050
rect 2737 -5154 2823 -5097
rect 2737 -5201 2755 -5154
rect 2809 -5201 2823 -5154
rect 2737 -5272 2823 -5201
rect -274 -5285 2823 -5272
rect -274 -5286 499 -5285
rect -274 -5335 -239 -5286
rect -176 -5287 18 -5286
rect -176 -5335 -111 -5287
rect -274 -5336 -111 -5335
rect -48 -5335 18 -5287
rect 81 -5287 370 -5286
rect 81 -5335 135 -5287
rect -48 -5336 135 -5335
rect 198 -5288 370 -5287
rect 198 -5336 247 -5288
rect -274 -5337 247 -5336
rect 310 -5335 370 -5288
rect 433 -5334 499 -5286
rect 562 -5286 1101 -5285
rect 562 -5334 616 -5286
rect 433 -5335 616 -5334
rect 679 -5287 972 -5286
rect 679 -5335 728 -5287
rect 310 -5336 728 -5335
rect 791 -5336 846 -5287
rect 909 -5335 972 -5287
rect 1035 -5334 1101 -5286
rect 1164 -5286 2823 -5285
rect 1164 -5334 1218 -5286
rect 1035 -5335 1218 -5334
rect 1281 -5287 2823 -5286
rect 1281 -5335 1330 -5287
rect 909 -5336 1330 -5335
rect 1393 -5336 1448 -5287
rect 1511 -5336 1571 -5287
rect 1634 -5336 1688 -5287
rect 1751 -5336 1809 -5287
rect 1872 -5336 1931 -5287
rect 1994 -5288 2513 -5287
rect 1994 -5336 2042 -5288
rect 310 -5337 2042 -5336
rect 2105 -5337 2161 -5288
rect 2224 -5337 2273 -5288
rect 2336 -5337 2394 -5288
rect 2457 -5336 2513 -5288
rect 2576 -5289 2739 -5287
rect 2576 -5336 2628 -5289
rect 2457 -5337 2628 -5336
rect -274 -5338 2628 -5337
rect 2691 -5336 2739 -5289
rect 2802 -5336 2823 -5287
rect 2691 -5338 2823 -5336
rect -274 -5352 2823 -5338
rect 3240 -2537 3333 -2475
rect 6359 -2457 6452 -2395
rect 6359 -2506 6374 -2457
rect 6437 -2506 6452 -2457
rect 3240 -2586 3255 -2537
rect 3318 -2586 3333 -2537
rect 3240 -2648 3333 -2586
rect 3240 -2697 3255 -2648
rect 3318 -2697 3333 -2648
rect 3240 -2759 3333 -2697
rect 6359 -2568 6452 -2506
rect 6359 -2617 6374 -2568
rect 6437 -2617 6452 -2568
rect 6359 -2679 6452 -2617
rect 6359 -2728 6374 -2679
rect 6437 -2728 6452 -2679
rect 3240 -2808 3255 -2759
rect 3318 -2808 3333 -2759
rect 3240 -2870 3333 -2808
rect 3240 -2919 3255 -2870
rect 3318 -2919 3333 -2870
rect 6359 -2790 6452 -2728
rect 3240 -2981 3333 -2919
rect 6359 -2839 6374 -2790
rect 6437 -2839 6452 -2790
rect 6359 -2901 6452 -2839
rect 3240 -3030 3255 -2981
rect 3318 -3030 3333 -2981
rect 3240 -3092 3333 -3030
rect 3240 -3141 3255 -3092
rect 3318 -3141 3333 -3092
rect 6359 -2950 6374 -2901
rect 6437 -2950 6452 -2901
rect 6359 -3012 6452 -2950
rect 6359 -3061 6374 -3012
rect 6437 -3061 6452 -3012
rect 3240 -3203 3333 -3141
rect 3240 -3252 3255 -3203
rect 3318 -3252 3333 -3203
rect 6359 -3123 6452 -3061
rect 3240 -3314 3333 -3252
rect 6359 -3172 6374 -3123
rect 6437 -3172 6452 -3123
rect 6359 -3234 6452 -3172
rect 3240 -3363 3255 -3314
rect 3318 -3363 3333 -3314
rect 3240 -3425 3333 -3363
rect 6359 -3283 6374 -3234
rect 6437 -3283 6452 -3234
rect 6359 -3345 6452 -3283
rect 6359 -3394 6374 -3345
rect 6437 -3394 6452 -3345
rect 3240 -3474 3255 -3425
rect 3318 -3474 3333 -3425
rect 3240 -3536 3333 -3474
rect 6359 -3456 6452 -3394
rect 3240 -3585 3255 -3536
rect 3318 -3585 3333 -3536
rect 6359 -3505 6374 -3456
rect 6437 -3505 6452 -3456
rect 3240 -3647 3333 -3585
rect 3240 -3696 3255 -3647
rect 3318 -3696 3333 -3647
rect 3240 -3758 3333 -3696
rect 6359 -3567 6452 -3505
rect 6359 -3616 6374 -3567
rect 6437 -3616 6452 -3567
rect 6359 -3678 6452 -3616
rect 6359 -3727 6374 -3678
rect 6437 -3727 6452 -3678
rect 3240 -3807 3255 -3758
rect 3318 -3807 3333 -3758
rect 3240 -3869 3333 -3807
rect 6359 -3789 6452 -3727
rect 3240 -3918 3255 -3869
rect 3318 -3918 3333 -3869
rect 3240 -3980 3333 -3918
rect 3240 -4029 3255 -3980
rect 3318 -4029 3333 -3980
rect 3240 -4091 3333 -4029
rect 3240 -4140 3255 -4091
rect 3318 -4140 3333 -4091
rect 3240 -4202 3333 -4140
rect 6359 -3838 6374 -3789
rect 6437 -3838 6452 -3789
rect 6359 -3900 6452 -3838
rect 6359 -3949 6374 -3900
rect 6437 -3949 6452 -3900
rect 6359 -4011 6452 -3949
rect 6359 -4060 6374 -4011
rect 6437 -4060 6452 -4011
rect 6359 -4122 6452 -4060
rect 3240 -4251 3255 -4202
rect 3318 -4251 3333 -4202
rect 3240 -4313 3333 -4251
rect 6359 -4171 6374 -4122
rect 6437 -4171 6452 -4122
rect 6359 -4233 6452 -4171
rect 3240 -4362 3255 -4313
rect 3318 -4362 3333 -4313
rect 3240 -4424 3333 -4362
rect 3240 -4473 3255 -4424
rect 3318 -4473 3333 -4424
rect 6359 -4282 6374 -4233
rect 6437 -4282 6452 -4233
rect 6359 -4344 6452 -4282
rect 6359 -4393 6374 -4344
rect 6437 -4393 6452 -4344
rect 3240 -4535 3333 -4473
rect 3240 -4584 3255 -4535
rect 3318 -4584 3333 -4535
rect 6359 -4455 6452 -4393
rect 3240 -4646 3333 -4584
rect 3240 -4695 3255 -4646
rect 3318 -4695 3333 -4646
rect 3240 -4757 3333 -4695
rect 3240 -4806 3255 -4757
rect 3318 -4806 3333 -4757
rect 3240 -4868 3333 -4806
rect 3240 -4917 3255 -4868
rect 3318 -4917 3333 -4868
rect 3240 -4979 3333 -4917
rect 3240 -5028 3255 -4979
rect 3318 -5028 3333 -4979
rect 3240 -5090 3333 -5028
rect 3240 -5139 3255 -5090
rect 3318 -5139 3333 -5090
rect 3240 -5201 3333 -5139
rect 3240 -5250 3255 -5201
rect 3318 -5250 3333 -5201
rect 6359 -4504 6374 -4455
rect 6437 -4504 6452 -4455
rect 6359 -4566 6452 -4504
rect 6359 -4615 6374 -4566
rect 6437 -4615 6452 -4566
rect 6359 -4677 6452 -4615
rect 6359 -4726 6374 -4677
rect 6437 -4726 6452 -4677
rect 6359 -4788 6452 -4726
rect 6359 -4837 6374 -4788
rect 6437 -4837 6452 -4788
rect 6359 -4899 6452 -4837
rect 6359 -4948 6374 -4899
rect 6437 -4948 6452 -4899
rect 6359 -5010 6452 -4948
rect 6359 -5059 6374 -5010
rect 6437 -5059 6452 -5010
rect 6359 -5121 6452 -5059
rect 6359 -5170 6374 -5121
rect 6437 -5170 6452 -5121
rect 3240 -5312 3333 -5250
rect 3240 -5361 3255 -5312
rect 3318 -5361 3333 -5312
rect 3240 -5423 3333 -5361
rect 3240 -5472 3255 -5423
rect 3318 -5472 3333 -5423
rect 3240 -5534 3333 -5472
rect 3240 -5583 3255 -5534
rect 3318 -5583 3333 -5534
rect 3240 -5645 3333 -5583
rect 3240 -5694 3255 -5645
rect 3318 -5694 3333 -5645
rect 3240 -5756 3333 -5694
rect 3240 -5805 3255 -5756
rect 3318 -5805 3333 -5756
rect 3240 -5867 3333 -5805
rect 6359 -5232 6452 -5170
rect 6359 -5281 6374 -5232
rect 6437 -5281 6452 -5232
rect 6359 -5343 6452 -5281
rect 6359 -5392 6374 -5343
rect 6437 -5392 6452 -5343
rect 6359 -5454 6452 -5392
rect 6359 -5503 6374 -5454
rect 6437 -5503 6452 -5454
rect 6359 -5565 6452 -5503
rect 6359 -5614 6374 -5565
rect 6437 -5614 6452 -5565
rect 6359 -5676 6452 -5614
rect 6359 -5725 6374 -5676
rect 6437 -5725 6452 -5676
rect 6359 -5787 6452 -5725
rect 6359 -5836 6374 -5787
rect 6437 -5836 6452 -5787
rect 3240 -5916 3255 -5867
rect 3318 -5916 3333 -5867
rect 3240 -5978 3333 -5916
rect 6359 -5898 6452 -5836
rect 3240 -6027 3255 -5978
rect 3318 -6027 3333 -5978
rect 6359 -5947 6374 -5898
rect 6437 -5947 6452 -5898
rect 6359 -6009 6452 -5947
rect 3240 -6089 3333 -6027
rect 3240 -6138 3255 -6089
rect 3318 -6138 3333 -6089
rect 3240 -6200 3333 -6138
rect 3240 -6249 3255 -6200
rect 3318 -6249 3333 -6200
rect 6359 -6058 6374 -6009
rect 6437 -6058 6452 -6009
rect 6359 -6120 6452 -6058
rect 6359 -6169 6374 -6120
rect 6437 -6169 6452 -6120
rect 3240 -6311 3333 -6249
rect 3240 -6360 3255 -6311
rect 3318 -6360 3333 -6311
rect 6359 -6231 6452 -6169
rect 3240 -6422 3333 -6360
rect 6359 -6280 6374 -6231
rect 6437 -6280 6452 -6231
rect 6359 -6342 6452 -6280
rect 3240 -6471 3255 -6422
rect 3318 -6471 3333 -6422
rect 3240 -6594 3333 -6471
rect 6359 -6391 6374 -6342
rect 6437 -6391 6452 -6342
rect 6359 -6453 6452 -6391
rect 6359 -6502 6374 -6453
rect 6437 -6502 6452 -6453
rect 3240 -6595 3435 -6594
rect 6359 -6595 6452 -6502
rect 3240 -6611 6452 -6595
rect 3240 -6660 3318 -6611
rect 3381 -6612 6452 -6611
rect 3381 -6660 3439 -6612
rect 3240 -6661 3439 -6660
rect 3502 -6661 3560 -6612
rect 3623 -6661 3681 -6612
rect 3744 -6661 3802 -6612
rect 3865 -6661 3923 -6612
rect 3986 -6661 4044 -6612
rect 4107 -6661 4165 -6612
rect 4228 -6661 4286 -6612
rect 4349 -6661 4407 -6612
rect 4470 -6661 4528 -6612
rect 4591 -6661 4649 -6612
rect 4712 -6661 4770 -6612
rect 4833 -6661 4891 -6612
rect 4954 -6661 5012 -6612
rect 5075 -6661 5133 -6612
rect 5196 -6661 5254 -6612
rect 5317 -6661 5375 -6612
rect 5438 -6661 5496 -6612
rect 5559 -6661 5617 -6612
rect 5680 -6661 5738 -6612
rect 5801 -6661 5859 -6612
rect 5922 -6661 5980 -6612
rect 6043 -6661 6101 -6612
rect 6164 -6661 6452 -6612
rect 3240 -6675 6452 -6661
rect 3240 -6677 3333 -6675
<< psubdiffcont >>
rect 2690 1920 2763 1974
rect 2834 1920 2907 1974
rect 2978 1920 3051 1974
rect 3122 1920 3195 1974
rect 3266 1920 3339 1974
rect 3410 1920 3483 1974
rect 3554 1920 3627 1974
rect 3698 1920 3771 1974
rect 3842 1920 3915 1974
rect 3986 1920 4059 1974
rect 4130 1920 4203 1974
rect 4274 1920 4347 1974
rect 4418 1920 4491 1974
rect 4562 1920 4635 1974
rect 4706 1920 4779 1974
rect 4850 1920 4923 1974
rect 4994 1920 5067 1974
rect 5138 1920 5211 1974
rect 5282 1920 5355 1974
rect 5426 1920 5499 1974
rect 5570 1920 5643 1974
rect 5714 1920 5787 1974
rect 5858 1920 5931 1974
rect 6002 1920 6075 1974
rect 6146 1920 6219 1974
rect 2678 1772 2751 1826
rect 6254 1800 6327 1854
rect 2678 1652 2751 1706
rect 2678 1532 2751 1586
rect 6254 1680 6327 1734
rect 6254 1560 6327 1614
rect 2678 1412 2751 1466
rect 2678 1292 2751 1346
rect 6254 1440 6327 1494
rect 6254 1320 6327 1374
rect 2678 1172 2751 1226
rect 6254 1200 6327 1254
rect 2678 1052 2751 1106
rect 2678 932 2751 986
rect 6254 1080 6327 1134
rect 6254 960 6327 1014
rect 2678 812 2751 866
rect 2678 692 2751 746
rect 6254 840 6327 894
rect 6254 720 6327 774
rect 2678 572 2751 626
rect 6254 600 6327 654
rect 2678 452 2751 506
rect 2678 332 2751 386
rect 6254 480 6327 534
rect 2678 212 2751 266
rect 6254 360 6327 414
rect 2678 92 2751 146
rect 6254 240 6327 294
rect 6254 120 6327 174
rect 2678 -28 2751 26
rect 2678 -148 2751 -94
rect 6254 0 6327 54
rect 2678 -268 2751 -214
rect 6254 -120 6327 -66
rect 6254 -240 6327 -186
rect 2678 -388 2751 -334
rect 2678 -508 2751 -454
rect 6254 -360 6327 -306
rect 6254 -480 6327 -426
rect 2678 -628 2751 -574
rect 2678 -748 2751 -694
rect 6254 -600 6327 -546
rect 6254 -720 6327 -666
rect 2678 -868 2751 -814
rect 6254 -840 6327 -786
rect 2678 -988 2751 -934
rect 2678 -1108 2751 -1054
rect 2678 -1228 2751 -1174
rect 6254 -960 6327 -906
rect 6254 -1080 6327 -1026
rect 2678 -1348 2751 -1294
rect 2678 -1468 2751 -1414
rect 6254 -1200 6327 -1146
rect 6254 -1320 6327 -1266
rect 6254 -1440 6327 -1386
rect 2681 -1618 2754 -1564
rect 2806 -1618 2879 -1564
rect 2931 -1618 3004 -1564
rect 3056 -1618 3129 -1564
rect 3181 -1618 3254 -1564
rect 3318 -1614 3381 -1565
rect 3439 -1615 3502 -1566
rect 3560 -1615 3623 -1566
rect 3681 -1615 3744 -1566
rect 3802 -1615 3865 -1566
rect 3923 -1615 3986 -1566
rect 4044 -1615 4107 -1566
rect 4165 -1615 4228 -1566
rect 4286 -1615 4349 -1566
rect 4407 -1615 4470 -1566
rect 4528 -1615 4591 -1566
rect 4649 -1615 4712 -1566
rect 4770 -1615 4833 -1566
rect 4891 -1615 4954 -1566
rect 5012 -1615 5075 -1566
rect 5133 -1615 5196 -1566
rect 5254 -1615 5317 -1566
rect 5375 -1615 5438 -1566
rect 5496 -1615 5559 -1566
rect 5617 -1615 5680 -1566
rect 5738 -1615 5801 -1566
rect 5859 -1615 5922 -1566
rect 5980 -1615 6043 -1566
rect 6101 -1615 6164 -1566
rect 6229 -1614 6292 -1565
rect 6375 -1633 6438 -1584
rect 3255 -1809 3318 -1760
rect 6375 -1740 6438 -1691
rect 3255 -1920 3318 -1871
rect 6374 -1840 6437 -1791
rect 3255 -2031 3318 -1982
rect 6374 -1951 6437 -1902
rect 6374 -2062 6437 -2013
rect 3255 -2142 3318 -2093
rect 3255 -2253 3318 -2204
rect 6374 -2173 6437 -2124
rect 3255 -2364 3318 -2315
rect 3255 -2475 3318 -2426
rect 6374 -2284 6437 -2235
rect 6374 -2395 6437 -2346
rect -236 -2598 -173 -2549
rect -108 -2599 -45 -2550
rect 21 -2598 84 -2549
rect 138 -2599 201 -2550
rect 250 -2600 313 -2551
rect 373 -2598 436 -2549
rect 502 -2597 565 -2548
rect 619 -2598 682 -2549
rect 731 -2599 794 -2550
rect 849 -2599 912 -2550
rect 975 -2598 1038 -2549
rect 1104 -2597 1167 -2548
rect 1221 -2598 1284 -2549
rect 1333 -2599 1396 -2550
rect 1451 -2599 1514 -2550
rect 1574 -2599 1637 -2550
rect 1691 -2599 1754 -2550
rect 1812 -2599 1875 -2550
rect 1934 -2599 1997 -2550
rect 2045 -2600 2108 -2551
rect 2164 -2600 2227 -2551
rect 2276 -2600 2339 -2551
rect 2397 -2600 2460 -2551
rect 2516 -2599 2579 -2550
rect 2631 -2601 2694 -2552
rect 2742 -2599 2805 -2550
rect -250 -2711 -196 -2664
rect -249 -2812 -195 -2765
rect -250 -2909 -196 -2862
rect -249 -3017 -195 -2970
rect -249 -3142 -195 -3095
rect 2753 -2697 2807 -2650
rect 2754 -2798 2808 -2751
rect 2753 -2895 2807 -2848
rect 2754 -3003 2808 -2956
rect 2754 -3128 2808 -3081
rect -248 -3256 -194 -3209
rect 2755 -3242 2809 -3195
rect -247 -3368 -193 -3321
rect -249 -3472 -195 -3425
rect -249 -3576 -195 -3529
rect 2756 -3354 2810 -3307
rect 2754 -3458 2808 -3411
rect -251 -3671 -197 -3624
rect 2754 -3562 2808 -3515
rect 2752 -3657 2806 -3610
rect -250 -3780 -196 -3733
rect -250 -3884 -196 -3837
rect 2753 -3766 2807 -3719
rect -252 -3979 -198 -3932
rect -251 -4089 -197 -4042
rect 2753 -3870 2807 -3823
rect 2751 -3965 2805 -3918
rect -251 -4193 -197 -4146
rect -253 -4288 -199 -4241
rect 2752 -4075 2806 -4028
rect 2752 -4179 2806 -4132
rect -250 -4389 -196 -4342
rect 2750 -4274 2804 -4227
rect -250 -4493 -196 -4446
rect -252 -4588 -198 -4541
rect 2753 -4375 2807 -4328
rect 2753 -4479 2807 -4432
rect 2751 -4574 2805 -4527
rect -251 -4698 -197 -4651
rect 2752 -4684 2806 -4637
rect -251 -4802 -197 -4755
rect -253 -4897 -199 -4850
rect 2752 -4788 2806 -4741
rect 2750 -4883 2804 -4836
rect -249 -5001 -195 -4954
rect -248 -5111 -194 -5064
rect 2754 -4987 2808 -4940
rect -248 -5215 -194 -5168
rect 2755 -5097 2809 -5050
rect 2755 -5201 2809 -5154
rect -239 -5335 -176 -5286
rect -111 -5336 -48 -5287
rect 18 -5335 81 -5286
rect 135 -5336 198 -5287
rect 247 -5337 310 -5288
rect 370 -5335 433 -5286
rect 499 -5334 562 -5285
rect 616 -5335 679 -5286
rect 728 -5336 791 -5287
rect 846 -5336 909 -5287
rect 972 -5335 1035 -5286
rect 1101 -5334 1164 -5285
rect 1218 -5335 1281 -5286
rect 1330 -5336 1393 -5287
rect 1448 -5336 1511 -5287
rect 1571 -5336 1634 -5287
rect 1688 -5336 1751 -5287
rect 1809 -5336 1872 -5287
rect 1931 -5336 1994 -5287
rect 2042 -5337 2105 -5288
rect 2161 -5337 2224 -5288
rect 2273 -5337 2336 -5288
rect 2394 -5337 2457 -5288
rect 2513 -5336 2576 -5287
rect 2628 -5338 2691 -5289
rect 2739 -5336 2802 -5287
rect 6374 -2506 6437 -2457
rect 3255 -2586 3318 -2537
rect 3255 -2697 3318 -2648
rect 6374 -2617 6437 -2568
rect 6374 -2728 6437 -2679
rect 3255 -2808 3318 -2759
rect 3255 -2919 3318 -2870
rect 6374 -2839 6437 -2790
rect 3255 -3030 3318 -2981
rect 3255 -3141 3318 -3092
rect 6374 -2950 6437 -2901
rect 6374 -3061 6437 -3012
rect 3255 -3252 3318 -3203
rect 6374 -3172 6437 -3123
rect 3255 -3363 3318 -3314
rect 6374 -3283 6437 -3234
rect 6374 -3394 6437 -3345
rect 3255 -3474 3318 -3425
rect 3255 -3585 3318 -3536
rect 6374 -3505 6437 -3456
rect 3255 -3696 3318 -3647
rect 6374 -3616 6437 -3567
rect 6374 -3727 6437 -3678
rect 3255 -3807 3318 -3758
rect 3255 -3918 3318 -3869
rect 3255 -4029 3318 -3980
rect 3255 -4140 3318 -4091
rect 6374 -3838 6437 -3789
rect 6374 -3949 6437 -3900
rect 6374 -4060 6437 -4011
rect 3255 -4251 3318 -4202
rect 6374 -4171 6437 -4122
rect 3255 -4362 3318 -4313
rect 3255 -4473 3318 -4424
rect 6374 -4282 6437 -4233
rect 6374 -4393 6437 -4344
rect 3255 -4584 3318 -4535
rect 3255 -4695 3318 -4646
rect 3255 -4806 3318 -4757
rect 3255 -4917 3318 -4868
rect 3255 -5028 3318 -4979
rect 3255 -5139 3318 -5090
rect 3255 -5250 3318 -5201
rect 6374 -4504 6437 -4455
rect 6374 -4615 6437 -4566
rect 6374 -4726 6437 -4677
rect 6374 -4837 6437 -4788
rect 6374 -4948 6437 -4899
rect 6374 -5059 6437 -5010
rect 6374 -5170 6437 -5121
rect 3255 -5361 3318 -5312
rect 3255 -5472 3318 -5423
rect 3255 -5583 3318 -5534
rect 3255 -5694 3318 -5645
rect 3255 -5805 3318 -5756
rect 6374 -5281 6437 -5232
rect 6374 -5392 6437 -5343
rect 6374 -5503 6437 -5454
rect 6374 -5614 6437 -5565
rect 6374 -5725 6437 -5676
rect 6374 -5836 6437 -5787
rect 3255 -5916 3318 -5867
rect 3255 -6027 3318 -5978
rect 6374 -5947 6437 -5898
rect 3255 -6138 3318 -6089
rect 3255 -6249 3318 -6200
rect 6374 -6058 6437 -6009
rect 6374 -6169 6437 -6120
rect 3255 -6360 3318 -6311
rect 6374 -6280 6437 -6231
rect 3255 -6471 3318 -6422
rect 6374 -6391 6437 -6342
rect 6374 -6502 6437 -6453
rect 3318 -6660 3381 -6611
rect 3439 -6661 3502 -6612
rect 3560 -6661 3623 -6612
rect 3681 -6661 3744 -6612
rect 3802 -6661 3865 -6612
rect 3923 -6661 3986 -6612
rect 4044 -6661 4107 -6612
rect 4165 -6661 4228 -6612
rect 4286 -6661 4349 -6612
rect 4407 -6661 4470 -6612
rect 4528 -6661 4591 -6612
rect 4649 -6661 4712 -6612
rect 4770 -6661 4833 -6612
rect 4891 -6661 4954 -6612
rect 5012 -6661 5075 -6612
rect 5133 -6661 5196 -6612
rect 5254 -6661 5317 -6612
rect 5375 -6661 5438 -6612
rect 5496 -6661 5559 -6612
rect 5617 -6661 5680 -6612
rect 5738 -6661 5801 -6612
rect 5859 -6661 5922 -6612
rect 5980 -6661 6043 -6612
rect 6101 -6661 6164 -6612
<< polysilicon >>
rect 3524 1782 3634 1795
rect 3524 1769 3542 1782
rect 3119 1710 3223 1724
rect 3119 1647 3146 1710
rect 3209 1647 3223 1710
rect 3119 1608 3223 1647
rect 3150 1606 3223 1608
rect 3480 1705 3542 1769
rect 3619 1705 3634 1782
rect 3480 1688 3634 1705
rect 3738 1769 3843 1783
rect 3738 1692 3752 1769
rect 3829 1760 3843 1769
rect 3829 1692 3879 1760
rect 3150 1559 3205 1606
rect 3480 1559 3535 1688
rect 3738 1678 3879 1692
rect 4161 1695 4247 1709
rect 4161 1684 4175 1695
rect 3820 1557 3879 1678
rect 4012 1647 4175 1684
rect 4012 1608 4112 1647
rect 4161 1637 4175 1647
rect 4233 1684 4247 1695
rect 4233 1637 4324 1684
rect 4161 1623 4324 1637
rect 4224 1608 4324 1623
rect 5007 1623 5107 1637
rect 5007 1576 5021 1623
rect 5093 1576 5107 1623
rect 5007 1542 5107 1576
rect 5559 1634 5659 1648
rect 5559 1584 5573 1634
rect 5645 1584 5659 1634
rect 5559 1542 5659 1584
rect 3482 1460 3526 1495
rect 2930 1397 3017 1411
rect 2930 1338 2944 1397
rect 3003 1387 3017 1397
rect 3003 1348 3224 1387
rect 3003 1338 3017 1348
rect 3461 1347 3556 1460
rect 3800 1449 3900 1499
rect 3671 1433 3900 1449
rect 3671 1419 3847 1433
rect 3660 1405 3847 1419
rect 3660 1347 3760 1405
rect 4795 1386 4895 1400
rect 2930 1324 3017 1338
rect 3482 1304 3526 1347
rect 3671 1304 3715 1347
rect 4795 1339 4809 1386
rect 4881 1339 4895 1386
rect 4795 1300 4895 1339
rect 5007 1300 5107 1394
rect 5347 1300 5447 1394
rect 5559 1300 5659 1395
rect 5899 1300 5999 1395
rect 5007 1145 5107 1195
rect 5357 1152 5419 1186
rect 5571 1152 5627 1188
rect 3864 1133 3964 1141
rect 4068 1133 4168 1140
rect 3864 1124 4168 1133
rect 4272 1124 4372 1140
rect 3864 1119 4372 1124
rect 3864 1071 3991 1119
rect 3067 1052 3155 1066
rect 3067 992 3081 1052
rect 3141 1044 3155 1052
rect 3977 1058 3991 1071
rect 4052 1068 4372 1119
rect 5007 1082 5241 1145
rect 4052 1058 4066 1068
rect 3977 1044 4066 1058
rect 3141 992 3190 1044
rect 5141 1022 5241 1082
rect 5351 1124 5447 1152
rect 5559 1124 5647 1152
rect 5899 1143 5999 1192
rect 5351 1039 5647 1124
rect 3067 978 3190 992
rect 3146 936 3190 978
rect 5150 969 5213 1022
rect 5351 1021 5445 1039
rect 5549 1022 5647 1039
rect 5753 1089 5999 1143
rect 5753 1022 5853 1089
rect 5562 1021 5647 1022
rect 5357 969 5419 1021
rect 5571 972 5627 1021
rect 5783 973 5837 1022
rect 3489 838 3545 865
rect 3460 824 3560 838
rect 3460 774 3474 824
rect 3546 816 3560 824
rect 3546 774 3706 816
rect 3460 760 3706 774
rect 3606 701 3706 760
rect 3814 812 3900 875
rect 4352 865 4411 885
rect 4012 812 4104 865
rect 4352 827 4452 865
rect 3814 790 4104 812
rect 3814 743 3828 790
rect 3897 743 4104 790
rect 3814 726 4104 743
rect 3814 702 3911 726
rect 4014 702 4104 726
rect 4218 768 4696 827
rect 4218 702 4318 768
rect 4637 714 4696 768
rect 4937 809 5037 823
rect 4937 757 4951 809
rect 5023 757 5037 809
rect 4937 720 5037 757
rect 5141 718 5241 814
rect 5345 719 5445 815
rect 5549 720 5649 815
rect 5753 720 5853 815
rect 3628 652 3684 701
rect 3814 637 3900 702
rect 4016 636 4104 702
rect 4254 651 4313 702
rect 4637 700 4772 714
rect 4637 639 4695 700
rect 4681 637 4695 639
rect 4758 637 4772 700
rect 4681 623 4772 637
rect 3282 501 3402 515
rect 3282 499 3296 501
rect 3197 445 3296 499
rect 3282 443 3296 445
rect 3354 499 3402 501
rect 4461 513 4505 538
rect 4461 499 4620 513
rect 3354 445 3502 499
rect 4461 445 4542 499
rect 3354 443 3368 445
rect 3282 429 3368 443
rect 4528 435 4542 445
rect 4606 435 4620 499
rect 4528 421 4620 435
rect 5141 463 5241 513
rect 5753 463 5853 513
rect 3854 414 3955 415
rect 5141 414 5853 463
rect 3854 361 4341 414
rect 3242 359 4341 361
rect 3242 306 3955 359
rect 3043 265 3135 279
rect 3043 201 3057 265
rect 3121 201 3135 265
rect 3043 176 3135 201
rect 3242 178 3343 306
rect 3446 222 3751 258
rect 3446 178 3546 222
rect 3650 178 3750 222
rect 3854 178 3955 306
rect 4286 355 4341 359
rect 4286 305 5501 355
rect 4058 290 4158 304
rect 4286 294 4608 305
rect 4058 236 4072 290
rect 4144 236 4158 290
rect 3063 131 3114 176
rect 3268 129 3323 178
rect 3868 144 3923 178
rect 4058 143 4158 236
rect 4509 142 4608 294
rect 4953 243 5040 257
rect 4953 231 4967 243
rect 4848 195 4967 231
rect 4849 184 4967 195
rect 5026 231 5040 243
rect 5026 230 5160 231
rect 5026 184 5161 230
rect 4849 170 5161 184
rect 4849 142 4949 170
rect 5061 142 5161 170
rect 5401 142 5501 305
rect 4532 95 4582 142
rect 5433 107 5483 142
rect 3276 -30 3330 7
rect 3687 -30 3741 19
rect 4540 -5 4592 42
rect 3242 -90 3341 -30
rect 2947 -120 3036 -106
rect 2947 -181 2961 -120
rect 3022 -121 3036 -120
rect 3022 -181 3115 -121
rect 3242 -144 3546 -90
rect 2947 -195 3115 -181
rect 3036 -200 3115 -195
rect 3446 -200 3546 -144
rect 3650 -94 3750 -30
rect 4509 -60 4609 -5
rect 3854 -94 3954 -93
rect 3650 -148 3954 -94
rect 4509 -112 4948 -60
rect 3854 -200 3954 -148
rect 4848 -174 4948 -112
rect 5095 -67 5152 45
rect 5612 -36 5713 3
rect 5095 -124 5489 -67
rect 5612 -82 5627 -36
rect 5699 -82 5713 -36
rect 5612 -96 5713 -82
rect 3058 -244 3102 -200
rect 3453 -249 3507 -200
rect 3882 -249 3936 -200
rect 4859 -207 4911 -174
rect 5432 -211 5489 -124
rect 3038 -479 3138 -408
rect 3242 -479 3342 -408
rect 3446 -411 3546 -408
rect 3650 -411 3750 -408
rect 3446 -460 3750 -411
rect 3446 -479 3546 -460
rect 3650 -479 3750 -460
rect 3854 -479 3954 -408
rect 4058 -409 4158 -395
rect 4058 -459 4072 -409
rect 4144 -459 4158 -409
rect 4508 -424 4608 -322
rect 4848 -344 4948 -322
rect 5060 -344 5160 -322
rect 4848 -395 5160 -344
rect 4848 -424 4948 -395
rect 5060 -424 5160 -395
rect 5400 -424 5500 -322
rect 5612 -329 5712 -315
rect 5612 -376 5626 -329
rect 5698 -376 5712 -329
rect 5612 -424 5712 -376
rect 4058 -479 4158 -459
rect 4540 -572 4588 -539
rect 4508 -620 4609 -572
rect 3243 -747 3342 -630
rect 4292 -636 4609 -620
rect 3869 -687 3922 -647
rect 4292 -684 4922 -636
rect 3854 -744 3954 -687
rect 4292 -744 4349 -684
rect 3695 -747 4349 -744
rect 3243 -800 4349 -747
rect 4874 -795 4922 -684
rect 5082 -639 5133 -556
rect 5082 -690 5500 -639
rect 5400 -750 5500 -690
rect 5423 -796 5474 -750
rect 3243 -801 3342 -800
rect 3650 -801 4349 -800
rect 3650 -857 3750 -801
rect 3666 -902 3713 -857
rect 4534 -897 4589 -847
rect 5411 -897 5466 -861
rect 3038 -1101 3138 -1049
rect 3277 -1064 3331 -1016
rect -4857 -1200 -4414 -1186
rect -4857 -1272 -4843 -1200
rect -4771 -1272 -4414 -1200
rect -4857 -1286 -4414 -1272
rect 3036 -1115 3141 -1101
rect 3036 -1192 3050 -1115
rect 3127 -1192 3141 -1115
rect 3036 -1206 3141 -1192
rect 3242 -1181 3342 -1064
rect 3545 -1065 3546 -1064
rect 3869 -1065 3923 -1023
rect 4508 -1049 4608 -897
rect 4848 -914 4948 -897
rect 5060 -914 5160 -897
rect 4848 -928 5160 -914
rect 4848 -976 4959 -928
rect 4945 -988 4959 -976
rect 5019 -976 5160 -928
rect 5019 -988 5033 -976
rect 4945 -1002 5033 -988
rect 4508 -1050 4619 -1049
rect 5400 -1050 5500 -897
rect 5612 -901 5712 -887
rect 5612 -950 5626 -901
rect 5698 -950 5712 -901
rect 5612 -964 5712 -950
rect 3446 -1068 3546 -1065
rect 3650 -1068 3750 -1065
rect 3446 -1130 3750 -1068
rect 3854 -1181 3954 -1065
rect 4058 -1072 4251 -1055
rect 4058 -1124 4170 -1072
rect 4236 -1124 4251 -1072
rect 4058 -1155 4251 -1124
rect 4508 -1105 5500 -1050
rect 3242 -1208 3954 -1181
rect 4508 -1208 4619 -1105
rect 3242 -1235 4619 -1208
rect 3854 -1308 4619 -1235
rect 3854 -1330 3954 -1308
rect 3854 -1402 3868 -1330
rect 3933 -1402 3954 -1330
rect 3854 -1416 3954 -1402
rect 3793 -1707 3893 -1670
rect 3793 -1756 3807 -1707
rect 3879 -1734 3893 -1707
rect 3879 -1756 5834 -1734
rect 3589 -1807 3689 -1770
rect 3589 -1856 3603 -1807
rect 3675 -1856 3689 -1807
rect 3589 -1870 3689 -1856
rect 3793 -1814 5834 -1756
rect 3793 -1862 3893 -1814
rect 4661 -1862 4761 -1814
rect 4865 -1862 4965 -1814
rect 5733 -1862 5833 -1814
rect 5937 -1819 6037 -1783
rect 5937 -1869 5951 -1819
rect 6023 -1869 6037 -1819
rect 5937 -1883 6037 -1869
rect 4125 -2112 4225 -2070
rect 4329 -2112 4429 -2066
rect 4125 -2122 4429 -2112
rect 5197 -2122 5297 -2070
rect 5401 -2122 5501 -2070
rect 3793 -2126 5833 -2122
rect 3793 -2184 4256 -2126
rect 4314 -2184 5833 -2126
rect 3793 -2188 5833 -2184
rect 3793 -2246 3893 -2188
rect 4242 -2198 4328 -2188
rect 4661 -2246 4761 -2188
rect 4865 -2246 4965 -2188
rect 5733 -2246 5833 -2188
rect 5937 -2449 6037 -2435
rect 4125 -2453 4426 -2450
rect 5200 -2453 5497 -2451
rect -643 -3092 -596 -3005
rect 228 -2790 2266 -2690
rect 21 -3051 121 -3037
rect 21 -3100 35 -3051
rect 107 -3100 121 -3051
rect 21 -3129 121 -3100
rect 228 -3173 325 -2790
rect 1093 -2845 1193 -2790
rect 1297 -2845 1397 -2790
rect 2166 -2848 2266 -2790
rect 556 -3053 860 -3050
rect 1628 -3053 1932 -3050
rect 556 -3129 861 -3053
rect 1093 -3129 1193 -3053
rect 1297 -3129 1397 -3053
rect 1628 -3129 1933 -3053
rect 2165 -3129 2265 -3053
rect 2369 -3063 2469 -3049
rect 2369 -3111 2383 -3063
rect 2455 -3111 2469 -3063
rect 2369 -3129 2469 -3111
rect 556 -3130 860 -3129
rect 1628 -3130 1932 -3129
rect 1629 -3131 1729 -3130
rect 1833 -3131 1932 -3130
rect 225 -3529 325 -3316
rect 761 -3385 861 -3293
rect 1629 -3385 1728 -3293
rect 760 -3453 1728 -3385
rect 1836 -3351 1933 -3266
rect 1836 -3365 2021 -3351
rect 1836 -3419 1938 -3365
rect 2007 -3419 2021 -3365
rect 1836 -3448 2021 -3419
rect 1044 -3529 1125 -3528
rect 21 -3547 121 -3533
rect 21 -3595 35 -3547
rect 107 -3595 121 -3547
rect 21 -3686 121 -3595
rect 225 -3543 1754 -3529
rect 225 -3590 851 -3543
rect 923 -3590 1754 -3543
rect 225 -3607 1754 -3590
rect 1857 -3563 1956 -3549
rect 225 -3661 325 -3607
rect 837 -3661 937 -3607
rect 1041 -3661 1141 -3607
rect 1653 -3661 1753 -3607
rect 1857 -3610 1871 -3563
rect 1942 -3610 1956 -3563
rect 1857 -3661 1956 -3610
rect 2189 -3568 2289 -3554
rect 2189 -3615 2203 -3568
rect 2275 -3615 2289 -3568
rect 2189 -3661 2289 -3615
rect 2393 -3568 2493 -3554
rect 2393 -3615 2407 -3568
rect 2479 -3615 2493 -3568
rect 2393 -3661 2493 -3615
rect 225 -3705 230 -3661
rect 428 -3913 528 -3867
rect 428 -3930 442 -3913
rect 226 -3960 442 -3930
rect 514 -3930 528 -3913
rect 633 -3930 733 -3868
rect 1245 -3930 1345 -3869
rect 1449 -3930 1549 -3869
rect 514 -3960 1753 -3930
rect 226 -3996 1753 -3960
rect 226 -4052 325 -3996
rect 837 -4050 937 -3996
rect 1041 -4050 1141 -3996
rect 1653 -4050 1753 -3996
rect 21 -4266 121 -4252
rect 21 -4315 35 -4266
rect 107 -4315 121 -4266
rect 21 -4345 121 -4315
rect 225 -4345 325 -4258
rect 429 -4263 529 -4258
rect 633 -4263 733 -4258
rect 429 -4345 733 -4263
rect 837 -4278 937 -4258
rect 1041 -4278 1141 -4258
rect 837 -4345 1141 -4278
rect 1245 -4339 1553 -4258
rect 1245 -4345 1345 -4339
rect 1449 -4345 1549 -4339
rect 1653 -4345 1753 -4258
rect 1857 -4265 1957 -4251
rect 1857 -4311 1871 -4265
rect 1943 -4311 1957 -4265
rect 1857 -4345 1957 -4311
rect 2189 -4274 2289 -4258
rect 2189 -4322 2203 -4274
rect 2275 -4322 2289 -4274
rect 2189 -4345 2289 -4322
rect 2393 -4271 2493 -4257
rect 2393 -4318 2407 -4271
rect 2479 -4318 2493 -4271
rect 2393 -4345 2493 -4318
rect 438 -4346 732 -4345
rect 846 -4361 1140 -4345
rect 633 -4601 733 -4552
rect 1245 -4601 1345 -4553
rect 165 -4615 1753 -4601
rect 165 -4687 179 -4615
rect 241 -4663 851 -4615
rect 923 -4663 1753 -4615
rect 241 -4669 1753 -4663
rect 241 -4687 325 -4669
rect 165 -4701 325 -4687
rect 225 -4730 325 -4701
rect 837 -4730 937 -4669
rect 1041 -4730 1141 -4669
rect 1653 -4730 1753 -4669
rect 21 -4983 121 -4915
rect 1461 -4938 1537 -4910
rect 429 -4966 529 -4938
rect 21 -5029 35 -4983
rect 107 -5029 121 -4983
rect 21 -5069 121 -5029
rect 373 -4980 529 -4966
rect 373 -5029 387 -4980
rect 459 -4989 529 -4980
rect 633 -4989 733 -4938
rect 1245 -4989 1345 -4938
rect 1449 -4980 1549 -4938
rect 1449 -4989 1487 -4980
rect 459 -5029 1487 -4989
rect 373 -5052 1487 -5029
rect 1535 -5052 1549 -4980
rect 1857 -4953 1957 -4938
rect 1857 -4999 1871 -4953
rect 1943 -4999 1957 -4953
rect 1857 -5039 1957 -4999
rect 2189 -4953 2289 -4938
rect 2189 -4999 2203 -4953
rect 2275 -4999 2289 -4953
rect 2189 -5039 2289 -4999
rect 2393 -4953 2493 -4938
rect 2393 -5003 2407 -4953
rect 2479 -5003 2493 -4953
rect 2393 -5039 2493 -5003
rect 373 -5066 1549 -5052
rect 3589 -2469 3689 -2453
rect 3589 -2518 3603 -2469
rect 3675 -2518 3689 -2469
rect 3589 -2536 3689 -2518
rect 3793 -2536 3893 -2453
rect 4125 -2528 4429 -2453
rect 4125 -2536 4225 -2528
rect 4329 -2536 4429 -2528
rect 4661 -2537 4761 -2454
rect 4865 -2536 4965 -2453
rect 5197 -2526 5501 -2453
rect 5197 -2536 5297 -2526
rect 5401 -2536 5501 -2526
rect 5733 -2536 5833 -2453
rect 5937 -2499 5951 -2449
rect 6023 -2499 6037 -2449
rect 5937 -2536 6037 -2499
rect 3741 -2796 3893 -2795
rect 4329 -2796 4429 -2744
rect 5197 -2796 5297 -2744
rect 3741 -2809 5833 -2796
rect 3741 -2860 3755 -2809
rect 3826 -2860 5833 -2809
rect 3741 -2867 5833 -2860
rect 3741 -2894 3893 -2867
rect 3793 -2921 3893 -2894
rect 4660 -2928 4761 -2867
rect 4864 -2934 4965 -2867
rect 5733 -2920 5833 -2867
rect 3589 -3118 3689 -3104
rect 3589 -3166 3603 -3118
rect 3675 -3166 3689 -3118
rect 3589 -3204 3689 -3166
rect 4125 -3176 4225 -3128
rect 4329 -3176 4429 -3128
rect 5197 -3176 5297 -3126
rect 5401 -3176 5501 -3127
rect 4125 -3192 5501 -3176
rect 4125 -3249 4245 -3192
rect 4305 -3249 5501 -3192
rect 5937 -3141 6037 -3127
rect 5937 -3187 5951 -3141
rect 6023 -3187 6037 -3141
rect 5937 -3201 6037 -3187
rect 4125 -3263 5501 -3249
rect 3561 -3422 3660 -3408
rect 3561 -3492 3576 -3422
rect 3646 -3445 3660 -3422
rect 3646 -3492 5321 -3445
rect 3561 -3506 5321 -3492
rect 3793 -3554 3893 -3506
rect 4405 -3554 4505 -3506
rect 4609 -3554 4709 -3506
rect 5221 -3554 5321 -3506
rect 5425 -3491 5525 -3473
rect 5425 -3541 5439 -3491
rect 5511 -3541 5525 -3491
rect 5425 -3555 5525 -3541
rect 5757 -3493 6060 -3479
rect 5757 -3540 5771 -3493
rect 5843 -3540 6060 -3493
rect 5757 -3555 6060 -3540
rect 5758 -3556 5857 -3555
rect 3505 -3762 3689 -3748
rect 3505 -3809 3519 -3762
rect 3590 -3809 3689 -3762
rect 3505 -3847 3689 -3809
rect 3997 -3812 4097 -3762
rect 4201 -3812 4301 -3762
rect 4813 -3812 4913 -3762
rect 5017 -3812 5117 -3762
rect 5560 -3812 5658 -3799
rect 3793 -3813 5658 -3812
rect 3793 -3883 5574 -3813
rect 5644 -3883 5658 -3813
rect 3793 -3885 5658 -3883
rect 3793 -3943 3893 -3885
rect 4405 -4151 4505 -3885
rect 4609 -4151 4709 -3885
rect 5221 -3943 5321 -3885
rect 5560 -3897 5658 -3885
rect 3589 -4166 3689 -4151
rect 3589 -4216 3603 -4166
rect 3675 -4216 3689 -4166
rect 3589 -4238 3689 -4216
rect 3793 -4238 3893 -4151
rect 3997 -4154 4097 -4151
rect 4201 -4154 4301 -4151
rect 3997 -4234 4301 -4154
rect 3997 -4238 4097 -4234
rect 4201 -4238 4301 -4234
rect 4405 -4236 4709 -4151
rect 4405 -4252 4505 -4236
rect 4609 -4238 4709 -4236
rect 4813 -4154 4913 -4151
rect 5017 -4154 5117 -4151
rect 4813 -4238 5117 -4154
rect 5221 -4238 5321 -4151
rect 5425 -4152 5525 -4138
rect 5425 -4203 5439 -4152
rect 5511 -4203 5525 -4152
rect 5425 -4238 5525 -4203
rect 5757 -4166 5857 -4151
rect 5757 -4216 5771 -4166
rect 5843 -4216 5857 -4166
rect 5757 -4238 5857 -4216
rect 5961 -4164 6061 -4150
rect 5961 -4211 5975 -4164
rect 6047 -4211 6061 -4164
rect 5961 -4238 6061 -4211
rect 3462 -4494 3551 -4483
rect 4201 -4494 4301 -4446
rect 4813 -4494 4913 -4446
rect 3462 -4497 5321 -4494
rect 3462 -4558 3476 -4497
rect 3537 -4558 5321 -4497
rect 3462 -4562 5321 -4558
rect 3462 -4572 3551 -4562
rect 3793 -4623 3893 -4562
rect 4096 -4831 4097 -4830
rect 3589 -4858 3688 -4831
rect 3589 -4914 3603 -4858
rect 3674 -4914 3688 -4858
rect 3589 -4950 3688 -4914
rect 3793 -4950 3892 -4831
rect 3997 -4844 4097 -4831
rect 4201 -4844 4301 -4831
rect 3997 -4943 4301 -4844
rect 3997 -4950 4097 -4943
rect 4201 -5208 4301 -4943
rect 4405 -4833 4505 -4562
rect 4609 -4833 4709 -4562
rect 5221 -4623 5321 -4562
rect 4405 -4926 4709 -4833
rect 4405 -4950 4505 -4926
rect 4609 -4950 4709 -4926
rect 4813 -4844 4913 -4831
rect 5017 -4844 5117 -4831
rect 4813 -4933 5117 -4844
rect 4813 -5208 4913 -4933
rect 5017 -4950 5117 -4933
rect 5221 -4950 5321 -4831
rect 5425 -4856 5525 -4831
rect 5425 -4907 5439 -4856
rect 5511 -4907 5525 -4856
rect 5425 -4950 5525 -4907
rect 5757 -4859 5857 -4831
rect 5757 -4908 5771 -4859
rect 5843 -4908 5857 -4859
rect 5757 -4950 5857 -4908
rect 5961 -4856 6061 -4831
rect 5961 -4903 5975 -4856
rect 6047 -4903 6061 -4856
rect 5961 -4950 6061 -4903
rect 5562 -5208 5658 -5194
rect 3793 -5276 5576 -5208
rect 5644 -5276 5658 -5208
rect 3589 -5554 3688 -5540
rect 3589 -5604 3603 -5554
rect 3674 -5604 3688 -5554
rect 3589 -5634 3688 -5604
rect 3793 -5835 3892 -5276
rect 4009 -5547 4301 -5542
rect 3997 -5616 4301 -5547
rect 3997 -5634 4097 -5616
rect 4201 -5634 4301 -5616
rect 4405 -5558 4505 -5276
rect 4609 -5558 4709 -5276
rect 4405 -5631 4709 -5558
rect 4095 -5635 4097 -5634
rect 4405 -5653 4505 -5631
rect 4609 -5644 4709 -5631
rect 4813 -5553 4913 -5547
rect 5017 -5553 5117 -5547
rect 4813 -5634 5117 -5553
rect 5221 -5832 5321 -5276
rect 5562 -5290 5658 -5276
rect 5425 -5559 5525 -5545
rect 5425 -5605 5439 -5559
rect 5511 -5605 5525 -5559
rect 5425 -5634 5525 -5605
rect 5757 -5552 5857 -5538
rect 5757 -5602 5771 -5552
rect 5843 -5602 5857 -5552
rect 5757 -5634 5857 -5602
rect 5961 -5551 6061 -5537
rect 5961 -5604 5975 -5551
rect 6047 -5604 6061 -5551
rect 5961 -5634 6061 -5604
rect 3456 -5889 3544 -5875
rect 3456 -5949 3470 -5889
rect 3530 -5891 3544 -5889
rect 4201 -5891 4301 -5842
rect 4813 -5891 4913 -5842
rect 3530 -5948 5321 -5891
rect 5515 -5925 5602 -5915
rect 3530 -5949 3544 -5948
rect 3456 -5963 3544 -5949
rect 3793 -6020 3893 -5948
rect 4405 -6019 4505 -5948
rect 4609 -6019 4709 -5948
rect 5221 -6019 5321 -5948
rect 5424 -5929 5602 -5925
rect 5424 -5988 5529 -5929
rect 5588 -5988 5602 -5929
rect 5424 -5992 5602 -5988
rect 5425 -6002 5602 -5992
rect 5755 -5962 6061 -5948
rect 5425 -6019 5526 -6002
rect 5755 -6011 5975 -5962
rect 6047 -6011 6061 -5962
rect 5755 -6018 6061 -6011
rect 5757 -6019 5857 -6018
rect 5961 -6025 6061 -6018
rect 3589 -6228 3689 -6214
rect 3589 -6280 3603 -6228
rect 3675 -6280 3689 -6228
rect 3589 -6314 3689 -6280
rect 3997 -6282 4097 -6227
rect 4201 -6282 4301 -6227
rect 4813 -6282 4913 -6226
rect 5017 -6282 5117 -6226
rect 5584 -6282 5678 -6272
rect 3997 -6286 5678 -6282
rect 3997 -6352 5598 -6286
rect 5664 -6352 5678 -6286
rect 3997 -6357 5678 -6352
rect 5584 -6366 5678 -6357
<< polycontact >>
rect 3146 1647 3209 1710
rect 3542 1705 3619 1782
rect 3752 1692 3829 1769
rect 4175 1637 4233 1695
rect 5021 1576 5093 1623
rect 5573 1584 5645 1634
rect 2944 1338 3003 1397
rect 4809 1339 4881 1386
rect 3081 992 3141 1052
rect 3991 1058 4052 1119
rect 3474 774 3546 824
rect 3828 743 3897 790
rect 4951 757 5023 809
rect 4695 637 4758 700
rect 3296 443 3354 501
rect 4542 435 4606 499
rect 3057 201 3121 265
rect 4072 236 4144 290
rect 4967 184 5026 243
rect 2961 -181 3022 -120
rect 5627 -82 5699 -36
rect 4072 -459 4144 -409
rect 5626 -376 5698 -329
rect -4843 -1272 -4771 -1200
rect 3050 -1192 3127 -1115
rect 4959 -988 5019 -928
rect 5626 -950 5698 -901
rect 4170 -1124 4236 -1072
rect 3868 -1402 3933 -1330
rect 3807 -1756 3879 -1707
rect 3603 -1856 3675 -1807
rect 5951 -1869 6023 -1819
rect 4256 -2184 4314 -2126
rect 35 -3100 107 -3051
rect 2383 -3111 2455 -3063
rect 1938 -3419 2007 -3365
rect 35 -3595 107 -3547
rect 851 -3590 923 -3543
rect 1871 -3610 1942 -3563
rect 2203 -3615 2275 -3568
rect 2407 -3615 2479 -3568
rect 442 -3960 514 -3913
rect 35 -4315 107 -4266
rect 1871 -4311 1943 -4265
rect 2203 -4322 2275 -4274
rect 2407 -4318 2479 -4271
rect 179 -4687 241 -4615
rect 851 -4663 923 -4615
rect 35 -5029 107 -4983
rect 387 -5029 459 -4980
rect 1487 -5052 1535 -4980
rect 1871 -4999 1943 -4953
rect 2203 -4999 2275 -4953
rect 2407 -5003 2479 -4953
rect 3603 -2518 3675 -2469
rect 5951 -2499 6023 -2449
rect 3755 -2860 3826 -2809
rect 3603 -3166 3675 -3118
rect 4245 -3249 4305 -3192
rect 5951 -3187 6023 -3141
rect 3576 -3492 3646 -3422
rect 5439 -3541 5511 -3491
rect 5771 -3540 5843 -3493
rect 3519 -3809 3590 -3762
rect 5574 -3883 5644 -3813
rect 3603 -4216 3675 -4166
rect 5439 -4203 5511 -4152
rect 5771 -4216 5843 -4166
rect 5975 -4211 6047 -4164
rect 3476 -4558 3537 -4497
rect 3603 -4914 3674 -4858
rect 5439 -4907 5511 -4856
rect 5771 -4908 5843 -4859
rect 5975 -4903 6047 -4856
rect 5576 -5276 5644 -5208
rect 3603 -5604 3674 -5554
rect 5439 -5605 5511 -5559
rect 5771 -5602 5843 -5552
rect 5975 -5604 6047 -5551
rect 3470 -5949 3530 -5889
rect 5529 -5988 5588 -5929
rect 5975 -6011 6047 -5962
rect 3603 -6280 3675 -6228
rect 5598 -6352 5664 -6286
<< metal1 >>
rect -2453 6690 -1670 6731
rect -2453 6561 -2381 6690
rect -2252 6561 -2101 6690
rect -1972 6561 -1815 6690
rect -1686 6561 -1670 6690
rect -2453 6544 -1670 6561
rect 5875 6549 6167 6577
rect 5875 6468 5895 6549
rect 5976 6548 6357 6549
rect 5976 6469 6068 6548
rect 6147 6469 6357 6548
rect 5976 6468 6357 6469
rect 5875 6431 6167 6468
rect 5880 5811 5996 5830
rect 5618 5730 5895 5811
rect 5976 5730 5996 5811
rect 5880 5724 5996 5730
rect 5638 5540 6233 5626
rect -5494 5092 -2371 5219
rect -3273 4876 -2364 5024
rect -5666 3848 -5181 3881
rect -5837 3847 -5337 3848
rect -5837 3724 -5652 3847
rect -5529 3724 -5337 3847
rect -5837 3723 -5337 3724
rect -5207 3723 -5181 3848
rect -5666 3696 -5181 3723
rect -3273 3126 -3125 4876
rect -2315 4785 -1674 4808
rect -2315 4656 -2304 4785
rect -2175 4656 -2083 4785
rect -1954 4656 -1825 4785
rect -1696 4656 -1674 4785
rect -2315 4641 -1674 4656
rect 5637 3897 5991 3906
rect 5633 3896 5991 3897
rect -2892 3811 -2731 3849
rect 5633 3814 5731 3896
rect 5813 3814 5894 3896
rect 5976 3814 5991 3896
rect 5633 3813 5991 3814
rect -2892 3684 -2874 3811
rect -2747 3684 -2731 3811
rect 5637 3805 5991 3813
rect -2892 3559 -2731 3684
rect 5634 3636 5831 3692
rect 5723 3599 5831 3636
rect -2892 3434 -2874 3559
rect -2749 3434 -2731 3559
rect -2892 3415 -2731 3434
rect -2875 3305 -2748 3415
rect -2875 3178 -2494 3305
rect -3273 2978 -2024 3126
rect -2172 2530 -2024 2978
rect 5775 2581 5831 3599
rect 3790 2525 5831 2581
rect 3790 2319 3846 2525
rect 4690 2344 5150 2359
rect 6147 2344 6233 5540
rect 4690 2343 6233 2344
rect 4690 2334 4865 2343
rect 3923 2319 4000 2330
rect -4196 2176 -4138 2303
rect 3790 2263 3933 2319
rect 3989 2263 4000 2319
rect 3923 2247 4000 2263
rect 4690 2269 4703 2334
rect 4766 2269 4865 2334
rect 4690 2259 4865 2269
rect 4949 2259 5063 2343
rect 5147 2259 6233 2343
rect 4690 2258 6233 2259
rect 4690 2246 5150 2258
rect 1930 2114 2220 2150
rect 1836 2113 2220 2114
rect 1836 2027 1937 2113
rect 2023 2111 2220 2113
rect 2023 2030 2130 2111
rect 2211 2030 2220 2111
rect 2023 2027 2220 2030
rect 1836 2026 2220 2027
rect 1930 2000 2220 2026
rect 6224 1999 6343 2000
rect 2654 1989 6367 1999
rect 2654 1974 6369 1989
rect 2654 1920 2690 1974
rect 2763 1920 2834 1974
rect 2907 1920 2978 1974
rect 3051 1920 3122 1974
rect 3195 1920 3266 1974
rect 3339 1920 3410 1974
rect 3483 1920 3554 1974
rect 3627 1920 3698 1974
rect 3771 1920 3842 1974
rect 3915 1920 3986 1974
rect 4059 1920 4130 1974
rect 4203 1920 4274 1974
rect 4347 1920 4418 1974
rect 4491 1920 4562 1974
rect 4635 1920 4706 1974
rect 4779 1920 4850 1974
rect 4923 1920 4994 1974
rect 5067 1920 5138 1974
rect 5211 1920 5282 1974
rect 5355 1920 5426 1974
rect 5499 1920 5570 1974
rect 5643 1920 5714 1974
rect 5787 1920 5858 1974
rect 5931 1920 6002 1974
rect 6075 1920 6146 1974
rect 6219 1920 6369 1974
rect 2654 1878 6369 1920
rect 2654 1826 2775 1878
rect 2654 1772 2678 1826
rect 2751 1772 2775 1826
rect 6223 1854 6369 1878
rect 2654 1706 2775 1772
rect 3524 1787 3636 1799
rect 3137 1712 3218 1719
rect 2654 1652 2678 1706
rect 2751 1652 2775 1706
rect -5300 1608 -5160 1626
rect -5300 1507 -5285 1608
rect -5184 1507 -5160 1608
rect -5300 1489 -5160 1507
rect 2654 1586 2775 1652
rect 2654 1532 2678 1586
rect 2751 1532 2775 1586
rect -5286 930 -5183 1489
rect 2654 1466 2775 1532
rect 3030 1710 3305 1712
rect 3030 1647 3146 1710
rect 3209 1677 3305 1710
rect 3371 1677 3429 1755
rect 3524 1700 3538 1787
rect 3625 1700 3636 1787
rect 3524 1688 3636 1700
rect 3743 1769 3838 1778
rect 5004 1775 5110 1818
rect 3743 1692 3752 1769
rect 3829 1692 3838 1769
rect 3743 1683 3838 1692
rect 3914 1756 4010 1771
rect 3914 1687 3928 1756
rect 3997 1687 4010 1756
rect 5004 1752 5019 1775
rect 3914 1686 4010 1687
rect 4166 1695 4242 1704
rect 5003 1701 5019 1752
rect 5092 1701 5110 1775
rect 4166 1686 4175 1695
rect 3914 1677 4175 1686
rect 3209 1647 3429 1677
rect 3030 1639 3429 1647
rect 3030 1499 3087 1639
rect 3137 1638 3429 1639
rect 3248 1619 3429 1638
rect 3932 1637 4175 1677
rect 4233 1686 4242 1695
rect 4233 1637 4406 1686
rect 3248 1506 3305 1619
rect 3371 1562 3429 1619
rect 3584 1621 3646 1635
rect 3584 1565 3587 1621
rect 3643 1565 3646 1621
rect 3584 1562 3646 1565
rect 3932 1631 4406 1637
rect 3716 1562 3769 1563
rect 3932 1562 3987 1631
rect 4166 1628 4242 1631
rect 3371 1511 3648 1562
rect 3712 1511 3987 1562
rect 4351 1558 4406 1631
rect 4683 1684 4786 1700
rect 4683 1623 4704 1684
rect 4765 1623 4786 1684
rect 4683 1610 4786 1623
rect 5003 1646 5110 1701
rect 3371 1500 3429 1511
rect 3584 1483 3646 1511
rect 2654 1412 2678 1466
rect 2751 1412 2775 1466
rect 3716 1412 3769 1511
rect 3932 1498 3987 1511
rect 4130 1503 4406 1558
rect 4351 1502 4406 1503
rect 2654 1346 2775 1412
rect -3986 1309 -3892 1310
rect -4078 1222 -3890 1309
rect 2654 1292 2678 1346
rect 2751 1292 2775 1346
rect 2935 1397 3012 1406
rect 2935 1338 2944 1397
rect 3003 1386 3012 1397
rect 3375 1386 3769 1412
rect 3003 1359 3769 1386
rect 4703 1396 4766 1610
rect 5003 1577 5016 1646
rect 5091 1623 5110 1646
rect 6223 1800 6254 1854
rect 6327 1800 6369 1854
rect 6223 1734 6369 1800
rect 6223 1680 6254 1734
rect 6327 1680 6369 1734
rect 5003 1576 5021 1577
rect 5093 1576 5110 1623
rect 5003 1564 5110 1576
rect 5564 1636 5656 1644
rect 5564 1634 5581 1636
rect 5643 1634 5656 1636
rect 5564 1584 5573 1634
rect 5645 1584 5656 1634
rect 5564 1574 5581 1584
rect 5643 1574 5656 1584
rect 5564 1559 5656 1574
rect 6223 1614 6369 1680
rect 6223 1560 6254 1614
rect 6327 1560 6369 1614
rect 4913 1403 4985 1506
rect 5128 1403 5191 1506
rect 4913 1396 5191 1403
rect 4703 1391 5191 1396
rect 4703 1386 5023 1391
rect 3003 1338 3428 1359
rect 2935 1334 3428 1338
rect 2935 1329 3098 1334
rect 2654 1226 2775 1292
rect -3986 1220 -3892 1222
rect -4058 966 -4012 1137
rect -2092 1028 -2034 1220
rect 2654 1172 2678 1226
rect 2751 1172 2775 1226
rect 3046 1182 3098 1329
rect 3251 1185 3303 1334
rect 3375 1183 3428 1334
rect 4703 1339 4809 1386
rect 4881 1339 5023 1386
rect 4703 1337 5023 1339
rect 5077 1390 5191 1391
rect 5077 1337 5192 1390
rect 5259 1380 5317 1501
rect 5469 1380 5527 1506
rect 5684 1380 5742 1503
rect 4703 1330 5191 1337
rect 3581 1193 3637 1309
rect 3784 1193 3837 1305
rect 3580 1189 3638 1193
rect 3578 1184 3646 1189
rect 3783 1184 3839 1193
rect 2654 1106 2775 1172
rect 3578 1128 3581 1184
rect 3637 1128 3646 1184
rect 3578 1116 3646 1128
rect 3772 1130 3784 1184
rect 3838 1171 3850 1184
rect 3993 1171 4043 1309
rect 3838 1130 4043 1171
rect 3772 1128 4043 1130
rect 3772 1121 4061 1128
rect 3772 1118 3850 1121
rect 3982 1120 4061 1121
rect 4197 1124 4247 1302
rect 4397 1132 4447 1308
rect 4703 1306 4766 1330
rect 4702 1193 4766 1306
rect 4913 1326 5191 1330
rect 4913 1198 4976 1326
rect 5128 1198 5191 1326
rect 5259 1322 5742 1380
rect 5259 1198 5317 1322
rect 5469 1203 5527 1322
rect 5684 1200 5742 1322
rect 5811 1398 5869 1498
rect 6023 1398 6081 1503
rect 5811 1389 6081 1398
rect 5811 1333 5932 1389
rect 5988 1333 6081 1389
rect 5811 1320 6081 1333
rect 4702 1132 4758 1193
rect 4397 1124 4764 1132
rect 4197 1120 4764 1124
rect 3982 1119 4764 1120
rect 2654 1052 2678 1106
rect 2751 1052 2775 1106
rect 3072 1060 3150 1061
rect 3031 1056 3150 1060
rect 3982 1058 3991 1119
rect 4052 1082 4764 1119
rect 5130 1089 5181 1198
rect 5690 1135 5739 1200
rect 5811 1195 5869 1320
rect 6023 1200 6081 1320
rect 6223 1494 6369 1560
rect 6223 1440 6254 1494
rect 6327 1440 6369 1494
rect 6223 1374 6369 1440
rect 6223 1320 6254 1374
rect 6327 1320 6369 1374
rect 6223 1254 6369 1320
rect 6223 1200 6254 1254
rect 6327 1200 6369 1254
rect 5687 1094 5747 1135
rect 6223 1134 6369 1200
rect 4052 1074 4447 1082
rect 4052 1058 4061 1074
rect 2654 986 2775 1052
rect 3030 1052 3640 1056
rect 3030 1006 3081 1052
rect 1455 966 1579 981
rect -5286 827 -4897 930
rect -4058 922 -2844 966
rect -4028 869 -2844 922
rect -543 965 1579 966
rect -543 870 1462 965
rect 1557 870 1579 965
rect -543 869 1579 870
rect 1455 853 1579 869
rect 2654 932 2678 986
rect 2751 932 2775 986
rect 2654 866 2775 932
rect 3031 992 3081 1006
rect 3141 1044 3640 1052
rect 3982 1049 4061 1058
rect 3141 1027 3650 1044
rect 3141 1006 3588 1027
rect 3141 992 3150 1006
rect 3031 983 3150 992
rect 3031 881 3083 983
rect 3251 881 3301 1006
rect 3372 875 3432 1006
rect 3576 966 3588 1006
rect 3649 966 3650 1027
rect 4258 1026 4547 1027
rect 4258 967 4270 1026
rect 4329 967 4547 1026
rect 4258 966 4338 967
rect 3576 958 3650 966
rect 3582 928 3650 958
rect 3582 927 3640 928
rect 3590 882 3640 927
rect 3711 883 4192 943
rect 4262 929 4330 966
rect 4262 928 4329 929
rect 4474 928 4547 967
rect 2654 812 2678 866
rect 2751 812 2775 866
rect 487 650 538 781
rect 895 585 945 771
rect 2654 746 2775 812
rect 3465 824 3555 833
rect 3465 805 3474 824
rect 2654 692 2678 746
rect 2751 692 2775 746
rect 3458 796 3474 805
rect 3458 723 3471 796
rect 3546 774 3555 824
rect 3884 823 3982 835
rect 3884 799 3900 823
rect 3544 765 3555 774
rect 3819 790 3900 799
rect 3544 723 3554 765
rect 3819 743 3828 790
rect 3897 754 3900 790
rect 3969 798 3982 823
rect 3969 754 3989 798
rect 3897 743 3989 754
rect 3819 735 3989 743
rect 4135 760 4190 883
rect 4269 882 4329 928
rect 4487 831 4547 928
rect 4702 831 4758 1082
rect 5130 1038 5522 1089
rect 5687 1045 5928 1094
rect 4487 776 4758 831
rect 4487 775 4544 776
rect 4602 775 4758 776
rect 4856 823 4912 983
rect 5061 831 5117 976
rect 5037 823 5117 831
rect 4856 822 5117 823
rect 4856 809 5039 822
rect 3819 734 3906 735
rect 3458 711 3554 723
rect 4135 705 4390 760
rect 4856 757 4951 809
rect 5023 757 5039 809
rect 4856 744 5039 757
rect 5102 744 5117 822
rect 4856 743 5117 744
rect 2654 626 2775 692
rect 2965 659 3024 661
rect 2654 572 2678 626
rect 2751 572 2775 626
rect 2962 645 3038 659
rect 2962 589 2971 645
rect 3027 589 3038 645
rect 2962 574 3038 589
rect 2654 506 2775 572
rect 2654 452 2678 506
rect 2751 452 2775 506
rect 2654 386 2775 452
rect 2654 332 2678 386
rect 2751 332 2775 386
rect 2654 266 2775 332
rect 2965 382 3024 574
rect 3123 497 3173 656
rect 3326 510 3376 679
rect 3925 672 3999 684
rect 3528 552 3582 659
rect 3287 501 3376 510
rect 3287 497 3296 501
rect 3123 447 3296 497
rect 3287 443 3296 447
rect 3354 497 3376 501
rect 3512 538 3588 552
rect 3512 497 3528 538
rect 3354 484 3528 497
rect 3582 484 3588 538
rect 3354 476 3588 484
rect 3735 490 3783 661
rect 3925 611 3928 672
rect 3989 611 3999 672
rect 4335 659 4390 705
rect 4675 708 4772 717
rect 3925 598 3999 611
rect 3936 543 3985 598
rect 4141 490 4189 657
rect 4335 548 4393 659
rect 4548 577 4598 656
rect 4675 629 4687 708
rect 4758 629 4772 708
rect 4675 619 4772 629
rect 3354 447 3586 476
rect 3354 443 3376 447
rect 3287 436 3376 443
rect 3735 442 4189 490
rect 4332 544 4408 548
rect 4545 544 4598 577
rect 4856 559 4912 743
rect 5037 735 5117 743
rect 5061 552 5117 735
rect 4332 539 4598 544
rect 4332 483 4342 539
rect 4398 508 4598 539
rect 5266 508 5322 978
rect 5471 666 5522 1038
rect 5461 656 5540 666
rect 5461 600 5471 656
rect 5527 600 5540 656
rect 5461 592 5540 600
rect 5471 557 5522 592
rect 4398 499 4615 508
rect 4398 494 4542 499
rect 4398 483 4408 494
rect 4332 472 4408 483
rect 3287 434 3363 436
rect 3735 382 3794 442
rect 4533 435 4542 494
rect 4606 435 4615 499
rect 5265 501 5346 508
rect 5670 501 5726 975
rect 5879 824 5928 1045
rect 6223 1080 6254 1134
rect 6327 1080 6369 1134
rect 6223 1014 6369 1080
rect 6223 960 6254 1014
rect 6327 960 6369 1014
rect 6223 894 6369 960
rect 6223 840 6254 894
rect 6327 840 6369 894
rect 5873 811 5941 824
rect 5873 755 5876 811
rect 5932 755 5941 811
rect 5873 742 5941 755
rect 6223 774 6369 840
rect 5265 499 5726 501
rect 5265 443 5278 499
rect 5334 445 5726 499
rect 5879 669 5928 742
rect 6223 720 6254 774
rect 6327 720 6369 774
rect 5334 443 5346 445
rect 5265 441 5346 443
rect 4533 426 4615 435
rect 2965 323 3794 382
rect 4529 319 5481 351
rect 5879 319 5931 669
rect 4063 290 4153 299
rect 4529 298 5931 319
rect 4063 279 4072 290
rect 2654 212 2678 266
rect 2751 212 2775 266
rect 3048 265 3130 274
rect 3048 256 3057 265
rect 2654 146 2775 212
rect -4529 109 -4127 146
rect -4529 11 -4486 109
rect -4391 100 -4127 109
rect -4391 11 -4263 100
rect -4529 4 -4263 11
rect -4162 4 -4127 100
rect -4529 -16 -4127 4
rect 2654 92 2678 146
rect 2751 92 2775 146
rect 2654 26 2775 92
rect 2654 -28 2678 26
rect 2751 -28 2775 26
rect 2960 201 3057 256
rect 3121 244 3130 265
rect 3121 201 3212 244
rect 3363 219 3828 269
rect 3363 217 3444 219
rect 2960 192 3212 201
rect 2960 15 3008 192
rect 2654 -94 2775 -28
rect 3164 -36 3212 192
rect 3350 205 3444 217
rect 3350 135 3362 205
rect 3432 135 3444 205
rect 3350 122 3444 135
rect 3778 133 3828 219
rect 3979 236 4072 279
rect 4144 236 4235 290
rect 3979 227 4235 236
rect -2913 -140 -2771 -94
rect 2654 -148 2678 -94
rect 2751 -148 2775 -94
rect 3147 -49 3228 -36
rect 3147 -105 3160 -49
rect 3216 -105 3228 -49
rect 3368 -65 3418 122
rect 3572 -56 3620 133
rect 3778 -48 3829 133
rect -3609 -319 -3562 -195
rect 2654 -214 2775 -148
rect 2952 -120 3031 -111
rect 3147 -117 3228 -105
rect 2952 -181 2961 -120
rect 3022 -181 3031 -120
rect 2952 -190 3031 -181
rect 2654 -268 2678 -214
rect 2751 -268 2775 -214
rect -2760 -375 -2714 -300
rect -2811 -421 -2714 -375
rect 2654 -334 2775 -268
rect 2654 -388 2678 -334
rect 2751 -388 2775 -334
rect 2962 -315 3010 -190
rect 3154 -235 3220 -223
rect 3154 -291 3158 -235
rect 3214 -291 3220 -235
rect 3154 -315 3220 -291
rect 2962 -316 3220 -315
rect 3369 -237 3417 -65
rect 3553 -68 3637 -56
rect 3553 -124 3568 -68
rect 3624 -124 3637 -68
rect 3553 -136 3637 -124
rect 3778 -237 3828 -48
rect 3979 -50 4031 227
rect 4185 16 4232 227
rect 4529 119 4582 298
rect 5428 267 5931 298
rect 6223 654 6369 720
rect 6223 600 6254 654
rect 6327 600 6369 654
rect 6223 534 6369 600
rect 6223 480 6254 534
rect 6327 480 6369 534
rect 6223 414 6369 480
rect 6223 360 6254 414
rect 6327 360 6369 414
rect 6223 294 6369 360
rect 4958 243 5035 252
rect 4958 184 4967 243
rect 5026 184 5035 243
rect 4958 181 4969 184
rect 5025 181 5035 184
rect 4958 175 5035 181
rect 4968 172 5026 175
rect 4490 118 4582 119
rect 4417 100 4582 118
rect 4417 97 4693 100
rect 4417 36 4421 97
rect 4482 44 4693 97
rect 5082 98 5164 108
rect 4764 93 5026 95
rect 5082 93 5094 98
rect 4482 42 4688 44
rect 4764 42 5094 93
rect 5150 93 5164 98
rect 5428 97 5481 267
rect 6223 240 6254 294
rect 6327 240 6369 294
rect 6223 174 6369 240
rect 6223 120 6254 174
rect 6327 120 6369 174
rect 5318 93 5580 97
rect 5739 93 5793 96
rect 5150 42 5239 93
rect 5318 45 5793 93
rect 5318 44 5580 45
rect 4482 36 4492 42
rect 4977 40 5239 42
rect 4417 22 4492 36
rect 5082 34 5164 40
rect 3966 -60 4045 -50
rect 3966 -116 3977 -60
rect 4033 -116 4045 -60
rect 5435 -102 5487 44
rect 5739 -27 5793 45
rect 5618 -28 5793 -27
rect 6223 54 6369 120
rect 6223 0 6254 54
rect 6327 0 6369 54
rect 5618 -36 5797 -28
rect 5618 -82 5627 -36
rect 5699 -82 5797 -36
rect 5618 -90 5797 -82
rect 6223 -66 6369 0
rect 5618 -91 5708 -90
rect 3966 -130 4045 -116
rect 5190 -154 5487 -102
rect 2962 -335 3215 -316
rect 2654 -454 2775 -388
rect 2654 -508 2678 -454
rect 2751 -508 2775 -454
rect 2654 -574 2775 -508
rect 2654 -628 2678 -574
rect 2751 -628 2775 -574
rect 2654 -694 2775 -628
rect 2961 -363 3215 -335
rect 2961 -642 3009 -363
rect 3167 -641 3213 -363
rect 3369 -642 3421 -237
rect 3572 -624 3622 -241
rect 3558 -634 3633 -624
rect 2654 -748 2678 -694
rect 2751 -748 2775 -694
rect 2654 -814 2775 -748
rect 2654 -868 2678 -814
rect 2751 -868 2775 -814
rect 3150 -782 3229 -770
rect 3150 -836 3161 -782
rect 3215 -836 3229 -782
rect 3150 -848 3229 -836
rect -1825 -1028 -1778 -927
rect 2654 -934 2775 -868
rect 2654 -988 2678 -934
rect 2751 -988 2775 -934
rect -5194 -1186 -4732 -1165
rect -6506 -1222 -6253 -1206
rect -6506 -1278 -6481 -1222
rect -6425 -1225 -6253 -1222
rect -6425 -1278 -6334 -1225
rect -6506 -1281 -6334 -1278
rect -6278 -1281 -6253 -1225
rect -6506 -1333 -6253 -1281
rect -6506 -1389 -6479 -1333
rect -6423 -1334 -6253 -1333
rect -6423 -1389 -6335 -1334
rect -6506 -1390 -6335 -1389
rect -6279 -1390 -6253 -1334
rect -6506 -1459 -6253 -1390
rect -5194 -1286 -5130 -1186
rect -5030 -1187 -4732 -1186
rect -5030 -1285 -4856 -1187
rect -4758 -1285 -4732 -1187
rect -3977 -1241 -3931 -1122
rect -5030 -1286 -4732 -1285
rect -5194 -1424 -4732 -1286
rect -3231 -1320 -3175 -1039
rect -3029 -1215 -2974 -1043
rect -2492 -1241 -2439 -1128
rect -1622 -1133 -1571 -1018
rect -2160 -1278 -2108 -1153
rect -5194 -1425 -4840 -1424
rect -5194 -1523 -5129 -1425
rect -5031 -1523 -4840 -1425
rect -5194 -1524 -4840 -1523
rect -4740 -1524 -4732 -1424
rect -5194 -1556 -4732 -1524
rect -2825 -1567 -2771 -1444
rect -1831 -1457 -1774 -1203
rect -1297 -1204 -1234 -1010
rect 2654 -1054 2775 -988
rect 2654 -1108 2678 -1054
rect 2751 -1108 2775 -1054
rect 2654 -1174 2775 -1108
rect 2964 -1100 3012 -906
rect 3165 -1100 3211 -848
rect 3369 -902 3417 -642
rect 3558 -688 3570 -634
rect 3624 -688 3633 -634
rect 3775 -642 3828 -237
rect 3962 -231 4061 -220
rect 3962 -232 4062 -231
rect 3962 -293 3973 -232
rect 4034 -293 4062 -232
rect 3962 -301 4062 -293
rect 3972 -302 4062 -301
rect 3558 -700 3633 -688
rect 3556 -789 3636 -777
rect 3556 -843 3569 -789
rect 3623 -843 3636 -789
rect 3556 -855 3636 -843
rect 3370 -903 3417 -902
rect 3370 -1020 3416 -903
rect 3573 -1020 3619 -855
rect 3778 -1022 3828 -642
rect 3981 -306 4062 -302
rect 3981 -400 4031 -306
rect 4186 -400 4233 -247
rect 3981 -409 4233 -400
rect 3981 -459 4072 -409
rect 4144 -459 4233 -409
rect 3981 -468 4233 -459
rect 3981 -646 4031 -468
rect 4186 -697 4233 -468
rect 4424 -336 4478 -221
rect 4637 -336 4691 -217
rect 4424 -390 4691 -336
rect 4424 -526 4478 -390
rect 4637 -618 4691 -390
rect 4767 -344 4819 -224
rect 4976 -344 5032 -224
rect 5190 -344 5242 -154
rect 5435 -155 5487 -154
rect 6223 -120 6254 -66
rect 6327 -120 6369 -66
rect 6223 -186 6369 -120
rect 5318 -342 5370 -220
rect 5531 -320 5583 -222
rect 5736 -320 5799 -216
rect 5531 -329 5799 -320
rect 5531 -342 5626 -329
rect 4767 -396 5244 -344
rect 5318 -376 5626 -342
rect 5698 -376 5799 -329
rect 5318 -385 5799 -376
rect 5318 -394 5583 -385
rect 4767 -526 4819 -396
rect 4976 -534 5032 -396
rect 5190 -526 5242 -396
rect 5318 -522 5370 -394
rect 5531 -467 5583 -394
rect 5527 -524 5583 -467
rect 4637 -630 4740 -618
rect 5527 -630 5581 -524
rect 5736 -527 5799 -385
rect 6223 -240 6254 -186
rect 6327 -240 6369 -186
rect 6223 -306 6369 -240
rect 6223 -360 6254 -306
rect 6327 -360 6369 -306
rect 6223 -426 6369 -360
rect 6223 -480 6254 -426
rect 6327 -480 6369 -426
rect 4637 -684 4672 -630
rect 4660 -686 4672 -684
rect 4728 -684 5581 -630
rect 6223 -546 6369 -480
rect 6223 -600 6254 -546
rect 6327 -600 6369 -546
rect 6223 -666 6369 -600
rect 4728 -686 4740 -684
rect 4660 -689 4740 -686
rect 4186 -744 4479 -697
rect 3966 -759 4044 -747
rect 3966 -813 3978 -759
rect 4032 -813 4044 -759
rect 4432 -792 4479 -744
rect 3966 -824 4044 -813
rect 3982 -891 4028 -824
rect 4417 -846 4698 -792
rect 4894 -793 4947 -684
rect 5186 -690 5306 -684
rect 6223 -720 6254 -666
rect 6327 -720 6369 -666
rect 6223 -786 6369 -720
rect 4765 -795 5027 -793
rect 5080 -794 5164 -787
rect 5080 -795 5095 -794
rect 4765 -846 5095 -795
rect 3982 -914 4029 -891
rect 3982 -1021 4030 -914
rect 2964 -1115 3211 -1100
rect 2964 -1170 3050 -1115
rect 2654 -1228 2678 -1174
rect 2751 -1228 2775 -1174
rect 3036 -1192 3050 -1170
rect 3127 -1172 3211 -1115
rect 3983 -1063 4030 -1021
rect 4186 -1063 4233 -904
rect 4557 -1053 4610 -846
rect 4977 -848 5095 -846
rect 5149 -795 5164 -794
rect 5311 -795 5581 -793
rect 5149 -848 5239 -795
rect 5311 -846 5592 -795
rect 5080 -855 5164 -848
rect 4950 -928 5028 -919
rect 4784 -930 4863 -928
rect 4784 -984 4796 -930
rect 4850 -934 4863 -930
rect 4950 -934 4959 -928
rect 4850 -980 4959 -934
rect 4850 -984 4863 -980
rect 4784 -995 4863 -984
rect 4950 -988 4959 -980
rect 5019 -988 5028 -928
rect 4950 -997 5028 -988
rect 5410 -1053 5463 -846
rect 5531 -892 5592 -846
rect 5742 -892 5794 -801
rect 5531 -893 5794 -892
rect 6223 -840 6254 -786
rect 6327 -840 6369 -786
rect 5531 -901 5800 -893
rect 5531 -950 5626 -901
rect 5698 -950 5800 -901
rect 5531 -957 5800 -950
rect 6223 -906 6369 -840
rect 5617 -959 5707 -957
rect 3983 -1072 4245 -1063
rect 3983 -1124 4170 -1072
rect 4236 -1124 4245 -1072
rect 4557 -1106 5463 -1053
rect 6223 -960 6254 -906
rect 6327 -960 6369 -906
rect 6223 -1026 6369 -960
rect 6223 -1080 6254 -1026
rect 6327 -1080 6369 -1026
rect 3983 -1129 4245 -1124
rect 3127 -1184 3227 -1172
rect 3127 -1192 3161 -1184
rect 3036 -1205 3161 -1192
rect -1623 -1349 -1572 -1250
rect 2654 -1294 2775 -1228
rect 3149 -1238 3161 -1205
rect 3215 -1190 3227 -1184
rect 3983 -1190 4029 -1129
rect 4161 -1133 4245 -1129
rect 6223 -1146 6369 -1080
rect 4661 -1186 4738 -1174
rect 4661 -1190 4673 -1186
rect 3215 -1236 4673 -1190
rect 3215 -1238 3227 -1236
rect 3149 -1250 3227 -1238
rect 4661 -1240 4673 -1236
rect 4727 -1240 4738 -1186
rect 4661 -1252 4738 -1240
rect 6223 -1200 6254 -1146
rect 6327 -1200 6369 -1146
rect 2654 -1348 2678 -1294
rect 2751 -1348 2775 -1294
rect 6223 -1266 6369 -1200
rect 2654 -1414 2775 -1348
rect 3853 -1330 3943 -1319
rect 3853 -1402 3868 -1330
rect 3933 -1402 3943 -1330
rect 3853 -1411 3943 -1402
rect 6223 -1320 6254 -1266
rect 6327 -1320 6369 -1266
rect 6223 -1386 6369 -1320
rect 2654 -1468 2678 -1414
rect 2751 -1468 2775 -1414
rect -552 -1582 -501 -1468
rect 2654 -1545 2775 -1468
rect 6223 -1440 6254 -1386
rect 6327 -1440 6369 -1386
rect 6223 -1545 6369 -1440
rect 2654 -1546 6369 -1545
rect 2654 -1547 6457 -1546
rect 2652 -1564 6457 -1547
rect 2652 -1618 2681 -1564
rect 2754 -1618 2806 -1564
rect 2879 -1618 2931 -1564
rect 3004 -1618 3056 -1564
rect 3129 -1618 3181 -1564
rect 3254 -1565 6457 -1564
rect 3254 -1614 3318 -1565
rect 3381 -1566 6229 -1565
rect 3381 -1614 3439 -1566
rect 3254 -1615 3439 -1614
rect 3502 -1615 3560 -1566
rect 3623 -1615 3681 -1566
rect 3744 -1615 3802 -1566
rect 3865 -1615 3923 -1566
rect 3986 -1615 4044 -1566
rect 4107 -1615 4165 -1566
rect 4228 -1615 4286 -1566
rect 4349 -1615 4407 -1566
rect 4470 -1615 4528 -1566
rect 4591 -1615 4649 -1566
rect 4712 -1615 4770 -1566
rect 4833 -1615 4891 -1566
rect 4954 -1615 5012 -1566
rect 5075 -1615 5133 -1566
rect 5196 -1615 5254 -1566
rect 5317 -1615 5375 -1566
rect 5438 -1615 5496 -1566
rect 5559 -1615 5617 -1566
rect 5680 -1615 5738 -1566
rect 5801 -1615 5859 -1566
rect 5922 -1615 5980 -1566
rect 6043 -1615 6101 -1566
rect 6164 -1614 6229 -1566
rect 6292 -1576 6457 -1565
rect 6292 -1584 6458 -1576
rect 6292 -1614 6375 -1584
rect 6164 -1615 6375 -1614
rect 3254 -1618 6375 -1615
rect 2652 -1631 6375 -1618
rect 2652 -1641 3339 -1631
rect -2285 -1846 -2235 -1669
rect 3231 -1760 3339 -1641
rect 6350 -1633 6375 -1631
rect 6438 -1633 6458 -1584
rect 3231 -1809 3255 -1760
rect 3318 -1809 3339 -1760
rect 3798 -1690 3888 -1678
rect 3798 -1758 3805 -1690
rect 3873 -1707 3888 -1690
rect 3879 -1756 3888 -1707
rect 6350 -1691 6458 -1633
rect 3873 -1758 3888 -1756
rect 3798 -1770 3888 -1758
rect 4990 -1783 5702 -1733
rect 3231 -1871 3339 -1809
rect 3594 -1807 3684 -1798
rect 3594 -1815 3603 -1807
rect 3524 -1827 3603 -1815
rect 3524 -1838 3536 -1827
rect 97 -2214 216 -1913
rect -6370 -2333 216 -2214
rect 97 -2522 216 -2333
rect 3231 -1920 3255 -1871
rect 3318 -1920 3339 -1871
rect 3231 -1982 3339 -1920
rect 3231 -2031 3255 -1982
rect 3318 -2031 3339 -1982
rect 3231 -2093 3339 -2031
rect 3513 -1883 3536 -1838
rect 3592 -1856 3603 -1827
rect 3675 -1838 3684 -1807
rect 3675 -1856 3972 -1838
rect 3592 -1883 3972 -1856
rect 3513 -1889 3972 -1883
rect 3513 -1895 3600 -1889
rect 3513 -2040 3564 -1895
rect 3718 -2030 3769 -1889
rect 3231 -2142 3255 -2093
rect 3318 -2142 3339 -2093
rect 3231 -2204 3339 -2142
rect 3920 -2126 3972 -1889
rect 4044 -1845 4127 -1836
rect 4786 -1841 4836 -1839
rect 4990 -1841 5040 -1783
rect 5463 -1830 5543 -1829
rect 5463 -1838 5475 -1830
rect 4254 -1845 4304 -1844
rect 4456 -1845 4506 -1844
rect 4044 -1901 4058 -1845
rect 4114 -1895 4506 -1845
rect 4114 -1901 4127 -1895
rect 4044 -1906 4127 -1901
rect 4048 -2030 4098 -1906
rect 4254 -2030 4304 -1895
rect 4456 -2032 4506 -1895
rect 4585 -1891 5040 -1841
rect 4585 -2026 4635 -1891
rect 4786 -2026 4836 -1891
rect 4990 -2022 5040 -1891
rect 5119 -1886 5475 -1838
rect 5531 -1837 5543 -1830
rect 5652 -1834 5702 -1783
rect 6350 -1740 6375 -1691
rect 6438 -1740 6458 -1691
rect 6350 -1791 6458 -1740
rect 5859 -1819 6111 -1810
rect 5859 -1834 5951 -1819
rect 5531 -1886 5578 -1837
rect 5119 -1888 5578 -1886
rect 5119 -1907 5169 -1888
rect 5117 -2031 5169 -1907
rect 5324 -2026 5374 -1888
rect 5463 -1896 5578 -1888
rect 5528 -2025 5578 -1896
rect 5652 -1869 5951 -1834
rect 6023 -1869 6111 -1819
rect 5652 -1878 6111 -1869
rect 5652 -1884 5910 -1878
rect 5652 -2015 5704 -1884
rect 4231 -2115 4325 -2106
rect 3920 -2178 4094 -2126
rect 3231 -2253 3255 -2204
rect 3318 -2253 3339 -2204
rect 3231 -2315 3339 -2253
rect 3231 -2364 3255 -2315
rect 3318 -2364 3339 -2315
rect 3231 -2426 3339 -2364
rect 3231 -2475 3255 -2426
rect 3318 -2475 3339 -2426
rect -280 -2548 2839 -2522
rect -280 -2549 502 -2548
rect -4412 -2595 -4232 -2562
rect -4412 -2733 -4396 -2595
rect -4258 -2733 -4232 -2595
rect -4412 -2857 -4232 -2733
rect -280 -2598 -236 -2549
rect -173 -2550 21 -2549
rect -173 -2598 -108 -2550
rect -280 -2599 -108 -2598
rect -45 -2598 21 -2550
rect 84 -2550 373 -2549
rect 84 -2598 138 -2550
rect -45 -2599 138 -2598
rect 201 -2551 373 -2550
rect 201 -2599 250 -2551
rect -280 -2600 250 -2599
rect 313 -2598 373 -2551
rect 436 -2597 502 -2549
rect 565 -2549 1104 -2548
rect 565 -2597 619 -2549
rect 436 -2598 619 -2597
rect 682 -2550 975 -2549
rect 682 -2598 731 -2550
rect 313 -2599 731 -2598
rect 794 -2599 849 -2550
rect 912 -2598 975 -2550
rect 1038 -2597 1104 -2549
rect 1167 -2549 2839 -2548
rect 1167 -2597 1221 -2549
rect 1038 -2598 1221 -2597
rect 1284 -2550 2839 -2549
rect 1284 -2598 1333 -2550
rect 912 -2599 1333 -2598
rect 1396 -2599 1451 -2550
rect 1514 -2599 1574 -2550
rect 1637 -2599 1691 -2550
rect 1754 -2599 1812 -2550
rect 1875 -2599 1934 -2550
rect 1997 -2551 2516 -2550
rect 1997 -2599 2045 -2551
rect 313 -2600 2045 -2599
rect 2108 -2600 2164 -2551
rect 2227 -2600 2276 -2551
rect 2339 -2600 2397 -2551
rect 2460 -2599 2516 -2551
rect 2579 -2552 2742 -2550
rect 2579 -2599 2631 -2552
rect 2460 -2600 2631 -2599
rect -280 -2601 2631 -2600
rect 2694 -2599 2742 -2552
rect 2805 -2599 2839 -2550
rect 2694 -2601 2839 -2599
rect -280 -2634 2839 -2601
rect -280 -2664 -170 -2634
rect -280 -2711 -250 -2664
rect -196 -2711 -170 -2664
rect -280 -2765 -170 -2711
rect 2724 -2650 2839 -2634
rect 2724 -2697 2753 -2650
rect 2807 -2697 2839 -2650
rect 1014 -2747 1068 -2744
rect -280 -2812 -249 -2765
rect -195 -2812 -170 -2765
rect -6301 -2858 -2458 -2857
rect -6301 -2994 -4395 -2858
rect -4259 -2874 -2458 -2858
rect -280 -2862 -170 -2812
rect -4259 -2885 -2356 -2874
rect -4259 -2886 -1667 -2885
rect -4259 -2966 -2482 -2886
rect -2399 -2966 -1667 -2886
rect -4259 -2967 -1667 -2966
rect -280 -2909 -250 -2862
rect -196 -2909 -170 -2862
rect 350 -2801 1068 -2747
rect 2724 -2751 2839 -2697
rect 2079 -2763 2155 -2752
rect -4259 -2979 -2356 -2967
rect -280 -2970 -170 -2909
rect -4259 -2994 -2458 -2979
rect -6301 -2995 -2458 -2994
rect -4412 -3023 -4232 -2995
rect -576 -3005 -473 -2992
rect -683 -3006 -473 -3005
rect -683 -3010 -569 -3006
rect -725 -3086 -569 -3010
rect -683 -3091 -569 -3086
rect -484 -3091 -473 -3006
rect -683 -3092 -473 -3091
rect -576 -3106 -473 -3092
rect -280 -3017 -249 -2970
rect -195 -3017 -170 -2970
rect -280 -3095 -170 -3017
rect -280 -3142 -249 -3095
rect -195 -3142 -170 -3095
rect -280 -3209 -170 -3142
rect -644 -3230 -557 -3221
rect -6335 -3311 -2063 -3230
rect -853 -3231 -557 -3230
rect -853 -3297 -634 -3231
rect -568 -3297 -557 -3231
rect -853 -3298 -557 -3297
rect -644 -3308 -557 -3298
rect -280 -3256 -248 -3209
rect -194 -3256 -170 -3209
rect -280 -3321 -170 -3256
rect -59 -3036 -5 -2887
rect 146 -3036 200 -2880
rect -59 -3051 200 -3036
rect -59 -3100 35 -3051
rect 107 -3052 200 -3051
rect 350 -3052 404 -2801
rect 107 -3100 404 -3052
rect -59 -3108 404 -3100
rect -59 -3113 200 -3108
rect -59 -3293 -5 -3113
rect 146 -3286 200 -3113
rect 350 -3213 404 -3108
rect 473 -3056 530 -2887
rect 677 -3056 731 -2892
rect 885 -3056 942 -2887
rect 473 -3113 942 -3056
rect 332 -3222 415 -3213
rect 332 -3279 346 -3222
rect 403 -3279 415 -3222
rect 332 -3284 415 -3279
rect 350 -3293 404 -3284
rect 473 -3294 530 -3113
rect -280 -3368 -247 -3321
rect -193 -3368 -170 -3321
rect -280 -3425 -170 -3368
rect -280 -3472 -249 -3425
rect -195 -3472 -170 -3425
rect 677 -3436 731 -3113
rect 885 -3284 942 -3113
rect 1014 -3128 1068 -2801
rect 1420 -2780 2155 -2763
rect 1420 -2817 2089 -2780
rect 1217 -3128 1271 -2947
rect 1420 -3128 1474 -2817
rect 2079 -2836 2089 -2817
rect 2145 -2836 2155 -2780
rect 2079 -2849 2155 -2836
rect 2724 -2798 2754 -2751
rect 2808 -2798 2839 -2751
rect 2724 -2848 2839 -2798
rect 1547 -3065 1601 -2890
rect 1757 -3050 1808 -2894
rect 1748 -3064 1824 -3050
rect 1748 -3065 1757 -3064
rect 1547 -3119 1757 -3065
rect 1014 -3182 1478 -3128
rect 1014 -3356 1068 -3182
rect 1217 -3353 1271 -3182
rect 1420 -3353 1474 -3182
rect 1547 -3296 1601 -3119
rect 1748 -3120 1757 -3119
rect 1813 -3065 1824 -3064
rect 1961 -3065 2014 -2891
rect 2088 -3055 2141 -2849
rect 2290 -3049 2343 -2892
rect 2496 -3049 2549 -2893
rect 2290 -3055 2549 -3049
rect 2088 -3063 2549 -3055
rect 1813 -3119 2017 -3065
rect 2088 -3108 2383 -3063
rect 1813 -3120 1824 -3119
rect 1748 -3132 1824 -3120
rect 1757 -3436 1808 -3132
rect 1961 -3291 2014 -3119
rect 2088 -3292 2141 -3108
rect 2290 -3111 2383 -3108
rect 2455 -3111 2549 -3063
rect 2290 -3125 2549 -3111
rect 2290 -3292 2343 -3125
rect 2496 -3293 2549 -3125
rect 2724 -2895 2753 -2848
rect 2807 -2895 2839 -2848
rect 2724 -2956 2839 -2895
rect 2724 -3003 2754 -2956
rect 2808 -3003 2839 -2956
rect 2724 -3081 2839 -3003
rect 2724 -3128 2754 -3081
rect 2808 -3128 2839 -3081
rect 2724 -3195 2839 -3128
rect 2724 -3242 2755 -3195
rect 2809 -3242 2839 -3195
rect 2724 -3307 2839 -3242
rect 1927 -3354 2023 -3344
rect 1927 -3365 1948 -3354
rect 2005 -3365 2023 -3354
rect 1927 -3419 1938 -3365
rect 2007 -3419 2023 -3365
rect 1927 -3434 2023 -3419
rect 2724 -3354 2756 -3307
rect 2810 -3354 2839 -3307
rect 2724 -3411 2839 -3354
rect -643 -3539 -642 -3480
rect -280 -3529 -170 -3472
rect -280 -3576 -249 -3529
rect -195 -3576 -170 -3529
rect 148 -3484 1833 -3436
rect 148 -3538 196 -3484
rect -2323 -3592 -2234 -3581
rect -2323 -3593 -1687 -3592
rect -2323 -3658 -2310 -3593
rect -2245 -3658 -1687 -3593
rect -2323 -3659 -1687 -3658
rect -280 -3624 -170 -3576
rect -2323 -3666 -2234 -3659
rect -280 -3671 -251 -3624
rect -197 -3671 -170 -3624
rect -280 -3733 -170 -3671
rect -2459 -3745 -2353 -3736
rect -2459 -3827 -2450 -3745
rect -2398 -3827 -2012 -3745
rect -280 -3780 -250 -3733
rect -196 -3780 -170 -3733
rect -2459 -3841 -2353 -3827
rect -280 -3837 -170 -3780
rect -57 -3547 196 -3538
rect -57 -3595 35 -3547
rect 107 -3595 196 -3547
rect 646 -3548 714 -3536
rect -57 -3604 196 -3595
rect -57 -3826 -6 -3604
rect 148 -3828 196 -3604
rect 347 -3549 714 -3548
rect 347 -3605 647 -3549
rect 703 -3605 714 -3549
rect 842 -3543 932 -3534
rect 842 -3590 851 -3543
rect 923 -3590 932 -3543
rect 842 -3599 932 -3590
rect 347 -3606 714 -3605
rect 347 -3817 405 -3606
rect 646 -3617 714 -3606
rect 663 -3648 714 -3617
rect 663 -3695 809 -3648
rect 558 -3771 607 -3703
rect 308 -3827 405 -3817
rect 544 -3783 616 -3771
rect -280 -3884 -250 -3837
rect -196 -3884 -170 -3837
rect -722 -3948 -517 -3884
rect -280 -3932 -170 -3884
rect -280 -3979 -252 -3932
rect -198 -3979 -170 -3932
rect -280 -4042 -170 -3979
rect -647 -4090 -547 -4078
rect -871 -4091 -547 -4090
rect -6309 -4179 -2048 -4098
rect -871 -4158 -630 -4091
rect -563 -4158 -547 -4091
rect -871 -4159 -547 -4158
rect -647 -4171 -547 -4159
rect -280 -4089 -251 -4042
rect -197 -4089 -170 -4042
rect 308 -3864 400 -3827
rect 544 -3837 556 -3783
rect 610 -3837 616 -3783
rect 544 -3850 616 -3837
rect 761 -3823 809 -3695
rect 308 -4031 355 -3864
rect 433 -3913 523 -3904
rect 433 -3960 442 -3913
rect 514 -3960 523 -3913
rect 433 -3969 523 -3960
rect 308 -4078 400 -4031
rect -280 -4146 -170 -4089
rect 150 -4090 197 -4089
rect -280 -4193 -251 -4146
rect -197 -4193 -170 -4146
rect -280 -4241 -170 -4193
rect -280 -4288 -253 -4241
rect -199 -4288 -170 -4241
rect -280 -4342 -170 -4288
rect -280 -4389 -250 -4342
rect -196 -4389 -170 -4342
rect -280 -4446 -170 -4389
rect -2322 -4462 -2233 -4459
rect -2322 -4463 -2092 -4462
rect -2322 -4530 -2310 -4463
rect -2243 -4529 -2092 -4463
rect -280 -4493 -250 -4446
rect -196 -4493 -170 -4446
rect -2243 -4530 -2233 -4529
rect -2322 -4544 -2233 -4530
rect -280 -4541 -170 -4493
rect -56 -4209 -9 -4095
rect 133 -4097 215 -4090
rect 133 -4154 146 -4097
rect 203 -4154 215 -4097
rect 133 -4165 215 -4154
rect -56 -4255 -8 -4209
rect 150 -4255 197 -4165
rect -56 -4266 197 -4255
rect -56 -4315 35 -4266
rect 107 -4315 197 -4266
rect -56 -4324 197 -4315
rect -56 -4507 -9 -4324
rect 150 -4503 197 -4324
rect -280 -4588 -252 -4541
rect -198 -4588 -170 -4541
rect -2476 -4601 -2361 -4591
rect -2476 -4602 -2359 -4601
rect -2476 -4684 -2450 -4602
rect -2398 -4684 -1955 -4602
rect -280 -4651 -170 -4588
rect -2476 -4685 -2359 -4684
rect -2476 -4698 -2361 -4685
rect -280 -4698 -251 -4651
rect -197 -4698 -170 -4651
rect -522 -4745 -447 -4733
rect -721 -4746 -447 -4745
rect -721 -4805 -517 -4746
rect -458 -4805 -447 -4746
rect -721 -4806 -447 -4805
rect -522 -4820 -447 -4806
rect -280 -4755 -170 -4698
rect 165 -4615 250 -4599
rect 165 -4618 179 -4615
rect 165 -4683 176 -4618
rect 165 -4687 179 -4683
rect 241 -4687 250 -4615
rect 165 -4699 250 -4687
rect -280 -4802 -251 -4755
rect -197 -4802 -170 -4755
rect -280 -4850 -170 -4802
rect -280 -4897 -253 -4850
rect -199 -4897 -170 -4850
rect -641 -4952 -549 -4940
rect -868 -4953 -549 -4952
rect -6287 -5039 -2110 -4967
rect -868 -5013 -630 -4953
rect -570 -5013 -549 -4953
rect -868 -5014 -549 -5013
rect -641 -5025 -549 -5014
rect -280 -4954 -170 -4897
rect -280 -5001 -249 -4954
rect -195 -5001 -170 -4954
rect -55 -4973 -6 -4775
rect 149 -4973 198 -4776
rect 353 -4896 400 -4078
rect 455 -4971 506 -3969
rect 556 -4211 603 -4022
rect 556 -4253 604 -4211
rect 556 -4265 671 -4253
rect 556 -4321 601 -4265
rect 657 -4321 671 -4265
rect 556 -4333 671 -4321
rect 556 -4507 603 -4333
rect 761 -4506 808 -3823
rect 724 -4553 808 -4506
rect 724 -4715 771 -4553
rect 863 -4606 911 -3599
rect 1033 -3634 1081 -3484
rect 1160 -3548 1233 -3535
rect 1160 -3606 1166 -3548
rect 1224 -3551 1233 -3548
rect 1224 -3603 1626 -3551
rect 1224 -3606 1233 -3603
rect 1160 -3619 1233 -3606
rect 966 -3682 1081 -3634
rect 966 -3903 1014 -3682
rect 1166 -3824 1218 -3619
rect 1365 -3781 1433 -3768
rect 966 -3951 1105 -3903
rect 1049 -3980 1105 -3951
rect 1049 -3993 1119 -3980
rect 1049 -4047 1054 -3993
rect 1108 -4047 1119 -3993
rect 1049 -4059 1119 -4047
rect 965 -4258 1012 -4096
rect 965 -4272 1049 -4258
rect 965 -4329 988 -4272
rect 1045 -4329 1049 -4272
rect 965 -4345 1049 -4329
rect 965 -4508 1012 -4345
rect 842 -4615 932 -4606
rect 842 -4663 851 -4615
rect 923 -4663 932 -4615
rect 842 -4672 932 -4663
rect 724 -4762 809 -4715
rect -280 -5064 -170 -5001
rect -56 -4983 200 -4973
rect -56 -5029 35 -4983
rect 107 -5029 200 -4983
rect -56 -5038 200 -5029
rect 372 -4980 506 -4971
rect 372 -5029 387 -4980
rect 459 -5029 506 -4980
rect 557 -4934 606 -4776
rect 761 -4898 808 -4762
rect 950 -4779 1030 -4774
rect 950 -4835 962 -4779
rect 1018 -4835 1030 -4779
rect 950 -4845 1030 -4835
rect 962 -4893 1018 -4845
rect 1170 -4896 1217 -3824
rect 1365 -3838 1368 -3781
rect 1425 -3838 1433 -3781
rect 1574 -3827 1626 -3603
rect 1785 -3554 1833 -3484
rect 2724 -3458 2754 -3411
rect 2808 -3458 2839 -3411
rect 2724 -3515 2839 -3458
rect 1985 -3554 2036 -3553
rect 1785 -3559 2036 -3554
rect 2112 -3559 2163 -3558
rect 1785 -3563 2569 -3559
rect 1785 -3610 1871 -3563
rect 1942 -3568 2569 -3563
rect 1942 -3610 2203 -3568
rect 1785 -3615 2203 -3610
rect 2275 -3615 2407 -3568
rect 2479 -3581 2569 -3568
rect 2724 -3562 2754 -3515
rect 2808 -3562 2839 -3515
rect 2479 -3615 2570 -3581
rect 1785 -3619 2570 -3615
rect 1785 -3827 1833 -3619
rect 1985 -3626 2570 -3619
rect 1985 -3823 2036 -3626
rect 2112 -3823 2163 -3626
rect 2316 -3825 2367 -3626
rect 2519 -3820 2570 -3626
rect 2724 -3610 2839 -3562
rect 2724 -3657 2752 -3610
rect 2806 -3657 2839 -3610
rect 2724 -3719 2839 -3657
rect 2724 -3766 2753 -3719
rect 2807 -3766 2839 -3719
rect 3231 -2537 3339 -2475
rect 3231 -2586 3255 -2537
rect 3318 -2586 3339 -2537
rect 3231 -2648 3339 -2586
rect 3231 -2697 3255 -2648
rect 3318 -2697 3339 -2648
rect 3231 -2759 3339 -2697
rect 3512 -2460 3561 -2293
rect 3717 -2460 3766 -2292
rect 3919 -2456 3968 -2289
rect 4042 -2294 4094 -2178
rect 4231 -2185 4244 -2115
rect 4314 -2185 4325 -2115
rect 4456 -2132 4505 -2032
rect 4456 -2181 4631 -2132
rect 5117 -2142 5166 -2031
rect 5653 -2131 5704 -2015
rect 5860 -2027 5910 -1884
rect 6061 -2030 6111 -1878
rect 6350 -1840 6374 -1791
rect 6437 -1840 6458 -1791
rect 6350 -1902 6458 -1840
rect 6350 -1951 6374 -1902
rect 6437 -1951 6458 -1902
rect 6350 -2013 6458 -1951
rect 4231 -2194 4325 -2185
rect 4042 -2402 4096 -2294
rect 3512 -2469 3766 -2460
rect 3512 -2518 3603 -2469
rect 3675 -2472 3766 -2469
rect 3862 -2469 3968 -2456
rect 3862 -2472 3875 -2469
rect 3675 -2518 3875 -2472
rect 3512 -2521 3875 -2518
rect 3512 -2527 3766 -2521
rect 3512 -2702 3561 -2527
rect 3717 -2701 3766 -2527
rect 3862 -2523 3875 -2521
rect 3929 -2472 3968 -2469
rect 4047 -2466 4096 -2402
rect 4253 -2466 4302 -2290
rect 4456 -2451 4505 -2287
rect 4419 -2463 4505 -2451
rect 4419 -2466 4431 -2463
rect 3929 -2521 3970 -2472
rect 4047 -2515 4431 -2466
rect 3929 -2523 3968 -2521
rect 3862 -2536 3968 -2523
rect 3919 -2698 3968 -2536
rect 4047 -2583 4096 -2515
rect 3231 -2808 3255 -2759
rect 3318 -2808 3339 -2759
rect 4045 -2703 4096 -2583
rect 4253 -2699 4302 -2515
rect 4419 -2517 4431 -2515
rect 4485 -2466 4505 -2463
rect 4485 -2515 4507 -2466
rect 4582 -2478 4631 -2181
rect 4990 -2191 5166 -2142
rect 5526 -2182 5704 -2131
rect 6350 -2062 6374 -2013
rect 6437 -2062 6458 -2013
rect 6350 -2124 6458 -2062
rect 6350 -2173 6374 -2124
rect 6437 -2173 6458 -2124
rect 4789 -2478 4838 -2286
rect 4990 -2478 5039 -2191
rect 5120 -2450 5170 -2289
rect 5116 -2462 5187 -2450
rect 4485 -2517 4505 -2515
rect 4419 -2529 4505 -2517
rect 4456 -2696 4505 -2529
rect 4582 -2527 5040 -2478
rect 5116 -2518 5122 -2462
rect 5178 -2475 5187 -2462
rect 5324 -2475 5373 -2291
rect 5526 -2429 5577 -2182
rect 6350 -2235 6458 -2173
rect 6350 -2284 6374 -2235
rect 6437 -2284 6458 -2235
rect 5526 -2475 5575 -2429
rect 5178 -2518 5575 -2475
rect 5116 -2524 5575 -2518
rect 5116 -2527 5187 -2524
rect 3231 -2870 3339 -2808
rect 3231 -2919 3255 -2870
rect 3318 -2919 3339 -2870
rect 3746 -2801 3846 -2789
rect 3746 -2809 3768 -2801
rect 3746 -2860 3755 -2809
rect 3746 -2868 3768 -2860
rect 3834 -2868 3846 -2801
rect 4045 -2807 4095 -2703
rect 4582 -2797 4631 -2527
rect 4789 -2695 4838 -2527
rect 3746 -2880 3846 -2868
rect 3918 -2857 4095 -2807
rect 4459 -2846 4631 -2797
rect 4990 -2816 5039 -2527
rect 5120 -2697 5169 -2527
rect 5324 -2700 5373 -2524
rect 5526 -2582 5575 -2524
rect 5655 -2450 5704 -2287
rect 5859 -2440 5908 -2288
rect 6064 -2440 6113 -2289
rect 5859 -2449 6113 -2440
rect 5655 -2463 5731 -2450
rect 5655 -2517 5666 -2463
rect 5720 -2466 5731 -2463
rect 5859 -2466 5951 -2449
rect 5720 -2499 5951 -2466
rect 6023 -2499 6113 -2449
rect 5720 -2515 6113 -2499
rect 5720 -2517 5731 -2515
rect 5655 -2529 5731 -2517
rect 5526 -2697 5581 -2582
rect 5655 -2696 5704 -2529
rect 5859 -2697 5908 -2515
rect 5531 -2804 5581 -2697
rect 6064 -2698 6113 -2515
rect 6350 -2346 6458 -2284
rect 6350 -2395 6374 -2346
rect 6437 -2395 6458 -2346
rect 6350 -2457 6458 -2395
rect 6350 -2506 6374 -2457
rect 6437 -2506 6458 -2457
rect 6350 -2568 6458 -2506
rect 6350 -2617 6374 -2568
rect 6437 -2617 6458 -2568
rect 6350 -2679 6458 -2617
rect 6350 -2728 6374 -2679
rect 6437 -2728 6458 -2679
rect 6350 -2790 6458 -2728
rect 3231 -2981 3339 -2919
rect 3231 -3030 3255 -2981
rect 3318 -3030 3339 -2981
rect 3231 -3092 3339 -3030
rect 3231 -3141 3255 -3092
rect 3318 -3141 3339 -3092
rect 3514 -3108 3564 -2965
rect 3716 -3089 3766 -2965
rect 3918 -3089 3968 -2857
rect 4048 -2909 4098 -2908
rect 4459 -2909 4508 -2846
rect 4990 -2865 5174 -2816
rect 5531 -2854 5707 -2804
rect 4048 -2958 4508 -2909
rect 4048 -3082 4098 -2958
rect 4045 -3089 4101 -3082
rect 4251 -3088 4301 -2958
rect 4457 -3072 4508 -2958
rect 4457 -3088 4507 -3072
rect 4586 -3089 4636 -2960
rect 4786 -3089 4836 -2965
rect 4992 -3089 5047 -2959
rect 5125 -2965 5174 -2865
rect 3716 -3108 3968 -3089
rect 3231 -3203 3339 -3141
rect 3511 -3118 3968 -3108
rect 3511 -3166 3603 -3118
rect 3675 -3139 3968 -3118
rect 4031 -3091 4117 -3089
rect 3675 -3166 3767 -3139
rect 4031 -3145 4046 -3091
rect 4100 -3145 4117 -3091
rect 4586 -3139 5047 -3089
rect 4031 -3160 4117 -3145
rect 3511 -3175 3767 -3166
rect 3231 -3252 3255 -3203
rect 3318 -3252 3339 -3203
rect 3231 -3314 3339 -3252
rect 4232 -3184 4326 -3180
rect 4232 -3257 4245 -3184
rect 4313 -3257 4326 -3184
rect 4997 -3205 5047 -3139
rect 5117 -3091 5174 -2965
rect 5326 -3091 5376 -2959
rect 5528 -3091 5578 -2963
rect 5117 -3141 5578 -3091
rect 5657 -3088 5707 -2854
rect 6350 -2839 6374 -2790
rect 6437 -2839 6458 -2790
rect 6350 -2901 6458 -2839
rect 6350 -2950 6374 -2901
rect 6437 -2950 6458 -2901
rect 5856 -3088 5906 -2962
rect 5657 -3097 5906 -3088
rect 5657 -3151 5762 -3097
rect 5816 -3132 5906 -3097
rect 6063 -3132 6113 -2960
rect 5816 -3141 6113 -3132
rect 5816 -3151 5951 -3141
rect 5657 -3165 5951 -3151
rect 5657 -3205 5707 -3165
rect 5861 -3187 5951 -3165
rect 6023 -3187 6113 -3141
rect 5861 -3195 6113 -3187
rect 5942 -3196 6113 -3195
rect 6350 -3012 6458 -2950
rect 6350 -3061 6374 -3012
rect 6437 -3061 6458 -3012
rect 6350 -3123 6458 -3061
rect 6350 -3172 6374 -3123
rect 6437 -3172 6458 -3123
rect 4997 -3255 5707 -3205
rect 6350 -3234 6458 -3172
rect 4232 -3269 4326 -3257
rect 3231 -3363 3255 -3314
rect 3318 -3363 3339 -3314
rect 6350 -3283 6374 -3234
rect 6437 -3283 6458 -3234
rect 6350 -3345 6458 -3283
rect 3231 -3425 3339 -3363
rect 4029 -3368 4115 -3358
rect 4029 -3388 4045 -3368
rect 3231 -3474 3255 -3425
rect 3318 -3474 3339 -3425
rect 3567 -3422 3655 -3413
rect 3567 -3438 3576 -3422
rect 3231 -3536 3339 -3474
rect 3559 -3440 3576 -3438
rect 3646 -3438 3655 -3422
rect 3715 -3424 4045 -3388
rect 4101 -3388 4115 -3368
rect 5064 -3385 5147 -3376
rect 5064 -3388 5078 -3385
rect 4101 -3424 5078 -3388
rect 3646 -3440 3665 -3438
rect 3559 -3500 3568 -3440
rect 3654 -3500 3665 -3440
rect 3559 -3511 3665 -3500
rect 3715 -3439 5078 -3424
rect 3231 -3585 3255 -3536
rect 3318 -3585 3339 -3536
rect 3231 -3647 3339 -3585
rect 3231 -3696 3255 -3647
rect 3318 -3696 3339 -3647
rect 3231 -3758 3339 -3696
rect 3512 -3708 3562 -3591
rect 3715 -3708 3766 -3439
rect 4314 -3498 4392 -3486
rect 3512 -3753 3766 -3708
rect 3919 -3499 4392 -3498
rect 3919 -3549 4326 -3499
rect 3919 -3720 3970 -3549
rect 4314 -3553 4326 -3549
rect 4380 -3553 4392 -3499
rect 4314 -3563 4392 -3553
rect 3231 -3766 3255 -3758
rect 2724 -3807 3255 -3766
rect 3318 -3807 3339 -3758
rect 2724 -3823 3339 -3807
rect 3510 -3759 3766 -3753
rect 3510 -3762 3599 -3759
rect 3510 -3809 3519 -3762
rect 3590 -3809 3599 -3762
rect 4123 -3805 4174 -3595
rect 4327 -3718 4379 -3563
rect 4530 -3711 4581 -3439
rect 5064 -3441 5078 -3439
rect 5134 -3388 5147 -3385
rect 5134 -3439 5400 -3388
rect 5134 -3441 5147 -3439
rect 5064 -3443 5147 -3441
rect 5349 -3482 5400 -3439
rect 6350 -3394 6374 -3345
rect 6437 -3394 6458 -3345
rect 6350 -3456 6458 -3394
rect 5349 -3483 5725 -3482
rect 5349 -3484 5730 -3483
rect 4730 -3494 4804 -3486
rect 5349 -3491 6138 -3484
rect 4730 -3498 5194 -3494
rect 4730 -3554 4738 -3498
rect 4794 -3545 5194 -3498
rect 4794 -3554 4804 -3545
rect 4730 -3567 4804 -3554
rect 4733 -3718 4785 -3567
rect 4938 -3597 4989 -3593
rect 4937 -3716 4989 -3597
rect 5143 -3713 5194 -3545
rect 5349 -3541 5439 -3491
rect 5511 -3493 6138 -3491
rect 5511 -3540 5771 -3493
rect 5843 -3540 6138 -3493
rect 5511 -3541 6138 -3540
rect 5349 -3549 6138 -3541
rect 5349 -3550 5730 -3549
rect 5349 -3716 5400 -3550
rect 5549 -3714 5600 -3550
rect 5679 -3714 5730 -3550
rect 5884 -3716 5935 -3549
rect 6087 -3715 6138 -3549
rect 6350 -3505 6374 -3456
rect 6437 -3505 6458 -3456
rect 6350 -3567 6458 -3505
rect 6350 -3616 6374 -3567
rect 6437 -3616 6458 -3567
rect 6350 -3678 6458 -3616
rect 3510 -3818 3599 -3809
rect 4110 -3814 4187 -3805
rect 4110 -3817 4122 -3814
rect 1365 -3850 1433 -3838
rect 1365 -3997 1432 -3984
rect 1365 -4053 1367 -3997
rect 1423 -4053 1432 -3997
rect 1365 -4067 1432 -4053
rect 1371 -4096 1420 -4067
rect 1371 -4569 1419 -4096
rect 1356 -4581 1427 -4569
rect 1356 -4635 1368 -4581
rect 1422 -4635 1427 -4581
rect 1356 -4647 1427 -4635
rect 557 -4946 716 -4934
rect 557 -5003 652 -4946
rect 709 -4955 716 -4946
rect 1369 -4955 1418 -4775
rect 1577 -4898 1624 -3827
rect 2724 -3870 2753 -3823
rect 2807 -3870 2839 -3823
rect 2724 -3918 2839 -3870
rect 2724 -3965 2751 -3918
rect 2805 -3965 2839 -3918
rect 2724 -4028 2839 -3965
rect 2724 -4075 2752 -4028
rect 2806 -4075 2839 -4028
rect 1780 -4112 1827 -4095
rect 1760 -4119 1842 -4112
rect 1760 -4176 1773 -4119
rect 1830 -4176 1842 -4119
rect 1760 -4183 1842 -4176
rect 1780 -4211 1827 -4183
rect 1780 -4256 1828 -4211
rect 1986 -4256 2033 -4095
rect 1779 -4265 2033 -4256
rect 2114 -4265 2161 -4097
rect 2318 -4262 2365 -4095
rect 2522 -4262 2569 -4091
rect 2318 -4265 2569 -4262
rect 1779 -4311 1871 -4265
rect 1943 -4271 2569 -4265
rect 1943 -4274 2407 -4271
rect 1943 -4311 2203 -4274
rect 1779 -4319 2203 -4311
rect 1780 -4321 2203 -4319
rect 1780 -4507 1827 -4321
rect 1986 -4322 2203 -4321
rect 2275 -4318 2407 -4274
rect 2479 -4318 2569 -4271
rect 2275 -4322 2569 -4318
rect 1986 -4330 2569 -4322
rect 1986 -4331 2365 -4330
rect 1986 -4507 2033 -4331
rect 2114 -4509 2161 -4331
rect 2318 -4507 2365 -4331
rect 2522 -4503 2569 -4330
rect 2724 -4132 2839 -4075
rect 2724 -4179 2752 -4132
rect 2806 -4179 2839 -4132
rect 2724 -4227 2839 -4179
rect 2724 -4274 2750 -4227
rect 2804 -4274 2839 -4227
rect 2724 -4328 2839 -4274
rect 2724 -4375 2753 -4328
rect 2807 -4375 2839 -4328
rect 2724 -4432 2839 -4375
rect 2724 -4479 2753 -4432
rect 2807 -4479 2839 -4432
rect 2724 -4527 2839 -4479
rect 2724 -4574 2751 -4527
rect 2805 -4574 2839 -4527
rect 2724 -4637 2839 -4574
rect 2724 -4684 2752 -4637
rect 2806 -4684 2839 -4637
rect 2724 -4741 2839 -4684
rect 1782 -4792 1831 -4777
rect 1764 -4795 1846 -4792
rect 1764 -4851 1777 -4795
rect 1833 -4851 1846 -4795
rect 1764 -4860 1846 -4851
rect 709 -5003 1418 -4955
rect 1782 -4943 1831 -4860
rect 1983 -4943 2034 -4757
rect 2111 -4943 2162 -4758
rect 2317 -4943 2368 -4758
rect 2521 -4943 2572 -4757
rect 1782 -4953 2572 -4943
rect 557 -5004 1418 -5003
rect 1478 -4977 1544 -4971
rect 1478 -4980 1638 -4977
rect 647 -5013 716 -5004
rect 372 -5032 506 -5029
rect 372 -5038 468 -5032
rect -280 -5111 -248 -5064
rect -194 -5111 -170 -5064
rect -280 -5168 -170 -5111
rect 149 -5110 198 -5038
rect 1478 -5052 1487 -4980
rect 1535 -4989 1638 -4980
rect 1535 -5043 1572 -4989
rect 1626 -5043 1638 -4989
rect 1535 -5052 1638 -5043
rect 1782 -4999 1871 -4953
rect 1943 -4999 2203 -4953
rect 2275 -4999 2407 -4953
rect 1782 -5003 2407 -4999
rect 2479 -5003 2572 -4953
rect 1782 -5008 2572 -5003
rect 2724 -4788 2752 -4741
rect 2806 -4788 2839 -4741
rect 2724 -4836 2839 -4788
rect 2724 -4883 2750 -4836
rect 2804 -4883 2839 -4836
rect 2724 -4940 2839 -4883
rect 2724 -4987 2754 -4940
rect 2808 -4987 2839 -4940
rect 1478 -5061 1544 -5052
rect 1782 -5110 1831 -5008
rect 2398 -5012 2488 -5008
rect 149 -5159 1831 -5110
rect 2724 -5050 2839 -4987
rect 2724 -5097 2755 -5050
rect 2809 -5097 2839 -5050
rect 2724 -5154 2839 -5097
rect -280 -5215 -248 -5168
rect -194 -5215 -170 -5168
rect -280 -5259 -170 -5215
rect 2724 -5201 2755 -5154
rect 2809 -5201 2839 -5154
rect 2724 -5259 2839 -5201
rect -280 -5285 2839 -5259
rect -280 -5286 499 -5285
rect -2326 -5312 -2231 -5307
rect -2326 -5313 -2048 -5312
rect -2326 -5380 -2310 -5313
rect -2243 -5379 -2048 -5313
rect -2243 -5380 -2231 -5379
rect -2326 -5391 -2231 -5380
rect -558 -5402 -477 -5322
rect -280 -5335 -239 -5286
rect -176 -5287 18 -5286
rect -176 -5335 -111 -5287
rect -280 -5336 -111 -5335
rect -48 -5335 18 -5287
rect 81 -5287 370 -5286
rect 81 -5335 135 -5287
rect -48 -5336 135 -5335
rect 198 -5288 370 -5287
rect 198 -5336 247 -5288
rect -280 -5337 247 -5336
rect 310 -5335 370 -5288
rect 433 -5334 499 -5286
rect 562 -5286 1101 -5285
rect 562 -5334 616 -5286
rect 433 -5335 616 -5334
rect 679 -5287 972 -5286
rect 679 -5335 728 -5287
rect 310 -5336 728 -5335
rect 791 -5336 846 -5287
rect 909 -5335 972 -5287
rect 1035 -5334 1101 -5286
rect 1164 -5286 2839 -5285
rect 1164 -5334 1218 -5286
rect 1035 -5335 1218 -5334
rect 1281 -5287 2839 -5286
rect 1281 -5335 1330 -5287
rect 909 -5336 1330 -5335
rect 1393 -5336 1448 -5287
rect 1511 -5336 1571 -5287
rect 1634 -5336 1688 -5287
rect 1751 -5336 1809 -5287
rect 1872 -5336 1931 -5287
rect 1994 -5288 2513 -5287
rect 1994 -5336 2042 -5288
rect 310 -5337 2042 -5336
rect 2105 -5337 2161 -5288
rect 2224 -5337 2273 -5288
rect 2336 -5337 2394 -5288
rect 2457 -5336 2513 -5288
rect 2576 -5289 2739 -5287
rect 2576 -5336 2628 -5289
rect 2457 -5337 2628 -5336
rect -280 -5338 2628 -5337
rect 2691 -5336 2739 -5289
rect 2802 -5336 2839 -5287
rect 2691 -5338 2839 -5336
rect -280 -5371 2839 -5338
rect 3231 -3869 3339 -3823
rect 3715 -3867 4122 -3817
rect 3231 -3918 3255 -3869
rect 3318 -3918 3339 -3869
rect 3231 -3980 3339 -3918
rect 3231 -4029 3255 -3980
rect 3318 -4029 3339 -3980
rect 3231 -4091 3339 -4029
rect 3231 -4140 3255 -4091
rect 3318 -4140 3339 -4091
rect 3231 -4202 3339 -4140
rect 3231 -4251 3255 -4202
rect 3318 -4251 3339 -4202
rect 3231 -4313 3339 -4251
rect 3231 -4362 3255 -4313
rect 3318 -4362 3339 -4313
rect 3231 -4424 3339 -4362
rect 3513 -4157 3565 -3992
rect 3716 -4157 3768 -3867
rect 4110 -3868 4122 -3867
rect 4176 -3868 4187 -3814
rect 4110 -3880 4187 -3868
rect 3513 -4166 3768 -4157
rect 3513 -4216 3603 -4166
rect 3675 -4216 3768 -4166
rect 3513 -4225 3768 -4216
rect 3513 -4402 3565 -4225
rect 3231 -4473 3255 -4424
rect 3318 -4473 3339 -4424
rect 3231 -4535 3339 -4473
rect 3231 -4584 3255 -4535
rect 3318 -4584 3339 -4535
rect 3456 -4489 3553 -4476
rect 3456 -4543 3468 -4489
rect 3545 -4543 3553 -4489
rect 3456 -4548 3476 -4543
rect 3467 -4558 3476 -4548
rect 3537 -4548 3553 -4543
rect 3537 -4558 3546 -4548
rect 3467 -4567 3546 -4558
rect 3716 -4553 3768 -4225
rect 3919 -4455 3971 -3988
rect 4327 -3990 4378 -3718
rect 4123 -4176 4175 -3995
rect 4113 -4188 4187 -4176
rect 4113 -4244 4122 -4188
rect 4178 -4244 4187 -4188
rect 4113 -4255 4187 -4244
rect 4123 -4405 4175 -4255
rect 4325 -4455 4378 -3990
rect 4517 -3949 4599 -3940
rect 4517 -4003 4530 -3949
rect 4584 -4003 4599 -3949
rect 4517 -4007 4599 -4003
rect 4733 -3981 4784 -3718
rect 4937 -3804 4988 -3716
rect 6350 -3727 6374 -3678
rect 6437 -3727 6458 -3678
rect 6350 -3789 6458 -3727
rect 4928 -3813 5009 -3804
rect 5565 -3806 5653 -3804
rect 4928 -3869 4941 -3813
rect 4997 -3817 5009 -3813
rect 5557 -3813 5662 -3806
rect 5557 -3816 5574 -3813
rect 5644 -3816 5662 -3813
rect 4997 -3867 5396 -3817
rect 4997 -3869 5009 -3867
rect 4928 -3878 5009 -3869
rect 4529 -4012 4585 -4007
rect 4530 -4399 4584 -4012
rect 3919 -4507 4378 -4455
rect 3231 -4646 3339 -4584
rect 3716 -4605 4176 -4553
rect 3231 -4695 3255 -4646
rect 3318 -4695 3339 -4646
rect 3231 -4757 3339 -4695
rect 3231 -4806 3255 -4757
rect 3318 -4806 3339 -4757
rect 3231 -4868 3339 -4806
rect 3512 -4849 3564 -4669
rect 3714 -4849 3766 -4669
rect 3231 -4917 3255 -4868
rect 3318 -4917 3339 -4868
rect 3231 -4979 3339 -4917
rect 3510 -4858 3766 -4849
rect 3510 -4914 3603 -4858
rect 3674 -4914 3766 -4858
rect 3510 -4923 3766 -4914
rect 3231 -5028 3255 -4979
rect 3318 -5028 3339 -4979
rect 3231 -5090 3339 -5028
rect 3231 -5139 3255 -5090
rect 3318 -5139 3339 -5090
rect 3512 -5112 3564 -4923
rect 3231 -5201 3339 -5139
rect 3231 -5250 3255 -5201
rect 3318 -5250 3339 -5201
rect 3231 -5312 3339 -5250
rect 3231 -5361 3255 -5312
rect 3318 -5361 3339 -5312
rect 3714 -5265 3766 -4923
rect 3918 -5160 3970 -4668
rect 4124 -4849 4176 -4605
rect 4325 -4667 4378 -4507
rect 4733 -4449 4785 -3981
rect 4937 -4165 4989 -3983
rect 4925 -4167 5007 -4165
rect 4925 -4223 4938 -4167
rect 4994 -4223 5007 -4167
rect 4925 -4225 5007 -4223
rect 4937 -4227 4994 -4225
rect 4937 -4393 4989 -4227
rect 5140 -4449 5192 -3983
rect 4733 -4501 5192 -4449
rect 5344 -4143 5396 -3867
rect 5557 -3891 5566 -3816
rect 5652 -3891 5662 -3816
rect 5557 -3903 5662 -3891
rect 6350 -3838 6374 -3789
rect 6437 -3838 6458 -3789
rect 6350 -3900 6458 -3838
rect 6350 -3949 6374 -3900
rect 6437 -3949 6458 -3900
rect 5550 -4143 5602 -3981
rect 5344 -4152 5602 -4143
rect 5344 -4203 5439 -4152
rect 5511 -4155 5602 -4152
rect 5677 -4153 5729 -3985
rect 5677 -4155 5818 -4153
rect 5881 -4155 5933 -3984
rect 6086 -4155 6138 -3985
rect 5511 -4162 6138 -4155
rect 5511 -4203 5761 -4162
rect 5817 -4164 6138 -4162
rect 5817 -4166 5975 -4164
rect 5344 -4212 5761 -4203
rect 4733 -4665 4785 -4501
rect 5344 -4552 5396 -4212
rect 5550 -4218 5761 -4212
rect 5843 -4211 5975 -4166
rect 6047 -4211 6138 -4164
rect 5843 -4216 6138 -4211
rect 5817 -4218 6138 -4216
rect 5550 -4220 6138 -4218
rect 5550 -4225 5933 -4220
rect 5550 -4391 5602 -4225
rect 5677 -4227 5818 -4225
rect 5677 -4395 5729 -4227
rect 5881 -4394 5933 -4225
rect 6086 -4395 6138 -4220
rect 6350 -4011 6458 -3949
rect 6350 -4060 6374 -4011
rect 6437 -4060 6458 -4011
rect 6350 -4122 6458 -4060
rect 6350 -4171 6374 -4122
rect 6437 -4171 6458 -4122
rect 6350 -4233 6458 -4171
rect 6350 -4282 6374 -4233
rect 6437 -4282 6458 -4233
rect 6350 -4344 6458 -4282
rect 6350 -4393 6374 -4344
rect 6437 -4393 6458 -4344
rect 4123 -4854 4181 -4849
rect 4324 -4854 4378 -4667
rect 4120 -4858 4190 -4854
rect 4323 -4855 4379 -4854
rect 4120 -4914 4124 -4858
rect 4180 -4914 4190 -4858
rect 4120 -4919 4190 -4914
rect 4311 -4863 4391 -4855
rect 4311 -4917 4324 -4863
rect 4378 -4917 4391 -4863
rect 4123 -4923 4181 -4919
rect 4311 -4920 4391 -4917
rect 4124 -5112 4176 -4923
rect 4323 -4926 4379 -4920
rect 4324 -5110 4378 -4926
rect 4326 -5160 4378 -5110
rect 3918 -5212 4378 -5160
rect 4529 -5265 4581 -4667
rect 4732 -4793 4785 -4665
rect 4939 -4604 5396 -4552
rect 6350 -4455 6458 -4393
rect 6350 -4504 6374 -4455
rect 6437 -4504 6458 -4455
rect 6350 -4566 6458 -4504
rect 4939 -4666 4991 -4604
rect 6350 -4615 6374 -4566
rect 6437 -4615 6458 -4566
rect 4732 -5160 4784 -4793
rect 4938 -4805 4991 -4666
rect 4938 -5109 4990 -4805
rect 5144 -4994 5196 -4667
rect 5346 -4846 5398 -4665
rect 5549 -4846 5601 -4666
rect 5678 -4846 5730 -4666
rect 5346 -4848 5730 -4846
rect 5886 -4847 5938 -4666
rect 6086 -4847 6138 -4663
rect 5882 -4848 6138 -4847
rect 5346 -4849 6138 -4848
rect 5333 -4856 6138 -4849
rect 5333 -4864 5439 -4856
rect 5333 -4918 5345 -4864
rect 5399 -4907 5439 -4864
rect 5511 -4859 5975 -4856
rect 5511 -4907 5771 -4859
rect 5399 -4908 5771 -4907
rect 5843 -4903 5975 -4859
rect 6047 -4903 6138 -4856
rect 5843 -4908 6138 -4903
rect 5399 -4912 6138 -4908
rect 5399 -4916 5938 -4912
rect 5399 -4918 5412 -4916
rect 5333 -4929 5412 -4918
rect 5346 -4991 5398 -4929
rect 5144 -5110 5200 -4994
rect 5346 -5108 5399 -4991
rect 5148 -5160 5200 -5110
rect 4732 -5212 5200 -5160
rect 5347 -5265 5399 -5108
rect 5549 -5109 5601 -4916
rect 5678 -4917 5938 -4916
rect 5678 -5109 5730 -4917
rect 5886 -5109 5938 -4917
rect 6086 -5106 6138 -4912
rect 6350 -4677 6458 -4615
rect 6350 -4726 6374 -4677
rect 6437 -4726 6458 -4677
rect 6350 -4788 6458 -4726
rect 6350 -4837 6374 -4788
rect 6437 -4837 6458 -4788
rect 6350 -4899 6458 -4837
rect 6350 -4948 6374 -4899
rect 6437 -4948 6458 -4899
rect 6350 -5010 6458 -4948
rect 6350 -5059 6374 -5010
rect 6437 -5059 6458 -5010
rect 6350 -5121 6458 -5059
rect 6350 -5170 6374 -5121
rect 6437 -5170 6458 -5121
rect 3714 -5317 5399 -5265
rect 5559 -5200 5662 -5185
rect 5559 -5267 5568 -5200
rect 5652 -5267 5662 -5200
rect 5559 -5276 5576 -5267
rect 5644 -5276 5662 -5267
rect 5559 -5279 5662 -5276
rect 6350 -5232 6458 -5170
rect 5567 -5285 5653 -5279
rect 6350 -5281 6374 -5232
rect 6437 -5281 6458 -5232
rect 3231 -5423 3339 -5361
rect 3231 -5472 3255 -5423
rect 3318 -5472 3339 -5423
rect -2463 -5492 -2356 -5486
rect -4255 -5574 -2450 -5492
rect -2398 -5574 -1999 -5492
rect -839 -5534 -454 -5479
rect 779 -5552 1133 -5497
rect 3231 -5534 3339 -5472
rect -4255 -5593 -2356 -5574
rect 3231 -5583 3255 -5534
rect 3318 -5583 3339 -5534
rect -4255 -5610 -2368 -5593
rect -5020 -5814 -4689 -5791
rect -6230 -5815 -4689 -5814
rect -6230 -5900 -4998 -5815
rect -5020 -5920 -4998 -5900
rect -4893 -5920 -4807 -5815
rect -5020 -5922 -4807 -5920
rect -4700 -5922 -4689 -5815
rect -5020 -5933 -4689 -5922
rect -5152 -6332 -4899 -6323
rect -6266 -6345 -4899 -6332
rect -6266 -6406 -5150 -6345
rect -5089 -6406 -4986 -6345
rect -6266 -6408 -4986 -6406
rect -4923 -6408 -4899 -6345
rect -6266 -6417 -4899 -6408
rect -5152 -6425 -4899 -6417
rect -5152 -6535 -4929 -6511
rect -6271 -6536 -5014 -6535
rect -6271 -6604 -5138 -6536
rect -5070 -6604 -5014 -6536
rect -6271 -6605 -5014 -6604
rect -4944 -6605 -4929 -6535
rect -6271 -6618 -4929 -6605
rect -5152 -6626 -4929 -6618
rect -4255 -7905 -4137 -5610
rect 3231 -5645 3339 -5583
rect 3231 -5694 3255 -5645
rect 3318 -5694 3339 -5645
rect 3231 -5756 3339 -5694
rect 3231 -5805 3255 -5756
rect 3318 -5805 3339 -5756
rect 3511 -5545 3564 -5379
rect 3716 -5545 3769 -5382
rect 3511 -5553 3769 -5545
rect 3511 -5554 3781 -5553
rect 3511 -5604 3603 -5554
rect 3674 -5562 3781 -5554
rect 3674 -5604 3716 -5562
rect 3511 -5613 3716 -5604
rect 3511 -5798 3564 -5613
rect 3706 -5616 3716 -5613
rect 3770 -5616 3781 -5562
rect 3706 -5626 3781 -5616
rect -2654 -5831 -2404 -5815
rect -761 -5827 -682 -5814
rect -2654 -5903 -2636 -5831
rect -2564 -5832 -2070 -5831
rect -2564 -5902 -2487 -5832
rect -2417 -5902 -2070 -5832
rect -869 -5881 -749 -5827
rect -695 -5881 -682 -5827
rect -761 -5893 -682 -5881
rect -2564 -5903 -2070 -5902
rect -623 -5903 -501 -5825
rect -2654 -5922 -2404 -5903
rect -623 -5949 -545 -5903
rect 968 -5906 1164 -5825
rect 3231 -5867 3339 -5805
rect 3231 -5916 3255 -5867
rect 3318 -5916 3339 -5867
rect 3231 -5978 3339 -5916
rect 3458 -5882 3539 -5872
rect 3458 -5944 3469 -5882
rect 3531 -5944 3539 -5882
rect 3458 -5949 3470 -5944
rect 3530 -5949 3539 -5944
rect 3461 -5958 3539 -5949
rect 3716 -5952 3769 -5626
rect 3919 -5844 3972 -5378
rect 4122 -5798 4175 -5317
rect 4328 -5569 4381 -5381
rect 4310 -5572 4388 -5569
rect 4310 -5628 4323 -5572
rect 4379 -5628 4388 -5572
rect 4310 -5637 4388 -5628
rect 4326 -5797 4381 -5637
rect 4326 -5844 4380 -5797
rect 4531 -5814 4584 -5378
rect 4733 -5563 4786 -5375
rect 4937 -5549 4990 -5317
rect 6350 -5343 6458 -5281
rect 4936 -5555 4992 -5549
rect 4924 -5558 5005 -5555
rect 4728 -5574 4800 -5563
rect 4728 -5630 4734 -5574
rect 4790 -5630 4800 -5574
rect 4924 -5612 4937 -5558
rect 4991 -5612 5005 -5558
rect 4924 -5617 5005 -5612
rect 4936 -5621 4992 -5617
rect 4728 -5641 4800 -5630
rect 4530 -5818 4586 -5814
rect 3919 -5897 4380 -5844
rect 4519 -5823 4597 -5818
rect 4519 -5877 4531 -5823
rect 4585 -5877 4597 -5823
rect 4519 -5885 4597 -5877
rect 4733 -5843 4786 -5641
rect 4937 -5789 4990 -5621
rect 5142 -5843 5195 -5374
rect 4530 -5886 4586 -5885
rect 4109 -5952 4189 -5943
rect 3231 -6027 3255 -5978
rect 3318 -6027 3339 -5978
rect 3716 -6005 4121 -5952
rect 4109 -6008 4121 -6005
rect 4177 -6008 4189 -5952
rect 4109 -6018 4189 -6008
rect 3231 -6089 3339 -6027
rect 3231 -6138 3255 -6089
rect 3318 -6138 3339 -6089
rect -2323 -6185 -2232 -6180
rect -2323 -6186 -2060 -6185
rect -2323 -6253 -2310 -6186
rect -2243 -6252 -2060 -6186
rect -2243 -6253 -2232 -6252
rect -2323 -6264 -2232 -6253
rect -1779 -7067 -1666 -6164
rect -838 -6253 -497 -6199
rect -131 -7060 -18 -6164
rect 780 -6258 1127 -6204
rect 1514 -7075 1627 -6164
rect 3231 -6193 3339 -6138
rect 2389 -6200 3339 -6193
rect 2389 -6247 3255 -6200
rect 3231 -6249 3255 -6247
rect 3318 -6249 3339 -6200
rect 3231 -6311 3339 -6249
rect 3512 -6217 3563 -6053
rect 3716 -6217 3767 -6056
rect 3512 -6228 3767 -6217
rect 3512 -6280 3603 -6228
rect 3675 -6280 3767 -6228
rect 3512 -6290 3767 -6280
rect 3920 -6230 3971 -6058
rect 4123 -6178 4177 -6018
rect 4329 -6057 4380 -5897
rect 4327 -6180 4380 -6057
rect 4733 -5896 5195 -5843
rect 5348 -5549 5401 -5376
rect 5550 -5549 5603 -5382
rect 5678 -5542 5731 -5384
rect 5882 -5542 5935 -5384
rect 6085 -5542 6138 -5383
rect 5678 -5549 6138 -5542
rect 5348 -5551 6138 -5549
rect 5348 -5552 5975 -5551
rect 5348 -5559 5771 -5552
rect 5348 -5605 5439 -5559
rect 5511 -5602 5771 -5559
rect 5843 -5602 5975 -5552
rect 5511 -5604 5975 -5602
rect 6047 -5604 6138 -5551
rect 5511 -5605 6138 -5604
rect 5348 -5612 6138 -5605
rect 5348 -5614 5731 -5612
rect 4329 -6230 4380 -6180
rect 3920 -6281 4380 -6230
rect 3512 -6291 3563 -6290
rect 3231 -6360 3255 -6311
rect 3318 -6360 3339 -6311
rect 3231 -6422 3339 -6360
rect 3716 -6328 3767 -6290
rect 4531 -6328 4582 -6058
rect 4733 -6060 4786 -5896
rect 5348 -5944 5401 -5614
rect 5550 -5789 5603 -5614
rect 5678 -5791 5731 -5614
rect 5882 -5613 6138 -5612
rect 5882 -5791 5935 -5613
rect 6085 -5790 6138 -5613
rect 6350 -5392 6374 -5343
rect 6437 -5392 6458 -5343
rect 6350 -5454 6458 -5392
rect 6350 -5503 6374 -5454
rect 6437 -5503 6458 -5454
rect 6350 -5565 6458 -5503
rect 6350 -5614 6374 -5565
rect 6437 -5614 6458 -5565
rect 6350 -5676 6458 -5614
rect 6350 -5725 6374 -5676
rect 6437 -5725 6458 -5676
rect 6350 -5787 6458 -5725
rect 6350 -5836 6374 -5787
rect 6437 -5836 6458 -5787
rect 6350 -5898 6458 -5836
rect 4926 -5953 5401 -5944
rect 4926 -6007 4938 -5953
rect 4992 -5997 5401 -5953
rect 5520 -5929 5601 -5920
rect 5520 -5988 5529 -5929
rect 5588 -5950 5601 -5929
rect 6350 -5947 6374 -5898
rect 6437 -5947 6458 -5898
rect 5588 -5962 6137 -5950
rect 5588 -5988 5975 -5962
rect 5520 -5997 5975 -5988
rect 4992 -6007 5004 -5997
rect 4926 -6019 5004 -6007
rect 5550 -6011 5975 -5997
rect 6047 -6011 6137 -5962
rect 4733 -6231 4789 -6060
rect 4938 -6185 4991 -6019
rect 5550 -6021 6137 -6011
rect 5349 -6056 5400 -6052
rect 5144 -6231 5195 -6058
rect 5347 -6179 5400 -6056
rect 5550 -6179 5601 -6021
rect 4733 -6282 5195 -6231
rect 5349 -6328 5400 -6179
rect 5679 -6183 5730 -6021
rect 3716 -6375 5400 -6328
rect 3716 -6379 4936 -6375
rect 3231 -6471 3255 -6422
rect 3318 -6471 3339 -6422
rect 4922 -6431 4936 -6379
rect 4992 -6379 5400 -6375
rect 4992 -6431 5005 -6379
rect 4922 -6437 5005 -6431
rect 5349 -6436 5400 -6379
rect 5561 -6286 5676 -6277
rect 5561 -6294 5598 -6286
rect 5561 -6363 5576 -6294
rect 5664 -6352 5676 -6286
rect 5645 -6363 5676 -6352
rect 5561 -6381 5676 -6363
rect 5883 -6436 5934 -6021
rect 6086 -6180 6137 -6021
rect 6350 -6009 6458 -5947
rect 6350 -6058 6374 -6009
rect 6437 -6058 6458 -6009
rect 6350 -6120 6458 -6058
rect 6350 -6169 6374 -6120
rect 6437 -6169 6458 -6120
rect 3231 -6591 3339 -6471
rect 5349 -6487 5934 -6436
rect 5883 -6489 5934 -6487
rect 6350 -6231 6458 -6169
rect 6350 -6280 6374 -6231
rect 6437 -6280 6458 -6231
rect 6350 -6342 6458 -6280
rect 6350 -6391 6374 -6342
rect 6437 -6391 6458 -6342
rect 6350 -6453 6458 -6391
rect 6350 -6502 6374 -6453
rect 6437 -6502 6458 -6453
rect 6350 -6591 6458 -6502
rect 3231 -6611 6461 -6591
rect 3231 -6660 3318 -6611
rect 3381 -6612 6461 -6611
rect 3381 -6660 3439 -6612
rect 3231 -6661 3439 -6660
rect 3502 -6661 3560 -6612
rect 3623 -6661 3681 -6612
rect 3744 -6661 3802 -6612
rect 3865 -6661 3923 -6612
rect 3986 -6661 4044 -6612
rect 4107 -6661 4165 -6612
rect 4228 -6661 4286 -6612
rect 4349 -6661 4407 -6612
rect 4470 -6661 4528 -6612
rect 4591 -6661 4649 -6612
rect 4712 -6661 4770 -6612
rect 4833 -6661 4891 -6612
rect 4954 -6661 5012 -6612
rect 5075 -6661 5133 -6612
rect 5196 -6661 5254 -6612
rect 5317 -6661 5375 -6612
rect 5438 -6661 5496 -6612
rect 5559 -6661 5617 -6612
rect 5680 -6661 5738 -6612
rect 5801 -6661 5859 -6612
rect 5922 -6661 5980 -6612
rect 6043 -6661 6101 -6612
rect 6164 -6661 6461 -6612
rect 3231 -6677 6461 -6661
rect 3231 -7072 3339 -6677
rect 6272 -6678 6461 -6677
rect -3839 -7368 -3532 -7333
rect -3839 -7456 -3822 -7368
rect -3734 -7369 -2830 -7368
rect -3734 -7455 -3638 -7369
rect -3552 -7455 -2830 -7369
rect -2553 -7416 -2507 -7293
rect -3734 -7456 -2830 -7455
rect -3839 -7472 -3532 -7456
rect -4255 -8023 -3568 -7905
rect -3686 -8178 -3568 -8023
rect -3690 -8198 -3330 -8178
rect -3690 -8299 -3675 -8198
rect -3574 -8299 -3330 -8198
rect -3690 -8329 -3330 -8299
rect -2327 -8216 -1628 -8190
rect -2327 -8217 -1777 -8216
rect -2327 -8222 -2006 -8217
rect -2327 -8344 -2276 -8222
rect -2141 -8339 -2006 -8222
rect -1871 -8338 -1777 -8217
rect -1642 -8338 -1628 -8216
rect -1871 -8339 -1628 -8338
rect -2141 -8344 -1628 -8339
rect -2327 -8367 -1628 -8344
rect -3067 -8644 -2850 -8574
rect -2164 -8999 -1783 -8916
rect -2601 -9819 -2555 -9786
rect -2261 -11457 -2256 -11452
rect -2329 -11503 -2256 -11457
rect -2261 -11508 -2256 -11503
rect -2194 -11508 -2189 -11452
rect -3469 -12152 -3160 -12130
rect -3700 -12153 -3160 -12152
rect -3700 -12246 -3459 -12153
rect -3366 -12155 -3160 -12153
rect -3366 -12245 -3283 -12155
rect -3193 -12245 -3160 -12155
rect -3366 -12246 -3160 -12245
rect -3700 -12247 -3160 -12246
rect -3469 -12274 -3160 -12247
rect -3490 -12385 -3139 -12343
rect -3565 -12386 -3266 -12385
rect -3565 -12387 -3479 -12386
rect -3714 -12472 -3479 -12387
rect -3393 -12472 -3266 -12386
rect -3714 -12473 -3266 -12472
rect -3178 -12473 -3139 -12385
rect -3490 -12515 -3139 -12473
<< via1 >>
rect -2381 6561 -2252 6690
rect -2101 6561 -1972 6690
rect -1815 6561 -1686 6690
rect 5895 6468 5976 6549
rect 6068 6469 6147 6548
rect 5895 5730 5976 5811
rect -5652 3724 -5529 3847
rect -5337 3723 -5207 3848
rect -2304 4656 -2175 4785
rect -2083 4656 -1954 4785
rect -1825 4656 -1696 4785
rect 5731 3814 5813 3896
rect 5894 3814 5976 3896
rect -2874 3684 -2747 3811
rect -2874 3434 -2749 3559
rect 3933 2263 3989 2319
rect 4703 2269 4766 2334
rect 4865 2259 4949 2343
rect 5063 2259 5147 2343
rect 1937 2027 2023 2113
rect 2130 2030 2211 2111
rect -5285 1507 -5184 1608
rect 3538 1782 3625 1787
rect 3538 1705 3542 1782
rect 3542 1705 3619 1782
rect 3619 1705 3625 1782
rect 3538 1700 3625 1705
rect 3759 1693 3825 1759
rect 3928 1687 3997 1756
rect 5019 1701 5092 1775
rect 3587 1565 3643 1621
rect 4704 1623 4765 1684
rect 5016 1623 5091 1646
rect 5016 1577 5021 1623
rect 5021 1577 5091 1623
rect 5581 1634 5643 1636
rect 5581 1584 5643 1634
rect 5581 1574 5643 1584
rect 5023 1337 5077 1391
rect 3581 1128 3637 1184
rect 3784 1130 3838 1184
rect 5932 1333 5988 1389
rect 1462 870 1557 965
rect 3588 966 3649 1027
rect 4270 967 4329 1026
rect 3471 774 3474 796
rect 3474 774 3544 796
rect 3471 723 3544 774
rect 3900 754 3969 823
rect 5039 744 5102 822
rect 2971 589 3027 645
rect 3528 484 3582 538
rect 3928 611 3989 672
rect 4687 700 4758 708
rect 4687 637 4695 700
rect 4695 637 4758 700
rect 4687 629 4758 637
rect 4342 483 4398 539
rect 5471 600 5527 656
rect 5876 755 5932 811
rect 5278 443 5334 499
rect -4486 11 -4391 109
rect -4263 4 -4162 100
rect 3362 135 3432 205
rect 3160 -105 3216 -49
rect 3158 -291 3214 -235
rect 3568 -124 3624 -68
rect 4969 184 5025 237
rect 4969 181 5025 184
rect 4421 36 4482 97
rect 5094 42 5150 98
rect 3977 -116 4033 -60
rect 3161 -836 3215 -782
rect -6481 -1278 -6425 -1222
rect -6334 -1281 -6278 -1225
rect -6479 -1389 -6423 -1333
rect -6335 -1390 -6279 -1334
rect -5130 -1286 -5030 -1186
rect -4856 -1200 -4758 -1187
rect -4856 -1272 -4843 -1200
rect -4843 -1272 -4771 -1200
rect -4771 -1272 -4758 -1200
rect -4856 -1285 -4758 -1272
rect -5129 -1523 -5031 -1425
rect -4840 -1524 -4740 -1424
rect 3570 -688 3624 -634
rect 3973 -293 4034 -232
rect 3569 -843 3623 -789
rect 4672 -686 4728 -630
rect 3978 -813 4032 -759
rect 5095 -848 5149 -794
rect 4796 -984 4850 -930
rect 3161 -1238 3215 -1184
rect 4673 -1240 4727 -1186
rect 3868 -1390 3928 -1330
rect 3805 -1707 3873 -1690
rect 3805 -1756 3807 -1707
rect 3807 -1756 3873 -1707
rect 3805 -1758 3873 -1756
rect 3536 -1883 3592 -1827
rect 4058 -1901 4114 -1845
rect 5475 -1886 5531 -1830
rect -4396 -2733 -4258 -2595
rect -4395 -2994 -4259 -2858
rect -2482 -2966 -2399 -2886
rect -569 -3091 -484 -3006
rect -634 -3297 -568 -3231
rect 346 -3279 403 -3222
rect 2089 -2836 2145 -2780
rect 1757 -3120 1813 -3064
rect 1948 -3365 2005 -3354
rect 1948 -3411 2005 -3365
rect -2310 -3658 -2245 -3593
rect -2450 -3827 -2398 -3745
rect 647 -3605 703 -3549
rect -630 -4158 -563 -4091
rect 556 -3837 610 -3783
rect -2310 -4530 -2243 -4463
rect 146 -4154 203 -4097
rect -2450 -4684 -2398 -4602
rect -517 -4805 -458 -4746
rect 176 -4683 179 -4618
rect 179 -4683 241 -4618
rect -630 -5013 -570 -4953
rect 601 -4321 657 -4265
rect 1166 -3606 1224 -3548
rect 1054 -4047 1108 -3993
rect 988 -4329 1045 -4272
rect 962 -4835 1018 -4779
rect 1368 -3838 1425 -3781
rect 4244 -2126 4314 -2115
rect 4244 -2184 4256 -2126
rect 4256 -2184 4314 -2126
rect 4244 -2185 4314 -2184
rect 3875 -2523 3929 -2469
rect 4431 -2517 4485 -2463
rect 5122 -2518 5178 -2462
rect 3768 -2809 3834 -2801
rect 3768 -2860 3826 -2809
rect 3826 -2860 3834 -2809
rect 3768 -2868 3834 -2860
rect 5666 -2517 5720 -2463
rect 4046 -3145 4100 -3091
rect 4245 -3192 4313 -3184
rect 4245 -3249 4305 -3192
rect 4305 -3249 4313 -3192
rect 4245 -3257 4313 -3249
rect 5762 -3151 5816 -3097
rect 4045 -3424 4101 -3368
rect 3568 -3492 3576 -3440
rect 3576 -3492 3646 -3440
rect 3646 -3492 3654 -3440
rect 3568 -3500 3654 -3492
rect 4326 -3553 4380 -3499
rect 5078 -3441 5134 -3385
rect 4738 -3554 4794 -3498
rect 1367 -4053 1423 -3997
rect 1368 -4635 1422 -4581
rect 652 -5003 709 -4946
rect 1773 -4176 1830 -4119
rect 1777 -4851 1833 -4795
rect 1572 -5043 1626 -4989
rect -2310 -5380 -2243 -5313
rect 4122 -3868 4176 -3814
rect 3468 -4497 3545 -4489
rect 3468 -4543 3476 -4497
rect 3476 -4543 3537 -4497
rect 3537 -4543 3545 -4497
rect 4122 -4244 4178 -4188
rect 4530 -4003 4584 -3949
rect 4941 -3869 4997 -3813
rect 4938 -4223 4994 -4167
rect 5566 -3883 5574 -3816
rect 5574 -3883 5644 -3816
rect 5644 -3883 5652 -3816
rect 5566 -3891 5652 -3883
rect 5761 -4166 5817 -4162
rect 5761 -4216 5771 -4166
rect 5771 -4216 5817 -4166
rect 5761 -4218 5817 -4216
rect 4124 -4914 4180 -4858
rect 4324 -4917 4378 -4863
rect 5345 -4918 5399 -4864
rect 5568 -5208 5652 -5200
rect 5568 -5267 5576 -5208
rect 5576 -5267 5644 -5208
rect 5644 -5267 5652 -5208
rect -2450 -5574 -2398 -5492
rect -4998 -5920 -4893 -5815
rect -4807 -5922 -4700 -5815
rect -5150 -6406 -5089 -6345
rect -4986 -6408 -4923 -6345
rect -5138 -6604 -5070 -6536
rect -5014 -6605 -4944 -6535
rect 3716 -5616 3770 -5562
rect -2636 -5903 -2564 -5831
rect -2487 -5902 -2417 -5832
rect -749 -5881 -695 -5827
rect 3469 -5889 3531 -5882
rect 3469 -5944 3470 -5889
rect 3470 -5944 3530 -5889
rect 3530 -5944 3531 -5889
rect 4323 -5628 4379 -5572
rect 4734 -5630 4790 -5574
rect 4937 -5612 4991 -5558
rect 4531 -5877 4585 -5823
rect 4121 -6008 4177 -5952
rect -2310 -6253 -2243 -6186
rect 4938 -6007 4992 -5953
rect 4936 -6431 4992 -6375
rect 5576 -6352 5598 -6294
rect 5598 -6352 5645 -6294
rect 5576 -6363 5645 -6352
rect -3822 -7456 -3734 -7368
rect -3638 -7455 -3552 -7369
rect -3675 -8299 -3574 -8198
rect -2276 -8344 -2141 -8222
rect -2006 -8339 -1871 -8217
rect -1777 -8338 -1642 -8216
rect -2256 -11510 -2194 -11449
rect -3459 -12246 -3366 -12153
rect -3283 -12245 -3193 -12155
rect -3479 -12472 -3393 -12386
rect -3266 -12473 -3178 -12385
<< metal2 >>
rect -2453 6690 -1670 6731
rect -2453 6561 -2381 6690
rect -2252 6561 -2101 6690
rect -1972 6561 -1815 6690
rect -1686 6561 -1670 6690
rect -2453 6544 -1670 6561
rect 5875 6549 6167 6577
rect 5875 6468 5895 6549
rect 5976 6548 6167 6549
rect 5976 6469 6068 6548
rect 6147 6469 6167 6548
rect 5976 6468 6167 6469
rect 5875 6431 6167 6468
rect 5895 5830 5976 6431
rect 5880 5811 5996 5830
rect 5880 5730 5895 5811
rect 5976 5730 5996 5811
rect 5880 5724 5996 5730
rect -2315 4785 -1674 4808
rect -2315 4656 -2304 4785
rect -2175 4656 -2083 4785
rect -1954 4656 -1825 4785
rect -1696 4656 -1674 4785
rect -2315 4641 -1674 4656
rect 5895 3906 5976 5724
rect 5637 3896 5991 3906
rect -5666 3848 -5181 3881
rect -2892 3848 -2731 3849
rect -5666 3847 -5337 3848
rect -5666 3724 -5652 3847
rect -5529 3724 -5337 3847
rect -5666 3723 -5337 3724
rect -5207 3811 -2731 3848
rect -5207 3723 -2874 3811
rect -5666 3696 -5181 3723
rect -2892 3684 -2874 3723
rect -2747 3684 -2731 3811
rect 5637 3814 5731 3896
rect 5813 3814 5894 3896
rect 5976 3814 5991 3896
rect 5637 3805 5991 3814
rect -2892 3559 -2731 3684
rect -2892 3434 -2874 3559
rect -2749 3434 -2731 3559
rect -2892 3415 -2731 3434
rect 2749 2499 6330 2580
rect 1930 2113 2220 2150
rect 1930 2027 1937 2113
rect 2023 2111 2220 2113
rect 2749 2111 2830 2499
rect 4690 2343 5150 2359
rect 4690 2334 4865 2343
rect 3923 2319 4000 2330
rect 3923 2263 3933 2319
rect 3989 2263 4000 2319
rect 3923 2247 4000 2263
rect 4690 2269 4703 2334
rect 4766 2269 4865 2334
rect 4690 2259 4865 2269
rect 4949 2259 5063 2343
rect 5147 2259 5150 2343
rect 2023 2030 2130 2111
rect 2211 2030 2830 2111
rect 2023 2027 2220 2030
rect 1930 2000 2220 2027
rect 3524 1787 3636 1799
rect 3524 1700 3538 1787
rect 3625 1700 3636 1787
rect 3933 1771 3989 2247
rect 4690 2246 5150 2259
rect 3524 1688 3636 1700
rect 3746 1759 3837 1769
rect 3746 1693 3759 1759
rect 3825 1693 3837 1759
rect 3746 1686 3837 1693
rect 3916 1756 4009 1771
rect 3916 1687 3928 1756
rect 3997 1687 4009 1756
rect 4703 1700 4766 2246
rect 6045 1986 6170 1998
rect 5004 1881 6053 1986
rect 6158 1881 6170 1986
rect 5004 1816 5109 1881
rect 6045 1862 6170 1881
rect 5004 1775 5110 1816
rect 5004 1752 5019 1775
rect 5003 1701 5019 1752
rect 5092 1701 5110 1775
rect 3916 1675 4009 1687
rect 4683 1684 4786 1700
rect -5300 1609 -5160 1626
rect -5924 1608 -5160 1609
rect -5924 1507 -5285 1608
rect -5184 1507 -5160 1608
rect 3575 1621 3651 1625
rect 3575 1565 3587 1621
rect 3643 1565 3839 1621
rect 3575 1563 3651 1565
rect -5924 1506 -5160 1507
rect -6506 -1222 -6253 -1206
rect -6506 -1278 -6481 -1222
rect -6425 -1225 -6253 -1222
rect -6425 -1278 -6334 -1225
rect -6506 -1281 -6334 -1278
rect -6278 -1281 -6253 -1225
rect -6506 -1333 -6253 -1281
rect -6506 -1389 -6479 -1333
rect -6423 -1334 -6253 -1333
rect -6423 -1389 -6335 -1334
rect -6506 -1390 -6335 -1389
rect -6279 -1390 -6253 -1334
rect -6506 -1459 -6253 -1390
rect -5924 -7332 -5821 1506
rect -5300 1489 -5160 1506
rect -5622 1191 -4398 1318
rect -5622 -7060 -5495 1191
rect 3578 1184 3649 1189
rect 3783 1186 3839 1565
rect 3933 1555 3989 1675
rect 4683 1623 4704 1684
rect 4765 1623 4786 1684
rect 4683 1610 4786 1623
rect 5003 1646 5110 1701
rect 5003 1577 5016 1646
rect 5091 1577 5110 1646
rect 5003 1564 5110 1577
rect 5564 1636 5656 1644
rect 5564 1574 5581 1636
rect 5643 1574 5656 1636
rect 5564 1559 5656 1574
rect 3933 1499 4535 1555
rect 2088 1128 3581 1184
rect 3637 1128 3649 1184
rect 1455 965 1579 981
rect 1455 870 1462 965
rect 1557 957 1579 965
rect 1557 877 1960 957
rect 1557 870 1579 877
rect 1455 853 1579 870
rect -4508 133 -4134 136
rect -4509 109 -4133 133
rect -4509 11 -4486 109
rect -4391 100 -4133 109
rect -4391 11 -4263 100
rect -4509 4 -4263 11
rect -4162 4 -4133 100
rect -4509 -10 -4133 4
rect -4509 -11 -4391 -10
rect -4262 -11 -4133 -10
rect -5194 -1186 -4732 -1165
rect -5194 -1286 -5130 -1186
rect -5030 -1286 -4857 -1186
rect -4757 -1286 -4732 -1186
rect -5194 -1424 -4732 -1286
rect -5194 -1524 -5130 -1424
rect -5030 -1524 -4840 -1424
rect -4740 -1524 -4732 -1424
rect -5194 -1556 -4732 -1524
rect 1880 -2080 1960 877
rect 2088 -864 2144 1128
rect 3578 1116 3649 1128
rect 3772 1184 3850 1186
rect 3772 1130 3784 1184
rect 3838 1130 3850 1184
rect 3772 1118 3850 1130
rect 3576 1027 3651 1044
rect 4259 1027 4337 1036
rect 3576 966 3588 1027
rect 3649 1026 4337 1027
rect 3649 967 4270 1026
rect 4329 967 4337 1026
rect 3649 966 4337 967
rect 3576 958 3719 966
rect 3458 796 3554 805
rect 3458 723 3471 796
rect 3544 723 3554 796
rect 3458 711 3554 723
rect 3658 672 3719 958
rect 4259 956 4337 966
rect 4479 878 4535 1499
rect 5013 1391 5093 1403
rect 5013 1337 5023 1391
rect 5077 1389 5093 1391
rect 5923 1389 6003 1398
rect 5077 1337 5932 1389
rect 5013 1333 5932 1337
rect 5988 1333 6003 1389
rect 5013 1326 5093 1333
rect 5923 1325 6003 1333
rect 3884 823 3982 835
rect 3884 754 3900 823
rect 3969 754 3982 823
rect 3884 743 3982 754
rect 4479 822 4963 878
rect 3925 672 3999 684
rect 2230 646 2318 662
rect 2962 646 3038 659
rect 2230 582 2244 646
rect 2308 645 3038 646
rect 2308 589 2971 645
rect 3027 589 3038 645
rect 3658 611 3928 672
rect 3989 611 3999 672
rect 3925 598 3999 611
rect 2308 582 3038 589
rect 2230 566 2318 582
rect 2962 574 3038 582
rect 3512 539 3588 552
rect 4332 539 4408 548
rect 4479 539 4535 822
rect 4907 811 4963 822
rect 5036 822 5107 835
rect 5036 811 5039 822
rect 4907 755 5039 811
rect 5036 744 5039 755
rect 5102 811 5107 822
rect 5873 811 5941 824
rect 5102 755 5876 811
rect 5932 755 5941 811
rect 5102 744 5107 755
rect 5036 732 5107 744
rect 5873 742 5941 755
rect 4675 708 4772 717
rect 4675 629 4686 708
rect 4759 629 4772 708
rect 4675 619 4772 629
rect 5461 656 5540 666
rect 5461 600 5471 656
rect 5527 600 5540 656
rect 5461 592 5540 600
rect 3512 538 4342 539
rect 2445 494 2553 495
rect 2445 471 2556 494
rect 3512 484 3528 538
rect 3582 484 4342 538
rect 3512 483 4342 484
rect 4398 483 4535 539
rect 5265 499 5345 508
rect 3512 476 3588 483
rect 4332 472 4408 483
rect 2445 401 2462 471
rect 2532 401 2556 471
rect 2445 391 2556 401
rect 5265 443 5278 499
rect 5334 443 5345 499
rect 5265 441 5345 443
rect 5265 394 5334 441
rect 2445 326 2554 391
rect 2445 257 2465 326
rect 2534 257 2554 326
rect 2445 168 2554 257
rect 2445 99 2465 168
rect 2534 99 2554 168
rect 2445 88 2554 99
rect 2715 338 5334 394
rect 2445 77 2553 88
rect 2208 -732 2293 -717
rect 2208 -802 2213 -732
rect 2283 -733 2293 -732
rect 2465 -733 2534 77
rect 2715 -401 2771 338
rect 4958 237 5034 250
rect 3350 205 3444 217
rect 3350 135 3362 205
rect 3432 135 3444 205
rect 3350 122 3444 135
rect 4795 181 4969 237
rect 5025 181 5034 237
rect 4417 97 4492 118
rect 4216 36 4421 97
rect 4482 36 4492 97
rect 3147 -49 3228 -36
rect 3147 -105 3160 -49
rect 3216 -105 3228 -49
rect 3553 -62 3637 -56
rect 3966 -60 4045 -50
rect 3553 -68 3905 -62
rect 3553 -71 3568 -68
rect 3147 -117 3228 -105
rect 3308 -124 3568 -71
rect 3624 -123 3905 -68
rect 3624 -124 3637 -123
rect 3308 -127 3637 -124
rect 3154 -235 3220 -223
rect 3308 -235 3364 -127
rect 3553 -136 3637 -127
rect 3149 -291 3158 -235
rect 3214 -291 3364 -235
rect 3844 -232 3905 -123
rect 3966 -116 3977 -60
rect 4033 -116 4045 -60
rect 3966 -130 4045 -116
rect 3962 -232 4061 -220
rect 4216 -232 4277 36
rect 4417 22 4492 36
rect 3154 -303 3220 -291
rect 3844 -293 3973 -232
rect 4034 -293 4277 -232
rect 3962 -301 4061 -293
rect 2600 -417 2771 -401
rect 2600 -473 2603 -417
rect 2659 -473 2771 -417
rect 2600 -486 2669 -473
rect 3558 -633 3633 -624
rect 4660 -630 4735 -618
rect 3558 -634 4035 -633
rect 3558 -688 3570 -634
rect 3624 -688 4035 -634
rect 3558 -689 4035 -688
rect 4660 -686 4672 -630
rect 4728 -686 4735 -630
rect 4660 -689 4735 -686
rect 3558 -700 3633 -689
rect 2283 -802 2534 -733
rect 3979 -747 4035 -689
rect 3966 -758 4044 -747
rect 3150 -781 3229 -770
rect 2208 -803 2352 -802
rect 2208 -813 2293 -803
rect 3150 -837 3160 -781
rect 3216 -837 3229 -781
rect 3150 -848 3229 -837
rect 3556 -788 3636 -777
rect 3556 -844 3568 -788
rect 3624 -844 3636 -788
rect 3966 -814 3977 -758
rect 4033 -814 4044 -758
rect 3966 -824 4044 -814
rect 3556 -855 3636 -844
rect 2074 -882 2174 -864
rect 2074 -938 2096 -882
rect 2152 -938 2174 -882
rect 2074 -954 2174 -938
rect 3149 -1184 3227 -1172
rect 4672 -1174 4728 -689
rect 4795 -928 4851 181
rect 4958 172 5034 181
rect 5082 98 5164 108
rect 5082 42 5094 98
rect 5150 42 5164 98
rect 5082 34 5164 42
rect 5094 -76 5150 34
rect 5471 -76 5527 592
rect 5094 -132 5527 -76
rect 5094 -787 5150 -132
rect 5080 -794 5164 -787
rect 5080 -848 5095 -794
rect 5149 -848 5164 -794
rect 5080 -855 5164 -848
rect 4784 -930 4863 -928
rect 4784 -984 4796 -930
rect 4784 -995 4801 -984
rect 4866 -995 4879 -930
rect 3149 -1238 3161 -1184
rect 3215 -1238 3227 -1184
rect 3149 -1250 3227 -1238
rect 4661 -1175 4738 -1174
rect 4661 -1186 4739 -1175
rect 4661 -1240 4673 -1186
rect 4727 -1240 4739 -1186
rect 3160 -1341 3216 -1250
rect 4661 -1252 4739 -1240
rect 640 -2160 1960 -2080
rect 2600 -1397 3216 -1341
rect 3853 -1330 3943 -1319
rect 3853 -1390 3866 -1330
rect 3928 -1390 3943 -1330
rect -4412 -2595 -4232 -2562
rect -4412 -2733 -4396 -2595
rect -4258 -2733 -4232 -2595
rect -4412 -2857 -4232 -2733
rect -4412 -2995 -4396 -2857
rect -4258 -2995 -4232 -2857
rect -2492 -2886 -2386 -2874
rect -2492 -2966 -2482 -2886
rect -2399 -2966 -2386 -2886
rect -2492 -2979 -2386 -2966
rect -4412 -3023 -4232 -2995
rect -3133 -3058 -2988 -3052
rect -3133 -3127 -3091 -3058
rect -3022 -3127 -2988 -3058
rect -3133 -3227 -2988 -3127
rect -3133 -3296 -3091 -3227
rect -3022 -3296 -2988 -3227
rect -3133 -3460 -2988 -3296
rect -3133 -3529 -3091 -3460
rect -3022 -3529 -2988 -3460
rect -3133 -3551 -2988 -3529
rect -3120 -3556 -2999 -3551
rect -3091 -4077 -3022 -3556
rect -2480 -3736 -2398 -2979
rect -576 -3005 -473 -2992
rect -643 -3092 -570 -3005
rect -483 -3092 -473 -3005
rect -576 -3106 -473 -3092
rect -644 -3230 -557 -3221
rect -644 -3298 -635 -3230
rect -567 -3298 -557 -3230
rect 332 -3222 415 -3213
rect 332 -3279 346 -3222
rect 403 -3279 415 -3222
rect 332 -3284 415 -3279
rect -644 -3308 -557 -3298
rect 346 -3308 415 -3284
rect 346 -3365 483 -3308
rect -2323 -3593 -2234 -3581
rect -2323 -3658 -2310 -3593
rect -2245 -3658 -2234 -3593
rect -2323 -3666 -2234 -3658
rect -2489 -3745 -2383 -3736
rect -2489 -3827 -2450 -3745
rect -2398 -3827 -2383 -3745
rect -2489 -3841 -2383 -3827
rect -3117 -4106 -2996 -4077
rect -3117 -4175 -3091 -4106
rect -3022 -4175 -2996 -4106
rect -3117 -4205 -2996 -4175
rect -2480 -4591 -2398 -3841
rect -2310 -4459 -2243 -3666
rect 426 -3781 483 -3365
rect 640 -3530 720 -2160
rect 2600 -2365 2656 -1397
rect 3853 -1411 3943 -1390
rect 4683 -1415 4739 -1252
rect 4058 -1471 4739 -1415
rect 3798 -1690 3888 -1678
rect 3706 -1758 3805 -1690
rect 3873 -1758 3888 -1690
rect 3706 -1770 3888 -1758
rect 3524 -1827 3600 -1815
rect 3524 -1883 3536 -1827
rect 3592 -1883 3601 -1827
rect 3524 -1895 3600 -1883
rect 1757 -2421 2656 -2365
rect 1757 -3050 1813 -2421
rect 2079 -2780 2155 -2752
rect 2079 -2836 2089 -2780
rect 2145 -2836 2155 -2780
rect 2079 -2849 2155 -2836
rect 3706 -2789 3774 -1770
rect 4058 -1836 4114 -1471
rect 5463 -1830 5543 -1821
rect 4044 -1845 4127 -1836
rect 4044 -1901 4058 -1845
rect 4114 -1901 4127 -1845
rect 5463 -1886 5475 -1830
rect 5531 -1886 5543 -1830
rect 5463 -1896 5543 -1886
rect 4044 -1906 4127 -1901
rect 3862 -2468 3933 -2456
rect 4058 -2468 4114 -1906
rect 4231 -2115 4325 -2106
rect 4231 -2185 4244 -2115
rect 4314 -2185 4325 -2115
rect 4231 -2194 4325 -2185
rect 3862 -2469 4114 -2468
rect 3862 -2523 3875 -2469
rect 3929 -2523 4114 -2469
rect 3862 -2524 4114 -2523
rect 3862 -2536 3933 -2524
rect 3706 -2801 3846 -2789
rect 3706 -2868 3768 -2801
rect 3834 -2868 3846 -2801
rect 3706 -2880 3846 -2868
rect 1748 -3064 1824 -3050
rect 1748 -3120 1757 -3064
rect 1813 -3120 1824 -3064
rect 1748 -3132 1824 -3120
rect 1927 -3354 2023 -3344
rect 1927 -3411 1948 -3354
rect 2005 -3411 2023 -3354
rect 3766 -3405 3828 -2880
rect 4031 -3091 4117 -3089
rect 4031 -3145 4046 -3091
rect 4100 -3145 4117 -3091
rect 4031 -3160 4117 -3145
rect 4244 -3110 4314 -2194
rect 4419 -2462 4488 -2451
rect 5116 -2462 5187 -2450
rect 4419 -2463 5122 -2462
rect 4419 -2517 4431 -2463
rect 4485 -2517 5122 -2463
rect 4419 -2518 5122 -2517
rect 5178 -2518 5187 -2462
rect 5475 -2462 5531 -1896
rect 5663 -2462 5731 -2450
rect 5475 -2463 5731 -2462
rect 5475 -2517 5666 -2463
rect 5720 -2517 5731 -2463
rect 5475 -2518 5731 -2517
rect 4419 -2529 4488 -2518
rect 5116 -2527 5187 -2518
rect 5663 -2529 5731 -2518
rect 5751 -3097 5827 -3088
rect 4045 -3358 4101 -3160
rect 4244 -3180 5649 -3110
rect 5751 -3151 5762 -3097
rect 5816 -3151 5827 -3097
rect 5751 -3165 5827 -3151
rect 4232 -3184 4326 -3180
rect 4232 -3257 4245 -3184
rect 4313 -3257 4326 -3184
rect 4232 -3269 4326 -3257
rect 1927 -3434 2023 -3411
rect 640 -3548 730 -3530
rect 1160 -3548 1233 -3535
rect 640 -3549 1166 -3548
rect 640 -3605 647 -3549
rect 703 -3605 1166 -3549
rect 640 -3606 1166 -3605
rect 1224 -3606 1233 -3548
rect 640 -3620 730 -3606
rect 1160 -3619 1233 -3606
rect 544 -3781 616 -3771
rect 1365 -3781 1433 -3768
rect 1534 -3781 1591 -3780
rect 257 -3783 1368 -3781
rect 257 -3837 556 -3783
rect 610 -3837 1368 -3783
rect 257 -3838 1368 -3837
rect 1425 -3838 1722 -3781
rect -1554 -3944 -1545 -3879
rect -1480 -3944 -1471 -3879
rect 257 -4015 314 -3838
rect 146 -4072 314 -4015
rect -647 -4090 -547 -4078
rect 146 -4090 215 -4072
rect -647 -4159 -631 -4090
rect -562 -4159 -547 -4090
rect -647 -4171 -547 -4159
rect 133 -4097 215 -4090
rect 133 -4154 146 -4097
rect 203 -4154 215 -4097
rect 133 -4165 215 -4154
rect -2322 -4463 -2233 -4459
rect -2322 -4530 -2310 -4463
rect -2243 -4530 -2233 -4463
rect -2322 -4544 -2233 -4530
rect -2506 -4602 -2391 -4591
rect -2506 -4684 -2450 -4602
rect -2398 -4684 -2391 -4602
rect -2506 -4698 -2391 -4684
rect -2480 -5486 -2398 -4698
rect -2310 -5307 -2243 -4544
rect 165 -4618 250 -4599
rect 165 -4683 176 -4618
rect 241 -4683 250 -4618
rect 165 -4699 250 -4683
rect -522 -4745 -447 -4733
rect -522 -4806 -518 -4745
rect -457 -4806 -447 -4745
rect -522 -4820 -447 -4806
rect -1844 -5022 -1725 -5019
rect -2002 -5039 -1725 -5022
rect -2002 -5124 -1986 -5039
rect -1896 -5043 -1725 -5039
rect -1896 -5124 -1826 -5043
rect -2002 -5129 -1826 -5124
rect -1740 -5044 -1725 -5043
rect -1446 -5044 -1363 -4938
rect -641 -4952 -549 -4940
rect -641 -5014 -631 -4952
rect -569 -5014 -549 -4952
rect 426 -4946 483 -3838
rect 544 -3850 616 -3838
rect 1365 -3850 1433 -3838
rect 1049 -3993 1119 -3980
rect 1049 -3997 1054 -3993
rect 671 -4047 1054 -3997
rect 1108 -3997 1119 -3993
rect 1365 -3997 1432 -3984
rect 1108 -4047 1367 -3997
rect 671 -4053 1367 -4047
rect 1423 -4053 1432 -3997
rect 671 -4253 727 -4053
rect 1049 -4059 1119 -4053
rect 1365 -4067 1432 -4053
rect 592 -4265 727 -4253
rect 592 -4321 601 -4265
rect 657 -4321 727 -4265
rect 980 -4272 1049 -4258
rect 1534 -4272 1591 -3838
rect 1665 -3968 1722 -3838
rect 1665 -4025 1830 -3968
rect 1773 -4112 1830 -4025
rect 1760 -4119 1842 -4112
rect 1760 -4176 1773 -4119
rect 1830 -4176 1842 -4119
rect 1760 -4183 1842 -4176
rect 1773 -4185 1830 -4183
rect 592 -4333 671 -4321
rect 979 -4329 988 -4272
rect 1045 -4329 1591 -4272
rect 980 -4345 1049 -4329
rect 1356 -4580 1427 -4569
rect 962 -4581 1833 -4580
rect 962 -4635 1368 -4581
rect 1422 -4635 1833 -4581
rect 962 -4636 1833 -4635
rect 962 -4774 1018 -4636
rect 1356 -4647 1427 -4636
rect 950 -4779 1030 -4774
rect 950 -4835 962 -4779
rect 1018 -4835 1030 -4779
rect 1777 -4792 1833 -4636
rect 950 -4845 1030 -4835
rect 1764 -4795 1846 -4792
rect 1764 -4851 1777 -4795
rect 1833 -4851 1846 -4795
rect 1764 -4860 1846 -4851
rect 647 -4946 716 -4934
rect 426 -5003 652 -4946
rect 709 -5003 718 -4946
rect 1569 -4983 1638 -4977
rect 1569 -4987 1653 -4983
rect 1948 -4987 2005 -3434
rect 3580 -3438 3828 -3405
rect 4029 -3368 4115 -3358
rect 4029 -3424 4045 -3368
rect 4101 -3424 4115 -3368
rect 4029 -3429 4115 -3424
rect 5064 -3385 5147 -3376
rect 4045 -3433 4101 -3429
rect 3554 -3440 3828 -3438
rect 3554 -3500 3568 -3440
rect 3654 -3467 3828 -3440
rect 5064 -3441 5078 -3385
rect 5134 -3441 5147 -3385
rect 5064 -3443 5147 -3441
rect 3654 -3500 3668 -3467
rect 4334 -3486 4390 -3485
rect 3554 -3512 3668 -3500
rect 4314 -3498 4401 -3486
rect 4730 -3498 4804 -3486
rect 4940 -3498 5014 -3482
rect 4314 -3499 4738 -3498
rect 3580 -4476 3642 -3512
rect 4314 -3553 4326 -3499
rect 4380 -3553 4738 -3499
rect 4314 -3554 4738 -3553
rect 4794 -3554 4948 -3498
rect 5004 -3554 5014 -3498
rect 4314 -3558 4401 -3554
rect 4314 -3563 4392 -3558
rect 4730 -3567 4804 -3554
rect 4940 -3568 5014 -3554
rect 4110 -3813 4187 -3805
rect 4928 -3813 5009 -3804
rect 4110 -3814 4941 -3813
rect 4110 -3868 4122 -3814
rect 4176 -3868 4941 -3814
rect 4110 -3869 4941 -3868
rect 4997 -3869 5009 -3813
rect 4110 -3880 4187 -3869
rect 4529 -3940 4585 -3869
rect 4928 -3878 5009 -3869
rect 4517 -3949 4599 -3940
rect 4517 -4003 4530 -3949
rect 4584 -4003 4599 -3949
rect 4517 -4007 4599 -4003
rect 5078 -4157 5134 -3443
rect 5579 -3806 5649 -3180
rect 5557 -3816 5662 -3806
rect 5557 -3891 5566 -3816
rect 5652 -3891 5662 -3816
rect 5557 -3903 5662 -3891
rect 4925 -4167 5134 -4157
rect 4113 -4188 4187 -4176
rect 4113 -4244 4122 -4188
rect 4178 -4244 4293 -4188
rect 4925 -4223 4938 -4167
rect 4994 -4213 5134 -4167
rect 4994 -4223 5006 -4213
rect 4925 -4227 5006 -4223
rect 4113 -4255 4293 -4244
rect 4237 -4397 4293 -4255
rect 4933 -4397 4989 -4227
rect 4237 -4453 5263 -4397
rect 3456 -4489 3642 -4476
rect 3456 -4543 3468 -4489
rect 3545 -4543 3642 -4489
rect 3456 -4548 3642 -4543
rect 1569 -4989 2005 -4987
rect 647 -5013 716 -5003
rect -641 -5025 -549 -5014
rect -1740 -5127 -1363 -5044
rect 1569 -5043 1572 -4989
rect 1626 -4996 2005 -4989
rect 1569 -5055 1580 -5043
rect 1573 -5060 1580 -5055
rect 1644 -5044 2005 -4996
rect 1644 -5060 1653 -5044
rect 1573 -5071 1653 -5060
rect -1740 -5129 -1725 -5127
rect -2002 -5135 -1725 -5129
rect -1844 -5141 -1725 -5135
rect -2326 -5313 -2231 -5307
rect -2326 -5380 -2310 -5313
rect -2243 -5380 -2231 -5313
rect -2326 -5391 -2231 -5380
rect -558 -5332 -477 -5322
rect 3349 -5332 3426 -5323
rect -2493 -5492 -2386 -5486
rect -2493 -5574 -2450 -5492
rect -2398 -5574 -2386 -5492
rect -2493 -5593 -2386 -5574
rect -5020 -5815 -4689 -5791
rect -5020 -5920 -4998 -5815
rect -4893 -5920 -4807 -5815
rect -5020 -5922 -4807 -5920
rect -4700 -5831 -2404 -5815
rect -4700 -5903 -2636 -5831
rect -2564 -5832 -2404 -5831
rect -2564 -5902 -2487 -5832
rect -2417 -5902 -2404 -5832
rect -2564 -5903 -2404 -5902
rect -4700 -5922 -2404 -5903
rect -5020 -5933 -4689 -5922
rect -2310 -6180 -2243 -5391
rect -558 -5392 -548 -5332
rect -488 -5392 3355 -5332
rect 3415 -5392 3426 -5332
rect -558 -5402 -477 -5392
rect 3349 -5402 3426 -5392
rect 3357 -5471 3436 -5459
rect -638 -5536 3361 -5471
rect 3426 -5536 3436 -5471
rect -638 -5600 -573 -5536
rect 3357 -5548 3436 -5536
rect -645 -5606 -573 -5600
rect -888 -5671 -573 -5606
rect 585 -5606 667 -5596
rect 585 -5671 595 -5606
rect 660 -5612 908 -5606
rect 660 -5671 961 -5612
rect 2250 -5671 2503 -5606
rect 2568 -5671 2577 -5606
rect 585 -5682 667 -5671
rect 897 -5681 961 -5671
rect 887 -5682 971 -5681
rect -809 -5826 -682 -5814
rect -809 -5882 -750 -5826
rect -694 -5882 -682 -5826
rect -809 -5893 -682 -5882
rect 564 -5885 573 -5818
rect 640 -5885 748 -5818
rect 2349 -5872 2421 -5823
rect 3580 -5872 3642 -4548
rect 4120 -4858 4193 -4854
rect 4013 -4914 4124 -4858
rect 4180 -4914 4193 -4858
rect 4013 -4919 4193 -4914
rect 4311 -4863 4391 -4855
rect 4311 -4917 4324 -4863
rect 4378 -4917 4391 -4863
rect 3706 -5561 3781 -5553
rect 4013 -5561 4069 -4919
rect 4311 -4920 4391 -4917
rect 5207 -4865 5263 -4453
rect 5333 -4864 5412 -4849
rect 5333 -4865 5345 -4864
rect 5207 -4918 5345 -4865
rect 5399 -4918 5412 -4864
rect 3706 -5562 4069 -5561
rect 3706 -5616 3716 -5562
rect 3770 -5616 4069 -5562
rect 4323 -5569 4379 -4920
rect 5207 -4921 5412 -4918
rect 5333 -4929 5412 -4921
rect 5576 -5185 5645 -3903
rect 5761 -4153 5817 -3165
rect 6249 -3498 6330 2499
rect 6249 -3554 6262 -3498
rect 6318 -3554 6330 -3498
rect 6249 -3602 6330 -3554
rect 6249 -3630 6262 -3602
rect 6250 -3658 6262 -3630
rect 6318 -3658 6330 -3602
rect 6250 -3670 6330 -3658
rect 5754 -4162 5825 -4153
rect 5752 -4218 5761 -4162
rect 5817 -4218 5826 -4162
rect 5754 -4228 5825 -4218
rect 5559 -5200 5662 -5185
rect 5559 -5267 5568 -5200
rect 5652 -5267 5662 -5200
rect 5559 -5279 5662 -5267
rect 4924 -5558 5113 -5555
rect 3706 -5617 4069 -5616
rect 4310 -5572 4388 -5569
rect 3706 -5626 3781 -5617
rect 4310 -5628 4323 -5572
rect 4379 -5574 4388 -5572
rect 4728 -5574 4800 -5563
rect 4379 -5628 4734 -5574
rect 4310 -5630 4734 -5628
rect 4790 -5630 4800 -5574
rect 4924 -5612 4937 -5558
rect 4991 -5612 5113 -5558
rect 4924 -5617 5112 -5612
rect 4310 -5637 4388 -5630
rect 4728 -5641 4800 -5630
rect 2349 -5882 3642 -5872
rect 2349 -5944 3469 -5882
rect 3531 -5944 3642 -5882
rect 4519 -5823 4597 -5818
rect 4519 -5877 4531 -5823
rect 4585 -5877 4597 -5823
rect 4519 -5885 4597 -5877
rect 3457 -5949 3539 -5944
rect 4109 -5952 4189 -5943
rect 4530 -5952 4586 -5885
rect 4926 -5952 4996 -5941
rect 4109 -6008 4121 -5952
rect 4177 -5953 4996 -5952
rect 4177 -6007 4938 -5953
rect 4992 -6007 4996 -5953
rect 4177 -6008 4996 -6007
rect 4109 -6018 4189 -6008
rect 4926 -6019 4996 -6008
rect -2323 -6186 -2232 -6180
rect -2323 -6253 -2310 -6186
rect -2243 -6253 -2232 -6186
rect -2323 -6264 -2232 -6253
rect -5152 -6345 -4899 -6323
rect -526 -6345 -463 -6067
rect -5152 -6406 -5150 -6345
rect -5089 -6406 -4986 -6345
rect -5152 -6408 -4986 -6406
rect -4923 -6408 -463 -6345
rect -5152 -6425 -4899 -6408
rect -5152 -6535 -4929 -6511
rect 1085 -6535 1143 -6025
rect 5056 -6366 5112 -5617
rect 5576 -6263 5645 -5279
rect 5573 -6273 5666 -6263
rect 5573 -6277 5589 -6273
rect 4922 -6375 5112 -6366
rect 4922 -6431 4936 -6375
rect 4992 -6431 5112 -6375
rect 5561 -6294 5589 -6277
rect 5654 -6277 5666 -6273
rect 5561 -6363 5576 -6294
rect 5654 -6338 5676 -6277
rect 5645 -6363 5676 -6338
rect 5561 -6381 5676 -6363
rect 4922 -6441 5112 -6431
rect -5152 -6536 -5014 -6535
rect -5152 -6604 -5138 -6536
rect -5070 -6604 -5014 -6536
rect -5152 -6605 -5014 -6604
rect -4944 -6605 1149 -6535
rect -5152 -6626 -4929 -6605
rect -3751 -6861 -2398 -6845
rect -3751 -6925 -2397 -6861
rect -3751 -7060 -3624 -6925
rect -5622 -7187 -3624 -7060
rect -2469 -7200 -2397 -6925
rect -2562 -7256 -2397 -7200
rect -2469 -7257 -2399 -7256
rect -5924 -7333 -3555 -7332
rect -5924 -7368 -3532 -7333
rect -5924 -7435 -3822 -7368
rect -3839 -7456 -3822 -7435
rect -3734 -7369 -3532 -7368
rect -3734 -7455 -3638 -7369
rect -3552 -7455 -3532 -7369
rect -3734 -7456 -3532 -7455
rect -3839 -7472 -3532 -7456
rect -3690 -8198 -3330 -8178
rect -3690 -8299 -3675 -8198
rect -3574 -8299 -3437 -8198
rect -3336 -8299 -3330 -8198
rect -3690 -8329 -3330 -8299
rect -2327 -8216 -1628 -8190
rect -2327 -8217 -1777 -8216
rect -2327 -8222 -2006 -8217
rect -2327 -8344 -2276 -8222
rect -2141 -8339 -2006 -8222
rect -1871 -8338 -1777 -8217
rect -1642 -8338 -1628 -8216
rect -1871 -8339 -1628 -8338
rect -2141 -8344 -1628 -8339
rect -2327 -8367 -1628 -8344
rect -2269 -11449 -2178 -11434
rect -2269 -11483 -2256 -11449
rect -2270 -11510 -2256 -11483
rect -2194 -11510 -2178 -11449
rect -2270 -11524 -2178 -11510
rect -3469 -12153 -3160 -12130
rect -3469 -12246 -3459 -12153
rect -3366 -12155 -3160 -12153
rect -2270 -12155 -2180 -11524
rect -3366 -12245 -3283 -12155
rect -3193 -12245 -2180 -12155
rect -1255 -11752 -1167 -11736
rect -1255 -11808 -1037 -11752
rect -3366 -12246 -3160 -12245
rect -3469 -12274 -3160 -12246
rect -3490 -12385 -3139 -12343
rect -1255 -12385 -1167 -11808
rect -3490 -12386 -3266 -12385
rect -3490 -12472 -3479 -12386
rect -3393 -12472 -3266 -12386
rect -3490 -12473 -3266 -12472
rect -3178 -12473 -1167 -12385
rect -3490 -12515 -3139 -12473
<< via2 >>
rect -2381 6561 -2252 6690
rect -2101 6561 -1972 6690
rect -1815 6561 -1686 6690
rect -2304 4656 -2175 4785
rect -2083 4656 -1954 4785
rect -1825 4656 -1696 4785
rect 3538 1700 3625 1787
rect 3759 1693 3825 1759
rect 6053 1881 6158 1986
rect -6481 -1278 -6425 -1222
rect -6334 -1281 -6278 -1225
rect -6479 -1389 -6423 -1333
rect -6335 -1390 -6279 -1334
rect 5581 1574 5643 1636
rect -4486 11 -4391 109
rect -4263 4 -4162 100
rect -5130 -1286 -5030 -1186
rect -4857 -1187 -4757 -1186
rect -4857 -1285 -4856 -1187
rect -4856 -1285 -4758 -1187
rect -4758 -1285 -4757 -1187
rect -4857 -1286 -4757 -1285
rect -5130 -1425 -5030 -1424
rect -5130 -1523 -5129 -1425
rect -5129 -1523 -5031 -1425
rect -5031 -1523 -5030 -1425
rect -5130 -1524 -5030 -1523
rect -4840 -1524 -4740 -1424
rect 3471 723 3544 796
rect 3900 754 3969 823
rect 2244 582 2308 646
rect 2971 589 3027 645
rect 4686 629 4687 708
rect 4687 629 4758 708
rect 4758 629 4759 708
rect 2462 401 2532 471
rect 2465 257 2534 326
rect 2465 99 2534 168
rect 2213 -802 2283 -732
rect 3362 135 3432 205
rect 3160 -105 3216 -49
rect 3568 -124 3624 -68
rect 3977 -116 4033 -60
rect 2603 -473 2659 -417
rect 3160 -782 3216 -781
rect 3160 -836 3161 -782
rect 3161 -836 3215 -782
rect 3215 -836 3216 -782
rect 3160 -837 3216 -836
rect 3568 -789 3624 -788
rect 3568 -843 3569 -789
rect 3569 -843 3623 -789
rect 3623 -843 3624 -789
rect 3568 -844 3624 -843
rect 3977 -759 4033 -758
rect 3977 -813 3978 -759
rect 3978 -813 4032 -759
rect 4032 -813 4033 -759
rect 3977 -814 4033 -813
rect 2096 -938 2152 -882
rect 4801 -984 4850 -930
rect 4850 -984 4866 -930
rect 4801 -995 4866 -984
rect 3866 -1390 3868 -1330
rect 3868 -1390 3928 -1330
rect -4396 -2733 -4258 -2595
rect -4396 -2858 -4258 -2857
rect -4396 -2994 -4395 -2858
rect -4395 -2994 -4259 -2858
rect -4259 -2994 -4258 -2858
rect -4396 -2995 -4258 -2994
rect -3091 -3127 -3022 -3058
rect -3091 -3296 -3022 -3227
rect -3091 -3529 -3022 -3460
rect -570 -3006 -483 -3005
rect -570 -3091 -569 -3006
rect -569 -3091 -484 -3006
rect -484 -3091 -483 -3006
rect -570 -3092 -483 -3091
rect -635 -3231 -567 -3230
rect -635 -3297 -634 -3231
rect -634 -3297 -568 -3231
rect -568 -3297 -567 -3231
rect -635 -3298 -567 -3297
rect -3091 -4175 -3022 -4106
rect 3536 -1883 3592 -1827
rect 2089 -2836 2145 -2780
rect -1545 -3944 -1480 -3879
rect -631 -4091 -562 -4090
rect -631 -4158 -630 -4091
rect -630 -4158 -563 -4091
rect -563 -4158 -562 -4091
rect -631 -4159 -562 -4158
rect 176 -4683 241 -4618
rect -518 -4746 -457 -4745
rect -518 -4805 -517 -4746
rect -517 -4805 -458 -4746
rect -458 -4805 -457 -4746
rect -518 -4806 -457 -4805
rect -1986 -5124 -1896 -5039
rect -1826 -5129 -1740 -5043
rect -631 -4953 -569 -4952
rect -631 -5013 -630 -4953
rect -630 -5013 -570 -4953
rect -570 -5013 -569 -4953
rect -631 -5014 -569 -5013
rect 4948 -3554 5004 -3498
rect 1580 -5043 1626 -4996
rect 1626 -5043 1644 -4996
rect 1580 -5060 1644 -5043
rect -548 -5392 -488 -5332
rect 3355 -5392 3415 -5332
rect 3361 -5536 3426 -5471
rect 595 -5671 660 -5606
rect 2503 -5671 2568 -5606
rect -750 -5827 -694 -5826
rect -750 -5881 -749 -5827
rect -749 -5881 -695 -5827
rect -695 -5881 -694 -5827
rect -750 -5882 -694 -5881
rect 573 -5885 640 -5818
rect 6262 -3554 6318 -3498
rect 6262 -3658 6318 -3602
rect 5589 -6294 5654 -6273
rect 5589 -6338 5645 -6294
rect 5645 -6338 5654 -6294
rect -3675 -8299 -3574 -8198
rect -3437 -8299 -3336 -8198
rect -2276 -8344 -2141 -8222
rect -2006 -8339 -1871 -8217
rect -1777 -8338 -1642 -8216
<< metal3 >>
rect -2453 6690 -1670 6731
rect -4391 6561 -2381 6690
rect -2252 6561 -2101 6690
rect -1972 6561 -1815 6690
rect -1686 6561 -1670 6690
rect -4391 4785 -4262 6561
rect -2453 6544 -1670 6561
rect -2315 4785 -1674 4808
rect -4391 4656 -2304 4785
rect -2175 4656 -2083 4785
rect -1954 4656 -1825 4785
rect -1696 4656 -1674 4785
rect -4391 136 -4262 4656
rect -2315 4641 -1674 4656
rect -3756 2769 5658 2861
rect -4508 133 -4134 136
rect -4509 109 -4133 133
rect -4509 11 -4486 109
rect -4391 100 -4133 109
rect -4391 11 -4263 100
rect -4509 4 -4263 11
rect -4162 4 -4133 100
rect -4509 -11 -4133 4
rect -5194 -1186 -4732 -1165
rect -5194 -1206 -5130 -1186
rect -6506 -1222 -5130 -1206
rect -6506 -1278 -6481 -1222
rect -6425 -1225 -5130 -1222
rect -6425 -1278 -6334 -1225
rect -6506 -1281 -6334 -1278
rect -6278 -1281 -5130 -1225
rect -6506 -1286 -5130 -1281
rect -5030 -1286 -4857 -1186
rect -4757 -1286 -4732 -1186
rect -6506 -1333 -4732 -1286
rect -6506 -1389 -6479 -1333
rect -6423 -1334 -4732 -1333
rect -6423 -1389 -6335 -1334
rect -6506 -1390 -6335 -1389
rect -6279 -1390 -4732 -1334
rect -6506 -1424 -4732 -1390
rect -6506 -1459 -5130 -1424
rect -5194 -1524 -5130 -1459
rect -5030 -1524 -4840 -1424
rect -4740 -1524 -4731 -1424
rect -5194 -1556 -4732 -1524
rect -4391 -2562 -4262 -11
rect -4412 -2595 -4232 -2562
rect -4412 -2733 -4396 -2595
rect -4258 -2733 -4232 -2595
rect -4412 -2857 -4232 -2733
rect -4412 -2995 -4396 -2857
rect -4258 -2995 -4232 -2857
rect -4412 -3023 -4232 -2995
rect -3756 -5043 -3664 2769
rect -3352 2558 4590 2643
rect -3352 -3868 -3267 2558
rect -3091 2303 4206 2372
rect -3091 -3052 -3022 2303
rect -171 1908 3839 1976
rect -2883 889 -1765 945
rect -171 251 -103 1908
rect 3551 1799 3638 1807
rect 3524 1787 3638 1799
rect 3524 1700 3538 1787
rect 3625 1700 3638 1787
rect 3771 1784 3839 1908
rect 3524 1688 3638 1700
rect 3551 1457 3638 1688
rect 3745 1759 3839 1784
rect 3745 1693 3759 1759
rect 3825 1693 3839 1759
rect 3745 1682 3839 1693
rect 3771 1681 3839 1682
rect -2000 183 -103 251
rect 609 1370 3638 1457
rect -3133 -3058 -2988 -3052
rect -3133 -3127 -3091 -3058
rect -3022 -3127 -2988 -3058
rect -3133 -3227 -2988 -3127
rect -3133 -3296 -3091 -3227
rect -3022 -3296 -2988 -3227
rect -3133 -3460 -2988 -3296
rect -2000 -3230 -1932 183
rect 609 -331 696 1370
rect 4137 1185 4206 2303
rect 3900 1116 4206 1185
rect 3900 835 3969 1116
rect 3884 823 3982 835
rect 3458 796 3554 819
rect 3458 723 3471 796
rect 3544 723 3554 796
rect 3884 754 3900 823
rect 3969 754 3982 823
rect 3884 743 3982 754
rect 3458 711 3554 723
rect 3468 685 3554 711
rect 4505 685 4590 2558
rect 5566 1644 5658 2769
rect 6045 1986 6170 1998
rect 6045 1881 6053 1986
rect 6158 1881 6170 1986
rect 6045 1862 6170 1881
rect 5564 1636 5658 1644
rect 5564 1574 5581 1636
rect 5643 1631 5658 1636
rect 5643 1574 5656 1631
rect 5564 1559 5656 1574
rect 4675 708 4772 717
rect 4675 685 4686 708
rect 2230 646 2318 662
rect 2230 582 2244 646
rect 2308 582 2318 646
rect 2230 566 2318 582
rect 2962 645 3038 659
rect 2962 589 2971 645
rect 3027 589 3038 645
rect 3468 629 4686 685
rect 4759 629 4772 708
rect 3468 619 4772 629
rect 3468 612 4686 619
rect 4505 607 4590 612
rect 2962 574 3038 589
rect -1797 -418 696 -331
rect -1797 -3000 -1710 -418
rect 2250 -481 2306 566
rect 2445 494 2553 495
rect 2445 471 2556 494
rect 2445 401 2462 471
rect 2532 401 3432 471
rect 2445 391 2556 401
rect 2445 326 2554 391
rect 2445 257 2465 326
rect 2534 257 2554 326
rect 2445 168 2554 257
rect 3362 217 3432 401
rect 2445 99 2465 168
rect 2534 99 2554 168
rect 3350 205 3444 217
rect 3350 135 3362 205
rect 3432 135 3444 205
rect 3350 122 3444 135
rect 2445 88 2554 99
rect 2445 77 2553 88
rect 3147 -49 3228 -36
rect 3147 -105 3160 -49
rect 3216 -105 3228 -49
rect 3147 -117 3228 -105
rect 3553 -68 3637 -56
rect 2600 -406 2669 -401
rect -1294 -537 2306 -481
rect 2362 -417 2669 -406
rect 2362 -462 2603 -417
rect -1294 -731 -1238 -537
rect 2208 -732 2293 -717
rect 543 -802 2213 -732
rect 2283 -802 2293 -732
rect 2208 -813 2293 -802
rect 2074 -882 2174 -864
rect 513 -938 2096 -882
rect 2152 -938 2174 -882
rect 2074 -954 2174 -938
rect 2362 -1620 2418 -462
rect 2595 -473 2603 -462
rect 2659 -473 2669 -417
rect 2600 -486 2669 -473
rect 3160 -770 3216 -117
rect 3553 -124 3568 -68
rect 3624 -124 3637 -68
rect 3553 -136 3637 -124
rect 3966 -60 4045 -50
rect 3966 -116 3977 -60
rect 4033 -116 4045 -60
rect 3966 -130 4045 -116
rect 3150 -781 3229 -770
rect 3568 -777 3624 -136
rect 3977 -747 4033 -130
rect 3966 -758 4044 -747
rect 3150 -837 3160 -781
rect 3216 -837 3229 -781
rect 3150 -848 3229 -837
rect 3556 -788 3636 -777
rect 3556 -844 3568 -788
rect 3624 -844 3636 -788
rect 3966 -814 3977 -758
rect 4033 -814 4044 -758
rect 3966 -824 4044 -814
rect 3556 -855 3636 -844
rect 3568 -1052 3624 -855
rect 4778 -926 4880 -920
rect 4778 -930 4881 -926
rect 4778 -995 4801 -930
rect 4866 -995 4881 -930
rect 4778 -1007 4881 -995
rect 496 -1676 2418 -1620
rect 3536 -1110 3624 -1052
rect 3536 -1815 3592 -1110
rect 3853 -1330 3943 -1319
rect 3853 -1390 3866 -1330
rect 3928 -1390 4550 -1330
rect 3853 -1411 3943 -1390
rect 3524 -1827 3600 -1815
rect 3524 -1883 3536 -1827
rect 3592 -1883 3600 -1827
rect 3524 -1895 3600 -1883
rect 2079 -2755 2155 -2752
rect 3535 -2755 3591 -1895
rect 2079 -2780 3591 -2755
rect 2079 -2836 2089 -2780
rect 2145 -2811 3591 -2780
rect 2145 -2836 2155 -2811
rect 2079 -2849 2155 -2836
rect -576 -3000 -473 -2992
rect -1797 -3005 -473 -3000
rect -1797 -3087 -570 -3005
rect -576 -3092 -570 -3087
rect -483 -3092 -473 -3005
rect -576 -3106 -473 -3092
rect -644 -3230 -557 -3221
rect -2000 -3298 -635 -3230
rect -567 -3298 -557 -3230
rect -644 -3308 -557 -3298
rect -3133 -3529 -3091 -3460
rect -3022 -3529 -2988 -3460
rect -3133 -3551 -2988 -3529
rect -3120 -3556 -2999 -3551
rect -3352 -3879 -1469 -3868
rect -3352 -3944 -1545 -3879
rect -1480 -3944 -1469 -3879
rect -3352 -3953 -1469 -3944
rect -759 -4073 -643 -4072
rect -759 -4077 -547 -4073
rect -3117 -4090 -547 -4077
rect -3117 -4106 -631 -4090
rect -3117 -4175 -3091 -4106
rect -3022 -4159 -631 -4106
rect -562 -4159 -547 -4090
rect -3022 -4169 -547 -4159
rect -3022 -4175 -2996 -4169
rect -759 -4172 -547 -4169
rect -759 -4175 -643 -4172
rect -3117 -4205 -2996 -4175
rect 165 -4618 250 -4599
rect 165 -4683 176 -4618
rect 241 -4683 250 -4618
rect 165 -4699 250 -4683
rect -522 -4745 -447 -4733
rect -1657 -4806 -518 -4745
rect -457 -4806 -447 -4745
rect -1844 -5022 -1725 -5019
rect -2002 -5039 -1725 -5022
rect -2002 -5043 -1986 -5039
rect -3756 -5124 -1986 -5043
rect -1896 -5043 -1725 -5039
rect -1896 -5124 -1826 -5043
rect -3756 -5129 -1826 -5124
rect -1740 -5129 -1725 -5043
rect -3756 -5132 -3664 -5129
rect -2002 -5135 -1725 -5129
rect -1844 -5141 -1725 -5135
rect -1657 -6578 -1596 -4806
rect -522 -4820 -447 -4806
rect -641 -4952 -549 -4940
rect -641 -4963 -631 -4952
rect -642 -5014 -631 -4963
rect -569 -5014 -549 -4952
rect -642 -5044 -549 -5014
rect -558 -5332 -477 -5322
rect -750 -5392 -548 -5332
rect -488 -5392 -477 -5332
rect -750 -5814 -694 -5392
rect -558 -5402 -477 -5392
rect -761 -5826 -682 -5814
rect -761 -5882 -750 -5826
rect -694 -5882 -682 -5826
rect -761 -5893 -682 -5882
rect 174 -5818 241 -4699
rect 1573 -4996 1653 -4983
rect 1573 -5000 1580 -4996
rect 595 -5060 1580 -5000
rect 1644 -5060 1653 -4996
rect 595 -5065 1653 -5060
rect 595 -5596 660 -5065
rect 1573 -5071 1653 -5065
rect 3349 -5332 3426 -5323
rect 4490 -5332 4550 -1390
rect 3349 -5392 3355 -5332
rect 3415 -5392 4550 -5332
rect 3349 -5402 3426 -5392
rect 3357 -5471 3436 -5459
rect 4816 -5471 4881 -1007
rect 6059 -3262 6152 1862
rect 6059 -3355 6485 -3262
rect 4940 -3498 5014 -3482
rect 6250 -3498 6330 -3490
rect 4940 -3554 4948 -3498
rect 5004 -3554 6262 -3498
rect 6318 -3554 6330 -3498
rect 4940 -3568 5014 -3554
rect 6250 -3602 6330 -3554
rect 6250 -3658 6262 -3602
rect 6318 -3658 6330 -3602
rect 6250 -3670 6330 -3658
rect 3357 -5536 3361 -5471
rect 3426 -5536 4881 -5471
rect 3357 -5548 3436 -5536
rect 585 -5606 667 -5596
rect 585 -5671 595 -5606
rect 660 -5671 667 -5606
rect 585 -5682 667 -5671
rect 2499 -5606 2581 -5592
rect 2499 -5671 2503 -5606
rect 2568 -5671 3185 -5606
rect 2499 -5682 2581 -5671
rect 568 -5818 646 -5807
rect 174 -5885 573 -5818
rect 640 -5885 646 -5818
rect 568 -5895 646 -5885
rect 3120 -6273 3185 -5671
rect 5573 -6273 5666 -6263
rect 3120 -6338 5589 -6273
rect 5654 -6338 5666 -6273
rect 5573 -6350 5666 -6338
rect 6392 -6578 6485 -3355
rect -1657 -6644 6485 -6578
rect -1655 -6671 6485 -6644
rect -3690 -8198 -3330 -8178
rect -2365 -8198 -1628 -8190
rect -3690 -8299 -3675 -8198
rect -3574 -8299 -3437 -8198
rect -3336 -8216 -1628 -8198
rect -3336 -8217 -1777 -8216
rect -3336 -8222 -2006 -8217
rect -3336 -8299 -2276 -8222
rect -3690 -8329 -3330 -8299
rect -2365 -8344 -2276 -8299
rect -2141 -8339 -2006 -8222
rect -1871 -8338 -1777 -8217
rect -1642 -8338 -1628 -8216
rect -1871 -8339 -1628 -8338
rect -2141 -8344 -1628 -8339
rect -2365 -8366 -1628 -8344
rect -2327 -8367 -1628 -8366
use Balance_Inverter  Balance_Inverter_0
timestamp 1694400330
transform 1 0 -2144 0 1 -6278
box -29 0 1503 813
use Balance_Inverter  Balance_Inverter_1
timestamp 1694400330
transform 1 0 -2144 0 1 -5410
box -29 0 1503 813
use Balance_Inverter  Balance_Inverter_2
timestamp 1694400330
transform 1 0 -2144 0 1 -4551
box -29 0 1503 813
use Balance_Inverter  Balance_Inverter_3
timestamp 1694400330
transform 1 0 -2144 0 1 -3683
box -29 0 1503 813
use Balance_Inverter  Balance_Inverter_4
timestamp 1694400330
transform 1 0 -526 0 1 -6278
box -29 0 1503 813
use Balance_Inverter  Balance_Inverter_5
timestamp 1694400330
transform 1 0 1083 0 1 -6278
box -29 0 1503 813
use CM_32  CM_32_0
timestamp 1693893072
transform 1 0 -2794 0 -1 -7230
box -356 -267 6929 4816
use CM_LSB_mod  CM_LSB_mod_0
timestamp 1693830637
transform 1 0 -1877 0 1 -1203
box -3789 -772 4358 3860
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_140
timestamp 1692803904
transform 1 0 4987 0 1 616
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_141
timestamp 1692803904
transform 1 0 5395 0 1 918
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_142
timestamp 1692803904
transform 1 0 3710 0 1 1244
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_143
timestamp 1692803904
transform 1 0 3174 0 1 1244
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_144
timestamp 1692803904
transform 1 0 5599 0 1 918
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_145
timestamp 1692803904
transform 1 0 5803 0 1 918
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_146
timestamp 1692803904
transform 1 0 3700 0 1 -961
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_147
timestamp 1692803904
transform 1 0 3860 0 1 598
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_148
timestamp 1692803904
transform 1 0 4064 0 1 598
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_149
timestamp 1692803904
transform 1 0 4268 0 1 598
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_150
timestamp 1692803904
transform 1 0 5191 0 1 616
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_151
timestamp 1692803904
transform 1 0 5395 0 1 616
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_152
timestamp 1692803904
transform 1 0 5599 0 1 616
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_153
timestamp 1692803904
transform 1 0 5803 0 1 616
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_154
timestamp 1692803904
transform 1 0 3506 0 1 1244
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_155
timestamp 1692803904
transform 1 0 3656 0 1 598
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_156
timestamp 1692803904
transform 1 0 5191 0 1 918
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_157
timestamp 1692803904
transform 1 0 3914 0 1 1244
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_158
timestamp 1692803904
transform 1 0 3452 0 1 598
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_159
timestamp 1692803904
transform 1 0 4472 0 1 598
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_160
timestamp 1692803904
transform 1 0 4987 0 1 918
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_161
timestamp 1692803904
transform 1 0 4322 0 1 1244
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_162
timestamp 1692803904
transform 1 0 4118 0 1 1244
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_163
timestamp 1692803904
transform 1 0 3248 0 1 598
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_164
timestamp 1692803904
transform 1 0 3904 0 1 -961
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_165
timestamp 1692803904
transform 1 0 3292 0 1 -961
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_166
timestamp 1692803904
transform 1 0 3496 0 1 -961
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_167
timestamp 1692803904
transform 1 0 3088 0 1 74
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_168
timestamp 1692803904
transform 1 0 3700 0 1 74
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_169
timestamp 1692803904
transform 1 0 3496 0 1 74
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_170
timestamp 1692803904
transform 1 0 3904 0 1 74
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_171
timestamp 1692803904
transform 1 0 3292 0 1 -304
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_172
timestamp 1692803904
transform 1 0 3496 0 1 -304
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_173
timestamp 1692803904
transform 1 0 3700 0 1 -304
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_174
timestamp 1692803904
transform 1 0 3904 0 1 -304
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_175
timestamp 1692803904
transform 1 0 3292 0 1 -583
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_176
timestamp 1692803904
transform 1 0 3496 0 1 -583
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_177
timestamp 1692803904
transform 1 0 3700 0 1 -583
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_178
timestamp 1692803904
transform 1 0 3904 0 1 -583
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_179
timestamp 1692803904
transform 1 0 3292 0 1 74
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_180
timestamp 1692803904
transform 1 0 3088 0 1 -961
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_181
timestamp 1692803904
transform 1 0 3088 0 1 -304
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_182
timestamp 1692803904
transform 1 0 3088 0 1 -583
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_183
timestamp 1692803904
transform 1 0 4108 0 1 74
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_184
timestamp 1692803904
transform 1 0 4108 0 1 -961
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_185
timestamp 1692803904
transform 1 0 4108 0 1 -304
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_186
timestamp 1692803904
transform 1 0 4108 0 1 -583
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_187
timestamp 1692803904
transform 1 0 71 0 1 -4834
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_188
timestamp 1692803904
transform 1 0 4379 0 1 -3024
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_189
timestamp 1692803904
transform 1 0 683 0 1 -4834
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_190
timestamp 1692803904
transform 1 0 4175 0 1 -3024
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_191
timestamp 1692803904
transform 1 0 5247 0 1 -3024
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_192
timestamp 1692803904
transform 1 0 4711 0 1 -3024
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_193
timestamp 1692803904
transform 1 0 4915 0 1 -3024
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_194
timestamp 1692803904
transform 1 0 5987 0 1 -3024
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_195
timestamp 1692803904
transform 1 0 5451 0 1 -3024
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_196
timestamp 1692803904
transform 1 0 5783 0 1 -3024
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_197
timestamp 1692803904
transform 1 0 71 0 1 -2949
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_198
timestamp 1692803904
transform 1 0 4379 0 1 -2640
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_199
timestamp 1692803904
transform 1 0 4175 0 1 -2640
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_200
timestamp 1692803904
transform 1 0 3843 0 1 -2640
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_201
timestamp 1692803904
transform 1 0 5247 0 1 -2640
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_202
timestamp 1692803904
transform 1 0 4915 0 1 -2640
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_203
timestamp 1692803904
transform 1 0 4711 0 1 -2640
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_204
timestamp 1692803904
transform 1 0 5987 0 1 -2640
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_205
timestamp 1692803904
transform 1 0 5783 0 1 -2640
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_206
timestamp 1692803904
transform 1 0 5451 0 1 -2640
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_207
timestamp 1692803904
transform 1 0 71 0 1 -3233
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_208
timestamp 1692803904
transform 1 0 3843 0 1 -3024
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_209
timestamp 1692803904
transform 1 0 479 0 1 -4834
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_210
timestamp 1692803904
transform 1 0 275 0 1 -4834
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_211
timestamp 1692803904
transform 1 0 887 0 1 -4834
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_212
timestamp 1692803904
transform 1 0 1091 0 1 -4834
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_213
timestamp 1692803904
transform 1 0 1295 0 1 -4834
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_214
timestamp 1692803904
transform 1 0 1499 0 1 -4834
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_215
timestamp 1692803904
transform 1 0 1703 0 1 -4834
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_216
timestamp 1692803904
transform 1 0 2443 0 1 -4834
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_217
timestamp 1692803904
transform 1 0 3639 0 1 -5054
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_218
timestamp 1692803904
transform 1 0 4455 0 1 -5054
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_219
timestamp 1692803904
transform 1 0 2239 0 1 -4834
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_220
timestamp 1692803904
transform 1 0 1907 0 1 -4834
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_221
timestamp 1692803904
transform 1 0 4047 0 1 -5054
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_222
timestamp 1692803904
transform 1 0 4251 0 1 -5054
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_223
timestamp 1692803904
transform 1 0 3843 0 1 -5054
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_224
timestamp 1692803904
transform 1 0 5271 0 1 -5054
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_225
timestamp 1692803904
transform 1 0 4659 0 1 -5054
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_226
timestamp 1692803904
transform 1 0 4863 0 1 -5054
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_227
timestamp 1692803904
transform 1 0 5067 0 1 -5054
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_228
timestamp 1692803904
transform 1 0 5807 0 1 -5054
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_229
timestamp 1692803904
transform 1 0 6011 0 1 -5054
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_230
timestamp 1692803904
transform 1 0 5475 0 1 -5054
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_232
timestamp 1692803904
transform 1 0 3843 0 1 -5443
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_233
timestamp 1692803904
transform 1 0 4047 0 1 -5443
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_234
timestamp 1692803904
transform 1 0 4251 0 1 -5443
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_235
timestamp 1692803904
transform 1 0 4455 0 1 -5443
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_236
timestamp 1692803904
transform 1 0 4659 0 1 -5443
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_237
timestamp 1692803904
transform 1 0 4863 0 1 -5443
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_238
timestamp 1692803904
transform 1 0 5067 0 1 -5443
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_239
timestamp 1692803904
transform 1 0 5271 0 1 -5443
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_240
timestamp 1692803904
transform 1 0 5475 0 1 -5443
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_241
timestamp 1692803904
transform 1 0 5807 0 1 -5443
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_242
timestamp 1692803904
transform 1 0 6011 0 1 -5443
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_243
timestamp 1692803904
transform 1 0 3639 0 1 -5738
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_244
timestamp 1692803904
transform 1 0 4251 0 1 -5738
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_245
timestamp 1692803904
transform 1 0 4455 0 1 -5738
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_246
timestamp 1692803904
transform 1 0 3843 0 1 -5738
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_247
timestamp 1692803904
transform 1 0 4047 0 1 -5738
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_248
timestamp 1692803904
transform 1 0 5067 0 1 -5738
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_249
timestamp 1692803904
transform 1 0 5271 0 1 -5738
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_250
timestamp 1692803904
transform 1 0 4659 0 1 -5738
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_251
timestamp 1692803904
transform 1 0 4863 0 1 -5738
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_252
timestamp 1692803904
transform 1 0 6011 0 1 -5738
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_253
timestamp 1692803904
transform 1 0 5475 0 1 -5738
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_254
timestamp 1692803904
transform 1 0 5807 0 1 -5738
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_255
timestamp 1692803904
transform 1 0 607 0 1 -3233
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_256
timestamp 1692803904
transform 1 0 811 0 1 -3233
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_257
timestamp 1692803904
transform 1 0 275 0 1 -3233
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_258
timestamp 1692803904
transform 1 0 1679 0 1 -3233
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_259
timestamp 1692803904
transform 1 0 1143 0 1 -3233
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_260
timestamp 1692803904
transform 1 0 1347 0 1 -3233
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_261
timestamp 1692803904
transform 1 0 2419 0 1 -3233
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_262
timestamp 1692803904
transform 1 0 2215 0 1 -3233
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_263
timestamp 1692803904
transform 1 0 1883 0 1 -3233
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_264
timestamp 1692803904
transform 1 0 607 0 1 -2949
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_265
timestamp 1692803904
transform 1 0 811 0 1 -2949
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_266
timestamp 1692803904
transform 1 0 275 0 1 -2949
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_267
timestamp 1692803904
transform 1 0 1679 0 1 -2949
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_268
timestamp 1692803904
transform 1 0 1143 0 1 -2949
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_269
timestamp 1692803904
transform 1 0 1347 0 1 -2949
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_270
timestamp 1692803904
transform 1 0 2215 0 1 -2949
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_271
timestamp 1692803904
transform 1 0 2419 0 1 -2949
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_272
timestamp 1692803904
transform 1 0 1883 0 1 -2949
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_273
timestamp 1692803904
transform 1 0 3639 0 1 -2640
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_274
timestamp 1692803904
transform 1 0 3639 0 1 -3024
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_275
timestamp 1692803904
transform 1 0 3639 0 1 -1966
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_276
timestamp 1692803904
transform 1 0 3843 0 1 -1966
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_277
timestamp 1692803904
transform 1 0 3639 0 1 -2350
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_278
timestamp 1692803904
transform 1 0 3843 0 1 -2350
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_279
timestamp 1692803904
transform 1 0 4711 0 1 -1966
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_280
timestamp 1692803904
transform 1 0 4175 0 1 -1966
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_281
timestamp 1692803904
transform 1 0 4379 0 1 -1966
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_282
timestamp 1692803904
transform 1 0 4711 0 1 -2350
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_283
timestamp 1692803904
transform 1 0 4175 0 1 -2350
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_284
timestamp 1692803904
transform 1 0 4379 0 1 -2350
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_285
timestamp 1692803904
transform 1 0 5451 0 1 -2350
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_286
timestamp 1692803904
transform 1 0 5451 0 1 -1966
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_287
timestamp 1692803904
transform 1 0 5247 0 1 -1966
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_288
timestamp 1692803904
transform 1 0 4915 0 1 -1966
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_289
timestamp 1692803904
transform 1 0 5247 0 1 -2350
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_290
timestamp 1692803904
transform 1 0 4915 0 1 -2350
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_291
timestamp 1692803904
transform 1 0 5783 0 1 -2350
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_292
timestamp 1692803904
transform 1 0 5783 0 1 -1966
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_293
timestamp 1692803904
transform 1 0 5987 0 1 -2350
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_294
timestamp 1692803904
transform 1 0 5987 0 1 -1966
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_295
timestamp 1692803904
transform 1 0 3639 0 1 -6123
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_296
timestamp 1692803904
transform 1 0 3843 0 1 -6123
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_297
timestamp 1692803904
transform 1 0 4047 0 1 -6123
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_298
timestamp 1692803904
transform 1 0 4455 0 1 -6123
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_299
timestamp 1692803904
transform 1 0 4659 0 1 -6123
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_300
timestamp 1692803904
transform 1 0 4251 0 1 -6123
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_301
timestamp 1692803904
transform 1 0 5067 0 1 -6123
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_302
timestamp 1692803904
transform 1 0 5271 0 1 -6123
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_303
timestamp 1692803904
transform 1 0 5475 0 1 -6123
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_304
timestamp 1692803904
transform 1 0 4863 0 1 -6123
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_305
timestamp 1692803904
transform 1 0 5807 0 1 -6123
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_306
timestamp 1692803904
transform 1 0 6011 0 1 -6123
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_307
timestamp 1692803904
transform 1 0 71 0 1 -4449
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_308
timestamp 1692803904
transform 1 0 71 0 1 -4154
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_309
timestamp 1692803904
transform 1 0 479 0 1 -4449
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_310
timestamp 1692803904
transform 1 0 275 0 1 -4449
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_311
timestamp 1692803904
transform 1 0 683 0 1 -4449
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_312
timestamp 1692803904
transform 1 0 887 0 1 -4449
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_313
timestamp 1692803904
transform 1 0 479 0 1 -4154
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_314
timestamp 1692803904
transform 1 0 275 0 1 -4154
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_315
timestamp 1692803904
transform 1 0 683 0 1 -4154
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_316
timestamp 1692803904
transform 1 0 887 0 1 -4154
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_317
timestamp 1692803904
transform 1 0 1091 0 1 -4449
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_318
timestamp 1692803904
transform 1 0 1295 0 1 -4449
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_319
timestamp 1692803904
transform 1 0 1499 0 1 -4449
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_320
timestamp 1692803904
transform 1 0 1703 0 1 -4449
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_321
timestamp 1692803904
transform 1 0 1091 0 1 -4154
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_322
timestamp 1692803904
transform 1 0 1295 0 1 -4154
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_323
timestamp 1692803904
transform 1 0 1499 0 1 -4154
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_324
timestamp 1692803904
transform 1 0 1703 0 1 -4154
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_325
timestamp 1692803904
transform 1 0 2239 0 1 -4449
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_326
timestamp 1692803904
transform 1 0 2443 0 1 -4449
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_327
timestamp 1692803904
transform 1 0 2239 0 1 -4154
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_328
timestamp 1692803904
transform 1 0 2443 0 1 -4154
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_329
timestamp 1692803904
transform 1 0 1907 0 1 -4449
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_330
timestamp 1692803904
transform 1 0 1907 0 1 -4154
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_331
timestamp 1692803904
transform 1 0 71 0 1 -3765
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_332
timestamp 1692803904
transform 1 0 479 0 1 -3765
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_333
timestamp 1692803904
transform 1 0 683 0 1 -3765
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_334
timestamp 1692803904
transform 1 0 887 0 1 -3765
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_335
timestamp 1692803904
transform 1 0 275 0 1 -3765
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_336
timestamp 1692803904
transform 1 0 1703 0 1 -3765
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_337
timestamp 1692803904
transform 1 0 1091 0 1 -3765
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_338
timestamp 1692803904
transform 1 0 1295 0 1 -3765
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_339
timestamp 1692803904
transform 1 0 1499 0 1 -3765
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_340
timestamp 1692803904
transform 1 0 2239 0 1 -3765
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_341
timestamp 1692803904
transform 1 0 2443 0 1 -3765
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_342
timestamp 1692803904
transform 1 0 1907 0 1 -3765
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_343
timestamp 1692803904
transform 1 0 3843 0 1 -4342
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_344
timestamp 1692803904
transform 1 0 3639 0 1 -4342
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_345
timestamp 1692803904
transform 1 0 4047 0 1 -4342
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_346
timestamp 1692803904
transform 1 0 3639 0 1 -4727
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_347
timestamp 1692803904
transform 1 0 3843 0 1 -4727
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_348
timestamp 1692803904
transform 1 0 4047 0 1 -4727
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_349
timestamp 1692803904
transform 1 0 4455 0 1 -4342
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_350
timestamp 1692803904
transform 1 0 4659 0 1 -4342
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_351
timestamp 1692803904
transform 1 0 4251 0 1 -4342
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_352
timestamp 1692803904
transform 1 0 4455 0 1 -4727
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_353
timestamp 1692803904
transform 1 0 4251 0 1 -4727
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_354
timestamp 1692803904
transform 1 0 4659 0 1 -4727
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_355
timestamp 1692803904
transform 1 0 5067 0 1 -4342
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_356
timestamp 1692803904
transform 1 0 5271 0 1 -4342
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_357
timestamp 1692803904
transform 1 0 5475 0 1 -4342
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_358
timestamp 1692803904
transform 1 0 4863 0 1 -4342
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_359
timestamp 1692803904
transform 1 0 4863 0 1 -4727
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_360
timestamp 1692803904
transform 1 0 5067 0 1 -4727
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_361
timestamp 1692803904
transform 1 0 5271 0 1 -4727
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_362
timestamp 1692803904
transform 1 0 5475 0 1 -4727
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_363
timestamp 1692803904
transform 1 0 5807 0 1 -4342
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_364
timestamp 1692803904
transform 1 0 6011 0 1 -4342
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_365
timestamp 1692803904
transform 1 0 5807 0 1 -4727
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_366
timestamp 1692803904
transform 1 0 6011 0 1 -4727
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_367
timestamp 1692803904
transform 1 0 3843 0 1 -4047
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_368
timestamp 1692803904
transform 1 0 3639 0 1 -4047
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_369
timestamp 1692803904
transform 1 0 4047 0 1 -4047
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_370
timestamp 1692803904
transform 1 0 3843 0 1 -3658
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_371
timestamp 1692803904
transform 1 0 3639 0 1 -3658
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_372
timestamp 1692803904
transform 1 0 4047 0 1 -3658
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_373
timestamp 1692803904
transform 1 0 4455 0 1 -4047
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_374
timestamp 1692803904
transform 1 0 4659 0 1 -4047
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_375
timestamp 1692803904
transform 1 0 4455 0 1 -3658
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_376
timestamp 1692803904
transform 1 0 4659 0 1 -3658
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_377
timestamp 1692803904
transform 1 0 4251 0 1 -4047
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_378
timestamp 1692803904
transform 1 0 4251 0 1 -3658
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_379
timestamp 1692803904
transform 1 0 5067 0 1 -4047
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_380
timestamp 1692803904
transform 1 0 4863 0 1 -4047
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_381
timestamp 1692803904
transform 1 0 5271 0 1 -4047
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_382
timestamp 1692803904
transform 1 0 5475 0 1 -4047
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_383
timestamp 1692803904
transform 1 0 5067 0 1 -3658
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_384
timestamp 1692803904
transform 1 0 4863 0 1 -3658
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_385
timestamp 1692803904
transform 1 0 5271 0 1 -3658
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_386
timestamp 1692803904
transform 1 0 5475 0 1 -3658
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_387
timestamp 1692803904
transform 1 0 5807 0 1 -4047
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_388
timestamp 1692803904
transform 1 0 6011 0 1 -4047
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_389
timestamp 1692803904
transform 1 0 5807 0 1 -3658
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_390
timestamp 1692803904
transform 1 0 6011 0 1 -3658
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_391
timestamp 1692803904
transform 1 0 3639 0 1 -5443
box -162 -128 162 128
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_0
timestamp 1692705520
transform 1 0 4402 0 1 906
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_1
timestamp 1692705520
transform 1 0 3850 0 1 1534
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_2
timestamp 1692705520
transform 1 0 3170 0 1 1534
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_3
timestamp 1692705520
transform 1 0 4559 0 1 68
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_4
timestamp 1692705520
transform 1 0 5397 0 1 1468
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_5
timestamp 1692705520
transform 1 0 5609 0 1 1468
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_6
timestamp 1692705520
transform 1 0 3510 0 1 906
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_7
timestamp 1692705520
transform 1 0 3850 0 1 906
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_8
timestamp 1692705520
transform 1 0 4062 0 1 906
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_9
timestamp 1692705520
transform 1 0 5949 0 1 1226
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_10
timestamp 1692705520
transform 1 0 4845 0 1 1226
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_11
timestamp 1692705520
transform 1 0 5397 0 1 1226
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_12
timestamp 1692705520
transform 1 0 5609 0 1 1226
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_13
timestamp 1692705520
transform 1 0 5949 0 1 1468
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_14
timestamp 1692705520
transform 1 0 3510 0 1 1534
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_15
timestamp 1692705520
transform 1 0 3170 0 1 906
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_16
timestamp 1692705520
transform 1 0 5057 0 1 1226
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_17
timestamp 1692705520
transform 1 0 5057 0 1 1468
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_18
timestamp 1692705520
transform 1 0 4274 0 1 1534
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_19
timestamp 1692705520
transform 1 0 4062 0 1 1534
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_20
timestamp 1692705520
transform 1 0 4845 0 1 1468
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_21
timestamp 1692705520
transform 1 0 4899 0 1 68
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_22
timestamp 1692705520
transform 1 0 5111 0 1 68
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_23
timestamp 1692705520
transform 1 0 5451 0 1 68
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_24
timestamp 1692705520
transform 1 0 4558 0 1 -823
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_25
timestamp 1692705520
transform 1 0 4898 0 1 -823
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_26
timestamp 1692705520
transform 1 0 5110 0 1 -823
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_27
timestamp 1692705520
transform 1 0 5450 0 1 -823
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_28
timestamp 1692705520
transform 1 0 4558 0 1 -248
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_29
timestamp 1692705520
transform 1 0 4898 0 1 -248
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_30
timestamp 1692705520
transform 1 0 5110 0 1 -248
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_31
timestamp 1692705520
transform 1 0 5450 0 1 -248
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_32
timestamp 1692705520
transform 1 0 4558 0 1 -498
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_33
timestamp 1692705520
transform 1 0 4898 0 1 -498
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_34
timestamp 1692705520
transform 1 0 5110 0 1 -498
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_35
timestamp 1692705520
transform 1 0 5450 0 1 -498
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_36
timestamp 1692705520
transform 1 0 5663 0 1 68
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_37
timestamp 1692705520
transform 1 0 5662 0 1 -248
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_38
timestamp 1692705520
transform 1 0 5662 0 1 -823
box -166 -101 166 101
use nmos_3p3_MGEAJ7  nmos_3p3_MGEAJ7_39
timestamp 1692705520
transform 1 0 5662 0 1 -498
box -166 -101 166 101
use TG  TG_0
timestamp 1692688075
transform -1 0 3090 0 1 4510
box -2664 -1529 5711 271
use TG  TG_1
timestamp 1692688075
transform -1 0 3075 0 1 6424
box -2664 -1529 5711 271
<< labels >>
flabel metal1 -2331 -4136 -2331 -4136 0 FreeSans 480 0 0 0 B2
port 5 nsew
flabel metal3 -583 -3049 -583 -3049 0 FreeSans 800 0 0 0 b1
port 16 nsew
flabel metal3 -659 -3269 -659 -3269 0 FreeSans 800 0 0 0 b1b
port 17 nsew
flabel metal1 -576 -3918 -576 -3918 0 FreeSans 800 0 0 0 b2
port 18 nsew
flabel metal3 -672 -4125 -672 -4125 0 FreeSans 800 0 0 0 b2b
port 19 nsew
flabel metal3 -575 -4773 -575 -4773 0 FreeSans 800 0 0 0 b3
port 20 nsew
flabel metal1 -687 -4981 -687 -4981 0 FreeSans 800 0 0 0 b3b
port 21 nsew
flabel metal2 -686 -5647 -686 -5647 0 FreeSans 800 0 0 0 b4
port 22 nsew
flabel via2 -732 -5856 -732 -5856 0 FreeSans 800 0 0 0 b4b
port 23 nsew
flabel metal2 914 -5634 914 -5634 0 FreeSans 800 0 0 0 b5
port 24 nsew
flabel polycontact 881 -4634 881 -4634 0 FreeSans 800 0 0 0 b5b
port 25 nsew
flabel via1 5606 -5237 5606 -5237 0 FreeSans 800 0 0 0 b6
port 26 nsew
flabel via1 3498 -5922 3498 -5922 0 FreeSans 800 0 0 0 b6b
port 27 nsew
flabel metal1 -1815 -966 -1815 -966 0 FreeSans 1600 0 0 0 OUT1
port 30 nsew
flabel metal1 -1267 -1164 -1267 -1164 0 FreeSans 1600 0 0 0 OUT2
port 31 nsew
flabel metal1 -521 -1514 -521 -1514 0 FreeSans 800 0 0 0 OUT3
port 32 nsew
flabel metal1 -2801 -1521 -2801 -1521 0 FreeSans 800 0 0 0 OUT4
port 33 nsew
flabel metal1 1365 913 1365 913 0 FreeSans 800 0 0 0 OUT5
port 34 nsew
flabel metal1 1883 2066 1883 2066 0 FreeSans 800 0 0 0 OUT6
port 35 nsew
flabel metal1 -1596 -1280 -1596 -1280 0 FreeSans 480 0 0 0 G2
port 37 nsew
flabel metal1 -1597 -1045 -1597 -1045 0 FreeSans 480 0 0 0 SD2_2
port 38 nsew
flabel metal1 -2132 -1191 -2132 -1191 0 FreeSans 480 0 0 0 SD2_3
port 41 nsew
flabel metal1 -2998 -1166 -2998 -1166 0 FreeSans 480 0 0 0 SD2_5
port 42 nsew
flabel metal1 -3956 -1167 -3955 -1167 0 FreeSans 480 0 0 0 SD2_1
port 43 nsew
flabel metal1 -2468 -1173 -2468 -1173 0 FreeSans 480 0 0 0 SD2_4
port 44 nsew
flabel metal1 -2744 -400 -2744 -400 0 FreeSans 480 0 0 0 G1_2
port 45 nsew
flabel metal1 -3586 -300 -3586 -300 0 FreeSans 480 0 0 0 SD1_1
port 46 nsew
flabel metal1 -2853 -121 -2853 -121 0 FreeSans 480 0 0 0 G1_1
port 48 nsew
flabel metal1 -4166 2293 -4166 2293 0 FreeSans 480 0 0 0 SD3_1
port 51 nsew
flabel metal1 919 608 919 608 0 FreeSans 1600 0 0 0 SDn_1
port 52 nsew
flabel metal1 -2066 1187 -2066 1187 0 FreeSans 1600 0 0 0 SDn_2
port 53 nsew
flabel metal1 -4044 1266 -4044 1266 0 FreeSans 800 0 0 0 IT
port 54 nsew
flabel metal1 -6267 -3278 -6267 -3278 0 FreeSans 1600 0 0 0 B1
port 59 nsew
flabel metal1 -6262 -4145 -6262 -4145 0 FreeSans 1600 0 0 0 B2
port 60 nsew
flabel metal1 -6226 -5008 -6226 -5008 0 FreeSans 1600 0 0 0 B3
port 61 nsew
flabel metal1 -6175 -5859 -6175 -5859 0 FreeSans 1600 0 0 0 B4
port 62 nsew
flabel metal1 -6214 -6374 -6214 -6374 0 FreeSans 1600 0 0 0 B5
port 63 nsew
flabel metal1 -6221 -6581 -6221 -6581 0 FreeSans 1600 0 0 0 B6
port 64 nsew
flabel metal1 -5413 5151 -5413 5151 0 FreeSans 1600 0 0 0 OUT-
port 65 nsew
flabel metal1 -5768 3776 -5768 3776 0 FreeSans 1600 0 0 0 OUT+
port 66 nsew
flabel metal1 -6318 -2271 -6318 -2271 0 FreeSans 1600 0 0 0 VSS
port 70 nsew
flabel metal1 -6240 -2941 -6240 -2941 0 FreeSans 1600 0 0 0 VDD
port 71 nsew
flabel metal1 -6371 -1324 -6371 -1324 0 FreeSans 1600 0 0 0 ITAIL
port 72 nsew
flabel metal1 -3633 -12206 -3633 -12206 0 FreeSans 1600 0 0 0 C32_D
port 74 nsew
flabel metal1 -3653 -12455 -3653 -12455 0 FreeSans 1600 0 0 0 C32_U
port 75 nsew
flabel metal1 6284 6502 6284 6502 0 FreeSans 1600 0 0 0 SEL_L
port 76 nsew
flabel metal1 -2531 -7305 -2531 -7305 0 FreeSans 800 0 0 0 SDc_1
port 77 nsew
flabel metal1 -2997 -8619 -2997 -8619 0 FreeSans 800 0 0 0 Gc_1
port 78 nsew
flabel metal1 -1980 -8955 -1980 -8955 0 FreeSans 800 0 0 0 Gc_2
port 79 nsew
flabel metal1 -2579 -9795 -2579 -9795 0 FreeSans 800 0 0 0 SDc_2
port 80 nsew
<< end >>
