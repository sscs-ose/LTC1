magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2208 -2120 3080 3120
<< nwell >>
rect -208 -120 1080 1120
<< mvpmos >>
rect 0 0 140 1000
rect 244 0 384 1000
rect 488 0 628 1000
rect 732 0 872 1000
<< mvpdiff >>
rect -88 987 0 1000
rect -88 941 -75 987
rect -29 941 0 987
rect -88 884 0 941
rect -88 838 -75 884
rect -29 838 0 884
rect -88 781 0 838
rect -88 735 -75 781
rect -29 735 0 781
rect -88 678 0 735
rect -88 632 -75 678
rect -29 632 0 678
rect -88 575 0 632
rect -88 529 -75 575
rect -29 529 0 575
rect -88 472 0 529
rect -88 426 -75 472
rect -29 426 0 472
rect -88 369 0 426
rect -88 323 -75 369
rect -29 323 0 369
rect -88 266 0 323
rect -88 220 -75 266
rect -29 220 0 266
rect -88 163 0 220
rect -88 117 -75 163
rect -29 117 0 163
rect -88 59 0 117
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 140 987 244 1000
rect 140 941 169 987
rect 215 941 244 987
rect 140 884 244 941
rect 140 838 169 884
rect 215 838 244 884
rect 140 781 244 838
rect 140 735 169 781
rect 215 735 244 781
rect 140 678 244 735
rect 140 632 169 678
rect 215 632 244 678
rect 140 575 244 632
rect 140 529 169 575
rect 215 529 244 575
rect 140 472 244 529
rect 140 426 169 472
rect 215 426 244 472
rect 140 369 244 426
rect 140 323 169 369
rect 215 323 244 369
rect 140 266 244 323
rect 140 220 169 266
rect 215 220 244 266
rect 140 163 244 220
rect 140 117 169 163
rect 215 117 244 163
rect 140 59 244 117
rect 140 13 169 59
rect 215 13 244 59
rect 140 0 244 13
rect 384 987 488 1000
rect 384 941 413 987
rect 459 941 488 987
rect 384 884 488 941
rect 384 838 413 884
rect 459 838 488 884
rect 384 781 488 838
rect 384 735 413 781
rect 459 735 488 781
rect 384 678 488 735
rect 384 632 413 678
rect 459 632 488 678
rect 384 575 488 632
rect 384 529 413 575
rect 459 529 488 575
rect 384 472 488 529
rect 384 426 413 472
rect 459 426 488 472
rect 384 369 488 426
rect 384 323 413 369
rect 459 323 488 369
rect 384 266 488 323
rect 384 220 413 266
rect 459 220 488 266
rect 384 163 488 220
rect 384 117 413 163
rect 459 117 488 163
rect 384 59 488 117
rect 384 13 413 59
rect 459 13 488 59
rect 384 0 488 13
rect 628 987 732 1000
rect 628 941 657 987
rect 703 941 732 987
rect 628 884 732 941
rect 628 838 657 884
rect 703 838 732 884
rect 628 781 732 838
rect 628 735 657 781
rect 703 735 732 781
rect 628 678 732 735
rect 628 632 657 678
rect 703 632 732 678
rect 628 575 732 632
rect 628 529 657 575
rect 703 529 732 575
rect 628 472 732 529
rect 628 426 657 472
rect 703 426 732 472
rect 628 369 732 426
rect 628 323 657 369
rect 703 323 732 369
rect 628 266 732 323
rect 628 220 657 266
rect 703 220 732 266
rect 628 163 732 220
rect 628 117 657 163
rect 703 117 732 163
rect 628 59 732 117
rect 628 13 657 59
rect 703 13 732 59
rect 628 0 732 13
rect 872 987 960 1000
rect 872 941 901 987
rect 947 941 960 987
rect 872 884 960 941
rect 872 838 901 884
rect 947 838 960 884
rect 872 781 960 838
rect 872 735 901 781
rect 947 735 960 781
rect 872 678 960 735
rect 872 632 901 678
rect 947 632 960 678
rect 872 575 960 632
rect 872 529 901 575
rect 947 529 960 575
rect 872 472 960 529
rect 872 426 901 472
rect 947 426 960 472
rect 872 369 960 426
rect 872 323 901 369
rect 947 323 960 369
rect 872 266 960 323
rect 872 220 901 266
rect 947 220 960 266
rect 872 163 960 220
rect 872 117 901 163
rect 947 117 960 163
rect 872 59 960 117
rect 872 13 901 59
rect 947 13 960 59
rect 872 0 960 13
<< mvpdiffc >>
rect -75 941 -29 987
rect -75 838 -29 884
rect -75 735 -29 781
rect -75 632 -29 678
rect -75 529 -29 575
rect -75 426 -29 472
rect -75 323 -29 369
rect -75 220 -29 266
rect -75 117 -29 163
rect -75 13 -29 59
rect 169 941 215 987
rect 169 838 215 884
rect 169 735 215 781
rect 169 632 215 678
rect 169 529 215 575
rect 169 426 215 472
rect 169 323 215 369
rect 169 220 215 266
rect 169 117 215 163
rect 169 13 215 59
rect 413 941 459 987
rect 413 838 459 884
rect 413 735 459 781
rect 413 632 459 678
rect 413 529 459 575
rect 413 426 459 472
rect 413 323 459 369
rect 413 220 459 266
rect 413 117 459 163
rect 413 13 459 59
rect 657 941 703 987
rect 657 838 703 884
rect 657 735 703 781
rect 657 632 703 678
rect 657 529 703 575
rect 657 426 703 472
rect 657 323 703 369
rect 657 220 703 266
rect 657 117 703 163
rect 657 13 703 59
rect 901 941 947 987
rect 901 838 947 884
rect 901 735 947 781
rect 901 632 947 678
rect 901 529 947 575
rect 901 426 947 472
rect 901 323 947 369
rect 901 220 947 266
rect 901 117 947 163
rect 901 13 947 59
<< polysilicon >>
rect 0 1000 140 1044
rect 244 1000 384 1044
rect 488 1000 628 1044
rect 732 1000 872 1044
rect 0 -44 140 0
rect 244 -44 384 0
rect 488 -44 628 0
rect 732 -44 872 0
<< metal1 >>
rect -75 987 -29 1000
rect -75 884 -29 941
rect -75 781 -29 838
rect -75 678 -29 735
rect -75 575 -29 632
rect -75 472 -29 529
rect -75 369 -29 426
rect -75 266 -29 323
rect -75 163 -29 220
rect -75 59 -29 117
rect -75 0 -29 13
rect 169 987 215 1000
rect 169 884 215 941
rect 169 781 215 838
rect 169 678 215 735
rect 169 575 215 632
rect 169 472 215 529
rect 169 369 215 426
rect 169 266 215 323
rect 169 163 215 220
rect 169 59 215 117
rect 169 0 215 13
rect 413 987 459 1000
rect 413 884 459 941
rect 413 781 459 838
rect 413 678 459 735
rect 413 575 459 632
rect 413 472 459 529
rect 413 369 459 426
rect 413 266 459 323
rect 413 163 459 220
rect 413 59 459 117
rect 413 0 459 13
rect 657 987 703 1000
rect 657 884 703 941
rect 657 781 703 838
rect 657 678 703 735
rect 657 575 703 632
rect 657 472 703 529
rect 657 369 703 426
rect 657 266 703 323
rect 657 163 703 220
rect 657 59 703 117
rect 657 0 703 13
rect 901 987 947 1000
rect 901 884 947 941
rect 901 781 947 838
rect 901 678 947 735
rect 901 575 947 632
rect 901 472 947 529
rect 901 369 947 426
rect 901 266 947 323
rect 901 163 947 220
rect 901 59 947 117
rect 901 0 947 13
<< labels >>
rlabel metal1 680 500 680 500 4 D
rlabel metal1 436 500 436 500 4 S
rlabel metal1 192 500 192 500 4 D
rlabel metal1 924 500 924 500 4 S
rlabel metal1 -52 500 -52 500 4 S
<< end >>
