* NGSPICE file created from therm_Dec_flat.ext - technology: gf180mcuC

.subckt therm_Dec_flat VDD VSS D1 D2 D4 D3 D5 D6 D7 B3 B2 B1
X0 a_268_n4206# B1.t0 OR_4.Inverter_0.IN VDD.t63 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X1 a_1557_n2284# B1.t1 OR_1.Inverter_0.IN VDD.t62 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X2 OR_3.OUT OR_3.Inverter_0.IN VDD.t16 VDD.t15 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X3 D2 INV_BUFF_1.Inverter_0.IN VSS.t19 VSS.t18 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X4 INV_BUFF_1.Inverter_0.IN AND_2.OUT VSS.t72 VSS.t71 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X5 a_268_215# B1.t2 VSS.t46 VSS.t45 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X6 OR_3.Inverter_0.IN B3.t0 VSS.t5 VSS.t4 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X7 AND_3.Inverter_0.IN B1.t3 VDD.t61 VDD.t60 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X8 VDD B2.t0 AND_1.Inverter_0.IN VDD.t4 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X9 a_268_n3244# B1.t4 OR_2.Inverter_0.IN VDD.t59 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X10 OR_1.Inverter_0.IN OR_1.B VSS.t23 VSS.t22 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X11 AND_0.OUT AND_0.Inverter_0.IN VSS.t1 VSS.t0 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X12 a_268_n2622# B2.t1 VSS.t21 VSS.t20 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X13 AND_2.OUT AND_2.Inverter_0.IN VSS.t54 VSS.t53 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X14 a_268_n1326# B2.t2 OR_0.Inverter_0.IN VDD.t74 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X15 OR_3.B OR_4.Inverter_0.IN VSS.t17 VSS.t16 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X16 OR_4.Inverter_0.IN B1.t5 a_268_n4206# VDD.t58 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X17 OR_1.Inverter_0.IN B1.t6 a_1557_n2284# VDD.t57 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X18 INV_BUFF_2.Inverter_0.IN AND_3.OUT VSS.t58 VSS.t57 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X19 INV_BUFF_5.Inverter_0.IN OR_2.OUT VSS.t68 VSS.t67 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X20 INV_BUFF_4.Inverter_0.IN OR_1.OUT VDD.t18 VDD.t17 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X21 OR_1.B AND_4.Inverter_0.IN VDD.t78 VDD.t77 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X22 D4 INV_BUFF_3.Inverter_0.IN VDD.t43 VDD.t42 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X23 INV_BUFF_6.Inverter_0.IN OR_3.OUT VSS.t60 VSS.t59 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X24 VDD OR_3.B a_1840_n4206# VDD.t12 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X25 AND_0.Inverter_0.IN AND_0.B a_1628_215# VSS.t50 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X26 AND_0.Inverter_0.IN B3.t1 VDD.t92 VDD.t91 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X27 OR_4.Inverter_0.IN B2.t3 VSS.t76 VSS.t75 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X28 a_268_n4206# B2.t4 VDD.t45 VDD.t44 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X29 OR_2.OUT OR_2.Inverter_0.IN VSS.t3 VSS.t2 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X30 INV_BUFF_3.Inverter_0.IN B1.t7 VSS.t44 VSS.t43 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X31 OR_2.Inverter_0.IN B1.t8 a_268_n3244# VDD.t56 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X32 D5 INV_BUFF_4.Inverter_0.IN VSS.t32 VSS.t31 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X33 VDD B3.t2 AND_4.Inverter_0.IN VDD.t93 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X34 AND_2.Inverter_0.IN B1.t9 VDD.t55 VDD.t54 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X35 INV_BUFF_1.Inverter_0.IN AND_2.OUT VDD.t102 VDD.t101 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X36 VDD B2.t5 AND_2.Inverter_0.IN VDD.t69 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X37 a_1840_n4206# B3.t3 OR_3.Inverter_0.IN VDD.t21 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X38 AND_3.B OR_0.Inverter_0.IN VSS.t64 VSS.t63 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X39 D2 INV_BUFF_1.Inverter_0.IN VDD.t28 VDD.t27 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X40 OR_1.OUT OR_1.Inverter_0.IN VSS.t74 VSS.t73 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X41 INV_BUFF_0.Inverter_0.IN AND_0.OUT VDD.t97 VDD.t96 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X42 D3 INV_BUFF_2.Inverter_0.IN VSS.t52 VSS.t51 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X43 OR_0.Inverter_0.IN B2.t6 a_268_n1326# VDD.t41 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X44 OR_2.Inverter_0.IN B2.t7 VSS.t28 VSS.t27 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X45 D7 INV_BUFF_6.Inverter_0.IN VSS.t66 VSS.t65 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X46 a_1557_n2284# OR_1.B VDD.t35 VDD.t34 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X47 AND_3.OUT AND_3.Inverter_0.IN VSS.t13 VSS.t12 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X48 VDD AND_3.B AND_3.Inverter_0.IN VDD.t38 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X49 a_268_n3244# B2.t8 VDD.t30 VDD.t29 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X50 AND_2.OUT AND_2.Inverter_0.IN VDD.t76 VDD.t75 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X51 a_1840_n4206# OR_3.B VDD.t11 VDD.t10 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X52 OR_0.Inverter_0.IN B3.t4 VSS.t15 VSS.t14 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X53 OR_3.B OR_4.Inverter_0.IN VDD.t26 VDD.t25 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X54 OR_1.Inverter_0.IN B1.t10 VSS.t42 VSS.t41 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X55 INV_BUFF_2.Inverter_0.IN AND_3.OUT VDD.t80 VDD.t79 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X56 a_268_n1326# B3.t5 VDD.t8 VDD.t7 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X57 INV_BUFF_5.Inverter_0.IN OR_2.OUT VDD.t90 VDD.t89 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X58 INV_BUFF_6.Inverter_0.IN OR_3.OUT VDD.t82 VDD.t81 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X59 D6 INV_BUFF_5.Inverter_0.IN VSS.t48 VSS.t47 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X60 OR_3.Inverter_0.IN B3.t6 a_1840_n4206# VDD.t9 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X61 a_1881_n1685# B1.t11 VSS.t40 VSS.t39 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X62 AND_1.Inverter_0.IN B2.t9 a_268_215# VSS.t80 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X63 AND_0.B AND_1.Inverter_0.IN VDD.t84 VDD.t83 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X64 AND_4.Inverter_0.IN B3.t7 a_268_n2622# VSS.t77 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X65 a_268_n724# B1.t12 VSS.t38 VSS.t37 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X66 AND_2.Inverter_0.IN B2.t10 a_268_n724# VSS.t49 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X67 AND_1.Inverter_0.IN B1.t13 VDD.t53 VDD.t52 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X68 OR_2.OUT OR_2.Inverter_0.IN VDD.t3 VDD.t2 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X69 INV_BUFF_3.Inverter_0.IN B1.t14 VDD.t51 VDD.t50 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X70 INV_BUFF_0.Inverter_0.IN AND_0.OUT VSS.t70 VSS.t69 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X71 D5 INV_BUFF_4.Inverter_0.IN VDD.t49 VDD.t48 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X72 D1 INV_BUFF_0.Inverter_0.IN VDD.t47 VDD.t46 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X73 AND_3.B OR_0.Inverter_0.IN VDD.t86 VDD.t85 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X74 OR_1.OUT OR_1.Inverter_0.IN VDD.t104 VDD.t103 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X75 D3 INV_BUFF_2.Inverter_0.IN VDD.t73 VDD.t72 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X76 D7 INV_BUFF_6.Inverter_0.IN VDD.t88 VDD.t87 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X77 AND_3.OUT AND_3.Inverter_0.IN VDD.t20 VDD.t19 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X78 OR_4.Inverter_0.IN B1.t15 VSS.t36 VSS.t35 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X79 a_1628_215# B3.t8 VSS.t79 VSS.t78 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X80 OR_3.OUT OR_3.Inverter_0.IN VSS.t9 VSS.t8 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X81 OR_3.Inverter_0.IN OR_3.B VSS.t7 VSS.t6 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X82 VDD B2.t11 a_268_n4206# VDD.t98 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X83 VDD AND_0.B AND_0.Inverter_0.IN VDD.t66 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X84 AND_0.B AND_1.Inverter_0.IN VSS.t62 VSS.t61 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X85 D6 INV_BUFF_5.Inverter_0.IN VDD.t65 VDD.t64 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X86 OR_2.Inverter_0.IN B1.t16 VSS.t34 VSS.t33 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X87 VDD OR_1.B a_1557_n2284# VDD.t31 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X88 D1 INV_BUFF_0.Inverter_0.IN VSS.t30 VSS.t29 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X89 VDD B2.t12 a_268_n3244# VDD.t105 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X90 AND_3.Inverter_0.IN AND_3.B a_1881_n1685# VSS.t24 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X91 OR_0.Inverter_0.IN B2.t13 VSS.t82 VSS.t81 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X92 INV_BUFF_4.Inverter_0.IN OR_1.OUT VSS.t11 VSS.t10 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X93 OR_1.B AND_4.Inverter_0.IN VSS.t56 VSS.t55 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X94 AND_4.Inverter_0.IN B2.t14 VDD.t37 VDD.t36 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X95 AND_0.OUT AND_0.Inverter_0.IN VDD.t1 VDD.t0 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X96 D4 INV_BUFF_3.Inverter_0.IN VSS.t26 VSS.t25 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X97 VDD B3.t9 a_268_n1326# VDD.t22 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
R0 B1.t6 B1.t1 44.4957
R1 B1.t8 B1.t4 44.4957
R2 B1.t5 B1.t0 44.4957
R3 B1 B1.n0 32.7242
R4 B1.n0 B1.t2 31.938
R5 B1.n1 B1.t12 31.938
R6 B1.n6 B1.t11 31.938
R7 B1.n7 B1.n6 31.598
R8 B1.n8 B1.t10 27.2239
R9 B1.n10 B1.t16 27.2239
R10 B1.n11 B1.t15 27.2239
R11 B1.n2 B1.n1 26.2635
R12 B1.n4 B1.t7 19.0247
R13 B1.n4 B1.t14 17.3935
R14 B1.n8 B1.t6 15.0244
R15 B1.n10 B1.t8 15.0244
R16 B1.n11 B1.t5 15.0244
R17 B1.n0 B1.t13 12.2541
R18 B1.n1 B1.t9 12.2541
R19 B1.n6 B1.t3 12.2541
R20 B1.n14 B1.n7 10.375
R21 B1.n13 B1.n9 10.1883
R22 B1.n5 B1 8.08376
R23 B1 B1.n10 5.30993
R24 B1 B1.n11 5.30993
R25 B1.n9 B1.n8 5.29037
R26 B1.n12 B1 5.05067
R27 B1.n3 B1.n2 4.96776
R28 B1 B1.n15 4.75904
R29 B1 B1.n4 4.15272
R30 B1.n12 B1 3.53829
R31 B1.n15 B1.n5 3.24798
R32 B1.n14 B1.n13 2.14814
R33 B1.n2 B1 1.79407
R34 B1.n15 B1.n14 1.28892
R35 B1.n13 B1.n12 1.14672
R36 B1.n9 B1 0.0200652
R37 B1.n5 B1.n3 0.0119745
R38 B1.n7 B1 0.0067069
R39 B1.n3 B1 0.00153448
R40 VDD.n4 VDD.t0 1130.33
R41 VDD.t10 VDD.t25 948.718
R42 VDD.t19 VDD.n32 943.129
R43 VDD.t101 VDD.n19 917.062
R44 VDD.t50 VDD.n16 917.062
R45 VDD.n30 VDD.t79 917.062
R46 VDD.n49 VDD.t17 917.062
R47 VDD.n66 VDD.t89 917.062
R48 VDD.t81 VDD.n81 917.062
R49 VDD.t96 VDD.n3 917.062
R50 VDD.n33 VDD.t38 870.938
R51 VDD.t66 VDD.n7 870.938
R52 VDD.t21 VDD.n83 826.923
R53 VDD.t63 VDD.n88 826.923
R54 VDD.n60 VDD.t34 598.292
R55 VDD.n52 VDD.n51 464.455
R56 VDD.n41 VDD.t41 448.719
R57 VDD.n59 VDD.t57 448.719
R58 VDD.n72 VDD.t56 448.719
R59 VDD.n84 VDD.t9 448.719
R60 VDD.n89 VDD.t58 448.719
R61 VDD.n12 VDD.t4 443.255
R62 VDD.n23 VDD.t69 443.255
R63 VDD.n38 VDD.t38 443.255
R64 VDD.n61 VDD.t93 443.255
R65 VDD.n8 VDD.t66 443.255
R66 VDD.t4 VDD.n10 432.548
R67 VDD.t69 VDD.n22 432.548
R68 VDD.t93 VDD.n60 432.548
R69 VDD.t74 VDD.n40 431.625
R70 VDD.n53 VDD.t62 431.625
R71 VDD.t59 VDD.n71 431.625
R72 VDD.n12 VDD.t52 421.842
R73 VDD.n23 VDD.t54 421.842
R74 VDD.t60 VDD.n38 421.842
R75 VDD.n61 VDD.t36 421.842
R76 VDD.n8 VDD.t91 421.842
R77 VDD.n41 VDD.t22 414.531
R78 VDD.t31 VDD.n59 414.531
R79 VDD.n72 VDD.t105 414.531
R80 VDD.n84 VDD.t12 414.531
R81 VDD.n89 VDD.t98 414.531
R82 VDD.n70 VDD.n69 407.034
R83 VDD.t41 VDD.t74 341.88
R84 VDD.t22 VDD.t7 341.88
R85 VDD.t62 VDD.t57 341.88
R86 VDD.t34 VDD.t31 341.88
R87 VDD.t56 VDD.t59 341.88
R88 VDD.t105 VDD.t29 341.88
R89 VDD.t9 VDD.t21 341.88
R90 VDD.t12 VDD.t10 341.88
R91 VDD.t58 VDD.t63 341.88
R92 VDD.t98 VDD.t44 341.88
R93 VDD.n60 VDD 316.474
R94 VDD.n22 VDD 315.707
R95 VDD VDD.n10 315.707
R96 VDD.n39 VDD.t60 254.819
R97 VDD.n53 VDD.n52 188.119
R98 VDD.n71 VDD.n70 181.667
R99 VDD VDD.n53 167.191
R100 VDD.n71 VDD 159.602
R101 VDD.n39 VDD.t85 151.409
R102 VDD.n40 VDD 120.737
R103 VDD.n10 VDD.t83 116.338
R104 VDD.n22 VDD.t75 116.338
R105 VDD.n60 VDD.t77 115.803
R106 VDD.n52 VDD.t103 76.7332
R107 VDD.n70 VDD.t2 69.9242
R108 VDD VDD.t50 46.5849
R109 VDD VDD.t101 46.5849
R110 VDD VDD.t81 46.5849
R111 VDD.n19 VDD.t27 40.2849
R112 VDD.n16 VDD.t42 40.2849
R113 VDD.n30 VDD.t72 40.2849
R114 VDD.n32 VDD.t79 40.2849
R115 VDD.n33 VDD.t19 40.2849
R116 VDD.n49 VDD.t48 40.2849
R117 VDD.n51 VDD.t17 40.2849
R118 VDD.n66 VDD.t64 40.2849
R119 VDD.n69 VDD.t89 40.2849
R120 VDD.n81 VDD.t87 40.2849
R121 VDD.n3 VDD.t46 40.2849
R122 VDD.n4 VDD.t96 40.2849
R123 VDD.n7 VDD.t0 40.2849
R124 VDD.n40 VDD.n39 36.9723
R125 VDD.n83 VDD.t15 36.3253
R126 VDD.n88 VDD.t25 36.3253
R127 VDD.n44 VDD.t8 6.61028
R128 VDD.n43 VDD.n26 6.61028
R129 VDD.n56 VDD.t35 6.61028
R130 VDD.n57 VDD.n55 6.61028
R131 VDD.n75 VDD.t30 6.61028
R132 VDD.n74 VDD.n64 6.61028
R133 VDD.n87 VDD.t11 6.61028
R134 VDD.n86 VDD.n78 6.61028
R135 VDD.n92 VDD.t45 6.61028
R136 VDD.n91 VDD.n76 6.61028
R137 VDD.n25 VDD.t55 6.57115
R138 VDD.n14 VDD.n13 6.57115
R139 VDD.n36 VDD.t61 6.57115
R140 VDD.n35 VDD.n28 6.57115
R141 VDD.n63 VDD.t37 6.57115
R142 VDD.n46 VDD.n45 6.57115
R143 VDD.n97 VDD.t53 6.57115
R144 VDD.n99 VDD.n11 6.57115
R145 VDD.n101 VDD.t92 6.57115
R146 VDD.n1 VDD.n0 6.57115
R147 VDD.n17 VDD.t51 6.40636
R148 VDD.n15 VDD.t43 6.40636
R149 VDD.n21 VDD.t76 6.40636
R150 VDD.n20 VDD.t102 6.40636
R151 VDD.n18 VDD.t28 6.40636
R152 VDD.n34 VDD.t20 6.40636
R153 VDD.n29 VDD.t80 6.40636
R154 VDD.n31 VDD.t73 6.40636
R155 VDD.n27 VDD.t86 6.40636
R156 VDD.n54 VDD.t104 6.40636
R157 VDD.n48 VDD.t18 6.40636
R158 VDD.n50 VDD.t49 6.40636
R159 VDD.n47 VDD.t78 6.40636
R160 VDD.n65 VDD.t3 6.40636
R161 VDD.n68 VDD.t90 6.40636
R162 VDD.n67 VDD.t65 6.40636
R163 VDD.n82 VDD.t82 6.40636
R164 VDD.n80 VDD.t88 6.40636
R165 VDD.n79 VDD.t16 6.40636
R166 VDD.n77 VDD.t26 6.40636
R167 VDD.n100 VDD.t84 6.40636
R168 VDD.n6 VDD.t1 6.40636
R169 VDD.n5 VDD.t97 6.40636
R170 VDD.n2 VDD.t47 6.40636
R171 VDD.n16 VDD 6.3005
R172 VDD.n19 VDD 6.3005
R173 VDD.n24 VDD.n23 6.3005
R174 VDD VDD.n33 6.3005
R175 VDD.n32 VDD 6.3005
R176 VDD VDD.n30 6.3005
R177 VDD.n38 VDD.n37 6.3005
R178 VDD.n42 VDD.n41 6.3005
R179 VDD.n51 VDD 6.3005
R180 VDD VDD.n49 6.3005
R181 VDD.n59 VDD.n58 6.3005
R182 VDD.n62 VDD.n61 6.3005
R183 VDD.n69 VDD 6.3005
R184 VDD VDD.n66 6.3005
R185 VDD.n73 VDD.n72 6.3005
R186 VDD.n81 VDD 6.3005
R187 VDD.n83 VDD 6.3005
R188 VDD.n85 VDD.n84 6.3005
R189 VDD.n88 VDD 6.3005
R190 VDD.n90 VDD.n89 6.3005
R191 VDD.n98 VDD.n12 6.3005
R192 VDD.n7 VDD 6.3005
R193 VDD VDD.n4 6.3005
R194 VDD.n3 VDD 6.3005
R195 VDD.n9 VDD.n8 6.3005
R196 VDD.n93 VDD.n92 5.17727
R197 VDD.n97 VDD.n96 5.11649
R198 VDD.n95 VDD.n44 3.66683
R199 VDD.n93 VDD.n75 3.65957
R200 VDD.n96 VDD.n25 3.65055
R201 VDD.n94 VDD.n63 3.64928
R202 VDD.n95 VDD.n94 1.52123
R203 VDD.n94 VDD.n93 1.47616
R204 VDD.n96 VDD.n95 1.46275
R205 VDD.n42 VDD.n27 0.567623
R206 VDD.n58 VDD.n54 0.567623
R207 VDD.n73 VDD.n65 0.567623
R208 VDD.n85 VDD.n79 0.567623
R209 VDD.n90 VDD.n77 0.567623
R210 VDD VDD.n17 0.522334
R211 VDD.n44 VDD.n43 0.291409
R212 VDD.n57 VDD.n56 0.291409
R213 VDD.n75 VDD.n74 0.291409
R214 VDD.n87 VDD.n86 0.291409
R215 VDD.n92 VDD.n91 0.291409
R216 VDD.n56 VDD 0.284603
R217 VDD.n36 VDD 0.246101
R218 VDD VDD.n87 0.240744
R219 VDD VDD.n82 0.23967
R220 VDD.n24 VDD.n14 0.219398
R221 VDD.n62 VDD.n46 0.219398
R222 VDD.n99 VDD.n98 0.219398
R223 VDD.n9 VDD.n1 0.219398
R224 VDD VDD.n20 0.213013
R225 VDD VDD.n5 0.198406
R226 VDD.n37 VDD.n35 0.186327
R227 VDD.n25 VDD 0.169059
R228 VDD.n63 VDD 0.169059
R229 VDD VDD.n97 0.169059
R230 VDD VDD.n101 0.169059
R231 VDD.n101 VDD 0.153042
R232 VDD.n21 VDD.n14 0.145855
R233 VDD.n47 VDD.n46 0.145855
R234 VDD.n100 VDD.n99 0.145855
R235 VDD.n6 VDD.n1 0.145855
R236 VDD VDD.n29 0.145264
R237 VDD VDD.n48 0.145264
R238 VDD.n68 VDD 0.145264
R239 VDD VDD.n36 0.143594
R240 VDD.n35 VDD.n34 0.126615
R241 VDD.n43 VDD 0.103227
R242 VDD VDD.n57 0.103227
R243 VDD.n74 VDD 0.103227
R244 VDD.n86 VDD 0.103227
R245 VDD.n91 VDD 0.103227
R246 VDD.n15 VDD 0.0641126
R247 VDD.n18 VDD 0.0641126
R248 VDD.n2 VDD 0.0641126
R249 VDD VDD.n31 0.0578113
R250 VDD VDD.n50 0.0578113
R251 VDD VDD.n67 0.0578113
R252 VDD.n80 VDD 0.0578113
R253 VDD VDD.n24 0.0432119
R254 VDD VDD.n62 0.0432119
R255 VDD.n98 VDD 0.0432119
R256 VDD VDD.n9 0.0432119
R257 VDD.n37 VDD 0.036759
R258 VDD VDD.n15 0.0353691
R259 VDD.n17 VDD 0.0353691
R260 VDD VDD.n18 0.0353691
R261 VDD.n20 VDD 0.0353691
R262 VDD VDD.n21 0.0353691
R263 VDD VDD.n47 0.0353691
R264 VDD VDD.n100 0.0353691
R265 VDD VDD.n2 0.0353691
R266 VDD.n5 VDD 0.0353691
R267 VDD VDD.n6 0.0353691
R268 VDD.n31 VDD 0.0319151
R269 VDD VDD.n29 0.0319151
R270 VDD.n34 VDD 0.0319151
R271 VDD VDD.n27 0.0319151
R272 VDD.n50 VDD 0.0319151
R273 VDD VDD.n48 0.0319151
R274 VDD.n54 VDD 0.0319151
R275 VDD.n67 VDD 0.0319151
R276 VDD VDD.n68 0.0319151
R277 VDD VDD.n65 0.0319151
R278 VDD VDD.n80 0.0319151
R279 VDD.n82 VDD 0.0319151
R280 VDD VDD.n79 0.0319151
R281 VDD VDD.n77 0.0319151
R282 VDD VDD.n42 0.00140909
R283 VDD.n58 VDD 0.00140909
R284 VDD VDD.n73 0.00140909
R285 VDD VDD.n85 0.00140909
R286 VDD VDD.n90 0.00140909
R287 VSS.n75 VSS.t51 21242.4
R288 VSS.n105 VSS.t75 6110.29
R289 VSS.t45 VSS.n108 4862.48
R290 VSS.n57 VSS.n38 4789.2
R291 VSS.n8 VSS.t4 4388.35
R292 VSS.t51 VSS.n74 4212.86
R293 VSS.t33 VSS.n99 3914.16
R294 VSS.n74 VSS.t29 3831.86
R295 VSS.n106 VSS.n105 3549.15
R296 VSS.n107 VSS.n106 3541.76
R297 VSS.n108 VSS.n107 3504.83
R298 VSS.n4 VSS.t59 3503.36
R299 VSS.n7 VSS.n6 3319.89
R300 VSS.n96 VSS.t2 3172.99
R301 VSS.t67 VSS.n95 3088.27
R302 VSS.n59 VSS.n58 3049.28
R303 VSS.n12 VSS.t6 3005.52
R304 VSS.n85 VSS.t22 2863.86
R305 VSS.n44 VSS.n43 2779.1
R306 VSS.n72 VSS.n71 2715.2
R307 VSS.n13 VSS.t35 2649.77
R308 VSS.n73 VSS.t69 2616.97
R309 VSS.n36 VSS.t57 2520.79
R310 VSS.n60 VSS.n59 2449.11
R311 VSS.n107 VSS.t14 2401.02
R312 VSS.n105 VSS.t27 2381.58
R313 VSS.t81 VSS.n24 2167.12
R314 VSS VSS.n13 2124.07
R315 VSS.t78 VSS.n63 1892.57
R316 VSS.n61 VSS.t80 1601.74
R317 VSS.t8 VSS.n7 1590.05
R318 VSS.n87 VSS.n86 1563.87
R319 VSS.n104 VSS.t35 1537.16
R320 VSS.n11 VSS.t4 1537.16
R321 VSS.t75 VSS.n104 1420.05
R322 VSS.t6 VSS.n11 1420.05
R323 VSS.n50 VSS.t49 1401.69
R324 VSS.n33 VSS.t24 1396.81
R325 VSS.n25 VSS.t81 1392.86
R326 VSS.n108 VSS.t37 1387.95
R327 VSS.n20 VSS.t39 1382.98
R328 VSS.n100 VSS.t33 1381.58
R329 VSS.n109 VSS.t45 1377.12
R330 VSS VSS.n24 1371.4
R331 VSS.n35 VSS.n34 1344.92
R332 VSS.n88 VSS.t77 1344.83
R333 VSS.n106 VSS.t20 1331.64
R334 VSS.n65 VSS.t50 1331.33
R335 VSS.n88 VSS.t20 1318.46
R336 VSS.n56 VSS 1305.2
R337 VSS.n25 VSS.t14 1286.73
R338 VSS.n100 VSS.t27 1276.32
R339 VSS.t53 VSS.n44 1250.59
R340 VSS.t71 VSS.n39 1189.96
R341 VSS.n84 VSS.t41 1154.82
R342 VSS.n62 VSS.n1 1117.8
R343 VSS.t22 VSS.n84 1066.84
R344 VSS.t73 VSS.n78 968.886
R345 VSS.n76 VSS.t10 943.018
R346 VSS.n33 VSS.n32 896.351
R347 VSS.n64 VSS.t78 835.341
R348 VSS.n85 VSS.t55 691.832
R349 VSS.n61 VSS.t61 683.788
R350 VSS.n34 VSS.t12 664.105
R351 VSS.n23 VSS.t63 603.342
R352 VSS.n70 VSS.n60 561.245
R353 VSS.n58 VSS.n57 524.581
R354 VSS.t31 VSS.n75 470.334
R355 VSS.n65 VSS.n64 469.88
R356 VSS.n80 VSS.n79 467.981
R357 VSS.n71 VSS.t0 465.135
R358 VSS.n12 VSS.t16 418.317
R359 VSS.n63 VSS.n62 391.567
R360 VSS.n62 VSS.n61 313.738
R361 VSS.n24 VSS.n23 218.083
R362 VSS.n56 VSS.n39 166.986
R363 VSS.n74 VSS.t25 147.327
R364 VSS.n86 VSS.n85 80.4465
R365 VSS.n13 VSS.n12 72.402
R366 VSS.n57 VSS.n56 60.938
R367 VSS.n51 VSS.n46 56.8118
R368 VSS.n32 VSS.n21 56.8118
R369 VSS.n89 VSS.n87 56.8118
R370 VSS.n110 VSS.n1 56.8118
R371 VSS.n69 VSS.n66 56.8118
R372 VSS.n58 VSS.t18 55.0191
R373 VSS.n4 VSS.t65 26.2102
R374 VSS.n6 VSS.t59 26.2102
R375 VSS.n8 VSS.t8 26.2102
R376 VSS.n43 VSS.t71 23.1596
R377 VSS.n45 VSS.t53 23.1596
R378 VSS.n95 VSS.t47 23.1048
R379 VSS.n96 VSS.t67 23.1048
R380 VSS.n99 VSS.t2 23.1048
R381 VSS.t29 VSS.n73 19.5788
R382 VSS.t69 VSS.n72 19.5788
R383 VSS.t0 VSS.n70 19.5788
R384 VSS.t51 VSS.n36 18.8593
R385 VSS.t57 VSS.n35 18.8593
R386 VSS.n40 VSS.t25 18.7505
R387 VSS.n38 VSS.t43 18.7505
R388 VSS.n93 VSS.t34 9.0005
R389 VSS.n101 VSS.t28 9.0005
R390 VSS.n82 VSS.t42 9.0005
R391 VSS.n83 VSS.t23 9.0005
R392 VSS.n10 VSS.t5 9.0005
R393 VSS.n2 VSS.t7 9.0005
R394 VSS.n15 VSS.t36 9.0005
R395 VSS.n103 VSS.t76 9.0005
R396 VSS.n27 VSS.t82 8.99388
R397 VSS.n26 VSS.t15 8.99388
R398 VSS.n41 VSS.t26 8.96939
R399 VSS.n42 VSS.t44 8.96939
R400 VSS.n55 VSS.t19 8.96939
R401 VSS.n54 VSS.t72 8.96939
R402 VSS.n53 VSS.t54 8.96939
R403 VSS.n94 VSS.t48 8.96939
R404 VSS.n97 VSS.t68 8.96939
R405 VSS.n98 VSS.t3 8.96939
R406 VSS.n77 VSS.t32 8.96939
R407 VSS.n18 VSS.t11 8.96939
R408 VSS.n81 VSS.t74 8.96939
R409 VSS.n17 VSS.t56 8.96939
R410 VSS.n112 VSS.t62 8.96939
R411 VSS.n5 VSS.t66 8.96939
R412 VSS.n3 VSS.t60 8.96939
R413 VSS.n9 VSS.t9 8.96939
R414 VSS.n14 VSS.t17 8.96939
R415 VSS.n37 VSS.t30 8.96939
R416 VSS.n67 VSS.t70 8.96939
R417 VSS.n68 VSS.t1 8.96939
R418 VSS.n19 VSS.t52 8.96383
R419 VSS.n22 VSS.t58 8.96383
R420 VSS.n31 VSS.t13 8.96383
R421 VSS.n28 VSS.t64 8.96383
R422 VSS.n76 VSS.t31 7.05549
R423 VSS.n78 VSS.t10 7.05549
R424 VSS.n80 VSS.t73 7.05549
R425 VSS.n49 VSS.t38 6.71411
R426 VSS.n29 VSS.t40 6.71411
R427 VSS.n91 VSS.t21 6.71411
R428 VSS.n47 VSS.t46 6.71411
R429 VSS.n113 VSS.t79 6.71411
R430 VSS VSS.n40 5.2005
R431 VSS VSS.n38 5.2005
R432 VSS VSS.n43 5.2005
R433 VSS.n36 VSS 5.2005
R434 VSS.n35 VSS 5.2005
R435 VSS VSS.n25 5.2005
R436 VSS.n84 VSS 5.2005
R437 VSS.n95 VSS 5.2005
R438 VSS VSS.n96 5.2005
R439 VSS.n99 VSS 5.2005
R440 VSS VSS.n100 5.2005
R441 VSS.n104 VSS 5.2005
R442 VSS.n11 VSS 5.2005
R443 VSS VSS.n4 5.2005
R444 VSS.n6 VSS 5.2005
R445 VSS VSS.n8 5.2005
R446 VSS VSS.n76 5.2005
R447 VSS.n78 VSS 5.2005
R448 VSS VSS.n80 5.2005
R449 VSS.n72 VSS 5.2005
R450 VSS.n73 VSS 5.2005
R451 VSS.n103 VSS.n102 4.22722
R452 VSS.n48 VSS.n47 4.19767
R453 VSS.n26 VSS.n16 2.81165
R454 VSS.n102 VSS.n101 2.77598
R455 VSS.n49 VSS.n48 2.64103
R456 VSS.n92 VSS.n91 2.63174
R457 VSS VSS.n46 2.6005
R458 VSS.n46 VSS.n45 2.6005
R459 VSS.n52 VSS.n51 2.6005
R460 VSS.n51 VSS.n50 2.6005
R461 VSS.n32 VSS 2.6005
R462 VSS.n30 VSS.n21 2.6005
R463 VSS.n21 VSS.n20 2.6005
R464 VSS.n90 VSS.n89 2.6005
R465 VSS.n89 VSS.n88 2.6005
R466 VSS.n87 VSS 2.6005
R467 VSS VSS.n1 2.6005
R468 VSS.n111 VSS.n110 2.6005
R469 VSS.n110 VSS.n109 2.6005
R470 VSS.n69 VSS 2.6005
R471 VSS.n70 VSS.n69 2.6005
R472 VSS.n66 VSS.n0 2.6005
R473 VSS.n66 VSS.n65 2.6005
R474 VSS.n102 VSS.n92 1.56038
R475 VSS.n48 VSS.n16 1.50617
R476 VSS.n92 VSS.n16 1.48074
R477 VSS VSS.n42 0.511827
R478 VSS.n98 VSS.n93 0.445721
R479 VSS.n82 VSS.n81 0.445721
R480 VSS.n10 VSS.n9 0.445721
R481 VSS.n15 VSS.n14 0.445721
R482 VSS.n28 VSS.n27 0.426856
R483 VSS.n83 VSS 0.42093
R484 VSS VSS.n2 0.417049
R485 VSS.n53 VSS.n52 0.400161
R486 VSS.n112 VSS.n111 0.400161
R487 VSS.n68 VSS.n0 0.400161
R488 VSS.n31 VSS.n30 0.396347
R489 VSS VSS.n3 0.382004
R490 VSS.n54 VSS 0.350146
R491 VSS.n90 VSS.n17 0.339273
R492 VSS.n34 VSS.n33 0.333763
R493 VSS VSS.n67 0.325456
R494 VSS.n29 VSS 0.311686
R495 VSS VSS.n97 0.262535
R496 VSS VSS.n18 0.262535
R497 VSS VSS.n22 0.251432
R498 VSS.n101 VSS 0.221916
R499 VSS VSS.n83 0.221916
R500 VSS VSS.n2 0.221916
R501 VSS VSS.n103 0.221916
R502 VSS VSS.n26 0.212534
R503 VSS VSS.n49 0.200331
R504 VSS VSS.n29 0.200331
R505 VSS.n47 VSS 0.200331
R506 VSS VSS.n113 0.200331
R507 VSS.n91 VSS 0.17014
R508 VSS.n113 VSS 0.157619
R509 VSS VSS.n93 0.100854
R510 VSS VSS.n82 0.100854
R511 VSS VSS.n10 0.100854
R512 VSS VSS.n15 0.100854
R513 VSS.n27 VSS 0.0966017
R514 VSS VSS.n41 0.0936858
R515 VSS.n55 VSS 0.0936858
R516 VSS.n94 VSS 0.0936858
R517 VSS VSS.n77 0.0936858
R518 VSS VSS.n5 0.0936858
R519 VSS VSS.n37 0.0936858
R520 VSS VSS.n19 0.0897373
R521 VSS.n41 VSS 0.0689956
R522 VSS.n42 VSS 0.0689956
R523 VSS VSS.n55 0.0689956
R524 VSS VSS.n54 0.0689956
R525 VSS VSS.n53 0.0689956
R526 VSS VSS.n94 0.0689956
R527 VSS.n97 VSS 0.0689956
R528 VSS VSS.n98 0.0689956
R529 VSS.n77 VSS 0.0689956
R530 VSS VSS.n18 0.0689956
R531 VSS.n81 VSS 0.0689956
R532 VSS VSS.n112 0.0689956
R533 VSS.n5 VSS 0.0689956
R534 VSS VSS.n3 0.0689956
R535 VSS.n9 VSS 0.0689956
R536 VSS.n14 VSS 0.0689956
R537 VSS.n37 VSS 0.0689956
R538 VSS.n67 VSS 0.0689956
R539 VSS VSS.n68 0.0689956
R540 VSS.n19 VSS 0.0660932
R541 VSS.n22 VSS 0.0660932
R542 VSS VSS.n31 0.0660932
R543 VSS VSS.n28 0.0660932
R544 VSS VSS.n17 0.0582612
R545 VSS.n52 VSS 0.0142288
R546 VSS.n30 VSS 0.0142288
R547 VSS.n111 VSS 0.0142288
R548 VSS VSS.n0 0.0142288
R549 VSS VSS.n90 0.0121547
R550 D2.n3 D2.n2 9.02722
R551 D2.n3 D2.n1 6.48941
R552 D2 D2.n0 2.25262
R553 D2 D2.n3 0.130713
R554 B3.t9 B3.t5 46.118
R555 B3.t6 B3.t3 44.4957
R556 B3 B3.n5 33.3896
R557 B3.n0 B3.t8 31.938
R558 B3.n1 B3.n0 31.598
R559 B3.n5 B3.t2 31.5469
R560 B3.n4 B3.t9 30.0142
R561 B3.n6 B3.t0 27.2239
R562 B3.n6 B3.t6 15.0244
R563 B3.n7 B3 13.5904
R564 B3.n5 B3.t7 12.6451
R565 B3.n4 B3.t4 12.341
R566 B3.n0 B3.t1 12.2541
R567 B3 B3.n6 5.30993
R568 B3.n3 B3.n1 4.77938
R569 B3 B3.n4 4.51075
R570 B3 B3.n8 3.35445
R571 B3.n8 B3 2.95504
R572 B3.n7 B3 2.9154
R573 B3.n3 B3.n2 2.26266
R574 B3.n8 B3.n7 1.42038
R575 B3 B3.n3 0.0126622
R576 B3.n1 B3 0.0067069
R577 B2.t12 B2.t8 46.118
R578 B2.t11 B2.t4 46.118
R579 B2.t6 B2.t2 44.4957
R580 B2 B2.n1 33.3896
R581 B2 B2.n0 33.3896
R582 B2 B2.n3 32.7242
R583 B2.n3 B2.t1 31.938
R584 B2.n1 B2.t5 31.5469
R585 B2.n0 B2.t0 31.5469
R586 B2.n4 B2.t12 30.0142
R587 B2.n5 B2.t11 30.0142
R588 B2.n2 B2.t13 27.2239
R589 B2.n2 B2.t6 15.0244
R590 B2.n1 B2.t10 12.6451
R591 B2.n0 B2.t9 12.6451
R592 B2.n4 B2.t7 12.341
R593 B2.n5 B2.t3 12.341
R594 B2.n3 B2.t14 12.2541
R595 B2 B2.n2 5.30993
R596 B2.n6 B2 4.75471
R597 B2 B2.n9 4.60259
R598 B2 B2.n4 4.51075
R599 B2 B2.n5 4.51075
R600 B2.n6 B2 3.24079
R601 B2.n8 B2 3.22985
R602 B2.n9 B2 3.2092
R603 B2.n7 B2 3.01142
R604 B2.n7 B2.n6 1.81841
R605 B2.n8 B2.n7 1.41293
R606 B2.n9 B2.n8 1.34865
R607 D4.n2 D4.n1 9.02722
R608 D4.n2 D4.n0 6.48941
R609 D4 D4.n2 0.130713
R610 D5.n2 D5.n1 9.02722
R611 D5.n2 D5.n0 6.48941
R612 D5 D5.n2 0.130713
R613 D3.n2 D3.n1 9.02722
R614 D3.n2 D3.n0 6.48941
R615 D3 D3.n2 0.130713
R616 D7.n2 D7.n1 9.02722
R617 D7.n2 D7.n0 6.48941
R618 D7 D7.n2 0.130713
R619 D6.n2 D6.n1 9.02722
R620 D6.n2 D6.n0 6.48941
R621 D6 D6.n2 0.130713
R622 D1.n2 D1.n1 9.02722
R623 D1.n2 D1.n0 6.48941
R624 D1 D1.n2 0.130713
C0 AND_0.B AND_1.Inverter_0.IN 0.114f
C1 B3 OR_2.OUT 0.00185f
C2 a_268_n1326# B2 0.166f
C3 OR_0.Inverter_0.IN B3 0.039f
C4 VDD OR_1.B 0.414f
C5 AND_1.Inverter_0.IN B2 0.124f
C6 a_268_n3244# VDD 0.893f
C7 INV_BUFF_2.Inverter_0.IN D3 0.114f
C8 OR_4.Inverter_0.IN B3 0.0848f
C9 AND_0.B INV_BUFF_0.Inverter_0.IN 2.46e-20
C10 VDD a_1881_n1685# 0.00253f
C11 a_268_n2622# VDD 0.00253f
C12 AND_4.Inverter_0.IN a_1557_n2284# 7.88e-20
C13 B3 a_268_215# 0.0154f
C14 a_268_n4206# B3 0.166f
C15 OR_1.Inverter_0.IN B1 0.261f
C16 VDD AND_2.Inverter_0.IN 0.581f
C17 INV_BUFF_2.Inverter_0.IN INV_BUFF_4.Inverter_0.IN 0.00203f
C18 OR_1.OUT INV_BUFF_4.Inverter_0.IN 0.126f
C19 B1 AND_2.OUT 0.0414f
C20 INV_BUFF_4.Inverter_0.IN OR_3.OUT 2.1e-19
C21 AND_0.B B3 0.168f
C22 B1 AND_0.OUT 4.92e-19
C23 a_268_n1326# AND_2.Inverter_0.IN 0.00344f
C24 INV_BUFF_5.Inverter_0.IN a_1557_n2284# 7.49e-19
C25 OR_1.Inverter_0.IN AND_3.Inverter_0.IN 0.00203f
C26 AND_1.Inverter_0.IN AND_2.Inverter_0.IN 0.00218f
C27 D3 AND_3.B 1.39e-20
C28 VDD a_268_n1326# 0.888f
C29 B1 AND_0.Inverter_0.IN 0.00652f
C30 B3 B2 2.98f
C31 B3 INV_BUFF_1.Inverter_0.IN 3.27e-21
C32 VDD AND_1.Inverter_0.IN 0.58f
C33 VDD OR_3.B 0.393f
C34 D3 D5 0.00346f
C35 VDD AND_3.OUT 0.417f
C36 OR_3.Inverter_0.IN OR_3.OUT 0.125f
C37 B1 OR_2.Inverter_0.IN 0.261f
C38 a_1840_n4206# OR_4.Inverter_0.IN 1.21e-19
C39 D7 VDD 0.123f
C40 INV_BUFF_2.Inverter_0.IN B1 1.19e-19
C41 D6 VDD 0.133f
C42 OR_1.OUT B1 2.74e-19
C43 B3 OR_1.B 0.00122f
C44 a_1840_n4206# a_268_n4206# 0.00394f
C45 a_268_n3244# B3 0.00418f
C46 INV_BUFF_4.Inverter_0.IN D5 0.114f
C47 B1 D4 1.31e-19
C48 VDD INV_BUFF_0.Inverter_0.IN 0.406f
C49 AND_0.OUT INV_BUFF_3.Inverter_0.IN 1.55e-19
C50 OR_1.Inverter_0.IN a_1557_n2284# 0.162f
C51 a_268_n2622# B3 0.155f
C52 B1 D2 0.252f
C53 OR_1.Inverter_0.IN AND_4.Inverter_0.IN 1.3e-19
C54 B3 AND_2.Inverter_0.IN 2.4e-19
C55 a_1557_n2284# AND_2.OUT 8.01e-21
C56 AND_0.Inverter_0.IN a_1628_215# 0.0608f
C57 VDD B3 1.87f
C58 B1 AND_3.B 0.184f
C59 INV_BUFF_2.Inverter_0.IN INV_BUFF_3.Inverter_0.IN 4.65e-20
C60 B1 OR_2.OUT 2.02e-19
C61 OR_3.Inverter_0.IN OR_4.Inverter_0.IN 3.8e-19
C62 D1 D2 0.00125f
C63 AND_3.Inverter_0.IN D2 0.00288f
C64 INV_BUFF_3.Inverter_0.IN D4 0.115f
C65 B1 OR_0.Inverter_0.IN 0.0875f
C66 OR_1.Inverter_0.IN INV_BUFF_5.Inverter_0.IN 4.57e-19
C67 B3 a_268_n1326# 0.0199f
C68 B1 D5 2.19e-20
C69 a_268_n724# B2 0.155f
C70 AND_1.Inverter_0.IN B3 0.0951f
C71 B3 OR_3.B 0.478f
C72 AND_3.B AND_3.Inverter_0.IN 0.129f
C73 B1 OR_4.Inverter_0.IN 0.258f
C74 INV_BUFF_3.Inverter_0.IN D2 0.0904f
C75 AND_4.Inverter_0.IN OR_2.Inverter_0.IN 4.83e-20
C76 B1 a_268_215# 0.00321f
C77 D7 B3 1.67e-20
C78 D6 B3 4.29e-19
C79 OR_0.Inverter_0.IN AND_3.Inverter_0.IN 9.03e-19
C80 B1 a_268_n4206# 0.164f
C81 B3 INV_BUFF_0.Inverter_0.IN 1.08e-19
C82 a_1557_n2284# D2 1.17e-19
C83 a_1840_n4206# VDD 0.901f
C84 B1 AND_0.B 0.00684f
C85 D3 VDD 0.123f
C86 a_268_n724# AND_2.Inverter_0.IN 0.0608f
C87 AND_3.B a_1557_n2284# 0.00203f
C88 a_1557_n2284# OR_2.OUT 0.00116f
C89 B1 INV_BUFF_1.Inverter_0.IN 0.0438f
C90 B1 B2 3.72f
C91 INV_BUFF_6.Inverter_0.IN OR_3.OUT 0.12f
C92 AND_0.B D1 1.24e-20
C93 a_1840_n4206# OR_3.B 0.0242f
C94 VDD a_268_n724# 0.00253f
C95 AND_0.B AND_3.Inverter_0.IN 6.34e-21
C96 VDD INV_BUFF_4.Inverter_0.IN 0.403f
C97 B1 OR_1.B 0.369f
C98 OR_0.Inverter_0.IN AND_4.Inverter_0.IN 1.29e-19
C99 D6 a_1840_n4206# 0.00231f
C100 a_268_n724# a_268_n1326# 0.00272f
C101 INV_BUFF_1.Inverter_0.IN AND_3.Inverter_0.IN 1.75e-19
C102 a_268_n3244# B1 0.202f
C103 B2 AND_3.Inverter_0.IN 4.44e-22
C104 B1 a_1881_n1685# 0.00178f
C105 a_268_n2622# B1 0.0192f
C106 AND_0.B a_1628_215# 0.155f
C107 OR_3.Inverter_0.IN VDD 0.308f
C108 INV_BUFF_5.Inverter_0.IN OR_2.OUT 0.126f
C109 AND_0.Inverter_0.IN AND_0.OUT 0.123f
C110 OR_1.Inverter_0.IN OR_1.OUT 0.128f
C111 AND_4.Inverter_0.IN a_268_n4206# 5.09e-20
C112 B1 AND_2.Inverter_0.IN 0.0761f
C113 a_1628_215# INV_BUFF_1.Inverter_0.IN 9.25e-20
C114 a_1881_n1685# AND_3.Inverter_0.IN 0.0608f
C115 B1 VDD 6.04f
C116 a_1840_n4206# B3 0.173f
C117 OR_3.Inverter_0.IN OR_3.B 0.044f
C118 OR_1.Inverter_0.IN D2 1.45e-19
C119 a_1557_n2284# B2 5.15e-20
C120 a_1557_n2284# INV_BUFF_1.Inverter_0.IN 5.66e-19
C121 B1 a_268_n1326# 0.19f
C122 D1 VDD 0.125f
C123 AND_4.Inverter_0.IN B2 0.0106f
C124 B1 OR_3.B 0.00152f
C125 VDD AND_3.Inverter_0.IN 0.587f
C126 B1 AND_1.Inverter_0.IN 0.0145f
C127 AND_2.OUT D2 6.79e-19
C128 B3 a_268_n724# 3.35e-19
C129 B1 AND_3.OUT 4.97e-19
C130 OR_1.Inverter_0.IN AND_3.B 2.75e-21
C131 AND_0.OUT D2 0.0036f
C132 OR_1.Inverter_0.IN OR_2.OUT 2.2e-19
C133 a_1557_n2284# OR_1.B 0.0242f
C134 D6 B1 1.71e-19
C135 AND_0.Inverter_0.IN D2 1.1e-19
C136 a_1557_n2284# a_1881_n1685# 0.00139f
C137 AND_4.Inverter_0.IN OR_1.B 0.12f
C138 AND_3.B AND_2.OUT 9.25e-20
C139 VDD INV_BUFF_3.Inverter_0.IN 0.405f
C140 a_268_n3244# AND_4.Inverter_0.IN 0.00236f
C141 INV_BUFF_2.Inverter_0.IN D4 8.69e-21
C142 AND_3.Inverter_0.IN AND_3.OUT 0.125f
C143 OR_1.OUT OR_3.OUT 8.94e-21
C144 VDD a_1628_215# 0.00253f
C145 OR_0.Inverter_0.IN AND_2.OUT 1.54e-19
C146 OR_3.Inverter_0.IN B3 0.261f
C147 a_268_n2622# AND_4.Inverter_0.IN 0.0608f
C148 AND_3.B AND_0.Inverter_0.IN 6.33e-21
C149 INV_BUFF_2.Inverter_0.IN D2 0.00112f
C150 OR_1.OUT D2 3.14e-20
C151 a_1557_n2284# VDD 0.91f
C152 D1 INV_BUFF_0.Inverter_0.IN 0.114f
C153 INV_BUFF_3.Inverter_0.IN AND_3.OUT 0.00147f
C154 AND_4.Inverter_0.IN AND_2.Inverter_0.IN 4.44e-19
C155 D2 D4 0.103f
C156 OR_2.Inverter_0.IN OR_2.OUT 0.128f
C157 AND_1.Inverter_0.IN a_1628_215# 1.61e-19
C158 B1 B3 0.657f
C159 INV_BUFF_2.Inverter_0.IN AND_3.B 2.9e-20
C160 AND_4.Inverter_0.IN VDD 0.586f
C161 OR_0.Inverter_0.IN OR_2.Inverter_0.IN 4.37e-19
C162 INV_BUFF_0.Inverter_0.IN INV_BUFF_3.Inverter_0.IN 1.22e-19
C163 OR_4.Inverter_0.IN OR_2.Inverter_0.IN 0.00209f
C164 AND_4.Inverter_0.IN a_268_n1326# 1.15e-19
C165 AND_0.B AND_2.OUT 6.53e-20
C166 AND_0.B AND_0.OUT 2.17e-19
C167 INV_BUFF_6.Inverter_0.IN VDD 0.402f
C168 D5 OR_3.OUT 1.89e-21
C169 AND_3.B D2 6.27e-19
C170 a_268_n4206# OR_2.Inverter_0.IN 0.00198f
C171 INV_BUFF_5.Inverter_0.IN VDD 0.407f
C172 INV_BUFF_1.Inverter_0.IN AND_2.OUT 0.121f
C173 AND_0.B AND_0.Inverter_0.IN 0.129f
C174 B2 AND_2.OUT 2.17e-19
C175 a_1840_n4206# OR_3.Inverter_0.IN 0.162f
C176 OR_1.Inverter_0.IN OR_1.B 0.0438f
C177 B3 a_1628_215# 0.00106f
C178 INV_BUFF_5.Inverter_0.IN OR_3.B 8.18e-19
C179 OR_1.B AND_2.OUT 7.77e-19
C180 OR_0.Inverter_0.IN AND_3.B 0.117f
C181 a_1840_n4206# B1 7.2e-19
C182 INV_BUFF_6.Inverter_0.IN D7 0.115f
C183 B2 OR_2.Inverter_0.IN 0.0387f
C184 a_1557_n2284# B3 9.19e-20
C185 INV_BUFF_5.Inverter_0.IN D6 0.115f
C186 OR_1.Inverter_0.IN VDD 0.313f
C187 AND_4.Inverter_0.IN B3 0.125f
C188 B1 a_268_n724# 0.00491f
C189 AND_0.B D2 3.27e-21
C190 AND_2.Inverter_0.IN AND_2.OUT 0.122f
C191 OR_1.B OR_2.Inverter_0.IN 1.01e-19
C192 B1 INV_BUFF_4.Inverter_0.IN 4.5e-20
C193 a_268_n3244# OR_2.Inverter_0.IN 0.162f
C194 VDD AND_2.OUT 0.416f
C195 VDD AND_0.OUT 0.437f
C196 B2 D2 1.19e-20
C197 INV_BUFF_1.Inverter_0.IN D2 0.117f
C198 OR_1.Inverter_0.IN OR_3.B 4.09e-20
C199 INV_BUFF_6.Inverter_0.IN B3 3.34e-20
C200 a_268_n4206# OR_4.Inverter_0.IN 0.159f
C201 INV_BUFF_5.Inverter_0.IN B3 1.06e-19
C202 VDD AND_0.Inverter_0.IN 0.584f
C203 AND_3.B B2 1.41e-19
C204 AND_3.B INV_BUFF_1.Inverter_0.IN 8.2e-20
C205 VDD OR_2.Inverter_0.IN 0.318f
C206 OR_0.Inverter_0.IN B2 0.259f
C207 INV_BUFF_4.Inverter_0.IN INV_BUFF_3.Inverter_0.IN 5.17e-21
C208 INV_BUFF_2.Inverter_0.IN VDD 0.405f
C209 OR_1.OUT VDD 0.415f
C210 AND_1.Inverter_0.IN AND_0.Inverter_0.IN 8.39e-19
C211 AND_3.B OR_1.B 2.76e-19
C212 OR_1.B OR_2.OUT 5.47e-19
C213 OR_4.Inverter_0.IN B2 0.0387f
C214 VDD D4 0.133f
C215 VDD OR_3.OUT 0.41f
C216 INV_BUFF_0.Inverter_0.IN AND_0.OUT 0.122f
C217 AND_2.Inverter_0.IN D2 1.92e-19
C218 a_268_215# B2 0.156f
C219 OR_0.Inverter_0.IN OR_1.B 7.97e-20
C220 AND_3.B a_1881_n1685# 0.155f
C221 a_268_n4206# B2 0.0229f
C222 OR_1.Inverter_0.IN B3 6.96e-20
C223 VDD D2 0.332f
C224 B1 AND_3.Inverter_0.IN 0.0138f
C225 INV_BUFF_2.Inverter_0.IN AND_3.OUT 0.126f
C226 OR_1.OUT AND_3.OUT 0.00203f
C227 OR_0.Inverter_0.IN a_1881_n1685# 1.94e-19
C228 INV_BUFF_5.Inverter_0.IN a_1840_n4206# 0.0055f
C229 AND_0.B INV_BUFF_1.Inverter_0.IN 0.00218f
C230 AND_0.B B2 2.17e-19
C231 B3 AND_2.OUT 0.00192f
C232 AND_3.B VDD 0.386f
C233 B3 AND_0.OUT 3.44e-19
C234 OR_0.Inverter_0.IN AND_2.Inverter_0.IN 5.03e-20
C235 a_268_n3244# a_268_n4206# 0.0248f
C236 VDD OR_2.OUT 0.419f
C237 B1 INV_BUFF_3.Inverter_0.IN 0.109f
C238 AND_3.OUT D2 0.00246f
C239 B1 a_1628_215# 0.00237f
C240 B2 INV_BUFF_1.Inverter_0.IN 2.31e-20
C241 OR_0.Inverter_0.IN VDD 0.317f
C242 VDD D5 0.126f
C243 INV_BUFF_0.Inverter_0.IN D4 1.37e-19
C244 B3 AND_0.Inverter_0.IN 0.0112f
C245 AND_3.B a_268_n1326# 1.6e-20
C246 OR_4.Inverter_0.IN VDD 0.312f
C247 B3 OR_2.Inverter_0.IN 0.00513f
C248 OR_3.B OR_2.OUT 8.19e-19
C249 AND_3.B AND_3.OUT 2.17e-19
C250 B1 a_1557_n2284# 0.185f
C251 OR_0.Inverter_0.IN a_268_n1326# 0.159f
C252 INV_BUFF_0.Inverter_0.IN D2 0.00435f
C253 VDD a_268_215# 0.00253f
C254 OR_1.B B2 1.57e-20
C255 a_268_n3244# B2 0.0242f
C256 a_268_n4206# VDD 0.886f
C257 D6 AND_3.B 2.46e-21
C258 OR_1.Inverter_0.IN a_1840_n4206# 4.48e-19
C259 B1 AND_4.Inverter_0.IN 0.0912f
C260 a_1881_n1685# B2 1.37e-21
C261 INV_BUFF_5.Inverter_0.IN OR_3.Inverter_0.IN 7.18e-20
C262 a_1881_n1685# INV_BUFF_1.Inverter_0.IN 7.61e-20
C263 OR_4.Inverter_0.IN OR_3.B 0.123f
C264 B3 OR_3.OUT 2.91e-19
C265 a_268_n2622# B2 0.00118f
C266 a_1557_n2284# AND_3.Inverter_0.IN 5.89e-19
C267 AND_1.Inverter_0.IN a_268_215# 0.0608f
C268 AND_0.B VDD 0.382f
C269 B2 AND_2.Inverter_0.IN 0.126f
C270 a_268_n4206# OR_3.B 2.16e-19
C271 INV_BUFF_5.Inverter_0.IN B1 0.00153f
C272 a_268_n2622# OR_1.B 4.07e-20
C273 VDD INV_BUFF_1.Inverter_0.IN 0.408f
C274 VDD B2 2.1f
C275 a_268_n2622# a_268_n3244# 0.00223f
C276 D7 VSS 0.206f
C277 INV_BUFF_6.Inverter_0.IN VSS 0.408f
C278 OR_3.OUT VSS 0.461f
C279 OR_3.Inverter_0.IN VSS 0.749f
C280 a_1840_n4206# VSS 0.139f
C281 OR_4.Inverter_0.IN VSS 0.751f
C282 a_268_n4206# VSS 0.0696f
C283 OR_3.B VSS 0.594f
C284 D6 VSS 0.197f
C285 INV_BUFF_5.Inverter_0.IN VSS 0.399f
C286 OR_2.OUT VSS 0.38f
C287 OR_2.Inverter_0.IN VSS 0.747f
C288 a_268_n3244# VSS 0.0886f
C289 a_268_n2622# VSS 0.188f
C290 D5 VSS 0.193f
C291 INV_BUFF_4.Inverter_0.IN VSS 0.401f
C292 OR_1.OUT VSS 0.382f
C293 OR_1.Inverter_0.IN VSS 0.74f
C294 a_1557_n2284# VSS 0.122f
C295 AND_4.Inverter_0.IN VSS 0.4f
C296 OR_1.B VSS 0.602f
C297 a_1881_n1685# VSS 0.188f
C298 D3 VSS 0.195f
C299 INV_BUFF_2.Inverter_0.IN VSS 0.402f
C300 AND_3.OUT VSS 0.383f
C301 AND_3.Inverter_0.IN VSS 0.386f
C302 AND_3.B VSS 0.524f
C303 OR_0.Inverter_0.IN VSS 0.758f
C304 a_268_n1326# VSS 0.0641f
C305 a_268_n724# VSS 0.191f
C306 D4 VSS 0.171f
C307 D2 VSS 0.662f
C308 INV_BUFF_3.Inverter_0.IN VSS 0.404f
C309 INV_BUFF_1.Inverter_0.IN VSS 0.393f
C310 AND_2.OUT VSS 0.437f
C311 AND_2.Inverter_0.IN VSS 0.4f
C312 a_1628_215# VSS 0.188f
C313 D1 VSS 0.187f
C314 a_268_215# VSS 0.188f
C315 INV_BUFF_0.Inverter_0.IN VSS 0.403f
C316 AND_0.OUT VSS 0.401f
C317 AND_0.Inverter_0.IN VSS 0.393f
C318 AND_0.B VSS 0.566f
C319 B3 VSS 5.78f
C320 AND_1.Inverter_0.IN VSS 0.403f
C321 B2 VSS 6.78f
C322 B1 VSS 6.58f
C323 VDD VSS 50.1f
C324 B2.t0 VSS 0.0775f
C325 B2.t9 VSS 0.0332f
C326 B2.n0 VSS 0.153f
C327 B2.t5 VSS 0.0775f
C328 B2.t10 VSS 0.0332f
C329 B2.n1 VSS 0.153f
C330 B2.t2 VSS 0.0965f
C331 B2.t6 VSS 0.132f
C332 B2.t13 VSS 0.0543f
C333 B2.n2 VSS 0.257f
C334 B2.t14 VSS 0.0323f
C335 B2.t1 VSS 0.0784f
C336 B2.n3 VSS 0.146f
C337 B2.t8 VSS 0.0936f
C338 B2.t12 VSS 0.162f
C339 B2.t7 VSS 0.0224f
C340 B2.n4 VSS 0.21f
C341 B2.t4 VSS 0.0936f
C342 B2.t11 VSS 0.162f
C343 B2.t3 VSS 0.0224f
C344 B2.n5 VSS 0.21f
C345 B2.n6 VSS 0.993f
C346 B2.n7 VSS 0.693f
C347 B2.n8 VSS 0.606f
C348 B2.n9 VSS 0.856f
C349 B3.t1 VSS 0.0107f
C350 B3.t8 VSS 0.026f
C351 B3.n0 VSS 0.0473f
C352 B3.n1 VSS 0.143f
C353 B3.n2 VSS 0.0213f
C354 B3.n3 VSS 0.261f
C355 B3.t5 VSS 0.031f
C356 B3.t9 VSS 0.0537f
C357 B3.t4 VSS 0.00742f
C358 B3.n4 VSS 0.0696f
C359 B3.t2 VSS 0.0257f
C360 B3.t7 VSS 0.011f
C361 B3.n5 VSS 0.0509f
C362 B3.t3 VSS 0.032f
C363 B3.t6 VSS 0.0438f
C364 B3.t0 VSS 0.018f
C365 B3.n6 VSS 0.0853f
C366 B3.n7 VSS 0.664f
C367 B3.n8 VSS 0.323f
C368 VDD.n0 VSS 0.0031f
C369 VDD.n1 VSS 0.0238f
C370 VDD.t0 VSS 0.0561f
C371 VDD.t97 VSS 0.003f
C372 VDD.t46 VSS 0.0485f
C373 VDD.t47 VSS 0.003f
C374 VDD.n2 VSS 0.0196f
C375 VDD.n3 VSS 0.0517f
C376 VDD.t96 VSS 0.0461f
C377 VDD.n4 VSS 0.0615f
C378 VDD.n5 VSS 0.0345f
C379 VDD.t1 VSS 0.003f
C380 VDD.n6 VSS 0.0246f
C381 VDD.n7 VSS 0.0518f
C382 VDD.t66 VSS 0.0754f
C383 VDD.t91 VSS 0.0767f
C384 VDD.n8 VSS 0.0685f
C385 VDD.n9 VSS 0.0281f
C386 VDD.t92 VSS 0.0031f
C387 VDD.t83 VSS 0.0428f
C388 VDD.n10 VSS 0.0455f
C389 VDD.t84 VSS 0.003f
C390 VDD.n11 VSS 0.0031f
C391 VDD.t4 VSS 0.0522f
C392 VDD.t52 VSS 0.0767f
C393 VDD.n12 VSS 0.0685f
C394 VDD.t53 VSS 0.0031f
C395 VDD.t55 VSS 0.0031f
C396 VDD.n13 VSS 0.0031f
C397 VDD.n14 VSS 0.0238f
C398 VDD.t102 VSS 0.003f
C399 VDD.t27 VSS 0.0485f
C400 VDD.t51 VSS 0.003f
C401 VDD.t42 VSS 0.0485f
C402 VDD.t43 VSS 0.003f
C403 VDD.n15 VSS 0.0196f
C404 VDD.n16 VSS 0.0517f
C405 VDD.t50 VSS 0.0528f
C406 VDD.n17 VSS 0.0341f
C407 VDD.t28 VSS 0.003f
C408 VDD.n18 VSS 0.0196f
C409 VDD.n19 VSS 0.0517f
C410 VDD.t101 VSS 0.0528f
C411 VDD.n20 VSS 0.0361f
C412 VDD.t76 VSS 0.003f
C413 VDD.n21 VSS 0.0246f
C414 VDD.t75 VSS 0.0428f
C415 VDD.n22 VSS 0.0455f
C416 VDD.t69 VSS 0.0522f
C417 VDD.t54 VSS 0.0767f
C418 VDD.n23 VSS 0.0685f
C419 VDD.n24 VSS 0.0281f
C420 VDD.n25 VSS 0.0432f
C421 VDD.t8 VSS 0.00314f
C422 VDD.n26 VSS 0.00314f
C423 VDD.t86 VSS 0.003f
C424 VDD.n27 VSS 0.0395f
C425 VDD.t85 VSS 0.0641f
C426 VDD.t38 VSS 0.0754f
C427 VDD.n28 VSS 0.0031f
C428 VDD.t20 VSS 0.003f
C429 VDD.t80 VSS 0.003f
C430 VDD.n29 VSS 0.0328f
C431 VDD.t79 VSS 0.0461f
C432 VDD.t73 VSS 0.003f
C433 VDD.t72 VSS 0.0485f
C434 VDD.n30 VSS 0.0517f
C435 VDD.n31 VSS 0.0208f
C436 VDD.n32 VSS 0.0529f
C437 VDD.t19 VSS 0.0473f
C438 VDD.n33 VSS 0.0518f
C439 VDD.n34 VSS 0.0264f
C440 VDD.n35 VSS 0.0268f
C441 VDD.t61 VSS 0.0031f
C442 VDD.n36 VSS 0.0304f
C443 VDD.n37 VSS 0.03f
C444 VDD.n38 VSS 0.0685f
C445 VDD.t60 VSS 0.0403f
C446 VDD.n39 VSS 0.0318f
C447 VDD.n40 VSS 0.0428f
C448 VDD.t74 VSS 0.0463f
C449 VDD.t41 VSS 0.0473f
C450 VDD.t7 VSS 0.0721f
C451 VDD.t22 VSS 0.0452f
C452 VDD.n41 VSS 0.0736f
C453 VDD.n42 VSS 0.0393f
C454 VDD.n43 VSS 0.0193f
C455 VDD.n44 VSS 0.0439f
C456 VDD.t37 VSS 0.0031f
C457 VDD.n45 VSS 0.0031f
C458 VDD.n46 VSS 0.0238f
C459 VDD.t78 VSS 0.003f
C460 VDD.n47 VSS 0.0246f
C461 VDD.t77 VSS 0.0422f
C462 VDD.t57 VSS 0.0473f
C463 VDD.t104 VSS 0.003f
C464 VDD.t18 VSS 0.003f
C465 VDD.n48 VSS 0.0328f
C466 VDD.t62 VSS 0.0463f
C467 VDD.t17 VSS 0.0461f
C468 VDD.t49 VSS 0.003f
C469 VDD.t48 VSS 0.0485f
C470 VDD.n49 VSS 0.0517f
C471 VDD.n50 VSS 0.0208f
C472 VDD.n51 VSS 0.0301f
C473 VDD.t103 VSS 0.041f
C474 VDD.n52 VSS 0.0334f
C475 VDD.n53 VSS 0.0433f
C476 VDD.n54 VSS 0.0395f
C477 VDD.n55 VSS 0.00314f
C478 VDD.t35 VSS 0.00314f
C479 VDD.n56 VSS 0.0278f
C480 VDD.n57 VSS 0.0193f
C481 VDD.n58 VSS 0.0393f
C482 VDD.n59 VSS 0.0736f
C483 VDD.t31 VSS 0.0452f
C484 VDD.t34 VSS 0.0562f
C485 VDD.n60 VSS 0.0817f
C486 VDD.t93 VSS 0.0522f
C487 VDD.t36 VSS 0.0767f
C488 VDD.n61 VSS 0.0685f
C489 VDD.n62 VSS 0.0281f
C490 VDD.n63 VSS 0.0433f
C491 VDD.t30 VSS 0.00314f
C492 VDD.n64 VSS 0.00314f
C493 VDD.t3 VSS 0.003f
C494 VDD.n65 VSS 0.0395f
C495 VDD.t2 VSS 0.0424f
C496 VDD.t89 VSS 0.0461f
C497 VDD.t65 VSS 0.003f
C498 VDD.t64 VSS 0.0485f
C499 VDD.n66 VSS 0.0517f
C500 VDD.n67 VSS 0.0208f
C501 VDD.t90 VSS 0.003f
C502 VDD.n68 VSS 0.0328f
C503 VDD.n69 VSS 0.0303f
C504 VDD.n70 VSS 0.0339f
C505 VDD.n71 VSS 0.0446f
C506 VDD.t59 VSS 0.0463f
C507 VDD.t56 VSS 0.0473f
C508 VDD.t29 VSS 0.0721f
C509 VDD.t105 VSS 0.0452f
C510 VDD.n72 VSS 0.0736f
C511 VDD.n73 VSS 0.0393f
C512 VDD.n74 VSS 0.0193f
C513 VDD.n75 VSS 0.0447f
C514 VDD.t45 VSS 0.00314f
C515 VDD.n76 VSS 0.00314f
C516 VDD.t26 VSS 0.003f
C517 VDD.n77 VSS 0.0395f
C518 VDD.t25 VSS 0.0685f
C519 VDD.t11 VSS 0.00314f
C520 VDD.n78 VSS 0.00314f
C521 VDD.t16 VSS 0.003f
C522 VDD.n79 VSS 0.0395f
C523 VDD.t15 VSS 0.0634f
C524 VDD.t82 VSS 0.003f
C525 VDD.t87 VSS 0.0485f
C526 VDD.t88 VSS 0.003f
C527 VDD.n80 VSS 0.0208f
C528 VDD.n81 VSS 0.0517f
C529 VDD.t81 VSS 0.0528f
C530 VDD.n82 VSS 0.0374f
C531 VDD.n83 VSS 0.0584f
C532 VDD.t21 VSS 0.0699f
C533 VDD.t9 VSS 0.0473f
C534 VDD.t10 VSS 0.0772f
C535 VDD.t12 VSS 0.0452f
C536 VDD.n84 VSS 0.0736f
C537 VDD.n85 VSS 0.0393f
C538 VDD.n86 VSS 0.0193f
C539 VDD.n87 VSS 0.0273f
C540 VDD.n88 VSS 0.0584f
C541 VDD.t63 VSS 0.0699f
C542 VDD.t58 VSS 0.0473f
C543 VDD.t44 VSS 0.0721f
C544 VDD.t98 VSS 0.0452f
C545 VDD.n89 VSS 0.0736f
C546 VDD.n90 VSS 0.0393f
C547 VDD.n91 VSS 0.0193f
C548 VDD.n92 VSS 0.0509f
C549 VDD.n93 VSS 0.0547f
C550 VDD.n94 VSS 0.0359f
C551 VDD.n95 VSS 0.0362f
C552 VDD.n96 VSS 0.051f
C553 VDD.n97 VSS 0.0495f
C554 VDD.n98 VSS 0.0281f
C555 VDD.n99 VSS 0.0238f
C556 VDD.n100 VSS 0.0246f
C557 VDD.n101 VSS 0.0207f
C558 B1.t13 VSS 0.022f
C559 B1.t2 VSS 0.0534f
C560 B1.n0 VSS 0.0995f
C561 B1.t9 VSS 0.022f
C562 B1.t12 VSS 0.0534f
C563 B1.n1 VSS 0.0887f
C564 B1.n2 VSS 0.0646f
C565 B1.n3 VSS 0.011f
C566 B1.t14 VSS 0.0325f
C567 B1.t7 VSS 0.0244f
C568 B1.n4 VSS 0.113f
C569 B1.n5 VSS 0.928f
C570 B1.t3 VSS 0.022f
C571 B1.t11 VSS 0.0534f
C572 B1.n6 VSS 0.0973f
C573 B1.n7 VSS 0.718f
C574 B1.t1 VSS 0.0657f
C575 B1.t6 VSS 0.0901f
C576 B1.t10 VSS 0.037f
C577 B1.n8 VSS 0.174f
C578 B1.n9 VSS 0.849f
C579 B1.t4 VSS 0.0657f
C580 B1.t8 VSS 0.0901f
C581 B1.t16 VSS 0.037f
C582 B1.n10 VSS 0.175f
C583 B1.t0 VSS 0.0657f
C584 B1.t5 VSS 0.0901f
C585 B1.t15 VSS 0.037f
C586 B1.n11 VSS 0.175f
C587 B1.n12 VSS 0.619f
C588 B1.n13 VSS 0.941f
C589 B1.n14 VSS 0.98f
C590 B1.n15 VSS 0.613f
.ends

