magic
tech gf180mcuC
magscale 1 10
timestamp 1694155832
<< metal1 >>
rect 659 1268 830 1465
rect 1227 1363 1460 1379
rect 1227 1343 1243 1363
rect 899 1302 1243 1343
rect 1304 1362 1460 1363
rect 1304 1302 1385 1362
rect 899 1301 1385 1302
rect 1446 1343 1460 1362
rect 1446 1301 1785 1343
rect 899 1274 1785 1301
rect 1860 1276 2029 1460
rect 660 -280 831 -83
rect 905 -124 1791 -82
rect 905 -151 1262 -124
rect 1242 -185 1262 -151
rect 1323 -185 1403 -124
rect 1464 -151 1791 -124
rect 1464 -185 1482 -151
rect 1242 -197 1482 -185
rect 1860 -268 2029 -84
<< via1 >>
rect 1243 1302 1304 1363
rect 1385 1301 1446 1362
rect 1262 -185 1323 -124
rect 1403 -185 1464 -124
<< metal2 >>
rect 1247 1379 1445 1853
rect 1227 1363 1460 1379
rect 1227 1302 1243 1363
rect 1304 1362 1460 1363
rect 1304 1302 1385 1362
rect 1227 1301 1385 1302
rect 1446 1301 1460 1362
rect 1227 1294 1460 1301
rect 1254 -108 1452 -106
rect 1242 -124 1482 -108
rect 1242 -185 1262 -124
rect 1323 -185 1403 -124
rect 1464 -185 1482 -124
rect 1242 -197 1482 -185
rect 1254 -709 1452 -197
use ppolyf_u_WRMTN3  ppolyf_u_WRMTN3_0
timestamp 1694155832
transform 1 0 1348 0 1 592
box -864 -933 864 933
<< labels >>
flabel metal2 1331 -609 1331 -609 0 FreeSans 640 0 0 0 r2
port 2 nsew
flabel metal1 731 1455 731 1455 0 FreeSans 640 0 0 0 VDD
port 4 nsew
flabel metal2 1342 1740 1342 1740 0 FreeSans 640 0 0 0 r1
port 0 nsew
<< end >>
