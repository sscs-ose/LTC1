magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1201 1019 1201
<< metal1 >>
rect -19 195 19 201
rect -19 -195 -13 195
rect 13 -195 19 195
rect -19 -201 19 -195
<< via1 >>
rect -13 -195 13 195
<< metal2 >>
rect -19 195 19 201
rect -19 -195 -13 195
rect 13 -195 19 195
rect -19 -201 19 -195
<< end >>
