magic
tech gf180mcuC
magscale 1 10
timestamp 1699883071
<< nwell >>
rect 5835 3822 5911 3898
rect 2398 3450 2474 3526
rect 4178 3450 4254 3526
rect 6022 3450 6098 3526
rect 7142 -1430 7218 -1422
<< nsubdiff >>
rect 1810 3684 1858 3756
rect 3622 3684 3670 3756
rect 5434 3684 5482 3756
rect 7246 3684 7294 3756
rect -2387 -3645 -2339 -3572
rect 1810 -3644 1858 -3572
rect 3622 -3644 3670 -3572
rect 5434 -3644 5482 -3572
rect 7246 -3644 7294 -3572
<< polysilicon >>
rect 2398 3456 2474 3512
rect 4178 3456 4254 3512
rect 6022 3456 6098 3512
rect 7144 -1364 7216 -1356
rect 7144 -1369 7218 -1364
rect 7144 -1415 7157 -1369
rect 7203 -1415 7218 -1369
rect 7144 -1420 7218 -1415
rect 7144 -1428 7216 -1420
<< metal1 >>
rect -2 7682 9643 7767
rect -2 7680 170 7682
rect -2 7608 29 7680
rect 96 7610 170 7680
rect 237 7610 9643 7682
rect 96 7608 9643 7610
rect -2 7545 9643 7608
rect -2 7541 165 7545
rect -2 7469 32 7541
rect 99 7473 165 7541
rect 232 7473 9643 7545
rect 99 7469 9643 7473
rect -2 7402 9643 7469
rect 84 7328 9020 7402
rect 8922 7193 8998 7205
rect 6619 7120 6651 7167
rect 8922 7141 8934 7193
rect 8986 7141 8998 7193
rect 8922 7129 8998 7141
rect 6619 7093 6728 7120
rect 2991 7029 3089 7050
rect 1212 6976 1310 6997
rect 1212 6907 1230 6976
rect 1292 6907 1310 6976
rect 2991 6960 3009 7029
rect 3071 6960 3089 7029
rect 2991 6940 3089 6960
rect 4806 7018 4904 7039
rect 4806 6949 4824 7018
rect 4886 6949 4904 7018
rect 4806 6929 4904 6949
rect 6619 7024 6640 7093
rect 6702 7024 6728 7093
rect 6619 6971 6728 7024
rect 1212 6887 1310 6907
rect 6619 6902 6641 6971
rect 6703 6902 6728 6971
rect 2991 6820 3089 6841
rect 2991 6751 3009 6820
rect 3071 6751 3089 6820
rect 2991 6731 3089 6751
rect 4807 6830 4905 6851
rect 4807 6761 4825 6830
rect 4887 6761 4905 6830
rect 4807 6741 4905 6761
rect 6619 6849 6728 6902
rect 6619 6780 6641 6849
rect 6703 6780 6728 6849
rect 6619 6756 6728 6780
rect 4806 6649 4904 6670
rect 1215 6602 1313 6623
rect 1215 6533 1233 6602
rect 1295 6533 1313 6602
rect 1215 6513 1313 6533
rect 2995 6588 3093 6609
rect 2995 6519 3013 6588
rect 3075 6519 3093 6588
rect 4806 6580 4824 6649
rect 4886 6580 4904 6649
rect 4806 6560 4904 6580
rect 2995 6499 3093 6519
rect 1215 6269 1313 6290
rect 1215 6200 1233 6269
rect 1295 6200 1313 6269
rect 1215 6180 1313 6200
rect 1886 5962 1962 5974
rect 1886 5959 1898 5962
rect 1772 5913 1898 5959
rect 1886 5910 1898 5913
rect 1950 5910 1962 5962
rect 1886 5898 1962 5910
rect 3698 5962 3774 5974
rect 3698 5910 3710 5962
rect 3762 5910 3774 5962
rect 3698 5898 3774 5910
rect 5510 5962 5586 5974
rect 5510 5910 5522 5962
rect 5574 5910 5586 5962
rect 5510 5898 5586 5910
rect 7322 5963 7398 5975
rect 7322 5911 7334 5963
rect 7386 5911 7398 5963
rect 7322 5899 7398 5911
rect 7629 4426 7725 4443
rect 7629 4353 7646 4426
rect 7709 4353 7725 4426
rect 7629 4336 7725 4353
rect 8271 4430 8367 4447
rect 8271 4357 8288 4430
rect 8351 4357 8367 4430
rect 8271 4340 8367 4357
rect 7630 4179 7726 4196
rect -4878 3998 -301 4123
rect 7630 4106 7647 4179
rect 7710 4106 7726 4179
rect 7630 4089 7726 4106
rect 8271 4170 8367 4187
rect 8271 4097 8288 4170
rect 8351 4097 8367 4170
rect 8271 4080 8367 4097
rect -4878 3930 -4589 3998
rect -4519 3930 -4465 3998
rect -4395 3930 -4341 3998
rect -4271 3930 -4217 3998
rect -4147 3930 -301 3998
rect -4878 3874 -301 3930
rect -4878 3806 -4589 3874
rect -4519 3806 -4465 3874
rect -4395 3806 -4341 3874
rect -4271 3806 -4217 3874
rect -4147 3806 -301 3874
rect 1381 3886 1457 3898
rect 1381 3834 1393 3886
rect 1445 3834 1457 3886
rect 1381 3822 1457 3834
rect 2211 3886 2287 3898
rect 2211 3834 2223 3886
rect 2275 3834 2287 3886
rect 2211 3822 2287 3834
rect 4023 3886 4099 3898
rect 4023 3834 4035 3886
rect 4087 3834 4099 3886
rect 4023 3822 4099 3834
rect 5835 3886 5911 3898
rect 5835 3834 5847 3886
rect 5899 3834 5911 3886
rect 5835 3822 5911 3834
rect -4878 3776 -301 3806
rect -4878 3700 22 3776
rect -4603 3696 -4533 3700
rect -845 3664 22 3700
rect 1194 3514 1270 3526
rect 1194 3462 1206 3514
rect 1258 3462 1270 3514
rect 1194 3450 1270 3462
rect 2398 3514 2474 3526
rect 2398 3462 2410 3514
rect 2462 3462 2474 3514
rect 2398 3450 2474 3462
rect 4178 3514 4254 3526
rect 4178 3462 4190 3514
rect 4242 3462 4254 3514
rect 4178 3450 4254 3462
rect 6022 3514 6098 3526
rect 6022 3462 6034 3514
rect 6086 3462 6098 3514
rect 6022 3450 6098 3462
rect 7349 3514 7425 3526
rect 7349 3462 7361 3514
rect 7413 3462 7425 3514
rect 7349 3450 7425 3462
rect -5127 3156 -4839 3202
rect -59 2633 17 2645
rect -59 2630 -47 2633
rect -626 2584 -47 2630
rect -59 2581 -47 2584
rect 5 2581 17 2633
rect -59 2569 17 2581
rect -181 2450 -105 2462
rect -181 2447 -169 2450
rect -673 2401 -169 2447
rect -181 2398 -169 2401
rect -117 2398 -105 2450
rect -181 2386 -105 2398
rect 1674 1659 1750 1671
rect -303 1622 -227 1634
rect -303 1619 -291 1622
rect -649 1573 -291 1619
rect -303 1570 -291 1573
rect -239 1570 -227 1622
rect 1674 1607 1686 1659
rect 1738 1607 1750 1659
rect 1674 1595 1750 1607
rect -303 1558 -227 1570
rect -59 1530 17 1542
rect -59 1478 -47 1530
rect 5 1527 17 1530
rect 5 1481 81 1527
rect 5 1478 17 1481
rect 3589 1481 3700 1527
rect -59 1466 17 1478
rect 7824 1249 7920 1266
rect 7824 1176 7841 1249
rect 7904 1176 7920 1249
rect 7824 1159 7920 1176
rect -5127 818 -4842 864
rect 7820 850 7916 867
rect 7820 777 7837 850
rect 7900 777 7916 850
rect 7820 760 7916 777
rect -425 740 -349 752
rect -425 737 -413 740
rect -540 691 -413 737
rect -425 688 -413 691
rect -361 688 -349 740
rect -425 676 -349 688
rect 7824 477 7920 494
rect 7824 404 7841 477
rect 7904 404 7920 477
rect 7824 387 7920 404
rect 5298 299 5374 311
rect 5298 247 5310 299
rect 5362 247 5374 299
rect 5298 235 5374 247
rect 9180 152 9643 7402
rect 8893 112 9643 152
rect 84 0 9643 112
rect 8893 -29 9643 0
rect 554 -150 630 -138
rect 554 -202 566 -150
rect 618 -202 630 -150
rect 554 -214 630 -202
rect 3038 -150 3114 -138
rect 3038 -202 3050 -150
rect 3102 -202 3114 -150
rect 3038 -214 3114 -202
rect 4818 -150 4894 -138
rect 4818 -202 4830 -150
rect 4882 -202 4894 -150
rect 4818 -214 4894 -202
rect 6662 -150 6738 -138
rect 6662 -202 6674 -150
rect 6726 -202 6738 -150
rect 6662 -214 6738 -202
rect 7349 -150 7425 -138
rect 7349 -202 7361 -150
rect 7413 -202 7425 -150
rect 7349 -214 7425 -202
rect -5126 -264 -4839 -218
rect 7822 -329 7918 -312
rect 7822 -402 7839 -329
rect 7902 -402 7918 -329
rect 7822 -419 7918 -402
rect 7826 -707 7922 -690
rect 7826 -780 7843 -707
rect 7906 -780 7922 -707
rect 7826 -797 7922 -780
rect -547 -970 -471 -958
rect -547 -973 -535 -970
rect -728 -1019 -535 -973
rect -547 -1022 -535 -1019
rect -483 -1022 -471 -970
rect -547 -1034 -471 -1022
rect 7824 -1094 7920 -1077
rect 7824 -1167 7841 -1094
rect 7904 -1167 7920 -1094
rect 7824 -1184 7920 -1167
rect -4683 -1394 -4175 -1357
rect -4683 -1434 -3953 -1394
rect -4683 -1502 -4610 -1434
rect -4540 -1436 -3953 -1434
rect -3901 -1436 -3653 -1394
rect -3601 -1436 -3353 -1394
rect -3301 -1436 -3053 -1394
rect -3001 -1436 -2753 -1394
rect -1138 -1394 -865 -1354
rect 7146 -1366 7214 -1358
rect -2701 -1436 -865 -1394
rect 7146 -1369 7154 -1366
rect 3589 -1415 3702 -1369
rect 7142 -1415 7154 -1369
rect 7146 -1418 7154 -1415
rect 7206 -1418 7214 -1366
rect 7146 -1426 7214 -1418
rect -4540 -1502 -865 -1436
rect -4683 -1558 -865 -1502
rect -4683 -1626 -4610 -1558
rect -4540 -1626 -4486 -1558
rect -4416 -1626 -4362 -1558
rect -4292 -1626 -865 -1558
rect -4683 -1682 -865 -1626
rect -4683 -1750 -4610 -1682
rect -4540 -1750 -4486 -1682
rect -4416 -1750 -4362 -1682
rect -4292 -1750 -865 -1682
rect -4683 -1837 -865 -1750
rect 1918 -3365 1994 -3353
rect 1918 -3417 1930 -3365
rect 1982 -3403 1994 -3365
rect 5542 -3365 5618 -3353
rect 1982 -3417 2001 -3403
rect 1918 -3429 2001 -3417
rect 5542 -3417 5554 -3365
rect 5606 -3402 5618 -3365
rect 5606 -3417 5625 -3402
rect 5542 -3429 5625 -3417
rect 1965 -3476 2001 -3429
rect 5597 -3474 5625 -3429
rect -4175 -3582 9082 -3552
rect -4175 -3634 -3953 -3582
rect -3901 -3634 -3653 -3582
rect -3601 -3634 -3353 -3582
rect -3301 -3634 -3053 -3582
rect -3001 -3634 -2753 -3582
rect -2701 -3634 9082 -3582
rect -4175 -3664 9082 -3634
rect 5033 -3740 5131 -3733
rect -2495 -3773 -2228 -3745
rect -2495 -3836 -2449 -3773
rect -2385 -3774 -2228 -3773
rect -2385 -3836 -2323 -3774
rect -2495 -3837 -2323 -3836
rect -2259 -3837 -2228 -3774
rect 5024 -3749 5167 -3740
rect -1159 -3814 -1083 -3802
rect -2495 -3852 -2228 -3837
rect -1488 -3841 -1393 -3823
rect -1488 -3905 -1473 -3841
rect -1411 -3905 -1393 -3841
rect -1159 -3866 -1147 -3814
rect -1095 -3866 -1083 -3814
rect -1159 -3878 -1083 -3866
rect 4013 -3814 4089 -3802
rect 4013 -3866 4025 -3814
rect 4077 -3866 4089 -3814
rect 5024 -3812 5047 -3749
rect 5116 -3812 5167 -3749
rect 5024 -3819 5167 -3812
rect 5033 -3825 5131 -3819
rect 4013 -3878 4089 -3866
rect -1488 -3919 -1393 -3905
rect -2490 -4056 -2238 -3964
rect -2489 -4329 -2237 -4237
rect -2490 -5142 -2238 -5050
rect -2485 -5445 -2233 -5353
rect -679 -5798 -603 -5786
rect -679 -5850 -667 -5798
rect -615 -5850 -603 -5798
rect -679 -5862 -603 -5850
rect -303 -5798 -227 -5786
rect 3518 -5798 3594 -5786
rect 8954 -5798 9030 -5786
rect -303 -5850 -291 -5798
rect -239 -5801 -227 -5798
rect -239 -5847 81 -5801
rect -239 -5850 -227 -5847
rect 1674 -5823 1750 -5811
rect -303 -5862 -227 -5850
rect 1674 -5875 1686 -5823
rect 1738 -5875 1750 -5823
rect 1674 -5887 1750 -5875
rect 1918 -5823 1994 -5811
rect 1918 -5875 1930 -5823
rect 1982 -5875 1994 -5823
rect 3518 -5850 3530 -5798
rect 3582 -5801 3594 -5798
rect 3582 -5847 3700 -5801
rect 5298 -5823 5374 -5811
rect 3582 -5850 3594 -5847
rect 3518 -5862 3594 -5850
rect 1918 -5887 1994 -5875
rect 5298 -5875 5310 -5823
rect 5362 -5875 5374 -5823
rect 5298 -5887 5374 -5875
rect 5542 -5823 5618 -5811
rect 5542 -5875 5554 -5823
rect 5606 -5875 5618 -5823
rect 8954 -5850 8966 -5798
rect 9018 -5850 9030 -5798
rect 8954 -5862 9030 -5850
rect 5542 -5887 5618 -5875
rect 7825 -6076 7921 -6059
rect 7825 -6149 7842 -6076
rect 7905 -6149 7921 -6076
rect 7825 -6166 7921 -6149
rect 7821 -6448 7917 -6431
rect 7821 -6521 7838 -6448
rect 7901 -6521 7917 -6448
rect 7821 -6538 7917 -6521
rect 7825 -6833 7921 -6816
rect 7825 -6906 7842 -6833
rect 7905 -6906 7921 -6833
rect 7825 -6923 7921 -6906
rect -3330 -6987 -3244 -6974
rect -3330 -7047 -3319 -6987
rect -3257 -7047 -3244 -6987
rect -3330 -7055 -3244 -7047
rect -3003 -7014 -2927 -7002
rect -3003 -7066 -2991 -7014
rect -2939 -7066 -2927 -7014
rect 7354 -7028 7430 -7016
rect -3003 -7078 -2927 -7066
rect 238 -7084 440 -7064
rect 238 -7149 256 -7084
rect 320 -7086 440 -7084
rect 7354 -7080 7366 -7028
rect 7418 -7080 7430 -7028
rect 320 -7149 378 -7086
rect 238 -7151 378 -7149
rect 7354 -7092 7430 -7080
rect 238 -7168 440 -7151
rect -4113 -7253 9020 -7216
rect 9180 -7253 9643 -29
rect -4391 -7616 9643 -7253
<< via1 >>
rect 29 7608 96 7680
rect 170 7610 237 7682
rect 32 7469 99 7541
rect 165 7473 232 7545
rect 8934 7141 8986 7193
rect 1230 6907 1292 6976
rect 3009 6960 3071 7029
rect 4824 6949 4886 7018
rect 6640 7024 6702 7093
rect 6641 6902 6703 6971
rect 3009 6751 3071 6820
rect 4825 6761 4887 6830
rect 6641 6780 6703 6849
rect 1233 6533 1295 6602
rect 3013 6519 3075 6588
rect 4824 6580 4886 6649
rect 1233 6200 1295 6269
rect 1898 5910 1950 5962
rect 3710 5910 3762 5962
rect 5522 5910 5574 5962
rect 7334 5911 7386 5963
rect 7646 4353 7709 4426
rect 8288 4357 8351 4430
rect 7647 4106 7710 4179
rect 8288 4097 8351 4170
rect -4589 3930 -4519 3998
rect -4465 3930 -4395 3998
rect -4341 3930 -4271 3998
rect -4217 3930 -4147 3998
rect -4589 3806 -4519 3874
rect -4465 3806 -4395 3874
rect -4341 3806 -4271 3874
rect -4217 3806 -4147 3874
rect 1393 3834 1445 3886
rect 2223 3834 2275 3886
rect 4035 3834 4087 3886
rect 5847 3834 5899 3886
rect 1206 3462 1258 3514
rect 2410 3462 2462 3514
rect 4190 3462 4242 3514
rect 6034 3462 6086 3514
rect 7361 3462 7413 3514
rect -2749 2839 -2697 2891
rect -2185 2839 -2133 2891
rect -1682 2839 -1630 2891
rect -47 2581 5 2633
rect -169 2398 -117 2450
rect -291 1570 -239 1622
rect 1686 1607 1738 1659
rect -47 1478 5 1530
rect 86 1478 138 1530
rect 3530 1478 3582 1530
rect 7154 1478 7206 1530
rect 8966 1478 9018 1530
rect -2748 1129 -2696 1181
rect -2184 1129 -2132 1181
rect -1681 1129 -1629 1181
rect 7841 1176 7904 1249
rect 7837 777 7900 850
rect -413 688 -361 740
rect 7841 404 7904 477
rect 5310 247 5362 299
rect 566 -202 618 -150
rect 3050 -202 3102 -150
rect 4830 -202 4882 -150
rect 6674 -202 6726 -150
rect 7361 -202 7413 -150
rect 7839 -402 7902 -329
rect -2748 -581 -2696 -529
rect -2184 -581 -2132 -529
rect -1681 -581 -1629 -529
rect 7843 -780 7906 -707
rect -535 -1022 -483 -970
rect 7841 -1167 7904 -1094
rect -4610 -1502 -4540 -1434
rect -3953 -1436 -3901 -1384
rect -3653 -1436 -3601 -1384
rect -3353 -1436 -3301 -1384
rect -3053 -1436 -3001 -1384
rect -2753 -1436 -2701 -1384
rect 86 -1418 138 -1366
rect 3530 -1418 3582 -1366
rect 7154 -1418 7206 -1366
rect 8966 -1418 9018 -1366
rect -4610 -1626 -4540 -1558
rect -4486 -1626 -4416 -1558
rect -4362 -1626 -4292 -1558
rect -4610 -1750 -4540 -1682
rect -4486 -1750 -4416 -1682
rect -4362 -1750 -4292 -1682
rect 1930 -3417 1982 -3365
rect 5554 -3417 5606 -3365
rect -3953 -3634 -3901 -3582
rect -3653 -3634 -3601 -3582
rect -3353 -3634 -3301 -3582
rect -3053 -3634 -3001 -3582
rect -2753 -3634 -2701 -3582
rect -2449 -3836 -2385 -3773
rect -2323 -3837 -2259 -3774
rect -1473 -3905 -1411 -3841
rect -1147 -3866 -1095 -3814
rect 4025 -3866 4077 -3814
rect 5047 -3812 5116 -3749
rect -4111 -5850 -4059 -5798
rect -667 -5850 -615 -5798
rect -291 -5850 -239 -5798
rect 86 -5850 138 -5798
rect 1686 -5875 1738 -5823
rect 1930 -5875 1982 -5823
rect 3530 -5850 3582 -5798
rect 5310 -5875 5362 -5823
rect 5554 -5875 5606 -5823
rect 7154 -5850 7206 -5798
rect 8966 -5850 9018 -5798
rect 7842 -6149 7905 -6076
rect 7838 -6521 7901 -6448
rect 7842 -6906 7905 -6833
rect -3319 -7047 -3257 -6987
rect -2991 -7066 -2939 -7014
rect 256 -7149 320 -7084
rect 7366 -7080 7418 -7028
rect 378 -7151 442 -7086
<< metal2 >>
rect 10 7682 260 7706
rect 10 7680 170 7682
rect 10 7608 29 7680
rect 96 7610 170 7680
rect 237 7610 260 7682
rect 96 7608 260 7610
rect 10 7545 260 7608
rect 10 7541 165 7545
rect 10 7469 32 7541
rect 99 7473 165 7541
rect 232 7473 260 7545
rect 99 7469 260 7473
rect 10 7448 260 7469
rect 550 7195 633 7208
rect 550 7139 564 7195
rect 620 7139 633 7195
rect 550 5832 633 7139
rect 8922 7195 8998 7205
rect 8922 7139 8932 7195
rect 8988 7139 8998 7195
rect 8922 7129 8998 7139
rect 6619 7103 6728 7120
rect 2988 7029 3098 7102
rect 1208 6976 1318 7022
rect 1208 6907 1230 6976
rect 1292 6907 1318 6976
rect 1208 6602 1318 6907
rect 1208 6533 1233 6602
rect 1295 6533 1318 6602
rect 1208 6269 1318 6533
rect 2988 6960 3009 7029
rect 3071 6960 3098 7029
rect 2988 6820 3098 6960
rect 2988 6751 3009 6820
rect 3071 6751 3098 6820
rect 2988 6588 3098 6751
rect 2988 6519 3013 6588
rect 3075 6519 3098 6588
rect 4803 7018 4913 7099
rect 4803 6949 4824 7018
rect 4886 6949 4913 7018
rect 4803 6830 4913 6949
rect 4803 6761 4825 6830
rect 4887 6761 4913 6830
rect 4803 6662 4913 6761
rect 6616 7093 6728 7103
rect 6616 7024 6640 7093
rect 6702 7024 6728 7093
rect 6616 6971 6728 7024
rect 6616 6902 6641 6971
rect 6703 6902 6728 6971
rect 6616 6862 6728 6902
rect 6616 6849 10244 6862
rect 6616 6780 6641 6849
rect 6703 6780 10244 6849
rect 6616 6752 10244 6780
rect 4803 6649 10233 6662
rect 4803 6580 4824 6649
rect 4886 6580 10233 6649
rect 4803 6552 10233 6580
rect 2988 6462 3098 6519
rect 2988 6352 10209 6462
rect 1208 6200 1233 6269
rect 1295 6262 1318 6269
rect 1295 6200 10198 6262
rect 1208 6152 10198 6200
rect 1886 5964 1962 5974
rect 1886 5908 1896 5964
rect 1952 5908 1962 5964
rect 1886 5898 1962 5908
rect 3698 5964 3774 5974
rect 3698 5908 3708 5964
rect 3764 5908 3774 5964
rect 3698 5898 3774 5908
rect 5510 5964 5586 5974
rect 5510 5908 5520 5964
rect 5576 5908 5586 5964
rect 5510 5898 5586 5908
rect 7322 5965 7398 5975
rect 7322 5909 7332 5965
rect 7388 5909 7398 5965
rect 7322 5899 7398 5909
rect 8939 5965 10207 5987
rect 8939 5909 8964 5965
rect 9020 5964 10207 5965
rect 9020 5909 9080 5964
rect 8939 5908 9080 5909
rect 9136 5908 10207 5964
rect 8939 5889 10207 5908
rect 437 5749 633 5832
rect 437 5216 520 5749
rect 437 5133 667 5216
rect 8947 5184 9035 5889
rect -4651 3998 -4048 4035
rect -4651 3930 -4589 3998
rect -4519 3930 -4465 3998
rect -4395 3930 -4341 3998
rect -4271 3930 -4217 3998
rect -4147 3930 -4048 3998
rect -4651 3874 -4048 3930
rect -4651 3806 -4589 3874
rect -4519 3806 -4465 3874
rect -4395 3806 -4341 3874
rect -4271 3806 -4217 3874
rect -4147 3806 -4048 3874
rect -4651 3701 -4048 3806
rect -4651 -1357 -4360 3701
rect 584 3109 667 5133
rect 8754 5096 9035 5184
rect 7629 4426 7725 4443
rect 7629 4353 7646 4426
rect 7709 4353 7725 4426
rect 7629 4336 7725 4353
rect 8271 4430 8367 4447
rect 8271 4357 8288 4430
rect 8351 4357 8367 4430
rect 8271 4340 8367 4357
rect 7630 4179 7726 4196
rect 7630 4106 7647 4179
rect 7710 4106 7726 4179
rect 7630 4089 7726 4106
rect 8271 4170 8367 4187
rect 8271 4097 8288 4170
rect 8351 4097 8367 4170
rect 8271 4080 8367 4097
rect 1381 3888 1457 3898
rect 1204 3886 1457 3888
rect 1204 3834 1393 3886
rect 1445 3834 1457 3886
rect 1204 3832 1457 3834
rect 1204 3526 1260 3832
rect 1381 3822 1457 3832
rect 2211 3888 2287 3898
rect 4023 3888 4099 3898
rect 4809 3888 5231 3898
rect 2211 3886 2464 3888
rect 2211 3834 2223 3886
rect 2275 3834 2464 3886
rect 2211 3832 2464 3834
rect 2211 3822 2287 3832
rect 2408 3526 2464 3832
rect 4023 3886 4244 3888
rect 4023 3834 4035 3886
rect 4087 3834 4244 3886
rect 4023 3832 4244 3834
rect 4023 3822 4099 3832
rect 4188 3526 4244 3832
rect 4809 3832 4828 3888
rect 4884 3832 5231 3888
rect 4809 3798 5231 3832
rect 5835 3888 5911 3898
rect 5835 3832 5845 3888
rect 5901 3832 5911 3888
rect 5835 3822 5911 3832
rect 1194 3514 1270 3526
rect 1194 3462 1206 3514
rect 1258 3462 1270 3514
rect 1194 3450 1270 3462
rect 2398 3514 2474 3526
rect 2398 3462 2410 3514
rect 2462 3462 2474 3514
rect 2398 3450 2474 3462
rect 4178 3514 4254 3526
rect 4178 3462 4190 3514
rect 4242 3462 4254 3514
rect 4178 3450 4254 3462
rect 544 2980 667 3109
rect -2761 2893 -2685 2903
rect -2761 2837 -2751 2893
rect -2695 2837 -2685 2893
rect -2761 2827 -2685 2837
rect -2197 2893 -2121 2903
rect -2197 2837 -2187 2893
rect -2131 2837 -2121 2893
rect -2197 2827 -2121 2837
rect -1694 2893 -1618 2903
rect -1694 2837 -1684 2893
rect -1628 2837 -1618 2893
rect -1694 2827 -1618 2837
rect -59 2633 17 2645
rect -59 2581 -47 2633
rect 5 2581 17 2633
rect -59 2569 17 2581
rect -181 2450 -105 2462
rect -181 2398 -169 2450
rect -117 2398 -105 2450
rect -181 2386 -105 2398
rect -303 1622 -227 1634
rect -303 1570 -291 1622
rect -239 1570 -227 1622
rect -303 1558 -227 1570
rect -2760 1183 -2684 1193
rect -2760 1127 -2750 1183
rect -2694 1127 -2684 1183
rect -2760 1117 -2684 1127
rect -2196 1183 -2120 1193
rect -2196 1127 -2186 1183
rect -2130 1127 -2120 1183
rect -2196 1117 -2120 1127
rect -1693 1183 -1617 1193
rect -1693 1127 -1683 1183
rect -1627 1127 -1617 1183
rect -1693 1117 -1617 1127
rect -425 740 -349 752
rect -425 688 -413 740
rect -361 688 -349 740
rect -425 676 -349 688
rect -2760 -527 -2684 -517
rect -2760 -583 -2750 -527
rect -2694 -583 -2684 -527
rect -2760 -593 -2684 -583
rect -2196 -527 -2120 -517
rect -2196 -583 -2186 -527
rect -2130 -583 -2120 -527
rect -2196 -593 -2120 -583
rect -1693 -527 -1617 -517
rect -1693 -583 -1683 -527
rect -1627 -583 -1617 -527
rect -1693 -593 -1617 -583
rect -4683 -1434 -4175 -1357
rect -4683 -1502 -4610 -1434
rect -4540 -1502 -4175 -1434
rect -4683 -1558 -4175 -1502
rect -4683 -1620 -4610 -1558
rect -4651 -1626 -4610 -1620
rect -4540 -1626 -4486 -1558
rect -4416 -1626 -4362 -1558
rect -4292 -1626 -4175 -1558
rect -4651 -1682 -4175 -1626
rect -4651 -1750 -4610 -1682
rect -4540 -1750 -4486 -1682
rect -4416 -1750 -4362 -1682
rect -4292 -1750 -4175 -1682
rect -4651 -1817 -4175 -1750
rect -3983 -1384 -3871 -1374
rect -3983 -1436 -3953 -1384
rect -3901 -1436 -3871 -1384
rect -3983 -1809 -3871 -1436
rect -3683 -1384 -3571 -1374
rect -3683 -1436 -3653 -1384
rect -3601 -1436 -3571 -1384
rect -3683 -1809 -3571 -1436
rect -3383 -1384 -3271 -1374
rect -3383 -1436 -3353 -1384
rect -3301 -1436 -3271 -1384
rect -3383 -1809 -3271 -1436
rect -3083 -1384 -2971 -1374
rect -3083 -1436 -3053 -1384
rect -3001 -1436 -2971 -1384
rect -3083 -1809 -2971 -1436
rect -2783 -1384 -2671 -1374
rect -2783 -1436 -2753 -1384
rect -2701 -1436 -2671 -1384
rect -2783 -1809 -2671 -1436
rect -4651 -2295 -4360 -1817
rect -3983 -1921 -2671 -1809
rect -3983 -2295 -3871 -1921
rect -3683 -2295 -3571 -1921
rect -3383 -2295 -3271 -1921
rect -3083 -2295 -2971 -1921
rect -2783 -2295 -2671 -1921
rect -4651 -2586 -2671 -2295
rect -3983 -3048 -3871 -2586
rect -3683 -3048 -3571 -2586
rect -3383 -3048 -3271 -2586
rect -3083 -3048 -2971 -2586
rect -2783 -3048 -2671 -2586
rect -3983 -3160 -2671 -3048
rect -3983 -3582 -3871 -3160
rect -3983 -3634 -3953 -3582
rect -3901 -3634 -3871 -3582
rect -3983 -3646 -3871 -3634
rect -3683 -3582 -3571 -3160
rect -3683 -3634 -3653 -3582
rect -3601 -3634 -3571 -3582
rect -3683 -3646 -3571 -3634
rect -3383 -3582 -3271 -3160
rect -3383 -3634 -3353 -3582
rect -3301 -3634 -3271 -3582
rect -3383 -3646 -3271 -3634
rect -3083 -3582 -2971 -3160
rect -3083 -3634 -3053 -3582
rect -3001 -3634 -2971 -3582
rect -3083 -3646 -2971 -3634
rect -2783 -3582 -2671 -3160
rect -2783 -3634 -2753 -3582
rect -2701 -3634 -2671 -3582
rect -2783 -3646 -2671 -3634
rect -2495 -3773 -2228 -3745
rect -2495 -3836 -2449 -3773
rect -2385 -3774 -2228 -3773
rect -2385 -3836 -2323 -3774
rect -2495 -3837 -2323 -3836
rect -2259 -3837 -2228 -3774
rect -1159 -3812 -1083 -3802
rect -2495 -3852 -2228 -3837
rect -1489 -3841 -1397 -3827
rect -1489 -3905 -1473 -3841
rect -1411 -3905 -1397 -3841
rect -1159 -3868 -1149 -3812
rect -1093 -3868 -1083 -3812
rect -1159 -3878 -1083 -3868
rect -1489 -3917 -1397 -3905
rect -669 -5786 -613 -776
rect -547 -970 -471 -958
rect -547 -1022 -535 -970
rect -483 -1022 -471 -970
rect -547 -1034 -471 -1022
rect -537 -5786 -481 -1034
rect -415 -3245 -359 676
rect -425 -3255 -349 -3245
rect -425 -3311 -415 -3255
rect -359 -3311 -349 -3255
rect -425 -3321 -349 -3311
rect -293 -5786 -237 1558
rect -171 -1354 -115 2386
rect -49 1542 7 2569
rect 544 2330 627 2980
rect 544 2247 792 2330
rect 5131 2319 5231 3798
rect 6022 3516 6098 3526
rect 6022 3460 6032 3516
rect 6088 3460 6098 3516
rect 6022 3450 6098 3460
rect 7349 3516 7425 3526
rect 7349 3460 7359 3516
rect 7415 3460 7425 3516
rect 7349 3450 7425 3460
rect 8754 2944 8842 5096
rect 8754 2856 8999 2944
rect -59 1530 17 1542
rect -59 1478 -47 1530
rect 5 1478 17 1530
rect -59 1466 17 1478
rect 74 1532 150 1542
rect 74 1476 84 1532
rect 140 1476 150 1532
rect 74 1466 150 1476
rect 84 -1354 140 1466
rect 709 -132 792 2247
rect 4969 2219 5231 2319
rect 1642 1673 1759 1687
rect 4969 1676 5069 2219
rect 1642 1659 1766 1673
rect 1642 1607 1686 1659
rect 1738 1607 1766 1659
rect 1642 1588 1766 1607
rect 1653 1574 1766 1588
rect 545 -150 792 -132
rect 545 -202 566 -150
rect 618 -202 792 -150
rect 545 -215 792 -202
rect -181 -1364 -105 -1354
rect -181 -1420 -171 -1364
rect -115 -1420 -105 -1364
rect -181 -1430 -105 -1420
rect 74 -1366 150 -1354
rect 74 -1418 86 -1366
rect 138 -1418 150 -1366
rect 74 -1430 150 -1418
rect 1671 -2059 1766 1574
rect 4804 1576 5069 1676
rect 3518 1530 3594 1542
rect 3518 1478 3530 1530
rect 3582 1478 3594 1530
rect 3518 1466 3594 1478
rect 3030 -150 3124 -127
rect 3030 -202 3050 -150
rect 3102 -202 3124 -150
rect 3030 -1508 3124 -202
rect 3528 -1354 3584 1466
rect 4804 -150 4904 1576
rect 8911 1551 8999 2856
rect 7142 1532 7218 1542
rect 7142 1476 7152 1532
rect 7208 1476 7218 1532
rect 7142 1466 7218 1476
rect 8911 1530 9046 1551
rect 8911 1478 8966 1530
rect 9018 1478 9046 1530
rect 4804 -202 4830 -150
rect 4882 -202 4904 -150
rect 4804 -222 4904 -202
rect 5286 299 5388 334
rect 5286 247 5310 299
rect 5362 247 5388 299
rect 3518 -1364 3594 -1354
rect 3518 -1420 3528 -1364
rect 3584 -1420 3594 -1364
rect 3518 -1430 3594 -1420
rect 3030 -1602 3435 -1508
rect 1502 -2154 1766 -2059
rect 1502 -5069 1597 -2154
rect 1910 -3365 2487 -3349
rect 1910 -3417 1930 -3365
rect 1982 -3417 2487 -3365
rect 1910 -3455 2487 -3417
rect 2381 -5034 2487 -3455
rect 1502 -5164 1759 -5069
rect -4123 -5796 -4047 -5786
rect -4123 -5852 -4113 -5796
rect -4057 -5852 -4047 -5796
rect -4123 -5862 -4047 -5852
rect -679 -5798 -603 -5786
rect -679 -5850 -667 -5798
rect -615 -5850 -603 -5798
rect -679 -5862 -603 -5850
rect -547 -5796 -471 -5786
rect -547 -5852 -537 -5796
rect -481 -5852 -471 -5796
rect -547 -5862 -471 -5852
rect -303 -5798 -227 -5786
rect -303 -5850 -291 -5798
rect -239 -5850 -227 -5798
rect -303 -5862 -227 -5850
rect 74 -5796 150 -5786
rect 74 -5852 84 -5796
rect 140 -5852 150 -5796
rect 74 -5862 150 -5852
rect 1664 -5823 1759 -5164
rect 2230 -5140 2487 -5034
rect 2230 -5795 2336 -5140
rect 3341 -5598 3435 -1602
rect 5286 -2053 5388 247
rect 6662 -148 6738 -138
rect 6662 -204 6672 -148
rect 6728 -204 6738 -148
rect 6662 -214 6738 -204
rect 7152 -1354 7208 1466
rect 8911 1463 9046 1478
rect 7824 1249 7920 1266
rect 7824 1176 7841 1249
rect 7904 1176 7920 1249
rect 7824 1159 7920 1176
rect 7820 850 7916 867
rect 7820 777 7837 850
rect 7900 777 7916 850
rect 7820 760 7916 777
rect 7824 477 7920 494
rect 7824 404 7841 477
rect 7904 404 7920 477
rect 7824 387 7920 404
rect 7349 -148 7425 -138
rect 7349 -204 7359 -148
rect 7415 -204 7425 -148
rect 7349 -214 7425 -204
rect 7822 -329 7918 -312
rect 7822 -402 7839 -329
rect 7902 -402 7918 -329
rect 7822 -419 7918 -402
rect 7826 -707 7922 -690
rect 7826 -780 7843 -707
rect 7906 -780 7922 -707
rect 7826 -797 7922 -780
rect 7824 -1094 7920 -1077
rect 7824 -1167 7841 -1094
rect 7904 -1167 7920 -1094
rect 7824 -1184 7920 -1167
rect 8911 -1352 8999 1463
rect 7142 -1366 7218 -1354
rect 7142 -1418 7154 -1366
rect 7206 -1418 7218 -1366
rect 7142 -1430 7218 -1418
rect 8911 -1366 9046 -1352
rect 8911 -1418 8966 -1366
rect 9018 -1418 9046 -1366
rect 5120 -2155 5388 -2053
rect 8911 -1440 9046 -1418
rect 5120 -2720 5222 -2155
rect 5120 -2822 5375 -2720
rect 3518 -3255 3594 -3245
rect 3518 -3311 3528 -3255
rect 3584 -3311 3594 -3255
rect 3518 -3321 3594 -3311
rect 1664 -5875 1686 -5823
rect 1738 -5875 1759 -5823
rect 1664 -5899 1759 -5875
rect 1906 -5823 2336 -5795
rect 1906 -5875 1930 -5823
rect 1982 -5875 2336 -5823
rect 1906 -5901 2336 -5875
rect 3028 -5692 3435 -5598
rect -3330 -6987 -3244 -6974
rect -3330 -7047 -3319 -6987
rect -3257 -7047 -3244 -6987
rect -3330 -7055 -3244 -7047
rect -3003 -7012 -2927 -7002
rect -3003 -7068 -2993 -7012
rect -2937 -7068 -2927 -7012
rect -3003 -7078 -2927 -7068
rect 3028 -7026 3122 -5692
rect 3528 -5786 3584 -3321
rect 5033 -3749 5131 -3733
rect 4013 -3812 4089 -3802
rect 4013 -3868 4023 -3812
rect 4079 -3868 4089 -3812
rect 5033 -3812 5047 -3749
rect 5116 -3812 5131 -3749
rect 5033 -3825 5131 -3812
rect 4013 -3878 4089 -3868
rect 5273 -4022 5375 -2822
rect 5537 -3365 5793 -3351
rect 5537 -3417 5554 -3365
rect 5606 -3417 5793 -3365
rect 5537 -3453 5793 -3417
rect 5130 -4124 5375 -4022
rect 5130 -5026 5232 -4124
rect 5691 -5011 5793 -3453
rect 4968 -5128 5232 -5026
rect 5530 -5113 5793 -5011
rect 4968 -5618 5070 -5128
rect 4968 -5720 5387 -5618
rect 3518 -5798 3594 -5786
rect 3518 -5850 3530 -5798
rect 3582 -5850 3594 -5798
rect 3518 -5862 3594 -5850
rect 5285 -5823 5387 -5720
rect 5285 -5875 5310 -5823
rect 5362 -5875 5387 -5823
rect 5285 -5906 5387 -5875
rect 5530 -5823 5632 -5113
rect 8911 -5781 8999 -1440
rect 5530 -5875 5554 -5823
rect 5606 -5875 5632 -5823
rect 7142 -5796 7218 -5786
rect 7142 -5852 7152 -5796
rect 7208 -5852 7218 -5796
rect 7142 -5862 7218 -5852
rect 8911 -5798 9049 -5781
rect 8911 -5850 8966 -5798
rect 9018 -5850 9049 -5798
rect 8911 -5869 9049 -5850
rect 5530 -5902 5632 -5875
rect 7825 -6076 7921 -6059
rect 7825 -6149 7842 -6076
rect 7905 -6149 7921 -6076
rect 7825 -6166 7921 -6149
rect 7821 -6448 7917 -6431
rect 7821 -6521 7838 -6448
rect 7901 -6521 7917 -6448
rect 7821 -6538 7917 -6521
rect 7825 -6833 7921 -6816
rect 7825 -6906 7842 -6833
rect 7905 -6906 7921 -6833
rect 7825 -6923 7921 -6906
rect 238 -7084 456 -7069
rect 238 -7149 256 -7084
rect 320 -7086 456 -7084
rect 320 -7149 378 -7086
rect 238 -7151 378 -7149
rect 442 -7151 456 -7086
rect 3028 -7082 3048 -7026
rect 3104 -7082 3122 -7026
rect 3028 -7099 3122 -7082
rect 7354 -7026 7430 -7016
rect 7354 -7082 7364 -7026
rect 7420 -7082 7430 -7026
rect 7354 -7092 7430 -7082
rect 238 -7167 456 -7151
<< via2 >>
rect 29 7608 96 7680
rect 170 7610 237 7682
rect 32 7469 99 7541
rect 165 7473 232 7545
rect 564 7139 620 7195
rect 8932 7193 8988 7195
rect 8932 7141 8934 7193
rect 8934 7141 8986 7193
rect 8986 7141 8988 7193
rect 8932 7139 8988 7141
rect 1896 5962 1952 5964
rect 1896 5910 1898 5962
rect 1898 5910 1950 5962
rect 1950 5910 1952 5962
rect 1896 5908 1952 5910
rect 3708 5962 3764 5964
rect 3708 5910 3710 5962
rect 3710 5910 3762 5962
rect 3762 5910 3764 5962
rect 3708 5908 3764 5910
rect 5520 5962 5576 5964
rect 5520 5910 5522 5962
rect 5522 5910 5574 5962
rect 5574 5910 5576 5962
rect 5520 5908 5576 5910
rect 7332 5963 7388 5965
rect 7332 5911 7334 5963
rect 7334 5911 7386 5963
rect 7386 5911 7388 5963
rect 7332 5909 7388 5911
rect 8964 5909 9020 5965
rect 9080 5908 9136 5964
rect 7646 4353 7709 4426
rect 8288 4357 8351 4430
rect 7647 4106 7710 4179
rect 8288 4097 8351 4170
rect 4828 3832 4884 3888
rect 5845 3886 5901 3888
rect 5845 3834 5847 3886
rect 5847 3834 5899 3886
rect 5899 3834 5901 3886
rect 5845 3832 5901 3834
rect -2751 2891 -2695 2893
rect -2751 2839 -2749 2891
rect -2749 2839 -2697 2891
rect -2697 2839 -2695 2891
rect -2751 2837 -2695 2839
rect -2187 2891 -2131 2893
rect -2187 2839 -2185 2891
rect -2185 2839 -2133 2891
rect -2133 2839 -2131 2891
rect -2187 2837 -2131 2839
rect -1684 2891 -1628 2893
rect -1684 2839 -1682 2891
rect -1682 2839 -1630 2891
rect -1630 2839 -1628 2891
rect -1684 2837 -1628 2839
rect -2750 1181 -2694 1183
rect -2750 1129 -2748 1181
rect -2748 1129 -2696 1181
rect -2696 1129 -2694 1181
rect -2750 1127 -2694 1129
rect -2186 1181 -2130 1183
rect -2186 1129 -2184 1181
rect -2184 1129 -2132 1181
rect -2132 1129 -2130 1181
rect -2186 1127 -2130 1129
rect -1683 1181 -1627 1183
rect -1683 1129 -1681 1181
rect -1681 1129 -1629 1181
rect -1629 1129 -1627 1181
rect -1683 1127 -1627 1129
rect -2750 -529 -2694 -527
rect -2750 -581 -2748 -529
rect -2748 -581 -2696 -529
rect -2696 -581 -2694 -529
rect -2750 -583 -2694 -581
rect -2186 -529 -2130 -527
rect -2186 -581 -2184 -529
rect -2184 -581 -2132 -529
rect -2132 -581 -2130 -529
rect -2186 -583 -2130 -581
rect -1683 -529 -1627 -527
rect -1683 -581 -1681 -529
rect -1681 -581 -1629 -529
rect -1629 -581 -1627 -529
rect -1683 -583 -1627 -581
rect -2449 -3836 -2385 -3773
rect -2323 -3837 -2259 -3774
rect -1473 -3905 -1411 -3841
rect -1149 -3814 -1093 -3812
rect -1149 -3866 -1147 -3814
rect -1147 -3866 -1095 -3814
rect -1095 -3866 -1093 -3814
rect -1149 -3868 -1093 -3866
rect -415 -3311 -359 -3255
rect 6032 3514 6088 3516
rect 6032 3462 6034 3514
rect 6034 3462 6086 3514
rect 6086 3462 6088 3514
rect 6032 3460 6088 3462
rect 7359 3514 7415 3516
rect 7359 3462 7361 3514
rect 7361 3462 7413 3514
rect 7413 3462 7415 3514
rect 7359 3460 7415 3462
rect 84 1530 140 1532
rect 84 1478 86 1530
rect 86 1478 138 1530
rect 138 1478 140 1530
rect 84 1476 140 1478
rect -171 -1420 -115 -1364
rect 7152 1530 7208 1532
rect 7152 1478 7154 1530
rect 7154 1478 7206 1530
rect 7206 1478 7208 1530
rect 7152 1476 7208 1478
rect 3528 -1366 3584 -1364
rect 3528 -1418 3530 -1366
rect 3530 -1418 3582 -1366
rect 3582 -1418 3584 -1366
rect 3528 -1420 3584 -1418
rect -4113 -5798 -4057 -5796
rect -4113 -5850 -4111 -5798
rect -4111 -5850 -4059 -5798
rect -4059 -5850 -4057 -5798
rect -4113 -5852 -4057 -5850
rect -537 -5852 -481 -5796
rect 84 -5798 140 -5796
rect 84 -5850 86 -5798
rect 86 -5850 138 -5798
rect 138 -5850 140 -5798
rect 84 -5852 140 -5850
rect 6672 -150 6728 -148
rect 6672 -202 6674 -150
rect 6674 -202 6726 -150
rect 6726 -202 6728 -150
rect 6672 -204 6728 -202
rect 7841 1176 7904 1249
rect 7837 777 7900 850
rect 7841 404 7904 477
rect 7359 -150 7415 -148
rect 7359 -202 7361 -150
rect 7361 -202 7413 -150
rect 7413 -202 7415 -150
rect 7359 -204 7415 -202
rect 7839 -402 7902 -329
rect 7843 -780 7906 -707
rect 7841 -1167 7904 -1094
rect 3528 -3311 3584 -3255
rect -3319 -7047 -3257 -6987
rect -2993 -7014 -2937 -7012
rect -2993 -7066 -2991 -7014
rect -2991 -7066 -2939 -7014
rect -2939 -7066 -2937 -7014
rect -2993 -7068 -2937 -7066
rect 4023 -3814 4079 -3812
rect 4023 -3866 4025 -3814
rect 4025 -3866 4077 -3814
rect 4077 -3866 4079 -3814
rect 4023 -3868 4079 -3866
rect 5047 -3812 5116 -3749
rect 7152 -5798 7208 -5796
rect 7152 -5850 7154 -5798
rect 7154 -5850 7206 -5798
rect 7206 -5850 7208 -5798
rect 7152 -5852 7208 -5850
rect 7842 -6149 7905 -6076
rect 7838 -6521 7901 -6448
rect 7842 -6906 7905 -6833
rect 256 -7149 320 -7084
rect 378 -7151 442 -7086
rect 3048 -7082 3104 -7026
rect 7364 -7028 7420 -7026
rect 7364 -7080 7366 -7028
rect 7366 -7080 7418 -7028
rect 7418 -7080 7420 -7028
rect 7364 -7082 7420 -7080
<< metal3 >>
rect -2215 7682 321 7757
rect -2215 7680 170 7682
rect -2215 7608 29 7680
rect 96 7610 170 7680
rect 237 7610 321 7682
rect 96 7608 321 7610
rect -2215 7545 321 7608
rect -2215 7541 165 7545
rect -2215 7469 32 7541
rect 99 7473 165 7541
rect 232 7473 321 7545
rect 99 7469 321 7473
rect -2215 7408 321 7469
rect -2215 6685 -2103 7408
rect -1712 6685 -1600 7408
rect 554 7195 630 7205
rect 8922 7195 8998 7205
rect 554 7139 564 7195
rect 620 7139 8932 7195
rect 8988 7139 8998 7195
rect 554 7129 630 7139
rect 8922 7129 8998 7139
rect -2215 6573 -1600 6685
rect -2215 5802 -2103 6573
rect -1712 5802 -1600 6573
rect 1886 5964 1962 5974
rect 3698 5964 3774 5974
rect 5510 5964 5586 5974
rect 7322 5965 7398 5975
rect 8939 5965 9171 5987
rect 7322 5964 7332 5965
rect 1886 5908 1896 5964
rect 1952 5908 3708 5964
rect 3764 5908 5520 5964
rect 5576 5909 7332 5964
rect 7388 5909 8964 5965
rect 9020 5964 9171 5965
rect 9020 5909 9080 5964
rect 5576 5908 7398 5909
rect 1886 5898 1962 5908
rect 3698 5898 3774 5908
rect 5510 5898 5586 5908
rect 7322 5899 7398 5908
rect 8939 5908 9080 5909
rect 9136 5908 9171 5964
rect 8939 5889 9171 5908
rect -2215 5690 -1600 5802
rect -2215 5175 -2103 5690
rect -1712 5175 -1600 5690
rect -2215 5063 -1600 5175
rect -2215 4581 -2103 5063
rect -1712 4581 -1600 5063
rect -2215 4469 -1600 4581
rect -2779 2893 -2667 2921
rect -2779 2837 -2751 2893
rect -2695 2837 -2667 2893
rect -2779 1183 -2667 2837
rect -2779 1127 -2750 1183
rect -2694 1127 -2667 1183
rect -2779 -527 -2667 1127
rect -2779 -583 -2750 -527
rect -2694 -583 -2667 -527
rect -2779 -611 -2667 -583
rect -2215 2893 -2103 4469
rect -2215 2837 -2187 2893
rect -2131 2837 -2103 2893
rect -2215 1183 -2103 2837
rect -2215 1127 -2186 1183
rect -2130 1127 -2103 1183
rect -2215 -527 -2103 1127
rect -2215 -583 -2186 -527
rect -2130 -583 -2103 -527
rect -2215 -1382 -2103 -583
rect -1712 2893 -1600 4469
rect 7628 4426 7737 4467
rect 7628 4353 7646 4426
rect 7709 4353 7737 4426
rect 7628 4311 7737 4353
rect 8257 4430 8378 4461
rect 8257 4357 8288 4430
rect 8351 4357 8378 4430
rect 8257 4311 8378 4357
rect 7628 4202 10259 4311
rect 7628 4179 7737 4202
rect 7628 4106 7647 4179
rect 7710 4106 7737 4179
rect 7628 4058 7737 4106
rect 8257 4170 8378 4202
rect 8257 4097 8288 4170
rect 8351 4097 8378 4170
rect 8257 4061 8378 4097
rect 4796 3888 5921 3910
rect 4796 3832 4828 3888
rect 4884 3832 5845 3888
rect 5901 3832 5921 3888
rect 4796 3812 5921 3832
rect 6022 3516 6098 3526
rect 7349 3516 7425 3526
rect 6022 3460 6032 3516
rect 6088 3460 7359 3516
rect 7415 3460 7425 3516
rect 6022 3450 6098 3460
rect 7349 3450 7425 3460
rect -1712 2837 -1684 2893
rect -1628 2837 -1600 2893
rect -1712 1183 -1600 2837
rect 74 1532 150 1542
rect 7142 1532 7218 1542
rect 74 1476 84 1532
rect 140 1476 7152 1532
rect 7208 1476 7218 1532
rect 74 1466 150 1476
rect 7142 1466 7218 1476
rect -1712 1127 -1683 1183
rect -1627 1127 -1600 1183
rect -1712 -527 -1600 1127
rect 7815 1249 7924 1395
rect 7815 1176 7841 1249
rect 7904 1176 7924 1249
rect 7815 984 7924 1176
rect 7815 875 10206 984
rect 7815 850 7924 875
rect 7815 777 7837 850
rect 7900 777 7924 850
rect 7815 477 7924 777
rect 7815 404 7841 477
rect 7904 404 7924 477
rect 7815 351 7924 404
rect 6662 -148 6738 -138
rect 7349 -148 7425 -138
rect 6662 -204 6672 -148
rect 6728 -204 7359 -148
rect 7415 -204 7425 -148
rect 6662 -214 6738 -204
rect 7349 -214 7425 -204
rect -1712 -583 -1683 -527
rect -1627 -583 -1600 -527
rect -1712 -1382 -1600 -583
rect 7822 -329 7931 -236
rect 7822 -402 7839 -329
rect 7902 -402 7931 -329
rect 7822 -684 7931 -402
rect 7822 -707 10163 -684
rect 7822 -780 7843 -707
rect 7906 -780 10163 -707
rect 7822 -793 10163 -780
rect 7822 -1094 7931 -793
rect 7822 -1167 7841 -1094
rect 7904 -1167 7931 -1094
rect 7822 -1227 7931 -1167
rect -181 -1364 -105 -1354
rect 3518 -1364 3594 -1354
rect -181 -1420 -171 -1364
rect -115 -1420 3528 -1364
rect 3584 -1420 3594 -1364
rect -181 -1430 -105 -1420
rect 3518 -1430 3594 -1420
rect -425 -3255 -349 -3245
rect 3518 -3255 3594 -3245
rect -425 -3311 -415 -3255
rect -359 -3311 3528 -3255
rect 3584 -3311 3594 -3255
rect -425 -3321 -349 -3311
rect 3518 -3321 3594 -3311
rect -4608 -3773 -2221 -3726
rect -4608 -3836 -2449 -3773
rect -2385 -3774 -2221 -3773
rect -2385 -3836 -2323 -3774
rect -4608 -3837 -2323 -3836
rect -2259 -3837 -2221 -3774
rect 5010 -3749 5142 -3725
rect 5010 -3783 5047 -3749
rect -4608 -3870 -2221 -3837
rect -1492 -3812 5047 -3783
rect 5116 -3812 5142 -3749
rect -1492 -3841 -1149 -3812
rect -1492 -3905 -1473 -3841
rect -1411 -3868 -1149 -3841
rect -1093 -3868 4023 -3812
rect 4079 -3868 5142 -3812
rect -1411 -3894 5142 -3868
rect -1411 -3905 -1373 -3894
rect -1492 -3928 -1373 -3905
rect -4123 -5796 -4047 -5786
rect -547 -5796 -471 -5786
rect -4123 -5852 -4113 -5796
rect -4057 -5852 -537 -5796
rect -481 -5852 -471 -5796
rect -4123 -5862 -4047 -5852
rect -547 -5862 -471 -5852
rect 74 -5796 150 -5786
rect 7142 -5796 7218 -5786
rect 74 -5852 84 -5796
rect 140 -5852 7152 -5796
rect 7208 -5852 7218 -5796
rect 74 -5862 150 -5852
rect 7142 -5862 7218 -5852
rect 7817 -6076 7926 -5967
rect 7817 -6149 7842 -6076
rect 7905 -6149 7926 -6076
rect 7817 -6424 7926 -6149
rect 7817 -6448 10022 -6424
rect 7817 -6521 7838 -6448
rect 7901 -6521 10022 -6448
rect 7817 -6533 10022 -6521
rect 7817 -6833 7926 -6533
rect 7817 -6906 7842 -6833
rect 7905 -6906 7926 -6833
rect 7817 -6959 7926 -6906
rect -3335 -6987 455 -6974
rect -3335 -7047 -3319 -6987
rect -3257 -7012 455 -6987
rect -3257 -7047 -2993 -7012
rect -3335 -7068 -2993 -7047
rect -2937 -7068 455 -7012
rect -3335 -7084 455 -7068
rect -3335 -7101 256 -7084
rect 227 -7149 256 -7101
rect 320 -7086 455 -7084
rect 320 -7149 378 -7086
rect 227 -7151 378 -7149
rect 442 -7151 455 -7086
rect 2995 -7026 7458 -6993
rect 2995 -7082 3048 -7026
rect 3104 -7082 7364 -7026
rect 7420 -7082 7458 -7026
rect 2995 -7115 7458 -7082
rect 227 -7169 455 -7151
use Non_Ovl_CLK_Gen_Layout  Non_Ovl_CLK_Gen_Layout_0 ~/GF180Projects/Tapeout/Magic/Non_Ovl_CLK_Gen
timestamp 1699883071
transform 1 0 -3619 0 1 -611
box -1478 -868 3162 980
use Non_Ovl_CLK_Gen_Layout  Non_Ovl_CLK_Gen_Layout_1
timestamp 1699883071
transform 1 0 -3619 0 1 2809
box -1478 -868 3162 980
use Non_Ovl_CLK_Gen_Layout  Non_Ovl_CLK_Gen_Layout_2
timestamp 1699883071
transform 1 0 -3619 0 -1 1211
box -1478 -868 3162 980
use Transmission_Gate_Layout_mux  Transmission_Gate_Layout_mux_0 ~/GF180Projects/Tapeout/Magic/Logic_Gates/Transmission_Gate2
timestamp 1699854221
transform -1 0 6920 0 1 -7056
box -350 -272 1471 3508
use Transmission_Gate_Layout_mux  Transmission_Gate_Layout_mux_1
timestamp 1699854221
transform 1 0 3996 0 1 -7056
box -350 -272 1471 3508
use Transmission_Gate_Layout_mux  Transmission_Gate_Layout_mux_2
timestamp 1699854221
transform -1 0 3296 0 1 -7056
box -350 -272 1471 3508
use Transmission_Gate_Layout_mux  Transmission_Gate_Layout_mux_3
timestamp 1699854221
transform 1 0 372 0 1 -7056
box -350 -272 1471 3508
use Transmission_Gate_Layout_mux  Transmission_Gate_Layout_mux_4
timestamp 1699854221
transform 1 0 3996 0 1 272
box -350 -272 1471 3508
use Transmission_Gate_Layout_mux  Transmission_Gate_Layout_mux_5
timestamp 1699854221
transform -1 0 6920 0 1 272
box -350 -272 1471 3508
use Transmission_Gate_Layout_mux  Transmission_Gate_Layout_mux_6
timestamp 1699854221
transform -1 0 3296 0 1 272
box -350 -272 1471 3508
use Transmission_Gate_Layout_mux  Transmission_Gate_Layout_mux_7
timestamp 1699854221
transform 1 0 372 0 1 272
box -350 -272 1471 3508
use Transmission_Gate_Layout_mux  Transmission_Gate_Layout_mux_8
timestamp 1699854221
transform -1 0 6920 0 -1 -160
box -350 -272 1471 3508
use Transmission_Gate_Layout_mux  Transmission_Gate_Layout_mux_9
timestamp 1699854221
transform 1 0 3996 0 -1 -160
box -350 -272 1471 3508
use Transmission_Gate_Layout_mux  Transmission_Gate_Layout_mux_10
timestamp 1699854221
transform -1 0 3296 0 -1 -160
box -350 -272 1471 3508
use Transmission_Gate_Layout_mux  Transmission_Gate_Layout_mux_11
timestamp 1699854221
transform 1 0 372 0 -1 -160
box -350 -272 1471 3508
use Transmission_Gate_Layout_mux  Transmission_Gate_Layout_mux_12
timestamp 1699854221
transform -1 0 -901 0 1 -7056
box -350 -272 1471 3508
use Transmission_Gate_Layout_mux  Transmission_Gate_Layout_mux_13
timestamp 1699854221
transform 1 0 -3825 0 1 -7056
box -350 -272 1471 3508
use Transmission_Gate_Layout_mux  Transmission_Gate_Layout_mux_14
timestamp 1699854221
transform -1 0 8732 0 1 -7056
box -350 -272 1471 3508
use Transmission_Gate_Layout_mux  Transmission_Gate_Layout_mux_15
timestamp 1699854221
transform 1 0 5808 0 -1 7168
box -350 -272 1471 3508
use Transmission_Gate_Layout_mux  Transmission_Gate_Layout_mux_16
timestamp 1699854221
transform 1 0 2184 0 -1 7168
box -350 -272 1471 3508
use Transmission_Gate_Layout_mux  Transmission_Gate_Layout_mux_17
timestamp 1699854221
transform 1 0 3996 0 -1 7168
box -350 -272 1471 3508
use Transmission_Gate_Layout_mux  Transmission_Gate_Layout_mux_18
timestamp 1699854221
transform -1 0 1484 0 -1 7168
box -350 -272 1471 3508
use Transmission_Gate_Layout_mux  Transmission_Gate_Layout_mux_19
timestamp 1699854221
transform 1 0 7620 0 -1 7168
box -350 -272 1471 3508
use Transmission_Gate_Layout_mux  Transmission_Gate_Layout_mux_20
timestamp 1699854221
transform -1 0 8732 0 1 272
box -350 -272 1471 3508
use Transmission_Gate_Layout_mux  Transmission_Gate_Layout_mux_21
timestamp 1699854221
transform -1 0 8732 0 -1 -160
box -350 -272 1471 3508
<< labels >>
flabel metal1 -5082 3176 -5082 3176 0 FreeSans 320 0 0 0 A1
port 15 nsew
flabel metal1 -5088 841 -5088 841 0 FreeSans 320 0 0 0 B1
port 16 nsew
flabel metal1 -5079 -243 -5079 -243 0 FreeSans 320 0 0 0 C1
port 18 nsew
flabel metal1 3634 7382 3634 7382 0 FreeSans 320 0 0 0 VSS
port 19 nsew
flabel metal1 1831 -3615 1831 -3615 0 FreeSans 320 0 0 0 VDD
port 20 nsew
flabel metal3 -4518 -3800 -4518 -3800 0 FreeSans 1600 0 0 0 OUT
port 38 nsew
flabel metal3 10198 4256 10198 4256 0 FreeSans 1600 0 0 0 IN4
port 39 nsew
flabel metal3 10152 924 10152 924 0 FreeSans 1600 0 0 0 IN8
port 40 nsew
flabel metal3 10109 -750 10109 -750 0 FreeSans 1600 0 0 0 IN6
port 41 nsew
flabel metal3 9968 -6479 9968 -6479 0 FreeSans 1600 0 0 0 IN3
port 42 nsew
flabel metal2 10186 6816 10186 6816 0 FreeSans 1600 0 0 0 IN5
port 43 nsew
flabel metal2 10157 6584 10157 6584 0 FreeSans 1600 0 0 0 IN7
port 44 nsew
flabel metal2 10131 6368 10131 6368 0 FreeSans 1600 0 0 0 IN1
port 45 nsew
flabel metal2 10085 6165 10085 6165 0 FreeSans 1600 0 0 0 IN2
port 46 nsew
flabel metal2 10166 5897 10166 5897 0 FreeSans 1600 0 0 0 EN
port 47 nsew
<< end >>
