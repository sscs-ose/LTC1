magic
tech gf180mcuC
magscale 1 10
timestamp 1694669706
<< nwell >>
rect 1154 -30 2214 91
rect 1486 -410 2205 -254
rect 1154 -580 2214 -410
rect 1486 -960 2205 -580
rect 1154 -1243 2214 -960
rect 1486 -1549 2205 -1243
<< pwell >>
rect 494 170 507 177
<< ndiff >>
rect 494 170 507 177
<< psubdiff >>
rect 355 -1492 533 -1453
rect 355 -1538 418 -1492
rect 464 -1538 533 -1492
rect 355 -1575 533 -1538
<< psubdiffcont >>
rect 418 -1538 464 -1492
<< polysilicon >>
rect 1736 615 1836 617
rect 1304 590 2083 615
rect 1304 544 1328 590
rect 1374 589 2083 590
rect 1374 544 1989 589
rect 1304 543 1989 544
rect 2035 543 2083 589
rect 1304 515 2083 543
rect 187 410 729 413
rect 158 394 729 410
rect 158 393 320 394
rect 158 347 174 393
rect 220 348 320 393
rect 366 348 729 394
rect 1532 370 1632 515
rect 220 347 729 348
rect 158 331 729 347
rect 1736 336 1836 515
rect 187 313 729 331
rect 313 256 416 313
rect 316 206 416 256
rect 520 212 620 313
rect 1328 76 1428 196
rect 1940 76 2040 198
rect 112 -29 212 54
rect 724 -29 824 56
rect 1301 49 2082 76
rect 1301 3 1332 49
rect 1378 48 2082 49
rect 1378 3 2003 48
rect 1301 2 2003 3
rect 2049 2 2082 48
rect 1301 -24 2082 2
rect 112 -42 824 -29
rect 112 -57 825 -42
rect 112 -103 130 -57
rect 176 -59 825 -57
rect 176 -103 764 -59
rect 112 -105 764 -103
rect 810 -105 825 -59
rect 112 -121 825 -105
rect 112 -129 824 -121
rect 316 -198 416 -129
rect 520 -200 620 -129
rect 1532 -142 1632 -24
rect 1736 -144 1836 -24
rect 112 -480 212 -384
rect 724 -480 824 -382
rect 1328 -445 1428 -294
rect 1940 -445 2040 -311
rect 1307 -471 2100 -445
rect 1307 -472 2037 -471
rect 112 -504 826 -480
rect 112 -550 132 -504
rect 178 -510 826 -504
rect 178 -550 762 -510
rect 112 -556 762 -550
rect 808 -556 826 -510
rect 1307 -518 1327 -472
rect 1373 -517 2037 -472
rect 2083 -517 2100 -471
rect 1373 -518 2100 -517
rect 1307 -545 2100 -518
rect 112 -580 826 -556
rect 112 -669 212 -580
rect 724 -663 824 -580
rect 1328 -680 1428 -545
rect 1940 -680 2040 -545
rect 316 -951 416 -860
rect 520 -951 620 -860
rect 112 -978 837 -951
rect 112 -983 762 -978
rect 112 -1029 130 -983
rect 176 -1024 762 -983
rect 808 -1024 837 -978
rect 176 -1029 837 -1024
rect 112 -1051 837 -1029
rect 1532 -1050 1632 -871
rect 1736 -1050 1836 -872
rect 112 -1151 212 -1051
rect 724 -1146 824 -1051
rect 1328 -1078 2057 -1050
rect 1328 -1081 1973 -1078
rect 1328 -1127 1346 -1081
rect 1392 -1124 1973 -1081
rect 2019 -1124 2057 -1078
rect 1392 -1127 2057 -1124
rect 1328 -1150 2057 -1127
rect 1328 -1169 2040 -1150
rect 1328 -1346 1428 -1169
rect 1940 -1344 2040 -1169
<< polycontact >>
rect 1328 544 1374 590
rect 1989 543 2035 589
rect 174 347 220 393
rect 320 348 366 394
rect 1332 3 1378 49
rect 2003 2 2049 48
rect 130 -103 176 -57
rect 764 -105 810 -59
rect 132 -550 178 -504
rect 762 -556 808 -510
rect 1327 -518 1373 -472
rect 2037 -517 2083 -471
rect 130 -1029 176 -983
rect 762 -1024 808 -978
rect 1346 -1127 1392 -1081
rect 1973 -1124 2019 -1078
<< metal1 >>
rect 1312 595 1389 607
rect 1312 540 1324 595
rect 1377 540 1389 595
rect 1312 528 1389 540
rect 1973 594 2050 606
rect 1973 539 1985 594
rect 2038 539 2050 594
rect 1973 527 2050 539
rect 158 398 235 410
rect 158 343 170 398
rect 223 343 235 398
rect 158 331 235 343
rect 304 399 381 411
rect 304 344 316 399
rect 369 344 381 399
rect 304 332 381 344
rect 1253 390 2115 436
rect 37 238 900 284
rect 37 70 83 238
rect 241 20 287 186
rect 649 185 650 186
rect 430 165 507 177
rect 430 113 442 165
rect 495 113 507 165
rect 430 101 507 113
rect 445 81 491 101
rect 649 20 696 185
rect 854 173 900 238
rect 1253 216 1299 390
rect 839 161 916 173
rect 839 109 851 161
rect 904 109 916 161
rect 839 97 916 109
rect 1457 164 1503 332
rect 1646 315 1723 332
rect 1646 263 1658 315
rect 1711 263 1723 315
rect 1646 251 1723 263
rect 1865 164 1911 332
rect 2061 325 2115 390
rect 2050 313 2127 325
rect 2050 261 2062 313
rect 2115 261 2127 313
rect 2050 249 2127 261
rect 2061 216 2115 249
rect 1457 118 1911 164
rect 854 76 900 97
rect 241 -26 696 20
rect 1316 54 1393 66
rect 1316 -1 1328 54
rect 1381 -1 1393 54
rect 1316 -13 1393 -1
rect 114 -52 191 -40
rect 114 -107 126 -52
rect 179 -107 191 -52
rect 114 -119 191 -107
rect 35 -242 81 -237
rect 21 -254 98 -242
rect 21 -306 33 -254
rect 86 -306 98 -254
rect 21 -318 98 -306
rect 35 -384 81 -318
rect -26 -430 81 -384
rect 241 -399 287 -26
rect 429 -264 506 -252
rect 429 -316 441 -264
rect 494 -316 506 -264
rect 429 -328 506 -316
rect 649 -399 696 -26
rect 748 -54 825 -42
rect 748 -109 760 -54
rect 813 -109 825 -54
rect 748 -121 825 -109
rect 1250 -177 1296 -173
rect 1238 -189 1315 -177
rect 854 -253 900 -233
rect 1238 -241 1250 -189
rect 1303 -241 1315 -189
rect 1238 -253 1315 -241
rect 839 -265 916 -253
rect 839 -317 851 -265
rect 904 -317 916 -265
rect 839 -329 916 -317
rect 1250 -324 1296 -253
rect -26 -625 20 -430
rect 241 -445 696 -399
rect 854 -387 900 -329
rect 1201 -370 1296 -324
rect 1457 -358 1503 118
rect 1646 -182 1723 -170
rect 1646 -234 1658 -182
rect 1711 -234 1723 -182
rect 1646 -246 1723 -234
rect 1865 -358 1911 118
rect 1987 53 2064 65
rect 1987 -2 1999 53
rect 2052 -2 2064 53
rect 1987 -14 2064 -2
rect 2053 -173 2130 -161
rect 2053 -225 2065 -173
rect 2118 -225 2130 -173
rect 2053 -237 2130 -225
rect 854 -433 958 -387
rect 116 -499 193 -487
rect 116 -554 128 -499
rect 181 -554 193 -499
rect 116 -566 193 -554
rect -26 -671 83 -625
rect 37 -724 83 -671
rect 19 -736 97 -724
rect 19 -790 31 -736
rect 85 -790 97 -736
rect 19 -802 97 -790
rect 37 -820 83 -802
rect 114 -978 191 -966
rect 114 -1033 126 -978
rect 179 -1033 191 -978
rect 114 -1045 191 -1033
rect 37 -1351 83 -1186
rect 241 -1299 287 -445
rect 429 -737 507 -725
rect 429 -791 441 -737
rect 495 -791 507 -737
rect 429 -803 507 -791
rect 411 -1215 482 -1203
rect 411 -1269 423 -1215
rect 477 -1269 482 -1215
rect 411 -1281 482 -1269
rect 649 -1293 696 -445
rect 746 -505 823 -493
rect 746 -560 758 -505
rect 811 -560 823 -505
rect 746 -572 823 -560
rect 912 -627 958 -433
rect 853 -673 958 -627
rect 1201 -649 1247 -370
rect 1457 -404 1911 -358
rect 2072 -343 2118 -237
rect 2072 -389 2199 -343
rect 1311 -467 1388 -455
rect 1311 -522 1323 -467
rect 1376 -522 1388 -467
rect 1311 -534 1388 -522
rect 853 -820 899 -673
rect 1201 -695 1299 -649
rect 1253 -744 1299 -695
rect 1238 -756 1315 -744
rect 1238 -808 1250 -756
rect 1303 -808 1315 -756
rect 1238 -820 1315 -808
rect 1253 -828 1299 -820
rect 746 -973 823 -961
rect 746 -1028 758 -973
rect 811 -1028 823 -973
rect 746 -1040 823 -1028
rect 1330 -1076 1407 -1064
rect 1330 -1131 1342 -1076
rect 1395 -1131 1407 -1076
rect 1330 -1143 1407 -1131
rect 853 -1197 899 -1186
rect 839 -1209 915 -1197
rect 839 -1262 851 -1209
rect 903 -1262 915 -1209
rect 839 -1274 915 -1262
rect 853 -1351 899 -1274
rect 37 -1397 908 -1351
rect 8 -1481 930 -1453
rect 8 -1541 84 -1481
rect 144 -1482 930 -1481
rect 144 -1541 229 -1482
rect 8 -1542 229 -1541
rect 289 -1492 930 -1482
rect 289 -1538 418 -1492
rect 464 -1538 930 -1492
rect 289 -1542 930 -1538
rect 8 -1575 930 -1542
rect 1253 -1559 1299 -1375
rect 1457 -1485 1503 -404
rect 1645 -733 1722 -721
rect 1645 -785 1657 -733
rect 1710 -785 1722 -733
rect 1645 -797 1722 -785
rect 1645 -1394 1722 -1382
rect 1645 -1446 1657 -1394
rect 1710 -1446 1722 -1394
rect 1645 -1458 1722 -1446
rect 1865 -1486 1911 -404
rect 2021 -466 2098 -454
rect 2021 -521 2033 -466
rect 2086 -521 2098 -466
rect 2021 -533 2098 -521
rect 2153 -598 2199 -389
rect 2069 -644 2199 -598
rect 2069 -828 2115 -644
rect 1957 -1073 2034 -1061
rect 1957 -1128 1969 -1073
rect 2022 -1128 2034 -1073
rect 1957 -1140 2034 -1128
rect 2070 -1389 2123 -1375
rect 2054 -1401 2125 -1389
rect 2054 -1453 2066 -1401
rect 2119 -1453 2125 -1401
rect 2054 -1465 2125 -1453
rect 2070 -1559 2123 -1465
rect 1253 -1605 2123 -1559
<< via1 >>
rect 1324 590 1377 595
rect 1324 544 1328 590
rect 1328 544 1374 590
rect 1374 544 1377 590
rect 1324 540 1377 544
rect 1985 589 2038 594
rect 1985 543 1989 589
rect 1989 543 2035 589
rect 2035 543 2038 589
rect 1985 539 2038 543
rect 170 393 223 398
rect 170 347 174 393
rect 174 347 220 393
rect 220 347 223 393
rect 170 343 223 347
rect 316 394 369 399
rect 316 348 320 394
rect 320 348 366 394
rect 366 348 369 394
rect 316 344 369 348
rect 442 113 495 165
rect 851 109 904 161
rect 1658 263 1711 315
rect 2062 261 2115 313
rect 1328 49 1381 54
rect 1328 3 1332 49
rect 1332 3 1378 49
rect 1378 3 1381 49
rect 1328 -1 1381 3
rect 126 -57 179 -52
rect 126 -103 130 -57
rect 130 -103 176 -57
rect 176 -103 179 -57
rect 126 -107 179 -103
rect 33 -306 86 -254
rect 441 -316 494 -264
rect 760 -59 813 -54
rect 760 -105 764 -59
rect 764 -105 810 -59
rect 810 -105 813 -59
rect 760 -109 813 -105
rect 1250 -241 1303 -189
rect 851 -317 904 -265
rect 1658 -234 1711 -182
rect 1999 48 2052 53
rect 1999 2 2003 48
rect 2003 2 2049 48
rect 2049 2 2052 48
rect 1999 -2 2052 2
rect 2065 -225 2118 -173
rect 128 -504 181 -499
rect 128 -550 132 -504
rect 132 -550 178 -504
rect 178 -550 181 -504
rect 128 -554 181 -550
rect 31 -790 85 -736
rect 126 -983 179 -978
rect 126 -1029 130 -983
rect 130 -1029 176 -983
rect 176 -1029 179 -983
rect 126 -1033 179 -1029
rect 441 -791 495 -737
rect 423 -1269 477 -1215
rect 758 -510 811 -505
rect 758 -556 762 -510
rect 762 -556 808 -510
rect 808 -556 811 -510
rect 758 -560 811 -556
rect 1323 -472 1376 -467
rect 1323 -518 1327 -472
rect 1327 -518 1373 -472
rect 1373 -518 1376 -472
rect 1323 -522 1376 -518
rect 1250 -808 1303 -756
rect 758 -978 811 -973
rect 758 -1024 762 -978
rect 762 -1024 808 -978
rect 808 -1024 811 -978
rect 758 -1028 811 -1024
rect 1342 -1081 1395 -1076
rect 1342 -1127 1346 -1081
rect 1346 -1127 1392 -1081
rect 1392 -1127 1395 -1081
rect 1342 -1131 1395 -1127
rect 851 -1262 903 -1209
rect 84 -1541 144 -1481
rect 229 -1542 289 -1482
rect 1657 -785 1710 -733
rect 1657 -1446 1710 -1394
rect 2033 -471 2086 -466
rect 2033 -517 2037 -471
rect 2037 -517 2083 -471
rect 2083 -517 2086 -471
rect 2033 -521 2086 -517
rect 1969 -1078 2022 -1073
rect 1969 -1124 1973 -1078
rect 1973 -1124 2019 -1078
rect 2019 -1124 2022 -1078
rect 1969 -1128 2022 -1124
rect 2066 -1453 2119 -1401
<< metal2 >>
rect 1312 596 1389 607
rect 1312 539 1322 596
rect 1378 539 1389 596
rect 1312 528 1389 539
rect 1973 595 2050 606
rect 1973 538 1983 595
rect 2039 538 2050 595
rect 1973 527 2050 538
rect 158 399 235 410
rect 158 342 168 399
rect 224 342 235 399
rect 158 331 235 342
rect 304 400 381 411
rect 304 343 314 400
rect 370 343 381 400
rect 304 332 381 343
rect 1655 400 2248 456
rect 1655 332 1711 400
rect 1646 323 1723 332
rect 1522 315 1724 323
rect 437 242 1050 299
rect 437 177 494 242
rect 430 170 507 177
rect 291 165 507 170
rect 839 168 916 173
rect 291 113 442 165
rect 495 113 507 165
rect 114 -51 191 -40
rect 114 -108 124 -51
rect 180 -108 191 -51
rect 114 -119 191 -108
rect 21 -249 98 -242
rect 291 -249 348 113
rect 430 101 507 113
rect 563 161 916 168
rect 563 110 851 161
rect 21 -254 348 -249
rect 563 -252 621 110
rect 839 109 851 110
rect 904 109 916 161
rect 839 97 916 109
rect 748 -53 825 -42
rect 748 -110 758 -53
rect 814 -110 825 -53
rect 748 -121 825 -110
rect 21 -306 33 -254
rect 86 -306 348 -254
rect 429 -264 621 -252
rect 21 -318 98 -306
rect 429 -316 441 -264
rect 494 -316 621 -264
rect 429 -319 621 -316
rect 839 -262 916 -253
rect 993 -262 1050 242
rect 1522 267 1658 315
rect 1316 55 1393 66
rect 1316 -2 1326 55
rect 1382 -2 1393 55
rect 1316 -13 1393 -2
rect 1238 -185 1315 -177
rect 1522 -185 1578 267
rect 1646 263 1658 267
rect 1711 267 1724 315
rect 2050 313 2127 325
rect 2050 307 2062 313
rect 1711 263 1723 267
rect 1646 251 1723 263
rect 1781 261 2062 307
rect 2115 261 2127 313
rect 1781 249 2127 261
rect 1781 242 2111 249
rect 1238 -189 1578 -185
rect 1238 -241 1250 -189
rect 1303 -241 1578 -189
rect 1646 -179 1723 -170
rect 1781 -179 1837 242
rect 1987 54 2064 65
rect 1987 -3 1997 54
rect 2053 -3 2064 54
rect 1987 -14 2064 -3
rect 1646 -182 1837 -179
rect 1646 -234 1658 -182
rect 1711 -234 1837 -182
rect 1646 -241 1837 -234
rect 2053 -173 2130 -161
rect 2192 -173 2248 400
rect 2053 -225 2065 -173
rect 2118 -225 2248 -173
rect 2053 -229 2248 -225
rect 2053 -237 2130 -229
rect 1238 -253 1315 -241
rect 1646 -246 1723 -241
rect 839 -265 1050 -262
rect 839 -317 851 -265
rect 904 -317 1050 -265
rect 839 -319 1050 -317
rect 429 -328 506 -319
rect 116 -498 193 -487
rect 116 -555 126 -498
rect 182 -555 193 -498
rect 116 -566 193 -555
rect 23 -724 83 -723
rect 19 -736 97 -724
rect 440 -725 497 -328
rect 839 -329 916 -319
rect 1311 -466 1388 -455
rect 746 -504 823 -493
rect 746 -561 756 -504
rect 812 -561 823 -504
rect 1311 -523 1321 -466
rect 1377 -523 1388 -466
rect 1311 -534 1388 -523
rect 746 -572 823 -561
rect 1653 -721 1709 -246
rect 2021 -465 2098 -454
rect 2021 -522 2031 -465
rect 2087 -522 2098 -465
rect 2021 -533 2098 -522
rect 1645 -722 1722 -721
rect 19 -790 31 -736
rect 85 -790 97 -736
rect 19 -802 97 -790
rect 429 -737 507 -725
rect 429 -791 441 -737
rect 495 -791 507 -737
rect 1645 -733 1725 -722
rect 19 -833 83 -802
rect 429 -803 507 -791
rect 1238 -756 1315 -744
rect -69 -893 83 -833
rect -69 -1216 -9 -893
rect 114 -977 191 -966
rect 114 -1034 124 -977
rect 180 -1034 191 -977
rect 114 -1045 191 -1034
rect 433 -988 491 -803
rect 1238 -808 1250 -756
rect 1303 -808 1315 -756
rect 1645 -785 1657 -733
rect 1710 -785 1725 -733
rect 1645 -797 1725 -785
rect 1238 -820 1315 -808
rect 1238 -867 1305 -820
rect 1147 -923 1305 -867
rect 746 -972 823 -961
rect 433 -1046 604 -988
rect 746 -1029 756 -972
rect 812 -1029 823 -972
rect 746 -1040 823 -1029
rect 411 -1215 482 -1203
rect 411 -1216 423 -1215
rect -69 -1269 423 -1216
rect 477 -1216 482 -1215
rect 546 -1208 604 -1046
rect 839 -1208 915 -1197
rect 546 -1209 915 -1208
rect 477 -1269 485 -1216
rect 546 -1262 851 -1209
rect 903 -1262 915 -1209
rect 546 -1266 915 -1262
rect -69 -1276 485 -1269
rect 839 -1274 915 -1266
rect -69 -1482 -9 -1276
rect 411 -1281 482 -1276
rect 1147 -1380 1203 -923
rect 1330 -1075 1407 -1064
rect 1330 -1132 1340 -1075
rect 1396 -1132 1407 -1075
rect 1330 -1143 1407 -1132
rect 1653 -1084 1725 -797
rect 1957 -1072 2034 -1061
rect 1653 -1156 1841 -1084
rect 1957 -1129 1967 -1072
rect 2023 -1129 2034 -1072
rect 1957 -1140 2034 -1129
rect 1777 -1181 1841 -1156
rect 1147 -1382 1711 -1380
rect 1147 -1394 1722 -1382
rect 1147 -1436 1657 -1394
rect 1645 -1446 1657 -1436
rect 1710 -1446 1722 -1394
rect 1645 -1458 1722 -1446
rect 1778 -1389 1841 -1181
rect 1778 -1401 2126 -1389
rect 1778 -1453 2066 -1401
rect 2119 -1453 2126 -1401
rect 1778 -1461 2126 -1453
rect 2054 -1465 2125 -1461
rect 66 -1481 303 -1469
rect 66 -1482 84 -1481
rect -69 -1541 84 -1482
rect 144 -1482 303 -1481
rect 144 -1541 229 -1482
rect -69 -1542 229 -1541
rect 289 -1542 303 -1482
rect 66 -1562 303 -1542
<< via2 >>
rect 1322 595 1378 596
rect 1322 540 1324 595
rect 1324 540 1377 595
rect 1377 540 1378 595
rect 1322 539 1378 540
rect 1983 594 2039 595
rect 1983 539 1985 594
rect 1985 539 2038 594
rect 2038 539 2039 594
rect 1983 538 2039 539
rect 168 398 224 399
rect 168 343 170 398
rect 170 343 223 398
rect 223 343 224 398
rect 168 342 224 343
rect 314 399 370 400
rect 314 344 316 399
rect 316 344 369 399
rect 369 344 370 399
rect 314 343 370 344
rect 124 -52 180 -51
rect 124 -107 126 -52
rect 126 -107 179 -52
rect 179 -107 180 -52
rect 124 -108 180 -107
rect 758 -54 814 -53
rect 758 -109 760 -54
rect 760 -109 813 -54
rect 813 -109 814 -54
rect 758 -110 814 -109
rect 1326 54 1382 55
rect 1326 -1 1328 54
rect 1328 -1 1381 54
rect 1381 -1 1382 54
rect 1326 -2 1382 -1
rect 1997 53 2053 54
rect 1997 -2 1999 53
rect 1999 -2 2052 53
rect 2052 -2 2053 53
rect 1997 -3 2053 -2
rect 126 -499 182 -498
rect 126 -554 128 -499
rect 128 -554 181 -499
rect 181 -554 182 -499
rect 126 -555 182 -554
rect 756 -505 812 -504
rect 756 -560 758 -505
rect 758 -560 811 -505
rect 811 -560 812 -505
rect 756 -561 812 -560
rect 1321 -467 1377 -466
rect 1321 -522 1323 -467
rect 1323 -522 1376 -467
rect 1376 -522 1377 -467
rect 1321 -523 1377 -522
rect 2031 -466 2087 -465
rect 2031 -521 2033 -466
rect 2033 -521 2086 -466
rect 2086 -521 2087 -466
rect 2031 -522 2087 -521
rect 124 -978 180 -977
rect 124 -1033 126 -978
rect 126 -1033 179 -978
rect 179 -1033 180 -978
rect 124 -1034 180 -1033
rect 756 -973 812 -972
rect 756 -1028 758 -973
rect 758 -1028 811 -973
rect 811 -1028 812 -973
rect 756 -1029 812 -1028
rect 1340 -1076 1396 -1075
rect 1340 -1131 1342 -1076
rect 1342 -1131 1395 -1076
rect 1395 -1131 1396 -1076
rect 1340 -1132 1396 -1131
rect 1967 -1073 2023 -1072
rect 1967 -1128 1969 -1073
rect 1969 -1128 2022 -1073
rect 2022 -1128 2023 -1073
rect 1967 -1129 2023 -1128
<< metal3 >>
rect 1301 596 2085 617
rect 1301 539 1322 596
rect 1378 595 2085 596
rect 1378 539 1983 595
rect 1301 538 1983 539
rect 2039 538 2085 595
rect 1301 517 2085 538
rect 95 400 821 413
rect 95 399 314 400
rect 95 342 168 399
rect 224 343 314 399
rect 370 398 821 400
rect 370 343 1071 398
rect 224 342 1071 343
rect 95 340 1071 342
rect 95 319 821 340
rect 108 -43 834 -29
rect -151 -51 834 -43
rect -151 -108 124 -51
rect 180 -53 834 -51
rect 180 -108 758 -53
rect -151 -110 758 -108
rect 814 -110 834 -53
rect -151 -120 834 -110
rect -151 -959 -74 -120
rect 108 -123 834 -120
rect 110 -498 836 -480
rect 110 -555 126 -498
rect 182 -504 836 -498
rect 182 -555 756 -504
rect 110 -561 756 -555
rect 812 -509 836 -504
rect 1013 -509 1071 340
rect 1300 55 2089 85
rect 1300 -2 1326 55
rect 1382 54 2089 55
rect 1382 -2 1997 54
rect 1300 -3 1997 -2
rect 2053 -3 2089 54
rect 1300 -25 2089 -3
rect 812 -561 1071 -509
rect 1305 -465 2104 -439
rect 1305 -466 2031 -465
rect 1305 -523 1321 -466
rect 1377 -522 2031 -466
rect 2087 -522 2104 -465
rect 1377 -523 2104 -522
rect 1305 -550 2104 -523
rect 110 -567 1071 -561
rect 110 -574 836 -567
rect 112 -959 839 -951
rect -151 -972 839 -959
rect -151 -977 756 -972
rect -151 -1034 124 -977
rect 180 -1029 756 -977
rect 812 -1029 839 -972
rect 180 -1034 839 -1029
rect -151 -1036 839 -1034
rect 112 -1051 839 -1036
rect 1321 -1072 2060 -1046
rect 1321 -1075 1967 -1072
rect 1321 -1132 1340 -1075
rect 1396 -1129 1967 -1075
rect 2023 -1129 2060 -1072
rect 1396 -1132 2060 -1129
rect 1321 -1181 2060 -1132
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_0
timestamp 1693898385
transform 1 0 774 0 1 -291
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_1
timestamp 1693898385
transform 1 0 162 0 1 -291
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_2
timestamp 1693898385
transform 1 0 366 0 1 -291
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_3
timestamp 1693898385
transform 1 0 570 0 1 -291
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_4
timestamp 1693898385
transform 1 0 774 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_5
timestamp 1693898385
transform 1 0 570 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_6
timestamp 1693898385
transform 1 0 366 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_7
timestamp 1693898385
transform 1 0 162 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_8
timestamp 1693898385
transform 1 0 774 0 1 -1244
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_9
timestamp 1693898385
transform 1 0 570 0 1 -1244
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_10
timestamp 1693898385
transform 1 0 366 0 1 -1244
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_11
timestamp 1693898385
transform 1 0 162 0 1 -1244
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_12
timestamp 1693898385
transform 1 0 774 0 1 -762
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_13
timestamp 1693898385
transform 1 0 570 0 1 -762
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_14
timestamp 1693898385
transform 1 0 366 0 1 -762
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_15
timestamp 1693898385
transform 1 0 162 0 1 -762
box -162 -128 162 128
use pmos_3p3_K82TLM  pmos_3p3_K82TLM_0
timestamp 1693898385
transform 1 0 1990 0 1 274
box -224 -190 224 190
use pmos_3p3_K82TLM  pmos_3p3_K82TLM_1
timestamp 1693898385
transform 1 0 1786 0 1 274
box -224 -190 224 190
use pmos_3p3_K82TLM  pmos_3p3_K82TLM_2
timestamp 1693898385
transform 1 0 1582 0 1 -220
box -224 -190 224 190
use pmos_3p3_K82TLM  pmos_3p3_K82TLM_3
timestamp 1693898385
transform 1 0 1582 0 1 274
box -224 -190 224 190
use pmos_3p3_K82TLM  pmos_3p3_K82TLM_4
timestamp 1693898385
transform 1 0 1378 0 1 -220
box -224 -190 224 190
use pmos_3p3_K82TLM  pmos_3p3_K82TLM_5
timestamp 1693898385
transform 1 0 1786 0 1 -220
box -224 -190 224 190
use pmos_3p3_K82TLM  pmos_3p3_K82TLM_6
timestamp 1693898385
transform 1 0 1990 0 1 -220
box -224 -190 224 190
use pmos_3p3_K82TLM  pmos_3p3_K82TLM_7
timestamp 1693898385
transform 1 0 1378 0 1 274
box -224 -190 224 190
use pmos_3p3_K82TLM  pmos_3p3_K82TLM_8
timestamp 1693898385
transform 1 0 1786 0 1 -1433
box -224 -190 224 190
use pmos_3p3_K82TLM  pmos_3p3_K82TLM_9
timestamp 1693898385
transform 1 0 1582 0 1 -770
box -224 -190 224 190
use pmos_3p3_K82TLM  pmos_3p3_K82TLM_10
timestamp 1693898385
transform 1 0 1378 0 1 -770
box -224 -190 224 190
use pmos_3p3_K82TLM  pmos_3p3_K82TLM_11
timestamp 1693898385
transform 1 0 1990 0 1 -770
box -224 -190 224 190
use pmos_3p3_K82TLM  pmos_3p3_K82TLM_12
timestamp 1693898385
transform 1 0 1582 0 1 -1433
box -224 -190 224 190
use pmos_3p3_K82TLM  pmos_3p3_K82TLM_13
timestamp 1693898385
transform 1 0 1378 0 1 -1433
box -224 -190 224 190
use pmos_3p3_K82TLM  pmos_3p3_K82TLM_14
timestamp 1693898385
transform 1 0 1990 0 1 -1433
box -224 -190 224 190
use pmos_3p3_K82TLM  pmos_3p3_K82TLM_15
timestamp 1693898385
transform 1 0 1786 0 1 -770
box -224 -190 224 190
<< end >>
