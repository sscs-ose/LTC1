magic
tech gf180mcuC
magscale 1 10
timestamp 1692792393
<< nwell >>
rect -2144 -3292 -1740 -2870
rect -1608 -3292 -784 -2870
rect -2144 -3311 -1940 -3292
rect -2144 -4160 -1740 -3738
rect -1608 -4160 -784 -3738
rect -2144 -4179 -1940 -4160
rect -2144 -5019 -1740 -4597
rect -1608 -5019 -784 -4597
rect -2144 -5038 -1940 -5019
rect -2144 -5887 -1740 -5465
rect -1608 -5887 -784 -5465
rect -526 -5887 -122 -5465
rect 10 -5887 834 -5465
rect 1083 -5887 1487 -5465
rect 1619 -5887 2443 -5465
rect -2144 -5906 -1940 -5887
rect -526 -5906 -322 -5887
rect 1083 -5906 1287 -5887
<< pwell >>
rect -1796 1418 2356 1674
rect 3119 1645 3133 1724
rect 3119 1635 3135 1645
rect 3938 1635 3986 1752
rect 3004 1433 4440 1635
rect 3461 1372 3556 1433
rect -1796 1115 2356 1371
rect 3012 1116 4484 1372
rect 4679 1367 6115 1569
rect 5093 1327 5130 1337
rect 5684 1327 5742 1367
rect 5811 1327 6081 1367
rect 4679 1125 6115 1327
rect 4167 1104 4275 1116
rect 4248 1070 4272 1071
rect 5688 1064 5690 1123
rect 5753 1046 5853 1125
rect -1796 676 2356 932
rect 3004 805 4568 1007
rect 4380 775 4452 805
rect 4825 790 5965 1046
rect 3086 470 4634 726
rect 4825 488 5965 744
rect -1796 0 2356 256
rect 3446 222 3751 258
rect 3446 202 3546 222
rect 3650 202 3750 222
rect 1343 -70 1599 0
rect 2926 -54 4270 202
rect 4393 -33 5829 169
rect -1796 -325 2356 -70
rect 3650 -148 3750 -54
rect -1796 -326 -860 -325
rect -852 -326 2356 -325
rect 2926 -432 4270 -176
rect 4392 -349 5828 -147
rect 3446 -455 3546 -432
rect 3650 -455 3750 -432
rect 3854 -455 3954 -432
rect 2926 -711 4270 -455
rect 4392 -486 5828 -397
rect 4392 -599 4724 -486
rect 4732 -599 5276 -486
rect 5284 -599 5828 -486
rect 4392 -742 4724 -722
rect 4732 -742 5276 -722
rect 5284 -742 5828 -722
rect -1796 -1118 2356 -862
rect 2926 -1089 4270 -833
rect 4392 -924 5828 -742
rect 3634 -1094 3651 -1089
rect -481 -1293 -381 -1244
rect 335 -1293 435 -1244
rect 947 -1293 1047 -1244
rect 1151 -1293 1251 -1244
rect 1763 -1293 1863 -1244
rect -1796 -1549 2356 -1293
rect 539 -1603 639 -1549
rect 743 -1603 843 -1549
rect 947 -1603 1047 -1549
rect 1151 -1603 1251 -1549
rect 1559 -1603 1659 -1549
rect 1763 -1603 1863 -1549
rect -1796 -1859 2356 -1603
rect 3589 -1838 3689 -1770
rect 3793 -1814 5834 -1734
rect 5937 -1838 6037 -1783
rect 3477 -2094 6149 -1838
rect 3477 -2478 6149 -2222
rect 4125 -2512 4429 -2478
rect 4661 -2512 4761 -2478
rect 4865 -2512 4965 -2478
rect 5197 -2512 5501 -2478
rect 5733 -2512 5833 -2478
rect 5937 -2512 6037 -2478
rect 3477 -2513 5613 -2512
rect 5621 -2513 6149 -2512
rect 3477 -2768 6149 -2513
rect 5613 -2769 5621 -2768
rect -91 -3077 2581 -2821
rect 556 -3105 860 -3077
rect 1628 -3105 1932 -3077
rect 2165 -3105 2265 -3077
rect -2086 -3535 -1798 -3337
rect -1608 -3535 -1320 -3341
rect -1072 -3535 -784 -3341
rect -91 -3361 437 -3105
rect 445 -3361 973 -3105
rect 981 -3361 1509 -3105
rect 1517 -3361 2045 -3105
rect 2053 -3361 2581 -3105
rect 3477 -3152 6149 -2896
rect 5751 -3165 5827 -3152
rect -91 -3893 2605 -3637
rect 3477 -3786 5637 -3530
rect 5645 -3786 6173 -3530
rect -2086 -4403 -1798 -4205
rect -1608 -4403 -1320 -4209
rect -1072 -4403 -784 -4209
rect -91 -4282 2605 -4026
rect 3477 -4175 5637 -3919
rect 5645 -4175 6173 -3919
rect 4512 -4214 4614 -4175
rect 5003 -4214 5006 -4213
rect 5961 -4214 6061 -4175
rect -91 -4577 2605 -4321
rect 3477 -4470 5637 -4214
rect 5645 -4470 6173 -4214
rect -91 -4962 2605 -4706
rect 3477 -4855 5637 -4599
rect 5645 -4855 6173 -4599
rect 557 -5004 559 -4962
rect -2086 -5262 -1798 -5064
rect -1608 -5262 -1320 -5068
rect -1072 -5262 -784 -5068
rect 3477 -5182 5637 -4926
rect 5645 -5182 6173 -4926
rect 3477 -5571 5637 -5315
rect 5645 -5571 6173 -5315
rect 3477 -5866 5637 -5610
rect 5645 -5866 6173 -5610
rect -2086 -6130 -1798 -5932
rect -1608 -6130 -1320 -5936
rect -1072 -6130 -784 -5936
rect -468 -6130 -180 -5932
rect 10 -6130 298 -5936
rect 546 -6130 834 -5936
rect 1141 -6130 1429 -5932
rect 1619 -6130 1907 -5936
rect 2155 -6130 2443 -5936
rect 3477 -6251 5637 -5995
rect 5645 -6251 6173 -5995
<< nmos >>
rect -1684 1486 -1584 1606
rect -1297 1486 -1197 1606
rect -1093 1486 -993 1606
rect -889 1486 -789 1606
rect -685 1486 -585 1606
rect -481 1486 -381 1606
rect -277 1486 -177 1606
rect -73 1486 27 1606
rect 131 1486 231 1606
rect 335 1486 435 1606
rect 539 1486 639 1606
rect 743 1486 843 1606
rect 947 1486 1047 1606
rect 1151 1486 1251 1606
rect 1355 1486 1455 1606
rect 1559 1486 1659 1606
rect 1763 1486 1863 1606
rect 2144 1486 2244 1606
rect 3120 1504 3220 1564
rect 3460 1504 3560 1564
rect 3800 1504 3900 1564
rect 4012 1504 4112 1564
rect 4224 1504 4324 1564
rect -1684 1183 -1584 1303
rect -1297 1183 -1197 1303
rect -1093 1183 -993 1303
rect -889 1183 -789 1303
rect -685 1183 -585 1303
rect -481 1183 -381 1303
rect -277 1183 -177 1303
rect -73 1183 27 1303
rect 131 1183 231 1303
rect 335 1183 435 1303
rect 539 1183 639 1303
rect 743 1183 843 1303
rect 947 1183 1047 1303
rect 1151 1183 1251 1303
rect 1355 1183 1455 1303
rect 1559 1183 1659 1303
rect 1763 1183 1863 1303
rect 2144 1183 2244 1303
rect 4795 1438 4895 1498
rect 5007 1438 5107 1498
rect 3124 1184 3224 1304
rect 3456 1184 3556 1304
rect 3660 1184 3760 1304
rect 3864 1184 3964 1304
rect 4068 1184 4168 1304
rect 4272 1184 4372 1304
rect 5347 1438 5447 1498
rect 5559 1438 5659 1498
rect 4795 1196 4895 1256
rect 5007 1196 5107 1256
rect 5899 1438 5999 1498
rect 5347 1196 5447 1256
rect 5559 1196 5659 1256
rect 3120 876 3220 936
rect -1684 744 -1584 864
rect -1297 744 -1197 864
rect -1093 744 -993 864
rect -889 744 -789 864
rect -685 744 -585 864
rect -481 744 -381 864
rect -277 744 -177 864
rect -73 744 27 864
rect 131 744 231 864
rect 335 744 435 864
rect 539 744 639 864
rect 743 744 843 864
rect 947 744 1047 864
rect 1151 744 1251 864
rect 1355 744 1455 864
rect 1559 744 1659 864
rect 1763 744 1863 864
rect 2144 744 2244 864
rect 3460 876 3560 936
rect 3800 876 3900 936
rect 4012 876 4112 936
rect 5899 1196 5999 1256
rect 4352 876 4452 936
rect 4937 858 5037 978
rect 5141 858 5241 978
rect 5345 858 5445 978
rect 5549 858 5649 978
rect 5753 858 5853 978
rect 3198 538 3298 658
rect 3402 538 3502 658
rect 3606 538 3706 658
rect 3810 538 3910 658
rect 4014 538 4114 658
rect 4218 538 4318 658
rect 4422 538 4522 658
rect 4937 556 5037 676
rect 5141 556 5241 676
rect 5345 556 5445 676
rect 5549 556 5649 676
rect 5753 556 5853 676
rect -1684 68 -1584 188
rect -1480 68 -1380 188
rect -1276 68 -1176 188
rect -1072 68 -972 188
rect -740 68 -640 188
rect -536 68 -436 188
rect -204 68 -104 188
rect 128 68 228 188
rect 332 68 432 188
rect 664 68 764 188
rect 996 68 1096 188
rect 1200 68 1300 188
rect 1532 68 1632 188
rect 1736 68 1836 188
rect 1940 68 2040 188
rect 2144 68 2244 188
rect 3038 14 3138 134
rect 3242 14 3342 134
rect 3446 14 3546 134
rect 3650 14 3750 134
rect 3854 14 3954 134
rect 4058 14 4158 134
rect 4509 38 4609 98
rect -1684 -258 -1584 -138
rect -1480 -258 -1380 -138
rect -1276 -258 -1176 -138
rect -1072 -258 -972 -138
rect -740 -258 -640 -138
rect -536 -258 -436 -138
rect -204 -258 -104 -138
rect 128 -258 228 -138
rect 332 -258 432 -138
rect 664 -258 764 -138
rect 996 -258 1096 -138
rect 1200 -258 1300 -138
rect 1532 -258 1632 -138
rect 1736 -258 1836 -138
rect 1940 -258 2040 -138
rect 2144 -258 2244 -138
rect 4849 38 4949 98
rect 5061 38 5161 98
rect 5401 38 5501 98
rect 5613 38 5713 98
rect 3038 -364 3138 -244
rect 3242 -364 3342 -244
rect 3446 -364 3546 -244
rect 3650 -364 3750 -244
rect 3854 -364 3954 -244
rect 4058 -364 4158 -244
rect 4508 -278 4608 -218
rect 4848 -278 4948 -218
rect 5060 -278 5160 -218
rect 5400 -278 5500 -218
rect 5612 -278 5712 -218
rect 3038 -643 3138 -523
rect 3242 -643 3342 -523
rect 3446 -643 3546 -523
rect 3650 -643 3750 -523
rect 3854 -643 3954 -523
rect 4058 -643 4158 -523
rect 4508 -528 4608 -468
rect 4848 -528 4948 -468
rect 5060 -528 5160 -468
rect 5400 -528 5500 -468
rect 5612 -528 5712 -468
rect -1684 -1050 -1584 -930
rect -1297 -1050 -1197 -930
rect -1093 -1050 -993 -930
rect -889 -1050 -789 -930
rect -685 -1050 -585 -930
rect -481 -1050 -381 -930
rect -277 -1050 -177 -930
rect -73 -1050 27 -930
rect 131 -1050 231 -930
rect 335 -1050 435 -930
rect 539 -1050 639 -930
rect 743 -1050 843 -930
rect 947 -1050 1047 -930
rect 1151 -1050 1251 -930
rect 1355 -1050 1455 -930
rect 1559 -1050 1659 -930
rect 1763 -1050 1863 -930
rect 2144 -1050 2244 -930
rect 4508 -853 4608 -793
rect 3038 -1021 3138 -901
rect 3242 -1021 3342 -901
rect 3446 -1021 3546 -901
rect 3650 -1021 3750 -901
rect 3854 -1021 3954 -901
rect 4058 -1021 4158 -901
rect 4848 -853 4948 -793
rect 5060 -853 5160 -793
rect 5400 -853 5500 -793
rect 5612 -853 5712 -793
rect -1684 -1481 -1584 -1361
rect -1297 -1481 -1197 -1361
rect -1093 -1481 -993 -1361
rect -889 -1481 -789 -1361
rect -685 -1481 -585 -1361
rect -481 -1481 -381 -1361
rect -277 -1481 -177 -1361
rect -73 -1481 27 -1361
rect 131 -1481 231 -1361
rect 335 -1481 435 -1361
rect 539 -1481 639 -1361
rect 743 -1481 843 -1361
rect 947 -1481 1047 -1361
rect 1151 -1481 1251 -1361
rect 1355 -1481 1455 -1361
rect 1559 -1481 1659 -1361
rect 1763 -1481 1863 -1361
rect 2144 -1481 2244 -1361
rect -1684 -1791 -1584 -1671
rect -1297 -1791 -1197 -1671
rect -1093 -1791 -993 -1671
rect -889 -1791 -789 -1671
rect -685 -1791 -585 -1671
rect -481 -1791 -381 -1671
rect -277 -1791 -177 -1671
rect -73 -1791 27 -1671
rect 131 -1791 231 -1671
rect 335 -1791 435 -1671
rect 539 -1791 639 -1671
rect 743 -1791 843 -1671
rect 947 -1791 1047 -1671
rect 1151 -1791 1251 -1671
rect 1355 -1791 1455 -1671
rect 1559 -1791 1659 -1671
rect 1763 -1791 1863 -1671
rect 2144 -1791 2244 -1671
rect 3589 -2026 3689 -1906
rect 3793 -2026 3893 -1906
rect 4125 -2026 4225 -1906
rect 4329 -2026 4429 -1906
rect 4661 -2026 4761 -1906
rect 4865 -2026 4965 -1906
rect 5197 -2026 5297 -1906
rect 5401 -2026 5501 -1906
rect 5733 -2026 5833 -1906
rect 5937 -2026 6037 -1906
rect 3589 -2410 3689 -2290
rect 3793 -2410 3893 -2290
rect 4125 -2410 4225 -2290
rect 4329 -2410 4429 -2290
rect 4661 -2410 4761 -2290
rect 4865 -2410 4965 -2290
rect 5197 -2410 5297 -2290
rect 5401 -2410 5501 -2290
rect 5733 -2410 5833 -2290
rect 5937 -2410 6037 -2290
rect 21 -3009 121 -2889
rect 225 -3009 325 -2889
rect 557 -3009 657 -2889
rect 761 -3009 861 -2889
rect 1093 -3009 1193 -2889
rect 1297 -3009 1397 -2889
rect 1629 -3009 1729 -2889
rect 1833 -3009 1933 -2889
rect 2165 -3009 2265 -2889
rect 2369 -3009 2469 -2889
rect 21 -3293 121 -3173
rect 225 -3293 325 -3173
rect 557 -3293 657 -3173
rect 761 -3293 861 -3173
rect 1093 -3293 1193 -3173
rect 1297 -3293 1397 -3173
rect 1629 -3293 1729 -3173
rect 1833 -3293 1933 -3173
rect 2165 -3293 2265 -3173
rect 2369 -3293 2469 -3173
rect -1970 -3461 -1914 -3411
rect -1492 -3460 -1436 -3416
rect -956 -3460 -900 -3416
rect 21 -3825 121 -3705
rect 225 -3825 325 -3705
rect 429 -3825 529 -3705
rect 633 -3825 733 -3705
rect 837 -3825 937 -3705
rect 1041 -3825 1141 -3705
rect 1245 -3825 1345 -3705
rect 1449 -3825 1549 -3705
rect 1653 -3825 1753 -3705
rect 1857 -3825 1957 -3705
rect 2189 -3825 2289 -3705
rect 2393 -3825 2493 -3705
rect -1970 -4329 -1914 -4279
rect -1492 -4328 -1436 -4284
rect 21 -4214 121 -4094
rect 225 -4214 325 -4094
rect 429 -4214 529 -4094
rect 633 -4214 733 -4094
rect 837 -4214 937 -4094
rect 1041 -4214 1141 -4094
rect 1245 -4214 1345 -4094
rect 1449 -4214 1549 -4094
rect 1653 -4214 1753 -4094
rect 1857 -4214 1957 -4094
rect 2189 -4214 2289 -4094
rect 2393 -4214 2493 -4094
rect -956 -4328 -900 -4284
rect 21 -4509 121 -4389
rect 225 -4509 325 -4389
rect 429 -4509 529 -4389
rect 633 -4509 733 -4389
rect 837 -4509 937 -4389
rect 1041 -4509 1141 -4389
rect 1245 -4509 1345 -4389
rect 1449 -4509 1549 -4389
rect 1653 -4509 1753 -4389
rect 1857 -4509 1957 -4389
rect 2189 -4509 2289 -4389
rect 2393 -4509 2493 -4389
rect 21 -4894 121 -4774
rect 225 -4894 325 -4774
rect 429 -4894 529 -4774
rect 633 -4894 733 -4774
rect 837 -4894 937 -4774
rect 1041 -4894 1141 -4774
rect 1245 -4894 1345 -4774
rect 1449 -4894 1549 -4774
rect 1653 -4894 1753 -4774
rect 1857 -4894 1957 -4774
rect 2189 -4894 2289 -4774
rect 2393 -4894 2493 -4774
rect -1970 -5188 -1914 -5138
rect -1492 -5187 -1436 -5143
rect -956 -5187 -900 -5143
rect 3589 -2700 3689 -2580
rect 3793 -2700 3893 -2580
rect 4125 -2700 4225 -2580
rect 4329 -2700 4429 -2580
rect 4661 -2700 4761 -2580
rect 4865 -2700 4965 -2580
rect 5197 -2700 5297 -2580
rect 5401 -2700 5501 -2580
rect 5733 -2700 5833 -2580
rect 5937 -2700 6037 -2580
rect 3589 -3084 3689 -2964
rect 3793 -3084 3893 -2964
rect 4125 -3084 4225 -2964
rect 4329 -3084 4429 -2964
rect 4661 -3084 4761 -2964
rect 4865 -3084 4965 -2964
rect 5197 -3084 5297 -2964
rect 5401 -3084 5501 -2964
rect 5733 -3084 5833 -2964
rect 5937 -3084 6037 -2964
rect 3589 -3718 3689 -3598
rect 3793 -3718 3893 -3598
rect 3997 -3718 4097 -3598
rect 4201 -3718 4301 -3598
rect 4405 -3718 4505 -3598
rect 4609 -3718 4709 -3598
rect 4813 -3718 4913 -3598
rect 5017 -3718 5117 -3598
rect 5221 -3718 5321 -3598
rect 5425 -3718 5525 -3598
rect 5757 -3718 5857 -3598
rect 5961 -3718 6061 -3598
rect 3589 -4107 3689 -3987
rect 3793 -4107 3893 -3987
rect 3997 -4107 4097 -3987
rect 4201 -4107 4301 -3987
rect 4405 -4107 4505 -3987
rect 4609 -4107 4709 -3987
rect 4813 -4107 4913 -3987
rect 5017 -4107 5117 -3987
rect 5221 -4107 5321 -3987
rect 5425 -4107 5525 -3987
rect 5757 -4107 5857 -3987
rect 5961 -4107 6061 -3987
rect 3589 -4402 3689 -4282
rect 3793 -4402 3893 -4282
rect 3997 -4402 4097 -4282
rect 4201 -4402 4301 -4282
rect 4405 -4402 4505 -4282
rect 4609 -4402 4709 -4282
rect 4813 -4402 4913 -4282
rect 5017 -4402 5117 -4282
rect 5221 -4402 5321 -4282
rect 5425 -4402 5525 -4282
rect 5757 -4402 5857 -4282
rect 5961 -4402 6061 -4282
rect 3589 -4787 3689 -4667
rect 3793 -4787 3893 -4667
rect 3997 -4787 4097 -4667
rect 4201 -4787 4301 -4667
rect 4405 -4787 4505 -4667
rect 4609 -4787 4709 -4667
rect 4813 -4787 4913 -4667
rect 5017 -4787 5117 -4667
rect 5221 -4787 5321 -4667
rect 5425 -4787 5525 -4667
rect 5757 -4787 5857 -4667
rect 5961 -4787 6061 -4667
rect 3589 -5114 3689 -4994
rect 3793 -5114 3893 -4994
rect 3997 -5114 4097 -4994
rect 4201 -5114 4301 -4994
rect 4405 -5114 4505 -4994
rect 4609 -5114 4709 -4994
rect 4813 -5114 4913 -4994
rect 5017 -5114 5117 -4994
rect 5221 -5114 5321 -4994
rect 5425 -5114 5525 -4994
rect 5757 -5114 5857 -4994
rect 5961 -5114 6061 -4994
rect 3589 -5503 3689 -5383
rect 3793 -5503 3893 -5383
rect 3997 -5503 4097 -5383
rect 4201 -5503 4301 -5383
rect 4405 -5503 4505 -5383
rect 4609 -5503 4709 -5383
rect 4813 -5503 4913 -5383
rect 5017 -5503 5117 -5383
rect 5221 -5503 5321 -5383
rect 5425 -5503 5525 -5383
rect 5757 -5503 5857 -5383
rect 5961 -5503 6061 -5383
rect 3589 -5798 3689 -5678
rect 3793 -5798 3893 -5678
rect 3997 -5798 4097 -5678
rect 4201 -5798 4301 -5678
rect 4405 -5798 4505 -5678
rect 4609 -5798 4709 -5678
rect 4813 -5798 4913 -5678
rect 5017 -5798 5117 -5678
rect 5221 -5798 5321 -5678
rect 5425 -5798 5525 -5678
rect 5757 -5798 5857 -5678
rect 5961 -5798 6061 -5678
rect -1970 -6056 -1914 -6006
rect -1492 -6055 -1436 -6011
rect -956 -6055 -900 -6011
rect -352 -6056 -296 -6006
rect 126 -6055 182 -6011
rect 662 -6055 718 -6011
rect 1257 -6056 1313 -6006
rect 1735 -6055 1791 -6011
rect 2271 -6055 2327 -6011
rect 3589 -6183 3689 -6063
rect 3793 -6183 3893 -6063
rect 3997 -6183 4097 -6063
rect 4201 -6183 4301 -6063
rect 4405 -6183 4505 -6063
rect 4609 -6183 4709 -6063
rect 4813 -6183 4913 -6063
rect 5017 -6183 5117 -6063
rect 5221 -6183 5321 -6063
rect 5425 -6183 5525 -6063
rect 5757 -6183 5857 -6063
rect 5961 -6183 6061 -6063
<< pmos >>
rect -1970 -3162 -1914 -3062
rect -1430 -3155 -1374 -3111
rect -1018 -3155 -962 -3111
rect -1970 -4030 -1914 -3930
rect -1430 -4023 -1374 -3979
rect -1018 -4023 -962 -3979
rect -1970 -4889 -1914 -4789
rect -1430 -4882 -1374 -4838
rect -1018 -4882 -962 -4838
rect -1970 -5757 -1914 -5657
rect -1430 -5750 -1374 -5706
rect -1018 -5750 -962 -5706
rect -352 -5757 -296 -5657
rect 188 -5750 244 -5706
rect 600 -5750 656 -5706
rect 1257 -5757 1313 -5657
rect 1797 -5750 1853 -5706
rect 2209 -5750 2265 -5706
<< ndiff >>
rect -1772 1593 -1684 1606
rect -1772 1499 -1759 1593
rect -1713 1499 -1684 1593
rect -1772 1486 -1684 1499
rect -1584 1593 -1496 1606
rect -1584 1499 -1555 1593
rect -1509 1499 -1496 1593
rect -1584 1486 -1496 1499
rect -1385 1593 -1297 1606
rect -1385 1499 -1372 1593
rect -1326 1499 -1297 1593
rect -1385 1486 -1297 1499
rect -1197 1593 -1093 1606
rect -1197 1499 -1168 1593
rect -1122 1499 -1093 1593
rect -1197 1486 -1093 1499
rect -993 1593 -889 1606
rect -993 1499 -964 1593
rect -918 1499 -889 1593
rect -993 1486 -889 1499
rect -789 1593 -685 1606
rect -789 1499 -760 1593
rect -714 1499 -685 1593
rect -789 1486 -685 1499
rect -585 1593 -481 1606
rect -585 1499 -556 1593
rect -510 1499 -481 1593
rect -585 1486 -481 1499
rect -381 1593 -277 1606
rect -381 1499 -352 1593
rect -306 1499 -277 1593
rect -381 1486 -277 1499
rect -177 1593 -73 1606
rect -177 1499 -148 1593
rect -102 1499 -73 1593
rect -177 1486 -73 1499
rect 27 1593 131 1606
rect 27 1499 56 1593
rect 102 1499 131 1593
rect 27 1486 131 1499
rect 231 1593 335 1606
rect 231 1499 260 1593
rect 306 1499 335 1593
rect 231 1486 335 1499
rect 435 1593 539 1606
rect 435 1499 464 1593
rect 510 1499 539 1593
rect 435 1486 539 1499
rect 639 1593 743 1606
rect 639 1499 668 1593
rect 714 1499 743 1593
rect 639 1486 743 1499
rect 843 1593 947 1606
rect 843 1499 872 1593
rect 918 1499 947 1593
rect 843 1486 947 1499
rect 1047 1593 1151 1606
rect 1047 1499 1076 1593
rect 1122 1499 1151 1593
rect 1047 1486 1151 1499
rect 1251 1593 1355 1606
rect 1251 1499 1280 1593
rect 1326 1499 1355 1593
rect 1251 1486 1355 1499
rect 1455 1593 1559 1606
rect 1455 1499 1484 1593
rect 1530 1499 1559 1593
rect 1455 1486 1559 1499
rect 1659 1593 1763 1606
rect 1659 1499 1688 1593
rect 1734 1499 1763 1593
rect 1659 1486 1763 1499
rect 1863 1593 1951 1606
rect 1863 1499 1892 1593
rect 1938 1499 1951 1593
rect 1863 1486 1951 1499
rect 2056 1593 2144 1606
rect 2056 1499 2069 1593
rect 2115 1499 2144 1593
rect 2056 1486 2144 1499
rect 2244 1593 2332 1606
rect 2244 1499 2273 1593
rect 2319 1499 2332 1593
rect 2244 1486 2332 1499
rect 3028 1564 3100 1570
rect 3240 1564 3312 1570
rect 3028 1557 3120 1564
rect 3028 1511 3041 1557
rect 3087 1511 3120 1557
rect 3028 1504 3120 1511
rect 3220 1557 3312 1564
rect 3220 1511 3253 1557
rect 3299 1511 3312 1557
rect 3220 1504 3312 1511
rect 3028 1498 3100 1504
rect 3240 1498 3312 1504
rect 3368 1564 3440 1570
rect 3580 1564 3652 1570
rect 3368 1557 3460 1564
rect 3368 1511 3381 1557
rect 3427 1511 3460 1557
rect 3368 1504 3460 1511
rect 3560 1557 3652 1564
rect 3560 1511 3593 1557
rect 3639 1511 3652 1557
rect 3560 1504 3652 1511
rect 3368 1498 3440 1504
rect 3580 1498 3652 1504
rect 3708 1564 3780 1570
rect 3920 1564 3992 1570
rect 4132 1564 4204 1570
rect 4344 1564 4416 1570
rect 3708 1557 3800 1564
rect 3708 1511 3721 1557
rect 3767 1511 3800 1557
rect 3708 1504 3800 1511
rect 3900 1557 4012 1564
rect 3900 1511 3933 1557
rect 3979 1511 4012 1557
rect 3900 1504 4012 1511
rect 4112 1557 4224 1564
rect 4112 1511 4145 1557
rect 4191 1511 4224 1557
rect 4112 1504 4224 1511
rect 4324 1557 4416 1564
rect 4324 1511 4357 1557
rect 4403 1511 4416 1557
rect 4324 1504 4416 1511
rect 3708 1498 3780 1504
rect -1772 1290 -1684 1303
rect -1772 1196 -1759 1290
rect -1713 1196 -1684 1290
rect -1772 1183 -1684 1196
rect -1584 1290 -1496 1303
rect -1584 1196 -1555 1290
rect -1509 1196 -1496 1290
rect -1584 1183 -1496 1196
rect -1385 1290 -1297 1303
rect -1385 1196 -1372 1290
rect -1326 1196 -1297 1290
rect -1385 1183 -1297 1196
rect -1197 1290 -1093 1303
rect -1197 1196 -1168 1290
rect -1122 1196 -1093 1290
rect -1197 1183 -1093 1196
rect -993 1290 -889 1303
rect -993 1196 -964 1290
rect -918 1196 -889 1290
rect -993 1183 -889 1196
rect -789 1290 -685 1303
rect -789 1196 -760 1290
rect -714 1196 -685 1290
rect -789 1183 -685 1196
rect -585 1290 -481 1303
rect -585 1196 -556 1290
rect -510 1196 -481 1290
rect -585 1183 -481 1196
rect -381 1290 -277 1303
rect -381 1196 -352 1290
rect -306 1196 -277 1290
rect -381 1183 -277 1196
rect -177 1290 -73 1303
rect -177 1196 -148 1290
rect -102 1196 -73 1290
rect -177 1183 -73 1196
rect 27 1290 131 1303
rect 27 1196 56 1290
rect 102 1196 131 1290
rect 27 1183 131 1196
rect 231 1290 335 1303
rect 231 1196 260 1290
rect 306 1196 335 1290
rect 231 1183 335 1196
rect 435 1290 539 1303
rect 435 1196 464 1290
rect 510 1196 539 1290
rect 435 1183 539 1196
rect 639 1290 743 1303
rect 639 1196 668 1290
rect 714 1196 743 1290
rect 639 1183 743 1196
rect 843 1290 947 1303
rect 843 1196 872 1290
rect 918 1196 947 1290
rect 843 1183 947 1196
rect 1047 1290 1151 1303
rect 1047 1196 1076 1290
rect 1122 1196 1151 1290
rect 1047 1183 1151 1196
rect 1251 1290 1355 1303
rect 1251 1196 1280 1290
rect 1326 1196 1355 1290
rect 1251 1183 1355 1196
rect 1455 1290 1559 1303
rect 1455 1196 1484 1290
rect 1530 1196 1559 1290
rect 1455 1183 1559 1196
rect 1659 1290 1763 1303
rect 1659 1196 1688 1290
rect 1734 1196 1763 1290
rect 1659 1183 1763 1196
rect 1863 1290 1951 1303
rect 1863 1196 1892 1290
rect 1938 1196 1951 1290
rect 1863 1183 1951 1196
rect 2056 1290 2144 1303
rect 2056 1196 2069 1290
rect 2115 1196 2144 1290
rect 2056 1183 2144 1196
rect 2244 1290 2332 1303
rect 2244 1196 2273 1290
rect 2319 1196 2332 1290
rect 2244 1183 2332 1196
rect 3920 1498 3992 1504
rect 4132 1498 4204 1504
rect 4344 1498 4416 1504
rect 4703 1498 4775 1504
rect 4915 1498 4987 1504
rect 5127 1498 5199 1504
rect 4703 1491 4795 1498
rect 4703 1445 4716 1491
rect 4762 1445 4795 1491
rect 4703 1438 4795 1445
rect 4895 1491 5007 1498
rect 4895 1445 4928 1491
rect 4974 1445 5007 1491
rect 4895 1438 5007 1445
rect 5107 1491 5199 1498
rect 5107 1445 5140 1491
rect 5186 1445 5199 1491
rect 5107 1438 5199 1445
rect 4703 1432 4775 1438
rect 4915 1432 4987 1438
rect 3036 1291 3124 1304
rect 3036 1197 3049 1291
rect 3095 1197 3124 1291
rect 3036 1184 3124 1197
rect 3224 1291 3312 1304
rect 3224 1197 3253 1291
rect 3299 1197 3312 1291
rect 3224 1184 3312 1197
rect 3368 1291 3456 1304
rect 3368 1197 3381 1291
rect 3427 1197 3456 1291
rect 3368 1184 3456 1197
rect 3556 1291 3660 1304
rect 3556 1197 3585 1291
rect 3631 1197 3660 1291
rect 3556 1184 3660 1197
rect 3760 1291 3864 1304
rect 3760 1197 3789 1291
rect 3835 1197 3864 1291
rect 3760 1184 3864 1197
rect 3964 1291 4068 1304
rect 3964 1197 3993 1291
rect 4039 1197 4068 1291
rect 3964 1184 4068 1197
rect 4168 1291 4272 1304
rect 4168 1197 4197 1291
rect 4243 1197 4272 1291
rect 4168 1184 4272 1197
rect 4372 1291 4460 1304
rect 4372 1197 4401 1291
rect 4447 1197 4460 1291
rect 4372 1184 4460 1197
rect 4703 1256 4775 1262
rect 4915 1256 4987 1262
rect 5127 1432 5199 1438
rect 5255 1498 5327 1504
rect 5467 1498 5539 1504
rect 5679 1498 5751 1504
rect 5255 1491 5347 1498
rect 5255 1445 5268 1491
rect 5314 1445 5347 1491
rect 5255 1438 5347 1445
rect 5447 1491 5559 1498
rect 5447 1445 5480 1491
rect 5526 1445 5559 1491
rect 5447 1438 5559 1445
rect 5659 1491 5751 1498
rect 5659 1445 5692 1491
rect 5738 1445 5751 1491
rect 5659 1438 5751 1445
rect 5255 1432 5327 1438
rect 5127 1256 5199 1262
rect 4703 1249 4795 1256
rect 4703 1203 4716 1249
rect 4762 1203 4795 1249
rect 4703 1196 4795 1203
rect 4895 1249 5007 1256
rect 4895 1203 4928 1249
rect 4974 1203 5007 1249
rect 4895 1196 5007 1203
rect 5107 1249 5199 1256
rect 5107 1203 5140 1249
rect 5186 1203 5199 1249
rect 5107 1196 5199 1203
rect 4703 1190 4775 1196
rect 4915 1190 4987 1196
rect 5127 1190 5199 1196
rect 5255 1256 5327 1262
rect 5467 1432 5539 1438
rect 5467 1256 5539 1262
rect 5679 1432 5751 1438
rect 5807 1498 5879 1504
rect 6019 1498 6091 1504
rect 5807 1491 5899 1498
rect 5807 1445 5820 1491
rect 5866 1445 5899 1491
rect 5807 1438 5899 1445
rect 5999 1491 6091 1498
rect 5999 1445 6032 1491
rect 6078 1445 6091 1491
rect 5999 1438 6091 1445
rect 5807 1432 5879 1438
rect 5679 1256 5751 1262
rect 5255 1249 5347 1256
rect 5255 1203 5268 1249
rect 5314 1203 5347 1249
rect 5255 1196 5347 1203
rect 5447 1249 5559 1256
rect 5447 1203 5480 1249
rect 5526 1203 5559 1249
rect 5447 1196 5559 1203
rect 5659 1249 5751 1256
rect 5659 1203 5692 1249
rect 5738 1203 5751 1249
rect 5659 1196 5751 1203
rect 5255 1190 5327 1196
rect 5467 1190 5539 1196
rect 3028 936 3100 942
rect 3240 936 3312 942
rect 3028 929 3120 936
rect 3028 883 3041 929
rect 3087 883 3120 929
rect 3028 876 3120 883
rect 3220 929 3312 936
rect 3220 883 3253 929
rect 3299 883 3312 929
rect 3220 876 3312 883
rect 3028 870 3100 876
rect -1772 851 -1684 864
rect -1772 757 -1759 851
rect -1713 757 -1684 851
rect -1772 744 -1684 757
rect -1584 851 -1496 864
rect -1584 757 -1555 851
rect -1509 757 -1496 851
rect -1584 744 -1496 757
rect -1385 851 -1297 864
rect -1385 757 -1372 851
rect -1326 757 -1297 851
rect -1385 744 -1297 757
rect -1197 851 -1093 864
rect -1197 757 -1168 851
rect -1122 757 -1093 851
rect -1197 744 -1093 757
rect -993 851 -889 864
rect -993 757 -964 851
rect -918 757 -889 851
rect -993 744 -889 757
rect -789 851 -685 864
rect -789 757 -760 851
rect -714 757 -685 851
rect -789 744 -685 757
rect -585 851 -481 864
rect -585 757 -556 851
rect -510 757 -481 851
rect -585 744 -481 757
rect -381 851 -277 864
rect -381 757 -352 851
rect -306 757 -277 851
rect -381 744 -277 757
rect -177 851 -73 864
rect -177 757 -148 851
rect -102 757 -73 851
rect -177 744 -73 757
rect 27 851 131 864
rect 27 757 56 851
rect 102 757 131 851
rect 27 744 131 757
rect 231 851 335 864
rect 231 757 260 851
rect 306 757 335 851
rect 231 744 335 757
rect 435 851 539 864
rect 435 757 464 851
rect 510 757 539 851
rect 435 744 539 757
rect 639 851 743 864
rect 639 757 668 851
rect 714 757 743 851
rect 639 744 743 757
rect 843 851 947 864
rect 843 757 872 851
rect 918 757 947 851
rect 843 744 947 757
rect 1047 851 1151 864
rect 1047 757 1076 851
rect 1122 757 1151 851
rect 1047 744 1151 757
rect 1251 851 1355 864
rect 1251 757 1280 851
rect 1326 757 1355 851
rect 1251 744 1355 757
rect 1455 851 1559 864
rect 1455 757 1484 851
rect 1530 757 1559 851
rect 1455 744 1559 757
rect 1659 851 1763 864
rect 1659 757 1688 851
rect 1734 757 1763 851
rect 1659 744 1763 757
rect 1863 851 1951 864
rect 1863 757 1892 851
rect 1938 757 1951 851
rect 1863 744 1951 757
rect 2056 851 2144 864
rect 2056 757 2069 851
rect 2115 757 2144 851
rect 2056 744 2144 757
rect 2244 851 2332 864
rect 2244 757 2273 851
rect 2319 757 2332 851
rect 2244 744 2332 757
rect 3240 870 3312 876
rect 3368 936 3440 942
rect 3580 936 3652 942
rect 3368 929 3460 936
rect 3368 883 3381 929
rect 3427 883 3460 929
rect 3368 876 3460 883
rect 3560 929 3652 936
rect 3560 883 3593 929
rect 3639 883 3652 929
rect 3560 876 3652 883
rect 3368 870 3440 876
rect 3580 870 3652 876
rect 3708 936 3780 942
rect 3920 936 3992 942
rect 4132 936 4204 942
rect 3708 929 3800 936
rect 3708 883 3721 929
rect 3767 883 3800 929
rect 3708 876 3800 883
rect 3900 929 4012 936
rect 3900 883 3933 929
rect 3979 883 4012 929
rect 3900 876 4012 883
rect 4112 929 4204 936
rect 4112 883 4145 929
rect 4191 883 4204 929
rect 4112 876 4204 883
rect 3708 870 3780 876
rect 3920 870 3992 876
rect 4132 870 4204 876
rect 4260 936 4332 942
rect 5679 1190 5751 1196
rect 5807 1256 5879 1262
rect 6019 1432 6091 1438
rect 6019 1256 6091 1262
rect 5807 1249 5899 1256
rect 5807 1203 5820 1249
rect 5866 1203 5899 1249
rect 5807 1196 5899 1203
rect 5999 1249 6091 1256
rect 5999 1203 6032 1249
rect 6078 1203 6091 1249
rect 5999 1196 6091 1203
rect 5807 1190 5879 1196
rect 6019 1190 6091 1196
rect 4849 965 4937 978
rect 4472 936 4544 942
rect 4260 929 4352 936
rect 4260 883 4273 929
rect 4319 883 4352 929
rect 4260 876 4352 883
rect 4452 929 4544 936
rect 4452 883 4485 929
rect 4531 883 4544 929
rect 4452 876 4544 883
rect 4260 870 4332 876
rect 4472 870 4544 876
rect 4849 871 4862 965
rect 4908 871 4937 965
rect 4849 858 4937 871
rect 5037 965 5141 978
rect 5037 871 5066 965
rect 5112 871 5141 965
rect 5037 858 5141 871
rect 5241 965 5345 978
rect 5241 871 5270 965
rect 5316 871 5345 965
rect 5241 858 5345 871
rect 5445 965 5549 978
rect 5445 871 5474 965
rect 5520 871 5549 965
rect 5445 858 5549 871
rect 5649 965 5753 978
rect 5649 871 5678 965
rect 5724 871 5753 965
rect 5649 858 5753 871
rect 5853 965 5941 978
rect 5853 871 5882 965
rect 5928 871 5941 965
rect 5853 858 5941 871
rect 3110 645 3198 658
rect 3110 551 3123 645
rect 3169 551 3198 645
rect 3110 538 3198 551
rect 3298 645 3402 658
rect 3298 551 3327 645
rect 3373 551 3402 645
rect 3298 538 3402 551
rect 3502 645 3606 658
rect 3502 551 3531 645
rect 3577 551 3606 645
rect 3502 538 3606 551
rect 3706 645 3810 658
rect 3706 551 3735 645
rect 3781 551 3810 645
rect 3706 538 3810 551
rect 3910 645 4014 658
rect 3910 551 3939 645
rect 3985 551 4014 645
rect 3910 538 4014 551
rect 4114 645 4218 658
rect 4114 551 4143 645
rect 4189 551 4218 645
rect 4114 538 4218 551
rect 4318 645 4422 658
rect 4318 551 4347 645
rect 4393 551 4422 645
rect 4318 538 4422 551
rect 4522 645 4610 658
rect 4522 551 4551 645
rect 4597 551 4610 645
rect 4849 663 4937 676
rect 4849 569 4862 663
rect 4908 569 4937 663
rect 4849 556 4937 569
rect 5037 663 5141 676
rect 5037 569 5066 663
rect 5112 569 5141 663
rect 5037 556 5141 569
rect 5241 663 5345 676
rect 5241 569 5270 663
rect 5316 569 5345 663
rect 5241 556 5345 569
rect 5445 663 5549 676
rect 5445 569 5474 663
rect 5520 569 5549 663
rect 5445 556 5549 569
rect 5649 663 5753 676
rect 5649 569 5678 663
rect 5724 569 5753 663
rect 5649 556 5753 569
rect 5853 663 5941 676
rect 5853 569 5882 663
rect 5928 569 5941 663
rect 5853 556 5941 569
rect 4522 538 4610 551
rect -1772 175 -1684 188
rect -1772 81 -1759 175
rect -1713 81 -1684 175
rect -1772 68 -1684 81
rect -1584 175 -1480 188
rect -1584 81 -1555 175
rect -1509 81 -1480 175
rect -1584 68 -1480 81
rect -1380 175 -1276 188
rect -1380 81 -1351 175
rect -1305 81 -1276 175
rect -1380 68 -1276 81
rect -1176 175 -1072 188
rect -1176 81 -1147 175
rect -1101 81 -1072 175
rect -1176 68 -1072 81
rect -972 175 -884 188
rect -972 81 -943 175
rect -897 81 -884 175
rect -972 68 -884 81
rect -828 175 -740 188
rect -828 81 -815 175
rect -769 81 -740 175
rect -828 68 -740 81
rect -640 175 -536 188
rect -640 81 -611 175
rect -565 81 -536 175
rect -640 68 -536 81
rect -436 175 -348 188
rect -436 81 -407 175
rect -361 81 -348 175
rect -436 68 -348 81
rect -292 175 -204 188
rect -292 81 -279 175
rect -233 81 -204 175
rect -292 68 -204 81
rect -104 175 -16 188
rect -104 81 -75 175
rect -29 81 -16 175
rect -104 68 -16 81
rect 40 175 128 188
rect 40 81 53 175
rect 99 81 128 175
rect 40 68 128 81
rect 228 175 332 188
rect 228 81 257 175
rect 303 81 332 175
rect 228 68 332 81
rect 432 175 520 188
rect 432 81 461 175
rect 507 81 520 175
rect 432 68 520 81
rect 576 175 664 188
rect 576 81 589 175
rect 635 81 664 175
rect 576 68 664 81
rect 764 175 852 188
rect 764 81 793 175
rect 839 81 852 175
rect 764 68 852 81
rect 908 175 996 188
rect 908 81 921 175
rect 967 81 996 175
rect 908 68 996 81
rect 1096 175 1200 188
rect 1096 81 1125 175
rect 1171 81 1200 175
rect 1096 68 1200 81
rect 1300 175 1388 188
rect 1300 81 1329 175
rect 1375 81 1388 175
rect 1300 68 1388 81
rect 1444 175 1532 188
rect 1444 81 1457 175
rect 1503 81 1532 175
rect 1444 68 1532 81
rect 1632 175 1736 188
rect 1632 81 1661 175
rect 1707 81 1736 175
rect 1632 68 1736 81
rect 1836 175 1940 188
rect 1836 81 1865 175
rect 1911 81 1940 175
rect 1836 68 1940 81
rect 2040 175 2144 188
rect 2040 81 2069 175
rect 2115 81 2144 175
rect 2040 68 2144 81
rect 2244 175 2332 188
rect 2244 81 2273 175
rect 2319 81 2332 175
rect 2244 68 2332 81
rect 2950 121 3038 134
rect 2950 27 2963 121
rect 3009 27 3038 121
rect 2950 14 3038 27
rect 3138 121 3242 134
rect 3138 27 3167 121
rect 3213 27 3242 121
rect 3138 14 3242 27
rect 3342 121 3446 134
rect 3342 27 3371 121
rect 3417 27 3446 121
rect 3342 14 3446 27
rect 3546 121 3650 134
rect 3546 27 3575 121
rect 3621 27 3650 121
rect 3546 14 3650 27
rect 3750 121 3854 134
rect 3750 27 3779 121
rect 3825 27 3854 121
rect 3750 14 3854 27
rect 3954 121 4058 134
rect 3954 27 3983 121
rect 4029 27 4058 121
rect 3954 14 4058 27
rect 4158 121 4246 134
rect 4158 27 4187 121
rect 4233 27 4246 121
rect 4417 98 4489 104
rect 4629 98 4701 104
rect 4417 91 4509 98
rect 4417 45 4430 91
rect 4476 45 4509 91
rect 4417 38 4509 45
rect 4609 91 4701 98
rect 4609 45 4642 91
rect 4688 45 4701 91
rect 4609 38 4701 45
rect 4417 32 4489 38
rect 4158 14 4246 27
rect -1772 -151 -1684 -138
rect -1772 -245 -1759 -151
rect -1713 -245 -1684 -151
rect -1772 -258 -1684 -245
rect -1584 -151 -1480 -138
rect -1584 -245 -1555 -151
rect -1509 -245 -1480 -151
rect -1584 -258 -1480 -245
rect -1380 -151 -1276 -138
rect -1380 -245 -1351 -151
rect -1305 -245 -1276 -151
rect -1380 -258 -1276 -245
rect -1176 -151 -1072 -138
rect -1176 -245 -1147 -151
rect -1101 -245 -1072 -151
rect -1176 -258 -1072 -245
rect -972 -151 -884 -138
rect -972 -245 -943 -151
rect -897 -245 -884 -151
rect -972 -258 -884 -245
rect -828 -151 -740 -138
rect -828 -245 -815 -151
rect -769 -245 -740 -151
rect -828 -258 -740 -245
rect -640 -151 -536 -138
rect -640 -245 -611 -151
rect -565 -245 -536 -151
rect -640 -258 -536 -245
rect -436 -151 -348 -138
rect -436 -245 -407 -151
rect -361 -245 -348 -151
rect -436 -258 -348 -245
rect -292 -151 -204 -138
rect -292 -245 -279 -151
rect -233 -245 -204 -151
rect -292 -258 -204 -245
rect -104 -151 -16 -138
rect -104 -245 -75 -151
rect -29 -245 -16 -151
rect -104 -258 -16 -245
rect 40 -151 128 -138
rect 40 -245 53 -151
rect 99 -245 128 -151
rect 40 -258 128 -245
rect 228 -151 332 -138
rect 228 -245 257 -151
rect 303 -245 332 -151
rect 228 -258 332 -245
rect 432 -151 520 -138
rect 432 -245 461 -151
rect 507 -245 520 -151
rect 432 -258 520 -245
rect 576 -151 664 -138
rect 576 -245 589 -151
rect 635 -245 664 -151
rect 576 -258 664 -245
rect 764 -151 852 -138
rect 764 -245 793 -151
rect 839 -245 852 -151
rect 764 -258 852 -245
rect 908 -151 996 -138
rect 908 -245 921 -151
rect 967 -245 996 -151
rect 908 -258 996 -245
rect 1096 -151 1200 -138
rect 1096 -245 1125 -151
rect 1171 -245 1200 -151
rect 1096 -258 1200 -245
rect 1300 -151 1388 -138
rect 1300 -245 1329 -151
rect 1375 -245 1388 -151
rect 1300 -258 1388 -245
rect 1444 -151 1532 -138
rect 1444 -245 1457 -151
rect 1503 -245 1532 -151
rect 1444 -258 1532 -245
rect 1632 -151 1736 -138
rect 1632 -245 1661 -151
rect 1707 -245 1736 -151
rect 1632 -258 1736 -245
rect 1836 -151 1940 -138
rect 1836 -245 1865 -151
rect 1911 -245 1940 -151
rect 1836 -258 1940 -245
rect 2040 -151 2144 -138
rect 2040 -245 2069 -151
rect 2115 -245 2144 -151
rect 2040 -258 2144 -245
rect 2244 -151 2332 -138
rect 2244 -245 2273 -151
rect 2319 -245 2332 -151
rect 2244 -258 2332 -245
rect 4629 32 4701 38
rect 4757 98 4829 104
rect 4969 98 5041 104
rect 5181 98 5253 104
rect 4757 91 4849 98
rect 4757 45 4770 91
rect 4816 45 4849 91
rect 4757 38 4849 45
rect 4949 91 5061 98
rect 4949 45 4982 91
rect 5028 45 5061 91
rect 4949 38 5061 45
rect 5161 91 5253 98
rect 5161 45 5194 91
rect 5240 45 5253 91
rect 5161 38 5253 45
rect 4757 32 4829 38
rect 4969 32 5041 38
rect 5181 32 5253 38
rect 5309 98 5381 104
rect 5521 98 5593 104
rect 5733 98 5805 104
rect 5309 91 5401 98
rect 5309 45 5322 91
rect 5368 45 5401 91
rect 5309 38 5401 45
rect 5501 91 5613 98
rect 5501 45 5534 91
rect 5580 45 5613 91
rect 5501 38 5613 45
rect 5713 91 5805 98
rect 5713 45 5746 91
rect 5792 45 5805 91
rect 5713 38 5805 45
rect 5309 32 5381 38
rect 5521 32 5593 38
rect 5733 32 5805 38
rect 4416 -218 4488 -212
rect 4628 -218 4700 -212
rect 4416 -225 4508 -218
rect 2950 -257 3038 -244
rect 2950 -351 2963 -257
rect 3009 -351 3038 -257
rect 2950 -364 3038 -351
rect 3138 -257 3242 -244
rect 3138 -351 3167 -257
rect 3213 -351 3242 -257
rect 3138 -364 3242 -351
rect 3342 -257 3446 -244
rect 3342 -351 3371 -257
rect 3417 -351 3446 -257
rect 3342 -364 3446 -351
rect 3546 -257 3650 -244
rect 3546 -351 3575 -257
rect 3621 -351 3650 -257
rect 3546 -364 3650 -351
rect 3750 -257 3854 -244
rect 3750 -351 3779 -257
rect 3825 -351 3854 -257
rect 3750 -364 3854 -351
rect 3954 -257 4058 -244
rect 3954 -351 3983 -257
rect 4029 -351 4058 -257
rect 3954 -364 4058 -351
rect 4158 -257 4246 -244
rect 4158 -351 4187 -257
rect 4233 -351 4246 -257
rect 4416 -271 4429 -225
rect 4475 -271 4508 -225
rect 4416 -278 4508 -271
rect 4608 -225 4700 -218
rect 4608 -271 4641 -225
rect 4687 -271 4700 -225
rect 4608 -278 4700 -271
rect 4416 -284 4488 -278
rect 4158 -364 4246 -351
rect 4416 -468 4488 -462
rect 4628 -284 4700 -278
rect 4756 -218 4828 -212
rect 4968 -218 5040 -212
rect 5180 -218 5252 -212
rect 4756 -225 4848 -218
rect 4756 -271 4769 -225
rect 4815 -271 4848 -225
rect 4756 -278 4848 -271
rect 4948 -225 5060 -218
rect 4948 -271 4981 -225
rect 5027 -271 5060 -225
rect 4948 -278 5060 -271
rect 5160 -225 5252 -218
rect 5160 -271 5193 -225
rect 5239 -271 5252 -225
rect 5160 -278 5252 -271
rect 4756 -284 4828 -278
rect 4968 -284 5040 -278
rect 5180 -284 5252 -278
rect 5308 -218 5380 -212
rect 5520 -218 5592 -212
rect 5732 -218 5804 -212
rect 5308 -225 5400 -218
rect 5308 -271 5321 -225
rect 5367 -271 5400 -225
rect 5308 -278 5400 -271
rect 5500 -225 5612 -218
rect 5500 -271 5533 -225
rect 5579 -271 5612 -225
rect 5500 -278 5612 -271
rect 5712 -225 5804 -218
rect 5712 -271 5745 -225
rect 5791 -271 5804 -225
rect 5712 -278 5804 -271
rect 5308 -284 5380 -278
rect 4628 -468 4700 -462
rect 4416 -475 4508 -468
rect 4416 -521 4429 -475
rect 4475 -521 4508 -475
rect 2950 -536 3038 -523
rect 2950 -630 2963 -536
rect 3009 -630 3038 -536
rect 2950 -643 3038 -630
rect 3138 -536 3242 -523
rect 3138 -630 3167 -536
rect 3213 -630 3242 -536
rect 3138 -643 3242 -630
rect 3342 -536 3446 -523
rect 3342 -630 3371 -536
rect 3417 -630 3446 -536
rect 3342 -643 3446 -630
rect 3546 -536 3650 -523
rect 3546 -630 3575 -536
rect 3621 -630 3650 -536
rect 3546 -643 3650 -630
rect 3750 -536 3854 -523
rect 3750 -630 3779 -536
rect 3825 -630 3854 -536
rect 3750 -643 3854 -630
rect 3954 -536 4058 -523
rect 3954 -630 3983 -536
rect 4029 -630 4058 -536
rect 3954 -643 4058 -630
rect 4158 -536 4246 -523
rect 4416 -528 4508 -521
rect 4608 -475 4700 -468
rect 4608 -521 4641 -475
rect 4687 -521 4700 -475
rect 4608 -528 4700 -521
rect 4416 -534 4488 -528
rect 4158 -630 4187 -536
rect 4233 -630 4246 -536
rect 4628 -534 4700 -528
rect 4756 -468 4828 -462
rect 4968 -468 5040 -462
rect 5180 -468 5252 -462
rect 4756 -475 4848 -468
rect 4756 -521 4769 -475
rect 4815 -521 4848 -475
rect 4756 -528 4848 -521
rect 4948 -475 5060 -468
rect 4948 -521 4981 -475
rect 5027 -521 5060 -475
rect 4948 -528 5060 -521
rect 5160 -475 5252 -468
rect 5160 -521 5193 -475
rect 5239 -521 5252 -475
rect 5160 -528 5252 -521
rect 4756 -534 4828 -528
rect 4968 -534 5040 -528
rect 5180 -534 5252 -528
rect 5308 -468 5380 -462
rect 5520 -284 5592 -278
rect 5732 -284 5804 -278
rect 5520 -468 5592 -462
rect 5732 -468 5804 -462
rect 5308 -475 5400 -468
rect 5308 -521 5321 -475
rect 5367 -521 5400 -475
rect 5308 -528 5400 -521
rect 5500 -475 5612 -468
rect 5500 -521 5533 -475
rect 5579 -521 5612 -475
rect 5500 -528 5612 -521
rect 5712 -475 5804 -468
rect 5712 -521 5745 -475
rect 5791 -521 5804 -475
rect 5712 -528 5804 -521
rect 5308 -534 5380 -528
rect 5520 -534 5592 -528
rect 5732 -534 5804 -528
rect 4158 -643 4246 -630
rect 4416 -793 4488 -787
rect 4628 -793 4700 -787
rect 4416 -800 4508 -793
rect -1772 -943 -1684 -930
rect -1772 -1037 -1759 -943
rect -1713 -1037 -1684 -943
rect -1772 -1050 -1684 -1037
rect -1584 -943 -1496 -930
rect -1584 -1037 -1555 -943
rect -1509 -1037 -1496 -943
rect -1584 -1050 -1496 -1037
rect -1385 -943 -1297 -930
rect -1385 -1037 -1372 -943
rect -1326 -1037 -1297 -943
rect -1385 -1050 -1297 -1037
rect -1197 -943 -1093 -930
rect -1197 -1037 -1168 -943
rect -1122 -1037 -1093 -943
rect -1197 -1050 -1093 -1037
rect -993 -943 -889 -930
rect -993 -1037 -964 -943
rect -918 -1037 -889 -943
rect -993 -1050 -889 -1037
rect -789 -943 -685 -930
rect -789 -1037 -760 -943
rect -714 -1037 -685 -943
rect -789 -1050 -685 -1037
rect -585 -943 -481 -930
rect -585 -1037 -556 -943
rect -510 -1037 -481 -943
rect -585 -1050 -481 -1037
rect -381 -943 -277 -930
rect -381 -1037 -352 -943
rect -306 -1037 -277 -943
rect -381 -1050 -277 -1037
rect -177 -943 -73 -930
rect -177 -1037 -148 -943
rect -102 -1037 -73 -943
rect -177 -1050 -73 -1037
rect 27 -943 131 -930
rect 27 -1037 56 -943
rect 102 -1037 131 -943
rect 27 -1050 131 -1037
rect 231 -943 335 -930
rect 231 -1037 260 -943
rect 306 -1037 335 -943
rect 231 -1050 335 -1037
rect 435 -943 539 -930
rect 435 -1037 464 -943
rect 510 -1037 539 -943
rect 435 -1050 539 -1037
rect 639 -943 743 -930
rect 639 -1037 668 -943
rect 714 -1037 743 -943
rect 639 -1050 743 -1037
rect 843 -943 947 -930
rect 843 -1037 872 -943
rect 918 -1037 947 -943
rect 843 -1050 947 -1037
rect 1047 -943 1151 -930
rect 1047 -1037 1076 -943
rect 1122 -1037 1151 -943
rect 1047 -1050 1151 -1037
rect 1251 -943 1355 -930
rect 1251 -1037 1280 -943
rect 1326 -1037 1355 -943
rect 1251 -1050 1355 -1037
rect 1455 -943 1559 -930
rect 1455 -1037 1484 -943
rect 1530 -1037 1559 -943
rect 1455 -1050 1559 -1037
rect 1659 -943 1763 -930
rect 1659 -1037 1688 -943
rect 1734 -1037 1763 -943
rect 1659 -1050 1763 -1037
rect 1863 -943 1951 -930
rect 1863 -1037 1892 -943
rect 1938 -1037 1951 -943
rect 1863 -1050 1951 -1037
rect 2056 -943 2144 -930
rect 2056 -1037 2069 -943
rect 2115 -1037 2144 -943
rect 2056 -1050 2144 -1037
rect 2244 -943 2332 -930
rect 2244 -1037 2273 -943
rect 2319 -1037 2332 -943
rect 2244 -1050 2332 -1037
rect 4416 -846 4429 -800
rect 4475 -846 4508 -800
rect 4416 -853 4508 -846
rect 4608 -800 4700 -793
rect 4608 -846 4641 -800
rect 4687 -846 4700 -800
rect 4608 -853 4700 -846
rect 4416 -859 4488 -853
rect 2950 -914 3038 -901
rect 2950 -1008 2963 -914
rect 3009 -1008 3038 -914
rect 2950 -1021 3038 -1008
rect 3138 -914 3242 -901
rect 3138 -1008 3167 -914
rect 3213 -1008 3242 -914
rect 3138 -1021 3242 -1008
rect 3342 -914 3446 -901
rect 3342 -1008 3371 -914
rect 3417 -1008 3446 -914
rect 3342 -1021 3446 -1008
rect 3546 -914 3650 -901
rect 3546 -1008 3575 -914
rect 3621 -1008 3650 -914
rect 3546 -1021 3650 -1008
rect 3750 -914 3854 -901
rect 3750 -1008 3779 -914
rect 3825 -1008 3854 -914
rect 3750 -1021 3854 -1008
rect 3954 -914 4058 -901
rect 3954 -1008 3983 -914
rect 4029 -1008 4058 -914
rect 3954 -1021 4058 -1008
rect 4158 -914 4246 -901
rect 4158 -1008 4187 -914
rect 4233 -1008 4246 -914
rect 4158 -1021 4246 -1008
rect 4628 -859 4700 -853
rect 4756 -793 4828 -787
rect 4968 -793 5040 -787
rect 5180 -793 5252 -787
rect 4756 -800 4848 -793
rect 4756 -846 4769 -800
rect 4815 -846 4848 -800
rect 4756 -853 4848 -846
rect 4948 -800 5060 -793
rect 4948 -846 4981 -800
rect 5027 -846 5060 -800
rect 4948 -853 5060 -846
rect 5160 -800 5252 -793
rect 5160 -846 5193 -800
rect 5239 -846 5252 -800
rect 5160 -853 5252 -846
rect 4756 -859 4828 -853
rect 4968 -859 5040 -853
rect 5180 -859 5252 -853
rect 5308 -793 5380 -787
rect 5520 -793 5592 -787
rect 5732 -793 5804 -787
rect 5308 -800 5400 -793
rect 5308 -846 5321 -800
rect 5367 -846 5400 -800
rect 5308 -853 5400 -846
rect 5500 -800 5612 -793
rect 5500 -846 5533 -800
rect 5579 -846 5612 -800
rect 5500 -853 5612 -846
rect 5712 -800 5804 -793
rect 5712 -846 5745 -800
rect 5791 -846 5804 -800
rect 5712 -853 5804 -846
rect 5308 -859 5380 -853
rect 5520 -859 5592 -853
rect 5732 -859 5804 -853
rect -1772 -1374 -1684 -1361
rect -1772 -1468 -1759 -1374
rect -1713 -1468 -1684 -1374
rect -1772 -1481 -1684 -1468
rect -1584 -1374 -1496 -1361
rect -1584 -1468 -1555 -1374
rect -1509 -1468 -1496 -1374
rect -1584 -1481 -1496 -1468
rect -1385 -1374 -1297 -1361
rect -1385 -1468 -1372 -1374
rect -1326 -1468 -1297 -1374
rect -1385 -1481 -1297 -1468
rect -1197 -1374 -1093 -1361
rect -1197 -1468 -1168 -1374
rect -1122 -1468 -1093 -1374
rect -1197 -1481 -1093 -1468
rect -993 -1374 -889 -1361
rect -993 -1468 -964 -1374
rect -918 -1468 -889 -1374
rect -993 -1481 -889 -1468
rect -789 -1374 -685 -1361
rect -789 -1468 -760 -1374
rect -714 -1468 -685 -1374
rect -789 -1481 -685 -1468
rect -585 -1374 -481 -1361
rect -585 -1468 -556 -1374
rect -510 -1468 -481 -1374
rect -585 -1481 -481 -1468
rect -381 -1374 -277 -1361
rect -381 -1468 -352 -1374
rect -306 -1468 -277 -1374
rect -381 -1481 -277 -1468
rect -177 -1374 -73 -1361
rect -177 -1468 -148 -1374
rect -102 -1468 -73 -1374
rect -177 -1481 -73 -1468
rect 27 -1374 131 -1361
rect 27 -1468 56 -1374
rect 102 -1468 131 -1374
rect 27 -1481 131 -1468
rect 231 -1374 335 -1361
rect 231 -1468 260 -1374
rect 306 -1468 335 -1374
rect 231 -1481 335 -1468
rect 435 -1374 539 -1361
rect 435 -1468 464 -1374
rect 510 -1468 539 -1374
rect 435 -1481 539 -1468
rect 639 -1374 743 -1361
rect 639 -1468 668 -1374
rect 714 -1468 743 -1374
rect 639 -1481 743 -1468
rect 843 -1374 947 -1361
rect 843 -1468 872 -1374
rect 918 -1468 947 -1374
rect 843 -1481 947 -1468
rect 1047 -1374 1151 -1361
rect 1047 -1468 1076 -1374
rect 1122 -1468 1151 -1374
rect 1047 -1481 1151 -1468
rect 1251 -1374 1355 -1361
rect 1251 -1468 1280 -1374
rect 1326 -1468 1355 -1374
rect 1251 -1481 1355 -1468
rect 1455 -1374 1559 -1361
rect 1455 -1468 1484 -1374
rect 1530 -1468 1559 -1374
rect 1455 -1481 1559 -1468
rect 1659 -1374 1763 -1361
rect 1659 -1468 1688 -1374
rect 1734 -1468 1763 -1374
rect 1659 -1481 1763 -1468
rect 1863 -1374 1951 -1361
rect 1863 -1468 1892 -1374
rect 1938 -1468 1951 -1374
rect 1863 -1481 1951 -1468
rect 2056 -1374 2144 -1361
rect 2056 -1468 2069 -1374
rect 2115 -1468 2144 -1374
rect 2056 -1481 2144 -1468
rect 2244 -1374 2332 -1361
rect 2244 -1468 2273 -1374
rect 2319 -1468 2332 -1374
rect 2244 -1481 2332 -1468
rect -1772 -1684 -1684 -1671
rect -1772 -1778 -1759 -1684
rect -1713 -1778 -1684 -1684
rect -1772 -1791 -1684 -1778
rect -1584 -1684 -1496 -1671
rect -1584 -1778 -1555 -1684
rect -1509 -1778 -1496 -1684
rect -1584 -1791 -1496 -1778
rect -1385 -1684 -1297 -1671
rect -1385 -1778 -1372 -1684
rect -1326 -1778 -1297 -1684
rect -1385 -1791 -1297 -1778
rect -1197 -1684 -1093 -1671
rect -1197 -1778 -1168 -1684
rect -1122 -1778 -1093 -1684
rect -1197 -1791 -1093 -1778
rect -993 -1684 -889 -1671
rect -993 -1778 -964 -1684
rect -918 -1778 -889 -1684
rect -993 -1791 -889 -1778
rect -789 -1684 -685 -1671
rect -789 -1778 -760 -1684
rect -714 -1778 -685 -1684
rect -789 -1791 -685 -1778
rect -585 -1684 -481 -1671
rect -585 -1778 -556 -1684
rect -510 -1778 -481 -1684
rect -585 -1791 -481 -1778
rect -381 -1684 -277 -1671
rect -381 -1778 -352 -1684
rect -306 -1778 -277 -1684
rect -381 -1791 -277 -1778
rect -177 -1684 -73 -1671
rect -177 -1778 -148 -1684
rect -102 -1778 -73 -1684
rect -177 -1791 -73 -1778
rect 27 -1684 131 -1671
rect 27 -1778 56 -1684
rect 102 -1778 131 -1684
rect 27 -1791 131 -1778
rect 231 -1684 335 -1671
rect 231 -1778 260 -1684
rect 306 -1778 335 -1684
rect 231 -1791 335 -1778
rect 435 -1684 539 -1671
rect 435 -1778 464 -1684
rect 510 -1778 539 -1684
rect 435 -1791 539 -1778
rect 639 -1684 743 -1671
rect 639 -1778 668 -1684
rect 714 -1778 743 -1684
rect 639 -1791 743 -1778
rect 843 -1684 947 -1671
rect 843 -1778 872 -1684
rect 918 -1778 947 -1684
rect 843 -1791 947 -1778
rect 1047 -1684 1151 -1671
rect 1047 -1778 1076 -1684
rect 1122 -1778 1151 -1684
rect 1047 -1791 1151 -1778
rect 1251 -1684 1355 -1671
rect 1251 -1778 1280 -1684
rect 1326 -1778 1355 -1684
rect 1251 -1791 1355 -1778
rect 1455 -1684 1559 -1671
rect 1455 -1778 1484 -1684
rect 1530 -1778 1559 -1684
rect 1455 -1791 1559 -1778
rect 1659 -1684 1763 -1671
rect 1659 -1778 1688 -1684
rect 1734 -1778 1763 -1684
rect 1659 -1791 1763 -1778
rect 1863 -1684 1951 -1671
rect 1863 -1778 1892 -1684
rect 1938 -1778 1951 -1684
rect 1863 -1791 1951 -1778
rect 2056 -1684 2144 -1671
rect 2056 -1778 2069 -1684
rect 2115 -1778 2144 -1684
rect 2056 -1791 2144 -1778
rect 2244 -1684 2332 -1671
rect 2244 -1778 2273 -1684
rect 2319 -1778 2332 -1684
rect 2244 -1791 2332 -1778
rect 3501 -1919 3589 -1906
rect 3501 -2013 3514 -1919
rect 3560 -2013 3589 -1919
rect 3501 -2026 3589 -2013
rect 3689 -1919 3793 -1906
rect 3689 -2013 3718 -1919
rect 3764 -2013 3793 -1919
rect 3689 -2026 3793 -2013
rect 3893 -1919 3981 -1906
rect 3893 -2013 3922 -1919
rect 3968 -2013 3981 -1919
rect 3893 -2026 3981 -2013
rect 4037 -1919 4125 -1906
rect 4037 -2013 4050 -1919
rect 4096 -2013 4125 -1919
rect 4037 -2026 4125 -2013
rect 4225 -1919 4329 -1906
rect 4225 -2013 4254 -1919
rect 4300 -2013 4329 -1919
rect 4225 -2026 4329 -2013
rect 4429 -1919 4517 -1906
rect 4429 -2013 4458 -1919
rect 4504 -2013 4517 -1919
rect 4429 -2026 4517 -2013
rect 4573 -1919 4661 -1906
rect 4573 -2013 4586 -1919
rect 4632 -2013 4661 -1919
rect 4573 -2026 4661 -2013
rect 4761 -1919 4865 -1906
rect 4761 -2013 4790 -1919
rect 4836 -2013 4865 -1919
rect 4761 -2026 4865 -2013
rect 4965 -1919 5053 -1906
rect 4965 -2013 4994 -1919
rect 5040 -2013 5053 -1919
rect 4965 -2026 5053 -2013
rect 5109 -1919 5197 -1906
rect 5109 -2013 5122 -1919
rect 5168 -2013 5197 -1919
rect 5109 -2026 5197 -2013
rect 5297 -1919 5401 -1906
rect 5297 -2013 5326 -1919
rect 5372 -2013 5401 -1919
rect 5297 -2026 5401 -2013
rect 5501 -1919 5589 -1906
rect 5501 -2013 5530 -1919
rect 5576 -2013 5589 -1919
rect 5501 -2026 5589 -2013
rect 5645 -1919 5733 -1906
rect 5645 -2013 5658 -1919
rect 5704 -2013 5733 -1919
rect 5645 -2026 5733 -2013
rect 5833 -1919 5937 -1906
rect 5833 -2013 5862 -1919
rect 5908 -2013 5937 -1919
rect 5833 -2026 5937 -2013
rect 6037 -1919 6125 -1906
rect 6037 -2013 6066 -1919
rect 6112 -2013 6125 -1919
rect 6037 -2026 6125 -2013
rect 3501 -2303 3589 -2290
rect 3501 -2397 3514 -2303
rect 3560 -2397 3589 -2303
rect 3501 -2410 3589 -2397
rect 3689 -2303 3793 -2290
rect 3689 -2397 3718 -2303
rect 3764 -2397 3793 -2303
rect 3689 -2410 3793 -2397
rect 3893 -2303 3981 -2290
rect 3893 -2397 3922 -2303
rect 3968 -2397 3981 -2303
rect 3893 -2410 3981 -2397
rect 4037 -2303 4125 -2290
rect 4037 -2397 4050 -2303
rect 4096 -2397 4125 -2303
rect 4037 -2410 4125 -2397
rect 4225 -2303 4329 -2290
rect 4225 -2397 4254 -2303
rect 4300 -2397 4329 -2303
rect 4225 -2410 4329 -2397
rect 4429 -2303 4517 -2290
rect 4429 -2397 4458 -2303
rect 4504 -2397 4517 -2303
rect 4429 -2410 4517 -2397
rect 4573 -2303 4661 -2290
rect 4573 -2397 4586 -2303
rect 4632 -2397 4661 -2303
rect 4573 -2410 4661 -2397
rect 4761 -2303 4865 -2290
rect 4761 -2397 4790 -2303
rect 4836 -2397 4865 -2303
rect 4761 -2410 4865 -2397
rect 4965 -2303 5053 -2290
rect 4965 -2397 4994 -2303
rect 5040 -2397 5053 -2303
rect 4965 -2410 5053 -2397
rect 5109 -2303 5197 -2290
rect 5109 -2397 5122 -2303
rect 5168 -2397 5197 -2303
rect 5109 -2410 5197 -2397
rect 5297 -2303 5401 -2290
rect 5297 -2397 5326 -2303
rect 5372 -2397 5401 -2303
rect 5297 -2410 5401 -2397
rect 5501 -2303 5589 -2290
rect 5501 -2397 5530 -2303
rect 5576 -2397 5589 -2303
rect 5501 -2410 5589 -2397
rect 5645 -2303 5733 -2290
rect 5645 -2397 5658 -2303
rect 5704 -2397 5733 -2303
rect 5645 -2410 5733 -2397
rect 5833 -2303 5937 -2290
rect 5833 -2397 5862 -2303
rect 5908 -2397 5937 -2303
rect 5833 -2410 5937 -2397
rect 6037 -2303 6125 -2290
rect 6037 -2397 6066 -2303
rect 6112 -2397 6125 -2303
rect 6037 -2410 6125 -2397
rect -67 -2902 21 -2889
rect -67 -2996 -54 -2902
rect -8 -2996 21 -2902
rect -67 -3009 21 -2996
rect 121 -2902 225 -2889
rect 121 -2996 150 -2902
rect 196 -2996 225 -2902
rect 121 -3009 225 -2996
rect 325 -2902 413 -2889
rect 325 -2996 354 -2902
rect 400 -2996 413 -2902
rect 325 -3009 413 -2996
rect 469 -2902 557 -2889
rect 469 -2996 482 -2902
rect 528 -2996 557 -2902
rect 469 -3009 557 -2996
rect 657 -2902 761 -2889
rect 657 -2996 686 -2902
rect 732 -2996 761 -2902
rect 657 -3009 761 -2996
rect 861 -2902 949 -2889
rect 861 -2996 890 -2902
rect 936 -2996 949 -2902
rect 861 -3009 949 -2996
rect 1005 -2902 1093 -2889
rect 1005 -2996 1018 -2902
rect 1064 -2996 1093 -2902
rect 1005 -3009 1093 -2996
rect 1193 -2902 1297 -2889
rect 1193 -2996 1222 -2902
rect 1268 -2996 1297 -2902
rect 1193 -3009 1297 -2996
rect 1397 -2902 1485 -2889
rect 1397 -2996 1426 -2902
rect 1472 -2996 1485 -2902
rect 1397 -3009 1485 -2996
rect 1541 -2902 1629 -2889
rect 1541 -2996 1554 -2902
rect 1600 -2996 1629 -2902
rect 1541 -3009 1629 -2996
rect 1729 -2902 1833 -2889
rect 1729 -2996 1758 -2902
rect 1804 -2996 1833 -2902
rect 1729 -3009 1833 -2996
rect 1933 -2902 2021 -2889
rect 1933 -2996 1962 -2902
rect 2008 -2996 2021 -2902
rect 1933 -3009 2021 -2996
rect 2077 -2902 2165 -2889
rect 2077 -2996 2090 -2902
rect 2136 -2996 2165 -2902
rect 2077 -3009 2165 -2996
rect 2265 -2902 2369 -2889
rect 2265 -2996 2294 -2902
rect 2340 -2996 2369 -2902
rect 2265 -3009 2369 -2996
rect 2469 -2902 2557 -2889
rect 2469 -2996 2498 -2902
rect 2544 -2996 2557 -2902
rect 2469 -3009 2557 -2996
rect -2062 -3411 -1990 -3400
rect -67 -3186 21 -3173
rect -67 -3280 -54 -3186
rect -8 -3280 21 -3186
rect -67 -3293 21 -3280
rect 121 -3186 225 -3173
rect 121 -3280 150 -3186
rect 196 -3280 225 -3186
rect 121 -3293 225 -3280
rect 325 -3186 413 -3173
rect 325 -3280 354 -3186
rect 400 -3280 413 -3186
rect 325 -3293 413 -3280
rect 469 -3186 557 -3173
rect 469 -3280 482 -3186
rect 528 -3280 557 -3186
rect 469 -3293 557 -3280
rect 657 -3186 761 -3173
rect 657 -3280 686 -3186
rect 732 -3280 761 -3186
rect 657 -3293 761 -3280
rect 861 -3186 949 -3173
rect 861 -3280 890 -3186
rect 936 -3280 949 -3186
rect 861 -3293 949 -3280
rect 1005 -3186 1093 -3173
rect 1005 -3280 1018 -3186
rect 1064 -3280 1093 -3186
rect 1005 -3293 1093 -3280
rect 1193 -3186 1297 -3173
rect 1193 -3280 1222 -3186
rect 1268 -3280 1297 -3186
rect 1193 -3293 1297 -3280
rect 1397 -3186 1485 -3173
rect 1397 -3280 1426 -3186
rect 1472 -3280 1485 -3186
rect 1397 -3293 1485 -3280
rect 1541 -3186 1629 -3173
rect 1541 -3280 1554 -3186
rect 1600 -3280 1629 -3186
rect 1541 -3293 1629 -3280
rect 1729 -3186 1833 -3173
rect 1729 -3280 1758 -3186
rect 1804 -3280 1833 -3186
rect 1729 -3293 1833 -3280
rect 1933 -3186 2021 -3173
rect 1933 -3280 1962 -3186
rect 2008 -3280 2021 -3186
rect 1933 -3293 2021 -3280
rect 2077 -3186 2165 -3173
rect 2077 -3280 2090 -3186
rect 2136 -3280 2165 -3186
rect 2077 -3293 2165 -3280
rect 2265 -3186 2369 -3173
rect 2265 -3280 2294 -3186
rect 2340 -3280 2369 -3186
rect 2265 -3293 2369 -3280
rect 2469 -3186 2557 -3173
rect 2469 -3280 2498 -3186
rect 2544 -3280 2557 -3186
rect 2469 -3293 2557 -3280
rect -1894 -3411 -1822 -3400
rect -2062 -3413 -1970 -3411
rect -2062 -3459 -2049 -3413
rect -2003 -3459 -1970 -3413
rect -2062 -3461 -1970 -3459
rect -1914 -3413 -1822 -3411
rect -1914 -3459 -1881 -3413
rect -1835 -3459 -1822 -3413
rect -1584 -3415 -1512 -3402
rect -1914 -3461 -1822 -3459
rect -2062 -3472 -1990 -3461
rect -1894 -3472 -1822 -3461
rect -1584 -3461 -1571 -3415
rect -1525 -3416 -1512 -3415
rect -1416 -3415 -1344 -3402
rect -1416 -3416 -1403 -3415
rect -1525 -3460 -1492 -3416
rect -1436 -3460 -1403 -3416
rect -1525 -3461 -1512 -3460
rect -1584 -3474 -1512 -3461
rect -1416 -3461 -1403 -3460
rect -1357 -3461 -1344 -3415
rect -1416 -3474 -1344 -3461
rect -1048 -3415 -976 -3402
rect -1048 -3461 -1035 -3415
rect -989 -3416 -976 -3415
rect -880 -3415 -808 -3402
rect -880 -3416 -867 -3415
rect -989 -3460 -956 -3416
rect -900 -3460 -867 -3416
rect -989 -3461 -976 -3460
rect -1048 -3474 -976 -3461
rect -880 -3461 -867 -3460
rect -821 -3461 -808 -3415
rect -880 -3474 -808 -3461
rect -67 -3718 21 -3705
rect -67 -3812 -54 -3718
rect -8 -3812 21 -3718
rect -67 -3825 21 -3812
rect 121 -3718 225 -3705
rect 121 -3812 150 -3718
rect 196 -3812 225 -3718
rect 121 -3825 225 -3812
rect 325 -3718 429 -3705
rect 325 -3812 354 -3718
rect 400 -3812 429 -3718
rect 325 -3825 429 -3812
rect 529 -3718 633 -3705
rect 529 -3812 558 -3718
rect 604 -3812 633 -3718
rect 529 -3825 633 -3812
rect 733 -3718 837 -3705
rect 733 -3812 762 -3718
rect 808 -3812 837 -3718
rect 733 -3825 837 -3812
rect 937 -3718 1041 -3705
rect 937 -3812 966 -3718
rect 1012 -3812 1041 -3718
rect 937 -3825 1041 -3812
rect 1141 -3718 1245 -3705
rect 1141 -3812 1170 -3718
rect 1216 -3812 1245 -3718
rect 1141 -3825 1245 -3812
rect 1345 -3718 1449 -3705
rect 1345 -3812 1374 -3718
rect 1420 -3812 1449 -3718
rect 1345 -3825 1449 -3812
rect 1549 -3718 1653 -3705
rect 1549 -3812 1578 -3718
rect 1624 -3812 1653 -3718
rect 1549 -3825 1653 -3812
rect 1753 -3718 1857 -3705
rect 1753 -3812 1782 -3718
rect 1828 -3812 1857 -3718
rect 1753 -3825 1857 -3812
rect 1957 -3718 2045 -3705
rect 1957 -3812 1986 -3718
rect 2032 -3812 2045 -3718
rect 1957 -3825 2045 -3812
rect 2101 -3718 2189 -3705
rect 2101 -3812 2114 -3718
rect 2160 -3812 2189 -3718
rect 2101 -3825 2189 -3812
rect 2289 -3718 2393 -3705
rect 2289 -3812 2318 -3718
rect 2364 -3812 2393 -3718
rect 2289 -3825 2393 -3812
rect 2493 -3718 2581 -3705
rect 2493 -3812 2522 -3718
rect 2568 -3812 2581 -3718
rect 2493 -3825 2581 -3812
rect -2062 -4279 -1990 -4268
rect -1894 -4279 -1822 -4268
rect -2062 -4281 -1970 -4279
rect -2062 -4327 -2049 -4281
rect -2003 -4327 -1970 -4281
rect -2062 -4329 -1970 -4327
rect -1914 -4281 -1822 -4279
rect -1914 -4327 -1881 -4281
rect -1835 -4327 -1822 -4281
rect -1584 -4283 -1512 -4270
rect -1914 -4329 -1822 -4327
rect -2062 -4340 -1990 -4329
rect -1894 -4340 -1822 -4329
rect -1584 -4329 -1571 -4283
rect -1525 -4284 -1512 -4283
rect -1416 -4283 -1344 -4270
rect -1416 -4284 -1403 -4283
rect -1525 -4328 -1492 -4284
rect -1436 -4328 -1403 -4284
rect -1525 -4329 -1512 -4328
rect -1584 -4342 -1512 -4329
rect -1416 -4329 -1403 -4328
rect -1357 -4329 -1344 -4283
rect -1416 -4342 -1344 -4329
rect -1048 -4283 -976 -4270
rect -1048 -4329 -1035 -4283
rect -989 -4284 -976 -4283
rect -67 -4107 21 -4094
rect -67 -4201 -54 -4107
rect -8 -4201 21 -4107
rect -67 -4214 21 -4201
rect 121 -4107 225 -4094
rect 121 -4201 150 -4107
rect 196 -4201 225 -4107
rect 121 -4214 225 -4201
rect 325 -4107 429 -4094
rect 325 -4201 354 -4107
rect 400 -4201 429 -4107
rect 325 -4214 429 -4201
rect 529 -4107 633 -4094
rect 529 -4201 558 -4107
rect 604 -4201 633 -4107
rect 529 -4214 633 -4201
rect 733 -4107 837 -4094
rect 733 -4201 762 -4107
rect 808 -4201 837 -4107
rect 733 -4214 837 -4201
rect 937 -4107 1041 -4094
rect 937 -4201 966 -4107
rect 1012 -4201 1041 -4107
rect 937 -4214 1041 -4201
rect 1141 -4107 1245 -4094
rect 1141 -4201 1170 -4107
rect 1216 -4201 1245 -4107
rect 1141 -4214 1245 -4201
rect 1345 -4107 1449 -4094
rect 1345 -4201 1374 -4107
rect 1420 -4201 1449 -4107
rect 1345 -4214 1449 -4201
rect 1549 -4107 1653 -4094
rect 1549 -4201 1578 -4107
rect 1624 -4201 1653 -4107
rect 1549 -4214 1653 -4201
rect 1753 -4107 1857 -4094
rect 1753 -4201 1782 -4107
rect 1828 -4201 1857 -4107
rect 1753 -4214 1857 -4201
rect 1957 -4107 2045 -4094
rect 1957 -4201 1986 -4107
rect 2032 -4201 2045 -4107
rect 1957 -4214 2045 -4201
rect 2101 -4107 2189 -4094
rect 2101 -4201 2114 -4107
rect 2160 -4201 2189 -4107
rect 2101 -4214 2189 -4201
rect 2289 -4107 2393 -4094
rect 2289 -4201 2318 -4107
rect 2364 -4201 2393 -4107
rect 2289 -4214 2393 -4201
rect 2493 -4107 2581 -4094
rect 2493 -4201 2522 -4107
rect 2568 -4201 2581 -4107
rect 2493 -4214 2581 -4201
rect -880 -4283 -808 -4270
rect -880 -4284 -867 -4283
rect -989 -4328 -956 -4284
rect -900 -4328 -867 -4284
rect -989 -4329 -976 -4328
rect -1048 -4342 -976 -4329
rect -880 -4329 -867 -4328
rect -821 -4329 -808 -4283
rect -880 -4342 -808 -4329
rect -67 -4402 21 -4389
rect -67 -4496 -54 -4402
rect -8 -4496 21 -4402
rect -67 -4509 21 -4496
rect 121 -4402 225 -4389
rect 121 -4496 150 -4402
rect 196 -4496 225 -4402
rect 121 -4509 225 -4496
rect 325 -4402 429 -4389
rect 325 -4496 354 -4402
rect 400 -4496 429 -4402
rect 325 -4509 429 -4496
rect 529 -4402 633 -4389
rect 529 -4496 558 -4402
rect 604 -4496 633 -4402
rect 529 -4509 633 -4496
rect 733 -4402 837 -4389
rect 733 -4496 762 -4402
rect 808 -4496 837 -4402
rect 733 -4509 837 -4496
rect 937 -4402 1041 -4389
rect 937 -4496 966 -4402
rect 1012 -4496 1041 -4402
rect 937 -4509 1041 -4496
rect 1141 -4402 1245 -4389
rect 1141 -4496 1170 -4402
rect 1216 -4496 1245 -4402
rect 1141 -4509 1245 -4496
rect 1345 -4402 1449 -4389
rect 1345 -4496 1374 -4402
rect 1420 -4496 1449 -4402
rect 1345 -4509 1449 -4496
rect 1549 -4402 1653 -4389
rect 1549 -4496 1578 -4402
rect 1624 -4496 1653 -4402
rect 1549 -4509 1653 -4496
rect 1753 -4402 1857 -4389
rect 1753 -4496 1782 -4402
rect 1828 -4496 1857 -4402
rect 1753 -4509 1857 -4496
rect 1957 -4402 2045 -4389
rect 1957 -4496 1986 -4402
rect 2032 -4496 2045 -4402
rect 1957 -4509 2045 -4496
rect 2101 -4402 2189 -4389
rect 2101 -4496 2114 -4402
rect 2160 -4496 2189 -4402
rect 2101 -4509 2189 -4496
rect 2289 -4402 2393 -4389
rect 2289 -4496 2318 -4402
rect 2364 -4496 2393 -4402
rect 2289 -4509 2393 -4496
rect 2493 -4402 2581 -4389
rect 2493 -4496 2522 -4402
rect 2568 -4496 2581 -4402
rect 2493 -4509 2581 -4496
rect -67 -4787 21 -4774
rect -67 -4881 -54 -4787
rect -8 -4881 21 -4787
rect -67 -4894 21 -4881
rect 121 -4787 225 -4774
rect 121 -4881 150 -4787
rect 196 -4881 225 -4787
rect 121 -4894 225 -4881
rect 325 -4787 429 -4774
rect 325 -4881 354 -4787
rect 400 -4881 429 -4787
rect 325 -4894 429 -4881
rect 529 -4787 633 -4774
rect 529 -4881 558 -4787
rect 604 -4881 633 -4787
rect 529 -4894 633 -4881
rect 733 -4787 837 -4774
rect 733 -4881 762 -4787
rect 808 -4881 837 -4787
rect 733 -4894 837 -4881
rect 937 -4787 1041 -4774
rect 937 -4881 966 -4787
rect 1012 -4881 1041 -4787
rect 937 -4894 1041 -4881
rect 1141 -4787 1245 -4774
rect 1141 -4881 1170 -4787
rect 1216 -4881 1245 -4787
rect 1141 -4894 1245 -4881
rect 1345 -4787 1449 -4774
rect 1345 -4881 1374 -4787
rect 1420 -4881 1449 -4787
rect 1345 -4894 1449 -4881
rect 1549 -4787 1653 -4774
rect 1549 -4881 1578 -4787
rect 1624 -4881 1653 -4787
rect 1549 -4894 1653 -4881
rect 1753 -4787 1857 -4774
rect 1753 -4881 1782 -4787
rect 1828 -4881 1857 -4787
rect 1753 -4894 1857 -4881
rect 1957 -4787 2045 -4774
rect 1957 -4881 1986 -4787
rect 2032 -4881 2045 -4787
rect 1957 -4894 2045 -4881
rect 2101 -4787 2189 -4774
rect 2101 -4881 2114 -4787
rect 2160 -4881 2189 -4787
rect 2101 -4894 2189 -4881
rect 2289 -4787 2393 -4774
rect 2289 -4881 2318 -4787
rect 2364 -4881 2393 -4787
rect 2289 -4894 2393 -4881
rect 2493 -4787 2581 -4774
rect 2493 -4881 2522 -4787
rect 2568 -4881 2581 -4787
rect 2493 -4894 2581 -4881
rect -2062 -5138 -1990 -5127
rect -1894 -5138 -1822 -5127
rect -2062 -5140 -1970 -5138
rect -2062 -5186 -2049 -5140
rect -2003 -5186 -1970 -5140
rect -2062 -5188 -1970 -5186
rect -1914 -5140 -1822 -5138
rect -1914 -5186 -1881 -5140
rect -1835 -5186 -1822 -5140
rect -1584 -5142 -1512 -5129
rect -1914 -5188 -1822 -5186
rect -2062 -5199 -1990 -5188
rect -1894 -5199 -1822 -5188
rect -1584 -5188 -1571 -5142
rect -1525 -5143 -1512 -5142
rect -1416 -5142 -1344 -5129
rect -1416 -5143 -1403 -5142
rect -1525 -5187 -1492 -5143
rect -1436 -5187 -1403 -5143
rect -1525 -5188 -1512 -5187
rect -1584 -5201 -1512 -5188
rect -1416 -5188 -1403 -5187
rect -1357 -5188 -1344 -5142
rect -1416 -5201 -1344 -5188
rect -1048 -5142 -976 -5129
rect -1048 -5188 -1035 -5142
rect -989 -5143 -976 -5142
rect -880 -5142 -808 -5129
rect -880 -5143 -867 -5142
rect -989 -5187 -956 -5143
rect -900 -5187 -867 -5143
rect -989 -5188 -976 -5187
rect -1048 -5201 -976 -5188
rect -880 -5188 -867 -5187
rect -821 -5188 -808 -5142
rect -880 -5201 -808 -5188
rect 3501 -2593 3589 -2580
rect 3501 -2687 3514 -2593
rect 3560 -2687 3589 -2593
rect 3501 -2700 3589 -2687
rect 3689 -2593 3793 -2580
rect 3689 -2687 3718 -2593
rect 3764 -2687 3793 -2593
rect 3689 -2700 3793 -2687
rect 3893 -2593 3981 -2580
rect 3893 -2687 3922 -2593
rect 3968 -2687 3981 -2593
rect 3893 -2700 3981 -2687
rect 4037 -2593 4125 -2580
rect 4037 -2687 4050 -2593
rect 4096 -2687 4125 -2593
rect 4037 -2700 4125 -2687
rect 4225 -2593 4329 -2580
rect 4225 -2687 4254 -2593
rect 4300 -2687 4329 -2593
rect 4225 -2700 4329 -2687
rect 4429 -2593 4517 -2580
rect 4429 -2687 4458 -2593
rect 4504 -2687 4517 -2593
rect 4429 -2700 4517 -2687
rect 4573 -2593 4661 -2580
rect 4573 -2687 4586 -2593
rect 4632 -2687 4661 -2593
rect 4573 -2700 4661 -2687
rect 4761 -2593 4865 -2580
rect 4761 -2687 4790 -2593
rect 4836 -2687 4865 -2593
rect 4761 -2700 4865 -2687
rect 4965 -2593 5053 -2580
rect 4965 -2687 4994 -2593
rect 5040 -2687 5053 -2593
rect 4965 -2700 5053 -2687
rect 5109 -2593 5197 -2580
rect 5109 -2687 5122 -2593
rect 5168 -2687 5197 -2593
rect 5109 -2700 5197 -2687
rect 5297 -2593 5401 -2580
rect 5297 -2687 5326 -2593
rect 5372 -2687 5401 -2593
rect 5297 -2700 5401 -2687
rect 5501 -2593 5589 -2580
rect 5501 -2687 5530 -2593
rect 5576 -2687 5589 -2593
rect 5501 -2700 5589 -2687
rect 5645 -2593 5733 -2580
rect 5645 -2687 5658 -2593
rect 5704 -2687 5733 -2593
rect 5645 -2700 5733 -2687
rect 5833 -2593 5937 -2580
rect 5833 -2687 5862 -2593
rect 5908 -2687 5937 -2593
rect 5833 -2700 5937 -2687
rect 6037 -2593 6125 -2580
rect 6037 -2687 6066 -2593
rect 6112 -2687 6125 -2593
rect 6037 -2700 6125 -2687
rect 3501 -2977 3589 -2964
rect 3501 -3071 3514 -2977
rect 3560 -3071 3589 -2977
rect 3501 -3084 3589 -3071
rect 3689 -2977 3793 -2964
rect 3689 -3071 3718 -2977
rect 3764 -3071 3793 -2977
rect 3689 -3084 3793 -3071
rect 3893 -2977 3981 -2964
rect 3893 -3071 3922 -2977
rect 3968 -3071 3981 -2977
rect 3893 -3084 3981 -3071
rect 4037 -2977 4125 -2964
rect 4037 -3071 4050 -2977
rect 4096 -3071 4125 -2977
rect 4037 -3084 4125 -3071
rect 4225 -2977 4329 -2964
rect 4225 -3071 4254 -2977
rect 4300 -3071 4329 -2977
rect 4225 -3084 4329 -3071
rect 4429 -2977 4517 -2964
rect 4429 -3071 4458 -2977
rect 4504 -3071 4517 -2977
rect 4429 -3084 4517 -3071
rect 4573 -2977 4661 -2964
rect 4573 -3071 4586 -2977
rect 4632 -3071 4661 -2977
rect 4573 -3084 4661 -3071
rect 4761 -2977 4865 -2964
rect 4761 -3071 4790 -2977
rect 4836 -3071 4865 -2977
rect 4761 -3084 4865 -3071
rect 4965 -2977 5053 -2964
rect 4965 -3071 4994 -2977
rect 5040 -3071 5053 -2977
rect 4965 -3084 5053 -3071
rect 5109 -2977 5197 -2964
rect 5109 -3071 5122 -2977
rect 5168 -3071 5197 -2977
rect 5109 -3084 5197 -3071
rect 5297 -2977 5401 -2964
rect 5297 -3071 5326 -2977
rect 5372 -3071 5401 -2977
rect 5297 -3084 5401 -3071
rect 5501 -2977 5589 -2964
rect 5501 -3071 5530 -2977
rect 5576 -3071 5589 -2977
rect 5501 -3084 5589 -3071
rect 5645 -2977 5733 -2964
rect 5645 -3071 5658 -2977
rect 5704 -3071 5733 -2977
rect 5645 -3084 5733 -3071
rect 5833 -2977 5937 -2964
rect 5833 -3071 5862 -2977
rect 5908 -3071 5937 -2977
rect 5833 -3084 5937 -3071
rect 6037 -2977 6125 -2964
rect 6037 -3071 6066 -2977
rect 6112 -3071 6125 -2977
rect 6037 -3084 6125 -3071
rect 3501 -3611 3589 -3598
rect 3501 -3705 3514 -3611
rect 3560 -3705 3589 -3611
rect 3501 -3718 3589 -3705
rect 3689 -3611 3793 -3598
rect 3689 -3705 3718 -3611
rect 3764 -3705 3793 -3611
rect 3689 -3718 3793 -3705
rect 3893 -3611 3997 -3598
rect 3893 -3705 3922 -3611
rect 3968 -3705 3997 -3611
rect 3893 -3718 3997 -3705
rect 4097 -3611 4201 -3598
rect 4097 -3705 4126 -3611
rect 4172 -3705 4201 -3611
rect 4097 -3718 4201 -3705
rect 4301 -3611 4405 -3598
rect 4301 -3705 4330 -3611
rect 4376 -3705 4405 -3611
rect 4301 -3718 4405 -3705
rect 4505 -3611 4609 -3598
rect 4505 -3705 4534 -3611
rect 4580 -3705 4609 -3611
rect 4505 -3718 4609 -3705
rect 4709 -3611 4813 -3598
rect 4709 -3705 4738 -3611
rect 4784 -3705 4813 -3611
rect 4709 -3718 4813 -3705
rect 4913 -3611 5017 -3598
rect 4913 -3705 4942 -3611
rect 4988 -3705 5017 -3611
rect 4913 -3718 5017 -3705
rect 5117 -3611 5221 -3598
rect 5117 -3705 5146 -3611
rect 5192 -3705 5221 -3611
rect 5117 -3718 5221 -3705
rect 5321 -3611 5425 -3598
rect 5321 -3705 5350 -3611
rect 5396 -3705 5425 -3611
rect 5321 -3718 5425 -3705
rect 5525 -3611 5613 -3598
rect 5525 -3705 5554 -3611
rect 5600 -3705 5613 -3611
rect 5525 -3718 5613 -3705
rect 5669 -3611 5757 -3598
rect 5669 -3705 5682 -3611
rect 5728 -3705 5757 -3611
rect 5669 -3718 5757 -3705
rect 5857 -3611 5961 -3598
rect 5857 -3705 5886 -3611
rect 5932 -3705 5961 -3611
rect 5857 -3718 5961 -3705
rect 6061 -3611 6149 -3598
rect 6061 -3705 6090 -3611
rect 6136 -3705 6149 -3611
rect 6061 -3718 6149 -3705
rect 3501 -4000 3589 -3987
rect 3501 -4094 3514 -4000
rect 3560 -4094 3589 -4000
rect 3501 -4107 3589 -4094
rect 3689 -4000 3793 -3987
rect 3689 -4094 3718 -4000
rect 3764 -4094 3793 -4000
rect 3689 -4107 3793 -4094
rect 3893 -4000 3997 -3987
rect 3893 -4094 3922 -4000
rect 3968 -4094 3997 -4000
rect 3893 -4107 3997 -4094
rect 4097 -4000 4201 -3987
rect 4097 -4094 4126 -4000
rect 4172 -4094 4201 -4000
rect 4097 -4107 4201 -4094
rect 4301 -4000 4405 -3987
rect 4301 -4094 4330 -4000
rect 4376 -4094 4405 -4000
rect 4301 -4107 4405 -4094
rect 4505 -4000 4609 -3987
rect 4505 -4094 4534 -4000
rect 4580 -4094 4609 -4000
rect 4505 -4107 4609 -4094
rect 4709 -4000 4813 -3987
rect 4709 -4094 4738 -4000
rect 4784 -4094 4813 -4000
rect 4709 -4107 4813 -4094
rect 4913 -4000 5017 -3987
rect 4913 -4094 4942 -4000
rect 4988 -4094 5017 -4000
rect 4913 -4107 5017 -4094
rect 5117 -4000 5221 -3987
rect 5117 -4094 5146 -4000
rect 5192 -4094 5221 -4000
rect 5117 -4107 5221 -4094
rect 5321 -4000 5425 -3987
rect 5321 -4094 5350 -4000
rect 5396 -4094 5425 -4000
rect 5321 -4107 5425 -4094
rect 5525 -4000 5613 -3987
rect 5525 -4094 5554 -4000
rect 5600 -4094 5613 -4000
rect 5525 -4107 5613 -4094
rect 5669 -4000 5757 -3987
rect 5669 -4094 5682 -4000
rect 5728 -4094 5757 -4000
rect 5669 -4107 5757 -4094
rect 5857 -4000 5961 -3987
rect 5857 -4094 5886 -4000
rect 5932 -4094 5961 -4000
rect 5857 -4107 5961 -4094
rect 6061 -4000 6149 -3987
rect 6061 -4094 6090 -4000
rect 6136 -4094 6149 -4000
rect 6061 -4107 6149 -4094
rect 3501 -4295 3589 -4282
rect 3501 -4389 3514 -4295
rect 3560 -4389 3589 -4295
rect 3501 -4402 3589 -4389
rect 3689 -4295 3793 -4282
rect 3689 -4389 3718 -4295
rect 3764 -4389 3793 -4295
rect 3689 -4402 3793 -4389
rect 3893 -4295 3997 -4282
rect 3893 -4389 3922 -4295
rect 3968 -4389 3997 -4295
rect 3893 -4402 3997 -4389
rect 4097 -4295 4201 -4282
rect 4097 -4389 4126 -4295
rect 4172 -4389 4201 -4295
rect 4097 -4402 4201 -4389
rect 4301 -4295 4405 -4282
rect 4301 -4389 4330 -4295
rect 4376 -4389 4405 -4295
rect 4301 -4402 4405 -4389
rect 4505 -4295 4609 -4282
rect 4505 -4389 4534 -4295
rect 4580 -4389 4609 -4295
rect 4505 -4402 4609 -4389
rect 4709 -4295 4813 -4282
rect 4709 -4389 4738 -4295
rect 4784 -4389 4813 -4295
rect 4709 -4402 4813 -4389
rect 4913 -4295 5017 -4282
rect 4913 -4389 4942 -4295
rect 4988 -4389 5017 -4295
rect 4913 -4402 5017 -4389
rect 5117 -4295 5221 -4282
rect 5117 -4389 5146 -4295
rect 5192 -4389 5221 -4295
rect 5117 -4402 5221 -4389
rect 5321 -4295 5425 -4282
rect 5321 -4389 5350 -4295
rect 5396 -4389 5425 -4295
rect 5321 -4402 5425 -4389
rect 5525 -4295 5613 -4282
rect 5525 -4389 5554 -4295
rect 5600 -4389 5613 -4295
rect 5525 -4402 5613 -4389
rect 5669 -4295 5757 -4282
rect 5669 -4389 5682 -4295
rect 5728 -4389 5757 -4295
rect 5669 -4402 5757 -4389
rect 5857 -4295 5961 -4282
rect 5857 -4389 5886 -4295
rect 5932 -4389 5961 -4295
rect 5857 -4402 5961 -4389
rect 6061 -4295 6149 -4282
rect 6061 -4389 6090 -4295
rect 6136 -4389 6149 -4295
rect 6061 -4402 6149 -4389
rect 3501 -4680 3589 -4667
rect 3501 -4774 3514 -4680
rect 3560 -4774 3589 -4680
rect 3501 -4787 3589 -4774
rect 3689 -4680 3793 -4667
rect 3689 -4774 3718 -4680
rect 3764 -4774 3793 -4680
rect 3689 -4787 3793 -4774
rect 3893 -4680 3997 -4667
rect 3893 -4774 3922 -4680
rect 3968 -4774 3997 -4680
rect 3893 -4787 3997 -4774
rect 4097 -4680 4201 -4667
rect 4097 -4774 4126 -4680
rect 4172 -4774 4201 -4680
rect 4097 -4787 4201 -4774
rect 4301 -4680 4405 -4667
rect 4301 -4774 4330 -4680
rect 4376 -4774 4405 -4680
rect 4301 -4787 4405 -4774
rect 4505 -4680 4609 -4667
rect 4505 -4774 4534 -4680
rect 4580 -4774 4609 -4680
rect 4505 -4787 4609 -4774
rect 4709 -4680 4813 -4667
rect 4709 -4774 4738 -4680
rect 4784 -4774 4813 -4680
rect 4709 -4787 4813 -4774
rect 4913 -4680 5017 -4667
rect 4913 -4774 4942 -4680
rect 4988 -4774 5017 -4680
rect 4913 -4787 5017 -4774
rect 5117 -4680 5221 -4667
rect 5117 -4774 5146 -4680
rect 5192 -4774 5221 -4680
rect 5117 -4787 5221 -4774
rect 5321 -4680 5425 -4667
rect 5321 -4774 5350 -4680
rect 5396 -4774 5425 -4680
rect 5321 -4787 5425 -4774
rect 5525 -4680 5613 -4667
rect 5525 -4774 5554 -4680
rect 5600 -4774 5613 -4680
rect 5525 -4787 5613 -4774
rect 5669 -4680 5757 -4667
rect 5669 -4774 5682 -4680
rect 5728 -4774 5757 -4680
rect 5669 -4787 5757 -4774
rect 5857 -4680 5961 -4667
rect 5857 -4774 5886 -4680
rect 5932 -4774 5961 -4680
rect 5857 -4787 5961 -4774
rect 6061 -4680 6149 -4667
rect 6061 -4774 6090 -4680
rect 6136 -4774 6149 -4680
rect 6061 -4787 6149 -4774
rect 3501 -5007 3589 -4994
rect 3501 -5101 3514 -5007
rect 3560 -5101 3589 -5007
rect 3501 -5114 3589 -5101
rect 3689 -5007 3793 -4994
rect 3689 -5101 3718 -5007
rect 3764 -5101 3793 -5007
rect 3689 -5114 3793 -5101
rect 3893 -5007 3997 -4994
rect 3893 -5101 3922 -5007
rect 3968 -5101 3997 -5007
rect 3893 -5114 3997 -5101
rect 4097 -5007 4201 -4994
rect 4097 -5101 4126 -5007
rect 4172 -5101 4201 -5007
rect 4097 -5114 4201 -5101
rect 4301 -5007 4405 -4994
rect 4301 -5101 4330 -5007
rect 4376 -5101 4405 -5007
rect 4301 -5114 4405 -5101
rect 4505 -5007 4609 -4994
rect 4505 -5101 4534 -5007
rect 4580 -5101 4609 -5007
rect 4505 -5114 4609 -5101
rect 4709 -5007 4813 -4994
rect 4709 -5101 4738 -5007
rect 4784 -5101 4813 -5007
rect 4709 -5114 4813 -5101
rect 4913 -5007 5017 -4994
rect 4913 -5101 4942 -5007
rect 4988 -5101 5017 -5007
rect 4913 -5114 5017 -5101
rect 5117 -5007 5221 -4994
rect 5117 -5101 5146 -5007
rect 5192 -5101 5221 -5007
rect 5117 -5114 5221 -5101
rect 5321 -5007 5425 -4994
rect 5321 -5101 5350 -5007
rect 5396 -5101 5425 -5007
rect 5321 -5114 5425 -5101
rect 5525 -5007 5613 -4994
rect 5525 -5101 5554 -5007
rect 5600 -5101 5613 -5007
rect 5525 -5114 5613 -5101
rect 5669 -5007 5757 -4994
rect 5669 -5101 5682 -5007
rect 5728 -5101 5757 -5007
rect 5669 -5114 5757 -5101
rect 5857 -5007 5961 -4994
rect 5857 -5101 5886 -5007
rect 5932 -5101 5961 -5007
rect 5857 -5114 5961 -5101
rect 6061 -5007 6149 -4994
rect 6061 -5101 6090 -5007
rect 6136 -5101 6149 -5007
rect 6061 -5114 6149 -5101
rect 3501 -5396 3589 -5383
rect 3501 -5490 3514 -5396
rect 3560 -5490 3589 -5396
rect 3501 -5503 3589 -5490
rect 3689 -5396 3793 -5383
rect 3689 -5490 3718 -5396
rect 3764 -5490 3793 -5396
rect 3689 -5503 3793 -5490
rect 3893 -5396 3997 -5383
rect 3893 -5490 3922 -5396
rect 3968 -5490 3997 -5396
rect 3893 -5503 3997 -5490
rect 4097 -5396 4201 -5383
rect 4097 -5490 4126 -5396
rect 4172 -5490 4201 -5396
rect 4097 -5503 4201 -5490
rect 4301 -5396 4405 -5383
rect 4301 -5490 4330 -5396
rect 4376 -5490 4405 -5396
rect 4301 -5503 4405 -5490
rect 4505 -5396 4609 -5383
rect 4505 -5490 4534 -5396
rect 4580 -5490 4609 -5396
rect 4505 -5503 4609 -5490
rect 4709 -5396 4813 -5383
rect 4709 -5490 4738 -5396
rect 4784 -5490 4813 -5396
rect 4709 -5503 4813 -5490
rect 4913 -5396 5017 -5383
rect 4913 -5490 4942 -5396
rect 4988 -5490 5017 -5396
rect 4913 -5503 5017 -5490
rect 5117 -5396 5221 -5383
rect 5117 -5490 5146 -5396
rect 5192 -5490 5221 -5396
rect 5117 -5503 5221 -5490
rect 5321 -5396 5425 -5383
rect 5321 -5490 5350 -5396
rect 5396 -5490 5425 -5396
rect 5321 -5503 5425 -5490
rect 5525 -5396 5613 -5383
rect 5525 -5490 5554 -5396
rect 5600 -5490 5613 -5396
rect 5525 -5503 5613 -5490
rect 5669 -5396 5757 -5383
rect 5669 -5490 5682 -5396
rect 5728 -5490 5757 -5396
rect 5669 -5503 5757 -5490
rect 5857 -5396 5961 -5383
rect 5857 -5490 5886 -5396
rect 5932 -5490 5961 -5396
rect 5857 -5503 5961 -5490
rect 6061 -5396 6149 -5383
rect 6061 -5490 6090 -5396
rect 6136 -5490 6149 -5396
rect 6061 -5503 6149 -5490
rect 3501 -5691 3589 -5678
rect 3501 -5785 3514 -5691
rect 3560 -5785 3589 -5691
rect 3501 -5798 3589 -5785
rect 3689 -5691 3793 -5678
rect 3689 -5785 3718 -5691
rect 3764 -5785 3793 -5691
rect 3689 -5798 3793 -5785
rect 3893 -5691 3997 -5678
rect 3893 -5785 3922 -5691
rect 3968 -5785 3997 -5691
rect 3893 -5798 3997 -5785
rect 4097 -5691 4201 -5678
rect 4097 -5785 4126 -5691
rect 4172 -5785 4201 -5691
rect 4097 -5798 4201 -5785
rect 4301 -5691 4405 -5678
rect 4301 -5785 4330 -5691
rect 4376 -5785 4405 -5691
rect 4301 -5798 4405 -5785
rect 4505 -5691 4609 -5678
rect 4505 -5785 4534 -5691
rect 4580 -5785 4609 -5691
rect 4505 -5798 4609 -5785
rect 4709 -5691 4813 -5678
rect 4709 -5785 4738 -5691
rect 4784 -5785 4813 -5691
rect 4709 -5798 4813 -5785
rect 4913 -5691 5017 -5678
rect 4913 -5785 4942 -5691
rect 4988 -5785 5017 -5691
rect 4913 -5798 5017 -5785
rect 5117 -5691 5221 -5678
rect 5117 -5785 5146 -5691
rect 5192 -5785 5221 -5691
rect 5117 -5798 5221 -5785
rect 5321 -5691 5425 -5678
rect 5321 -5785 5350 -5691
rect 5396 -5785 5425 -5691
rect 5321 -5798 5425 -5785
rect 5525 -5691 5613 -5678
rect 5525 -5785 5554 -5691
rect 5600 -5785 5613 -5691
rect 5525 -5798 5613 -5785
rect 5669 -5691 5757 -5678
rect 5669 -5785 5682 -5691
rect 5728 -5785 5757 -5691
rect 5669 -5798 5757 -5785
rect 5857 -5691 5961 -5678
rect 5857 -5785 5886 -5691
rect 5932 -5785 5961 -5691
rect 5857 -5798 5961 -5785
rect 6061 -5691 6149 -5678
rect 6061 -5785 6090 -5691
rect 6136 -5785 6149 -5691
rect 6061 -5798 6149 -5785
rect -2062 -6006 -1990 -5995
rect -1894 -6006 -1822 -5995
rect -2062 -6008 -1970 -6006
rect -2062 -6054 -2049 -6008
rect -2003 -6054 -1970 -6008
rect -2062 -6056 -1970 -6054
rect -1914 -6008 -1822 -6006
rect -1914 -6054 -1881 -6008
rect -1835 -6054 -1822 -6008
rect -1584 -6010 -1512 -5997
rect -1914 -6056 -1822 -6054
rect -2062 -6067 -1990 -6056
rect -1894 -6067 -1822 -6056
rect -1584 -6056 -1571 -6010
rect -1525 -6011 -1512 -6010
rect -1416 -6010 -1344 -5997
rect -1416 -6011 -1403 -6010
rect -1525 -6055 -1492 -6011
rect -1436 -6055 -1403 -6011
rect -1525 -6056 -1512 -6055
rect -1584 -6069 -1512 -6056
rect -1416 -6056 -1403 -6055
rect -1357 -6056 -1344 -6010
rect -1416 -6069 -1344 -6056
rect -1048 -6010 -976 -5997
rect -1048 -6056 -1035 -6010
rect -989 -6011 -976 -6010
rect -880 -6010 -808 -5997
rect -880 -6011 -867 -6010
rect -989 -6055 -956 -6011
rect -900 -6055 -867 -6011
rect -989 -6056 -976 -6055
rect -1048 -6069 -976 -6056
rect -880 -6056 -867 -6055
rect -821 -6056 -808 -6010
rect -880 -6069 -808 -6056
rect -444 -6006 -372 -5995
rect -276 -6006 -204 -5995
rect -444 -6008 -352 -6006
rect -444 -6054 -431 -6008
rect -385 -6054 -352 -6008
rect -444 -6056 -352 -6054
rect -296 -6008 -204 -6006
rect -296 -6054 -263 -6008
rect -217 -6054 -204 -6008
rect 34 -6010 106 -5997
rect -296 -6056 -204 -6054
rect -444 -6067 -372 -6056
rect -276 -6067 -204 -6056
rect 34 -6056 47 -6010
rect 93 -6011 106 -6010
rect 202 -6010 274 -5997
rect 202 -6011 215 -6010
rect 93 -6055 126 -6011
rect 182 -6055 215 -6011
rect 93 -6056 106 -6055
rect 34 -6069 106 -6056
rect 202 -6056 215 -6055
rect 261 -6056 274 -6010
rect 202 -6069 274 -6056
rect 570 -6010 642 -5997
rect 570 -6056 583 -6010
rect 629 -6011 642 -6010
rect 738 -6010 810 -5997
rect 738 -6011 751 -6010
rect 629 -6055 662 -6011
rect 718 -6055 751 -6011
rect 629 -6056 642 -6055
rect 570 -6069 642 -6056
rect 738 -6056 751 -6055
rect 797 -6056 810 -6010
rect 738 -6069 810 -6056
rect 1165 -6006 1237 -5995
rect 1333 -6006 1405 -5995
rect 1165 -6008 1257 -6006
rect 1165 -6054 1178 -6008
rect 1224 -6054 1257 -6008
rect 1165 -6056 1257 -6054
rect 1313 -6008 1405 -6006
rect 1313 -6054 1346 -6008
rect 1392 -6054 1405 -6008
rect 1643 -6010 1715 -5997
rect 1313 -6056 1405 -6054
rect 1165 -6067 1237 -6056
rect 1333 -6067 1405 -6056
rect 1643 -6056 1656 -6010
rect 1702 -6011 1715 -6010
rect 1811 -6010 1883 -5997
rect 1811 -6011 1824 -6010
rect 1702 -6055 1735 -6011
rect 1791 -6055 1824 -6011
rect 1702 -6056 1715 -6055
rect 1643 -6069 1715 -6056
rect 1811 -6056 1824 -6055
rect 1870 -6056 1883 -6010
rect 1811 -6069 1883 -6056
rect 2179 -6010 2251 -5997
rect 2179 -6056 2192 -6010
rect 2238 -6011 2251 -6010
rect 2347 -6010 2419 -5997
rect 2347 -6011 2360 -6010
rect 2238 -6055 2271 -6011
rect 2327 -6055 2360 -6011
rect 2238 -6056 2251 -6055
rect 2179 -6069 2251 -6056
rect 2347 -6056 2360 -6055
rect 2406 -6056 2419 -6010
rect 2347 -6069 2419 -6056
rect 3501 -6076 3589 -6063
rect 3501 -6170 3514 -6076
rect 3560 -6170 3589 -6076
rect 3501 -6183 3589 -6170
rect 3689 -6076 3793 -6063
rect 3689 -6170 3718 -6076
rect 3764 -6170 3793 -6076
rect 3689 -6183 3793 -6170
rect 3893 -6076 3997 -6063
rect 3893 -6170 3922 -6076
rect 3968 -6170 3997 -6076
rect 3893 -6183 3997 -6170
rect 4097 -6076 4201 -6063
rect 4097 -6170 4126 -6076
rect 4172 -6170 4201 -6076
rect 4097 -6183 4201 -6170
rect 4301 -6076 4405 -6063
rect 4301 -6170 4330 -6076
rect 4376 -6170 4405 -6076
rect 4301 -6183 4405 -6170
rect 4505 -6076 4609 -6063
rect 4505 -6170 4534 -6076
rect 4580 -6170 4609 -6076
rect 4505 -6183 4609 -6170
rect 4709 -6076 4813 -6063
rect 4709 -6170 4738 -6076
rect 4784 -6170 4813 -6076
rect 4709 -6183 4813 -6170
rect 4913 -6076 5017 -6063
rect 4913 -6170 4942 -6076
rect 4988 -6170 5017 -6076
rect 4913 -6183 5017 -6170
rect 5117 -6076 5221 -6063
rect 5117 -6170 5146 -6076
rect 5192 -6170 5221 -6076
rect 5117 -6183 5221 -6170
rect 5321 -6076 5425 -6063
rect 5321 -6170 5350 -6076
rect 5396 -6170 5425 -6076
rect 5321 -6183 5425 -6170
rect 5525 -6076 5613 -6063
rect 5525 -6170 5554 -6076
rect 5600 -6170 5613 -6076
rect 5525 -6183 5613 -6170
rect 5669 -6076 5757 -6063
rect 5669 -6170 5682 -6076
rect 5728 -6170 5757 -6076
rect 5669 -6183 5757 -6170
rect 5857 -6076 5961 -6063
rect 5857 -6170 5886 -6076
rect 5932 -6170 5961 -6076
rect 5857 -6183 5961 -6170
rect 6061 -6076 6149 -6063
rect 6061 -6170 6090 -6076
rect 6136 -6170 6149 -6076
rect 6061 -6183 6149 -6170
<< pdiff >>
rect -2058 -3075 -1970 -3062
rect -2058 -3149 -2045 -3075
rect -1999 -3149 -1970 -3075
rect -2058 -3162 -1970 -3149
rect -1914 -3075 -1826 -3062
rect -1914 -3149 -1885 -3075
rect -1839 -3149 -1826 -3075
rect -1914 -3162 -1826 -3149
rect -1522 -3110 -1450 -3097
rect -1522 -3156 -1509 -3110
rect -1463 -3111 -1450 -3110
rect -1354 -3110 -1282 -3097
rect -1354 -3111 -1341 -3110
rect -1463 -3155 -1430 -3111
rect -1374 -3155 -1341 -3111
rect -1463 -3156 -1450 -3155
rect -1522 -3169 -1450 -3156
rect -1354 -3156 -1341 -3155
rect -1295 -3156 -1282 -3110
rect -1354 -3169 -1282 -3156
rect -1110 -3110 -1038 -3097
rect -1110 -3156 -1097 -3110
rect -1051 -3111 -1038 -3110
rect -942 -3110 -870 -3097
rect -942 -3111 -929 -3110
rect -1051 -3155 -1018 -3111
rect -962 -3155 -929 -3111
rect -1051 -3156 -1038 -3155
rect -1110 -3169 -1038 -3156
rect -942 -3156 -929 -3155
rect -883 -3156 -870 -3110
rect -942 -3169 -870 -3156
rect -2058 -3943 -1970 -3930
rect -2058 -4017 -2045 -3943
rect -1999 -4017 -1970 -3943
rect -2058 -4030 -1970 -4017
rect -1914 -3943 -1826 -3930
rect -1914 -4017 -1885 -3943
rect -1839 -4017 -1826 -3943
rect -1914 -4030 -1826 -4017
rect -1522 -3978 -1450 -3965
rect -1522 -4024 -1509 -3978
rect -1463 -3979 -1450 -3978
rect -1354 -3978 -1282 -3965
rect -1354 -3979 -1341 -3978
rect -1463 -4023 -1430 -3979
rect -1374 -4023 -1341 -3979
rect -1463 -4024 -1450 -4023
rect -1522 -4037 -1450 -4024
rect -1354 -4024 -1341 -4023
rect -1295 -4024 -1282 -3978
rect -1354 -4037 -1282 -4024
rect -1110 -3978 -1038 -3965
rect -1110 -4024 -1097 -3978
rect -1051 -3979 -1038 -3978
rect -942 -3978 -870 -3965
rect -942 -3979 -929 -3978
rect -1051 -4023 -1018 -3979
rect -962 -4023 -929 -3979
rect -1051 -4024 -1038 -4023
rect -1110 -4037 -1038 -4024
rect -942 -4024 -929 -4023
rect -883 -4024 -870 -3978
rect -942 -4037 -870 -4024
rect -2058 -4802 -1970 -4789
rect -2058 -4876 -2045 -4802
rect -1999 -4876 -1970 -4802
rect -2058 -4889 -1970 -4876
rect -1914 -4802 -1826 -4789
rect -1914 -4876 -1885 -4802
rect -1839 -4876 -1826 -4802
rect -1914 -4889 -1826 -4876
rect -1522 -4837 -1450 -4824
rect -1522 -4883 -1509 -4837
rect -1463 -4838 -1450 -4837
rect -1354 -4837 -1282 -4824
rect -1354 -4838 -1341 -4837
rect -1463 -4882 -1430 -4838
rect -1374 -4882 -1341 -4838
rect -1463 -4883 -1450 -4882
rect -1522 -4896 -1450 -4883
rect -1354 -4883 -1341 -4882
rect -1295 -4883 -1282 -4837
rect -1354 -4896 -1282 -4883
rect -1110 -4837 -1038 -4824
rect -1110 -4883 -1097 -4837
rect -1051 -4838 -1038 -4837
rect -942 -4837 -870 -4824
rect -942 -4838 -929 -4837
rect -1051 -4882 -1018 -4838
rect -962 -4882 -929 -4838
rect -1051 -4883 -1038 -4882
rect -1110 -4896 -1038 -4883
rect -942 -4883 -929 -4882
rect -883 -4883 -870 -4837
rect -942 -4896 -870 -4883
rect -2058 -5670 -1970 -5657
rect -2058 -5744 -2045 -5670
rect -1999 -5744 -1970 -5670
rect -2058 -5757 -1970 -5744
rect -1914 -5670 -1826 -5657
rect -1914 -5744 -1885 -5670
rect -1839 -5744 -1826 -5670
rect -1914 -5757 -1826 -5744
rect -1522 -5705 -1450 -5692
rect -1522 -5751 -1509 -5705
rect -1463 -5706 -1450 -5705
rect -1354 -5705 -1282 -5692
rect -1354 -5706 -1341 -5705
rect -1463 -5750 -1430 -5706
rect -1374 -5750 -1341 -5706
rect -1463 -5751 -1450 -5750
rect -1522 -5764 -1450 -5751
rect -1354 -5751 -1341 -5750
rect -1295 -5751 -1282 -5705
rect -1354 -5764 -1282 -5751
rect -1110 -5705 -1038 -5692
rect -1110 -5751 -1097 -5705
rect -1051 -5706 -1038 -5705
rect -440 -5670 -352 -5657
rect -942 -5705 -870 -5692
rect -942 -5706 -929 -5705
rect -1051 -5750 -1018 -5706
rect -962 -5750 -929 -5706
rect -1051 -5751 -1038 -5750
rect -1110 -5764 -1038 -5751
rect -942 -5751 -929 -5750
rect -883 -5751 -870 -5705
rect -942 -5764 -870 -5751
rect -440 -5744 -427 -5670
rect -381 -5744 -352 -5670
rect -440 -5757 -352 -5744
rect -296 -5670 -208 -5657
rect -296 -5744 -267 -5670
rect -221 -5744 -208 -5670
rect -296 -5757 -208 -5744
rect 96 -5705 168 -5692
rect 96 -5751 109 -5705
rect 155 -5706 168 -5705
rect 264 -5705 336 -5692
rect 264 -5706 277 -5705
rect 155 -5750 188 -5706
rect 244 -5750 277 -5706
rect 155 -5751 168 -5750
rect 96 -5764 168 -5751
rect 264 -5751 277 -5750
rect 323 -5751 336 -5705
rect 264 -5764 336 -5751
rect 508 -5705 580 -5692
rect 508 -5751 521 -5705
rect 567 -5706 580 -5705
rect 1169 -5670 1257 -5657
rect 676 -5705 748 -5692
rect 676 -5706 689 -5705
rect 567 -5750 600 -5706
rect 656 -5750 689 -5706
rect 567 -5751 580 -5750
rect 508 -5764 580 -5751
rect 676 -5751 689 -5750
rect 735 -5751 748 -5705
rect 676 -5764 748 -5751
rect 1169 -5744 1182 -5670
rect 1228 -5744 1257 -5670
rect 1169 -5757 1257 -5744
rect 1313 -5670 1401 -5657
rect 1313 -5744 1342 -5670
rect 1388 -5744 1401 -5670
rect 1313 -5757 1401 -5744
rect 1705 -5705 1777 -5692
rect 1705 -5751 1718 -5705
rect 1764 -5706 1777 -5705
rect 1873 -5705 1945 -5692
rect 1873 -5706 1886 -5705
rect 1764 -5750 1797 -5706
rect 1853 -5750 1886 -5706
rect 1764 -5751 1777 -5750
rect 1705 -5764 1777 -5751
rect 1873 -5751 1886 -5750
rect 1932 -5751 1945 -5705
rect 1873 -5764 1945 -5751
rect 2117 -5705 2189 -5692
rect 2117 -5751 2130 -5705
rect 2176 -5706 2189 -5705
rect 2285 -5705 2357 -5692
rect 2285 -5706 2298 -5705
rect 2176 -5750 2209 -5706
rect 2265 -5750 2298 -5706
rect 2176 -5751 2189 -5750
rect 2117 -5764 2189 -5751
rect 2285 -5751 2298 -5750
rect 2344 -5751 2357 -5705
rect 2285 -5764 2357 -5751
<< ndiffc >>
rect -1759 1499 -1713 1593
rect -1555 1499 -1509 1593
rect -1372 1499 -1326 1593
rect -1168 1499 -1122 1593
rect -964 1499 -918 1593
rect -760 1499 -714 1593
rect -556 1499 -510 1593
rect -352 1499 -306 1593
rect -148 1499 -102 1593
rect 56 1499 102 1593
rect 260 1499 306 1593
rect 464 1499 510 1593
rect 668 1499 714 1593
rect 872 1499 918 1593
rect 1076 1499 1122 1593
rect 1280 1499 1326 1593
rect 1484 1499 1530 1593
rect 1688 1499 1734 1593
rect 1892 1499 1938 1593
rect 2069 1499 2115 1593
rect 2273 1499 2319 1593
rect 3041 1511 3087 1557
rect 3253 1511 3299 1557
rect 3381 1511 3427 1557
rect 3593 1511 3639 1557
rect 3721 1511 3767 1557
rect 3933 1511 3979 1557
rect 4145 1511 4191 1557
rect 4357 1511 4403 1557
rect -1759 1196 -1713 1290
rect -1555 1196 -1509 1290
rect -1372 1196 -1326 1290
rect -1168 1196 -1122 1290
rect -964 1196 -918 1290
rect -760 1196 -714 1290
rect -556 1196 -510 1290
rect -352 1196 -306 1290
rect -148 1196 -102 1290
rect 56 1196 102 1290
rect 260 1196 306 1290
rect 464 1196 510 1290
rect 668 1196 714 1290
rect 872 1196 918 1290
rect 1076 1196 1122 1290
rect 1280 1196 1326 1290
rect 1484 1196 1530 1290
rect 1688 1196 1734 1290
rect 1892 1196 1938 1290
rect 2069 1196 2115 1290
rect 2273 1196 2319 1290
rect 4716 1445 4762 1491
rect 4928 1445 4974 1491
rect 5140 1445 5186 1491
rect 3049 1197 3095 1291
rect 3253 1197 3299 1291
rect 3381 1197 3427 1291
rect 3585 1197 3631 1291
rect 3789 1197 3835 1291
rect 3993 1197 4039 1291
rect 4197 1197 4243 1291
rect 4401 1197 4447 1291
rect 5268 1445 5314 1491
rect 5480 1445 5526 1491
rect 5692 1445 5738 1491
rect 4716 1203 4762 1249
rect 4928 1203 4974 1249
rect 5140 1203 5186 1249
rect 5820 1445 5866 1491
rect 6032 1445 6078 1491
rect 5268 1203 5314 1249
rect 5480 1203 5526 1249
rect 5692 1203 5738 1249
rect 3041 883 3087 929
rect 3253 883 3299 929
rect -1759 757 -1713 851
rect -1555 757 -1509 851
rect -1372 757 -1326 851
rect -1168 757 -1122 851
rect -964 757 -918 851
rect -760 757 -714 851
rect -556 757 -510 851
rect -352 757 -306 851
rect -148 757 -102 851
rect 56 757 102 851
rect 260 757 306 851
rect 464 757 510 851
rect 668 757 714 851
rect 872 757 918 851
rect 1076 757 1122 851
rect 1280 757 1326 851
rect 1484 757 1530 851
rect 1688 757 1734 851
rect 1892 757 1938 851
rect 2069 757 2115 851
rect 2273 757 2319 851
rect 3381 883 3427 929
rect 3593 883 3639 929
rect 3721 883 3767 929
rect 3933 883 3979 929
rect 4145 883 4191 929
rect 5820 1203 5866 1249
rect 6032 1203 6078 1249
rect 4273 883 4319 929
rect 4485 883 4531 929
rect 4862 871 4908 965
rect 5066 871 5112 965
rect 5270 871 5316 965
rect 5474 871 5520 965
rect 5678 871 5724 965
rect 5882 871 5928 965
rect 3123 551 3169 645
rect 3327 551 3373 645
rect 3531 551 3577 645
rect 3735 551 3781 645
rect 3939 551 3985 645
rect 4143 551 4189 645
rect 4347 551 4393 645
rect 4551 551 4597 645
rect 4862 569 4908 663
rect 5066 569 5112 663
rect 5270 569 5316 663
rect 5474 569 5520 663
rect 5678 569 5724 663
rect 5882 569 5928 663
rect -1759 81 -1713 175
rect -1555 81 -1509 175
rect -1351 81 -1305 175
rect -1147 81 -1101 175
rect -943 81 -897 175
rect -815 81 -769 175
rect -611 81 -565 175
rect -407 81 -361 175
rect -279 81 -233 175
rect -75 81 -29 175
rect 53 81 99 175
rect 257 81 303 175
rect 461 81 507 175
rect 589 81 635 175
rect 793 81 839 175
rect 921 81 967 175
rect 1125 81 1171 175
rect 1329 81 1375 175
rect 1457 81 1503 175
rect 1661 81 1707 175
rect 1865 81 1911 175
rect 2069 81 2115 175
rect 2273 81 2319 175
rect 2963 27 3009 121
rect 3167 27 3213 121
rect 3371 27 3417 121
rect 3575 27 3621 121
rect 3779 27 3825 121
rect 3983 27 4029 121
rect 4187 27 4233 121
rect 4430 45 4476 91
rect 4642 45 4688 91
rect -1759 -245 -1713 -151
rect -1555 -245 -1509 -151
rect -1351 -245 -1305 -151
rect -1147 -245 -1101 -151
rect -943 -245 -897 -151
rect -815 -245 -769 -151
rect -611 -245 -565 -151
rect -407 -245 -361 -151
rect -279 -245 -233 -151
rect -75 -245 -29 -151
rect 53 -245 99 -151
rect 257 -245 303 -151
rect 461 -245 507 -151
rect 589 -245 635 -151
rect 793 -245 839 -151
rect 921 -245 967 -151
rect 1125 -245 1171 -151
rect 1329 -245 1375 -151
rect 1457 -245 1503 -151
rect 1661 -245 1707 -151
rect 1865 -245 1911 -151
rect 2069 -245 2115 -151
rect 2273 -245 2319 -151
rect 4770 45 4816 91
rect 4982 45 5028 91
rect 5194 45 5240 91
rect 5322 45 5368 91
rect 5534 45 5580 91
rect 5746 45 5792 91
rect 2963 -351 3009 -257
rect 3167 -351 3213 -257
rect 3371 -351 3417 -257
rect 3575 -351 3621 -257
rect 3779 -351 3825 -257
rect 3983 -351 4029 -257
rect 4187 -351 4233 -257
rect 4429 -271 4475 -225
rect 4641 -271 4687 -225
rect 4769 -271 4815 -225
rect 4981 -271 5027 -225
rect 5193 -271 5239 -225
rect 5321 -271 5367 -225
rect 5533 -271 5579 -225
rect 5745 -271 5791 -225
rect 4429 -521 4475 -475
rect 2963 -630 3009 -536
rect 3167 -630 3213 -536
rect 3371 -630 3417 -536
rect 3575 -630 3621 -536
rect 3779 -630 3825 -536
rect 3983 -630 4029 -536
rect 4641 -521 4687 -475
rect 4187 -630 4233 -536
rect 4769 -521 4815 -475
rect 4981 -521 5027 -475
rect 5193 -521 5239 -475
rect 5321 -521 5367 -475
rect 5533 -521 5579 -475
rect 5745 -521 5791 -475
rect -1759 -1037 -1713 -943
rect -1555 -1037 -1509 -943
rect -1372 -1037 -1326 -943
rect -1168 -1037 -1122 -943
rect -964 -1037 -918 -943
rect -760 -1037 -714 -943
rect -556 -1037 -510 -943
rect -352 -1037 -306 -943
rect -148 -1037 -102 -943
rect 56 -1037 102 -943
rect 260 -1037 306 -943
rect 464 -1037 510 -943
rect 668 -1037 714 -943
rect 872 -1037 918 -943
rect 1076 -1037 1122 -943
rect 1280 -1037 1326 -943
rect 1484 -1037 1530 -943
rect 1688 -1037 1734 -943
rect 1892 -1037 1938 -943
rect 2069 -1037 2115 -943
rect 2273 -1037 2319 -943
rect 4429 -846 4475 -800
rect 4641 -846 4687 -800
rect 2963 -1008 3009 -914
rect 3167 -1008 3213 -914
rect 3371 -1008 3417 -914
rect 3575 -1008 3621 -914
rect 3779 -1008 3825 -914
rect 3983 -1008 4029 -914
rect 4187 -1008 4233 -914
rect 4769 -846 4815 -800
rect 4981 -846 5027 -800
rect 5193 -846 5239 -800
rect 5321 -846 5367 -800
rect 5533 -846 5579 -800
rect 5745 -846 5791 -800
rect -1759 -1468 -1713 -1374
rect -1555 -1468 -1509 -1374
rect -1372 -1468 -1326 -1374
rect -1168 -1468 -1122 -1374
rect -964 -1468 -918 -1374
rect -760 -1468 -714 -1374
rect -556 -1468 -510 -1374
rect -352 -1468 -306 -1374
rect -148 -1468 -102 -1374
rect 56 -1468 102 -1374
rect 260 -1468 306 -1374
rect 464 -1468 510 -1374
rect 668 -1468 714 -1374
rect 872 -1468 918 -1374
rect 1076 -1468 1122 -1374
rect 1280 -1468 1326 -1374
rect 1484 -1468 1530 -1374
rect 1688 -1468 1734 -1374
rect 1892 -1468 1938 -1374
rect 2069 -1468 2115 -1374
rect 2273 -1468 2319 -1374
rect -1759 -1778 -1713 -1684
rect -1555 -1778 -1509 -1684
rect -1372 -1778 -1326 -1684
rect -1168 -1778 -1122 -1684
rect -964 -1778 -918 -1684
rect -760 -1778 -714 -1684
rect -556 -1778 -510 -1684
rect -352 -1778 -306 -1684
rect -148 -1778 -102 -1684
rect 56 -1778 102 -1684
rect 260 -1778 306 -1684
rect 464 -1778 510 -1684
rect 668 -1778 714 -1684
rect 872 -1778 918 -1684
rect 1076 -1778 1122 -1684
rect 1280 -1778 1326 -1684
rect 1484 -1778 1530 -1684
rect 1688 -1778 1734 -1684
rect 1892 -1778 1938 -1684
rect 2069 -1778 2115 -1684
rect 2273 -1778 2319 -1684
rect 3514 -2013 3560 -1919
rect 3718 -2013 3764 -1919
rect 3922 -2013 3968 -1919
rect 4050 -2013 4096 -1919
rect 4254 -2013 4300 -1919
rect 4458 -2013 4504 -1919
rect 4586 -2013 4632 -1919
rect 4790 -2013 4836 -1919
rect 4994 -2013 5040 -1919
rect 5122 -2013 5168 -1919
rect 5326 -2013 5372 -1919
rect 5530 -2013 5576 -1919
rect 5658 -2013 5704 -1919
rect 5862 -2013 5908 -1919
rect 6066 -2013 6112 -1919
rect 3514 -2397 3560 -2303
rect 3718 -2397 3764 -2303
rect 3922 -2397 3968 -2303
rect 4050 -2397 4096 -2303
rect 4254 -2397 4300 -2303
rect 4458 -2397 4504 -2303
rect 4586 -2397 4632 -2303
rect 4790 -2397 4836 -2303
rect 4994 -2397 5040 -2303
rect 5122 -2397 5168 -2303
rect 5326 -2397 5372 -2303
rect 5530 -2397 5576 -2303
rect 5658 -2397 5704 -2303
rect 5862 -2397 5908 -2303
rect 6066 -2397 6112 -2303
rect -54 -2996 -8 -2902
rect 150 -2996 196 -2902
rect 354 -2996 400 -2902
rect 482 -2996 528 -2902
rect 686 -2996 732 -2902
rect 890 -2996 936 -2902
rect 1018 -2996 1064 -2902
rect 1222 -2996 1268 -2902
rect 1426 -2996 1472 -2902
rect 1554 -2996 1600 -2902
rect 1758 -2996 1804 -2902
rect 1962 -2996 2008 -2902
rect 2090 -2996 2136 -2902
rect 2294 -2996 2340 -2902
rect 2498 -2996 2544 -2902
rect -54 -3280 -8 -3186
rect 150 -3280 196 -3186
rect 354 -3280 400 -3186
rect 482 -3280 528 -3186
rect 686 -3280 732 -3186
rect 890 -3280 936 -3186
rect 1018 -3280 1064 -3186
rect 1222 -3280 1268 -3186
rect 1426 -3280 1472 -3186
rect 1554 -3280 1600 -3186
rect 1758 -3280 1804 -3186
rect 1962 -3280 2008 -3186
rect 2090 -3280 2136 -3186
rect 2294 -3280 2340 -3186
rect 2498 -3280 2544 -3186
rect -2049 -3459 -2003 -3413
rect -1881 -3459 -1835 -3413
rect -1571 -3461 -1525 -3415
rect -1403 -3461 -1357 -3415
rect -1035 -3461 -989 -3415
rect -867 -3461 -821 -3415
rect -54 -3812 -8 -3718
rect 150 -3812 196 -3718
rect 354 -3812 400 -3718
rect 558 -3812 604 -3718
rect 762 -3812 808 -3718
rect 966 -3812 1012 -3718
rect 1170 -3812 1216 -3718
rect 1374 -3812 1420 -3718
rect 1578 -3812 1624 -3718
rect 1782 -3812 1828 -3718
rect 1986 -3812 2032 -3718
rect 2114 -3812 2160 -3718
rect 2318 -3812 2364 -3718
rect 2522 -3812 2568 -3718
rect -2049 -4327 -2003 -4281
rect -1881 -4327 -1835 -4281
rect -1571 -4329 -1525 -4283
rect -1403 -4329 -1357 -4283
rect -1035 -4329 -989 -4283
rect -54 -4201 -8 -4107
rect 150 -4201 196 -4107
rect 354 -4201 400 -4107
rect 558 -4201 604 -4107
rect 762 -4201 808 -4107
rect 966 -4201 1012 -4107
rect 1170 -4201 1216 -4107
rect 1374 -4201 1420 -4107
rect 1578 -4201 1624 -4107
rect 1782 -4201 1828 -4107
rect 1986 -4201 2032 -4107
rect 2114 -4201 2160 -4107
rect 2318 -4201 2364 -4107
rect 2522 -4201 2568 -4107
rect -867 -4329 -821 -4283
rect -54 -4496 -8 -4402
rect 150 -4496 196 -4402
rect 354 -4496 400 -4402
rect 558 -4496 604 -4402
rect 762 -4496 808 -4402
rect 966 -4496 1012 -4402
rect 1170 -4496 1216 -4402
rect 1374 -4496 1420 -4402
rect 1578 -4496 1624 -4402
rect 1782 -4496 1828 -4402
rect 1986 -4496 2032 -4402
rect 2114 -4496 2160 -4402
rect 2318 -4496 2364 -4402
rect 2522 -4496 2568 -4402
rect -54 -4881 -8 -4787
rect 150 -4881 196 -4787
rect 354 -4881 400 -4787
rect 558 -4881 604 -4787
rect 762 -4881 808 -4787
rect 966 -4881 1012 -4787
rect 1170 -4881 1216 -4787
rect 1374 -4881 1420 -4787
rect 1578 -4881 1624 -4787
rect 1782 -4881 1828 -4787
rect 1986 -4881 2032 -4787
rect 2114 -4881 2160 -4787
rect 2318 -4881 2364 -4787
rect 2522 -4881 2568 -4787
rect -2049 -5186 -2003 -5140
rect -1881 -5186 -1835 -5140
rect -1571 -5188 -1525 -5142
rect -1403 -5188 -1357 -5142
rect -1035 -5188 -989 -5142
rect -867 -5188 -821 -5142
rect 3514 -2687 3560 -2593
rect 3718 -2687 3764 -2593
rect 3922 -2687 3968 -2593
rect 4050 -2687 4096 -2593
rect 4254 -2687 4300 -2593
rect 4458 -2687 4504 -2593
rect 4586 -2687 4632 -2593
rect 4790 -2687 4836 -2593
rect 4994 -2687 5040 -2593
rect 5122 -2687 5168 -2593
rect 5326 -2687 5372 -2593
rect 5530 -2687 5576 -2593
rect 5658 -2687 5704 -2593
rect 5862 -2687 5908 -2593
rect 6066 -2687 6112 -2593
rect 3514 -3071 3560 -2977
rect 3718 -3071 3764 -2977
rect 3922 -3071 3968 -2977
rect 4050 -3071 4096 -2977
rect 4254 -3071 4300 -2977
rect 4458 -3071 4504 -2977
rect 4586 -3071 4632 -2977
rect 4790 -3071 4836 -2977
rect 4994 -3071 5040 -2977
rect 5122 -3071 5168 -2977
rect 5326 -3071 5372 -2977
rect 5530 -3071 5576 -2977
rect 5658 -3071 5704 -2977
rect 5862 -3071 5908 -2977
rect 6066 -3071 6112 -2977
rect 3514 -3705 3560 -3611
rect 3718 -3705 3764 -3611
rect 3922 -3705 3968 -3611
rect 4126 -3705 4172 -3611
rect 4330 -3705 4376 -3611
rect 4534 -3705 4580 -3611
rect 4738 -3705 4784 -3611
rect 4942 -3705 4988 -3611
rect 5146 -3705 5192 -3611
rect 5350 -3705 5396 -3611
rect 5554 -3705 5600 -3611
rect 5682 -3705 5728 -3611
rect 5886 -3705 5932 -3611
rect 6090 -3705 6136 -3611
rect 3514 -4094 3560 -4000
rect 3718 -4094 3764 -4000
rect 3922 -4094 3968 -4000
rect 4126 -4094 4172 -4000
rect 4330 -4094 4376 -4000
rect 4534 -4094 4580 -4000
rect 4738 -4094 4784 -4000
rect 4942 -4094 4988 -4000
rect 5146 -4094 5192 -4000
rect 5350 -4094 5396 -4000
rect 5554 -4094 5600 -4000
rect 5682 -4094 5728 -4000
rect 5886 -4094 5932 -4000
rect 6090 -4094 6136 -4000
rect 3514 -4389 3560 -4295
rect 3718 -4389 3764 -4295
rect 3922 -4389 3968 -4295
rect 4126 -4389 4172 -4295
rect 4330 -4389 4376 -4295
rect 4534 -4389 4580 -4295
rect 4738 -4389 4784 -4295
rect 4942 -4389 4988 -4295
rect 5146 -4389 5192 -4295
rect 5350 -4389 5396 -4295
rect 5554 -4389 5600 -4295
rect 5682 -4389 5728 -4295
rect 5886 -4389 5932 -4295
rect 6090 -4389 6136 -4295
rect 3514 -4774 3560 -4680
rect 3718 -4774 3764 -4680
rect 3922 -4774 3968 -4680
rect 4126 -4774 4172 -4680
rect 4330 -4774 4376 -4680
rect 4534 -4774 4580 -4680
rect 4738 -4774 4784 -4680
rect 4942 -4774 4988 -4680
rect 5146 -4774 5192 -4680
rect 5350 -4774 5396 -4680
rect 5554 -4774 5600 -4680
rect 5682 -4774 5728 -4680
rect 5886 -4774 5932 -4680
rect 6090 -4774 6136 -4680
rect 3514 -5101 3560 -5007
rect 3718 -5101 3764 -5007
rect 3922 -5101 3968 -5007
rect 4126 -5101 4172 -5007
rect 4330 -5101 4376 -5007
rect 4534 -5101 4580 -5007
rect 4738 -5101 4784 -5007
rect 4942 -5101 4988 -5007
rect 5146 -5101 5192 -5007
rect 5350 -5101 5396 -5007
rect 5554 -5101 5600 -5007
rect 5682 -5101 5728 -5007
rect 5886 -5101 5932 -5007
rect 6090 -5101 6136 -5007
rect 3514 -5490 3560 -5396
rect 3718 -5490 3764 -5396
rect 3922 -5490 3968 -5396
rect 4126 -5490 4172 -5396
rect 4330 -5490 4376 -5396
rect 4534 -5490 4580 -5396
rect 4738 -5490 4784 -5396
rect 4942 -5490 4988 -5396
rect 5146 -5490 5192 -5396
rect 5350 -5490 5396 -5396
rect 5554 -5490 5600 -5396
rect 5682 -5490 5728 -5396
rect 5886 -5490 5932 -5396
rect 6090 -5490 6136 -5396
rect 3514 -5785 3560 -5691
rect 3718 -5785 3764 -5691
rect 3922 -5785 3968 -5691
rect 4126 -5785 4172 -5691
rect 4330 -5785 4376 -5691
rect 4534 -5785 4580 -5691
rect 4738 -5785 4784 -5691
rect 4942 -5785 4988 -5691
rect 5146 -5785 5192 -5691
rect 5350 -5785 5396 -5691
rect 5554 -5785 5600 -5691
rect 5682 -5785 5728 -5691
rect 5886 -5785 5932 -5691
rect 6090 -5785 6136 -5691
rect -2049 -6054 -2003 -6008
rect -1881 -6054 -1835 -6008
rect -1571 -6056 -1525 -6010
rect -1403 -6056 -1357 -6010
rect -1035 -6056 -989 -6010
rect -867 -6056 -821 -6010
rect -431 -6054 -385 -6008
rect -263 -6054 -217 -6008
rect 47 -6056 93 -6010
rect 215 -6056 261 -6010
rect 583 -6056 629 -6010
rect 751 -6056 797 -6010
rect 1178 -6054 1224 -6008
rect 1346 -6054 1392 -6008
rect 1656 -6056 1702 -6010
rect 1824 -6056 1870 -6010
rect 2192 -6056 2238 -6010
rect 2360 -6056 2406 -6010
rect 3514 -6170 3560 -6076
rect 3718 -6170 3764 -6076
rect 3922 -6170 3968 -6076
rect 4126 -6170 4172 -6076
rect 4330 -6170 4376 -6076
rect 4534 -6170 4580 -6076
rect 4738 -6170 4784 -6076
rect 4942 -6170 4988 -6076
rect 5146 -6170 5192 -6076
rect 5350 -6170 5396 -6076
rect 5554 -6170 5600 -6076
rect 5682 -6170 5728 -6076
rect 5886 -6170 5932 -6076
rect 6090 -6170 6136 -6076
<< pdiffc >>
rect -2045 -3149 -1999 -3075
rect -1885 -3149 -1839 -3075
rect -1509 -3156 -1463 -3110
rect -1341 -3156 -1295 -3110
rect -1097 -3156 -1051 -3110
rect -929 -3156 -883 -3110
rect -2045 -4017 -1999 -3943
rect -1885 -4017 -1839 -3943
rect -1509 -4024 -1463 -3978
rect -1341 -4024 -1295 -3978
rect -1097 -4024 -1051 -3978
rect -929 -4024 -883 -3978
rect -2045 -4876 -1999 -4802
rect -1885 -4876 -1839 -4802
rect -1509 -4883 -1463 -4837
rect -1341 -4883 -1295 -4837
rect -1097 -4883 -1051 -4837
rect -929 -4883 -883 -4837
rect -2045 -5744 -1999 -5670
rect -1885 -5744 -1839 -5670
rect -1509 -5751 -1463 -5705
rect -1341 -5751 -1295 -5705
rect -1097 -5751 -1051 -5705
rect -929 -5751 -883 -5705
rect -427 -5744 -381 -5670
rect -267 -5744 -221 -5670
rect 109 -5751 155 -5705
rect 277 -5751 323 -5705
rect 521 -5751 567 -5705
rect 689 -5751 735 -5705
rect 1182 -5744 1228 -5670
rect 1342 -5744 1388 -5670
rect 1718 -5751 1764 -5705
rect 1886 -5751 1932 -5705
rect 2130 -5751 2176 -5705
rect 2298 -5751 2344 -5705
<< psubdiff >>
rect -1235 2008 1843 2027
rect -1235 1938 -1191 2008
rect 1787 1938 1843 2008
rect -1235 1916 1843 1938
rect 2665 1988 6316 1990
rect 2665 1986 6334 1988
rect 2665 1974 6353 1986
rect 2665 1920 2690 1974
rect 2763 1920 2834 1974
rect 2907 1920 2978 1974
rect 3051 1920 3122 1974
rect 3195 1920 3266 1974
rect 3339 1920 3410 1974
rect 3483 1920 3554 1974
rect 3627 1920 3698 1974
rect 3771 1920 3842 1974
rect 3915 1920 3986 1974
rect 4059 1920 4130 1974
rect 4203 1920 4274 1974
rect 4347 1920 4418 1974
rect 4491 1920 4562 1974
rect 4635 1920 4706 1974
rect 4779 1920 4850 1974
rect 4923 1920 4994 1974
rect 5067 1920 5138 1974
rect 5211 1920 5282 1974
rect 5355 1920 5426 1974
rect 5499 1920 5570 1974
rect 5643 1920 5714 1974
rect 5787 1920 5858 1974
rect 5931 1920 6002 1974
rect 6075 1920 6146 1974
rect 6219 1920 6353 1974
rect 2665 1892 6353 1920
rect 2665 1826 2764 1892
rect 2665 1772 2678 1826
rect 2751 1772 2764 1826
rect 6231 1854 6353 1892
rect 6231 1800 6254 1854
rect 6327 1800 6353 1854
rect 2665 1706 2764 1772
rect 2665 1652 2678 1706
rect 2751 1652 2764 1706
rect 2665 1586 2764 1652
rect 6231 1734 6353 1800
rect 2665 1532 2678 1586
rect 2751 1532 2764 1586
rect 2665 1466 2764 1532
rect 2665 1412 2678 1466
rect 2751 1412 2764 1466
rect 6231 1680 6254 1734
rect 6327 1680 6353 1734
rect 2665 1346 2764 1412
rect 2665 1292 2678 1346
rect 2751 1292 2764 1346
rect 2665 1226 2764 1292
rect 2665 1172 2678 1226
rect 2751 1172 2764 1226
rect 6231 1614 6353 1680
rect 6231 1560 6254 1614
rect 6327 1560 6353 1614
rect 2665 1106 2764 1172
rect 2665 1052 2678 1106
rect 2751 1052 2764 1106
rect 2665 986 2764 1052
rect 2665 932 2678 986
rect 2751 932 2764 986
rect 2665 866 2764 932
rect 2665 812 2678 866
rect 2751 812 2764 866
rect 2665 746 2764 812
rect 2665 692 2678 746
rect 2751 692 2764 746
rect 2665 626 2764 692
rect 6231 1494 6353 1560
rect 6231 1440 6254 1494
rect 6327 1440 6353 1494
rect 6231 1374 6353 1440
rect 6231 1320 6254 1374
rect 6327 1320 6353 1374
rect 6231 1254 6353 1320
rect 6231 1200 6254 1254
rect 6327 1200 6353 1254
rect 6231 1134 6353 1200
rect 6231 1080 6254 1134
rect 6327 1080 6353 1134
rect 6231 1014 6353 1080
rect 6231 960 6254 1014
rect 6327 960 6353 1014
rect 6231 894 6353 960
rect 2665 572 2678 626
rect 2751 572 2764 626
rect -876 511 1629 537
rect -876 436 -801 511
rect 1521 436 1629 511
rect -876 413 1629 436
rect 2665 506 2764 572
rect 6231 840 6254 894
rect 6327 840 6353 894
rect 6231 774 6353 840
rect 6231 720 6254 774
rect 6327 720 6353 774
rect 6231 654 6353 720
rect 6231 600 6254 654
rect 6327 600 6353 654
rect 2665 452 2678 506
rect 2751 452 2764 506
rect 2665 386 2764 452
rect 2665 332 2678 386
rect 2751 332 2764 386
rect 6231 534 6353 600
rect 6231 480 6254 534
rect 6327 480 6353 534
rect 6231 414 6353 480
rect 2665 266 2764 332
rect 2665 212 2678 266
rect 2751 212 2764 266
rect 2665 146 2764 212
rect 2665 92 2678 146
rect 2751 92 2764 146
rect 6231 360 6254 414
rect 6327 360 6353 414
rect 2665 26 2764 92
rect 2665 -28 2678 26
rect 2751 -28 2764 26
rect 2665 -94 2764 -28
rect 2665 -148 2678 -94
rect 2751 -148 2764 -94
rect 2665 -214 2764 -148
rect 2665 -268 2678 -214
rect 2751 -268 2764 -214
rect 6231 294 6353 360
rect 6231 240 6254 294
rect 6327 240 6353 294
rect 6231 174 6353 240
rect 6231 120 6254 174
rect 6327 120 6353 174
rect 6231 54 6353 120
rect 2665 -334 2764 -268
rect 2665 -388 2678 -334
rect 2751 -388 2764 -334
rect 2665 -454 2764 -388
rect 2665 -508 2678 -454
rect 2751 -508 2764 -454
rect 2665 -574 2764 -508
rect 6231 0 6254 54
rect 6327 0 6353 54
rect 6231 -66 6353 0
rect 6231 -120 6254 -66
rect 6327 -120 6353 -66
rect 6231 -186 6353 -120
rect -764 -603 1707 -578
rect -764 -681 -656 -603
rect 1599 -681 1707 -603
rect -764 -706 1707 -681
rect 2665 -628 2678 -574
rect 2751 -628 2764 -574
rect 2665 -694 2764 -628
rect 6231 -240 6254 -186
rect 6327 -240 6353 -186
rect 6231 -306 6353 -240
rect 6231 -360 6254 -306
rect 6327 -360 6353 -306
rect 6231 -426 6353 -360
rect 6231 -480 6254 -426
rect 6327 -480 6353 -426
rect 6231 -546 6353 -480
rect 2665 -748 2678 -694
rect 2751 -748 2764 -694
rect 2665 -814 2764 -748
rect 6231 -600 6254 -546
rect 6327 -600 6353 -546
rect 2665 -868 2678 -814
rect 2751 -868 2764 -814
rect 2665 -934 2764 -868
rect 2665 -988 2678 -934
rect 2751 -988 2764 -934
rect 2665 -1054 2764 -988
rect 2665 -1108 2678 -1054
rect 2751 -1108 2764 -1054
rect 2665 -1174 2764 -1108
rect 2665 -1228 2678 -1174
rect 2751 -1228 2764 -1174
rect 6231 -666 6353 -600
rect 6231 -720 6254 -666
rect 6327 -720 6353 -666
rect 6231 -786 6353 -720
rect 6231 -840 6254 -786
rect 6327 -840 6353 -786
rect 6231 -906 6353 -840
rect 6231 -960 6254 -906
rect 6327 -960 6353 -906
rect 6231 -1026 6353 -960
rect 6231 -1080 6254 -1026
rect 6327 -1080 6353 -1026
rect 2665 -1294 2764 -1228
rect 2665 -1348 2678 -1294
rect 2751 -1348 2764 -1294
rect 2665 -1414 2764 -1348
rect 2665 -1468 2678 -1414
rect 2751 -1468 2764 -1414
rect 6231 -1146 6353 -1080
rect 6231 -1200 6254 -1146
rect 6327 -1200 6353 -1146
rect 6231 -1266 6353 -1200
rect 6231 -1320 6254 -1266
rect 6327 -1320 6353 -1266
rect 6231 -1386 6353 -1320
rect 2665 -1550 2764 -1468
rect 6231 -1440 6254 -1386
rect 6327 -1440 6353 -1386
rect 3241 -1549 3435 -1548
rect 6231 -1549 6353 -1440
rect 3241 -1550 6452 -1549
rect 2665 -1564 6452 -1550
rect 2665 -1578 2681 -1564
rect 2667 -1618 2681 -1578
rect 2754 -1618 2806 -1564
rect 2879 -1618 2931 -1564
rect 3004 -1618 3056 -1564
rect 3129 -1618 3181 -1564
rect 3254 -1565 6452 -1564
rect 3254 -1614 3318 -1565
rect 3381 -1566 6229 -1565
rect 3381 -1614 3439 -1566
rect 3254 -1615 3439 -1614
rect 3502 -1615 3560 -1566
rect 3623 -1615 3681 -1566
rect 3744 -1615 3802 -1566
rect 3865 -1615 3923 -1566
rect 3986 -1615 4044 -1566
rect 4107 -1615 4165 -1566
rect 4228 -1615 4286 -1566
rect 4349 -1615 4407 -1566
rect 4470 -1615 4528 -1566
rect 4591 -1615 4649 -1566
rect 4712 -1615 4770 -1566
rect 4833 -1615 4891 -1566
rect 4954 -1615 5012 -1566
rect 5075 -1615 5133 -1566
rect 5196 -1615 5254 -1566
rect 5317 -1615 5375 -1566
rect 5438 -1615 5496 -1566
rect 5559 -1615 5617 -1566
rect 5680 -1615 5738 -1566
rect 5801 -1615 5859 -1566
rect 5922 -1615 5980 -1566
rect 6043 -1615 6101 -1566
rect 6164 -1614 6229 -1566
rect 6292 -1584 6452 -1565
rect 6292 -1614 6375 -1584
rect 6164 -1615 6375 -1614
rect 3254 -1618 6375 -1615
rect 2667 -1629 6375 -1618
rect 2667 -1635 3333 -1629
rect 3240 -1760 3333 -1635
rect 6360 -1633 6375 -1629
rect 6438 -1633 6452 -1584
rect 3240 -1809 3255 -1760
rect 3318 -1809 3333 -1760
rect 6360 -1691 6452 -1633
rect 6360 -1719 6375 -1691
rect 3240 -1871 3333 -1809
rect 3240 -1920 3255 -1871
rect 3318 -1920 3333 -1871
rect 6359 -1740 6375 -1719
rect 6438 -1740 6452 -1691
rect 6359 -1791 6452 -1740
rect 6359 -1840 6374 -1791
rect 6437 -1840 6452 -1791
rect 6359 -1902 6452 -1840
rect 3240 -1982 3333 -1920
rect -1189 -2029 1828 -2013
rect -1189 -2080 -1162 -2029
rect 1713 -2080 1828 -2029
rect -1189 -2094 1828 -2080
rect 3240 -2031 3255 -1982
rect 3318 -2031 3333 -1982
rect 6359 -1951 6374 -1902
rect 6437 -1951 6452 -1902
rect 6359 -2013 6452 -1951
rect 3240 -2093 3333 -2031
rect 3240 -2142 3255 -2093
rect 3318 -2142 3333 -2093
rect 6359 -2062 6374 -2013
rect 6437 -2062 6452 -2013
rect 3240 -2204 3333 -2142
rect 3240 -2253 3255 -2204
rect 3318 -2253 3333 -2204
rect 3240 -2315 3333 -2253
rect 6359 -2124 6452 -2062
rect 6359 -2173 6374 -2124
rect 6437 -2173 6452 -2124
rect 6359 -2235 6452 -2173
rect 6359 -2284 6374 -2235
rect 6437 -2284 6452 -2235
rect 3240 -2364 3255 -2315
rect 3318 -2364 3333 -2315
rect 3240 -2426 3333 -2364
rect 6359 -2346 6452 -2284
rect 6359 -2395 6374 -2346
rect 6437 -2395 6452 -2346
rect 3240 -2475 3255 -2426
rect 3318 -2475 3333 -2426
rect -274 -2548 2823 -2535
rect -274 -2549 502 -2548
rect -274 -2598 -236 -2549
rect -173 -2550 21 -2549
rect -173 -2598 -108 -2550
rect -274 -2599 -108 -2598
rect -45 -2598 21 -2550
rect 84 -2550 373 -2549
rect 84 -2598 138 -2550
rect -45 -2599 138 -2598
rect 201 -2551 373 -2550
rect 201 -2599 250 -2551
rect -274 -2600 250 -2599
rect 313 -2598 373 -2551
rect 436 -2597 502 -2549
rect 565 -2549 1104 -2548
rect 565 -2597 619 -2549
rect 436 -2598 619 -2597
rect 682 -2550 975 -2549
rect 682 -2598 731 -2550
rect 313 -2599 731 -2598
rect 794 -2599 849 -2550
rect 912 -2598 975 -2550
rect 1038 -2597 1104 -2549
rect 1167 -2549 2823 -2548
rect 1167 -2597 1221 -2549
rect 1038 -2598 1221 -2597
rect 1284 -2550 2823 -2549
rect 1284 -2598 1333 -2550
rect 912 -2599 1333 -2598
rect 1396 -2599 1451 -2550
rect 1514 -2599 1574 -2550
rect 1637 -2599 1691 -2550
rect 1754 -2599 1812 -2550
rect 1875 -2599 1934 -2550
rect 1997 -2551 2516 -2550
rect 1997 -2599 2045 -2551
rect 313 -2600 2045 -2599
rect 2108 -2600 2164 -2551
rect 2227 -2600 2276 -2551
rect 2339 -2600 2397 -2551
rect 2460 -2599 2516 -2551
rect 2579 -2552 2742 -2550
rect 2579 -2599 2631 -2552
rect 2460 -2600 2631 -2599
rect -274 -2601 2631 -2600
rect 2694 -2599 2742 -2552
rect 2805 -2599 2823 -2550
rect 2694 -2601 2823 -2599
rect -274 -2615 2823 -2601
rect -274 -2664 -180 -2615
rect -274 -2711 -250 -2664
rect -196 -2711 -180 -2664
rect 2737 -2650 2823 -2615
rect -274 -2765 -180 -2711
rect -274 -2812 -249 -2765
rect -195 -2812 -180 -2765
rect -274 -2862 -180 -2812
rect -274 -2909 -250 -2862
rect -196 -2909 -180 -2862
rect 2737 -2697 2753 -2650
rect 2807 -2697 2823 -2650
rect 2737 -2751 2823 -2697
rect 2737 -2798 2754 -2751
rect 2808 -2798 2823 -2751
rect 2737 -2848 2823 -2798
rect -274 -2970 -180 -2909
rect -274 -3017 -249 -2970
rect -195 -3017 -180 -2970
rect 2737 -2895 2753 -2848
rect 2807 -2895 2823 -2848
rect 2737 -2956 2823 -2895
rect 2737 -3003 2754 -2956
rect 2808 -3003 2823 -2956
rect -274 -3095 -180 -3017
rect -274 -3142 -249 -3095
rect -195 -3142 -180 -3095
rect -274 -3209 -180 -3142
rect 2737 -3081 2823 -3003
rect 2737 -3128 2754 -3081
rect 2808 -3128 2823 -3081
rect -274 -3256 -248 -3209
rect -194 -3256 -180 -3209
rect -274 -3321 -180 -3256
rect 2737 -3195 2823 -3128
rect 2737 -3242 2755 -3195
rect 2809 -3242 2823 -3195
rect -274 -3368 -247 -3321
rect -193 -3368 -180 -3321
rect -274 -3425 -180 -3368
rect -274 -3472 -249 -3425
rect -195 -3472 -180 -3425
rect -274 -3529 -180 -3472
rect -274 -3576 -249 -3529
rect -195 -3576 -180 -3529
rect 2737 -3307 2823 -3242
rect 2737 -3354 2756 -3307
rect 2810 -3354 2823 -3307
rect 2737 -3411 2823 -3354
rect 2737 -3458 2754 -3411
rect 2808 -3458 2823 -3411
rect 2737 -3515 2823 -3458
rect -2118 -3605 -1770 -3592
rect -2118 -3654 -2099 -3605
rect -1790 -3654 -1770 -3605
rect -2118 -3669 -1770 -3654
rect -1586 -3603 -815 -3588
rect -1586 -3649 -1567 -3603
rect -838 -3649 -815 -3603
rect -1586 -3664 -815 -3649
rect -274 -3624 -180 -3576
rect -274 -3671 -251 -3624
rect -197 -3671 -180 -3624
rect -274 -3733 -180 -3671
rect 2737 -3562 2754 -3515
rect 2808 -3562 2823 -3515
rect 2737 -3610 2823 -3562
rect 2737 -3657 2752 -3610
rect 2806 -3657 2823 -3610
rect -274 -3780 -250 -3733
rect -196 -3780 -180 -3733
rect -274 -3837 -180 -3780
rect 2737 -3719 2823 -3657
rect 2737 -3766 2753 -3719
rect 2807 -3766 2823 -3719
rect 2737 -3823 2823 -3766
rect -274 -3884 -250 -3837
rect -196 -3884 -180 -3837
rect -274 -3932 -180 -3884
rect -274 -3979 -252 -3932
rect -198 -3979 -180 -3932
rect -274 -4042 -180 -3979
rect -274 -4089 -251 -4042
rect -197 -4089 -180 -4042
rect 2737 -3870 2753 -3823
rect 2807 -3870 2823 -3823
rect 2737 -3918 2823 -3870
rect -274 -4146 -180 -4089
rect 2737 -3965 2751 -3918
rect 2805 -3965 2823 -3918
rect 2737 -4028 2823 -3965
rect 2737 -4075 2752 -4028
rect 2806 -4075 2823 -4028
rect -274 -4193 -251 -4146
rect -197 -4193 -180 -4146
rect -274 -4241 -180 -4193
rect 2737 -4132 2823 -4075
rect 2737 -4179 2752 -4132
rect 2806 -4179 2823 -4132
rect -274 -4288 -253 -4241
rect -199 -4288 -180 -4241
rect -274 -4342 -180 -4288
rect -274 -4389 -250 -4342
rect -196 -4389 -180 -4342
rect 2737 -4227 2823 -4179
rect 2737 -4274 2750 -4227
rect 2804 -4274 2823 -4227
rect 2737 -4328 2823 -4274
rect 2737 -4375 2753 -4328
rect 2807 -4375 2823 -4328
rect -274 -4446 -180 -4389
rect -2118 -4473 -1770 -4460
rect -2118 -4522 -2099 -4473
rect -1790 -4522 -1770 -4473
rect -2118 -4537 -1770 -4522
rect -1586 -4471 -815 -4456
rect -1586 -4517 -1567 -4471
rect -838 -4517 -815 -4471
rect -1586 -4532 -815 -4517
rect -274 -4493 -250 -4446
rect -196 -4493 -180 -4446
rect -274 -4541 -180 -4493
rect 2737 -4432 2823 -4375
rect 2737 -4479 2753 -4432
rect 2807 -4479 2823 -4432
rect -274 -4588 -252 -4541
rect -198 -4588 -180 -4541
rect -274 -4651 -180 -4588
rect 2737 -4527 2823 -4479
rect 2737 -4574 2751 -4527
rect 2805 -4574 2823 -4527
rect -274 -4698 -251 -4651
rect -197 -4698 -180 -4651
rect -274 -4755 -180 -4698
rect -274 -4802 -251 -4755
rect -197 -4802 -180 -4755
rect 2737 -4637 2823 -4574
rect 2737 -4684 2752 -4637
rect 2806 -4684 2823 -4637
rect 2737 -4741 2823 -4684
rect -274 -4850 -180 -4802
rect -274 -4897 -253 -4850
rect -199 -4897 -180 -4850
rect 2737 -4788 2752 -4741
rect 2806 -4788 2823 -4741
rect 2737 -4836 2823 -4788
rect 2737 -4883 2750 -4836
rect 2804 -4883 2823 -4836
rect -274 -4954 -180 -4897
rect -274 -5001 -249 -4954
rect -195 -5001 -180 -4954
rect -274 -5064 -180 -5001
rect -274 -5111 -248 -5064
rect -194 -5111 -180 -5064
rect 2737 -4940 2823 -4883
rect 2737 -4987 2754 -4940
rect 2808 -4987 2823 -4940
rect 2737 -5050 2823 -4987
rect -274 -5168 -180 -5111
rect -274 -5215 -248 -5168
rect -194 -5215 -180 -5168
rect -274 -5272 -180 -5215
rect 2737 -5097 2755 -5050
rect 2809 -5097 2823 -5050
rect 2737 -5154 2823 -5097
rect 2737 -5201 2755 -5154
rect 2809 -5201 2823 -5154
rect 2737 -5272 2823 -5201
rect -274 -5285 2823 -5272
rect -274 -5286 499 -5285
rect -2118 -5332 -1770 -5319
rect -2118 -5381 -2099 -5332
rect -1790 -5381 -1770 -5332
rect -2118 -5396 -1770 -5381
rect -1586 -5330 -815 -5315
rect -1586 -5376 -1567 -5330
rect -838 -5376 -815 -5330
rect -274 -5335 -239 -5286
rect -176 -5287 18 -5286
rect -176 -5335 -111 -5287
rect -274 -5336 -111 -5335
rect -48 -5335 18 -5287
rect 81 -5287 370 -5286
rect 81 -5335 135 -5287
rect -48 -5336 135 -5335
rect 198 -5288 370 -5287
rect 198 -5336 247 -5288
rect -274 -5337 247 -5336
rect 310 -5335 370 -5288
rect 433 -5334 499 -5286
rect 562 -5286 1101 -5285
rect 562 -5334 616 -5286
rect 433 -5335 616 -5334
rect 679 -5287 972 -5286
rect 679 -5335 728 -5287
rect 310 -5336 728 -5335
rect 791 -5336 846 -5287
rect 909 -5335 972 -5287
rect 1035 -5334 1101 -5286
rect 1164 -5286 2823 -5285
rect 1164 -5334 1218 -5286
rect 1035 -5335 1218 -5334
rect 1281 -5287 2823 -5286
rect 1281 -5335 1330 -5287
rect 909 -5336 1330 -5335
rect 1393 -5336 1448 -5287
rect 1511 -5336 1571 -5287
rect 1634 -5336 1688 -5287
rect 1751 -5336 1809 -5287
rect 1872 -5336 1931 -5287
rect 1994 -5288 2513 -5287
rect 1994 -5336 2042 -5288
rect 310 -5337 2042 -5336
rect 2105 -5337 2161 -5288
rect 2224 -5337 2273 -5288
rect 2336 -5337 2394 -5288
rect 2457 -5336 2513 -5288
rect 2576 -5289 2739 -5287
rect 2576 -5336 2628 -5289
rect 2457 -5337 2628 -5336
rect -274 -5338 2628 -5337
rect 2691 -5336 2739 -5289
rect 2802 -5336 2823 -5287
rect 2691 -5338 2823 -5336
rect -274 -5352 2823 -5338
rect 3240 -2537 3333 -2475
rect 3240 -2586 3255 -2537
rect 3318 -2586 3333 -2537
rect 6359 -2457 6452 -2395
rect 6359 -2506 6374 -2457
rect 6437 -2506 6452 -2457
rect 6359 -2568 6452 -2506
rect 3240 -2648 3333 -2586
rect 3240 -2697 3255 -2648
rect 3318 -2697 3333 -2648
rect 3240 -2759 3333 -2697
rect 6359 -2617 6374 -2568
rect 6437 -2617 6452 -2568
rect 6359 -2679 6452 -2617
rect 3240 -2808 3255 -2759
rect 3318 -2808 3333 -2759
rect 3240 -2870 3333 -2808
rect 3240 -2919 3255 -2870
rect 3318 -2919 3333 -2870
rect 6359 -2728 6374 -2679
rect 6437 -2728 6452 -2679
rect 6359 -2790 6452 -2728
rect 3240 -2981 3333 -2919
rect 6359 -2839 6374 -2790
rect 6437 -2839 6452 -2790
rect 6359 -2901 6452 -2839
rect 6359 -2950 6374 -2901
rect 6437 -2950 6452 -2901
rect 3240 -3030 3255 -2981
rect 3318 -3030 3333 -2981
rect 3240 -3092 3333 -3030
rect 6359 -3012 6452 -2950
rect 6359 -3061 6374 -3012
rect 6437 -3061 6452 -3012
rect 3240 -3141 3255 -3092
rect 3318 -3141 3333 -3092
rect 3240 -3203 3333 -3141
rect 3240 -3252 3255 -3203
rect 3318 -3252 3333 -3203
rect 3240 -3314 3333 -3252
rect 6359 -3123 6452 -3061
rect 6359 -3172 6374 -3123
rect 6437 -3172 6452 -3123
rect 6359 -3234 6452 -3172
rect 3240 -3363 3255 -3314
rect 3318 -3363 3333 -3314
rect 3240 -3425 3333 -3363
rect 6359 -3283 6374 -3234
rect 6437 -3283 6452 -3234
rect 6359 -3345 6452 -3283
rect 6359 -3394 6374 -3345
rect 6437 -3394 6452 -3345
rect 3240 -3474 3255 -3425
rect 3318 -3474 3333 -3425
rect 3240 -3536 3333 -3474
rect 6359 -3456 6452 -3394
rect 3240 -3585 3255 -3536
rect 3318 -3585 3333 -3536
rect 3240 -3647 3333 -3585
rect 6359 -3505 6374 -3456
rect 6437 -3505 6452 -3456
rect 6359 -3567 6452 -3505
rect 3240 -3696 3255 -3647
rect 3318 -3696 3333 -3647
rect 3240 -3758 3333 -3696
rect 6359 -3616 6374 -3567
rect 6437 -3616 6452 -3567
rect 6359 -3678 6452 -3616
rect 3240 -3807 3255 -3758
rect 3318 -3807 3333 -3758
rect 3240 -3869 3333 -3807
rect 6359 -3727 6374 -3678
rect 6437 -3727 6452 -3678
rect 6359 -3789 6452 -3727
rect 3240 -3918 3255 -3869
rect 3318 -3918 3333 -3869
rect 3240 -3980 3333 -3918
rect 3240 -4029 3255 -3980
rect 3318 -4029 3333 -3980
rect 6359 -3838 6374 -3789
rect 6437 -3838 6452 -3789
rect 6359 -3900 6452 -3838
rect 6359 -3949 6374 -3900
rect 6437 -3949 6452 -3900
rect 3240 -4091 3333 -4029
rect 3240 -4140 3255 -4091
rect 3318 -4140 3333 -4091
rect 6359 -4011 6452 -3949
rect 6359 -4060 6374 -4011
rect 6437 -4060 6452 -4011
rect 3240 -4202 3333 -4140
rect 3240 -4251 3255 -4202
rect 3318 -4251 3333 -4202
rect 3240 -4313 3333 -4251
rect 6359 -4122 6452 -4060
rect 6359 -4171 6374 -4122
rect 6437 -4171 6452 -4122
rect 6359 -4233 6452 -4171
rect 6359 -4282 6374 -4233
rect 6437 -4282 6452 -4233
rect 3240 -4362 3255 -4313
rect 3318 -4362 3333 -4313
rect 3240 -4424 3333 -4362
rect 6359 -4344 6452 -4282
rect 6359 -4393 6374 -4344
rect 6437 -4393 6452 -4344
rect 3240 -4473 3255 -4424
rect 3318 -4473 3333 -4424
rect 3240 -4535 3333 -4473
rect 3240 -4584 3255 -4535
rect 3318 -4584 3333 -4535
rect 6359 -4455 6452 -4393
rect 3240 -4646 3333 -4584
rect 3240 -4695 3255 -4646
rect 3318 -4695 3333 -4646
rect 6359 -4504 6374 -4455
rect 6437 -4504 6452 -4455
rect 6359 -4566 6452 -4504
rect 6359 -4615 6374 -4566
rect 6437 -4615 6452 -4566
rect 3240 -4757 3333 -4695
rect 3240 -4806 3255 -4757
rect 3318 -4806 3333 -4757
rect 6359 -4677 6452 -4615
rect 6359 -4726 6374 -4677
rect 6437 -4726 6452 -4677
rect 3240 -4868 3333 -4806
rect 3240 -4917 3255 -4868
rect 3318 -4917 3333 -4868
rect 3240 -4979 3333 -4917
rect 3240 -5028 3255 -4979
rect 3318 -5028 3333 -4979
rect 6359 -4788 6452 -4726
rect 6359 -4837 6374 -4788
rect 6437 -4837 6452 -4788
rect 6359 -4899 6452 -4837
rect 6359 -4948 6374 -4899
rect 6437 -4948 6452 -4899
rect 3240 -5090 3333 -5028
rect 3240 -5139 3255 -5090
rect 3318 -5139 3333 -5090
rect 6359 -5010 6452 -4948
rect 6359 -5059 6374 -5010
rect 6437 -5059 6452 -5010
rect 3240 -5201 3333 -5139
rect 3240 -5250 3255 -5201
rect 3318 -5250 3333 -5201
rect 6359 -5121 6452 -5059
rect 6359 -5170 6374 -5121
rect 6437 -5170 6452 -5121
rect 3240 -5312 3333 -5250
rect -1586 -5391 -815 -5376
rect 3240 -5361 3255 -5312
rect 3318 -5361 3333 -5312
rect 3240 -5423 3333 -5361
rect 6359 -5232 6452 -5170
rect 6359 -5281 6374 -5232
rect 6437 -5281 6452 -5232
rect 6359 -5343 6452 -5281
rect 3240 -5472 3255 -5423
rect 3318 -5472 3333 -5423
rect 3240 -5534 3333 -5472
rect 6359 -5392 6374 -5343
rect 6437 -5392 6452 -5343
rect 6359 -5454 6452 -5392
rect 6359 -5503 6374 -5454
rect 6437 -5503 6452 -5454
rect 3240 -5583 3255 -5534
rect 3318 -5583 3333 -5534
rect 3240 -5645 3333 -5583
rect 3240 -5694 3255 -5645
rect 3318 -5694 3333 -5645
rect 6359 -5565 6452 -5503
rect 6359 -5614 6374 -5565
rect 6437 -5614 6452 -5565
rect 6359 -5676 6452 -5614
rect 3240 -5756 3333 -5694
rect 3240 -5805 3255 -5756
rect 3318 -5805 3333 -5756
rect 6359 -5725 6374 -5676
rect 6437 -5725 6452 -5676
rect 6359 -5787 6452 -5725
rect 3240 -5867 3333 -5805
rect 3240 -5916 3255 -5867
rect 3318 -5916 3333 -5867
rect 3240 -5978 3333 -5916
rect 6359 -5836 6374 -5787
rect 6437 -5836 6452 -5787
rect 6359 -5898 6452 -5836
rect 3240 -6027 3255 -5978
rect 3318 -6027 3333 -5978
rect 3240 -6089 3333 -6027
rect 6359 -5947 6374 -5898
rect 6437 -5947 6452 -5898
rect 6359 -6009 6452 -5947
rect 6359 -6058 6374 -6009
rect 6437 -6058 6452 -6009
rect 3240 -6138 3255 -6089
rect 3318 -6138 3333 -6089
rect -2118 -6200 -1770 -6187
rect -2118 -6249 -2099 -6200
rect -1790 -6249 -1770 -6200
rect -2118 -6264 -1770 -6249
rect -1586 -6198 -815 -6183
rect -1586 -6244 -1567 -6198
rect -838 -6244 -815 -6198
rect -1586 -6259 -815 -6244
rect -500 -6200 -152 -6187
rect -500 -6249 -481 -6200
rect -172 -6249 -152 -6200
rect -500 -6264 -152 -6249
rect 32 -6198 803 -6183
rect 32 -6244 51 -6198
rect 780 -6244 803 -6198
rect 32 -6259 803 -6244
rect 1109 -6200 1457 -6187
rect 1109 -6249 1128 -6200
rect 1437 -6249 1457 -6200
rect 1109 -6264 1457 -6249
rect 1641 -6198 2412 -6183
rect 1641 -6244 1660 -6198
rect 2389 -6244 2412 -6198
rect 1641 -6259 2412 -6244
rect 3240 -6200 3333 -6138
rect 6359 -6120 6452 -6058
rect 6359 -6169 6374 -6120
rect 6437 -6169 6452 -6120
rect 3240 -6249 3255 -6200
rect 3318 -6249 3333 -6200
rect 3240 -6311 3333 -6249
rect 3240 -6360 3255 -6311
rect 3318 -6360 3333 -6311
rect 6359 -6231 6452 -6169
rect 3240 -6422 3333 -6360
rect 6359 -6280 6374 -6231
rect 6437 -6280 6452 -6231
rect 6359 -6342 6452 -6280
rect 3240 -6471 3255 -6422
rect 3318 -6471 3333 -6422
rect 3240 -6594 3333 -6471
rect 6359 -6391 6374 -6342
rect 6437 -6391 6452 -6342
rect 6359 -6453 6452 -6391
rect 6359 -6502 6374 -6453
rect 6437 -6502 6452 -6453
rect 3240 -6595 3435 -6594
rect 6359 -6595 6452 -6502
rect 3240 -6611 6452 -6595
rect 3240 -6660 3318 -6611
rect 3381 -6612 6452 -6611
rect 3381 -6660 3439 -6612
rect 3240 -6661 3439 -6660
rect 3502 -6661 3560 -6612
rect 3623 -6661 3681 -6612
rect 3744 -6661 3802 -6612
rect 3865 -6661 3923 -6612
rect 3986 -6661 4044 -6612
rect 4107 -6661 4165 -6612
rect 4228 -6661 4286 -6612
rect 4349 -6661 4407 -6612
rect 4470 -6661 4528 -6612
rect 4591 -6661 4649 -6612
rect 4712 -6661 4770 -6612
rect 4833 -6661 4891 -6612
rect 4954 -6661 5012 -6612
rect 5075 -6661 5133 -6612
rect 5196 -6661 5254 -6612
rect 5317 -6661 5375 -6612
rect 5438 -6661 5496 -6612
rect 5559 -6661 5617 -6612
rect 5680 -6661 5738 -6612
rect 5801 -6661 5859 -6612
rect 5922 -6661 5980 -6612
rect 6043 -6661 6101 -6612
rect 6164 -6661 6452 -6612
rect 3240 -6675 6452 -6661
rect 3240 -6677 3333 -6675
<< nsubdiff >>
rect -2104 -2914 -1812 -2897
rect -2104 -2965 -2084 -2914
rect -1834 -2965 -1812 -2914
rect -2104 -2982 -1812 -2965
rect -1580 -2909 -817 -2894
rect -1580 -2955 -1551 -2909
rect -839 -2955 -817 -2909
rect -1580 -2968 -817 -2955
rect -2104 -3782 -1812 -3765
rect -2104 -3833 -2084 -3782
rect -1834 -3833 -1812 -3782
rect -2104 -3850 -1812 -3833
rect -1580 -3777 -817 -3762
rect -1580 -3823 -1551 -3777
rect -839 -3823 -817 -3777
rect -1580 -3836 -817 -3823
rect -2104 -4641 -1812 -4624
rect -2104 -4692 -2084 -4641
rect -1834 -4692 -1812 -4641
rect -2104 -4709 -1812 -4692
rect -1580 -4636 -817 -4621
rect -1580 -4682 -1551 -4636
rect -839 -4682 -817 -4636
rect -1580 -4695 -817 -4682
rect -2104 -5509 -1812 -5492
rect -2104 -5560 -2084 -5509
rect -1834 -5560 -1812 -5509
rect -2104 -5577 -1812 -5560
rect -1580 -5504 -817 -5489
rect -1580 -5550 -1551 -5504
rect -839 -5550 -817 -5504
rect -1580 -5563 -817 -5550
rect -486 -5509 -194 -5492
rect -486 -5560 -466 -5509
rect -216 -5560 -194 -5509
rect -486 -5577 -194 -5560
rect 38 -5504 801 -5489
rect 38 -5550 67 -5504
rect 779 -5550 801 -5504
rect 38 -5563 801 -5550
rect 1123 -5509 1415 -5492
rect 1123 -5560 1143 -5509
rect 1393 -5560 1415 -5509
rect 1123 -5577 1415 -5560
rect 1647 -5504 2410 -5489
rect 1647 -5550 1676 -5504
rect 2388 -5550 2410 -5504
rect 1647 -5563 2410 -5550
<< psubdiffcont >>
rect -1191 1938 1787 2008
rect 2690 1920 2763 1974
rect 2834 1920 2907 1974
rect 2978 1920 3051 1974
rect 3122 1920 3195 1974
rect 3266 1920 3339 1974
rect 3410 1920 3483 1974
rect 3554 1920 3627 1974
rect 3698 1920 3771 1974
rect 3842 1920 3915 1974
rect 3986 1920 4059 1974
rect 4130 1920 4203 1974
rect 4274 1920 4347 1974
rect 4418 1920 4491 1974
rect 4562 1920 4635 1974
rect 4706 1920 4779 1974
rect 4850 1920 4923 1974
rect 4994 1920 5067 1974
rect 5138 1920 5211 1974
rect 5282 1920 5355 1974
rect 5426 1920 5499 1974
rect 5570 1920 5643 1974
rect 5714 1920 5787 1974
rect 5858 1920 5931 1974
rect 6002 1920 6075 1974
rect 6146 1920 6219 1974
rect 2678 1772 2751 1826
rect 6254 1800 6327 1854
rect 2678 1652 2751 1706
rect 2678 1532 2751 1586
rect 2678 1412 2751 1466
rect 6254 1680 6327 1734
rect 2678 1292 2751 1346
rect 2678 1172 2751 1226
rect 6254 1560 6327 1614
rect 2678 1052 2751 1106
rect 2678 932 2751 986
rect 2678 812 2751 866
rect 2678 692 2751 746
rect 6254 1440 6327 1494
rect 6254 1320 6327 1374
rect 6254 1200 6327 1254
rect 6254 1080 6327 1134
rect 6254 960 6327 1014
rect 2678 572 2751 626
rect -801 436 1521 511
rect 6254 840 6327 894
rect 6254 720 6327 774
rect 6254 600 6327 654
rect 2678 452 2751 506
rect 2678 332 2751 386
rect 6254 480 6327 534
rect 2678 212 2751 266
rect 2678 92 2751 146
rect 6254 360 6327 414
rect 2678 -28 2751 26
rect 2678 -148 2751 -94
rect 2678 -268 2751 -214
rect 6254 240 6327 294
rect 6254 120 6327 174
rect 2678 -388 2751 -334
rect 2678 -508 2751 -454
rect 6254 0 6327 54
rect 6254 -120 6327 -66
rect -656 -681 1599 -603
rect 2678 -628 2751 -574
rect 6254 -240 6327 -186
rect 6254 -360 6327 -306
rect 6254 -480 6327 -426
rect 2678 -748 2751 -694
rect 6254 -600 6327 -546
rect 2678 -868 2751 -814
rect 2678 -988 2751 -934
rect 2678 -1108 2751 -1054
rect 2678 -1228 2751 -1174
rect 6254 -720 6327 -666
rect 6254 -840 6327 -786
rect 6254 -960 6327 -906
rect 6254 -1080 6327 -1026
rect 2678 -1348 2751 -1294
rect 2678 -1468 2751 -1414
rect 6254 -1200 6327 -1146
rect 6254 -1320 6327 -1266
rect 6254 -1440 6327 -1386
rect 2681 -1618 2754 -1564
rect 2806 -1618 2879 -1564
rect 2931 -1618 3004 -1564
rect 3056 -1618 3129 -1564
rect 3181 -1618 3254 -1564
rect 3318 -1614 3381 -1565
rect 3439 -1615 3502 -1566
rect 3560 -1615 3623 -1566
rect 3681 -1615 3744 -1566
rect 3802 -1615 3865 -1566
rect 3923 -1615 3986 -1566
rect 4044 -1615 4107 -1566
rect 4165 -1615 4228 -1566
rect 4286 -1615 4349 -1566
rect 4407 -1615 4470 -1566
rect 4528 -1615 4591 -1566
rect 4649 -1615 4712 -1566
rect 4770 -1615 4833 -1566
rect 4891 -1615 4954 -1566
rect 5012 -1615 5075 -1566
rect 5133 -1615 5196 -1566
rect 5254 -1615 5317 -1566
rect 5375 -1615 5438 -1566
rect 5496 -1615 5559 -1566
rect 5617 -1615 5680 -1566
rect 5738 -1615 5801 -1566
rect 5859 -1615 5922 -1566
rect 5980 -1615 6043 -1566
rect 6101 -1615 6164 -1566
rect 6229 -1614 6292 -1565
rect 6375 -1633 6438 -1584
rect 3255 -1809 3318 -1760
rect 3255 -1920 3318 -1871
rect 6375 -1740 6438 -1691
rect 6374 -1840 6437 -1791
rect -1162 -2080 1713 -2029
rect 3255 -2031 3318 -1982
rect 6374 -1951 6437 -1902
rect 3255 -2142 3318 -2093
rect 6374 -2062 6437 -2013
rect 3255 -2253 3318 -2204
rect 6374 -2173 6437 -2124
rect 6374 -2284 6437 -2235
rect 3255 -2364 3318 -2315
rect 6374 -2395 6437 -2346
rect 3255 -2475 3318 -2426
rect -236 -2598 -173 -2549
rect -108 -2599 -45 -2550
rect 21 -2598 84 -2549
rect 138 -2599 201 -2550
rect 250 -2600 313 -2551
rect 373 -2598 436 -2549
rect 502 -2597 565 -2548
rect 619 -2598 682 -2549
rect 731 -2599 794 -2550
rect 849 -2599 912 -2550
rect 975 -2598 1038 -2549
rect 1104 -2597 1167 -2548
rect 1221 -2598 1284 -2549
rect 1333 -2599 1396 -2550
rect 1451 -2599 1514 -2550
rect 1574 -2599 1637 -2550
rect 1691 -2599 1754 -2550
rect 1812 -2599 1875 -2550
rect 1934 -2599 1997 -2550
rect 2045 -2600 2108 -2551
rect 2164 -2600 2227 -2551
rect 2276 -2600 2339 -2551
rect 2397 -2600 2460 -2551
rect 2516 -2599 2579 -2550
rect 2631 -2601 2694 -2552
rect 2742 -2599 2805 -2550
rect -250 -2711 -196 -2664
rect -249 -2812 -195 -2765
rect -250 -2909 -196 -2862
rect 2753 -2697 2807 -2650
rect 2754 -2798 2808 -2751
rect -249 -3017 -195 -2970
rect 2753 -2895 2807 -2848
rect 2754 -3003 2808 -2956
rect -249 -3142 -195 -3095
rect 2754 -3128 2808 -3081
rect -248 -3256 -194 -3209
rect 2755 -3242 2809 -3195
rect -247 -3368 -193 -3321
rect -249 -3472 -195 -3425
rect -249 -3576 -195 -3529
rect 2756 -3354 2810 -3307
rect 2754 -3458 2808 -3411
rect -2099 -3654 -1790 -3605
rect -1567 -3649 -838 -3603
rect -251 -3671 -197 -3624
rect 2754 -3562 2808 -3515
rect 2752 -3657 2806 -3610
rect -250 -3780 -196 -3733
rect 2753 -3766 2807 -3719
rect -250 -3884 -196 -3837
rect -252 -3979 -198 -3932
rect -251 -4089 -197 -4042
rect 2753 -3870 2807 -3823
rect 2751 -3965 2805 -3918
rect 2752 -4075 2806 -4028
rect -251 -4193 -197 -4146
rect 2752 -4179 2806 -4132
rect -253 -4288 -199 -4241
rect -250 -4389 -196 -4342
rect 2750 -4274 2804 -4227
rect 2753 -4375 2807 -4328
rect -2099 -4522 -1790 -4473
rect -1567 -4517 -838 -4471
rect -250 -4493 -196 -4446
rect 2753 -4479 2807 -4432
rect -252 -4588 -198 -4541
rect 2751 -4574 2805 -4527
rect -251 -4698 -197 -4651
rect -251 -4802 -197 -4755
rect 2752 -4684 2806 -4637
rect -253 -4897 -199 -4850
rect 2752 -4788 2806 -4741
rect 2750 -4883 2804 -4836
rect -249 -5001 -195 -4954
rect -248 -5111 -194 -5064
rect 2754 -4987 2808 -4940
rect -248 -5215 -194 -5168
rect 2755 -5097 2809 -5050
rect 2755 -5201 2809 -5154
rect -2099 -5381 -1790 -5332
rect -1567 -5376 -838 -5330
rect -239 -5335 -176 -5286
rect -111 -5336 -48 -5287
rect 18 -5335 81 -5286
rect 135 -5336 198 -5287
rect 247 -5337 310 -5288
rect 370 -5335 433 -5286
rect 499 -5334 562 -5285
rect 616 -5335 679 -5286
rect 728 -5336 791 -5287
rect 846 -5336 909 -5287
rect 972 -5335 1035 -5286
rect 1101 -5334 1164 -5285
rect 1218 -5335 1281 -5286
rect 1330 -5336 1393 -5287
rect 1448 -5336 1511 -5287
rect 1571 -5336 1634 -5287
rect 1688 -5336 1751 -5287
rect 1809 -5336 1872 -5287
rect 1931 -5336 1994 -5287
rect 2042 -5337 2105 -5288
rect 2161 -5337 2224 -5288
rect 2273 -5337 2336 -5288
rect 2394 -5337 2457 -5288
rect 2513 -5336 2576 -5287
rect 2628 -5338 2691 -5289
rect 2739 -5336 2802 -5287
rect 3255 -2586 3318 -2537
rect 6374 -2506 6437 -2457
rect 3255 -2697 3318 -2648
rect 6374 -2617 6437 -2568
rect 3255 -2808 3318 -2759
rect 3255 -2919 3318 -2870
rect 6374 -2728 6437 -2679
rect 6374 -2839 6437 -2790
rect 6374 -2950 6437 -2901
rect 3255 -3030 3318 -2981
rect 6374 -3061 6437 -3012
rect 3255 -3141 3318 -3092
rect 3255 -3252 3318 -3203
rect 6374 -3172 6437 -3123
rect 3255 -3363 3318 -3314
rect 6374 -3283 6437 -3234
rect 6374 -3394 6437 -3345
rect 3255 -3474 3318 -3425
rect 3255 -3585 3318 -3536
rect 6374 -3505 6437 -3456
rect 3255 -3696 3318 -3647
rect 6374 -3616 6437 -3567
rect 3255 -3807 3318 -3758
rect 6374 -3727 6437 -3678
rect 3255 -3918 3318 -3869
rect 3255 -4029 3318 -3980
rect 6374 -3838 6437 -3789
rect 6374 -3949 6437 -3900
rect 3255 -4140 3318 -4091
rect 6374 -4060 6437 -4011
rect 3255 -4251 3318 -4202
rect 6374 -4171 6437 -4122
rect 6374 -4282 6437 -4233
rect 3255 -4362 3318 -4313
rect 6374 -4393 6437 -4344
rect 3255 -4473 3318 -4424
rect 3255 -4584 3318 -4535
rect 3255 -4695 3318 -4646
rect 6374 -4504 6437 -4455
rect 6374 -4615 6437 -4566
rect 3255 -4806 3318 -4757
rect 6374 -4726 6437 -4677
rect 3255 -4917 3318 -4868
rect 3255 -5028 3318 -4979
rect 6374 -4837 6437 -4788
rect 6374 -4948 6437 -4899
rect 3255 -5139 3318 -5090
rect 6374 -5059 6437 -5010
rect 3255 -5250 3318 -5201
rect 6374 -5170 6437 -5121
rect 3255 -5361 3318 -5312
rect 6374 -5281 6437 -5232
rect 3255 -5472 3318 -5423
rect 6374 -5392 6437 -5343
rect 6374 -5503 6437 -5454
rect 3255 -5583 3318 -5534
rect 3255 -5694 3318 -5645
rect 6374 -5614 6437 -5565
rect 3255 -5805 3318 -5756
rect 6374 -5725 6437 -5676
rect 3255 -5916 3318 -5867
rect 6374 -5836 6437 -5787
rect 3255 -6027 3318 -5978
rect 6374 -5947 6437 -5898
rect 6374 -6058 6437 -6009
rect 3255 -6138 3318 -6089
rect -2099 -6249 -1790 -6200
rect -1567 -6244 -838 -6198
rect -481 -6249 -172 -6200
rect 51 -6244 780 -6198
rect 1128 -6249 1437 -6200
rect 1660 -6244 2389 -6198
rect 6374 -6169 6437 -6120
rect 3255 -6249 3318 -6200
rect 3255 -6360 3318 -6311
rect 6374 -6280 6437 -6231
rect 3255 -6471 3318 -6422
rect 6374 -6391 6437 -6342
rect 6374 -6502 6437 -6453
rect 3318 -6660 3381 -6611
rect 3439 -6661 3502 -6612
rect 3560 -6661 3623 -6612
rect 3681 -6661 3744 -6612
rect 3802 -6661 3865 -6612
rect 3923 -6661 3986 -6612
rect 4044 -6661 4107 -6612
rect 4165 -6661 4228 -6612
rect 4286 -6661 4349 -6612
rect 4407 -6661 4470 -6612
rect 4528 -6661 4591 -6612
rect 4649 -6661 4712 -6612
rect 4770 -6661 4833 -6612
rect 4891 -6661 4954 -6612
rect 5012 -6661 5075 -6612
rect 5133 -6661 5196 -6612
rect 5254 -6661 5317 -6612
rect 5375 -6661 5438 -6612
rect 5496 -6661 5559 -6612
rect 5617 -6661 5680 -6612
rect 5738 -6661 5801 -6612
rect 5859 -6661 5922 -6612
rect 5980 -6661 6043 -6612
rect 6101 -6661 6164 -6612
<< nsubdiffcont >>
rect -2084 -2965 -1834 -2914
rect -1551 -2955 -839 -2909
rect -2084 -3833 -1834 -3782
rect -1551 -3823 -839 -3777
rect -2084 -4692 -1834 -4641
rect -1551 -4682 -839 -4636
rect -2084 -5560 -1834 -5509
rect -1551 -5550 -839 -5504
rect -466 -5560 -216 -5509
rect 67 -5550 779 -5504
rect 1143 -5560 1393 -5509
rect 1676 -5550 2388 -5504
<< polysilicon >>
rect -1297 1744 1863 1745
rect -1684 1728 -1584 1742
rect -1684 1656 -1658 1728
rect -1598 1656 -1584 1728
rect -1684 1606 -1584 1656
rect -1297 1709 1864 1744
rect -1297 1606 -1197 1709
rect -1093 1606 -993 1650
rect -889 1606 -789 1650
rect -685 1606 -585 1709
rect -481 1606 -381 1709
rect -277 1606 -177 1650
rect -73 1606 27 1650
rect 131 1606 231 1709
rect 335 1606 435 1709
rect 539 1606 639 1650
rect 743 1606 843 1650
rect 947 1606 1047 1709
rect 1151 1606 1251 1709
rect 1764 1650 1864 1709
rect 3524 1782 3634 1795
rect 3524 1769 3542 1782
rect 1355 1606 1455 1650
rect 1559 1606 1659 1650
rect 1763 1606 1863 1650
rect 2144 1606 2244 1650
rect 3119 1710 3223 1724
rect 3119 1647 3146 1710
rect 3209 1647 3223 1710
rect 3119 1608 3223 1647
rect 3480 1705 3542 1769
rect 3619 1705 3634 1782
rect 3480 1688 3634 1705
rect 3738 1769 3843 1783
rect 3738 1692 3752 1769
rect 3829 1760 3843 1769
rect 3829 1692 3879 1760
rect 3480 1608 3535 1688
rect 3738 1678 3879 1692
rect 4161 1695 4247 1709
rect 4161 1684 4175 1695
rect 3820 1608 3879 1678
rect 4012 1647 4175 1684
rect 3120 1606 3223 1608
rect -1684 1303 -1584 1486
rect -1297 1303 -1197 1486
rect -1093 1303 -993 1486
rect -889 1303 -789 1486
rect -685 1303 -585 1486
rect -481 1303 -381 1486
rect -277 1303 -177 1486
rect -73 1303 27 1486
rect 131 1303 231 1486
rect 335 1303 435 1486
rect 539 1303 639 1486
rect 743 1303 843 1486
rect 947 1303 1047 1486
rect 1151 1303 1251 1486
rect 1355 1303 1455 1486
rect 1559 1303 1659 1486
rect 1763 1303 1863 1486
rect 2144 1418 2244 1486
rect 2144 1370 2158 1418
rect 2230 1370 2244 1418
rect 2144 1303 2244 1370
rect 3120 1564 3220 1606
rect 3120 1460 3220 1504
rect 3460 1564 3560 1608
rect 3460 1460 3560 1504
rect 3800 1564 3900 1608
rect 4012 1564 4112 1647
rect 4161 1637 4175 1647
rect 4233 1684 4247 1695
rect 4233 1637 4324 1684
rect 4161 1623 4324 1637
rect 4224 1564 4324 1623
rect 5007 1623 5107 1637
rect 5007 1576 5021 1623
rect 5093 1576 5107 1623
rect 2930 1397 3017 1411
rect 2930 1338 2944 1397
rect 3003 1387 3017 1397
rect 3003 1348 3224 1387
rect 3461 1348 3556 1460
rect 3800 1449 3900 1504
rect 4012 1460 4112 1504
rect 4224 1460 4324 1504
rect 4795 1498 4895 1542
rect 5007 1498 5107 1576
rect 5559 1634 5659 1648
rect 5559 1584 5573 1634
rect 5645 1584 5659 1634
rect 3671 1433 3900 1449
rect 3671 1419 3847 1433
rect 3003 1338 3017 1348
rect 2930 1324 3017 1338
rect 3124 1304 3224 1348
rect 3456 1304 3556 1348
rect 3660 1405 3847 1419
rect 3660 1304 3760 1405
rect 4795 1386 4895 1438
rect 3864 1304 3964 1348
rect 4068 1304 4168 1348
rect 4272 1304 4372 1348
rect 4795 1339 4809 1386
rect 4881 1339 4895 1386
rect -1684 1139 -1584 1183
rect -1297 1141 -1197 1183
rect -1684 1033 -1584 1047
rect -1684 961 -1670 1033
rect -1598 961 -1584 1033
rect -1684 864 -1584 961
rect -1297 1005 -1196 1141
rect -1093 1091 -993 1183
rect -889 1091 -789 1183
rect -685 1139 -585 1183
rect -481 1139 -381 1183
rect -277 1091 -177 1183
rect -73 1091 27 1183
rect 131 1139 231 1183
rect 335 1139 435 1183
rect 539 1091 639 1183
rect 743 1091 843 1183
rect 947 1139 1047 1183
rect 1151 1139 1251 1183
rect 1355 1091 1455 1183
rect 1559 1091 1659 1183
rect 1763 1139 1863 1183
rect 2144 1139 2244 1183
rect 4795 1256 4895 1339
rect 5007 1256 5107 1438
rect 5347 1498 5447 1542
rect 5559 1498 5659 1584
rect 2435 1102 2522 1116
rect 2435 1091 2449 1102
rect -1093 1054 2449 1091
rect 2435 1043 2449 1054
rect 2508 1043 2522 1102
rect 2435 1029 2522 1043
rect 3124 1140 3224 1184
rect 3456 1140 3556 1184
rect 3660 1140 3760 1184
rect 3864 1133 3964 1184
rect 4068 1133 4168 1184
rect 3864 1124 4168 1133
rect 4272 1124 4372 1184
rect 4795 1152 4895 1196
rect 3864 1119 4372 1124
rect 3864 1071 3991 1119
rect -1297 966 1863 1005
rect -1297 864 -1197 966
rect -1093 864 -993 908
rect -889 864 -789 908
rect -685 864 -585 966
rect -481 864 -381 966
rect -277 864 -177 908
rect -73 864 27 908
rect 131 864 231 966
rect 335 864 435 966
rect 539 864 639 908
rect 743 864 843 908
rect 947 864 1047 966
rect 1151 864 1251 966
rect 1355 864 1455 908
rect 1559 864 1659 908
rect 1763 864 1863 966
rect 2144 984 2244 998
rect 2144 935 2158 984
rect 2230 935 2244 984
rect 2144 864 2244 935
rect 3067 1052 3155 1066
rect 3067 992 3081 1052
rect 3141 1044 3155 1052
rect 3977 1058 3991 1071
rect 4052 1068 4372 1119
rect 5007 1145 5107 1196
rect 5347 1256 5447 1438
rect 5559 1256 5659 1438
rect 5899 1498 5999 1542
rect 5347 1152 5447 1196
rect 5007 1082 5241 1145
rect 4052 1058 4066 1068
rect 3977 1044 4066 1058
rect 3141 992 3190 1044
rect 3067 980 3190 992
rect 3067 978 3220 980
rect 3120 936 3220 978
rect 3120 832 3220 876
rect 3460 936 3560 980
rect 3460 824 3560 876
rect 3800 936 3900 980
rect 4012 936 4112 980
rect 3800 832 3900 876
rect 3460 774 3474 824
rect 3546 816 3560 824
rect 3546 774 3706 816
rect 3460 760 3706 774
rect -1684 700 -1584 744
rect -1297 619 -1197 744
rect -1296 324 -1197 619
rect -1093 647 -993 744
rect -889 647 -789 744
rect -685 700 -585 744
rect -481 700 -381 744
rect -277 647 -177 744
rect -73 647 27 744
rect 131 700 231 744
rect 335 700 435 744
rect 539 647 639 744
rect 743 701 843 744
rect 742 700 843 701
rect 947 700 1047 744
rect 1151 700 1251 744
rect 742 647 842 700
rect 1355 647 1455 744
rect 1559 647 1659 744
rect 1763 700 1863 744
rect 2144 700 2244 744
rect 2431 652 2519 666
rect 2431 647 2445 652
rect -1093 597 2445 647
rect 2431 592 2445 597
rect 2505 592 2519 652
rect 2431 578 2519 592
rect 3198 658 3298 702
rect 3402 658 3502 702
rect 3606 658 3706 760
rect 3814 812 3900 832
rect 4012 832 4112 876
rect 4352 936 4452 980
rect 4937 978 5037 1022
rect 5141 978 5241 1082
rect 5351 1124 5447 1152
rect 5559 1152 5659 1196
rect 5899 1256 5999 1438
rect 5559 1124 5647 1152
rect 5899 1143 5999 1196
rect 5351 1039 5647 1124
rect 5351 1022 5445 1039
rect 5345 978 5445 1022
rect 5549 1022 5647 1039
rect 5753 1089 5999 1143
rect 5549 978 5649 1022
rect 5753 978 5853 1089
rect 4012 812 4104 832
rect 4352 827 4452 876
rect 3814 790 4104 812
rect 3814 743 3828 790
rect 3897 743 4104 790
rect 3814 726 4104 743
rect 3814 702 3911 726
rect 4014 702 4104 726
rect 4218 768 4696 827
rect 3810 658 3910 702
rect 4014 658 4114 702
rect 4218 658 4318 768
rect 4637 714 4696 768
rect 4937 809 5037 858
rect 4937 757 4951 809
rect 5023 757 5037 809
rect 4422 658 4522 702
rect 4637 700 4772 714
rect 4637 639 4695 700
rect 4681 637 4695 639
rect 4758 637 4772 700
rect 4937 676 5037 757
rect 5141 676 5241 858
rect 5345 676 5445 858
rect 5549 676 5649 858
rect 5753 676 5853 858
rect 4681 623 4772 637
rect 3198 515 3298 538
rect 3402 515 3502 538
rect 3198 501 3502 515
rect 3198 499 3296 501
rect 3197 445 3296 499
rect 3282 443 3296 445
rect 3354 445 3502 501
rect 3606 494 3706 538
rect 3810 494 3910 538
rect 4014 494 4114 538
rect 4218 494 4318 538
rect 4422 513 4522 538
rect 4422 499 4620 513
rect 4937 512 5037 556
rect 4422 494 4542 499
rect 4461 445 4542 494
rect 3354 443 3368 445
rect 3282 429 3368 443
rect 4528 435 4542 445
rect 4606 435 4620 499
rect 4528 421 4620 435
rect 5141 463 5241 556
rect 5345 512 5445 556
rect 5549 512 5649 556
rect 5753 463 5853 556
rect 3854 414 3955 415
rect 5141 414 5853 463
rect 3854 361 4341 414
rect -1684 288 2244 324
rect -1684 188 -1584 288
rect -1480 188 -1380 232
rect -1276 188 -1176 232
rect -1072 188 -972 288
rect -740 188 -640 288
rect -204 283 764 288
rect -536 188 -436 232
rect -204 188 -104 283
rect 128 188 228 232
rect 332 188 432 232
rect 663 229 764 283
rect 1200 280 2244 288
rect 664 188 764 229
rect 996 188 1096 232
rect 1200 188 1300 280
rect 1532 188 1632 280
rect 1736 188 1836 232
rect 1940 188 2040 232
rect 2144 188 2244 280
rect 3242 359 4341 361
rect 3242 306 3955 359
rect 3043 265 3135 279
rect 3043 201 3057 265
rect 3121 201 3135 265
rect 3043 178 3135 201
rect 3242 178 3343 306
rect 3446 222 3751 258
rect 3038 134 3138 178
rect 3242 134 3342 178
rect 3446 134 3546 222
rect 3650 134 3750 222
rect 3854 178 3955 306
rect 4286 355 4341 359
rect 4286 305 5501 355
rect 4058 290 4158 304
rect 4286 294 4608 305
rect 4058 236 4072 290
rect 4144 236 4158 290
rect 3854 134 3954 178
rect 4058 134 4158 236
rect 4509 142 4608 294
rect 4953 243 5040 257
rect 4953 231 4967 243
rect 4848 195 4967 231
rect 4849 184 4967 195
rect 5026 231 5040 243
rect 5026 230 5160 231
rect 5026 184 5161 230
rect 4849 170 5161 184
rect -1684 -138 -1584 68
rect -1480 -138 -1380 68
rect -1276 -138 -1176 68
rect -1072 -138 -972 68
rect -740 -138 -640 68
rect -536 -138 -436 68
rect -204 27 -104 68
rect 128 27 228 68
rect -204 -4 228 27
rect -204 -42 109 -4
rect 45 -61 109 -42
rect 175 -61 228 -4
rect 45 -79 228 -61
rect -204 -138 -104 -94
rect 128 -138 228 -79
rect 332 -9 432 68
rect 664 24 764 68
rect 332 -81 346 -9
rect 403 -81 432 -9
rect 332 -138 432 -81
rect 664 -138 764 -94
rect 996 -138 1096 68
rect 1200 -138 1300 68
rect 1532 -138 1632 68
rect 1736 -138 1836 68
rect 1940 -138 2040 68
rect 2144 -138 2244 68
rect 4509 98 4609 142
rect 3038 -30 3138 14
rect 3242 -30 3342 14
rect 3446 -30 3546 14
rect 3242 -90 3341 -30
rect 2947 -120 3036 -106
rect 2947 -181 2961 -120
rect 3022 -121 3036 -120
rect 3022 -181 3115 -121
rect 3242 -144 3546 -90
rect 2947 -195 3115 -181
rect 3036 -200 3115 -195
rect -1684 -430 -1584 -258
rect -1480 -353 -1380 -258
rect -1276 -353 -1176 -258
rect -1072 -302 -972 -258
rect -740 -302 -640 -258
rect -536 -353 -436 -258
rect -1480 -354 -436 -353
rect -204 -354 -104 -258
rect 128 -302 228 -258
rect 332 -354 432 -258
rect -1480 -356 432 -354
rect 664 -356 764 -258
rect 996 -352 1096 -258
rect 1200 -302 1300 -258
rect 1532 -302 1632 -258
rect 1736 -352 1836 -258
rect 1940 -352 2040 -258
rect 2144 -302 2244 -258
rect 3038 -244 3138 -200
rect 3242 -244 3342 -200
rect 3446 -244 3546 -144
rect 3650 -94 3750 14
rect 3854 -30 3954 14
rect 4058 -30 4158 14
rect 4509 -60 4609 38
rect 4849 98 4949 170
rect 5061 98 5161 170
rect 4849 -6 4949 38
rect 5061 -6 5161 38
rect 5401 98 5501 305
rect 5613 98 5713 142
rect 5401 -6 5501 38
rect 5613 3 5713 38
rect 3854 -94 3954 -93
rect 3650 -148 3954 -94
rect 4509 -112 4948 -60
rect 3650 -244 3750 -200
rect 3854 -244 3954 -148
rect 4058 -244 4158 -200
rect 4508 -218 4608 -174
rect 2438 -350 2517 -336
rect 2438 -352 2452 -350
rect 996 -356 2452 -352
rect -1480 -399 2452 -356
rect 2438 -401 2452 -399
rect 2503 -401 2517 -350
rect 2438 -415 2517 -401
rect -1684 -502 -1670 -430
rect -1598 -502 -1584 -430
rect -1684 -516 -1584 -502
rect 3038 -523 3138 -364
rect 3242 -523 3342 -364
rect 3446 -411 3546 -364
rect 3650 -411 3750 -364
rect 3446 -460 3750 -411
rect 3446 -523 3546 -460
rect 3650 -523 3750 -460
rect 3854 -523 3954 -364
rect 4058 -409 4158 -364
rect 4058 -459 4072 -409
rect 4144 -459 4158 -409
rect 4058 -523 4158 -459
rect 4508 -468 4608 -278
rect 4848 -218 4948 -112
rect 5095 -67 5152 -6
rect 5612 -36 5713 3
rect 5095 -124 5489 -67
rect 5612 -82 5627 -36
rect 5699 -82 5713 -36
rect 5612 -96 5713 -82
rect 5432 -174 5489 -124
rect 5060 -218 5160 -174
rect 4848 -344 4948 -278
rect 5060 -344 5160 -278
rect 5400 -218 5500 -174
rect 5612 -218 5712 -174
rect 4848 -395 5160 -344
rect 4508 -572 4608 -528
rect 4848 -468 4948 -395
rect 5060 -468 5160 -395
rect 4848 -572 4948 -528
rect 5060 -572 5160 -528
rect 5400 -468 5500 -278
rect 5612 -329 5712 -278
rect 5612 -376 5626 -329
rect 5698 -376 5712 -329
rect 5612 -468 5712 -376
rect 5400 -572 5500 -528
rect 5612 -572 5712 -528
rect 4508 -620 4609 -572
rect 4292 -636 4609 -620
rect 3038 -687 3138 -643
rect 3242 -687 3342 -643
rect 3446 -687 3546 -643
rect 3650 -687 3750 -643
rect -1442 -748 -1197 -734
rect -1684 -824 -1584 -810
rect -1684 -871 -1670 -824
rect -1598 -871 -1584 -824
rect -1442 -820 -1428 -748
rect -1356 -800 -1197 -748
rect -1356 -820 1863 -800
rect -1442 -834 1863 -820
rect -1684 -930 -1584 -871
rect -1297 -836 1863 -834
rect -1297 -930 -1197 -836
rect -1093 -930 -993 -886
rect -889 -930 -789 -886
rect -685 -930 -585 -836
rect -481 -930 -381 -836
rect -277 -930 -177 -886
rect -73 -930 27 -886
rect 131 -930 231 -836
rect 335 -930 435 -836
rect 539 -930 639 -886
rect 743 -930 843 -886
rect 947 -930 1047 -836
rect 1151 -930 1251 -836
rect 1355 -930 1455 -886
rect 1559 -930 1659 -886
rect 1763 -930 1863 -836
rect 2144 -813 2244 -794
rect 2144 -885 2158 -813
rect 2230 -885 2244 -813
rect 2144 -930 2244 -885
rect 3243 -747 3342 -687
rect 3854 -744 3954 -643
rect 4058 -687 4158 -643
rect 4292 -684 4922 -636
rect 4292 -744 4349 -684
rect 3695 -747 4349 -744
rect 3243 -800 4349 -747
rect 4874 -749 4922 -684
rect 5082 -639 5133 -572
rect 5082 -690 5500 -639
rect 3243 -801 3342 -800
rect 3650 -801 4349 -800
rect 4508 -793 4608 -749
rect 3038 -901 3138 -857
rect 3242 -901 3342 -857
rect 3446 -901 3546 -857
rect 3650 -901 3750 -801
rect 3854 -901 3954 -857
rect 4058 -901 4158 -857
rect -1684 -1094 -1584 -1050
rect -1297 -1229 -1197 -1050
rect -1093 -1144 -993 -1050
rect -889 -1144 -789 -1050
rect -685 -1094 -585 -1050
rect -481 -1094 -381 -1050
rect -277 -1094 -177 -1050
rect -278 -1144 -178 -1094
rect -73 -1144 27 -1050
rect 131 -1094 231 -1050
rect 335 -1094 435 -1050
rect 539 -1144 639 -1050
rect 743 -1144 843 -1050
rect 947 -1094 1047 -1050
rect 1151 -1094 1251 -1050
rect 1355 -1094 1455 -1050
rect 1354 -1144 1454 -1094
rect 1559 -1144 1659 -1050
rect 1763 -1094 1863 -1050
rect 2144 -1094 2244 -1050
rect 3038 -1101 3138 -1021
rect 2432 -1132 2521 -1118
rect 2432 -1144 2446 -1132
rect -1093 -1181 2446 -1144
rect 2432 -1193 2446 -1181
rect 2507 -1144 2521 -1132
rect 2507 -1181 2523 -1144
rect 2507 -1193 2521 -1181
rect 2432 -1207 2521 -1193
rect 3036 -1115 3141 -1101
rect 3036 -1192 3050 -1115
rect 3127 -1192 3141 -1115
rect 3036 -1206 3141 -1192
rect 3242 -1181 3342 -1021
rect 3446 -1068 3546 -1021
rect 3650 -1068 3750 -1021
rect 3446 -1130 3750 -1068
rect 3854 -1181 3954 -1021
rect 4058 -1055 4158 -1021
rect 4508 -1049 4608 -853
rect 4848 -793 4948 -749
rect 5060 -793 5160 -749
rect 4848 -914 4948 -853
rect 5060 -914 5160 -853
rect 5400 -793 5500 -690
rect 5612 -793 5712 -749
rect 4848 -928 5160 -914
rect 4848 -976 4959 -928
rect 4945 -988 4959 -976
rect 5019 -976 5160 -928
rect 5019 -988 5033 -976
rect 4945 -1002 5033 -988
rect 4508 -1050 4619 -1049
rect 5400 -1050 5500 -853
rect 5612 -901 5712 -853
rect 5612 -950 5626 -901
rect 5698 -950 5712 -901
rect 5612 -964 5712 -950
rect 4058 -1072 4251 -1055
rect 4058 -1124 4170 -1072
rect 4236 -1124 4251 -1072
rect 4058 -1155 4251 -1124
rect 4508 -1105 5500 -1050
rect -1297 -1269 1863 -1229
rect -1684 -1361 -1584 -1317
rect -1297 -1361 -1197 -1269
rect -1093 -1361 -993 -1317
rect -889 -1361 -789 -1317
rect -685 -1361 -585 -1269
rect -481 -1361 -381 -1269
rect -277 -1361 -177 -1317
rect -73 -1361 27 -1317
rect 131 -1361 231 -1269
rect 335 -1361 435 -1269
rect 539 -1361 639 -1317
rect 743 -1361 843 -1317
rect 947 -1361 1047 -1269
rect 1151 -1361 1251 -1269
rect 1355 -1361 1455 -1317
rect 1559 -1361 1659 -1317
rect 1763 -1361 1863 -1269
rect 3242 -1208 3954 -1181
rect 4508 -1208 4619 -1105
rect 3242 -1235 4619 -1208
rect 2144 -1361 2244 -1317
rect 3854 -1308 4619 -1235
rect 3854 -1330 3954 -1308
rect 3854 -1402 3868 -1330
rect 3933 -1402 3954 -1330
rect 3854 -1416 3954 -1402
rect -1684 -1547 -1584 -1481
rect -1684 -1619 -1670 -1547
rect -1598 -1619 -1584 -1547
rect -1684 -1671 -1584 -1619
rect -1297 -1671 -1197 -1481
rect -1093 -1671 -993 -1481
rect -889 -1671 -789 -1481
rect -685 -1671 -585 -1481
rect -481 -1671 -381 -1481
rect -277 -1671 -177 -1481
rect -73 -1671 27 -1481
rect 131 -1671 231 -1481
rect 335 -1671 435 -1481
rect 539 -1671 639 -1481
rect 743 -1671 843 -1481
rect 947 -1671 1047 -1481
rect 1151 -1671 1251 -1481
rect 1355 -1671 1455 -1481
rect 1559 -1671 1659 -1481
rect 1763 -1671 1863 -1481
rect 2144 -1538 2244 -1481
rect 2144 -1584 2158 -1538
rect 2230 -1584 2244 -1538
rect 2144 -1671 2244 -1584
rect -1684 -1835 -1584 -1791
rect -1297 -1835 -1197 -1791
rect -1093 -1884 -993 -1791
rect -889 -1884 -789 -1791
rect -685 -1835 -585 -1791
rect -481 -1835 -381 -1791
rect -277 -1884 -177 -1791
rect -73 -1884 27 -1791
rect 131 -1835 231 -1791
rect 335 -1835 435 -1791
rect 539 -1884 639 -1791
rect 743 -1884 843 -1791
rect 947 -1835 1047 -1791
rect 1151 -1835 1251 -1791
rect 1355 -1884 1455 -1791
rect 1559 -1884 1659 -1791
rect 1763 -1835 1863 -1791
rect 2144 -1835 2244 -1791
rect 3793 -1707 3893 -1670
rect 3793 -1756 3807 -1707
rect 3879 -1734 3893 -1707
rect 3879 -1756 5834 -1734
rect 2437 -1873 2523 -1859
rect 2437 -1884 2451 -1873
rect -1093 -1920 2451 -1884
rect 2437 -1931 2451 -1920
rect 2509 -1931 2523 -1873
rect 2437 -1945 2523 -1931
rect 3589 -1807 3689 -1770
rect 3589 -1856 3603 -1807
rect 3675 -1856 3689 -1807
rect 3589 -1906 3689 -1856
rect 3793 -1814 5834 -1756
rect 3793 -1906 3893 -1814
rect 4125 -1906 4225 -1862
rect 4329 -1906 4429 -1862
rect 4661 -1906 4761 -1814
rect 4865 -1906 4965 -1814
rect 5197 -1906 5297 -1862
rect 5401 -1906 5501 -1862
rect 5733 -1906 5833 -1814
rect 5937 -1819 6037 -1783
rect 5937 -1869 5951 -1819
rect 6023 -1869 6037 -1819
rect 5937 -1906 6037 -1869
rect 3589 -2070 3689 -2026
rect 3793 -2070 3893 -2026
rect 4125 -2112 4225 -2026
rect 4329 -2112 4429 -2026
rect 4661 -2070 4761 -2026
rect 4865 -2070 4965 -2026
rect 4125 -2122 4429 -2112
rect 5197 -2122 5297 -2026
rect 5401 -2122 5501 -2026
rect 5733 -2070 5833 -2026
rect 5937 -2070 6037 -2026
rect 3793 -2126 5833 -2122
rect 3793 -2184 4256 -2126
rect 4314 -2184 5833 -2126
rect 3793 -2188 5833 -2184
rect 3589 -2290 3689 -2246
rect 3793 -2290 3893 -2188
rect 4242 -2198 4328 -2188
rect 4125 -2290 4225 -2246
rect 4329 -2290 4429 -2246
rect 4661 -2290 4761 -2188
rect 4865 -2290 4965 -2188
rect 5197 -2290 5297 -2246
rect 5401 -2290 5501 -2246
rect 5733 -2290 5833 -2188
rect 5937 -2290 6037 -2246
rect 228 -2790 2266 -2690
rect 228 -2845 325 -2790
rect 21 -2889 121 -2845
rect 225 -2889 325 -2845
rect 557 -2889 657 -2845
rect 761 -2889 861 -2845
rect 1093 -2889 1193 -2790
rect 1297 -2889 1397 -2790
rect 2166 -2845 2266 -2790
rect 1629 -2889 1729 -2845
rect 1833 -2889 1933 -2845
rect 2165 -2848 2266 -2845
rect 2165 -2889 2265 -2848
rect 2369 -2889 2469 -2845
rect -1970 -3062 -1914 -3018
rect -732 -3019 -596 -3005
rect -732 -3025 -719 -3019
rect -1430 -3111 -1374 -3067
rect -1018 -3077 -719 -3025
rect -1970 -3224 -1914 -3162
rect -1430 -3210 -1374 -3155
rect -1018 -3111 -962 -3077
rect -732 -3079 -719 -3077
rect -656 -3079 -596 -3019
rect -732 -3092 -596 -3079
rect -1018 -3199 -962 -3155
rect 21 -3051 121 -3009
rect 21 -3100 35 -3051
rect 107 -3100 121 -3051
rect 225 -3053 325 -3009
rect 557 -3050 657 -3009
rect 761 -3050 861 -3009
rect 21 -3173 121 -3100
rect 228 -3129 325 -3053
rect 225 -3173 325 -3129
rect 556 -3130 861 -3050
rect 557 -3173 657 -3130
rect 761 -3173 861 -3130
rect 1093 -3173 1193 -3009
rect 1297 -3173 1397 -3009
rect 1629 -3050 1729 -3009
rect 1833 -3050 1933 -3009
rect 1628 -3130 1933 -3050
rect 1629 -3173 1729 -3130
rect 1833 -3173 1933 -3130
rect 2165 -3173 2265 -3009
rect 2369 -3063 2469 -3009
rect 2369 -3111 2383 -3063
rect 2455 -3111 2469 -3063
rect 2369 -3173 2469 -3111
rect -2029 -3238 -1914 -3224
rect -2029 -3297 -2015 -3238
rect -1952 -3297 -1914 -3238
rect -1441 -3223 -1352 -3210
rect -1441 -3283 -1428 -3223
rect -1365 -3283 -1352 -3223
rect -1441 -3297 -1352 -3283
rect -2029 -3311 -1914 -3297
rect -1970 -3411 -1914 -3311
rect 21 -3337 121 -3293
rect -1731 -3382 -1642 -3368
rect -1731 -3442 -1718 -3382
rect -1655 -3442 -1642 -3382
rect -1731 -3455 -1642 -3442
rect -1970 -3505 -1914 -3461
rect -1693 -3504 -1648 -3455
rect -1492 -3416 -1436 -3372
rect -1492 -3504 -1436 -3460
rect -956 -3416 -900 -3372
rect -1693 -3551 -1436 -3504
rect -956 -3495 -900 -3460
rect -730 -3477 -641 -3463
rect -730 -3495 -717 -3477
rect -956 -3537 -717 -3495
rect -654 -3537 -641 -3477
rect -956 -3541 -641 -3537
rect -730 -3550 -641 -3541
rect 225 -3529 325 -3293
rect 557 -3337 657 -3293
rect 761 -3385 861 -3293
rect 1093 -3337 1193 -3293
rect 1297 -3337 1397 -3293
rect 1629 -3337 1729 -3293
rect 1833 -3337 1933 -3293
rect 2165 -3337 2265 -3293
rect 2369 -3337 2469 -3293
rect 1629 -3385 1728 -3337
rect 760 -3453 1728 -3385
rect 1836 -3351 1933 -3337
rect 1836 -3365 2021 -3351
rect 1836 -3419 1938 -3365
rect 2007 -3419 2021 -3365
rect 1836 -3448 2021 -3419
rect 1044 -3529 1125 -3528
rect 21 -3547 121 -3533
rect 21 -3595 35 -3547
rect 107 -3595 121 -3547
rect 21 -3705 121 -3595
rect 225 -3543 1754 -3529
rect 225 -3590 851 -3543
rect 923 -3590 1754 -3543
rect 225 -3607 1754 -3590
rect 1857 -3563 1956 -3549
rect 225 -3705 325 -3607
rect 429 -3705 529 -3661
rect 633 -3705 733 -3661
rect 837 -3705 937 -3607
rect 1041 -3705 1141 -3607
rect 1245 -3705 1345 -3661
rect 1449 -3705 1549 -3661
rect 1653 -3705 1753 -3607
rect 1857 -3610 1871 -3563
rect 1942 -3610 1956 -3563
rect 1857 -3661 1956 -3610
rect 2189 -3568 2289 -3554
rect 2189 -3615 2203 -3568
rect 2275 -3615 2289 -3568
rect 1857 -3705 1957 -3661
rect 2189 -3705 2289 -3615
rect 2393 -3568 2493 -3554
rect 2393 -3615 2407 -3568
rect 2479 -3615 2493 -3568
rect 2393 -3705 2493 -3615
rect -1970 -3930 -1914 -3886
rect -732 -3887 -643 -3873
rect -732 -3893 -719 -3887
rect -1430 -3979 -1374 -3935
rect -1018 -3945 -719 -3893
rect -1970 -4092 -1914 -4030
rect -1430 -4078 -1374 -4023
rect -1018 -3979 -962 -3945
rect -732 -3947 -719 -3945
rect -656 -3947 -643 -3887
rect -732 -3960 -643 -3947
rect 21 -3869 121 -3825
rect 225 -3869 325 -3825
rect 429 -3867 529 -3825
rect 428 -3869 529 -3867
rect 428 -3913 528 -3869
rect 428 -3930 442 -3913
rect -1018 -4067 -962 -4023
rect -2029 -4106 -1914 -4092
rect -2029 -4165 -2015 -4106
rect -1952 -4165 -1914 -4106
rect -1441 -4091 -1352 -4078
rect -1441 -4151 -1428 -4091
rect -1365 -4151 -1352 -4091
rect -1441 -4165 -1352 -4151
rect 226 -3960 442 -3930
rect 514 -3930 528 -3913
rect 633 -3930 733 -3825
rect 837 -3869 937 -3825
rect 1041 -3869 1141 -3825
rect 1245 -3930 1345 -3825
rect 1449 -3930 1549 -3825
rect 1653 -3869 1753 -3825
rect 1857 -3869 1957 -3825
rect 2189 -3869 2289 -3825
rect 2393 -3869 2493 -3825
rect 514 -3960 1753 -3930
rect 226 -3996 1753 -3960
rect 226 -4050 325 -3996
rect 21 -4094 121 -4050
rect 225 -4094 325 -4050
rect 429 -4094 529 -4050
rect 633 -4094 733 -4050
rect 837 -4094 937 -3996
rect 1041 -4094 1141 -3996
rect 1245 -4094 1345 -4050
rect 1449 -4094 1549 -4050
rect 1653 -4094 1753 -3996
rect 1857 -4094 1957 -4050
rect 2189 -4094 2289 -4050
rect 2393 -4094 2493 -4050
rect -2029 -4179 -1914 -4165
rect -1970 -4279 -1914 -4179
rect -1731 -4250 -1642 -4236
rect -1731 -4310 -1718 -4250
rect -1655 -4310 -1642 -4250
rect -1731 -4323 -1642 -4310
rect -1970 -4373 -1914 -4329
rect -1693 -4372 -1648 -4323
rect -1492 -4284 -1436 -4240
rect -1492 -4372 -1436 -4328
rect -956 -4284 -900 -4240
rect -1693 -4419 -1436 -4372
rect -956 -4363 -900 -4328
rect -730 -4345 -641 -4331
rect -730 -4363 -717 -4345
rect -956 -4405 -717 -4363
rect -654 -4405 -641 -4345
rect -956 -4409 -641 -4405
rect -730 -4418 -641 -4409
rect 21 -4266 121 -4214
rect 21 -4315 35 -4266
rect 107 -4315 121 -4266
rect 21 -4389 121 -4315
rect 225 -4389 325 -4214
rect 429 -4263 529 -4214
rect 633 -4263 733 -4214
rect 429 -4346 733 -4263
rect 429 -4389 529 -4346
rect 633 -4389 733 -4346
rect 837 -4278 937 -4214
rect 1041 -4278 1141 -4214
rect 837 -4361 1141 -4278
rect 837 -4389 937 -4361
rect 1041 -4389 1141 -4361
rect 1245 -4258 1345 -4214
rect 1449 -4258 1549 -4214
rect 1245 -4339 1553 -4258
rect 1245 -4389 1345 -4339
rect 1449 -4389 1549 -4339
rect 1653 -4389 1753 -4214
rect 1857 -4265 1957 -4214
rect 1857 -4311 1871 -4265
rect 1943 -4311 1957 -4265
rect 1857 -4389 1957 -4311
rect 2189 -4274 2289 -4214
rect 2189 -4322 2203 -4274
rect 2275 -4322 2289 -4274
rect 2189 -4389 2289 -4322
rect 2393 -4271 2493 -4214
rect 2393 -4318 2407 -4271
rect 2479 -4318 2493 -4271
rect 2393 -4389 2493 -4318
rect 21 -4553 121 -4509
rect 225 -4553 325 -4509
rect 429 -4553 529 -4509
rect 633 -4601 733 -4509
rect 837 -4553 937 -4509
rect 1041 -4553 1141 -4509
rect 1245 -4601 1345 -4509
rect 1449 -4553 1549 -4509
rect 1653 -4553 1753 -4509
rect 1857 -4553 1957 -4509
rect 2189 -4553 2289 -4509
rect 2393 -4553 2493 -4509
rect -1970 -4789 -1914 -4745
rect -732 -4746 -643 -4732
rect -732 -4752 -719 -4746
rect -1430 -4838 -1374 -4794
rect -1018 -4804 -719 -4752
rect -1970 -4951 -1914 -4889
rect -1430 -4937 -1374 -4882
rect -1018 -4838 -962 -4804
rect -732 -4806 -719 -4804
rect -656 -4806 -643 -4746
rect -732 -4819 -643 -4806
rect 165 -4615 1753 -4601
rect 165 -4687 179 -4615
rect 241 -4663 851 -4615
rect 923 -4663 1753 -4615
rect 241 -4669 1753 -4663
rect 241 -4687 325 -4669
rect 165 -4701 325 -4687
rect 21 -4774 121 -4730
rect 225 -4774 325 -4701
rect 429 -4774 529 -4730
rect 633 -4774 733 -4730
rect 837 -4774 937 -4669
rect 1041 -4774 1141 -4669
rect 1245 -4774 1345 -4730
rect 1449 -4774 1549 -4730
rect 1653 -4774 1753 -4669
rect 1857 -4774 1957 -4730
rect 2189 -4774 2289 -4730
rect 2393 -4774 2493 -4730
rect -1018 -4926 -962 -4882
rect -2029 -4965 -1914 -4951
rect -2029 -5024 -2015 -4965
rect -1952 -5024 -1914 -4965
rect -1441 -4950 -1352 -4937
rect -1441 -5010 -1428 -4950
rect -1365 -5010 -1352 -4950
rect -1441 -5024 -1352 -5010
rect -2029 -5038 -1914 -5024
rect -1970 -5138 -1914 -5038
rect -1731 -5109 -1642 -5095
rect -1731 -5169 -1718 -5109
rect -1655 -5169 -1642 -5109
rect -1731 -5182 -1642 -5169
rect -1970 -5232 -1914 -5188
rect -1693 -5231 -1648 -5182
rect -1492 -5143 -1436 -5099
rect -1492 -5231 -1436 -5187
rect -956 -5143 -900 -5099
rect 21 -4983 121 -4894
rect 225 -4938 325 -4894
rect 429 -4966 529 -4894
rect 21 -5029 35 -4983
rect 107 -5029 121 -4983
rect 21 -5069 121 -5029
rect 373 -4980 529 -4966
rect 373 -5029 387 -4980
rect 459 -4989 529 -4980
rect 633 -4989 733 -4894
rect 837 -4938 937 -4894
rect 1041 -4938 1141 -4894
rect 1245 -4989 1345 -4894
rect 1449 -4980 1549 -4894
rect 1653 -4938 1753 -4894
rect 1449 -4989 1487 -4980
rect 459 -5029 1487 -4989
rect 373 -5052 1487 -5029
rect 1535 -5052 1549 -4980
rect 1857 -4953 1957 -4894
rect 1857 -4999 1871 -4953
rect 1943 -4999 1957 -4953
rect 1857 -5039 1957 -4999
rect 2189 -4953 2289 -4894
rect 2189 -4999 2203 -4953
rect 2275 -4999 2289 -4953
rect 2189 -5039 2289 -4999
rect 2393 -4953 2493 -4894
rect 2393 -5003 2407 -4953
rect 2479 -5003 2493 -4953
rect 2393 -5039 2493 -5003
rect 373 -5066 1549 -5052
rect -1693 -5278 -1436 -5231
rect -956 -5222 -900 -5187
rect -730 -5204 -641 -5190
rect -730 -5222 -717 -5204
rect -956 -5264 -717 -5222
rect -654 -5264 -641 -5204
rect -956 -5268 -641 -5264
rect -730 -5277 -641 -5268
rect 3589 -2469 3689 -2410
rect 3589 -2518 3603 -2469
rect 3675 -2518 3689 -2469
rect 3589 -2580 3689 -2518
rect 3793 -2580 3893 -2410
rect 4125 -2450 4225 -2410
rect 4329 -2450 4429 -2410
rect 4125 -2528 4429 -2450
rect 4125 -2580 4225 -2528
rect 4329 -2580 4429 -2528
rect 4661 -2580 4761 -2410
rect 4865 -2580 4965 -2410
rect 5197 -2451 5297 -2410
rect 5401 -2451 5501 -2410
rect 5197 -2526 5501 -2451
rect 5197 -2580 5297 -2526
rect 5401 -2580 5501 -2526
rect 5733 -2580 5833 -2410
rect 5937 -2449 6037 -2410
rect 5937 -2499 5951 -2449
rect 6023 -2499 6037 -2449
rect 5937 -2580 6037 -2499
rect 3589 -2744 3689 -2700
rect 3793 -2744 3893 -2700
rect 4125 -2744 4225 -2700
rect 3741 -2796 3893 -2795
rect 4329 -2796 4429 -2700
rect 4661 -2744 4761 -2700
rect 4865 -2744 4965 -2700
rect 5197 -2796 5297 -2700
rect 5401 -2744 5501 -2700
rect 5733 -2744 5833 -2700
rect 5937 -2744 6037 -2700
rect 3741 -2809 5833 -2796
rect 3741 -2860 3755 -2809
rect 3826 -2860 5833 -2809
rect 3741 -2867 5833 -2860
rect 3741 -2894 3893 -2867
rect 3589 -2964 3689 -2920
rect 3793 -2964 3893 -2894
rect 4125 -2964 4225 -2920
rect 4329 -2964 4429 -2920
rect 4660 -2928 4761 -2867
rect 4661 -2964 4761 -2928
rect 4864 -2934 4965 -2867
rect 4865 -2964 4965 -2934
rect 5197 -2964 5297 -2920
rect 5401 -2964 5501 -2920
rect 5733 -2964 5833 -2867
rect 5937 -2964 6037 -2920
rect 3589 -3118 3689 -3084
rect 3589 -3166 3603 -3118
rect 3675 -3166 3689 -3118
rect 3793 -3128 3893 -3084
rect 3589 -3204 3689 -3166
rect 4125 -3176 4225 -3084
rect 4329 -3176 4429 -3084
rect 4661 -3128 4761 -3084
rect 4865 -3128 4965 -3084
rect 5197 -3176 5297 -3084
rect 5401 -3176 5501 -3084
rect 5733 -3128 5833 -3084
rect 4125 -3192 5501 -3176
rect 4125 -3249 4245 -3192
rect 4305 -3249 5501 -3192
rect 5937 -3141 6037 -3084
rect 5937 -3187 5951 -3141
rect 6023 -3187 6037 -3141
rect 5937 -3201 6037 -3187
rect 4125 -3263 5501 -3249
rect 3561 -3422 3660 -3408
rect 3561 -3492 3576 -3422
rect 3646 -3445 3660 -3422
rect 3646 -3492 5321 -3445
rect 3561 -3506 5321 -3492
rect 3589 -3598 3689 -3554
rect 3793 -3598 3893 -3506
rect 3997 -3598 4097 -3554
rect 4201 -3598 4301 -3554
rect 4405 -3598 4505 -3506
rect 4609 -3598 4709 -3506
rect 4813 -3598 4913 -3554
rect 5017 -3598 5117 -3554
rect 5221 -3598 5321 -3506
rect 5425 -3491 5525 -3473
rect 5425 -3541 5439 -3491
rect 5511 -3541 5525 -3491
rect 5425 -3598 5525 -3541
rect 5757 -3493 6060 -3479
rect 5757 -3540 5771 -3493
rect 5843 -3540 6060 -3493
rect 5757 -3554 6060 -3540
rect 5757 -3555 6061 -3554
rect 5757 -3598 5857 -3555
rect 5961 -3598 6061 -3555
rect 3589 -3748 3689 -3718
rect 3505 -3762 3689 -3748
rect 3793 -3762 3893 -3718
rect 3505 -3809 3519 -3762
rect 3590 -3809 3689 -3762
rect 3505 -3847 3689 -3809
rect 3997 -3812 4097 -3718
rect 4201 -3812 4301 -3718
rect 4405 -3762 4505 -3718
rect 4609 -3762 4709 -3718
rect 4813 -3812 4913 -3718
rect 5017 -3812 5117 -3718
rect 5221 -3762 5321 -3718
rect 5425 -3762 5525 -3718
rect 5757 -3762 5857 -3718
rect 5961 -3762 6061 -3718
rect 5560 -3812 5658 -3799
rect 3793 -3813 5658 -3812
rect 3793 -3883 5574 -3813
rect 5644 -3883 5658 -3813
rect 3793 -3885 5658 -3883
rect 3589 -3987 3689 -3943
rect 3793 -3987 3893 -3885
rect 3997 -3987 4097 -3943
rect 4201 -3987 4301 -3943
rect 4405 -3987 4505 -3885
rect 4609 -3987 4709 -3885
rect 4813 -3987 4913 -3943
rect 5017 -3987 5117 -3943
rect 5221 -3987 5321 -3885
rect 5560 -3897 5658 -3885
rect 5425 -3987 5525 -3943
rect 5757 -3987 5857 -3943
rect 5961 -3987 6061 -3943
rect 3589 -4166 3689 -4107
rect 3589 -4216 3603 -4166
rect 3675 -4216 3689 -4166
rect 3589 -4282 3689 -4216
rect 3793 -4282 3893 -4107
rect 3997 -4154 4097 -4107
rect 4201 -4154 4301 -4107
rect 3997 -4234 4301 -4154
rect 3997 -4282 4097 -4234
rect 4201 -4282 4301 -4234
rect 4405 -4151 4505 -4107
rect 4609 -4151 4709 -4107
rect 4405 -4236 4709 -4151
rect 4405 -4282 4505 -4236
rect 4609 -4282 4709 -4236
rect 4813 -4154 4913 -4107
rect 5017 -4154 5117 -4107
rect 4813 -4238 5117 -4154
rect 4813 -4282 4913 -4238
rect 5017 -4282 5117 -4238
rect 5221 -4282 5321 -4107
rect 5425 -4152 5525 -4107
rect 5425 -4203 5439 -4152
rect 5511 -4203 5525 -4152
rect 5425 -4282 5525 -4203
rect 5757 -4166 5857 -4107
rect 5757 -4216 5771 -4166
rect 5843 -4216 5857 -4166
rect 5757 -4282 5857 -4216
rect 5961 -4164 6061 -4107
rect 5961 -4211 5975 -4164
rect 6047 -4211 6061 -4164
rect 5961 -4282 6061 -4211
rect 3589 -4446 3689 -4402
rect 3793 -4446 3893 -4402
rect 3997 -4446 4097 -4402
rect 3462 -4494 3551 -4483
rect 4201 -4494 4301 -4402
rect 4405 -4446 4505 -4402
rect 4609 -4446 4709 -4402
rect 4813 -4494 4913 -4402
rect 5017 -4446 5117 -4402
rect 5221 -4446 5321 -4402
rect 5425 -4446 5525 -4402
rect 5757 -4446 5857 -4402
rect 5961 -4446 6061 -4402
rect 3462 -4497 5321 -4494
rect 3462 -4558 3476 -4497
rect 3537 -4558 5321 -4497
rect 3462 -4562 5321 -4558
rect 3462 -4572 3551 -4562
rect 3589 -4667 3689 -4623
rect 3793 -4667 3893 -4562
rect 3997 -4667 4097 -4623
rect 4201 -4667 4301 -4623
rect 4405 -4667 4505 -4562
rect 4609 -4667 4709 -4562
rect 4813 -4667 4913 -4623
rect 5017 -4667 5117 -4623
rect 5221 -4667 5321 -4562
rect 5425 -4667 5525 -4623
rect 5757 -4667 5857 -4623
rect 5961 -4667 6061 -4623
rect 3589 -4831 3689 -4787
rect 3793 -4831 3893 -4787
rect 3589 -4858 3688 -4831
rect 3589 -4914 3603 -4858
rect 3674 -4914 3688 -4858
rect 3589 -4950 3688 -4914
rect 3793 -4950 3892 -4831
rect 3997 -4844 4097 -4787
rect 4201 -4844 4301 -4787
rect 3997 -4943 4301 -4844
rect 3589 -4994 3689 -4950
rect 3793 -4994 3893 -4950
rect 3997 -4994 4097 -4943
rect 4201 -4994 4301 -4943
rect 4405 -4833 4505 -4787
rect 4609 -4833 4709 -4787
rect 4405 -4926 4709 -4833
rect 4405 -4994 4505 -4926
rect 4609 -4994 4709 -4926
rect 4813 -4844 4913 -4787
rect 5017 -4844 5117 -4787
rect 4813 -4933 5117 -4844
rect 4813 -4994 4913 -4933
rect 5017 -4994 5117 -4933
rect 5221 -4994 5321 -4787
rect 5425 -4856 5525 -4787
rect 5425 -4907 5439 -4856
rect 5511 -4907 5525 -4856
rect 5425 -4994 5525 -4907
rect 5757 -4859 5857 -4787
rect 5757 -4908 5771 -4859
rect 5843 -4908 5857 -4859
rect 5757 -4994 5857 -4908
rect 5961 -4856 6061 -4787
rect 5961 -4903 5975 -4856
rect 6047 -4903 6061 -4856
rect 5961 -4994 6061 -4903
rect 3589 -5158 3689 -5114
rect 3793 -5158 3893 -5114
rect 3997 -5158 4097 -5114
rect 4201 -5208 4301 -5114
rect 4405 -5158 4505 -5114
rect 4609 -5158 4709 -5114
rect 4813 -5208 4913 -5114
rect 5017 -5158 5117 -5114
rect 5221 -5158 5321 -5114
rect 5425 -5158 5525 -5114
rect 5757 -5158 5857 -5114
rect 5961 -5158 6061 -5114
rect 5562 -5208 5658 -5194
rect 3793 -5276 5576 -5208
rect 5644 -5276 5658 -5208
rect 3793 -5339 3892 -5276
rect 3589 -5383 3689 -5339
rect 3793 -5383 3893 -5339
rect 3997 -5383 4097 -5339
rect 4201 -5383 4301 -5339
rect 4405 -5383 4505 -5276
rect 4609 -5383 4709 -5276
rect 4813 -5383 4913 -5339
rect 5017 -5383 5117 -5339
rect 5221 -5383 5321 -5276
rect 5562 -5290 5658 -5276
rect 5425 -5383 5525 -5339
rect 5757 -5383 5857 -5339
rect 5961 -5383 6061 -5339
rect -1970 -5657 -1914 -5613
rect -732 -5614 -643 -5600
rect -732 -5620 -719 -5614
rect -1430 -5706 -1374 -5662
rect -1018 -5672 -719 -5620
rect -1970 -5819 -1914 -5757
rect -1430 -5805 -1374 -5750
rect -1018 -5706 -962 -5672
rect -732 -5674 -719 -5672
rect -656 -5674 -643 -5614
rect -352 -5657 -296 -5613
rect 886 -5614 975 -5600
rect 886 -5620 899 -5614
rect -732 -5687 -643 -5674
rect -1018 -5794 -962 -5750
rect 188 -5706 244 -5662
rect 600 -5672 899 -5620
rect -2029 -5833 -1914 -5819
rect -2029 -5892 -2015 -5833
rect -1952 -5892 -1914 -5833
rect -1441 -5818 -1352 -5805
rect -1441 -5878 -1428 -5818
rect -1365 -5878 -1352 -5818
rect -352 -5819 -296 -5757
rect 188 -5805 244 -5750
rect 600 -5706 656 -5672
rect 886 -5674 899 -5672
rect 962 -5674 975 -5614
rect 1257 -5657 1313 -5613
rect 2495 -5614 2584 -5600
rect 2495 -5620 2508 -5614
rect 886 -5687 975 -5674
rect 600 -5794 656 -5750
rect 1797 -5706 1853 -5662
rect 2209 -5672 2508 -5620
rect -1441 -5892 -1352 -5878
rect -411 -5833 -296 -5819
rect -411 -5892 -397 -5833
rect -334 -5892 -296 -5833
rect 177 -5818 266 -5805
rect 177 -5878 190 -5818
rect 253 -5878 266 -5818
rect 1257 -5819 1313 -5757
rect 1797 -5805 1853 -5750
rect 2209 -5706 2265 -5672
rect 2495 -5674 2508 -5672
rect 2571 -5674 2584 -5614
rect 2495 -5687 2584 -5674
rect 2209 -5794 2265 -5750
rect 3589 -5547 3689 -5503
rect 3793 -5547 3893 -5503
rect 3997 -5542 4097 -5503
rect 4201 -5542 4301 -5503
rect 3589 -5554 3688 -5547
rect 3589 -5604 3603 -5554
rect 3674 -5604 3688 -5554
rect 3589 -5634 3688 -5604
rect 3793 -5634 3892 -5547
rect 3997 -5616 4301 -5542
rect 3589 -5678 3689 -5634
rect 3793 -5678 3893 -5634
rect 3997 -5678 4097 -5616
rect 4201 -5678 4301 -5616
rect 4405 -5558 4505 -5503
rect 4609 -5558 4709 -5503
rect 4405 -5631 4709 -5558
rect 4405 -5678 4505 -5631
rect 4609 -5678 4709 -5631
rect 4813 -5553 4913 -5503
rect 5017 -5553 5117 -5503
rect 4813 -5634 5117 -5553
rect 4813 -5678 4913 -5634
rect 5017 -5678 5117 -5634
rect 5221 -5678 5321 -5503
rect 5425 -5559 5525 -5503
rect 5425 -5605 5439 -5559
rect 5511 -5605 5525 -5559
rect 5425 -5678 5525 -5605
rect 5757 -5552 5857 -5503
rect 5757 -5602 5771 -5552
rect 5843 -5602 5857 -5552
rect 5757 -5678 5857 -5602
rect 5961 -5551 6061 -5503
rect 5961 -5604 5975 -5551
rect 6047 -5604 6061 -5551
rect 5961 -5678 6061 -5604
rect 177 -5892 266 -5878
rect 1198 -5833 1313 -5819
rect 1198 -5892 1212 -5833
rect 1275 -5892 1313 -5833
rect 1786 -5818 1875 -5805
rect 1786 -5878 1799 -5818
rect 1862 -5878 1875 -5818
rect 1786 -5892 1875 -5878
rect 3589 -5842 3689 -5798
rect 3793 -5842 3893 -5798
rect 3997 -5842 4097 -5798
rect -2029 -5906 -1914 -5892
rect -411 -5906 -296 -5892
rect 1198 -5906 1313 -5892
rect -1970 -6006 -1914 -5906
rect -1731 -5977 -1642 -5963
rect -1731 -6037 -1718 -5977
rect -1655 -6037 -1642 -5977
rect -1731 -6050 -1642 -6037
rect -1970 -6100 -1914 -6056
rect -1693 -6099 -1648 -6050
rect -1492 -6011 -1436 -5967
rect -1492 -6099 -1436 -6055
rect -956 -6011 -900 -5967
rect -1693 -6146 -1436 -6099
rect -956 -6090 -900 -6055
rect -352 -6006 -296 -5906
rect -113 -5977 -24 -5963
rect -113 -6037 -100 -5977
rect -37 -6037 -24 -5977
rect -113 -6050 -24 -6037
rect -730 -6072 -641 -6058
rect -730 -6090 -717 -6072
rect -956 -6132 -717 -6090
rect -654 -6132 -641 -6072
rect -352 -6100 -296 -6056
rect -75 -6099 -30 -6050
rect 126 -6011 182 -5967
rect 126 -6099 182 -6055
rect 662 -6011 718 -5967
rect -956 -6136 -641 -6132
rect -730 -6145 -641 -6136
rect -75 -6146 182 -6099
rect 662 -6090 718 -6055
rect 1257 -6006 1313 -5906
rect 1496 -5977 1585 -5963
rect 1496 -6037 1509 -5977
rect 1572 -6037 1585 -5977
rect 1496 -6050 1585 -6037
rect 888 -6072 977 -6058
rect 888 -6090 901 -6072
rect 662 -6132 901 -6090
rect 964 -6132 977 -6072
rect 1257 -6100 1313 -6056
rect 1534 -6099 1579 -6050
rect 1735 -6011 1791 -5967
rect 1735 -6099 1791 -6055
rect 2271 -6011 2327 -5967
rect 3456 -5889 3544 -5875
rect 3456 -5949 3470 -5889
rect 3530 -5891 3544 -5889
rect 4201 -5891 4301 -5798
rect 4405 -5842 4505 -5798
rect 4609 -5842 4709 -5798
rect 4813 -5891 4913 -5798
rect 5017 -5842 5117 -5798
rect 5221 -5842 5321 -5798
rect 5425 -5842 5525 -5798
rect 5757 -5842 5857 -5798
rect 5961 -5842 6061 -5798
rect 3530 -5948 5321 -5891
rect 5515 -5925 5602 -5915
rect 3530 -5949 3544 -5948
rect 3456 -5963 3544 -5949
rect 662 -6136 977 -6132
rect 888 -6145 977 -6136
rect 1534 -6146 1791 -6099
rect 2271 -6090 2327 -6055
rect 2497 -6072 2586 -6058
rect 2497 -6090 2510 -6072
rect 2271 -6132 2510 -6090
rect 2573 -6132 2586 -6072
rect 2271 -6136 2586 -6132
rect 2497 -6145 2586 -6136
rect 3589 -6063 3689 -6019
rect 3793 -6063 3893 -5948
rect 3997 -6063 4097 -6019
rect 4201 -6063 4301 -6019
rect 4405 -6063 4505 -5948
rect 4609 -6063 4709 -5948
rect 4813 -6063 4913 -6019
rect 5017 -6063 5117 -6019
rect 5221 -6063 5321 -5948
rect 5424 -5929 5602 -5925
rect 5424 -5988 5529 -5929
rect 5588 -5988 5602 -5929
rect 5424 -5992 5602 -5988
rect 5425 -6002 5602 -5992
rect 5755 -5962 6061 -5948
rect 5425 -6019 5526 -6002
rect 5755 -6011 5975 -5962
rect 6047 -6011 6061 -5962
rect 5755 -6018 6061 -6011
rect 5425 -6063 5525 -6019
rect 5757 -6063 5857 -6018
rect 5961 -6063 6061 -6018
rect 3589 -6228 3689 -6183
rect 3793 -6227 3893 -6183
rect 3589 -6280 3603 -6228
rect 3675 -6280 3689 -6228
rect 3589 -6314 3689 -6280
rect 3997 -6282 4097 -6183
rect 4201 -6282 4301 -6183
rect 4405 -6227 4505 -6183
rect 4609 -6227 4709 -6183
rect 4813 -6282 4913 -6183
rect 5017 -6282 5117 -6183
rect 5221 -6227 5321 -6183
rect 5425 -6227 5525 -6183
rect 5757 -6227 5857 -6183
rect 5961 -6227 6061 -6183
rect 5584 -6282 5678 -6272
rect 3997 -6286 5678 -6282
rect 3997 -6352 5598 -6286
rect 5664 -6352 5678 -6286
rect 3997 -6357 5678 -6352
rect 5584 -6366 5678 -6357
<< polycontact >>
rect -1658 1656 -1598 1728
rect 3146 1647 3209 1710
rect 3542 1705 3619 1782
rect 3752 1692 3829 1769
rect 2158 1370 2230 1418
rect 4175 1637 4233 1695
rect 5021 1576 5093 1623
rect 2944 1338 3003 1397
rect 5573 1584 5645 1634
rect 4809 1339 4881 1386
rect -1670 961 -1598 1033
rect 2449 1043 2508 1102
rect 2158 935 2230 984
rect 3081 992 3141 1052
rect 3991 1058 4052 1119
rect 3474 774 3546 824
rect 2445 592 2505 652
rect 3828 743 3897 790
rect 4951 757 5023 809
rect 4695 637 4758 700
rect 3296 443 3354 501
rect 4542 435 4606 499
rect 3057 201 3121 265
rect 4072 236 4144 290
rect 4967 184 5026 243
rect 109 -61 175 -4
rect 346 -81 403 -9
rect 2961 -181 3022 -120
rect 2452 -401 2503 -350
rect -1670 -502 -1598 -430
rect 4072 -459 4144 -409
rect 5627 -82 5699 -36
rect 5626 -376 5698 -329
rect -1670 -871 -1598 -824
rect -1428 -820 -1356 -748
rect 2158 -885 2230 -813
rect 2446 -1193 2507 -1132
rect 3050 -1192 3127 -1115
rect 4959 -988 5019 -928
rect 5626 -950 5698 -901
rect 4170 -1124 4236 -1072
rect 3868 -1402 3933 -1330
rect -1670 -1619 -1598 -1547
rect 2158 -1584 2230 -1538
rect 3807 -1756 3879 -1707
rect 2451 -1931 2509 -1873
rect 3603 -1856 3675 -1807
rect 5951 -1869 6023 -1819
rect 4256 -2184 4314 -2126
rect -719 -3079 -656 -3019
rect 35 -3100 107 -3051
rect 2383 -3111 2455 -3063
rect -2015 -3297 -1952 -3238
rect -1428 -3283 -1365 -3223
rect -1718 -3442 -1655 -3382
rect -717 -3537 -654 -3477
rect 1938 -3419 2007 -3365
rect 35 -3595 107 -3547
rect 851 -3590 923 -3543
rect 1871 -3610 1942 -3563
rect 2203 -3615 2275 -3568
rect 2407 -3615 2479 -3568
rect -719 -3947 -656 -3887
rect -2015 -4165 -1952 -4106
rect -1428 -4151 -1365 -4091
rect 442 -3960 514 -3913
rect -1718 -4310 -1655 -4250
rect -717 -4405 -654 -4345
rect 35 -4315 107 -4266
rect 1871 -4311 1943 -4265
rect 2203 -4322 2275 -4274
rect 2407 -4318 2479 -4271
rect -719 -4806 -656 -4746
rect 179 -4687 241 -4615
rect 851 -4663 923 -4615
rect -2015 -5024 -1952 -4965
rect -1428 -5010 -1365 -4950
rect -1718 -5169 -1655 -5109
rect 35 -5029 107 -4983
rect 387 -5029 459 -4980
rect 1487 -5052 1535 -4980
rect 1871 -4999 1943 -4953
rect 2203 -4999 2275 -4953
rect 2407 -5003 2479 -4953
rect -717 -5264 -654 -5204
rect 3603 -2518 3675 -2469
rect 5951 -2499 6023 -2449
rect 3755 -2860 3826 -2809
rect 3603 -3166 3675 -3118
rect 4245 -3249 4305 -3192
rect 5951 -3187 6023 -3141
rect 3576 -3492 3646 -3422
rect 5439 -3541 5511 -3491
rect 5771 -3540 5843 -3493
rect 3519 -3809 3590 -3762
rect 5574 -3883 5644 -3813
rect 3603 -4216 3675 -4166
rect 5439 -4203 5511 -4152
rect 5771 -4216 5843 -4166
rect 5975 -4211 6047 -4164
rect 3476 -4558 3537 -4497
rect 3603 -4914 3674 -4858
rect 5439 -4907 5511 -4856
rect 5771 -4908 5843 -4859
rect 5975 -4903 6047 -4856
rect 5576 -5276 5644 -5208
rect -719 -5674 -656 -5614
rect -2015 -5892 -1952 -5833
rect -1428 -5878 -1365 -5818
rect 899 -5674 962 -5614
rect -397 -5892 -334 -5833
rect 190 -5878 253 -5818
rect 2508 -5674 2571 -5614
rect 3603 -5604 3674 -5554
rect 5439 -5605 5511 -5559
rect 5771 -5602 5843 -5552
rect 5975 -5604 6047 -5551
rect 1212 -5892 1275 -5833
rect 1799 -5878 1862 -5818
rect -1718 -6037 -1655 -5977
rect -100 -6037 -37 -5977
rect -717 -6132 -654 -6072
rect 1509 -6037 1572 -5977
rect 901 -6132 964 -6072
rect 3470 -5949 3530 -5889
rect 2510 -6132 2573 -6072
rect 5529 -5988 5588 -5929
rect 5975 -6011 6047 -5962
rect 3603 -6280 3675 -6228
rect 5598 -6352 5664 -6286
<< metal1 >>
rect 4691 2334 4779 2347
rect 3923 2319 4000 2330
rect 3790 2263 3933 2319
rect 3989 2263 4000 2319
rect 3923 2247 4000 2263
rect 4691 2269 4703 2334
rect 4766 2333 4779 2334
rect 4766 2270 4886 2333
rect 4766 2269 4779 2270
rect 4691 2252 4779 2269
rect -1365 2008 1976 2051
rect -1365 1938 -1191 2008
rect 1787 1938 1976 2008
rect 6224 1999 6343 2000
rect -1365 1901 -14 1938
rect 42 1901 1976 1938
rect -1365 1881 1976 1901
rect 2654 1989 6367 1999
rect 2654 1974 6369 1989
rect 2654 1920 2690 1974
rect 2763 1920 2834 1974
rect 2907 1920 2978 1974
rect 3051 1920 3122 1974
rect 3195 1920 3266 1974
rect 3339 1920 3410 1974
rect 3483 1920 3554 1974
rect 3627 1920 3698 1974
rect 3771 1920 3842 1974
rect 3915 1920 3986 1974
rect 4059 1920 4130 1974
rect 4203 1920 4274 1974
rect 4347 1920 4418 1974
rect 4491 1920 4562 1974
rect 4635 1920 4706 1974
rect 4779 1920 4850 1974
rect 4923 1920 4994 1974
rect 5067 1920 5138 1974
rect 5211 1920 5282 1974
rect 5355 1920 5426 1974
rect 5499 1920 5570 1974
rect 5643 1920 5714 1974
rect 5787 1920 5858 1974
rect 5931 1920 6002 1974
rect 6075 1920 6146 1974
rect 6219 1920 6369 1974
rect 2654 1878 6369 1920
rect -1973 1786 -1062 1834
rect -1973 -1247 -1925 1786
rect -1667 1728 -1589 1737
rect -1667 1656 -1658 1728
rect -1598 1717 -1589 1728
rect -1110 1717 -1062 1786
rect 2654 1826 2775 1878
rect 2654 1772 2678 1826
rect 2751 1772 2775 1826
rect 6223 1854 6369 1878
rect 6223 1800 6254 1854
rect 6327 1800 6369 1854
rect -1598 1656 -1508 1717
rect -1667 1647 -1508 1656
rect -1557 1609 -1508 1647
rect -1172 1663 -711 1717
rect -1761 1593 -1712 1607
rect -1761 1499 -1759 1593
rect -1713 1499 -1712 1593
rect -1761 1439 -1712 1499
rect -1557 1593 -1507 1609
rect -1557 1499 -1555 1593
rect -1509 1499 -1507 1593
rect -1557 1490 -1507 1499
rect -1774 1432 -1697 1439
rect -1556 1437 -1507 1490
rect -1375 1593 -1321 1604
rect -1375 1499 -1372 1593
rect -1326 1499 -1321 1593
rect -1375 1437 -1321 1499
rect -1172 1593 -1118 1663
rect -765 1604 -711 1663
rect -354 1660 103 1714
rect 463 1668 921 1709
rect 1274 1687 1738 1709
rect 2654 1706 2775 1772
rect 3524 1787 3636 1799
rect 3137 1712 3218 1719
rect 463 1666 922 1668
rect -964 1601 -918 1604
rect -1172 1499 -1168 1593
rect -1122 1499 -1118 1593
rect -1556 1432 -1311 1437
rect -1774 1427 -1311 1432
rect -1774 1373 -1763 1427
rect -1709 1425 -1311 1427
rect -1709 1388 -1375 1425
rect -1709 1383 -1506 1388
rect -1709 1373 -1697 1383
rect -1774 1360 -1697 1373
rect -1761 1290 -1712 1360
rect -1761 1196 -1759 1290
rect -1713 1196 -1712 1290
rect -1761 1179 -1712 1196
rect -1556 1290 -1507 1383
rect -1384 1371 -1375 1388
rect -1321 1371 -1311 1425
rect -1384 1362 -1311 1371
rect -1556 1196 -1555 1290
rect -1509 1196 -1507 1290
rect -1556 1180 -1507 1196
rect -1375 1290 -1321 1362
rect -1375 1196 -1372 1290
rect -1326 1196 -1321 1290
rect -1375 1185 -1321 1196
rect -1172 1290 -1118 1499
rect -968 1593 -914 1601
rect -968 1499 -964 1593
rect -918 1499 -914 1593
rect -968 1431 -914 1499
rect -766 1593 -711 1604
rect -766 1499 -760 1593
rect -714 1499 -711 1593
rect -978 1418 -905 1431
rect -978 1364 -968 1418
rect -914 1364 -905 1418
rect -978 1356 -905 1364
rect -1172 1196 -1168 1290
rect -1122 1196 -1118 1290
rect -1172 1182 -1118 1196
rect -968 1290 -914 1356
rect -968 1196 -964 1290
rect -918 1196 -914 1290
rect -968 1182 -914 1196
rect -766 1290 -711 1499
rect -766 1196 -760 1290
rect -714 1196 -711 1290
rect -560 1593 -506 1623
rect -354 1603 -300 1660
rect -148 1603 -102 1604
rect -560 1499 -556 1593
rect -510 1499 -506 1593
rect -560 1290 -506 1499
rect -560 1242 -556 1290
rect -766 1185 -711 1196
rect -965 1112 -916 1182
rect -1272 1063 -916 1112
rect -765 1121 -711 1185
rect -572 1233 -556 1242
rect -510 1242 -506 1290
rect -355 1593 -300 1603
rect -355 1499 -352 1593
rect -306 1499 -300 1593
rect -355 1290 -300 1499
rect -154 1593 -100 1603
rect -154 1499 -148 1593
rect -102 1499 -100 1593
rect -154 1431 -100 1499
rect 49 1593 103 1660
rect 461 1655 922 1666
rect 49 1499 56 1593
rect 102 1499 103 1593
rect 260 1593 306 1604
rect -157 1419 -97 1431
rect -157 1363 -156 1419
rect -100 1363 -97 1419
rect -157 1351 -97 1363
rect -510 1233 -490 1242
rect -572 1177 -559 1233
rect -503 1177 -490 1233
rect -355 1196 -352 1290
rect -306 1196 -300 1290
rect -355 1184 -300 1196
rect -154 1290 -100 1351
rect -154 1196 -148 1290
rect -102 1196 -100 1290
rect -154 1184 -100 1196
rect 49 1290 103 1499
rect 49 1196 56 1290
rect 102 1196 103 1290
rect 254 1499 260 1527
rect 461 1593 517 1655
rect 306 1499 308 1527
rect 254 1290 308 1499
rect 254 1238 260 1290
rect -572 1175 -490 1177
rect -354 1121 -300 1184
rect -765 1067 -300 1121
rect 49 1125 103 1196
rect 241 1237 260 1238
rect 306 1238 308 1290
rect 461 1499 464 1593
rect 510 1499 517 1593
rect 668 1593 714 1604
rect 461 1290 517 1499
rect 664 1499 668 1527
rect 867 1593 922 1655
rect 1274 1655 1740 1687
rect 714 1499 718 1527
rect 664 1431 718 1499
rect 867 1499 872 1593
rect 918 1499 922 1593
rect 1076 1593 1122 1604
rect 660 1419 721 1431
rect 660 1363 662 1419
rect 718 1363 721 1419
rect 660 1351 721 1363
rect 306 1237 322 1238
rect 241 1180 253 1237
rect 310 1180 322 1237
rect 461 1196 464 1290
rect 510 1196 517 1290
rect 461 1186 517 1196
rect 241 1179 322 1180
rect 463 1125 517 1186
rect 664 1290 718 1351
rect 664 1196 668 1290
rect 714 1196 718 1290
rect 664 1182 718 1196
rect 867 1290 922 1499
rect 867 1196 872 1290
rect 918 1196 922 1290
rect 1071 1499 1076 1527
rect 1274 1593 1329 1655
rect 1122 1499 1125 1527
rect 1071 1290 1125 1499
rect 1071 1246 1076 1290
rect 867 1184 922 1196
rect 1058 1245 1076 1246
rect 1122 1246 1125 1290
rect 1274 1499 1280 1593
rect 1326 1499 1329 1593
rect 1484 1593 1530 1604
rect 1274 1290 1329 1499
rect 1477 1499 1484 1527
rect 1684 1593 1740 1655
rect 2654 1652 2678 1706
rect 2751 1652 2775 1706
rect 1892 1597 1938 1604
rect 2069 1597 2115 1604
rect 2273 1600 2319 1604
rect 1530 1499 1531 1527
rect 1477 1431 1531 1499
rect 1684 1499 1688 1593
rect 1734 1499 1740 1593
rect 1474 1419 1539 1431
rect 1474 1363 1477 1419
rect 1533 1363 1539 1419
rect 1474 1351 1539 1363
rect 1122 1245 1138 1246
rect 1058 1189 1070 1245
rect 1126 1189 1138 1245
rect 1058 1188 1138 1189
rect 1274 1196 1280 1290
rect 1326 1196 1329 1290
rect 1071 1185 1125 1188
rect 49 1071 517 1125
rect 867 1128 921 1184
rect 1274 1182 1329 1196
rect 1477 1290 1531 1351
rect 1477 1196 1484 1290
rect 1530 1196 1531 1290
rect 1477 1186 1531 1196
rect 1684 1290 1740 1499
rect 1684 1196 1688 1290
rect 1734 1196 1740 1290
rect 1888 1593 1942 1597
rect 1888 1499 1892 1593
rect 1938 1499 1942 1593
rect 1888 1419 1942 1499
rect 2066 1593 2119 1597
rect 2066 1499 2069 1593
rect 2115 1499 2119 1593
rect 2066 1432 2119 1499
rect 2271 1593 2323 1600
rect 2271 1499 2273 1593
rect 2319 1499 2323 1593
rect 2271 1432 2323 1499
rect 2066 1419 2323 1432
rect 1888 1418 2323 1419
rect 1888 1370 2158 1418
rect 2230 1370 2323 1418
rect 1888 1369 2323 1370
rect 1888 1290 1942 1369
rect 1888 1256 1892 1290
rect 1875 1250 1892 1256
rect 1484 1185 1530 1186
rect 1684 1185 1740 1196
rect 1874 1248 1892 1250
rect 1938 1256 1942 1290
rect 2066 1356 2323 1369
rect 2066 1290 2119 1356
rect 1938 1248 1955 1256
rect 1874 1192 1886 1248
rect 1942 1192 1955 1248
rect 1874 1191 1955 1192
rect 2066 1196 2069 1290
rect 2115 1196 2119 1290
rect 1874 1190 1952 1191
rect 1888 1185 1942 1190
rect 1684 1184 1738 1185
rect 1274 1128 1328 1182
rect 2066 1180 2119 1196
rect 2271 1290 2323 1356
rect 2271 1196 2273 1290
rect 2319 1196 2323 1290
rect 2271 1183 2323 1196
rect 2654 1586 2775 1652
rect 2654 1532 2678 1586
rect 2751 1532 2775 1586
rect 2654 1466 2775 1532
rect 3030 1710 3305 1712
rect 3030 1647 3146 1710
rect 3209 1677 3305 1710
rect 3371 1677 3429 1755
rect 3524 1700 3538 1787
rect 3625 1700 3636 1787
rect 3524 1688 3636 1700
rect 3743 1769 3838 1778
rect 3743 1692 3752 1769
rect 3829 1692 3838 1769
rect 3743 1683 3838 1692
rect 3914 1756 4010 1771
rect 3914 1687 3928 1756
rect 3997 1687 4010 1756
rect 6223 1734 6369 1800
rect 3914 1686 4010 1687
rect 4166 1695 4242 1704
rect 4166 1686 4175 1695
rect 3914 1677 4175 1686
rect 3209 1647 3429 1677
rect 3030 1639 3429 1647
rect 3030 1557 3087 1639
rect 3137 1638 3429 1639
rect 3248 1619 3429 1638
rect 3932 1637 4175 1677
rect 4233 1686 4242 1695
rect 4233 1637 4406 1686
rect 3248 1557 3305 1619
rect 3371 1562 3429 1619
rect 3584 1621 3646 1635
rect 3584 1565 3587 1621
rect 3643 1565 3646 1621
rect 3584 1562 3646 1565
rect 3932 1631 4406 1637
rect 3716 1562 3769 1563
rect 3932 1562 3987 1631
rect 4166 1628 4242 1631
rect 3371 1557 3648 1562
rect 3712 1557 3987 1562
rect 4351 1558 4406 1631
rect 4683 1684 4786 1700
rect 4683 1623 4704 1684
rect 4765 1623 4786 1684
rect 6223 1680 6254 1734
rect 6327 1680 6369 1734
rect 4683 1610 4786 1623
rect 5010 1643 5104 1651
rect 5010 1623 5034 1643
rect 4130 1557 4406 1558
rect 3030 1511 3041 1557
rect 3087 1511 3098 1557
rect 3242 1511 3253 1557
rect 3299 1511 3310 1557
rect 3370 1511 3381 1557
rect 3427 1511 3593 1557
rect 3639 1511 3650 1557
rect 3710 1511 3721 1557
rect 3767 1511 3933 1557
rect 3979 1511 3990 1557
rect 4130 1511 4145 1557
rect 4191 1511 4357 1557
rect 4403 1511 4414 1557
rect 3030 1499 3087 1511
rect 3248 1506 3305 1511
rect 3371 1500 3429 1511
rect 3584 1483 3646 1511
rect 2654 1412 2678 1466
rect 2751 1412 2775 1466
rect 3716 1412 3769 1511
rect 3932 1498 3987 1511
rect 4130 1503 4406 1511
rect 4351 1502 4406 1503
rect 2654 1346 2775 1412
rect 2654 1292 2678 1346
rect 2751 1292 2775 1346
rect 2935 1397 3012 1406
rect 2935 1338 2944 1397
rect 3003 1386 3012 1397
rect 3375 1386 3769 1412
rect 3003 1359 3769 1386
rect 4703 1491 4766 1610
rect 5010 1576 5021 1623
rect 5095 1582 5104 1643
rect 5093 1576 5104 1582
rect 5010 1569 5104 1576
rect 5564 1636 5656 1644
rect 5564 1634 5581 1636
rect 5643 1634 5656 1636
rect 5564 1584 5573 1634
rect 5645 1584 5656 1634
rect 5564 1574 5581 1584
rect 5643 1574 5656 1584
rect 5012 1567 5102 1569
rect 5564 1559 5656 1574
rect 6223 1614 6369 1680
rect 6223 1560 6254 1614
rect 6327 1560 6369 1614
rect 4913 1491 4985 1506
rect 4703 1445 4716 1491
rect 4762 1445 4773 1491
rect 4913 1445 4928 1491
rect 4974 1445 4985 1491
rect 4703 1396 4766 1445
rect 4913 1403 4985 1445
rect 5128 1491 5191 1506
rect 5259 1491 5317 1501
rect 5469 1491 5527 1506
rect 5684 1491 5742 1503
rect 5811 1491 5869 1498
rect 6023 1491 6081 1503
rect 6223 1494 6369 1560
rect 5128 1445 5140 1491
rect 5186 1445 5197 1491
rect 5257 1445 5268 1491
rect 5314 1445 5325 1491
rect 5469 1445 5480 1491
rect 5526 1445 5537 1491
rect 5681 1445 5692 1491
rect 5738 1445 5749 1491
rect 5809 1445 5820 1491
rect 5866 1445 5877 1491
rect 6021 1445 6032 1491
rect 6078 1445 6089 1491
rect 5128 1403 5191 1445
rect 4913 1396 5191 1403
rect 4703 1391 5191 1396
rect 4703 1386 5023 1391
rect 3003 1338 3428 1359
rect 2935 1334 3428 1338
rect 2935 1329 3098 1334
rect 2654 1226 2775 1292
rect 867 1074 1328 1128
rect 2654 1172 2678 1226
rect 2751 1172 2775 1226
rect 3046 1291 3098 1329
rect 3046 1197 3049 1291
rect 3095 1197 3098 1291
rect 3046 1182 3098 1197
rect 3251 1291 3303 1334
rect 3251 1197 3253 1291
rect 3299 1197 3303 1291
rect 3251 1185 3303 1197
rect 3375 1291 3428 1334
rect 4703 1339 4809 1386
rect 4881 1339 5023 1386
rect 4703 1337 5023 1339
rect 5077 1390 5191 1391
rect 5077 1337 5192 1390
rect 5259 1380 5317 1445
rect 5469 1380 5527 1445
rect 5684 1380 5742 1445
rect 4703 1330 5191 1337
rect 3375 1197 3381 1291
rect 3427 1197 3428 1291
rect 3375 1183 3428 1197
rect 3581 1291 3637 1309
rect 3581 1197 3585 1291
rect 3631 1197 3637 1291
rect 3581 1193 3637 1197
rect 3784 1291 3837 1305
rect 3784 1197 3789 1291
rect 3835 1197 3837 1291
rect 3784 1193 3837 1197
rect 3993 1291 4043 1309
rect 4039 1197 4043 1291
rect 3580 1189 3638 1193
rect 3578 1184 3646 1189
rect 3783 1184 3839 1193
rect 2440 1102 2517 1111
rect -1679 1033 -1589 1042
rect -1679 961 -1670 1033
rect -1598 1021 -1589 1033
rect -1598 961 -1508 1021
rect -1679 952 -1508 961
rect -1758 862 -1709 869
rect -1759 851 -1709 862
rect -1713 757 -1709 851
rect -1759 746 -1709 757
rect -1758 694 -1709 746
rect -1557 851 -1508 952
rect -1377 987 -1319 1000
rect -1377 933 -1375 987
rect -1321 933 -1319 987
rect -1377 921 -1319 933
rect -1557 757 -1555 851
rect -1509 757 -1508 851
rect -1557 694 -1508 757
rect -1373 851 -1324 921
rect -1373 757 -1372 851
rect -1326 757 -1324 851
rect -1373 694 -1324 757
rect -1874 645 -1324 694
rect -1874 -1067 -1826 645
rect -1272 565 -1223 1063
rect 2440 1043 2449 1102
rect 2508 1043 2517 1102
rect 2440 1034 2517 1043
rect 2654 1106 2775 1172
rect 3578 1128 3581 1184
rect 3637 1128 3646 1184
rect 3578 1116 3646 1128
rect 3772 1130 3784 1184
rect 3838 1171 3850 1184
rect 3993 1171 4043 1197
rect 3838 1130 4043 1171
rect 3772 1128 4043 1130
rect 4197 1291 4247 1302
rect 4243 1197 4247 1291
rect 3772 1121 4061 1128
rect 3772 1118 3850 1121
rect 3982 1120 4061 1121
rect 4197 1124 4247 1197
rect 4397 1291 4447 1308
rect 4703 1306 4766 1330
rect 4397 1197 4401 1291
rect 4397 1132 4447 1197
rect 4702 1249 4766 1306
rect 4913 1326 5191 1330
rect 4913 1249 4976 1326
rect 5128 1249 5191 1326
rect 5259 1322 5742 1380
rect 5259 1249 5317 1322
rect 5469 1249 5527 1322
rect 5684 1249 5742 1322
rect 5811 1398 5869 1445
rect 6023 1398 6081 1445
rect 5811 1389 6081 1398
rect 5811 1333 5932 1389
rect 5988 1333 6081 1389
rect 5811 1320 6081 1333
rect 5811 1249 5869 1320
rect 6023 1249 6081 1320
rect 6223 1440 6254 1494
rect 6327 1440 6369 1494
rect 6223 1374 6369 1440
rect 6223 1320 6254 1374
rect 6327 1320 6369 1374
rect 6223 1254 6369 1320
rect 4702 1203 4716 1249
rect 4762 1203 4773 1249
rect 4913 1203 4928 1249
rect 4974 1203 4985 1249
rect 5128 1203 5140 1249
rect 5186 1203 5197 1249
rect 5257 1203 5268 1249
rect 5314 1203 5325 1249
rect 5469 1203 5480 1249
rect 5526 1203 5537 1249
rect 5681 1203 5692 1249
rect 5738 1203 5749 1249
rect 5809 1203 5820 1249
rect 5866 1203 5877 1249
rect 6021 1203 6032 1249
rect 6078 1203 6089 1249
rect 4702 1193 4766 1203
rect 4913 1198 4976 1203
rect 5128 1198 5191 1203
rect 5259 1198 5317 1203
rect 5684 1200 5742 1203
rect 4702 1132 4758 1193
rect 4397 1124 4764 1132
rect 4197 1120 4764 1124
rect 3982 1119 4764 1120
rect 2654 1052 2678 1106
rect 2751 1052 2775 1106
rect 3072 1060 3150 1061
rect 3031 1056 3150 1060
rect 3982 1058 3991 1119
rect 4052 1082 4764 1119
rect 5130 1089 5181 1198
rect 5690 1135 5739 1200
rect 5811 1195 5869 1203
rect 6023 1200 6081 1203
rect 6223 1200 6254 1254
rect 6327 1200 6369 1254
rect 5687 1094 5747 1135
rect 6223 1134 6369 1200
rect 4052 1074 4447 1082
rect 4052 1058 4061 1074
rect -564 988 -499 1001
rect -1169 909 -712 959
rect -564 932 -559 988
rect -503 932 -499 988
rect 244 988 319 998
rect -564 917 -499 932
rect -358 925 104 977
rect -1169 851 -1119 909
rect -1169 757 -1168 851
rect -1122 757 -1119 851
rect -1169 738 -1119 757
rect -967 862 -919 863
rect -967 851 -918 862
rect -967 757 -964 851
rect -967 746 -918 757
rect -764 851 -712 909
rect -764 757 -760 851
rect -714 757 -712 851
rect -1354 564 -1034 565
rect -967 564 -919 746
rect -764 687 -712 757
rect -561 851 -505 917
rect -561 757 -556 851
rect -510 757 -505 851
rect -561 738 -505 757
rect -358 851 -306 925
rect -358 757 -352 851
rect -358 687 -306 757
rect -764 635 -306 687
rect -151 851 -100 863
rect -151 757 -148 851
rect -102 757 -100 851
rect -151 564 -100 757
rect 52 851 104 925
rect 244 932 253 988
rect 309 932 319 988
rect 1066 988 1127 1002
rect 244 922 319 932
rect 462 981 512 982
rect 462 934 919 981
rect 52 757 56 851
rect 102 757 104 851
rect 52 677 104 757
rect 256 851 307 922
rect 256 757 260 851
rect 306 757 307 851
rect 256 739 307 757
rect 462 851 512 934
rect 462 757 464 851
rect 510 757 512 851
rect 462 677 512 757
rect 52 628 512 677
rect 664 851 718 863
rect 664 757 668 851
rect 714 757 718 851
rect 664 564 718 757
rect 869 851 919 934
rect 1066 932 1067 988
rect 1123 932 1127 988
rect 1066 920 1127 932
rect 1276 946 1736 998
rect 869 757 872 851
rect 918 757 919 851
rect 869 746 919 757
rect 1075 851 1122 920
rect 1075 757 1076 851
rect 869 680 916 746
rect 1075 742 1122 757
rect 1276 851 1328 946
rect 1276 757 1280 851
rect 1326 757 1328 851
rect 1276 680 1328 757
rect 869 633 1328 680
rect 1484 851 1532 866
rect 1530 757 1532 851
rect 1484 564 1532 757
rect 1684 851 1736 946
rect 1873 988 1955 999
rect 1873 932 1886 988
rect 1942 932 1955 988
rect 1873 925 1955 932
rect 2066 984 2239 998
rect 2066 935 2158 984
rect 2230 935 2239 984
rect 1889 922 1942 925
rect 1684 757 1688 851
rect 1734 757 1736 851
rect 1684 689 1736 757
rect 1890 851 1942 922
rect 1890 757 1892 851
rect 1938 757 1942 851
rect 1890 727 1942 757
rect 2066 921 2239 935
rect 2066 851 2118 921
rect 2066 757 2069 851
rect 2115 757 2118 851
rect 2066 727 2118 757
rect 2273 851 2326 866
rect 2319 757 2326 851
rect 2273 727 2326 757
rect 1671 677 1743 689
rect 1671 623 1683 677
rect 1737 623 1743 677
rect 1890 675 2326 727
rect 2452 661 2504 1034
rect 2654 986 2775 1052
rect 3030 1052 3640 1056
rect 3030 1006 3081 1052
rect 2654 932 2678 986
rect 2751 932 2775 986
rect 2654 866 2775 932
rect 3031 992 3081 1006
rect 3141 1044 3640 1052
rect 3982 1049 4061 1058
rect 3141 1027 3650 1044
rect 3141 1006 3588 1027
rect 3141 992 3150 1006
rect 3031 983 3150 992
rect 3031 929 3083 983
rect 3251 929 3301 1006
rect 3372 929 3432 1006
rect 3576 966 3588 1006
rect 3649 966 3650 1027
rect 4258 1026 4547 1027
rect 4258 967 4270 1026
rect 4329 967 4547 1026
rect 4258 966 4338 967
rect 3576 958 3650 966
rect 3582 929 3650 958
rect 3711 929 4192 943
rect 4262 929 4330 966
rect 3030 883 3041 929
rect 3087 883 3098 929
rect 3242 883 3253 929
rect 3299 883 3310 929
rect 3370 883 3381 929
rect 3427 883 3438 929
rect 3582 883 3593 929
rect 3639 883 3650 929
rect 3710 883 3721 929
rect 3767 883 3933 929
rect 3979 883 4145 929
rect 4191 883 4202 929
rect 4262 883 4273 929
rect 4319 883 4330 929
rect 4474 929 4547 967
rect 4474 883 4485 929
rect 4531 883 4547 929
rect 3031 881 3083 883
rect 3251 881 3301 883
rect 3372 875 3432 883
rect 3590 882 3640 883
rect 2654 812 2678 866
rect 2751 812 2775 866
rect 2654 746 2775 812
rect 3465 824 3555 833
rect 3465 805 3474 824
rect 2654 692 2678 746
rect 2751 692 2775 746
rect 3458 796 3474 805
rect 3458 723 3471 796
rect 3546 774 3555 824
rect 3884 823 3982 835
rect 3884 799 3900 823
rect 3544 765 3555 774
rect 3819 790 3900 799
rect 3544 723 3554 765
rect 3819 743 3828 790
rect 3897 754 3900 790
rect 3969 798 3982 823
rect 3969 754 3989 798
rect 3897 743 3989 754
rect 3819 735 3989 743
rect 4135 760 4190 883
rect 4269 882 4329 883
rect 4487 831 4547 883
rect 4702 831 4758 1082
rect 5130 1038 5522 1089
rect 5687 1045 5928 1094
rect 4487 776 4758 831
rect 4487 775 4544 776
rect 4602 775 4758 776
rect 4856 965 4912 983
rect 4856 871 4862 965
rect 4908 871 4912 965
rect 4856 823 4912 871
rect 5061 965 5117 976
rect 5061 871 5066 965
rect 5112 871 5117 965
rect 5061 831 5117 871
rect 5037 823 5117 831
rect 4856 822 5117 823
rect 4856 809 5039 822
rect 3819 734 3906 735
rect 3458 711 3554 723
rect 4135 705 4390 760
rect 4856 757 4951 809
rect 5023 757 5039 809
rect 4856 744 5039 757
rect 5102 744 5117 822
rect 4856 743 5117 744
rect 1671 611 1743 623
rect 2436 652 2514 661
rect 2436 592 2445 652
rect 2505 592 2514 652
rect 2436 583 2514 592
rect 2654 626 2775 692
rect 2965 659 3024 661
rect 1711 564 1913 565
rect -1354 511 1913 564
rect -1354 436 -801 511
rect 1521 436 1913 511
rect -1354 381 1913 436
rect -1776 259 -1695 271
rect -1776 205 -1762 259
rect -1708 205 -1695 259
rect -1776 193 -1695 205
rect -1760 175 -1711 193
rect -1760 81 -1759 175
rect -1713 81 -1711 175
rect -1760 -151 -1711 81
rect -1559 175 -1503 190
rect -1559 81 -1555 175
rect -1509 81 -1503 175
rect -1559 -7 -1503 81
rect -1354 175 -1298 381
rect -1354 81 -1351 175
rect -1305 81 -1298 175
rect -1568 -16 -1494 -7
rect -1568 -72 -1559 -16
rect -1503 -72 -1494 -16
rect -1568 -80 -1494 -72
rect -1560 -81 -1502 -80
rect -1760 -245 -1759 -151
rect -1713 -245 -1711 -151
rect -1760 -317 -1711 -245
rect -1559 -151 -1503 -81
rect -1559 -245 -1555 -151
rect -1509 -245 -1503 -151
rect -1559 -261 -1503 -245
rect -1354 -151 -1298 81
rect -1152 175 -1097 186
rect -1152 81 -1147 175
rect -1101 81 -1097 175
rect -1152 -4 -1097 81
rect -948 175 -894 187
rect -948 81 -943 175
rect -897 81 -894 175
rect -1158 -16 -1085 -4
rect -1158 -72 -1150 -16
rect -1094 -72 -1085 -16
rect -1158 -81 -1085 -72
rect -1354 -245 -1351 -151
rect -1305 -245 -1298 -151
rect -1354 -261 -1298 -245
rect -1152 -151 -1097 -81
rect -1152 -245 -1147 -151
rect -1101 -245 -1097 -151
rect -1152 -260 -1097 -245
rect -948 -151 -894 81
rect -948 -245 -943 -151
rect -897 -245 -894 -151
rect -948 -317 -894 -245
rect -1760 -366 -894 -317
rect -818 175 -766 191
rect -818 81 -815 175
rect -769 81 -766 175
rect -818 -151 -766 81
rect -615 175 -562 190
rect -615 81 -611 175
rect -565 81 -562 175
rect -615 -9 -562 81
rect -408 175 -358 381
rect 37 320 108 332
rect 37 266 49 320
rect 103 266 108 320
rect 37 253 108 266
rect -408 81 -407 175
rect -361 81 -358 175
rect -625 -26 -545 -9
rect -625 -80 -615 -26
rect -561 -80 -545 -26
rect -625 -94 -545 -80
rect -818 -245 -815 -151
rect -769 -245 -766 -151
rect -818 -404 -766 -245
rect -615 -151 -562 -94
rect -615 -245 -611 -151
rect -565 -245 -562 -151
rect -615 -263 -562 -245
rect -408 -151 -358 81
rect -408 -245 -407 -151
rect -361 -245 -358 -151
rect -833 -412 -751 -404
rect -1679 -430 -1589 -421
rect -1679 -502 -1670 -430
rect -1598 -502 -1589 -430
rect -833 -466 -819 -412
rect -765 -466 -751 -412
rect -833 -476 -751 -466
rect -1679 -511 -1589 -502
rect -1671 -598 -1596 -511
rect -408 -549 -358 -245
rect -283 175 -231 188
rect -283 81 -279 175
rect -233 81 -231 175
rect -283 -151 -231 81
rect -81 175 -25 190
rect -81 81 -75 175
rect -29 81 -25 175
rect -81 16 -25 81
rect 52 175 99 253
rect 52 81 53 175
rect 52 72 99 81
rect 53 70 99 72
rect 255 175 306 187
rect 255 81 257 175
rect 303 81 306 175
rect 255 70 306 81
rect 458 175 516 381
rect 458 81 461 175
rect 507 81 516 175
rect -92 13 -22 16
rect -92 -41 -80 13
rect -26 -41 -22 13
rect -92 -55 -22 -41
rect 46 -4 186 8
rect 46 -61 109 -4
rect 175 -61 186 -4
rect 46 -78 186 -61
rect 254 -9 412 0
rect -283 -245 -279 -151
rect -233 -245 -231 -151
rect -283 -268 -231 -245
rect -81 -151 -29 -135
rect -81 -245 -75 -151
rect -298 -271 -218 -268
rect -298 -325 -284 -271
rect -230 -325 -218 -271
rect -298 -331 -218 -325
rect -81 -323 -29 -245
rect 46 -151 103 -78
rect 46 -245 53 -151
rect 99 -245 103 -151
rect 46 -258 103 -245
rect 254 -81 346 -9
rect 403 -81 412 -9
rect 254 -90 412 -81
rect 254 -151 305 -90
rect 254 -245 257 -151
rect 303 -245 305 -151
rect 254 -259 305 -245
rect 458 -151 516 81
rect 580 175 643 193
rect 580 81 589 175
rect 635 81 643 175
rect 580 18 643 81
rect 791 175 841 223
rect 791 81 793 175
rect 839 81 841 175
rect 576 14 650 18
rect 576 -42 583 14
rect 639 -42 650 14
rect 576 -55 650 -42
rect 458 -245 461 -151
rect 507 -245 516 -151
rect 458 -323 516 -245
rect 585 -151 638 -131
rect 585 -245 589 -151
rect 635 -245 638 -151
rect 585 -323 638 -245
rect 791 -151 841 81
rect 791 -245 793 -151
rect 839 -245 841 -151
rect 791 -258 841 -245
rect 917 175 972 381
rect 917 81 921 175
rect 967 81 972 175
rect 917 -151 972 81
rect 1118 175 1175 190
rect 1118 81 1125 175
rect 1171 81 1175 175
rect 1118 -32 1175 81
rect 1325 175 1376 209
rect 1325 81 1329 175
rect 1375 81 1376 175
rect 1099 -41 1180 -32
rect 1099 -97 1115 -41
rect 1171 -97 1180 -41
rect 1099 -106 1180 -97
rect 917 -245 921 -151
rect 967 -245 972 -151
rect -81 -369 638 -323
rect 785 -270 858 -258
rect 917 -264 972 -245
rect 1118 -151 1175 -106
rect 1118 -245 1125 -151
rect 1171 -245 1175 -151
rect 1118 -260 1175 -245
rect 1325 -151 1376 81
rect 1325 -245 1329 -151
rect 1375 -245 1376 -151
rect 785 -326 789 -270
rect 845 -326 858 -270
rect 785 -339 858 -326
rect -81 -370 -28 -369
rect 1325 -372 1376 -245
rect 1453 175 1505 192
rect 1453 81 1457 175
rect 1503 81 1505 175
rect 1453 -151 1505 81
rect 1658 175 1710 189
rect 1658 81 1661 175
rect 1707 81 1710 175
rect 1658 15 1710 81
rect 1861 175 1913 381
rect 2268 260 2341 273
rect 2268 204 2278 260
rect 2334 204 2341 260
rect 1861 81 1865 175
rect 1911 81 1913 175
rect 1644 10 1725 15
rect 1644 -46 1657 10
rect 1713 -46 1725 10
rect 1644 -55 1725 -46
rect 1453 -245 1457 -151
rect 1503 -245 1505 -151
rect 1453 -301 1505 -245
rect 1658 -151 1710 -55
rect 1658 -245 1661 -151
rect 1707 -245 1710 -151
rect 1658 -262 1710 -245
rect 1861 -151 1913 81
rect 2065 175 2117 188
rect 2268 185 2341 204
rect 2065 81 2069 175
rect 2115 81 2117 175
rect 2065 23 2117 81
rect 2270 175 2321 185
rect 2270 81 2273 175
rect 2319 81 2321 175
rect 2059 10 2132 23
rect 2059 -46 2067 10
rect 2123 -46 2132 10
rect 2059 -58 2132 -46
rect 1861 -245 1865 -151
rect 1911 -245 1913 -151
rect 1861 -258 1913 -245
rect 2065 -151 2117 -58
rect 2065 -245 2069 -151
rect 2115 -245 2117 -151
rect 2065 -263 2117 -245
rect 2270 -151 2321 81
rect 2270 -245 2273 -151
rect 2319 -245 2321 -151
rect 1453 -337 1589 -301
rect 2270 -337 2321 -245
rect 2445 -335 2509 583
rect 2654 572 2678 626
rect 2751 572 2775 626
rect 2962 645 3038 659
rect 2962 589 2971 645
rect 3027 589 3038 645
rect 2962 574 3038 589
rect 3123 645 3173 656
rect 2654 506 2775 572
rect 2654 452 2678 506
rect 2751 452 2775 506
rect 2654 386 2775 452
rect 2654 332 2678 386
rect 2751 332 2775 386
rect 2654 266 2775 332
rect 2965 382 3024 574
rect 3169 551 3173 645
rect 3123 497 3173 551
rect 3326 645 3376 679
rect 3925 672 3999 684
rect 3326 551 3327 645
rect 3373 551 3376 645
rect 3528 645 3582 659
rect 3528 552 3531 645
rect 3326 510 3376 551
rect 3287 501 3376 510
rect 3287 497 3296 501
rect 3123 447 3296 497
rect 3287 443 3296 447
rect 3354 497 3376 501
rect 3512 551 3531 552
rect 3577 552 3582 645
rect 3735 645 3783 661
rect 3577 551 3588 552
rect 3512 538 3588 551
rect 3512 497 3528 538
rect 3354 484 3528 497
rect 3582 484 3588 538
rect 3354 476 3588 484
rect 3781 551 3783 645
rect 3925 611 3928 672
rect 3989 611 3999 672
rect 4335 659 4390 705
rect 4675 708 4772 717
rect 3925 598 3939 611
rect 3735 490 3783 551
rect 3936 551 3939 598
rect 3985 598 3999 611
rect 4141 645 4189 657
rect 3936 543 3985 551
rect 3939 540 3985 543
rect 4141 551 4143 645
rect 4141 490 4189 551
rect 4335 645 4393 659
rect 4335 551 4347 645
rect 4548 645 4598 656
rect 4548 577 4551 645
rect 4335 548 4393 551
rect 4545 551 4551 577
rect 4597 551 4598 645
rect 4675 629 4687 708
rect 4758 629 4772 708
rect 4675 619 4772 629
rect 4856 663 4912 743
rect 5037 735 5117 743
rect 4856 569 4862 663
rect 4908 569 4912 663
rect 4856 559 4912 569
rect 5061 663 5117 735
rect 5061 569 5066 663
rect 5112 569 5117 663
rect 4862 558 4908 559
rect 5061 552 5117 569
rect 5266 965 5322 978
rect 5266 871 5270 965
rect 5316 871 5322 965
rect 5266 663 5322 871
rect 5471 965 5522 1038
rect 5678 975 5724 976
rect 5471 871 5474 965
rect 5520 871 5522 965
rect 5471 666 5522 871
rect 5670 965 5726 975
rect 5670 871 5678 965
rect 5724 871 5726 965
rect 5266 569 5270 663
rect 5316 569 5322 663
rect 5461 663 5540 666
rect 5461 656 5474 663
rect 5520 656 5540 663
rect 5461 600 5471 656
rect 5527 600 5540 656
rect 5461 592 5474 600
rect 3354 447 3586 476
rect 3354 443 3376 447
rect 3287 436 3376 443
rect 3735 442 4189 490
rect 4332 544 4408 548
rect 4545 544 4598 551
rect 4332 539 4598 544
rect 4332 483 4342 539
rect 4398 508 4598 539
rect 5266 508 5322 569
rect 5471 569 5474 592
rect 5520 592 5540 600
rect 5670 663 5726 871
rect 5879 965 5928 1045
rect 5879 871 5882 965
rect 5879 824 5928 871
rect 6223 1080 6254 1134
rect 6327 1080 6369 1134
rect 6223 1014 6369 1080
rect 6223 960 6254 1014
rect 6327 960 6369 1014
rect 6223 894 6369 960
rect 6223 840 6254 894
rect 6327 840 6369 894
rect 5873 811 5941 824
rect 5873 755 5876 811
rect 5932 755 5941 811
rect 5873 742 5941 755
rect 6223 774 6369 840
rect 5520 569 5522 592
rect 5471 557 5522 569
rect 5670 569 5678 663
rect 5724 569 5726 663
rect 4398 499 4615 508
rect 4398 494 4542 499
rect 4398 483 4408 494
rect 4332 472 4408 483
rect 3287 434 3363 436
rect 3735 382 3794 442
rect 4533 435 4542 494
rect 4606 435 4615 499
rect 5265 501 5346 508
rect 5670 501 5726 569
rect 5265 499 5726 501
rect 5265 443 5278 499
rect 5334 445 5726 499
rect 5879 669 5928 742
rect 6223 720 6254 774
rect 6327 720 6369 774
rect 5879 663 5931 669
rect 5879 569 5882 663
rect 5928 569 5931 663
rect 5334 443 5346 445
rect 5265 441 5346 443
rect 4533 426 4615 435
rect 2965 323 3794 382
rect 4529 319 5481 351
rect 5879 319 5931 569
rect 4063 290 4153 299
rect 4529 298 5931 319
rect 4063 279 4072 290
rect 2654 212 2678 266
rect 2751 212 2775 266
rect 3048 265 3130 274
rect 3048 256 3057 265
rect 2654 146 2775 212
rect 2654 92 2678 146
rect 2751 92 2775 146
rect 2654 26 2775 92
rect 2654 -28 2678 26
rect 2751 -28 2775 26
rect 2960 201 3057 256
rect 3121 244 3130 265
rect 3121 201 3212 244
rect 3363 219 3828 269
rect 3363 217 3444 219
rect 2960 192 3212 201
rect 2960 132 3008 192
rect 3164 132 3212 192
rect 3350 205 3444 217
rect 3350 135 3362 205
rect 3432 135 3444 205
rect 2960 121 3009 132
rect 2960 27 2963 121
rect 2960 16 3009 27
rect 3164 121 3213 132
rect 3350 122 3444 135
rect 3778 133 3828 219
rect 3979 236 4072 279
rect 4144 236 4235 290
rect 3979 227 4235 236
rect 3572 132 3620 133
rect 3164 27 3167 121
rect 3164 16 3213 27
rect 3368 121 3418 122
rect 3368 27 3371 121
rect 3417 27 3418 121
rect 2960 15 3008 16
rect 2654 -94 2775 -28
rect 3164 -36 3212 16
rect 2654 -148 2678 -94
rect 2751 -148 2775 -94
rect 3147 -49 3228 -36
rect 3147 -105 3160 -49
rect 3216 -105 3228 -49
rect 3368 -65 3418 27
rect 3572 121 3621 132
rect 3572 27 3575 121
rect 3572 16 3621 27
rect 3778 121 3829 133
rect 3778 27 3779 121
rect 3825 27 3829 121
rect 3572 -56 3620 16
rect 3778 -48 3829 27
rect 3979 121 4031 227
rect 3979 27 3983 121
rect 4029 27 4031 121
rect 2654 -214 2775 -148
rect 2952 -120 3031 -111
rect 3147 -117 3228 -105
rect 2952 -181 2961 -120
rect 3022 -181 3031 -120
rect 2952 -190 3031 -181
rect 2654 -268 2678 -214
rect 2751 -268 2775 -214
rect 2654 -334 2775 -268
rect 1453 -353 2321 -337
rect 1325 -382 1409 -372
rect 1325 -438 1341 -382
rect 1397 -438 1409 -382
rect 1537 -389 2321 -353
rect 2438 -350 2518 -335
rect 2438 -401 2452 -350
rect 2503 -401 2518 -350
rect 2438 -414 2518 -401
rect 2654 -388 2678 -334
rect 2751 -388 2775 -334
rect 2962 -257 3010 -190
rect 2962 -335 2963 -257
rect 1325 -439 1409 -438
rect -1671 -673 -1348 -598
rect -1435 -739 -1348 -673
rect -1250 -603 1947 -549
rect -1250 -681 -656 -603
rect 1599 -615 1947 -603
rect 1599 -677 2373 -615
rect 1599 -681 1947 -677
rect -1437 -748 -1347 -739
rect -1679 -822 -1589 -815
rect -1437 -820 -1428 -748
rect -1356 -820 -1347 -748
rect -1250 -750 1947 -681
rect 2300 -718 2373 -677
rect 2300 -720 2384 -718
rect -1679 -824 -1512 -822
rect -1679 -871 -1670 -824
rect -1598 -871 -1512 -824
rect -1437 -829 -1347 -820
rect -1679 -878 -1512 -871
rect -1679 -880 -1325 -878
rect -1558 -926 -1325 -880
rect -1760 -943 -1711 -929
rect -1760 -1037 -1759 -943
rect -1713 -1037 -1711 -943
rect -1760 -1064 -1711 -1037
rect -1558 -943 -1509 -926
rect -1558 -1037 -1555 -943
rect -1558 -1064 -1509 -1037
rect -1760 -1067 -1509 -1064
rect -1874 -1115 -1509 -1067
rect -1373 -943 -1325 -926
rect -1168 -935 -1122 -932
rect -1373 -1037 -1372 -943
rect -1326 -1037 -1325 -943
rect -1373 -1090 -1325 -1037
rect -1175 -943 -1117 -935
rect -1175 -1037 -1168 -943
rect -1122 -1037 -1117 -943
rect -1385 -1104 -1311 -1090
rect -1385 -1158 -1376 -1104
rect -1322 -1158 -1311 -1104
rect -1385 -1172 -1311 -1158
rect -1175 -1104 -1117 -1037
rect -968 -943 -912 -750
rect -968 -1037 -964 -943
rect -918 -1037 -912 -943
rect -968 -1056 -912 -1037
rect -765 -883 -299 -826
rect -765 -943 -708 -883
rect -556 -935 -510 -932
rect -765 -1037 -760 -943
rect -714 -1037 -708 -943
rect -765 -1104 -708 -1037
rect -562 -943 -507 -935
rect -562 -1037 -556 -943
rect -510 -1037 -507 -943
rect -562 -1091 -507 -1037
rect -356 -943 -299 -883
rect -356 -1037 -352 -943
rect -306 -1037 -299 -943
rect -1175 -1161 -708 -1104
rect -566 -1103 -503 -1091
rect -566 -1159 -561 -1103
rect -505 -1159 -503 -1103
rect -356 -1098 -299 -1037
rect -148 -943 -100 -750
rect -102 -1037 -100 -943
rect -148 -1052 -100 -1037
rect 50 -884 516 -827
rect 50 -943 107 -884
rect 260 -934 306 -932
rect 50 -1037 56 -943
rect 102 -1037 107 -943
rect 50 -1098 107 -1037
rect 255 -943 307 -934
rect 255 -1037 260 -943
rect 306 -1037 307 -943
rect 255 -1091 307 -1037
rect 459 -943 516 -884
rect 459 -1037 464 -943
rect 510 -1037 516 -943
rect -356 -1155 107 -1098
rect 253 -1103 316 -1091
rect -566 -1171 -503 -1159
rect 253 -1159 256 -1103
rect 312 -1159 316 -1103
rect 459 -1100 516 -1037
rect 663 -943 715 -750
rect 663 -1037 668 -943
rect 714 -1037 715 -943
rect 663 -1048 715 -1037
rect 870 -870 1328 -813
rect 870 -943 927 -870
rect 1076 -934 1122 -932
rect 870 -1037 872 -943
rect 918 -1037 927 -943
rect 870 -1100 927 -1037
rect 1075 -943 1124 -934
rect 1075 -1037 1076 -943
rect 1122 -1037 1124 -943
rect 1075 -1091 1124 -1037
rect 1271 -943 1328 -870
rect 1271 -1037 1280 -943
rect 1326 -1037 1328 -943
rect 459 -1157 927 -1100
rect 1066 -1103 1131 -1091
rect 253 -1171 316 -1159
rect 1066 -1159 1071 -1103
rect 1127 -1159 1131 -1103
rect 1271 -1094 1328 -1037
rect 1483 -943 1531 -750
rect 2300 -780 2312 -720
rect 2372 -780 2384 -720
rect 2300 -793 2384 -780
rect 1668 -803 1750 -798
rect 1668 -859 1681 -803
rect 1737 -859 1750 -803
rect 2149 -813 2239 -804
rect 2149 -815 2158 -813
rect 1668 -870 1750 -859
rect 2049 -869 2158 -815
rect 1483 -1037 1484 -943
rect 1530 -1037 1531 -943
rect 1483 -1046 1531 -1037
rect 1681 -930 1737 -870
rect 1886 -885 2158 -869
rect 2230 -885 2239 -813
rect 1886 -894 2239 -885
rect 1886 -928 2118 -894
rect 1681 -943 1740 -930
rect 1681 -1037 1688 -943
rect 1734 -1037 1740 -943
rect 1484 -1048 1530 -1046
rect 1681 -1094 1740 -1037
rect 1886 -943 1945 -928
rect 1886 -1037 1892 -943
rect 1938 -1037 1945 -943
rect 1886 -1091 1945 -1037
rect 2058 -943 2118 -928
rect 2058 -1037 2069 -943
rect 2115 -1037 2118 -943
rect 2058 -1059 2118 -1037
rect 2270 -943 2329 -929
rect 2270 -1037 2273 -943
rect 2319 -1037 2329 -943
rect 1271 -1151 1740 -1094
rect 1885 -1103 1953 -1091
rect 1066 -1171 1131 -1159
rect 1885 -1159 1894 -1103
rect 1950 -1159 1953 -1103
rect 1885 -1171 1953 -1159
rect 2058 -1114 2117 -1059
rect 2270 -1114 2329 -1037
rect 2058 -1173 2329 -1114
rect 2445 -1123 2507 -414
rect 2654 -454 2775 -388
rect 2654 -508 2678 -454
rect 2751 -508 2775 -454
rect 2654 -574 2775 -508
rect 2654 -628 2678 -574
rect 2751 -628 2775 -574
rect 2654 -694 2775 -628
rect 2961 -351 2963 -335
rect 3009 -315 3010 -257
rect 3154 -235 3220 -223
rect 3154 -291 3158 -235
rect 3214 -291 3220 -235
rect 3154 -315 3167 -291
rect 3009 -351 3167 -315
rect 3213 -316 3220 -291
rect 3369 -237 3417 -65
rect 3553 -68 3637 -56
rect 3553 -124 3568 -68
rect 3624 -124 3637 -68
rect 3553 -136 3637 -124
rect 3778 -237 3828 -48
rect 3979 -50 4031 27
rect 4185 132 4232 227
rect 4185 121 4233 132
rect 4185 27 4187 121
rect 4529 119 4582 298
rect 5428 267 5931 298
rect 6223 654 6369 720
rect 6223 600 6254 654
rect 6327 600 6369 654
rect 6223 534 6369 600
rect 6223 480 6254 534
rect 6327 480 6369 534
rect 6223 414 6369 480
rect 6223 360 6254 414
rect 6327 360 6369 414
rect 6223 294 6369 360
rect 4958 243 5035 252
rect 4958 184 4967 243
rect 5026 184 5035 243
rect 4958 181 4969 184
rect 5025 181 5035 184
rect 4958 175 5035 181
rect 4968 172 5026 175
rect 4490 118 4582 119
rect 4185 16 4233 27
rect 4417 100 4582 118
rect 4417 97 4693 100
rect 4417 36 4421 97
rect 4482 91 4693 97
rect 5082 98 5164 108
rect 4764 93 5026 95
rect 5082 93 5094 98
rect 4764 91 5094 93
rect 4482 45 4642 91
rect 4688 45 4699 91
rect 4759 45 4770 91
rect 4816 45 4982 91
rect 5028 45 5094 91
rect 4482 44 4693 45
rect 4482 42 4688 44
rect 4764 42 5094 45
rect 5150 93 5164 98
rect 5428 97 5481 267
rect 6223 240 6254 294
rect 6327 240 6369 294
rect 6223 174 6369 240
rect 6223 120 6254 174
rect 6327 120 6369 174
rect 5318 93 5580 97
rect 5739 93 5793 96
rect 5150 91 5239 93
rect 5318 91 5793 93
rect 5150 45 5194 91
rect 5240 45 5251 91
rect 5311 45 5322 91
rect 5368 45 5534 91
rect 5580 45 5746 91
rect 5792 45 5803 91
rect 6223 54 6369 120
rect 5150 42 5239 45
rect 5318 44 5580 45
rect 4482 36 4492 42
rect 4977 40 5239 42
rect 4417 22 4492 36
rect 5082 34 5164 40
rect 3966 -60 4045 -50
rect 3966 -116 3977 -60
rect 4033 -116 4045 -60
rect 5435 -102 5487 44
rect 5739 -27 5793 45
rect 5618 -28 5793 -27
rect 6223 0 6254 54
rect 6327 0 6369 54
rect 5618 -36 5797 -28
rect 5618 -82 5627 -36
rect 5699 -82 5797 -36
rect 5618 -90 5797 -82
rect 6223 -66 6369 0
rect 5618 -91 5708 -90
rect 3966 -130 4045 -116
rect 5190 -154 5487 -102
rect 3369 -257 3421 -237
rect 3213 -351 3215 -316
rect 2961 -363 3215 -351
rect 3369 -351 3371 -257
rect 3417 -351 3421 -257
rect 2961 -536 3009 -363
rect 2961 -630 2963 -536
rect 2961 -642 3009 -630
rect 3167 -536 3213 -363
rect 3167 -641 3213 -630
rect 3369 -536 3421 -351
rect 3369 -630 3371 -536
rect 3417 -630 3421 -536
rect 3572 -257 3622 -241
rect 3572 -351 3575 -257
rect 3621 -351 3622 -257
rect 3572 -536 3622 -351
rect 3572 -624 3575 -536
rect 3369 -642 3421 -630
rect 3558 -630 3575 -624
rect 3621 -624 3622 -536
rect 3775 -257 3828 -237
rect 3775 -351 3779 -257
rect 3825 -351 3828 -257
rect 3962 -231 4061 -220
rect 4424 -225 4478 -221
rect 4637 -225 4691 -217
rect 4767 -225 4819 -224
rect 4976 -225 5032 -224
rect 5190 -225 5242 -154
rect 5435 -155 5487 -154
rect 6223 -120 6254 -66
rect 6327 -120 6369 -66
rect 6223 -186 6369 -120
rect 5318 -225 5370 -220
rect 5531 -225 5583 -222
rect 5736 -225 5799 -216
rect 3962 -232 4062 -231
rect 3962 -293 3973 -232
rect 4034 -293 4062 -232
rect 4187 -247 4233 -246
rect 3962 -301 3983 -293
rect 3972 -302 3983 -301
rect 3775 -536 3828 -351
rect 3621 -630 3633 -624
rect 3558 -634 3633 -630
rect 2654 -748 2678 -694
rect 2751 -748 2775 -694
rect 2654 -814 2775 -748
rect 2654 -868 2678 -814
rect 2751 -868 2775 -814
rect 3150 -782 3229 -770
rect 3150 -836 3161 -782
rect 3215 -836 3229 -782
rect 3150 -848 3229 -836
rect 2654 -934 2775 -868
rect 3165 -903 3211 -848
rect 3369 -902 3417 -642
rect 3558 -688 3570 -634
rect 3624 -688 3633 -634
rect 3775 -630 3779 -536
rect 3825 -630 3828 -536
rect 3775 -642 3828 -630
rect 3558 -700 3633 -688
rect 3556 -789 3636 -777
rect 3556 -843 3569 -789
rect 3623 -843 3636 -789
rect 3556 -855 3636 -843
rect 2654 -988 2678 -934
rect 2751 -988 2775 -934
rect 2654 -1054 2775 -988
rect 2963 -906 3009 -903
rect 2963 -914 3012 -906
rect 3009 -1008 3012 -914
rect 2963 -1019 3012 -1008
rect 2654 -1108 2678 -1054
rect 2751 -1108 2775 -1054
rect 2437 -1132 2516 -1123
rect 2437 -1193 2446 -1132
rect 2507 -1193 2516 -1132
rect 2437 -1202 2516 -1193
rect 2654 -1174 2775 -1108
rect 2964 -1100 3012 -1019
rect 3165 -914 3213 -903
rect 3165 -1008 3167 -914
rect 3165 -1019 3213 -1008
rect 3370 -914 3417 -902
rect 3370 -1008 3371 -914
rect 3370 -1019 3417 -1008
rect 3573 -903 3619 -855
rect 3573 -914 3621 -903
rect 3573 -1008 3575 -914
rect 3573 -1019 3621 -1008
rect 3778 -914 3828 -642
rect 3981 -351 3983 -302
rect 4029 -306 4062 -293
rect 4186 -257 4233 -247
rect 4029 -351 4031 -306
rect 3981 -400 4031 -351
rect 4186 -351 4187 -257
rect 4418 -271 4429 -225
rect 4475 -271 4486 -225
rect 4630 -271 4641 -225
rect 4687 -271 4698 -225
rect 4758 -271 4769 -225
rect 4815 -271 4826 -225
rect 4970 -271 4981 -225
rect 5027 -271 5038 -225
rect 5182 -271 5193 -225
rect 5239 -271 5250 -225
rect 5310 -271 5321 -225
rect 5367 -271 5378 -225
rect 5522 -271 5533 -225
rect 5579 -271 5590 -225
rect 5734 -271 5745 -225
rect 5791 -271 5802 -225
rect 6223 -240 6254 -186
rect 6327 -240 6369 -186
rect 4186 -400 4233 -351
rect 3981 -409 4233 -400
rect 3981 -459 4072 -409
rect 4144 -459 4233 -409
rect 3981 -468 4233 -459
rect 3981 -536 4031 -468
rect 3981 -630 3983 -536
rect 4029 -630 4031 -536
rect 3981 -646 4031 -630
rect 4186 -536 4233 -468
rect 4424 -336 4478 -271
rect 4637 -336 4691 -271
rect 4424 -390 4691 -336
rect 4424 -475 4478 -390
rect 4637 -475 4691 -390
rect 4767 -344 4819 -271
rect 4976 -344 5032 -271
rect 5190 -344 5242 -271
rect 5318 -342 5370 -271
rect 5531 -320 5583 -271
rect 5736 -320 5799 -271
rect 5531 -329 5799 -320
rect 5531 -342 5626 -329
rect 4767 -396 5244 -344
rect 5318 -376 5626 -342
rect 5698 -376 5799 -329
rect 5318 -385 5799 -376
rect 5318 -394 5583 -385
rect 4767 -475 4819 -396
rect 4976 -475 5032 -396
rect 5190 -475 5242 -396
rect 5318 -475 5370 -394
rect 5531 -467 5583 -394
rect 5527 -475 5583 -467
rect 5736 -475 5799 -385
rect 6223 -306 6369 -240
rect 6223 -360 6254 -306
rect 6327 -360 6369 -306
rect 6223 -426 6369 -360
rect 4418 -521 4429 -475
rect 4475 -521 4486 -475
rect 4630 -521 4641 -475
rect 4687 -521 4698 -475
rect 4758 -521 4769 -475
rect 4815 -521 4826 -475
rect 4970 -521 4981 -475
rect 5027 -521 5038 -475
rect 5182 -521 5193 -475
rect 5239 -521 5250 -475
rect 5310 -521 5321 -475
rect 5367 -521 5378 -475
rect 5522 -521 5533 -475
rect 5579 -521 5590 -475
rect 5734 -521 5745 -475
rect 5791 -521 5802 -475
rect 6223 -480 6254 -426
rect 6327 -480 6369 -426
rect 4424 -526 4478 -521
rect 4186 -630 4187 -536
rect 4186 -697 4233 -630
rect 4637 -618 4691 -521
rect 4767 -526 4819 -521
rect 4976 -534 5032 -521
rect 5190 -526 5242 -521
rect 5318 -522 5370 -521
rect 5527 -524 5583 -521
rect 4637 -630 4740 -618
rect 5527 -630 5581 -524
rect 5736 -527 5799 -521
rect 4637 -684 4672 -630
rect 4660 -686 4672 -684
rect 4728 -684 5581 -630
rect 6223 -546 6369 -480
rect 6223 -600 6254 -546
rect 6327 -600 6369 -546
rect 6223 -666 6369 -600
rect 4728 -686 4740 -684
rect 4660 -689 4740 -686
rect 4186 -744 4479 -697
rect 3966 -759 4044 -747
rect 3966 -813 3978 -759
rect 4032 -813 4044 -759
rect 4432 -792 4479 -744
rect 3966 -824 4044 -813
rect 4417 -800 4698 -792
rect 4894 -793 4947 -684
rect 5186 -690 5306 -684
rect 6223 -720 6254 -666
rect 6327 -720 6369 -666
rect 6223 -786 6369 -720
rect 4765 -795 5027 -793
rect 5080 -794 5164 -787
rect 5080 -795 5095 -794
rect 4765 -800 5095 -795
rect 3778 -1008 3779 -914
rect 3825 -1008 3828 -914
rect 3165 -1100 3211 -1019
rect 3370 -1020 3416 -1019
rect 3573 -1020 3619 -1019
rect 3778 -1022 3828 -1008
rect 3982 -891 4028 -824
rect 4417 -846 4429 -800
rect 4475 -846 4641 -800
rect 4687 -846 4698 -800
rect 4758 -846 4769 -800
rect 4815 -846 4981 -800
rect 5027 -846 5095 -800
rect 3982 -914 4029 -891
rect 4187 -904 4233 -903
rect 4186 -914 4233 -904
rect 3982 -1008 3983 -914
rect 4029 -1008 4030 -914
rect 3982 -1021 4030 -1008
rect 2964 -1115 3211 -1100
rect 2964 -1170 3050 -1115
rect -1973 -1295 1736 -1247
rect -1762 -1374 -1709 -1362
rect -1762 -1468 -1759 -1374
rect -1713 -1468 -1709 -1374
rect -1762 -1538 -1709 -1468
rect -1559 -1374 -1506 -1358
rect -1559 -1468 -1555 -1374
rect -1509 -1468 -1506 -1374
rect -1559 -1538 -1506 -1468
rect -1373 -1374 -1325 -1360
rect -1373 -1468 -1372 -1374
rect -1326 -1468 -1325 -1374
rect -1373 -1532 -1325 -1468
rect -1169 -1374 -1121 -1295
rect -1169 -1468 -1168 -1374
rect -1122 -1468 -1121 -1374
rect -1762 -1547 -1506 -1538
rect -1762 -1548 -1670 -1547
rect -1762 -1604 -1756 -1548
rect -1700 -1604 -1670 -1548
rect -1762 -1619 -1670 -1604
rect -1598 -1559 -1506 -1547
rect -1388 -1544 -1310 -1532
rect -1388 -1559 -1376 -1544
rect -1598 -1598 -1376 -1559
rect -1322 -1598 -1310 -1544
rect -1598 -1607 -1310 -1598
rect -1598 -1619 -1506 -1607
rect -1388 -1611 -1310 -1607
rect -1762 -1628 -1506 -1619
rect -1762 -1684 -1709 -1628
rect -1762 -1778 -1759 -1684
rect -1713 -1778 -1709 -1684
rect -1762 -1793 -1709 -1778
rect -1559 -1684 -1506 -1628
rect -1559 -1778 -1555 -1684
rect -1509 -1778 -1506 -1684
rect -1559 -1789 -1506 -1778
rect -1373 -1684 -1325 -1611
rect -1373 -1778 -1372 -1684
rect -1326 -1778 -1325 -1684
rect -1373 -1791 -1325 -1778
rect -1169 -1684 -1121 -1468
rect -1169 -1778 -1168 -1684
rect -1122 -1778 -1121 -1684
rect -1169 -1791 -1121 -1778
rect -965 -1374 -917 -1362
rect -965 -1468 -964 -1374
rect -918 -1468 -917 -1374
rect -965 -1684 -917 -1468
rect -965 -1778 -964 -1684
rect -918 -1778 -917 -1684
rect -965 -1990 -917 -1778
rect -762 -1374 -714 -1295
rect -762 -1468 -760 -1374
rect -762 -1684 -714 -1468
rect -557 -1374 -509 -1362
rect -352 -1363 -304 -1295
rect -557 -1468 -556 -1374
rect -510 -1468 -509 -1374
rect -557 -1531 -509 -1468
rect -353 -1374 -304 -1363
rect -148 -1365 -102 -1363
rect -353 -1468 -352 -1374
rect -306 -1468 -304 -1374
rect -564 -1543 -505 -1531
rect -564 -1599 -562 -1543
rect -506 -1599 -505 -1543
rect -564 -1611 -505 -1599
rect -762 -1778 -760 -1684
rect -762 -1791 -714 -1778
rect -557 -1684 -509 -1611
rect -557 -1778 -556 -1684
rect -510 -1778 -509 -1684
rect -557 -1793 -509 -1778
rect -353 -1684 -304 -1468
rect -353 -1778 -352 -1684
rect -306 -1778 -304 -1684
rect -353 -1794 -304 -1778
rect -149 -1374 -101 -1365
rect -149 -1468 -148 -1374
rect -102 -1468 -101 -1374
rect -149 -1684 -101 -1468
rect -149 -1778 -148 -1684
rect -102 -1778 -101 -1684
rect -149 -1990 -101 -1778
rect 54 -1374 102 -1295
rect 54 -1468 56 -1374
rect 54 -1684 102 -1468
rect 259 -1374 307 -1361
rect 464 -1363 512 -1295
rect 873 -1362 921 -1295
rect 259 -1468 260 -1374
rect 306 -1468 307 -1374
rect 259 -1531 307 -1468
rect 463 -1374 512 -1363
rect 463 -1468 464 -1374
rect 510 -1468 512 -1374
rect 463 -1479 512 -1468
rect 666 -1374 714 -1362
rect 666 -1468 668 -1374
rect 252 -1543 315 -1531
rect 252 -1599 255 -1543
rect 311 -1599 315 -1543
rect 252 -1612 315 -1599
rect 54 -1778 56 -1684
rect 54 -1792 102 -1778
rect 259 -1684 307 -1612
rect 259 -1778 260 -1684
rect 306 -1778 307 -1684
rect 259 -1792 307 -1778
rect 463 -1684 511 -1479
rect 463 -1778 464 -1684
rect 510 -1778 511 -1684
rect 463 -1794 511 -1778
rect 666 -1684 714 -1468
rect 666 -1778 668 -1684
rect 666 -1990 714 -1778
rect 871 -1374 921 -1362
rect 871 -1468 872 -1374
rect 918 -1468 921 -1374
rect 871 -1484 921 -1468
rect 1075 -1374 1123 -1360
rect 1075 -1468 1076 -1374
rect 1122 -1468 1123 -1374
rect 871 -1684 919 -1484
rect 1075 -1531 1123 -1468
rect 1279 -1374 1327 -1295
rect 1688 -1361 1736 -1295
rect 1484 -1364 1530 -1363
rect 1279 -1468 1280 -1374
rect 1326 -1468 1327 -1374
rect 1066 -1543 1130 -1531
rect 1066 -1599 1071 -1543
rect 1127 -1599 1130 -1543
rect 1066 -1611 1130 -1599
rect 871 -1778 872 -1684
rect 918 -1778 919 -1684
rect 871 -1793 919 -1778
rect 1075 -1684 1123 -1611
rect 1075 -1778 1076 -1684
rect 1122 -1778 1123 -1684
rect 1075 -1791 1123 -1778
rect 1279 -1684 1327 -1468
rect 1279 -1778 1280 -1684
rect 1326 -1778 1327 -1684
rect 1279 -1792 1327 -1778
rect 1483 -1374 1531 -1364
rect 1483 -1468 1484 -1374
rect 1530 -1468 1531 -1374
rect 1483 -1684 1531 -1468
rect 1483 -1778 1484 -1684
rect 1530 -1778 1531 -1684
rect 1483 -1990 1531 -1778
rect 1687 -1374 1736 -1361
rect 1687 -1468 1688 -1374
rect 1734 -1468 1736 -1374
rect 1687 -1479 1736 -1468
rect 1891 -1374 1939 -1361
rect 1891 -1468 1892 -1374
rect 1938 -1468 1939 -1374
rect 1687 -1684 1735 -1479
rect 1891 -1531 1939 -1468
rect 2067 -1374 2115 -1361
rect 2067 -1468 2069 -1374
rect 2067 -1524 2115 -1468
rect 2272 -1374 2320 -1362
rect 2272 -1468 2273 -1374
rect 2319 -1468 2320 -1374
rect 2272 -1524 2320 -1468
rect 1883 -1536 1950 -1531
rect 2067 -1536 2320 -1524
rect 1883 -1538 2320 -1536
rect 1883 -1543 2158 -1538
rect 1883 -1599 1885 -1543
rect 1941 -1583 2158 -1543
rect 1941 -1599 1950 -1583
rect 1883 -1612 1950 -1599
rect 2067 -1584 2158 -1583
rect 2230 -1584 2320 -1538
rect 2067 -1597 2320 -1584
rect 1687 -1778 1688 -1684
rect 1734 -1778 1735 -1684
rect 1687 -1792 1735 -1778
rect 1891 -1684 1939 -1612
rect 1891 -1778 1892 -1684
rect 1938 -1778 1939 -1684
rect 1891 -1792 1939 -1778
rect 2067 -1684 2115 -1597
rect 2067 -1778 2069 -1684
rect 2067 -1792 2115 -1778
rect 2272 -1684 2320 -1597
rect 2272 -1778 2273 -1684
rect 2319 -1778 2320 -1684
rect 2272 -1793 2320 -1778
rect 2451 -1864 2510 -1202
rect 2654 -1228 2678 -1174
rect 2751 -1228 2775 -1174
rect 3036 -1192 3050 -1170
rect 3127 -1172 3211 -1115
rect 3983 -1063 4030 -1021
rect 4186 -1008 4187 -914
rect 4186 -1063 4233 -1008
rect 4557 -1053 4610 -846
rect 4977 -848 5095 -846
rect 5149 -795 5164 -794
rect 5311 -795 5581 -793
rect 5149 -800 5239 -795
rect 5311 -800 5592 -795
rect 5149 -846 5193 -800
rect 5239 -846 5250 -800
rect 5310 -846 5321 -800
rect 5367 -846 5533 -800
rect 5579 -846 5592 -800
rect 5734 -846 5745 -800
rect 5791 -846 5802 -800
rect 6223 -840 6254 -786
rect 6327 -840 6369 -786
rect 5149 -848 5239 -846
rect 5080 -855 5164 -848
rect 4950 -928 5028 -919
rect 4784 -930 4863 -928
rect 4784 -984 4796 -930
rect 4850 -934 4863 -930
rect 4950 -934 4959 -928
rect 4850 -980 4959 -934
rect 4850 -984 4863 -980
rect 4784 -995 4863 -984
rect 4950 -988 4959 -980
rect 5019 -988 5028 -928
rect 4950 -997 5028 -988
rect 5410 -1053 5463 -846
rect 5531 -892 5592 -846
rect 5742 -892 5794 -846
rect 5531 -893 5794 -892
rect 5531 -901 5800 -893
rect 5531 -950 5626 -901
rect 5698 -950 5800 -901
rect 5531 -957 5800 -950
rect 6223 -906 6369 -840
rect 5617 -959 5707 -957
rect 3983 -1072 4245 -1063
rect 3983 -1124 4170 -1072
rect 4236 -1124 4245 -1072
rect 4557 -1106 5463 -1053
rect 6223 -960 6254 -906
rect 6327 -960 6369 -906
rect 6223 -1026 6369 -960
rect 6223 -1080 6254 -1026
rect 6327 -1080 6369 -1026
rect 3983 -1129 4245 -1124
rect 3127 -1184 3227 -1172
rect 3127 -1192 3161 -1184
rect 3036 -1205 3161 -1192
rect 2654 -1294 2775 -1228
rect 3149 -1238 3161 -1205
rect 3215 -1190 3227 -1184
rect 3983 -1190 4029 -1129
rect 4161 -1133 4245 -1129
rect 6223 -1146 6369 -1080
rect 4661 -1186 4738 -1174
rect 4661 -1190 4673 -1186
rect 3215 -1236 4673 -1190
rect 3215 -1238 3227 -1236
rect 3149 -1250 3227 -1238
rect 4661 -1240 4673 -1236
rect 4727 -1240 4738 -1186
rect 4661 -1252 4738 -1240
rect 6223 -1200 6254 -1146
rect 6327 -1200 6369 -1146
rect 2654 -1348 2678 -1294
rect 2751 -1348 2775 -1294
rect 6223 -1266 6369 -1200
rect 2654 -1414 2775 -1348
rect 3853 -1330 3943 -1319
rect 3853 -1402 3868 -1330
rect 3933 -1402 3943 -1330
rect 3853 -1411 3943 -1402
rect 6223 -1320 6254 -1266
rect 6327 -1320 6369 -1266
rect 6223 -1386 6369 -1320
rect 2654 -1468 2678 -1414
rect 2751 -1468 2775 -1414
rect 2654 -1545 2775 -1468
rect 6223 -1440 6254 -1386
rect 6327 -1440 6369 -1386
rect 6223 -1545 6369 -1440
rect 2654 -1546 6369 -1545
rect 2654 -1547 6457 -1546
rect 2652 -1564 6457 -1547
rect 2652 -1618 2681 -1564
rect 2754 -1618 2806 -1564
rect 2879 -1618 2931 -1564
rect 3004 -1618 3056 -1564
rect 3129 -1618 3181 -1564
rect 3254 -1565 6457 -1564
rect 3254 -1614 3318 -1565
rect 3381 -1566 6229 -1565
rect 3381 -1614 3439 -1566
rect 3254 -1615 3439 -1614
rect 3502 -1615 3560 -1566
rect 3623 -1615 3681 -1566
rect 3744 -1615 3802 -1566
rect 3865 -1615 3923 -1566
rect 3986 -1615 4044 -1566
rect 4107 -1615 4165 -1566
rect 4228 -1615 4286 -1566
rect 4349 -1615 4407 -1566
rect 4470 -1615 4528 -1566
rect 4591 -1615 4649 -1566
rect 4712 -1615 4770 -1566
rect 4833 -1615 4891 -1566
rect 4954 -1615 5012 -1566
rect 5075 -1615 5133 -1566
rect 5196 -1615 5254 -1566
rect 5317 -1615 5375 -1566
rect 5438 -1615 5496 -1566
rect 5559 -1615 5617 -1566
rect 5680 -1615 5738 -1566
rect 5801 -1615 5859 -1566
rect 5922 -1615 5980 -1566
rect 6043 -1615 6101 -1566
rect 6164 -1614 6229 -1566
rect 6292 -1576 6457 -1565
rect 6292 -1584 6458 -1576
rect 6292 -1614 6375 -1584
rect 6164 -1615 6375 -1614
rect 3254 -1618 6375 -1615
rect 2652 -1631 6375 -1618
rect 2652 -1641 3339 -1631
rect 3231 -1760 3339 -1641
rect 6350 -1633 6375 -1631
rect 6438 -1633 6458 -1584
rect 3231 -1809 3255 -1760
rect 3318 -1809 3339 -1760
rect 3798 -1690 3888 -1678
rect 3798 -1758 3805 -1690
rect 3873 -1707 3888 -1690
rect 3879 -1756 3888 -1707
rect 6350 -1691 6458 -1633
rect 3873 -1758 3888 -1756
rect 3798 -1770 3888 -1758
rect 4990 -1783 5702 -1733
rect 2442 -1873 2518 -1864
rect 2442 -1931 2451 -1873
rect 2509 -1931 2518 -1873
rect 2442 -1940 2518 -1931
rect 3231 -1871 3339 -1809
rect 3594 -1807 3684 -1798
rect 3594 -1815 3603 -1807
rect 3524 -1827 3603 -1815
rect 3524 -1838 3536 -1827
rect 3231 -1920 3255 -1871
rect 3318 -1920 3339 -1871
rect 3231 -1982 3339 -1920
rect -1374 -2014 2012 -1990
rect -1374 -2029 1939 -2014
rect -1374 -2080 -1162 -2029
rect 1713 -2076 1939 -2029
rect 2001 -2076 2012 -2014
rect 1713 -2080 2012 -2076
rect -1374 -2117 2012 -2080
rect 3231 -2031 3255 -1982
rect 3318 -2031 3339 -1982
rect 3231 -2093 3339 -2031
rect 3513 -1883 3536 -1838
rect 3592 -1856 3603 -1827
rect 3675 -1838 3684 -1807
rect 3675 -1856 3972 -1838
rect 3592 -1883 3972 -1856
rect 3513 -1889 3972 -1883
rect 3513 -1895 3600 -1889
rect 3513 -1919 3564 -1895
rect 3513 -2013 3514 -1919
rect 3560 -2013 3564 -1919
rect 3513 -2040 3564 -2013
rect 3718 -1919 3769 -1889
rect 3764 -2013 3769 -1919
rect 3718 -2030 3769 -2013
rect 3920 -1919 3972 -1889
rect 4044 -1845 4127 -1836
rect 4786 -1841 4836 -1839
rect 4990 -1841 5040 -1783
rect 5463 -1830 5543 -1829
rect 5463 -1838 5475 -1830
rect 4254 -1845 4304 -1844
rect 4456 -1845 4506 -1844
rect 4044 -1901 4058 -1845
rect 4114 -1895 4506 -1845
rect 4114 -1901 4127 -1895
rect 4044 -1906 4127 -1901
rect 3920 -2013 3922 -1919
rect 3968 -2013 3972 -1919
rect 476 -2522 534 -2117
rect 3231 -2142 3255 -2093
rect 3318 -2142 3339 -2093
rect 3231 -2204 3339 -2142
rect 3920 -2126 3972 -2013
rect 4048 -1919 4098 -1906
rect 4048 -2013 4050 -1919
rect 4096 -2013 4098 -1919
rect 4048 -2030 4098 -2013
rect 4254 -1919 4304 -1895
rect 4300 -2013 4304 -1919
rect 4254 -2030 4304 -2013
rect 4456 -1919 4506 -1895
rect 4456 -2013 4458 -1919
rect 4504 -2013 4506 -1919
rect 4456 -2032 4506 -2013
rect 4585 -1891 5040 -1841
rect 4585 -1919 4635 -1891
rect 4585 -2013 4586 -1919
rect 4632 -2013 4635 -1919
rect 4585 -2026 4635 -2013
rect 4786 -1919 4836 -1891
rect 4786 -2013 4790 -1919
rect 4786 -2026 4836 -2013
rect 4990 -1919 5040 -1891
rect 5119 -1886 5475 -1838
rect 5531 -1837 5543 -1830
rect 5652 -1834 5702 -1783
rect 6350 -1740 6375 -1691
rect 6438 -1740 6458 -1691
rect 6350 -1791 6458 -1740
rect 5859 -1819 6111 -1810
rect 5859 -1834 5951 -1819
rect 5531 -1886 5578 -1837
rect 5119 -1888 5578 -1886
rect 5119 -1907 5169 -1888
rect 4990 -2013 4994 -1919
rect 4990 -2022 5040 -2013
rect 4994 -2024 5040 -2022
rect 5117 -1919 5169 -1907
rect 5117 -2013 5122 -1919
rect 5168 -2013 5169 -1919
rect 5117 -2031 5169 -2013
rect 5324 -1919 5374 -1888
rect 5463 -1896 5578 -1888
rect 5324 -2013 5326 -1919
rect 5372 -2013 5374 -1919
rect 5324 -2026 5374 -2013
rect 5528 -1919 5578 -1896
rect 5528 -2013 5530 -1919
rect 5576 -2013 5578 -1919
rect 5528 -2025 5578 -2013
rect 5652 -1869 5951 -1834
rect 6023 -1869 6111 -1819
rect 5652 -1878 6111 -1869
rect 5652 -1884 5910 -1878
rect 5652 -1919 5704 -1884
rect 5652 -2013 5658 -1919
rect 5652 -2015 5704 -2013
rect 4231 -2115 4325 -2106
rect 3920 -2178 4094 -2126
rect 3231 -2253 3255 -2204
rect 3318 -2253 3339 -2204
rect 3231 -2315 3339 -2253
rect 3514 -2293 3560 -2292
rect 3231 -2364 3255 -2315
rect 3318 -2364 3339 -2315
rect 3231 -2426 3339 -2364
rect 3231 -2475 3255 -2426
rect 3318 -2475 3339 -2426
rect -280 -2548 2839 -2522
rect -280 -2549 502 -2548
rect -280 -2598 -236 -2549
rect -173 -2550 21 -2549
rect -173 -2598 -108 -2550
rect -280 -2599 -108 -2598
rect -45 -2598 21 -2550
rect 84 -2550 373 -2549
rect 84 -2598 138 -2550
rect -45 -2599 138 -2598
rect 201 -2551 373 -2550
rect 201 -2599 250 -2551
rect -280 -2600 250 -2599
rect 313 -2598 373 -2551
rect 436 -2597 502 -2549
rect 565 -2549 1104 -2548
rect 565 -2597 619 -2549
rect 436 -2598 619 -2597
rect 682 -2550 975 -2549
rect 682 -2598 731 -2550
rect 313 -2599 731 -2598
rect 794 -2599 849 -2550
rect 912 -2598 975 -2550
rect 1038 -2597 1104 -2549
rect 1167 -2549 2839 -2548
rect 1167 -2597 1221 -2549
rect 1038 -2598 1221 -2597
rect 1284 -2550 2839 -2549
rect 1284 -2598 1333 -2550
rect 912 -2599 1333 -2598
rect 1396 -2599 1451 -2550
rect 1514 -2599 1574 -2550
rect 1637 -2599 1691 -2550
rect 1754 -2599 1812 -2550
rect 1875 -2599 1934 -2550
rect 1997 -2551 2516 -2550
rect 1997 -2599 2045 -2551
rect 313 -2600 2045 -2599
rect 2108 -2600 2164 -2551
rect 2227 -2600 2276 -2551
rect 2339 -2600 2397 -2551
rect 2460 -2599 2516 -2551
rect 2579 -2552 2742 -2550
rect 2579 -2599 2631 -2552
rect 2460 -2600 2631 -2599
rect -280 -2601 2631 -2600
rect 2694 -2599 2742 -2552
rect 2805 -2599 2839 -2550
rect 2694 -2601 2839 -2599
rect -280 -2634 2839 -2601
rect -280 -2664 -170 -2634
rect -280 -2711 -250 -2664
rect -196 -2711 -170 -2664
rect -280 -2765 -170 -2711
rect 2724 -2650 2839 -2634
rect 2724 -2697 2753 -2650
rect 2807 -2697 2839 -2650
rect 1014 -2747 1068 -2744
rect -280 -2812 -249 -2765
rect -195 -2812 -170 -2765
rect -280 -2862 -170 -2812
rect -2492 -2885 -2356 -2874
rect -2144 -2885 -784 -2870
rect -2492 -2886 -784 -2885
rect -2492 -2966 -2482 -2886
rect -2399 -2909 -784 -2886
rect -2399 -2914 -1551 -2909
rect -2399 -2965 -2084 -2914
rect -1834 -2955 -1551 -2914
rect -839 -2955 -784 -2909
rect -1834 -2965 -784 -2955
rect -2399 -2966 -784 -2965
rect -2492 -2967 -784 -2966
rect -2492 -2979 -2356 -2967
rect -2144 -2983 -784 -2967
rect -280 -2909 -250 -2862
rect -196 -2909 -170 -2862
rect 350 -2801 1068 -2747
rect 2724 -2751 2839 -2697
rect 2079 -2763 2155 -2752
rect -280 -2970 -170 -2909
rect -2068 -3075 -1998 -2983
rect -2068 -3149 -2045 -3075
rect -1999 -3149 -1998 -3075
rect -2068 -3164 -1998 -3149
rect -1886 -3075 -1822 -3062
rect -1886 -3149 -1885 -3075
rect -1839 -3149 -1822 -3075
rect -1704 -3069 -1617 -3051
rect -1704 -3134 -1691 -3069
rect -1626 -3107 -1617 -3069
rect -1626 -3110 -1452 -3107
rect -1626 -3134 -1509 -3110
rect -1704 -3136 -1509 -3134
rect -2290 -3238 -1940 -3230
rect -2290 -3285 -2015 -3238
rect -2290 -3311 -2142 -3285
rect -2167 -3343 -2142 -3311
rect -2084 -3297 -2015 -3285
rect -1952 -3297 -1940 -3238
rect -2084 -3311 -1940 -3297
rect -1886 -3265 -1822 -3149
rect -1698 -3156 -1509 -3136
rect -1463 -3156 -1452 -3110
rect -1698 -3158 -1452 -3156
rect -1354 -3110 -1283 -2983
rect -1354 -3156 -1341 -3110
rect -1295 -3156 -1283 -3110
rect -1354 -3158 -1283 -3156
rect -1109 -3110 -1038 -2983
rect -576 -3005 -473 -2992
rect -732 -3006 -473 -3005
rect -732 -3019 -569 -3006
rect -732 -3079 -719 -3019
rect -656 -3079 -569 -3019
rect -732 -3091 -569 -3079
rect -484 -3091 -473 -3006
rect -732 -3092 -473 -3091
rect -576 -3106 -473 -3092
rect -280 -3017 -249 -2970
rect -195 -3017 -170 -2970
rect -280 -3095 -170 -3017
rect -1109 -3156 -1097 -3110
rect -1051 -3156 -1038 -3110
rect -1109 -3158 -1038 -3156
rect -940 -3110 -809 -3109
rect -940 -3156 -929 -3110
rect -883 -3156 -809 -3110
rect -940 -3158 -809 -3156
rect -1698 -3178 -1513 -3158
rect -2084 -3343 -2070 -3311
rect -2167 -3346 -2070 -3343
rect -1886 -3312 -1685 -3265
rect -2071 -3413 -1990 -3408
rect -1886 -3413 -1822 -3312
rect -1732 -3368 -1685 -3312
rect -1732 -3382 -1642 -3368
rect -1732 -3396 -1718 -3382
rect -2071 -3459 -2049 -3413
rect -2003 -3459 -1990 -3413
rect -1892 -3459 -1881 -3413
rect -1835 -3459 -1822 -3413
rect -1731 -3442 -1718 -3396
rect -1655 -3442 -1642 -3382
rect -1731 -3455 -1642 -3442
rect -1584 -3415 -1513 -3178
rect -1441 -3223 -1352 -3210
rect -1441 -3283 -1428 -3223
rect -1365 -3283 -1352 -3223
rect -1441 -3297 -1352 -3283
rect -878 -3227 -809 -3158
rect -280 -3142 -249 -3095
rect -195 -3142 -170 -3095
rect -280 -3209 -170 -3142
rect -878 -3286 -869 -3227
rect -817 -3230 -809 -3227
rect -626 -3230 -536 -3219
rect -817 -3286 -617 -3230
rect -878 -3298 -617 -3286
rect -549 -3298 -536 -3230
rect -878 -3415 -809 -3298
rect -626 -3313 -536 -3298
rect -280 -3256 -248 -3209
rect -194 -3256 -170 -3209
rect -2071 -3570 -1990 -3459
rect -1886 -3460 -1822 -3459
rect -1584 -3461 -1571 -3415
rect -1525 -3461 -1513 -3415
rect -1584 -3462 -1513 -3461
rect -1415 -3461 -1403 -3415
rect -1357 -3461 -1343 -3415
rect -1415 -3570 -1343 -3461
rect -1047 -3461 -1035 -3415
rect -989 -3461 -977 -3415
rect -1047 -3570 -977 -3461
rect -878 -3461 -867 -3415
rect -821 -3461 -809 -3415
rect -878 -3462 -809 -3461
rect -280 -3321 -170 -3256
rect -59 -2902 -5 -2887
rect -59 -2996 -54 -2902
rect -8 -2996 -5 -2902
rect -59 -3036 -5 -2996
rect 146 -2902 200 -2880
rect 146 -2996 150 -2902
rect 196 -2996 200 -2902
rect 146 -3036 200 -2996
rect -59 -3051 200 -3036
rect -59 -3100 35 -3051
rect 107 -3052 200 -3051
rect 350 -2902 404 -2801
rect 350 -2996 354 -2902
rect 400 -2996 404 -2902
rect 350 -3052 404 -2996
rect 107 -3100 404 -3052
rect -59 -3108 404 -3100
rect -59 -3113 200 -3108
rect -59 -3186 -5 -3113
rect -59 -3280 -54 -3186
rect -8 -3280 -5 -3186
rect -59 -3293 -5 -3280
rect 146 -3186 200 -3113
rect 146 -3280 150 -3186
rect 196 -3280 200 -3186
rect 350 -3186 404 -3108
rect 350 -3213 354 -3186
rect 146 -3286 200 -3280
rect 332 -3222 354 -3213
rect 400 -3213 404 -3186
rect 473 -2902 530 -2887
rect 686 -2892 732 -2891
rect 473 -2996 482 -2902
rect 528 -2996 530 -2902
rect 473 -3056 530 -2996
rect 677 -2902 732 -2892
rect 677 -2996 686 -2902
rect 677 -3007 732 -2996
rect 885 -2902 942 -2887
rect 885 -2996 890 -2902
rect 936 -2996 942 -2902
rect 677 -3056 731 -3007
rect 885 -3056 942 -2996
rect 473 -3113 942 -3056
rect 473 -3186 530 -3113
rect 400 -3222 415 -3213
rect 332 -3279 346 -3222
rect 403 -3279 415 -3222
rect 332 -3280 354 -3279
rect 400 -3280 415 -3279
rect 332 -3284 415 -3280
rect 473 -3280 482 -3186
rect 528 -3280 530 -3186
rect 150 -3291 196 -3286
rect 350 -3293 404 -3284
rect 473 -3294 530 -3280
rect 677 -3175 731 -3113
rect 677 -3186 732 -3175
rect 677 -3280 686 -3186
rect 677 -3291 732 -3280
rect 885 -3186 942 -3113
rect 885 -3280 890 -3186
rect 936 -3280 942 -3186
rect 885 -3284 942 -3280
rect 1014 -2902 1068 -2801
rect 1420 -2780 2155 -2763
rect 1420 -2817 2089 -2780
rect 1014 -2996 1018 -2902
rect 1064 -2996 1068 -2902
rect 1222 -2902 1268 -2891
rect 1014 -3128 1068 -2996
rect 1217 -2996 1222 -2947
rect 1420 -2902 1474 -2817
rect 2079 -2836 2089 -2817
rect 2145 -2836 2155 -2780
rect 2079 -2849 2155 -2836
rect 2724 -2798 2754 -2751
rect 2808 -2798 2839 -2751
rect 2724 -2848 2839 -2798
rect 1268 -2996 1271 -2947
rect 1217 -3128 1271 -2996
rect 1420 -2996 1426 -2902
rect 1472 -2996 1474 -2902
rect 1420 -3128 1474 -2996
rect 1547 -2902 1601 -2890
rect 1758 -2894 1804 -2891
rect 1547 -2996 1554 -2902
rect 1600 -2996 1601 -2902
rect 1547 -3065 1601 -2996
rect 1757 -2902 1808 -2894
rect 1757 -2996 1758 -2902
rect 1804 -2996 1808 -2902
rect 1757 -3050 1808 -2996
rect 1961 -2902 2014 -2891
rect 1961 -2996 1962 -2902
rect 2008 -2996 2014 -2902
rect 1748 -3064 1824 -3050
rect 1748 -3065 1757 -3064
rect 1547 -3119 1757 -3065
rect 1014 -3182 1478 -3128
rect 1014 -3186 1068 -3182
rect 1014 -3280 1018 -3186
rect 1064 -3280 1068 -3186
rect 890 -3291 936 -3284
rect -280 -3368 -247 -3321
rect -193 -3368 -170 -3321
rect -280 -3425 -170 -3368
rect -730 -3477 -641 -3463
rect -730 -3537 -717 -3477
rect -654 -3537 -641 -3477
rect -730 -3550 -641 -3537
rect -280 -3472 -249 -3425
rect -195 -3472 -170 -3425
rect 677 -3436 731 -3291
rect 1014 -3356 1068 -3280
rect 1217 -3186 1271 -3182
rect 1217 -3280 1222 -3186
rect 1268 -3280 1271 -3186
rect 1217 -3353 1271 -3280
rect 1420 -3186 1474 -3182
rect 1420 -3280 1426 -3186
rect 1472 -3280 1474 -3186
rect 1420 -3353 1474 -3280
rect 1547 -3186 1601 -3119
rect 1748 -3120 1757 -3119
rect 1813 -3065 1824 -3064
rect 1961 -3065 2014 -2996
rect 2088 -2902 2141 -2849
rect 2294 -2892 2340 -2891
rect 2088 -2996 2090 -2902
rect 2136 -2996 2141 -2902
rect 2088 -3055 2141 -2996
rect 2290 -2902 2343 -2892
rect 2498 -2893 2544 -2891
rect 2290 -2996 2294 -2902
rect 2340 -2996 2343 -2902
rect 2290 -3049 2343 -2996
rect 2496 -2902 2549 -2893
rect 2496 -2996 2498 -2902
rect 2544 -2996 2549 -2902
rect 2496 -3049 2549 -2996
rect 2290 -3055 2549 -3049
rect 2088 -3063 2549 -3055
rect 1813 -3119 2017 -3065
rect 2088 -3108 2383 -3063
rect 1813 -3120 1824 -3119
rect 1748 -3132 1824 -3120
rect 1547 -3280 1554 -3186
rect 1600 -3280 1601 -3186
rect 1547 -3296 1601 -3280
rect 1757 -3186 1808 -3132
rect 1757 -3280 1758 -3186
rect 1804 -3280 1808 -3186
rect 1757 -3436 1808 -3280
rect 1961 -3186 2014 -3119
rect 1961 -3280 1962 -3186
rect 2008 -3280 2014 -3186
rect 1961 -3291 2014 -3280
rect 2088 -3186 2141 -3108
rect 2088 -3280 2090 -3186
rect 2136 -3280 2141 -3186
rect 2088 -3292 2141 -3280
rect 2290 -3111 2383 -3108
rect 2455 -3111 2549 -3063
rect 2290 -3125 2549 -3111
rect 2290 -3186 2343 -3125
rect 2290 -3280 2294 -3186
rect 2340 -3280 2343 -3186
rect 2290 -3292 2343 -3280
rect 2496 -3186 2549 -3125
rect 2496 -3280 2498 -3186
rect 2544 -3280 2549 -3186
rect 2496 -3293 2549 -3280
rect 2724 -2895 2753 -2848
rect 2807 -2895 2839 -2848
rect 2724 -2956 2839 -2895
rect 2724 -3003 2754 -2956
rect 2808 -3003 2839 -2956
rect 2724 -3081 2839 -3003
rect 2724 -3128 2754 -3081
rect 2808 -3128 2839 -3081
rect 2724 -3195 2839 -3128
rect 2724 -3242 2755 -3195
rect 2809 -3242 2839 -3195
rect 2724 -3307 2839 -3242
rect 1927 -3354 2023 -3344
rect 1927 -3365 1948 -3354
rect 2005 -3365 2023 -3354
rect 1927 -3419 1938 -3365
rect 2007 -3419 2023 -3365
rect 1927 -3434 2023 -3419
rect 2724 -3354 2756 -3307
rect 2810 -3354 2839 -3307
rect 2724 -3411 2839 -3354
rect -280 -3529 -170 -3472
rect -2323 -3592 -2234 -3581
rect -2144 -3592 -784 -3570
rect -2323 -3593 -784 -3592
rect -2323 -3658 -2310 -3593
rect -2245 -3603 -784 -3593
rect -2245 -3605 -1567 -3603
rect -2245 -3654 -2099 -3605
rect -1790 -3649 -1567 -3605
rect -838 -3649 -784 -3603
rect -1790 -3654 -784 -3649
rect -2245 -3658 -784 -3654
rect -2323 -3659 -784 -3658
rect -2323 -3666 -2234 -3659
rect -2144 -3683 -784 -3659
rect -280 -3576 -249 -3529
rect -195 -3576 -170 -3529
rect 148 -3484 1833 -3436
rect 148 -3538 196 -3484
rect -280 -3624 -170 -3576
rect -280 -3671 -251 -3624
rect -197 -3671 -170 -3624
rect -280 -3733 -170 -3671
rect -2459 -3745 -2353 -3736
rect -2144 -3745 -784 -3738
rect -2459 -3827 -2450 -3745
rect -2398 -3777 -784 -3745
rect -2398 -3782 -1551 -3777
rect -2398 -3827 -2084 -3782
rect -2459 -3841 -2353 -3827
rect -2144 -3833 -2084 -3827
rect -1834 -3823 -1551 -3782
rect -839 -3823 -784 -3777
rect -1834 -3833 -784 -3823
rect -2144 -3851 -784 -3833
rect -280 -3780 -250 -3733
rect -196 -3780 -170 -3733
rect -280 -3837 -170 -3780
rect -57 -3547 196 -3538
rect -57 -3595 35 -3547
rect 107 -3595 196 -3547
rect 646 -3548 714 -3536
rect -57 -3604 196 -3595
rect -57 -3718 -6 -3604
rect -57 -3812 -54 -3718
rect -8 -3812 -6 -3718
rect -57 -3826 -6 -3812
rect 148 -3718 196 -3604
rect 148 -3812 150 -3718
rect 148 -3828 196 -3812
rect 347 -3549 714 -3548
rect 347 -3605 647 -3549
rect 703 -3605 714 -3549
rect 842 -3543 932 -3534
rect 842 -3590 851 -3543
rect 923 -3590 932 -3543
rect 842 -3599 932 -3590
rect 347 -3606 714 -3605
rect 347 -3718 405 -3606
rect 646 -3617 714 -3606
rect 663 -3648 714 -3617
rect 663 -3695 809 -3648
rect 347 -3812 354 -3718
rect 400 -3812 405 -3718
rect 558 -3718 607 -3703
rect 347 -3817 405 -3812
rect 308 -3827 405 -3817
rect 544 -3783 558 -3771
rect 604 -3771 607 -3718
rect 761 -3718 809 -3695
rect 604 -3783 616 -3771
rect -2068 -3943 -1998 -3851
rect -2068 -4017 -2045 -3943
rect -1999 -4017 -1998 -3943
rect -2068 -4032 -1998 -4017
rect -1886 -3943 -1822 -3930
rect -1886 -4017 -1885 -3943
rect -1839 -4017 -1822 -3943
rect -1704 -3937 -1617 -3919
rect -1704 -4002 -1691 -3937
rect -1626 -3975 -1617 -3937
rect -1626 -3978 -1452 -3975
rect -1626 -4002 -1509 -3978
rect -1704 -4004 -1509 -4002
rect -2340 -4106 -1940 -4098
rect -2340 -4153 -2015 -4106
rect -2340 -4179 -2142 -4153
rect -2167 -4211 -2142 -4179
rect -2084 -4165 -2015 -4153
rect -1952 -4165 -1940 -4106
rect -2084 -4179 -1940 -4165
rect -1886 -4133 -1822 -4017
rect -1698 -4024 -1509 -4004
rect -1463 -4024 -1452 -3978
rect -1698 -4026 -1452 -4024
rect -1354 -3978 -1283 -3851
rect -1354 -4024 -1341 -3978
rect -1295 -4024 -1283 -3978
rect -1354 -4026 -1283 -4024
rect -1109 -3978 -1038 -3851
rect -732 -3884 -643 -3873
rect -486 -3884 -404 -3872
rect -732 -3885 -404 -3884
rect -732 -3887 -475 -3885
rect -732 -3947 -719 -3887
rect -656 -3947 -475 -3887
rect -413 -3947 -404 -3885
rect -732 -3948 -404 -3947
rect -732 -3960 -643 -3948
rect -486 -3960 -404 -3948
rect -280 -3884 -250 -3837
rect -196 -3884 -170 -3837
rect -280 -3932 -170 -3884
rect -1109 -4024 -1097 -3978
rect -1051 -4024 -1038 -3978
rect -1109 -4026 -1038 -4024
rect -940 -3978 -809 -3977
rect -940 -4024 -929 -3978
rect -883 -4024 -809 -3978
rect -940 -4026 -809 -4024
rect -1698 -4046 -1513 -4026
rect -2084 -4211 -2070 -4179
rect -2167 -4214 -2070 -4211
rect -1886 -4180 -1685 -4133
rect -2071 -4281 -1990 -4276
rect -1886 -4281 -1822 -4180
rect -1732 -4236 -1685 -4180
rect -1732 -4250 -1642 -4236
rect -1732 -4264 -1718 -4250
rect -2071 -4327 -2049 -4281
rect -2003 -4327 -1990 -4281
rect -1892 -4327 -1881 -4281
rect -1835 -4327 -1822 -4281
rect -1731 -4310 -1718 -4264
rect -1655 -4310 -1642 -4250
rect -1731 -4323 -1642 -4310
rect -1584 -4283 -1513 -4046
rect -1441 -4091 -1352 -4078
rect -1441 -4151 -1428 -4091
rect -1365 -4151 -1352 -4091
rect -1441 -4165 -1352 -4151
rect -878 -4090 -809 -4026
rect -280 -3979 -252 -3932
rect -198 -3979 -170 -3932
rect -280 -4042 -170 -3979
rect -647 -4090 -547 -4078
rect -878 -4091 -547 -4090
rect -878 -4095 -630 -4091
rect -878 -4154 -869 -4095
rect -817 -4154 -630 -4095
rect -878 -4158 -630 -4154
rect -563 -4158 -547 -4091
rect -878 -4159 -547 -4158
rect -878 -4283 -809 -4159
rect -647 -4171 -547 -4159
rect -280 -4089 -251 -4042
rect -197 -4089 -170 -4042
rect 308 -3864 400 -3827
rect 544 -3837 556 -3783
rect 610 -3837 616 -3783
rect 544 -3850 616 -3837
rect 761 -3812 762 -3718
rect 808 -3812 809 -3718
rect 761 -3823 809 -3812
rect 308 -4031 355 -3864
rect 433 -3913 523 -3904
rect 433 -3960 442 -3913
rect 514 -3960 523 -3913
rect 433 -3969 523 -3960
rect 308 -4078 400 -4031
rect -280 -4146 -170 -4089
rect 150 -4090 197 -4089
rect -2071 -4438 -1990 -4327
rect -1886 -4328 -1822 -4327
rect -1584 -4329 -1571 -4283
rect -1525 -4329 -1513 -4283
rect -1584 -4330 -1513 -4329
rect -1415 -4329 -1403 -4283
rect -1357 -4329 -1343 -4283
rect -1415 -4438 -1343 -4329
rect -1047 -4329 -1035 -4283
rect -989 -4329 -977 -4283
rect -1047 -4438 -977 -4329
rect -878 -4329 -867 -4283
rect -821 -4329 -809 -4283
rect -878 -4330 -809 -4329
rect -280 -4193 -251 -4146
rect -197 -4193 -170 -4146
rect -280 -4241 -170 -4193
rect -280 -4288 -253 -4241
rect -199 -4288 -170 -4241
rect -730 -4345 -641 -4331
rect -730 -4405 -717 -4345
rect -654 -4405 -641 -4345
rect -730 -4418 -641 -4405
rect -280 -4342 -170 -4288
rect -280 -4389 -250 -4342
rect -196 -4389 -170 -4342
rect -2322 -4462 -2233 -4459
rect -2144 -4462 -784 -4438
rect -2322 -4463 -784 -4462
rect -2322 -4530 -2310 -4463
rect -2243 -4471 -784 -4463
rect -2243 -4473 -1567 -4471
rect -2243 -4522 -2099 -4473
rect -1790 -4517 -1567 -4473
rect -838 -4517 -784 -4471
rect -1790 -4522 -784 -4517
rect -2243 -4529 -784 -4522
rect -2243 -4530 -2233 -4529
rect -2322 -4544 -2233 -4530
rect -2144 -4551 -784 -4529
rect -280 -4446 -170 -4389
rect -280 -4493 -250 -4446
rect -196 -4493 -170 -4446
rect -280 -4541 -170 -4493
rect -56 -4096 -9 -4095
rect -56 -4107 -8 -4096
rect -56 -4201 -54 -4107
rect 133 -4097 215 -4090
rect 133 -4154 146 -4097
rect 203 -4154 215 -4097
rect 133 -4165 150 -4154
rect -56 -4255 -8 -4201
rect 196 -4165 215 -4154
rect 353 -4107 400 -4078
rect 196 -4201 197 -4165
rect 150 -4255 197 -4201
rect -56 -4266 197 -4255
rect -56 -4315 35 -4266
rect 107 -4315 197 -4266
rect -56 -4324 197 -4315
rect -56 -4391 -9 -4324
rect -56 -4402 -8 -4391
rect -56 -4496 -54 -4402
rect -56 -4507 -8 -4496
rect 150 -4402 197 -4324
rect 196 -4496 197 -4402
rect 150 -4503 197 -4496
rect 353 -4201 354 -4107
rect 353 -4402 400 -4201
rect 353 -4496 354 -4402
rect 150 -4507 196 -4503
rect -280 -4588 -252 -4541
rect -198 -4588 -170 -4541
rect -2476 -4601 -2361 -4591
rect -2476 -4602 -2359 -4601
rect -2144 -4602 -784 -4597
rect -2476 -4684 -2450 -4602
rect -2398 -4636 -784 -4602
rect -2398 -4641 -1551 -4636
rect -2398 -4684 -2084 -4641
rect -2476 -4685 -2359 -4684
rect -2476 -4698 -2361 -4685
rect -2144 -4692 -2084 -4684
rect -1834 -4682 -1551 -4641
rect -839 -4682 -784 -4636
rect -1834 -4692 -784 -4682
rect -2144 -4710 -784 -4692
rect -280 -4651 -170 -4588
rect -280 -4698 -251 -4651
rect -197 -4698 -170 -4651
rect -2068 -4802 -1998 -4710
rect -2068 -4876 -2045 -4802
rect -1999 -4876 -1998 -4802
rect -2068 -4891 -1998 -4876
rect -1886 -4802 -1822 -4789
rect -1886 -4876 -1885 -4802
rect -1839 -4876 -1822 -4802
rect -1704 -4796 -1617 -4778
rect -1704 -4861 -1691 -4796
rect -1626 -4834 -1617 -4796
rect -1626 -4837 -1452 -4834
rect -1626 -4861 -1509 -4837
rect -1704 -4863 -1509 -4861
rect -2144 -4965 -1940 -4957
rect -2144 -4967 -2015 -4965
rect -2331 -5012 -2015 -4967
rect -2331 -5039 -2142 -5012
rect -2167 -5070 -2142 -5039
rect -2084 -5024 -2015 -5012
rect -1952 -5024 -1940 -4965
rect -2084 -5038 -1940 -5024
rect -1886 -4992 -1822 -4876
rect -1698 -4883 -1509 -4863
rect -1463 -4883 -1452 -4837
rect -1698 -4885 -1452 -4883
rect -1354 -4837 -1283 -4710
rect -1354 -4883 -1341 -4837
rect -1295 -4883 -1283 -4837
rect -1354 -4885 -1283 -4883
rect -1109 -4837 -1038 -4710
rect -732 -4745 -643 -4732
rect -522 -4745 -447 -4733
rect -732 -4746 -447 -4745
rect -732 -4806 -719 -4746
rect -656 -4805 -517 -4746
rect -458 -4805 -447 -4746
rect -656 -4806 -447 -4805
rect -732 -4819 -643 -4806
rect -522 -4820 -447 -4806
rect -280 -4755 -170 -4698
rect 165 -4615 250 -4599
rect 165 -4618 179 -4615
rect 165 -4683 176 -4618
rect 165 -4687 179 -4683
rect 241 -4687 250 -4615
rect 165 -4699 250 -4687
rect -280 -4802 -251 -4755
rect -197 -4802 -170 -4755
rect -1109 -4883 -1097 -4837
rect -1051 -4883 -1038 -4837
rect -1109 -4885 -1038 -4883
rect -940 -4837 -809 -4836
rect -940 -4883 -929 -4837
rect -883 -4883 -809 -4837
rect -940 -4885 -809 -4883
rect -1698 -4905 -1513 -4885
rect -2084 -5070 -2070 -5038
rect -2167 -5073 -2070 -5070
rect -1886 -5039 -1685 -4992
rect -2071 -5140 -1990 -5135
rect -1886 -5140 -1822 -5039
rect -1732 -5095 -1685 -5039
rect -1732 -5109 -1642 -5095
rect -1732 -5123 -1718 -5109
rect -2071 -5186 -2049 -5140
rect -2003 -5186 -1990 -5140
rect -1892 -5186 -1881 -5140
rect -1835 -5186 -1822 -5140
rect -1731 -5169 -1718 -5123
rect -1655 -5169 -1642 -5109
rect -1731 -5182 -1642 -5169
rect -1584 -5142 -1513 -4905
rect -1441 -4950 -1352 -4937
rect -1441 -5010 -1428 -4950
rect -1365 -5010 -1352 -4950
rect -1441 -5024 -1352 -5010
rect -878 -4952 -809 -4885
rect -280 -4850 -170 -4802
rect -280 -4897 -253 -4850
rect -199 -4897 -170 -4850
rect -641 -4952 -549 -4940
rect -878 -4953 -549 -4952
rect -878 -4954 -630 -4953
rect -878 -5013 -869 -4954
rect -817 -5013 -630 -4954
rect -570 -5013 -549 -4953
rect -878 -5014 -549 -5013
rect -878 -5142 -809 -5014
rect -641 -5025 -549 -5014
rect -280 -4954 -170 -4897
rect -280 -5001 -249 -4954
rect -195 -5001 -170 -4954
rect -55 -4787 -6 -4775
rect -55 -4881 -54 -4787
rect -8 -4881 -6 -4787
rect -55 -4973 -6 -4881
rect 149 -4787 198 -4776
rect 149 -4881 150 -4787
rect 196 -4881 198 -4787
rect 149 -4973 198 -4881
rect 353 -4787 400 -4496
rect 353 -4881 354 -4787
rect 353 -4896 400 -4881
rect 455 -4971 506 -3969
rect 556 -4096 603 -4022
rect 556 -4107 604 -4096
rect 556 -4201 558 -4107
rect 556 -4253 604 -4201
rect 761 -4107 808 -3823
rect 761 -4201 762 -4107
rect 556 -4265 671 -4253
rect 556 -4321 601 -4265
rect 657 -4321 671 -4265
rect 556 -4333 671 -4321
rect 556 -4391 603 -4333
rect 556 -4402 604 -4391
rect 556 -4496 558 -4402
rect 556 -4507 604 -4496
rect 761 -4402 808 -4201
rect 761 -4496 762 -4402
rect 761 -4506 808 -4496
rect 724 -4553 808 -4506
rect 724 -4715 771 -4553
rect 863 -4606 911 -3599
rect 1033 -3634 1081 -3484
rect 1160 -3548 1233 -3535
rect 1160 -3606 1166 -3548
rect 1224 -3551 1233 -3548
rect 1224 -3603 1626 -3551
rect 1224 -3606 1233 -3603
rect 1160 -3619 1233 -3606
rect 966 -3682 1081 -3634
rect 966 -3718 1014 -3682
rect 1012 -3812 1014 -3718
rect 966 -3903 1014 -3812
rect 1166 -3718 1218 -3619
rect 1166 -3812 1170 -3718
rect 1216 -3812 1218 -3718
rect 1374 -3718 1420 -3707
rect 1166 -3824 1218 -3812
rect 1365 -3781 1374 -3768
rect 1574 -3718 1626 -3603
rect 1785 -3554 1833 -3484
rect 2724 -3458 2754 -3411
rect 2808 -3458 2839 -3411
rect 2724 -3515 2839 -3458
rect 1985 -3554 2036 -3553
rect 1785 -3559 2036 -3554
rect 2112 -3559 2163 -3558
rect 1785 -3563 2569 -3559
rect 1785 -3610 1871 -3563
rect 1942 -3568 2569 -3563
rect 1942 -3610 2203 -3568
rect 1785 -3615 2203 -3610
rect 2275 -3615 2407 -3568
rect 2479 -3581 2569 -3568
rect 2724 -3562 2754 -3515
rect 2808 -3562 2839 -3515
rect 2479 -3615 2570 -3581
rect 1785 -3619 2570 -3615
rect 1785 -3707 1833 -3619
rect 1420 -3781 1433 -3768
rect 966 -3951 1105 -3903
rect 1049 -3980 1105 -3951
rect 1049 -3993 1119 -3980
rect 1049 -4047 1054 -3993
rect 1108 -4047 1119 -3993
rect 1049 -4059 1119 -4047
rect 965 -4107 1012 -4096
rect 965 -4201 966 -4107
rect 965 -4258 1012 -4201
rect 1170 -4107 1217 -3824
rect 1365 -3838 1368 -3781
rect 1425 -3838 1433 -3781
rect 1574 -3812 1578 -3718
rect 1624 -3812 1626 -3718
rect 1574 -3827 1626 -3812
rect 1782 -3718 1833 -3707
rect 1828 -3812 1833 -3718
rect 1782 -3823 1833 -3812
rect 1985 -3626 2570 -3619
rect 1985 -3718 2036 -3626
rect 1985 -3812 1986 -3718
rect 2032 -3812 2036 -3718
rect 1985 -3823 2036 -3812
rect 2112 -3718 2163 -3626
rect 2112 -3812 2114 -3718
rect 2160 -3812 2163 -3718
rect 2112 -3823 2163 -3812
rect 2316 -3718 2367 -3626
rect 2316 -3812 2318 -3718
rect 2364 -3812 2367 -3718
rect 1785 -3827 1833 -3823
rect 2316 -3825 2367 -3812
rect 2519 -3718 2570 -3626
rect 2519 -3812 2522 -3718
rect 2568 -3812 2570 -3718
rect 2519 -3820 2570 -3812
rect 2724 -3610 2839 -3562
rect 2724 -3657 2752 -3610
rect 2806 -3657 2839 -3610
rect 2724 -3719 2839 -3657
rect 2724 -3766 2753 -3719
rect 2807 -3766 2839 -3719
rect 3231 -2537 3339 -2475
rect 3231 -2586 3255 -2537
rect 3318 -2586 3339 -2537
rect 3231 -2648 3339 -2586
rect 3231 -2697 3255 -2648
rect 3318 -2697 3339 -2648
rect 3231 -2759 3339 -2697
rect 3512 -2303 3561 -2293
rect 3512 -2397 3514 -2303
rect 3560 -2397 3561 -2303
rect 3512 -2460 3561 -2397
rect 3717 -2303 3766 -2292
rect 3717 -2397 3718 -2303
rect 3764 -2397 3766 -2303
rect 3717 -2460 3766 -2397
rect 3919 -2303 3968 -2289
rect 3919 -2397 3922 -2303
rect 3919 -2456 3968 -2397
rect 4042 -2292 4094 -2178
rect 4231 -2185 4244 -2115
rect 4314 -2185 4325 -2115
rect 4456 -2132 4505 -2032
rect 4456 -2181 4631 -2132
rect 5117 -2142 5166 -2031
rect 5653 -2131 5704 -2015
rect 5860 -1919 5910 -1884
rect 5860 -2013 5862 -1919
rect 5908 -2013 5910 -1919
rect 5860 -2027 5910 -2013
rect 6061 -1908 6111 -1878
rect 6350 -1840 6374 -1791
rect 6437 -1840 6458 -1791
rect 6350 -1902 6458 -1840
rect 6061 -1919 6112 -1908
rect 6061 -2013 6066 -1919
rect 6061 -2024 6112 -2013
rect 6350 -1951 6374 -1902
rect 6437 -1951 6458 -1902
rect 6350 -2013 6458 -1951
rect 6061 -2030 6111 -2024
rect 4231 -2194 4325 -2185
rect 4042 -2303 4096 -2292
rect 4042 -2397 4050 -2303
rect 4042 -2402 4096 -2397
rect 3512 -2469 3766 -2460
rect 3512 -2518 3603 -2469
rect 3675 -2472 3766 -2469
rect 3862 -2469 3968 -2456
rect 3862 -2472 3875 -2469
rect 3675 -2518 3875 -2472
rect 3512 -2521 3875 -2518
rect 3512 -2527 3766 -2521
rect 3512 -2593 3561 -2527
rect 3512 -2687 3514 -2593
rect 3560 -2687 3561 -2593
rect 3512 -2702 3561 -2687
rect 3717 -2593 3766 -2527
rect 3862 -2523 3875 -2521
rect 3929 -2472 3968 -2469
rect 4047 -2466 4096 -2402
rect 4253 -2303 4302 -2290
rect 4253 -2397 4254 -2303
rect 4300 -2397 4302 -2303
rect 4253 -2466 4302 -2397
rect 4456 -2303 4505 -2287
rect 4456 -2397 4458 -2303
rect 4504 -2397 4505 -2303
rect 4456 -2451 4505 -2397
rect 4419 -2463 4505 -2451
rect 4419 -2466 4431 -2463
rect 3929 -2521 3970 -2472
rect 4047 -2515 4431 -2466
rect 3929 -2523 3968 -2521
rect 3862 -2536 3968 -2523
rect 3717 -2687 3718 -2593
rect 3764 -2687 3766 -2593
rect 3717 -2701 3766 -2687
rect 3919 -2593 3968 -2536
rect 4047 -2583 4096 -2515
rect 3919 -2687 3922 -2593
rect 3919 -2698 3968 -2687
rect 4045 -2593 4096 -2583
rect 4045 -2687 4050 -2593
rect 3231 -2808 3255 -2759
rect 3318 -2808 3339 -2759
rect 4045 -2703 4096 -2687
rect 4253 -2593 4302 -2515
rect 4419 -2517 4431 -2515
rect 4485 -2466 4505 -2463
rect 4582 -2292 4631 -2181
rect 4990 -2191 5166 -2142
rect 5526 -2182 5704 -2131
rect 6350 -2062 6374 -2013
rect 6437 -2062 6458 -2013
rect 6350 -2124 6458 -2062
rect 6350 -2173 6374 -2124
rect 6437 -2173 6458 -2124
rect 4582 -2303 4632 -2292
rect 4582 -2397 4586 -2303
rect 4582 -2408 4632 -2397
rect 4789 -2303 4838 -2286
rect 4789 -2397 4790 -2303
rect 4836 -2397 4838 -2303
rect 4485 -2515 4507 -2466
rect 4582 -2478 4631 -2408
rect 4789 -2478 4838 -2397
rect 4990 -2292 5039 -2191
rect 4990 -2303 5040 -2292
rect 4990 -2397 4994 -2303
rect 4990 -2408 5040 -2397
rect 5120 -2303 5170 -2289
rect 5120 -2397 5122 -2303
rect 5168 -2397 5170 -2303
rect 4990 -2478 5039 -2408
rect 5120 -2450 5170 -2397
rect 5324 -2303 5373 -2291
rect 5324 -2397 5326 -2303
rect 5372 -2397 5373 -2303
rect 5116 -2462 5187 -2450
rect 4485 -2517 4505 -2515
rect 4419 -2529 4505 -2517
rect 4253 -2687 4254 -2593
rect 4300 -2687 4302 -2593
rect 4253 -2699 4302 -2687
rect 4456 -2593 4505 -2529
rect 4456 -2687 4458 -2593
rect 4504 -2687 4505 -2593
rect 4456 -2696 4505 -2687
rect 4582 -2527 5040 -2478
rect 5116 -2518 5122 -2462
rect 5178 -2475 5187 -2462
rect 5324 -2475 5373 -2397
rect 5526 -2303 5577 -2182
rect 6350 -2235 6458 -2173
rect 6350 -2284 6374 -2235
rect 6437 -2284 6458 -2235
rect 5526 -2397 5530 -2303
rect 5576 -2397 5577 -2303
rect 5526 -2429 5577 -2397
rect 5655 -2303 5704 -2287
rect 5655 -2397 5658 -2303
rect 5526 -2475 5575 -2429
rect 5178 -2518 5575 -2475
rect 5116 -2524 5575 -2518
rect 5116 -2527 5187 -2524
rect 4582 -2582 4631 -2527
rect 4582 -2593 4632 -2582
rect 4582 -2687 4586 -2593
rect 4458 -2698 4504 -2696
rect 4582 -2698 4632 -2687
rect 4789 -2593 4838 -2527
rect 4789 -2687 4790 -2593
rect 4836 -2687 4838 -2593
rect 4789 -2695 4838 -2687
rect 4990 -2582 5039 -2527
rect 4990 -2593 5040 -2582
rect 4990 -2687 4994 -2593
rect 4790 -2698 4836 -2695
rect 4990 -2698 5040 -2687
rect 5120 -2593 5169 -2527
rect 5120 -2687 5122 -2593
rect 5168 -2687 5169 -2593
rect 5120 -2697 5169 -2687
rect 5324 -2593 5373 -2524
rect 5324 -2687 5326 -2593
rect 5372 -2687 5373 -2593
rect 5122 -2698 5168 -2697
rect 3231 -2870 3339 -2808
rect 3231 -2919 3255 -2870
rect 3318 -2919 3339 -2870
rect 3746 -2801 3846 -2789
rect 3746 -2809 3768 -2801
rect 3746 -2860 3755 -2809
rect 3746 -2868 3768 -2860
rect 3834 -2868 3846 -2801
rect 4045 -2807 4095 -2703
rect 4582 -2797 4631 -2698
rect 3746 -2880 3846 -2868
rect 3918 -2857 4095 -2807
rect 4459 -2846 4631 -2797
rect 4990 -2816 5039 -2698
rect 5324 -2700 5373 -2687
rect 5526 -2582 5575 -2524
rect 5655 -2450 5704 -2397
rect 5859 -2303 5908 -2288
rect 5859 -2397 5862 -2303
rect 5859 -2440 5908 -2397
rect 6064 -2303 6113 -2289
rect 6064 -2397 6066 -2303
rect 6112 -2397 6113 -2303
rect 6064 -2440 6113 -2397
rect 5859 -2449 6113 -2440
rect 5655 -2463 5731 -2450
rect 5655 -2517 5666 -2463
rect 5720 -2466 5731 -2463
rect 5859 -2466 5951 -2449
rect 5720 -2499 5951 -2466
rect 6023 -2499 6113 -2449
rect 5720 -2515 6113 -2499
rect 5720 -2517 5731 -2515
rect 5655 -2529 5731 -2517
rect 5526 -2593 5581 -2582
rect 5526 -2687 5530 -2593
rect 5576 -2687 5581 -2593
rect 5526 -2697 5581 -2687
rect 5655 -2593 5704 -2529
rect 5655 -2687 5658 -2593
rect 5655 -2696 5704 -2687
rect 5530 -2698 5581 -2697
rect 5658 -2698 5704 -2696
rect 5859 -2593 5908 -2515
rect 5859 -2687 5862 -2593
rect 5859 -2697 5908 -2687
rect 5862 -2698 5908 -2697
rect 6064 -2593 6113 -2515
rect 6064 -2687 6066 -2593
rect 6112 -2687 6113 -2593
rect 6064 -2698 6113 -2687
rect 6350 -2346 6458 -2284
rect 6350 -2395 6374 -2346
rect 6437 -2395 6458 -2346
rect 6350 -2457 6458 -2395
rect 6350 -2506 6374 -2457
rect 6437 -2506 6458 -2457
rect 6350 -2568 6458 -2506
rect 6350 -2617 6374 -2568
rect 6437 -2617 6458 -2568
rect 6350 -2679 6458 -2617
rect 5531 -2804 5581 -2698
rect 6350 -2728 6374 -2679
rect 6437 -2728 6458 -2679
rect 6350 -2790 6458 -2728
rect 3231 -2981 3339 -2919
rect 3231 -3030 3255 -2981
rect 3318 -3030 3339 -2981
rect 3231 -3092 3339 -3030
rect 3231 -3141 3255 -3092
rect 3318 -3141 3339 -3092
rect 3514 -2977 3564 -2965
rect 3560 -3071 3564 -2977
rect 3514 -3108 3564 -3071
rect 3716 -2977 3766 -2965
rect 3716 -3071 3718 -2977
rect 3764 -3071 3766 -2977
rect 3716 -3089 3766 -3071
rect 3918 -2977 3968 -2857
rect 3918 -3071 3922 -2977
rect 3918 -3089 3968 -3071
rect 4048 -2909 4098 -2908
rect 4459 -2909 4508 -2846
rect 4990 -2865 5174 -2816
rect 5531 -2854 5707 -2804
rect 4048 -2958 4508 -2909
rect 4048 -2977 4098 -2958
rect 4048 -3071 4050 -2977
rect 4096 -3071 4098 -2977
rect 4048 -3082 4098 -3071
rect 4251 -2977 4301 -2958
rect 4251 -3071 4254 -2977
rect 4300 -3071 4301 -2977
rect 4045 -3089 4101 -3082
rect 4251 -3088 4301 -3071
rect 4457 -2977 4508 -2958
rect 4457 -3071 4458 -2977
rect 4504 -3071 4508 -2977
rect 4457 -3072 4508 -3071
rect 4586 -2977 4636 -2960
rect 4632 -3071 4636 -2977
rect 4457 -3088 4507 -3072
rect 4586 -3089 4636 -3071
rect 4786 -2977 4836 -2965
rect 4786 -3071 4790 -2977
rect 4786 -3089 4836 -3071
rect 4992 -2977 5047 -2959
rect 5125 -2965 5174 -2865
rect 4992 -3071 4994 -2977
rect 5040 -3071 5047 -2977
rect 4992 -3089 5047 -3071
rect 3716 -3108 3968 -3089
rect 3231 -3203 3339 -3141
rect 3511 -3118 3968 -3108
rect 3511 -3166 3603 -3118
rect 3675 -3139 3968 -3118
rect 4031 -3091 4117 -3089
rect 3675 -3166 3767 -3139
rect 4031 -3145 4046 -3091
rect 4100 -3145 4117 -3091
rect 4586 -3139 5047 -3089
rect 4031 -3160 4117 -3145
rect 3511 -3175 3767 -3166
rect 3231 -3252 3255 -3203
rect 3318 -3252 3339 -3203
rect 3231 -3314 3339 -3252
rect 4232 -3184 4326 -3180
rect 4232 -3257 4245 -3184
rect 4313 -3257 4326 -3184
rect 4997 -3205 5047 -3139
rect 5117 -2977 5174 -2965
rect 5117 -3071 5122 -2977
rect 5168 -3071 5174 -2977
rect 5117 -3091 5174 -3071
rect 5326 -2977 5376 -2959
rect 5372 -3071 5376 -2977
rect 5326 -3091 5376 -3071
rect 5528 -2977 5578 -2963
rect 5528 -3071 5530 -2977
rect 5576 -3071 5578 -2977
rect 5528 -3091 5578 -3071
rect 5117 -3141 5578 -3091
rect 5657 -2977 5707 -2854
rect 6350 -2839 6374 -2790
rect 6437 -2839 6458 -2790
rect 6350 -2901 6458 -2839
rect 6350 -2950 6374 -2901
rect 6437 -2950 6458 -2901
rect 5657 -3071 5658 -2977
rect 5704 -3071 5707 -2977
rect 5657 -3088 5707 -3071
rect 5856 -2966 5906 -2962
rect 5856 -2977 5908 -2966
rect 5856 -3071 5862 -2977
rect 5856 -3082 5908 -3071
rect 6063 -2977 6113 -2960
rect 6063 -3071 6066 -2977
rect 6112 -3071 6113 -2977
rect 5856 -3088 5906 -3082
rect 5657 -3097 5906 -3088
rect 5657 -3151 5762 -3097
rect 5816 -3132 5906 -3097
rect 6063 -3132 6113 -3071
rect 5816 -3141 6113 -3132
rect 5816 -3151 5951 -3141
rect 5657 -3165 5951 -3151
rect 5657 -3205 5707 -3165
rect 5861 -3187 5951 -3165
rect 6023 -3187 6113 -3141
rect 5861 -3195 6113 -3187
rect 5942 -3196 6113 -3195
rect 6350 -3012 6458 -2950
rect 6350 -3061 6374 -3012
rect 6437 -3061 6458 -3012
rect 6350 -3123 6458 -3061
rect 6350 -3172 6374 -3123
rect 6437 -3172 6458 -3123
rect 4997 -3255 5707 -3205
rect 6350 -3234 6458 -3172
rect 4232 -3269 4326 -3257
rect 3231 -3363 3255 -3314
rect 3318 -3363 3339 -3314
rect 6350 -3283 6374 -3234
rect 6437 -3283 6458 -3234
rect 6350 -3345 6458 -3283
rect 3231 -3425 3339 -3363
rect 4029 -3368 4115 -3358
rect 4029 -3388 4045 -3368
rect 3231 -3474 3255 -3425
rect 3318 -3474 3339 -3425
rect 3567 -3422 3655 -3413
rect 3567 -3438 3576 -3422
rect 3231 -3536 3339 -3474
rect 3559 -3440 3576 -3438
rect 3646 -3438 3655 -3422
rect 3715 -3424 4045 -3388
rect 4101 -3388 4115 -3368
rect 5064 -3385 5147 -3376
rect 5064 -3388 5078 -3385
rect 4101 -3424 5078 -3388
rect 3646 -3440 3665 -3438
rect 3559 -3500 3568 -3440
rect 3654 -3500 3665 -3440
rect 3559 -3511 3665 -3500
rect 3715 -3439 5078 -3424
rect 3231 -3585 3255 -3536
rect 3318 -3585 3339 -3536
rect 3231 -3647 3339 -3585
rect 3231 -3696 3255 -3647
rect 3318 -3696 3339 -3647
rect 3231 -3758 3339 -3696
rect 3512 -3611 3562 -3591
rect 3512 -3705 3514 -3611
rect 3560 -3705 3562 -3611
rect 3512 -3708 3562 -3705
rect 3715 -3611 3766 -3439
rect 4314 -3498 4392 -3486
rect 3715 -3705 3718 -3611
rect 3764 -3705 3766 -3611
rect 3715 -3708 3766 -3705
rect 3512 -3753 3766 -3708
rect 3919 -3499 4392 -3498
rect 3919 -3549 4326 -3499
rect 3919 -3611 3970 -3549
rect 4314 -3553 4326 -3549
rect 4380 -3553 4392 -3499
rect 4314 -3563 4392 -3553
rect 3919 -3705 3922 -3611
rect 3968 -3705 3970 -3611
rect 3919 -3720 3970 -3705
rect 4123 -3611 4174 -3595
rect 4123 -3705 4126 -3611
rect 4172 -3705 4174 -3611
rect 3231 -3766 3255 -3758
rect 2724 -3807 3255 -3766
rect 3318 -3807 3339 -3758
rect 2522 -3823 2568 -3820
rect 2724 -3823 3339 -3807
rect 3510 -3759 3766 -3753
rect 3510 -3762 3599 -3759
rect 3510 -3809 3519 -3762
rect 3590 -3809 3599 -3762
rect 4123 -3805 4174 -3705
rect 4327 -3611 4379 -3563
rect 4327 -3705 4330 -3611
rect 4376 -3705 4379 -3611
rect 4327 -3718 4379 -3705
rect 4530 -3611 4581 -3439
rect 5064 -3441 5078 -3439
rect 5134 -3388 5147 -3385
rect 5134 -3439 5400 -3388
rect 5134 -3441 5147 -3439
rect 5064 -3443 5147 -3441
rect 5349 -3482 5400 -3439
rect 6350 -3394 6374 -3345
rect 6437 -3394 6458 -3345
rect 6350 -3456 6458 -3394
rect 5349 -3483 5725 -3482
rect 5349 -3484 5730 -3483
rect 4730 -3494 4804 -3486
rect 5349 -3491 6138 -3484
rect 4730 -3498 5194 -3494
rect 4730 -3554 4738 -3498
rect 4794 -3545 5194 -3498
rect 4794 -3554 4804 -3545
rect 4730 -3567 4804 -3554
rect 4530 -3705 4534 -3611
rect 4580 -3705 4581 -3611
rect 4530 -3711 4581 -3705
rect 4733 -3611 4785 -3567
rect 4938 -3597 4989 -3593
rect 4733 -3705 4738 -3611
rect 4784 -3705 4785 -3611
rect 4534 -3716 4580 -3711
rect 4733 -3718 4785 -3705
rect 4937 -3611 4989 -3597
rect 4937 -3705 4942 -3611
rect 4988 -3705 4989 -3611
rect 4937 -3716 4989 -3705
rect 5143 -3611 5194 -3545
rect 5143 -3705 5146 -3611
rect 5192 -3705 5194 -3611
rect 5143 -3713 5194 -3705
rect 5349 -3541 5439 -3491
rect 5511 -3493 6138 -3491
rect 5511 -3540 5771 -3493
rect 5843 -3540 6138 -3493
rect 5511 -3541 6138 -3540
rect 5349 -3549 6138 -3541
rect 5349 -3550 5730 -3549
rect 5349 -3611 5400 -3550
rect 5349 -3705 5350 -3611
rect 5396 -3705 5400 -3611
rect 5146 -3716 5192 -3713
rect 5349 -3716 5400 -3705
rect 5549 -3611 5600 -3550
rect 5549 -3705 5554 -3611
rect 5549 -3714 5600 -3705
rect 5679 -3611 5730 -3550
rect 5679 -3705 5682 -3611
rect 5728 -3705 5730 -3611
rect 5679 -3714 5730 -3705
rect 5884 -3611 5935 -3549
rect 5884 -3705 5886 -3611
rect 5932 -3705 5935 -3611
rect 5554 -3716 5600 -3714
rect 5682 -3716 5728 -3714
rect 5884 -3716 5935 -3705
rect 6087 -3611 6138 -3549
rect 6087 -3705 6090 -3611
rect 6136 -3705 6138 -3611
rect 6087 -3715 6138 -3705
rect 6350 -3505 6374 -3456
rect 6437 -3505 6458 -3456
rect 6350 -3567 6458 -3505
rect 6350 -3616 6374 -3567
rect 6437 -3616 6458 -3567
rect 6350 -3678 6458 -3616
rect 6090 -3716 6136 -3715
rect 3510 -3818 3599 -3809
rect 4110 -3814 4187 -3805
rect 4110 -3817 4122 -3814
rect 1365 -3850 1433 -3838
rect 1365 -3997 1432 -3984
rect 1365 -4053 1367 -3997
rect 1423 -4053 1432 -3997
rect 1365 -4067 1432 -4053
rect 1216 -4201 1217 -4107
rect 965 -4272 1049 -4258
rect 965 -4329 988 -4272
rect 1045 -4329 1049 -4272
rect 965 -4345 1049 -4329
rect 965 -4402 1012 -4345
rect 965 -4496 966 -4402
rect 965 -4508 1012 -4496
rect 1170 -4402 1217 -4201
rect 1216 -4496 1217 -4402
rect 842 -4615 932 -4606
rect 842 -4663 851 -4615
rect 923 -4663 932 -4615
rect 842 -4672 932 -4663
rect 724 -4762 809 -4715
rect -2071 -5297 -1990 -5186
rect -1886 -5187 -1822 -5186
rect -1584 -5188 -1571 -5142
rect -1525 -5188 -1513 -5142
rect -1584 -5189 -1513 -5188
rect -1415 -5188 -1403 -5142
rect -1357 -5188 -1343 -5142
rect -1415 -5297 -1343 -5188
rect -1047 -5188 -1035 -5142
rect -989 -5188 -977 -5142
rect -1047 -5297 -977 -5188
rect -878 -5188 -867 -5142
rect -821 -5188 -809 -5142
rect -878 -5189 -809 -5188
rect -280 -5064 -170 -5001
rect -56 -4983 200 -4973
rect -56 -5029 35 -4983
rect 107 -5029 200 -4983
rect -56 -5038 200 -5029
rect 372 -4980 506 -4971
rect 372 -5029 387 -4980
rect 459 -5029 506 -4980
rect 557 -4787 606 -4776
rect 557 -4881 558 -4787
rect 604 -4881 606 -4787
rect 557 -4934 606 -4881
rect 761 -4787 808 -4762
rect 761 -4881 762 -4787
rect 950 -4779 1030 -4774
rect 950 -4835 962 -4779
rect 1018 -4835 1030 -4779
rect 950 -4845 966 -4835
rect 761 -4898 808 -4881
rect 962 -4881 966 -4845
rect 1012 -4845 1030 -4835
rect 1170 -4787 1217 -4496
rect 1371 -4107 1420 -4067
rect 1371 -4201 1374 -4107
rect 1371 -4212 1420 -4201
rect 1577 -4107 1624 -3827
rect 2724 -3870 2753 -3823
rect 2807 -3870 2839 -3823
rect 2724 -3918 2839 -3870
rect 2724 -3965 2751 -3918
rect 2805 -3965 2839 -3918
rect 2724 -4028 2839 -3965
rect 2724 -4075 2752 -4028
rect 2806 -4075 2839 -4028
rect 1577 -4201 1578 -4107
rect 1780 -4096 1827 -4095
rect 1780 -4107 1828 -4096
rect 1780 -4112 1782 -4107
rect 1760 -4119 1782 -4112
rect 1986 -4107 2033 -4095
rect 1828 -4119 1842 -4112
rect 1760 -4176 1773 -4119
rect 1830 -4176 1842 -4119
rect 1760 -4183 1782 -4176
rect 1371 -4391 1419 -4212
rect 1371 -4402 1420 -4391
rect 1371 -4496 1374 -4402
rect 1371 -4507 1420 -4496
rect 1577 -4402 1624 -4201
rect 1780 -4201 1782 -4183
rect 1828 -4183 1842 -4176
rect 1780 -4256 1828 -4201
rect 2032 -4201 2033 -4107
rect 1986 -4256 2033 -4201
rect 1779 -4265 2033 -4256
rect 2114 -4097 2160 -4096
rect 2114 -4107 2161 -4097
rect 2160 -4201 2161 -4107
rect 2114 -4265 2161 -4201
rect 2318 -4107 2365 -4095
rect 2364 -4201 2365 -4107
rect 2318 -4262 2365 -4201
rect 2522 -4107 2569 -4091
rect 2568 -4201 2569 -4107
rect 2522 -4262 2569 -4201
rect 2318 -4265 2569 -4262
rect 1779 -4311 1871 -4265
rect 1943 -4271 2569 -4265
rect 1943 -4274 2407 -4271
rect 1943 -4311 2203 -4274
rect 1779 -4319 2203 -4311
rect 1577 -4496 1578 -4402
rect 1371 -4569 1419 -4507
rect 1356 -4581 1427 -4569
rect 1356 -4635 1368 -4581
rect 1422 -4635 1427 -4581
rect 1356 -4647 1427 -4635
rect 1012 -4881 1018 -4845
rect 962 -4893 1018 -4881
rect 1216 -4881 1217 -4787
rect 1170 -4896 1217 -4881
rect 1369 -4776 1418 -4775
rect 1369 -4787 1420 -4776
rect 1369 -4881 1374 -4787
rect 1369 -4892 1420 -4881
rect 1577 -4787 1624 -4496
rect 1780 -4321 2203 -4319
rect 1780 -4391 1827 -4321
rect 1986 -4322 2203 -4321
rect 2275 -4318 2407 -4274
rect 2479 -4318 2569 -4271
rect 2275 -4322 2569 -4318
rect 1986 -4330 2569 -4322
rect 1986 -4331 2365 -4330
rect 1780 -4402 1828 -4391
rect 1780 -4496 1782 -4402
rect 1780 -4507 1828 -4496
rect 1986 -4402 2033 -4331
rect 2032 -4496 2033 -4402
rect 1986 -4507 2033 -4496
rect 2114 -4402 2161 -4331
rect 2160 -4496 2161 -4402
rect 2114 -4509 2161 -4496
rect 2318 -4402 2365 -4331
rect 2364 -4496 2365 -4402
rect 2318 -4507 2365 -4496
rect 2522 -4402 2569 -4330
rect 2568 -4496 2569 -4402
rect 2522 -4503 2569 -4496
rect 2724 -4132 2839 -4075
rect 2724 -4179 2752 -4132
rect 2806 -4179 2839 -4132
rect 2724 -4227 2839 -4179
rect 2724 -4274 2750 -4227
rect 2804 -4274 2839 -4227
rect 2724 -4328 2839 -4274
rect 2724 -4375 2753 -4328
rect 2807 -4375 2839 -4328
rect 2724 -4432 2839 -4375
rect 2724 -4479 2753 -4432
rect 2807 -4479 2839 -4432
rect 2522 -4507 2568 -4503
rect 2724 -4527 2839 -4479
rect 2724 -4574 2751 -4527
rect 2805 -4574 2839 -4527
rect 2724 -4637 2839 -4574
rect 2724 -4684 2752 -4637
rect 2806 -4684 2839 -4637
rect 2724 -4741 2839 -4684
rect 1577 -4881 1578 -4787
rect 1782 -4777 1828 -4776
rect 1782 -4787 1831 -4777
rect 1764 -4795 1782 -4792
rect 1828 -4792 1831 -4787
rect 1983 -4787 2034 -4757
rect 1828 -4795 1846 -4792
rect 1764 -4851 1777 -4795
rect 1833 -4851 1846 -4795
rect 1764 -4860 1782 -4851
rect 557 -4946 716 -4934
rect 557 -5003 652 -4946
rect 709 -4955 716 -4946
rect 1369 -4955 1418 -4892
rect 1577 -4898 1624 -4881
rect 1828 -4860 1846 -4851
rect 1828 -4881 1831 -4860
rect 709 -5003 1418 -4955
rect 1782 -4943 1831 -4881
rect 1983 -4881 1986 -4787
rect 2032 -4881 2034 -4787
rect 1983 -4943 2034 -4881
rect 2111 -4787 2162 -4758
rect 2111 -4881 2114 -4787
rect 2160 -4881 2162 -4787
rect 2111 -4943 2162 -4881
rect 2317 -4787 2368 -4758
rect 2317 -4881 2318 -4787
rect 2364 -4881 2368 -4787
rect 2317 -4943 2368 -4881
rect 2521 -4787 2572 -4757
rect 2521 -4881 2522 -4787
rect 2568 -4881 2572 -4787
rect 2521 -4943 2572 -4881
rect 1782 -4953 2572 -4943
rect 557 -5004 1418 -5003
rect 1478 -4977 1544 -4971
rect 1478 -4980 1638 -4977
rect 647 -5013 716 -5004
rect 372 -5032 506 -5029
rect 372 -5038 468 -5032
rect -280 -5111 -248 -5064
rect -194 -5111 -170 -5064
rect -280 -5168 -170 -5111
rect 149 -5110 198 -5038
rect 1478 -5052 1487 -4980
rect 1535 -4989 1638 -4980
rect 1535 -5043 1572 -4989
rect 1626 -5043 1638 -4989
rect 1535 -5052 1638 -5043
rect 1782 -4999 1871 -4953
rect 1943 -4999 2203 -4953
rect 2275 -4999 2407 -4953
rect 1782 -5003 2407 -4999
rect 2479 -5003 2572 -4953
rect 1782 -5008 2572 -5003
rect 2724 -4788 2752 -4741
rect 2806 -4788 2839 -4741
rect 2724 -4836 2839 -4788
rect 2724 -4883 2750 -4836
rect 2804 -4883 2839 -4836
rect 2724 -4940 2839 -4883
rect 2724 -4987 2754 -4940
rect 2808 -4987 2839 -4940
rect 1478 -5061 1544 -5052
rect 1782 -5110 1831 -5008
rect 2398 -5012 2488 -5008
rect 149 -5159 1831 -5110
rect 2724 -5050 2839 -4987
rect 2724 -5097 2755 -5050
rect 2809 -5097 2839 -5050
rect 2724 -5154 2839 -5097
rect -730 -5204 -641 -5190
rect -730 -5264 -717 -5204
rect -654 -5264 -641 -5204
rect -730 -5277 -641 -5264
rect -280 -5215 -248 -5168
rect -194 -5215 -170 -5168
rect -280 -5259 -170 -5215
rect 2724 -5201 2755 -5154
rect 2809 -5201 2839 -5154
rect 2724 -5259 2839 -5201
rect -280 -5285 2839 -5259
rect -280 -5286 499 -5285
rect -2326 -5312 -2231 -5307
rect -2144 -5312 -784 -5297
rect -2326 -5313 -784 -5312
rect -2326 -5380 -2310 -5313
rect -2243 -5330 -784 -5313
rect -2243 -5332 -1567 -5330
rect -2243 -5379 -2099 -5332
rect -2243 -5380 -2231 -5379
rect -2326 -5391 -2231 -5380
rect -2144 -5381 -2099 -5379
rect -1790 -5376 -1567 -5332
rect -838 -5376 -784 -5330
rect -1790 -5381 -784 -5376
rect -2144 -5410 -784 -5381
rect -558 -5402 -477 -5322
rect -280 -5335 -239 -5286
rect -176 -5287 18 -5286
rect -176 -5335 -111 -5287
rect -280 -5336 -111 -5335
rect -48 -5335 18 -5287
rect 81 -5287 370 -5286
rect 81 -5335 135 -5287
rect -48 -5336 135 -5335
rect 198 -5288 370 -5287
rect 198 -5336 247 -5288
rect -280 -5337 247 -5336
rect 310 -5335 370 -5288
rect 433 -5334 499 -5286
rect 562 -5286 1101 -5285
rect 562 -5334 616 -5286
rect 433 -5335 616 -5334
rect 679 -5287 972 -5286
rect 679 -5335 728 -5287
rect 310 -5336 728 -5335
rect 791 -5336 846 -5287
rect 909 -5335 972 -5287
rect 1035 -5334 1101 -5286
rect 1164 -5286 2839 -5285
rect 1164 -5334 1218 -5286
rect 1035 -5335 1218 -5334
rect 1281 -5287 2839 -5286
rect 1281 -5335 1330 -5287
rect 909 -5336 1330 -5335
rect 1393 -5336 1448 -5287
rect 1511 -5336 1571 -5287
rect 1634 -5336 1688 -5287
rect 1751 -5336 1809 -5287
rect 1872 -5336 1931 -5287
rect 1994 -5288 2513 -5287
rect 1994 -5336 2042 -5288
rect 310 -5337 2042 -5336
rect 2105 -5337 2161 -5288
rect 2224 -5337 2273 -5288
rect 2336 -5337 2394 -5288
rect 2457 -5336 2513 -5288
rect 2576 -5289 2739 -5287
rect 2576 -5336 2628 -5289
rect 2457 -5337 2628 -5336
rect -280 -5338 2628 -5337
rect 2691 -5336 2739 -5289
rect 2802 -5336 2839 -5287
rect 2691 -5338 2839 -5336
rect -280 -5371 2839 -5338
rect 3231 -3869 3339 -3823
rect 3715 -3867 4122 -3817
rect 3231 -3918 3255 -3869
rect 3318 -3918 3339 -3869
rect 3231 -3980 3339 -3918
rect 3231 -4029 3255 -3980
rect 3318 -4029 3339 -3980
rect 3514 -3992 3560 -3989
rect 3231 -4091 3339 -4029
rect 3231 -4140 3255 -4091
rect 3318 -4140 3339 -4091
rect 3231 -4202 3339 -4140
rect 3231 -4251 3255 -4202
rect 3318 -4251 3339 -4202
rect 3231 -4313 3339 -4251
rect 3231 -4362 3255 -4313
rect 3318 -4362 3339 -4313
rect 3231 -4424 3339 -4362
rect 3513 -4000 3565 -3992
rect 3513 -4094 3514 -4000
rect 3560 -4094 3565 -4000
rect 3513 -4157 3565 -4094
rect 3716 -4000 3768 -3867
rect 4110 -3868 4122 -3867
rect 4176 -3868 4187 -3814
rect 4110 -3880 4187 -3868
rect 3716 -4094 3718 -4000
rect 3764 -4094 3768 -4000
rect 3716 -4157 3768 -4094
rect 3513 -4166 3768 -4157
rect 3513 -4216 3603 -4166
rect 3675 -4216 3768 -4166
rect 3513 -4225 3768 -4216
rect 3513 -4295 3565 -4225
rect 3513 -4389 3514 -4295
rect 3560 -4389 3565 -4295
rect 3513 -4402 3565 -4389
rect 3716 -4295 3768 -4225
rect 3716 -4389 3718 -4295
rect 3764 -4389 3768 -4295
rect 3231 -4473 3255 -4424
rect 3318 -4473 3339 -4424
rect 3231 -4535 3339 -4473
rect 3231 -4584 3255 -4535
rect 3318 -4584 3339 -4535
rect 3456 -4489 3553 -4476
rect 3456 -4543 3468 -4489
rect 3545 -4543 3553 -4489
rect 3456 -4548 3476 -4543
rect 3467 -4558 3476 -4548
rect 3537 -4548 3553 -4543
rect 3537 -4558 3546 -4548
rect 3467 -4567 3546 -4558
rect 3716 -4553 3768 -4389
rect 3919 -4000 3971 -3988
rect 4126 -3995 4172 -3989
rect 4327 -3990 4378 -3718
rect 3919 -4094 3922 -4000
rect 3968 -4094 3971 -4000
rect 3919 -4295 3971 -4094
rect 4123 -4000 4175 -3995
rect 4123 -4094 4126 -4000
rect 4172 -4094 4175 -4000
rect 4123 -4176 4175 -4094
rect 4325 -4000 4378 -3990
rect 4325 -4094 4330 -4000
rect 4376 -4094 4378 -4000
rect 4517 -3949 4599 -3940
rect 4517 -4003 4530 -3949
rect 4584 -4003 4599 -3949
rect 4517 -4007 4534 -4003
rect 4529 -4012 4534 -4007
rect 4113 -4188 4187 -4176
rect 4113 -4244 4122 -4188
rect 4178 -4244 4187 -4188
rect 4113 -4255 4187 -4244
rect 3919 -4389 3922 -4295
rect 3968 -4389 3971 -4295
rect 3919 -4455 3971 -4389
rect 4123 -4295 4175 -4255
rect 4123 -4389 4126 -4295
rect 4172 -4389 4175 -4295
rect 4123 -4405 4175 -4389
rect 4325 -4295 4378 -4094
rect 4325 -4389 4330 -4295
rect 4376 -4389 4378 -4295
rect 4325 -4455 4378 -4389
rect 4530 -4094 4534 -4012
rect 4580 -4007 4599 -4003
rect 4733 -3981 4784 -3718
rect 4937 -3804 4988 -3716
rect 6350 -3727 6374 -3678
rect 6437 -3727 6458 -3678
rect 6350 -3789 6458 -3727
rect 4928 -3813 5009 -3804
rect 5565 -3806 5653 -3804
rect 4928 -3869 4941 -3813
rect 4997 -3817 5009 -3813
rect 5557 -3813 5662 -3806
rect 5557 -3816 5574 -3813
rect 5644 -3816 5662 -3813
rect 4997 -3867 5396 -3817
rect 4997 -3869 5009 -3867
rect 4928 -3878 5009 -3869
rect 4733 -4000 4785 -3981
rect 4580 -4012 4585 -4007
rect 4580 -4094 4584 -4012
rect 4530 -4295 4584 -4094
rect 4530 -4389 4534 -4295
rect 4580 -4389 4584 -4295
rect 4530 -4399 4584 -4389
rect 4733 -4094 4738 -4000
rect 4784 -4094 4785 -4000
rect 4733 -4295 4785 -4094
rect 4937 -4000 4989 -3983
rect 4937 -4094 4942 -4000
rect 4988 -4094 4989 -4000
rect 4937 -4165 4989 -4094
rect 5140 -4000 5192 -3983
rect 5140 -4094 5146 -4000
rect 4925 -4167 5007 -4165
rect 4925 -4223 4938 -4167
rect 4994 -4223 5007 -4167
rect 4925 -4225 5007 -4223
rect 4733 -4389 4738 -4295
rect 4784 -4389 4785 -4295
rect 4534 -4400 4580 -4399
rect 3919 -4507 4378 -4455
rect 3231 -4646 3339 -4584
rect 3716 -4605 4176 -4553
rect 3231 -4695 3255 -4646
rect 3318 -4695 3339 -4646
rect 3231 -4757 3339 -4695
rect 3231 -4806 3255 -4757
rect 3318 -4806 3339 -4757
rect 3231 -4868 3339 -4806
rect 3512 -4680 3564 -4669
rect 3512 -4774 3514 -4680
rect 3560 -4774 3564 -4680
rect 3512 -4849 3564 -4774
rect 3714 -4680 3766 -4669
rect 3714 -4774 3718 -4680
rect 3764 -4774 3766 -4680
rect 3714 -4849 3766 -4774
rect 3231 -4917 3255 -4868
rect 3318 -4917 3339 -4868
rect 3231 -4979 3339 -4917
rect 3510 -4858 3766 -4849
rect 3510 -4914 3603 -4858
rect 3674 -4914 3766 -4858
rect 3510 -4923 3766 -4914
rect 3231 -5028 3255 -4979
rect 3318 -5028 3339 -4979
rect 3231 -5090 3339 -5028
rect 3231 -5139 3255 -5090
rect 3318 -5139 3339 -5090
rect 3512 -5007 3564 -4923
rect 3512 -5101 3514 -5007
rect 3560 -5101 3564 -5007
rect 3512 -5112 3564 -5101
rect 3714 -5007 3766 -4923
rect 3714 -5101 3718 -5007
rect 3764 -5101 3766 -5007
rect 3231 -5201 3339 -5139
rect 3231 -5250 3255 -5201
rect 3318 -5250 3339 -5201
rect 3231 -5312 3339 -5250
rect 3231 -5361 3255 -5312
rect 3318 -5361 3339 -5312
rect 3714 -5265 3766 -5101
rect 3918 -4680 3970 -4668
rect 3918 -4774 3922 -4680
rect 3968 -4774 3970 -4680
rect 3918 -5007 3970 -4774
rect 4124 -4680 4176 -4605
rect 4325 -4667 4378 -4507
rect 4733 -4449 4785 -4389
rect 4937 -4227 4994 -4225
rect 4937 -4295 4989 -4227
rect 4937 -4389 4942 -4295
rect 4988 -4389 4989 -4295
rect 4937 -4393 4989 -4389
rect 5140 -4295 5192 -4094
rect 5140 -4389 5146 -4295
rect 4942 -4400 4988 -4393
rect 5140 -4449 5192 -4389
rect 4733 -4501 5192 -4449
rect 5344 -4000 5396 -3867
rect 5557 -3891 5566 -3816
rect 5652 -3891 5662 -3816
rect 5557 -3903 5662 -3891
rect 6350 -3838 6374 -3789
rect 6437 -3838 6458 -3789
rect 6350 -3900 6458 -3838
rect 6350 -3949 6374 -3900
rect 6437 -3949 6458 -3900
rect 5344 -4094 5350 -4000
rect 5344 -4143 5396 -4094
rect 5550 -4000 5602 -3981
rect 5550 -4094 5554 -4000
rect 5600 -4094 5602 -4000
rect 5550 -4143 5602 -4094
rect 5344 -4152 5602 -4143
rect 5344 -4203 5439 -4152
rect 5511 -4155 5602 -4152
rect 5677 -4000 5729 -3985
rect 5677 -4094 5682 -4000
rect 5728 -4094 5729 -4000
rect 5677 -4153 5729 -4094
rect 5881 -4000 5933 -3984
rect 5881 -4094 5886 -4000
rect 5932 -4094 5933 -4000
rect 5677 -4155 5818 -4153
rect 5881 -4155 5933 -4094
rect 6086 -4000 6138 -3985
rect 6086 -4094 6090 -4000
rect 6136 -4094 6138 -4000
rect 6086 -4155 6138 -4094
rect 5511 -4162 6138 -4155
rect 5511 -4203 5761 -4162
rect 5817 -4164 6138 -4162
rect 5817 -4166 5975 -4164
rect 5344 -4212 5761 -4203
rect 5344 -4295 5396 -4212
rect 5344 -4389 5350 -4295
rect 4733 -4665 4785 -4501
rect 5344 -4552 5396 -4389
rect 5550 -4218 5761 -4212
rect 5843 -4211 5975 -4166
rect 6047 -4211 6138 -4164
rect 5843 -4216 6138 -4211
rect 5817 -4218 6138 -4216
rect 5550 -4220 6138 -4218
rect 5550 -4225 5933 -4220
rect 5550 -4295 5602 -4225
rect 5550 -4389 5554 -4295
rect 5600 -4389 5602 -4295
rect 5550 -4391 5602 -4389
rect 5677 -4227 5818 -4225
rect 5677 -4295 5729 -4227
rect 5677 -4389 5682 -4295
rect 5728 -4389 5729 -4295
rect 5554 -4400 5600 -4391
rect 5677 -4395 5729 -4389
rect 5881 -4295 5933 -4225
rect 5881 -4389 5886 -4295
rect 5932 -4389 5933 -4295
rect 5881 -4394 5933 -4389
rect 6086 -4295 6138 -4220
rect 6086 -4389 6090 -4295
rect 6136 -4389 6138 -4295
rect 5682 -4400 5728 -4395
rect 5886 -4400 5932 -4394
rect 6086 -4395 6138 -4389
rect 6350 -4011 6458 -3949
rect 6350 -4060 6374 -4011
rect 6437 -4060 6458 -4011
rect 6350 -4122 6458 -4060
rect 6350 -4171 6374 -4122
rect 6437 -4171 6458 -4122
rect 6350 -4233 6458 -4171
rect 6350 -4282 6374 -4233
rect 6437 -4282 6458 -4233
rect 6350 -4344 6458 -4282
rect 6350 -4393 6374 -4344
rect 6437 -4393 6458 -4344
rect 6090 -4400 6136 -4395
rect 4124 -4774 4126 -4680
rect 4172 -4774 4176 -4680
rect 4124 -4849 4176 -4774
rect 4324 -4680 4378 -4667
rect 4324 -4774 4330 -4680
rect 4376 -4774 4378 -4680
rect 4123 -4854 4181 -4849
rect 4324 -4854 4378 -4774
rect 4529 -4680 4581 -4667
rect 4529 -4774 4534 -4680
rect 4580 -4774 4581 -4680
rect 4120 -4858 4190 -4854
rect 4323 -4855 4379 -4854
rect 4120 -4914 4124 -4858
rect 4180 -4914 4190 -4858
rect 4120 -4919 4190 -4914
rect 4311 -4863 4391 -4855
rect 4311 -4917 4324 -4863
rect 4378 -4917 4391 -4863
rect 4123 -4923 4181 -4919
rect 4311 -4920 4391 -4917
rect 3918 -5101 3922 -5007
rect 3968 -5101 3970 -5007
rect 3918 -5160 3970 -5101
rect 4124 -5007 4176 -4923
rect 4323 -4926 4379 -4920
rect 4124 -5101 4126 -5007
rect 4172 -5101 4176 -5007
rect 4124 -5112 4176 -5101
rect 4324 -5007 4378 -4926
rect 4324 -5101 4330 -5007
rect 4376 -5101 4378 -5007
rect 4324 -5110 4378 -5101
rect 4326 -5160 4378 -5110
rect 3918 -5212 4378 -5160
rect 4529 -5007 4581 -4774
rect 4529 -5101 4534 -5007
rect 4580 -5101 4581 -5007
rect 4529 -5265 4581 -5101
rect 4732 -4680 4785 -4665
rect 4939 -4604 5396 -4552
rect 6350 -4455 6458 -4393
rect 6350 -4504 6374 -4455
rect 6437 -4504 6458 -4455
rect 6350 -4566 6458 -4504
rect 4939 -4666 4991 -4604
rect 6350 -4615 6374 -4566
rect 6437 -4615 6458 -4566
rect 4732 -4774 4738 -4680
rect 4784 -4774 4785 -4680
rect 4732 -4793 4785 -4774
rect 4938 -4680 4991 -4666
rect 4938 -4774 4942 -4680
rect 4988 -4774 4991 -4680
rect 4732 -5007 4784 -4793
rect 4732 -5101 4738 -5007
rect 4732 -5160 4784 -5101
rect 4938 -4805 4991 -4774
rect 5144 -4680 5196 -4667
rect 5144 -4774 5146 -4680
rect 5192 -4774 5196 -4680
rect 4938 -5007 4990 -4805
rect 4938 -5101 4942 -5007
rect 4988 -5101 4990 -5007
rect 4938 -5109 4990 -5101
rect 5144 -4994 5196 -4774
rect 5346 -4680 5398 -4665
rect 5346 -4774 5350 -4680
rect 5396 -4774 5398 -4680
rect 5346 -4846 5398 -4774
rect 5549 -4680 5601 -4666
rect 5549 -4774 5554 -4680
rect 5600 -4774 5601 -4680
rect 5549 -4846 5601 -4774
rect 5678 -4680 5730 -4666
rect 5678 -4774 5682 -4680
rect 5728 -4774 5730 -4680
rect 5678 -4846 5730 -4774
rect 5346 -4848 5730 -4846
rect 5886 -4680 5938 -4666
rect 5932 -4774 5938 -4680
rect 5886 -4847 5938 -4774
rect 6086 -4680 6138 -4663
rect 6086 -4774 6090 -4680
rect 6136 -4774 6138 -4680
rect 6086 -4847 6138 -4774
rect 5882 -4848 6138 -4847
rect 5346 -4849 6138 -4848
rect 5333 -4856 6138 -4849
rect 5333 -4864 5439 -4856
rect 5333 -4918 5345 -4864
rect 5399 -4907 5439 -4864
rect 5511 -4859 5975 -4856
rect 5511 -4907 5771 -4859
rect 5399 -4908 5771 -4907
rect 5843 -4903 5975 -4859
rect 6047 -4903 6138 -4856
rect 5843 -4908 6138 -4903
rect 5399 -4912 6138 -4908
rect 5399 -4916 5938 -4912
rect 5399 -4918 5412 -4916
rect 5333 -4929 5412 -4918
rect 5346 -4991 5398 -4929
rect 5144 -5007 5200 -4994
rect 5144 -5101 5146 -5007
rect 5192 -5101 5200 -5007
rect 4942 -5112 4988 -5109
rect 5144 -5110 5200 -5101
rect 5346 -5007 5399 -4991
rect 5346 -5101 5350 -5007
rect 5396 -5101 5399 -5007
rect 5346 -5108 5399 -5101
rect 5146 -5112 5200 -5110
rect 5148 -5160 5200 -5112
rect 4732 -5212 5200 -5160
rect 5347 -5265 5399 -5108
rect 5549 -5007 5601 -4916
rect 5549 -5101 5554 -5007
rect 5600 -5101 5601 -5007
rect 5549 -5109 5601 -5101
rect 5678 -4917 5938 -4916
rect 5678 -5007 5730 -4917
rect 5678 -5101 5682 -5007
rect 5728 -5101 5730 -5007
rect 5678 -5109 5730 -5101
rect 5886 -5007 5938 -4917
rect 5932 -5101 5938 -5007
rect 5886 -5109 5938 -5101
rect 6086 -5007 6138 -4912
rect 6086 -5101 6090 -5007
rect 6136 -5101 6138 -5007
rect 6086 -5106 6138 -5101
rect 6350 -4677 6458 -4615
rect 6350 -4726 6374 -4677
rect 6437 -4726 6458 -4677
rect 6350 -4788 6458 -4726
rect 6350 -4837 6374 -4788
rect 6437 -4837 6458 -4788
rect 6350 -4899 6458 -4837
rect 6350 -4948 6374 -4899
rect 6437 -4948 6458 -4899
rect 6350 -5010 6458 -4948
rect 6350 -5059 6374 -5010
rect 6437 -5059 6458 -5010
rect 5554 -5112 5600 -5109
rect 5682 -5112 5728 -5109
rect 5886 -5112 5932 -5109
rect 6090 -5112 6136 -5106
rect 6350 -5121 6458 -5059
rect 6350 -5170 6374 -5121
rect 6437 -5170 6458 -5121
rect 3714 -5317 5399 -5265
rect 5559 -5200 5662 -5185
rect 5559 -5267 5568 -5200
rect 5652 -5267 5662 -5200
rect 5559 -5276 5576 -5267
rect 5644 -5276 5662 -5267
rect 5559 -5279 5662 -5276
rect 6350 -5232 6458 -5170
rect 5567 -5285 5653 -5279
rect 6350 -5281 6374 -5232
rect 6437 -5281 6458 -5232
rect 3231 -5423 3339 -5361
rect -2144 -5479 -784 -5465
rect -526 -5479 834 -5465
rect -2463 -5492 -2356 -5486
rect -2144 -5492 834 -5479
rect -2463 -5574 -2450 -5492
rect -2398 -5497 834 -5492
rect 1083 -5497 2443 -5465
rect -2398 -5504 2443 -5497
rect -2398 -5509 -1551 -5504
rect -2398 -5560 -2084 -5509
rect -1834 -5550 -1551 -5509
rect -839 -5509 67 -5504
rect -839 -5534 -466 -5509
rect -839 -5550 -784 -5534
rect -1834 -5560 -784 -5550
rect -2398 -5574 -784 -5560
rect -2463 -5593 -2356 -5574
rect -2144 -5578 -784 -5574
rect -526 -5560 -466 -5534
rect -216 -5550 67 -5509
rect 779 -5509 1676 -5504
rect 779 -5550 1143 -5509
rect -216 -5552 1143 -5550
rect -216 -5560 834 -5552
rect -526 -5578 834 -5560
rect 1083 -5560 1143 -5552
rect 1393 -5550 1676 -5509
rect 2388 -5550 2443 -5504
rect 1393 -5560 2443 -5550
rect 1083 -5578 2443 -5560
rect 3231 -5472 3255 -5423
rect 3318 -5472 3339 -5423
rect 3231 -5534 3339 -5472
rect -2068 -5670 -1998 -5578
rect -2068 -5744 -2045 -5670
rect -1999 -5744 -1998 -5670
rect -2068 -5759 -1998 -5744
rect -1886 -5670 -1822 -5657
rect -1886 -5744 -1885 -5670
rect -1839 -5744 -1822 -5670
rect -1704 -5664 -1617 -5646
rect -1704 -5729 -1691 -5664
rect -1626 -5702 -1617 -5664
rect -1626 -5705 -1452 -5702
rect -1626 -5729 -1509 -5705
rect -1704 -5731 -1509 -5729
rect -2144 -5831 -1940 -5825
rect -2278 -5833 -1940 -5831
rect -2278 -5880 -2015 -5833
rect -2278 -5903 -2142 -5880
rect -2167 -5938 -2142 -5903
rect -2084 -5892 -2015 -5880
rect -1952 -5892 -1940 -5833
rect -2084 -5906 -1940 -5892
rect -1886 -5860 -1822 -5744
rect -1698 -5751 -1509 -5731
rect -1463 -5751 -1452 -5705
rect -1698 -5753 -1452 -5751
rect -1354 -5705 -1283 -5578
rect -1354 -5751 -1341 -5705
rect -1295 -5751 -1283 -5705
rect -1354 -5753 -1283 -5751
rect -1109 -5705 -1038 -5578
rect -732 -5614 -643 -5600
rect -732 -5674 -719 -5614
rect -656 -5674 -643 -5614
rect -732 -5687 -643 -5674
rect -450 -5670 -380 -5578
rect -1109 -5751 -1097 -5705
rect -1051 -5751 -1038 -5705
rect -1109 -5753 -1038 -5751
rect -940 -5705 -809 -5704
rect -940 -5751 -929 -5705
rect -883 -5751 -809 -5705
rect -940 -5753 -809 -5751
rect -1698 -5773 -1513 -5753
rect -2084 -5938 -2070 -5906
rect -2167 -5941 -2070 -5938
rect -1886 -5907 -1685 -5860
rect -2071 -6008 -1990 -6003
rect -1886 -6008 -1822 -5907
rect -1732 -5963 -1685 -5907
rect -1732 -5977 -1642 -5963
rect -1732 -5991 -1718 -5977
rect -2071 -6054 -2049 -6008
rect -2003 -6054 -1990 -6008
rect -1892 -6054 -1881 -6008
rect -1835 -6054 -1822 -6008
rect -1731 -6037 -1718 -5991
rect -1655 -6037 -1642 -5977
rect -1731 -6050 -1642 -6037
rect -1584 -6010 -1513 -5773
rect -1441 -5818 -1352 -5805
rect -1441 -5878 -1428 -5818
rect -1365 -5878 -1352 -5818
rect -1441 -5892 -1352 -5878
rect -878 -5822 -809 -5753
rect -450 -5744 -427 -5670
rect -381 -5744 -380 -5670
rect -450 -5759 -380 -5744
rect -268 -5670 -204 -5657
rect -268 -5744 -267 -5670
rect -221 -5744 -204 -5670
rect -86 -5664 1 -5646
rect -86 -5729 -73 -5664
rect -8 -5702 1 -5664
rect -8 -5705 166 -5702
rect -8 -5729 109 -5705
rect -86 -5731 109 -5729
rect -878 -5881 -869 -5822
rect -817 -5827 -809 -5822
rect -761 -5827 -682 -5814
rect -817 -5881 -749 -5827
rect -695 -5881 -682 -5827
rect -878 -6010 -809 -5881
rect -761 -5893 -682 -5881
rect -623 -5833 -322 -5825
rect -623 -5880 -397 -5833
rect -623 -5938 -524 -5880
rect -466 -5892 -397 -5880
rect -334 -5892 -322 -5833
rect -466 -5906 -322 -5892
rect -268 -5860 -204 -5744
rect -80 -5751 109 -5731
rect 155 -5751 166 -5705
rect -80 -5753 166 -5751
rect 264 -5705 335 -5578
rect 264 -5751 277 -5705
rect 323 -5751 335 -5705
rect 264 -5753 335 -5751
rect 509 -5705 580 -5578
rect 886 -5614 975 -5600
rect 886 -5674 899 -5614
rect 962 -5674 975 -5614
rect 886 -5687 975 -5674
rect 1159 -5670 1229 -5578
rect 509 -5751 521 -5705
rect 567 -5751 580 -5705
rect 509 -5753 580 -5751
rect 678 -5705 809 -5704
rect 678 -5751 689 -5705
rect 735 -5751 809 -5705
rect 678 -5753 809 -5751
rect -80 -5773 105 -5753
rect -466 -5938 -452 -5906
rect -623 -5941 -452 -5938
rect -268 -5907 -67 -5860
rect -623 -5949 -545 -5941
rect -2071 -6165 -1990 -6054
rect -1886 -6055 -1822 -6054
rect -1584 -6056 -1571 -6010
rect -1525 -6056 -1513 -6010
rect -1584 -6057 -1513 -6056
rect -1415 -6056 -1403 -6010
rect -1357 -6056 -1343 -6010
rect -1415 -6165 -1343 -6056
rect -1047 -6056 -1035 -6010
rect -989 -6056 -977 -6010
rect -1047 -6165 -977 -6056
rect -878 -6056 -867 -6010
rect -821 -6056 -809 -6010
rect -878 -6057 -809 -6056
rect -453 -6008 -372 -6003
rect -268 -6008 -204 -5907
rect -114 -5963 -67 -5907
rect -114 -5977 -24 -5963
rect -114 -5991 -100 -5977
rect -453 -6054 -431 -6008
rect -385 -6054 -372 -6008
rect -274 -6054 -263 -6008
rect -217 -6054 -204 -6008
rect -113 -6037 -100 -5991
rect -37 -6037 -24 -5977
rect -113 -6050 -24 -6037
rect 34 -6010 105 -5773
rect 177 -5818 266 -5805
rect 177 -5878 190 -5818
rect 253 -5878 266 -5818
rect 177 -5892 266 -5878
rect 740 -5822 809 -5753
rect 1159 -5744 1182 -5670
rect 1228 -5744 1229 -5670
rect 1159 -5759 1229 -5744
rect 1341 -5670 1405 -5657
rect 1341 -5744 1342 -5670
rect 1388 -5744 1405 -5670
rect 1523 -5664 1610 -5646
rect 1523 -5729 1536 -5664
rect 1601 -5702 1610 -5664
rect 1601 -5705 1775 -5702
rect 1601 -5729 1718 -5705
rect 1523 -5731 1718 -5729
rect 740 -5881 749 -5822
rect 801 -5881 809 -5822
rect 740 -6010 809 -5881
rect 968 -5833 1287 -5825
rect 968 -5880 1212 -5833
rect 968 -5906 1085 -5880
rect 1060 -5938 1085 -5906
rect 1143 -5892 1212 -5880
rect 1275 -5892 1287 -5833
rect 1143 -5906 1287 -5892
rect 1341 -5860 1405 -5744
rect 1529 -5751 1718 -5731
rect 1764 -5751 1775 -5705
rect 1529 -5753 1775 -5751
rect 1873 -5705 1944 -5578
rect 1873 -5751 1886 -5705
rect 1932 -5751 1944 -5705
rect 1873 -5753 1944 -5751
rect 2118 -5705 2189 -5578
rect 3231 -5583 3255 -5534
rect 3318 -5583 3339 -5534
rect 2495 -5614 2584 -5600
rect 2495 -5674 2508 -5614
rect 2571 -5674 2584 -5614
rect 2495 -5687 2584 -5674
rect 3231 -5645 3339 -5583
rect 3231 -5694 3255 -5645
rect 3318 -5694 3339 -5645
rect 2118 -5751 2130 -5705
rect 2176 -5751 2189 -5705
rect 2118 -5753 2189 -5751
rect 2287 -5705 2418 -5704
rect 2287 -5751 2298 -5705
rect 2344 -5751 2418 -5705
rect 2287 -5753 2418 -5751
rect 1529 -5773 1714 -5753
rect 1143 -5938 1157 -5906
rect 1060 -5941 1157 -5938
rect 1341 -5907 1542 -5860
rect -730 -6072 -641 -6058
rect -730 -6132 -717 -6072
rect -654 -6132 -641 -6072
rect -730 -6145 -641 -6132
rect -453 -6165 -372 -6054
rect -268 -6055 -204 -6054
rect 34 -6056 47 -6010
rect 93 -6056 105 -6010
rect 34 -6057 105 -6056
rect 203 -6056 215 -6010
rect 261 -6056 275 -6010
rect 203 -6165 275 -6056
rect 571 -6056 583 -6010
rect 629 -6056 641 -6010
rect 571 -6165 641 -6056
rect 740 -6056 751 -6010
rect 797 -6056 809 -6010
rect 740 -6057 809 -6056
rect 1156 -6008 1237 -6003
rect 1341 -6008 1405 -5907
rect 1495 -5963 1542 -5907
rect 1495 -5977 1585 -5963
rect 1495 -5991 1509 -5977
rect 1156 -6054 1178 -6008
rect 1224 -6054 1237 -6008
rect 1335 -6054 1346 -6008
rect 1392 -6054 1405 -6008
rect 1496 -6037 1509 -5991
rect 1572 -6037 1585 -5977
rect 1496 -6050 1585 -6037
rect 1643 -6010 1714 -5773
rect 1786 -5818 1875 -5805
rect 1786 -5878 1799 -5818
rect 1862 -5878 1875 -5818
rect 1786 -5892 1875 -5878
rect 2349 -5822 2418 -5753
rect 2349 -5881 2358 -5822
rect 2410 -5881 2418 -5822
rect 2349 -6010 2418 -5881
rect 888 -6072 977 -6058
rect 888 -6132 901 -6072
rect 964 -6132 977 -6072
rect 888 -6145 977 -6132
rect 1156 -6165 1237 -6054
rect 1341 -6055 1405 -6054
rect 1643 -6056 1656 -6010
rect 1702 -6056 1714 -6010
rect 1643 -6057 1714 -6056
rect 1812 -6056 1824 -6010
rect 1870 -6056 1884 -6010
rect 1812 -6165 1884 -6056
rect 2180 -6056 2192 -6010
rect 2238 -6056 2250 -6010
rect 2180 -6165 2250 -6056
rect 2349 -6056 2360 -6010
rect 2406 -6056 2418 -6010
rect 2349 -6057 2418 -6056
rect 3231 -5756 3339 -5694
rect 3231 -5805 3255 -5756
rect 3318 -5805 3339 -5756
rect 3511 -5396 3564 -5379
rect 3511 -5490 3514 -5396
rect 3560 -5490 3564 -5396
rect 3511 -5545 3564 -5490
rect 3716 -5396 3769 -5382
rect 3716 -5490 3718 -5396
rect 3764 -5490 3769 -5396
rect 3716 -5545 3769 -5490
rect 3511 -5553 3769 -5545
rect 3919 -5396 3972 -5378
rect 3919 -5490 3922 -5396
rect 3968 -5490 3972 -5396
rect 3511 -5554 3781 -5553
rect 3511 -5604 3603 -5554
rect 3674 -5562 3781 -5554
rect 3674 -5604 3716 -5562
rect 3511 -5613 3716 -5604
rect 3511 -5691 3564 -5613
rect 3706 -5616 3716 -5613
rect 3770 -5616 3781 -5562
rect 3706 -5626 3781 -5616
rect 3511 -5785 3514 -5691
rect 3560 -5785 3564 -5691
rect 3511 -5798 3564 -5785
rect 3716 -5691 3769 -5626
rect 3716 -5785 3718 -5691
rect 3764 -5785 3769 -5691
rect 3231 -5867 3339 -5805
rect 3231 -5916 3255 -5867
rect 3318 -5916 3339 -5867
rect 3231 -5978 3339 -5916
rect 3458 -5882 3539 -5872
rect 3458 -5944 3469 -5882
rect 3531 -5944 3539 -5882
rect 3458 -5949 3470 -5944
rect 3530 -5949 3539 -5944
rect 3461 -5958 3539 -5949
rect 3716 -5952 3769 -5785
rect 3919 -5691 3972 -5490
rect 3919 -5785 3922 -5691
rect 3968 -5785 3972 -5691
rect 3919 -5844 3972 -5785
rect 4122 -5396 4175 -5317
rect 4122 -5490 4126 -5396
rect 4172 -5490 4175 -5396
rect 4122 -5691 4175 -5490
rect 4328 -5396 4381 -5381
rect 4328 -5490 4330 -5396
rect 4376 -5490 4381 -5396
rect 4328 -5569 4381 -5490
rect 4531 -5396 4584 -5378
rect 4531 -5490 4534 -5396
rect 4580 -5490 4584 -5396
rect 4310 -5572 4388 -5569
rect 4310 -5628 4323 -5572
rect 4379 -5628 4388 -5572
rect 4310 -5637 4388 -5628
rect 4122 -5785 4126 -5691
rect 4172 -5785 4175 -5691
rect 4122 -5798 4175 -5785
rect 4326 -5691 4381 -5637
rect 4326 -5785 4330 -5691
rect 4376 -5785 4381 -5691
rect 4326 -5797 4381 -5785
rect 4531 -5691 4584 -5490
rect 4733 -5396 4786 -5375
rect 4733 -5490 4738 -5396
rect 4784 -5490 4786 -5396
rect 4733 -5563 4786 -5490
rect 4937 -5396 4990 -5317
rect 6350 -5343 6458 -5281
rect 4937 -5490 4942 -5396
rect 4988 -5490 4990 -5396
rect 4937 -5549 4990 -5490
rect 5142 -5396 5195 -5374
rect 5142 -5490 5146 -5396
rect 5192 -5490 5195 -5396
rect 4936 -5555 4992 -5549
rect 4924 -5558 5005 -5555
rect 4728 -5574 4800 -5563
rect 4728 -5630 4734 -5574
rect 4790 -5630 4800 -5574
rect 4924 -5612 4937 -5558
rect 4991 -5612 5005 -5558
rect 4924 -5617 5005 -5612
rect 4936 -5621 4992 -5617
rect 4728 -5641 4800 -5630
rect 4531 -5785 4534 -5691
rect 4580 -5785 4584 -5691
rect 4326 -5844 4380 -5797
rect 4531 -5814 4584 -5785
rect 4733 -5691 4786 -5641
rect 4733 -5785 4738 -5691
rect 4784 -5785 4786 -5691
rect 4530 -5818 4586 -5814
rect 3919 -5897 4380 -5844
rect 4519 -5823 4597 -5818
rect 4519 -5877 4531 -5823
rect 4585 -5877 4597 -5823
rect 4519 -5885 4597 -5877
rect 4733 -5843 4786 -5785
rect 4937 -5691 4990 -5621
rect 4937 -5785 4942 -5691
rect 4988 -5785 4990 -5691
rect 4937 -5789 4990 -5785
rect 5142 -5691 5195 -5490
rect 5142 -5785 5146 -5691
rect 5192 -5785 5195 -5691
rect 4942 -5796 4988 -5789
rect 5142 -5843 5195 -5785
rect 4530 -5886 4586 -5885
rect 4109 -5952 4189 -5943
rect 3231 -6027 3255 -5978
rect 3318 -6027 3339 -5978
rect 3716 -6005 4121 -5952
rect 4109 -6008 4121 -6005
rect 4177 -6008 4189 -5952
rect 4109 -6018 4189 -6008
rect 2497 -6072 2586 -6058
rect 2497 -6132 2510 -6072
rect 2573 -6132 2586 -6072
rect 2497 -6145 2586 -6132
rect 3231 -6089 3339 -6027
rect 3231 -6138 3255 -6089
rect 3318 -6138 3339 -6089
rect -2323 -6185 -2232 -6180
rect -2144 -6185 -784 -6165
rect -2323 -6186 -784 -6185
rect -2323 -6253 -2310 -6186
rect -2243 -6198 -784 -6186
rect -2243 -6200 -1567 -6198
rect -2243 -6249 -2099 -6200
rect -1790 -6244 -1567 -6200
rect -838 -6199 -784 -6198
rect -526 -6198 834 -6165
rect -526 -6199 51 -6198
rect -838 -6200 51 -6199
rect -838 -6244 -481 -6200
rect -1790 -6249 -481 -6244
rect -172 -6244 51 -6200
rect 780 -6204 834 -6198
rect 1083 -6193 2443 -6165
rect 3231 -6193 3339 -6138
rect 1083 -6198 3339 -6193
rect 1083 -6200 1660 -6198
rect 1083 -6204 1128 -6200
rect 780 -6244 1128 -6204
rect -172 -6249 1128 -6244
rect 1437 -6244 1660 -6200
rect 2389 -6200 3339 -6198
rect 2389 -6244 3255 -6200
rect 1437 -6247 3255 -6244
rect 1437 -6249 2443 -6247
rect -2243 -6252 2443 -6249
rect -2243 -6253 -2232 -6252
rect -2323 -6264 -2232 -6253
rect -2144 -6253 2443 -6252
rect -2144 -6278 -784 -6253
rect -526 -6258 2443 -6253
rect -526 -6278 834 -6258
rect 1083 -6278 2443 -6258
rect 3231 -6249 3255 -6247
rect 3318 -6249 3339 -6200
rect 3231 -6311 3339 -6249
rect 3512 -6076 3563 -6053
rect 3512 -6170 3514 -6076
rect 3560 -6170 3563 -6076
rect 3512 -6217 3563 -6170
rect 3716 -6076 3767 -6056
rect 3716 -6170 3718 -6076
rect 3764 -6170 3767 -6076
rect 3716 -6217 3767 -6170
rect 3512 -6228 3767 -6217
rect 3512 -6280 3603 -6228
rect 3675 -6280 3767 -6228
rect 3512 -6290 3767 -6280
rect 3920 -6076 3971 -6058
rect 3920 -6170 3922 -6076
rect 3968 -6170 3971 -6076
rect 3920 -6230 3971 -6170
rect 4123 -6076 4177 -6018
rect 4329 -6057 4380 -5897
rect 4123 -6170 4126 -6076
rect 4172 -6170 4177 -6076
rect 4123 -6178 4177 -6170
rect 4327 -6076 4380 -6057
rect 4733 -5896 5195 -5843
rect 5348 -5396 5401 -5376
rect 5348 -5490 5350 -5396
rect 5396 -5490 5401 -5396
rect 5348 -5549 5401 -5490
rect 5550 -5396 5603 -5382
rect 5550 -5490 5554 -5396
rect 5600 -5490 5603 -5396
rect 5550 -5549 5603 -5490
rect 5678 -5396 5731 -5384
rect 5678 -5490 5682 -5396
rect 5728 -5490 5731 -5396
rect 5678 -5542 5731 -5490
rect 5882 -5396 5935 -5384
rect 5882 -5490 5886 -5396
rect 5932 -5490 5935 -5396
rect 5882 -5542 5935 -5490
rect 6085 -5396 6138 -5383
rect 6085 -5490 6090 -5396
rect 6136 -5490 6138 -5396
rect 6085 -5542 6138 -5490
rect 5678 -5549 6138 -5542
rect 5348 -5551 6138 -5549
rect 5348 -5552 5975 -5551
rect 5348 -5559 5771 -5552
rect 5348 -5605 5439 -5559
rect 5511 -5602 5771 -5559
rect 5843 -5602 5975 -5552
rect 5511 -5604 5975 -5602
rect 6047 -5604 6138 -5551
rect 5511 -5605 6138 -5604
rect 5348 -5612 6138 -5605
rect 5348 -5614 5731 -5612
rect 5348 -5691 5401 -5614
rect 5348 -5785 5350 -5691
rect 5396 -5785 5401 -5691
rect 4327 -6170 4330 -6076
rect 4376 -6170 4380 -6076
rect 4126 -6181 4172 -6178
rect 4327 -6180 4380 -6170
rect 4329 -6230 4380 -6180
rect 3920 -6281 4380 -6230
rect 4531 -6076 4582 -6058
rect 4531 -6170 4534 -6076
rect 4580 -6170 4582 -6076
rect 3512 -6291 3563 -6290
rect 3231 -6360 3255 -6311
rect 3318 -6360 3339 -6311
rect 3231 -6422 3339 -6360
rect 3716 -6328 3767 -6290
rect 4531 -6328 4582 -6170
rect 4733 -6060 4786 -5896
rect 5348 -5944 5401 -5785
rect 5550 -5691 5603 -5614
rect 5550 -5785 5554 -5691
rect 5600 -5785 5603 -5691
rect 5550 -5789 5603 -5785
rect 5678 -5691 5731 -5614
rect 5678 -5785 5682 -5691
rect 5728 -5785 5731 -5691
rect 5554 -5796 5600 -5789
rect 5678 -5791 5731 -5785
rect 5882 -5613 6138 -5612
rect 5882 -5691 5935 -5613
rect 5882 -5785 5886 -5691
rect 5932 -5785 5935 -5691
rect 5882 -5791 5935 -5785
rect 6085 -5691 6138 -5613
rect 6085 -5785 6090 -5691
rect 6136 -5785 6138 -5691
rect 6085 -5790 6138 -5785
rect 6350 -5392 6374 -5343
rect 6437 -5392 6458 -5343
rect 6350 -5454 6458 -5392
rect 6350 -5503 6374 -5454
rect 6437 -5503 6458 -5454
rect 6350 -5565 6458 -5503
rect 6350 -5614 6374 -5565
rect 6437 -5614 6458 -5565
rect 6350 -5676 6458 -5614
rect 6350 -5725 6374 -5676
rect 6437 -5725 6458 -5676
rect 6350 -5787 6458 -5725
rect 5682 -5796 5728 -5791
rect 5886 -5796 5932 -5791
rect 6090 -5796 6136 -5790
rect 6350 -5836 6374 -5787
rect 6437 -5836 6458 -5787
rect 6350 -5898 6458 -5836
rect 4926 -5953 5401 -5944
rect 4926 -6007 4938 -5953
rect 4992 -5997 5401 -5953
rect 5520 -5929 5601 -5920
rect 5520 -5988 5529 -5929
rect 5588 -5950 5601 -5929
rect 6350 -5947 6374 -5898
rect 6437 -5947 6458 -5898
rect 5588 -5962 6137 -5950
rect 5588 -5988 5975 -5962
rect 5520 -5997 5975 -5988
rect 4992 -6007 5004 -5997
rect 4926 -6019 5004 -6007
rect 5550 -6011 5975 -5997
rect 6047 -6011 6137 -5962
rect 4733 -6076 4789 -6060
rect 4733 -6170 4738 -6076
rect 4784 -6170 4789 -6076
rect 4733 -6231 4789 -6170
rect 4938 -6076 4991 -6019
rect 5550 -6021 6137 -6011
rect 5349 -6056 5400 -6052
rect 4938 -6170 4942 -6076
rect 4988 -6170 4991 -6076
rect 4938 -6185 4991 -6170
rect 5144 -6076 5195 -6058
rect 5144 -6170 5146 -6076
rect 5192 -6170 5195 -6076
rect 5144 -6231 5195 -6170
rect 5347 -6076 5400 -6056
rect 5347 -6170 5350 -6076
rect 5396 -6170 5400 -6076
rect 5347 -6179 5400 -6170
rect 5550 -6076 5601 -6021
rect 5550 -6170 5554 -6076
rect 5600 -6170 5601 -6076
rect 5550 -6179 5601 -6170
rect 5679 -6076 5730 -6021
rect 5679 -6170 5682 -6076
rect 5728 -6170 5730 -6076
rect 4733 -6282 5195 -6231
rect 5349 -6328 5400 -6179
rect 5554 -6181 5600 -6179
rect 5679 -6183 5730 -6170
rect 5883 -6076 5934 -6021
rect 5883 -6170 5886 -6076
rect 5932 -6170 5934 -6076
rect 3716 -6375 5400 -6328
rect 3716 -6379 4936 -6375
rect 3231 -6471 3255 -6422
rect 3318 -6471 3339 -6422
rect 4922 -6431 4936 -6379
rect 4992 -6379 5400 -6375
rect 4992 -6431 5005 -6379
rect 4922 -6437 5005 -6431
rect 5349 -6436 5400 -6379
rect 5561 -6286 5676 -6277
rect 5561 -6294 5598 -6286
rect 5561 -6363 5576 -6294
rect 5664 -6352 5676 -6286
rect 5645 -6363 5676 -6352
rect 5561 -6381 5676 -6363
rect 5883 -6436 5934 -6170
rect 6086 -6076 6137 -6021
rect 6086 -6170 6090 -6076
rect 6136 -6170 6137 -6076
rect 6086 -6180 6137 -6170
rect 6350 -6009 6458 -5947
rect 6350 -6058 6374 -6009
rect 6437 -6058 6458 -6009
rect 6350 -6120 6458 -6058
rect 6350 -6169 6374 -6120
rect 6437 -6169 6458 -6120
rect 6090 -6181 6136 -6180
rect 3231 -6591 3339 -6471
rect 5349 -6487 5934 -6436
rect 5883 -6489 5934 -6487
rect 6350 -6231 6458 -6169
rect 6350 -6280 6374 -6231
rect 6437 -6280 6458 -6231
rect 6350 -6342 6458 -6280
rect 6350 -6391 6374 -6342
rect 6437 -6391 6458 -6342
rect 6350 -6453 6458 -6391
rect 6350 -6502 6374 -6453
rect 6437 -6502 6458 -6453
rect 6350 -6591 6458 -6502
rect 3231 -6611 6461 -6591
rect 3231 -6660 3318 -6611
rect 3381 -6612 6461 -6611
rect 3381 -6660 3439 -6612
rect 3231 -6661 3439 -6660
rect 3502 -6661 3560 -6612
rect 3623 -6661 3681 -6612
rect 3744 -6661 3802 -6612
rect 3865 -6661 3923 -6612
rect 3986 -6661 4044 -6612
rect 4107 -6661 4165 -6612
rect 4228 -6661 4286 -6612
rect 4349 -6661 4407 -6612
rect 4470 -6661 4528 -6612
rect 4591 -6661 4649 -6612
rect 4712 -6661 4770 -6612
rect 4833 -6661 4891 -6612
rect 4954 -6661 5012 -6612
rect 5075 -6661 5133 -6612
rect 5196 -6661 5254 -6612
rect 5317 -6661 5375 -6612
rect 5438 -6661 5496 -6612
rect 5559 -6661 5617 -6612
rect 5680 -6661 5738 -6612
rect 5801 -6661 5859 -6612
rect 5922 -6661 5980 -6612
rect 6043 -6661 6101 -6612
rect 6164 -6661 6461 -6612
rect 3231 -6677 6461 -6661
rect 6272 -6678 6461 -6677
<< via1 >>
rect 3933 2263 3989 2319
rect 4703 2269 4766 2334
rect -14 1938 42 1957
rect -14 1901 42 1938
rect -1763 1373 -1709 1427
rect -1375 1371 -1321 1425
rect -968 1364 -914 1418
rect -156 1363 -100 1419
rect -559 1196 -556 1233
rect -556 1196 -510 1233
rect -510 1196 -503 1233
rect -559 1177 -503 1196
rect 662 1363 718 1419
rect 253 1196 260 1237
rect 260 1196 306 1237
rect 306 1196 310 1237
rect 253 1180 310 1196
rect 1477 1363 1533 1419
rect 1070 1196 1076 1245
rect 1076 1196 1122 1245
rect 1122 1196 1126 1245
rect 1070 1189 1126 1196
rect 1886 1196 1892 1248
rect 1892 1196 1938 1248
rect 1938 1196 1942 1248
rect 1886 1192 1942 1196
rect 3538 1782 3625 1787
rect 3538 1705 3542 1782
rect 3542 1705 3619 1782
rect 3619 1705 3625 1782
rect 3538 1700 3625 1705
rect 3759 1693 3825 1759
rect 3928 1687 3997 1756
rect 3587 1565 3643 1621
rect 4704 1623 4765 1684
rect 5034 1623 5095 1643
rect 5034 1582 5093 1623
rect 5093 1582 5095 1623
rect 5581 1634 5643 1636
rect 5581 1584 5643 1634
rect 5581 1574 5643 1584
rect 5023 1337 5077 1391
rect -1375 933 -1321 987
rect 3581 1128 3637 1184
rect 3784 1130 3838 1184
rect 5932 1333 5988 1389
rect -559 932 -503 988
rect 253 932 309 988
rect 1067 932 1123 988
rect 1886 932 1942 988
rect 1683 623 1737 677
rect 3588 966 3649 1027
rect 4270 967 4329 1026
rect 3471 774 3474 796
rect 3474 774 3544 796
rect 3471 723 3544 774
rect 3900 754 3969 823
rect 5039 744 5102 822
rect -1762 205 -1708 259
rect -1559 -72 -1503 -16
rect -1150 -72 -1094 -16
rect 49 266 103 320
rect -615 -80 -561 -26
rect -819 -466 -765 -412
rect -80 -41 -26 13
rect -284 -325 -230 -271
rect 583 -42 639 14
rect 1115 -97 1171 -41
rect 789 -326 845 -270
rect 2278 204 2334 260
rect 1657 -46 1713 10
rect 2067 -46 2123 10
rect 2971 589 3027 645
rect 3528 484 3582 538
rect 3928 645 3989 672
rect 3928 611 3939 645
rect 3939 611 3985 645
rect 3985 611 3989 645
rect 4687 700 4758 708
rect 4687 637 4695 700
rect 4695 637 4758 700
rect 4687 629 4758 637
rect 5471 600 5474 656
rect 5474 600 5520 656
rect 5520 600 5527 656
rect 4342 483 4398 539
rect 5876 755 5932 811
rect 5278 443 5334 499
rect 3362 135 3432 205
rect 3160 -105 3216 -49
rect 1341 -438 1397 -382
rect -1376 -1158 -1322 -1104
rect -561 -1159 -505 -1103
rect 256 -1159 312 -1103
rect 1071 -1159 1127 -1103
rect 2312 -780 2372 -720
rect 1681 -859 1737 -803
rect 1894 -1159 1950 -1103
rect 3158 -257 3214 -235
rect 3158 -291 3167 -257
rect 3167 -291 3213 -257
rect 3213 -291 3214 -257
rect 3568 -124 3624 -68
rect 4969 184 5025 237
rect 4969 181 5025 184
rect 4421 91 4482 97
rect 4421 45 4430 91
rect 4430 45 4476 91
rect 4476 45 4482 91
rect 4421 36 4482 45
rect 5094 42 5150 98
rect 3977 -116 4033 -60
rect 3973 -257 4034 -232
rect 3973 -293 3983 -257
rect 3983 -293 4029 -257
rect 4029 -293 4034 -257
rect 3161 -836 3215 -782
rect 3570 -688 3624 -634
rect 3569 -843 3623 -789
rect 4672 -686 4728 -630
rect 3978 -813 4032 -759
rect -1756 -1604 -1700 -1548
rect -1376 -1598 -1322 -1544
rect -562 -1599 -506 -1543
rect 255 -1599 311 -1543
rect 1071 -1599 1127 -1543
rect 1885 -1599 1941 -1543
rect 5095 -848 5149 -794
rect 4796 -984 4850 -930
rect 3161 -1238 3215 -1184
rect 4673 -1240 4727 -1186
rect 3868 -1390 3928 -1330
rect 3805 -1707 3873 -1690
rect 3805 -1756 3807 -1707
rect 3807 -1756 3873 -1707
rect 3805 -1758 3873 -1756
rect 1939 -2076 2001 -2014
rect 3536 -1883 3592 -1827
rect 4058 -1901 4114 -1845
rect 5475 -1886 5531 -1830
rect -2482 -2966 -2399 -2886
rect -1691 -3134 -1626 -3069
rect -2142 -3343 -2084 -3285
rect -719 -3079 -656 -3019
rect -569 -3091 -484 -3006
rect -1428 -3283 -1365 -3223
rect -869 -3286 -817 -3227
rect -617 -3298 -549 -3230
rect 346 -3279 354 -3222
rect 354 -3279 400 -3222
rect 400 -3279 403 -3222
rect 2089 -2836 2145 -2780
rect -717 -3537 -654 -3477
rect 1757 -3120 1813 -3064
rect 1948 -3365 2005 -3354
rect 1948 -3411 2005 -3365
rect -2310 -3658 -2245 -3593
rect -2450 -3827 -2398 -3745
rect 647 -3605 703 -3549
rect -1691 -4002 -1626 -3937
rect -2142 -4211 -2084 -4153
rect -719 -3947 -656 -3887
rect -475 -3947 -413 -3885
rect -1428 -4151 -1365 -4091
rect -869 -4154 -817 -4095
rect -630 -4158 -563 -4091
rect 556 -3812 558 -3783
rect 558 -3812 604 -3783
rect 604 -3812 610 -3783
rect 556 -3837 610 -3812
rect -717 -4405 -654 -4345
rect -2310 -4530 -2243 -4463
rect 146 -4107 203 -4097
rect 146 -4154 150 -4107
rect 150 -4154 196 -4107
rect 196 -4154 203 -4107
rect -2450 -4684 -2398 -4602
rect -1691 -4861 -1626 -4796
rect -2142 -5070 -2084 -5012
rect -719 -4806 -656 -4746
rect -517 -4805 -458 -4746
rect 176 -4683 179 -4618
rect 179 -4683 241 -4618
rect -1428 -5010 -1365 -4950
rect -869 -5013 -817 -4954
rect -630 -5013 -570 -4953
rect 601 -4321 657 -4265
rect 1166 -3606 1224 -3548
rect 1054 -4047 1108 -3993
rect 1368 -3812 1374 -3781
rect 1374 -3812 1420 -3781
rect 1420 -3812 1425 -3781
rect 1368 -3838 1425 -3812
rect 4244 -2126 4314 -2115
rect 4244 -2184 4256 -2126
rect 4256 -2184 4314 -2126
rect 4244 -2185 4314 -2184
rect 3875 -2523 3929 -2469
rect 4431 -2517 4485 -2463
rect 5122 -2518 5178 -2462
rect 3768 -2809 3834 -2801
rect 3768 -2860 3826 -2809
rect 3826 -2860 3834 -2809
rect 3768 -2868 3834 -2860
rect 5666 -2517 5720 -2463
rect 4046 -3145 4100 -3091
rect 4245 -3192 4313 -3184
rect 4245 -3249 4305 -3192
rect 4305 -3249 4313 -3192
rect 4245 -3257 4313 -3249
rect 5762 -3151 5816 -3097
rect 4045 -3424 4101 -3368
rect 3568 -3492 3576 -3440
rect 3576 -3492 3646 -3440
rect 3646 -3492 3654 -3440
rect 3568 -3500 3654 -3492
rect 4326 -3553 4380 -3499
rect 5078 -3441 5134 -3385
rect 4738 -3554 4794 -3498
rect 1367 -4053 1423 -3997
rect 988 -4329 1045 -4272
rect 962 -4787 1018 -4779
rect 962 -4835 966 -4787
rect 966 -4835 1012 -4787
rect 1012 -4835 1018 -4787
rect 1773 -4176 1782 -4119
rect 1782 -4176 1828 -4119
rect 1828 -4176 1830 -4119
rect 1368 -4635 1422 -4581
rect 1777 -4851 1782 -4795
rect 1782 -4851 1828 -4795
rect 1828 -4851 1833 -4795
rect 652 -5003 709 -4946
rect 1572 -5043 1626 -4989
rect -717 -5264 -654 -5204
rect -2310 -5380 -2243 -5313
rect 4122 -3868 4176 -3814
rect 3468 -4497 3545 -4489
rect 3468 -4543 3476 -4497
rect 3476 -4543 3537 -4497
rect 3537 -4543 3545 -4497
rect 4530 -4000 4584 -3949
rect 4530 -4003 4534 -4000
rect 4534 -4003 4580 -4000
rect 4580 -4003 4584 -4000
rect 4122 -4244 4178 -4188
rect 4941 -3869 4997 -3813
rect 4938 -4223 4994 -4167
rect 5566 -3883 5574 -3816
rect 5574 -3883 5644 -3816
rect 5644 -3883 5652 -3816
rect 5566 -3891 5652 -3883
rect 5761 -4166 5817 -4162
rect 5761 -4216 5771 -4166
rect 5771 -4216 5817 -4166
rect 5761 -4218 5817 -4216
rect 4124 -4914 4180 -4858
rect 4324 -4917 4378 -4863
rect 5345 -4918 5399 -4864
rect 5568 -5208 5652 -5200
rect 5568 -5267 5576 -5208
rect 5576 -5267 5644 -5208
rect 5644 -5267 5652 -5208
rect -2450 -5574 -2398 -5492
rect -1691 -5729 -1626 -5664
rect -2142 -5938 -2084 -5880
rect -719 -5674 -656 -5614
rect -1428 -5878 -1365 -5818
rect -73 -5729 -8 -5664
rect -869 -5881 -817 -5822
rect -749 -5881 -695 -5827
rect -524 -5938 -466 -5880
rect 899 -5674 962 -5614
rect 190 -5878 253 -5818
rect 1536 -5729 1601 -5664
rect 749 -5881 801 -5822
rect 1085 -5938 1143 -5880
rect 2508 -5674 2571 -5614
rect -717 -6132 -654 -6072
rect 1799 -5878 1862 -5818
rect 2358 -5881 2410 -5822
rect 901 -6132 964 -6072
rect 3716 -5616 3770 -5562
rect 3469 -5889 3531 -5882
rect 3469 -5944 3470 -5889
rect 3470 -5944 3530 -5889
rect 3530 -5944 3531 -5889
rect 4323 -5628 4379 -5572
rect 4734 -5630 4790 -5574
rect 4937 -5612 4991 -5558
rect 4531 -5877 4585 -5823
rect 4121 -6008 4177 -5952
rect 2510 -6132 2573 -6072
rect -2310 -6253 -2243 -6186
rect 4938 -6007 4992 -5953
rect 4936 -6431 4992 -6375
rect 5576 -6352 5598 -6294
rect 5598 -6352 5645 -6294
rect 5576 -6363 5645 -6352
<< metal2 >>
rect 4691 2334 4779 2347
rect 3923 2319 4000 2330
rect 3923 2263 3933 2319
rect 3989 2263 4000 2319
rect 3923 2247 4000 2263
rect 4691 2269 4703 2334
rect 4766 2269 4779 2334
rect 4691 2252 4779 2269
rect -21 1957 50 1971
rect -21 1901 -14 1957
rect 42 1901 50 1957
rect -21 1897 50 1901
rect -1774 1428 -1697 1439
rect -1904 1427 -1697 1428
rect -1904 1373 -1763 1427
rect -1709 1373 -1697 1427
rect -1904 1372 -1697 1373
rect -1904 -1548 -1848 1372
rect -1774 1360 -1697 1372
rect -1384 1426 -1311 1437
rect -1384 1425 -1178 1426
rect -1384 1371 -1375 1425
rect -1321 1371 -1178 1425
rect -1384 1370 -1178 1371
rect -1384 1362 -1311 1370
rect -1234 1166 -1178 1370
rect -978 1419 -904 1431
rect -158 1419 -97 1431
rect -14 1419 42 1897
rect 3524 1787 3636 1799
rect 3524 1700 3538 1787
rect 3625 1700 3636 1787
rect 3933 1771 3989 2247
rect 3524 1688 3636 1700
rect 3746 1759 3837 1769
rect 3746 1693 3759 1759
rect 3825 1693 3837 1759
rect 3746 1686 3837 1693
rect 3916 1756 4009 1771
rect 3916 1687 3928 1756
rect 3997 1687 4009 1756
rect 4703 1700 4766 2252
rect 3916 1675 4009 1687
rect 4683 1684 4786 1700
rect 3575 1621 3651 1625
rect 3575 1565 3587 1621
rect 3643 1565 3839 1621
rect 3575 1563 3651 1565
rect 660 1419 721 1431
rect 1474 1419 1542 1431
rect -978 1418 -156 1419
rect -978 1364 -968 1418
rect -914 1364 -156 1418
rect -978 1363 -156 1364
rect -100 1363 662 1419
rect 718 1363 1477 1419
rect 1533 1363 1542 1419
rect -978 1351 -904 1363
rect -158 1351 -97 1363
rect 660 1351 721 1363
rect 1474 1351 1542 1363
rect 1874 1256 1942 1257
rect 1070 1248 1126 1254
rect 1874 1248 1955 1256
rect -572 1233 -490 1242
rect -572 1177 -559 1233
rect -503 1177 -490 1233
rect -572 1166 -490 1177
rect 241 1237 323 1246
rect 241 1180 253 1237
rect 310 1180 323 1237
rect 241 1166 323 1180
rect 1058 1245 1138 1248
rect 1058 1189 1070 1245
rect 1126 1189 1138 1245
rect 1058 1166 1138 1189
rect 1874 1192 1886 1248
rect 1942 1192 1955 1248
rect 1874 1166 1955 1192
rect 3578 1184 3649 1189
rect 3783 1186 3839 1565
rect 3933 1555 3989 1675
rect 4683 1623 4704 1684
rect 4765 1623 4786 1684
rect 4683 1610 4786 1623
rect 5010 1643 5104 1651
rect 5010 1582 5034 1643
rect 5095 1582 5104 1643
rect 5010 1569 5104 1582
rect 5564 1636 5656 1644
rect 5564 1574 5581 1636
rect 5643 1574 5656 1636
rect 5564 1559 5656 1574
rect 3933 1499 4535 1555
rect -1234 1110 1955 1166
rect 2566 1128 3581 1184
rect 3637 1128 3649 1184
rect -1385 988 -1314 1000
rect -564 988 -499 1001
rect 244 988 319 998
rect 1063 988 1127 1002
rect 1873 988 1955 999
rect -1385 987 -559 988
rect -1385 933 -1375 987
rect -1321 933 -559 987
rect -1385 932 -559 933
rect -503 932 253 988
rect 309 932 1067 988
rect 1123 932 1886 988
rect 1942 932 1955 988
rect -1385 921 -1314 932
rect -564 917 -499 932
rect 244 922 319 932
rect 1063 920 1127 932
rect 1873 923 1955 932
rect 1671 678 1743 689
rect 1671 677 2476 678
rect 1671 623 1683 677
rect 1737 623 2476 677
rect 1671 622 2476 623
rect 1671 611 1743 622
rect 2140 476 2265 484
rect 2140 460 2153 476
rect -1747 404 2153 460
rect -1747 271 -1691 404
rect 2140 389 2153 404
rect 2240 460 2265 476
rect 2240 389 2317 460
rect 2140 378 2317 389
rect -1776 259 -1691 271
rect -1776 205 -1762 259
rect -1708 205 -1691 259
rect 37 321 108 332
rect 2010 321 2078 331
rect 37 320 2012 321
rect 37 266 49 320
rect 103 266 2012 320
rect 37 265 2012 266
rect 2068 265 2078 321
rect 37 253 108 265
rect 2010 255 2078 265
rect 2261 273 2317 378
rect 2261 260 2341 273
rect -1776 198 -1691 205
rect 2261 204 2278 260
rect 2334 204 2343 260
rect -1776 193 -1695 198
rect 2261 187 2341 204
rect 2268 185 2341 187
rect -907 90 1713 146
rect -1568 -16 -1494 -7
rect -1158 -16 -1085 -4
rect -907 -16 -851 90
rect -92 14 -22 16
rect 575 14 651 18
rect 1657 15 1713 90
rect -92 13 583 14
rect -1568 -72 -1559 -16
rect -1503 -72 -1150 -16
rect -1094 -72 -851 -16
rect -625 -25 -545 -9
rect -625 -26 -350 -25
rect -1568 -81 -1494 -72
rect -1158 -81 -1085 -72
rect -625 -80 -615 -26
rect -561 -80 -350 -26
rect -92 -41 -80 13
rect -26 -41 583 13
rect -92 -42 583 -41
rect 639 -42 651 14
rect 1647 10 1725 15
rect 2059 10 2132 23
rect 1099 -41 1180 -32
rect -92 -55 -22 -42
rect 575 -55 651 -42
rect -625 -81 -350 -80
rect -625 -94 -545 -81
rect -406 -128 -350 -81
rect 837 -97 1115 -41
rect 1171 -97 1180 -41
rect 1647 -46 1657 10
rect 1713 -46 2067 10
rect 2123 -46 2132 10
rect 1647 -55 1725 -46
rect 2059 -58 2132 -46
rect 837 -128 893 -97
rect 1099 -106 1180 -97
rect -406 -184 893 -128
rect -300 -270 -216 -258
rect 785 -270 858 -258
rect -300 -271 789 -270
rect -300 -325 -284 -271
rect -230 -325 789 -271
rect -300 -326 789 -325
rect 845 -326 858 -270
rect -300 -342 -216 -326
rect 785 -339 858 -326
rect 1325 -382 1409 -372
rect -827 -412 -753 -404
rect -827 -466 -819 -412
rect -765 -417 -753 -412
rect 1325 -417 1341 -382
rect -765 -438 1341 -417
rect 1397 -417 1409 -382
rect 2273 -417 2345 -407
rect 1397 -438 2283 -417
rect -765 -466 2283 -438
rect -827 -473 2283 -466
rect 2339 -473 2345 -417
rect -827 -481 -753 -473
rect 2273 -486 2345 -473
rect 2420 -605 2476 622
rect 2566 327 2622 1128
rect 3578 1116 3649 1128
rect 3772 1184 3850 1186
rect 3772 1130 3784 1184
rect 3838 1130 3850 1184
rect 3772 1118 3850 1130
rect 3576 1027 3651 1044
rect 4259 1027 4337 1036
rect 3576 966 3588 1027
rect 3649 1026 4337 1027
rect 3649 967 4270 1026
rect 4329 967 4337 1026
rect 3649 966 4337 967
rect 3576 958 3719 966
rect 3458 796 3554 805
rect 3458 723 3471 796
rect 3544 723 3554 796
rect 3458 711 3554 723
rect 3658 672 3719 958
rect 4259 956 4337 966
rect 4479 878 4535 1499
rect 5013 1391 5093 1403
rect 5013 1337 5023 1391
rect 5077 1389 5093 1391
rect 5923 1389 6003 1398
rect 5077 1337 5932 1389
rect 5013 1333 5932 1337
rect 5988 1333 6003 1389
rect 5013 1326 5093 1333
rect 5923 1325 6003 1333
rect 3884 823 3982 835
rect 3884 754 3900 823
rect 3969 754 3982 823
rect 3884 743 3982 754
rect 4479 822 4963 878
rect 3925 672 3999 684
rect 2962 645 3038 659
rect 2962 589 2971 645
rect 3027 589 3038 645
rect 3658 611 3928 672
rect 3989 611 3999 672
rect 3925 598 3999 611
rect 2962 574 3038 589
rect 3512 539 3588 552
rect 4332 539 4408 548
rect 4479 539 4535 822
rect 4907 811 4963 822
rect 5036 822 5107 835
rect 5036 811 5039 822
rect 4907 755 5039 811
rect 5036 744 5039 755
rect 5102 811 5107 822
rect 5873 811 5941 824
rect 5102 755 5876 811
rect 5932 755 5941 811
rect 5102 744 5107 755
rect 5036 732 5107 744
rect 5873 742 5941 755
rect 4675 708 4772 717
rect 4675 629 4686 708
rect 4759 629 4772 708
rect 4675 619 4772 629
rect 5461 656 5540 666
rect 5461 600 5471 656
rect 5527 600 5540 656
rect 5461 592 5540 600
rect 3512 538 4342 539
rect 3512 484 3528 538
rect 3582 484 4342 538
rect 3512 483 4342 484
rect 4398 483 4535 539
rect 5265 499 5345 508
rect 3512 476 3588 483
rect 4332 472 4408 483
rect 5265 443 5278 499
rect 5334 443 5345 499
rect 5265 441 5345 443
rect 5265 394 5334 441
rect 2715 338 5334 394
rect 2561 321 2632 327
rect 2561 265 2566 321
rect 2622 265 2632 321
rect 2561 254 2632 265
rect 2715 -401 2771 338
rect 4958 237 5034 250
rect 3350 205 3444 217
rect 3350 135 3362 205
rect 3432 135 3444 205
rect 3350 122 3444 135
rect 4795 181 4969 237
rect 5025 181 5034 237
rect 4417 97 4492 118
rect 4216 36 4421 97
rect 4482 36 4492 97
rect 3147 -49 3228 -36
rect 3147 -105 3160 -49
rect 3216 -105 3228 -49
rect 3553 -62 3637 -56
rect 3966 -60 4045 -50
rect 3553 -68 3905 -62
rect 3553 -71 3568 -68
rect 3147 -117 3228 -105
rect 3308 -124 3568 -71
rect 3624 -123 3905 -68
rect 3624 -124 3637 -123
rect 3308 -127 3637 -124
rect 3154 -235 3220 -223
rect 3308 -235 3364 -127
rect 3553 -136 3637 -127
rect 3149 -291 3158 -235
rect 3214 -291 3364 -235
rect 3844 -232 3905 -123
rect 3966 -116 3977 -60
rect 4033 -116 4045 -60
rect 3966 -130 4045 -116
rect 3962 -232 4061 -220
rect 4216 -232 4277 36
rect 4417 22 4492 36
rect 3154 -303 3220 -291
rect 3844 -293 3973 -232
rect 4034 -293 4277 -232
rect 3962 -301 4061 -293
rect 2600 -417 2771 -401
rect 2600 -473 2603 -417
rect 2659 -473 2771 -417
rect 2600 -486 2669 -473
rect 1681 -661 2476 -605
rect 3558 -633 3633 -624
rect 4660 -630 4735 -618
rect 3558 -634 4035 -633
rect 1681 -798 1737 -661
rect 3558 -688 3570 -634
rect 3624 -688 4035 -634
rect 3558 -689 4035 -688
rect 4660 -686 4672 -630
rect 4728 -686 4735 -630
rect 4660 -689 4735 -686
rect 3558 -700 3633 -689
rect 2300 -720 2384 -718
rect 2300 -780 2312 -720
rect 2372 -780 2384 -720
rect 3979 -747 4035 -689
rect 3966 -758 4044 -747
rect 2300 -793 2384 -780
rect 3150 -781 3229 -770
rect 1671 -803 1750 -798
rect 1671 -859 1681 -803
rect 1737 -859 1750 -803
rect 1671 -870 1750 -859
rect -1385 -1103 -1311 -1090
rect -566 -1103 -503 -1091
rect 253 -1103 316 -1091
rect 559 -1103 627 -1092
rect 1066 -1103 1131 -1092
rect 1885 -1103 1959 -1091
rect -1385 -1104 -561 -1103
rect -1385 -1158 -1376 -1104
rect -1322 -1158 -561 -1104
rect -1385 -1159 -561 -1158
rect -505 -1159 256 -1103
rect 312 -1159 564 -1103
rect 620 -1159 1071 -1103
rect 1127 -1159 1894 -1103
rect 1950 -1159 1959 -1103
rect -1385 -1172 -1311 -1159
rect -566 -1171 -503 -1159
rect 253 -1171 316 -1159
rect 559 -1163 627 -1159
rect 1066 -1171 1131 -1159
rect 1885 -1171 1959 -1159
rect -1762 -1548 -1687 -1542
rect -1904 -1604 -1756 -1548
rect -1700 -1604 -1687 -1548
rect -1762 -1608 -1687 -1604
rect -1388 -1543 -1310 -1532
rect -564 -1543 -503 -1531
rect 252 -1543 315 -1531
rect 1066 -1543 1130 -1531
rect 1883 -1543 1950 -1531
rect -1388 -1544 -562 -1543
rect -1388 -1598 -1376 -1544
rect -1322 -1598 -562 -1544
rect -1388 -1599 -562 -1598
rect -506 -1599 255 -1543
rect 311 -1599 1071 -1543
rect 1127 -1599 1885 -1543
rect 1941 -1599 1950 -1543
rect -1388 -1611 -1310 -1599
rect -564 -1611 -503 -1599
rect 252 -1612 315 -1599
rect 1066 -1608 1130 -1599
rect 1796 -1612 1950 -1599
rect -292 -2219 -204 -2209
rect -292 -2283 -280 -2219
rect -216 -2283 -204 -2219
rect 1796 -2213 1852 -1612
rect 1937 -2014 2012 -2002
rect 2311 -2014 2373 -793
rect 3150 -837 3160 -781
rect 3216 -837 3229 -781
rect 3150 -848 3229 -837
rect 3556 -788 3636 -777
rect 3556 -844 3568 -788
rect 3624 -844 3636 -788
rect 3966 -814 3977 -758
rect 4033 -814 4044 -758
rect 3966 -824 4044 -814
rect 3556 -855 3636 -844
rect 3149 -1184 3227 -1172
rect 4672 -1174 4728 -689
rect 4795 -928 4851 181
rect 4958 172 5034 181
rect 5082 98 5164 108
rect 5082 42 5094 98
rect 5150 42 5164 98
rect 5082 34 5164 42
rect 5094 -76 5150 34
rect 5471 -76 5527 592
rect 5094 -132 5527 -76
rect 5094 -787 5150 -132
rect 5080 -794 5164 -787
rect 5080 -848 5095 -794
rect 5149 -848 5164 -794
rect 5080 -855 5164 -848
rect 4784 -930 4863 -928
rect 4784 -984 4796 -930
rect 4784 -995 4801 -984
rect 4866 -995 4879 -930
rect 3149 -1238 3161 -1184
rect 3215 -1238 3227 -1184
rect 3149 -1250 3227 -1238
rect 4661 -1175 4738 -1174
rect 4661 -1186 4739 -1175
rect 4661 -1240 4673 -1186
rect 4727 -1240 4739 -1186
rect 3160 -1341 3216 -1250
rect 4661 -1252 4739 -1240
rect 1937 -2076 1939 -2014
rect 2001 -2076 2373 -2014
rect 2600 -1397 3216 -1341
rect 3853 -1330 3943 -1319
rect 3853 -1390 3866 -1330
rect 3928 -1390 3943 -1330
rect 1937 -2093 2012 -2076
rect 2398 -2213 2466 -2203
rect 1796 -2269 2401 -2213
rect 2457 -2269 2466 -2213
rect 2398 -2281 2466 -2269
rect -292 -2287 -204 -2283
rect -2492 -2886 -2386 -2874
rect -2492 -2966 -2482 -2886
rect -2399 -2966 -2386 -2886
rect -2492 -2979 -2386 -2966
rect -2480 -3736 -2398 -2979
rect -576 -3005 -473 -2992
rect -732 -3011 -570 -3005
rect -1691 -3019 -570 -3011
rect -1691 -3051 -719 -3019
rect -1704 -3069 -719 -3051
rect -1704 -3134 -1691 -3069
rect -1626 -3076 -719 -3069
rect -1626 -3134 -1614 -3076
rect -732 -3079 -719 -3076
rect -656 -3079 -570 -3019
rect -732 -3092 -570 -3079
rect -483 -3092 -473 -3005
rect -576 -3106 -473 -3092
rect -1704 -3136 -1614 -3134
rect -1441 -3223 -1352 -3210
rect -2167 -3285 -2070 -3268
rect -2167 -3343 -2142 -3285
rect -2084 -3343 -2070 -3285
rect -1441 -3283 -1428 -3223
rect -1365 -3227 -805 -3223
rect -1365 -3283 -869 -3227
rect -1441 -3286 -869 -3283
rect -817 -3286 -805 -3227
rect -1441 -3290 -805 -3286
rect -626 -3230 -536 -3219
rect -1441 -3297 -1352 -3290
rect -626 -3298 -617 -3230
rect -549 -3298 -536 -3230
rect -626 -3313 -536 -3298
rect -2167 -3346 -2070 -3343
rect -2142 -3481 -2084 -3346
rect -730 -3477 -641 -3463
rect -730 -3481 -717 -3477
rect -2142 -3537 -717 -3481
rect -654 -3537 -641 -3477
rect -2142 -3539 -641 -3537
rect -772 -3545 -641 -3539
rect -730 -3550 -641 -3545
rect -2323 -3593 -2234 -3581
rect -2323 -3658 -2310 -3593
rect -2245 -3658 -2234 -3593
rect -2323 -3666 -2234 -3658
rect -2489 -3745 -2383 -3736
rect -2489 -3827 -2450 -3745
rect -2398 -3827 -2383 -3745
rect -2489 -3841 -2383 -3827
rect -2480 -4591 -2398 -3841
rect -2310 -4459 -2243 -3666
rect -732 -3879 -643 -3873
rect -1691 -3887 -643 -3879
rect -1691 -3919 -719 -3887
rect -1704 -3937 -719 -3919
rect -1704 -4002 -1691 -3937
rect -1626 -3944 -719 -3937
rect -1626 -4002 -1614 -3944
rect -732 -3947 -719 -3944
rect -656 -3947 -643 -3887
rect -732 -3960 -643 -3947
rect -486 -3884 -404 -3872
rect -280 -3884 -216 -2287
rect 2600 -2365 2656 -1397
rect 3853 -1411 3943 -1390
rect 4683 -1415 4739 -1252
rect 4058 -1471 4739 -1415
rect 3798 -1690 3888 -1678
rect 3706 -1758 3805 -1690
rect 3873 -1758 3888 -1690
rect 3706 -1770 3888 -1758
rect 3524 -1827 3600 -1815
rect 3524 -1883 3536 -1827
rect 3592 -1883 3601 -1827
rect 3524 -1895 3600 -1883
rect 1757 -2421 2656 -2365
rect 1757 -3050 1813 -2421
rect 2079 -2780 2155 -2752
rect 2079 -2836 2089 -2780
rect 2145 -2836 2155 -2780
rect 2079 -2849 2155 -2836
rect 3706 -2789 3774 -1770
rect 4058 -1836 4114 -1471
rect 5463 -1830 5543 -1821
rect 4044 -1845 4127 -1836
rect 4044 -1901 4058 -1845
rect 4114 -1901 4127 -1845
rect 5463 -1886 5475 -1830
rect 5531 -1886 5543 -1830
rect 5463 -1896 5543 -1886
rect 4044 -1906 4127 -1901
rect 3862 -2468 3933 -2456
rect 4058 -2468 4114 -1906
rect 4231 -2115 4325 -2106
rect 4231 -2185 4244 -2115
rect 4314 -2185 4325 -2115
rect 4231 -2194 4325 -2185
rect 3862 -2469 4114 -2468
rect 3862 -2523 3875 -2469
rect 3929 -2523 4114 -2469
rect 3862 -2524 4114 -2523
rect 3862 -2536 3933 -2524
rect 3706 -2801 3846 -2789
rect 3706 -2868 3768 -2801
rect 3834 -2868 3846 -2801
rect 3706 -2880 3846 -2868
rect 1748 -3064 1824 -3050
rect 1748 -3120 1757 -3064
rect 1813 -3120 1824 -3064
rect 1748 -3132 1824 -3120
rect 332 -3222 415 -3213
rect 332 -3279 346 -3222
rect 403 -3279 415 -3222
rect 332 -3284 415 -3279
rect 346 -3308 415 -3284
rect 346 -3365 483 -3308
rect 426 -3781 483 -3365
rect 1927 -3354 2023 -3344
rect 1927 -3411 1948 -3354
rect 2005 -3411 2023 -3354
rect 3766 -3405 3828 -2880
rect 4031 -3091 4117 -3089
rect 4031 -3145 4046 -3091
rect 4100 -3145 4117 -3091
rect 4031 -3160 4117 -3145
rect 4244 -3110 4314 -2194
rect 4419 -2462 4488 -2451
rect 5116 -2462 5187 -2450
rect 4419 -2463 5122 -2462
rect 4419 -2517 4431 -2463
rect 4485 -2517 5122 -2463
rect 4419 -2518 5122 -2517
rect 5178 -2518 5187 -2462
rect 5475 -2462 5531 -1896
rect 5663 -2462 5731 -2450
rect 5475 -2463 5731 -2462
rect 5475 -2517 5666 -2463
rect 5720 -2517 5731 -2463
rect 5475 -2518 5731 -2517
rect 4419 -2529 4488 -2518
rect 5116 -2527 5187 -2518
rect 5663 -2529 5731 -2518
rect 5751 -3097 5827 -3088
rect 4045 -3358 4101 -3160
rect 4244 -3180 5649 -3110
rect 5751 -3151 5762 -3097
rect 5816 -3151 5827 -3097
rect 5751 -3165 5827 -3151
rect 4232 -3184 4326 -3180
rect 4232 -3257 4245 -3184
rect 4313 -3257 4326 -3184
rect 4232 -3269 4326 -3257
rect 1927 -3434 2023 -3411
rect 642 -3544 727 -3534
rect 642 -3549 660 -3544
rect 716 -3548 727 -3544
rect 1160 -3548 1233 -3535
rect 642 -3605 647 -3549
rect 716 -3600 1166 -3548
rect 703 -3605 1166 -3600
rect 642 -3606 1166 -3605
rect 1224 -3606 1233 -3548
rect 642 -3618 727 -3606
rect 1160 -3619 1233 -3606
rect 544 -3781 616 -3771
rect 1365 -3781 1433 -3768
rect 1534 -3781 1591 -3780
rect -486 -3885 -216 -3884
rect -486 -3947 -475 -3885
rect -413 -3947 -216 -3885
rect -486 -3948 -216 -3947
rect 257 -3783 1368 -3781
rect 257 -3837 556 -3783
rect 610 -3837 1368 -3783
rect 257 -3838 1368 -3837
rect 1425 -3838 1722 -3781
rect -486 -3960 -404 -3948
rect -1704 -4004 -1614 -4002
rect 257 -4015 314 -3838
rect 146 -4072 314 -4015
rect -1441 -4091 -1352 -4078
rect -647 -4090 -547 -4078
rect 146 -4090 215 -4072
rect -2167 -4153 -2070 -4136
rect -2167 -4211 -2142 -4153
rect -2084 -4211 -2070 -4153
rect -1441 -4151 -1428 -4091
rect -1365 -4095 -805 -4091
rect -1365 -4151 -869 -4095
rect -1441 -4154 -869 -4151
rect -817 -4154 -805 -4095
rect -1441 -4158 -805 -4154
rect -1441 -4165 -1352 -4158
rect -647 -4159 -631 -4090
rect -562 -4159 -547 -4090
rect -647 -4171 -547 -4159
rect 133 -4097 215 -4090
rect 133 -4154 146 -4097
rect 203 -4154 215 -4097
rect 133 -4165 215 -4154
rect -2167 -4214 -2070 -4211
rect -2142 -4349 -2084 -4214
rect -730 -4345 -641 -4331
rect -730 -4349 -717 -4345
rect -2142 -4405 -717 -4349
rect -654 -4405 -641 -4345
rect -2142 -4407 -641 -4405
rect -772 -4413 -641 -4407
rect -730 -4418 -641 -4413
rect -2322 -4463 -2233 -4459
rect -2322 -4530 -2310 -4463
rect -2243 -4530 -2233 -4463
rect -2322 -4544 -2233 -4530
rect -2506 -4602 -2391 -4591
rect -2506 -4684 -2450 -4602
rect -2398 -4684 -2391 -4602
rect -2506 -4698 -2391 -4684
rect -2480 -5486 -2398 -4698
rect -2310 -5307 -2243 -4544
rect 165 -4618 250 -4599
rect 165 -4683 176 -4618
rect 241 -4683 250 -4618
rect 165 -4699 250 -4683
rect -732 -4738 -643 -4732
rect -1691 -4746 -643 -4738
rect -1691 -4778 -719 -4746
rect -1704 -4796 -719 -4778
rect -1704 -4861 -1691 -4796
rect -1626 -4803 -719 -4796
rect -1626 -4861 -1614 -4803
rect -732 -4806 -719 -4803
rect -656 -4806 -643 -4746
rect -732 -4819 -643 -4806
rect -522 -4745 -447 -4733
rect -522 -4806 -518 -4745
rect -457 -4806 -447 -4745
rect -522 -4820 -447 -4806
rect -1704 -4863 -1614 -4861
rect -1441 -4950 -1352 -4937
rect -2167 -5012 -2070 -4995
rect -2167 -5070 -2142 -5012
rect -2084 -5070 -2070 -5012
rect -1441 -5010 -1428 -4950
rect -1365 -4954 -805 -4950
rect -1365 -5010 -869 -4954
rect -1441 -5013 -869 -5010
rect -817 -5013 -805 -4954
rect -1441 -5017 -805 -5013
rect -641 -4952 -549 -4940
rect -641 -5014 -631 -4952
rect -569 -5014 -549 -4952
rect 426 -4946 483 -3838
rect 544 -3850 616 -3838
rect 1365 -3850 1433 -3838
rect 1049 -3993 1119 -3980
rect 1049 -3997 1054 -3993
rect 671 -4047 1054 -3997
rect 1108 -3997 1119 -3993
rect 1365 -3997 1432 -3984
rect 1108 -4047 1367 -3997
rect 671 -4053 1367 -4047
rect 1423 -4053 1432 -3997
rect 671 -4253 727 -4053
rect 1049 -4059 1119 -4053
rect 1365 -4067 1432 -4053
rect 592 -4265 727 -4253
rect 592 -4321 601 -4265
rect 657 -4321 727 -4265
rect 980 -4272 1049 -4258
rect 1534 -4272 1591 -3838
rect 1665 -3968 1722 -3838
rect 1665 -4025 1830 -3968
rect 1773 -4112 1830 -4025
rect 1760 -4119 1842 -4112
rect 1760 -4176 1773 -4119
rect 1830 -4176 1842 -4119
rect 1760 -4183 1842 -4176
rect 1773 -4185 1830 -4183
rect 592 -4333 671 -4321
rect 979 -4329 988 -4272
rect 1045 -4329 1591 -4272
rect 980 -4345 1049 -4329
rect 1356 -4580 1427 -4569
rect 962 -4581 1833 -4580
rect 962 -4635 1368 -4581
rect 1422 -4635 1833 -4581
rect 962 -4636 1833 -4635
rect 962 -4774 1018 -4636
rect 1356 -4647 1427 -4636
rect 950 -4779 1030 -4774
rect 950 -4835 962 -4779
rect 1018 -4835 1030 -4779
rect 1777 -4792 1833 -4636
rect 950 -4845 1030 -4835
rect 1764 -4795 1846 -4792
rect 1764 -4851 1777 -4795
rect 1833 -4851 1846 -4795
rect 1764 -4860 1846 -4851
rect 647 -4946 716 -4934
rect 426 -5003 652 -4946
rect 709 -5003 718 -4946
rect 1569 -4983 1638 -4977
rect 1569 -4987 1653 -4983
rect 1948 -4987 2005 -3434
rect 3580 -3438 3828 -3405
rect 4029 -3368 4115 -3358
rect 4029 -3424 4045 -3368
rect 4101 -3424 4115 -3368
rect 4029 -3429 4115 -3424
rect 5064 -3385 5147 -3376
rect 4045 -3433 4101 -3429
rect 3554 -3440 3828 -3438
rect 3554 -3500 3568 -3440
rect 3654 -3467 3828 -3440
rect 5064 -3441 5078 -3385
rect 5134 -3441 5147 -3385
rect 5064 -3443 5147 -3441
rect 3654 -3500 3668 -3467
rect 4334 -3486 4390 -3485
rect 3554 -3512 3668 -3500
rect 4314 -3494 4401 -3486
rect 4314 -3499 4334 -3494
rect 4390 -3498 4401 -3494
rect 4730 -3498 4804 -3486
rect 3580 -4476 3642 -3512
rect 4314 -3553 4326 -3499
rect 4390 -3550 4738 -3498
rect 4380 -3553 4738 -3550
rect 4314 -3554 4738 -3553
rect 4794 -3554 4804 -3498
rect 4314 -3558 4401 -3554
rect 4314 -3563 4392 -3558
rect 4730 -3567 4804 -3554
rect 4110 -3813 4187 -3805
rect 4928 -3813 5009 -3804
rect 4110 -3814 4941 -3813
rect 4110 -3868 4122 -3814
rect 4176 -3868 4941 -3814
rect 4110 -3869 4941 -3868
rect 4997 -3869 5009 -3813
rect 4110 -3880 4187 -3869
rect 4529 -3940 4585 -3869
rect 4928 -3878 5009 -3869
rect 4517 -3949 4599 -3940
rect 4517 -4003 4530 -3949
rect 4584 -4003 4599 -3949
rect 4517 -4007 4599 -4003
rect 5078 -4157 5134 -3443
rect 5579 -3806 5649 -3180
rect 5557 -3816 5662 -3806
rect 5557 -3891 5566 -3816
rect 5652 -3891 5662 -3816
rect 5557 -3903 5662 -3891
rect 4925 -4167 5134 -4157
rect 4113 -4188 4187 -4176
rect 4113 -4244 4122 -4188
rect 4178 -4244 4293 -4188
rect 4925 -4223 4938 -4167
rect 4994 -4213 5134 -4167
rect 4994 -4223 5006 -4213
rect 4925 -4227 5006 -4223
rect 4113 -4255 4293 -4244
rect 4237 -4397 4293 -4255
rect 4933 -4397 4989 -4227
rect 4237 -4453 5263 -4397
rect 3456 -4489 3642 -4476
rect 3456 -4543 3468 -4489
rect 3545 -4543 3642 -4489
rect 3456 -4548 3642 -4543
rect 1569 -4989 2005 -4987
rect 647 -5013 716 -5003
rect -1441 -5024 -1352 -5017
rect -641 -5025 -549 -5014
rect 1569 -5043 1572 -4989
rect 1626 -4996 2005 -4989
rect 1569 -5055 1580 -5043
rect -2167 -5073 -2070 -5070
rect 1573 -5060 1580 -5055
rect 1644 -5044 2005 -4996
rect 1644 -5060 1653 -5044
rect 1573 -5071 1653 -5060
rect -2142 -5208 -2084 -5073
rect -730 -5204 -641 -5190
rect -730 -5208 -717 -5204
rect -2142 -5264 -717 -5208
rect -654 -5264 -641 -5204
rect -2142 -5266 -641 -5264
rect -772 -5272 -641 -5266
rect -730 -5277 -641 -5272
rect -2326 -5313 -2231 -5307
rect -2326 -5380 -2310 -5313
rect -2243 -5380 -2231 -5313
rect -2326 -5391 -2231 -5380
rect -558 -5332 -477 -5322
rect 3349 -5332 3426 -5323
rect -2493 -5492 -2386 -5486
rect -2493 -5574 -2450 -5492
rect -2398 -5574 -2386 -5492
rect -2493 -5593 -2386 -5574
rect -2310 -6180 -2243 -5391
rect -558 -5392 -548 -5332
rect -488 -5392 3355 -5332
rect 3415 -5392 3426 -5332
rect -558 -5402 -477 -5392
rect 3349 -5402 3426 -5392
rect 3357 -5471 3436 -5459
rect -638 -5536 3361 -5471
rect 3426 -5536 3436 -5471
rect -638 -5600 -573 -5536
rect 3357 -5548 3436 -5536
rect -732 -5606 -573 -5600
rect 585 -5606 667 -5596
rect 886 -5606 975 -5600
rect 2495 -5606 2584 -5600
rect -1691 -5614 -573 -5606
rect -1691 -5646 -719 -5614
rect -1704 -5664 -719 -5646
rect -1704 -5729 -1691 -5664
rect -1626 -5671 -719 -5664
rect -1626 -5729 -1614 -5671
rect -732 -5674 -719 -5671
rect -656 -5671 -573 -5614
rect -73 -5646 595 -5606
rect -86 -5664 595 -5646
rect -656 -5674 -643 -5671
rect -732 -5687 -643 -5674
rect -1704 -5731 -1614 -5729
rect -86 -5729 -73 -5664
rect -8 -5671 595 -5664
rect 660 -5614 975 -5606
rect 660 -5671 899 -5614
rect -8 -5729 4 -5671
rect 585 -5682 667 -5671
rect 886 -5674 899 -5671
rect 962 -5674 975 -5614
rect 1536 -5646 2503 -5606
rect 2568 -5614 2584 -5606
rect 886 -5687 975 -5674
rect 1523 -5664 2503 -5646
rect -86 -5731 4 -5729
rect 1523 -5729 1536 -5664
rect 1601 -5671 2503 -5664
rect 1601 -5729 1613 -5671
rect 2495 -5674 2508 -5671
rect 2571 -5674 2584 -5614
rect 2495 -5687 2584 -5674
rect 1523 -5731 1613 -5729
rect -1441 -5818 -1352 -5805
rect -809 -5818 -682 -5814
rect -2167 -5880 -2070 -5863
rect -2167 -5938 -2142 -5880
rect -2084 -5938 -2070 -5880
rect -1441 -5878 -1428 -5818
rect -1365 -5822 -682 -5818
rect -1365 -5878 -869 -5822
rect -1441 -5881 -869 -5878
rect -817 -5826 -682 -5822
rect -817 -5881 -750 -5826
rect -1441 -5882 -750 -5881
rect -694 -5882 -682 -5826
rect 177 -5818 266 -5805
rect 1786 -5818 1875 -5805
rect -1441 -5885 -682 -5882
rect -1441 -5892 -1352 -5885
rect -809 -5893 -682 -5885
rect -549 -5880 -452 -5863
rect -2167 -5941 -2070 -5938
rect -549 -5938 -524 -5880
rect -466 -5938 -452 -5880
rect 177 -5878 190 -5818
rect 253 -5878 573 -5818
rect 177 -5885 573 -5878
rect 640 -5822 813 -5818
rect 640 -5881 749 -5822
rect 801 -5881 813 -5822
rect 640 -5885 813 -5881
rect 1060 -5880 1157 -5863
rect 177 -5892 266 -5885
rect -549 -5941 -452 -5938
rect 1060 -5938 1085 -5880
rect 1143 -5938 1157 -5880
rect 1786 -5878 1799 -5818
rect 1862 -5822 2422 -5818
rect 1862 -5878 2358 -5822
rect 1786 -5881 2358 -5878
rect 2410 -5872 2422 -5822
rect 3580 -5872 3642 -4548
rect 4120 -4858 4193 -4854
rect 4013 -4914 4124 -4858
rect 4180 -4914 4193 -4858
rect 4013 -4919 4193 -4914
rect 4311 -4863 4391 -4855
rect 4311 -4917 4324 -4863
rect 4378 -4917 4391 -4863
rect 3706 -5561 3781 -5553
rect 4013 -5561 4069 -4919
rect 4311 -4920 4391 -4917
rect 5207 -4865 5263 -4453
rect 5333 -4864 5412 -4849
rect 5333 -4865 5345 -4864
rect 5207 -4918 5345 -4865
rect 5399 -4918 5412 -4864
rect 3706 -5562 4069 -5561
rect 3706 -5616 3716 -5562
rect 3770 -5616 4069 -5562
rect 4323 -5569 4379 -4920
rect 5207 -4921 5412 -4918
rect 5333 -4929 5412 -4921
rect 5576 -5185 5645 -3903
rect 5761 -4153 5817 -3165
rect 5754 -4162 5825 -4153
rect 5752 -4218 5761 -4162
rect 5817 -4218 5826 -4162
rect 5754 -4228 5825 -4218
rect 5559 -5200 5662 -5185
rect 5559 -5267 5568 -5200
rect 5652 -5267 5662 -5200
rect 5559 -5279 5662 -5267
rect 4924 -5558 5113 -5555
rect 3706 -5617 4069 -5616
rect 4310 -5572 4388 -5569
rect 3706 -5626 3781 -5617
rect 4310 -5628 4323 -5572
rect 4379 -5574 4388 -5572
rect 4728 -5574 4800 -5563
rect 4379 -5628 4734 -5574
rect 4310 -5630 4734 -5628
rect 4790 -5630 4800 -5574
rect 4924 -5612 4937 -5558
rect 4991 -5612 5113 -5558
rect 4924 -5617 5112 -5612
rect 4310 -5637 4388 -5630
rect 4728 -5641 4800 -5630
rect 2410 -5881 3642 -5872
rect 1786 -5882 3642 -5881
rect 1786 -5885 3469 -5882
rect 1786 -5892 1875 -5885
rect 1060 -5941 1157 -5938
rect -2142 -6076 -2084 -5941
rect -730 -6072 -641 -6058
rect -730 -6076 -717 -6072
rect -2142 -6132 -717 -6076
rect -654 -6132 -641 -6072
rect -2142 -6134 -641 -6132
rect -524 -6076 -466 -5941
rect 888 -6072 977 -6058
rect 888 -6076 901 -6072
rect -524 -6132 901 -6076
rect 964 -6132 977 -6072
rect -524 -6134 977 -6132
rect 1085 -6076 1143 -5941
rect 2349 -5944 3469 -5885
rect 3531 -5944 3642 -5882
rect 4519 -5823 4597 -5818
rect 4519 -5877 4531 -5823
rect 4585 -5877 4597 -5823
rect 4519 -5885 4597 -5877
rect 3457 -5949 3539 -5944
rect 4109 -5952 4189 -5943
rect 4530 -5952 4586 -5885
rect 4926 -5952 4996 -5941
rect 4109 -6008 4121 -5952
rect 4177 -5953 4996 -5952
rect 4177 -6007 4938 -5953
rect 4992 -6007 4996 -5953
rect 4177 -6008 4996 -6007
rect 4109 -6018 4189 -6008
rect 4926 -6019 4996 -6008
rect 2497 -6072 2586 -6058
rect 2497 -6076 2510 -6072
rect 1085 -6132 2510 -6076
rect 2573 -6132 2586 -6072
rect 1085 -6134 2586 -6132
rect -772 -6140 -641 -6134
rect 846 -6140 977 -6134
rect 2455 -6140 2586 -6134
rect -730 -6145 -641 -6140
rect 888 -6145 977 -6140
rect 2497 -6145 2586 -6140
rect -2323 -6186 -2232 -6180
rect -2323 -6253 -2310 -6186
rect -2243 -6253 -2232 -6186
rect -2323 -6264 -2232 -6253
rect 5056 -6366 5112 -5617
rect 5576 -6263 5645 -5279
rect 5573 -6273 5666 -6263
rect 5573 -6277 5589 -6273
rect 4922 -6375 5112 -6366
rect 4922 -6431 4936 -6375
rect 4992 -6431 5112 -6375
rect 5561 -6294 5589 -6277
rect 5654 -6277 5666 -6273
rect 5561 -6363 5576 -6294
rect 5654 -6338 5676 -6277
rect 5645 -6363 5676 -6338
rect 5561 -6381 5676 -6363
rect 4922 -6441 5112 -6431
<< via2 >>
rect 3538 1700 3625 1787
rect 3759 1693 3825 1759
rect 5034 1582 5095 1643
rect 5581 1574 5643 1636
rect 2153 389 2240 476
rect 2012 265 2068 321
rect 583 -42 639 14
rect 2283 -473 2339 -417
rect 3471 723 3544 796
rect 3900 754 3969 823
rect 2971 589 3027 645
rect 4686 629 4687 708
rect 4687 629 4758 708
rect 4758 629 4759 708
rect 2566 265 2622 321
rect 3362 135 3432 205
rect 3160 -105 3216 -49
rect 3568 -124 3624 -68
rect 3977 -116 4033 -60
rect 2603 -473 2659 -417
rect 564 -1159 620 -1103
rect -280 -2283 -216 -2219
rect 3160 -782 3216 -781
rect 3160 -836 3161 -782
rect 3161 -836 3215 -782
rect 3215 -836 3216 -782
rect 3160 -837 3216 -836
rect 3568 -789 3624 -788
rect 3568 -843 3569 -789
rect 3569 -843 3623 -789
rect 3623 -843 3624 -789
rect 3568 -844 3624 -843
rect 3977 -759 4033 -758
rect 3977 -813 3978 -759
rect 3978 -813 4032 -759
rect 4032 -813 4033 -759
rect 3977 -814 4033 -813
rect 4801 -984 4850 -930
rect 4850 -984 4866 -930
rect 4801 -995 4866 -984
rect 3866 -1390 3868 -1330
rect 3868 -1390 3928 -1330
rect 2401 -2269 2457 -2213
rect -570 -3006 -483 -3005
rect -570 -3091 -569 -3006
rect -569 -3091 -484 -3006
rect -484 -3091 -483 -3006
rect -570 -3092 -483 -3091
rect -617 -3298 -549 -3230
rect 3536 -1883 3592 -1827
rect 2089 -2836 2145 -2780
rect 660 -3549 716 -3544
rect 660 -3600 703 -3549
rect 703 -3600 716 -3549
rect -631 -4091 -562 -4090
rect -631 -4158 -630 -4091
rect -630 -4158 -563 -4091
rect -563 -4158 -562 -4091
rect -631 -4159 -562 -4158
rect 176 -4683 241 -4618
rect -518 -4746 -457 -4745
rect -518 -4805 -517 -4746
rect -517 -4805 -458 -4746
rect -458 -4805 -457 -4746
rect -518 -4806 -457 -4805
rect -631 -4953 -569 -4952
rect -631 -5013 -630 -4953
rect -630 -5013 -570 -4953
rect -570 -5013 -569 -4953
rect -631 -5014 -569 -5013
rect 4334 -3499 4390 -3494
rect 4334 -3550 4380 -3499
rect 4380 -3550 4390 -3499
rect 1580 -5043 1626 -4996
rect 1626 -5043 1644 -4996
rect 1580 -5060 1644 -5043
rect -548 -5392 -488 -5332
rect 3355 -5392 3415 -5332
rect 3361 -5536 3426 -5471
rect 595 -5671 660 -5606
rect 2503 -5614 2568 -5606
rect 2503 -5671 2508 -5614
rect 2508 -5671 2568 -5614
rect -750 -5827 -694 -5826
rect -750 -5881 -749 -5827
rect -749 -5881 -695 -5827
rect -695 -5881 -694 -5827
rect -750 -5882 -694 -5881
rect 573 -5885 640 -5818
rect 5589 -6294 5654 -6273
rect 5589 -6338 5645 -6294
rect 5645 -6338 5654 -6294
<< metal3 >>
rect -2254 2106 5643 2168
rect -2254 -5044 -2192 2106
rect -2129 1944 5095 2005
rect -2129 -4745 -2068 1944
rect 3524 1787 3636 1799
rect -1137 1700 3538 1787
rect 3625 1700 3636 1787
rect -1137 -3000 -1050 1700
rect 3524 1688 3636 1700
rect 3746 1759 3837 1769
rect 3746 1693 3759 1759
rect 3825 1693 3837 1759
rect 3746 1686 3837 1693
rect 3756 1562 3824 1686
rect 5034 1651 5095 1944
rect 5010 1643 5104 1651
rect 5581 1644 5643 2106
rect 5010 1582 5034 1643
rect 5095 1582 5104 1643
rect 5010 1569 5104 1582
rect 5564 1636 5656 1644
rect 5564 1574 5581 1636
rect 5643 1574 5656 1636
rect -891 1494 3824 1562
rect 5564 1559 5656 1574
rect -891 -2815 -823 1494
rect -509 973 3969 1042
rect -509 -2456 -440 973
rect 3900 835 3969 973
rect 3884 823 3982 835
rect -280 796 3554 819
rect -280 754 3471 796
rect -280 -2209 -215 754
rect 3458 723 3471 754
rect 3544 723 3554 796
rect 3884 754 3900 823
rect 3969 754 3982 823
rect 3884 743 3982 754
rect 3458 711 3554 723
rect 3468 685 3554 711
rect 4675 708 4772 717
rect 4675 685 4686 708
rect 2962 645 3038 659
rect 583 589 2971 645
rect 3027 589 3038 645
rect 3468 629 4686 685
rect 4759 629 4772 708
rect 3468 619 4772 629
rect 3468 612 4686 619
rect 583 25 639 589
rect 2962 574 3038 589
rect 2153 484 2240 485
rect 2140 476 2265 484
rect 2140 389 2153 476
rect 2240 471 2265 476
rect 2240 401 3432 471
rect 2240 389 2265 401
rect 2140 378 2265 389
rect 2010 321 2078 331
rect 2561 321 2632 327
rect 2010 265 2012 321
rect 2068 265 2566 321
rect 2622 265 2632 321
rect 2010 255 2078 265
rect 2561 254 2632 265
rect 3362 217 3432 401
rect 3350 205 3444 217
rect 3350 135 3362 205
rect 3432 135 3444 205
rect 3350 122 3444 135
rect 574 14 652 25
rect 574 -42 583 14
rect 639 -42 652 14
rect 574 -54 652 -42
rect 3147 -49 3228 -36
rect 574 -55 651 -54
rect 3147 -105 3160 -49
rect 3216 -105 3228 -49
rect 3147 -117 3228 -105
rect 3553 -68 3637 -56
rect 2273 -417 2345 -407
rect 2600 -417 2669 -401
rect 2273 -473 2283 -417
rect 2339 -473 2603 -417
rect 2659 -473 2669 -417
rect 2273 -486 2345 -473
rect 2600 -486 2669 -473
rect 3160 -770 3216 -117
rect 3553 -124 3568 -68
rect 3624 -124 3637 -68
rect 3553 -136 3637 -124
rect 3966 -60 4045 -50
rect 3966 -116 3977 -60
rect 4033 -116 4045 -60
rect 3966 -130 4045 -116
rect 3150 -781 3229 -770
rect 3568 -777 3624 -136
rect 3977 -747 4033 -130
rect 3966 -758 4044 -747
rect 3150 -837 3160 -781
rect 3216 -837 3229 -781
rect 3150 -848 3229 -837
rect 3556 -788 3636 -777
rect 3556 -844 3568 -788
rect 3624 -844 3636 -788
rect 3966 -814 3977 -758
rect 4033 -814 4044 -758
rect 3966 -824 4044 -814
rect 3556 -855 3636 -844
rect 559 -1103 627 -1092
rect 559 -1159 564 -1103
rect 620 -1159 627 -1103
rect 3568 -1110 3624 -855
rect 559 -1163 627 -1159
rect -292 -2219 -204 -2209
rect -292 -2283 -280 -2219
rect -216 -2283 -204 -2219
rect -292 -2287 -204 -2283
rect -509 -2525 -198 -2456
rect -891 -2883 -347 -2815
rect -576 -3000 -473 -2992
rect -1137 -3005 -473 -3000
rect -1137 -3087 -570 -3005
rect -576 -3092 -570 -3087
rect -483 -3092 -473 -3005
rect -576 -3106 -473 -3092
rect -626 -3230 -536 -3219
rect -415 -3230 -347 -2883
rect -626 -3298 -617 -3230
rect -549 -3298 -347 -3230
rect -626 -3313 -536 -3298
rect -267 -3596 -198 -2525
rect -631 -3665 -198 -3596
rect 564 -3534 620 -1163
rect 2089 -1166 3624 -1110
rect 4801 -930 4867 -920
rect 4866 -995 4867 -930
rect 2089 -2752 2145 -1166
rect 3536 -1815 3592 -1166
rect 4801 -1274 4866 -995
rect 3853 -1330 3943 -1319
rect 3853 -1390 3866 -1330
rect 3928 -1390 4550 -1330
rect 3853 -1411 3943 -1390
rect 3524 -1827 3600 -1815
rect 3524 -1883 3536 -1827
rect 3592 -1883 3600 -1827
rect 3524 -1895 3600 -1883
rect 2398 -2213 2466 -2203
rect 2398 -2269 2401 -2213
rect 2457 -2269 3107 -2213
rect 2398 -2281 2466 -2269
rect 2079 -2780 2155 -2752
rect 2079 -2836 2089 -2780
rect 2145 -2836 2155 -2780
rect 2079 -2849 2155 -2836
rect 3051 -3494 3107 -2269
rect 4317 -3494 4401 -3486
rect 564 -3544 727 -3534
rect 564 -3600 660 -3544
rect 716 -3600 727 -3544
rect 3051 -3550 4334 -3494
rect 4390 -3550 4401 -3494
rect 4317 -3558 4401 -3550
rect 643 -3616 727 -3600
rect -631 -4078 -562 -3665
rect -647 -4090 -547 -4078
rect -647 -4159 -631 -4090
rect -562 -4159 -547 -4090
rect -647 -4171 -547 -4159
rect 165 -4618 250 -4599
rect 165 -4683 176 -4618
rect 241 -4683 250 -4618
rect 165 -4699 250 -4683
rect -522 -4745 -447 -4733
rect -2129 -4806 -518 -4745
rect -457 -4806 -447 -4745
rect -522 -4820 -447 -4806
rect -641 -4952 -549 -4940
rect -641 -4963 -631 -4952
rect -642 -5014 -631 -4963
rect -569 -5014 -549 -4952
rect -642 -5044 -549 -5014
rect -2254 -5106 -549 -5044
rect -558 -5332 -477 -5322
rect -750 -5392 -548 -5332
rect -488 -5392 -477 -5332
rect -750 -5814 -694 -5392
rect -558 -5402 -477 -5392
rect -761 -5826 -682 -5814
rect -761 -5882 -750 -5826
rect -694 -5882 -682 -5826
rect -761 -5893 -682 -5882
rect 174 -5818 241 -4699
rect 1573 -4996 1653 -4983
rect 1573 -5000 1580 -4996
rect 595 -5060 1580 -5000
rect 1644 -5060 1653 -4996
rect 595 -5065 1653 -5060
rect 595 -5596 660 -5065
rect 1573 -5071 1653 -5065
rect 3349 -5332 3426 -5323
rect 4490 -5332 4550 -1390
rect 3349 -5392 3355 -5332
rect 3415 -5392 4550 -5332
rect 4636 -1339 4866 -1274
rect 3349 -5402 3426 -5392
rect 3357 -5471 3436 -5459
rect 4636 -5471 4701 -1339
rect 3357 -5536 3361 -5471
rect 3426 -5536 4701 -5471
rect 3357 -5548 3436 -5536
rect 585 -5606 667 -5596
rect 585 -5671 595 -5606
rect 660 -5671 667 -5606
rect 585 -5682 667 -5671
rect 2499 -5606 2581 -5592
rect 2499 -5671 2503 -5606
rect 2568 -5671 3185 -5606
rect 2499 -5682 2581 -5671
rect 568 -5818 646 -5807
rect 174 -5885 573 -5818
rect 640 -5885 646 -5818
rect 568 -5895 646 -5885
rect 3120 -6273 3185 -5671
rect 5573 -6273 5666 -6263
rect 3120 -6338 5589 -6273
rect 5654 -6338 5666 -6273
rect 5573 -6350 5666 -6338
<< labels >>
flabel metal1 -1936 -2934 -1936 -2934 0 FreeSans 480 0 0 0 VDD
port 3 nsew
flabel metal1 -2277 -3266 -2277 -3266 0 FreeSans 480 0 0 0 B1
port 4 nsew
flabel metal1 -2331 -4136 -2331 -4136 0 FreeSans 480 0 0 0 B2
port 5 nsew
flabel metal1 -2324 -5010 -2324 -5010 0 FreeSans 480 0 0 0 B3
port 6 nsew
flabel metal1 -2211 -5869 -2211 -5869 0 FreeSans 480 0 0 0 B4
port 7 nsew
flabel metal1 -590 -5894 -590 -5894 0 FreeSans 480 0 0 0 B5
port 8 nsew
flabel metal1 1006 -5871 1006 -5871 0 FreeSans 480 0 0 0 B6
port 9 nsew
flabel metal1 78 -55 78 -55 0 FreeSans 480 0 0 0 ITAIL
port 10 nsew
flabel psubdiffcont 249 -2054 249 -2054 0 FreeSans 480 0 0 0 VSS
port 13 nsew
flabel metal1 4832 2302 4832 2302 0 FreeSans 480 0 0 0 OUT-
port 14 nsew
flabel metal1 3830 2291 3830 2291 0 FreeSans 480 0 0 0 OUT+
port 15 nsew
flabel nsubdiffcont -1212 -5531 -1212 -5531 0 FreeSans 640 0 0 0 Balance_Inverter_0.VDD
flabel psubdiffcont -1204 -6214 -1204 -6214 0 FreeSans 640 0 0 0 Balance_Inverter_0.VSS
flabel via1 -697 -5635 -697 -5635 0 FreeSans 640 0 0 0 Balance_Inverter_0.OUT
flabel via1 -845 -5861 -845 -5861 0 FreeSans 640 0 0 0 Balance_Inverter_0.OUT_B
flabel via1 -2118 -5916 -2118 -5916 0 FreeSans 640 0 0 0 Balance_Inverter_0.VIN
flabel nsubdiffcont -1959 -5534 -1959 -5534 0 FreeSans 640 0 0 0 Balance_Inverter_0.Inverter_0.VDD
flabel psubdiffcont -1945 -6226 -1945 -6226 0 FreeSans 640 0 0 0 Balance_Inverter_0.Inverter_0.VSS
flabel metal1 -2121 -5865 -2121 -5865 0 FreeSans 640 0 0 0 Balance_Inverter_0.Inverter_0.IN
flabel metal1 -1754 -5892 -1754 -5892 0 FreeSans 640 0 0 0 Balance_Inverter_0.Inverter_0.OUT
flabel nsubdiffcont 406 -5531 406 -5531 0 FreeSans 640 0 0 0 Balance_Inverter_4.VDD
flabel psubdiffcont 414 -6214 414 -6214 0 FreeSans 640 0 0 0 Balance_Inverter_4.VSS
flabel via1 921 -5635 921 -5635 0 FreeSans 640 0 0 0 Balance_Inverter_4.OUT
flabel via1 773 -5861 773 -5861 0 FreeSans 640 0 0 0 Balance_Inverter_4.OUT_B
flabel via1 -500 -5916 -500 -5916 0 FreeSans 640 0 0 0 Balance_Inverter_4.VIN
flabel nsubdiffcont -341 -5534 -341 -5534 0 FreeSans 640 0 0 0 Balance_Inverter_4.Inverter_0.VDD
flabel psubdiffcont -327 -6226 -327 -6226 0 FreeSans 640 0 0 0 Balance_Inverter_4.Inverter_0.VSS
flabel metal1 -503 -5865 -503 -5865 0 FreeSans 640 0 0 0 Balance_Inverter_4.Inverter_0.IN
flabel metal1 -136 -5892 -136 -5892 0 FreeSans 640 0 0 0 Balance_Inverter_4.Inverter_0.OUT
flabel nsubdiffcont 2015 -5531 2015 -5531 0 FreeSans 640 0 0 0 Balance_Inverter_5.VDD
flabel psubdiffcont 2023 -6214 2023 -6214 0 FreeSans 640 0 0 0 Balance_Inverter_5.VSS
flabel via1 2530 -5635 2530 -5635 0 FreeSans 640 0 0 0 Balance_Inverter_5.OUT
flabel via1 2382 -5861 2382 -5861 0 FreeSans 640 0 0 0 Balance_Inverter_5.OUT_B
flabel via1 1109 -5916 1109 -5916 0 FreeSans 640 0 0 0 Balance_Inverter_5.VIN
flabel nsubdiffcont 1268 -5534 1268 -5534 0 FreeSans 640 0 0 0 Balance_Inverter_5.Inverter_0.VDD
flabel psubdiffcont 1282 -6226 1282 -6226 0 FreeSans 640 0 0 0 Balance_Inverter_5.Inverter_0.VSS
flabel metal1 1106 -5865 1106 -5865 0 FreeSans 640 0 0 0 Balance_Inverter_5.Inverter_0.IN
flabel metal1 1473 -5892 1473 -5892 0 FreeSans 640 0 0 0 Balance_Inverter_5.Inverter_0.OUT
flabel nsubdiffcont -1212 -4663 -1212 -4663 0 FreeSans 640 0 0 0 Balance_Inverter_1.VDD
flabel psubdiffcont -1204 -5346 -1204 -5346 0 FreeSans 640 0 0 0 Balance_Inverter_1.VSS
flabel via1 -697 -4767 -697 -4767 0 FreeSans 640 0 0 0 Balance_Inverter_1.OUT
flabel via1 -845 -4993 -845 -4993 0 FreeSans 640 0 0 0 Balance_Inverter_1.OUT_B
flabel via1 -2118 -5048 -2118 -5048 0 FreeSans 640 0 0 0 Balance_Inverter_1.VIN
flabel nsubdiffcont -1959 -4666 -1959 -4666 0 FreeSans 640 0 0 0 Balance_Inverter_1.Inverter_0.VDD
flabel psubdiffcont -1945 -5358 -1945 -5358 0 FreeSans 640 0 0 0 Balance_Inverter_1.Inverter_0.VSS
flabel metal1 -2121 -4997 -2121 -4997 0 FreeSans 640 0 0 0 Balance_Inverter_1.Inverter_0.IN
flabel metal1 -1754 -5024 -1754 -5024 0 FreeSans 640 0 0 0 Balance_Inverter_1.Inverter_0.OUT
flabel nsubdiffcont -1212 -3804 -1212 -3804 0 FreeSans 640 0 0 0 Balance_Inverter_2.VDD
flabel psubdiffcont -1204 -4487 -1204 -4487 0 FreeSans 640 0 0 0 Balance_Inverter_2.VSS
flabel via1 -697 -3908 -697 -3908 0 FreeSans 640 0 0 0 Balance_Inverter_2.OUT
flabel via1 -845 -4134 -845 -4134 0 FreeSans 640 0 0 0 Balance_Inverter_2.OUT_B
flabel via1 -2118 -4189 -2118 -4189 0 FreeSans 640 0 0 0 Balance_Inverter_2.VIN
flabel nsubdiffcont -1959 -3807 -1959 -3807 0 FreeSans 640 0 0 0 Balance_Inverter_2.Inverter_0.VDD
flabel psubdiffcont -1945 -4499 -1945 -4499 0 FreeSans 640 0 0 0 Balance_Inverter_2.Inverter_0.VSS
flabel metal1 -2121 -4138 -2121 -4138 0 FreeSans 640 0 0 0 Balance_Inverter_2.Inverter_0.IN
flabel metal1 -1754 -4165 -1754 -4165 0 FreeSans 640 0 0 0 Balance_Inverter_2.Inverter_0.OUT
flabel nsubdiffcont -1212 -2936 -1212 -2936 0 FreeSans 640 0 0 0 Balance_Inverter_3.VDD
flabel psubdiffcont -1204 -3619 -1204 -3619 0 FreeSans 640 0 0 0 Balance_Inverter_3.VSS
flabel via1 -697 -3040 -697 -3040 0 FreeSans 640 0 0 0 Balance_Inverter_3.OUT
flabel via1 -845 -3266 -845 -3266 0 FreeSans 640 0 0 0 Balance_Inverter_3.OUT_B
flabel via1 -2118 -3321 -2118 -3321 0 FreeSans 640 0 0 0 Balance_Inverter_3.VIN
flabel nsubdiffcont -1959 -2939 -1959 -2939 0 FreeSans 640 0 0 0 Balance_Inverter_3.Inverter_0.VDD
flabel psubdiffcont -1945 -3631 -1945 -3631 0 FreeSans 640 0 0 0 Balance_Inverter_3.Inverter_0.VSS
flabel metal1 -2121 -3270 -2121 -3270 0 FreeSans 640 0 0 0 Balance_Inverter_3.Inverter_0.IN
flabel metal1 -1754 -3297 -1754 -3297 0 FreeSans 640 0 0 0 Balance_Inverter_3.Inverter_0.OUT
<< end >>
