magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1123 -1045 1123 1045
<< metal1 >>
rect -123 39 123 45
rect -123 -39 -117 39
rect 117 -39 123 39
rect -123 -45 123 -39
<< via1 >>
rect -117 -39 117 39
<< metal2 >>
rect -123 39 123 45
rect -123 -39 -117 39
rect 117 -39 123 39
rect -123 -45 123 -39
<< end >>
