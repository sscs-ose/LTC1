* NGSPICE file created from LSBs_magic_flat.ext - technology: gf180mcuC

.subckt pex_LSBs_magic VDD VSS B1 B2 B3 B4 B5 B6 ITAIL OUT+ OUT- OUT1 OUT2 OUT3 OUT4 OUT5 OUT6 
X0 OUT+.t119 OUT+.t118 OUT+.t119 VSS.t148 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X1 Balance_Inverter_5.Inverter_0.OUT B6.t0 VDD.t4 VDD.t3 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X2 SD3_1 SDn_2.t24 VSS.t168 VSS.t154 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X3 OUT-.t90 b6.t2 OUT-.t90 VSS.t39 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X4 OUT+.t117 OUT+.t116 OUT+.t117 VSS.t147 nfet_03v3 ad=94.8f pd=0.92u as=0 ps=0 w=0.3u l=0.5u
X5 OUT6 IT.t24 SD3_1.t62 VSS.t283 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X6 OUT+.t145 b6b.t2 OUT+.t145 VSS.t89 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X7 OUT+.t115 OUT+.t114 OUT+.t115 VSS.t138 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X8 OUT+ b2.t2 OUT2.t4 VSS.t230 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X9 SD3_1 IT.t25 OUT6.t37 VSS.t254 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X10 OUT- b5b.t2 OUT5.t31 VSS.t186 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X11 VSS G2.t3 SD2_5.t11 VSS.t13 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X12 SD3_1 SDn_2.t25 VSS.t170 VSS.t169 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X13 OUT+.t113 OUT+.t112 OUT+.t113 VSS.t112 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X14 OUT+ b5.t2 OUT5.t44 VSS.t200 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X15 OUT- b4b.t2 OUT4.t21 VSS.t210 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X16 OUT6 IT.t26 SD3_1.t0 VSS.t36 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X17 OUT6 b6b.t3 OUT-.t37 VSS.t16 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X18 OUT6 b6.t3 OUT+.t12 VSS.t16 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X19 OUT+.t161 b5b.t3 OUT+.t161 VSS.t201 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X20 OUT- b2b.t2 OUT2.t1 VSS.t42 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X21 SD3_1 IT.t27 OUT6.t35 VSS.t37 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X22 OUT-.t179 OUT-.t178 OUT-.t179 VSS.t67 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X23 b1b B1.t0 VSS.t218 VSS.t217 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X24 SD2_5 ITAIL.t2 OUT4.t10 VSS.t113 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X25 OUT- b6b.t4 OUT6.t46 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X26 OUT+.t111 OUT+.t110 OUT+.t111 VSS.t144 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X27 VSS Balance_Inverter_5.Inverter_0.OUT b6.t0 VSS.t319 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X28 SDn_1 IT.t28 OUT5.t7 VSS.t38 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X29 SDn_2 SDn_2.t14 VSS.t88 VSS.t87 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X30 OUT5 b5.t3 OUT+.t142 VSS.t194 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X31 OUT+ b3.t2 OUT3.t4 VSS.t70 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X32 VSS SDn_2.t27 SD3_1.t59 VSS.t171 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X33 OUT+ b6.t4 OUT6.t91 VSS.t21 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X34 OUT-.t177 OUT-.t176 OUT-.t177 VSS.t111 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X35 b2b b2.t3 VDD.t60 VDD.t59 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X36 OUT6 IT.t29 SD3_1.t8 VSS.t130 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X37 SD3_1 IT.t30 OUT6.t33 VSS.t131 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X38 OUT- b6b.t5 OUT6.t4 VSS.t41 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X39 OUT+.t109 OUT+.t108 OUT+.t109 VSS.t146 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X40 OUT-.t175 OUT-.t174 OUT-.t175 VSS.t91 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X41 OUT-.t173 OUT-.t172 OUT-.t173 VSS.t136 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X42 OUT4 b4.t2 OUT+.t125 VSS.t182 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X43 SD3_1 IT.t31 OUT6.t32 VSS.t132 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X44 OUT-.t171 OUT-.t170 OUT-.t171 VSS.t174 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X45 SD3_1 IT.t32 OUT6.t31 VSS.t149 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X46 SD2_1 G2.t4 VSS.t236 VSS.t208 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X47 OUT6 b6.t5 OUT+.t168 VSS.t18 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X48 OUT-.t72 b4.t3 OUT-.t72 VSS.t227 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X49 OUT6 IT.t33 SD3_1.t15 VSS.t150 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X50 SDn_2 IT.t14 IT.t15 VSS.t83 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X51 OUT- b6b.t6 OUT6.t5 VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X52 OUT-.t73 b4.t4 OUT-.t73 VSS.t287 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X53 IT G1_2.t24 SD1_1.t7 VDD.t19 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X54 OUT-.t57 b2.t4 OUT-.t57 VSS.t231 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X55 OUT- b6b.t7 OUT6.t2 VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X56 VSS G2.t5 SD2_4.t3 VSS.t73 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X57 OUT+.t107 OUT+.t106 OUT+.t107 VSS.t93 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X58 OUT6 b6.t6 OUT+.t169 VSS.t17 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X59 OUT6 IT.t34 SD3_1.t16 VSS.t151 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X60 OUT+.t105 OUT+.t104 OUT+.t105 VSS.t93 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X61 VSS SDn_2.t28 SDn_1.t31 VSS.t239 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X62 G1_1 G1_2.t12 G1_2.t13 VDD.t48 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X63 OUT-.t34 b5.t4 OUT-.t34 VSS.t199 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X64 OUT4 ITAIL.t3 SD2_5.t15 VSS.t318 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X65 OUT+.t103 OUT+.t102 OUT+.t103 VSS.t91 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X66 OUT-.t169 OUT-.t168 OUT-.t169 VSS.t91 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X67 OUT-.t167 OUT-.t166 OUT-.t167 VSS.t138 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X68 OUT6 b6b.t8 OUT-.t3 VSS.t18 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X69 OUT6 b6.t7 OUT+.t186 VSS.t18 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X70 OUT+.t178 b6b.t9 OUT+.t178 VSS.t72 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X71 SD2_1 ITAIL.t4 G1_2.t23 VSS.t119 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X72 VSS SDn_2.t29 SD3_1.t58 VSS.t242 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X73 G1_2 G1_2.t4 G1_1.t6 VDD.t17 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X74 Balance_Inverter_1.Inverter_0.OUT B3.t0 VDD.t41 VDD.t40 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X75 OUT+ b6.t8 OUT6.t87 VSS.t21 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X76 OUT+.t155 b4b.t3 OUT+.t155 VSS.t215 nfet_03v3 ad=0.16p pd=1.64u as=0 ps=0 w=0.3u l=0.5u
X77 OUT+ b4.t5 OUT4.t0 VSS.t26 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X78 OUT-.t89 b6.t9 OUT-.t89 VSS.t129 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X79 OUT+.t101 OUT+.t100 OUT+.t101 VSS.t138 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X80 OUT- b6b.t10 OUT6.t93 VSS.t41 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X81 OUT+.t99 OUT+.t98 OUT+.t99 VSS.t93 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X82 OUT5 b5b.t4 OUT-.t58 VSS.t190 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X83 VSS SDn_2.t30 SD3_1.t57 VSS.t245 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X84 G1_2 ITAIL.t5 SD2_1.t11 VSS.t108 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X85 OUT6 IT.t35 SD3_1.t11 VSS.t133 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X86 OUT-.t35 b5.t5 OUT-.t35 VSS.t196 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X87 SD1_1 G1_2.t26 IT.t17 VDD.t20 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X88 SDn_1 SDn_2.t31 VSS.t248 VSS.t38 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X89 OUT5 b5.t6 OUT+.t140 VSS.t29 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X90 VDD G1_1.t24 SD1_1.t10 VDD.t26 pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X91 SD3_1 IT.t36 OUT6.t27 VSS.t134 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X92 VSS SDn_2.t32 SDn_1.t29 VSS.t124 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X93 OUT-.t165 OUT-.t164 OUT-.t165 VSS.t80 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X94 OUT-.t163 OUT-.t162 OUT-.t163 VSS.t79 nfet_03v3 ad=94.8f pd=0.92u as=0 ps=0 w=0.3u l=0.5u
X95 OUT5 b5b.t5 OUT-.t59 VSS.t194 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X96 OUT-.t32 b5.t7 OUT-.t32 VSS.t198 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X97 OUT+ b6.t10 OUT6.t86 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X98 OUT6 IT.t37 SD3_1.t13 VSS.t135 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X99 SDn_1 IT.t38 OUT5.t6 VSS.t152 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X100 G1_2 G1_2.t2 G1_1.t5 VDD.t35 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X101 OUT+ b6.t11 OUT6.t85 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X102 OUT+.t127 b6b.t11 OUT+.t127 VSS.t90 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X103 OUT+.t97 OUT+.t96 OUT+.t97 VSS.t82 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X104 VDD b3b.t2 b3.t0 VDD.t69 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X105 VSS G2.t6 SD2_5.t10 VSS.t10 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X106 OUT6 b6b.t12 OUT-.t22 VSS.t19 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X107 VSS Balance_Inverter_0.Inverter_0.OUT b4.t0 VSS.t183 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X108 OUT+.t95 OUT+.t94 OUT+.t95 VSS.t81 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X109 OUT6 IT.t39 SD3_1.t17 VSS.t153 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X110 OUT+.t93 OUT+.t92 OUT+.t93 VSS.t111 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X111 VSS G2.t7 SD2_5.t9 VSS.t13 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X112 SD3_1 IT.t40 OUT6.t24 VSS.t154 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X113 VSS SDn_2.t33 SDn_1.t28 VSS.t251 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X114 OUT5 b5b.t6 OUT-.t60 VSS.t28 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X115 VDD G1_1.t22 G1_1.t23 VDD.t42 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X116 OUT+.t91 OUT+.t90 OUT+.t91 VSS.t111 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X117 OUT- b1b.t2 OUT1.t1 VSS.t216 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X118 SD3_1 SDn_2.t34 VSS.t255 VSS.t254 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X119 OUT6 b6b.t13 OUT-.t64 VSS.t17 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X120 OUT3 ITAIL.t6 SD2_4.t7 VSS.t107 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X121 SDn_1 IT.t41 OUT5.t5 VSS.t261 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X122 OUT-.t88 b6.t12 OUT-.t88 VSS.t72 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X123 SD3_1 IT.t42 OUT6.t23 VSS.t306 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X124 OUT-.t33 b5.t8 OUT-.t33 VSS.t195 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X125 VSS SDn_2.t35 SD3_1.t55 VSS.t36 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X126 SDn_1 IT.t43 OUT5.t4 VSS.t308 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X127 SD1_1 G1_1.t25 VDD.t30 VDD.t29 pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X128 SD3_1 SDn_2.t36 VSS.t258 VSS.t37 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X129 OUT+.t171 b3b.t3 OUT+.t171 VSS.t280 nfet_03v3 ad=94.8f pd=0.92u as=0 ps=0 w=0.3u l=0.5u
X130 OUT5 b5b.t7 OUT-.t27 VSS.t190 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X131 OUT+.t89 OUT+.t88 OUT+.t89 VSS.t109 nfet_03v3 ad=94.8f pd=0.92u as=0 ps=0 w=0.3u l=0.5u
X132 VSS SDn_2.t37 SDn_1.t27 VSS.t49 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X133 OUT5 b5.t9 OUT+.t139 VSS.t29 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X134 OUT6 b6.t13 OUT+.t26 VSS.t19 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X135 OUT6 b6b.t14 OUT-.t65 VSS.t19 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X136 SD3_1 SDn_2.t38 VSS.t53 VSS.t52 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X137 OUT+.t156 b4b.t4 OUT+.t156 VSS.t181 nfet_03v3 ad=0 pd=0 as=94.8f ps=0.92u w=0.3u l=0.5u
X138 VSS SDn_2.t39 SDn_1.t26 VSS.t54 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X139 OUT-.t87 b6.t14 OUT-.t87 VSS.t17 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X140 OUT- b5b.t8 OUT5.t26 VSS.t191 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X141 SDn_1 SDn_2.t40 VSS.t58 VSS.t57 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X142 OUT-.t6 b4.t6 OUT-.t6 VSS.t27 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X143 VSS SDn_2.t41 SD3_1.t52 VSS.t130 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X144 OUT-.t86 b6.t15 OUT-.t86 VSS.t90 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X145 OUT+.t87 OUT+.t86 OUT+.t87 VSS.t82 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X146 G1_1 G1_1.t20 VDD.t76 VDD.t75 pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X147 OUT+ b5.t10 OUT5.t40 VSS.t197 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X148 OUT+.t166 b6b.t15 OUT+.t166 VSS.t39 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X149 SD2_5 G2.t8 VSS.t207 VSS.t5 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X150 SD2_1 G2.t9 VSS.t209 VSS.t208 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X151 SDn_2 SDn_2.t12 VSS.t86 VSS.t85 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X152 OUT-.t85 b6.t16 OUT-.t85 VSS.t40 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X153 OUT-.t84 b6.t17 OUT-.t84 VSS.t89 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X154 OUT-.t161 OUT-.t160 OUT-.t161 VSS.t315 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X155 OUT5 b5b.t9 OUT-.t7 VSS.t28 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X156 VSS Balance_Inverter_2.Inverter_0.OUT b2.t1 VSS.t114 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X157 Balance_Inverter_3.Inverter_0.OUT B1.t1 VSS.t161 VSS.t160 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X158 VSS SDn_2.t43 SD3_1.t51 VSS.t122 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X159 VSS G2.t10 SD2_1.t5 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X160 SD3_1 SDn_2.t44 VSS.t292 VSS.t132 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X161 OUT-.t83 b6.t18 OUT-.t83 VSS.t187 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X162 OUT-.t159 OUT-.t158 OUT-.t159 VSS.t112 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X163 OUT5 IT.t44 SDn_1.t11 VSS.t251 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X164 OUT- b6b.t16 OUT6.t56 VSS.t21 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X165 SD2_3 G2.t11 VSS.t214 VSS.t213 nfet_03v3 ad=0.264p pd=2.08u as=0.264p ps=2.08u w=0.6u l=0.5u
X166 VSS G2.t12 SD2_4.t2 VSS.t73 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X167 OUT- b6b.t17 OUT6.t59 VSS.t21 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X168 SDn_2 SDn_2.t10 VSS.t84 VSS.t83 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X169 OUT-.t15 b3.t3 OUT-.t15 VSS.t71 nfet_03v3 ad=0.16p pd=1.64u as=0 ps=0 w=0.3u l=0.5u
X170 OUT+ b6.t19 OUT6.t83 VSS.t41 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X171 OUT4 b4b.t5 OUT-.t44 VSS.t180 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X172 OUT+ b6.t20 OUT6.t82 VSS.t41 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X173 OUT-.t157 OUT-.t156 OUT-.t157 VSS.t81 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X174 OUT6 b6b.t18 OUT-.t69 VSS.t16 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X175 OUT6 b6b.t19 OUT-.t16 VSS.t17 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X176 SDn_2 IT.t12 IT.t13 VSS.t178 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X177 OUT+.t85 OUT+.t84 OUT+.t85 VSS.t145 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X178 G2 ITAIL.t0 ITAIL.t1 VSS.t45 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X179 OUT4 ITAIL.t7 SD2_5.t14 VSS.t318 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X180 VSS SDn_2.t46 SD3_1.t49 VSS.t151 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X181 VDD b1b.t3 b1.t1 VDD.t54 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X182 OUT+.t158 b4b.t6 OUT+.t158 VSS.t35 nfet_03v3 ad=0.16p pd=1.64u as=0 ps=0 w=0.3u l=0.5u
X183 SDn_1 SDn_2.t47 VSS.t262 VSS.t261 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X184 SD1_1 G1_2.t28 IT.t18 VDD.t36 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X185 OUT+.t159 b4b.t7 OUT+.t159 VSS.t219 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X186 b5b b5.t11 VDD.t53 VDD.t52 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X187 G1_1 G1_1.t18 VDD.t8 VDD.t7 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X188 SDn_1 IT.t45 OUT5.t3 VSS.t57 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X189 OUT+ b6.t21 OUT6.t81 VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X190 VSS G2.t13 SD2_3.t0 VSS.t76 nfet_03v3 ad=0.264p pd=2.08u as=0.264p ps=2.08u w=0.6u l=0.5u
X191 OUT+.t21 b6b.t20 OUT+.t21 VSS.t40 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X192 OUT-.t155 OUT-.t154 OUT-.t155 VSS.t93 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X193 SD2_5 ITAIL.t8 OUT4.t11 VSS.t104 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X194 G1_2 ITAIL.t9 SD2_1.t10 VSS.t108 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X195 SD3_1 SDn_2.t48 VSS.t263 VSS.t126 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X196 OUT5 b5.t12 OUT+.t138 VSS.t190 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X197 SD2_5 G2.t14 VSS.t156 VSS.t155 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X198 OUT+.t150 b6b.t21 OUT+.t150 VSS.t187 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X199 OUT5 b5b.t10 OUT-.t8 VSS.t29 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X200 VDD G1_1.t16 G1_1.t17 VDD.t10 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X201 OUT6 IT.t46 SD3_1.t20 VSS.t245 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X202 VSS SDn_2.t49 SD3_1.t47 VSS.t133 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X203 b5b B5.t0 VSS.t222 VSS.t221 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X204 OUT+.t148 b5b.t11 OUT+.t148 VSS.t202 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X205 OUT+.t160 b4b.t8 OUT+.t160 VSS.t220 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X206 SD3_1 SDn_2.t50 VSS.t266 VSS.t134 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X207 VSS SDn_2.t8 SDn_2.t9 VSS.t165 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X208 VSS G2.t15 SD2_5.t6 VSS.t10 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X209 b3b b3.t4 VDD.t14 VDD.t13 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X210 OUT+.t149 b5b.t12 OUT+.t149 VSS.t203 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X211 SD1_1 G1_1.t28 VDD.t87 VDD.t86 pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X212 OUT+.t146 b5b.t13 OUT+.t146 VSS.t29 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X213 VSS SDn_2.t6 SDn_2.t7 VSS.t162 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X214 OUT-.t153 OUT-.t152 OUT-.t153 VSS.t82 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X215 OUT-.t19 b4.t7 OUT-.t19 VSS.t117 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X216 SD3_1 SDn_2.t51 VSS.t303 VSS.t302 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X217 VDD b4b.t9 b4.t1 VDD.t83 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X218 OUT- b6b.t22 OUT6.t47 VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X219 OUT+ b6.t22 OUT6.t80 VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X220 VDD G1_1.t29 SD1_1.t15 VDD.t88 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X221 Balance_Inverter_0.Inverter_0.OUT B4.t0 VSS.t323 VSS.t322 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X222 OUT-.t151 OUT-.t150 OUT-.t151 VSS.t81 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X223 OUT4 b4.t8 OUT+.t25 VSS.t118 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X224 OUT+.t83 OUT+.t82 OUT+.t83 VSS.t93 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X225 OUT5 b5.t13 OUT+.t143 VSS.t28 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X226 OUT3 ITAIL.t10 SD2_4.t6 VSS.t107 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X227 SD1_1 G1_2.t29 IT.t19 VDD.t37 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X228 VSS SDn_2.t52 SD3_1.t44 VSS.t153 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X229 OUT-.t149 OUT-.t148 OUT-.t149 VSS.t93 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X230 OUT+.t147 b5b.t14 OUT+.t147 VSS.t201 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X231 OUT+.t81 OUT+.t80 OUT+.t81 VSS.t91 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X232 SD1_1 G1_1.t30 VDD.t39 VDD.t38 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X233 OUT6 b6.t23 OUT+.t0 VSS.t16 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X234 OUT4 b4b.t10 OUT-.t94 VSS.t182 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X235 OUT+.t14 b2b.t3 OUT+.t14 VSS.t43 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X236 OUT6 b6b.t23 OUT-.t42 VSS.t18 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X237 OUT+.t79 OUT+.t78 OUT+.t79 VSS.t144 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X238 SD3_1 SDn_2.t53 VSS.t307 VSS.t306 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X239 G1_2 ITAIL.t11 SD2_1.t9 VSS.t105 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X240 OUT- b4b.t11 OUT4.t18 VSS.t26 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X241 VDD G1_1.t14 G1_1.t15 VDD.t92 pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X242 OUT- b6b.t24 OUT6.t49 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X243 b4b B4.t1 VSS.t311 VSS.t310 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X244 SDn_1 SDn_2.t54 VSS.t309 VSS.t308 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X245 OUT+ b4.t9 OUT4.t1 VSS.t32 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X246 G1_1 G1_1.t12 VDD.t6 VDD.t5 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X247 OUT5 IT.t47 SDn_1.t9 VSS.t97 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X248 SDn_1 SDn_2.t55 VSS.t268 VSS.t125 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X249 OUT-.t14 b3.t5 OUT-.t14 VSS.t68 nfet_03v3 ad=94.8f pd=0.92u as=0 ps=0 w=0.3u l=0.5u
X250 OUT1 b1.t2 OUT+.t120 VSS.t159 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X251 OUT-.t147 OUT-.t146 OUT-.t147 VSS.t140 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X252 OUT5 IT.t48 SDn_1.t8 VSS.t124 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X253 OUT5 IT.t49 SDn_1.t7 VSS.t54 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X254 VDD b5b.t15 b5.t1 VDD.t49 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X255 OUT-.t145 OUT-.t144 OUT-.t145 VSS.t111 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X256 OUT5 IT.t50 SDn_1.t6 VSS.t128 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X257 OUT6 b6.t24 OUT+.t1 VSS.t17 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X258 OUT-.t9 b4.t10 OUT-.t9 VSS.t33 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X259 VSS SDn_2.t56 SD3_1.t42 VSS.t269 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X260 OUT- b5b.t16 OUT5.t23 VSS.t186 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X261 OUT6 b6.t25 OUT+.t189 VSS.t17 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X262 SD3_1 IT.t51 OUT6.t21 VSS.t52 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X263 SD1_1 G1_2.t30 IT.t20 VDD.t57 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X264 OUT+ b5.t14 OUT5.t47 VSS.t200 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X265 OUT+.t77 OUT+.t76 OUT+.t77 VSS.t80 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X266 SD2_5 G2.t16 VSS.t6 VSS.t5 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X267 OUT6 IT.t52 SD3_1.t7 VSS.t94 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X268 OUT-.t71 b4.t11 OUT-.t71 VSS.t267 nfet_03v3 ad=0 pd=0 as=94.8f ps=0.92u w=0.3u l=0.5u
X269 SDn_2 IT.t10 IT.t11 VSS.t85 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X270 OUT+.t75 OUT+.t74 OUT+.t75 VSS.t143 nfet_03v3 ad=0 pd=0 as=94.8f ps=0.92u w=0.3u l=0.5u
X271 OUT+.t73 OUT+.t72 OUT+.t73 VSS.t142 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X272 OUT3 b3.t6 OUT+.t16 VSS.t69 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X273 SD3_1 IT.t53 OUT6.t19 VSS.t102 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X274 VSS G2.t17 SD2_1.t4 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X275 OUT+ b6.t26 OUT6.t76 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X276 OUT- b6b.t25 OUT6.t41 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X277 Balance_Inverter_2.Inverter_0.OUT B2.t0 VSS.t226 VSS.t225 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X278 SDn_1 SDn_2.t57 VSS.t272 VSS.t152 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X279 SD2_3 ITAIL.t12 OUT2.t5 VSS.t213 nfet_03v3 ad=0.264p pd=2.08u as=0.264p ps=2.08u w=0.6u l=0.5u
X280 OUT+.t122 b6b.t26 OUT+.t122 VSS.t129 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X281 OUT+.t19 b6b.t27 OUT+.t19 VSS.t72 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X282 OUT6 IT.t54 SD3_1.t3 VSS.t122 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X283 SDn_1 IT.t55 OUT5.t2 VSS.t123 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X284 OUT-.t143 OUT-.t142 OUT-.t143 VSS.t93 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X285 OUT+.t71 OUT+.t70 OUT+.t71 VSS.t111 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X286 OUT-.t141 OUT-.t140 OUT-.t141 VSS.t111 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X287 OUT+.t20 b6b.t28 OUT+.t20 VSS.t17 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X288 IT IT.t8 SDn_2.t18 VSS.t175 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X289 SD2_2 ITAIL.t13 OUT1.t2 VSS.t45 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X290 IT IT.t6 SDn_2.t17 VSS.t162 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X291 SDn_1 IT.t58 OUT5.t1 VSS.t125 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X292 OUT-.t139 OUT-.t138 OUT-.t139 VSS.t328 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X293 Balance_Inverter_4.Inverter_0.OUT B5.t1 VSS.t224 VSS.t223 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X294 OUT4 ITAIL.t14 SD2_5.t1 VSS.t106 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X295 OUT+.t188 b3b.t4 OUT+.t188 VSS.t24 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X296 OUT6 b6.t27 OUT+.t170 VSS.t16 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X297 b2b B2.t1 VSS.t279 VSS.t278 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X298 OUT-.t36 b5.t15 OUT-.t36 VSS.t199 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X299 b1b b1.t3 VDD.t78 VDD.t77 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X300 OUT+.t163 b4b.t12 OUT+.t163 VSS.t227 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X301 SDn_1 SDn_2.t58 VSS.t274 VSS.t273 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X302 OUT-.t82 b6.t28 OUT-.t82 VSS.t39 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X303 SD3_1 SDn_2.t59 VSS.t276 VSS.t275 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X304 OUT+.t23 b6b.t29 OUT+.t23 VSS.t89 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X305 OUT-.t137 OUT-.t136 OUT-.t137 VSS.t91 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X306 OUT-.t135 OUT-.t134 OUT-.t135 VSS.t136 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X307 SDn_1 SDn_2.t60 VSS.t277 VSS.t123 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X308 OUT-.t133 OUT-.t132 OUT-.t133 VSS.t145 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X309 OUT6 b6.t29 OUT+.t2 VSS.t18 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X310 OUT6 b6.t30 OUT+.t3 VSS.t19 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X311 OUT+.t69 OUT+.t68 OUT+.t69 VSS.t80 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X312 OUT+.t67 OUT+.t66 OUT+.t67 VSS.t112 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X313 OUT- b4b.t13 OUT4.t17 VSS.t228 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X314 OUT2 ITAIL.t15 SD2_3.t2 VSS.t76 nfet_03v3 ad=0.264p pd=2.08u as=0.264p ps=2.08u w=0.6u l=0.5u
X315 OUT+.t24 b6b.t30 OUT+.t24 VSS.t90 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X316 OUT+ b6.t31 OUT6.t72 VSS.t21 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X317 OUT+.t65 OUT+.t64 OUT+.t65 VSS.t138 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X318 OUT+.t63 OUT+.t62 OUT+.t63 VSS.t81 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X319 OUT+ b5.t16 OUT5.t38 VSS.t191 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X320 SD2_5 ITAIL.t16 OUT4.t3 VSS.t104 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X321 OUT+.t61 OUT+.t60 OUT+.t61 VSS.t81 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X322 OUT- b6b.t31 OUT6.t94 VSS.t41 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X323 Balance_Inverter_3.Inverter_0.OUT B1.t2 VDD.t62 VDD.t61 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X324 OUT- b5b.t17 OUT5.t22 VSS.t197 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X325 SD2_5 G2.t18 VSS.t192 VSS.t155 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X326 VSS SDn_2.t61 SD3_1.t40 VSS.t293 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X327 SD2_4 G2.t19 VSS.t193 VSS.t62 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X328 SD3_1 IT.t59 OUT6.t17 VSS.t126 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X329 OUT-.t31 b5.t17 OUT-.t31 VSS.t198 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X330 OUT-.t81 b6.t32 OUT-.t81 VSS.t129 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X331 OUT+.t59 OUT+.t58 OUT+.t59 VSS.t141 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X332 OUT+.t57 OUT+.t56 OUT+.t57 VSS.t93 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X333 OUT-.t131 OUT-.t130 OUT-.t131 VSS.t138 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X334 OUT- b3b.t5 OUT3.t11 VSS.t23 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X335 OUT-.t129 OUT-.t128 OUT-.t129 VSS.t92 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X336 SD3_1 IT.t60 OUT6.t16 VSS.t127 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X337 VSS Balance_Inverter_4.Inverter_0.OUT b5.t0 VSS.t46 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X338 b4b b4.t12 VDD.t64 VDD.t63 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X339 OUT- b6b.t32 OUT6.t95 VSS.t21 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X340 OUT+ b6.t33 OUT6.t71 VSS.t21 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X341 OUT+ b6.t34 OUT6.t70 VSS.t41 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X342 OUT- b6b.t33 OUT6.t39 VSS.t41 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X343 OUT+.t55 OUT+.t54 OUT+.t55 VSS.t92 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X344 SD3_1 IT.t61 OUT6.t15 VSS.t302 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X345 OUT+.t175 b3b.t6 OUT+.t175 VSS.t280 nfet_03v3 ad=94.8f pd=0.92u as=0 ps=0 w=0.3u l=0.5u
X346 VSS G2.t20 SD2_1.t3 VSS.t64 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X347 SDn_2 SDn_2.t4 VSS.t179 VSS.t178 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X348 VSS SDn_2.t63 SDn_1.t18 VSS.t296 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X349 OUT-.t127 OUT-.t126 OUT-.t127 VSS.t91 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X350 OUT+.t164 b4b.t14 OUT+.t164 VSS.t229 nfet_03v3 ad=0 pd=0 as=94.8f ps=0.92u w=0.3u l=0.5u
X351 G1_2 ITAIL.t17 SD2_1.t8 VSS.t105 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X352 OUT+ b5.t18 OUT5.t39 VSS.t191 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X353 G1_1 G1_2.t10 G1_2.t11 VDD.t9 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X354 OUT6 b6.t35 OUT+.t157 VSS.t18 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X355 OUT5 b5b.t18 OUT-.t67 VSS.t194 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X356 IT G1_2.t31 SD1_1.t2 VDD.t58 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X357 OUT-.t80 b6.t36 OUT-.t80 VSS.t40 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X358 OUT4 b4b.t15 OUT-.t51 VSS.t34 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X359 OUT4 b4.t13 OUT+.t124 VSS.t180 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X360 Balance_Inverter_0.Inverter_0.OUT B4.t2 VDD.t74 VDD.t73 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X361 OUT- b5b.t19 OUT5.t20 VSS.t197 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X362 SD2_1 ITAIL.t18 G1_2.t18 VSS.t30 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X363 OUT-.t125 OUT-.t124 OUT-.t125 VSS.t174 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X364 OUT+.t53 OUT+.t52 OUT+.t53 VSS.t140 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X365 OUT+.t51 OUT+.t50 OUT+.t51 VSS.t137 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X366 SD2_1 G2.t21 VSS.t206 VSS.t0 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X367 OUT6 b6b.t34 OUT-.t18 VSS.t19 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X368 OUT-.t79 b6.t37 OUT-.t79 VSS.t187 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X369 VSS SDn_2.t64 SD3_1.t39 VSS.t299 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X370 VSS Balance_Inverter_1.Inverter_0.OUT b3.t1 VSS.t325 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X371 b6b B6.t1 VSS.t334 VSS.t333 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X372 OUT+.t15 b2b.t4 OUT+.t15 VSS.t44 nfet_03v3 ad=0 pd=0 as=94.8f ps=0.92u w=0.3u l=0.5u
X373 OUT6 b6b.t35 OUT-.t46 VSS.t16 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X374 OUT6 IT.t62 SD3_1.t28 VSS.t269 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X375 OUT6 b6b.t36 OUT-.t47 VSS.t16 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X376 G1_1 G1_2.t8 G1_2.t9 VDD.t47 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X377 OUT-.t123 OUT-.t122 OUT-.t123 VSS.t80 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X378 OUT-.t121 OUT-.t120 OUT-.t121 VSS.t110 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X379 VSS G2.t1 G2.t2 VSS.t2 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X380 VSS SDn_2.t65 SD3_1.t38 VSS.t94 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X381 VSS SDn_2.t66 SDn_1.t17 VSS.t97 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X382 SD3_1 SDn_2.t67 VSS.t101 VSS.t100 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X383 OUT-.t21 b4.t14 OUT-.t21 VSS.t181 nfet_03v3 ad=0 pd=0 as=94.8f ps=0.92u w=0.3u l=0.5u
X384 OUT-.t96 b3.t7 OUT-.t96 VSS.t71 nfet_03v3 ad=0.16p pd=1.64u as=0 ps=0 w=0.3u l=0.5u
X385 SD3_1 SDn_2.t68 VSS.t103 VSS.t102 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X386 SD2_4 ITAIL.t19 OUT3.t7 VSS.t31 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X387 OUT- b6b.t37 OUT6.t52 VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X388 OUT3 b3b.t7 OUT-.t74 VSS.t314 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X389 IT G1_2.t32 SD1_1.t1 VDD.t91 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X390 OUT+.t49 OUT+.t48 OUT+.t49 VSS.t93 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X391 Balance_Inverter_5.Inverter_0.OUT B6.t2 VSS.t317 VSS.t316 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X392 OUT4 ITAIL.t20 SD2_5.t2 VSS.t106 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X393 OUT6 b6b.t38 OUT-.t49 VSS.t17 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X394 OUT3 b3.t8 OUT+.t179 VSS.t69 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X395 OUT+.t123 b1b.t4 OUT+.t123 VSS.t43 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X396 OUT-.t30 b5.t19 OUT-.t30 VSS.t196 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X397 SD3_1 IT.t63 OUT6.t13 VSS.t275 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X398 VSS SDn_2.t69 SDn_1.t16 VSS.t128 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X399 VSS SDn_2.t70 SD3_1.t35 VSS.t283 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X400 OUT-.t26 b2.t5 OUT-.t26 VSS.t188 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X401 VSS Balance_Inverter_3.Inverter_0.OUT b1.t0 VSS.t59 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X402 Balance_Inverter_4.Inverter_0.OUT B5.t2 VDD.t66 VDD.t65 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X403 OUT-.t78 b6.t38 OUT-.t78 VSS.t72 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X404 OUT6 b6b.t39 OUT-.t55 VSS.t19 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X405 OUT+ b4.t15 OUT4.t12 VSS.t228 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X406 OUT+ b5.t20 OUT5.t36 VSS.t186 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X407 OUT5 IT.t64 SDn_1.t3 VSS.t49 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X408 OUT-.t119 OUT-.t118 OUT-.t119 VSS.t109 nfet_03v3 ad=94.8f pd=0.92u as=0 ps=0 w=0.3u l=0.5u
X409 SD3_1 IT.t65 OUT6.t12 VSS.t169 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X410 OUT+.t47 OUT+.t46 OUT+.t47 VSS.t44 nfet_03v3 ad=0 pd=0 as=94.8f ps=0.92u w=0.3u l=0.5u
X411 OUT- b5b.t20 OUT5.t19 VSS.t200 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X412 OUT6 b6.t39 OUT+.t6 VSS.t17 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X413 OUT- b5b.t21 OUT5.t18 VSS.t191 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X414 SD2_4 G2.t22 VSS.t63 VSS.t62 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X415 OUT6 b6b.t40 OUT-.t56 VSS.t17 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X416 Balance_Inverter_2.Inverter_0.OUT B2.t2 VDD.t68 VDD.t67 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X417 OUT+ b3.t9 OUT3.t1 VSS.t70 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X418 OUT+ b5.t21 OUT5.t37 VSS.t197 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X419 OUT+.t45 OUT+.t44 OUT+.t45 VSS.t91 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X420 OUT+ b4.t16 OUT4.t13 VSS.t210 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X421 OUT+.t167 b5b.t22 OUT+.t167 VSS.t202 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X422 OUT6 IT.t66 SD3_1.t26 VSS.t293 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X423 OUT+.t43 OUT+.t42 OUT+.t43 VSS.t91 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X424 OUT-.t29 b5.t22 OUT-.t29 VSS.t195 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X425 OUT+ b6.t40 OUT6.t67 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X426 OUT6 b6b.t41 OUT-.t24 VSS.t18 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X427 OUT6 b6b.t42 OUT-.t25 VSS.t18 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X428 SD2_5 ITAIL.t21 OUT4.t6 VSS.t113 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X429 IT IT.t4 SDn_2.t16 VSS.t324 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X430 OUT+.t151 b5b.t23 OUT+.t151 VSS.t203 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X431 OUT+.t41 OUT+.t40 OUT+.t41 VSS.t139 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X432 OUT6 IT.t68 SD3_1.t22 VSS.t171 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X433 OUT+.t152 b5b.t24 OUT+.t152 VSS.t29 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X434 OUT4 b4.t17 OUT+.t9 VSS.t34 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X435 VSS SDn_2.t2 SDn_2.t3 VSS.t175 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X436 OUT+.t39 OUT+.t38 OUT+.t39 VSS.t111 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X437 OUT-.t77 b6.t41 OUT-.t77 VSS.t90 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X438 SD3_1 SDn_2.t71 VSS.t286 VSS.t131 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X439 SD3_1 SDn_2.t72 VSS.t335 VSS.t127 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X440 OUT4 b4b.t16 OUT-.t52 VSS.t118 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X441 OUT+ b6.t42 OUT6.t66 VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X442 OUT-.t117 OUT-.t116 OUT-.t117 VSS.t81 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X443 OUT-.t115 OUT-.t114 OUT-.t115 VSS.t67 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X444 OUT-.t113 OUT-.t112 OUT-.t113 VSS.t93 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X445 VDD b2b.t5 b2.t0 VDD.t0 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X446 VDD G1_1.t10 G1_1.t11 VDD.t31 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X447 VSS G2.t23 SD2_1.t1 VSS.t64 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X448 SD3_1 SDn_2.t73 VSS.t336 VSS.t149 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X449 OUT5 b5.t23 OUT+.t132 VSS.t190 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X450 OUT+.t37 OUT+.t36 OUT+.t37 VSS.t136 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X451 VDD G1_1.t32 SD1_1.t8 VDD.t21 pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X452 OUT- b3b.t8 OUT3.t0 VSS.t23 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X453 OUT+ b5.t24 OUT5.t33 VSS.t186 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X454 OUT5 b5b.t25 OUT-.t182 VSS.t29 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X455 VSS SDn_2.t74 SD3_1.t31 VSS.t150 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X456 OUT-.t41 b3.t10 OUT-.t41 VSS.t68 nfet_03v3 ad=94.8f pd=0.92u as=0 ps=0 w=0.3u l=0.5u
X457 G1_2 G1_2.t14 G1_1.t2 VDD.t72 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X458 OUT- b5b.t26 OUT5.t16 VSS.t200 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X459 SD2_1 ITAIL.t22 G1_2.t17 VSS.t30 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X460 G1_1 G1_2.t6 G1_2.t7 VDD.t18 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X461 SD2_1 G2.t24 VSS.t1 VSS.t0 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X462 OUT2 b2b.t6 OUT-.t5 VSS.t25 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X463 VDD b6b.t43 b6.t1 VDD.t95 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X464 OUT-.t10 b4.t18 OUT-.t10 VSS.t35 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X465 OUT-.t76 b6.t43 OUT-.t76 VSS.t17 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X466 SDn_2 IT.t2 IT.t3 VSS.t87 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X467 OUT-.t111 OUT-.t110 OUT-.t111 VSS.t82 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X468 OUT+.t191 b6b.t44 OUT+.t191 VSS.t129 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X469 OUT+.t35 OUT+.t34 OUT+.t35 VSS.t81 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X470 OUT-.t109 OUT-.t108 OUT-.t109 VSS.t81 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X471 OUT-.t107 OUT-.t106 OUT-.t107 VSS.t93 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X472 G1_1 G1_1.t8 VDD.t46 VDD.t45 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X473 OUT5 b5.t25 OUT+.t131 VSS.t28 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X474 OUT+.t10 b6b.t45 OUT+.t10 VSS.t39 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X475 b6b b6.t44 VDD.t16 VDD.t15 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X476 OUT6 IT.t69 SD3_1.t23 VSS.t299 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X477 OUT-.t75 b6.t45 OUT-.t75 VSS.t89 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X478 Balance_Inverter_1.Inverter_0.OUT B3.t1 VSS.t121 VSS.t120 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X479 VSS G2.t25 SD2_2.t0 VSS.t2 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X480 OUT- b4b.t17 OUT4.t14 VSS.t32 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X481 OUT+.t33 OUT+.t32 OUT+.t33 VSS.t138 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X482 OUT+.t31 OUT+.t30 OUT+.t31 VSS.t137 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X483 IT IT.t0 SDn_2.t20 VSS.t165 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X484 OUT-.t91 b1.t4 OUT-.t91 VSS.t231 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X485 OUT-.t105 OUT-.t104 OUT-.t105 VSS.t112 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X486 OUT6 IT.t71 SD3_1.t24 VSS.t242 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X487 OUT+.t11 b6b.t46 OUT+.t11 VSS.t40 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X488 SDn_1 IT.t72 OUT5.t0 VSS.t273 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X489 OUT- b6b.t47 OUT6.t0 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X490 SD2_4 ITAIL.t23 OUT3.t6 VSS.t31 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X491 SD1_1 G1_1.t34 VDD.t25 VDD.t24 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X492 IT G1_2.t34 SD1_1.t0 VDD.t79 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X493 OUT- b6b.t48 OUT6.t1 VSS.t21 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X494 OUT+.t29 OUT+.t28 OUT+.t29 VSS.t136 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X495 SD3_1 IT.t73 OUT6.t7 VSS.t100 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X496 OUT6 b6.t46 OUT+.t174 VSS.t19 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X497 SD2_1 ITAIL.t24 G1_2.t16 VSS.t119 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X498 OUT6 b6.t47 OUT+.t22 VSS.t19 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X499 b3b B3.t2 VSS.t313 VSS.t312 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X500 OUT2 b2.t6 OUT+.t128 VSS.t189 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X501 OUT+.t4 b3b.t9 OUT+.t4 VSS.t24 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X502 OUT+ b6.t48 OUT6.t63 VSS.t41 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X503 OUT+ b6.t49 OUT6.t62 VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X504 OUT+.t176 b6b.t49 OUT+.t176 VSS.t187 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X505 OUT-.t103 OUT-.t102 OUT-.t103 VSS.t111 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X506 OUT-.t101 OUT-.t100 OUT-.t101 VSS.t93 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X507 OUT5 IT.t74 SDn_1.t1 VSS.t296 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X508 OUT-.t99 OUT-.t98 OUT-.t99 VSS.t148 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X509 OUT+.t162 b4b.t18 OUT+.t162 VSS.t117 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X510 OUT6 b6.t50 OUT+.t121 VSS.t16 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X511 VSS SDn_2.t75 SD3_1.t30 VSS.t135 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X512 OUT5 b5.t26 OUT+.t129 VSS.t194 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X513 OUT5 IT.t75 SDn_1.t0 VSS.t239 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X514 G1_2 G1_2.t0 G1_1.t0 VDD.t34 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X515 VDD G1_1.t35 SD1_1.t13 VDD.t80 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X516 OUT+.t177 b6b.t50 OUT+.t177 VSS.t17 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X517 OUT3 b3b.t10 OUT-.t93 VSS.t314 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X518 VSS SDn_2.t0 SDn_2.t1 VSS.t324 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
R0 OUT+.n3 OUT+.t58 37.0108
R1 OUT+.n1 OUT+.t46 22.8811
R2 OUT+.t84 OUT+.t52 20.3675
R3 OUT+.n238 OUT+.t84 19.9024
R4 OUT+.n17 OUT+.t40 15.8102
R5 OUT+.n9 OUT+.t108 15.18
R6 OUT+.n52 OUT+.t112 14.2205
R7 OUT+.n160 OUT+.t98 13.7825
R8 OUT+.n276 OUT+.t116 13.576
R9 OUT+.n45 OUT+.t66 12.9065
R10 OUT+.n35 OUT+.t56 12.6145
R11 OUT+.n290 OUT+.t30 12.1915
R12 OUT+.n63 OUT+.t42 11.9725
R13 OUT+.n96 OUT+.t70 11.7535
R14 OUT+.n190 OUT+.t86 11.7535
R15 OUT+.n93 OUT+.t34 11.6805
R16 OUT+.n75 OUT+.t82 11.6643
R17 OUT+.n203 OUT+.t114 11.5345
R18 OUT+.n248 OUT+.t88 11.5195
R19 OUT+.n212 OUT+.t100 11.4615
R20 OUT+.n101 OUT+.t102 11.3885
R21 OUT+.n59 OUT+.t60 11.2425
R22 OUT+.n179 OUT+.t28 11.2425
R23 OUT+.n119 OUT+.t104 11.0235
R24 OUT+.n55 OUT+.t90 11.0235
R25 OUT+.n185 OUT+.t68 11.0235
R26 OUT+.n254 OUT+.t118 10.8775
R27 OUT+.n226 OUT+.t110 10.6585
R28 OUT+.n119 OUT+.t48 10.5125
R29 OUT+.n55 OUT+.t38 10.5125
R30 OUT+.n185 OUT+.t76 10.5125
R31 OUT+.n17 OUT+.t72 10.5049
R32 OUT+.n1 OUT+.t74 10.3852
R33 OUT+.n59 OUT+.t94 10.2935
R34 OUT+.n179 OUT+.t36 10.2935
R35 OUT+.n101 OUT+.t44 10.1475
R36 OUT+.n226 OUT+.t78 10.0745
R37 OUT+.n203 OUT+.t32 10.0015
R38 OUT+.n75 OUT+.t106 9.96832
R39 OUT+.n290 OUT+.t50 9.8555
R40 OUT+.n93 OUT+.t62 9.8555
R41 OUT+.n96 OUT+.t92 9.7825
R42 OUT+.n190 OUT+.t96 9.7825
R43 OUT+.n63 OUT+.t80 9.5635
R44 OUT+.n254 OUT+.t54 9.4905
R45 OUT+.n212 OUT+.t64 9.2715
R46 OUT+.n273 OUT+.t156 8.57704
R47 OUT+.n250 OUT+.t163 8.55673
R48 OUT+.n26 OUT+.t171 8.53705
R49 OUT+.n27 OUT+.t175 8.4005
R50 OUT+.n274 OUT+.t164 8.4005
R51 OUT+.n232 OUT+.n231 8.22813
R52 OUT+.n265 OUT+.t155 7.8755
R53 OUT+.n235 OUT+.n234 6.39076
R54 OUT+.n116 OUT+.n113 6.15786
R55 OUT+.n99 OUT+.t71 6.14541
R56 OUT+.n143 OUT+.t43 6.14358
R57 OUT+.n152 OUT+.t127 6.12228
R58 OUT+.n153 OUT+.t24 6.1112
R59 OUT+.n98 OUT+.t93 6.10805
R60 OUT+.n142 OUT+.t81 6.10723
R61 OUT+.n187 OUT+.t69 6.10646
R62 OUT+.n187 OUT+.t77 6.09305
R63 OUT+.n229 OUT+.t149 6.09276
R64 OUT+.n144 OUT+.t91 6.07954
R65 OUT+.n4 OUT+.t120 6.07748
R66 OUT+.n144 OUT+.t39 6.06396
R67 OUT+.n161 OUT+.t99 6.02733
R68 OUT+.n221 OUT+.t161 5.9655
R69 OUT+.n29 OUT+.n28 5.8805
R70 OUT+.n285 OUT+.n30 5.8805
R71 OUT+.n157 OUT+.t191 5.8805
R72 OUT+.n38 OUT+.t122 5.8805
R73 OUT+.n37 OUT+.t177 5.8805
R74 OUT+.n148 OUT+.t150 5.8805
R75 OUT+.n49 OUT+.t176 5.8805
R76 OUT+.n222 OUT+.t147 5.8805
R77 OUT+.n217 OUT+.t152 5.8805
R78 OUT+.n230 OUT+.t151 5.8805
R79 OUT+.n244 OUT+.n243 5.68489
R80 OUT+.n154 OUT+.n153 5.58414
R81 OUT+.n6 OUT+.t123 5.2505
R82 OUT+.n6 OUT+.t47 5.2505
R83 OUT+.n23 OUT+.t4 5.2505
R84 OUT+.n22 OUT+.t188 5.2505
R85 OUT+.n247 OUT+.t89 5.2505
R86 OUT+.n277 OUT+.t160 5.2505
R87 OUT+.n277 OUT+.t117 5.2505
R88 OUT+.n271 OUT+.t162 5.2505
R89 OUT+.n270 OUT+.t159 5.2505
R90 OUT+.n146 OUT+.n145 4.78361
R91 OUT+.n168 OUT+.n165 4.65832
R92 OUT+.n232 OUT+.n161 4.51156
R93 OUT+.n208 OUT+.n168 4.34231
R94 OUT+.n251 OUT+.t158 4.18308
R95 OUT+.n209 OUT+.t146 4.1532
R96 OUT+.n2 OUT+.n1 4.0005
R97 OUT+.n18 OUT+.n17 4.0005
R98 OUT+.n292 OUT+.n290 4.0005
R99 OUT+.n255 OUT+.n254 4.0005
R100 OUT+.n77 OUT+.n75 4.0005
R101 OUT+.n94 OUT+.n93 4.0005
R102 OUT+.n97 OUT+.n96 4.0005
R103 OUT+.n102 OUT+.n101 4.0005
R104 OUT+.n121 OUT+.n119 4.0005
R105 OUT+.n141 OUT+.n63 4.0005
R106 OUT+.n60 OUT+.n59 4.0005
R107 OUT+.n180 OUT+.n179 4.0005
R108 OUT+.n186 OUT+.n185 4.0005
R109 OUT+.n191 OUT+.n190 4.0005
R110 OUT+.n205 OUT+.n203 4.0005
R111 OUT+.n214 OUT+.n212 4.0005
R112 OUT+.n227 OUT+.n226 4.0005
R113 OUT+.n198 OUT+.n177 3.7799
R114 OUT+.n138 OUT+.n137 3.71391
R115 OUT+.n68 OUT+.n67 3.66911
R116 OUT+.n87 OUT+.n84 3.65144
R117 OUT+.n240 OUT+.n237 3.61617
R118 OUT+.n284 OUT+.n268 3.54956
R119 OUT+.n294 OUT+.n286 3.54793
R120 OUT+.n21 OUT+.n20 3.53029
R121 OUT+.n289 OUT+.n288 3.47675
R122 OUT+.n168 OUT+.n167 3.46146
R123 OUT+.n220 OUT+.n162 3.44883
R124 OUT+.n184 OUT+.n183 3.43965
R125 OUT+.n116 OUT+.n115 3.42587
R126 OUT+.n289 OUT+.n287 3.42532
R127 OUT+.n182 OUT+.n181 3.42241
R128 OUT+.n128 OUT+.n127 3.41469
R129 OUT+.n124 OUT+.n70 3.40991
R130 OUT+.n177 OUT+.n176 3.39679
R131 OUT+.n177 OUT+.n174 3.39572
R132 OUT+.n10 OUT+.t14 3.39531
R133 OUT+.n194 OUT+.n193 3.39468
R134 OUT+.n206 OUT+.n202 3.38986
R135 OUT+.n151 OUT+.n42 3.38009
R136 OUT+.n155 OUT+.n40 3.38009
R137 OUT+.n79 OUT+.n78 3.37228
R138 OUT+.n109 OUT+.n108 3.3721
R139 OUT+.n244 OUT+.n235 3.36946
R140 OUT+.n151 OUT+.n43 3.36356
R141 OUT+.n155 OUT+.n39 3.36356
R142 OUT+.n95 OUT+.n91 3.36276
R143 OUT+.n256 OUT+.n246 3.3575
R144 OUT+.n272 OUT+.n271 3.35621
R145 OUT+.n61 OUT+.n57 3.353
R146 OUT+.n215 OUT+.n211 3.3505
R147 OUT+.n272 OUT+.n270 3.34657
R148 OUT+.n61 OUT+.n56 3.33742
R149 OUT+.n228 OUT+.n224 3.3339
R150 OUT+.n103 OUT+.n89 3.3305
R151 OUT+.n111 OUT+.n82 3.3267
R152 OUT+.n228 OUT+.n223 3.32031
R153 OUT+.n95 OUT+.n90 3.31861
R154 OUT+.n36 OUT+.n34 3.31162
R155 OUT+.n19 OUT+.n16 3.3089
R156 OUT+ OUT+.n296 3.30598
R157 OUT+.n25 OUT+.n23 3.29947
R158 OUT+.n46 OUT+.n44 3.2981
R159 OUT+.n215 OUT+.n210 3.2955
R160 OUT+.n54 OUT+.n53 3.28884
R161 OUT+.n25 OUT+.n22 3.28705
R162 OUT+.n159 OUT+.n33 3.28638
R163 OUT+.n20 OUT+.n15 3.27572
R164 OUT+.n220 OUT+.n163 3.2355
R165 OUT+.n10 OUT+.t15 3.1617
R166 OUT+.n7 OUT+.n6 3.15377
R167 OUT+.n13 OUT+.n12 3.1505
R168 OUT+.n249 OUT+.n247 3.1505
R169 OUT+.n138 OUT+.n135 3.1505
R170 OUT+.n106 OUT+.n105 3.1505
R171 OUT+.n87 OUT+.n86 3.1505
R172 OUT+.n112 OUT+.n80 3.1505
R173 OUT+.n117 OUT+.n74 3.1505
R174 OUT+.n118 OUT+.n72 3.1505
R175 OUT+.n123 OUT+.n71 3.1505
R176 OUT+.n131 OUT+.n130 3.1505
R177 OUT+.n139 OUT+.n133 3.1505
R178 OUT+.n278 OUT+.n277 3.1505
R179 OUT+.n259 OUT+.n258 3.14382
R180 OUT+.n3 OUT+.t59 2.93148
R181 OUT+.n128 OUT+.n125 2.89661
R182 OUT+.n125 OUT+.n124 2.89194
R183 OUT+.n111 OUT+.n110 2.89154
R184 OUT+.n110 OUT+.n109 2.88693
R185 OUT+.n199 OUT+.n172 2.76701
R186 OUT+.n200 OUT+.n170 2.76641
R187 OUT+.n12 OUT+.t109 2.7305
R188 OUT+.n12 OUT+.n11 2.7305
R189 OUT+.n15 OUT+.t128 2.7305
R190 OUT+.n15 OUT+.t41 2.7305
R191 OUT+.n16 OUT+.t73 2.7305
R192 OUT+.n288 OUT+.t179 2.7305
R193 OUT+.n288 OUT+.t31 2.7305
R194 OUT+.n287 OUT+.t16 2.7305
R195 OUT+.n287 OUT+.t51 2.7305
R196 OUT+.n258 OUT+.t55 2.7305
R197 OUT+.n258 OUT+.n257 2.7305
R198 OUT+.n246 OUT+.t119 2.7305
R199 OUT+.n246 OUT+.n245 2.7305
R200 OUT+.n234 OUT+.t9 2.7305
R201 OUT+.n234 OUT+.n233 2.7305
R202 OUT+.n34 OUT+.t57 2.7305
R203 OUT+.n133 OUT+.n132 2.7305
R204 OUT+.n135 OUT+.t186 2.7305
R205 OUT+.n135 OUT+.n134 2.7305
R206 OUT+.n137 OUT+.t168 2.7305
R207 OUT+.n137 OUT+.n136 2.7305
R208 OUT+.n130 OUT+.n129 2.7305
R209 OUT+.n71 OUT+.t169 2.7305
R210 OUT+.n71 OUT+.t49 2.7305
R211 OUT+.n72 OUT+.t189 2.7305
R212 OUT+.n72 OUT+.t105 2.7305
R213 OUT+.n74 OUT+.t12 2.7305
R214 OUT+.n74 OUT+.n73 2.7305
R215 OUT+.n78 OUT+.t1 2.7305
R216 OUT+.n78 OUT+.t107 2.7305
R217 OUT+.n80 OUT+.t6 2.7305
R218 OUT+.n80 OUT+.t83 2.7305
R219 OUT+.n105 OUT+.t103 2.7305
R220 OUT+.n105 OUT+.n104 2.7305
R221 OUT+.n89 OUT+.t45 2.7305
R222 OUT+.n89 OUT+.n88 2.7305
R223 OUT+.n91 OUT+.t35 2.7305
R224 OUT+.n90 OUT+.t63 2.7305
R225 OUT+.n108 OUT+.t2 2.7305
R226 OUT+.n108 OUT+.n107 2.7305
R227 OUT+.n84 OUT+.t174 2.7305
R228 OUT+.n84 OUT+.n83 2.7305
R229 OUT+.n86 OUT+.t26 2.7305
R230 OUT+.n86 OUT+.n85 2.7305
R231 OUT+.n82 OUT+.t0 2.7305
R232 OUT+.n82 OUT+.n81 2.7305
R233 OUT+.n115 OUT+.t121 2.7305
R234 OUT+.n115 OUT+.n114 2.7305
R235 OUT+.n70 OUT+.t170 2.7305
R236 OUT+.n70 OUT+.n69 2.7305
R237 OUT+.n67 OUT+.t22 2.7305
R238 OUT+.n67 OUT+.n66 2.7305
R239 OUT+.n65 OUT+.t3 2.7305
R240 OUT+.n65 OUT+.n64 2.7305
R241 OUT+.n127 OUT+.t157 2.7305
R242 OUT+.n127 OUT+.n126 2.7305
R243 OUT+.n57 OUT+.t61 2.7305
R244 OUT+.n56 OUT+.t95 2.7305
R245 OUT+.n53 OUT+.t113 2.7305
R246 OUT+.n44 OUT+.t67 2.7305
R247 OUT+.n43 OUT+.t10 2.7305
R248 OUT+.n42 OUT+.t166 2.7305
R249 OUT+.n40 OUT+.t178 2.7305
R250 OUT+.n39 OUT+.t19 2.7305
R251 OUT+.n33 OUT+.t20 2.7305
R252 OUT+.n163 OUT+.t148 2.7305
R253 OUT+.n162 OUT+.t167 2.7305
R254 OUT+.n165 OUT+.t131 2.7305
R255 OUT+.n165 OUT+.n164 2.7305
R256 OUT+.n167 OUT+.t132 2.7305
R257 OUT+.n167 OUT+.n166 2.7305
R258 OUT+.n170 OUT+.t138 2.7305
R259 OUT+.n170 OUT+.n169 2.7305
R260 OUT+.n172 OUT+.t143 2.7305
R261 OUT+.n172 OUT+.n171 2.7305
R262 OUT+.n174 OUT+.t129 2.7305
R263 OUT+.n174 OUT+.n173 2.7305
R264 OUT+.n176 OUT+.t142 2.7305
R265 OUT+.n176 OUT+.n175 2.7305
R266 OUT+.n196 OUT+.t97 2.7305
R267 OUT+.n196 OUT+.n195 2.7305
R268 OUT+.n183 OUT+.t29 2.7305
R269 OUT+.n181 OUT+.t37 2.7305
R270 OUT+.n193 OUT+.t87 2.7305
R271 OUT+.n193 OUT+.n192 2.7305
R272 OUT+.n201 OUT+.t140 2.7305
R273 OUT+.n201 OUT+.t33 2.7305
R274 OUT+.n202 OUT+.t139 2.7305
R275 OUT+.n202 OUT+.t115 2.7305
R276 OUT+.n211 OUT+.t101 2.7305
R277 OUT+.n210 OUT+.t65 2.7305
R278 OUT+.n224 OUT+.t111 2.7305
R279 OUT+.n223 OUT+.t79 2.7305
R280 OUT+.n243 OUT+.t124 2.7305
R281 OUT+.n243 OUT+.n242 2.7305
R282 OUT+.n236 OUT+.t125 2.7305
R283 OUT+.n236 OUT+.t85 2.7305
R284 OUT+.n237 OUT+.t25 2.7305
R285 OUT+.n237 OUT+.t53 2.7305
R286 OUT+.n0 OUT+.t75 2.57389
R287 OUT+.n110 OUT+.n87 2.57097
R288 OUT+.n48 OUT+.n47 2.50602
R289 OUT+.n147 OUT+.n51 2.47399
R290 OUT+.n296 OUT+.n8 2.32319
R291 OUT+.n251 OUT+.n250 2.25866
R292 OUT+.n21 OUT+.n14 2.2505
R293 OUT+.n294 OUT+.n293 2.2505
R294 OUT+.n296 OUT+.n295 2.11341
R295 OUT+.n62 OUT+.n55 2.10931
R296 OUT+.n2 OUT+.n0 2.10014
R297 OUT+.n47 OUT+.t11 2.02309
R298 OUT+.n51 OUT+.t21 2.0096
R299 OUT+.n209 OUT+.n208 1.9401
R300 OUT+.n198 OUT+.n197 1.89913
R301 OUT+.n207 OUT+.n201 1.84038
R302 OUT+.n241 OUT+.n236 1.83827
R303 OUT+.n68 OUT+.n65 1.83747
R304 OUT+.n51 OUT+.t145 1.81249
R305 OUT+.n47 OUT+.t23 1.80341
R306 OUT+.n244 OUT+.n241 1.72491
R307 OUT+.n13 OUT+.n10 1.67253
R308 OUT+.n208 OUT+.n207 1.65485
R309 OUT+.n235 OUT+.n232 1.60321
R310 OUT+.n218 OUT+.n217 1.6005
R311 OUT+.n265 OUT+.n264 1.50139
R312 OUT+.n197 OUT+.n196 1.42583
R313 OUT+.n231 OUT+.n222 1.29515
R314 OUT+.n118 OUT+.n117 1.283
R315 OUT+.n139 OUT+.n138 1.27582
R316 OUT+.n200 OUT+.n199 1.25824
R317 OUT+.n285 OUT+.n284 1.24838
R318 OUT+.n262 OUT+.n261 1.12395
R319 OUT+.n125 OUT+.n68 1.10964
R320 OUT+.n279 OUT+.n275 1.0955
R321 OUT+.n112 OUT+.n111 1.0351
R322 OUT+.n124 OUT+.n123 1.01651
R323 OUT+.n131 OUT+.n128 1.00696
R324 OUT+.n109 OUT+.n106 0.988998
R325 OUT+.n264 OUT+.n263 0.978718
R326 OUT+.n149 OUT+.n148 0.907373
R327 OUT+.n295 OUT+.n294 0.898066
R328 OUT+.n252 OUT+.n251 0.886808
R329 OUT+.n38 OUT+.n37 0.828076
R330 OUT+.n50 OUT+.n49 0.810602
R331 OUT+.n5 OUT+.n4 0.78333
R332 OUT+.n158 OUT+.n157 0.782551
R333 OUT+.n29 OUT+.n27 0.779029
R334 OUT+.n262 OUT+.n244 0.727459
R335 OUT+.n275 OUT+.n274 0.713635
R336 OUT+.n295 OUT+.n21 0.659429
R337 OUT+.n159 OUT+.n158 0.489391
R338 OUT+.n37 OUT+.n36 0.4343
R339 OUT+.n283 OUT+.n282 0.4055
R340 OUT+.n156 OUT+.n155 0.378867
R341 OUT+.n151 OUT+.n150 0.37152
R342 OUT+.n260 OUT+.n259 0.352867
R343 OUT+.n239 OUT+.n238 0.345125
R344 OUT+.n4 OUT+.n3 0.34121
R345 OUT+.n278 OUT+.n276 0.339348
R346 OUT+.n221 OUT+.n220 0.338833
R347 OUT+.n220 OUT+.n219 0.338833
R348 OUT+.n26 OUT+.n25 0.334121
R349 OUT+.n284 OUT+.n283 0.33333
R350 OUT+.n229 OUT+.n228 0.330157
R351 OUT+.n25 OUT+.n24 0.326362
R352 OUT+.n273 OUT+.n272 0.318962
R353 OUT+.n272 OUT+.n269 0.317231
R354 OUT+.n216 OUT+.n215 0.316523
R355 OUT+.n48 OUT+.n46 0.311122
R356 OUT+.n155 OUT+.n154 0.306316
R357 OUT+.n20 OUT+.n19 0.305311
R358 OUT+.n8 OUT+.n2 0.300773
R359 OUT+.n219 OUT+.n218 0.298833
R360 OUT+.n222 OUT+.n221 0.298833
R361 OUT+.n152 OUT+.n151 0.296214
R362 OUT+.n7 OUT+.n5 0.291543
R363 OUT+.n286 OUT+.n285 0.280577
R364 OUT+.n14 OUT+.n9 0.2705
R365 OUT+.n117 OUT+.n116 0.260555
R366 OUT+.n249 OUT+.n248 0.251632
R367 OUT+.n199 OUT+.n198 0.245769
R368 OUT+.n113 OUT+.n112 0.243546
R369 OUT+.n286 OUT+.n29 0.227418
R370 OUT+.n156 OUT+.n38 0.225986
R371 OUT+.n140 OUT+.n139 0.2255
R372 OUT+.n150 OUT+.n50 0.224402
R373 OUT+.n253 OUT+.n252 0.220713
R374 OUT+.n231 OUT+.n230 0.218864
R375 OUT+.n106 OUT+.n103 0.211066
R376 OUT+.n157 OUT+.n156 0.204718
R377 OUT+.n122 OUT+.n118 0.203
R378 OUT+.n150 OUT+.n149 0.20194
R379 OUT+.n216 OUT+.n209 0.200502
R380 OUT+.n54 OUT+.n52 0.191791
R381 OUT+.n123 OUT+.n122 0.190885
R382 OUT+.n208 OUT+.n200 0.187837
R383 OUT+.n8 OUT+.n7 0.187108
R384 OUT+.n49 OUT+.n48 0.185692
R385 OUT+.n207 OUT+.n206 0.185073
R386 OUT+.n230 OUT+.n229 0.1805
R387 OUT+.n240 OUT+.n239 0.172786
R388 OUT+.n217 OUT+.n216 0.172167
R389 OUT+.n250 OUT+.n249 0.167221
R390 OUT+.n140 OUT+.n131 0.166654
R391 OUT+.n274 OUT+.n273 0.166654
R392 OUT+.n197 OUT+.n194 0.164383
R393 OUT+.n259 OUT+.n256 0.155767
R394 OUT+.n36 OUT+.n35 0.153345
R395 OUT+.n27 OUT+.n26 0.149466
R396 OUT+.n160 OUT+.n159 0.149123
R397 OUT+.n194 OUT+.n191 0.143115
R398 OUT+.n188 OUT+.n187 0.142318
R399 OUT+.n61 OUT+.n60 0.141929
R400 OUT+.n100 OUT+.n99 0.141731
R401 OUT+.n102 OUT+.n100 0.140346
R402 OUT+.n103 OUT+.n102 0.140346
R403 OUT+.n60 OUT+.n58 0.140346
R404 OUT+.n187 OUT+.n186 0.139591
R405 OUT+.n141 OUT+.n140 0.137457
R406 OUT+.n122 OUT+.n121 0.136824
R407 OUT+.n256 OUT+.n255 0.1355
R408 OUT+.n180 OUT+.n178 0.1355
R409 OUT+.n205 OUT+.n204 0.134848
R410 OUT+.n255 OUT+.n253 0.134176
R411 OUT+.n77 OUT+.n76 0.134176
R412 OUT+.n206 OUT+.n205 0.133543
R413 OUT+.n121 OUT+.n120 0.132853
R414 OUT+.n46 OUT+.n45 0.132817
R415 OUT+.n95 OUT+.n94 0.131063
R416 OUT+.n97 OUT+.n95 0.129886
R417 OUT+.n62 OUT+.n61 0.128884
R418 OUT+.n144 OUT+.n143 0.12855
R419 OUT+.n94 OUT+.n92 0.127261
R420 OUT+.n147 OUT+.n146 0.125565
R421 OUT+.n279 OUT+.n278 0.124462
R422 OUT+.n227 OUT+.n225 0.122474
R423 OUT+.n228 OUT+.n227 0.122474
R424 OUT+.n214 OUT+.n213 0.12089
R425 OUT+.n215 OUT+.n214 0.119721
R426 OUT+.n292 OUT+.n291 0.116375
R427 OUT+.n148 OUT+.n147 0.1157
R428 OUT+.n281 OUT+.n280 0.113979
R429 OUT+.n191 OUT+.n189 0.109885
R430 OUT+.n186 OUT+.n184 0.108227
R431 OUT+.n182 OUT+.n180 0.103735
R432 OUT+.n145 OUT+.n144 0.102011
R433 OUT+.n142 OUT+.n141 0.0983261
R434 OUT+.n98 OUT+.n97 0.0982143
R435 OUT+.n293 OUT+.n292 0.093875
R436 OUT+.n79 OUT+.n77 0.0905
R437 OUT+.n14 OUT+.n13 0.0851915
R438 OUT+.n146 OUT+.n54 0.0829875
R439 OUT+.n268 OUT+.n267 0.068
R440 OUT+.n241 OUT+.n240 0.063158
R441 OUT+.n282 OUT+.n281 0.0450426
R442 OUT+.n161 OUT+.n160 0.0442269
R443 OUT+.n263 OUT+.n262 0.0385186
R444 OUT+.n19 OUT+.n18 0.0321216
R445 OUT+.n145 OUT+.n62 0.0305639
R446 OUT+.n267 OUT+.n266 0.0301053
R447 OUT+.n154 OUT+.n41 0.0258846
R448 OUT+.n143 OUT+.n142 0.0212692
R449 OUT+.n189 OUT+.n188 0.017734
R450 OUT+.n261 OUT+.n260 0.0169634
R451 OUT+.n113 OUT+.n79 0.0147857
R452 OUT+.n153 OUT+.n152 0.0131761
R453 OUT+.n264 OUT+.n32 0.00905914
R454 OUT+.n99 OUT+.n98 0.00899057
R455 OUT+.n293 OUT+.n289 0.008375
R456 OUT+.n282 OUT+.n279 0.00559434
R457 OUT+.n184 OUT+.n182 0.00432979
R458 OUT+.n32 OUT+.n31 0.002375
R459 OUT+.n266 OUT+.n265 0.00168421
R460 VSS.t278 VSS.n944 2045.19
R461 VSS.t312 VSS.n940 2003.92
R462 VSS.t217 VSS.n948 2003.92
R463 VSS.n1000 VSS 1757.65
R464 VSS.n884 VSS.t183 1708.91
R465 VSS VSS.n1000 1677.99
R466 VSS.n1000 VSS 1677.99
R467 VSS.n886 VSS.t114 1561.78
R468 VSS.n883 VSS.t325 1530.27
R469 VSS.n885 VSS.t59 1530.27
R470 VSS.n884 VSS.n883 1500.56
R471 VSS.n887 VSS.n886 1436.69
R472 VSS.n887 VSS.n885 1407.7
R473 VSS.t221 VSS.n1010 1129.9
R474 VSS.n877 VSS.t310 1129.9
R475 VSS.n868 VSS.t333 1129.9
R476 VSS.t310 VSS.n876 1121.68
R477 VSS.n1011 VSS.t221 1101.14
R478 VSS.n875 VSS.n874 1092.92
R479 VSS.n1013 VSS.n1012 1092.92
R480 VSS.n1010 VSS.t46 1072.38
R481 VSS.t183 VSS.n877 1072.38
R482 VSS.t319 VSS.n868 1072.38
R483 VSS.n949 VSS.t278 1070.94
R484 VSS.n949 VSS.t312 1049.33
R485 VSS.n949 VSS.t217 1049.33
R486 VSS.n1012 VSS.t319 862.832
R487 VSS VSS.n873 797.03
R488 VSS VSS.n1014 797.03
R489 VSS VSS.n879 797.03
R490 VSS.n876 VSS.n875 530.025
R491 VSS.n1013 VSS.n1011 513.591
R492 VSS.n1000 VSS.n887 268.024
R493 VSS.n147 VSS.n146 220.651
R494 VSS.n1000 VSS.n884 157.843
R495 VSS.n142 VSS.t169 98.195
R496 VSS.n88 VSS.t123 93.4051
R497 VSS.n132 VSS.t154 88.6151
R498 VSS.t38 VSS.t254 86.2201
R499 VSS.t49 VSS.t94 86.2201
R500 VSS.n1000 VSS.n999 86.0069
R501 VSS.n75 VSS.t245 83.8251
R502 VSS.t134 VSS.t87 76.6401
R503 VSS.n85 VSS.t128 74.2452
R504 VSS.n959 VSS.n958 73.6511
R505 VSS.n1313 VSS.t126 69.4552
R506 VSS.n352 VSS.t145 68.8564
R507 VSS.n112 VSS.t133 67.0602
R508 VSS.n141 VSS.t122 67.0602
R509 VSS.n41 VSS.t152 65.8627
R510 VSS.n343 VSS.t189 64.9218
R511 VSS.n963 VSS.t76 64.2774
R512 VSS.n71 VSS.t302 62.2702
R513 VSS.n310 VSS.t267 61.9708
R514 VSS.n973 VSS.t7 57.8594
R515 VSS.n118 VSS.t171 57.4802
R516 VSS.n135 VSS.t269 57.4802
R517 VSS.n82 VSS.t57 55.0852
R518 VSS.n950 VSS.n949 55.0085
R519 VSS.n968 VSS.t155 54.2106
R520 VSS.n295 VSS.t71 54.1016
R521 VSS.n979 VSS.n978 53.1681
R522 VSS.n298 VSS.t70 52.1343
R523 VSS.t280 VSS.t79 52.1343
R524 VSS.t33 VSS.t24 52.1343
R525 VSS.n968 VSS.t318 52.1256
R526 VSS.n325 VSS.t188 51.1506
R527 VSS.n1315 VSS.t150 50.2953
R528 VSS.n973 VSS.t0 48.4768
R529 VSS.n331 VSS.t328 47.216
R530 VSS.n38 VSS.t54 46.7028
R531 VSS.n127 VSS.t165 45.5053
R532 VSS.n974 VSS.t30 44.3068
R533 VSS.t139 VSS.t228 43.2814
R534 VSS.t182 VSS.t142 43.2814
R535 VSS.n313 VSS.t137 42.2977
R536 VSS.n969 VSS.t13 40.6581
R537 VSS.n316 VSS.t174 40.3304
R538 VSS.n334 VSS.t44 39.3467
R539 VSS.n322 VSS.t215 38.3631
R540 VSS.n653 VSS.t72 38.1825
R541 VSS.n934 VSS.t113 36.241
R542 VSS.n113 VSS.t131 35.9253
R543 VSS.n80 VSS.t49 35.9253
R544 VSS.n138 VSS.t275 35.9253
R545 VSS.n660 VSS.t16 35.5939
R546 VSS.n1137 VSS.t82 35.5939
R547 VSS.n634 VSS.t181 34.9467
R548 VSS.n972 VSS.t108 34.9243
R549 VSS.n1203 VSS.t5 34.2996
R550 VSS.n625 VSS.t91 33.6524
R551 VSS.n958 VSS.t45 33.478
R552 VSS.n1250 VSS.t208 33.0053
R553 VSS.n666 VSS.t26 32.3581
R554 VSS.n1256 VSS.t198 31.711
R555 VSS.n1317 VSS.t127 31.1354
R556 VSS.n128 VSS.t242 31.1354
R557 VSS.n675 VSS.t93 31.0638
R558 VSS.n215 VSS.n214 31.0638
R559 VSS.n226 VSS.n225 30.4167
R560 VSS.n905 VSS.t2 29.4607
R561 VSS.n628 VSS.t227 28.4752
R562 VSS.n950 VSS.n938 28.4752
R563 VSS.n999 VSS.t73 28.1481
R564 VSS.n36 VSS.t261 27.5429
R565 VSS.n970 VSS.t104 27.1056
R566 VSS.n313 VSS.t68 26.5592
R567 VSS.n221 VSS.t194 26.5338
R568 VSS.n187 VSS.t153 26.3454
R569 VSS.n117 VSS.t132 26.3454
R570 VSS.n56 VSS.t178 26.3454
R571 VSS.n136 VSS.t306 26.3454
R572 VSS.n210 VSS.t199 25.8866
R573 VSS.n1215 VSS.t195 25.8866
R574 VSS.n337 VSS.t210 25.5756
R575 VSS.n340 VSS.t216 23.6082
R576 VSS.n1268 VSS.t106 23.298
R577 VSS.t117 VSS.t21 22.6508
R578 VSS.t105 VSS.t197 22.0037
R579 VSS.n105 VSS.t135 21.5554
R580 VSS.n1329 VSS.t239 21.5554
R581 VSS.n663 VSS.t148 21.3565
R582 VSS.n657 VSS.n656 20.7094
R583 VSS.n949 VSS.t62 20.5066
R584 VSS.n646 VSS.t40 20.0622
R585 VSS.n663 VSS.t22 18.1208
R586 VSS.n1285 VSS.t144 18.1208
R587 VSS.n228 VSS.t200 18.1208
R588 VSS.n938 VSS.t107 18.1208
R589 VSS.n325 VSS.t146 17.7063
R590 VSS.n337 VSS.t42 17.7063
R591 VSS.n678 VSS.t32 16.8265
R592 VSS.n123 VSS.t324 16.7654
R593 VSS.n77 VSS.t38 16.7654
R594 VSS.n310 VSS.t69 16.7227
R595 VSS.t81 VSS.t112 15.5322
R596 VSS.t187 VSS.t111 15.5322
R597 VSS.t20 VSS.t90 15.5322
R598 VSS.n637 VSS.t18 15.5322
R599 VSS.t203 VSS.t80 15.5322
R600 VSS.t191 VSS.t196 15.5322
R601 VSS.n226 VSS.t186 15.5322
R602 VSS.n1221 VSS.t64 15.5322
R603 VSS.n1000 VSS.t225 14.7111
R604 VSS.n966 VSS.t31 14.5955
R605 VSS.n1000 VSS.t120 14.4262
R606 VSS.n1000 VSS.t160 14.4262
R607 VSS.n124 VSS.t83 14.3704
R608 VSS.n646 VSS.t19 13.5907
R609 VSS.n660 VSS.t129 13.5907
R610 VSS.n241 VSS.n240 13.5907
R611 VSS.t97 VSS.t52 13.1729
R612 VSS.t261 VSS.t283 13.1729
R613 VSS.t54 VSS.t37 13.1729
R614 VSS.t131 VSS.t124 13.1729
R615 VSS.t293 VSS.t273 13.1729
R616 VSS.n1131 VSS.t203 12.9436
R617 VSS.n244 VSS.t138 12.2964
R618 VSS.n1311 VSS.t162 11.9754
R619 VSS.n1320 VSS.t151 11.9754
R620 VSS.n316 VSS.t219 11.8044
R621 VSS.n328 VSS.t315 11.8044
R622 VSS.n352 VSS.t67 11.8044
R623 VSS.t89 VSS.t117 11.0021
R624 VSS.n653 VSS.t41 11.0021
R625 VSS.n1243 VSS.t28 11.0021
R626 VSS.n304 VSS.t220 10.8207
R627 VSS.n656 VSS.t143 10.8207
R628 VSS.n1292 VSS.t296 10.778
R629 VSS.n1142 VSS.t191 10.3549
R630 VSS.t328 VSS.t92 9.83706
R631 VSS.t210 VSS.t110 9.83706
R632 VSS.t42 VSS.t43 9.83706
R633 VSS.t216 VSS.t180 9.83706
R634 VSS.t228 VSS.t159 9.83706
R635 VSS.n349 VSS.t182 9.83706
R636 VSS.n258 VSS.t136 9.70779
R637 VSS.n102 VSS.t100 9.58046
R638 VSS.n939 VSS.t313 9.48597
R639 VSS.n943 VSS.t279 9.48597
R640 VSS.n947 VSS.t218 9.48597
R641 VSS.n1006 VSS.t311 9.33385
R642 VSS.n871 VSS.t222 9.33385
R643 VSS.n1017 VSS.t334 9.33385
R644 VSS.n882 VSS.n881 9.32914
R645 VSS.n942 VSS.n941 9.32914
R646 VSS.n946 VSS.n945 9.32914
R647 VSS.n1004 VSS.n878 9.32914
R648 VSS.n1008 VSS.n872 9.32914
R649 VSS.n1015 VSS.n869 9.32914
R650 VSS.n619 VSS.t187 9.06064
R651 VSS.n622 VSS.t109 9.06064
R652 VSS.n631 VSS.t20 9.06064
R653 VSS.n216 VSS.t201 9.06064
R654 VSS.n1001 VSS.t121 8.96939
R655 VSS.n888 VSS.t226 8.96939
R656 VSS.n889 VSS.t161 8.96939
R657 VSS.n1003 VSS.t323 8.96939
R658 VSS.n1007 VSS.t224 8.96939
R659 VSS.n870 VSS.t317 8.96939
R660 VSS.n934 VSS.n933 8.41348
R661 VSS.n1294 VSS.t125 8.38296
R662 VSS.n34 VSS.t97 8.38296
R663 VSS.n672 VSS.t34 7.76633
R664 VSS.n208 VSS.n207 7.76633
R665 VSS.n1348 VSS.t170 7.64137
R666 VSS.n1313 VSS.t85 7.18547
R667 VSS.n54 VSS.t175 7.18547
R668 VSS.n1322 VSS.t149 7.18547
R669 VSS.n64 VSS.t299 7.18547
R670 VSS.n1197 VSS.t10 7.11918
R671 VSS.n893 VSS.n892 7.09117
R672 VSS.n301 VSS.t314 6.88609
R673 VSS.n27 VSS.n26 6.51634
R674 VSS.n669 VSS.t17 6.47203
R675 VSS.n896 VSS.t193 6.41395
R676 VSS.n1327 VSS.t88 6.41267
R677 VSS.n1291 VSS.n98 6.41267
R678 VSS.n1307 VSS.t274 6.41267
R679 VSS.n1310 VSS.n95 6.41267
R680 VSS.n1328 VSS.n92 6.41267
R681 VSS.n1347 VSS.t277 6.41267
R682 VSS.n893 VSS.t214 6.26682
R683 VSS.n873 VSS.t223 6.09694
R684 VSS.n879 VSS.t322 6.09694
R685 VSS.n1014 VSS.t316 6.09694
R686 VSS.t143 VSS.t230 5.90244
R687 VSS.n346 VSS.t139 5.90244
R688 VSS.n1287 VSS.n205 5.89743
R689 VSS.n920 VSS.n919 5.8805
R690 VSS.n922 VSS.n921 5.8805
R691 VSS.n894 VSS.n891 5.8805
R692 VSS.n895 VSS.n890 5.8805
R693 VSS.n896 VSS.t63 5.8805
R694 VSS.n213 VSS.n212 5.82487
R695 VSS.n1228 VSS.t105 5.82487
R696 VSS.n954 VSS.t213 5.35691
R697 VSS.n940 VSS.n939 5.2005
R698 VSS.n944 VSS.n943 5.2005
R699 VSS.n1005 VSS.n877 5.2005
R700 VSS.n1010 VSS.n1009 5.2005
R701 VSS.n1016 VSS.n868 5.2005
R702 VSS.n948 VSS.n947 5.2005
R703 VSS.n906 VSS.n905 5.2005
R704 VSS.n29 VSS.n28 5.2005
R705 VSS.n32 VSS.n31 5.2005
R706 VSS.n35 VSS.n34 5.2005
R707 VSS.n37 VSS.n36 5.2005
R708 VSS.n39 VSS.n38 5.2005
R709 VSS.n42 VSS.n41 5.2005
R710 VSS.n45 VSS.n44 5.2005
R711 VSS.n47 VSS.n46 5.2005
R712 VSS.n50 VSS.n49 5.2005
R713 VSS.n52 VSS.n51 5.2005
R714 VSS.n55 VSS.n54 5.2005
R715 VSS.n57 VSS.n56 5.2005
R716 VSS.n60 VSS.n59 5.2005
R717 VSS.n62 VSS.n61 5.2005
R718 VSS.n65 VSS.n64 5.2005
R719 VSS.n67 VSS.n66 5.2005
R720 VSS.n70 VSS.n69 5.2005
R721 VSS.n73 VSS.n72 5.2005
R722 VSS.n76 VSS.n75 5.2005
R723 VSS.n78 VSS.n77 5.2005
R724 VSS.n81 VSS.n80 5.2005
R725 VSS.n83 VSS.n82 5.2005
R726 VSS.n86 VSS.n85 5.2005
R727 VSS.n89 VSS.n88 5.2005
R728 VSS.n1293 VSS.n1292 5.2005
R729 VSS.n1295 VSS.n1294 5.2005
R730 VSS.n1297 VSS.n1296 5.2005
R731 VSS.n1299 VSS.n1298 5.2005
R732 VSS.n1302 VSS.n1301 5.2005
R733 VSS.n1304 VSS.n1303 5.2005
R734 VSS.n1306 VSS.n1305 5.2005
R735 VSS.n1309 VSS.n1308 5.2005
R736 VSS.n1312 VSS.n1311 5.2005
R737 VSS.n1314 VSS.n1313 5.2005
R738 VSS.n1316 VSS.n1315 5.2005
R739 VSS.n1318 VSS.n1317 5.2005
R740 VSS.n1321 VSS.n1320 5.2005
R741 VSS.n1323 VSS.n1322 5.2005
R742 VSS.n1325 VSS.n1324 5.2005
R743 VSS.n1327 VSS.n1326 5.2005
R744 VSS.n1330 VSS.n1329 5.2005
R745 VSS.n1332 VSS.n1331 5.2005
R746 VSS.n1334 VSS.n1333 5.2005
R747 VSS.n1337 VSS.n1336 5.2005
R748 VSS.n1340 VSS.n1339 5.2005
R749 VSS.n1342 VSS.n1341 5.2005
R750 VSS.n1344 VSS.n1343 5.2005
R751 VSS.n1346 VSS.n1345 5.2005
R752 VSS.n197 VSS.n99 5.2005
R753 VSS.n196 VSS.n100 5.2005
R754 VSS.n195 VSS.n101 5.2005
R755 VSS.n184 VSS.n102 5.2005
R756 VSS.n182 VSS.n105 5.2005
R757 VSS.n181 VSS.n106 5.2005
R758 VSS.n180 VSS.n107 5.2005
R759 VSS.n179 VSS.n108 5.2005
R760 VSS.n177 VSS.n111 5.2005
R761 VSS.n176 VSS.n112 5.2005
R762 VSS.n175 VSS.n113 5.2005
R763 VSS.n173 VSS.n116 5.2005
R764 VSS.n172 VSS.n117 5.2005
R765 VSS.n171 VSS.n118 5.2005
R766 VSS.n170 VSS.n119 5.2005
R767 VSS.n168 VSS.n122 5.2005
R768 VSS.n167 VSS.n123 5.2005
R769 VSS.n166 VSS.n124 5.2005
R770 VSS.n164 VSS.n127 5.2005
R771 VSS.n163 VSS.t134 5.2005
R772 VSS.n162 VSS.n128 5.2005
R773 VSS.n159 VSS.n131 5.2005
R774 VSS.n157 VSS.n132 5.2005
R775 VSS.n155 VSS.n135 5.2005
R776 VSS.n154 VSS.n136 5.2005
R777 VSS.n153 VSS.n137 5.2005
R778 VSS.n152 VSS.n138 5.2005
R779 VSS.n150 VSS.n141 5.2005
R780 VSS.n149 VSS.n142 5.2005
R781 VSS.n189 VSS.n187 5.2005
R782 VSS.n148 VSS.n143 5.2005
R783 VSS.n983 VSS.n982 5.2005
R784 VSS.n981 VSS.n980 5.2005
R785 VSS.n145 VSS.n144 5.2005
R786 VSS.n985 VSS.n979 5.2005
R787 VSS.n986 VSS.n977 5.2005
R788 VSS.n987 VSS.n976 5.2005
R789 VSS.n988 VSS.n975 5.2005
R790 VSS.n989 VSS.n974 5.2005
R791 VSS.n990 VSS.n973 5.2005
R792 VSS.n991 VSS.n972 5.2005
R793 VSS.n992 VSS.n971 5.2005
R794 VSS.n993 VSS.n970 5.2005
R795 VSS.n994 VSS.n969 5.2005
R796 VSS.n995 VSS.n968 5.2005
R797 VSS.n996 VSS.n967 5.2005
R798 VSS.n997 VSS.n966 5.2005
R799 VSS.n999 VSS.n998 5.2005
R800 VSS.n964 VSS.n963 5.2005
R801 VSS.n962 VSS.n961 5.2005
R802 VSS.n960 VSS.n959 5.2005
R803 VSS.n957 VSS.n956 5.2005
R804 VSS.n955 VSS.n954 5.2005
R805 VSS.n953 VSS.n952 5.2005
R806 VSS.n951 VSS.n950 5.2005
R807 VSS.n937 VSS.n936 5.2005
R808 VSS.n935 VSS.n934 5.2005
R809 VSS.n231 VSS.n230 5.2005
R810 VSS.n1276 VSS.n229 5.2005
R811 VSS.n1277 VSS.n228 5.2005
R812 VSS.n1278 VSS.n227 5.2005
R813 VSS.n1279 VSS.n226 5.2005
R814 VSS.n1280 VSS.n224 5.2005
R815 VSS.n1281 VSS.n219 5.2005
R816 VSS.n1282 VSS.n215 5.2005
R817 VSS.n1283 VSS.n213 5.2005
R818 VSS.n1284 VSS.n208 5.2005
R819 VSS.n116 VSS.t293 4.79048
R820 VSS.n137 VSS.t130 4.79048
R821 VSS.t41 VSS.n652 4.69176
R822 VSS.n640 VSS.t89 4.53057
R823 VSS.n219 VSS.n218 4.53057
R824 VSS.n189 VSS.n188 4.5005
R825 VSS.t159 VSS.t231 3.93512
R826 VSS.t67 VSS.t141 3.93512
R827 VSS.n741 VSS.t118 3.88342
R828 VSS.n224 VSS.n223 3.88342
R829 VSS.n916 VSS.n915 3.78833
R830 VSS.n204 VSS.n203 3.78833
R831 VSS.n84 VSS.n3 3.7355
R832 VSS.n74 VSS.n7 3.7355
R833 VSS.n63 VSS.n11 3.7355
R834 VSS.n53 VSS.n15 3.7355
R835 VSS.n43 VSS.n19 3.7355
R836 VSS.n33 VSS.n23 3.7355
R837 VSS.n901 VSS.n900 3.71473
R838 VSS.n30 VSS.n25 3.7042
R839 VSS.n40 VSS.n21 3.7042
R840 VSS.n48 VSS.n17 3.7042
R841 VSS.n58 VSS.n13 3.7042
R842 VSS.n68 VSS.n9 3.7042
R843 VSS.n79 VSS.n5 3.7042
R844 VSS.n87 VSS.n1 3.7042
R845 VSS.n1300 VSS.n97 3.68267
R846 VSS.n1319 VSS.n94 3.68267
R847 VSS.n1338 VSS.n91 3.68267
R848 VSS.n911 VSS.n910 3.67443
R849 VSS.n889 VSS.n880 3.65208
R850 VSS.n151 VSS.n140 3.64941
R851 VSS.n156 VSS.n134 3.64941
R852 VSS.n160 VSS.n130 3.64941
R853 VSS.n165 VSS.n126 3.64941
R854 VSS.n169 VSS.n121 3.64941
R855 VSS.n174 VSS.n115 3.64941
R856 VSS.n178 VSS.n110 3.64941
R857 VSS.n183 VSS.n104 3.64941
R858 VSS.n1003 VSS.n1002 3.64802
R859 VSS.n916 VSS.n913 3.1505
R860 VSS.n911 VSS.n908 3.1505
R861 VSS.n204 VSS.n201 3.1505
R862 VSS.n901 VSS.n898 3.1505
R863 VSS.n301 VSS.t280 2.95147
R864 VSS.n140 VSS.t276 2.7305
R865 VSS.n140 VSS.n139 2.7305
R866 VSS.n134 VSS.t168 2.7305
R867 VSS.n134 VSS.n133 2.7305
R868 VSS.n130 VSS.t303 2.7305
R869 VSS.n130 VSS.n129 2.7305
R870 VSS.n126 VSS.t336 2.7305
R871 VSS.n126 VSS.n125 2.7305
R872 VSS.n121 VSS.t263 2.7305
R873 VSS.n121 VSS.n120 2.7305
R874 VSS.n115 VSS.t286 2.7305
R875 VSS.n115 VSS.n114 2.7305
R876 VSS.n110 VSS.t53 2.7305
R877 VSS.n110 VSS.n109 2.7305
R878 VSS.n104 VSS.t101 2.7305
R879 VSS.n104 VSS.n103 2.7305
R880 VSS.n913 VSS.t1 2.7305
R881 VSS.n913 VSS.n912 2.7305
R882 VSS.n915 VSS.t206 2.7305
R883 VSS.n915 VSS.n914 2.7305
R884 VSS.n910 VSS.t156 2.7305
R885 VSS.n910 VSS.n909 2.7305
R886 VSS.n908 VSS.t192 2.7305
R887 VSS.n908 VSS.n907 2.7305
R888 VSS.n201 VSS.t209 2.7305
R889 VSS.n201 VSS.n200 2.7305
R890 VSS.n203 VSS.t236 2.7305
R891 VSS.n203 VSS.n202 2.7305
R892 VSS.n900 VSS.t207 2.7305
R893 VSS.n900 VSS.n899 2.7305
R894 VSS.n898 VSS.t6 2.7305
R895 VSS.n898 VSS.n897 2.7305
R896 VSS.n25 VSS.t103 2.7305
R897 VSS.n25 VSS.n24 2.7305
R898 VSS.n21 VSS.t258 2.7305
R899 VSS.n21 VSS.n20 2.7305
R900 VSS.n17 VSS.t292 2.7305
R901 VSS.n17 VSS.n16 2.7305
R902 VSS.n13 VSS.t335 2.7305
R903 VSS.n13 VSS.n12 2.7305
R904 VSS.n9 VSS.t266 2.7305
R905 VSS.n9 VSS.n8 2.7305
R906 VSS.n5 VSS.t255 2.7305
R907 VSS.n5 VSS.n4 2.7305
R908 VSS.n1 VSS.t307 2.7305
R909 VSS.n1 VSS.n0 2.7305
R910 VSS.n3 VSS.t58 2.7305
R911 VSS.n3 VSS.n2 2.7305
R912 VSS.n7 VSS.t309 2.7305
R913 VSS.n7 VSS.n6 2.7305
R914 VSS.n11 VSS.t84 2.7305
R915 VSS.n11 VSS.n10 2.7305
R916 VSS.n15 VSS.t86 2.7305
R917 VSS.n15 VSS.n14 2.7305
R918 VSS.n19 VSS.t272 2.7305
R919 VSS.n19 VSS.n18 2.7305
R920 VSS.n23 VSS.t268 2.7305
R921 VSS.n23 VSS.n22 2.7305
R922 VSS.n97 VSS.t262 2.7305
R923 VSS.n97 VSS.n96 2.7305
R924 VSS.n94 VSS.t179 2.7305
R925 VSS.n94 VSS.n93 2.7305
R926 VSS.n91 VSS.t248 2.7305
R927 VSS.n91 VSS.n90 2.7305
R928 VSS.n570 VSS.n569 2.63579
R929 VSS.n530 VSS.n458 2.6255
R930 VSS.n529 VSS.n460 2.60377
R931 VSS.n251 VSS.n248 2.60285
R932 VSS.n192 VSS.n191 2.60175
R933 VSS.n191 VSS.n190 2.601
R934 VSS.n412 VSS.n411 2.6005
R935 VSS.n410 VSS.n409 2.6005
R936 VSS.n403 VSS.n402 2.6005
R937 VSS.n401 VSS.n400 2.6005
R938 VSS.n398 VSS.n397 2.6005
R939 VSS.n396 VSS.n395 2.6005
R940 VSS.n393 VSS.n392 2.6005
R941 VSS.n391 VSS.n390 2.6005
R942 VSS.n388 VSS.n387 2.6005
R943 VSS.n386 VSS.n385 2.6005
R944 VSS.n383 VSS.n382 2.6005
R945 VSS.n381 VSS.n380 2.6005
R946 VSS.n378 VSS.n377 2.6005
R947 VSS.n376 VSS.n375 2.6005
R948 VSS.n374 VSS.n373 2.6005
R949 VSS.n372 VSS.n371 2.6005
R950 VSS.n370 VSS.n369 2.6005
R951 VSS.n368 VSS.n367 2.6005
R952 VSS.n366 VSS.n365 2.6005
R953 VSS.n536 VSS.n535 2.6005
R954 VSS.n535 VSS.n534 2.6005
R955 VSS.n533 VSS.n532 2.6005
R956 VSS.n532 VSS.n531 2.6005
R957 VSS.n297 VSS.n296 2.6005
R958 VSS.n296 VSS.n295 2.6005
R959 VSS.n300 VSS.n299 2.6005
R960 VSS.n299 VSS.n298 2.6005
R961 VSS.n303 VSS.n302 2.6005
R962 VSS.n302 VSS.n301 2.6005
R963 VSS.n306 VSS.n305 2.6005
R964 VSS.n305 VSS.n304 2.6005
R965 VSS.n309 VSS.n308 2.6005
R966 VSS.n308 VSS.n307 2.6005
R967 VSS.n312 VSS.n311 2.6005
R968 VSS.n311 VSS.n310 2.6005
R969 VSS.n315 VSS.n314 2.6005
R970 VSS.n314 VSS.n313 2.6005
R971 VSS.n318 VSS.n317 2.6005
R972 VSS.n317 VSS.n316 2.6005
R973 VSS.n321 VSS.n320 2.6005
R974 VSS.n320 VSS.n319 2.6005
R975 VSS.n324 VSS.n323 2.6005
R976 VSS.n323 VSS.n322 2.6005
R977 VSS.n327 VSS.n326 2.6005
R978 VSS.n326 VSS.n325 2.6005
R979 VSS.n330 VSS.n329 2.6005
R980 VSS.n329 VSS.n328 2.6005
R981 VSS.n333 VSS.n332 2.6005
R982 VSS.n332 VSS.n331 2.6005
R983 VSS.n336 VSS.n335 2.6005
R984 VSS.n335 VSS.n334 2.6005
R985 VSS.n339 VSS.n338 2.6005
R986 VSS.n338 VSS.n337 2.6005
R987 VSS.n342 VSS.n341 2.6005
R988 VSS.n341 VSS.n340 2.6005
R989 VSS.n345 VSS.n344 2.6005
R990 VSS.n344 VSS.n343 2.6005
R991 VSS.n348 VSS.n347 2.6005
R992 VSS.n347 VSS.n346 2.6005
R993 VSS.n351 VSS.n350 2.6005
R994 VSS.n350 VSS.n349 2.6005
R995 VSS.n354 VSS.n353 2.6005
R996 VSS.n353 VSS.n352 2.6005
R997 VSS.n357 VSS.n356 2.6005
R998 VSS.n356 VSS.n355 2.6005
R999 VSS.n360 VSS.n359 2.6005
R1000 VSS.n359 VSS.n358 2.6005
R1001 VSS.n364 VSS.n363 2.6005
R1002 VSS.n363 VSS.n362 2.6005
R1003 VSS.n538 VSS.n537 2.6005
R1004 VSS.n540 VSS.n539 2.6005
R1005 VSS.n542 VSS.n541 2.6005
R1006 VSS.n544 VSS.n543 2.6005
R1007 VSS.n546 VSS.n545 2.6005
R1008 VSS.n548 VSS.n547 2.6005
R1009 VSS.n550 VSS.n549 2.6005
R1010 VSS.n553 VSS.n552 2.6005
R1011 VSS.n555 VSS.n554 2.6005
R1012 VSS.n558 VSS.n557 2.6005
R1013 VSS.n560 VSS.n559 2.6005
R1014 VSS.n563 VSS.n562 2.6005
R1015 VSS.n565 VSS.n564 2.6005
R1016 VSS.n568 VSS.n567 2.6005
R1017 VSS.n571 VSS.n570 2.6005
R1018 VSS.n573 VSS.n572 2.6005
R1019 VSS.n576 VSS.n575 2.6005
R1020 VSS.n578 VSS.n577 2.6005
R1021 VSS.n585 VSS.n584 2.6005
R1022 VSS.n793 VSS.n792 2.6005
R1023 VSS.n796 VSS.n795 2.6005
R1024 VSS.n795 VSS.n794 2.6005
R1025 VSS.n799 VSS.n798 2.6005
R1026 VSS.n798 VSS.n797 2.6005
R1027 VSS.n802 VSS.n801 2.6005
R1028 VSS.n801 VSS.n800 2.6005
R1029 VSS.n805 VSS.n804 2.6005
R1030 VSS.n804 VSS.n803 2.6005
R1031 VSS.n808 VSS.n807 2.6005
R1032 VSS.n807 VSS.n806 2.6005
R1033 VSS.n811 VSS.n810 2.6005
R1034 VSS.n810 VSS.n809 2.6005
R1035 VSS.n814 VSS.n813 2.6005
R1036 VSS.n813 VSS.n812 2.6005
R1037 VSS.n817 VSS.n816 2.6005
R1038 VSS.n816 VSS.n815 2.6005
R1039 VSS.n820 VSS.n819 2.6005
R1040 VSS.n819 VSS.n818 2.6005
R1041 VSS.n823 VSS.n822 2.6005
R1042 VSS.n822 VSS.n821 2.6005
R1043 VSS.n826 VSS.n825 2.6005
R1044 VSS.n825 VSS.n824 2.6005
R1045 VSS.n829 VSS.n828 2.6005
R1046 VSS.n828 VSS.n827 2.6005
R1047 VSS.n832 VSS.n831 2.6005
R1048 VSS.n831 VSS.n830 2.6005
R1049 VSS.n835 VSS.n834 2.6005
R1050 VSS.n834 VSS.n833 2.6005
R1051 VSS.n838 VSS.n837 2.6005
R1052 VSS.n837 VSS.n836 2.6005
R1053 VSS.n841 VSS.n840 2.6005
R1054 VSS.n840 VSS.n839 2.6005
R1055 VSS.n844 VSS.n843 2.6005
R1056 VSS.n843 VSS.n842 2.6005
R1057 VSS.n847 VSS.n846 2.6005
R1058 VSS.n846 VSS.n845 2.6005
R1059 VSS.n850 VSS.n849 2.6005
R1060 VSS.n849 VSS.n848 2.6005
R1061 VSS.n853 VSS.n852 2.6005
R1062 VSS.n852 VSS.n851 2.6005
R1063 VSS.n856 VSS.n855 2.6005
R1064 VSS.n855 VSS.n854 2.6005
R1065 VSS.n859 VSS.n858 2.6005
R1066 VSS.n858 VSS.n857 2.6005
R1067 VSS.n764 VSS.n763 2.6005
R1068 VSS.n767 VSS.n766 2.6005
R1069 VSS.n769 VSS.n768 2.6005
R1070 VSS.n772 VSS.n771 2.6005
R1071 VSS.n774 VSS.n773 2.6005
R1072 VSS.n777 VSS.n776 2.6005
R1073 VSS.n779 VSS.n778 2.6005
R1074 VSS.n782 VSS.n781 2.6005
R1075 VSS.n784 VSS.n783 2.6005
R1076 VSS.n788 VSS.n787 2.6005
R1077 VSS.n862 VSS.n861 2.6005
R1078 VSS.n864 VSS.n863 2.6005
R1079 VSS.n867 VSS.n866 2.6005
R1080 VSS.n1021 VSS.n1020 2.6005
R1081 VSS.n1024 VSS.n1023 2.6005
R1082 VSS.n1027 VSS.n1026 2.6005
R1083 VSS.n1030 VSS.n1029 2.6005
R1084 VSS.n1033 VSS.n1032 2.6005
R1085 VSS.n1037 VSS.n1036 2.6005
R1086 VSS.n791 VSS.n790 2.6005
R1087 VSS.n790 VSS.n789 2.6005
R1088 VSS.n1264 VSS.n1263 2.6005
R1089 VSS.n1263 VSS.n1262 2.6005
R1090 VSS.n248 VSS.n247 2.6005
R1091 VSS.n1139 VSS.n1138 2.6005
R1092 VSS.n1138 VSS.n1137 2.6005
R1093 VSS.n212 VSS.n211 2.6005
R1094 VSS.n1144 VSS.n1143 2.6005
R1095 VSS.n1143 VSS.n1142 2.6005
R1096 VSS.n1238 VSS.n1237 2.6005
R1097 VSS.n1239 VSS.n1238 2.6005
R1098 VSS.n1236 VSS.n1235 2.6005
R1099 VSS.n1235 VSS.n1234 2.6005
R1100 VSS.n1233 VSS.n1232 2.6005
R1101 VSS.n1124 VSS.n1123 2.6005
R1102 VSS.n1123 VSS.n1122 2.6005
R1103 VSS.n233 VSS.n232 2.6005
R1104 VSS.n1146 VSS.n1145 2.6005
R1105 VSS.n1148 VSS.n1147 2.6005
R1106 VSS.n1150 VSS.n1149 2.6005
R1107 VSS.n1152 VSS.n1151 2.6005
R1108 VSS.n1154 VSS.n1153 2.6005
R1109 VSS.n1156 VSS.n1155 2.6005
R1110 VSS.n1158 VSS.n1157 2.6005
R1111 VSS.n1160 VSS.n1159 2.6005
R1112 VSS.n1162 VSS.n1161 2.6005
R1113 VSS.n1164 VSS.n1163 2.6005
R1114 VSS.n1166 VSS.n1165 2.6005
R1115 VSS.n1168 VSS.n1167 2.6005
R1116 VSS.n1170 VSS.n1169 2.6005
R1117 VSS.n1172 VSS.n1171 2.6005
R1118 VSS.n1174 VSS.n1173 2.6005
R1119 VSS.n1176 VSS.n1175 2.6005
R1120 VSS.n1178 VSS.n1177 2.6005
R1121 VSS.n1180 VSS.n1179 2.6005
R1122 VSS.n1182 VSS.n1181 2.6005
R1123 VSS.n1184 VSS.n1183 2.6005
R1124 VSS.n1186 VSS.n1185 2.6005
R1125 VSS.n1188 VSS.n1187 2.6005
R1126 VSS.n1193 VSS.n1192 2.6005
R1127 VSS.n235 VSS.n234 2.6005
R1128 VSS.n254 VSS.n253 2.6005
R1129 VSS.n253 VSS.n252 2.6005
R1130 VSS.n246 VSS.n245 2.6005
R1131 VSS.n245 VSS.n244 2.6005
R1132 VSS.n239 VSS.n238 2.6005
R1133 VSS.n238 VSS.n237 2.6005
R1134 VSS.n243 VSS.n242 2.6005
R1135 VSS.n242 VSS.n241 2.6005
R1136 VSS.n1267 VSS.n1266 2.6005
R1137 VSS.n1266 VSS.n1265 2.6005
R1138 VSS.n1270 VSS.n1269 2.6005
R1139 VSS.n1269 VSS.n1268 2.6005
R1140 VSS.n260 VSS.n259 2.6005
R1141 VSS.n259 VSS.n258 2.6005
R1142 VSS.n263 VSS.n262 2.6005
R1143 VSS.n262 VSS.n261 2.6005
R1144 VSS.n265 VSS.n264 2.6005
R1145 VSS.n267 VSS.n266 2.6005
R1146 VSS.n223 VSS.n222 2.6005
R1147 VSS.n257 VSS.n256 2.6005
R1148 VSS.n256 VSS.n255 2.6005
R1149 VSS.n270 VSS.n269 2.6005
R1150 VSS.n269 VSS.n268 2.6005
R1151 VSS.n210 VSS.n209 2.6005
R1152 VSS.n273 VSS.n272 2.6005
R1153 VSS.n1242 VSS.n1241 2.6005
R1154 VSS.n1241 VSS.n1240 2.6005
R1155 VSS.n1245 VSS.n1244 2.6005
R1156 VSS.n1244 VSS.n1243 2.6005
R1157 VSS.n218 VSS.n217 2.6005
R1158 VSS.n1248 VSS.n1247 2.6005
R1159 VSS.n1252 VSS.n1251 2.6005
R1160 VSS.n1251 VSS.n1250 2.6005
R1161 VSS.n1255 VSS.n1254 2.6005
R1162 VSS.n1254 VSS.n1253 2.6005
R1163 VSS.n1258 VSS.n1257 2.6005
R1164 VSS.n1257 VSS.n1256 2.6005
R1165 VSS.n1261 VSS.n1260 2.6005
R1166 VSS.n1260 VSS.n1259 2.6005
R1167 VSS.n250 VSS.n249 2.6005
R1168 VSS.n275 VSS.n274 2.6005
R1169 VSS.n277 VSS.n276 2.6005
R1170 VSS.n279 VSS.n278 2.6005
R1171 VSS.n281 VSS.n280 2.6005
R1172 VSS.n283 VSS.n282 2.6005
R1173 VSS.n285 VSS.n284 2.6005
R1174 VSS.n287 VSS.n286 2.6005
R1175 VSS.n290 VSS.n289 2.6005
R1176 VSS.n292 VSS.n291 2.6005
R1177 VSS.n294 VSS.n293 2.6005
R1178 VSS.n1077 VSS.n1076 2.6005
R1179 VSS.n1079 VSS.n1078 2.6005
R1180 VSS.n1081 VSS.n1080 2.6005
R1181 VSS.n1084 VSS.n1083 2.6005
R1182 VSS.n1086 VSS.n1085 2.6005
R1183 VSS.n1088 VSS.n1087 2.6005
R1184 VSS.n1092 VSS.n1091 2.6005
R1185 VSS.n1094 VSS.n1093 2.6005
R1186 VSS.n1096 VSS.n1095 2.6005
R1187 VSS.n1101 VSS.n1100 2.6005
R1188 VSS.n1104 VSS.n1103 2.6005
R1189 VSS.n1103 VSS.n1102 2.6005
R1190 VSS.n1106 VSS.n1105 2.6005
R1191 VSS.n1108 VSS.n1107 2.6005
R1192 VSS.n1115 VSS.n1114 2.6005
R1193 VSS.n1214 VSS.n1213 2.6005
R1194 VSS.n1213 VSS.n1212 2.6005
R1195 VSS.n1202 VSS.n1201 2.6005
R1196 VSS.n1201 VSS.n1200 2.6005
R1197 VSS.n1211 VSS.n1210 2.6005
R1198 VSS.n1210 VSS.n1209 2.6005
R1199 VSS.n1217 VSS.n1216 2.6005
R1200 VSS.n1216 VSS.n1215 2.6005
R1201 VSS.n1220 VSS.n1219 2.6005
R1202 VSS.n1219 VSS.n1218 2.6005
R1203 VSS.n1223 VSS.n1222 2.6005
R1204 VSS.n1222 VSS.n1221 2.6005
R1205 VSS.n1226 VSS.n1225 2.6005
R1206 VSS.n1225 VSS.n1224 2.6005
R1207 VSS.n221 VSS.n220 2.6005
R1208 VSS.n1231 VSS.n1230 2.6005
R1209 VSS.n1230 VSS.n1229 2.6005
R1210 VSS.n1118 VSS.n1117 2.6005
R1211 VSS.n1117 VSS.n1116 2.6005
R1212 VSS.n1121 VSS.n1120 2.6005
R1213 VSS.n1120 VSS.n1119 2.6005
R1214 VSS.n1127 VSS.n1126 2.6005
R1215 VSS.n1126 VSS.n1125 2.6005
R1216 VSS.n1130 VSS.n1129 2.6005
R1217 VSS.n1129 VSS.n1128 2.6005
R1218 VSS.n1134 VSS.n1133 2.6005
R1219 VSS.n1133 VSS.n1132 2.6005
R1220 VSS.n1136 VSS.n1135 2.6005
R1221 VSS.n1208 VSS.n1207 2.6005
R1222 VSS.n1207 VSS.n1206 2.6005
R1223 VSS.n1205 VSS.n1204 2.6005
R1224 VSS.n1204 VSS.n1203 2.6005
R1225 VSS.n1199 VSS.n1198 2.6005
R1226 VSS.n1198 VSS.n1197 2.6005
R1227 VSS.n1196 VSS.n1195 2.6005
R1228 VSS.n1195 VSS.n1194 2.6005
R1229 VSS.n732 VSS.n731 2.6005
R1230 VSS.n729 VSS.n728 2.6005
R1231 VSS.n726 VSS.n725 2.6005
R1232 VSS.n723 VSS.n722 2.6005
R1233 VSS.n720 VSS.n719 2.6005
R1234 VSS.n717 VSS.n716 2.6005
R1235 VSS.n714 VSS.n713 2.6005
R1236 VSS.n711 VSS.n710 2.6005
R1237 VSS.n708 VSS.n707 2.6005
R1238 VSS.n705 VSS.n704 2.6005
R1239 VSS.n702 VSS.n701 2.6005
R1240 VSS.n699 VSS.n698 2.6005
R1241 VSS.n696 VSS.n695 2.6005
R1242 VSS.n694 VSS.n693 2.6005
R1243 VSS.n692 VSS.n691 2.6005
R1244 VSS.n690 VSS.n689 2.6005
R1245 VSS.n688 VSS.n687 2.6005
R1246 VSS.n455 VSS.n454 2.6005
R1247 VSS.n454 VSS.n453 2.6005
R1248 VSS.n452 VSS.n451 2.6005
R1249 VSS.n451 VSS.n450 2.6005
R1250 VSS.n449 VSS.n448 2.6005
R1251 VSS.n448 VSS.n447 2.6005
R1252 VSS.n445 VSS.n444 2.6005
R1253 VSS.n444 VSS.n443 2.6005
R1254 VSS.n442 VSS.n441 2.6005
R1255 VSS.n441 VSS.n440 2.6005
R1256 VSS.n439 VSS.n438 2.6005
R1257 VSS.n435 VSS.n434 2.6005
R1258 VSS.n432 VSS.n431 2.6005
R1259 VSS.n429 VSS.n428 2.6005
R1260 VSS.n426 VSS.n425 2.6005
R1261 VSS.n423 VSS.n422 2.6005
R1262 VSS.n420 VSS.n419 2.6005
R1263 VSS.n417 VSS.n416 2.6005
R1264 VSS.n415 VSS.n414 2.6005
R1265 VSS.n588 VSS.n587 2.6005
R1266 VSS.n590 VSS.n589 2.6005
R1267 VSS.n593 VSS.n592 2.6005
R1268 VSS.n595 VSS.n594 2.6005
R1269 VSS.n598 VSS.n597 2.6005
R1270 VSS.n600 VSS.n599 2.6005
R1271 VSS.n603 VSS.n602 2.6005
R1272 VSS.n605 VSS.n604 2.6005
R1273 VSS.n609 VSS.n608 2.6005
R1274 VSS.n685 VSS.n684 2.6005
R1275 VSS.n684 VSS.n683 2.6005
R1276 VSS.n680 VSS.n679 2.6005
R1277 VSS.n679 VSS.n678 2.6005
R1278 VSS.n677 VSS.n676 2.6005
R1279 VSS.n676 VSS.n675 2.6005
R1280 VSS.n674 VSS.n673 2.6005
R1281 VSS.n673 VSS.n672 2.6005
R1282 VSS.n671 VSS.n670 2.6005
R1283 VSS.n670 VSS.n669 2.6005
R1284 VSS.n668 VSS.n667 2.6005
R1285 VSS.n667 VSS.n666 2.6005
R1286 VSS.n665 VSS.n664 2.6005
R1287 VSS.n664 VSS.n663 2.6005
R1288 VSS.n662 VSS.n661 2.6005
R1289 VSS.n661 VSS.n660 2.6005
R1290 VSS.n659 VSS.n658 2.6005
R1291 VSS.n658 VSS.n657 2.6005
R1292 VSS.n655 VSS.n654 2.6005
R1293 VSS.n654 VSS.n653 2.6005
R1294 VSS.n651 VSS.n650 2.6005
R1295 VSS.n650 VSS.n649 2.6005
R1296 VSS.n648 VSS.n647 2.6005
R1297 VSS.n647 VSS.n646 2.6005
R1298 VSS.n645 VSS.n644 2.6005
R1299 VSS.n644 VSS.n643 2.6005
R1300 VSS.n642 VSS.n641 2.6005
R1301 VSS.n641 VSS.n640 2.6005
R1302 VSS.n639 VSS.n638 2.6005
R1303 VSS.n638 VSS.n637 2.6005
R1304 VSS.n636 VSS.n635 2.6005
R1305 VSS.n635 VSS.n634 2.6005
R1306 VSS.n633 VSS.n632 2.6005
R1307 VSS.n632 VSS.n631 2.6005
R1308 VSS.n630 VSS.n629 2.6005
R1309 VSS.n629 VSS.n628 2.6005
R1310 VSS.n627 VSS.n626 2.6005
R1311 VSS.n626 VSS.n625 2.6005
R1312 VSS.n624 VSS.n623 2.6005
R1313 VSS.n623 VSS.n622 2.6005
R1314 VSS.n621 VSS.n620 2.6005
R1315 VSS.n620 VSS.n619 2.6005
R1316 VSS.n618 VSS.n617 2.6005
R1317 VSS.n617 VSS.n616 2.6005
R1318 VSS.n615 VSS.n614 2.6005
R1319 VSS.n614 VSS.t81 2.6005
R1320 VSS.n613 VSS.n612 2.6005
R1321 VSS.n612 VSS.n611 2.6005
R1322 VSS.n458 VSS.n457 2.6005
R1323 VSS.n528 VSS.n527 2.6005
R1324 VSS.n526 VSS.n525 2.6005
R1325 VSS.n512 VSS.n511 2.6005
R1326 VSS.n510 VSS.n509 2.6005
R1327 VSS.n507 VSS.n506 2.6005
R1328 VSS.n504 VSS.n503 2.6005
R1329 VSS.n502 VSS.n501 2.6005
R1330 VSS.n499 VSS.n498 2.6005
R1331 VSS.n497 VSS.n496 2.6005
R1332 VSS.n494 VSS.n493 2.6005
R1333 VSS.n492 VSS.n491 2.6005
R1334 VSS.n489 VSS.n488 2.6005
R1335 VSS.n487 VSS.n486 2.6005
R1336 VSS.n484 VSS.n483 2.6005
R1337 VSS.n482 VSS.n481 2.6005
R1338 VSS.n480 VSS.n479 2.6005
R1339 VSS.n478 VSS.n477 2.6005
R1340 VSS.n476 VSS.n475 2.6005
R1341 VSS.n474 VSS.n473 2.6005
R1342 VSS.n472 VSS.n471 2.6005
R1343 VSS.n470 VSS.n469 2.6005
R1344 VSS.n468 VSS.n467 2.6005
R1345 VSS.n466 VSS.n465 2.6005
R1346 VSS.n464 VSS.n463 2.6005
R1347 VSS.n462 VSS.n461 2.6005
R1348 VSS.n746 VSS.n745 2.6005
R1349 VSS.n748 VSS.n747 2.6005
R1350 VSS.n750 VSS.n749 2.6005
R1351 VSS.n752 VSS.n751 2.6005
R1352 VSS.n754 VSS.n753 2.6005
R1353 VSS.n756 VSS.n755 2.6005
R1354 VSS.n758 VSS.n757 2.6005
R1355 VSS.n760 VSS.n759 2.6005
R1356 VSS.n762 VSS.n761 2.6005
R1357 VSS.n734 VSS.n733 2.6005
R1358 VSS.n1039 VSS.n1038 2.6005
R1359 VSS.n1041 VSS.n1040 2.6005
R1360 VSS.n1043 VSS.n1042 2.6005
R1361 VSS.n1045 VSS.n1044 2.6005
R1362 VSS.n1047 VSS.n1046 2.6005
R1363 VSS.n1050 VSS.n1049 2.6005
R1364 VSS.n1052 VSS.n1051 2.6005
R1365 VSS.n1055 VSS.n1054 2.6005
R1366 VSS.n1057 VSS.n1056 2.6005
R1367 VSS.n1060 VSS.n1059 2.6005
R1368 VSS.n1062 VSS.n1061 2.6005
R1369 VSS.n1065 VSS.n1064 2.6005
R1370 VSS.n1067 VSS.n1066 2.6005
R1371 VSS.n1070 VSS.n1069 2.6005
R1372 VSS.n1072 VSS.n1071 2.6005
R1373 VSS.n744 VSS.n743 2.6005
R1374 VSS.n1274 VSS.n1273 2.6005
R1375 VSS.n1273 VSS.n1272 2.6005
R1376 VSS.n450 VSS.t140 2.58911
R1377 VSS.n1002 VSS.n1001 2.50665
R1378 VSS.n888 VSS.n880 2.50664
R1379 VSS.n1292 VSS.t102 2.39549
R1380 VSS.n31 VSS.t36 2.39549
R1381 VSS.n72 VSS.n71 2.39549
R1382 VSS.n1331 VSS.t308 2.39549
R1383 VSS.n75 VSS.t251 2.39549
R1384 VSS.n1336 VSS.n1335 2.39549
R1385 VSS.n419 VSS.n418 2.33733
R1386 VSS.n422 VSS.n421 2.33733
R1387 VSS.n425 VSS.n424 2.33733
R1388 VSS.n428 VSS.n427 2.33733
R1389 VSS.n431 VSS.n430 2.33733
R1390 VSS.n434 VSS.n433 2.33733
R1391 VSS.n698 VSS.n697 2.31748
R1392 VSS.n701 VSS.n700 2.31748
R1393 VSS.n704 VSS.n703 2.31748
R1394 VSS.n707 VSS.n706 2.31748
R1395 VSS.n710 VSS.n709 2.31748
R1396 VSS.n713 VSS.n712 2.31748
R1397 VSS.n716 VSS.n715 2.31748
R1398 VSS.n719 VSS.n718 2.31748
R1399 VSS.n722 VSS.n721 2.31748
R1400 VSS.n725 VSS.n724 2.31748
R1401 VSS.n728 VSS.n727 2.31748
R1402 VSS.n1032 VSS.n1031 2.31748
R1403 VSS.n1029 VSS.n1028 2.31748
R1404 VSS.n1026 VSS.n1025 2.31748
R1405 VSS.n1023 VSS.n1022 2.31748
R1406 VSS.n1020 VSS.n1019 2.31748
R1407 VSS.n866 VSS.n865 2.31748
R1408 VSS.n189 VSS.n186 2.15773
R1409 VSS.n875 VSS.n873 2.1063
R1410 VSS.n1014 VSS.n1013 2.1063
R1411 VSS.n1000 VSS.n879 2.1063
R1412 VSS.t24 VSS.t23 1.96781
R1413 VSS.t44 VSS.t25 1.96781
R1414 VSS.n1132 VSS.n1131 1.94196
R1415 VSS.n207 VSS.n206 1.94196
R1416 VSS.n212 VSS.n210 1.94196
R1417 VSS.n1142 VSS.n1141 1.94196
R1418 VSS.n1240 VSS.n1239 1.94196
R1419 VSS.n218 VSS.n216 1.94196
R1420 VSS.n1229 VSS.n1228 1.94196
R1421 VSS.n223 VSS.n221 1.94196
R1422 VSS.n1206 VSS.t29 1.94196
R1423 VSS.n448 VSS.n446 1.7198
R1424 VSS.n552 VSS.n551 1.70459
R1425 VSS.n557 VSS.n556 1.70459
R1426 VSS.n562 VSS.n561 1.70459
R1427 VSS.n567 VSS.n566 1.70459
R1428 VSS.n575 VSS.n574 1.70459
R1429 VSS.n584 VSS.n583 1.70459
R1430 VSS.n597 VSS.n596 1.70459
R1431 VSS.n602 VSS.n601 1.70459
R1432 VSS.n608 VSS.n607 1.70459
R1433 VSS.n409 VSS.n408 1.61305
R1434 VSS.n400 VSS.n399 1.61305
R1435 VSS.n395 VSS.n394 1.61305
R1436 VSS.n390 VSS.n389 1.61305
R1437 VSS.n385 VSS.n384 1.61305
R1438 VSS.n380 VSS.n379 1.61305
R1439 VSS.n289 VSS.n288 1.61162
R1440 VSS.n1076 VSS.n1075 1.61162
R1441 VSS.n1083 VSS.n1082 1.61162
R1442 VSS.n1091 VSS.n1090 1.61162
R1443 VSS.n1100 VSS.n1099 1.61162
R1444 VSS.n1114 VSS.n1113 1.61162
R1445 VSS.n766 VSS.n765 1.60368
R1446 VSS.n771 VSS.n770 1.60357
R1447 VSS.n776 VSS.n775 1.60357
R1448 VSS.n781 VSS.n780 1.60357
R1449 VSS.n787 VSS.n786 1.60357
R1450 VSS.n506 VSS.n505 1.60357
R1451 VSS.n501 VSS.n500 1.60357
R1452 VSS.n496 VSS.n495 1.60357
R1453 VSS.n491 VSS.n490 1.60357
R1454 VSS.n486 VSS.n485 1.60357
R1455 VSS.n1049 VSS.n1048 1.60357
R1456 VSS.n1054 VSS.n1053 1.60357
R1457 VSS.n1059 VSS.n1058 1.60357
R1458 VSS.n1064 VSS.n1063 1.60357
R1459 VSS.n1069 VSS.n1068 1.60357
R1460 VSS.n743 VSS.n742 1.60357
R1461 VSS.n460 VSS.n459 1.58772
R1462 VSS.n1192 VSS.n1191 1.55656
R1463 VSS.n1018 VSS.n1017 1.49543
R1464 VSS.n587 VSS.n586 1.45409
R1465 VSS.n592 VSS.n591 1.45409
R1466 VSS.n741 VSS.n737 1.44276
R1467 VSS.n741 VSS.n738 1.44276
R1468 VSS.n741 VSS.n739 1.44276
R1469 VSS.n1348 VSS.n1347 1.43392
R1470 VSS.n684 VSS.n682 1.38322
R1471 VSS.n414 VSS.n413 1.35581
R1472 VSS.n438 VSS.n437 1.35567
R1473 VSS.n1036 VSS.n1035 1.34579
R1474 VSS.n525 VSS.n524 1.34565
R1475 VSS.n509 VSS.n508 1.34565
R1476 VSS.n731 VSS.n730 1.34565
R1477 VSS.n861 VSS.n860 1.34565
R1478 VSS.n1291 VSS.n1290 1.34093
R1479 VSS.n224 VSS.t202 1.29481
R1480 VSS.n227 VSS.t190 1.29481
R1481 VSS.n1215 VSS.t119 1.29481
R1482 VSS.n682 VSS.n681 1.28007
R1483 VSS.n1286 VSS.n1285 1.22876
R1484 VSS.n1002 VSS.n880 1.11085
R1485 VSS.t79 VSS.t147 0.984156
R1486 VSS.t220 VSS.t33 0.984156
R1487 VSS.t267 VSS.t229 0.984156
R1488 VSS.t219 VSS.t287 0.984156
R1489 VSS.t215 VSS.t27 0.984156
R1490 VSS.n917 VSS.n916 0.96262
R1491 VSS.n1035 VSS.n1034 0.838098
R1492 VSS.n741 VSS.n740 0.838098
R1493 VSS.n524 VSS.n523 0.837901
R1494 VSS.n437 VSS.n436 0.83122
R1495 VSS.n965 VSS.n922 0.7259
R1496 VSS.n1007 VSS.n1006 0.702093
R1497 VSS.n871 VSS.n870 0.687093
R1498 VSS.n984 VSS.n983 0.673934
R1499 VSS.n29 VSS.n27 0.661796
R1500 VSS.t227 VSS.t39 0.647653
R1501 VSS.n649 VSS.t35 0.647653
R1502 VSS.n1112 VSS.n1109 0.647653
R1503 VSS.n1112 VSS.n1111 0.647653
R1504 VSS.n1098 VSS.n1097 0.647653
R1505 VSS.n1239 VSS.n215 0.647653
R1506 VSS.n1190 VSS.n1189 0.647653
R1507 VSS.n928 VSS.n925 0.647653
R1508 VSS.n931 VSS.n928 0.647653
R1509 VSS.n932 VSS.n931 0.647653
R1510 VSS.n933 VSS.n932 0.647653
R1511 VSS.n148 VSS.n147 0.644436
R1512 VSS.n1074 VSS.n1073 0.619447
R1513 VSS.n147 VSS.n145 0.609948
R1514 VSS.n922 VSS.n920 0.5873
R1515 VSS.n199 VSS.n197 0.569951
R1516 VSS.n928 VSS.n927 0.523462
R1517 VSS.n928 VSS.n926 0.523462
R1518 VSS.n925 VSS.n923 0.523222
R1519 VSS.n931 VSS.n930 0.523222
R1520 VSS.n931 VSS.n929 0.523222
R1521 VSS.n1191 VSS.n1190 0.523222
R1522 VSS.n895 VSS.n894 0.506362
R1523 VSS.n786 VSS.n785 0.499715
R1524 VSS.n523 VSS.n522 0.499715
R1525 VSS.n523 VSS.n521 0.499715
R1526 VSS.n523 VSS.n520 0.499715
R1527 VSS.n523 VSS.n519 0.499715
R1528 VSS.n523 VSS.n518 0.499715
R1529 VSS.n523 VSS.n517 0.499715
R1530 VSS.n523 VSS.n516 0.499715
R1531 VSS.n523 VSS.n515 0.499715
R1532 VSS.n523 VSS.n514 0.499715
R1533 VSS.n523 VSS.n513 0.499715
R1534 VSS.n741 VSS.n735 0.499715
R1535 VSS.n741 VSS.n736 0.499715
R1536 VSS.n742 VSS.n741 0.499715
R1537 VSS.n1090 VSS.n1089 0.49569
R1538 VSS.n1099 VSS.n1098 0.49569
R1539 VSS.n1113 VSS.n1112 0.49569
R1540 VSS.n408 VSS.n407 0.494977
R1541 VSS.n407 VSS.n406 0.494977
R1542 VSS.n407 VSS.n405 0.494977
R1543 VSS.n407 VSS.n404 0.494977
R1544 VSS.n205 VSS.n204 0.491587
R1545 VSS.n925 VSS.n924 0.466933
R1546 VSS.n903 VSS.n902 0.4638
R1547 VSS.n918 VSS.n917 0.46349
R1548 VSS.n920 VSS.n918 0.4559
R1549 VSS VSS.n882 0.451296
R1550 VSS.n942 VSS 0.451296
R1551 VSS.n946 VSS 0.451296
R1552 VSS.n1004 VSS 0.451296
R1553 VSS.n1008 VSS 0.451296
R1554 VSS.n1015 VSS 0.451296
R1555 VSS.n582 VSS.n581 0.449449
R1556 VSS.n582 VSS.n580 0.449206
R1557 VSS.n582 VSS.n579 0.449206
R1558 VSS.n583 VSS.n582 0.449206
R1559 VSS.n607 VSS.n606 0.449206
R1560 VSS.n1111 VSS.n1110 0.440691
R1561 VSS.n902 VSS.n901 0.438385
R1562 VSS.n199 VSS.n198 0.432926
R1563 VSS.n191 VSS.n189 0.426383
R1564 VSS.n363 VSS.n361 0.424742
R1565 VSS.n1290 VSS.n199 0.421958
R1566 VSS.n903 VSS.n896 0.4145
R1567 VSS.n917 VSS.n911 0.407107
R1568 VSS.n1286 VSS.n1284 0.406886
R1569 VSS.n904 VSS.n895 0.393086
R1570 VSS.n918 VSS.n906 0.36591
R1571 VSS.n791 VSS.n788 0.358535
R1572 VSS.n1289 VSS.n1288 0.300993
R1573 VSS.n1287 VSS.n1286 0.296642
R1574 VSS.n1275 VSS 0.244029
R1575 VSS.n149 VSS.n148 0.242079
R1576 VSS.n1290 VSS.n1289 0.236806
R1577 VSS.n894 VSS.n893 0.230155
R1578 VSS.n904 VSS.n903 0.225254
R1579 VSS VSS.n1274 0.210752
R1580 VSS VSS.n1348 0.183461
R1581 VSS.n985 VSS.n984 0.177572
R1582 VSS.n862 VSS.n859 0.166798
R1583 VSS.n688 VSS.n686 0.1605
R1584 VSS.n530 VSS.n529 0.159151
R1585 VSS.n1006 VSS.n1005 0.152624
R1586 VSS.n1009 VSS.n871 0.152624
R1587 VSS.n1017 VSS.n1016 0.152624
R1588 VSS VSS.n882 0.139881
R1589 VSS VSS.n942 0.139881
R1590 VSS VSS.n946 0.139881
R1591 VSS VSS.n1004 0.139881
R1592 VSS VSS.n1008 0.139881
R1593 VSS VSS.n1015 0.139881
R1594 VSS.n615 VSS.n613 0.127128
R1595 VSS.n618 VSS.n615 0.127128
R1596 VSS.n621 VSS.n618 0.127128
R1597 VSS.n624 VSS.n621 0.127128
R1598 VSS.n627 VSS.n624 0.127128
R1599 VSS.n630 VSS.n627 0.127128
R1600 VSS.n633 VSS.n630 0.127128
R1601 VSS.n636 VSS.n633 0.127128
R1602 VSS.n639 VSS.n636 0.127128
R1603 VSS.n642 VSS.n639 0.127128
R1604 VSS.n645 VSS.n642 0.127128
R1605 VSS.n648 VSS.n645 0.127128
R1606 VSS.n651 VSS.n648 0.127128
R1607 VSS.n655 VSS.n651 0.127128
R1608 VSS.n659 VSS.n655 0.127128
R1609 VSS.n662 VSS.n659 0.127128
R1610 VSS.n665 VSS.n662 0.127128
R1611 VSS.n668 VSS.n665 0.127128
R1612 VSS.n671 VSS.n668 0.127128
R1613 VSS.n674 VSS.n671 0.127128
R1614 VSS.n677 VSS.n674 0.127128
R1615 VSS.n680 VSS.n677 0.127128
R1616 VSS.n685 VSS.n680 0.127128
R1617 VSS.n793 VSS.n791 0.127128
R1618 VSS.n796 VSS.n793 0.127128
R1619 VSS.n799 VSS.n796 0.127128
R1620 VSS.n802 VSS.n799 0.127128
R1621 VSS.n805 VSS.n802 0.127128
R1622 VSS.n808 VSS.n805 0.127128
R1623 VSS.n811 VSS.n808 0.127128
R1624 VSS.n814 VSS.n811 0.127128
R1625 VSS.n817 VSS.n814 0.127128
R1626 VSS.n820 VSS.n817 0.127128
R1627 VSS.n823 VSS.n820 0.127128
R1628 VSS.n826 VSS.n823 0.127128
R1629 VSS.n829 VSS.n826 0.127128
R1630 VSS.n832 VSS.n829 0.127128
R1631 VSS.n835 VSS.n832 0.127128
R1632 VSS.n838 VSS.n835 0.127128
R1633 VSS.n841 VSS.n838 0.127128
R1634 VSS.n844 VSS.n841 0.127128
R1635 VSS.n847 VSS.n844 0.127128
R1636 VSS.n850 VSS.n847 0.127128
R1637 VSS.n853 VSS.n850 0.127128
R1638 VSS.n856 VSS.n853 0.127128
R1639 VSS.n859 VSS.n856 0.127128
R1640 VSS.n197 VSS.n196 0.121553
R1641 VSS.n196 VSS.n195 0.121553
R1642 VSS.n182 VSS.n181 0.121553
R1643 VSS.n181 VSS.n180 0.121553
R1644 VSS.n180 VSS.n179 0.121553
R1645 VSS.n177 VSS.n176 0.121553
R1646 VSS.n176 VSS.n175 0.121553
R1647 VSS.n173 VSS.n172 0.121553
R1648 VSS.n172 VSS.n171 0.121553
R1649 VSS.n171 VSS.n170 0.121553
R1650 VSS.n168 VSS.n167 0.121553
R1651 VSS.n167 VSS.n166 0.121553
R1652 VSS.n164 VSS.n163 0.121553
R1653 VSS.n163 VSS.n162 0.121553
R1654 VSS.n162 VSS.n161 0.121553
R1655 VSS.n159 VSS.n158 0.121553
R1656 VSS.n158 VSS.n157 0.121553
R1657 VSS.n155 VSS.n154 0.121553
R1658 VSS.n154 VSS.n153 0.121553
R1659 VSS.n153 VSS.n152 0.121553
R1660 VSS.n150 VSS.n149 0.121553
R1661 VSS.n983 VSS.n981 0.121553
R1662 VSS.n1284 VSS.n1283 0.121553
R1663 VSS.n1283 VSS.n1282 0.121553
R1664 VSS.n1282 VSS.n1281 0.121553
R1665 VSS.n1281 VSS.n1280 0.121553
R1666 VSS.n1280 VSS.n1279 0.121553
R1667 VSS.n1279 VSS.n1278 0.121553
R1668 VSS.n1278 VSS.n1277 0.121553
R1669 VSS.n1277 VSS.n1276 0.121553
R1670 VSS.n935 VSS.n231 0.121553
R1671 VSS.n937 VSS.n935 0.121553
R1672 VSS.n951 VSS.n937 0.121553
R1673 VSS.n953 VSS.n951 0.121553
R1674 VSS.n955 VSS.n953 0.121553
R1675 VSS.n957 VSS.n955 0.121553
R1676 VSS.n960 VSS.n957 0.121553
R1677 VSS.n962 VSS.n960 0.121553
R1678 VSS.n964 VSS.n962 0.121553
R1679 VSS.n998 VSS.n997 0.121553
R1680 VSS.n997 VSS.n996 0.121553
R1681 VSS.n996 VSS.n995 0.121553
R1682 VSS.n995 VSS.n994 0.121553
R1683 VSS.n994 VSS.n993 0.121553
R1684 VSS.n993 VSS.n992 0.121553
R1685 VSS.n992 VSS.n991 0.121553
R1686 VSS.n991 VSS.n990 0.121553
R1687 VSS.n990 VSS.n989 0.121553
R1688 VSS.n989 VSS.n988 0.121553
R1689 VSS.n988 VSS.n987 0.121553
R1690 VSS.n987 VSS.n986 0.121553
R1691 VSS.n986 VSS.n985 0.121553
R1692 VSS.n178 VSS.n177 0.118395
R1693 VSS.n455 VSS.n452 0.117688
R1694 VSS.n452 VSS.n449 0.117688
R1695 VSS.n449 VSS.n445 0.117688
R1696 VSS.n37 VSS.n35 0.116289
R1697 VSS.n39 VSS.n37 0.116289
R1698 VSS.n47 VSS.n45 0.116289
R1699 VSS.n52 VSS.n50 0.116289
R1700 VSS.n57 VSS.n55 0.116289
R1701 VSS.n62 VSS.n60 0.116289
R1702 VSS.n67 VSS.n65 0.116289
R1703 VSS.n73 VSS.n70 0.116289
R1704 VSS.n78 VSS.n76 0.116289
R1705 VSS.n83 VSS.n81 0.116289
R1706 VSS.n1295 VSS.n1293 0.116289
R1707 VSS.n1297 VSS.n1295 0.116289
R1708 VSS.n1299 VSS.n1297 0.116289
R1709 VSS.n1304 VSS.n1302 0.116289
R1710 VSS.n1306 VSS.n1304 0.116289
R1711 VSS.n1314 VSS.n1312 0.116289
R1712 VSS.n1316 VSS.n1314 0.116289
R1713 VSS.n1318 VSS.n1316 0.116289
R1714 VSS.n1323 VSS.n1321 0.116289
R1715 VSS.n1325 VSS.n1323 0.116289
R1716 VSS.n1327 VSS.n1325 0.116289
R1717 VSS.n1332 VSS.n1330 0.116289
R1718 VSS.n1334 VSS.n1332 0.116289
R1719 VSS.n1337 VSS.n1334 0.116289
R1720 VSS.n1342 VSS.n1340 0.116289
R1721 VSS.n1344 VSS.n1342 0.116289
R1722 VSS.n1346 VSS.n1344 0.116289
R1723 VSS.n1307 VSS.n1306 0.115763
R1724 VSS.n185 VSS.n184 0.115237
R1725 VSS.n442 VSS.n439 0.11207
R1726 VSS.n48 VSS.n47 0.109974
R1727 VSS.n81 VSS.n79 0.107868
R1728 VSS.n536 VSS.n533 0.107607
R1729 VSS.n300 VSS.n297 0.107607
R1730 VSS.n303 VSS.n300 0.107607
R1731 VSS.n306 VSS.n303 0.107607
R1732 VSS.n309 VSS.n306 0.107607
R1733 VSS.n312 VSS.n309 0.107607
R1734 VSS.n315 VSS.n312 0.107607
R1735 VSS.n318 VSS.n315 0.107607
R1736 VSS.n321 VSS.n318 0.107607
R1737 VSS.n324 VSS.n321 0.107607
R1738 VSS.n327 VSS.n324 0.107607
R1739 VSS.n330 VSS.n327 0.107607
R1740 VSS.n333 VSS.n330 0.107607
R1741 VSS.n336 VSS.n333 0.107607
R1742 VSS.n339 VSS.n336 0.107607
R1743 VSS.n342 VSS.n339 0.107607
R1744 VSS.n345 VSS.n342 0.107607
R1745 VSS.n348 VSS.n345 0.107607
R1746 VSS.n351 VSS.n348 0.107607
R1747 VSS.n354 VSS.n351 0.107607
R1748 VSS.n357 VSS.n354 0.107607
R1749 VSS.n360 VSS.n357 0.107607
R1750 VSS.n364 VSS.n360 0.107607
R1751 VSS.n169 VSS.n168 0.106816
R1752 VSS.n1118 VSS.n1115 0.10537
R1753 VSS.n246 VSS.n243 0.104161
R1754 VSS.n1227 VSS.n1226 0.104161
R1755 VSS.n1214 VSS.n1211 0.104161
R1756 VSS.n1202 VSS.n1199 0.104161
R1757 VSS.n1252 VSS.n1249 0.104161
R1758 VSS.n1267 VSS.n1264 0.104161
R1759 VSS.n243 VSS.n239 0.103357
R1760 VSS.n1199 VSS.n1196 0.103357
R1761 VSS.n1150 VSS.n1148 0.102773
R1762 VSS.n1226 VSS.n1223 0.10175
R1763 VSS.n1255 VSS.n1252 0.10175
R1764 VSS.n1237 VSS.n1236 0.0993393
R1765 VSS.n1211 VSS.n1208 0.0993393
R1766 VSS.n1245 VSS.n1242 0.0993393
R1767 VSS.n1270 VSS.n1267 0.0993393
R1768 VSS.n1140 VSS.n1139 0.0985357
R1769 VSS.n271 VSS.n270 0.0985357
R1770 VSS.n281 VSS.n279 0.0983261
R1771 VSS.n1130 VSS.n1127 0.0977321
R1772 VSS.n1144 VSS.n1140 0.0977321
R1773 VSS.n263 VSS.n260 0.0977321
R1774 VSS.n273 VSS.n271 0.0977321
R1775 VSS.n538 VSS.n536 0.0963383
R1776 VSS.n1127 VSS.n1124 0.096125
R1777 VSS.n1136 VSS.n1134 0.096125
R1778 VSS.n260 VSS.n257 0.096125
R1779 VSS.n267 VSS.n265 0.096125
R1780 VSS.n965 VSS.n964 0.0957632
R1781 VSS.n613 VSS.n610 0.0957326
R1782 VSS.n1236 VSS.n1233 0.0953214
R1783 VSS.n1223 VSS.n1220 0.0953214
R1784 VSS.n1246 VSS.n1245 0.0953214
R1785 VSS.n1258 VSS.n1255 0.0953214
R1786 VSS.n160 VSS.n159 0.0952368
R1787 VSS.n1237 VSS.n1144 0.0945179
R1788 VSS.n1231 VSS.n1227 0.0945179
R1789 VSS.n1217 VSS.n1214 0.0945179
R1790 VSS.n1205 VSS.n1202 0.0945179
R1791 VSS.n1242 VSS.n273 0.0945179
R1792 VSS.n1249 VSS.n1248 0.0945179
R1793 VSS.n1264 VSS.n1261 0.0945179
R1794 VSS.n1152 VSS.n1150 0.0937727
R1795 VSS.n157 VSS.n156 0.0931316
R1796 VSS.n526 VSS.n512 0.093
R1797 VSS.n512 VSS.n510 0.093
R1798 VSS.n510 VSS.n507 0.093
R1799 VSS.n507 VSS.n504 0.093
R1800 VSS.n504 VSS.n502 0.093
R1801 VSS.n502 VSS.n499 0.093
R1802 VSS.n499 VSS.n497 0.093
R1803 VSS.n497 VSS.n494 0.093
R1804 VSS.n494 VSS.n492 0.093
R1805 VSS.n492 VSS.n489 0.093
R1806 VSS.n489 VSS.n487 0.093
R1807 VSS.n487 VSS.n484 0.093
R1808 VSS.n484 VSS.n482 0.093
R1809 VSS.n482 VSS.n480 0.093
R1810 VSS.n480 VSS.n478 0.093
R1811 VSS.n478 VSS.n476 0.093
R1812 VSS.n476 VSS.n474 0.093
R1813 VSS.n474 VSS.n472 0.093
R1814 VSS.n472 VSS.n470 0.093
R1815 VSS.n470 VSS.n468 0.093
R1816 VSS.n468 VSS.n466 0.093
R1817 VSS.n466 VSS.n464 0.093
R1818 VSS.n464 VSS.n462 0.093
R1819 VSS.n748 VSS.n746 0.093
R1820 VSS.n750 VSS.n748 0.093
R1821 VSS.n752 VSS.n750 0.093
R1822 VSS.n754 VSS.n752 0.093
R1823 VSS.n756 VSS.n754 0.093
R1824 VSS.n758 VSS.n756 0.093
R1825 VSS.n760 VSS.n758 0.093
R1826 VSS.n762 VSS.n760 0.093
R1827 VSS.n764 VSS.n762 0.093
R1828 VSS.n767 VSS.n764 0.093
R1829 VSS.n769 VSS.n767 0.093
R1830 VSS.n772 VSS.n769 0.093
R1831 VSS.n774 VSS.n772 0.093
R1832 VSS.n777 VSS.n774 0.093
R1833 VSS.n779 VSS.n777 0.093
R1834 VSS.n782 VSS.n779 0.093
R1835 VSS.n784 VSS.n782 0.093
R1836 VSS.n788 VSS.n784 0.093
R1837 VSS.n690 VSS.n688 0.093
R1838 VSS.n692 VSS.n690 0.093
R1839 VSS.n694 VSS.n692 0.093
R1840 VSS.n696 VSS.n694 0.093
R1841 VSS.n699 VSS.n696 0.093
R1842 VSS.n702 VSS.n699 0.093
R1843 VSS.n705 VSS.n702 0.093
R1844 VSS.n708 VSS.n705 0.093
R1845 VSS.n711 VSS.n708 0.093
R1846 VSS.n714 VSS.n711 0.093
R1847 VSS.n717 VSS.n714 0.093
R1848 VSS.n720 VSS.n717 0.093
R1849 VSS.n723 VSS.n720 0.093
R1850 VSS.n726 VSS.n723 0.093
R1851 VSS.n729 VSS.n726 0.093
R1852 VSS.n732 VSS.n729 0.093
R1853 VSS.n734 VSS.n732 0.093
R1854 VSS.n744 VSS.n734 0.093
R1855 VSS.n1072 VSS.n1070 0.093
R1856 VSS.n1070 VSS.n1067 0.093
R1857 VSS.n1067 VSS.n1065 0.093
R1858 VSS.n1065 VSS.n1062 0.093
R1859 VSS.n1062 VSS.n1060 0.093
R1860 VSS.n1060 VSS.n1057 0.093
R1861 VSS.n1057 VSS.n1055 0.093
R1862 VSS.n1055 VSS.n1052 0.093
R1863 VSS.n1052 VSS.n1050 0.093
R1864 VSS.n1050 VSS.n1047 0.093
R1865 VSS.n1047 VSS.n1045 0.093
R1866 VSS.n1045 VSS.n1043 0.093
R1867 VSS.n1043 VSS.n1041 0.093
R1868 VSS.n1041 VSS.n1039 0.093
R1869 VSS.n1039 VSS.n1037 0.093
R1870 VSS.n1037 VSS.n1033 0.093
R1871 VSS.n1033 VSS.n1030 0.093
R1872 VSS.n1030 VSS.n1027 0.093
R1873 VSS.n1027 VSS.n1024 0.093
R1874 VSS.n1024 VSS.n1021 0.093
R1875 VSS.n867 VSS.n864 0.093
R1876 VSS.n864 VSS.n862 0.093
R1877 VSS.n1124 VSS.n1121 0.0929107
R1878 VSS.n257 VSS.n254 0.0929107
R1879 VSS.n195 VSS.n194 0.0923636
R1880 VSS.n1154 VSS.n1152 0.0921364
R1881 VSS.n45 VSS.n43 0.0915526
R1882 VSS.n65 VSS.n63 0.0910263
R1883 VSS.n87 VSS.n86 0.0910263
R1884 VSS.n1168 VSS.n1166 0.0905
R1885 VSS.n1180 VSS.n1178 0.0905
R1886 VSS.n1188 VSS.n1186 0.0905
R1887 VSS.n1134 VSS.n1130 0.0905
R1888 VSS.n1233 VSS.n1231 0.0905
R1889 VSS.n1220 VSS.n1217 0.0905
R1890 VSS.n1208 VSS.n1205 0.0905
R1891 VSS.n265 VSS.n263 0.0905
R1892 VSS.n1248 VSS.n1246 0.0905
R1893 VSS.n1261 VSS.n1258 0.0905
R1894 VSS.n368 VSS.n366 0.0897562
R1895 VSS.n370 VSS.n368 0.0897562
R1896 VSS.n372 VSS.n370 0.0897562
R1897 VSS.n374 VSS.n372 0.0897562
R1898 VSS.n376 VSS.n374 0.0897562
R1899 VSS.n378 VSS.n376 0.0897562
R1900 VSS.n381 VSS.n378 0.0897562
R1901 VSS.n383 VSS.n381 0.0897562
R1902 VSS.n386 VSS.n383 0.0897562
R1903 VSS.n388 VSS.n386 0.0897562
R1904 VSS.n391 VSS.n388 0.0897562
R1905 VSS.n393 VSS.n391 0.0897562
R1906 VSS.n396 VSS.n393 0.0897562
R1907 VSS.n398 VSS.n396 0.0897562
R1908 VSS.n401 VSS.n398 0.0897562
R1909 VSS.n403 VSS.n401 0.0897562
R1910 VSS.n410 VSS.n403 0.0897562
R1911 VSS.n412 VSS.n410 0.0897562
R1912 VSS.n415 VSS.n412 0.0897562
R1913 VSS.n417 VSS.n415 0.0897562
R1914 VSS.n420 VSS.n417 0.0897562
R1915 VSS.n423 VSS.n420 0.0897562
R1916 VSS.n426 VSS.n423 0.0897562
R1917 VSS.n429 VSS.n426 0.0897562
R1918 VSS.n432 VSS.n429 0.0897562
R1919 VSS.n435 VSS.n432 0.0897562
R1920 VSS.n439 VSS.n435 0.0897562
R1921 VSS.n283 VSS.n281 0.0897174
R1922 VSS.n1139 VSS.n1136 0.0896964
R1923 VSS.n270 VSS.n267 0.0896964
R1924 VSS.n1162 VSS.n1160 0.0896818
R1925 VSS.n42 VSS.n40 0.0889211
R1926 VSS.n1148 VSS.n1146 0.0888636
R1927 VSS.n1021 VSS.n1018 0.0888333
R1928 VSS.n285 VSS.n283 0.0881522
R1929 VSS.n1275 VSS.n231 0.0873421
R1930 VSS.n86 VSS.n84 0.0868158
R1931 VSS.n1081 VSS.n1079 0.086587
R1932 VSS.n1096 VSS.n1094 0.086587
R1933 VSS.n1108 VSS.n1106 0.086587
R1934 VSS.n294 VSS.n292 0.0858043
R1935 VSS.n1156 VSS.n1154 0.0855909
R1936 VSS.n1158 VSS.n1156 0.0855909
R1937 VSS.n1164 VSS.n1162 0.0855909
R1938 VSS.n1170 VSS.n1168 0.0855909
R1939 VSS.n1176 VSS.n1174 0.0855909
R1940 VSS.n1182 VSS.n1180 0.0855909
R1941 VSS.n1186 VSS.n1184 0.0855909
R1942 VSS.n1193 VSS.n1188 0.0855909
R1943 VSS.n279 VSS.n277 0.0850217
R1944 VSS.n528 VSS.n526 0.0838333
R1945 VSS.n151 VSS.n150 0.0836579
R1946 VSS.n235 VSS.n233 0.0831364
R1947 VSS.n1174 VSS.n1172 0.0831364
R1948 VSS.n1302 VSS.n1300 0.0831316
R1949 VSS.n1073 VSS.n1072 0.083
R1950 VSS.n458 VSS.n456 0.0828529
R1951 VSS.n1321 VSS.n1319 0.0826053
R1952 VSS.n610 VSS.n609 0.0824863
R1953 VSS.n287 VSS.n285 0.0818913
R1954 VSS.n290 VSS.n287 0.0818913
R1955 VSS.n1084 VSS.n1081 0.0818913
R1956 VSS.n1092 VSS.n1088 0.0818913
R1957 VSS.n1101 VSS.n1096 0.0818913
R1958 VSS.n1106 VSS.n1104 0.0818913
R1959 VSS.n1115 VSS.n1108 0.0818913
R1960 VSS.n166 VSS.n165 0.0815526
R1961 VSS.n1088 VSS.n1086 0.0795435
R1962 VSS.n1340 VSS.n1338 0.0783947
R1963 VSS.n1160 VSS.n1158 0.0782273
R1964 VSS.n1166 VSS.n1164 0.0782273
R1965 VSS.n1172 VSS.n1170 0.0782273
R1966 VSS.n1178 VSS.n1176 0.0782273
R1967 VSS.n1184 VSS.n1182 0.0782273
R1968 VSS.n277 VSS.n275 0.076413
R1969 VSS.n58 VSS.n57 0.0762895
R1970 VSS.n251 VSS.n250 0.0756304
R1971 VSS.n238 VSS.n236 0.0749681
R1972 VSS.n292 VSS.n290 0.0748478
R1973 VSS.n1079 VSS.n1077 0.0748478
R1974 VSS.n1086 VSS.n1084 0.0748478
R1975 VSS.n1094 VSS.n1092 0.0748478
R1976 VSS.n1104 VSS.n1101 0.0748478
R1977 VSS.n540 VSS.n538 0.0744726
R1978 VSS.n542 VSS.n540 0.0744726
R1979 VSS.n544 VSS.n542 0.0744726
R1980 VSS.n546 VSS.n544 0.0744726
R1981 VSS.n548 VSS.n546 0.0744726
R1982 VSS.n550 VSS.n548 0.0744726
R1983 VSS.n553 VSS.n550 0.0744726
R1984 VSS.n555 VSS.n553 0.0744726
R1985 VSS.n558 VSS.n555 0.0744726
R1986 VSS.n560 VSS.n558 0.0744726
R1987 VSS.n563 VSS.n560 0.0744726
R1988 VSS.n565 VSS.n563 0.0744726
R1989 VSS.n568 VSS.n565 0.0744726
R1990 VSS.n571 VSS.n568 0.0744726
R1991 VSS.n573 VSS.n571 0.0744726
R1992 VSS.n576 VSS.n573 0.0744726
R1993 VSS.n578 VSS.n576 0.0744726
R1994 VSS.n585 VSS.n578 0.0744726
R1995 VSS.n588 VSS.n585 0.0744726
R1996 VSS.n590 VSS.n588 0.0744726
R1997 VSS.n593 VSS.n590 0.0744726
R1998 VSS.n595 VSS.n593 0.0744726
R1999 VSS.n598 VSS.n595 0.0744726
R2000 VSS.n600 VSS.n598 0.0744726
R2001 VSS.n603 VSS.n600 0.0744726
R2002 VSS.n605 VSS.n603 0.0744726
R2003 VSS.n609 VSS.n605 0.0744726
R2004 VSS.n70 VSS.n68 0.0741842
R2005 VSS.n1328 VSS.n1327 0.0720789
R2006 VSS.n529 VSS.n528 0.0713333
R2007 VSS.n175 VSS.n174 0.0699737
R2008 VSS.n1001 VSS 0.0689956
R2009 VSS VSS.n888 0.0689956
R2010 VSS VSS.n889 0.0689956
R2011 VSS VSS.n1003 0.0689956
R2012 VSS VSS.n1007 0.0689956
R2013 VSS VSS.n870 0.0689956
R2014 VSS.n1196 VSS.n1193 0.0689789
R2015 VSS.n366 VSS.n364 0.068186
R2016 VSS.n1310 VSS.n1309 0.0678684
R2017 VSS.n445 VSS.n442 0.0648001
R2018 VSS.n74 VSS.n73 0.0636579
R2019 VSS.n183 VSS.n182 0.0636579
R2020 VSS.n906 VSS.n904 0.062959
R2021 VSS.n1288 VSS.n1287 0.0624089
R2022 VSS.n30 VSS.n29 0.0615526
R2023 VSS.n239 VSS.n235 0.0607533
R2024 VSS.n53 VSS.n52 0.0594474
R2025 VSS.n33 VSS.n32 0.058921
R2026 VSS.n184 VSS.n183 0.0583947
R2027 VSS.n35 VSS.n33 0.0578684
R2028 VSS.n55 VSS.n53 0.0573421
R2029 VSS.n32 VSS.n30 0.0552368
R2030 VSS.n1121 VSS.n1118 0.05508
R2031 VSS.n76 VSS.n74 0.0531316
R2032 VSS.n1271 VSS.n1270 0.0527321
R2033 VSS.n174 VSS.n173 0.052079
R2034 VSS.n254 VSS.n251 0.0503214
R2035 VSS.n1293 VSS.n1291 0.0494474
R2036 VSS.n1312 VSS.n1310 0.0489211
R2037 VSS.n1330 VSS.n1328 0.0447105
R2038 VSS.n68 VSS.n67 0.0426053
R2039 VSS.n1074 VSS.n294 0.0411957
R2040 VSS.n1077 VSS.n1074 0.0411957
R2041 VSS.n60 VSS.n58 0.0405
R2042 VSS.n165 VSS.n164 0.0405
R2043 VSS.n1338 VSS.n1337 0.0383947
R2044 VSS.n152 VSS.n151 0.0383947
R2045 VSS.n1271 VSS.n246 0.0366607
R2046 VSS.n1276 VSS.n1275 0.0347105
R2047 VSS.n1319 VSS.n1318 0.0341842
R2048 VSS.n1300 VSS.n1299 0.0336579
R2049 VSS.n84 VSS.n83 0.0299737
R2050 VSS.n156 VSS.n155 0.0289211
R2051 VSS.n40 VSS.n39 0.0278684
R2052 VSS.n161 VSS.n160 0.0268158
R2053 VSS.n998 VSS.n965 0.0262895
R2054 VSS.n63 VSS.n62 0.0257632
R2055 VSS.n89 VSS.n87 0.0257632
R2056 VSS.n610 VSS.n530 0.0257083
R2057 VSS.n43 VSS.n42 0.0252368
R2058 VSS.n193 VSS.n192 0.0231316
R2059 VSS.n170 VSS.n169 0.0152368
R2060 VSS.n686 VSS.n685 0.0151318
R2061 VSS.n686 VSS.n455 0.013625
R2062 VSS.n194 VSS.n193 0.013217
R2063 VSS.n1073 VSS.n744 0.0105
R2064 VSS.n79 VSS.n78 0.00892105
R2065 VSS VSS.n89 0.00892105
R2066 VSS.n50 VSS.n48 0.00681579
R2067 VSS.n192 VSS.n185 0.00681579
R2068 VSS.n1347 VSS.n1346 0.00471053
R2069 VSS.n1018 VSS.n867 0.00466667
R2070 VSS.n179 VSS.n178 0.00365789
R2071 VSS.n1274 VSS.n1271 0.00276891
R2072 VSS.n939 VSS 0.00129646
R2073 VSS.n943 VSS 0.00129646
R2074 VSS.n947 VSS 0.00129646
R2075 VSS.n1005 VSS 0.00129646
R2076 VSS.n1009 VSS 0.00129646
R2077 VSS.n1016 VSS 0.00129646
R2078 VSS.n1309 VSS.n1307 0.00102632
R2079 B6 B6.t1 48.6474
R2080 B6.n0 B6.t2 19.0247
R2081 B6.n0 B6.t0 17.3935
R2082 B6.n1 B6.n0 4.12942
R2083 B6.n1 B6 2.25699
R2084 B6 B6.n1 0.0067069
R2085 VDD.n1 VDD.t54 490.522
R2086 VDD.n5 VDD.t0 490.522
R2087 VDD.n10 VDD.t69 490.522
R2088 VDD.n27 VDD.t83 490.522
R2089 VDD.n22 VDD.t49 490.522
R2090 VDD.n17 VDD.t95 490.522
R2091 VDD.n1 VDD.t77 485.783
R2092 VDD.n5 VDD.t59 485.783
R2093 VDD.n10 VDD.t13 485.783
R2094 VDD.n27 VDD.t63 485.783
R2095 VDD.n22 VDD.t52 485.783
R2096 VDD.n17 VDD.t15 485.783
R2097 VDD VDD.t67 432.043
R2098 VDD VDD.t40 432.043
R2099 VDD VDD.t3 432.043
R2100 VDD VDD.t65 432.043
R2101 VDD VDD.t73 432.043
R2102 VDD VDD.t61 432.043
R2103 VDD.n135 VDD.n134 345.764
R2104 VDD.n120 VDD.t47 166.102
R2105 VDD.n135 VDD.t21 161.018
R2106 VDD.n106 VDD.t34 159.322
R2107 VDD.n122 VDD.t35 155.933
R2108 VDD.n137 VDD.t36 150.847
R2109 VDD.n104 VDD.t18 149.154
R2110 VDD.n124 VDD.t75 145.763
R2111 VDD.n139 VDD.t19 140.679
R2112 VDD.n102 VDD.t10 138.983
R2113 VDD.n45 VDD.t26 135.114
R2114 VDD.n141 VDD.t24 130.508
R2115 VDD.n117 VDD.t42 118.865
R2116 VDD.n46 VDD.t37 118.644
R2117 VDD.n88 VDD.t17 118.644
R2118 VDD.n115 VDD.t5 111.865
R2119 VDD.n155 VDD.t20 110.169
R2120 VDD.n48 VDD.t79 108.475
R2121 VDD.n86 VDD.t9 108.475
R2122 VDD.n157 VDD.t58 100.001
R2123 VDD.n50 VDD.t38 98.3056
R2124 VDD.n84 VDD.t31 98.3056
R2125 VDD.n93 VDD.t45 98.3056
R2126 VDD.n158 VDD.t86 89.831
R2127 VDD.n53 VDD.t80 88.1361
R2128 VDD.n55 VDD.t57 77.9666
R2129 VDD.n70 VDD.t72 77.9666
R2130 VDD.n57 VDD.t91 67.7971
R2131 VDD.n68 VDD.t48 67.7971
R2132 VDD.n75 VDD.t7 67.7971
R2133 VDD.n59 VDD.t29 57.6276
R2134 VDD.n66 VDD.t92 57.6276
R2135 VDD.n149 VDD.t88 52.5429
R2136 VDD.n6 VDD.t60 9.56883
R2137 VDD.n11 VDD.t14 9.56883
R2138 VDD.n18 VDD.t16 9.56883
R2139 VDD.n2 VDD.t78 9.56883
R2140 VDD.n7 VDD.n4 9.47246
R2141 VDD.n12 VDD.n9 9.47246
R2142 VDD.n19 VDD.n16 9.47246
R2143 VDD.n24 VDD.n15 9.47246
R2144 VDD.n21 VDD.t53 9.47246
R2145 VDD.n29 VDD.n14 9.47246
R2146 VDD.n26 VDD.t64 9.47246
R2147 VDD.n3 VDD.n0 9.47246
R2148 VDD.n65 VDD.n64 8.30127
R2149 VDD.n126 VDD.t76 7.67003
R2150 VDD.n8 VDD.t68 6.40636
R2151 VDD.n13 VDD.t41 6.40636
R2152 VDD.n20 VDD.t4 6.40636
R2153 VDD.n25 VDD.t66 6.40636
R2154 VDD.n30 VDD.t74 6.40636
R2155 VDD.n165 VDD.t62 6.40636
R2156 VDD.n6 VDD.n5 6.3005
R2157 VDD.n11 VDD.n10 6.3005
R2158 VDD.n18 VDD.n17 6.3005
R2159 VDD.n23 VDD.n22 6.3005
R2160 VDD.n28 VDD.n27 6.3005
R2161 VDD.n150 VDD.n149 6.3005
R2162 VDD.n134 VDD.n133 6.3005
R2163 VDD.n118 VDD.n115 6.3005
R2164 VDD.n94 VDD.n93 6.3005
R2165 VDD.n76 VDD.n75 6.3005
R2166 VDD.n47 VDD.n46 6.3005
R2167 VDD.n49 VDD.n48 6.3005
R2168 VDD.n51 VDD.n50 6.3005
R2169 VDD.n54 VDD.n53 6.3005
R2170 VDD.n56 VDD.n55 6.3005
R2171 VDD.n58 VDD.n57 6.3005
R2172 VDD.n60 VDD.n59 6.3005
R2173 VDD.n63 VDD.n62 6.3005
R2174 VDD.n67 VDD.n66 6.3005
R2175 VDD.n69 VDD.n68 6.3005
R2176 VDD.n71 VDD.n70 6.3005
R2177 VDD.n85 VDD.n84 6.3005
R2178 VDD.n87 VDD.n86 6.3005
R2179 VDD.n89 VDD.n88 6.3005
R2180 VDD.n103 VDD.n102 6.3005
R2181 VDD.n105 VDD.n104 6.3005
R2182 VDD.n107 VDD.n106 6.3005
R2183 VDD.n121 VDD.n120 6.3005
R2184 VDD.n123 VDD.n122 6.3005
R2185 VDD.n125 VDD.n124 6.3005
R2186 VDD.n136 VDD.n135 6.3005
R2187 VDD.n138 VDD.n137 6.3005
R2188 VDD.n140 VDD.n139 6.3005
R2189 VDD.n142 VDD.n141 6.3005
R2190 VDD.n160 VDD.n157 6.3005
R2191 VDD.n159 VDD.n158 6.3005
R2192 VDD.n2 VDD.n1 6.3005
R2193 VDD.n159 VDD.t87 6.18063
R2194 VDD.n45 VDD.n44 6.10984
R2195 VDD.n40 VDD.n39 6.09557
R2196 VDD.n61 VDD.t30 6.09557
R2197 VDD.n114 VDD.n113 4.98502
R2198 VDD.n164 VDD.n163 4.7945
R2199 VDD.n133 VDD.n132 4.5005
R2200 VDD.n94 VDD.n92 4.5005
R2201 VDD.n76 VDD.n74 4.5005
R2202 VDD.n150 VDD.n148 4.5005
R2203 VDD.n101 VDD.n100 4.26092
R2204 VDD.n83 VDD.n82 4.24066
R2205 VDD.n156 VDD.n155 3.70778
R2206 VDD.n31 VDD.n30 3.57624
R2207 VDD.n100 VDD.n99 3.2271
R2208 VDD.n82 VDD.n81 3.20234
R2209 VDD.n113 VDD.n112 3.17695
R2210 VDD.n164 VDD.n32 3.16881
R2211 VDD.n96 VDD.n95 3.15175
R2212 VDD.n130 VDD.n129 3.15175
R2213 VDD.n78 VDD.n77 3.15175
R2214 VDD.n111 VDD.n110 3.15175
R2215 VDD.n152 VDD.n151 3.15175
R2216 VDD.n130 VDD.n41 3.151
R2217 VDD.n79 VDD.n78 3.151
R2218 VDD.n151 VDD.n147 3.151
R2219 VDD.n110 VDD.n109 3.151
R2220 VDD.n97 VDD.n96 3.151
R2221 VDD.n144 VDD.n38 3.06224
R2222 VDD.n52 VDD.n43 3.06224
R2223 VDD.n38 VDD.t25 3.03383
R2224 VDD.n38 VDD.n37 3.03383
R2225 VDD.n43 VDD.t39 3.03383
R2226 VDD.n43 VDD.n42 3.03383
R2227 VDD.n113 VDD.t6 2.69573
R2228 VDD.n82 VDD.t8 2.66058
R2229 VDD.n31 VDD.n13 2.63002
R2230 VDD.n32 VDD.n8 2.62915
R2231 VDD.n100 VDD.t46 2.62483
R2232 VDD.n119 VDD.n118 2.62147
R2233 VDD.n163 VDD.n34 2.3203
R2234 VDD.n163 VDD.n162 2.31907
R2235 VDD.n76 VDD.n73 1.88512
R2236 VDD.n118 VDD.n116 1.83127
R2237 VDD.n133 VDD.n131 1.77742
R2238 VDD.n94 VDD.n91 1.56204
R2239 VDD.n162 VDD.n161 1.49872
R2240 VDD.n96 VDD.n94 1.12174
R2241 VDD.n32 VDD.n31 0.911065
R2242 VDD.n26 VDD.n25 0.742062
R2243 VDD.n21 VDD.n20 0.727335
R2244 VDD.n133 VDD.n130 0.724621
R2245 VDD.n151 VDD.n150 0.59316
R2246 VDD.n78 VDD.n76 0.525399
R2247 VDD VDD.n7 0.510235
R2248 VDD VDD.n12 0.510235
R2249 VDD VDD.n19 0.510235
R2250 VDD VDD.n24 0.510235
R2251 VDD VDD.n29 0.510235
R2252 VDD VDD.n3 0.491916
R2253 VDD.n118 VDD.n117 0.415309
R2254 VDD.n165 VDD.n164 0.394447
R2255 VDD.n47 VDD.n45 0.115744
R2256 VDD.n49 VDD.n47 0.115744
R2257 VDD.n51 VDD.n49 0.115744
R2258 VDD.n56 VDD.n54 0.115744
R2259 VDD.n58 VDD.n56 0.115744
R2260 VDD.n60 VDD.n58 0.115744
R2261 VDD.n69 VDD.n67 0.115744
R2262 VDD.n71 VDD.n69 0.115744
R2263 VDD.n87 VDD.n85 0.115744
R2264 VDD.n89 VDD.n87 0.115744
R2265 VDD.n105 VDD.n103 0.115744
R2266 VDD.n107 VDD.n105 0.115744
R2267 VDD.n123 VDD.n121 0.115744
R2268 VDD.n125 VDD.n123 0.115744
R2269 VDD.n138 VDD.n136 0.115744
R2270 VDD.n140 VDD.n138 0.115744
R2271 VDD.n142 VDD.n140 0.115744
R2272 VDD.n160 VDD.n159 0.115744
R2273 VDD.n72 VDD.n71 0.109159
R2274 VDD.n161 VDD.n160 0.108104
R2275 VDD.n121 VDD.n119 0.106804
R2276 VDD.n90 VDD.n89 0.105866
R2277 VDD.n108 VDD.n107 0.0970854
R2278 VDD.n23 VDD.n21 0.0968717
R2279 VDD.n28 VDD.n26 0.0968717
R2280 VDD VDD.n40 0.0959878
R2281 VDD.n103 VDD.n101 0.0957073
R2282 VDD.n126 VDD.n125 0.0953491
R2283 VDD.n85 VDD.n83 0.0913202
R2284 VDD.n52 VDD.n51 0.0883049
R2285 VDD.n7 VDD 0.0857212
R2286 VDD.n12 VDD 0.0857212
R2287 VDD.n19 VDD 0.0857212
R2288 VDD.n24 VDD 0.0857212
R2289 VDD.n29 VDD 0.0857212
R2290 VDD.n3 VDD 0.0857212
R2291 VDD.n143 VDD.n142 0.085561
R2292 VDD.n67 VDD.n65 0.0789756
R2293 VDD.n61 VDD.n60 0.0751341
R2294 VDD.n65 VDD.n63 0.0723902
R2295 VDD.n154 VDD.n153 0.0690976
R2296 VDD.n8 VDD 0.0594381
R2297 VDD.n13 VDD 0.0594381
R2298 VDD.n20 VDD 0.0594381
R2299 VDD.n25 VDD 0.0594381
R2300 VDD.n30 VDD 0.0594381
R2301 VDD VDD.n165 0.0594381
R2302 VDD.n63 VDD.n61 0.0411098
R2303 VDD.n36 VDD.n35 0.0282397
R2304 VDD.n54 VDD.n52 0.027939
R2305 VDD.n156 VDD.n154 0.0251951
R2306 VDD.n153 VDD.n152 0.0224512
R2307 VDD.n111 VDD.n108 0.0191585
R2308 VDD.n80 VDD.n79 0.018061
R2309 VDD.n129 VDD.n127 0.0153171
R2310 VDD.n98 VDD.n97 0.0147683
R2311 VDD VDD.n6 0.0140398
R2312 VDD VDD.n11 0.0140398
R2313 VDD VDD.n18 0.0140398
R2314 VDD VDD.n23 0.0140398
R2315 VDD VDD.n28 0.0140398
R2316 VDD VDD.n2 0.0140398
R2317 VDD.n144 VDD.n143 0.0136707
R2318 VDD.n128 VDD 0.013122
R2319 VDD.n97 VDD.n90 0.010378
R2320 VDD.n161 VDD.n156 0.0100485
R2321 VDD.n129 VDD.n128 0.00982927
R2322 VDD.n83 VDD.n80 0.00933668
R2323 VDD.n145 VDD.n144 0.00928049
R2324 VDD.n119 VDD.n114 0.00876098
R2325 VDD.n101 VDD.n98 0.00824116
R2326 VDD.n127 VDD.n126 0.00805275
R2327 VDD.n34 VDD.n33 0.00728082
R2328 VDD.n79 VDD.n72 0.00708537
R2329 VDD.n146 VDD.n145 0.00653659
R2330 VDD.n136 VDD.n40 0.00434146
R2331 VDD.n152 VDD.n146 0.00269512
R2332 VDD.n114 VDD.n111 0.00214634
R2333 VDD.n162 VDD.n36 0.00111644
R2334 SDn_2.n34 SDn_2.n33 133.643
R2335 SDn_2.n42 SDn_2.n41 48.6672
R2336 SDn_2.n69 SDn_2.n68 47.4505
R2337 SDn_2.n3 SDn_2.t52 35.1054
R2338 SDn_2.n62 SDn_2.t63 34.0104
R2339 SDn_2.n72 SDn_2.n71 21.2922
R2340 SDn_2.n63 SDn_2.n62 21.0894
R2341 SDn_2.n64 SDn_2.n63 21.0894
R2342 SDn_2.n65 SDn_2.n64 21.0894
R2343 SDn_2.n66 SDn_2.n65 21.0894
R2344 SDn_2.n67 SDn_2.n66 21.0894
R2345 SDn_2.n68 SDn_2.n67 21.0894
R2346 SDn_2.n70 SDn_2.n69 21.0894
R2347 SDn_2.n72 SDn_2.n70 21.0894
R2348 SDn_2.n44 SDn_2.n43 21.0894
R2349 SDn_2.n4 SDn_2.n3 21.0894
R2350 SDn_2.n5 SDn_2.n4 21.0894
R2351 SDn_2.n6 SDn_2.n5 21.0894
R2352 SDn_2.n7 SDn_2.n6 21.0894
R2353 SDn_2.n8 SDn_2.n7 21.0894
R2354 SDn_2.n9 SDn_2.n8 21.0894
R2355 SDn_2.n10 SDn_2.n9 21.0894
R2356 SDn_2.n11 SDn_2.n10 21.0894
R2357 SDn_2.n12 SDn_2.n11 21.0894
R2358 SDn_2.n13 SDn_2.n12 21.0894
R2359 SDn_2.n14 SDn_2.n13 21.0894
R2360 SDn_2.n15 SDn_2.n14 21.0894
R2361 SDn_2.n16 SDn_2.n15 21.0894
R2362 SDn_2.n17 SDn_2.n16 21.0894
R2363 SDn_2.n18 SDn_2.n17 21.0894
R2364 SDn_2.n19 SDn_2.n18 21.0894
R2365 SDn_2.n20 SDn_2.n19 21.0894
R2366 SDn_2.n21 SDn_2.n20 21.0894
R2367 SDn_2.n22 SDn_2.n21 21.0894
R2368 SDn_2.n23 SDn_2.n22 21.0894
R2369 SDn_2.n24 SDn_2.n23 21.0894
R2370 SDn_2.n25 SDn_2.n24 21.0894
R2371 SDn_2.n26 SDn_2.n25 21.0894
R2372 SDn_2.n27 SDn_2.n26 21.0894
R2373 SDn_2.n28 SDn_2.n27 21.0894
R2374 SDn_2.n29 SDn_2.n28 21.0894
R2375 SDn_2.n30 SDn_2.n29 21.0894
R2376 SDn_2.n31 SDn_2.n30 21.0894
R2377 SDn_2.n32 SDn_2.n31 21.0894
R2378 SDn_2.n33 SDn_2.n32 21.0894
R2379 SDn_2.n35 SDn_2.n34 21.0894
R2380 SDn_2.n36 SDn_2.n35 21.0894
R2381 SDn_2.n37 SDn_2.n36 21.0894
R2382 SDn_2.n38 SDn_2.n37 21.0894
R2383 SDn_2.n39 SDn_2.n38 21.0894
R2384 SDn_2.n40 SDn_2.n39 21.0894
R2385 SDn_2.n41 SDn_2.n40 21.0894
R2386 SDn_2.n45 SDn_2.n42 21.0894
R2387 SDn_2.n45 SDn_2.n44 21.0894
R2388 SDn_2.n3 SDn_2.t67 14.7465
R2389 SDn_2.n4 SDn_2.t75 14.7465
R2390 SDn_2.n7 SDn_2.t38 14.7465
R2391 SDn_2.n8 SDn_2.t70 14.7465
R2392 SDn_2.n11 SDn_2.t71 14.7465
R2393 SDn_2.n12 SDn_2.t61 14.7465
R2394 SDn_2.n15 SDn_2.t48 14.7465
R2395 SDn_2.n16 SDn_2.t74 14.7465
R2396 SDn_2.n19 SDn_2.t73 14.7465
R2397 SDn_2.n20 SDn_2.t64 14.7465
R2398 SDn_2.n23 SDn_2.t51 14.7465
R2399 SDn_2.n24 SDn_2.t30 14.7465
R2400 SDn_2.n27 SDn_2.t24 14.7465
R2401 SDn_2.n28 SDn_2.t56 14.7465
R2402 SDn_2.n31 SDn_2.t59 14.7465
R2403 SDn_2.n32 SDn_2.t43 14.7465
R2404 SDn_2.n62 SDn_2.t55 14.3815
R2405 SDn_2.n63 SDn_2.t66 14.3815
R2406 SDn_2.n66 SDn_2.t57 14.3815
R2407 SDn_2.n67 SDn_2.t32 14.3815
R2408 SDn_2.n70 SDn_2.t12 14.3815
R2409 SDn_2.n44 SDn_2.t10 14.3815
R2410 SDn_2.n35 SDn_2.t69 14.3815
R2411 SDn_2.n36 SDn_2.t40 14.3815
R2412 SDn_2.n39 SDn_2.t33 14.3815
R2413 SDn_2.n40 SDn_2.t54 14.3815
R2414 SDn_2.n5 SDn_2.t68 14.0165
R2415 SDn_2.n6 SDn_2.t35 14.0165
R2416 SDn_2.n9 SDn_2.t36 14.0165
R2417 SDn_2.n10 SDn_2.t49 14.0165
R2418 SDn_2.n13 SDn_2.t44 14.0165
R2419 SDn_2.n14 SDn_2.t27 14.0165
R2420 SDn_2.n17 SDn_2.t72 14.0165
R2421 SDn_2.n18 SDn_2.t46 14.0165
R2422 SDn_2.n21 SDn_2.t50 14.0165
R2423 SDn_2.n22 SDn_2.t29 14.0165
R2424 SDn_2.n25 SDn_2.t34 14.0165
R2425 SDn_2.n26 SDn_2.t65 14.0165
R2426 SDn_2.n29 SDn_2.t53 14.0165
R2427 SDn_2.n30 SDn_2.t41 14.0165
R2428 SDn_2.n33 SDn_2.t25 14.0165
R2429 SDn_2.n69 SDn_2.t6 12.9916
R2430 SDn_2.n71 SDn_2.t4 12.9916
R2431 SDn_2.n43 SDn_2.t0 12.9916
R2432 SDn_2.n64 SDn_2.t47 12.9215
R2433 SDn_2.n65 SDn_2.t39 12.9215
R2434 SDn_2.n68 SDn_2.t58 12.9215
R2435 SDn_2.n34 SDn_2.t60 12.9215
R2436 SDn_2.n37 SDn_2.t37 12.9215
R2437 SDn_2.n38 SDn_2.t31 12.9215
R2438 SDn_2.n41 SDn_2.t28 12.9215
R2439 SDn_2.n42 SDn_2.t14 12.9215
R2440 SDn_2.n74 SDn_2.t2 10.7743
R2441 SDn_2.n47 SDn_2.t8 10.7743
R2442 SDn_2.n75 SDn_2.n73 3.54502
R2443 SDn_2.n48 SDn_2.n46 3.54477
R2444 SDn_2.n75 SDn_2.n74 3.50535
R2445 SDn_2.n48 SDn_2.n47 3.50535
R2446 SDn_2.n59 SDn_2.n56 3.07598
R2447 SDn_2.n85 SDn_2.n52 3.01065
R2448 SDn_2.n54 SDn_2.n53 2.90221
R2449 SDn_2.n82 SDn_2.n81 2.90214
R2450 SDn_2.n77 SDn_2.n76 2.88451
R2451 SDn_2.n49 SDn_2.n2 2.88438
R2452 SDn_2.n61 SDn_2.n60 2.87834
R2453 SDn_2.n56 SDn_2.n55 2.87828
R2454 SDn_2.n58 SDn_2.n57 2.87828
R2455 SDn_2.n52 SDn_2.n51 2.82902
R2456 SDn_2.n50 SDn_2.n1 2.76772
R2457 SDn_2.n78 SDn_2.n61 2.75462
R2458 SDn_2.n1 SDn_2.t20 2.7305
R2459 SDn_2.n1 SDn_2.n0 2.7305
R2460 SDn_2.n90 SDn_2.t9 2.7305
R2461 SDn_2.n90 SDn_2.n89 2.7305
R2462 SDn_2.n59 SDn_2.n58 2.50797
R2463 SDn_2.n80 SDn_2.n54 2.50522
R2464 SDn_2.n52 SDn_2.t1 2.49942
R2465 SDn_2.n58 SDn_2.t17 2.43824
R2466 SDn_2.n56 SDn_2.t7 2.43824
R2467 SDn_2.n61 SDn_2.t18 2.4382
R2468 SDn_2.n82 SDn_2.t16 2.40701
R2469 SDn_2.n54 SDn_2.t3 2.40696
R2470 SDn_2.n78 SDn_2.n77 2.35277
R2471 SDn_2.n50 SDn_2.n49 2.3515
R2472 SDn_2.n84 SDn_2.n83 2.24989
R2473 SDn_2.n93 SDn_2.n92 1.50283
R2474 SDn_2.n91 SDn_2.n90 1.42666
R2475 SDn_2.n83 SDn_2.n82 1.0106
R2476 SDn_2.n46 SDn_2.n45 0.967483
R2477 SDn_2.n73 SDn_2.n72 0.96743
R2478 SDn_2.n84 SDn_2.n80 0.610728
R2479 SDn_2.n79 SDn_2.n59 0.564953
R2480 SDn_2.n87 SDn_2.n86 0.560976
R2481 SDn_2.n79 SDn_2.n78 0.141929
R2482 SDn_2.n91 SDn_2 0.140162
R2483 SDn_2.n88 SDn_2.n50 0.119429
R2484 SDn_2.n88 SDn_2.n87 0.0205
R2485 SDn_2.n86 SDn_2.n85 0.0171667
R2486 SDn_2.n92 SDn_2.n91 0.0135282
R2487 SDn_2.n80 SDn_2.n79 0.013514
R2488 SDn_2.n85 SDn_2.n84 0.0109989
R2489 SDn_2.n93 SDn_2.n88 0.00943873
R2490 SDn_2.n49 SDn_2.n48 0.0045
R2491 SDn_2 SDn_2.n93 0.00355856
R2492 SDn_2.n77 SDn_2.n75 0.0025
R2493 SD3_1.n97 SD3_1.n7 3.48971
R2494 SD3_1.n109 SD3_1.n3 3.48281
R2495 SD3_1.n56 SD3_1.n55 3.07792
R2496 SD3_1.n85 SD3_1.n27 3.07726
R2497 SD3_1.n88 SD3_1.n22 3.07632
R2498 SD3_1.n120 SD3_1.n117 3.07564
R2499 SD3_1.n76 SD3_1.n42 3.0732
R2500 SD3_1.n82 SD3_1.n32 3.07118
R2501 SD3_1.n79 SD3_1.n37 3.06982
R2502 SD3_1.n70 SD3_1.n44 3.06866
R2503 SD3_1.n91 SD3_1.n17 3.06533
R2504 SD3_1.n64 SD3_1.n49 3.06484
R2505 SD3_1 SD3_1.n1 3.06384
R2506 SD3_1.n58 SD3_1.n51 3.05987
R2507 SD3_1.n100 SD3_1.n5 3.05915
R2508 SD3_1.n94 SD3_1.n12 3.05307
R2509 SD3_1.n12 SD3_1.n11 2.90211
R2510 SD3_1.n102 SD3_1.n101 2.90208
R2511 SD3_1.n119 SD3_1.t51 2.7305
R2512 SD3_1.n119 SD3_1.n118 2.7305
R2513 SD3_1.n117 SD3_1.t3 2.7305
R2514 SD3_1.n117 SD3_1.n116 2.7305
R2515 SD3_1.n106 SD3_1.t42 2.7305
R2516 SD3_1.n106 SD3_1.n105 2.7305
R2517 SD3_1.n9 SD3_1.t57 2.7305
R2518 SD3_1.n9 SD3_1.n8 2.7305
R2519 SD3_1.n14 SD3_1.t24 2.7305
R2520 SD3_1.n14 SD3_1.n13 2.7305
R2521 SD3_1.n19 SD3_1.t39 2.7305
R2522 SD3_1.n19 SD3_1.n18 2.7305
R2523 SD3_1.n24 SD3_1.t16 2.7305
R2524 SD3_1.n24 SD3_1.n23 2.7305
R2525 SD3_1.n29 SD3_1.t31 2.7305
R2526 SD3_1.n29 SD3_1.n28 2.7305
R2527 SD3_1.n34 SD3_1.t22 2.7305
R2528 SD3_1.n34 SD3_1.n33 2.7305
R2529 SD3_1.n39 SD3_1.t40 2.7305
R2530 SD3_1.n39 SD3_1.n38 2.7305
R2531 SD3_1.n73 SD3_1.t11 2.7305
R2532 SD3_1.n73 SD3_1.n72 2.7305
R2533 SD3_1.n46 SD3_1.t35 2.7305
R2534 SD3_1.n46 SD3_1.n45 2.7305
R2535 SD3_1.n66 SD3_1.t0 2.7305
R2536 SD3_1.n66 SD3_1.n65 2.7305
R2537 SD3_1.n60 SD3_1.t30 2.7305
R2538 SD3_1.n60 SD3_1.n59 2.7305
R2539 SD3_1.n53 SD3_1.t17 2.7305
R2540 SD3_1.n53 SD3_1.n52 2.7305
R2541 SD3_1.n55 SD3_1.t44 2.7305
R2542 SD3_1.n55 SD3_1.n54 2.7305
R2543 SD3_1.n51 SD3_1.t13 2.7305
R2544 SD3_1.n51 SD3_1.n50 2.7305
R2545 SD3_1.n49 SD3_1.t55 2.7305
R2546 SD3_1.n49 SD3_1.n48 2.7305
R2547 SD3_1.n44 SD3_1.t62 2.7305
R2548 SD3_1.n44 SD3_1.n43 2.7305
R2549 SD3_1.n42 SD3_1.t47 2.7305
R2550 SD3_1.n42 SD3_1.n41 2.7305
R2551 SD3_1.n37 SD3_1.t26 2.7305
R2552 SD3_1.n37 SD3_1.n36 2.7305
R2553 SD3_1.n32 SD3_1.t59 2.7305
R2554 SD3_1.n32 SD3_1.n31 2.7305
R2555 SD3_1.n27 SD3_1.t15 2.7305
R2556 SD3_1.n27 SD3_1.n26 2.7305
R2557 SD3_1.n22 SD3_1.t49 2.7305
R2558 SD3_1.n22 SD3_1.n21 2.7305
R2559 SD3_1.n17 SD3_1.t23 2.7305
R2560 SD3_1.n17 SD3_1.n16 2.7305
R2561 SD3_1.n7 SD3_1.t20 2.7305
R2562 SD3_1.n7 SD3_1.n6 2.7305
R2563 SD3_1.n5 SD3_1.t38 2.7305
R2564 SD3_1.n5 SD3_1.n4 2.7305
R2565 SD3_1.n3 SD3_1.t28 2.7305
R2566 SD3_1.n3 SD3_1.n2 2.7305
R2567 SD3_1.n1 SD3_1.t52 2.7305
R2568 SD3_1.n1 SD3_1.n0 2.7305
R2569 SD3_1.n112 SD3_1.t8 2.7305
R2570 SD3_1.n112 SD3_1.n111 2.7305
R2571 SD3_1.n56 SD3_1.n53 2.5571
R2572 SD3_1.n120 SD3_1.n119 2.55706
R2573 SD3_1.n102 SD3_1.t7 2.40707
R2574 SD3_1.n12 SD3_1.t58 2.40704
R2575 SD3_1.n108 SD3_1.n107 2.24937
R2576 SD3_1.n104 SD3_1.n103 2.24505
R2577 SD3_1.n62 SD3_1.n61 2.24478
R2578 SD3_1.n68 SD3_1.n67 2.24478
R2579 SD3_1.n75 SD3_1.n74 1.49476
R2580 SD3_1.n87 SD3_1.n25 1.49463
R2581 SD3_1.n115 SD3_1.n114 1.49463
R2582 SD3_1.n81 SD3_1.n35 1.49463
R2583 SD3_1.n90 SD3_1.n20 1.49463
R2584 SD3_1.n69 SD3_1.n47 1.49439
R2585 SD3_1.n84 SD3_1.n30 1.49439
R2586 SD3_1.n78 SD3_1.n40 1.49439
R2587 SD3_1.n93 SD3_1.n15 1.49439
R2588 SD3_1.n96 SD3_1.n10 1.49439
R2589 SD3_1.n40 SD3_1.n39 1.43788
R2590 SD3_1.n74 SD3_1.n73 1.43788
R2591 SD3_1.n10 SD3_1.n9 1.43741
R2592 SD3_1.n25 SD3_1.n24 1.43741
R2593 SD3_1.n30 SD3_1.n29 1.43741
R2594 SD3_1.n47 SD3_1.n46 1.43741
R2595 SD3_1.n20 SD3_1.n19 1.43705
R2596 SD3_1.n107 SD3_1.n106 1.43694
R2597 SD3_1.n35 SD3_1.n34 1.43694
R2598 SD3_1.n67 SD3_1.n66 1.43694
R2599 SD3_1.n15 SD3_1.n14 1.43673
R2600 SD3_1.n61 SD3_1.n60 1.43673
R2601 SD3_1.n113 SD3_1.n112 1.42872
R2602 SD3_1.n103 SD3_1.n102 1.01023
R2603 SD3_1.n108 SD3_1.n104 0.593824
R2604 SD3_1.n57 SD3_1.n56 0.593282
R2605 SD3_1.n69 SD3_1.n68 0.586829
R2606 SD3_1.n99 SD3_1.n98 0.583544
R2607 SD3_1.n63 SD3_1.n62 0.581823
R2608 SD3_1.n78 SD3_1.n77 0.579925
R2609 SD3_1.n121 SD3_1.n120 0.577695
R2610 SD3_1.n93 SD3_1.n92 0.577272
R2611 SD3_1.n84 SD3_1.n83 0.576023
R2612 SD3_1.n90 SD3_1.n89 0.575664
R2613 SD3_1.n96 SD3_1.n95 0.575142
R2614 SD3_1.n81 SD3_1.n80 0.573011
R2615 SD3_1.n87 SD3_1.n86 0.572285
R2616 SD3_1.n115 SD3_1.n110 0.571741
R2617 SD3_1.n75 SD3_1.n71 0.569825
R2618 SD3_1.n113 SD3_1 0.0644679
R2619 SD3_1.n71 SD3_1.n70 0.0254398
R2620 SD3_1.n92 SD3_1.n91 0.0254398
R2621 SD3_1 SD3_1.n121 0.0243554
R2622 SD3_1.n80 SD3_1.n79 0.0232711
R2623 SD3_1.n98 SD3_1.n97 0.0232711
R2624 SD3_1.n110 SD3_1.n109 0.0232711
R2625 SD3_1.n88 SD3_1.n87 0.0218667
R2626 SD3_1.n86 SD3_1.n85 0.0211024
R2627 SD3_1.n95 SD3_1.n94 0.0211024
R2628 SD3_1.n82 SD3_1.n81 0.0200598
R2629 SD3_1.n77 SD3_1.n76 0.0200181
R2630 SD3_1.n76 SD3_1.n75 0.0190332
R2631 SD3_1.n83 SD3_1.n82 0.0189337
R2632 SD3_1.n85 SD3_1.n84 0.0186111
R2633 SD3_1.n94 SD3_1.n93 0.0178882
R2634 SD3_1.n89 SD3_1.n88 0.0178494
R2635 SD3_1.n58 SD3_1.n57 0.0166884
R2636 SD3_1.n68 SD3_1.n64 0.0166884
R2637 SD3_1.n79 SD3_1.n78 0.0157195
R2638 SD3_1.n97 SD3_1.n96 0.0157195
R2639 SD3_1.n62 SD3_1.n58 0.0156041
R2640 SD3_1.n64 SD3_1.n63 0.0156041
R2641 SD3_1.n104 SD3_1.n100 0.0150649
R2642 SD3_1 SD3_1.n115 0.0143027
R2643 SD3_1.n70 SD3_1.n69 0.0142737
R2644 SD3_1.n91 SD3_1.n90 0.0135538
R2645 SD3_1.n114 SD3_1.n113 0.00977503
R2646 SD3_1.n109 SD3_1.n108 0.00641934
R2647 SD3_1.n100 SD3_1.n99 0.00592169
R2648 b6.n8 b6.n7 64.4419
R2649 b6.n31 b6.n24 51.1109
R2650 b6.n25 b6.t44 50.6807
R2651 b6.n23 b6.n22 49.8352
R2652 b6.n35 b6.t24 47.9333
R2653 b6.n5 b6.t14 40.2611
R2654 b6.n0 b6.t37 39.8961
R2655 b6.n43 b6.n42 33.0652
R2656 b6.n44 b6.n43 31.6402
R2657 b6.n20 b6.n19 30.5682
R2658 b6.n4 b6.n3 26.0261
R2659 b6.n2 b6.n1 25.6611
R2660 b6.n11 b6.t6 24.8545
R2661 b6.n22 b6.t42 24.5042
R2662 b6.n7 b6.t2 23.0349
R2663 b6.t24 b6.t39 21.6159
R2664 b6.t10 b6.t26 21.5355
R2665 b6.t6 b6.t25 21.5355
R2666 b6.t40 b6.t11 21.5355
R2667 b6.t14 b6.t43 21.1705
R2668 b6.t37 b6.t18 21.1705
R2669 b6.t17 b6.t45 21.1705
R2670 b6.t36 b6.t16 21.1705
R2671 b6.n9 b6.t32 18.5039
R2672 b6.n36 b6.t19 14.6735
R2673 b6.n39 b6.t46 14.6735
R2674 b6.n43 b6.t10 14.6735
R2675 b6.n13 b6.t48 14.4545
R2676 b6.n16 b6.t30 14.4545
R2677 b6.n19 b6.t40 14.4545
R2678 b6.n22 b6.t23 14.3815
R2679 b6.n23 b6.t4 14.3815
R2680 b6.n24 b6.t29 14.3815
R2681 b6.n7 b6.t15 14.3085
R2682 b6.n8 b6.t12 14.3085
R2683 b6.n2 b6.t17 14.2355
R2684 b6.n3 b6.t36 14.2355
R2685 b6.n11 b6.t49 13.9435
R2686 b6.n12 b6.t27 13.9435
R2687 b6.n17 b6.t8 13.9435
R2688 b6.n18 b6.t35 13.9435
R2689 b6.n0 b6.t28 13.7975
R2690 b6.n1 b6.t41 13.7975
R2691 b6.n35 b6.t50 13.7245
R2692 b6.n42 b6.t31 13.7245
R2693 b6.n5 b6.t9 13.4325
R2694 b6.n4 b6.t38 13.4325
R2695 b6.n33 b6.t22 12.1915
R2696 b6.n34 b6.t3 12.1915
R2697 b6.n40 b6.t5 12.0455
R2698 b6.t31 b6.n41 12.0455
R2699 b6.n40 b6.t7 11.8265
R2700 b6.n41 b6.t33 11.8265
R2701 b6.n33 b6.t21 11.6805
R2702 b6.t50 b6.n34 11.6805
R2703 b6.n27 b6.t1 11.6029
R2704 b6.n1 b6.n0 11.5035
R2705 b6.n3 b6.n2 11.5035
R2706 b6.n36 b6.n35 11.1652
R2707 b6.n39 b6.n36 11.1652
R2708 b6.n42 b6.n39 11.1652
R2709 b6.t46 b6.n38 11.0965
R2710 b6.n14 b6.t20 10.8045
R2711 b6.n15 b6.t47 10.8045
R2712 b6.t30 b6.n15 10.7315
R2713 b6.n37 b6.t34 10.4395
R2714 b6.n38 b6.t13 10.4395
R2715 b6.n38 b6.n37 10.4005
R2716 b6.n12 b6.n11 10.4005
R2717 b6.n13 b6.n12 10.4005
R2718 b6.n16 b6.n13 10.4005
R2719 b6.n17 b6.n16 10.4005
R2720 b6.n18 b6.n17 10.4005
R2721 b6.n19 b6.n18 10.4005
R2722 b6.n24 b6.n23 10.1232
R2723 b6.n27 b6.t0 9.49371
R2724 b6.n15 b6.n14 8.93226
R2725 b6.n41 b6.n40 8.53084
R2726 b6.n34 b6.n33 7.66919
R2727 b6.n31 b6.n30 6.19053
R2728 b6.n6 b6.n5 5.28339
R2729 b6.n10 b6.n6 5.02841
R2730 b6.n9 b6.n8 4.53153
R2731 b6.n29 b6.n28 4.5305
R2732 b6.n10 b6.n9 3.85224
R2733 b6.n6 b6.n4 3.74655
R2734 b6.n28 b6.n27 3.63044
R2735 b6.n20 b6.n10 2.50672
R2736 b6.n29 b6.n26 2.2505
R2737 b6.n21 b6.n20 1.74245
R2738 b6.n46 b6.n45 1.50779
R2739 b6.n46 b6.n31 1.35684
R2740 b6.n28 b6 0.0263621
R2741 b6 b6.n21 0.0166901
R2742 b6 b6.n26 0.00567241
R2743 b6.n26 b6.n25 0.00360345
R2744 b6.n45 b6.n32 0.00355446
R2745 b6.n30 b6.n29 0.0035
R2746 b6.n45 b6.n44 0.00227316
R2747 b6 b6.n46 0.00137379
R2748 OUT-.n261 OUT-.t160 27.5082
R2749 OUT-.n160 OUT-.t102 18.6921
R2750 OUT-.n86 OUT-.t166 18.1625
R2751 OUT-.n32 OUT-.t146 17.9053
R2752 OUT-.n22 OUT-.t128 17.7975
R2753 OUT-.n30 OUT-.t98 17.7975
R2754 OUT-.n107 OUT-.t150 17.3759
R2755 OUT-.n51 OUT-.t152 17.0653
R2756 OUT-.n192 OUT-.t100 16.8013
R2757 OUT-.n46 OUT-.t172 16.6295
R2758 OUT-.n48 OUT-.t122 16.6295
R2759 OUT-.n62 OUT-.t130 16.5565
R2760 OUT-.n33 OUT-.t132 16.0963
R2761 OUT-.n162 OUT-.t136 15.9834
R2762 OUT-.n262 OUT-.t120 15.5061
R2763 OUT-.n268 OUT-.t178 14.8228
R2764 OUT-.n65 OUT-.t134 14.5125
R2765 OUT-.n256 OUT-.t114 14.3746
R2766 OUT-.n67 OUT-.t164 14.3665
R2767 OUT-.n70 OUT-.t110 14.3665
R2768 OUT-.n111 OUT-.t126 14.3665
R2769 OUT-.n171 OUT-.t112 13.5635
R2770 OUT-.n119 OUT-.t116 12.7025
R2771 OUT-.n130 OUT-.t174 12.5565
R2772 OUT-.n125 OUT-.t144 12.4105
R2773 OUT-.n143 OUT-.t154 12.3279
R2774 OUT-.n206 OUT-.t104 12.1185
R2775 OUT-.n143 OUT-.t148 11.6643
R2776 OUT-.n125 OUT-.t140 11.4615
R2777 OUT-.n130 OUT-.t168 11.3155
R2778 OUT-.n119 OUT-.t108 11.1695
R2779 OUT-.n227 OUT-.t142 10.6585
R2780 OUT-.n10 OUT-.t118 10.5855
R2781 OUT-.n227 OUT-.t106 10.5125
R2782 OUT-.n107 OUT-.t176 10.2935
R2783 OUT-.n251 OUT-.t170 9.9285
R2784 OUT-.n160 OUT-.t156 9.9285
R2785 OUT-.n99 OUT-.n98 9.56292
R2786 OUT-.n37 OUT-.n35 9.14299
R2787 OUT-.n206 OUT-.t158 9.0525
R2788 OUT-.n245 OUT-.t96 8.54636
R2789 OUT-.n239 OUT-.t21 8.54439
R2790 OUT-.n245 OUT-.t15 8.50912
R2791 OUT-.n275 OUT-.t125 8.4005
R2792 OUT-.n273 OUT-.t171 8.4005
R2793 OUT-.n251 OUT-.t124 7.7385
R2794 OUT-.n10 OUT-.t162 7.6655
R2795 OUT-.n262 OUT-.n261 7.06268
R2796 OUT-.n26 OUT-.n25 6.58106
R2797 OUT-.n127 OUT-.t145 6.17646
R2798 OUT-.n128 OUT-.t141 6.14704
R2799 OUT-.n209 OUT-.t83 6.12938
R2800 OUT-.n265 OUT-.t161 6.1271
R2801 OUT-.n49 OUT-.t123 6.12579
R2802 OUT-.n210 OUT-.t79 6.11154
R2803 OUT-.n224 OUT-.t87 6.07519
R2804 OUT-.n68 OUT-.t165 6.07285
R2805 OUT-.n224 OUT-.t76 6.07152
R2806 OUT-.n198 OUT-.t88 6.03932
R2807 OUT-.n177 OUT-.n174 6.02244
R2808 OUT-.n223 OUT-.t89 6.00521
R2809 OUT-.n248 OUT-.n247 5.9303
R2810 OUT-.n220 OUT-.t80 5.8805
R2811 OUT-.n199 OUT-.t85 5.8805
R2812 OUT-.n213 OUT-.t77 5.8805
R2813 OUT-.n211 OUT-.n210 5.74421
R2814 OUT- OUT-.n275 5.73903
R2815 OUT-.n258 OUT-.n257 5.5964
R2816 OUT-.n7 OUT-.t19 5.2505
R2817 OUT-.n15 OUT-.t72 5.2505
R2818 OUT-.n15 OUT-.t119 5.2505
R2819 OUT-.n12 OUT-.t9 5.2505
R2820 OUT-.n12 OUT-.t163 5.2505
R2821 OUT-.n1 OUT-.t14 5.2505
R2822 OUT-.n0 OUT-.t41 5.2505
R2823 OUT-.n195 OUT-.n194 5.06613
R2824 OUT-.n261 OUT-.t138 4.3805
R2825 OUT-.n234 OUT-.t6 4.36508
R2826 OUT-.n256 OUT-.t115 4.29173
R2827 OUT-.n268 OUT-.t179 4.22806
R2828 OUT-.n269 OUT-.t57 4.20189
R2829 OUT-.n234 OUT-.t10 4.201
R2830 OUT-.n271 OUT-.t26 4.15013
R2831 OUT-.n257 OUT-.t91 4.1302
R2832 OUT-.n120 OUT-.n119 4.0005
R2833 OUT-.n126 OUT-.n125 4.0005
R2834 OUT-.n131 OUT-.n130 4.0005
R2835 OUT-.n145 OUT-.n143 4.0005
R2836 OUT-.n161 OUT-.n160 4.0005
R2837 OUT-.n108 OUT-.n107 4.0005
R2838 OUT-.n207 OUT-.n206 4.0005
R2839 OUT-.n229 OUT-.n227 4.0005
R2840 OUT-.n11 OUT-.n10 4.0005
R2841 OUT-.n252 OUT-.n251 4.0005
R2842 OUT-.n263 OUT-.n262 4.0005
R2843 OUT-.n187 OUT-.n186 3.74421
R2844 OUT-.n141 OUT-.n138 3.71646
R2845 OUT-.n21 OUT-.n18 3.6527
R2846 OUT-.n153 OUT-.n152 3.65144
R2847 OUT-.n189 OUT-.n188 3.64267
R2848 OUT-.n75 OUT-.n74 3.62822
R2849 OUT-.n233 OUT-.n100 3.57702
R2850 OUT-.n270 OUT-.n267 3.57312
R2851 OUT-.n187 OUT-.n181 3.55437
R2852 OUT-.n190 OUT-.n103 3.53697
R2853 OUT-.n173 OUT-.n169 3.51226
R2854 OUT-.n167 OUT-.n159 3.50854
R2855 OUT-.n117 OUT-.n116 3.47247
R2856 OUT-.n232 OUT-.n231 3.47027
R2857 OUT-.n106 OUT-.t177 3.46533
R2858 OUT-.n87 OUT-.n85 3.45237
R2859 OUT-.n124 OUT-.n123 3.44226
R2860 OUT-.n186 OUT-.n183 3.42242
R2861 OUT-.n52 OUT-.n44 3.41785
R2862 OUT-.n122 OUT-.n121 3.41123
R2863 OUT-.n63 OUT-.n61 3.40581
R2864 OUT-.n134 OUT-.n133 3.40419
R2865 OUT-.n82 OUT-.n81 3.40162
R2866 OUT-.n47 OUT-.n45 3.39579
R2867 OUT-.n177 OUT-.n176 3.39116
R2868 OUT-.n240 OUT-.n6 3.38977
R2869 OUT-.n117 OUT-.n114 3.38766
R2870 OUT-.n218 OUT-.n200 3.3856
R2871 OUT-.n208 OUT-.n204 3.38009
R2872 OUT-.n98 OUT-.n41 3.37847
R2873 OUT-.n82 OUT-.n79 3.36743
R2874 OUT-.n264 OUT-.n253 3.3665
R2875 OUT-.n146 OUT-.n142 3.36165
R2876 OUT-.n218 OUT-.n201 3.35805
R2877 OUT-.n230 OUT-.n226 3.35805
R2878 OUT-.n6 OUT-.t73 3.35317
R2879 OUT-.n230 OUT-.n225 3.35254
R2880 OUT-.n186 OUT-.n185 3.34851
R2881 OUT-.n66 OUT-.n64 3.34285
R2882 OUT-.n112 OUT-.n105 3.34109
R2883 OUT-.n240 OUT-.n239 3.33961
R2884 OUT-.n13 OUT-.n12 3.33223
R2885 OUT-.n91 OUT-.n88 3.32708
R2886 OUT-.n71 OUT-.n63 3.31948
R2887 OUT-.n260 OUT-.n259 3.31879
R2888 OUT-.n172 OUT-.n170 3.31638
R2889 OUT-.n208 OUT-.n203 3.31581
R2890 OUT-.n197 OUT-.n196 3.3125
R2891 OUT-.n271 OUT-.n270 3.29517
R2892 OUT-.n250 OUT-.n0 3.29336
R2893 OUT-.n212 OUT-.n202 3.2909
R2894 OUT-.n222 OUT-.n101 3.2783
R2895 OUT-.n83 OUT-.n82 3.27278
R2896 OUT-.n258 OUT-.n255 3.26657
R2897 OUT-.n249 OUT-.n1 3.23175
R2898 OUT-.n6 OUT-.t71 3.20968
R2899 OUT-.n235 OUT-.n233 3.20101
R2900 OUT-.n93 OUT-.n92 3.1505
R2901 OUT-.n76 OUT-.n58 3.1505
R2902 OUT-.n77 OUT-.n56 3.1505
R2903 OUT-.n84 OUT-.n54 3.1505
R2904 OUT-.n97 OUT-.n42 3.1505
R2905 OUT-.n35 OUT-.n34 3.1505
R2906 OUT-.n37 OUT-.n36 3.1505
R2907 OUT-.n21 OUT-.n20 3.1505
R2908 OUT-.n25 OUT-.n24 3.1505
R2909 OUT-.n29 OUT-.n28 3.1505
R2910 OUT-.n193 OUT-.n191 3.1505
R2911 OUT-.n148 OUT-.n147 3.1505
R2912 OUT-.n153 OUT-.n150 3.1505
R2913 OUT-.n141 OUT-.n140 3.1505
R2914 OUT-.n166 OUT-.n165 3.1505
R2915 OUT-.n178 OUT-.n157 3.1505
R2916 OUT-.n180 OUT-.n136 3.1505
R2917 OUT-.n16 OUT-.n15 3.1505
R2918 OUT-.n238 OUT-.n7 3.1505
R2919 OUT-.n242 OUT-.n3 3.1505
R2920 OUT-.n26 OUT-.n21 3.14562
R2921 OUT-.n83 OUT-.n77 2.93789
R2922 OUT-.n241 OUT-.n240 2.82033
R2923 OUT-.n84 OUT-.n83 2.75648
R2924 OUT-.n3 OUT-.t74 2.7305
R2925 OUT-.n3 OUT-.n2 2.7305
R2926 OUT-.n41 OUT-.t36 2.7305
R2927 OUT-.n41 OUT-.t35 2.7305
R2928 OUT-.n42 OUT-.t34 2.7305
R2929 OUT-.n42 OUT-.t30 2.7305
R2930 OUT-.n85 OUT-.t8 2.7305
R2931 OUT-.n85 OUT-.t167 2.7305
R2932 OUT-.n92 OUT-.t32 2.7305
R2933 OUT-.n92 OUT-.t29 2.7305
R2934 OUT-.n88 OUT-.t31 2.7305
R2935 OUT-.n88 OUT-.t33 2.7305
R2936 OUT-.n54 OUT-.t59 2.7305
R2937 OUT-.n54 OUT-.n53 2.7305
R2938 OUT-.n79 OUT-.t58 2.7305
R2939 OUT-.n79 OUT-.n78 2.7305
R2940 OUT-.n81 OUT-.t27 2.7305
R2941 OUT-.n81 OUT-.n80 2.7305
R2942 OUT-.n56 OUT-.t60 2.7305
R2943 OUT-.n56 OUT-.n55 2.7305
R2944 OUT-.n58 OUT-.t7 2.7305
R2945 OUT-.n58 OUT-.n57 2.7305
R2946 OUT-.n74 OUT-.t67 2.7305
R2947 OUT-.n74 OUT-.n73 2.7305
R2948 OUT-.n60 OUT-.t111 2.7305
R2949 OUT-.n60 OUT-.n59 2.7305
R2950 OUT-.n61 OUT-.t182 2.7305
R2951 OUT-.n61 OUT-.t131 2.7305
R2952 OUT-.n64 OUT-.t135 2.7305
R2953 OUT-.n44 OUT-.t153 2.7305
R2954 OUT-.n44 OUT-.n43 2.7305
R2955 OUT-.n45 OUT-.t173 2.7305
R2956 OUT-.n36 OUT-.t52 2.7305
R2957 OUT-.n36 OUT-.t147 2.7305
R2958 OUT-.n34 OUT-.t94 2.7305
R2959 OUT-.n34 OUT-.t133 2.7305
R2960 OUT-.n28 OUT-.t99 2.7305
R2961 OUT-.n28 OUT-.n27 2.7305
R2962 OUT-.n18 OUT-.t44 2.7305
R2963 OUT-.n18 OUT-.n17 2.7305
R2964 OUT-.n20 OUT-.t51 2.7305
R2965 OUT-.n20 OUT-.n19 2.7305
R2966 OUT-.n24 OUT-.t129 2.7305
R2967 OUT-.n24 OUT-.n23 2.7305
R2968 OUT-.n191 OUT-.t16 2.7305
R2969 OUT-.n191 OUT-.t101 2.7305
R2970 OUT-.n114 OUT-.t42 2.7305
R2971 OUT-.n114 OUT-.n113 2.7305
R2972 OUT-.n116 OUT-.t25 2.7305
R2973 OUT-.n116 OUT-.n115 2.7305
R2974 OUT-.n183 OUT-.t69 2.7305
R2975 OUT-.n183 OUT-.n182 2.7305
R2976 OUT-.n185 OUT-.t47 2.7305
R2977 OUT-.n185 OUT-.n184 2.7305
R2978 OUT-.n121 OUT-.t109 2.7305
R2979 OUT-.n123 OUT-.t117 2.7305
R2980 OUT-.n133 OUT-.t169 2.7305
R2981 OUT-.n133 OUT-.n132 2.7305
R2982 OUT-.n136 OUT-.t175 2.7305
R2983 OUT-.n136 OUT-.n135 2.7305
R2984 OUT-.n147 OUT-.t49 2.7305
R2985 OUT-.n147 OUT-.t155 2.7305
R2986 OUT-.n142 OUT-.t56 2.7305
R2987 OUT-.n142 OUT-.t149 2.7305
R2988 OUT-.n152 OUT-.t37 2.7305
R2989 OUT-.n152 OUT-.n151 2.7305
R2990 OUT-.n150 OUT-.t46 2.7305
R2991 OUT-.n150 OUT-.n149 2.7305
R2992 OUT-.n138 OUT-.t65 2.7305
R2993 OUT-.n138 OUT-.n137 2.7305
R2994 OUT-.n140 OUT-.t22 2.7305
R2995 OUT-.n140 OUT-.n139 2.7305
R2996 OUT-.n157 OUT-.t24 2.7305
R2997 OUT-.n157 OUT-.n156 2.7305
R2998 OUT-.n169 OUT-.t18 2.7305
R2999 OUT-.n169 OUT-.n168 2.7305
R3000 OUT-.n170 OUT-.t64 2.7305
R3001 OUT-.n170 OUT-.t113 2.7305
R3002 OUT-.n165 OUT-.t157 2.7305
R3003 OUT-.n165 OUT-.t103 2.7305
R3004 OUT-.n159 OUT-.t137 2.7305
R3005 OUT-.n159 OUT-.n158 2.7305
R3006 OUT-.n176 OUT-.t3 2.7305
R3007 OUT-.n176 OUT-.n175 2.7305
R3008 OUT-.n105 OUT-.t127 2.7305
R3009 OUT-.n105 OUT-.n104 2.7305
R3010 OUT-.n103 OUT-.t55 2.7305
R3011 OUT-.n103 OUT-.n102 2.7305
R3012 OUT-.n196 OUT-.t81 2.7305
R3013 OUT-.n204 OUT-.t105 2.7305
R3014 OUT-.n203 OUT-.t159 2.7305
R3015 OUT-.n202 OUT-.t82 2.7305
R3016 OUT-.n201 OUT-.t75 2.7305
R3017 OUT-.n200 OUT-.t84 2.7305
R3018 OUT-.n101 OUT-.t78 2.7305
R3019 OUT-.n226 OUT-.t143 2.7305
R3020 OUT-.n225 OUT-.t107 2.7305
R3021 OUT-.n5 OUT-.t93 2.7305
R3022 OUT-.n5 OUT-.n4 2.7305
R3023 OUT-.n255 OUT-.n254 2.7305
R3024 OUT-.n259 OUT-.t121 2.7305
R3025 OUT-.n253 OUT-.t139 2.7305
R3026 OUT-.n267 OUT-.t5 2.7305
R3027 OUT-.n267 OUT-.n266 2.7305
R3028 OUT-.n29 OUT-.n26 2.56342
R3029 OUT-.n76 OUT-.n75 2.52272
R3030 OUT-.n270 OUT-.n269 2.48586
R3031 OUT-.n188 OUT-.n117 2.2505
R3032 OUT-.n232 OUT-.n223 2.2505
R3033 OUT-.n215 OUT-.t90 2.05255
R3034 OUT-.n75 OUT-.n72 2.04187
R3035 OUT-.n216 OUT-.n215 1.94696
R3036 OUT-.n233 OUT-.n232 1.93866
R3037 OUT-.n108 OUT-.n106 1.85121
R3038 OUT-.n215 OUT-.t86 1.76935
R3039 OUT-.n167 OUT-.n166 1.59579
R3040 OUT-.n100 OUT-.n99 1.54309
R3041 OUT-.n173 OUT-.n172 1.50579
R3042 OUT-.n241 OUT-.n5 1.43159
R3043 OUT-.n72 OUT-.n60 1.42496
R3044 OUT-.n106 OUT-.t151 1.39688
R3045 OUT-.n96 OUT-.n95 1.35988
R3046 OUT-.n236 OUT-.n16 1.25562
R3047 OUT-.n94 OUT-.n87 1.04863
R3048 OUT-.n272 OUT-.n271 1.04839
R3049 OUT-.n243 OUT-.n242 1.04638
R3050 OUT-.n154 OUT-.n148 1.02685
R3051 OUT-.n180 OUT-.n179 1.02681
R3052 OUT-.n190 OUT-.n189 0.955153
R3053 OUT-.n194 OUT-.n193 0.945859
R3054 OUT-.n221 OUT-.n220 0.84268
R3055 OUT-.n214 OUT-.n213 0.840053
R3056 OUT-.n194 OUT-.n190 0.823637
R3057 OUT-.n174 OUT-.n167 0.68553
R3058 OUT-.n174 OUT-.n173 0.681061
R3059 OUT-.n199 OUT-.n198 0.672487
R3060 OUT-.n179 OUT-.n155 0.661654
R3061 OUT-.n155 OUT-.n154 0.658192
R3062 OUT-.n95 OUT-.n94 0.61175
R3063 OUT-.n95 OUT-.n84 0.563
R3064 OUT-.n77 OUT-.n76 0.549186
R3065 OUT-.n189 OUT-.n112 0.532045
R3066 OUT-.n213 OUT-.n212 0.505815
R3067 OUT-.n222 OUT-.n221 0.4919
R3068 OUT-.n257 OUT-.n256 0.482612
R3069 OUT-.n242 OUT-.n241 0.481551
R3070 OUT-.n269 OUT-.n268 0.460088
R3071 OUT-.n272 OUT-.n265 0.4595
R3072 OUT-.n197 OUT-.n195 0.44352
R3073 OUT-.n25 OUT-.n22 0.421942
R3074 OUT-.n235 OUT-.n234 0.420112
R3075 OUT-.n219 OUT-.n218 0.380704
R3076 OUT-.n94 OUT-.n93 0.377076
R3077 OUT-.n193 OUT-.n192 0.374377
R3078 OUT-.n218 OUT-.n217 0.369684
R3079 OUT-.n155 OUT-.n141 0.365692
R3080 OUT-.n35 OUT-.n33 0.364915
R3081 OUT-.n97 OUT-.n96 0.358735
R3082 OUT-.n236 OUT-.n235 0.355045
R3083 OUT-.n38 OUT-.n37 0.344664
R3084 OUT-.n264 OUT-.n263 0.332093
R3085 OUT-.n91 OUT-.n89 0.3305
R3086 OUT-.n265 OUT-.n264 0.3299
R3087 OUT-.n223 OUT-.n222 0.326814
R3088 OUT-.n14 OUT-.n8 0.324154
R3089 OUT-.n91 OUT-.n90 0.321026
R3090 OUT-.n260 OUT-.n258 0.3083
R3091 OUT-.n98 OUT-.n40 0.2905
R3092 OUT-.n198 OUT-.n197 0.287031
R3093 OUT-.n188 OUT-.n187 0.280143
R3094 OUT-.n98 OUT-.n39 0.272167
R3095 OUT-.n212 OUT-.n211 0.266717
R3096 OUT-.n181 OUT-.n180 0.266607
R3097 OUT-.n31 OUT-.n30 0.265864
R3098 OUT-.n209 OUT-.n208 0.264402
R3099 OUT-.n164 OUT-.n163 0.259092
R3100 OUT-.n154 OUT-.n153 0.258613
R3101 OUT-.n179 OUT-.n178 0.258613
R3102 OUT-.n231 OUT-.n230 0.255409
R3103 OUT-.n217 OUT-.n214 0.233471
R3104 OUT-.n220 OUT-.n219 0.233471
R3105 OUT-.n148 OUT-.n146 0.227231
R3106 OUT-.n98 OUT-.n97 0.226104
R3107 OUT-.n178 OUT-.n177 0.223476
R3108 OUT-.n16 OUT-.n14 0.221668
R3109 OUT-.n219 OUT-.n199 0.20592
R3110 OUT-.n217 OUT-.n216 0.20592
R3111 OUT-.n93 OUT-.n91 0.198742
R3112 OUT-.n274 OUT-.n273 0.194429
R3113 OUT-.n31 OUT-.n29 0.193426
R3114 OUT-.n237 OUT-.n236 0.185594
R3115 OUT-.n273 OUT-.n272 0.185121
R3116 OUT-.n239 OUT-.n238 0.183725
R3117 OUT-.n96 OUT-.n52 0.182375
R3118 OUT-.n166 OUT-.n164 0.1805
R3119 OUT-.n72 OUT-.n71 0.180219
R3120 OUT-.n69 OUT-.n68 0.177731
R3121 OUT-.n110 OUT-.n109 0.172572
R3122 OUT-.n275 OUT-.n274 0.1505
R3123 OUT-.n11 OUT-.n9 0.145885
R3124 OUT-.n244 OUT-.n243 0.143357
R3125 OUT-.n67 OUT-.n66 0.143115
R3126 OUT-.n68 OUT-.n67 0.143115
R3127 OUT-.n63 OUT-.n62 0.141731
R3128 OUT-.n238 OUT-.n237 0.141474
R3129 OUT-.n70 OUT-.n69 0.140346
R3130 OUT-.n71 OUT-.n70 0.140346
R3131 OUT-.n120 OUT-.n118 0.140346
R3132 OUT-.n247 OUT-.n246 0.138962
R3133 OUT-.n229 OUT-.n228 0.138858
R3134 OUT-.n87 OUT-.n86 0.138227
R3135 OUT-.n47 OUT-.n46 0.137515
R3136 OUT-.n48 OUT-.n47 0.137515
R3137 OUT-.n49 OUT-.n48 0.137515
R3138 OUT-.n230 OUT-.n229 0.137515
R3139 OUT-.n66 OUT-.n65 0.136734
R3140 OUT-.n50 OUT-.n49 0.136172
R3141 OUT-.n109 OUT-.n108 0.135487
R3142 OUT-.n52 OUT-.n51 0.134808
R3143 OUT-.n112 OUT-.n111 0.134176
R3144 OUT-.n129 OUT-.n128 0.132929
R3145 OUT-.n111 OUT-.n110 0.131529
R3146 OUT-.n164 OUT-.n161 0.131063
R3147 OUT-.n163 OUT-.n162 0.131063
R3148 OUT-.n252 OUT-.n250 0.129461
R3149 OUT-.n131 OUT-.n129 0.129071
R3150 OUT-.n248 OUT-.n244 0.127903
R3151 OUT-.n172 OUT-.n171 0.126253
R3152 OUT-.n208 OUT-.n207 0.1253
R3153 OUT-.n146 OUT-.n145 0.124554
R3154 OUT-.n145 OUT-.n144 0.122122
R3155 OUT-.n207 OUT-.n205 0.1217
R3156 OUT-.n51 OUT-.n50 0.120473
R3157 OUT-.n100 OUT-.n31 0.119848
R3158 OUT-.n249 OUT-.n248 0.118552
R3159 OUT-.n13 OUT-.n11 0.109885
R3160 OUT-.n274 OUT-.n252 0.108227
R3161 OUT-.n247 OUT-.n245 0.106654
R3162 OUT-.n122 OUT-.n120 0.101577
R3163 OUT-.n127 OUT-.n126 0.100935
R3164 OUT-.n126 OUT-.n124 0.0983261
R3165 OUT-.n263 OUT-.n260 0.0860738
R3166 OUT-.n99 OUT-.n38 0.0846936
R3167 OUT-.n134 OUT-.n131 0.0815
R3168 OUT-.n38 OUT-.n32 0.0527857
R3169 OUT-.n231 OUT-.n224 0.046625
R3170 OUT-.n14 OUT-.n13 0.0264615
R3171 OUT-.n181 OUT-.n134 0.0141364
R3172 OUT-.n250 OUT-.n249 0.00634416
R3173 OUT-.n124 OUT-.n122 0.00532143
R3174 OUT-.n128 OUT-.n127 0.00396154
R3175 OUT-.n210 OUT-.n209 0.00168421
R3176 IT.n80 IT.n79 132.385
R3177 IT.n74 IT.n73 131.189
R3178 IT.n0 IT.t39 117.838
R3179 IT.n54 IT.n53 108.54
R3180 IT.n59 IT.n58 106.138
R3181 IT.n48 IT.n47 105.632
R3182 IT.n14 IT.n13 105.126
R3183 IT.n108 IT.n107 104.26
R3184 IT.n37 IT.n36 103.823
R3185 IT.n72 IT.n71 103.823
R3186 IT.n2 IT.n1 103.823
R3187 IT.n4 IT.n3 103.823
R3188 IT.n6 IT.n5 103.823
R3189 IT.n8 IT.n7 103.823
R3190 IT.n10 IT.n9 103.823
R3191 IT.n12 IT.n11 103.823
R3192 IT.n31 IT.n30 103.823
R3193 IT.n29 IT.n28 103.823
R3194 IT.n27 IT.n26 103.823
R3195 IT.n25 IT.n24 103.823
R3196 IT.n23 IT.n22 103.823
R3197 IT.n41 IT.n40 103.823
R3198 IT.n50 IT.n49 103.823
R3199 IT.n63 IT.n62 36.3254
R3200 IT.n71 IT.t58 34.7404
R3201 IT.n52 IT.n50 33.2561
R3202 IT.n42 IT.n41 22.0563
R3203 IT.n38 IT.n37 21.6519
R3204 IT.n73 IT.n72 21.0894
R3205 IT.n107 IT.n106 21.0894
R3206 IT.n1 IT.n0 21.0894
R3207 IT.n3 IT.n2 21.0894
R3208 IT.n5 IT.n4 21.0894
R3209 IT.n7 IT.n6 21.0894
R3210 IT.n9 IT.n8 21.0894
R3211 IT.n11 IT.n10 21.0894
R3212 IT.n13 IT.n12 21.0894
R3213 IT.n32 IT.n31 21.0894
R3214 IT.n30 IT.n29 21.0894
R3215 IT.n28 IT.n27 21.0894
R3216 IT.n26 IT.n25 21.0894
R3217 IT.n24 IT.n23 21.0894
R3218 IT.n22 IT.n21 21.0894
R3219 IT.n40 IT.n39 21.0894
R3220 IT.n49 IT.n48 21.0894
R3221 IT.n0 IT.t53 14.0165
R3222 IT.n1 IT.t26 14.0165
R3223 IT.n2 IT.t27 14.0165
R3224 IT.n3 IT.t35 14.0165
R3225 IT.n4 IT.t31 14.0165
R3226 IT.n5 IT.t68 14.0165
R3227 IT.n6 IT.t60 14.0165
R3228 IT.n7 IT.t34 14.0165
R3229 IT.n8 IT.t36 14.0165
R3230 IT.n9 IT.t71 14.0165
R3231 IT.n10 IT.t25 14.0165
R3232 IT.n11 IT.t52 14.0165
R3233 IT.n12 IT.t42 14.0165
R3234 IT.n13 IT.t29 14.0165
R3235 IT.n31 IT.t63 14.0165
R3236 IT.n30 IT.t62 14.0165
R3237 IT.n29 IT.t40 14.0165
R3238 IT.n28 IT.t46 14.0165
R3239 IT.n27 IT.t61 14.0165
R3240 IT.n26 IT.t69 14.0165
R3241 IT.n25 IT.t32 14.0165
R3242 IT.n24 IT.t33 14.0165
R3243 IT.n23 IT.t59 14.0165
R3244 IT.n22 IT.t66 14.0165
R3245 IT.n21 IT.t30 14.0165
R3246 IT.n39 IT.t24 14.0165
R3247 IT.n40 IT.t51 14.0165
R3248 IT.n41 IT.t37 14.0165
R3249 IT.n107 IT.t64 13.7245
R3250 IT.n106 IT.t28 13.7245
R3251 IT.n62 IT.t75 13.7245
R3252 IT.n48 IT.t41 13.7245
R3253 IT.n49 IT.t49 13.7245
R3254 IT.n50 IT.t72 13.7245
R3255 IT.n37 IT.t45 13.6515
R3256 IT.n36 IT.t44 13.6515
R3257 IT.n79 IT.t43 13.6515
R3258 IT.n71 IT.t47 13.6515
R3259 IT.n72 IT.t38 13.6515
R3260 IT.n73 IT.t48 13.6515
R3261 IT.n108 IT.t55 13.2848
R3262 IT.n38 IT.t50 13.0378
R3263 IT.n81 IT.t14 12.6295
R3264 IT.n80 IT.t0 12.6295
R3265 IT.n54 IT.t12 12.5565
R3266 IT.n58 IT.t4 12.5565
R3267 IT.n75 IT.t8 12.3375
R3268 IT.n74 IT.t10 12.3375
R3269 IT.n59 IT.t2 12.1915
R3270 IT.n47 IT.t74 10.8639
R3271 IT.n43 IT.t73 10.4542
R3272 IT.n20 IT.t54 10.4093
R3273 IT.n52 IT.n51 10.1427
R3274 IT.n16 IT.t65 9.3445
R3275 IT.n53 IT.t6 7.7385
R3276 IT.n57 IT.n56 7.45611
R3277 IT.n100 IT.n99 7.24501
R3278 IT.n53 IT.n52 6.3515
R3279 IT.n64 IT.t3 6.33405
R3280 IT.n47 IT.n46 6.07308
R3281 IT.n82 IT.n80 4.63315
R3282 IT.n67 IT.n63 4.5005
R3283 IT.n57 IT.n54 4.33237
R3284 IT.n76 IT.n74 4.19412
R3285 IT.n82 IT.n81 4.03194
R3286 IT.n58 IT.n57 4.01149
R3287 IT.n76 IT.n75 3.88348
R3288 IT.n99 IT.n96 3.67213
R3289 IT.n90 IT.n38 3.64368
R3290 IT.n44 IT.n42 3.54502
R3291 IT.n44 IT.n43 3.51942
R3292 IT.n86 IT.n85 3.43549
R3293 IT.n77 IT.n70 3.41085
R3294 IT.n35 IT.n18 3.14528
R3295 IT.n96 IT.t19 3.03383
R3296 IT.n96 IT.n95 3.03383
R3297 IT.n98 IT.t20 3.03383
R3298 IT.n98 IT.n97 3.03383
R3299 IT.n94 IT.t18 3.03383
R3300 IT.n94 IT.n93 3.03383
R3301 IT.n92 IT.t17 3.03383
R3302 IT.n92 IT.n91 3.03383
R3303 IT.n18 IT.n17 2.88564
R3304 IT.n46 IT.n45 2.88451
R3305 IT.n109 IT.n108 2.8819
R3306 IT.n100 IT.n94 2.82159
R3307 IT.n101 IT.n92 2.82159
R3308 IT.n99 IT.n98 2.81922
R3309 IT.n85 IT.t15 2.7305
R3310 IT.n85 IT.n84 2.7305
R3311 IT.n70 IT.t11 2.7305
R3312 IT.n70 IT.n69 2.7305
R3313 IT.n56 IT.t13 2.7305
R3314 IT.n56 IT.n55 2.7305
R3315 IT.n17 IT.n16 2.3365
R3316 IT.n35 IT.n34 2.25242
R3317 IT.n87 IT.n86 2.24675
R3318 IT.n15 IT.n14 2.23635
R3319 IT.n34 IT.n33 2.12238
R3320 IT.n77 IT.n76 2.11998
R3321 IT.n33 IT.n32 2.1175
R3322 IT.n61 IT.n60 1.90845
R3323 IT.n102 IT.n101 1.44061
R3324 IT.n78 IT.n77 1.3863
R3325 IT.n83 IT.n82 1.32705
R3326 IT.n33 IT.n20 1.21129
R3327 IT.n68 IT.n67 1.13148
R3328 IT.n90 IT.n89 1.01644
R3329 IT.n110 IT.n104 0.927254
R3330 IT.n60 IT.n59 0.747091
R3331 IT.n103 IT.n35 0.710424
R3332 IT.n63 IT.n61 0.581182
R3333 IT.n101 IT.n100 0.525071
R3334 IT.n103 IT.n102 0.400171
R3335 IT.n89 IT.n68 0.286359
R3336 IT.n89 IT.n88 0.166826
R3337 IT.n102 IT.n90 0.0964132
R3338 IT.n105 IT 0.0795
R3339 IT.n109 IT.n105 0.0275
R3340 IT.n65 IT.n64 0.0250455
R3341 IT.n86 IT.n83 0.0151731
R3342 IT.n104 IT.n103 0.0133571
R3343 IT.n88 IT.n87 0.00905634
R3344 IT.n34 IT.n19 0.00457413
R3345 IT.n67 IT.n66 0.00356818
R3346 IT.n66 IT.n65 0.00356818
R3347 IT IT.n110 0.00340389
R3348 IT.n46 IT.n44 0.0025
R3349 IT.n110 IT.n109 0.00159453
R3350 IT.n18 IT.n15 0.0015
R3351 IT.n87 IT.n78 0.000816901
R3352 OUT6 OUT6.n94 18.695
R3353 OUT6.n126 OUT6.t12 6.52669
R3354 OUT6.n141 OUT6.n95 6.10941
R3355 OUT6.n72 OUT6.n71 4.24612
R3356 OUT6.n50 OUT6.n49 4.22703
R3357 OUT6.n93 OUT6.n92 4.04138
R3358 OUT6.n28 OUT6.n1 3.99956
R3359 OUT6.n83 OUT6.n80 3.71646
R3360 OUT6.n16 OUT6.n13 3.70904
R3361 OUT6.n23 OUT6.n20 3.66108
R3362 OUT6.n39 OUT6.n36 3.66108
R3363 OUT6.n67 OUT6.n64 3.65144
R3364 OUT6.n55 OUT6.n52 3.65144
R3365 OUT6.n126 OUT6.n125 3.52028
R3366 OUT6.n128 OUT6.n121 3.52028
R3367 OUT6.n130 OUT6.n117 3.52028
R3368 OUT6.n132 OUT6.n113 3.52028
R3369 OUT6.n134 OUT6.n109 3.52028
R3370 OUT6.n136 OUT6.n105 3.52028
R3371 OUT6.n138 OUT6.n101 3.52028
R3372 OUT6.n140 OUT6.n97 3.52028
R3373 OUT6.n58 OUT6.n43 3.40302
R3374 OUT6.n75 OUT6.n60 3.40023
R3375 OUT6.n139 OUT6.n99 3.37941
R3376 OUT6.n137 OUT6.n103 3.37941
R3377 OUT6.n135 OUT6.n107 3.37941
R3378 OUT6.n133 OUT6.n111 3.37941
R3379 OUT6.n131 OUT6.n115 3.37941
R3380 OUT6.n129 OUT6.n119 3.37941
R3381 OUT6.n127 OUT6.n123 3.37941
R3382 OUT6.n85 OUT6.n76 3.32729
R3383 OUT6.n16 OUT6.n15 3.1505
R3384 OUT6.n17 OUT6.n11 3.1505
R3385 OUT6.n18 OUT6.n9 3.1505
R3386 OUT6.n23 OUT6.n22 3.1505
R3387 OUT6.n26 OUT6.n5 3.1505
R3388 OUT6.n25 OUT6.n7 3.1505
R3389 OUT6.n27 OUT6.n3 3.1505
R3390 OUT6.n39 OUT6.n38 3.1505
R3391 OUT6.n67 OUT6.n66 3.1505
R3392 OUT6.n72 OUT6.n69 3.1505
R3393 OUT6.n74 OUT6.n62 3.1505
R3394 OUT6.n50 OUT6.n47 3.1505
R3395 OUT6.n55 OUT6.n54 3.1505
R3396 OUT6.n57 OUT6.n45 3.1505
R3397 OUT6.n83 OUT6.n82 3.1505
R3398 OUT6.n84 OUT6.n78 3.1505
R3399 OUT6.n86 OUT6.n41 3.1505
R3400 OUT6.n89 OUT6.n32 3.1505
R3401 OUT6.n88 OUT6.n34 3.1505
R3402 OUT6.n90 OUT6.n30 3.1505
R3403 OUT6.n76 OUT6.n58 2.88513
R3404 OUT6.n94 OUT6.n93 2.83512
R3405 OUT6.n1 OUT6.t46 2.7305
R3406 OUT6.n1 OUT6.n0 2.7305
R3407 OUT6.n3 OUT6.t87 2.7305
R3408 OUT6.n3 OUT6.n2 2.7305
R3409 OUT6.n7 OUT6.t59 2.7305
R3410 OUT6.n7 OUT6.n6 2.7305
R3411 OUT6.n5 OUT6.t1 2.7305
R3412 OUT6.n5 OUT6.n4 2.7305
R3413 OUT6.n9 OUT6.t71 2.7305
R3414 OUT6.n9 OUT6.n8 2.7305
R3415 OUT6.n11 OUT6.t72 2.7305
R3416 OUT6.n11 OUT6.n10 2.7305
R3417 OUT6.n15 OUT6.t49 2.7305
R3418 OUT6.n15 OUT6.n14 2.7305
R3419 OUT6.n13 OUT6.t41 2.7305
R3420 OUT6.n13 OUT6.n12 2.7305
R3421 OUT6.n20 OUT6.t67 2.7305
R3422 OUT6.n20 OUT6.n19 2.7305
R3423 OUT6.n22 OUT6.t85 2.7305
R3424 OUT6.n22 OUT6.n21 2.7305
R3425 OUT6.n30 OUT6.t93 2.7305
R3426 OUT6.n30 OUT6.n29 2.7305
R3427 OUT6.n34 OUT6.t82 2.7305
R3428 OUT6.n34 OUT6.n33 2.7305
R3429 OUT6.n32 OUT6.t63 2.7305
R3430 OUT6.n32 OUT6.n31 2.7305
R3431 OUT6.n36 OUT6.t52 2.7305
R3432 OUT6.n36 OUT6.n35 2.7305
R3433 OUT6.n38 OUT6.t2 2.7305
R3434 OUT6.n38 OUT6.n37 2.7305
R3435 OUT6.n41 OUT6.t39 2.7305
R3436 OUT6.n41 OUT6.n40 2.7305
R3437 OUT6.n60 OUT6.t83 2.7305
R3438 OUT6.n60 OUT6.n59 2.7305
R3439 OUT6.n62 OUT6.t70 2.7305
R3440 OUT6.n62 OUT6.n61 2.7305
R3441 OUT6.n64 OUT6.t5 2.7305
R3442 OUT6.n64 OUT6.n63 2.7305
R3443 OUT6.n66 OUT6.t47 2.7305
R3444 OUT6.n66 OUT6.n65 2.7305
R3445 OUT6.n69 OUT6.t4 2.7305
R3446 OUT6.n69 OUT6.n68 2.7305
R3447 OUT6.n71 OUT6.t66 2.7305
R3448 OUT6.n71 OUT6.n70 2.7305
R3449 OUT6.n43 OUT6.t56 2.7305
R3450 OUT6.n43 OUT6.n42 2.7305
R3451 OUT6.n45 OUT6.t95 2.7305
R3452 OUT6.n45 OUT6.n44 2.7305
R3453 OUT6.n47 OUT6.t91 2.7305
R3454 OUT6.n47 OUT6.n46 2.7305
R3455 OUT6.n49 OUT6.t0 2.7305
R3456 OUT6.n49 OUT6.n48 2.7305
R3457 OUT6.n52 OUT6.t86 2.7305
R3458 OUT6.n52 OUT6.n51 2.7305
R3459 OUT6.n54 OUT6.t76 2.7305
R3460 OUT6.n54 OUT6.n53 2.7305
R3461 OUT6.n78 OUT6.t94 2.7305
R3462 OUT6.n78 OUT6.n77 2.7305
R3463 OUT6.n80 OUT6.t80 2.7305
R3464 OUT6.n80 OUT6.n79 2.7305
R3465 OUT6.n82 OUT6.t81 2.7305
R3466 OUT6.n82 OUT6.n81 2.7305
R3467 OUT6.n92 OUT6.t62 2.7305
R3468 OUT6.n92 OUT6.n91 2.7305
R3469 OUT6.n99 OUT6.t19 2.7305
R3470 OUT6.n99 OUT6.n98 2.7305
R3471 OUT6.n103 OUT6.t35 2.7305
R3472 OUT6.n103 OUT6.n102 2.7305
R3473 OUT6.n107 OUT6.t32 2.7305
R3474 OUT6.n107 OUT6.n106 2.7305
R3475 OUT6.n111 OUT6.t16 2.7305
R3476 OUT6.n111 OUT6.n110 2.7305
R3477 OUT6.n115 OUT6.t27 2.7305
R3478 OUT6.n115 OUT6.n114 2.7305
R3479 OUT6.n119 OUT6.t37 2.7305
R3480 OUT6.n119 OUT6.n118 2.7305
R3481 OUT6.n123 OUT6.t23 2.7305
R3482 OUT6.n123 OUT6.n122 2.7305
R3483 OUT6.n125 OUT6.t13 2.7305
R3484 OUT6.n125 OUT6.n124 2.7305
R3485 OUT6.n121 OUT6.t24 2.7305
R3486 OUT6.n121 OUT6.n120 2.7305
R3487 OUT6.n117 OUT6.t15 2.7305
R3488 OUT6.n117 OUT6.n116 2.7305
R3489 OUT6.n113 OUT6.t31 2.7305
R3490 OUT6.n113 OUT6.n112 2.7305
R3491 OUT6.n109 OUT6.t17 2.7305
R3492 OUT6.n109 OUT6.n108 2.7305
R3493 OUT6.n105 OUT6.t33 2.7305
R3494 OUT6.n105 OUT6.n104 2.7305
R3495 OUT6.n101 OUT6.t21 2.7305
R3496 OUT6.n101 OUT6.n100 2.7305
R3497 OUT6.n97 OUT6.t7 2.7305
R3498 OUT6.n97 OUT6.n96 2.7305
R3499 OUT6.n76 OUT6.n75 2.2505
R3500 OUT6.n94 OUT6.n28 2.2505
R3501 OUT6.n17 OUT6.n16 1.08037
R3502 OUT6.n84 OUT6.n83 1.06999
R3503 OUT6.n24 OUT6.n23 0.890115
R3504 OUT6.n56 OUT6.n55 0.87333
R3505 OUT6.n87 OUT6.n39 0.853769
R3506 OUT6.n73 OUT6.n67 0.827481
R3507 OUT6.n27 OUT6.n26 0.682695
R3508 OUT6.n90 OUT6.n89 0.681139
R3509 OUT6.n18 OUT6.n17 0.564306
R3510 OUT6.n26 OUT6.n25 0.511077
R3511 OUT6.n89 OUT6.n88 0.501443
R3512 OUT6.n73 OUT6.n72 0.438262
R3513 OUT6.n141 OUT6.n140 0.417773
R3514 OUT6.n140 OUT6.n139 0.417773
R3515 OUT6.n139 OUT6.n138 0.417773
R3516 OUT6.n138 OUT6.n137 0.417773
R3517 OUT6.n137 OUT6.n136 0.417773
R3518 OUT6.n136 OUT6.n135 0.417773
R3519 OUT6.n135 OUT6.n134 0.417773
R3520 OUT6.n134 OUT6.n133 0.417773
R3521 OUT6.n133 OUT6.n132 0.417773
R3522 OUT6.n132 OUT6.n131 0.417773
R3523 OUT6.n131 OUT6.n130 0.417773
R3524 OUT6.n130 OUT6.n129 0.417773
R3525 OUT6.n129 OUT6.n128 0.417773
R3526 OUT6.n128 OUT6.n127 0.417773
R3527 OUT6.n127 OUT6.n126 0.417773
R3528 OUT6.n87 OUT6.n86 0.416349
R3529 OUT6.n24 OUT6.n18 0.389629
R3530 OUT6.n56 OUT6.n50 0.380241
R3531 OUT6.n85 OUT6.n84 0.257226
R3532 OUT6.n86 OUT6.n85 0.253149
R3533 OUT6.n88 OUT6.n87 0.236538
R3534 OUT6.n74 OUT6.n73 0.220379
R3535 OUT6.n58 OUT6.n57 0.213967
R3536 OUT6.n75 OUT6.n74 0.208465
R3537 OUT6.n28 OUT6.n27 0.207865
R3538 OUT6.n25 OUT6.n24 0.185692
R3539 OUT6.n57 OUT6.n56 0.178802
R3540 OUT6.n93 OUT6.n90 0.164923
R3541 OUT6 OUT6.n141 0.133455
R3542 b6b.n0 b6b.t49 84.0965
R3543 b6b.n17 b6b.t4 74.5586
R3544 b6b.n2 b6b.n1 70.0805
R3545 b6b.n19 b6b.n18 61.2726
R3546 b6b.n7 b6b.t21 58.8447
R3547 b6b.n40 b6b.t47 54.2651
R3548 b6b.n23 b6b.t25 47.5922
R3549 b6b.n13 b6b.n12 45.3788
R3550 b6b.n46 b6b.n45 39.4461
R3551 b6b.n47 b6b.n46 37.6576
R3552 b6b.n31 b6b.n30 33.0652
R3553 b6b.n32 b6b.n31 32.8101
R3554 b6b.n12 b6b.n9 26.5717
R3555 b6b.t40 b6b.t38 23.9755
R3556 b6b.t25 b6b.t24 23.8715
R3557 b6b.n8 b6b.n7 23.854
R3558 b6b.n20 b6b.n19 22.5861
R3559 b6b b6b.t43 19.4018
R3560 b6b.n41 b6b.t34 14.8195
R3561 b6b.n42 b6b.t5 14.8195
R3562 b6b.n46 b6b.t13 14.8195
R3563 b6b.n24 b6b.t14 14.5275
R3564 b6b.n27 b6b.t33 14.5275
R3565 b6b.n31 b6b.t40 14.5275
R3566 b6b.n7 b6b.t11 14.0165
R3567 b6b.n12 b6b.t9 14.0165
R3568 b6b.n0 b6b.t29 14.0165
R3569 b6b.n1 b6b.t46 14.0165
R3570 b6b.n2 b6b.t28 14.0165
R3571 b6b.n8 b6b.t2 13.9428
R3572 b6b.n23 b6b.t17 13.5785
R3573 b6b.n30 b6b.t36 13.5785
R3574 b6b.n13 b6b.t50 13.4138
R3575 b6b.n9 b6b.n8 13.3558
R3576 b6b.n41 b6b.n40 13.3198
R3577 b6b.n42 b6b.n41 13.3198
R3578 b6b.n45 b6b.n42 13.3198
R3579 b6b.n40 b6b.t32 13.2865
R3580 b6b.n45 b6b.t3 13.2865
R3581 b6b.n17 b6b.t39 13.2865
R3582 b6b.n18 b6b.t10 13.2865
R3583 b6b.n19 b6b.t19 13.2865
R3584 b6b.n25 b6b.t12 12.7025
R3585 b6b.n26 b6b.t31 12.7025
R3586 b6b.n18 b6b.n17 12.4464
R3587 b6b.n43 b6b.t22 11.6075
R3588 b6b.t3 b6b.n44 11.6075
R3589 b6b.t33 b6b.n26 11.1695
R3590 b6b.n27 b6b.n24 11.1652
R3591 b6b.n24 b6b.n23 11.1652
R3592 b6b.n30 b6b.n27 11.1652
R3593 b6b.n38 b6b.t41 11.0235
R3594 b6b.n39 b6b.t16 11.0235
R3595 b6b.n5 b6b.t45 11.0235
R3596 b6b.t11 b6b.n6 11.0235
R3597 b6b.n10 b6b.t26 11.0235
R3598 b6b.t9 b6b.n11 11.0235
R3599 b6b.n21 b6b.t23 10.8775
R3600 b6b.n22 b6b.t48 10.8775
R3601 b6b.n28 b6b.t7 10.8045
R3602 b6b.t36 b6b.n29 10.8045
R3603 b6b.n28 b6b.t37 10.7315
R3604 b6b.n29 b6b.t18 10.7315
R3605 b6b.n21 b6b.t42 10.6585
R3606 b6b.t17 b6b.n22 10.6585
R3607 b6b.n38 b6b.t8 10.5125
R3608 b6b.t32 b6b.n39 10.5125
R3609 b6b.n44 b6b.n43 10.26
R3610 b6b.n5 b6b.t15 10.1475
R3611 b6b.n6 b6b.t30 10.1475
R3612 b6b.n10 b6b.t44 10.1475
R3613 b6b.n11 b6b.t27 10.1475
R3614 b6b.n6 b6b.n5 10.1232
R3615 b6b.n43 b6b.t6 9.9285
R3616 b6b.n44 b6b.t35 9.9285
R3617 b6b.n11 b6b.n10 9.73383
R3618 b6b.n36 b6b.n34 9.49418
R3619 b6b.n1 b6b.n0 9.4905
R3620 b6b.n29 b6b.n28 9.4905
R3621 b6b.n36 b6b.n35 9.40022
R3622 b6b.n39 b6b.n38 9.37334
R3623 b6b.n22 b6b.n21 9.0386
R3624 b6b.n26 b6b.n25 8.16394
R3625 b6b.n3 b6b.n2 7.52054
R3626 b6b.n9 b6b.t20 7.0085
R3627 b6b.n49 b6b.n48 4.53085
R3628 b6b.n37 b6b.n36 2.2505
R3629 b6b.n14 b6b.n13 2.13621
R3630 b6b.n33 b6b.n32 2.04965
R3631 b6b.n15 b6b.n14 1.5034
R3632 b6b.n32 b6b.n20 1.40687
R3633 b6b.n49 b6b.n37 1.33542
R3634 b6b.n47 b6b.n33 1.12144
R3635 b6b.n20 b6b.n16 1.00188
R3636 b6b b6b.n49 0.0343961
R3637 b6b.n15 b6b.n3 0.0197857
R3638 b6b.n16 b6b.n15 0.0191429
R3639 b6b b6b.n33 0.0120079
R3640 b6b.n14 b6b.n4 0.00265339
R3641 b6b.n48 b6b.n47 0.00259302
R3642 b6b.n37 b6b 0.00192857
R3643 b2.n0 b2.t3 49.5502
R3644 b2.n10 b2.n9 44.2287
R3645 b2.n9 b2.t2 22.1139
R3646 b2.n12 b2.n10 21.2987
R3647 b2.n6 b2.t6 19.8669
R3648 b2.n11 b2.t1 9.49371
R3649 b2.n11 b2.t0 9.3756
R3650 b2.n4 b2.t4 7.0085
R3651 b2.n10 b2.n8 4.66598
R3652 b2.n8 b2.n7 4.5005
R3653 b2.n12 b2.n11 2.53871
R3654 b2 b2.n0 2.25981
R3655 b2.n9 b2.t5 2.1905
R3656 b2 b2.n12 1.11809
R3657 b2.n5 b2.n4 0.8035
R3658 b2.n6 b2.n5 0.8035
R3659 b2.n7 b2.n6 0.2195
R3660 b2.n0 b2 0.14127
R3661 b2.n3 b2.n2 0.0340106
R3662 b2.n8 b2.n1 0.00371429
R3663 b2.n8 b2.n3 0.00145745
R3664 OUT2.n6 OUT2.n5 17.8839
R3665 OUT2 OUT2.t5 6.00764
R3666 OUT2.n7 OUT2.n0 5.8805
R3667 OUT2.n5 OUT2.n2 4.04862
R3668 OUT2.n7 OUT2.n6 3.51222
R3669 OUT2.n5 OUT2.n4 3.38961
R3670 OUT2.n2 OUT2.t4 2.7305
R3671 OUT2.n2 OUT2.n1 2.7305
R3672 OUT2.n4 OUT2.t1 2.7305
R3673 OUT2.n4 OUT2.n3 2.7305
R3674 OUT2.n6 OUT2 2.31942
R3675 OUT2 OUT2.n7 0.068
R3676 b5b.t24 b5b.n11 75.0723
R3677 b5b.n10 b5b.t23 72.0525
R3678 b5b.n13 b5b.t21 62.2995
R3679 b5b.n14 b5b.n12 47.9184
R3680 b5b.n7 b5b.t8 47.5922
R3681 b5b.n18 b5b.n17 36.7152
R3682 b5b.n12 b5b.t13 24.4555
R3683 b5b.t13 b5b.t24 21.0034
R3684 b5b.t22 b5b.t11 20.7325
R3685 b5b.t14 b5b.t3 20.7325
R3686 b5b.t23 b5b.t12 20.7325
R3687 b5b.n19 b5b.t15 19.1982
R3688 b5b.n11 b5b.n10 14.8925
R3689 b5b.n8 b5b.t18 14.5275
R3690 b5b.n19 b5b.n18 14.5057
R3691 b5b.n13 b5b.t5 14.3815
R3692 b5b.n12 b5b.t10 14.3815
R3693 b5b.n14 b5b.t2 14.3815
R3694 b5b.n15 b5b.t16 14.2355
R3695 b5b.n7 b5b.t19 13.5785
R3696 b5b.n17 b5b.t7 13.5785
R3697 b5b.n11 b5b.t22 11.6075
R3698 b5b.n10 b5b.t14 11.6075
R3699 b5b.n8 b5b.n7 11.1652
R3700 b5b.n17 b5b.n16 11.1652
R3701 b5b.n16 b5b.n8 11.1652
R3702 b5b.n3 b5b.t20 11.0235
R3703 b5b.n4 b5b.t4 11.0235
R3704 b5b.n5 b5b.t9 10.9505
R3705 b5b.t19 b5b.n6 10.9505
R3706 b5b.n5 b5b.t6 10.5855
R3707 b5b.n6 b5b.t17 10.5855
R3708 b5b.n3 b5b.t26 10.5125
R3709 b5b.t7 b5b.n4 10.5125
R3710 b5b.n14 b5b.n13 9.73383
R3711 b5b.n18 b5b.t25 9.7095
R3712 b5b.n2 b5b.n0 9.49418
R3713 b5b.n2 b5b.n1 9.40022
R3714 b5b.n6 b5b.n5 9.37334
R3715 b5b.n4 b5b.n3 9.14749
R3716 b5b b5b.n14 6.02162
R3717 b5b.n15 b5b 4.0055
R3718 b5b b5b.n2 2.25319
R3719 b5b.n16 b5b.n15 0.2925
R3720 b5b b5b.n19 0.224828
R3721 b5b.n16 b5b.n9 0.0735
R3722 OUT5.n65 OUT5.n64 11.1462
R3723 OUT5 OUT5.n46 9.06769
R3724 OUT5.n57 OUT5.n56 6.90515
R3725 OUT5.n62 OUT5.t2 6.48993
R3726 OUT5.n65 OUT5.t0 6.12071
R3727 OUT5.n69 OUT5.n47 6.11137
R3728 OUT5.n42 OUT5.n41 3.88773
R3729 OUT5.n8 OUT5.n7 3.88773
R3730 OUT5.n19 OUT5.n18 3.88773
R3731 OUT5.n31 OUT5.n30 3.80786
R3732 OUT5.n57 OUT5.n55 3.54767
R3733 OUT5.n62 OUT5.n61 3.46159
R3734 OUT5.n66 OUT5.n53 3.46159
R3735 OUT5.n68 OUT5.n49 3.46159
R3736 OUT5.n63 OUT5.n59 3.38137
R3737 OUT5.n67 OUT5.n51 3.38137
R3738 OUT5.n42 OUT5.n39 3.1505
R3739 OUT5.n43 OUT5.n37 3.1505
R3740 OUT5.n44 OUT5.n35 3.1505
R3741 OUT5.n31 OUT5.n28 3.1505
R3742 OUT5.n32 OUT5.n26 3.1505
R3743 OUT5.n33 OUT5.n24 3.1505
R3744 OUT5.n8 OUT5.n5 3.1505
R3745 OUT5.n9 OUT5.n3 3.1505
R3746 OUT5.n10 OUT5.n1 3.1505
R3747 OUT5.n20 OUT5.n14 3.1505
R3748 OUT5.n19 OUT5.n16 3.1505
R3749 OUT5.n21 OUT5.n12 3.1505
R3750 OUT5.n46 OUT5.n22 3.00524
R3751 OUT5.n59 OUT5.t7 2.7305
R3752 OUT5.n59 OUT5.n58 2.7305
R3753 OUT5.n61 OUT5.t3 2.7305
R3754 OUT5.n61 OUT5.n60 2.7305
R3755 OUT5.n55 OUT5.t4 2.7305
R3756 OUT5.n55 OUT5.n54 2.7305
R3757 OUT5.n35 OUT5.t44 2.7305
R3758 OUT5.n35 OUT5.n34 2.7305
R3759 OUT5.n37 OUT5.t19 2.7305
R3760 OUT5.n37 OUT5.n36 2.7305
R3761 OUT5.n39 OUT5.t16 2.7305
R3762 OUT5.n39 OUT5.n38 2.7305
R3763 OUT5.n41 OUT5.t47 2.7305
R3764 OUT5.n41 OUT5.n40 2.7305
R3765 OUT5.n24 OUT5.t31 2.7305
R3766 OUT5.n24 OUT5.n23 2.7305
R3767 OUT5.n26 OUT5.t36 2.7305
R3768 OUT5.n26 OUT5.n25 2.7305
R3769 OUT5.n28 OUT5.t33 2.7305
R3770 OUT5.n28 OUT5.n27 2.7305
R3771 OUT5.n30 OUT5.t23 2.7305
R3772 OUT5.n30 OUT5.n29 2.7305
R3773 OUT5.n1 OUT5.t18 2.7305
R3774 OUT5.n1 OUT5.n0 2.7305
R3775 OUT5.n3 OUT5.t38 2.7305
R3776 OUT5.n3 OUT5.n2 2.7305
R3777 OUT5.n5 OUT5.t39 2.7305
R3778 OUT5.n5 OUT5.n4 2.7305
R3779 OUT5.n7 OUT5.t26 2.7305
R3780 OUT5.n7 OUT5.n6 2.7305
R3781 OUT5.n12 OUT5.t37 2.7305
R3782 OUT5.n12 OUT5.n11 2.7305
R3783 OUT5.n18 OUT5.t40 2.7305
R3784 OUT5.n18 OUT5.n17 2.7305
R3785 OUT5.n16 OUT5.t20 2.7305
R3786 OUT5.n16 OUT5.n15 2.7305
R3787 OUT5.n14 OUT5.t22 2.7305
R3788 OUT5.n14 OUT5.n13 2.7305
R3789 OUT5.n51 OUT5.t5 2.7305
R3790 OUT5.n51 OUT5.n50 2.7305
R3791 OUT5.n53 OUT5.t6 2.7305
R3792 OUT5.n53 OUT5.n52 2.7305
R3793 OUT5.n49 OUT5.t1 2.7305
R3794 OUT5.n49 OUT5.n48 2.7305
R3795 OUT5.n46 OUT5.n45 2.2555
R3796 OUT5.n22 OUT5.n10 0.916077
R3797 OUT5.n44 OUT5.n43 0.826683
R3798 OUT5.n33 OUT5.n32 0.74308
R3799 OUT5.n21 OUT5.n20 0.73453
R3800 OUT5.n10 OUT5.n9 0.733978
R3801 OUT5.n45 OUT5.n44 0.698412
R3802 OUT5.n43 OUT5.n42 0.565394
R3803 OUT5.n32 OUT5.n31 0.565394
R3804 OUT5.n9 OUT5.n8 0.565394
R3805 OUT5.n20 OUT5.n19 0.565394
R3806 OUT5.n64 OUT5.n63 0.379057
R3807 OUT5.n63 OUT5.n62 0.379057
R3808 OUT5.n69 OUT5.n68 0.379057
R3809 OUT5.n68 OUT5.n67 0.379057
R3810 OUT5.n67 OUT5.n66 0.379057
R3811 OUT5.n45 OUT5.n33 0.376378
R3812 OUT5.n66 OUT5.n65 0.370706
R3813 OUT5.n22 OUT5.n21 0.304973
R3814 OUT5 OUT5.n69 0.136892
R3815 OUT5.n64 OUT5.n57 0.00235567
R3816 G2.n1 G2.n0 102.993
R3817 G2.n3 G2.n2 101.566
R3818 G2.n6 G2.n5 99.4048
R3819 G2.n8 G2.n7 99.4048
R3820 G2.n10 G2.n4 70.7294
R3821 G2.n9 G2.n8 39.5325
R3822 G2.n10 G2.n9 39.4595
R3823 G2.n4 G2.n3 37.7091
R3824 G2.n0 G2.t10 29.4988
R3825 G2.n5 G2.t4 29.1477
R3826 G2.t10 G2.t17 23.7985
R3827 G2.t21 G2.t24 23.7985
R3828 G2.t3 G2.t7 23.7985
R3829 G2.t14 G2.t18 23.7985
R3830 G2.t5 G2.t12 23.7985
R3831 G2.t4 G2.t9 23.7985
R3832 G2.t20 G2.t23 23.7985
R3833 G2.t8 G2.t16 23.7985
R3834 G2.t6 G2.t15 23.7985
R3835 G2.t19 G2.t22 23.7985
R3836 G2.n2 G2.n1 16.5048
R3837 G2.n7 G2.n6 16.1537
R3838 G2.n9 G2.t11 13.1405
R3839 G2.n4 G2.t13 13.0675
R3840 G2.t1 G2.n10 13.0675
R3841 G2.n0 G2.t21 12.9945
R3842 G2.n1 G2.t3 12.9945
R3843 G2.n2 G2.t14 12.9945
R3844 G2.n3 G2.t5 12.9945
R3845 G2.n5 G2.t20 12.9945
R3846 G2.n6 G2.t8 12.9945
R3847 G2.n7 G2.t6 12.9945
R3848 G2.n8 G2.t19 12.9945
R3849 G2.n11 G2.t25 12.6295
R3850 G2.n11 G2.t1 11.1695
R3851 G2.n14 G2.n11 4.0005
R3852 G2 G2.n13 3.34309
R3853 G2.n13 G2.t2 2.7305
R3854 G2.n13 G2.n12 2.7305
R3855 G2.n14 G2 0.0935
R3856 G2 G2.n14 0.0065
R3857 SD2_5 SD2_5.n10 4.78409
R3858 SD2_5.n4 SD2_5.n3 3.44212
R3859 SD2_5.n9 SD2_5.n8 3.43911
R3860 SD2_5.n15 SD2_5.n12 3.41246
R3861 SD2_5.n20 SD2_5.n19 3.38757
R3862 SD2_5.n15 SD2_5.n14 3.38387
R3863 SD2_5.n4 SD2_5.n1 3.38278
R3864 SD2_5.n9 SD2_5.n6 3.38274
R3865 SD2_5 SD2_5.n17 3.29941
R3866 SD2_5.n10 SD2_5.n4 2.87871
R3867 SD2_5.n21 SD2_5.n15 2.87758
R3868 SD2_5.n17 SD2_5.t14 2.7305
R3869 SD2_5.n17 SD2_5.n16 2.7305
R3870 SD2_5.n12 SD2_5.t9 2.7305
R3871 SD2_5.n12 SD2_5.n11 2.7305
R3872 SD2_5.n14 SD2_5.t11 2.7305
R3873 SD2_5.n14 SD2_5.n13 2.7305
R3874 SD2_5.n6 SD2_5.t6 2.7305
R3875 SD2_5.n6 SD2_5.n5 2.7305
R3876 SD2_5.n8 SD2_5.t10 2.7305
R3877 SD2_5.n8 SD2_5.n7 2.7305
R3878 SD2_5.n1 SD2_5.t2 2.7305
R3879 SD2_5.n1 SD2_5.n0 2.7305
R3880 SD2_5.n3 SD2_5.t1 2.7305
R3881 SD2_5.n3 SD2_5.n2 2.7305
R3882 SD2_5.n19 SD2_5.t15 2.7305
R3883 SD2_5.n19 SD2_5.n18 2.7305
R3884 SD2_5.n10 SD2_5.n9 2.2505
R3885 SD2_5.n21 SD2_5.n20 2.2505
R3886 SD2_5.n20 SD2_5 0.116906
R3887 SD2_5 SD2_5.n21 0.00283766
R3888 b5.t19 b5.t7 109.68
R3889 b5 b5.t11 51.8095
R3890 b5.n14 b5.n13 48.5408
R3891 b5.n11 b5.t6 28.2458
R3892 b5.n4 b5.t16 25.4465
R3893 b5.t6 b5.t9 21.5355
R3894 b5.t16 b5.t18 21.5355
R3895 b5.n16 b5.t4 20.3746
R3896 b5.n4 b5.t13 14.4545
R3897 b5.n5 b5.t21 14.4545
R3898 b5.n10 b5.t12 14.4545
R3899 b5.n11 b5.n10 14.398
R3900 b5.n13 b5.t23 14.1625
R3901 b5.n14 b5.t10 14.1625
R3902 b5.t26 b5.n6 13.9435
R3903 b5.n9 b5.t20 13.9435
R3904 b5.n12 b5.n11 13.9116
R3905 b5.n13 b5.n12 13.5102
R3906 b5.n15 b5.t25 13.2865
R3907 b5.n7 b5.t26 12.1185
R3908 b5.t20 b5.n8 12.1185
R3909 b5.n5 b5.n4 11.5035
R3910 b5.n9 b5.n6 11.5035
R3911 b5.n6 b5.n5 11.5035
R3912 b5.n10 b5.n9 11.5035
R3913 b5.n15 b5.n14 10.7362
R3914 b5.n0 b5.t22 10.4395
R3915 b5.t7 b5.n1 10.4395
R3916 b5.n2 b5.t19 10.4395
R3917 b5.t4 b5.n3 10.4395
R3918 b5.n2 b5.t5 10.2935
R3919 b5.n0 b5.t8 10.2935
R3920 b5.n1 b5.t17 10.2935
R3921 b5.n3 b5.t15 10.2935
R3922 b5.n12 b5.t14 9.6365
R3923 b5.n17 b5.t0 9.49371
R3924 b5.n1 b5.n0 9.4905
R3925 b5.n3 b5.n2 9.4905
R3926 b5.n7 b5.t3 9.4175
R3927 b5.n8 b5.t24 9.4175
R3928 b5.n17 b5.t1 9.3756
R3929 b5.n8 b5.n7 9.14749
R3930 b5.n18 b5.n16 5.49961
R3931 b5.n16 b5.n15 5.23946
R3932 b5.n11 b5.t2 4.3805
R3933 b5.n18 b5.n17 3.24728
R3934 b5 b5.n18 0.374557
R3935 b4b.n3 b4b.t8 135.346
R3936 b4b.n6 b4b.t12 122.275
R3937 b4b.n7 b4b.t16 87.2463
R3938 b4b.n2 b4b.t10 86.6191
R3939 b4b.n3 b4b.n2 75.3342
R3940 b4b.t12 b4b.t4 68.4445
R3941 b4b.t7 b4b.t3 56.6204
R3942 b4b.n8 b4b.n6 52.2803
R3943 b4b.t10 b4b.t13 41.8693
R3944 b4b.n9 b4b.n8 32.8633
R3945 b4b b4b.t9 19.4226
R3946 b4b.t3 b4b.n3 18.8389
R3947 b4b.n2 b4b.t2 18.7955
R3948 b4b.n6 b4b.t6 18.4057
R3949 b4b.n7 b4b.t11 18.0315
R3950 b4b.n5 b4b.n4 16.0319
R3951 b4b.n1 b4b.n0 15.4944
R3952 b4b.n0 b4b.t15 10.7315
R3953 b4b.n1 b4b.t17 10.7315
R3954 b4b.n0 b4b.t5 9.6365
R3955 b4b.t13 b4b.n1 9.6365
R3956 b4b.n18 b4b.n13 9.49418
R3957 b4b.n17 b4b.n16 9.39762
R3958 b4b.n4 b4b.t18 9.3445
R3959 b4b.n4 b4b.t7 8.9065
R3960 b4b.n5 b4b.t14 8.9065
R3961 b4b.t4 b4b.n5 7.1545
R3962 b4b.n12 b4b.n11 4.5005
R3963 b4b.n8 b4b.n7 3.6505
R3964 b4b.n17 b4b.n15 2.37493
R3965 b4b.n19 b4b.n18 2.2505
R3966 b4b.n19 b4b.n12 0.113387
R3967 b4b.n14 b4b.n12 0.0210063
R3968 b4b.n15 b4b.n14 0.0118924
R3969 b4b.n11 b4b.n9 0.0112067
R3970 b4b b4b.n19 0.00318657
R3971 b4b.n18 b4b.n17 0.0031087
R3972 b4b.n11 b4b.n10 0.0021391
R3973 b4b.n10 b4b 0.00213881
R3974 OUT4.n31 OUT4.n30 15.3782
R3975 OUT4.n32 OUT4.n31 8.93169
R3976 OUT4.n5 OUT4.t10 6.44473
R3977 OUT4.n2 OUT4.n0 6.42383
R3978 OUT4.n2 OUT4.n1 5.8805
R3979 OUT4.n33 OUT4.t11 5.8805
R3980 OUT4.n32 OUT4.t3 5.8805
R3981 OUT4.n6 OUT4.n4 5.8805
R3982 OUT4.n7 OUT4.n3 5.8805
R3983 OUT4.n5 OUT4.t6 5.8805
R3984 OUT4.n27 OUT4.n26 3.85309
R3985 OUT4.n16 OUT4.n15 3.82489
R3986 OUT4.n17 OUT4.n11 3.1505
R3987 OUT4.n16 OUT4.n13 3.1505
R3988 OUT4.n18 OUT4.n9 3.1505
R3989 OUT4.n28 OUT4.n22 3.1505
R3990 OUT4.n27 OUT4.n24 3.1505
R3991 OUT4.n29 OUT4.n20 3.1505
R3992 OUT4.n9 OUT4.t21 2.7305
R3993 OUT4.n9 OUT4.n8 2.7305
R3994 OUT4.n13 OUT4.t0 2.7305
R3995 OUT4.n13 OUT4.n12 2.7305
R3996 OUT4.n11 OUT4.t13 2.7305
R3997 OUT4.n11 OUT4.n10 2.7305
R3998 OUT4.n15 OUT4.t18 2.7305
R3999 OUT4.n15 OUT4.n14 2.7305
R4000 OUT4.n20 OUT4.t12 2.7305
R4001 OUT4.n20 OUT4.n19 2.7305
R4002 OUT4.n24 OUT4.t14 2.7305
R4003 OUT4.n24 OUT4.n23 2.7305
R4004 OUT4.n22 OUT4.t17 2.7305
R4005 OUT4.n22 OUT4.n21 2.7305
R4006 OUT4.n26 OUT4.t1 2.7305
R4007 OUT4.n26 OUT4.n25 2.7305
R4008 OUT4.n31 OUT4.n7 2.72598
R4009 OUT4.n6 OUT4.n5 1.79955
R4010 OUT4 OUT4.n33 1.70642
R4011 OUT4.n30 OUT4.n18 1.02158
R4012 OUT4.n29 OUT4.n28 0.689162
R4013 OUT4.n18 OUT4.n17 0.669768
R4014 OUT4.n33 OUT4.n32 0.599276
R4015 OUT4.n7 OUT4.n6 0.575794
R4016 OUT4.n28 OUT4.n27 0.483385
R4017 OUT4.n17 OUT4.n16 0.474274
R4018 OUT4.n30 OUT4.n29 0.132857
R4019 OUT4 OUT4.n2 0.0205
R4020 b2b b2b.n2 33.3766
R4021 b2b b2b.t5 19.4226
R4022 b2b.n0 b2b.t6 13.1296
R4023 b2b.n1 b2b.t3 10.5977
R4024 b2b.n0 b2b.t4 10.5411
R4025 b2b.n5 b2b.n3 9.44853
R4026 b2b.n5 b2b.n4 9.35588
R4027 b2b.n2 b2b.t2 9.19699
R4028 b2b.n1 b2b.n0 8.57376
R4029 b2b.n6 b2b 3.36483
R4030 b2b b2b.n6 2.25319
R4031 b2b.n2 b2b.n1 0.226273
R4032 b2b.n6 b2b.n5 0.00180435
R4033 B1 B1.t0 48.6474
R4034 B1.n0 B1.t1 19.0247
R4035 B1.n0 B1.t2 17.3935
R4036 B1.n1 B1.n0 4.12942
R4037 B1.n1 B1 2.25699
R4038 B1 B1.n1 0.0067069
R4039 b1b b1b.n5 37.091
R4040 b1b.n3 b1b.t2 26.9594
R4041 b1b b1b.t3 19.4226
R4042 b1b.n5 b1b.n2 9.59479
R4043 b1b.n7 b1b.n0 9.49418
R4044 b1b.n6 b1b.n1 9.39109
R4045 b1b.n4 b1b.n3 7.55447
R4046 b1b.n3 b1b.n2 4.95899
R4047 b1b.n6 b1b 3.31968
R4048 b1b.t4 b1b.n2 2.79883
R4049 b1b b1b.n7 2.25319
R4050 b1b.n5 b1b.n4 1.68928
R4051 b1b.n4 b1b.t4 0.678302
R4052 b1b.n7 b1b.n6 0.00963044
R4053 ITAIL.n12 ITAIL.n7 333.663
R4054 ITAIL.n8 ITAIL.t22 116.817
R4055 ITAIL.n10 ITAIL.n9 103.823
R4056 ITAIL.n3 ITAIL.t17 97.648
R4057 ITAIL.n7 ITAIL.n6 90.8936
R4058 ITAIL.n12 ITAIL.n11 88.6306
R4059 ITAIL.n5 ITAIL.n4 84.9459
R4060 ITAIL.n9 ITAIL.n8 48.8699
R4061 ITAIL.n11 ITAIL.n10 47.0449
R4062 ITAIL.n4 ITAIL.n3 38.4914
R4063 ITAIL.n6 ITAIL.n5 38.4914
R4064 ITAIL ITAIL.t15 27.414
R4065 ITAIL.t22 ITAIL.t18 23.7985
R4066 ITAIL.t9 ITAIL.t5 23.7985
R4067 ITAIL.t16 ITAIL.t8 23.7985
R4068 ITAIL.t7 ITAIL.t3 23.7985
R4069 ITAIL.t23 ITAIL.t19 23.7985
R4070 ITAIL.t17 ITAIL.t11 23.7985
R4071 ITAIL.t4 ITAIL.t24 23.7985
R4072 ITAIL.t20 ITAIL.t14 23.7985
R4073 ITAIL.t2 ITAIL.t21 23.7985
R4074 ITAIL.t10 ITAIL.t6 23.7985
R4075 ITAIL.n8 ITAIL.t9 12.9945
R4076 ITAIL.n9 ITAIL.t16 12.9945
R4077 ITAIL.n10 ITAIL.t7 12.9945
R4078 ITAIL.n11 ITAIL.t23 12.9945
R4079 ITAIL.t15 ITAIL.n12 12.7755
R4080 ITAIL.n3 ITAIL.t4 12.7025
R4081 ITAIL.n4 ITAIL.t20 12.7025
R4082 ITAIL.n5 ITAIL.t2 12.7025
R4083 ITAIL.n6 ITAIL.t10 12.7025
R4084 ITAIL.n7 ITAIL.t12 10.8045
R4085 ITAIL.n0 ITAIL.t0 8.6875
R4086 ITAIL.n0 ITAIL.t13 7.3735
R4087 ITAIL.n1 ITAIL.t1 6.06997
R4088 ITAIL ITAIL.n2 4.95899
R4089 ITAIL.n2 ITAIL.n1 4.07166
R4090 ITAIL.n2 ITAIL.n0 2.47975
R4091 ITAIL.n1 ITAIL 0.00782558
R4092 SDn_1.n38 SDn_1.n35 4.73161
R4093 SDn_1.n34 SDn_1.n33 3.08659
R4094 SDn_1.n41 SDn_1.n40 3.04854
R4095 SDn_1.n25 SDn_1.n10 3.04726
R4096 SDn_1.n17 SDn_1.n16 3.04688
R4097 SDn_1.n52 SDn_1.n6 3.04375
R4098 SDn_1.n43 SDn_1.n8 3.04171
R4099 SDn_1.n19 SDn_1.n12 3.03541
R4100 SDn_1.n40 SDn_1.n39 2.9021
R4101 SDn_1.n4 SDn_1.t1 2.7305
R4102 SDn_1.n4 SDn_1.n3 2.7305
R4103 SDn_1.n49 SDn_1.t17 2.7305
R4104 SDn_1.n49 SDn_1.n48 2.7305
R4105 SDn_1.n45 SDn_1.t7 2.7305
R4106 SDn_1.n45 SDn_1.n44 2.7305
R4107 SDn_1.n37 SDn_1.t29 2.7305
R4108 SDn_1.n37 SDn_1.n36 2.7305
R4109 SDn_1.n31 SDn_1.t0 2.7305
R4110 SDn_1.n31 SDn_1.n30 2.7305
R4111 SDn_1.n27 SDn_1.t28 2.7305
R4112 SDn_1.n27 SDn_1.n26 2.7305
R4113 SDn_1.n21 SDn_1.t3 2.7305
R4114 SDn_1.n21 SDn_1.n20 2.7305
R4115 SDn_1.n14 SDn_1.t16 2.7305
R4116 SDn_1.n14 SDn_1.n13 2.7305
R4117 SDn_1.n16 SDn_1.t6 2.7305
R4118 SDn_1.n16 SDn_1.n15 2.7305
R4119 SDn_1.n12 SDn_1.t27 2.7305
R4120 SDn_1.n12 SDn_1.n11 2.7305
R4121 SDn_1.n10 SDn_1.t11 2.7305
R4122 SDn_1.n10 SDn_1.n9 2.7305
R4123 SDn_1.n33 SDn_1.t31 2.7305
R4124 SDn_1.n33 SDn_1.n32 2.7305
R4125 SDn_1.n8 SDn_1.t26 2.7305
R4126 SDn_1.n8 SDn_1.n7 2.7305
R4127 SDn_1.n6 SDn_1.t9 2.7305
R4128 SDn_1.n6 SDn_1.n5 2.7305
R4129 SDn_1.n1 SDn_1.t18 2.7305
R4130 SDn_1.n1 SDn_1.n0 2.7305
R4131 SDn_1.n17 SDn_1.n14 2.56247
R4132 SDn_1.n38 SDn_1.n37 2.56221
R4133 SDn_1.n34 SDn_1.n31 2.562
R4134 SDn_1.n54 SDn_1.n4 2.55991
R4135 SDn_1.n40 SDn_1.t8 2.40706
R4136 SDn_1.n51 SDn_1.n50 1.49447
R4137 SDn_1.n23 SDn_1.n22 1.49447
R4138 SDn_1.n29 SDn_1.n28 1.49423
R4139 SDn_1.n47 SDn_1.n46 1.49423
R4140 SDn_1.n50 SDn_1.n49 1.43787
R4141 SDn_1.n28 SDn_1.n27 1.43765
R4142 SDn_1.n46 SDn_1.n45 1.43732
R4143 SDn_1.n22 SDn_1.n21 1.437
R4144 SDn_1.n2 SDn_1.n1 1.4264
R4145 SDn_1.n55 SDn_1.n2 1.14083
R4146 SDn_1.n51 SDn_1.n47 0.58072
R4147 SDn_1.n18 SDn_1.n17 0.575838
R4148 SDn_1.n24 SDn_1.n23 0.574178
R4149 SDn_1.n54 SDn_1.n53 0.566624
R4150 SDn_1.n35 SDn_1.n29 0.554675
R4151 SDn_1.n42 SDn_1.n41 0.513212
R4152 SDn_1.n55 SDn_1.n54 0.482617
R4153 SDn_1.n2 SDn_1 0.157421
R4154 SDn_1.n19 SDn_1.n18 0.0271667
R4155 SDn_1.n53 SDn_1.n52 0.0249444
R4156 SDn_1.n47 SDn_1.n43 0.0212506
R4157 SDn_1.n25 SDn_1.n24 0.0205
R4158 SDn_1.n29 SDn_1.n25 0.0201395
R4159 SDn_1.n43 SDn_1.n42 0.0193889
R4160 SDn_1.n52 SDn_1.n51 0.0153623
R4161 SDn_1.n23 SDn_1.n19 0.0134755
R4162 SDn_1.n35 SDn_1.n34 0.0132059
R4163 SDn_1 SDn_1.n55 0.00682738
R4164 SDn_1.n41 SDn_1.n38 0.00579412
R4165 b3.t8 b3.t2 102.266
R4166 b3.n0 b3.t4 49.5502
R4167 b3 b3.t5 34.9792
R4168 b3.t9 b3.t7 28.703
R4169 b3.t10 b3.t6 26.4242
R4170 b3.t2 b3.t9 22.0465
R4171 b3.t6 b3.t8 22.0465
R4172 b3.t7 b3.t3 17.6665
R4173 b3.t5 b3.t10 17.6665
R4174 b3.n1 b3.t1 9.49371
R4175 b3.n1 b3.t0 9.3756
R4176 b3 b3.n1 3.6563
R4177 b3.n0 b3 3.36711
R4178 b3 b3.n0 2.25981
R4179 OUT3.n14 OUT3.n10 19.1949
R4180 OUT3.n13 OUT3.n11 6.45579
R4181 OUT3.n15 OUT3.n14 6.06989
R4182 OUT3.n13 OUT3.n12 5.8805
R4183 OUT3.n16 OUT3.t6 5.8805
R4184 OUT3.n15 OUT3.t7 5.8805
R4185 OUT3.n4 OUT3.n1 3.63586
R4186 OUT3.n9 OUT3.n6 3.63586
R4187 OUT3.n4 OUT3.n3 3.1505
R4188 OUT3.n9 OUT3.n8 3.1505
R4189 OUT3.n1 OUT3.t1 2.7305
R4190 OUT3.n1 OUT3.n0 2.7305
R4191 OUT3.n3 OUT3.t4 2.7305
R4192 OUT3.n3 OUT3.n2 2.7305
R4193 OUT3.n6 OUT3.t11 2.7305
R4194 OUT3.n6 OUT3.n5 2.7305
R4195 OUT3.n8 OUT3.t0 2.7305
R4196 OUT3.n8 OUT3.n7 2.7305
R4197 OUT3.n14 OUT3 2.39886
R4198 OUT3.n10 OUT3.n4 0.804767
R4199 OUT3.n16 OUT3.n15 0.564731
R4200 OUT3 OUT3.n13 0.199912
R4201 OUT3.n10 OUT3.n9 0.190191
R4202 OUT3 OUT3.n16 0.0558846
R4203 b4.n3 b4.n0 485.19
R4204 b4.n7 b4.n6 79.2611
R4205 b4.n1 b4.t10 65.6295
R4206 b4.n5 b4.t8 64.5576
R4207 b4.t13 b4.t15 62.9752
R4208 b4.t7 b4.n7 62.5658
R4209 b4.n10 b4.t12 51.8002
R4210 b4.t16 b4.t13 41.6538
R4211 b4.t17 b4.t9 32.3937
R4212 b4.t8 b4.t2 20.3675
R4213 b4.t5 b4.t16 20.3675
R4214 b4.n6 b4.n5 20.0889
R4215 b4.t18 b4.t6 18.2505
R4216 b4 b4.n9 17.3009
R4217 b4.t10 b4.t3 16.0605
R4218 b4.n8 b4.t14 15.7355
R4219 b4.n6 b4.t5 13.8705
R4220 b4.n4 b4.t4 13.2149
R4221 b4.n8 b4.t7 10.1176
R4222 b4.n5 b4.t17 10.0015
R4223 b4.n11 b4.t0 9.49371
R4224 b4.n11 b4.t1 9.3756
R4225 b4.n2 b4.n1 8.61736
R4226 b4.n4 b4.n3 8.26992
R4227 b4.n9 b4.n8 5.77524
R4228 b4.n7 b4.t18 5.4025
R4229 b4.n3 b4.n2 4.86717
R4230 b4.n9 b4.n4 4.43773
R4231 b4 b4.n11 3.6563
R4232 b4.n1 b4.n0 2.03842
R4233 b4.t11 b4.n0 1.91942
R4234 b4.n2 b4.t11 0.122167
R4235 b4 b4.n10 0.00981034
R4236 b4.n10 b4 0.00256897
R4237 SD2_1 SD2_1.n20 9.24575
R4238 SD2_1.n19 SD2_1.n18 3.45039
R4239 SD2_1.n14 SD2_1.n13 3.44985
R4240 SD2_1.n9 SD2_1.n8 3.44969
R4241 SD2_1.n4 SD2_1.n3 3.44925
R4242 SD2_1.n14 SD2_1.n11 3.4367
R4243 SD2_1.n19 SD2_1.n16 3.43615
R4244 SD2_1.n4 SD2_1.n1 3.43133
R4245 SD2_1 SD2_1.n6 3.3305
R4246 SD2_1.n20 SD2_1.n19 2.87896
R4247 SD2_1 SD2_1.n4 2.8298
R4248 SD2_1.n6 SD2_1.t10 2.7305
R4249 SD2_1.n6 SD2_1.n5 2.7305
R4250 SD2_1.n11 SD2_1.t1 2.7305
R4251 SD2_1.n11 SD2_1.n10 2.7305
R4252 SD2_1.n13 SD2_1.t3 2.7305
R4253 SD2_1.n13 SD2_1.n12 2.7305
R4254 SD2_1.n16 SD2_1.t8 2.7305
R4255 SD2_1.n16 SD2_1.n15 2.7305
R4256 SD2_1.n18 SD2_1.t9 2.7305
R4257 SD2_1.n18 SD2_1.n17 2.7305
R4258 SD2_1.n1 SD2_1.t4 2.7305
R4259 SD2_1.n1 SD2_1.n0 2.7305
R4260 SD2_1.n3 SD2_1.t5 2.7305
R4261 SD2_1.n3 SD2_1.n2 2.7305
R4262 SD2_1.n8 SD2_1.t11 2.7305
R4263 SD2_1.n8 SD2_1.n7 2.7305
R4264 SD2_1.n20 SD2_1.n14 2.25147
R4265 SD2_1 SD2_1.n9 2.2505
R4266 SD2_1.n9 SD2_1 0.100126
R4267 G1_2.n6 G1_2.n2 147.578
R4268 G1_2.n17 G1_2.n16 142.844
R4269 G1_2.n15 G1_2.n14 101.016
R4270 G1_2.n1 G1_2.n0 101.016
R4271 G1_2.n5 G1_2.n4 101.016
R4272 G1_2.n13 G1_2.n12 101.016
R4273 G1_2.n14 G1_2.t29 33.5864
R4274 G1_2.n0 G1_2.t31 33.5864
R4275 G1_2.n16 G1_2.n15 20.5194
R4276 G1_2.n2 G1_2.n1 20.5194
R4277 G1_2.n6 G1_2.n5 20.5194
R4278 G1_2.n4 G1_2.n3 20.5194
R4279 G1_2.n12 G1_2.n11 20.5194
R4280 G1_2.n17 G1_2.n13 20.5194
R4281 G1_2.n14 G1_2.t34 13.0675
R4282 G1_2.n15 G1_2.t30 13.0675
R4283 G1_2.n16 G1_2.t32 13.0675
R4284 G1_2.n0 G1_2.t26 13.0675
R4285 G1_2.n1 G1_2.t24 13.0675
R4286 G1_2.n2 G1_2.t28 13.0675
R4287 G1_2.n5 G1_2.t8 13.0675
R4288 G1_2.n4 G1_2.t0 13.0675
R4289 G1_2.n3 G1_2.t6 13.0675
R4290 G1_2.n11 G1_2.t4 13.0675
R4291 G1_2.n12 G1_2.t10 13.0675
R4292 G1_2.n13 G1_2.t14 13.0675
R4293 G1_2.n9 G1_2.t12 8.3225
R4294 G1_2.n47 G1_2.t2 8.1765
R4295 G1_2.n43 G1_2.n41 6.51833
R4296 G1_2.n37 G1_2.t23 6.51833
R4297 G1_2.n45 G1_2.t17 5.8805
R4298 G1_2.n44 G1_2.t18 5.8805
R4299 G1_2.n43 G1_2.n42 5.8805
R4300 G1_2.n39 G1_2.n35 5.8805
R4301 G1_2.n38 G1_2.n36 5.8805
R4302 G1_2.n37 G1_2.t16 5.8805
R4303 G1_2.n46 G1_2.n45 5.81863
R4304 G1_2.n40 G1_2.n39 5.52662
R4305 G1_2.n49 G1_2.n48 4.5005
R4306 G1_2.n46 G1_2.n40 4.28996
R4307 G1_2.n8 G1_2.n7 3.53359
R4308 G1_2.n33 G1_2.n18 3.50535
R4309 G1_2.n20 G1_2.t13 3.03383
R4310 G1_2.n20 G1_2.n19 3.03383
R4311 G1_2.n22 G1_2.t11 3.03383
R4312 G1_2.n22 G1_2.n21 3.03383
R4313 G1_2.n24 G1_2.t7 3.03383
R4314 G1_2.n24 G1_2.n23 3.03383
R4315 G1_2.n26 G1_2.t9 3.03383
R4316 G1_2.n26 G1_2.n25 3.03383
R4317 G1_2.n34 G1_2.n10 2.88425
R4318 G1_2.n30 G1_2.n22 2.8392
R4319 G1_2.n29 G1_2.n24 2.8392
R4320 G1_2.n31 G1_2.n20 2.80007
R4321 G1_2.n28 G1_2.n26 2.80007
R4322 G1_2.n40 G1_2.n34 2.5439
R4323 G1_2.n10 G1_2.n9 2.1905
R4324 G1_2.n44 G1_2.n43 2.07441
R4325 G1_2.n48 G1_2.n47 2.0445
R4326 G1_2.n38 G1_2.n37 2.0118
R4327 G1_2.n49 G1_2.n46 1.80063
R4328 G1_2.n30 G1_2.n29 1.59702
R4329 G1_2.n31 G1_2.n30 1.58339
R4330 G1_2.n29 G1_2.n28 1.58339
R4331 G1_2.n7 G1_2.n6 1.15481
R4332 G1_2.n18 G1_2.n17 1.06529
R4333 G1_2.n45 G1_2.n44 0.638326
R4334 G1_2.n39 G1_2.n38 0.638326
R4335 G1_2.n32 G1_2.n31 0.0932273
R4336 G1_2 G1_2.n27 0.0876818
R4337 G1_2.n33 G1_2.n32 0.0305
R4338 G1_2.n27 G1_2.n8 0.0265
R4339 G1_2.n28 G1_2 0.0100455
R4340 G1_2 G1_2.n8 0.0085
R4341 G1_2.n34 G1_2.n33 0.0055
R4342 G1_2 G1_2.n49 0.0025
R4343 SD1_1.n15 SD1_1.n14 7.78572
R4344 SD1_1.n9 SD1_1.n8 3.20235
R4345 SD1_1.n17 SD1_1.n16 3.17681
R4346 SD1_1.n1 SD1_1.t8 3.03383
R4347 SD1_1.n1 SD1_1.n0 3.03383
R4348 SD1_1.n22 SD1_1.t7 3.03383
R4349 SD1_1.n22 SD1_1.n21 3.03383
R4350 SD1_1.n19 SD1_1.t15 3.03383
R4351 SD1_1.n19 SD1_1.n18 3.03383
R4352 SD1_1.n13 SD1_1.t1 3.03383
R4353 SD1_1.n13 SD1_1.n12 3.03383
R4354 SD1_1.n5 SD1_1.t13 3.03383
R4355 SD1_1.n5 SD1_1.n4 3.03383
R4356 SD1_1.n7 SD1_1.t0 3.03383
R4357 SD1_1.n7 SD1_1.n6 3.03383
R4358 SD1_1.n20 SD1_1.n17 2.97146
R4359 SD1_1.n10 SD1_1.n9 2.94829
R4360 SD1_1.n10 SD1_1.n7 2.75112
R4361 SD1_1.n17 SD1_1.t2 2.69498
R4362 SD1_1.n9 SD1_1.t10 2.66057
R4363 SD1_1.n14 SD1_1.n13 2.38615
R4364 SD1_1.n23 SD1_1.n22 2.37424
R4365 SD1_1.n20 SD1_1.n19 2.37412
R4366 SD1_1.n11 SD1_1.n5 2.37207
R4367 SD1_1.n2 SD1_1.n1 1.63787
R4368 SD1_1.n15 SD1_1.n3 1.12886
R4369 SD1_1.n23 SD1_1.n20 0.626727
R4370 SD1_1.n11 SD1_1.n10 0.613463
R4371 SD1_1.n14 SD1_1.n11 0.609042
R4372 SD1_1.n24 SD1_1.n23 0.584266
R4373 SD1_1.n2 SD1_1 0.0568907
R4374 SD1_1 SD1_1.n24 0.0265
R4375 SD1_1.n3 SD1_1.n2 0.0213805
R4376 SD1_1 SD1_1.n15 0.00686644
R4377 SD2_4.n10 SD2_4.n4 5.11704
R4378 SD2_4.n4 SD2_4.n1 3.44424
R4379 SD2_4.n9 SD2_4.n8 3.37323
R4380 SD2_4.n4 SD2_4.n3 3.33687
R4381 SD2_4 SD2_4.n6 3.31692
R4382 SD2_4.n6 SD2_4.t2 2.7305
R4383 SD2_4.n6 SD2_4.n5 2.7305
R4384 SD2_4.n1 SD2_4.t6 2.7305
R4385 SD2_4.n1 SD2_4.n0 2.7305
R4386 SD2_4.n3 SD2_4.t7 2.7305
R4387 SD2_4.n3 SD2_4.n2 2.7305
R4388 SD2_4.n8 SD2_4.t3 2.7305
R4389 SD2_4.n8 SD2_4.n7 2.7305
R4390 SD2_4.n10 SD2_4.n9 2.2505
R4391 SD2_4.n9 SD2_4 0.116226
R4392 SD2_4 SD2_4.n10 0.00261765
R4393 G1_1.n27 G1_1.t24 113.573
R4394 G1_1.n17 G1_1.t28 113.573
R4395 G1_1.n29 G1_1.n28 101.016
R4396 G1_1.n19 G1_1.n18 101.016
R4397 G1_1.n21 G1_1.n20 101.016
R4398 G1_1.n23 G1_1.n22 101.016
R4399 G1_1.n25 G1_1.n24 101.016
R4400 G1_1.n30 G1_1.n26 101.016
R4401 G1_1.n20 G1_1.n19 67.0816
R4402 G1_1.n30 G1_1.n29 62.3464
R4403 G1_1.n28 G1_1.n27 20.5194
R4404 G1_1.n18 G1_1.n17 20.5194
R4405 G1_1.n22 G1_1.n21 20.5194
R4406 G1_1.n24 G1_1.n23 20.5194
R4407 G1_1.n26 G1_1.n25 20.5194
R4408 G1_1.n27 G1_1.t30 12.5565
R4409 G1_1.n28 G1_1.t35 12.5565
R4410 G1_1.n29 G1_1.t25 12.5565
R4411 G1_1.n17 G1_1.t29 12.5565
R4412 G1_1.n18 G1_1.t34 12.5565
R4413 G1_1.n19 G1_1.t32 12.5565
R4414 G1_1.n21 G1_1.t22 12.5565
R4415 G1_1.n22 G1_1.t12 12.5565
R4416 G1_1.n23 G1_1.t16 12.5565
R4417 G1_1.n24 G1_1.t8 12.5565
R4418 G1_1.n25 G1_1.t10 12.5565
R4419 G1_1.n26 G1_1.t18 12.5565
R4420 G1_1.n0 G1_1.t20 10.2935
R4421 G1_1.n31 G1_1.t14 10.2935
R4422 G1_1.n32 G1_1.n31 4.12693
R4423 G1_1 G1_1.n0 4.0015
R4424 G1_1.n2 G1_1.t5 3.03383
R4425 G1_1.n2 G1_1.n1 3.03383
R4426 G1_1.n16 G1_1.t15 3.03383
R4427 G1_1.n16 G1_1.n15 3.03383
R4428 G1_1.n4 G1_1.t23 3.03383
R4429 G1_1.n4 G1_1.n3 3.03383
R4430 G1_1.n6 G1_1.t0 3.03383
R4431 G1_1.n6 G1_1.n5 3.03383
R4432 G1_1.n8 G1_1.t17 3.03383
R4433 G1_1.n8 G1_1.n7 3.03383
R4434 G1_1.n10 G1_1.t6 3.03383
R4435 G1_1.n10 G1_1.n9 3.03383
R4436 G1_1.n12 G1_1.t11 3.03383
R4437 G1_1.n12 G1_1.n11 3.03383
R4438 G1_1.n14 G1_1.t2 3.03383
R4439 G1_1.n14 G1_1.n13 3.03383
R4440 G1_1.n38 G1_1.n4 2.82159
R4441 G1_1.n37 G1_1.n6 2.82159
R4442 G1_1.n36 G1_1.n8 2.82159
R4443 G1_1.n35 G1_1.n10 2.82159
R4444 G1_1.n34 G1_1.n12 2.82159
R4445 G1_1.n33 G1_1.n14 2.82159
R4446 G1_1.n39 G1_1.n2 2.78833
R4447 G1_1.n32 G1_1.n16 2.78833
R4448 G1_1.n20 G1_1.n0 2.2635
R4449 G1_1.n31 G1_1.n30 2.2635
R4450 G1_1.n34 G1_1.n33 0.798761
R4451 G1_1.n35 G1_1.n34 0.798761
R4452 G1_1.n36 G1_1.n35 0.798761
R4453 G1_1.n37 G1_1.n36 0.798761
R4454 G1_1.n38 G1_1.n37 0.798761
R4455 G1_1.n33 G1_1.n32 0.786618
R4456 G1_1 G1_1.n38 0.626587
R4457 G1_1.n39 G1_1 0.160531
R4458 G1_1 G1_1.n39 0.0949286
R4459 B3 B3.t2 48.6474
R4460 B3.n0 B3.t1 19.0247
R4461 B3.n0 B3.t0 17.3935
R4462 B3.n1 B3.n0 4.12942
R4463 B3.n1 B3 2.25699
R4464 B3 B3.n1 0.0067069
R4465 b3b.n6 b3b.t3 36.6929
R4466 b3b.t5 b3b.t8 22.0465
R4467 b3b.t7 b3b.t10 22.0465
R4468 b3b.n6 b3b.t2 18.6988
R4469 b3b.t9 b3b.t4 17.6665
R4470 b3b.t3 b3b.t6 17.6665
R4471 b3b.n4 b3b.t5 12.209
R4472 b3b.n5 b3b.t7 12.0202
R4473 b3b.t6 b3b.n5 11.1473
R4474 b3b.n4 b3b.t9 10.8684
R4475 b3b.n1 b3b.n0 9.49288
R4476 b3b.n3 b3b.n2 9.40022
R4477 b3b.n5 b3b.n4 8.7605
R4478 b3b b3b.n3 2.25319
R4479 b3b b3b.n6 0.681545
R4480 b3b.n1 b3b 0.177597
R4481 b3b.n3 b3b.n1 0.00180435
R4482 OUT1 OUT1.n1 24.2283
R4483 OUT1 OUT1.t2 5.96093
R4484 OUT1.n1 OUT1.t1 2.7305
R4485 OUT1.n1 OUT1.n0 2.7305
R4486 SD2_3.n3 SD2_3.n2 6.50095
R4487 SD2_3.n2 SD2_3.n0 6.4673
R4488 SD2_3 SD2_3.t2 6.08127
R4489 SD2_3.n3 SD2_3.t0 5.8805
R4490 SD2_3.n2 SD2_3.n1 5.8805
R4491 SD2_3 SD2_3.n3 0.291269
R4492 b1.n4 b1.t3 50.6785
R4493 b1.n1 b1.n0 41.4888
R4494 b1 b1.n3 33.4868
R4495 b1.n1 b1.t2 17.9739
R4496 b1.n5 b1.t0 9.49371
R4497 b1.n5 b1.t1 9.3756
R4498 b1.n3 b1.n0 6.4245
R4499 b1.t4 b1.n0 4.50217
R4500 b1 b1.n5 3.6563
R4501 b1.n3 b1.n2 2.47632
R4502 b1.n2 b1.n1 1.66454
R4503 b1.n4 b1 0.858629
R4504 b1.n2 b1.t4 0.254192
R4505 b1 b1.n4 0.0800215
R4506 B5 B5.t0 48.6474
R4507 B5.n0 B5.t1 19.0247
R4508 B5.n0 B5.t2 17.3935
R4509 B5.n1 B5.n0 4.12942
R4510 B5.n1 B5 2.25699
R4511 B5 B5.n1 0.0067069
R4512 B4 B4.t1 48.6474
R4513 B4.n0 B4.t0 19.0247
R4514 B4.n0 B4.t2 17.3935
R4515 B4.n1 B4.n0 4.12942
R4516 B4.n1 B4 2.25699
R4517 B4 B4.n1 0.0067069
R4518 B2 B2.t1 48.6474
R4519 B2.n0 B2.t0 19.0247
R4520 B2.n0 B2.t2 17.3935
R4521 B2.n1 B2.n0 4.12942
R4522 B2.n1 B2 2.25699
R4523 B2 B2.n1 0.0067069
R4524 SD2_2 SD2_2.n1 3.20344
R4525 SD2_2.n1 SD2_2.t0 2.7305
R4526 SD2_2.n1 SD2_2.n0 2.7305
C0 OUT2 ITAIL 0.148f
C1 b1b b5b 0.00116f
C2 b1 b5 7.09e-19
C3 b3 b6 0.638f
C4 b2 SD2_5 0.0557f
C5 OUT1 SD2_2 0.037f
C6 OUT3 G2 0.131f
C7 b2b SD2_1 0.0528f
C8 G1_1 G1_2 2.47f
C9 b4 OUT4 0.286f
C10 Balance_Inverter_5.Inverter_0.OUT OUT- 2.36e-19
C11 OUT5 B2 1.94e-19
C12 b4b m1_n558_n5402# 0.0175f
C13 b4b B5 0.0998f
C14 SD2_1 SD2_5 0.0861f
C15 G2 SD2_4 0.162f
C16 b4b B3 0.0144f
C17 b4 b5 0.473f
C18 OUT4 b6b 0.0011f
C19 ITAIL SD2_3 0.0655f
C20 OUT5 OUT+ 1.49f
C21 Balance_Inverter_4.Inverter_0.OUT B6 8.24e-19
C22 B5 Balance_Inverter_5.Inverter_0.OUT 0.00124f
C23 B4 Balance_Inverter_4.Inverter_0.OUT 0.00122f
C24 Balance_Inverter_0.Inverter_0.OUT B5 8.09e-19
C25 B3 Balance_Inverter_0.Inverter_0.OUT 0.00299f
C26 Balance_Inverter_1.Inverter_0.OUT B4 5.37e-20
C27 B1 Balance_Inverter_2.Inverter_0.OUT 0.00299f
C28 B2 Balance_Inverter_1.Inverter_0.OUT 0.00207f
C29 Balance_Inverter_2.Inverter_0.OUT B3 5.45e-20
C30 Balance_Inverter_3.Inverter_0.OUT B2 5.37e-20
C31 b6 b5b 0.0019f
C32 b6b b5 0.0482f
C33 Balance_Inverter_4.Inverter_0.OUT OUT+ 3.2e-20
C34 VDD b1 0.945f
C35 SDn_2 b2 0.0229f
C36 OUT6 SDn_1 0.0272f
C37 VDD b4 1.22f
C38 b1b b3b 1.73e-19
C39 b1 OUT1 0.14f
C40 SD3_1 OUT5 0.0124f
C41 IT b2b 0.267f
C42 b1 OUT- 0.294f
C43 b1 SD1_1 0.136f
C44 VDD b6b 0.316f
C45 b1b OUT4 0.0382f
C46 SDn_1 OUT2 0.00105f
C47 b2 OUT3 0.0568f
C48 b3b G1_1 0.00976f
C49 OUT5 b4b 0.00918f
C50 OUT1 b4 5.52e-19
C51 b4 OUT- 1.52f
C52 OUT5 Balance_Inverter_5.Inverter_0.OUT 7.09e-20
C53 b2 SD2_4 1.72e-19
C54 b1 B1 0.0809f
C55 b3 b5b 0.0547f
C56 OUT2 G2 0.0518f
C57 OUT3 SD2_1 1.08f
C58 b2b SD2_5 0.0626f
C59 b1b b5 5.92e-19
C60 G1_1 OUT4 2.54e-19
C61 b6b OUT- 2.62f
C62 b4b Balance_Inverter_4.Inverter_0.OUT 0.0129f
C63 b4b Balance_Inverter_1.Inverter_0.OUT 1.07e-19
C64 b4 m1_n558_n5402# 1.3e-19
C65 b4 B5 0.0558f
C66 b4 B3 0.138f
C67 G2 SD2_3 0.0979f
C68 G1_2 b5b 2.13e-19
C69 SD2_1 SD2_4 0.00298f
C70 ITAIL SD2_2 0.00992f
C71 Balance_Inverter_4.Inverter_0.OUT Balance_Inverter_5.Inverter_0.OUT 3.48e-19
C72 Balance_Inverter_0.Inverter_0.OUT Balance_Inverter_4.Inverter_0.OUT 3.46e-19
C73 Balance_Inverter_1.Inverter_0.OUT Balance_Inverter_0.Inverter_0.OUT 0.00437f
C74 Balance_Inverter_2.Inverter_0.OUT Balance_Inverter_1.Inverter_0.OUT 0.00442f
C75 Balance_Inverter_3.Inverter_0.OUT Balance_Inverter_2.Inverter_0.OUT 0.00437f
C76 b6 b5 0.0112f
C77 G2 OUT+ 0.00111f
C78 IT SDn_2 4.09f
C79 VDD b1b 0.595f
C80 b1 OUT5 0.0759f
C81 b1b OUT1 0.0235f
C82 VDD G1_1 8.11f
C83 b3 b3b 0.982f
C84 IT OUT3 4.23e-20
C85 SDn_2 b2b 0.105f
C86 SD3_1 SDn_1 0.297f
C87 OUT6 b2 0.323f
C88 b1b OUT- 0.131f
C89 OUT1 G1_1 5.82e-19
C90 b1 ITAIL 0.0202f
C91 b3b G1_2 0.0816f
C92 OUT5 b4 4.5e-19
C93 b2b OUT3 0.00957f
C94 b2 OUT2 0.0421f
C95 b1b SD1_1 0.223f
C96 VDD b6 0.567f
C97 G1_1 OUT- 4.07e-20
C98 b1 Balance_Inverter_3.Inverter_0.OUT 0.221f
C99 G1_2 OUT4 2.09f
C100 OUT3 SD2_5 0.182f
C101 b2b SD2_4 0.00446f
C102 G1_1 SD1_1 0.279f
C103 b3b b5b 0.0105f
C104 b2 SD2_3 1.08e-19
C105 b1b B1 0.257f
C106 OUT2 SD2_1 0.00162f
C107 b3 b5 0.0495f
C108 b6 OUT- 3.42f
C109 b4 Balance_Inverter_4.Inverter_0.OUT 0.00897f
C110 b4 Balance_Inverter_1.Inverter_0.OUT 0.00255f
C111 b2 B2 0.0869f
C112 G2 SD2_2 0.0436f
C113 SD2_1 SD2_3 8.03e-19
C114 SD2_5 SD2_4 0.31f
C115 b2 OUT+ 0.78f
C116 b5b b5 1.92f
C117 SD2_1 OUT+ 0.00903f
C118 IT OUT6 0.783f
C119 VDD b3 0.75f
C120 b1b OUT5 0.204f
C121 IT OUT2 0.093f
C122 OUT6 b2b 0.323f
C123 SD3_1 b2 0.167f
C124 b1 SDn_1 0.129f
C125 VDD G1_2 3.63f
C126 b3 OUT- 0.749f
C127 b2 b4b 0.0522f
C128 b1 G2 0.0266f
C129 b2b OUT2 0.0772f
C130 OUT1 G1_2 0.0347f
C131 b3b OUT4 0.0472f
C132 OUT5 G1_1 0.0268f
C133 VDD b5b 0.38f
C134 b1b ITAIL 0.0195f
C135 G1_2 OUT- 8.68e-23
C136 b1b Balance_Inverter_3.Inverter_0.OUT 0.0252f
C137 b3 m1_n558_n5402# 0.00587f
C138 b3 B5 0.0272f
C139 b2 Balance_Inverter_2.Inverter_0.OUT 0.224f
C140 b3 B3 0.0937f
C141 OUT3 SD2_4 0.373f
C142 b2b SD2_3 0.00175f
C143 b3b b5 4.52e-19
C144 G1_2 SD1_1 0.646f
C145 OUT2 SD2_5 0.363f
C146 b5b OUT- 1.25f
C147 b2b B2 0.288f
C148 IT OUT+ 4.29e-19
C149 SD2_5 SD2_3 0.0442f
C150 b2b OUT+ 0.469f
C151 b5b m1_n558_n5402# 2.68e-20
C152 b5b B5 0.169f
C153 b5b B3 0.0015f
C154 b5b B1 0.0019f
C155 VDD b3b 0.926f
C156 IT SD3_1 1.01f
C157 SDn_2 OUT6 1.22f
C158 b1b SDn_1 0.132f
C159 SDn_2 OUT2 0.0016f
C160 SD3_1 b2b 0.576f
C161 OUT6 OUT3 0.00428f
C162 VDD OUT4 0.00148f
C163 b1 b2 0.0351f
C164 b3 OUT5 3.51e-19
C165 b3b OUT- 0.211f
C166 b2 b4 0.0116f
C167 b3b SD1_1 0.0957f
C168 b2b b4b 0.033f
C169 OUT1 OUT4 1.78f
C170 VDD b5 0.754f
C171 SDn_1 G1_1 0.00119f
C172 b1 SD2_1 0.0946f
C173 OUT3 OUT2 0.265f
C174 b1b G2 0.0135f
C175 OUT5 G1_2 0.0345f
C176 OUT4 OUT- 0.841f
C177 b3 Balance_Inverter_4.Inverter_0.OUT 0.00594f
C178 b3 Balance_Inverter_1.Inverter_0.OUT 0.228f
C179 b3b m1_n558_n5402# 0.00129f
C180 b2b Balance_Inverter_2.Inverter_0.OUT 0.0239f
C181 b3b B3 0.531f
C182 OUT4 SD1_1 0.0013f
C183 OUT5 b5b 1.6f
C184 b3b B1 1.29e-19
C185 OUT2 SD2_4 0.281f
C186 OUT3 SD2_3 0.401f
C187 G1_2 ITAIL 0.404f
C188 b5 OUT- 2.15f
C189 SD2_4 SD2_3 0.461f
C190 SD2_5 SD2_2 0.0175f
C191 ITAIL b5b 9.45e-19
C192 b5b Balance_Inverter_4.Inverter_0.OUT 0.00753f
C193 OUT3 OUT+ 1.43f
C194 b5 m1_n558_n5402# 1.27e-20
C195 b5 B5 0.0874f
C196 b5 B3 1.07e-19
C197 VDD OUT1 0.0376f
C198 IT b1 0.2f
C199 SDn_2 SD3_1 0.716f
C200 VDD OUT- 0.00913f
C201 b1 b2b 0.0403f
C202 VDD SD1_1 1.94f
C203 b3b OUT5 0.0251f
C204 b1b b2 0.0845f
C205 OUT1 OUT- 0.257f
C206 VDD m1_n558_n5402# 0.0568f
C207 VDD B5 0.282f
C208 SDn_1 G1_2 5.13e-19
C209 OUT3 b4b 0.0594f
C210 OUT5 OUT4 0.0458f
C211 OUT1 SD1_1 5.9e-19
C212 VDD B1 0.411f
C213 b2 G1_1 0.0077f
C214 b3b ITAIL 0.0199f
C215 b1b SD2_1 0.0398f
C216 b2b b4 9.46e-20
C217 VDD B3 0.38f
C218 b1 SD2_5 0.0356f
C219 OUT6 B6 2.15e-19
C220 b3b Balance_Inverter_1.Inverter_0.OUT 0.0887f
C221 OUT4 ITAIL 0.346f
C222 OUT2 SD2_3 0.16f
C223 OUT5 b5 1.49f
C224 G1_2 G2 0.192f
C225 B5 OUT- 2.65e-20
C226 B1 OUT- 7.92e-19
C227 B3 OUT- 1.23e-19
C228 OUT6 OUT+ 5.15f
C229 G2 b5b 0.00908f
C230 b5 Balance_Inverter_4.Inverter_0.OUT 0.219f
C231 OUT2 OUT+ 0.798f
C232 B6 OUT+ 1.53e-19
C233 B2 OUT+ 0.0069f
C234 VDD OUT5 0.163f
C235 SDn_2 b1 0.0286f
C236 OUT6 SD3_1 3.97f
C237 IT b1b 0.316f
C238 b1b b2b 1.03f
C239 OUT1 OUT5 0.551f
C240 VDD ITAIL 0.0217f
C241 b3 b2 0.0682f
C242 OUT6 b4b 0.19f
C243 b3b SDn_1 0.11f
C244 IT G1_1 0.374f
C245 b1 OUT3 0.0392f
C246 OUT5 OUT- 2.33f
C247 VDD Balance_Inverter_4.Inverter_0.OUT 0.14f
C248 VDD Balance_Inverter_1.Inverter_0.OUT 0.153f
C249 VDD Balance_Inverter_3.Inverter_0.OUT 0.154f
C250 OUT1 ITAIL 0.168f
C251 OUT3 b4 0.1f
C252 b3b G2 0.0142f
C253 b2 G1_2 0.045f
C254 OUT2 b4b 0.107f
C255 b1b SD2_5 0.0386f
C256 b1 SD2_4 0.0372f
C257 OUT5 SD1_1 0.0778f
C258 b2b G1_1 0.0281f
C259 ITAIL OUT- 1.71e-20
C260 Balance_Inverter_4.Inverter_0.OUT OUT- 0.00136f
C261 Balance_Inverter_3.Inverter_0.OUT OUT- 4.26e-21
C262 OUT4 G2 0.246f
C263 OUT3 b6b 3.6e-21
C264 OUT2 SD2_2 0.00234f
C265 G1_2 SD2_1 0.906f
C266 OUT5 B1 3.74e-21
C267 b4b B6 9.34e-20
C268 b4b B4 0.2f
C269 SD2_1 b5b 0.00393f
C270 B6 Balance_Inverter_5.Inverter_0.OUT 0.158f
C271 B5 Balance_Inverter_4.Inverter_0.OUT 0.159f
C272 B4 Balance_Inverter_0.Inverter_0.OUT 0.158f
C273 B3 Balance_Inverter_1.Inverter_0.OUT 0.139f
C274 B2 Balance_Inverter_2.Inverter_0.OUT 0.158f
C275 B1 Balance_Inverter_3.Inverter_0.OUT 0.158f
C276 b4b OUT+ 1.18f
C277 Balance_Inverter_5.Inverter_0.OUT OUT+ 3.93e-21
C278 Balance_Inverter_2.Inverter_0.OUT OUT+ 3.09e-21
C279 OUT6 b1 0.0167f
C280 SDn_2 b1b 0.0933f
C281 VDD SDn_1 0.00435f
C282 b3 b2b 0.127f
C283 b3b b2 3.71f
C284 SDn_2 G1_1 0.0117f
C285 OUT1 SDn_1 0.00609f
C286 b1 OUT2 1.07f
C287 VDD G2 0.0272f
C288 b1b OUT3 0.0345f
C289 OUT6 b4 0.282f
C290 IT G1_2 2.95f
C291 b2b G1_2 0.0676f
C292 b3b SD2_1 0.0885f
C293 OUT1 G2 0.0299f
C294 b1b SD2_4 0.0374f
C295 b1 SD2_3 0.0369f
C296 OUT3 G1_1 5.54e-20
C297 OUT6 b6b 1.29f
C298 b2 OUT4 0.0745f
C299 OUT2 b4 0.00657f
C300 OUT5 ITAIL 0.0132f
C301 SDn_1 SD1_1 0.0889f
C302 G2 OUT- 2.86e-20
C303 b4b Balance_Inverter_5.Inverter_0.OUT 1.27e-19
C304 b4b Balance_Inverter_0.Inverter_0.OUT 0.00424f
C305 b2b b5b 4.11e-19
C306 b2 b5 0.00157f
C307 G1_2 SD2_5 0.00259f
C308 OUT4 SD2_1 0.0612f
C309 b4 B6 0.049f
C310 b1 OUT+ 0.119f
C311 b4 B4 0.0688f
C312 SD2_1 b5 0.0012f
C313 G2 B1 4.42e-19
C314 b6b B6 0.209f
C315 b4 OUT+ 1.31f
C316 b6b OUT+ 2.58f
C317 OUT6 b1b 0.199f
C318 VDD b2 0.825f
C319 IT b3b 0.294f
C320 SD3_1 b1 0.00977f
C321 OUT5 SDn_1 2.14f
C322 IT OUT4 0.00118f
C323 b1b OUT2 0.0214f
C324 VDD SD2_1 0.127f
C325 b3 OUT3 0.139f
C326 b3b b2b 0.132f
C327 b1 b4b 5.58e-20
C328 OUT1 b2 0.0236f
C329 b2 OUT- 0.551f
C330 OUT2 G1_1 0.0171f
C331 b4b b4 4.11f
C332 b1b SD2_3 0.0345f
C333 b3b SD2_5 0.00858f
C334 b2b OUT4 0.056f
C335 b1 SD2_2 0.00207f
C336 OUT6 b6 1.42f
C337 b2 SD1_1 0.0595f
C338 OUT3 G1_2 0.0268f
C339 OUT1 SD2_1 0.023f
C340 OUT5 G2 0.0135f
C341 SD2_1 OUT- 7.37e-19
C342 b4 Balance_Inverter_5.Inverter_0.OUT 0.00832f
C343 b4 Balance_Inverter_0.Inverter_0.OUT 0.219f
C344 b2b b5 0.00104f
C345 G1_2 SD2_4 2.28e-19
C346 b2 B1 0.166f
C347 OUT3 b5b 0.00986f
C348 ITAIL G2 1.17f
C349 OUT4 SD2_5 1.05f
C350 b4b b6b 0.235f
C351 G2 Balance_Inverter_3.Inverter_0.OUT 4.19e-20
C352 b1b OUT+ 0.255f
C353 b6b Balance_Inverter_5.Inverter_0.OUT 0.00445f
C354 SD2_1 B1 0.00396f
C355 b6 B6 0.0742f
C356 G1_1 OUT+ 8.45e-19
C357 b6 OUT+ 2.79f
C358 VDD IT 1.49f
C359 OUT6 b3 0.847f
C360 SDn_2 b3b 0.0371f
C361 IT OUT1 0.00193f
C362 SD3_1 b1b 0.272f
C363 VDD b2b 0.696f
C364 IT OUT- 2.35e-20
C365 b3 OUT2 4.2e-20
C366 b3b OUT3 0.111f
C367 VDD SD2_5 1.38e-19
C368 b1b b4b 0.00121f
C369 OUT1 b2b 0.00657f
C370 OUT5 b2 0.0264f
C371 IT SD1_1 2.13f
C372 b1 b4 1.1e-19
C373 b2b OUT- 0.406f
C374 OUT2 G1_2 0.273f
C375 b4b G1_1 5.38e-19
C376 b2 ITAIL 0.00991f
C377 OUT5 SD2_1 0.0727f
C378 OUT3 OUT4 1.33f
C379 b2b SD1_1 0.0397f
C380 b3b SD2_4 9.52e-20
C381 OUT1 SD2_5 0.548f
C382 b3 B6 0.0254f
C383 b3 B2 0.164f
C384 b2 Balance_Inverter_3.Inverter_0.OUT 0.00628f
C385 b3 B4 0.0697f
C386 G1_2 SD2_3 8.28e-20
C387 b4 b6b 0.286f
C388 b2b B3 0.00249f
C389 ITAIL SD2_1 0.159f
C390 OUT4 SD2_4 0.00348f
C391 OUT3 b5 0.00482f
C392 b4b b6 0.213f
C393 b2b B1 0.011f
C394 SD2_1 Balance_Inverter_3.Inverter_0.OUT 5.32e-19
C395 b3 OUT+ 0.534f
C396 b6 Balance_Inverter_5.Inverter_0.OUT 0.22f
C397 b5b B6 0.0464f
C398 b5b B2 6.52e-21
C399 G1_2 OUT+ 3.98e-19
C400 b5b OUT+ 1.39f
C401 VDD SDn_2 0.0496f
C402 b1 b1b 2.47f
C403 VDD OUT3 4.91e-20
C404 OUT6 b3b 0.219f
C405 SDn_2 OUT1 4.33e-19
C406 IT OUT5 1.02f
C407 OUT1 OUT3 0.223f
C408 OUT5 b2b 0.164f
C409 b1 G1_1 0.0912f
C410 b3 b4b 0.202f
C411 SDn_2 SD1_1 0.0268f
C412 SDn_1 b2 0.0994f
C413 IT ITAIL 0.0238f
C414 OUT3 OUT- 0.7f
C415 b3 Balance_Inverter_5.Inverter_0.OUT 0.00522f
C416 b3 Balance_Inverter_0.Inverter_0.OUT 0.0159f
C417 b3 Balance_Inverter_2.Inverter_0.OUT 0.00384f
C418 OUT2 OUT4 1.26f
C419 OUT3 SD1_1 1.31e-19
C420 b2 G2 0.021f
C421 b3b SD2_3 6.42e-20
C422 OUT1 SD2_4 0.00368f
C423 b2b ITAIL 0.0175f
C424 b2b Balance_Inverter_1.Inverter_0.OUT 0.00182f
C425 b3b B4 0.00452f
C426 b2b Balance_Inverter_3.Inverter_0.OUT 0.00219f
C427 b3b B2 0.0246f
C428 OUT4 SD2_3 0.00229f
C429 OUT3 B1 3.71e-20
C430 ITAIL SD2_5 0.265f
C431 G2 SD2_1 0.214f
C432 b4b b5b 0.11f
C433 b4 b6 0.783f
C434 b3b OUT+ 0.244f
C435 b5b Balance_Inverter_5.Inverter_0.OUT 0.0132f
C436 b6b b6 3.11f
C437 b5 B6 0.0134f
C438 b5 B2 4.82e-19
C439 OUT4 OUT+ 0.815f
C440 b5 OUT+ 1.33f
C441 b1 b3 6.43e-19
C442 SD3_1 b3b 0.162f
C443 OUT6 OUT1 0.0634f
C444 SDn_2 OUT5 0.926f
C445 VDD OUT2 0.0816f
C446 IT SDn_1 1.02f
C447 OUT6 OUT- 6.47f
C448 SDn_1 b2b 0.111f
C449 b1 G1_2 0.25f
C450 b3 b4 0.305f
C451 OUT1 OUT2 0.352f
C452 OUT5 OUT3 0.0882f
C453 b1b G1_1 0.0784f
C454 IT G2 0.00126f
C455 b3b b4b 0.0222f
C456 OUT2 OUT- 0.471f
C457 VDD B6 0.284f
C458 VDD B4 0.29f
C459 VDD B2 0.375f
C460 b3b Balance_Inverter_0.Inverter_0.OUT 0.00272f
C461 b3b Balance_Inverter_2.Inverter_0.OUT 0.00135f
C462 b2b G2 0.0204f
C463 OUT2 SD1_1 0.0494f
C464 b2 SD2_1 0.0523f
C465 b1 b5b 9.41e-19
C466 b3 b6b 0.0399f
C467 OUT1 SD2_3 0.00462f
C468 OUT3 ITAIL 0.128f
C469 b4b OUT4 0.224f
C470 VDD OUT+ 0.00687f
C471 B6 OUT- 0.00132f
C472 B2 OUT- 1.01e-20
C473 ITAIL SD2_4 0.124f
C474 b4b b5 0.154f
C475 G2 SD2_5 0.248f
C476 b4 b5b 0.0441f
C477 OUT1 OUT+ 0.172f
C478 OUT- OUT+ 15.8f
C479 b5 Balance_Inverter_5.Inverter_0.OUT 0.00537f
C480 b6b b5b 0.00479f
C481 B5 B6 0.0375f
C482 B3 B4 0.0325f
C483 B4 B5 0.0331f
C484 B2 B3 0.0158f
C485 SD1_1 OUT+ 5.17e-20
C486 B1 B2 0.0325f
C487 B1 OUT+ 0.00379f
C488 VDD b4b 0.428f
C489 OUT6 OUT5 0.0131f
C490 IT b2 0.161f
C491 SDn_2 SDn_1 0.586f
C492 b1 b3b 1.42e-19
C493 b1b b3 3.65e-19
C494 VDD Balance_Inverter_5.Inverter_0.OUT 0.14f
C495 VDD Balance_Inverter_2.Inverter_0.OUT 0.154f
C496 VDD Balance_Inverter_0.Inverter_0.OUT 0.14f
C497 b3b b4 0.00815f
C498 OUT5 OUT2 0.0703f
C499 b1 OUT4 0.103f
C500 IT SD2_1 0.00647f
C501 b2 b2b 4.83f
C502 OUT1 b4b 4.44e-19
C503 b1b G1_2 0.0867f
C504 b4b OUT- 1.34f
C505 OUT+ VSS 18.7f
C506 OUT- VSS 20.4f
C507 m1_n558_n5402# VSS 0.0572f $ **FLOATING
C508 Balance_Inverter_5.Inverter_0.OUT VSS 0.552f
C509 B6 VSS 1.37f
C510 Balance_Inverter_4.Inverter_0.OUT VSS 0.553f
C511 B5 VSS 1.34f
C512 Balance_Inverter_0.Inverter_0.OUT VSS 0.564f
C513 B4 VSS 1.49f
C514 Balance_Inverter_1.Inverter_0.OUT VSS 0.55f
C515 B3 VSS 1.2f
C516 Balance_Inverter_2.Inverter_0.OUT VSS 0.549f
C517 B2 VSS 1.22f
C518 Balance_Inverter_3.Inverter_0.OUT VSS 0.551f
C519 B1 VSS 1.12f
C520 b5 VSS 6.56f
C521 b5b VSS 7.46f
C522 b6 VSS 13.7f
C523 b6b VSS 14.4f
C524 SD2_2 VSS 0.0529f
C525 SD2_3 VSS 1.08f
C526 SD2_4 VSS 0.57f
C527 SD2_5 VSS 1.01f
C528 SD2_1 VSS 2.64f
C529 G2 VSS 7.64f
C530 ITAIL VSS 7.81f
C531 SD1_1 VSS 0.746f
C532 OUT4 VSS 3.18f
C533 G1_2 VSS 5.35f
C534 G1_1 VSS 1.57f
C535 b4 VSS 6.37f
C536 b4b VSS 8.37f
C537 OUT2 VSS 1.58f
C538 OUT3 VSS 1.84f
C539 b2b VSS 5.9f
C540 b2 VSS 3.51f
C541 SDn_1 VSS 2.33f
C542 OUT5 VSS 4.71f
C543 OUT1 VSS 1.3f
C544 b3b VSS 5.91f
C545 b3 VSS 8.03f
C546 b1b VSS 4f
C547 b1 VSS 4.5f
C548 SD3_1 VSS 3.94f
C549 OUT6 VSS 11.3f
C550 SDn_2 VSS 16.2f
C551 IT VSS 29.6f
C552 VDD VSS 35.9f
C553 b1.n0 VSS 0.00429f
C554 b1.t2 VSS 0.0263f
C555 b1.n1 VSS 0.0245f
C556 b1.t4 VSS 0.0025f
C557 b1.n2 VSS 0.00755f
C558 b1.n3 VSS 0.38f
C559 b1.t3 VSS 0.0221f
C560 b1.n4 VSS 0.112f
C561 b1.t0 VSS 0.00677f
C562 b1.t1 VSS 0.00536f
C563 b1.n5 VSS 0.116f
C564 b3b.n0 VSS 0.00469f
C565 b3b.n1 VSS 0.0325f
C566 b3b.n2 VSS 0.00523f
C567 b3b.n3 VSS 0.0274f
C568 b3b.t2 VSS 0.00861f
C569 b3b.t4 VSS 0.0172f
C570 b3b.t9 VSS 0.0312f
C571 b3b.t8 VSS 0.0269f
C572 b3b.t5 VSS 0.0376f
C573 b3b.n4 VSS 0.0308f
C574 b3b.t10 VSS 0.0269f
C575 b3b.t7 VSS 0.0375f
C576 b3b.n5 VSS 0.031f
C577 b3b.t6 VSS 0.0311f
C578 b3b.t3 VSS 1.01f
C579 b3b.n6 VSS 2.26f
C580 G1_1.t20 VSS 0.109f
C581 G1_1.n0 VSS 0.108f
C582 G1_1.t5 VSS 0.0392f
C583 G1_1.n1 VSS 0.0392f
C584 G1_1.n2 VSS 0.0826f
C585 G1_1.t23 VSS 0.0392f
C586 G1_1.n3 VSS 0.0392f
C587 G1_1.n4 VSS 0.0837f
C588 G1_1.t0 VSS 0.0392f
C589 G1_1.n5 VSS 0.0392f
C590 G1_1.n6 VSS 0.0837f
C591 G1_1.t17 VSS 0.0392f
C592 G1_1.n7 VSS 0.0392f
C593 G1_1.n8 VSS 0.0837f
C594 G1_1.t6 VSS 0.0392f
C595 G1_1.n9 VSS 0.0392f
C596 G1_1.n10 VSS 0.0837f
C597 G1_1.t11 VSS 0.0392f
C598 G1_1.n11 VSS 0.0392f
C599 G1_1.n12 VSS 0.0837f
C600 G1_1.t2 VSS 0.0392f
C601 G1_1.n13 VSS 0.0392f
C602 G1_1.n14 VSS 0.0837f
C603 G1_1.t15 VSS 0.0392f
C604 G1_1.n15 VSS 0.0392f
C605 G1_1.n16 VSS 0.0826f
C606 G1_1.t28 VSS 0.352f
C607 G1_1.t29 VSS 0.128f
C608 G1_1.n17 VSS 0.303f
C609 G1_1.t34 VSS 0.128f
C610 G1_1.n18 VSS 0.275f
C611 G1_1.t32 VSS 0.128f
C612 G1_1.n19 VSS 0.33f
C613 G1_1.n20 VSS 0.242f
C614 G1_1.t22 VSS 0.128f
C615 G1_1.n21 VSS 0.275f
C616 G1_1.t12 VSS 0.128f
C617 G1_1.n22 VSS 0.275f
C618 G1_1.t16 VSS 0.128f
C619 G1_1.n23 VSS 0.275f
C620 G1_1.t8 VSS 0.128f
C621 G1_1.n24 VSS 0.275f
C622 G1_1.t10 VSS 0.128f
C623 G1_1.n25 VSS 0.275f
C624 G1_1.t18 VSS 0.128f
C625 G1_1.n26 VSS 0.275f
C626 G1_1.t24 VSS 0.353f
C627 G1_1.t30 VSS 0.128f
C628 G1_1.n27 VSS 0.303f
C629 G1_1.t35 VSS 0.128f
C630 G1_1.n28 VSS 0.275f
C631 G1_1.t25 VSS 0.128f
C632 G1_1.n29 VSS 0.325f
C633 G1_1.n30 VSS 0.236f
C634 G1_1.t14 VSS 0.109f
C635 G1_1.n31 VSS 0.111f
C636 G1_1.n32 VSS 0.353f
C637 G1_1.n33 VSS 0.328f
C638 G1_1.n34 VSS 0.33f
C639 G1_1.n35 VSS 0.33f
C640 G1_1.n36 VSS 0.33f
C641 G1_1.n37 VSS 0.33f
C642 G1_1.n38 VSS 0.304f
C643 G1_1.n39 VSS 0.148f
C644 SD1_1.t8 VSS 0.0112f
C645 SD1_1.n0 VSS 0.0112f
C646 SD1_1.n1 VSS 0.0224f
C647 SD1_1.n2 VSS 0.00497f
C648 SD1_1.n3 VSS 0.022f
C649 SD1_1.t13 VSS 0.0112f
C650 SD1_1.n4 VSS 0.0112f
C651 SD1_1.n5 VSS 0.0297f
C652 SD1_1.t0 VSS 0.0112f
C653 SD1_1.n6 VSS 0.0112f
C654 SD1_1.n7 VSS 0.0308f
C655 SD1_1.n8 VSS 0.0121f
C656 SD1_1.t10 VSS 0.0103f
C657 SD1_1.n9 VSS 0.0453f
C658 SD1_1.n10 VSS 0.143f
C659 SD1_1.n11 VSS 0.094f
C660 SD1_1.t1 VSS 0.0112f
C661 SD1_1.n12 VSS 0.0112f
C662 SD1_1.n13 VSS 0.0337f
C663 SD1_1.n14 VSS 0.559f
C664 SD1_1.n15 VSS 0.506f
C665 SD1_1.t2 VSS 0.0104f
C666 SD1_1.n16 VSS 0.012f
C667 SD1_1.n17 VSS 0.0519f
C668 SD1_1.t15 VSS 0.0112f
C669 SD1_1.n18 VSS 0.0112f
C670 SD1_1.n19 VSS 0.0347f
C671 SD1_1.n20 VSS 0.153f
C672 SD1_1.t7 VSS 0.0112f
C673 SD1_1.n21 VSS 0.0112f
C674 SD1_1.n22 VSS 0.0347f
C675 SD1_1.n23 VSS 0.0988f
C676 SD1_1.n24 VSS 0.0438f
C677 G1_2.t31 VSS 0.143f
C678 G1_2.t26 VSS 0.0827f
C679 G1_2.n0 VSS 0.212f
C680 G1_2.t24 VSS 0.0827f
C681 G1_2.n1 VSS 0.174f
C682 G1_2.t28 VSS 0.0827f
C683 G1_2.n2 VSS 0.208f
C684 G1_2.t8 VSS 0.0827f
C685 G1_2.t0 VSS 0.0827f
C686 G1_2.t6 VSS 0.0827f
C687 G1_2.n3 VSS 0.174f
C688 G1_2.n4 VSS 0.174f
C689 G1_2.n5 VSS 0.174f
C690 G1_2.n6 VSS 0.149f
C691 G1_2.n7 VSS 0.00736f
C692 G1_2.n8 VSS 0.012f
C693 G1_2.t12 VSS 0.0572f
C694 G1_2.n9 VSS 0.0564f
C695 G1_2.n10 VSS 0.0239f
C696 G1_2.t4 VSS 0.0827f
C697 G1_2.n11 VSS 0.174f
C698 G1_2.t10 VSS 0.0827f
C699 G1_2.n12 VSS 0.174f
C700 G1_2.t14 VSS 0.0827f
C701 G1_2.n13 VSS 0.174f
C702 G1_2.t29 VSS 0.143f
C703 G1_2.t34 VSS 0.0827f
C704 G1_2.n14 VSS 0.212f
C705 G1_2.t30 VSS 0.0827f
C706 G1_2.n15 VSS 0.174f
C707 G1_2.t32 VSS 0.0827f
C708 G1_2.n16 VSS 0.204f
C709 G1_2.n17 VSS 0.146f
C710 G1_2.n18 VSS 0.00327f
C711 G1_2.t13 VSS 0.0244f
C712 G1_2.n19 VSS 0.0244f
C713 G1_2.n20 VSS 0.0517f
C714 G1_2.t11 VSS 0.0244f
C715 G1_2.n21 VSS 0.0244f
C716 G1_2.n22 VSS 0.0525f
C717 G1_2.t7 VSS 0.0244f
C718 G1_2.n23 VSS 0.0244f
C719 G1_2.n24 VSS 0.0525f
C720 G1_2.t9 VSS 0.0244f
C721 G1_2.n25 VSS 0.0244f
C722 G1_2.n26 VSS 0.0517f
C723 G1_2.n27 VSS 0.0312f
C724 G1_2.n28 VSS 0.209f
C725 G1_2.n29 VSS 0.354f
C726 G1_2.n30 VSS 0.354f
C727 G1_2.n31 VSS 0.225f
C728 G1_2.n32 VSS 0.0327f
C729 G1_2.n33 VSS 0.0123f
C730 G1_2.n34 VSS 0.0413f
C731 G1_2.n35 VSS 0.0557f
C732 G1_2.n36 VSS 0.0557f
C733 G1_2.t23 VSS 0.0661f
C734 G1_2.t16 VSS 0.0557f
C735 G1_2.n37 VSS 0.376f
C736 G1_2.n38 VSS 0.279f
C737 G1_2.n39 VSS 0.434f
C738 G1_2.n40 VSS 1.28f
C739 G1_2.t17 VSS 0.0557f
C740 G1_2.t18 VSS 0.0557f
C741 G1_2.n41 VSS 0.0661f
C742 G1_2.n42 VSS 0.0557f
C743 G1_2.n43 VSS 0.381f
C744 G1_2.n44 VSS 0.285f
C745 G1_2.n45 VSS 0.463f
C746 G1_2.n46 VSS 1.32f
C747 G1_2.t2 VSS 0.0564f
C748 G1_2.n47 VSS 0.0548f
C749 G1_2.n48 VSS 0.0228f
C750 G1_2.n49 VSS 0.0395f
C751 b4.n0 VSS 0.00816f
C752 b4.t11 VSS 0.00241f
C753 b4.t3 VSS 0.0268f
C754 b4.t10 VSS 0.098f
C755 b4.n1 VSS 0.0545f
C756 b4.n2 VSS 0.0155f
C757 b4.n3 VSS 0.0276f
C758 b4.t4 VSS 0.0233f
C759 b4.n4 VSS 0.11f
C760 b4.t14 VSS 0.0271f
C761 b4.t6 VSS 0.031f
C762 b4.t18 VSS 0.0453f
C763 b4.t2 VSS 0.0435f
C764 b4.t8 VSS 0.114f
C765 b4.t9 VSS 0.0607f
C766 b4.t17 VSS 0.0754f
C767 b4.n5 VSS 0.0752f
C768 b4.t15 VSS 0.0612f
C769 b4.t13 VSS 0.125f
C770 b4.t16 VSS 0.107f
C771 b4.t5 VSS 0.0655f
C772 b4.n6 VSS 0.102f
C773 b4.n7 VSS 0.124f
C774 b4.t7 VSS 0.0762f
C775 b4.n8 VSS 0.0623f
C776 b4.n9 VSS 1.11f
C777 b4.t12 VSS 0.0309f
C778 b4.n10 VSS 0.0606f
C779 b4.t0 VSS 0.00966f
C780 b4.t1 VSS 0.00765f
C781 b4.n11 VSS 0.165f
C782 SDn_1.t18 VSS 0.00812f
C783 SDn_1.n0 VSS 0.00812f
C784 SDn_1.n1 VSS 0.0163f
C785 SDn_1.n2 VSS 0.0188f
C786 SDn_1.t1 VSS 0.00812f
C787 SDn_1.n3 VSS 0.00812f
C788 SDn_1.n4 VSS 0.0223f
C789 SDn_1.t9 VSS 0.00812f
C790 SDn_1.n5 VSS 0.00812f
C791 SDn_1.n6 VSS 0.0284f
C792 SDn_1.t26 VSS 0.00812f
C793 SDn_1.n7 VSS 0.00812f
C794 SDn_1.n8 VSS 0.0296f
C795 SDn_1.t11 VSS 0.00812f
C796 SDn_1.n9 VSS 0.00812f
C797 SDn_1.n10 VSS 0.0297f
C798 SDn_1.t27 VSS 0.00812f
C799 SDn_1.n11 VSS 0.00812f
C800 SDn_1.n12 VSS 0.0296f
C801 SDn_1.t16 VSS 0.00812f
C802 SDn_1.n13 VSS 0.00812f
C803 SDn_1.n14 VSS 0.0223f
C804 SDn_1.t6 VSS 0.00812f
C805 SDn_1.n15 VSS 0.00812f
C806 SDn_1.n16 VSS 0.0298f
C807 SDn_1.n17 VSS 0.109f
C808 SDn_1.n18 VSS 0.0306f
C809 SDn_1.n19 VSS 0.0658f
C810 SDn_1.t3 VSS 0.00812f
C811 SDn_1.n20 VSS 0.00812f
C812 SDn_1.n21 VSS 0.0163f
C813 SDn_1.n22 VSS 0.0137f
C814 SDn_1.n23 VSS 0.0292f
C815 SDn_1.n24 VSS 0.03f
C816 SDn_1.n25 VSS 0.066f
C817 SDn_1.t28 VSS 0.00812f
C818 SDn_1.n26 VSS 0.00812f
C819 SDn_1.n27 VSS 0.0163f
C820 SDn_1.n28 VSS 0.0137f
C821 SDn_1.n29 VSS 0.0293f
C822 SDn_1.t0 VSS 0.00812f
C823 SDn_1.n30 VSS 0.00812f
C824 SDn_1.n31 VSS 0.0223f
C825 SDn_1.t31 VSS 0.00812f
C826 SDn_1.n32 VSS 0.00812f
C827 SDn_1.n33 VSS 0.0305f
C828 SDn_1.n34 VSS 0.078f
C829 SDn_1.n35 VSS 0.249f
C830 SDn_1.t29 VSS 0.00812f
C831 SDn_1.n36 VSS 0.00812f
C832 SDn_1.n37 VSS 0.0223f
C833 SDn_1.n38 VSS 0.232f
C834 SDn_1.n39 VSS 0.00883f
C835 SDn_1.t8 VSS 0.00751f
C836 SDn_1.n40 VSS 0.0324f
C837 SDn_1.n41 VSS 0.0943f
C838 SDn_1.n42 VSS 0.0294f
C839 SDn_1.n43 VSS 0.0654f
C840 SDn_1.t7 VSS 0.00812f
C841 SDn_1.n44 VSS 0.00812f
C842 SDn_1.n45 VSS 0.0163f
C843 SDn_1.n46 VSS 0.0137f
C844 SDn_1.n47 VSS 0.0324f
C845 SDn_1.t17 VSS 0.00812f
C846 SDn_1.n48 VSS 0.00812f
C847 SDn_1.n49 VSS 0.0163f
C848 SDn_1.n50 VSS 0.0137f
C849 SDn_1.n51 VSS 0.0317f
C850 SDn_1.n52 VSS 0.065f
C851 SDn_1.n53 VSS 0.0308f
C852 SDn_1.n54 VSS 0.0689f
C853 SDn_1.n55 VSS 0.0319f
C854 b1b.n0 VSS 0.0068f
C855 b1b.n1 VSS 0.00755f
C856 b1b.n2 VSS 0.00752f
C857 b1b.t2 VSS 0.0405f
C858 b1b.n3 VSS 0.0317f
C859 b1b.t4 VSS 0.00448f
C860 b1b.n4 VSS 0.00585f
C861 b1b.n5 VSS 0.5f
C862 b1b.n6 VSS 0.0854f
C863 b1b.n7 VSS 0.0389f
C864 b1b.t3 VSS 0.0157f
C865 b2b.t4 VSS 0.0158f
C866 b2b.t6 VSS 0.0295f
C867 b2b.n0 VSS 0.0536f
C868 b2b.t3 VSS 0.0156f
C869 b2b.n1 VSS 0.0317f
C870 b2b.t2 VSS 0.0292f
C871 b2b.n2 VSS 1.55f
C872 b2b.n3 VSS 0.00819f
C873 b2b.n4 VSS 0.00916f
C874 b2b.n5 VSS 0.0899f
C875 b2b.n6 VSS 0.0691f
C876 b2b.t5 VSS 0.0194f
C877 OUT4.n0 VSS 0.0146f
C878 OUT4.n1 VSS 0.0124f
C879 OUT4.n2 VSS 0.0464f
C880 OUT4.n3 VSS 0.0124f
C881 OUT4.n4 VSS 0.0124f
C882 OUT4.t10 VSS 0.0147f
C883 OUT4.t6 VSS 0.0124f
C884 OUT4.n5 VSS 0.0986f
C885 OUT4.n6 VSS 0.0701f
C886 OUT4.n7 VSS 0.0384f
C887 OUT4.t21 VSS 0.00542f
C888 OUT4.n8 VSS 0.00542f
C889 OUT4.n9 VSS 0.0108f
C890 OUT4.t13 VSS 0.00542f
C891 OUT4.n10 VSS 0.00542f
C892 OUT4.n11 VSS 0.0108f
C893 OUT4.t0 VSS 0.00542f
C894 OUT4.n12 VSS 0.00542f
C895 OUT4.n13 VSS 0.0108f
C896 OUT4.t18 VSS 0.00542f
C897 OUT4.n14 VSS 0.00542f
C898 OUT4.n15 VSS 0.0147f
C899 OUT4.n16 VSS 0.0475f
C900 OUT4.n17 VSS 0.0297f
C901 OUT4.n18 VSS 0.0433f
C902 OUT4.t12 VSS 0.00542f
C903 OUT4.n19 VSS 0.00542f
C904 OUT4.n20 VSS 0.0108f
C905 OUT4.t17 VSS 0.00542f
C906 OUT4.n21 VSS 0.00542f
C907 OUT4.n22 VSS 0.0108f
C908 OUT4.t14 VSS 0.00542f
C909 OUT4.n23 VSS 0.00542f
C910 OUT4.n24 VSS 0.0108f
C911 OUT4.t1 VSS 0.00542f
C912 OUT4.n25 VSS 0.00542f
C913 OUT4.n26 VSS 0.0145f
C914 OUT4.n27 VSS 0.0454f
C915 OUT4.n28 VSS 0.0289f
C916 OUT4.n29 VSS 0.0203f
C917 OUT4.n30 VSS 0.366f
C918 OUT4.n31 VSS 0.678f
C919 OUT4.t3 VSS 0.0124f
C920 OUT4.n32 VSS 0.188f
C921 OUT4.t11 VSS 0.0124f
C922 OUT4.n33 VSS 0.0613f
C923 b4b.t5 VSS 0.0217f
C924 b4b.t15 VSS 0.0237f
C925 b4b.n0 VSS 0.0437f
C926 b4b.t17 VSS 0.0237f
C927 b4b.n1 VSS 0.0437f
C928 b4b.t13 VSS 0.0821f
C929 b4b.t10 VSS 0.161f
C930 b4b.t2 VSS 0.0386f
C931 b4b.n2 VSS 0.151f
C932 b4b.t8 VSS 0.112f
C933 b4b.n3 VSS 0.16f
C934 b4b.t3 VSS 0.0986f
C935 b4b.t7 VSS 0.0817f
C936 b4b.t18 VSS 0.0132f
C937 b4b.n4 VSS 0.0407f
C938 b4b.t14 VSS 0.0124f
C939 b4b.n5 VSS 0.0367f
C940 b4b.t4 VSS 0.0738f
C941 b4b.t12 VSS 0.184f
C942 b4b.t6 VSS 0.0298f
C943 b4b.n6 VSS 0.222f
C944 b4b.t16 VSS 0.0976f
C945 b4b.t11 VSS 0.0369f
C946 b4b.n7 VSS 0.0917f
C947 b4b.n8 VSS 0.74f
C948 b4b.n9 VSS 1.15f
C949 b4b.n11 VSS 0.00307f
C950 b4b.n12 VSS 0.0118f
C951 b4b.n13 VSS 0.00771f
C952 b4b.n14 VSS 0.00293f
C953 b4b.n15 VSS 0.0103f
C954 b4b.n16 VSS 0.00858f
C955 b4b.n17 VSS 0.0672f
C956 b4b.n18 VSS 0.0436f
C957 b4b.n19 VSS 0.00866f
C958 b4b.t9 VSS 0.0178f
C959 b5.t11 VSS 0.0191f
C960 b5.t5 VSS 0.0149f
C961 b5.t8 VSS 0.0149f
C962 b5.t22 VSS 0.0151f
C963 b5.n0 VSS 0.0315f
C964 b5.t17 VSS 0.0149f
C965 b5.n1 VSS 0.0317f
C966 b5.t7 VSS 0.0953f
C967 b5.t19 VSS 0.0951f
C968 b5.n2 VSS 0.0315f
C969 b5.t15 VSS 0.0149f
C970 b5.n3 VSS 0.0317f
C971 b5.t4 VSS 0.0607f
C972 b5.t25 VSS 0.0185f
C973 b5.t14 VSS 0.0142f
C974 b5.t9 VSS 0.0282f
C975 b5.t6 VSS 0.0571f
C976 b5.t18 VSS 0.0282f
C977 b5.t16 VSS 0.0546f
C978 b5.t13 VSS 0.0198f
C979 b5.n4 VSS 0.05f
C980 b5.t21 VSS 0.0198f
C981 b5.n5 VSS 0.0346f
C982 b5.n6 VSS 0.034f
C983 b5.t26 VSS 0.0308f
C984 b5.t3 VSS 0.0139f
C985 b5.n7 VSS 0.0329f
C986 b5.t24 VSS 0.0139f
C987 b5.n8 VSS 0.0329f
C988 b5.t20 VSS 0.0308f
C989 b5.n9 VSS 0.034f
C990 b5.t12 VSS 0.0198f
C991 b5.n10 VSS 0.0369f
C992 b5.t2 VSS 0.00794f
C993 b5.n11 VSS 0.133f
C994 b5.n12 VSS 0.0778f
C995 b5.t23 VSS 0.0195f
C996 b5.n13 VSS 0.0673f
C997 b5.t10 VSS 0.0195f
C998 b5.n14 VSS 0.0654f
C999 b5.n15 VSS 0.0344f
C1000 b5.n16 VSS 0.365f
C1001 b5.t0 VSS 0.00597f
C1002 b5.t1 VSS 0.00472f
C1003 b5.n17 VSS 0.0923f
C1004 b5.n18 VSS 0.168f
C1005 OUT5.t18 VSS 0.00776f
C1006 OUT5.n0 VSS 0.00776f
C1007 OUT5.n1 VSS 0.0155f
C1008 OUT5.t38 VSS 0.00776f
C1009 OUT5.n2 VSS 0.00776f
C1010 OUT5.n3 VSS 0.0155f
C1011 OUT5.t39 VSS 0.00776f
C1012 OUT5.n4 VSS 0.00776f
C1013 OUT5.n5 VSS 0.0155f
C1014 OUT5.t26 VSS 0.00776f
C1015 OUT5.n6 VSS 0.00776f
C1016 OUT5.n7 VSS 0.0212f
C1017 OUT5.n8 VSS 0.0641f
C1018 OUT5.n9 VSS 0.0398f
C1019 OUT5.n10 VSS 0.0603f
C1020 OUT5.t37 VSS 0.00776f
C1021 OUT5.n11 VSS 0.00776f
C1022 OUT5.n12 VSS 0.0155f
C1023 OUT5.t22 VSS 0.00776f
C1024 OUT5.n13 VSS 0.00776f
C1025 OUT5.n14 VSS 0.0155f
C1026 OUT5.t20 VSS 0.00776f
C1027 OUT5.n15 VSS 0.00776f
C1028 OUT5.n16 VSS 0.0155f
C1029 OUT5.t40 VSS 0.00776f
C1030 OUT5.n17 VSS 0.00776f
C1031 OUT5.n18 VSS 0.0212f
C1032 OUT5.n19 VSS 0.0639f
C1033 OUT5.n20 VSS 0.0398f
C1034 OUT5.n21 VSS 0.0354f
C1035 OUT5.n22 VSS 0.0695f
C1036 OUT5.t31 VSS 0.00776f
C1037 OUT5.n23 VSS 0.00776f
C1038 OUT5.n24 VSS 0.0155f
C1039 OUT5.t36 VSS 0.00776f
C1040 OUT5.n25 VSS 0.00776f
C1041 OUT5.n26 VSS 0.0155f
C1042 OUT5.t33 VSS 0.00776f
C1043 OUT5.n27 VSS 0.00776f
C1044 OUT5.n28 VSS 0.0155f
C1045 OUT5.t23 VSS 0.00776f
C1046 OUT5.n29 VSS 0.00776f
C1047 OUT5.n30 VSS 0.0214f
C1048 OUT5.n31 VSS 0.0726f
C1049 OUT5.n32 VSS 0.0399f
C1050 OUT5.n33 VSS 0.0376f
C1051 OUT5.t44 VSS 0.00776f
C1052 OUT5.n34 VSS 0.00776f
C1053 OUT5.n35 VSS 0.0155f
C1054 OUT5.t19 VSS 0.00776f
C1055 OUT5.n36 VSS 0.00776f
C1056 OUT5.n37 VSS 0.0155f
C1057 OUT5.t16 VSS 0.00776f
C1058 OUT5.n38 VSS 0.00776f
C1059 OUT5.n39 VSS 0.0155f
C1060 OUT5.t47 VSS 0.00776f
C1061 OUT5.n40 VSS 0.00776f
C1062 OUT5.n41 VSS 0.0212f
C1063 OUT5.n42 VSS 0.0639f
C1064 OUT5.n43 VSS 0.0491f
C1065 OUT5.n44 VSS 0.0609f
C1066 OUT5.n45 VSS 0.0593f
C1067 OUT5.n46 VSS 0.856f
C1068 OUT5.n47 VSS 0.0185f
C1069 OUT5.t1 VSS 0.00776f
C1070 OUT5.n48 VSS 0.00776f
C1071 OUT5.n49 VSS 0.0169f
C1072 OUT5.t5 VSS 0.00776f
C1073 OUT5.n50 VSS 0.00776f
C1074 OUT5.n51 VSS 0.0164f
C1075 OUT5.t6 VSS 0.00776f
C1076 OUT5.n52 VSS 0.00776f
C1077 OUT5.n53 VSS 0.0169f
C1078 OUT5.t4 VSS 0.00776f
C1079 OUT5.n54 VSS 0.00776f
C1080 OUT5.n55 VSS 0.0175f
C1081 OUT5.n56 VSS 0.0247f
C1082 OUT5.n57 VSS 0.103f
C1083 OUT5.t7 VSS 0.00776f
C1084 OUT5.n58 VSS 0.00776f
C1085 OUT5.n59 VSS 0.0164f
C1086 OUT5.t3 VSS 0.00776f
C1087 OUT5.n60 VSS 0.00776f
C1088 OUT5.n61 VSS 0.0169f
C1089 OUT5.t2 VSS 0.0237f
C1090 OUT5.n62 VSS 0.205f
C1091 OUT5.n63 VSS 0.118f
C1092 OUT5.n64 VSS 0.272f
C1093 OUT5.t0 VSS 0.0186f
C1094 OUT5.n65 VSS 0.265f
C1095 OUT5.n66 VSS 0.121f
C1096 OUT5.n67 VSS 0.118f
C1097 OUT5.n68 VSS 0.122f
C1098 OUT5.n69 VSS 0.0949f
C1099 b2.t3 VSS 0.0437f
C1100 b2.n0 VSS 0.0996f
C1101 b2.n1 VSS 0.00542f
C1102 b2.n2 VSS 0.0111f
C1103 b2.n3 VSS 0.00733f
C1104 b2.t6 VSS 0.0659f
C1105 b2.t4 VSS 0.0147f
C1106 b2.n4 VSS 0.0232f
C1107 b2.n5 VSS 0.00477f
C1108 b2.n6 VSS 0.0497f
C1109 b2.n7 VSS 0.0115f
C1110 b2.n8 VSS 0.115f
C1111 b2.t5 VSS 4.33e-19
C1112 b2.t2 VSS 0.0732f
C1113 b2.n9 VSS 0.143f
C1114 b2.n10 VSS 4.25f
C1115 b2.t1 VSS 0.015f
C1116 b2.t0 VSS 0.0119f
C1117 b2.n11 VSS 0.202f
C1118 b2.n12 VSS 3.18f
C1119 b6b.t49 VSS 0.18f
C1120 b6b.t29 VSS 0.0418f
C1121 b6b.n0 VSS 0.209f
C1122 b6b.t46 VSS 0.0418f
C1123 b6b.n1 VSS 0.181f
C1124 b6b.t28 VSS 0.0418f
C1125 b6b.n2 VSS 0.221f
C1126 b6b.n3 VSS 0.333f
C1127 b6b.n4 VSS 0.0159f
C1128 b6b.t20 VSS 0.0239f
C1129 b6b.t21 VSS 0.123f
C1130 b6b.t15 VSS 0.0319f
C1131 b6b.t45 VSS 0.0342f
C1132 b6b.n5 VSS 0.0687f
C1133 b6b.t30 VSS 0.0319f
C1134 b6b.n6 VSS 0.0687f
C1135 b6b.t11 VSS 0.0641f
C1136 b6b.n7 VSS 0.163f
C1137 b6b.t2 VSS 0.0419f
C1138 b6b.n8 VSS 0.0996f
C1139 b6b.n9 VSS 0.102f
C1140 b6b.t44 VSS 0.0319f
C1141 b6b.t26 VSS 0.0342f
C1142 b6b.n10 VSS 0.0693f
C1143 b6b.t27 VSS 0.0319f
C1144 b6b.n11 VSS 0.0693f
C1145 b6b.t9 VSS 0.0641f
C1146 b6b.n12 VSS 0.143f
C1147 b6b.t50 VSS 0.0407f
C1148 b6b.n13 VSS 0.124f
C1149 b6b.n14 VSS 0.0214f
C1150 b6b.n15 VSS 0.0155f
C1151 b6b.n16 VSS 0.0961f
C1152 b6b.t4 VSS 0.125f
C1153 b6b.t39 VSS 0.04f
C1154 b6b.n17 VSS 0.134f
C1155 b6b.t10 VSS 0.04f
C1156 b6b.n18 VSS 0.116f
C1157 b6b.t19 VSS 0.04f
C1158 b6b.n19 VSS 0.131f
C1159 b6b.n20 VSS 0.299f
C1160 b6b.t24 VSS 0.0671f
C1161 b6b.t25 VSS 0.16f
C1162 b6b.t23 VSS 0.0338f
C1163 b6b.t42 VSS 0.0332f
C1164 b6b.n21 VSS 0.0714f
C1165 b6b.t48 VSS 0.0338f
C1166 b6b.n22 VSS 0.0714f
C1167 b6b.t17 VSS 0.062f
C1168 b6b.n23 VSS 0.127f
C1169 b6b.t14 VSS 0.0658f
C1170 b6b.n24 VSS 0.0763f
C1171 b6b.t12 VSS 0.0385f
C1172 b6b.n25 VSS 0.0791f
C1173 b6b.t31 VSS 0.0385f
C1174 b6b.n26 VSS 0.0791f
C1175 b6b.t33 VSS 0.0658f
C1176 b6b.n27 VSS 0.0763f
C1177 b6b.t37 VSS 0.0334f
C1178 b6b.t7 VSS 0.0336f
C1179 b6b.n28 VSS 0.0706f
C1180 b6b.t18 VSS 0.0334f
C1181 b6b.n29 VSS 0.0706f
C1182 b6b.t36 VSS 0.0624f
C1183 b6b.n30 VSS 0.0998f
C1184 b6b.t38 VSS 0.0668f
C1185 b6b.t40 VSS 0.098f
C1186 b6b.n31 VSS 0.131f
C1187 b6b.n32 VSS 0.398f
C1188 b6b.n33 VSS 0.178f
C1189 b6b.n34 VSS 0.0109f
C1190 b6b.n35 VSS 0.0121f
C1191 b6b.n36 VSS 0.125f
C1192 b6b.t43 VSS 0.0249f
C1193 b6b.n37 VSS 0.156f
C1194 b6b.t47 VSS 0.103f
C1195 b6b.t41 VSS 0.0342f
C1196 b6b.t8 VSS 0.0329f
C1197 b6b.n38 VSS 0.0708f
C1198 b6b.t16 VSS 0.0342f
C1199 b6b.n39 VSS 0.0708f
C1200 b6b.t32 VSS 0.0609f
C1201 b6b.n40 VSS 0.111f
C1202 b6b.t34 VSS 0.0439f
C1203 b6b.n41 VSS 0.0709f
C1204 b6b.t5 VSS 0.0439f
C1205 b6b.n42 VSS 0.0709f
C1206 b6b.t6 VSS 0.0314f
C1207 b6b.t22 VSS 0.0357f
C1208 b6b.n43 VSS 0.0695f
C1209 b6b.t35 VSS 0.0314f
C1210 b6b.n44 VSS 0.0695f
C1211 b6b.t3 VSS 0.0637f
C1212 b6b.n45 VSS 0.0883f
C1213 b6b.t13 VSS 0.0439f
C1214 b6b.n46 VSS 0.114f
C1215 b6b.n47 VSS 0.0618f
C1216 b6b.n48 VSS 0.0113f
C1217 b6b.n49 VSS 0.148f
C1218 OUT6.t46 VSS 0.0153f
C1219 OUT6.n0 VSS 0.0153f
C1220 OUT6.n1 VSS 0.0472f
C1221 OUT6.t87 VSS 0.0153f
C1222 OUT6.n2 VSS 0.0153f
C1223 OUT6.n3 VSS 0.0306f
C1224 OUT6.t1 VSS 0.0153f
C1225 OUT6.n4 VSS 0.0153f
C1226 OUT6.n5 VSS 0.0306f
C1227 OUT6.t59 VSS 0.0153f
C1228 OUT6.n6 VSS 0.0153f
C1229 OUT6.n7 VSS 0.0306f
C1230 OUT6.t71 VSS 0.0153f
C1231 OUT6.n8 VSS 0.0153f
C1232 OUT6.n9 VSS 0.0306f
C1233 OUT6.t72 VSS 0.0153f
C1234 OUT6.n10 VSS 0.0153f
C1235 OUT6.n11 VSS 0.0306f
C1236 OUT6.t41 VSS 0.0153f
C1237 OUT6.n12 VSS 0.0153f
C1238 OUT6.n13 VSS 0.0391f
C1239 OUT6.t49 VSS 0.0153f
C1240 OUT6.n14 VSS 0.0153f
C1241 OUT6.n15 VSS 0.0306f
C1242 OUT6.n16 VSS 0.18f
C1243 OUT6.n17 VSS 0.128f
C1244 OUT6.n18 VSS 0.0713f
C1245 OUT6.t67 VSS 0.0153f
C1246 OUT6.n19 VSS 0.0153f
C1247 OUT6.n20 VSS 0.0381f
C1248 OUT6.t85 VSS 0.0153f
C1249 OUT6.n21 VSS 0.0153f
C1250 OUT6.n22 VSS 0.0306f
C1251 OUT6.n23 VSS 0.155f
C1252 OUT6.n24 VSS 0.116f
C1253 OUT6.n25 VSS 0.0513f
C1254 OUT6.n26 VSS 0.0866f
C1255 OUT6.n27 VSS 0.0651f
C1256 OUT6.n28 VSS 0.159f
C1257 OUT6.t93 VSS 0.0153f
C1258 OUT6.n29 VSS 0.0153f
C1259 OUT6.n30 VSS 0.0306f
C1260 OUT6.t63 VSS 0.0153f
C1261 OUT6.n31 VSS 0.0153f
C1262 OUT6.n32 VSS 0.0306f
C1263 OUT6.t82 VSS 0.0153f
C1264 OUT6.n33 VSS 0.0153f
C1265 OUT6.n34 VSS 0.0306f
C1266 OUT6.t52 VSS 0.0153f
C1267 OUT6.n35 VSS 0.0153f
C1268 OUT6.n36 VSS 0.0379f
C1269 OUT6.t2 VSS 0.0153f
C1270 OUT6.n37 VSS 0.0153f
C1271 OUT6.n38 VSS 0.0306f
C1272 OUT6.n39 VSS 0.151f
C1273 OUT6.t39 VSS 0.0153f
C1274 OUT6.n40 VSS 0.0153f
C1275 OUT6.n41 VSS 0.0306f
C1276 OUT6.t56 VSS 0.0153f
C1277 OUT6.n42 VSS 0.0153f
C1278 OUT6.n43 VSS 0.0334f
C1279 OUT6.t95 VSS 0.0153f
C1280 OUT6.n44 VSS 0.0153f
C1281 OUT6.n45 VSS 0.0306f
C1282 OUT6.t91 VSS 0.0153f
C1283 OUT6.n46 VSS 0.0153f
C1284 OUT6.n47 VSS 0.0306f
C1285 OUT6.t0 VSS 0.0153f
C1286 OUT6.n48 VSS 0.0153f
C1287 OUT6.n49 VSS 0.0561f
C1288 OUT6.n50 VSS 0.194f
C1289 OUT6.t86 VSS 0.0153f
C1290 OUT6.n51 VSS 0.0153f
C1291 OUT6.n52 VSS 0.0383f
C1292 OUT6.t76 VSS 0.0153f
C1293 OUT6.n53 VSS 0.0153f
C1294 OUT6.n54 VSS 0.0306f
C1295 OUT6.n55 VSS 0.159f
C1296 OUT6.n56 VSS 0.118f
C1297 OUT6.n57 VSS 0.0307f
C1298 OUT6.n58 VSS 0.0983f
C1299 OUT6.t83 VSS 0.0153f
C1300 OUT6.n59 VSS 0.0153f
C1301 OUT6.n60 VSS 0.0332f
C1302 OUT6.t70 VSS 0.0153f
C1303 OUT6.n61 VSS 0.0153f
C1304 OUT6.n62 VSS 0.0306f
C1305 OUT6.t5 VSS 0.0153f
C1306 OUT6.n63 VSS 0.0153f
C1307 OUT6.n64 VSS 0.0382f
C1308 OUT6.t47 VSS 0.0153f
C1309 OUT6.n65 VSS 0.0153f
C1310 OUT6.n66 VSS 0.0306f
C1311 OUT6.n67 VSS 0.155f
C1312 OUT6.t4 VSS 0.0153f
C1313 OUT6.n68 VSS 0.0153f
C1314 OUT6.n69 VSS 0.0306f
C1315 OUT6.t66 VSS 0.0153f
C1316 OUT6.n70 VSS 0.0153f
C1317 OUT6.n71 VSS 0.0565f
C1318 OUT6.n72 VSS 0.192f
C1319 OUT6.n73 VSS 0.114f
C1320 OUT6.n74 VSS 0.0358f
C1321 OUT6.n75 VSS 0.0816f
C1322 OUT6.n76 VSS 0.298f
C1323 OUT6.t94 VSS 0.0153f
C1324 OUT6.n77 VSS 0.0153f
C1325 OUT6.n78 VSS 0.0306f
C1326 OUT6.t80 VSS 0.0153f
C1327 OUT6.n79 VSS 0.0153f
C1328 OUT6.n80 VSS 0.0392f
C1329 OUT6.t81 VSS 0.0153f
C1330 OUT6.n81 VSS 0.0153f
C1331 OUT6.n82 VSS 0.0306f
C1332 OUT6.n83 VSS 0.175f
C1333 OUT6.n84 VSS 0.107f
C1334 OUT6.n85 VSS 0.0896f
C1335 OUT6.n86 VSS 0.053f
C1336 OUT6.n87 VSS 0.114f
C1337 OUT6.n88 VSS 0.0564f
C1338 OUT6.n89 VSS 0.0876f
C1339 OUT6.n90 VSS 0.061f
C1340 OUT6.t62 VSS 0.0153f
C1341 OUT6.n91 VSS 0.0153f
C1342 OUT6.n92 VSS 0.0491f
C1343 OUT6.n93 VSS 0.181f
C1344 OUT6.n94 VSS 2.19f
C1345 OUT6.n95 VSS 0.0365f
C1346 OUT6.t7 VSS 0.0153f
C1347 OUT6.n96 VSS 0.0153f
C1348 OUT6.n97 VSS 0.0342f
C1349 OUT6.t19 VSS 0.0153f
C1350 OUT6.n98 VSS 0.0153f
C1351 OUT6.n99 VSS 0.0324f
C1352 OUT6.t21 VSS 0.0153f
C1353 OUT6.n100 VSS 0.0153f
C1354 OUT6.n101 VSS 0.0342f
C1355 OUT6.t35 VSS 0.0153f
C1356 OUT6.n102 VSS 0.0153f
C1357 OUT6.n103 VSS 0.0324f
C1358 OUT6.t33 VSS 0.0153f
C1359 OUT6.n104 VSS 0.0153f
C1360 OUT6.n105 VSS 0.0342f
C1361 OUT6.t32 VSS 0.0153f
C1362 OUT6.n106 VSS 0.0153f
C1363 OUT6.n107 VSS 0.0324f
C1364 OUT6.t17 VSS 0.0153f
C1365 OUT6.n108 VSS 0.0153f
C1366 OUT6.n109 VSS 0.0342f
C1367 OUT6.t16 VSS 0.0153f
C1368 OUT6.n110 VSS 0.0153f
C1369 OUT6.n111 VSS 0.0324f
C1370 OUT6.t31 VSS 0.0153f
C1371 OUT6.n112 VSS 0.0153f
C1372 OUT6.n113 VSS 0.0342f
C1373 OUT6.t27 VSS 0.0153f
C1374 OUT6.n114 VSS 0.0153f
C1375 OUT6.n115 VSS 0.0324f
C1376 OUT6.t15 VSS 0.0153f
C1377 OUT6.n116 VSS 0.0153f
C1378 OUT6.n117 VSS 0.0342f
C1379 OUT6.t37 VSS 0.0153f
C1380 OUT6.n118 VSS 0.0153f
C1381 OUT6.n119 VSS 0.0324f
C1382 OUT6.t24 VSS 0.0153f
C1383 OUT6.n120 VSS 0.0153f
C1384 OUT6.n121 VSS 0.0342f
C1385 OUT6.t23 VSS 0.0153f
C1386 OUT6.n122 VSS 0.0153f
C1387 OUT6.n123 VSS 0.0324f
C1388 OUT6.t13 VSS 0.0153f
C1389 OUT6.n124 VSS 0.0153f
C1390 OUT6.n125 VSS 0.0342f
C1391 OUT6.t12 VSS 0.0462f
C1392 OUT6.n126 VSS 0.371f
C1393 OUT6.n127 VSS 0.214f
C1394 OUT6.n128 VSS 0.228f
C1395 OUT6.n129 VSS 0.214f
C1396 OUT6.n130 VSS 0.228f
C1397 OUT6.n131 VSS 0.214f
C1398 OUT6.n132 VSS 0.228f
C1399 OUT6.n133 VSS 0.214f
C1400 OUT6.n134 VSS 0.228f
C1401 OUT6.n135 VSS 0.214f
C1402 OUT6.n136 VSS 0.228f
C1403 OUT6.n137 VSS 0.214f
C1404 OUT6.n138 VSS 0.228f
C1405 OUT6.n139 VSS 0.214f
C1406 OUT6.n140 VSS 0.228f
C1407 OUT6.n141 VSS 0.171f
C1408 IT.t39 VSS 0.0574f
C1409 IT.t53 VSS 0.0219f
C1410 IT.n0 VSS 0.0488f
C1411 IT.t26 VSS 0.0219f
C1412 IT.n1 VSS 0.044f
C1413 IT.t27 VSS 0.0219f
C1414 IT.n2 VSS 0.044f
C1415 IT.t35 VSS 0.0219f
C1416 IT.n3 VSS 0.044f
C1417 IT.t31 VSS 0.0219f
C1418 IT.n4 VSS 0.044f
C1419 IT.t68 VSS 0.0219f
C1420 IT.n5 VSS 0.044f
C1421 IT.t60 VSS 0.0219f
C1422 IT.n6 VSS 0.044f
C1423 IT.t34 VSS 0.0219f
C1424 IT.n7 VSS 0.044f
C1425 IT.t36 VSS 0.0219f
C1426 IT.n8 VSS 0.044f
C1427 IT.t71 VSS 0.0219f
C1428 IT.n9 VSS 0.044f
C1429 IT.t25 VSS 0.0219f
C1430 IT.n10 VSS 0.044f
C1431 IT.t52 VSS 0.0219f
C1432 IT.n11 VSS 0.044f
C1433 IT.t42 VSS 0.0219f
C1434 IT.n12 VSS 0.044f
C1435 IT.t29 VSS 0.0219f
C1436 IT.n13 VSS 0.0443f
C1437 IT.n14 VSS 0.0244f
C1438 IT.n15 VSS 0.00799f
C1439 IT.t65 VSS 0.0156f
C1440 IT.n16 VSS 0.0156f
C1441 IT.n17 VSS 0.0063f
C1442 IT.n18 VSS 0.0358f
C1443 IT.n19 VSS 0.00831f
C1444 IT.t54 VSS 0.0172f
C1445 IT.n20 VSS 0.0148f
C1446 IT.t63 VSS 0.0219f
C1447 IT.t62 VSS 0.0219f
C1448 IT.t40 VSS 0.0219f
C1449 IT.t46 VSS 0.0219f
C1450 IT.t61 VSS 0.0219f
C1451 IT.t69 VSS 0.0219f
C1452 IT.t32 VSS 0.0219f
C1453 IT.t33 VSS 0.0219f
C1454 IT.t59 VSS 0.0219f
C1455 IT.t66 VSS 0.0219f
C1456 IT.t30 VSS 0.0219f
C1457 IT.n21 VSS 0.044f
C1458 IT.n22 VSS 0.044f
C1459 IT.n23 VSS 0.044f
C1460 IT.n24 VSS 0.044f
C1461 IT.n25 VSS 0.044f
C1462 IT.n26 VSS 0.044f
C1463 IT.n27 VSS 0.044f
C1464 IT.n28 VSS 0.044f
C1465 IT.n29 VSS 0.044f
C1466 IT.n30 VSS 0.044f
C1467 IT.n31 VSS 0.044f
C1468 IT.n32 VSS 0.00995f
C1469 IT.n33 VSS 0.00589f
C1470 IT.n34 VSS 0.00754f
C1471 IT.n35 VSS 0.234f
C1472 IT.t45 VSS 0.0214f
C1473 IT.t44 VSS 0.0214f
C1474 IT.n36 VSS 0.0435f
C1475 IT.n37 VSS 0.0437f
C1476 IT.t50 VSS 0.0208f
C1477 IT.n38 VSS 0.0347f
C1478 IT.t6 VSS 0.0135f
C1479 IT.t24 VSS 0.0219f
C1480 IT.n39 VSS 0.044f
C1481 IT.t51 VSS 0.0219f
C1482 IT.n40 VSS 0.044f
C1483 IT.t37 VSS 0.0219f
C1484 IT.n41 VSS 0.0444f
C1485 IT.n42 VSS 0.00964f
C1486 IT.t73 VSS 0.0173f
C1487 IT.n43 VSS 0.0146f
C1488 IT.n44 VSS 0.00811f
C1489 IT.n45 VSS 0.00588f
C1490 IT.n46 VSS 0.108f
C1491 IT.t74 VSS 0.0179f
C1492 IT.n47 VSS 0.131f
C1493 IT.t41 VSS 0.0215f
C1494 IT.n48 VSS 0.044f
C1495 IT.t49 VSS 0.0215f
C1496 IT.n49 VSS 0.0436f
C1497 IT.t72 VSS 0.0215f
C1498 IT.n50 VSS 0.0462f
C1499 IT.n51 VSS 0.0293f
C1500 IT.n52 VSS 0.0447f
C1501 IT.n53 VSS 0.0461f
C1502 IT.t12 VSS 0.0199f
C1503 IT.n54 VSS 0.0472f
C1504 IT.t13 VSS 0.0061f
C1505 IT.n55 VSS 0.0061f
C1506 IT.n56 VSS 0.0332f
C1507 IT.n57 VSS 0.0264f
C1508 IT.t4 VSS 0.0199f
C1509 IT.n58 VSS 0.0461f
C1510 IT.t2 VSS 0.0195f
C1511 IT.n59 VSS 0.043f
C1512 IT.n60 VSS 0.00275f
C1513 IT.n61 VSS 0.00258f
C1514 IT.t75 VSS 0.0215f
C1515 IT.n62 VSS 0.0464f
C1516 IT.n63 VSS 0.012f
C1517 IT.t3 VSS 0.0153f
C1518 IT.n64 VSS 0.0266f
C1519 IT.n65 VSS 0.0205f
C1520 IT.n66 VSS 5.16e-19
C1521 IT.n67 VSS 0.00604f
C1522 IT.n68 VSS 0.179f
C1523 IT.t11 VSS 0.0061f
C1524 IT.n69 VSS 0.0061f
C1525 IT.n70 VSS 0.0131f
C1526 IT.t10 VSS 0.0196f
C1527 IT.t58 VSS 0.0369f
C1528 IT.t47 VSS 0.0214f
C1529 IT.n71 VSS 0.0535f
C1530 IT.t38 VSS 0.0214f
C1531 IT.n72 VSS 0.0435f
C1532 IT.t48 VSS 0.0214f
C1533 IT.n73 VSS 0.0483f
C1534 IT.n74 VSS 0.0511f
C1535 IT.t8 VSS 0.0196f
C1536 IT.n75 VSS 0.0462f
C1537 IT.n76 VSS 0.00957f
C1538 IT.n77 VSS 0.0908f
C1539 IT.n78 VSS 0.46f
C1540 IT.t43 VSS 0.0214f
C1541 IT.n79 VSS 0.0485f
C1542 IT.t0 VSS 0.02f
C1543 IT.n80 VSS 0.0503f
C1544 IT.t14 VSS 0.02f
C1545 IT.n81 VSS 0.0454f
C1546 IT.n82 VSS 0.00842f
C1547 IT.n83 VSS 0.0128f
C1548 IT.t15 VSS 0.0061f
C1549 IT.n84 VSS 0.0061f
C1550 IT.n85 VSS 0.0132f
C1551 IT.n86 VSS 0.0224f
C1552 IT.n87 VSS 0.00777f
C1553 IT.n88 VSS 0.119f
C1554 IT.n89 VSS 0.455f
C1555 IT.n90 VSS 0.281f
C1556 IT.t17 VSS 0.0061f
C1557 IT.n91 VSS 0.0061f
C1558 IT.n92 VSS 0.013f
C1559 IT.t18 VSS 0.0061f
C1560 IT.n93 VSS 0.0061f
C1561 IT.n94 VSS 0.013f
C1562 IT.t19 VSS 0.0061f
C1563 IT.n95 VSS 0.0061f
C1564 IT.n96 VSS 0.0328f
C1565 IT.t20 VSS 0.0061f
C1566 IT.n97 VSS 0.0061f
C1567 IT.n98 VSS 0.013f
C1568 IT.n99 VSS 0.362f
C1569 IT.n100 VSS 0.521f
C1570 IT.n101 VSS 0.595f
C1571 IT.n102 VSS 1.23f
C1572 IT.n103 VSS 0.183f
C1573 IT.n104 VSS 0.0156f
C1574 IT.n105 VSS 0.00906f
C1575 IT.t64 VSS 0.0215f
C1576 IT.t28 VSS 0.0215f
C1577 IT.n106 VSS 0.0436f
C1578 IT.n107 VSS 0.0437f
C1579 IT.t55 VSS 0.0209f
C1580 IT.n108 VSS 0.0436f
C1581 IT.n109 VSS 0.00264f
C1582 IT.n110 VSS 3.2e-19
C1583 OUT-.t125 VSS 0.0246f
C1584 OUT-.t41 VSS 0.0246f
C1585 OUT-.n0 VSS 0.0203f
C1586 OUT-.t14 VSS 0.0249f
C1587 OUT-.n1 VSS 0.0199f
C1588 OUT-.t74 VSS 0.0147f
C1589 OUT-.n2 VSS 0.0147f
C1590 OUT-.n3 VSS 0.0294f
C1591 OUT-.t93 VSS 0.0147f
C1592 OUT-.n4 VSS 0.0147f
C1593 OUT-.n5 VSS 0.0295f
C1594 OUT-.t71 VSS 0.028f
C1595 OUT-.t73 VSS 0.0314f
C1596 OUT-.n6 VSS 0.124f
C1597 OUT-.t21 VSS 0.025f
C1598 OUT-.t19 VSS 0.0254f
C1599 OUT-.n7 VSS 0.0193f
C1600 OUT-.n8 VSS 0.11f
C1601 OUT-.n9 VSS 0.123f
C1602 OUT-.t162 VSS 0.0181f
C1603 OUT-.t118 VSS 0.0275f
C1604 OUT-.n10 VSS 0.0588f
C1605 OUT-.n11 VSS 0.0281f
C1606 OUT-.t163 VSS 0.025f
C1607 OUT-.t9 VSS 0.0251f
C1608 OUT-.n12 VSS 0.0202f
C1609 OUT-.n13 VSS 0.0417f
C1610 OUT-.n14 VSS 0.0405f
C1611 OUT-.t119 VSS 0.0253f
C1612 OUT-.t72 VSS 0.0252f
C1613 OUT-.n15 VSS 0.0193f
C1614 OUT-.n16 VSS 0.119f
C1615 OUT-.t44 VSS 0.0147f
C1616 OUT-.n17 VSS 0.0147f
C1617 OUT-.n18 VSS 0.0359f
C1618 OUT-.t51 VSS 0.0147f
C1619 OUT-.n19 VSS 0.0147f
C1620 OUT-.n20 VSS 0.0294f
C1621 OUT-.n21 VSS 0.13f
C1622 OUT-.t128 VSS 0.0664f
C1623 OUT-.n22 VSS 0.189f
C1624 OUT-.t129 VSS 0.0521f
C1625 OUT-.n23 VSS 0.0147f
C1626 OUT-.n24 VSS 0.0294f
C1627 OUT-.n25 VSS 0.153f
C1628 OUT-.n26 VSS 0.352f
C1629 OUT-.t99 VSS 0.0495f
C1630 OUT-.n27 VSS 0.0147f
C1631 OUT-.n28 VSS 0.0294f
C1632 OUT-.n29 VSS 0.0653f
C1633 OUT-.t98 VSS 0.0816f
C1634 OUT-.n30 VSS 0.156f
C1635 OUT-.n31 VSS 0.0554f
C1636 OUT-.t146 VSS 0.0689f
C1637 OUT-.n32 VSS 0.178f
C1638 OUT-.t132 VSS 0.059f
C1639 OUT-.n33 VSS 0.174f
C1640 OUT-.t94 VSS 0.0147f
C1641 OUT-.t133 VSS 0.0514f
C1642 OUT-.n34 VSS 0.0294f
C1643 OUT-.n35 VSS 0.21f
C1644 OUT-.t52 VSS 0.0147f
C1645 OUT-.t147 VSS 0.0514f
C1646 OUT-.n36 VSS 0.0294f
C1647 OUT-.n37 VSS 0.239f
C1648 OUT-.n38 VSS 0.0489f
C1649 OUT-.n39 VSS 0.144f
C1650 OUT-.n40 VSS 0.148f
C1651 OUT-.t36 VSS 0.0496f
C1652 OUT-.t35 VSS 0.0496f
C1653 OUT-.n41 VSS 0.0313f
C1654 OUT-.t34 VSS 0.0496f
C1655 OUT-.t30 VSS 0.0496f
C1656 OUT-.n42 VSS 0.0294f
C1657 OUT-.t153 VSS 0.0506f
C1658 OUT-.n43 VSS 0.0147f
C1659 OUT-.n44 VSS 0.0318f
C1660 OUT-.t123 VSS 0.05f
C1661 OUT-.t173 VSS 0.0518f
C1662 OUT-.n45 VSS 0.0316f
C1663 OUT-.t172 VSS 0.0623f
C1664 OUT-.n46 VSS 0.159f
C1665 OUT-.n47 VSS 0.0777f
C1666 OUT-.t122 VSS 0.0623f
C1667 OUT-.n48 VSS 0.0767f
C1668 OUT-.n49 VSS 0.0934f
C1669 OUT-.n50 VSS 0.105f
C1670 OUT-.t152 VSS 0.0633f
C1671 OUT-.n51 VSS 0.0741f
C1672 OUT-.n52 VSS 0.0791f
C1673 OUT-.t59 VSS 0.0147f
C1674 OUT-.n53 VSS 0.0147f
C1675 OUT-.n54 VSS 0.0294f
C1676 OUT-.t60 VSS 0.0147f
C1677 OUT-.n55 VSS 0.0147f
C1678 OUT-.n56 VSS 0.0294f
C1679 OUT-.t7 VSS 0.0147f
C1680 OUT-.n57 VSS 0.0147f
C1681 OUT-.n58 VSS 0.0294f
C1682 OUT-.t111 VSS 0.0497f
C1683 OUT-.n59 VSS 0.0147f
C1684 OUT-.n60 VSS 0.0294f
C1685 OUT-.t182 VSS 0.0147f
C1686 OUT-.t131 VSS 0.0519f
C1687 OUT-.n61 VSS 0.0316f
C1688 OUT-.t130 VSS 0.065f
C1689 OUT-.n62 VSS 0.166f
C1690 OUT-.n63 VSS 0.281f
C1691 OUT-.t165 VSS 0.0496f
C1692 OUT-.t135 VSS 0.0515f
C1693 OUT-.n64 VSS 0.0312f
C1694 OUT-.t134 VSS 0.0587f
C1695 OUT-.n65 VSS 0.16f
C1696 OUT-.n66 VSS 0.0738f
C1697 OUT-.t164 VSS 0.0585f
C1698 OUT-.n67 VSS 0.077f
C1699 OUT-.n68 VSS 0.0945f
C1700 OUT-.n69 VSS 0.0944f
C1701 OUT-.t110 VSS 0.0585f
C1702 OUT-.n70 VSS 0.0764f
C1703 OUT-.n71 VSS 0.249f
C1704 OUT-.n72 VSS 0.0824f
C1705 OUT-.t67 VSS 0.0147f
C1706 OUT-.n73 VSS 0.0147f
C1707 OUT-.n74 VSS 0.0728f
C1708 OUT-.n75 VSS 0.321f
C1709 OUT-.n76 VSS 0.0832f
C1710 OUT-.n77 VSS 0.0871f
C1711 OUT-.t58 VSS 0.0147f
C1712 OUT-.n78 VSS 0.0147f
C1713 OUT-.n79 VSS 0.0301f
C1714 OUT-.t27 VSS 0.0147f
C1715 OUT-.n80 VSS 0.0147f
C1716 OUT-.n81 VSS 0.0315f
C1717 OUT-.n82 VSS 0.136f
C1718 OUT-.n83 VSS 0.284f
C1719 OUT-.n84 VSS 0.126f
C1720 OUT-.t8 VSS 0.0147f
C1721 OUT-.t167 VSS 0.0525f
C1722 OUT-.n85 VSS 0.0322f
C1723 OUT-.t166 VSS 0.0672f
C1724 OUT-.n86 VSS 0.17f
C1725 OUT-.n87 VSS 0.139f
C1726 OUT-.t31 VSS 0.0495f
C1727 OUT-.t33 VSS 0.0495f
C1728 OUT-.n88 VSS 0.0309f
C1729 OUT-.n89 VSS 0.155f
C1730 OUT-.n90 VSS 0.158f
C1731 OUT-.n91 VSS 0.111f
C1732 OUT-.t32 VSS 0.0495f
C1733 OUT-.t29 VSS 0.0497f
C1734 OUT-.n92 VSS 0.0294f
C1735 OUT-.n93 VSS 0.0447f
C1736 OUT-.n94 VSS 0.135f
C1737 OUT-.n95 VSS 0.157f
C1738 OUT-.n96 VSS 0.121f
C1739 OUT-.n97 VSS 0.0405f
C1740 OUT-.n98 VSS 0.565f
C1741 OUT-.n99 VSS 0.562f
C1742 OUT-.n100 VSS 0.226f
C1743 OUT-.t78 VSS 0.0481f
C1744 OUT-.n101 VSS 0.0303f
C1745 OUT-.t80 VSS 0.0481f
C1746 OUT-.t85 VSS 0.0481f
C1747 OUT-.t55 VSS 0.0147f
C1748 OUT-.n102 VSS 0.0147f
C1749 OUT-.n103 VSS 0.0335f
C1750 OUT-.t127 VSS 0.0495f
C1751 OUT-.n104 VSS 0.0147f
C1752 OUT-.n105 VSS 0.0309f
C1753 OUT-.t177 VSS 0.0561f
C1754 OUT-.t151 VSS 0.0536f
C1755 OUT-.n106 VSS 0.0377f
C1756 OUT-.t150 VSS 0.0822f
C1757 OUT-.t176 VSS 0.0407f
C1758 OUT-.n107 VSS 0.0976f
C1759 OUT-.n108 VSS 0.192f
C1760 OUT-.n109 VSS 0.0917f
C1761 OUT-.n110 VSS 0.0907f
C1762 OUT-.t126 VSS 0.0559f
C1763 OUT-.n111 VSS 0.0707f
C1764 OUT-.n112 VSS 0.104f
C1765 OUT-.t42 VSS 0.0147f
C1766 OUT-.n113 VSS 0.0147f
C1767 OUT-.n114 VSS 0.0317f
C1768 OUT-.t25 VSS 0.0147f
C1769 OUT-.n115 VSS 0.0147f
C1770 OUT-.n116 VSS 0.0323f
C1771 OUT-.n117 VSS 0.102f
C1772 OUT-.t141 VSS 0.0503f
C1773 OUT-.n118 VSS 0.144f
C1774 OUT-.t108 VSS 0.0435f
C1775 OUT-.t116 VSS 0.0485f
C1776 OUT-.n119 VSS 0.077f
C1777 OUT-.n120 VSS 0.0266f
C1778 OUT-.t109 VSS 0.0497f
C1779 OUT-.n121 VSS 0.0319f
C1780 OUT-.n122 VSS 0.062f
C1781 OUT-.t117 VSS 0.0499f
C1782 OUT-.n123 VSS 0.0322f
C1783 OUT-.n124 VSS 0.065f
C1784 OUT-.t140 VSS 0.0445f
C1785 OUT-.t144 VSS 0.0475f
C1786 OUT-.n125 VSS 0.077f
C1787 OUT-.n126 VSS 0.0247f
C1788 OUT-.t145 VSS 0.0505f
C1789 OUT-.n127 VSS 0.0813f
C1790 OUT-.n128 VSS 0.0839f
C1791 OUT-.n129 VSS 0.153f
C1792 OUT-.t168 VSS 0.044f
C1793 OUT-.t174 VSS 0.048f
C1794 OUT-.n130 VSS 0.077f
C1795 OUT-.n131 VSS 0.0269f
C1796 OUT-.t169 VSS 0.0497f
C1797 OUT-.n132 VSS 0.0147f
C1798 OUT-.n133 VSS 0.0319f
C1799 OUT-.n134 VSS 0.0636f
C1800 OUT-.t175 VSS 0.0499f
C1801 OUT-.n135 VSS 0.0147f
C1802 OUT-.n136 VSS 0.0294f
C1803 OUT-.t65 VSS 0.0147f
C1804 OUT-.n137 VSS 0.0147f
C1805 OUT-.n138 VSS 0.0377f
C1806 OUT-.t22 VSS 0.0147f
C1807 OUT-.n139 VSS 0.0147f
C1808 OUT-.n140 VSS 0.0294f
C1809 OUT-.n141 VSS 0.112f
C1810 OUT-.t56 VSS 0.0147f
C1811 OUT-.t149 VSS 0.0497f
C1812 OUT-.n142 VSS 0.0312f
C1813 OUT-.t148 VSS 0.045f
C1814 OUT-.t154 VSS 0.0471f
C1815 OUT-.n143 VSS 0.0763f
C1816 OUT-.n144 VSS 0.147f
C1817 OUT-.n145 VSS 0.0352f
C1818 OUT-.n146 VSS 0.0851f
C1819 OUT-.t49 VSS 0.0147f
C1820 OUT-.t155 VSS 0.0499f
C1821 OUT-.n147 VSS 0.0294f
C1822 OUT-.n148 VSS 0.0927f
C1823 OUT-.t46 VSS 0.0147f
C1824 OUT-.n149 VSS 0.0147f
C1825 OUT-.n150 VSS 0.0294f
C1826 OUT-.t37 VSS 0.0147f
C1827 OUT-.n151 VSS 0.0147f
C1828 OUT-.n152 VSS 0.0365f
C1829 OUT-.n153 VSS 0.1f
C1830 OUT-.n154 VSS 0.147f
C1831 OUT-.n155 VSS 0.119f
C1832 OUT-.t24 VSS 0.0147f
C1833 OUT-.n156 VSS 0.0147f
C1834 OUT-.n157 VSS 0.0294f
C1835 OUT-.t137 VSS 0.0499f
C1836 OUT-.n158 VSS 0.0147f
C1837 OUT-.n159 VSS 0.0336f
C1838 OUT-.t102 VSS 0.0819f
C1839 OUT-.t156 VSS 0.0395f
C1840 OUT-.n160 VSS 0.092f
C1841 OUT-.n161 VSS 0.111f
C1842 OUT-.t136 VSS 0.074f
C1843 OUT-.n162 VSS 0.141f
C1844 OUT-.n163 VSS 0.105f
C1845 OUT-.n164 VSS 0.0635f
C1846 OUT-.t157 VSS 0.051f
C1847 OUT-.t103 VSS 0.0494f
C1848 OUT-.n165 VSS 0.0294f
C1849 OUT-.n166 VSS 0.125f
C1850 OUT-.n167 VSS 0.231f
C1851 OUT-.t18 VSS 0.0147f
C1852 OUT-.n168 VSS 0.0147f
C1853 OUT-.n169 VSS 0.0335f
C1854 OUT-.t64 VSS 0.0147f
C1855 OUT-.t113 VSS 0.051f
C1856 OUT-.n170 VSS 0.0307f
C1857 OUT-.t112 VSS 0.0558f
C1858 OUT-.n171 VSS 0.155f
C1859 OUT-.n172 VSS 0.172f
C1860 OUT-.n173 VSS 0.21f
C1861 OUT-.n174 VSS 0.287f
C1862 OUT-.t3 VSS 0.0147f
C1863 OUT-.n175 VSS 0.0147f
C1864 OUT-.n176 VSS 0.0315f
C1865 OUT-.n177 VSS 0.232f
C1866 OUT-.n178 VSS 0.0359f
C1867 OUT-.n179 VSS 0.147f
C1868 OUT-.n180 VSS 0.0969f
C1869 OUT-.n181 VSS 0.0713f
C1870 OUT-.t69 VSS 0.0147f
C1871 OUT-.n182 VSS 0.0147f
C1872 OUT-.n183 VSS 0.0319f
C1873 OUT-.t47 VSS 0.0147f
C1874 OUT-.n184 VSS 0.0147f
C1875 OUT-.n185 VSS 0.0312f
C1876 OUT-.n186 VSS 0.168f
C1877 OUT-.n187 VSS 0.448f
C1878 OUT-.n188 VSS 0.244f
C1879 OUT-.n189 VSS 0.165f
C1880 OUT-.n190 VSS 0.181f
C1881 OUT-.t16 VSS 0.0147f
C1882 OUT-.t101 VSS 0.0488f
C1883 OUT-.n191 VSS 0.0294f
C1884 OUT-.t100 VSS 0.073f
C1885 OUT-.n192 VSS 0.171f
C1886 OUT-.n193 VSS 0.0992f
C1887 OUT-.n194 VSS 0.199f
C1888 OUT-.n195 VSS 0.144f
C1889 OUT-.t81 VSS 0.0481f
C1890 OUT-.n196 VSS 0.0306f
C1891 OUT-.n197 VSS 0.0891f
C1892 OUT-.t88 VSS 0.0491f
C1893 OUT-.n198 VSS 0.112f
C1894 OUT-.n199 VSS 0.0769f
C1895 OUT-.t84 VSS 0.0481f
C1896 OUT-.n200 VSS 0.0314f
C1897 OUT-.t75 VSS 0.0481f
C1898 OUT-.n201 VSS 0.0309f
C1899 OUT-.t82 VSS 0.0497f
C1900 OUT-.n202 VSS 0.0304f
C1901 OUT-.t79 VSS 0.0499f
C1902 OUT-.t159 VSS 0.0493f
C1903 OUT-.n203 VSS 0.0306f
C1904 OUT-.t105 VSS 0.0498f
C1905 OUT-.n204 VSS 0.0312f
C1906 OUT-.n205 VSS 0.133f
C1907 OUT-.t158 VSS 0.0367f
C1908 OUT-.t104 VSS 0.0466f
C1909 OUT-.n206 VSS 0.0683f
C1910 OUT-.n207 VSS 0.0362f
C1911 OUT-.n208 VSS 0.113f
C1912 OUT-.t83 VSS 0.05f
C1913 OUT-.n209 VSS 0.0831f
C1914 OUT-.n210 VSS 0.193f
C1915 OUT-.n211 VSS 0.209f
C1916 OUT-.n212 VSS 0.084f
C1917 OUT-.t77 VSS 0.0481f
C1918 OUT-.n213 VSS 0.114f
C1919 OUT-.n214 VSS 0.0904f
C1920 OUT-.t90 VSS 0.0715f
C1921 OUT-.t86 VSS 0.0545f
C1922 OUT-.n215 VSS 0.145f
C1923 OUT-.n216 VSS 0.226f
C1924 OUT-.n217 VSS 0.057f
C1925 OUT-.n218 VSS 0.126f
C1926 OUT-.n219 VSS 0.0572f
C1927 OUT-.n220 VSS 0.0904f
C1928 OUT-.n221 VSS 0.112f
C1929 OUT-.n222 VSS 0.0861f
C1930 OUT-.t89 VSS 0.049f
C1931 OUT-.n223 VSS 0.0859f
C1932 OUT-.t87 VSS 0.0495f
C1933 OUT-.t76 VSS 0.0494f
C1934 OUT-.n224 VSS 0.122f
C1935 OUT-.t107 VSS 0.0495f
C1936 OUT-.n225 VSS 0.0309f
C1937 OUT-.t143 VSS 0.0496f
C1938 OUT-.n226 VSS 0.031f
C1939 OUT-.t106 VSS 0.0414f
C1940 OUT-.t142 VSS 0.0419f
C1941 OUT-.n227 VSS 0.0683f
C1942 OUT-.n228 VSS 0.132f
C1943 OUT-.n229 VSS 0.0323f
C1944 OUT-.n230 VSS 0.112f
C1945 OUT-.n231 VSS 0.0771f
C1946 OUT-.n232 VSS 0.364f
C1947 OUT-.n233 VSS 0.349f
C1948 OUT-.t6 VSS 0.0403f
C1949 OUT-.t10 VSS 0.0358f
C1950 OUT-.n234 VSS 0.206f
C1951 OUT-.n235 VSS 0.122f
C1952 OUT-.n236 VSS 0.142f
C1953 OUT-.n237 VSS 0.074f
C1954 OUT-.n238 VSS 0.0254f
C1955 OUT-.n239 VSS 0.0969f
C1956 OUT-.n240 VSS 0.475f
C1957 OUT-.n241 VSS 0.163f
C1958 OUT-.n242 VSS 0.111f
C1959 OUT-.n243 VSS 0.107f
C1960 OUT-.n244 VSS 0.0885f
C1961 OUT-.t15 VSS 0.0335f
C1962 OUT-.t96 VSS 0.0339f
C1963 OUT-.n245 VSS 0.111f
C1964 OUT-.n246 VSS 0.116f
C1965 OUT-.n247 VSS 0.176f
C1966 OUT-.n248 VSS 0.176f
C1967 OUT-.n249 VSS 0.0535f
C1968 OUT-.n250 VSS 0.0532f
C1969 OUT-.t124 VSS 0.0184f
C1970 OUT-.t170 VSS 0.0254f
C1971 OUT-.n251 VSS 0.057f
C1972 OUT-.n252 VSS 0.0274f
C1973 OUT-.t171 VSS 0.0246f
C1974 OUT-.t161 VSS 0.05f
C1975 OUT-.t139 VSS 0.0294f
C1976 OUT-.n253 VSS 0.0312f
C1977 OUT-.n254 VSS 0.0147f
C1978 OUT-.n255 VSS 0.0302f
C1979 OUT-.t114 VSS 0.0442f
C1980 OUT-.t115 VSS 0.0354f
C1981 OUT-.n256 VSS 0.257f
C1982 OUT-.t91 VSS 0.0328f
C1983 OUT-.n257 VSS 0.222f
C1984 OUT-.n258 VSS 0.165f
C1985 OUT-.t121 VSS 0.0294f
C1986 OUT-.n259 VSS 0.0307f
C1987 OUT-.n260 VSS 0.0668f
C1988 OUT-.t138 VSS 0.0217f
C1989 OUT-.t160 VSS 0.083f
C1990 OUT-.n261 VSS 0.103f
C1991 OUT-.t120 VSS 0.0601f
C1992 OUT-.n262 VSS 0.0714f
C1993 OUT-.n263 VSS 0.0422f
C1994 OUT-.n264 VSS 0.0812f
C1995 OUT-.n265 VSS 0.119f
C1996 OUT-.t5 VSS 0.0147f
C1997 OUT-.n266 VSS 0.0147f
C1998 OUT-.n267 VSS 0.0734f
C1999 OUT-.t57 VSS 0.0341f
C2000 OUT-.t178 VSS 0.04f
C2001 OUT-.t179 VSS 0.0341f
C2002 OUT-.n268 VSS 0.203f
C2003 OUT-.n269 VSS 0.162f
C2004 OUT-.n270 VSS 0.404f
C2005 OUT-.t26 VSS 0.0333f
C2006 OUT-.n271 VSS 0.243f
C2007 OUT-.n272 VSS 0.145f
C2008 OUT-.n273 VSS 0.05f
C2009 OUT-.n274 VSS 0.0482f
C2010 OUT-.n275 VSS 0.233f
C2011 b6.t38 VSS 0.0391f
C2012 b6.t18 VSS 0.0583f
C2013 b6.t37 VSS 0.136f
C2014 b6.t28 VSS 0.04f
C2015 b6.n0 VSS 0.113f
C2016 b6.t41 VSS 0.04f
C2017 b6.n1 VSS 0.0863f
C2018 b6.t45 VSS 0.0583f
C2019 b6.t17 VSS 0.0878f
C2020 b6.n2 VSS 0.0874f
C2021 b6.t16 VSS 0.0583f
C2022 b6.t36 VSS 0.0878f
C2023 b6.n3 VSS 0.088f
C2024 b6.n4 VSS 0.081f
C2025 b6.t9 VSS 0.0391f
C2026 b6.t43 VSS 0.0583f
C2027 b6.t14 VSS 0.137f
C2028 b6.n5 VSS 0.11f
C2029 b6.n6 VSS 0.0655f
C2030 b6.t2 VSS 0.0668f
C2031 b6.t15 VSS 0.0413f
C2032 b6.n7 VSS 0.23f
C2033 b6.t12 VSS 0.0413f
C2034 b6.n8 VSS 0.181f
C2035 b6.t32 VSS 0.0546f
C2036 b6.n9 VSS 0.0701f
C2037 b6.n10 VSS 0.566f
C2038 b6.t25 VSS 0.0592f
C2039 b6.t6 VSS 0.116f
C2040 b6.t49 VSS 0.0404f
C2041 b6.n11 VSS 0.112f
C2042 b6.t27 VSS 0.0404f
C2043 b6.n12 VSS 0.0751f
C2044 b6.t48 VSS 0.0625f
C2045 b6.n13 VSS 0.0767f
C2046 b6.t20 VSS 0.0326f
C2047 b6.n14 VSS 0.0694f
C2048 b6.t47 VSS 0.0326f
C2049 b6.n15 VSS 0.0694f
C2050 b6.t30 VSS 0.0625f
C2051 b6.n16 VSS 0.0767f
C2052 b6.t8 VSS 0.0404f
C2053 b6.n17 VSS 0.0751f
C2054 b6.t35 VSS 0.0404f
C2055 b6.n18 VSS 0.0751f
C2056 b6.t11 VSS 0.0592f
C2057 b6.t40 VSS 0.0892f
C2058 b6.n19 VSS 0.107f
C2059 b6.n20 VSS 0.53f
C2060 b6.n21 VSS 0.175f
C2061 b6.t42 VSS 0.0676f
C2062 b6.t23 VSS 0.0415f
C2063 b6.n22 VSS 0.17f
C2064 b6.t4 VSS 0.0415f
C2065 b6.n23 VSS 0.133f
C2066 b6.t29 VSS 0.0415f
C2067 b6.n24 VSS 0.136f
C2068 b6.t44 VSS 0.0383f
C2069 b6.n25 VSS 0.0935f
C2070 b6.n26 VSS 0.00126f
C2071 b6.t0 VSS 0.0125f
C2072 b6.t1 VSS 0.00523f
C2073 b6.n27 VSS 0.203f
C2074 b6.n28 VSS 0.201f
C2075 b6.n29 VSS 0.0122f
C2076 b6.n30 VSS 0.532f
C2077 b6.n31 VSS 0.673f
C2078 b6.n32 VSS 0.0166f
C2079 b6.t39 VSS 0.059f
C2080 b6.t24 VSS 0.149f
C2081 b6.t22 VSS 0.036f
C2082 b6.t21 VSS 0.0348f
C2083 b6.n33 VSS 0.0778f
C2084 b6.t3 VSS 0.036f
C2085 b6.n34 VSS 0.0778f
C2086 b6.t50 VSS 0.063f
C2087 b6.n35 VSS 0.124f
C2088 b6.t19 VSS 0.0639f
C2089 b6.n36 VSS 0.0743f
C2090 b6.t34 VSS 0.0317f
C2091 b6.n37 VSS 0.0671f
C2092 b6.t13 VSS 0.0317f
C2093 b6.n38 VSS 0.0671f
C2094 b6.t46 VSS 0.0639f
C2095 b6.n39 VSS 0.0743f
C2096 b6.t7 VSS 0.0351f
C2097 b6.t5 VSS 0.0357f
C2098 b6.n40 VSS 0.076f
C2099 b6.t33 VSS 0.0351f
C2100 b6.n41 VSS 0.076f
C2101 b6.t31 VSS 0.0639f
C2102 b6.n42 VSS 0.0971f
C2103 b6.t26 VSS 0.0592f
C2104 b6.t10 VSS 0.0898f
C2105 b6.n43 VSS 0.125f
C2106 b6.n44 VSS 0.0708f
C2107 b6.n46 VSS 0.139f
C2108 SD3_1.t52 VSS 0.00898f
C2109 SD3_1.n0 VSS 0.00898f
C2110 SD3_1.n1 VSS 0.0372f
C2111 SD3_1.t28 VSS 0.00898f
C2112 SD3_1.n2 VSS 0.00898f
C2113 SD3_1.n3 VSS 0.0342f
C2114 SD3_1.t38 VSS 0.00898f
C2115 SD3_1.n4 VSS 0.00898f
C2116 SD3_1.n5 VSS 0.0371f
C2117 SD3_1.t20 VSS 0.00898f
C2118 SD3_1.n6 VSS 0.00898f
C2119 SD3_1.n7 VSS 0.0343f
C2120 SD3_1.t57 VSS 0.00898f
C2121 SD3_1.n8 VSS 0.00898f
C2122 SD3_1.n9 VSS 0.018f
C2123 SD3_1.n10 VSS 0.0222f
C2124 SD3_1.n11 VSS 0.00975f
C2125 SD3_1.t58 VSS 0.0083f
C2126 SD3_1.n12 VSS 0.0363f
C2127 SD3_1.t24 VSS 0.00898f
C2128 SD3_1.n13 VSS 0.00898f
C2129 SD3_1.n14 VSS 0.018f
C2130 SD3_1.n15 VSS 0.0161f
C2131 SD3_1.t23 VSS 0.00898f
C2132 SD3_1.n16 VSS 0.00898f
C2133 SD3_1.n17 VSS 0.0372f
C2134 SD3_1.t39 VSS 0.00898f
C2135 SD3_1.n18 VSS 0.00898f
C2136 SD3_1.n19 VSS 0.018f
C2137 SD3_1.n20 VSS 0.0161f
C2138 SD3_1.t49 VSS 0.00898f
C2139 SD3_1.n21 VSS 0.00898f
C2140 SD3_1.n22 VSS 0.0342f
C2141 SD3_1.t16 VSS 0.00898f
C2142 SD3_1.n23 VSS 0.00898f
C2143 SD3_1.n24 VSS 0.018f
C2144 SD3_1.n25 VSS 0.0222f
C2145 SD3_1.t15 VSS 0.00898f
C2146 SD3_1.n26 VSS 0.00898f
C2147 SD3_1.n27 VSS 0.0342f
C2148 SD3_1.t31 VSS 0.00898f
C2149 SD3_1.n28 VSS 0.00898f
C2150 SD3_1.n29 VSS 0.018f
C2151 SD3_1.n30 VSS 0.0222f
C2152 SD3_1.t59 VSS 0.00898f
C2153 SD3_1.n31 VSS 0.00898f
C2154 SD3_1.n32 VSS 0.034f
C2155 SD3_1.t22 VSS 0.00898f
C2156 SD3_1.n33 VSS 0.00898f
C2157 SD3_1.n34 VSS 0.018f
C2158 SD3_1.n35 VSS 0.0161f
C2159 SD3_1.t26 VSS 0.00898f
C2160 SD3_1.n36 VSS 0.00898f
C2161 SD3_1.n37 VSS 0.0377f
C2162 SD3_1.t40 VSS 0.00898f
C2163 SD3_1.n38 VSS 0.00898f
C2164 SD3_1.n39 VSS 0.0181f
C2165 SD3_1.n40 VSS 0.0229f
C2166 SD3_1.t47 VSS 0.00898f
C2167 SD3_1.n41 VSS 0.00898f
C2168 SD3_1.n42 VSS 0.0375f
C2169 SD3_1.t62 VSS 0.00898f
C2170 SD3_1.n43 VSS 0.00898f
C2171 SD3_1.n44 VSS 0.0373f
C2172 SD3_1.t35 VSS 0.00898f
C2173 SD3_1.n45 VSS 0.00898f
C2174 SD3_1.n46 VSS 0.018f
C2175 SD3_1.n47 VSS 0.0222f
C2176 SD3_1.t55 VSS 0.00898f
C2177 SD3_1.n48 VSS 0.00898f
C2178 SD3_1.n49 VSS 0.034f
C2179 SD3_1.t13 VSS 0.00898f
C2180 SD3_1.n50 VSS 0.00898f
C2181 SD3_1.n51 VSS 0.0374f
C2182 SD3_1.t17 VSS 0.00898f
C2183 SD3_1.n52 VSS 0.00898f
C2184 SD3_1.n53 VSS 0.0251f
C2185 SD3_1.t44 VSS 0.00898f
C2186 SD3_1.n54 VSS 0.00898f
C2187 SD3_1.n55 VSS 0.0343f
C2188 SD3_1.n56 VSS 0.125f
C2189 SD3_1.n57 VSS 0.0341f
C2190 SD3_1.n58 VSS 0.0788f
C2191 SD3_1.t30 VSS 0.00898f
C2192 SD3_1.n59 VSS 0.00898f
C2193 SD3_1.n60 VSS 0.018f
C2194 SD3_1.n61 VSS 0.0161f
C2195 SD3_1.n62 VSS 0.0333f
C2196 SD3_1.n63 VSS 0.0332f
C2197 SD3_1.n64 VSS 0.0762f
C2198 SD3_1.t0 VSS 0.00898f
C2199 SD3_1.n65 VSS 0.00898f
C2200 SD3_1.n66 VSS 0.018f
C2201 SD3_1.n67 VSS 0.0161f
C2202 SD3_1.n68 VSS 0.0338f
C2203 SD3_1.n69 VSS 0.0336f
C2204 SD3_1.n70 VSS 0.0792f
C2205 SD3_1.n71 VSS 0.0337f
C2206 SD3_1.t11 VSS 0.00898f
C2207 SD3_1.n72 VSS 0.00898f
C2208 SD3_1.n73 VSS 0.0181f
C2209 SD3_1.n74 VSS 0.0229f
C2210 SD3_1.n75 VSS 0.0339f
C2211 SD3_1.n76 VSS 0.0792f
C2212 SD3_1.n77 VSS 0.0333f
C2213 SD3_1.n78 VSS 0.0335f
C2214 SD3_1.n79 VSS 0.0793f
C2215 SD3_1.n80 VSS 0.0337f
C2216 SD3_1.n81 VSS 0.034f
C2217 SD3_1.n82 VSS 0.0758f
C2218 SD3_1.n83 VSS 0.0332f
C2219 SD3_1.n84 VSS 0.0338f
C2220 SD3_1.n85 VSS 0.0765f
C2221 SD3_1.n86 VSS 0.0333f
C2222 SD3_1.n87 VSS 0.0343f
C2223 SD3_1.n88 VSS 0.0762f
C2224 SD3_1.n89 VSS 0.033f
C2225 SD3_1.n90 VSS 0.033f
C2226 SD3_1.n91 VSS 0.079f
C2227 SD3_1.n92 VSS 0.034f
C2228 SD3_1.n93 VSS 0.0337f
C2229 SD3_1.n94 VSS 0.0733f
C2230 SD3_1.n95 VSS 0.0335f
C2231 SD3_1.n96 VSS 0.0332f
C2232 SD3_1.n97 VSS 0.0764f
C2233 SD3_1.n98 VSS 0.0342f
C2234 SD3_1.n99 VSS 0.0346f
C2235 SD3_1.n100 VSS 0.0761f
C2236 SD3_1.n101 VSS 0.00975f
C2237 SD3_1.t7 VSS 0.0083f
C2238 SD3_1.n102 VSS 0.0179f
C2239 SD3_1.n103 VSS 0.0161f
C2240 SD3_1.n104 VSS 0.0341f
C2241 SD3_1.t42 VSS 0.00898f
C2242 SD3_1.n105 VSS 0.00898f
C2243 SD3_1.n106 VSS 0.018f
C2244 SD3_1.n107 VSS 0.0161f
C2245 SD3_1.n108 VSS 0.0354f
C2246 SD3_1.n109 VSS 0.0739f
C2247 SD3_1.n110 VSS 0.0336f
C2248 SD3_1.t8 VSS 0.00898f
C2249 SD3_1.n111 VSS 0.00898f
C2250 SD3_1.n112 VSS 0.018f
C2251 SD3_1.n113 VSS 0.00381f
C2252 SD3_1.n114 VSS 0.0166f
C2253 SD3_1.n115 VSS 0.0329f
C2254 SD3_1.t3 VSS 0.00898f
C2255 SD3_1.n116 VSS 0.00898f
C2256 SD3_1.n117 VSS 0.0375f
C2257 SD3_1.t51 VSS 0.00898f
C2258 SD3_1.n118 VSS 0.00898f
C2259 SD3_1.n119 VSS 0.0251f
C2260 SD3_1.n120 VSS 0.126f
C2261 SD3_1.n121 VSS 0.034f
C2262 SDn_2.t20 VSS 0.00634f
C2263 SDn_2.n0 VSS 0.00634f
C2264 SDn_2.n1 VSS 0.0186f
C2265 SDn_2.n2 VSS 0.00621f
C2266 SDn_2.t52 VSS 0.039f
C2267 SDn_2.t67 VSS 0.0238f
C2268 SDn_2.n3 VSS 0.0426f
C2269 SDn_2.t75 VSS 0.0238f
C2270 SDn_2.n4 VSS 0.0318f
C2271 SDn_2.t68 VSS 0.0228f
C2272 SDn_2.n5 VSS 0.0308f
C2273 SDn_2.t35 VSS 0.0228f
C2274 SDn_2.n6 VSS 0.0308f
C2275 SDn_2.t38 VSS 0.0238f
C2276 SDn_2.n7 VSS 0.0318f
C2277 SDn_2.t70 VSS 0.0238f
C2278 SDn_2.n8 VSS 0.0318f
C2279 SDn_2.t36 VSS 0.0228f
C2280 SDn_2.n9 VSS 0.0308f
C2281 SDn_2.t49 VSS 0.0228f
C2282 SDn_2.n10 VSS 0.0308f
C2283 SDn_2.t71 VSS 0.0238f
C2284 SDn_2.n11 VSS 0.0318f
C2285 SDn_2.t61 VSS 0.0238f
C2286 SDn_2.n12 VSS 0.0318f
C2287 SDn_2.t44 VSS 0.0228f
C2288 SDn_2.n13 VSS 0.0308f
C2289 SDn_2.t27 VSS 0.0228f
C2290 SDn_2.n14 VSS 0.0308f
C2291 SDn_2.t48 VSS 0.0238f
C2292 SDn_2.n15 VSS 0.0318f
C2293 SDn_2.t74 VSS 0.0238f
C2294 SDn_2.n16 VSS 0.0318f
C2295 SDn_2.t72 VSS 0.0228f
C2296 SDn_2.n17 VSS 0.0308f
C2297 SDn_2.t46 VSS 0.0228f
C2298 SDn_2.n18 VSS 0.0308f
C2299 SDn_2.t73 VSS 0.0238f
C2300 SDn_2.n19 VSS 0.0318f
C2301 SDn_2.t64 VSS 0.0238f
C2302 SDn_2.n20 VSS 0.0318f
C2303 SDn_2.t50 VSS 0.0228f
C2304 SDn_2.n21 VSS 0.0308f
C2305 SDn_2.t29 VSS 0.0228f
C2306 SDn_2.n22 VSS 0.0308f
C2307 SDn_2.t51 VSS 0.0238f
C2308 SDn_2.n23 VSS 0.0318f
C2309 SDn_2.t30 VSS 0.0238f
C2310 SDn_2.n24 VSS 0.0318f
C2311 SDn_2.t34 VSS 0.0228f
C2312 SDn_2.n25 VSS 0.0308f
C2313 SDn_2.t65 VSS 0.0228f
C2314 SDn_2.n26 VSS 0.0308f
C2315 SDn_2.t24 VSS 0.0238f
C2316 SDn_2.n27 VSS 0.0318f
C2317 SDn_2.t56 VSS 0.0238f
C2318 SDn_2.n28 VSS 0.0318f
C2319 SDn_2.t53 VSS 0.0228f
C2320 SDn_2.n29 VSS 0.0308f
C2321 SDn_2.t41 VSS 0.0228f
C2322 SDn_2.n30 VSS 0.0308f
C2323 SDn_2.t59 VSS 0.0238f
C2324 SDn_2.n31 VSS 0.0318f
C2325 SDn_2.t43 VSS 0.0238f
C2326 SDn_2.n32 VSS 0.0318f
C2327 SDn_2.t25 VSS 0.0228f
C2328 SDn_2.n33 VSS 0.253f
C2329 SDn_2.t60 VSS 0.0212f
C2330 SDn_2.n34 VSS 0.171f
C2331 SDn_2.t69 VSS 0.0233f
C2332 SDn_2.n35 VSS 0.0313f
C2333 SDn_2.t40 VSS 0.0233f
C2334 SDn_2.n36 VSS 0.0313f
C2335 SDn_2.t37 VSS 0.0212f
C2336 SDn_2.n37 VSS 0.0292f
C2337 SDn_2.t31 VSS 0.0212f
C2338 SDn_2.n38 VSS 0.0292f
C2339 SDn_2.t33 VSS 0.0233f
C2340 SDn_2.n39 VSS 0.0313f
C2341 SDn_2.t54 VSS 0.0233f
C2342 SDn_2.n40 VSS 0.0313f
C2343 SDn_2.t28 VSS 0.0212f
C2344 SDn_2.n41 VSS 0.0342f
C2345 SDn_2.t14 VSS 0.0212f
C2346 SDn_2.n42 VSS 0.0342f
C2347 SDn_2.t0 VSS 0.0212f
C2348 SDn_2.n43 VSS 0.0291f
C2349 SDn_2.t10 VSS 0.0233f
C2350 SDn_2.n44 VSS 0.0313f
C2351 SDn_2.n45 VSS 0.0143f
C2352 SDn_2.t8 VSS 0.0184f
C2353 SDn_2.n47 VSS 0.0157f
C2354 SDn_2.n48 VSS 0.00861f
C2355 SDn_2.n49 VSS 0.00856f
C2356 SDn_2.n50 VSS 0.0645f
C2357 SDn_2.t1 VSS 0.00602f
C2358 SDn_2.n51 VSS 0.0067f
C2359 SDn_2.n52 VSS 0.0265f
C2360 SDn_2.t3 VSS 0.00586f
C2361 SDn_2.n53 VSS 0.00689f
C2362 SDn_2.n54 VSS 0.021f
C2363 SDn_2.n55 VSS 0.00683f
C2364 SDn_2.t7 VSS 0.00591f
C2365 SDn_2.n56 VSS 0.0241f
C2366 SDn_2.n57 VSS 0.00683f
C2367 SDn_2.t17 VSS 0.00591f
C2368 SDn_2.n58 VSS 0.0182f
C2369 SDn_2.n59 VSS 0.0756f
C2370 SDn_2.n60 VSS 0.00683f
C2371 SDn_2.t18 VSS 0.00591f
C2372 SDn_2.n61 VSS 0.0202f
C2373 SDn_2.t63 VSS 0.037f
C2374 SDn_2.t55 VSS 0.0233f
C2375 SDn_2.n62 VSS 0.0409f
C2376 SDn_2.t66 VSS 0.0233f
C2377 SDn_2.n63 VSS 0.0313f
C2378 SDn_2.t47 VSS 0.0212f
C2379 SDn_2.n64 VSS 0.0292f
C2380 SDn_2.t39 VSS 0.0212f
C2381 SDn_2.n65 VSS 0.0292f
C2382 SDn_2.t57 VSS 0.0233f
C2383 SDn_2.n66 VSS 0.0313f
C2384 SDn_2.t32 VSS 0.0233f
C2385 SDn_2.n67 VSS 0.0313f
C2386 SDn_2.t58 VSS 0.0212f
C2387 SDn_2.n68 VSS 0.034f
C2388 SDn_2.t6 VSS 0.0212f
C2389 SDn_2.n69 VSS 0.0338f
C2390 SDn_2.t12 VSS 0.0233f
C2391 SDn_2.n70 VSS 0.0313f
C2392 SDn_2.t4 VSS 0.0212f
C2393 SDn_2.n71 VSS 0.0291f
C2394 SDn_2.n72 VSS 0.0143f
C2395 SDn_2.t2 VSS 0.0184f
C2396 SDn_2.n74 VSS 0.0157f
C2397 SDn_2.n75 VSS 0.00842f
C2398 SDn_2.n76 VSS 0.00621f
C2399 SDn_2.n77 VSS 0.00877f
C2400 SDn_2.n78 VSS 0.0639f
C2401 SDn_2.n79 VSS 0.0297f
C2402 SDn_2.n80 VSS 0.0298f
C2403 SDn_2.n81 VSS 0.00689f
C2404 SDn_2.t16 VSS 0.00586f
C2405 SDn_2.n82 VSS 0.0126f
C2406 SDn_2.n83 VSS 0.00937f
C2407 SDn_2.n84 VSS 0.0254f
C2408 SDn_2.n85 VSS 0.0472f
C2409 SDn_2.n86 VSS 0.0224f
C2410 SDn_2.n87 VSS 0.0225f
C2411 SDn_2.n88 VSS 0.00636f
C2412 SDn_2.t9 VSS 0.00634f
C2413 SDn_2.n89 VSS 0.00634f
C2414 SDn_2.n90 VSS 0.0127f
C2415 SDn_2.n91 VSS 0.00567f
C2416 SDn_2.n92 VSS 0.0102f
C2417 SDn_2.n93 VSS 5.1e-19
C2418 VDD.n0 VSS 0.00271f
C2419 VDD.t78 VSS 0.00323f
C2420 VDD.t77 VSS 0.122f
C2421 VDD.t54 VSS 0.123f
C2422 VDD.n1 VSS 0.108f
C2423 VDD.n2 VSS 0.0853f
C2424 VDD.n3 VSS 0.0531f
C2425 VDD.t61 VSS 0.0984f
C2426 VDD.t62 VSS 0.00516f
C2427 VDD.t68 VSS 0.00516f
C2428 VDD.n4 VSS 0.00271f
C2429 VDD.t60 VSS 0.00323f
C2430 VDD.t59 VSS 0.122f
C2431 VDD.t0 VSS 0.123f
C2432 VDD.n5 VSS 0.108f
C2433 VDD.n6 VSS 0.0853f
C2434 VDD.n7 VSS 0.0544f
C2435 VDD.t67 VSS 0.0984f
C2436 VDD.n8 VSS 0.0545f
C2437 VDD.t41 VSS 0.00516f
C2438 VDD.n9 VSS 0.00271f
C2439 VDD.t14 VSS 0.00323f
C2440 VDD.t13 VSS 0.122f
C2441 VDD.t69 VSS 0.123f
C2442 VDD.n10 VSS 0.108f
C2443 VDD.n11 VSS 0.0853f
C2444 VDD.n12 VSS 0.0544f
C2445 VDD.t40 VSS 0.0984f
C2446 VDD.n13 VSS 0.0559f
C2447 VDD.t74 VSS 0.00516f
C2448 VDD.n14 VSS 0.00271f
C2449 VDD.t64 VSS 0.00271f
C2450 VDD.t66 VSS 0.00516f
C2451 VDD.n15 VSS 0.00271f
C2452 VDD.t53 VSS 0.00271f
C2453 VDD.t4 VSS 0.00516f
C2454 VDD.n16 VSS 0.00271f
C2455 VDD.t16 VSS 0.00323f
C2456 VDD.t15 VSS 0.122f
C2457 VDD.t95 VSS 0.123f
C2458 VDD.n17 VSS 0.108f
C2459 VDD.n18 VSS 0.0853f
C2460 VDD.n19 VSS 0.0544f
C2461 VDD.t3 VSS 0.0984f
C2462 VDD.n20 VSS 0.0426f
C2463 VDD.n21 VSS 0.0529f
C2464 VDD.t52 VSS 0.122f
C2465 VDD.t49 VSS 0.123f
C2466 VDD.n22 VSS 0.108f
C2467 VDD.n23 VSS 0.0339f
C2468 VDD.n24 VSS 0.0544f
C2469 VDD.t65 VSS 0.0984f
C2470 VDD.n25 VSS 0.0428f
C2471 VDD.n26 VSS 0.0532f
C2472 VDD.t63 VSS 0.122f
C2473 VDD.t83 VSS 0.123f
C2474 VDD.n27 VSS 0.108f
C2475 VDD.n28 VSS 0.0339f
C2476 VDD.n29 VSS 0.0544f
C2477 VDD.t73 VSS 0.0984f
C2478 VDD.n30 VSS 0.0666f
C2479 VDD.n31 VSS 0.107f
C2480 VDD.n32 VSS 0.0994f
C2481 VDD.n33 VSS 0.0124f
C2482 VDD.n34 VSS 0.0124f
C2483 VDD.n35 VSS 0.0147f
C2484 VDD.n36 VSS 0.00316f
C2485 VDD.t25 VSS 0.00293f
C2486 VDD.n37 VSS 0.00293f
C2487 VDD.n38 VSS 0.00701f
C2488 VDD.n39 VSS 0.00702f
C2489 VDD.n40 VSS 0.0296f
C2490 VDD.n41 VSS 0.0127f
C2491 VDD.t30 VSS 0.00702f
C2492 VDD.t39 VSS 0.00293f
C2493 VDD.n42 VSS 0.00293f
C2494 VDD.n43 VSS 0.00701f
C2495 VDD.n44 VSS 0.00711f
C2496 VDD.t26 VSS 0.0634f
C2497 VDD.n45 VSS 0.166f
C2498 VDD.t37 VSS 0.0582f
C2499 VDD.n46 VSS 0.0633f
C2500 VDD.n47 VSS 0.0391f
C2501 VDD.t79 VSS 0.0582f
C2502 VDD.n48 VSS 0.0633f
C2503 VDD.n49 VSS 0.0391f
C2504 VDD.t38 VSS 0.0582f
C2505 VDD.n50 VSS 0.0633f
C2506 VDD.n51 VSS 0.0353f
C2507 VDD.n52 VSS 0.0278f
C2508 VDD.t80 VSS 0.0582f
C2509 VDD.n53 VSS 0.0633f
C2510 VDD.n54 VSS 0.0268f
C2511 VDD.t57 VSS 0.0582f
C2512 VDD.n55 VSS 0.0633f
C2513 VDD.n56 VSS 0.0391f
C2514 VDD.t91 VSS 0.0582f
C2515 VDD.n57 VSS 0.0633f
C2516 VDD.n58 VSS 0.0391f
C2517 VDD.t29 VSS 0.0582f
C2518 VDD.n59 VSS 0.0633f
C2519 VDD.n60 VSS 0.0334f
C2520 VDD.n61 VSS 0.0318f
C2521 VDD.n62 VSS 0.122f
C2522 VDD.n63 VSS 0.0226f
C2523 VDD.n64 VSS 0.0171f
C2524 VDD.n65 VSS 0.0435f
C2525 VDD.t92 VSS 0.076f
C2526 VDD.n66 VSS 0.0633f
C2527 VDD.n67 VSS 0.034f
C2528 VDD.t48 VSS 0.0582f
C2529 VDD.n68 VSS 0.0633f
C2530 VDD.n69 VSS 0.0391f
C2531 VDD.t72 VSS 0.0582f
C2532 VDD.n70 VSS 0.0633f
C2533 VDD.n71 VSS 0.0382f
C2534 VDD.n72 VSS 0.0162f
C2535 VDD.n73 VSS 0.00445f
C2536 VDD.n74 VSS 0.0422f
C2537 VDD.t7 VSS 0.0549f
C2538 VDD.n75 VSS 0.0144f
C2539 VDD.n76 VSS 0.00354f
C2540 VDD.n77 VSS 0.0128f
C2541 VDD.n78 VSS 0.00441f
C2542 VDD.n79 VSS 0.00396f
C2543 VDD.n80 VSS 0.00421f
C2544 VDD.n81 VSS 0.00316f
C2545 VDD.t8 VSS 0.0027f
C2546 VDD.n82 VSS 0.0195f
C2547 VDD.n83 VSS 0.0289f
C2548 VDD.t31 VSS 0.0494f
C2549 VDD.n84 VSS 0.0633f
C2550 VDD.n85 VSS 0.0358f
C2551 VDD.t9 VSS 0.0582f
C2552 VDD.n86 VSS 0.0633f
C2553 VDD.n87 VSS 0.0391f
C2554 VDD.t17 VSS 0.0582f
C2555 VDD.n88 VSS 0.0633f
C2556 VDD.n89 VSS 0.0378f
C2557 VDD.n90 VSS 0.0162f
C2558 VDD.n91 VSS 0.00346f
C2559 VDD.n92 VSS 0.0355f
C2560 VDD.t45 VSS 0.0533f
C2561 VDD.n93 VSS 0.0211f
C2562 VDD.n94 VSS 0.0031f
C2563 VDD.n95 VSS 0.0127f
C2564 VDD.n96 VSS 0.00593f
C2565 VDD.n97 VSS 0.00391f
C2566 VDD.n98 VSS 0.00369f
C2567 VDD.n99 VSS 0.00319f
C2568 VDD.t46 VSS 0.00268f
C2569 VDD.n100 VSS 0.0198f
C2570 VDD.n101 VSS 0.0297f
C2571 VDD.t10 VSS 0.051f
C2572 VDD.n102 VSS 0.0633f
C2573 VDD.n103 VSS 0.0364f
C2574 VDD.t18 VSS 0.0582f
C2575 VDD.n104 VSS 0.0633f
C2576 VDD.n105 VSS 0.0391f
C2577 VDD.t34 VSS 0.0582f
C2578 VDD.n106 VSS 0.0633f
C2579 VDD.n107 VSS 0.0365f
C2580 VDD.n108 VSS 0.0162f
C2581 VDD.n109 VSS 0.0152f
C2582 VDD.n110 VSS 0.00467f
C2583 VDD.n111 VSS 0.0034f
C2584 VDD.n112 VSS 0.00314f
C2585 VDD.t6 VSS 0.00272f
C2586 VDD.n113 VSS 0.0235f
C2587 VDD.n114 VSS 0.0167f
C2588 VDD.t5 VSS 0.0488f
C2589 VDD.n115 VSS 0.0277f
C2590 VDD.n116 VSS 0.0044f
C2591 VDD.t42 VSS 0.0492f
C2592 VDD.n117 VSS 0.0326f
C2593 VDD.n118 VSS 0.00336f
C2594 VDD.n119 VSS 0.0143f
C2595 VDD.t47 VSS 0.0582f
C2596 VDD.n120 VSS 0.0633f
C2597 VDD.n121 VSS 0.038f
C2598 VDD.t35 VSS 0.0582f
C2599 VDD.n122 VSS 0.0633f
C2600 VDD.n123 VSS 0.0391f
C2601 VDD.t75 VSS 0.0508f
C2602 VDD.n124 VSS 0.0633f
C2603 VDD.n125 VSS 0.0363f
C2604 VDD.t76 VSS 0.0155f
C2605 VDD.n126 VSS 0.0391f
C2606 VDD.n127 VSS 0.0037f
C2607 VDD.n128 VSS 0.00308f
C2608 VDD.n129 VSS 0.00393f
C2609 VDD.n130 VSS 0.00496f
C2610 VDD.n131 VSS 0.00423f
C2611 VDD.n132 VSS 0.0344f
C2612 VDD.n133 VSS 0.00325f
C2613 VDD.n134 VSS 0.0613f
C2614 VDD.t21 VSS 0.0582f
C2615 VDD.n135 VSS 0.0897f
C2616 VDD.n136 VSS 0.0235f
C2617 VDD.t36 VSS 0.0582f
C2618 VDD.n137 VSS 0.0633f
C2619 VDD.n138 VSS 0.0391f
C2620 VDD.t19 VSS 0.0582f
C2621 VDD.n139 VSS 0.0633f
C2622 VDD.n140 VSS 0.0391f
C2623 VDD.t24 VSS 0.0571f
C2624 VDD.n141 VSS 0.0633f
C2625 VDD.n142 VSS 0.0349f
C2626 VDD.n143 VSS 0.0138f
C2627 VDD.n144 VSS 0.0147f
C2628 VDD.n145 VSS 0.00208f
C2629 VDD.n146 VSS 0.00116f
C2630 VDD.n147 VSS 0.0128f
C2631 VDD.n148 VSS 0.0369f
C2632 VDD.t88 VSS 0.0472f
C2633 VDD.n149 VSS 0.0197f
C2634 VDD.n150 VSS 0.00842f
C2635 VDD.n151 VSS 0.0039f
C2636 VDD.n152 VSS 0.00399f
C2637 VDD.n153 VSS 0.0127f
C2638 VDD.n154 VSS 0.0131f
C2639 VDD.t20 VSS 0.0582f
C2640 VDD.n155 VSS 0.0633f
C2641 VDD.n156 VSS 0.0137f
C2642 VDD.t58 VSS 0.0582f
C2643 VDD.n157 VSS 0.0633f
C2644 VDD.t86 VSS 0.139f
C2645 VDD.n158 VSS 0.0633f
C2646 VDD.t87 VSS 0.00766f
C2647 VDD.n159 VSS 0.0806f
C2648 VDD.n160 VSS 0.0382f
C2649 VDD.n161 VSS 0.0137f
C2650 VDD.n162 VSS 0.0103f
C2651 VDD.n163 VSS 0.436f
C2652 VDD.n164 VSS 0.419f
C2653 VDD.n165 VSS 0.0381f
C2654 OUT+.t75 VSS 0.0202f
C2655 OUT+.n0 VSS 0.0333f
C2656 OUT+.t74 VSS 0.0243f
C2657 OUT+.t46 VSS 0.0428f
C2658 OUT+.n1 VSS 0.0687f
C2659 OUT+.n2 VSS 0.134f
C2660 OUT+.t59 VSS 0.0568f
C2661 OUT+.t58 VSS 0.0666f
C2662 OUT+.n3 VSS 0.177f
C2663 OUT+.t120 VSS 0.0288f
C2664 OUT+.n4 VSS 0.149f
C2665 OUT+.n5 VSS 0.0853f
C2666 OUT+.t47 VSS 0.0167f
C2667 OUT+.t123 VSS 0.0202f
C2668 OUT+.n6 VSS 0.0159f
C2669 OUT+.n7 VSS 0.0364f
C2670 OUT+.n8 VSS 0.0629f
C2671 OUT+.t108 VSS 0.0573f
C2672 OUT+.n9 VSS 0.109f
C2673 OUT+.t15 VSS 0.0227f
C2674 OUT+.t14 VSS 0.0278f
C2675 OUT+.n10 VSS 0.092f
C2676 OUT+.t109 VSS 0.0403f
C2677 OUT+.n11 VSS 0.0121f
C2678 OUT+.n12 VSS 0.0242f
C2679 OUT+.n13 VSS 0.157f
C2680 OUT+.n14 VSS 0.0358f
C2681 OUT+.t128 VSS 0.0121f
C2682 OUT+.t41 VSS 0.0242f
C2683 OUT+.n15 VSS 0.025f
C2684 OUT+.t73 VSS 0.0437f
C2685 OUT+.n16 VSS 0.0254f
C2686 OUT+.t40 VSS 0.0505f
C2687 OUT+.t72 VSS 0.0434f
C2688 OUT+.n17 VSS 0.0705f
C2689 OUT+.n18 VSS 0.086f
C2690 OUT+.n19 VSS 0.0568f
C2691 OUT+.n20 VSS 0.102f
C2692 OUT+.n21 VSS 0.211f
C2693 OUT+.t171 VSS 0.0207f
C2694 OUT+.t188 VSS 0.0207f
C2695 OUT+.n22 VSS 0.0166f
C2696 OUT+.t4 VSS 0.0207f
C2697 OUT+.n23 VSS 0.0166f
C2698 OUT+.n24 VSS 0.103f
C2699 OUT+.n25 VSS 0.098f
C2700 OUT+.n26 VSS 0.0782f
C2701 OUT+.t175 VSS 0.0202f
C2702 OUT+.n27 VSS 0.0711f
C2703 OUT+.n28 VSS 0.0276f
C2704 OUT+.n29 VSS 0.0726f
C2705 OUT+.n30 VSS 0.0276f
C2706 OUT+.t155 VSS 0.027f
C2707 OUT+.n31 VSS 0.0148f
C2708 OUT+.n32 VSS 0.00522f
C2709 OUT+.t99 VSS 0.0405f
C2710 OUT+.t20 VSS 0.0397f
C2711 OUT+.n33 VSS 0.025f
C2712 OUT+.t191 VSS 0.0397f
C2713 OUT+.t122 VSS 0.0397f
C2714 OUT+.t177 VSS 0.0397f
C2715 OUT+.t57 VSS 0.0418f
C2716 OUT+.n34 VSS 0.0252f
C2717 OUT+.t56 VSS 0.044f
C2718 OUT+.n35 VSS 0.121f
C2719 OUT+.n36 VSS 0.0685f
C2720 OUT+.n37 VSS 0.0897f
C2721 OUT+.n38 VSS 0.0756f
C2722 OUT+.t19 VSS 0.0407f
C2723 OUT+.n39 VSS 0.0256f
C2724 OUT+.t178 VSS 0.0408f
C2725 OUT+.n40 VSS 0.0258f
C2726 OUT+.n41 VSS 0.0976f
C2727 OUT+.t24 VSS 0.0411f
C2728 OUT+.t166 VSS 0.0397f
C2729 OUT+.n42 VSS 0.0258f
C2730 OUT+.t10 VSS 0.0397f
C2731 OUT+.n43 VSS 0.0256f
C2732 OUT+.t67 VSS 0.0418f
C2733 OUT+.n44 VSS 0.0251f
C2734 OUT+.t66 VSS 0.0445f
C2735 OUT+.n45 VSS 0.118f
C2736 OUT+.n46 VSS 0.0616f
C2737 OUT+.t23 VSS 0.0456f
C2738 OUT+.t11 VSS 0.0567f
C2739 OUT+.n47 VSS 0.17f
C2740 OUT+.n48 VSS 0.215f
C2741 OUT+.t176 VSS 0.0397f
C2742 OUT+.n49 VSS 0.075f
C2743 OUT+.n50 VSS 0.0762f
C2744 OUT+.t150 VSS 0.0397f
C2745 OUT+.t21 VSS 0.0555f
C2746 OUT+.t145 VSS 0.0457f
C2747 OUT+.n51 VSS 0.168f
C2748 OUT+.t112 VSS 0.045f
C2749 OUT+.n52 VSS 0.123f
C2750 OUT+.t113 VSS 0.0423f
C2751 OUT+.n53 VSS 0.0251f
C2752 OUT+.n54 VSS 0.0564f
C2753 OUT+.t38 VSS 0.0341f
C2754 OUT+.t90 VSS 0.0355f
C2755 OUT+.n55 VSS 0.0572f
C2756 OUT+.t95 VSS 0.0408f
C2757 OUT+.n56 VSS 0.0255f
C2758 OUT+.t61 VSS 0.0409f
C2759 OUT+.n57 VSS 0.0255f
C2760 OUT+.n58 VSS 0.112f
C2761 OUT+.t94 VSS 0.0335f
C2762 OUT+.t60 VSS 0.0361f
C2763 OUT+.n59 VSS 0.0572f
C2764 OUT+.n60 VSS 0.0257f
C2765 OUT+.n61 VSS 0.0925f
C2766 OUT+.n62 VSS 0.0159f
C2767 OUT+.t39 VSS 0.0408f
C2768 OUT+.t91 VSS 0.0408f
C2769 OUT+.t80 VSS 0.0316f
C2770 OUT+.t42 VSS 0.038f
C2771 OUT+.n63 VSS 0.0572f
C2772 OUT+.t3 VSS 0.0121f
C2773 OUT+.n64 VSS 0.0121f
C2774 OUT+.n65 VSS 0.0242f
C2775 OUT+.t22 VSS 0.0121f
C2776 OUT+.n66 VSS 0.0121f
C2777 OUT+.n67 VSS 0.0305f
C2778 OUT+.n68 VSS 0.0996f
C2779 OUT+.t170 VSS 0.0121f
C2780 OUT+.n69 VSS 0.0121f
C2781 OUT+.n70 VSS 0.0262f
C2782 OUT+.t169 VSS 0.0121f
C2783 OUT+.t49 VSS 0.0407f
C2784 OUT+.n71 VSS 0.0242f
C2785 OUT+.t189 VSS 0.0121f
C2786 OUT+.t105 VSS 0.0409f
C2787 OUT+.n72 VSS 0.0242f
C2788 OUT+.t12 VSS 0.0121f
C2789 OUT+.n73 VSS 0.0121f
C2790 OUT+.n74 VSS 0.0242f
C2791 OUT+.t106 VSS 0.0326f
C2792 OUT+.t82 VSS 0.0371f
C2793 OUT+.n75 VSS 0.0568f
C2794 OUT+.n76 VSS 0.117f
C2795 OUT+.n77 VSS 0.0223f
C2796 OUT+.t1 VSS 0.0121f
C2797 OUT+.t107 VSS 0.0407f
C2798 OUT+.n78 VSS 0.0259f
C2799 OUT+.n79 VSS 0.0503f
C2800 OUT+.t6 VSS 0.0121f
C2801 OUT+.t83 VSS 0.041f
C2802 OUT+.n80 VSS 0.0242f
C2803 OUT+.t0 VSS 0.0121f
C2804 OUT+.n81 VSS 0.0121f
C2805 OUT+.n82 VSS 0.0254f
C2806 OUT+.t174 VSS 0.0121f
C2807 OUT+.n83 VSS 0.0121f
C2808 OUT+.n84 VSS 0.0302f
C2809 OUT+.t26 VSS 0.0121f
C2810 OUT+.n85 VSS 0.0121f
C2811 OUT+.n86 VSS 0.0242f
C2812 OUT+.n87 VSS 0.104f
C2813 OUT+.t45 VSS 0.0407f
C2814 OUT+.n88 VSS 0.0121f
C2815 OUT+.n89 VSS 0.0255f
C2816 OUT+.t63 VSS 0.0406f
C2817 OUT+.n90 VSS 0.0253f
C2818 OUT+.t35 VSS 0.0409f
C2819 OUT+.n91 VSS 0.0256f
C2820 OUT+.n92 VSS 0.114f
C2821 OUT+.t62 VSS 0.0324f
C2822 OUT+.t34 VSS 0.0372f
C2823 OUT+.n93 VSS 0.0572f
C2824 OUT+.n94 VSS 0.0279f
C2825 OUT+.n95 VSS 0.0936f
C2826 OUT+.t92 VSS 0.0322f
C2827 OUT+.t70 VSS 0.0374f
C2828 OUT+.n96 VSS 0.0572f
C2829 OUT+.n97 VSS 0.024f
C2830 OUT+.t93 VSS 0.0411f
C2831 OUT+.n98 VSS 0.0624f
C2832 OUT+.t71 VSS 0.0413f
C2833 OUT+.n99 VSS 0.0671f
C2834 OUT+.n100 VSS 0.119f
C2835 OUT+.t44 VSS 0.0332f
C2836 OUT+.t102 VSS 0.0364f
C2837 OUT+.n101 VSS 0.0572f
C2838 OUT+.n102 VSS 0.0255f
C2839 OUT+.n103 VSS 0.0662f
C2840 OUT+.t103 VSS 0.0409f
C2841 OUT+.n104 VSS 0.0121f
C2842 OUT+.n105 VSS 0.0242f
C2843 OUT+.n106 VSS 0.0762f
C2844 OUT+.t2 VSS 0.0121f
C2845 OUT+.n107 VSS 0.0121f
C2846 OUT+.n108 VSS 0.026f
C2847 OUT+.n109 VSS 0.128f
C2848 OUT+.n110 VSS 0.214f
C2849 OUT+.n111 VSS 0.127f
C2850 OUT+.n112 VSS 0.0812f
C2851 OUT+.n113 VSS 0.148f
C2852 OUT+.t121 VSS 0.0121f
C2853 OUT+.n114 VSS 0.0121f
C2854 OUT+.n115 VSS 0.0265f
C2855 OUT+.n116 VSS 0.198f
C2856 OUT+.n117 VSS 0.0961f
C2857 OUT+.n118 VSS 0.0911f
C2858 OUT+.t48 VSS 0.0341f
C2859 OUT+.t104 VSS 0.0355f
C2860 OUT+.n119 VSS 0.0572f
C2861 OUT+.n120 VSS 0.113f
C2862 OUT+.n121 VSS 0.0268f
C2863 OUT+.n122 VSS 0.0433f
C2864 OUT+.n123 VSS 0.0717f
C2865 OUT+.n124 VSS 0.127f
C2866 OUT+.n125 VSS 0.214f
C2867 OUT+.t157 VSS 0.0121f
C2868 OUT+.n126 VSS 0.0121f
C2869 OUT+.n127 VSS 0.0263f
C2870 OUT+.n128 VSS 0.126f
C2871 OUT+.n129 VSS 0.0121f
C2872 OUT+.n130 VSS 0.0242f
C2873 OUT+.n131 VSS 0.0699f
C2874 OUT+.n132 VSS 0.0121f
C2875 OUT+.n133 VSS 0.0242f
C2876 OUT+.t186 VSS 0.0121f
C2877 OUT+.n134 VSS 0.0121f
C2878 OUT+.n135 VSS 0.0242f
C2879 OUT+.t168 VSS 0.0121f
C2880 OUT+.n136 VSS 0.0121f
C2881 OUT+.n137 VSS 0.0308f
C2882 OUT+.n138 VSS 0.151f
C2883 OUT+.n139 VSS 0.092f
C2884 OUT+.n140 VSS 0.0438f
C2885 OUT+.n141 VSS 0.0241f
C2886 OUT+.t81 VSS 0.0411f
C2887 OUT+.n142 VSS 0.0629f
C2888 OUT+.t43 VSS 0.0412f
C2889 OUT+.n143 VSS 0.0656f
C2890 OUT+.n144 VSS 0.118f
C2891 OUT+.n145 VSS 0.181f
C2892 OUT+.n146 VSS 0.118f
C2893 OUT+.n147 VSS 0.215f
C2894 OUT+.n148 VSS 0.0723f
C2895 OUT+.n149 VSS 0.073f
C2896 OUT+.n150 VSS 0.0469f
C2897 OUT+.n151 VSS 0.0999f
C2898 OUT+.t127 VSS 0.0411f
C2899 OUT+.n152 VSS 0.0682f
C2900 OUT+.n153 VSS 0.145f
C2901 OUT+.n154 VSS 0.115f
C2902 OUT+.n155 VSS 0.101f
C2903 OUT+.n156 VSS 0.047f
C2904 OUT+.n157 VSS 0.077f
C2905 OUT+.n158 VSS 0.0957f
C2906 OUT+.n159 VSS 0.0664f
C2907 OUT+.t98 VSS 0.0467f
C2908 OUT+.n160 VSS 0.0609f
C2909 OUT+.n161 VSS 0.0851f
C2910 OUT+.t147 VSS 0.0397f
C2911 OUT+.t161 VSS 0.0403f
C2912 OUT+.t167 VSS 0.0397f
C2913 OUT+.n162 VSS 0.025f
C2914 OUT+.t148 VSS 0.0403f
C2915 OUT+.n163 VSS 0.025f
C2916 OUT+.t152 VSS 0.0397f
C2917 OUT+.t146 VSS 0.0341f
C2918 OUT+.t131 VSS 0.0121f
C2919 OUT+.n164 VSS 0.0121f
C2920 OUT+.n165 VSS 0.0547f
C2921 OUT+.t132 VSS 0.0121f
C2922 OUT+.n166 VSS 0.0121f
C2923 OUT+.n167 VSS 0.0271f
C2924 OUT+.n168 VSS 0.286f
C2925 OUT+.t138 VSS 0.0121f
C2926 OUT+.n169 VSS 0.0121f
C2927 OUT+.n170 VSS 0.0356f
C2928 OUT+.t143 VSS 0.0121f
C2929 OUT+.n171 VSS 0.0121f
C2930 OUT+.n172 VSS 0.0348f
C2931 OUT+.t129 VSS 0.0121f
C2932 OUT+.n173 VSS 0.0121f
C2933 OUT+.n174 VSS 0.0259f
C2934 OUT+.t142 VSS 0.0121f
C2935 OUT+.n175 VSS 0.0121f
C2936 OUT+.n176 VSS 0.0259f
C2937 OUT+.n177 VSS 0.136f
C2938 OUT+.t77 VSS 0.0408f
C2939 OUT+.t69 VSS 0.0409f
C2940 OUT+.n178 VSS 0.106f
C2941 OUT+.t36 VSS 0.0335f
C2942 OUT+.t28 VSS 0.0361f
C2943 OUT+.n179 VSS 0.0572f
C2944 OUT+.n180 VSS 0.0237f
C2945 OUT+.t37 VSS 0.0408f
C2946 OUT+.n181 VSS 0.0261f
C2947 OUT+.n182 VSS 0.0452f
C2948 OUT+.t29 VSS 0.0409f
C2949 OUT+.n183 VSS 0.0262f
C2950 OUT+.n184 VSS 0.0463f
C2951 OUT+.t76 VSS 0.0341f
C2952 OUT+.t68 VSS 0.0355f
C2953 OUT+.n185 VSS 0.0572f
C2954 OUT+.n186 VSS 0.0232f
C2955 OUT+.n187 VSS 0.114f
C2956 OUT+.n188 VSS 0.0638f
C2957 OUT+.n189 VSS 0.058f
C2958 OUT+.t96 VSS 0.0322f
C2959 OUT+.t86 VSS 0.0374f
C2960 OUT+.n190 VSS 0.0572f
C2961 OUT+.n191 VSS 0.0229f
C2962 OUT+.t87 VSS 0.0414f
C2963 OUT+.n192 VSS 0.0121f
C2964 OUT+.n193 VSS 0.0258f
C2965 OUT+.n194 VSS 0.0604f
C2966 OUT+.t97 VSS 0.0412f
C2967 OUT+.n195 VSS 0.0121f
C2968 OUT+.n196 VSS 0.0242f
C2969 OUT+.n197 VSS 0.0617f
C2970 OUT+.n198 VSS 0.315f
C2971 OUT+.n199 VSS 0.137f
C2972 OUT+.n200 VSS 0.134f
C2973 OUT+.t140 VSS 0.0121f
C2974 OUT+.t33 VSS 0.0407f
C2975 OUT+.n201 VSS 0.0242f
C2976 OUT+.t139 VSS 0.0121f
C2977 OUT+.t115 VSS 0.041f
C2978 OUT+.n202 VSS 0.0256f
C2979 OUT+.t32 VSS 0.0328f
C2980 OUT+.t114 VSS 0.0368f
C2981 OUT+.n203 VSS 0.0572f
C2982 OUT+.n204 VSS 0.108f
C2983 OUT+.n205 VSS 0.0274f
C2984 OUT+.n206 VSS 0.0598f
C2985 OUT+.n207 VSS 0.0704f
C2986 OUT+.n208 VSS 0.47f
C2987 OUT+.n209 VSS 0.087f
C2988 OUT+.t65 VSS 0.0405f
C2989 OUT+.n210 VSS 0.0252f
C2990 OUT+.t101 VSS 0.0409f
C2991 OUT+.n211 VSS 0.0256f
C2992 OUT+.t64 VSS 0.0308f
C2993 OUT+.t100 VSS 0.0366f
C2994 OUT+.n212 VSS 0.0551f
C2995 OUT+.n213 VSS 0.117f
C2996 OUT+.n214 VSS 0.0306f
C2997 OUT+.n215 VSS 0.106f
C2998 OUT+.n216 VSS 0.0513f
C2999 OUT+.n217 VSS 0.13f
C3000 OUT+.n218 VSS 0.138f
C3001 OUT+.n219 VSS 0.0948f
C3002 OUT+.n220 VSS 0.105f
C3003 OUT+.n221 VSS 0.0951f
C3004 OUT+.n222 VSS 0.118f
C3005 OUT+.t151 VSS 0.0397f
C3006 OUT+.t149 VSS 0.041f
C3007 OUT+.t79 VSS 0.0406f
C3008 OUT+.n223 VSS 0.0253f
C3009 OUT+.t111 VSS 0.0408f
C3010 OUT+.n224 VSS 0.0255f
C3011 OUT+.n225 VSS 0.114f
C3012 OUT+.t78 VSS 0.033f
C3013 OUT+.t110 VSS 0.0345f
C3014 OUT+.n226 VSS 0.0551f
C3015 OUT+.n227 VSS 0.0304f
C3016 OUT+.n228 VSS 0.103f
C3017 OUT+.n229 VSS 0.0862f
C3018 OUT+.n230 VSS 0.0382f
C3019 OUT+.n231 VSS 0.261f
C3020 OUT+.n232 VSS 0.549f
C3021 OUT+.t9 VSS 0.0121f
C3022 OUT+.n233 VSS 0.0121f
C3023 OUT+.n234 VSS 0.0533f
C3024 OUT+.n235 VSS 0.318f
C3025 OUT+.t125 VSS 0.0121f
C3026 OUT+.t85 VSS 0.0397f
C3027 OUT+.n236 VSS 0.0242f
C3028 OUT+.t25 VSS 0.0121f
C3029 OUT+.t53 VSS 0.0451f
C3030 OUT+.n237 VSS 0.0283f
C3031 OUT+.t52 VSS 0.0603f
C3032 OUT+.t84 VSS 0.106f
C3033 OUT+.n238 VSS 0.108f
C3034 OUT+.n239 VSS 0.0825f
C3035 OUT+.n240 VSS 0.0647f
C3036 OUT+.n241 VSS 0.0554f
C3037 OUT+.t124 VSS 0.0121f
C3038 OUT+.n242 VSS 0.0121f
C3039 OUT+.n243 VSS 0.0498f
C3040 OUT+.n244 VSS 0.242f
C3041 OUT+.t119 VSS 0.0397f
C3042 OUT+.n245 VSS 0.0121f
C3043 OUT+.n246 VSS 0.0256f
C3044 OUT+.t89 VSS 0.0213f
C3045 OUT+.n247 VSS 0.0159f
C3046 OUT+.t88 VSS 0.0266f
C3047 OUT+.n248 VSS 0.108f
C3048 OUT+.n249 VSS 0.0391f
C3049 OUT+.t163 VSS 0.0207f
C3050 OUT+.n250 VSS 0.191f
C3051 OUT+.t158 VSS 0.0274f
C3052 OUT+.n251 VSS 0.241f
C3053 OUT+.n252 VSS 0.0734f
C3054 OUT+.n253 VSS 0.0702f
C3055 OUT+.t54 VSS 0.0314f
C3056 OUT+.t118 VSS 0.0351f
C3057 OUT+.n254 VSS 0.0541f
C3058 OUT+.n255 VSS 0.0268f
C3059 OUT+.n256 VSS 0.0615f
C3060 OUT+.t55 VSS 0.0406f
C3061 OUT+.n257 VSS 0.0121f
C3062 OUT+.n258 VSS 0.0242f
C3063 OUT+.n259 VSS 0.0102f
C3064 OUT+.n260 VSS 0.0162f
C3065 OUT+.n261 VSS 0.01f
C3066 OUT+.n262 VSS 0.0769f
C3067 OUT+.n263 VSS 0.0956f
C3068 OUT+.n264 VSS 0.0898f
C3069 OUT+.n265 VSS 0.0227f
C3070 OUT+.n266 VSS 0.00964f
C3071 OUT+.n267 VSS 0.0121f
C3072 OUT+.n268 VSS 0.119f
C3073 OUT+.t164 VSS 0.0202f
C3074 OUT+.t156 VSS 0.0207f
C3075 OUT+.n269 VSS 0.09f
C3076 OUT+.t159 VSS 0.0207f
C3077 OUT+.n270 VSS 0.0169f
C3078 OUT+.t162 VSS 0.0207f
C3079 OUT+.n271 VSS 0.0171f
C3080 OUT+.n272 VSS 0.0979f
C3081 OUT+.n273 VSS 0.068f
C3082 OUT+.n274 VSS 0.0647f
C3083 OUT+.n275 VSS 0.0606f
C3084 OUT+.t116 VSS 0.0323f
C3085 OUT+.n276 VSS 0.12f
C3086 OUT+.t117 VSS 0.0202f
C3087 OUT+.t160 VSS 0.0205f
C3088 OUT+.n277 VSS 0.0159f
C3089 OUT+.n278 VSS 0.0251f
C3090 OUT+.n279 VSS 0.00865f
C3091 OUT+.n280 VSS 0.0369f
C3092 OUT+.n281 VSS 5.95e-19
C3093 OUT+.n282 VSS 0.00798f
C3094 OUT+.n283 VSS 0.0211f
C3095 OUT+.n284 VSS 0.268f
C3096 OUT+.n285 VSS 0.105f
C3097 OUT+.n286 VSS 0.074f
C3098 OUT+.t16 VSS 0.0121f
C3099 OUT+.t51 VSS 0.0406f
C3100 OUT+.n287 VSS 0.0264f
C3101 OUT+.t179 VSS 0.0121f
C3102 OUT+.t31 VSS 0.041f
C3103 OUT+.n288 VSS 0.0273f
C3104 OUT+.n289 VSS 0.0844f
C3105 OUT+.t50 VSS 0.0324f
C3106 OUT+.t30 VSS 0.0386f
C3107 OUT+.n290 VSS 0.0586f
C3108 OUT+.n291 VSS 0.124f
C3109 OUT+.n292 VSS 0.0288f
C3110 OUT+.n293 VSS 0.014f
C3111 OUT+.n294 VSS 0.244f
C3112 OUT+.n295 VSS 0.263f
C3113 OUT+.n296 VSS 0.29f
.ends

