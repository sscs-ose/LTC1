magic
tech gf180mcuC
magscale 1 10
timestamp 1699939503
<< pwell >>
rect -503 -1107 2693 998
rect -503 -1110 2662 -1107
<< psubdiff >>
rect -453 868 2643 885
rect -453 822 -437 868
rect -391 822 -339 868
rect -293 822 -241 868
rect -195 822 -143 868
rect -97 822 -33 868
rect 13 822 65 868
rect 111 822 163 868
rect 209 822 261 868
rect 307 822 359 868
rect 405 822 457 868
rect 503 822 555 868
rect 601 822 653 868
rect 699 822 751 868
rect 797 822 849 868
rect 895 822 947 868
rect 993 822 1045 868
rect 1091 822 1143 868
rect 1189 822 1241 868
rect 1287 822 1339 868
rect 1385 822 1437 868
rect 1483 822 1535 868
rect 1581 822 1633 868
rect 1679 822 1731 868
rect 1777 822 1829 868
rect 1875 822 1927 868
rect 1973 822 2025 868
rect 2071 822 2123 868
rect 2169 822 2221 868
rect 2267 822 2319 868
rect 2365 822 2417 868
rect 2463 822 2580 868
rect 2626 822 2643 868
rect -453 805 2643 822
rect -453 770 -374 805
rect -453 724 -437 770
rect -391 724 -374 770
rect -453 672 -374 724
rect -453 626 -437 672
rect -391 626 -374 672
rect -453 574 -374 626
rect -453 528 -437 574
rect -391 528 -374 574
rect -453 476 -374 528
rect -453 430 -437 476
rect -391 430 -374 476
rect -453 378 -374 430
rect -453 332 -437 378
rect -391 332 -374 378
rect -453 280 -374 332
rect -453 234 -437 280
rect -391 234 -374 280
rect -453 182 -374 234
rect -453 136 -437 182
rect -391 136 -374 182
rect -453 84 -374 136
rect -453 38 -437 84
rect -391 38 -374 84
rect -453 -14 -374 38
rect 2563 770 2643 805
rect 2563 724 2580 770
rect 2626 724 2643 770
rect 2563 672 2643 724
rect 2563 626 2580 672
rect 2626 626 2643 672
rect 2563 574 2643 626
rect 2563 528 2580 574
rect 2626 528 2643 574
rect 2563 476 2643 528
rect 2563 430 2580 476
rect 2626 430 2643 476
rect 2563 378 2643 430
rect 2563 332 2580 378
rect 2626 332 2643 378
rect 2563 280 2643 332
rect 2563 234 2580 280
rect 2626 234 2643 280
rect 2563 182 2643 234
rect 2563 136 2580 182
rect 2626 136 2643 182
rect 2563 84 2643 136
rect 2563 38 2580 84
rect 2626 38 2643 84
rect -453 -60 -437 -14
rect -391 -60 -374 -14
rect -453 -112 -374 -60
rect -453 -158 -437 -112
rect -391 -158 -374 -112
rect -453 -210 -374 -158
rect -453 -256 -437 -210
rect -391 -256 -374 -210
rect 2563 -14 2643 38
rect 2563 -60 2580 -14
rect 2626 -60 2643 -14
rect -453 -308 -374 -256
rect -453 -354 -437 -308
rect -391 -354 -374 -308
rect 2563 -112 2643 -60
rect 2563 -158 2580 -112
rect 2626 -158 2643 -112
rect 2563 -210 2643 -158
rect 2563 -256 2580 -210
rect 2626 -256 2643 -210
rect 2563 -308 2643 -256
rect -453 -406 -374 -354
rect -453 -452 -437 -406
rect -391 -452 -374 -406
rect -453 -504 -374 -452
rect -453 -550 -437 -504
rect -391 -550 -374 -504
rect -453 -602 -374 -550
rect -453 -648 -437 -602
rect -391 -648 -374 -602
rect -453 -700 -374 -648
rect -453 -746 -437 -700
rect -391 -746 -374 -700
rect -453 -798 -374 -746
rect -453 -844 -437 -798
rect -391 -844 -374 -798
rect -453 -896 -374 -844
rect -453 -942 -437 -896
rect -391 -942 -374 -896
rect -453 -977 -374 -942
rect 2563 -354 2580 -308
rect 2626 -354 2643 -308
rect 2563 -406 2643 -354
rect 2563 -452 2580 -406
rect 2626 -452 2643 -406
rect 2563 -504 2643 -452
rect 2563 -550 2580 -504
rect 2626 -550 2643 -504
rect 2563 -602 2643 -550
rect 2563 -648 2580 -602
rect 2626 -648 2643 -602
rect 2563 -700 2643 -648
rect 2563 -746 2580 -700
rect 2626 -746 2643 -700
rect 2563 -798 2643 -746
rect 2563 -844 2580 -798
rect 2626 -844 2643 -798
rect 2563 -896 2643 -844
rect 2563 -942 2580 -896
rect 2626 -942 2643 -896
rect 2563 -977 2643 -942
rect -453 -994 2643 -977
rect -453 -1040 -437 -994
rect -391 -1040 -339 -994
rect -293 -1040 -241 -994
rect -195 -1040 -143 -994
rect -97 -1040 -33 -994
rect 13 -1040 65 -994
rect 111 -1040 163 -994
rect 209 -1040 261 -994
rect 307 -1040 359 -994
rect 405 -1040 457 -994
rect 503 -1040 555 -994
rect 601 -1040 653 -994
rect 699 -1040 751 -994
rect 797 -1040 849 -994
rect 895 -1040 947 -994
rect 993 -1040 1045 -994
rect 1091 -1040 1143 -994
rect 1189 -1040 1241 -994
rect 1287 -1040 1339 -994
rect 1385 -1040 1437 -994
rect 1483 -1040 1535 -994
rect 1581 -1040 1633 -994
rect 1679 -1040 1731 -994
rect 1777 -1040 1829 -994
rect 1875 -1040 1927 -994
rect 1973 -1040 2025 -994
rect 2071 -1040 2123 -994
rect 2169 -1040 2221 -994
rect 2267 -1040 2319 -994
rect 2365 -1040 2417 -994
rect 2463 -1040 2580 -994
rect 2626 -1040 2643 -994
rect -453 -1057 2643 -1040
<< psubdiffcont >>
rect -437 822 -391 868
rect -339 822 -293 868
rect -241 822 -195 868
rect -143 822 -97 868
rect -33 822 13 868
rect 65 822 111 868
rect 163 822 209 868
rect 261 822 307 868
rect 359 822 405 868
rect 457 822 503 868
rect 555 822 601 868
rect 653 822 699 868
rect 751 822 797 868
rect 849 822 895 868
rect 947 822 993 868
rect 1045 822 1091 868
rect 1143 822 1189 868
rect 1241 822 1287 868
rect 1339 822 1385 868
rect 1437 822 1483 868
rect 1535 822 1581 868
rect 1633 822 1679 868
rect 1731 822 1777 868
rect 1829 822 1875 868
rect 1927 822 1973 868
rect 2025 822 2071 868
rect 2123 822 2169 868
rect 2221 822 2267 868
rect 2319 822 2365 868
rect 2417 822 2463 868
rect 2580 822 2626 868
rect -437 724 -391 770
rect -437 626 -391 672
rect -437 528 -391 574
rect -437 430 -391 476
rect -437 332 -391 378
rect -437 234 -391 280
rect -437 136 -391 182
rect -437 38 -391 84
rect 2580 724 2626 770
rect 2580 626 2626 672
rect 2580 528 2626 574
rect 2580 430 2626 476
rect 2580 332 2626 378
rect 2580 234 2626 280
rect 2580 136 2626 182
rect 2580 38 2626 84
rect -437 -60 -391 -14
rect -437 -158 -391 -112
rect -437 -256 -391 -210
rect 2580 -60 2626 -14
rect -437 -354 -391 -308
rect 2580 -158 2626 -112
rect 2580 -256 2626 -210
rect -437 -452 -391 -406
rect -437 -550 -391 -504
rect -437 -648 -391 -602
rect -437 -746 -391 -700
rect -437 -844 -391 -798
rect -437 -942 -391 -896
rect 2580 -354 2626 -308
rect 2580 -452 2626 -406
rect 2580 -550 2626 -504
rect 2580 -648 2626 -602
rect 2580 -746 2626 -700
rect 2580 -844 2626 -798
rect 2580 -942 2626 -896
rect -437 -1040 -391 -994
rect -339 -1040 -293 -994
rect -241 -1040 -195 -994
rect -143 -1040 -97 -994
rect -33 -1040 13 -994
rect 65 -1040 111 -994
rect 163 -1040 209 -994
rect 261 -1040 307 -994
rect 359 -1040 405 -994
rect 457 -1040 503 -994
rect 555 -1040 601 -994
rect 653 -1040 699 -994
rect 751 -1040 797 -994
rect 849 -1040 895 -994
rect 947 -1040 993 -994
rect 1045 -1040 1091 -994
rect 1143 -1040 1189 -994
rect 1241 -1040 1287 -994
rect 1339 -1040 1385 -994
rect 1437 -1040 1483 -994
rect 1535 -1040 1581 -994
rect 1633 -1040 1679 -994
rect 1731 -1040 1777 -994
rect 1829 -1040 1875 -994
rect 1927 -1040 1973 -994
rect 2025 -1040 2071 -994
rect 2123 -1040 2169 -994
rect 2221 -1040 2267 -994
rect 2319 -1040 2365 -994
rect 2417 -1040 2463 -994
rect 2580 -1040 2626 -994
<< polysilicon >>
rect -222 -61 -121 25
rect 29 24 214 34
rect 318 24 705 33
rect 869 24 1273 33
rect 1420 24 1810 33
rect 29 -18 2070 24
rect -303 -121 -47 -61
rect 29 -64 57 -18
rect 103 -64 392 -18
rect 438 -64 631 -18
rect 677 -64 969 -18
rect 1015 -19 1521 -18
rect 1015 -64 1186 -19
rect 29 -65 1186 -64
rect 1232 -64 1521 -19
rect 1567 -64 1715 -18
rect 1761 -64 2070 -18
rect 1232 -65 2070 -64
rect 29 -66 2070 -65
rect 29 -82 132 -66
rect 364 -82 467 -66
rect 603 -82 706 -66
rect 941 -82 1044 -66
rect 1158 -83 1261 -66
rect 1493 -82 1596 -66
rect 1687 -82 1790 -66
rect 2304 -74 2405 30
rect -303 -167 -289 -121
rect -243 -123 -47 -121
rect -243 -167 -125 -123
rect -303 -169 -125 -167
rect -79 -169 -47 -123
rect -303 -242 -47 -169
rect 2227 -137 2483 -74
rect 2227 -183 2245 -137
rect 2291 -183 2397 -137
rect 2443 -183 2483 -137
rect 29 -225 132 -209
rect 389 -225 492 -209
rect -222 -322 -121 -242
rect 29 -271 57 -225
rect 103 -271 417 -225
rect 463 -226 492 -225
rect 599 -225 702 -209
rect 961 -225 1064 -210
rect 1156 -225 1259 -209
rect 1495 -225 1598 -209
rect 1703 -225 1806 -209
rect 599 -226 627 -225
rect 463 -271 627 -226
rect 673 -226 1184 -225
rect 673 -271 989 -226
rect 29 -272 989 -271
rect 1035 -271 1184 -226
rect 1230 -271 1523 -225
rect 1569 -271 1731 -225
rect 1777 -271 2073 -225
rect 2227 -255 2483 -183
rect 1035 -272 2073 -271
rect 29 -315 2073 -272
rect 29 -325 214 -315
rect 318 -326 712 -315
rect 869 -325 1288 -315
rect 1420 -325 1847 -315
rect 2304 -317 2405 -255
<< polycontact >>
rect 57 -64 103 -18
rect 392 -64 438 -18
rect 631 -64 677 -18
rect 969 -64 1015 -18
rect 1186 -65 1232 -19
rect 1521 -64 1567 -18
rect 1715 -64 1761 -18
rect -289 -167 -243 -121
rect -125 -169 -79 -123
rect 2245 -183 2291 -137
rect 2397 -183 2443 -137
rect 57 -271 103 -225
rect 417 -271 463 -225
rect 627 -271 673 -225
rect 989 -272 1035 -226
rect 1184 -271 1230 -225
rect 1523 -271 1569 -225
rect 1731 -271 1777 -225
<< metal1 >>
rect -453 868 2643 885
rect -453 822 -437 868
rect -391 822 -339 868
rect -293 822 -241 868
rect -195 822 -143 868
rect -97 822 -33 868
rect 13 822 65 868
rect 111 822 163 868
rect 209 822 261 868
rect 307 822 359 868
rect 405 822 457 868
rect 503 822 555 868
rect 601 822 653 868
rect 699 822 751 868
rect 797 822 849 868
rect 895 822 947 868
rect 993 822 1045 868
rect 1091 822 1143 868
rect 1189 822 1241 868
rect 1287 822 1339 868
rect 1385 822 1437 868
rect 1483 822 1535 868
rect 1581 822 1633 868
rect 1679 822 1731 868
rect 1777 822 1829 868
rect 1875 822 1927 868
rect 1973 822 2025 868
rect 2071 822 2123 868
rect 2169 822 2221 868
rect 2267 822 2319 868
rect 2365 822 2417 868
rect 2463 822 2580 868
rect 2626 822 2643 868
rect -453 805 2643 822
rect -453 770 -374 805
rect -453 724 -437 770
rect -391 724 -374 770
rect -453 672 -374 724
rect -453 626 -437 672
rect -391 626 -374 672
rect -453 574 -374 626
rect -453 528 -437 574
rect -391 528 -374 574
rect -303 530 -241 805
rect -453 476 -374 528
rect -453 430 -437 476
rect -391 430 -374 476
rect -453 378 -374 430
rect -453 332 -437 378
rect -391 332 -374 378
rect -453 280 -374 332
rect -453 234 -437 280
rect -391 234 -374 280
rect -453 182 -374 234
rect -453 136 -437 182
rect -391 136 -374 182
rect -453 84 -374 136
rect -453 38 -437 84
rect -391 38 -374 84
rect -453 -14 -374 38
rect -453 -60 -437 -14
rect -391 -60 -374 -14
rect -453 -112 -374 -60
rect -301 -61 -244 530
rect -103 523 -41 805
rect -98 -61 -41 523
rect 12 604 517 713
rect 12 64 103 604
rect -453 -158 -437 -112
rect -391 -158 -374 -112
rect -453 -210 -374 -158
rect -453 -256 -437 -210
rect -391 -256 -374 -210
rect -303 -121 -41 -61
rect 29 -14 132 -2
rect 29 -70 52 -14
rect 108 -70 132 -14
rect 29 -82 132 -70
rect -303 -167 -289 -121
rect -243 -123 -41 -121
rect -243 -167 -125 -123
rect -303 -169 -125 -167
rect -79 -169 -41 -123
rect -303 -242 -41 -169
rect -453 -308 -374 -256
rect -453 -354 -437 -308
rect -391 -354 -374 -308
rect -453 -406 -374 -354
rect -453 -452 -437 -406
rect -391 -452 -374 -406
rect -453 -504 -374 -452
rect -453 -550 -437 -504
rect -391 -550 -374 -504
rect -453 -602 -374 -550
rect -453 -648 -437 -602
rect -391 -648 -374 -602
rect -453 -700 -374 -648
rect -453 -746 -437 -700
rect -391 -746 -374 -700
rect -301 -730 -244 -242
rect -453 -798 -374 -746
rect -453 -844 -437 -798
rect -391 -844 -374 -798
rect -453 -896 -374 -844
rect -453 -942 -437 -896
rect -391 -942 -374 -896
rect -453 -977 -374 -942
rect -306 -977 -244 -730
rect -98 -747 -41 -242
rect 29 -221 132 -209
rect 29 -277 52 -221
rect 108 -277 132 -221
rect 29 -289 132 -277
rect -103 -977 -41 -747
rect 21 -977 113 -349
rect 214 -835 316 548
rect 426 68 517 604
rect 563 604 1068 713
rect 563 64 654 604
rect 364 -14 467 -2
rect 364 -70 387 -14
rect 443 -70 467 -14
rect 364 -82 467 -70
rect 603 -14 706 -2
rect 603 -70 626 -14
rect 682 -70 706 -14
rect 603 -82 706 -70
rect 389 -221 492 -209
rect 389 -277 412 -221
rect 468 -277 492 -221
rect 389 -289 492 -277
rect 599 -221 702 -209
rect 599 -277 622 -221
rect 678 -277 702 -221
rect 599 -289 702 -277
rect 419 -977 520 -343
rect 572 -977 664 -349
rect 765 -835 867 548
rect 977 68 1068 604
rect 1114 604 1619 713
rect 1114 64 1205 604
rect 941 -14 1044 -2
rect 941 -70 964 -14
rect 1020 -70 1044 -14
rect 941 -82 1044 -70
rect 1158 -15 1261 -3
rect 1158 -71 1181 -15
rect 1237 -71 1261 -15
rect 1158 -83 1261 -71
rect 961 -222 1064 -210
rect 961 -278 984 -222
rect 1040 -278 1064 -222
rect 961 -290 1064 -278
rect 1156 -221 1259 -209
rect 1156 -277 1179 -221
rect 1235 -277 1259 -221
rect 1156 -289 1259 -277
rect 970 -977 1071 -343
rect 1123 -977 1215 -349
rect 1316 -835 1418 548
rect 1528 68 1619 604
rect 1665 604 2170 713
rect 1665 64 1756 604
rect 1493 -14 1596 -2
rect 1493 -70 1516 -14
rect 1572 -70 1596 -14
rect 1493 -82 1596 -70
rect 1687 -14 1790 -2
rect 1687 -70 1710 -14
rect 1766 -70 1790 -14
rect 1687 -82 1790 -70
rect 1495 -221 1598 -209
rect 1495 -277 1518 -221
rect 1574 -277 1598 -221
rect 1495 -289 1598 -277
rect 1703 -221 1806 -209
rect 1703 -277 1726 -221
rect 1782 -277 1806 -221
rect 1703 -289 1806 -277
rect 1521 -977 1622 -343
rect 1674 -977 1766 -349
rect 1867 -835 1969 548
rect 2079 68 2170 604
rect 2221 521 2283 805
rect 2431 526 2493 805
rect 2563 770 2643 805
rect 2563 724 2580 770
rect 2626 724 2643 770
rect 2563 672 2643 724
rect 2563 626 2580 672
rect 2626 626 2643 672
rect 2563 574 2643 626
rect 2563 528 2580 574
rect 2626 528 2643 574
rect 2222 -74 2279 521
rect 2431 -74 2488 526
rect 2222 -137 2488 -74
rect 2222 -183 2245 -137
rect 2291 -183 2397 -137
rect 2443 -183 2488 -137
rect 2222 -255 2488 -183
rect 2072 -977 2173 -343
rect 2222 -750 2279 -255
rect 2431 -741 2488 -255
rect 2563 476 2643 528
rect 2563 430 2580 476
rect 2626 430 2643 476
rect 2563 378 2643 430
rect 2563 332 2580 378
rect 2626 332 2643 378
rect 2563 280 2643 332
rect 2563 234 2580 280
rect 2626 234 2643 280
rect 2563 182 2643 234
rect 2563 136 2580 182
rect 2626 136 2643 182
rect 2563 84 2643 136
rect 2563 38 2580 84
rect 2626 38 2643 84
rect 2563 -14 2643 38
rect 2563 -60 2580 -14
rect 2626 -60 2643 -14
rect 2563 -112 2643 -60
rect 2563 -158 2580 -112
rect 2626 -158 2643 -112
rect 2563 -210 2643 -158
rect 2563 -256 2580 -210
rect 2626 -256 2643 -210
rect 2563 -308 2643 -256
rect 2563 -354 2580 -308
rect 2626 -354 2643 -308
rect 2563 -406 2643 -354
rect 2563 -452 2580 -406
rect 2626 -452 2643 -406
rect 2563 -504 2643 -452
rect 2563 -550 2580 -504
rect 2626 -550 2643 -504
rect 2563 -602 2643 -550
rect 2563 -648 2580 -602
rect 2626 -648 2643 -602
rect 2563 -700 2643 -648
rect 2221 -977 2283 -750
rect 2431 -977 2493 -741
rect 2563 -746 2580 -700
rect 2626 -746 2643 -700
rect 2563 -798 2643 -746
rect 2563 -844 2580 -798
rect 2626 -844 2643 -798
rect 2563 -896 2643 -844
rect 2563 -942 2580 -896
rect 2626 -942 2643 -896
rect 2563 -977 2643 -942
rect -453 -994 2643 -977
rect -453 -1040 -437 -994
rect -391 -1040 -339 -994
rect -293 -1040 -241 -994
rect -195 -1040 -143 -994
rect -97 -1040 -33 -994
rect 13 -1040 65 -994
rect 111 -1040 163 -994
rect 209 -1040 261 -994
rect 307 -1040 359 -994
rect 405 -1040 457 -994
rect 503 -1040 555 -994
rect 601 -1040 653 -994
rect 699 -1040 751 -994
rect 797 -1040 849 -994
rect 895 -1040 947 -994
rect 993 -1040 1045 -994
rect 1091 -1040 1143 -994
rect 1189 -1040 1241 -994
rect 1287 -1040 1339 -994
rect 1385 -1040 1437 -994
rect 1483 -1040 1535 -994
rect 1581 -1040 1633 -994
rect 1679 -1040 1731 -994
rect 1777 -1040 1829 -994
rect 1875 -1040 1927 -994
rect 1973 -1040 2025 -994
rect 2071 -1040 2123 -994
rect 2169 -1040 2221 -994
rect 2267 -1040 2319 -994
rect 2365 -1040 2417 -994
rect 2463 -1040 2580 -994
rect 2626 -1040 2643 -994
rect -453 -1057 2643 -1040
rect 419 -1060 520 -1057
<< via1 >>
rect 52 -18 108 -14
rect 52 -64 57 -18
rect 57 -64 103 -18
rect 103 -64 108 -18
rect 52 -70 108 -64
rect 52 -225 108 -221
rect 52 -271 57 -225
rect 57 -271 103 -225
rect 103 -271 108 -225
rect 52 -277 108 -271
rect 387 -18 443 -14
rect 387 -64 392 -18
rect 392 -64 438 -18
rect 438 -64 443 -18
rect 387 -70 443 -64
rect 626 -18 682 -14
rect 626 -64 631 -18
rect 631 -64 677 -18
rect 677 -64 682 -18
rect 626 -70 682 -64
rect 412 -225 468 -221
rect 412 -271 417 -225
rect 417 -271 463 -225
rect 463 -271 468 -225
rect 412 -277 468 -271
rect 622 -225 678 -221
rect 622 -271 627 -225
rect 627 -271 673 -225
rect 673 -271 678 -225
rect 622 -277 678 -271
rect 964 -18 1020 -14
rect 964 -64 969 -18
rect 969 -64 1015 -18
rect 1015 -64 1020 -18
rect 964 -70 1020 -64
rect 1181 -19 1237 -15
rect 1181 -65 1186 -19
rect 1186 -65 1232 -19
rect 1232 -65 1237 -19
rect 1181 -71 1237 -65
rect 984 -226 1040 -222
rect 984 -272 989 -226
rect 989 -272 1035 -226
rect 1035 -272 1040 -226
rect 984 -278 1040 -272
rect 1179 -225 1235 -221
rect 1179 -271 1184 -225
rect 1184 -271 1230 -225
rect 1230 -271 1235 -225
rect 1179 -277 1235 -271
rect 1516 -18 1572 -14
rect 1516 -64 1521 -18
rect 1521 -64 1567 -18
rect 1567 -64 1572 -18
rect 1516 -70 1572 -64
rect 1710 -18 1766 -14
rect 1710 -64 1715 -18
rect 1715 -64 1761 -18
rect 1761 -64 1766 -18
rect 1710 -70 1766 -64
rect 1518 -225 1574 -221
rect 1518 -271 1523 -225
rect 1523 -271 1569 -225
rect 1569 -271 1574 -225
rect 1518 -277 1574 -271
rect 1726 -225 1782 -221
rect 1726 -271 1731 -225
rect 1731 -271 1777 -225
rect 1777 -271 1782 -225
rect 1726 -277 1782 -271
<< metal2 >>
rect -658 -14 2073 -2
rect -658 -70 52 -14
rect 108 -70 387 -14
rect 443 -70 626 -14
rect 682 -70 964 -14
rect 1020 -15 1516 -14
rect 1020 -70 1181 -15
rect -658 -71 1181 -70
rect 1237 -70 1516 -15
rect 1572 -70 1710 -14
rect 1766 -70 2073 -14
rect 1237 -71 2073 -70
rect -658 -82 2073 -71
rect 1158 -83 1261 -82
rect -680 -221 2073 -209
rect -680 -277 52 -221
rect 108 -277 412 -221
rect 468 -277 622 -221
rect 678 -222 1179 -221
rect 678 -277 984 -222
rect -680 -278 984 -277
rect 1040 -277 1179 -222
rect 1235 -277 1518 -221
rect 1574 -277 1726 -221
rect 1782 -277 2073 -221
rect 1040 -278 2073 -277
rect -680 -289 2073 -278
rect 961 -290 1064 -289
use nfet_03v3_CT75PZ  nfet_03v3_CT75PZ_0
timestamp 1699925801
transform 1 0 1919 0 1 -599
box -264 -308 264 308
use nfet_03v3_CT75PZ  nfet_03v3_CT75PZ_1
timestamp 1699925801
transform 1 0 1919 0 1 308
box -264 -308 264 308
use nfet_03v3_CT75PZ  nfet_03v3_CT75PZ_2
timestamp 1699925801
transform 1 0 266 0 1 308
box -264 -308 264 308
use nfet_03v3_CT75PZ  nfet_03v3_CT75PZ_3
timestamp 1699925801
transform 1 0 266 0 1 -599
box -264 -308 264 308
use nfet_03v3_CT75PZ  nfet_03v3_CT75PZ_4
timestamp 1699925801
transform 1 0 817 0 1 -599
box -264 -308 264 308
use nfet_03v3_CT75PZ  nfet_03v3_CT75PZ_5
timestamp 1699925801
transform 1 0 817 0 1 308
box -264 -308 264 308
use nfet_03v3_CT75PZ  nfet_03v3_CT75PZ_6
timestamp 1699925801
transform 1 0 1368 0 1 -599
box -264 -308 264 308
use nfet_03v3_CT75PZ  nfet_03v3_CT75PZ_7
timestamp 1699925801
transform 1 0 1368 0 1 308
box -264 -308 264 308
use nfet_03v3_CTB5PZ  nfet_03v3_CTB5PZ_0
timestamp 1699938072
transform 1 0 -170 0 1 -600
box -162 -308 162 308
use nfet_03v3_CTB5PZ  nfet_03v3_CTB5PZ_1
timestamp 1699938072
transform 1 0 -170 0 1 308
box -162 -308 162 308
use nfet_03v3_CTB5PZ  nfet_03v3_CTB5PZ_2
timestamp 1699938072
transform 1 0 2354 0 1 -599
box -162 -308 162 308
use nfet_03v3_CTB5PZ  nfet_03v3_CTB5PZ_3
timestamp 1699938072
transform 1 0 2356 0 1 310
box -162 -308 162 308
<< labels >>
flabel metal1 38 657 38 657 0 FreeSans 480 0 0 0 IBIAS_BUF1
port 9 nsew
flabel metal1 724 639 724 639 0 FreeSans 480 0 0 0 IBIAS_BUF2
port 10 nsew
flabel metal1 1380 660 1380 660 0 FreeSans 480 0 0 0 IBIAS_FILTER
port 11 nsew
flabel metal1 1890 676 1890 676 0 FreeSans 480 0 0 0 IBIAS_PGA
port 13 nsew
flabel metal2 -627 -52 -627 -52 0 FreeSans 800 0 0 0 G_SINK_UP
port 14 nsew
flabel metal2 -617 -252 -617 -252 0 FreeSans 800 0 0 0 G_SINK_DOWN
port 16 nsew
flabel metal1 244 -1007 244 -1007 0 FreeSans 800 0 0 0 VSS
port 18 nsew
<< end >>
