magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2000 -2989 3784 2579
<< nwell >>
rect 0 466 1784 579
rect 985 -78 988 86
<< pwell >>
rect 830 -861 954 -501
<< psubdiff >>
rect 783 -926 980 -908
rect 783 -972 859 -926
rect 905 -972 980 -926
rect 783 -989 980 -972
<< nsubdiff >>
rect 634 538 880 552
rect 634 492 714 538
rect 760 492 880 538
rect 634 476 880 492
<< psubdiffcont >>
rect 859 -972 905 -926
<< nsubdiffcont >>
rect 714 492 760 538
<< polysilicon >>
rect 174 381 718 419
rect 1066 382 1610 420
rect 174 86 286 118
rect 78 13 286 86
rect 78 -33 95 13
rect 141 -33 286 13
rect 78 -78 286 -33
rect 174 -96 286 -78
rect 390 -96 502 118
rect 606 -100 718 114
rect 1066 86 1178 107
rect 985 18 1178 86
rect 985 -28 999 18
rect 1045 -28 1178 18
rect 985 -78 1178 -28
rect 1066 -97 1178 -78
rect 1282 -95 1394 109
rect 1498 -91 1610 113
rect 174 -537 286 -370
rect 390 -536 502 -369
rect 606 -534 718 -367
rect 1066 -534 1178 -367
rect 1282 -532 1394 -365
rect 1498 -532 1610 -365
rect 174 -864 718 -827
rect 1066 -864 1610 -827
<< polycontact >>
rect 95 -33 141 13
rect 999 -28 1045 18
<< metal1 >>
rect 84 538 1700 552
rect 84 492 714 538
rect 760 492 1700 538
rect 84 476 1700 492
rect 99 344 145 476
rect 99 173 147 344
rect 315 297 361 352
rect 298 284 376 297
rect 298 232 311 284
rect 363 232 376 284
rect 298 219 376 232
rect 99 132 268 173
rect 101 127 268 132
rect 74 16 157 25
rect 39 14 157 16
rect 39 -35 89 14
rect 74 -38 89 -35
rect 141 -38 157 14
rect 74 -51 157 -38
rect 99 -242 145 -124
rect 222 -242 268 127
rect 99 -288 268 -242
rect 99 -344 145 -288
rect 99 -908 145 -571
rect 315 -629 361 219
rect 531 -344 577 476
rect 747 296 793 352
rect 991 344 1037 476
rect 991 340 1038 344
rect 732 283 810 296
rect 732 231 745 283
rect 797 231 810 283
rect 732 218 810 231
rect 747 20 793 218
rect 992 197 1038 340
rect 1207 312 1253 352
rect 1191 299 1269 312
rect 1191 247 1204 299
rect 1256 247 1269 299
rect 1191 234 1269 247
rect 992 151 1159 197
rect 988 20 1056 29
rect 747 18 1056 20
rect 747 -28 999 18
rect 1045 -28 1056 18
rect 747 -32 1056 -28
rect 301 -642 378 -629
rect 301 -694 313 -642
rect 365 -694 378 -642
rect 301 -706 378 -694
rect 315 -791 361 -706
rect 531 -908 577 -571
rect 747 -636 793 -32
rect 988 -39 1056 -32
rect 991 -255 1037 -124
rect 1113 -255 1159 151
rect 991 -301 1159 -255
rect 991 -344 1037 -301
rect 732 -649 809 -636
rect 732 -701 744 -649
rect 796 -701 809 -649
rect 732 -713 809 -701
rect 747 -791 793 -713
rect 991 -908 1037 -571
rect 1207 -622 1253 234
rect 1423 -344 1469 476
rect 1639 310 1685 352
rect 1625 297 1703 310
rect 1625 245 1638 297
rect 1690 245 1703 297
rect 1625 232 1703 245
rect 1639 3 1685 232
rect 1639 -43 1781 3
rect 1192 -635 1269 -622
rect 1192 -687 1204 -635
rect 1256 -687 1269 -635
rect 1192 -699 1269 -687
rect 1207 -791 1253 -699
rect 1423 -908 1469 -571
rect 1639 -622 1685 -43
rect 1625 -635 1702 -622
rect 1625 -687 1637 -635
rect 1689 -687 1702 -635
rect 1625 -699 1702 -687
rect 1639 -791 1685 -699
rect 77 -926 1708 -908
rect 77 -972 859 -926
rect 905 -972 1708 -926
rect 77 -989 1708 -972
<< via1 >>
rect 311 232 363 284
rect 89 13 141 14
rect 89 -33 95 13
rect 95 -33 141 13
rect 89 -38 141 -33
rect 745 231 797 283
rect 1204 247 1256 299
rect 313 -694 365 -642
rect 744 -701 796 -649
rect 1638 245 1690 297
rect 1204 -687 1256 -635
rect 1637 -687 1689 -635
<< metal2 >>
rect 1191 299 1269 312
rect 298 287 376 297
rect 732 287 810 296
rect 298 284 810 287
rect 298 232 311 284
rect 363 283 810 284
rect 363 232 745 283
rect 298 231 745 232
rect 797 231 810 283
rect 1191 247 1204 299
rect 1256 297 1269 299
rect 1625 297 1703 310
rect 1256 247 1638 297
rect 1191 245 1638 247
rect 1690 245 1703 297
rect 1191 237 1703 245
rect 1191 234 1269 237
rect 1625 232 1703 237
rect 298 228 810 231
rect 298 219 376 228
rect 732 218 810 228
rect 74 14 157 25
rect 74 -38 89 14
rect 141 -38 157 14
rect 74 -51 157 -38
rect 301 -638 378 -629
rect 1192 -632 1269 -622
rect 1625 -632 1702 -622
rect 1192 -635 1702 -632
rect 732 -638 809 -636
rect 301 -642 809 -638
rect 301 -694 313 -642
rect 365 -649 809 -642
rect 365 -694 744 -649
rect 301 -696 744 -694
rect 301 -706 378 -696
rect 732 -701 744 -696
rect 796 -701 809 -649
rect 1192 -687 1204 -635
rect 1256 -687 1637 -635
rect 1689 -687 1702 -635
rect 1192 -690 1702 -687
rect 1192 -699 1269 -690
rect 1625 -699 1702 -690
rect 732 -713 809 -701
use nmos_3p3_G2UGVV  nmos_3p3_G2UGVV_0
timestamp 1713185578
transform 1 0 1338 0 1 -681
box -384 -180 384 180
use nmos_3p3_G2UGVV  nmos_3p3_G2UGVV_1
timestamp 1713185578
transform 1 0 446 0 1 -681
box -384 -180 384 180
use pmos_3p3_VRY6F7  pmos_3p3_VRY6F7_0
timestamp 1713185578
transform 1 0 446 0 1 -234
box -446 -242 446 242
use pmos_3p3_VRY6F7  pmos_3p3_VRY6F7_1
timestamp 1713185578
transform 1 0 1338 0 1 -234
box -446 -242 446 242
use pmos_3p3_VRY6F7  pmos_3p3_VRY6F7_2
timestamp 1713185578
transform 1 0 446 0 1 242
box -446 -242 446 242
use pmos_3p3_VRY6F7  pmos_3p3_VRY6F7_3
timestamp 1713185578
transform 1 0 1338 0 1 242
box -446 -242 446 242
<< labels >>
flabel nsubdiffcont 739 513 739 513 0 FreeSans 750 0 0 0 VDD
flabel psubdiffcont 882 -950 882 -950 0 FreeSans 750 0 0 0 VSS
<< end >>
