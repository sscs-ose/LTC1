magic
tech gf180mcuC
magscale 1 10
timestamp 1699683674
<< nwell >>
rect 2921 3726 5203 5254
rect 2921 3708 4519 3726
rect 4565 3708 5203 3726
rect 2921 1776 5203 3708
rect 7 -1916 5203 1776
rect 11377 2207 16573 2622
rect 11377 2150 12041 2207
rect 12087 2150 16573 2207
rect 11377 1193 16573 2150
rect 11377 1174 12314 1193
rect 12391 1174 13210 1193
rect 13287 1174 16573 1193
rect 11377 128 16573 1174
rect 11377 -52 13210 128
rect 13286 -52 16573 128
rect 11377 -272 16573 -52
rect 11377 -452 13498 -272
rect 13574 -452 16573 -272
rect 11377 -889 16573 -452
rect 11377 -890 13208 -889
rect 11377 -904 12313 -890
rect 12391 -903 13208 -890
rect 13286 -903 16573 -889
rect 12391 -904 16573 -903
rect 11377 -1916 16573 -904
rect 32106 -1815 40498 3099
rect 41802 -1815 50194 3099
rect 51498 -1815 59890 3099
rect 61194 -1815 65450 3099
rect 17590 -4251 31432 -3346
rect 17590 -4297 24268 -4251
rect 24352 -4297 31432 -4251
rect 386 -7140 4588 -4308
rect 17590 -5008 27456 -4297
rect 17590 -5012 26706 -5008
rect 26994 -5012 27456 -5008
rect 17590 -5291 27456 -5012
rect 17590 -5383 26256 -5291
rect 26732 -5383 27456 -5291
rect 27652 -5383 31432 -4297
rect 17590 -5429 26452 -5383
rect 26536 -5429 31432 -5383
rect 17590 -6206 31432 -5429
rect 17590 -6208 26994 -6206
rect 17590 -6223 27172 -6208
rect 27174 -6223 31432 -6206
rect 17590 -6269 26452 -6223
rect 26536 -6269 31432 -6223
rect 386 -7212 1327 -7140
rect 1399 -7212 4588 -7140
rect 386 -7758 4588 -7212
rect 17590 -7353 31432 -6269
rect 17590 -7490 23624 -7353
rect 23632 -7490 23812 -7353
rect 23820 -7355 31432 -7353
rect 23820 -7401 24262 -7355
rect 24548 -7401 31432 -7355
rect 23820 -7490 31432 -7401
rect 17590 -8218 31432 -7490
<< pwell >>
rect 8782 -5810 8858 -5760
rect 9827 -6689 10007 -6660
<< psubdiff >>
rect 5763 5508 8091 5521
rect 5763 5462 5776 5508
rect 5822 5462 5870 5508
rect 5916 5462 5964 5508
rect 6010 5462 6058 5508
rect 6104 5462 6152 5508
rect 6198 5462 6246 5508
rect 6292 5462 6340 5508
rect 6386 5462 6434 5508
rect 6480 5462 6528 5508
rect 6574 5462 6622 5508
rect 6668 5462 6716 5508
rect 6762 5462 6810 5508
rect 6856 5462 6904 5508
rect 6950 5462 6998 5508
rect 7044 5462 7092 5508
rect 7138 5462 7186 5508
rect 7232 5462 7280 5508
rect 7326 5462 7374 5508
rect 7420 5462 7468 5508
rect 7514 5462 7562 5508
rect 7608 5462 7656 5508
rect 7702 5462 7750 5508
rect 7796 5462 7844 5508
rect 7890 5462 7938 5508
rect 7984 5462 8032 5508
rect 8078 5462 8091 5508
rect 5763 5449 8091 5462
rect 5763 5414 5835 5449
rect 5763 5368 5776 5414
rect 5822 5368 5835 5414
rect 5763 5320 5835 5368
rect 5763 5274 5776 5320
rect 5822 5274 5835 5320
rect 5763 5226 5835 5274
rect 5763 5180 5776 5226
rect 5822 5180 5835 5226
rect 5763 5132 5835 5180
rect 5763 5086 5776 5132
rect 5822 5086 5835 5132
rect 5763 5038 5835 5086
rect 5763 4992 5776 5038
rect 5822 4992 5835 5038
rect 5763 4944 5835 4992
rect 5763 4898 5776 4944
rect 5822 4898 5835 4944
rect 5763 4850 5835 4898
rect 5763 4804 5776 4850
rect 5822 4804 5835 4850
rect 5763 4756 5835 4804
rect 5763 4710 5776 4756
rect 5822 4710 5835 4756
rect 5763 4662 5835 4710
rect 5763 4616 5776 4662
rect 5822 4616 5835 4662
rect 5763 4568 5835 4616
rect 5763 4522 5776 4568
rect 5822 4522 5835 4568
rect 8019 5414 8091 5449
rect 8019 5368 8032 5414
rect 8078 5368 8091 5414
rect 8019 5320 8091 5368
rect 8019 5274 8032 5320
rect 8078 5274 8091 5320
rect 8019 5226 8091 5274
rect 8019 5180 8032 5226
rect 8078 5180 8091 5226
rect 8019 5132 8091 5180
rect 8019 5086 8032 5132
rect 8078 5086 8091 5132
rect 8019 5038 8091 5086
rect 8019 4992 8032 5038
rect 8078 4992 8091 5038
rect 8019 4944 8091 4992
rect 8019 4898 8032 4944
rect 8078 4898 8091 4944
rect 8019 4850 8091 4898
rect 8019 4804 8032 4850
rect 8078 4804 8091 4850
rect 8019 4756 8091 4804
rect 8019 4710 8032 4756
rect 8078 4710 8091 4756
rect 8019 4662 8091 4710
rect 8019 4616 8032 4662
rect 8078 4616 8091 4662
rect 8019 4568 8091 4616
rect 5763 4474 5835 4522
rect 5763 4428 5776 4474
rect 5822 4428 5835 4474
rect 5763 4380 5835 4428
rect 5763 4334 5776 4380
rect 5822 4334 5835 4380
rect 5763 4286 5835 4334
rect 5763 4240 5776 4286
rect 5822 4240 5835 4286
rect 8019 4522 8032 4568
rect 8078 4522 8091 4568
rect 8019 4474 8091 4522
rect 8019 4428 8032 4474
rect 8078 4428 8091 4474
rect 8019 4380 8091 4428
rect 8019 4334 8032 4380
rect 8078 4334 8091 4380
rect 8019 4286 8091 4334
rect 5763 4192 5835 4240
rect 5763 4146 5776 4192
rect 5822 4146 5835 4192
rect 5763 4098 5835 4146
rect 5763 4052 5776 4098
rect 5822 4052 5835 4098
rect 5763 4004 5835 4052
rect 5763 3958 5776 4004
rect 5822 3958 5835 4004
rect 5763 3910 5835 3958
rect 5763 3864 5776 3910
rect 5822 3864 5835 3910
rect 5763 3816 5835 3864
rect 5763 3770 5776 3816
rect 5822 3770 5835 3816
rect 5763 3722 5835 3770
rect 5763 3676 5776 3722
rect 5822 3676 5835 3722
rect 8019 4240 8032 4286
rect 8078 4240 8091 4286
rect 8019 4192 8091 4240
rect 8019 4146 8032 4192
rect 8078 4146 8091 4192
rect 8019 4098 8091 4146
rect 8019 4052 8032 4098
rect 8078 4052 8091 4098
rect 8019 4004 8091 4052
rect 8019 3958 8032 4004
rect 8078 3958 8091 4004
rect 8019 3910 8091 3958
rect 8019 3864 8032 3910
rect 8078 3864 8091 3910
rect 8019 3816 8091 3864
rect 8019 3770 8032 3816
rect 8078 3770 8091 3816
rect 8019 3722 8091 3770
rect 5763 3628 5835 3676
rect 5763 3582 5776 3628
rect 5822 3582 5835 3628
rect 5763 3534 5835 3582
rect 5763 3488 5776 3534
rect 5822 3488 5835 3534
rect 5763 3440 5835 3488
rect 5763 3394 5776 3440
rect 5822 3394 5835 3440
rect 8019 3676 8032 3722
rect 8078 3676 8091 3722
rect 8019 3628 8091 3676
rect 8019 3582 8032 3628
rect 8078 3582 8091 3628
rect 8019 3534 8091 3582
rect 8019 3488 8032 3534
rect 8078 3488 8091 3534
rect 8019 3440 8091 3488
rect 5763 3346 5835 3394
rect 5763 3291 5776 3346
rect 5822 3291 5835 3346
rect 5763 3243 5835 3291
rect 5763 3197 5776 3243
rect 5822 3197 5835 3243
rect 5763 3149 5835 3197
rect 5763 3103 5776 3149
rect 5822 3103 5835 3149
rect 5763 3055 5835 3103
rect 5763 3009 5776 3055
rect 5822 3009 5835 3055
rect 5763 2961 5835 3009
rect 5763 2915 5776 2961
rect 5822 2915 5835 2961
rect 5763 2867 5835 2915
rect 5763 2821 5776 2867
rect 5822 2821 5835 2867
rect 5763 2773 5835 2821
rect 8019 3394 8032 3440
rect 8078 3394 8091 3440
rect 8019 3346 8091 3394
rect 8019 3291 8032 3346
rect 8078 3291 8091 3346
rect 8019 3243 8091 3291
rect 8019 3197 8032 3243
rect 8078 3197 8091 3243
rect 8019 3149 8091 3197
rect 8019 3103 8032 3149
rect 8078 3103 8091 3149
rect 8019 3055 8091 3103
rect 8019 3009 8032 3055
rect 8078 3009 8091 3055
rect 8019 2961 8091 3009
rect 8019 2915 8032 2961
rect 8078 2915 8091 2961
rect 8019 2867 8091 2915
rect 8019 2821 8032 2867
rect 8078 2821 8091 2867
rect 5763 2727 5776 2773
rect 5822 2727 5835 2773
rect 5763 2679 5835 2727
rect 5763 2633 5776 2679
rect 5822 2633 5835 2679
rect 5763 2585 5835 2633
rect 5763 2539 5776 2585
rect 5822 2539 5835 2585
rect 5763 2491 5835 2539
rect 8019 2773 8091 2821
rect 8019 2727 8032 2773
rect 8078 2727 8091 2773
rect 8019 2679 8091 2727
rect 8019 2633 8032 2679
rect 8078 2633 8091 2679
rect 8019 2585 8091 2633
rect 17637 4611 20717 4624
rect 17637 4565 17650 4611
rect 17696 4565 17744 4611
rect 17790 4565 17838 4611
rect 17884 4565 17932 4611
rect 17978 4565 18026 4611
rect 18072 4565 18120 4611
rect 18166 4565 18214 4611
rect 18260 4565 18308 4611
rect 18354 4565 18402 4611
rect 18448 4565 18496 4611
rect 18542 4565 18590 4611
rect 18636 4565 18684 4611
rect 18730 4565 18778 4611
rect 18824 4565 18872 4611
rect 18918 4565 18966 4611
rect 19012 4565 19060 4611
rect 19106 4565 19154 4611
rect 19200 4565 19248 4611
rect 19294 4565 19342 4611
rect 19388 4565 19436 4611
rect 19482 4565 19530 4611
rect 19576 4565 19624 4611
rect 19670 4565 19718 4611
rect 19764 4565 19812 4611
rect 19858 4565 19906 4611
rect 19952 4565 20000 4611
rect 20046 4565 20094 4611
rect 20140 4565 20188 4611
rect 20234 4565 20282 4611
rect 20328 4565 20376 4611
rect 20422 4565 20470 4611
rect 20516 4565 20564 4611
rect 20610 4565 20658 4611
rect 20704 4565 20717 4611
rect 17637 4552 20717 4565
rect 17637 4517 17709 4552
rect 17637 4471 17650 4517
rect 17696 4471 17709 4517
rect 17637 4423 17709 4471
rect 17637 4377 17650 4423
rect 17696 4377 17709 4423
rect 17637 4329 17709 4377
rect 17637 4283 17650 4329
rect 17696 4283 17709 4329
rect 17637 4235 17709 4283
rect 20645 4517 20717 4552
rect 20645 4471 20658 4517
rect 20704 4471 20717 4517
rect 20645 4423 20717 4471
rect 20645 4377 20658 4423
rect 20704 4377 20717 4423
rect 20645 4329 20717 4377
rect 20645 4283 20658 4329
rect 20704 4283 20717 4329
rect 17637 4189 17650 4235
rect 17696 4189 17709 4235
rect 17637 4141 17709 4189
rect 20645 4235 20717 4283
rect 20645 4189 20658 4235
rect 20704 4189 20717 4235
rect 17637 4095 17650 4141
rect 17696 4095 17709 4141
rect 17637 4047 17709 4095
rect 17637 4001 17650 4047
rect 17696 4001 17709 4047
rect 20645 4141 20717 4189
rect 20645 4095 20658 4141
rect 20704 4095 20717 4141
rect 20645 4047 20717 4095
rect 17637 3953 17709 4001
rect 17637 3907 17650 3953
rect 17696 3907 17709 3953
rect 17637 3859 17709 3907
rect 17637 3813 17650 3859
rect 17696 3813 17709 3859
rect 17637 3765 17709 3813
rect 17637 3719 17650 3765
rect 17696 3719 17709 3765
rect 17637 3671 17709 3719
rect 17637 3625 17650 3671
rect 17696 3625 17709 3671
rect 17637 3577 17709 3625
rect 17637 3531 17650 3577
rect 17696 3531 17709 3577
rect 17637 3483 17709 3531
rect 17637 3437 17650 3483
rect 17696 3437 17709 3483
rect 17637 3389 17709 3437
rect 20645 4001 20658 4047
rect 20704 4001 20717 4047
rect 20645 3953 20717 4001
rect 20645 3907 20658 3953
rect 20704 3907 20717 3953
rect 20645 3859 20717 3907
rect 20645 3813 20658 3859
rect 20704 3813 20717 3859
rect 20645 3765 20717 3813
rect 20645 3719 20658 3765
rect 20704 3719 20717 3765
rect 20645 3671 20717 3719
rect 20645 3625 20658 3671
rect 20704 3625 20717 3671
rect 20645 3577 20717 3625
rect 20645 3531 20658 3577
rect 20704 3531 20717 3577
rect 20645 3483 20717 3531
rect 20645 3437 20658 3483
rect 20704 3437 20717 3483
rect 17637 3343 17650 3389
rect 17696 3343 17709 3389
rect 17637 3295 17709 3343
rect 17637 3249 17650 3295
rect 17696 3249 17709 3295
rect 17637 3201 17709 3249
rect 20645 3389 20717 3437
rect 20645 3343 20658 3389
rect 20704 3343 20717 3389
rect 17637 3155 17650 3201
rect 17696 3155 17709 3201
rect 17637 3107 17709 3155
rect 17637 3061 17650 3107
rect 17696 3061 17709 3107
rect 17637 3013 17709 3061
rect 17637 2967 17650 3013
rect 17696 2967 17709 3013
rect 17637 2919 17709 2967
rect 17637 2873 17650 2919
rect 17696 2873 17709 2919
rect 17637 2825 17709 2873
rect 17637 2779 17650 2825
rect 17696 2779 17709 2825
rect 17637 2731 17709 2779
rect 17637 2685 17650 2731
rect 17696 2685 17709 2731
rect 17637 2637 17709 2685
rect 8019 2539 8032 2585
rect 8078 2539 8091 2585
rect 5763 2445 5776 2491
rect 5822 2445 5835 2491
rect 5763 2397 5835 2445
rect 5763 2351 5776 2397
rect 5822 2351 5835 2397
rect 5763 2303 5835 2351
rect 5763 2257 5776 2303
rect 5822 2257 5835 2303
rect 5763 2209 5835 2257
rect 5763 2163 5776 2209
rect 5822 2163 5835 2209
rect 5763 2115 5835 2163
rect 5763 2069 5776 2115
rect 5822 2069 5835 2115
rect 5763 2021 5835 2069
rect 5763 1975 5776 2021
rect 5822 1975 5835 2021
rect 5763 1927 5835 1975
rect 8019 2491 8091 2539
rect 8019 2445 8032 2491
rect 8078 2445 8091 2491
rect 8019 2397 8091 2445
rect 8019 2351 8032 2397
rect 8078 2351 8091 2397
rect 8019 2303 8091 2351
rect 8019 2257 8032 2303
rect 8078 2257 8091 2303
rect 8019 2209 8091 2257
rect 8019 2163 8032 2209
rect 8078 2163 8091 2209
rect 8019 2115 8091 2163
rect 8019 2069 8032 2115
rect 8078 2069 8091 2115
rect 8019 2034 8091 2069
rect 8019 2021 10817 2034
rect 8019 1975 8032 2021
rect 8078 1975 8126 2021
rect 8172 1975 8220 2021
rect 8266 1975 8314 2021
rect 8360 1975 8408 2021
rect 8454 1975 8502 2021
rect 8548 1975 8596 2021
rect 8642 1975 8690 2021
rect 8736 1975 8784 2021
rect 8830 1975 8878 2021
rect 8924 1975 8972 2021
rect 9018 1975 9066 2021
rect 9112 1975 9160 2021
rect 9206 1975 9254 2021
rect 9300 1975 9348 2021
rect 9394 1975 9442 2021
rect 9488 1975 9536 2021
rect 9582 1975 9630 2021
rect 9676 1975 9724 2021
rect 9770 1975 9818 2021
rect 9864 1975 9912 2021
rect 9958 1975 10006 2021
rect 10052 1975 10100 2021
rect 10146 1975 10194 2021
rect 10240 1975 10288 2021
rect 10334 1975 10382 2021
rect 10428 1975 10476 2021
rect 10522 1975 10570 2021
rect 10616 1975 10664 2021
rect 10710 1975 10758 2021
rect 10804 1975 10817 2021
rect 8019 1962 10817 1975
rect 5763 1881 5776 1927
rect 5822 1881 5835 1927
rect 5763 1833 5835 1881
rect 5763 1787 5776 1833
rect 5822 1787 5835 1833
rect 5763 1739 5835 1787
rect 5763 1693 5776 1739
rect 5822 1693 5835 1739
rect 5763 1645 5835 1693
rect 8019 1927 8091 1962
rect 8019 1881 8032 1927
rect 8078 1881 8091 1927
rect 8019 1833 8091 1881
rect 8019 1787 8032 1833
rect 8078 1787 8091 1833
rect 8019 1739 8091 1787
rect 8019 1693 8032 1739
rect 8078 1693 8091 1739
rect 5763 1599 5776 1645
rect 5822 1599 5835 1645
rect 5763 1551 5835 1599
rect 5763 1505 5776 1551
rect 5822 1505 5835 1551
rect 5763 1457 5835 1505
rect 5763 1411 5776 1457
rect 5822 1411 5835 1457
rect 5763 1363 5835 1411
rect 5763 1317 5776 1363
rect 5822 1317 5835 1363
rect 5763 1269 5835 1317
rect 5763 1223 5776 1269
rect 5822 1223 5835 1269
rect 5763 1175 5835 1223
rect 5763 1129 5776 1175
rect 5822 1129 5835 1175
rect 5763 1081 5835 1129
rect 8019 1645 8091 1693
rect 8019 1599 8032 1645
rect 8078 1599 8091 1645
rect 8019 1551 8091 1599
rect 8019 1505 8032 1551
rect 8078 1505 8091 1551
rect 8019 1457 8091 1505
rect 8019 1411 8032 1457
rect 8078 1411 8091 1457
rect 8019 1363 8091 1411
rect 8019 1317 8032 1363
rect 8078 1317 8091 1363
rect 8019 1269 8091 1317
rect 8019 1223 8032 1269
rect 8078 1223 8091 1269
rect 8019 1175 8091 1223
rect 8019 1129 8032 1175
rect 8078 1129 8091 1175
rect 5763 1035 5776 1081
rect 5822 1035 5835 1081
rect 5763 987 5835 1035
rect 5763 941 5776 987
rect 5822 941 5835 987
rect 5763 893 5835 941
rect 5763 847 5776 893
rect 5822 847 5835 893
rect 5763 799 5835 847
rect 8019 1081 8091 1129
rect 8019 1035 8032 1081
rect 8078 1035 8091 1081
rect 10745 1927 10817 1962
rect 10745 1881 10758 1927
rect 10804 1881 10817 1927
rect 10745 1833 10817 1881
rect 10745 1787 10758 1833
rect 10804 1787 10817 1833
rect 10745 1739 10817 1787
rect 10745 1693 10758 1739
rect 10804 1693 10817 1739
rect 10745 1645 10817 1693
rect 10745 1599 10758 1645
rect 10804 1599 10817 1645
rect 10745 1551 10817 1599
rect 10745 1505 10758 1551
rect 10804 1505 10817 1551
rect 10745 1457 10817 1505
rect 10745 1411 10758 1457
rect 10804 1411 10817 1457
rect 10745 1363 10817 1411
rect 10745 1317 10758 1363
rect 10804 1317 10817 1363
rect 10745 1269 10817 1317
rect 10745 1223 10758 1269
rect 10804 1223 10817 1269
rect 10745 1175 10817 1223
rect 10745 1129 10758 1175
rect 10804 1129 10817 1175
rect 10745 1081 10817 1129
rect 8019 987 8091 1035
rect 8019 941 8032 987
rect 8078 941 8091 987
rect 8019 893 8091 941
rect 8019 847 8032 893
rect 8078 847 8091 893
rect 5763 753 5776 799
rect 5822 753 5835 799
rect 5763 705 5835 753
rect 5763 659 5776 705
rect 5822 659 5835 705
rect 5763 611 5835 659
rect 5763 565 5776 611
rect 5822 565 5835 611
rect 5763 517 5835 565
rect 5763 471 5776 517
rect 5822 471 5835 517
rect 5763 423 5835 471
rect 5763 377 5776 423
rect 5822 377 5835 423
rect 5763 329 5835 377
rect 5763 283 5776 329
rect 5822 283 5835 329
rect 5763 235 5835 283
rect 5763 189 5776 235
rect 5822 189 5835 235
rect 8019 799 8091 847
rect 8019 753 8032 799
rect 8078 753 8091 799
rect 10745 1035 10758 1081
rect 10804 1035 10817 1081
rect 10745 987 10817 1035
rect 10745 941 10758 987
rect 10804 941 10817 987
rect 10745 893 10817 941
rect 10745 847 10758 893
rect 10804 847 10817 893
rect 10745 799 10817 847
rect 8019 705 8091 753
rect 8019 659 8032 705
rect 8078 659 8091 705
rect 8019 611 8091 659
rect 8019 565 8032 611
rect 8078 565 8091 611
rect 8019 517 8091 565
rect 8019 471 8032 517
rect 8078 471 8091 517
rect 8019 423 8091 471
rect 8019 377 8032 423
rect 8078 377 8091 423
rect 8019 329 8091 377
rect 8019 283 8032 329
rect 8078 283 8091 329
rect 8019 235 8091 283
rect 5763 141 5835 189
rect 5763 95 5776 141
rect 5822 95 5835 141
rect 5763 47 5835 95
rect 5763 1 5776 47
rect 5822 1 5835 47
rect 5763 -47 5835 1
rect 5763 -93 5776 -47
rect 5822 -93 5835 -47
rect 8019 189 8032 235
rect 8078 189 8091 235
rect 10745 753 10758 799
rect 10804 753 10817 799
rect 10745 705 10817 753
rect 10745 659 10758 705
rect 10804 659 10817 705
rect 10745 611 10817 659
rect 10745 565 10758 611
rect 10804 565 10817 611
rect 10745 517 10817 565
rect 10745 471 10758 517
rect 10804 471 10817 517
rect 10745 423 10817 471
rect 10745 377 10758 423
rect 10804 377 10817 423
rect 10745 329 10817 377
rect 10745 283 10758 329
rect 10804 283 10817 329
rect 10745 235 10817 283
rect 8019 141 8091 189
rect 8019 95 8032 141
rect 8078 95 8091 141
rect 8019 47 8091 95
rect 8019 1 8032 47
rect 8078 1 8091 47
rect 8019 -47 8091 1
rect 5763 -141 5835 -93
rect 5763 -187 5776 -141
rect 5822 -187 5835 -141
rect 5763 -235 5835 -187
rect 5763 -281 5776 -235
rect 5822 -281 5835 -235
rect 5763 -329 5835 -281
rect 5763 -375 5776 -329
rect 5822 -375 5835 -329
rect 5763 -423 5835 -375
rect 5763 -469 5776 -423
rect 5822 -469 5835 -423
rect 5763 -517 5835 -469
rect 5763 -563 5776 -517
rect 5822 -563 5835 -517
rect 5763 -611 5835 -563
rect 5763 -657 5776 -611
rect 5822 -657 5835 -611
rect 8019 -93 8032 -47
rect 8078 -93 8091 -47
rect 10745 189 10758 235
rect 10804 189 10817 235
rect 10745 141 10817 189
rect 10745 95 10758 141
rect 10804 95 10817 141
rect 10745 47 10817 95
rect 10745 1 10758 47
rect 10804 1 10817 47
rect 10745 -47 10817 1
rect 8019 -141 8091 -93
rect 8019 -187 8032 -141
rect 8078 -187 8091 -141
rect 8019 -235 8091 -187
rect 8019 -281 8032 -235
rect 8078 -281 8091 -235
rect 8019 -329 8091 -281
rect 8019 -375 8032 -329
rect 8078 -375 8091 -329
rect 8019 -423 8091 -375
rect 8019 -469 8032 -423
rect 8078 -469 8091 -423
rect 8019 -517 8091 -469
rect 8019 -563 8032 -517
rect 8078 -563 8091 -517
rect 8019 -611 8091 -563
rect 5763 -705 5835 -657
rect 5763 -751 5776 -705
rect 5822 -751 5835 -705
rect 5763 -799 5835 -751
rect 5763 -845 5776 -799
rect 5822 -845 5835 -799
rect 8019 -657 8032 -611
rect 8078 -657 8091 -611
rect 10745 -93 10758 -47
rect 10804 -93 10817 -47
rect 10745 -141 10817 -93
rect 10745 -187 10758 -141
rect 10804 -187 10817 -141
rect 10745 -235 10817 -187
rect 10745 -281 10758 -235
rect 10804 -281 10817 -235
rect 10745 -329 10817 -281
rect 10745 -375 10758 -329
rect 10804 -375 10817 -329
rect 10745 -423 10817 -375
rect 10745 -469 10758 -423
rect 10804 -469 10817 -423
rect 10745 -517 10817 -469
rect 10745 -563 10758 -517
rect 10804 -563 10817 -517
rect 10745 -611 10817 -563
rect 8019 -705 8091 -657
rect 5763 -893 5835 -845
rect 5763 -939 5776 -893
rect 5822 -939 5835 -893
rect 8019 -751 8032 -705
rect 8078 -751 8091 -705
rect 8019 -799 8091 -751
rect 8019 -845 8032 -799
rect 8078 -845 8091 -799
rect 10745 -657 10758 -611
rect 10804 -657 10817 -611
rect 10745 -705 10817 -657
rect 10745 -751 10758 -705
rect 10804 -751 10817 -705
rect 8019 -893 8091 -845
rect 5763 -987 5835 -939
rect 5763 -1033 5776 -987
rect 5822 -1033 5835 -987
rect 5763 -1081 5835 -1033
rect 5763 -1127 5776 -1081
rect 5822 -1127 5835 -1081
rect 5763 -1175 5835 -1127
rect 5763 -1221 5776 -1175
rect 5822 -1221 5835 -1175
rect 5763 -1269 5835 -1221
rect 5763 -1315 5776 -1269
rect 5822 -1315 5835 -1269
rect 5763 -1363 5835 -1315
rect 5763 -1409 5776 -1363
rect 5822 -1409 5835 -1363
rect 5763 -1457 5835 -1409
rect 5763 -1503 5776 -1457
rect 5822 -1503 5835 -1457
rect 5763 -1551 5835 -1503
rect 5763 -1597 5776 -1551
rect 5822 -1597 5835 -1551
rect 5763 -1645 5835 -1597
rect 5763 -1691 5776 -1645
rect 5822 -1691 5835 -1645
rect 5763 -1739 5835 -1691
rect 5763 -1785 5776 -1739
rect 5822 -1785 5835 -1739
rect 5763 -1820 5835 -1785
rect 8019 -939 8032 -893
rect 8078 -939 8091 -893
rect 10745 -799 10817 -751
rect 10745 -845 10758 -799
rect 10804 -845 10817 -799
rect 10745 -893 10817 -845
rect 8019 -987 8091 -939
rect 8019 -1033 8032 -987
rect 8078 -1033 8091 -987
rect 8019 -1081 8091 -1033
rect 8019 -1127 8032 -1081
rect 8078 -1127 8091 -1081
rect 8019 -1175 8091 -1127
rect 8019 -1221 8032 -1175
rect 8078 -1221 8091 -1175
rect 8019 -1269 8091 -1221
rect 8019 -1315 8032 -1269
rect 8078 -1315 8091 -1269
rect 8019 -1363 8091 -1315
rect 8019 -1409 8032 -1363
rect 8078 -1409 8091 -1363
rect 8019 -1457 8091 -1409
rect 8019 -1503 8032 -1457
rect 8078 -1503 8091 -1457
rect 8019 -1551 8091 -1503
rect 8019 -1597 8032 -1551
rect 8078 -1597 8091 -1551
rect 8019 -1645 8091 -1597
rect 8019 -1691 8032 -1645
rect 8078 -1691 8091 -1645
rect 8019 -1739 8091 -1691
rect 8019 -1785 8032 -1739
rect 8078 -1785 8091 -1739
rect 8019 -1820 8091 -1785
rect 10745 -939 10758 -893
rect 10804 -939 10817 -893
rect 10745 -987 10817 -939
rect 10745 -1033 10758 -987
rect 10804 -1033 10817 -987
rect 10745 -1081 10817 -1033
rect 10745 -1127 10758 -1081
rect 10804 -1127 10817 -1081
rect 10745 -1175 10817 -1127
rect 10745 -1221 10758 -1175
rect 10804 -1221 10817 -1175
rect 10745 -1269 10817 -1221
rect 10745 -1315 10758 -1269
rect 10804 -1315 10817 -1269
rect 10745 -1363 10817 -1315
rect 10745 -1409 10758 -1363
rect 10804 -1409 10817 -1363
rect 10745 -1457 10817 -1409
rect 10745 -1503 10758 -1457
rect 10804 -1503 10817 -1457
rect 10745 -1551 10817 -1503
rect 10745 -1597 10758 -1551
rect 10804 -1597 10817 -1551
rect 10745 -1645 10817 -1597
rect 10745 -1691 10758 -1645
rect 10804 -1691 10817 -1645
rect 10745 -1739 10817 -1691
rect 10745 -1785 10758 -1739
rect 10804 -1785 10817 -1739
rect 10745 -1820 10817 -1785
rect 5763 -1833 10817 -1820
rect 5763 -1879 5776 -1833
rect 5822 -1879 5870 -1833
rect 5916 -1879 5964 -1833
rect 6010 -1879 6058 -1833
rect 6104 -1879 6152 -1833
rect 6198 -1879 6246 -1833
rect 6292 -1879 6340 -1833
rect 6386 -1879 6434 -1833
rect 6480 -1879 6528 -1833
rect 6574 -1879 6622 -1833
rect 6668 -1879 6716 -1833
rect 6762 -1879 6810 -1833
rect 6856 -1879 6904 -1833
rect 6950 -1879 6998 -1833
rect 7044 -1879 7092 -1833
rect 7138 -1879 7186 -1833
rect 7232 -1879 7280 -1833
rect 7326 -1879 7374 -1833
rect 7420 -1879 7468 -1833
rect 7514 -1879 7562 -1833
rect 7608 -1879 7656 -1833
rect 7702 -1879 7750 -1833
rect 7796 -1879 7844 -1833
rect 7890 -1879 7938 -1833
rect 7984 -1879 8032 -1833
rect 8078 -1879 8126 -1833
rect 8172 -1879 8220 -1833
rect 8266 -1879 8314 -1833
rect 8360 -1879 8408 -1833
rect 8454 -1879 8502 -1833
rect 8548 -1879 8596 -1833
rect 8642 -1879 8690 -1833
rect 8736 -1879 8784 -1833
rect 8830 -1879 8878 -1833
rect 8924 -1879 8972 -1833
rect 9018 -1879 9066 -1833
rect 9112 -1879 9160 -1833
rect 9206 -1879 9254 -1833
rect 9300 -1879 9348 -1833
rect 9394 -1879 9442 -1833
rect 9488 -1879 9536 -1833
rect 9582 -1879 9630 -1833
rect 9676 -1879 9724 -1833
rect 9770 -1879 9818 -1833
rect 9864 -1879 9912 -1833
rect 9958 -1879 10006 -1833
rect 10052 -1879 10100 -1833
rect 10146 -1879 10194 -1833
rect 10240 -1879 10288 -1833
rect 10334 -1879 10382 -1833
rect 10428 -1879 10476 -1833
rect 10522 -1879 10570 -1833
rect 10616 -1879 10664 -1833
rect 10710 -1879 10758 -1833
rect 10804 -1879 10817 -1833
rect 5763 -1892 10817 -1879
rect 17637 2591 17650 2637
rect 17696 2591 17709 2637
rect 17637 2543 17709 2591
rect 17637 2497 17650 2543
rect 17696 2497 17709 2543
rect 17637 2449 17709 2497
rect 17637 2403 17650 2449
rect 17696 2403 17709 2449
rect 17637 2355 17709 2403
rect 17637 2309 17650 2355
rect 17696 2309 17709 2355
rect 17637 2261 17709 2309
rect 17637 2215 17650 2261
rect 17696 2215 17709 2261
rect 17637 2167 17709 2215
rect 17637 2121 17650 2167
rect 17696 2121 17709 2167
rect 17637 2073 17709 2121
rect 17637 2027 17650 2073
rect 17696 2027 17709 2073
rect 17637 1979 17709 2027
rect 17637 1933 17650 1979
rect 17696 1933 17709 1979
rect 17637 1885 17709 1933
rect 17637 1839 17650 1885
rect 17696 1839 17709 1885
rect 17637 1791 17709 1839
rect 17637 1745 17650 1791
rect 17696 1745 17709 1791
rect 17637 1697 17709 1745
rect 17637 1651 17650 1697
rect 17696 1651 17709 1697
rect 17637 1603 17709 1651
rect 17637 1557 17650 1603
rect 17696 1557 17709 1603
rect 17637 1509 17709 1557
rect 17637 1463 17650 1509
rect 17696 1463 17709 1509
rect 17637 1415 17709 1463
rect 17637 1369 17650 1415
rect 17696 1369 17709 1415
rect 17637 1321 17709 1369
rect 17637 1275 17650 1321
rect 17696 1275 17709 1321
rect 17637 1227 17709 1275
rect 17637 1181 17650 1227
rect 17696 1181 17709 1227
rect 17637 1133 17709 1181
rect 17637 1087 17650 1133
rect 17696 1087 17709 1133
rect 17637 1039 17709 1087
rect 17637 993 17650 1039
rect 17696 993 17709 1039
rect 17637 945 17709 993
rect 17637 899 17650 945
rect 17696 899 17709 945
rect 17637 851 17709 899
rect 17637 805 17650 851
rect 17696 805 17709 851
rect 17637 757 17709 805
rect 17637 711 17650 757
rect 17696 711 17709 757
rect 17637 663 17709 711
rect 17637 617 17650 663
rect 17696 617 17709 663
rect 17637 569 17709 617
rect 17637 523 17650 569
rect 17696 523 17709 569
rect 17637 475 17709 523
rect 17637 429 17650 475
rect 17696 429 17709 475
rect 17637 381 17709 429
rect 17637 335 17650 381
rect 17696 335 17709 381
rect 17637 287 17709 335
rect 17637 241 17650 287
rect 17696 241 17709 287
rect 17637 193 17709 241
rect 17637 147 17650 193
rect 17696 147 17709 193
rect 17637 99 17709 147
rect 17637 53 17650 99
rect 17696 53 17709 99
rect 17637 5 17709 53
rect 17637 -41 17650 5
rect 17696 -41 17709 5
rect 17637 -89 17709 -41
rect 17637 -135 17650 -89
rect 17696 -135 17709 -89
rect 17637 -183 17709 -135
rect 17637 -229 17650 -183
rect 17696 -229 17709 -183
rect 17637 -277 17709 -229
rect 17637 -323 17650 -277
rect 17696 -323 17709 -277
rect 17637 -371 17709 -323
rect 17637 -417 17650 -371
rect 17696 -417 17709 -371
rect 17637 -465 17709 -417
rect 20645 3295 20717 3343
rect 20645 3249 20658 3295
rect 20704 3249 20717 3295
rect 17637 -511 17650 -465
rect 17696 -511 17709 -465
rect 17637 -559 17709 -511
rect 20645 3201 20717 3249
rect 20645 3155 20658 3201
rect 20704 3155 20717 3201
rect 20645 3107 20717 3155
rect 20645 3061 20658 3107
rect 20704 3061 20717 3107
rect 20645 3013 20717 3061
rect 20645 2967 20658 3013
rect 20704 2967 20717 3013
rect 20645 2919 20717 2967
rect 20645 2873 20658 2919
rect 20704 2873 20717 2919
rect 20645 2825 20717 2873
rect 20645 2779 20658 2825
rect 20704 2779 20717 2825
rect 20645 2731 20717 2779
rect 20645 2685 20658 2731
rect 20704 2685 20717 2731
rect 20645 2637 20717 2685
rect 20645 2591 20658 2637
rect 20704 2591 20717 2637
rect 20645 2543 20717 2591
rect 20645 2497 20658 2543
rect 20704 2497 20717 2543
rect 20645 2449 20717 2497
rect 20645 2403 20658 2449
rect 20704 2403 20717 2449
rect 20645 2355 20717 2403
rect 20645 2309 20658 2355
rect 20704 2309 20717 2355
rect 20645 2261 20717 2309
rect 20645 2215 20658 2261
rect 20704 2215 20717 2261
rect 20645 2167 20717 2215
rect 20645 2121 20658 2167
rect 20704 2121 20717 2167
rect 20645 2073 20717 2121
rect 20645 2027 20658 2073
rect 20704 2027 20717 2073
rect 20645 1979 20717 2027
rect 20645 1933 20658 1979
rect 20704 1933 20717 1979
rect 20645 1885 20717 1933
rect 20645 1839 20658 1885
rect 20704 1839 20717 1885
rect 20645 1791 20717 1839
rect 20645 1745 20658 1791
rect 20704 1745 20717 1791
rect 20645 1697 20717 1745
rect 20645 1651 20658 1697
rect 20704 1651 20717 1697
rect 20645 1603 20717 1651
rect 20645 1557 20658 1603
rect 20704 1557 20717 1603
rect 20645 1509 20717 1557
rect 20645 1463 20658 1509
rect 20704 1463 20717 1509
rect 20645 1415 20717 1463
rect 20645 1369 20658 1415
rect 20704 1369 20717 1415
rect 20645 1321 20717 1369
rect 20645 1275 20658 1321
rect 20704 1275 20717 1321
rect 20645 1227 20717 1275
rect 20645 1181 20658 1227
rect 20704 1181 20717 1227
rect 20645 1133 20717 1181
rect 20645 1087 20658 1133
rect 20704 1087 20717 1133
rect 20645 1039 20717 1087
rect 20645 993 20658 1039
rect 20704 993 20717 1039
rect 20645 945 20717 993
rect 20645 899 20658 945
rect 20704 899 20717 945
rect 20645 851 20717 899
rect 20645 805 20658 851
rect 20704 805 20717 851
rect 20645 757 20717 805
rect 20645 711 20658 757
rect 20704 711 20717 757
rect 20645 663 20717 711
rect 20645 617 20658 663
rect 20704 617 20717 663
rect 20645 569 20717 617
rect 20645 523 20658 569
rect 20704 523 20717 569
rect 20645 475 20717 523
rect 20645 429 20658 475
rect 20704 429 20717 475
rect 20645 381 20717 429
rect 20645 335 20658 381
rect 20704 335 20717 381
rect 20645 287 20717 335
rect 20645 241 20658 287
rect 20704 241 20717 287
rect 20645 193 20717 241
rect 20645 147 20658 193
rect 20704 147 20717 193
rect 20645 99 20717 147
rect 20645 53 20658 99
rect 20704 53 20717 99
rect 20645 5 20717 53
rect 20645 -41 20658 5
rect 20704 -41 20717 5
rect 20645 -89 20717 -41
rect 20645 -135 20658 -89
rect 20704 -135 20717 -89
rect 20645 -183 20717 -135
rect 20645 -229 20658 -183
rect 20704 -229 20717 -183
rect 20645 -277 20717 -229
rect 20645 -323 20658 -277
rect 20704 -323 20717 -277
rect 20645 -371 20717 -323
rect 20645 -417 20658 -371
rect 20704 -417 20717 -371
rect 17637 -605 17650 -559
rect 17696 -605 17709 -559
rect 17637 -653 17709 -605
rect 20645 -465 20717 -417
rect 20645 -511 20658 -465
rect 20704 -511 20717 -465
rect 20645 -559 20717 -511
rect 20645 -605 20658 -559
rect 20704 -605 20717 -559
rect 17637 -699 17650 -653
rect 17696 -699 17709 -653
rect 17637 -747 17709 -699
rect 17637 -793 17650 -747
rect 17696 -793 17709 -747
rect 17637 -841 17709 -793
rect 17637 -887 17650 -841
rect 17696 -887 17709 -841
rect 17637 -935 17709 -887
rect 17637 -981 17650 -935
rect 17696 -981 17709 -935
rect 17637 -1029 17709 -981
rect 17637 -1075 17650 -1029
rect 17696 -1075 17709 -1029
rect 17637 -1123 17709 -1075
rect 17637 -1169 17650 -1123
rect 17696 -1169 17709 -1123
rect 17637 -1217 17709 -1169
rect 17637 -1263 17650 -1217
rect 17696 -1263 17709 -1217
rect 20645 -653 20717 -605
rect 20645 -699 20658 -653
rect 20704 -699 20717 -653
rect 20645 -747 20717 -699
rect 20645 -793 20658 -747
rect 20704 -793 20717 -747
rect 20645 -841 20717 -793
rect 20645 -887 20658 -841
rect 20704 -887 20717 -841
rect 20645 -935 20717 -887
rect 20645 -981 20658 -935
rect 20704 -981 20717 -935
rect 20645 -1029 20717 -981
rect 20645 -1075 20658 -1029
rect 20704 -1075 20717 -1029
rect 20645 -1123 20717 -1075
rect 20645 -1169 20658 -1123
rect 20704 -1169 20717 -1123
rect 20645 -1217 20717 -1169
rect 17637 -1311 17709 -1263
rect 17637 -1357 17650 -1311
rect 17696 -1357 17709 -1311
rect 17637 -1405 17709 -1357
rect 20645 -1263 20658 -1217
rect 20704 -1263 20717 -1217
rect 20645 -1311 20717 -1263
rect 20645 -1357 20658 -1311
rect 20704 -1357 20717 -1311
rect 17637 -1451 17650 -1405
rect 17696 -1451 17709 -1405
rect 17637 -1499 17709 -1451
rect 20645 -1405 20717 -1357
rect 20645 -1451 20658 -1405
rect 20704 -1451 20717 -1405
rect 17637 -1545 17650 -1499
rect 17696 -1545 17709 -1499
rect 17637 -1593 17709 -1545
rect 17637 -1639 17650 -1593
rect 17696 -1639 17709 -1593
rect 17637 -1687 17709 -1639
rect 17637 -1733 17650 -1687
rect 17696 -1733 17709 -1687
rect 17637 -1768 17709 -1733
rect 20645 -1499 20717 -1451
rect 20645 -1545 20658 -1499
rect 20704 -1545 20717 -1499
rect 20645 -1593 20717 -1545
rect 20645 -1639 20658 -1593
rect 20704 -1639 20717 -1593
rect 20645 -1687 20717 -1639
rect 20645 -1733 20658 -1687
rect 20704 -1733 20717 -1687
rect 20645 -1768 20717 -1733
rect 17637 -1781 20717 -1768
rect 17637 -1827 17650 -1781
rect 17696 -1827 17744 -1781
rect 17790 -1827 17838 -1781
rect 17884 -1827 17932 -1781
rect 17978 -1827 18026 -1781
rect 18072 -1827 18120 -1781
rect 18166 -1827 18214 -1781
rect 18260 -1827 18308 -1781
rect 18354 -1827 18402 -1781
rect 18448 -1827 18496 -1781
rect 18542 -1827 18590 -1781
rect 18636 -1827 18684 -1781
rect 18730 -1827 18778 -1781
rect 18824 -1827 18872 -1781
rect 18918 -1827 18966 -1781
rect 19012 -1827 19060 -1781
rect 19106 -1827 19154 -1781
rect 19200 -1827 19248 -1781
rect 19294 -1827 19342 -1781
rect 19388 -1827 19436 -1781
rect 19482 -1827 19530 -1781
rect 19576 -1827 19624 -1781
rect 19670 -1827 19718 -1781
rect 19764 -1827 19812 -1781
rect 19858 -1827 19906 -1781
rect 19952 -1827 20000 -1781
rect 20046 -1827 20094 -1781
rect 20140 -1827 20188 -1781
rect 20234 -1827 20282 -1781
rect 20328 -1827 20376 -1781
rect 20422 -1827 20470 -1781
rect 20516 -1827 20564 -1781
rect 20610 -1827 20658 -1781
rect 20704 -1827 20717 -1781
rect 17637 -1840 20717 -1827
rect 22789 4611 25869 4624
rect 22789 4565 22802 4611
rect 22848 4565 22896 4611
rect 22942 4565 22990 4611
rect 23036 4565 23084 4611
rect 23130 4565 23178 4611
rect 23224 4565 23272 4611
rect 23318 4565 23366 4611
rect 23412 4565 23460 4611
rect 23506 4565 23554 4611
rect 23600 4565 23648 4611
rect 23694 4565 23742 4611
rect 23788 4565 23836 4611
rect 23882 4565 23930 4611
rect 23976 4565 24024 4611
rect 24070 4565 24118 4611
rect 24164 4565 24212 4611
rect 24258 4565 24306 4611
rect 24352 4565 24400 4611
rect 24446 4565 24494 4611
rect 24540 4565 24588 4611
rect 24634 4565 24682 4611
rect 24728 4565 24776 4611
rect 24822 4565 24870 4611
rect 24916 4565 24964 4611
rect 25010 4565 25058 4611
rect 25104 4565 25152 4611
rect 25198 4565 25246 4611
rect 25292 4565 25340 4611
rect 25386 4565 25434 4611
rect 25480 4565 25528 4611
rect 25574 4565 25622 4611
rect 25668 4565 25716 4611
rect 25762 4565 25810 4611
rect 25856 4565 25869 4611
rect 22789 4552 25869 4565
rect 22789 4517 22861 4552
rect 22789 4471 22802 4517
rect 22848 4471 22861 4517
rect 22789 4423 22861 4471
rect 22789 4377 22802 4423
rect 22848 4377 22861 4423
rect 22789 4329 22861 4377
rect 22789 4283 22802 4329
rect 22848 4283 22861 4329
rect 22789 4235 22861 4283
rect 25797 4517 25869 4552
rect 25797 4471 25810 4517
rect 25856 4471 25869 4517
rect 25797 4423 25869 4471
rect 25797 4377 25810 4423
rect 25856 4377 25869 4423
rect 25797 4329 25869 4377
rect 25797 4283 25810 4329
rect 25856 4283 25869 4329
rect 22789 4189 22802 4235
rect 22848 4189 22861 4235
rect 22789 4141 22861 4189
rect 25797 4235 25869 4283
rect 25797 4189 25810 4235
rect 25856 4189 25869 4235
rect 22789 4095 22802 4141
rect 22848 4095 22861 4141
rect 22789 4047 22861 4095
rect 22789 4001 22802 4047
rect 22848 4001 22861 4047
rect 25797 4141 25869 4189
rect 25797 4095 25810 4141
rect 25856 4095 25869 4141
rect 25797 4047 25869 4095
rect 22789 3953 22861 4001
rect 22789 3907 22802 3953
rect 22848 3907 22861 3953
rect 22789 3859 22861 3907
rect 22789 3813 22802 3859
rect 22848 3813 22861 3859
rect 22789 3765 22861 3813
rect 22789 3719 22802 3765
rect 22848 3719 22861 3765
rect 22789 3671 22861 3719
rect 22789 3625 22802 3671
rect 22848 3625 22861 3671
rect 22789 3577 22861 3625
rect 22789 3531 22802 3577
rect 22848 3531 22861 3577
rect 22789 3483 22861 3531
rect 22789 3437 22802 3483
rect 22848 3437 22861 3483
rect 22789 3389 22861 3437
rect 25797 4001 25810 4047
rect 25856 4001 25869 4047
rect 25797 3953 25869 4001
rect 25797 3907 25810 3953
rect 25856 3907 25869 3953
rect 25797 3859 25869 3907
rect 25797 3813 25810 3859
rect 25856 3813 25869 3859
rect 25797 3765 25869 3813
rect 25797 3719 25810 3765
rect 25856 3719 25869 3765
rect 25797 3671 25869 3719
rect 25797 3625 25810 3671
rect 25856 3625 25869 3671
rect 25797 3577 25869 3625
rect 25797 3531 25810 3577
rect 25856 3531 25869 3577
rect 25797 3483 25869 3531
rect 25797 3437 25810 3483
rect 25856 3437 25869 3483
rect 22789 3343 22802 3389
rect 22848 3343 22861 3389
rect 22789 3295 22861 3343
rect 22789 3249 22802 3295
rect 22848 3249 22861 3295
rect 22789 3201 22861 3249
rect 25797 3389 25869 3437
rect 25797 3343 25810 3389
rect 25856 3343 25869 3389
rect 22789 3155 22802 3201
rect 22848 3155 22861 3201
rect 22789 3107 22861 3155
rect 22789 3061 22802 3107
rect 22848 3061 22861 3107
rect 22789 3013 22861 3061
rect 22789 2967 22802 3013
rect 22848 2967 22861 3013
rect 22789 2919 22861 2967
rect 22789 2873 22802 2919
rect 22848 2873 22861 2919
rect 22789 2825 22861 2873
rect 22789 2779 22802 2825
rect 22848 2779 22861 2825
rect 22789 2731 22861 2779
rect 22789 2685 22802 2731
rect 22848 2685 22861 2731
rect 22789 2637 22861 2685
rect 22789 2591 22802 2637
rect 22848 2591 22861 2637
rect 22789 2543 22861 2591
rect 22789 2497 22802 2543
rect 22848 2497 22861 2543
rect 22789 2449 22861 2497
rect 22789 2403 22802 2449
rect 22848 2403 22861 2449
rect 22789 2355 22861 2403
rect 22789 2309 22802 2355
rect 22848 2309 22861 2355
rect 22789 2261 22861 2309
rect 22789 2215 22802 2261
rect 22848 2215 22861 2261
rect 22789 2167 22861 2215
rect 22789 2121 22802 2167
rect 22848 2121 22861 2167
rect 22789 2073 22861 2121
rect 22789 2027 22802 2073
rect 22848 2027 22861 2073
rect 22789 1979 22861 2027
rect 22789 1933 22802 1979
rect 22848 1933 22861 1979
rect 22789 1885 22861 1933
rect 22789 1839 22802 1885
rect 22848 1839 22861 1885
rect 22789 1791 22861 1839
rect 22789 1745 22802 1791
rect 22848 1745 22861 1791
rect 22789 1697 22861 1745
rect 22789 1651 22802 1697
rect 22848 1651 22861 1697
rect 22789 1603 22861 1651
rect 22789 1557 22802 1603
rect 22848 1557 22861 1603
rect 22789 1509 22861 1557
rect 22789 1463 22802 1509
rect 22848 1463 22861 1509
rect 22789 1415 22861 1463
rect 22789 1369 22802 1415
rect 22848 1369 22861 1415
rect 22789 1321 22861 1369
rect 22789 1275 22802 1321
rect 22848 1275 22861 1321
rect 22789 1227 22861 1275
rect 22789 1181 22802 1227
rect 22848 1181 22861 1227
rect 22789 1133 22861 1181
rect 22789 1087 22802 1133
rect 22848 1087 22861 1133
rect 22789 1039 22861 1087
rect 22789 993 22802 1039
rect 22848 993 22861 1039
rect 22789 945 22861 993
rect 22789 899 22802 945
rect 22848 899 22861 945
rect 22789 851 22861 899
rect 22789 805 22802 851
rect 22848 805 22861 851
rect 22789 757 22861 805
rect 22789 711 22802 757
rect 22848 711 22861 757
rect 22789 663 22861 711
rect 22789 617 22802 663
rect 22848 617 22861 663
rect 22789 569 22861 617
rect 22789 523 22802 569
rect 22848 523 22861 569
rect 22789 475 22861 523
rect 22789 429 22802 475
rect 22848 429 22861 475
rect 22789 381 22861 429
rect 22789 335 22802 381
rect 22848 335 22861 381
rect 22789 287 22861 335
rect 22789 241 22802 287
rect 22848 241 22861 287
rect 22789 193 22861 241
rect 22789 147 22802 193
rect 22848 147 22861 193
rect 22789 99 22861 147
rect 22789 53 22802 99
rect 22848 53 22861 99
rect 22789 5 22861 53
rect 22789 -41 22802 5
rect 22848 -41 22861 5
rect 22789 -89 22861 -41
rect 22789 -135 22802 -89
rect 22848 -135 22861 -89
rect 22789 -183 22861 -135
rect 22789 -229 22802 -183
rect 22848 -229 22861 -183
rect 22789 -277 22861 -229
rect 22789 -323 22802 -277
rect 22848 -323 22861 -277
rect 22789 -371 22861 -323
rect 22789 -417 22802 -371
rect 22848 -417 22861 -371
rect 22789 -465 22861 -417
rect 25797 3295 25869 3343
rect 25797 3249 25810 3295
rect 25856 3249 25869 3295
rect 22789 -511 22802 -465
rect 22848 -511 22861 -465
rect 22789 -559 22861 -511
rect 25797 3201 25869 3249
rect 25797 3155 25810 3201
rect 25856 3155 25869 3201
rect 25797 3107 25869 3155
rect 25797 3061 25810 3107
rect 25856 3061 25869 3107
rect 25797 3013 25869 3061
rect 25797 2967 25810 3013
rect 25856 2967 25869 3013
rect 25797 2919 25869 2967
rect 25797 2873 25810 2919
rect 25856 2873 25869 2919
rect 25797 2825 25869 2873
rect 25797 2779 25810 2825
rect 25856 2779 25869 2825
rect 25797 2731 25869 2779
rect 25797 2685 25810 2731
rect 25856 2685 25869 2731
rect 25797 2637 25869 2685
rect 25797 2591 25810 2637
rect 25856 2591 25869 2637
rect 25797 2543 25869 2591
rect 25797 2497 25810 2543
rect 25856 2497 25869 2543
rect 25797 2449 25869 2497
rect 25797 2403 25810 2449
rect 25856 2403 25869 2449
rect 25797 2355 25869 2403
rect 25797 2309 25810 2355
rect 25856 2309 25869 2355
rect 25797 2261 25869 2309
rect 25797 2215 25810 2261
rect 25856 2215 25869 2261
rect 25797 2167 25869 2215
rect 25797 2121 25810 2167
rect 25856 2121 25869 2167
rect 25797 2073 25869 2121
rect 25797 2027 25810 2073
rect 25856 2027 25869 2073
rect 25797 1979 25869 2027
rect 25797 1933 25810 1979
rect 25856 1933 25869 1979
rect 25797 1885 25869 1933
rect 25797 1839 25810 1885
rect 25856 1839 25869 1885
rect 25797 1791 25869 1839
rect 25797 1745 25810 1791
rect 25856 1745 25869 1791
rect 25797 1697 25869 1745
rect 25797 1651 25810 1697
rect 25856 1651 25869 1697
rect 25797 1603 25869 1651
rect 25797 1557 25810 1603
rect 25856 1557 25869 1603
rect 25797 1509 25869 1557
rect 25797 1463 25810 1509
rect 25856 1463 25869 1509
rect 25797 1415 25869 1463
rect 25797 1369 25810 1415
rect 25856 1369 25869 1415
rect 25797 1321 25869 1369
rect 25797 1275 25810 1321
rect 25856 1275 25869 1321
rect 25797 1227 25869 1275
rect 25797 1181 25810 1227
rect 25856 1181 25869 1227
rect 25797 1133 25869 1181
rect 25797 1087 25810 1133
rect 25856 1087 25869 1133
rect 25797 1039 25869 1087
rect 25797 993 25810 1039
rect 25856 993 25869 1039
rect 25797 945 25869 993
rect 25797 899 25810 945
rect 25856 899 25869 945
rect 25797 851 25869 899
rect 25797 805 25810 851
rect 25856 805 25869 851
rect 25797 757 25869 805
rect 25797 711 25810 757
rect 25856 711 25869 757
rect 25797 663 25869 711
rect 25797 617 25810 663
rect 25856 617 25869 663
rect 25797 569 25869 617
rect 25797 523 25810 569
rect 25856 523 25869 569
rect 25797 475 25869 523
rect 25797 429 25810 475
rect 25856 429 25869 475
rect 25797 381 25869 429
rect 25797 335 25810 381
rect 25856 335 25869 381
rect 25797 287 25869 335
rect 25797 241 25810 287
rect 25856 241 25869 287
rect 25797 193 25869 241
rect 25797 147 25810 193
rect 25856 147 25869 193
rect 25797 99 25869 147
rect 25797 53 25810 99
rect 25856 53 25869 99
rect 25797 5 25869 53
rect 25797 -41 25810 5
rect 25856 -41 25869 5
rect 25797 -89 25869 -41
rect 25797 -135 25810 -89
rect 25856 -135 25869 -89
rect 25797 -183 25869 -135
rect 25797 -229 25810 -183
rect 25856 -229 25869 -183
rect 25797 -277 25869 -229
rect 25797 -323 25810 -277
rect 25856 -323 25869 -277
rect 25797 -371 25869 -323
rect 25797 -417 25810 -371
rect 25856 -417 25869 -371
rect 22789 -605 22802 -559
rect 22848 -605 22861 -559
rect 22789 -653 22861 -605
rect 25797 -465 25869 -417
rect 25797 -511 25810 -465
rect 25856 -511 25869 -465
rect 25797 -559 25869 -511
rect 25797 -605 25810 -559
rect 25856 -605 25869 -559
rect 22789 -699 22802 -653
rect 22848 -699 22861 -653
rect 22789 -747 22861 -699
rect 22789 -793 22802 -747
rect 22848 -793 22861 -747
rect 22789 -841 22861 -793
rect 22789 -887 22802 -841
rect 22848 -887 22861 -841
rect 22789 -935 22861 -887
rect 22789 -981 22802 -935
rect 22848 -981 22861 -935
rect 22789 -1029 22861 -981
rect 22789 -1075 22802 -1029
rect 22848 -1075 22861 -1029
rect 22789 -1123 22861 -1075
rect 22789 -1169 22802 -1123
rect 22848 -1169 22861 -1123
rect 22789 -1217 22861 -1169
rect 22789 -1263 22802 -1217
rect 22848 -1263 22861 -1217
rect 25797 -653 25869 -605
rect 25797 -699 25810 -653
rect 25856 -699 25869 -653
rect 25797 -747 25869 -699
rect 25797 -793 25810 -747
rect 25856 -793 25869 -747
rect 25797 -841 25869 -793
rect 25797 -887 25810 -841
rect 25856 -887 25869 -841
rect 25797 -935 25869 -887
rect 25797 -981 25810 -935
rect 25856 -981 25869 -935
rect 25797 -1029 25869 -981
rect 25797 -1075 25810 -1029
rect 25856 -1075 25869 -1029
rect 25797 -1123 25869 -1075
rect 25797 -1169 25810 -1123
rect 25856 -1169 25869 -1123
rect 25797 -1217 25869 -1169
rect 22789 -1311 22861 -1263
rect 22789 -1357 22802 -1311
rect 22848 -1357 22861 -1311
rect 22789 -1405 22861 -1357
rect 25797 -1263 25810 -1217
rect 25856 -1263 25869 -1217
rect 25797 -1311 25869 -1263
rect 25797 -1357 25810 -1311
rect 25856 -1357 25869 -1311
rect 22789 -1451 22802 -1405
rect 22848 -1451 22861 -1405
rect 22789 -1499 22861 -1451
rect 25797 -1405 25869 -1357
rect 25797 -1451 25810 -1405
rect 25856 -1451 25869 -1405
rect 22789 -1545 22802 -1499
rect 22848 -1545 22861 -1499
rect 22789 -1593 22861 -1545
rect 22789 -1639 22802 -1593
rect 22848 -1639 22861 -1593
rect 22789 -1687 22861 -1639
rect 22789 -1733 22802 -1687
rect 22848 -1733 22861 -1687
rect 22789 -1768 22861 -1733
rect 25797 -1499 25869 -1451
rect 25797 -1545 25810 -1499
rect 25856 -1545 25869 -1499
rect 25797 -1593 25869 -1545
rect 25797 -1639 25810 -1593
rect 25856 -1639 25869 -1593
rect 25797 -1687 25869 -1639
rect 25797 -1733 25810 -1687
rect 25856 -1733 25869 -1687
rect 25797 -1768 25869 -1733
rect 22789 -1781 25869 -1768
rect 22789 -1827 22802 -1781
rect 22848 -1827 22896 -1781
rect 22942 -1827 22990 -1781
rect 23036 -1827 23084 -1781
rect 23130 -1827 23178 -1781
rect 23224 -1827 23272 -1781
rect 23318 -1827 23366 -1781
rect 23412 -1827 23460 -1781
rect 23506 -1827 23554 -1781
rect 23600 -1827 23648 -1781
rect 23694 -1827 23742 -1781
rect 23788 -1827 23836 -1781
rect 23882 -1827 23930 -1781
rect 23976 -1827 24024 -1781
rect 24070 -1827 24118 -1781
rect 24164 -1827 24212 -1781
rect 24258 -1827 24306 -1781
rect 24352 -1827 24400 -1781
rect 24446 -1827 24494 -1781
rect 24540 -1827 24588 -1781
rect 24634 -1827 24682 -1781
rect 24728 -1827 24776 -1781
rect 24822 -1827 24870 -1781
rect 24916 -1827 24964 -1781
rect 25010 -1827 25058 -1781
rect 25104 -1827 25152 -1781
rect 25198 -1827 25246 -1781
rect 25292 -1827 25340 -1781
rect 25386 -1827 25434 -1781
rect 25480 -1827 25528 -1781
rect 25574 -1827 25622 -1781
rect 25668 -1827 25716 -1781
rect 25762 -1827 25810 -1781
rect 25856 -1827 25869 -1781
rect 22789 -1840 25869 -1827
rect 26758 4611 29838 4624
rect 26758 4565 26771 4611
rect 26817 4565 26865 4611
rect 26911 4565 26959 4611
rect 27005 4565 27053 4611
rect 27099 4565 27147 4611
rect 27193 4565 27241 4611
rect 27287 4565 27335 4611
rect 27381 4565 27429 4611
rect 27475 4565 27523 4611
rect 27569 4565 27617 4611
rect 27663 4565 27711 4611
rect 27757 4565 27805 4611
rect 27851 4565 27899 4611
rect 27945 4565 27993 4611
rect 28039 4565 28087 4611
rect 28133 4565 28181 4611
rect 28227 4565 28275 4611
rect 28321 4565 28369 4611
rect 28415 4565 28463 4611
rect 28509 4565 28557 4611
rect 28603 4565 28651 4611
rect 28697 4565 28745 4611
rect 28791 4565 28839 4611
rect 28885 4565 28933 4611
rect 28979 4565 29027 4611
rect 29073 4565 29121 4611
rect 29167 4565 29215 4611
rect 29261 4565 29309 4611
rect 29355 4565 29403 4611
rect 29449 4565 29497 4611
rect 29543 4565 29591 4611
rect 29637 4565 29685 4611
rect 29731 4565 29779 4611
rect 29825 4565 29838 4611
rect 26758 4552 29838 4565
rect 26758 4517 26830 4552
rect 26758 4471 26771 4517
rect 26817 4471 26830 4517
rect 26758 4423 26830 4471
rect 26758 4377 26771 4423
rect 26817 4377 26830 4423
rect 26758 4329 26830 4377
rect 26758 4283 26771 4329
rect 26817 4283 26830 4329
rect 26758 4235 26830 4283
rect 29766 4517 29838 4552
rect 29766 4471 29779 4517
rect 29825 4471 29838 4517
rect 29766 4423 29838 4471
rect 29766 4377 29779 4423
rect 29825 4377 29838 4423
rect 29766 4329 29838 4377
rect 29766 4283 29779 4329
rect 29825 4283 29838 4329
rect 26758 4189 26771 4235
rect 26817 4189 26830 4235
rect 26758 4141 26830 4189
rect 29766 4235 29838 4283
rect 29766 4189 29779 4235
rect 29825 4189 29838 4235
rect 26758 4095 26771 4141
rect 26817 4095 26830 4141
rect 26758 4047 26830 4095
rect 26758 4001 26771 4047
rect 26817 4001 26830 4047
rect 29766 4141 29838 4189
rect 29766 4095 29779 4141
rect 29825 4095 29838 4141
rect 29766 4047 29838 4095
rect 26758 3953 26830 4001
rect 26758 3907 26771 3953
rect 26817 3907 26830 3953
rect 26758 3859 26830 3907
rect 26758 3813 26771 3859
rect 26817 3813 26830 3859
rect 26758 3765 26830 3813
rect 26758 3719 26771 3765
rect 26817 3719 26830 3765
rect 26758 3671 26830 3719
rect 26758 3625 26771 3671
rect 26817 3625 26830 3671
rect 26758 3577 26830 3625
rect 26758 3531 26771 3577
rect 26817 3531 26830 3577
rect 26758 3483 26830 3531
rect 26758 3437 26771 3483
rect 26817 3437 26830 3483
rect 26758 3389 26830 3437
rect 29766 4001 29779 4047
rect 29825 4001 29838 4047
rect 29766 3953 29838 4001
rect 29766 3907 29779 3953
rect 29825 3907 29838 3953
rect 29766 3859 29838 3907
rect 29766 3813 29779 3859
rect 29825 3813 29838 3859
rect 29766 3765 29838 3813
rect 29766 3719 29779 3765
rect 29825 3719 29838 3765
rect 29766 3671 29838 3719
rect 29766 3625 29779 3671
rect 29825 3625 29838 3671
rect 29766 3577 29838 3625
rect 29766 3531 29779 3577
rect 29825 3531 29838 3577
rect 29766 3483 29838 3531
rect 29766 3437 29779 3483
rect 29825 3437 29838 3483
rect 26758 3343 26771 3389
rect 26817 3343 26830 3389
rect 26758 3295 26830 3343
rect 26758 3249 26771 3295
rect 26817 3249 26830 3295
rect 26758 3201 26830 3249
rect 29766 3389 29838 3437
rect 29766 3343 29779 3389
rect 29825 3343 29838 3389
rect 26758 3155 26771 3201
rect 26817 3155 26830 3201
rect 26758 3107 26830 3155
rect 26758 3061 26771 3107
rect 26817 3061 26830 3107
rect 26758 3013 26830 3061
rect 26758 2967 26771 3013
rect 26817 2967 26830 3013
rect 26758 2919 26830 2967
rect 26758 2873 26771 2919
rect 26817 2873 26830 2919
rect 26758 2825 26830 2873
rect 26758 2779 26771 2825
rect 26817 2779 26830 2825
rect 26758 2731 26830 2779
rect 26758 2685 26771 2731
rect 26817 2685 26830 2731
rect 26758 2637 26830 2685
rect 26758 2591 26771 2637
rect 26817 2591 26830 2637
rect 26758 2543 26830 2591
rect 26758 2497 26771 2543
rect 26817 2497 26830 2543
rect 26758 2449 26830 2497
rect 26758 2403 26771 2449
rect 26817 2403 26830 2449
rect 26758 2355 26830 2403
rect 26758 2309 26771 2355
rect 26817 2309 26830 2355
rect 26758 2261 26830 2309
rect 26758 2215 26771 2261
rect 26817 2215 26830 2261
rect 26758 2167 26830 2215
rect 26758 2121 26771 2167
rect 26817 2121 26830 2167
rect 26758 2073 26830 2121
rect 26758 2027 26771 2073
rect 26817 2027 26830 2073
rect 26758 1979 26830 2027
rect 26758 1933 26771 1979
rect 26817 1933 26830 1979
rect 26758 1885 26830 1933
rect 26758 1839 26771 1885
rect 26817 1839 26830 1885
rect 26758 1791 26830 1839
rect 26758 1745 26771 1791
rect 26817 1745 26830 1791
rect 26758 1697 26830 1745
rect 26758 1651 26771 1697
rect 26817 1651 26830 1697
rect 26758 1603 26830 1651
rect 26758 1557 26771 1603
rect 26817 1557 26830 1603
rect 26758 1509 26830 1557
rect 26758 1463 26771 1509
rect 26817 1463 26830 1509
rect 26758 1415 26830 1463
rect 26758 1369 26771 1415
rect 26817 1369 26830 1415
rect 26758 1321 26830 1369
rect 26758 1275 26771 1321
rect 26817 1275 26830 1321
rect 26758 1227 26830 1275
rect 26758 1181 26771 1227
rect 26817 1181 26830 1227
rect 26758 1133 26830 1181
rect 26758 1087 26771 1133
rect 26817 1087 26830 1133
rect 26758 1039 26830 1087
rect 26758 993 26771 1039
rect 26817 993 26830 1039
rect 26758 945 26830 993
rect 26758 899 26771 945
rect 26817 899 26830 945
rect 26758 851 26830 899
rect 26758 805 26771 851
rect 26817 805 26830 851
rect 26758 757 26830 805
rect 26758 711 26771 757
rect 26817 711 26830 757
rect 26758 663 26830 711
rect 26758 617 26771 663
rect 26817 617 26830 663
rect 26758 569 26830 617
rect 26758 523 26771 569
rect 26817 523 26830 569
rect 26758 475 26830 523
rect 26758 429 26771 475
rect 26817 429 26830 475
rect 26758 381 26830 429
rect 26758 335 26771 381
rect 26817 335 26830 381
rect 26758 287 26830 335
rect 26758 241 26771 287
rect 26817 241 26830 287
rect 26758 193 26830 241
rect 26758 147 26771 193
rect 26817 147 26830 193
rect 26758 99 26830 147
rect 26758 53 26771 99
rect 26817 53 26830 99
rect 26758 5 26830 53
rect 26758 -41 26771 5
rect 26817 -41 26830 5
rect 26758 -89 26830 -41
rect 26758 -135 26771 -89
rect 26817 -135 26830 -89
rect 26758 -183 26830 -135
rect 26758 -229 26771 -183
rect 26817 -229 26830 -183
rect 26758 -277 26830 -229
rect 26758 -323 26771 -277
rect 26817 -323 26830 -277
rect 26758 -371 26830 -323
rect 26758 -417 26771 -371
rect 26817 -417 26830 -371
rect 26758 -465 26830 -417
rect 29766 3295 29838 3343
rect 29766 3249 29779 3295
rect 29825 3249 29838 3295
rect 26758 -511 26771 -465
rect 26817 -511 26830 -465
rect 26758 -559 26830 -511
rect 29766 3201 29838 3249
rect 29766 3155 29779 3201
rect 29825 3155 29838 3201
rect 29766 3107 29838 3155
rect 29766 3061 29779 3107
rect 29825 3061 29838 3107
rect 29766 3013 29838 3061
rect 29766 2967 29779 3013
rect 29825 2967 29838 3013
rect 29766 2919 29838 2967
rect 29766 2873 29779 2919
rect 29825 2873 29838 2919
rect 29766 2825 29838 2873
rect 29766 2779 29779 2825
rect 29825 2779 29838 2825
rect 29766 2731 29838 2779
rect 29766 2685 29779 2731
rect 29825 2685 29838 2731
rect 29766 2637 29838 2685
rect 29766 2591 29779 2637
rect 29825 2591 29838 2637
rect 29766 2543 29838 2591
rect 29766 2497 29779 2543
rect 29825 2497 29838 2543
rect 29766 2449 29838 2497
rect 29766 2403 29779 2449
rect 29825 2403 29838 2449
rect 29766 2355 29838 2403
rect 29766 2309 29779 2355
rect 29825 2309 29838 2355
rect 29766 2261 29838 2309
rect 29766 2215 29779 2261
rect 29825 2215 29838 2261
rect 29766 2167 29838 2215
rect 29766 2121 29779 2167
rect 29825 2121 29838 2167
rect 29766 2073 29838 2121
rect 29766 2027 29779 2073
rect 29825 2027 29838 2073
rect 29766 1979 29838 2027
rect 29766 1933 29779 1979
rect 29825 1933 29838 1979
rect 29766 1885 29838 1933
rect 29766 1839 29779 1885
rect 29825 1839 29838 1885
rect 29766 1791 29838 1839
rect 29766 1745 29779 1791
rect 29825 1745 29838 1791
rect 29766 1697 29838 1745
rect 29766 1651 29779 1697
rect 29825 1651 29838 1697
rect 29766 1603 29838 1651
rect 29766 1557 29779 1603
rect 29825 1557 29838 1603
rect 29766 1509 29838 1557
rect 29766 1463 29779 1509
rect 29825 1463 29838 1509
rect 29766 1415 29838 1463
rect 29766 1369 29779 1415
rect 29825 1369 29838 1415
rect 29766 1321 29838 1369
rect 29766 1275 29779 1321
rect 29825 1275 29838 1321
rect 29766 1227 29838 1275
rect 29766 1181 29779 1227
rect 29825 1181 29838 1227
rect 29766 1133 29838 1181
rect 29766 1087 29779 1133
rect 29825 1087 29838 1133
rect 29766 1039 29838 1087
rect 29766 993 29779 1039
rect 29825 993 29838 1039
rect 29766 945 29838 993
rect 29766 899 29779 945
rect 29825 899 29838 945
rect 29766 851 29838 899
rect 29766 805 29779 851
rect 29825 805 29838 851
rect 29766 757 29838 805
rect 29766 711 29779 757
rect 29825 711 29838 757
rect 29766 663 29838 711
rect 29766 617 29779 663
rect 29825 617 29838 663
rect 29766 569 29838 617
rect 29766 523 29779 569
rect 29825 523 29838 569
rect 29766 475 29838 523
rect 29766 429 29779 475
rect 29825 429 29838 475
rect 29766 381 29838 429
rect 29766 335 29779 381
rect 29825 335 29838 381
rect 29766 287 29838 335
rect 29766 241 29779 287
rect 29825 241 29838 287
rect 29766 193 29838 241
rect 29766 147 29779 193
rect 29825 147 29838 193
rect 29766 99 29838 147
rect 29766 53 29779 99
rect 29825 53 29838 99
rect 29766 5 29838 53
rect 29766 -41 29779 5
rect 29825 -41 29838 5
rect 29766 -89 29838 -41
rect 29766 -135 29779 -89
rect 29825 -135 29838 -89
rect 29766 -183 29838 -135
rect 29766 -229 29779 -183
rect 29825 -229 29838 -183
rect 29766 -277 29838 -229
rect 29766 -323 29779 -277
rect 29825 -323 29838 -277
rect 29766 -371 29838 -323
rect 29766 -417 29779 -371
rect 29825 -417 29838 -371
rect 26758 -605 26771 -559
rect 26817 -605 26830 -559
rect 26758 -653 26830 -605
rect 29766 -465 29838 -417
rect 29766 -511 29779 -465
rect 29825 -511 29838 -465
rect 29766 -559 29838 -511
rect 29766 -605 29779 -559
rect 29825 -605 29838 -559
rect 26758 -699 26771 -653
rect 26817 -699 26830 -653
rect 26758 -747 26830 -699
rect 26758 -793 26771 -747
rect 26817 -793 26830 -747
rect 26758 -841 26830 -793
rect 26758 -887 26771 -841
rect 26817 -887 26830 -841
rect 26758 -935 26830 -887
rect 26758 -981 26771 -935
rect 26817 -981 26830 -935
rect 26758 -1029 26830 -981
rect 26758 -1075 26771 -1029
rect 26817 -1075 26830 -1029
rect 26758 -1123 26830 -1075
rect 26758 -1169 26771 -1123
rect 26817 -1169 26830 -1123
rect 26758 -1217 26830 -1169
rect 26758 -1263 26771 -1217
rect 26817 -1263 26830 -1217
rect 29766 -653 29838 -605
rect 29766 -699 29779 -653
rect 29825 -699 29838 -653
rect 29766 -747 29838 -699
rect 29766 -793 29779 -747
rect 29825 -793 29838 -747
rect 29766 -841 29838 -793
rect 29766 -887 29779 -841
rect 29825 -887 29838 -841
rect 29766 -935 29838 -887
rect 29766 -981 29779 -935
rect 29825 -981 29838 -935
rect 29766 -1029 29838 -981
rect 29766 -1075 29779 -1029
rect 29825 -1075 29838 -1029
rect 29766 -1123 29838 -1075
rect 29766 -1169 29779 -1123
rect 29825 -1169 29838 -1123
rect 29766 -1217 29838 -1169
rect 26758 -1311 26830 -1263
rect 26758 -1357 26771 -1311
rect 26817 -1357 26830 -1311
rect 26758 -1405 26830 -1357
rect 29766 -1263 29779 -1217
rect 29825 -1263 29838 -1217
rect 29766 -1311 29838 -1263
rect 29766 -1357 29779 -1311
rect 29825 -1357 29838 -1311
rect 26758 -1451 26771 -1405
rect 26817 -1451 26830 -1405
rect 26758 -1499 26830 -1451
rect 29766 -1405 29838 -1357
rect 29766 -1451 29779 -1405
rect 29825 -1451 29838 -1405
rect 26758 -1545 26771 -1499
rect 26817 -1545 26830 -1499
rect 26758 -1593 26830 -1545
rect 26758 -1639 26771 -1593
rect 26817 -1639 26830 -1593
rect 26758 -1687 26830 -1639
rect 26758 -1733 26771 -1687
rect 26817 -1733 26830 -1687
rect 26758 -1768 26830 -1733
rect 29766 -1499 29838 -1451
rect 29766 -1545 29779 -1499
rect 29825 -1545 29838 -1499
rect 29766 -1593 29838 -1545
rect 29766 -1639 29779 -1593
rect 29825 -1639 29838 -1593
rect 29766 -1687 29838 -1639
rect 29766 -1733 29779 -1687
rect 29825 -1733 29838 -1687
rect 29766 -1768 29838 -1733
rect 26758 -1781 29838 -1768
rect 26758 -1827 26771 -1781
rect 26817 -1827 26865 -1781
rect 26911 -1827 26959 -1781
rect 27005 -1827 27053 -1781
rect 27099 -1827 27147 -1781
rect 27193 -1827 27241 -1781
rect 27287 -1827 27335 -1781
rect 27381 -1827 27429 -1781
rect 27475 -1827 27523 -1781
rect 27569 -1827 27617 -1781
rect 27663 -1827 27711 -1781
rect 27757 -1827 27805 -1781
rect 27851 -1827 27899 -1781
rect 27945 -1827 27993 -1781
rect 28039 -1827 28087 -1781
rect 28133 -1827 28181 -1781
rect 28227 -1827 28275 -1781
rect 28321 -1827 28369 -1781
rect 28415 -1827 28463 -1781
rect 28509 -1827 28557 -1781
rect 28603 -1827 28651 -1781
rect 28697 -1827 28745 -1781
rect 28791 -1827 28839 -1781
rect 28885 -1827 28933 -1781
rect 28979 -1827 29027 -1781
rect 29073 -1827 29121 -1781
rect 29167 -1827 29215 -1781
rect 29261 -1827 29309 -1781
rect 29355 -1827 29403 -1781
rect 29449 -1827 29497 -1781
rect 29543 -1827 29591 -1781
rect 29637 -1827 29685 -1781
rect 29731 -1827 29779 -1781
rect 29825 -1827 29838 -1781
rect 26758 -1840 29838 -1827
rect 6435 -3039 9609 -3026
rect 6435 -3085 6448 -3039
rect 6494 -3085 6542 -3039
rect 6588 -3085 6636 -3039
rect 6682 -3085 6730 -3039
rect 6776 -3085 6824 -3039
rect 6870 -3085 6918 -3039
rect 6964 -3085 7012 -3039
rect 7058 -3085 7106 -3039
rect 7152 -3085 7200 -3039
rect 7246 -3085 7294 -3039
rect 7340 -3085 7388 -3039
rect 7434 -3085 7482 -3039
rect 7528 -3085 7576 -3039
rect 7622 -3085 7670 -3039
rect 7716 -3085 7764 -3039
rect 7810 -3085 7858 -3039
rect 7904 -3085 7952 -3039
rect 7998 -3085 8046 -3039
rect 8092 -3085 8140 -3039
rect 8186 -3085 8234 -3039
rect 8280 -3085 8328 -3039
rect 8374 -3085 8422 -3039
rect 8468 -3085 8516 -3039
rect 8562 -3085 8610 -3039
rect 8656 -3085 8704 -3039
rect 8750 -3085 8798 -3039
rect 8844 -3085 8892 -3039
rect 8938 -3085 8986 -3039
rect 9032 -3085 9080 -3039
rect 9126 -3085 9174 -3039
rect 9220 -3085 9268 -3039
rect 9314 -3085 9362 -3039
rect 9408 -3085 9456 -3039
rect 9502 -3085 9550 -3039
rect 9596 -3085 9609 -3039
rect 6435 -3098 9609 -3085
rect 6435 -3133 6507 -3098
rect 6435 -3179 6448 -3133
rect 6494 -3179 6507 -3133
rect 6435 -3227 6507 -3179
rect 9537 -3133 9609 -3098
rect 9537 -3179 9550 -3133
rect 9596 -3179 9609 -3133
rect 6435 -3273 6448 -3227
rect 6494 -3273 6507 -3227
rect 6435 -3321 6507 -3273
rect 6435 -3367 6448 -3321
rect 6494 -3367 6507 -3321
rect 6435 -3415 6507 -3367
rect 6435 -3461 6448 -3415
rect 6494 -3461 6507 -3415
rect 9537 -3227 9609 -3179
rect 9537 -3273 9550 -3227
rect 9596 -3273 9609 -3227
rect 9537 -3321 9609 -3273
rect 9537 -3367 9550 -3321
rect 9596 -3367 9609 -3321
rect 9537 -3415 9609 -3367
rect 6435 -3509 6507 -3461
rect 6435 -3555 6448 -3509
rect 6494 -3555 6507 -3509
rect 6435 -3603 6507 -3555
rect 6435 -3649 6448 -3603
rect 6494 -3649 6507 -3603
rect 9537 -3461 9550 -3415
rect 9596 -3461 9609 -3415
rect 9537 -3509 9609 -3461
rect 9537 -3555 9550 -3509
rect 9596 -3555 9609 -3509
rect 9537 -3603 9609 -3555
rect 6435 -3697 6507 -3649
rect 6435 -3743 6448 -3697
rect 6494 -3743 6507 -3697
rect 6435 -3791 6507 -3743
rect 6435 -3837 6448 -3791
rect 6494 -3837 6507 -3791
rect 6435 -3885 6507 -3837
rect 6435 -3931 6448 -3885
rect 6494 -3931 6507 -3885
rect 6435 -3979 6507 -3931
rect 6435 -4025 6448 -3979
rect 6494 -4025 6507 -3979
rect 6435 -4073 6507 -4025
rect 6435 -4119 6448 -4073
rect 6494 -4119 6507 -4073
rect 6435 -4167 6507 -4119
rect 6435 -4213 6448 -4167
rect 6494 -4213 6507 -4167
rect 6435 -4261 6507 -4213
rect 6435 -4307 6448 -4261
rect 6494 -4307 6507 -4261
rect 6435 -4355 6507 -4307
rect 6435 -4401 6448 -4355
rect 6494 -4401 6507 -4355
rect 6435 -4449 6507 -4401
rect 6435 -4495 6448 -4449
rect 6494 -4495 6507 -4449
rect 6435 -4543 6507 -4495
rect 6435 -4589 6448 -4543
rect 6494 -4589 6507 -4543
rect 6435 -4637 6507 -4589
rect 6435 -4683 6448 -4637
rect 6494 -4683 6507 -4637
rect 6435 -4731 6507 -4683
rect 6435 -4777 6448 -4731
rect 6494 -4777 6507 -4731
rect 6435 -4825 6507 -4777
rect 6435 -4871 6448 -4825
rect 6494 -4871 6507 -4825
rect 6435 -4919 6507 -4871
rect 6435 -4965 6448 -4919
rect 6494 -4965 6507 -4919
rect 6435 -5013 6507 -4965
rect 6435 -5059 6448 -5013
rect 6494 -5059 6507 -5013
rect 6435 -5107 6507 -5059
rect 6435 -5153 6448 -5107
rect 6494 -5153 6507 -5107
rect 6435 -5201 6507 -5153
rect 6435 -5247 6448 -5201
rect 6494 -5247 6507 -5201
rect 6435 -5295 6507 -5247
rect 6435 -5341 6448 -5295
rect 6494 -5341 6507 -5295
rect 6435 -5389 6507 -5341
rect 6435 -5435 6448 -5389
rect 6494 -5435 6507 -5389
rect 6435 -5483 6507 -5435
rect 6435 -5529 6448 -5483
rect 6494 -5529 6507 -5483
rect 6435 -5577 6507 -5529
rect 6435 -5623 6448 -5577
rect 6494 -5623 6507 -5577
rect 6435 -5671 6507 -5623
rect 6435 -5717 6448 -5671
rect 6494 -5717 6507 -5671
rect 6435 -5765 6507 -5717
rect 6435 -5811 6448 -5765
rect 6494 -5811 6507 -5765
rect 6435 -5859 6507 -5811
rect 6435 -5905 6448 -5859
rect 6494 -5905 6507 -5859
rect 6435 -5953 6507 -5905
rect 6435 -5999 6448 -5953
rect 6494 -5999 6507 -5953
rect 6435 -6047 6507 -5999
rect 6435 -6093 6448 -6047
rect 6494 -6093 6507 -6047
rect 6435 -6141 6507 -6093
rect 9537 -3649 9550 -3603
rect 9596 -3649 9609 -3603
rect 9537 -3697 9609 -3649
rect 9537 -3743 9550 -3697
rect 9596 -3743 9609 -3697
rect 9537 -3791 9609 -3743
rect 9537 -3837 9550 -3791
rect 9596 -3837 9609 -3791
rect 9537 -3885 9609 -3837
rect 9537 -3931 9550 -3885
rect 9596 -3931 9609 -3885
rect 9537 -3979 9609 -3931
rect 9537 -4025 9550 -3979
rect 9596 -4025 9609 -3979
rect 9537 -4073 9609 -4025
rect 9537 -4119 9550 -4073
rect 9596 -4119 9609 -4073
rect 9537 -4167 9609 -4119
rect 9537 -4213 9550 -4167
rect 9596 -4213 9609 -4167
rect 9537 -4261 9609 -4213
rect 9537 -4307 9550 -4261
rect 9596 -4307 9609 -4261
rect 9537 -4355 9609 -4307
rect 9537 -4401 9550 -4355
rect 9596 -4401 9609 -4355
rect 9537 -4449 9609 -4401
rect 9537 -4495 9550 -4449
rect 9596 -4495 9609 -4449
rect 9537 -4543 9609 -4495
rect 9537 -4589 9550 -4543
rect 9596 -4589 9609 -4543
rect 9537 -4637 9609 -4589
rect 9537 -4683 9550 -4637
rect 9596 -4683 9609 -4637
rect 9537 -4731 9609 -4683
rect 9537 -4777 9550 -4731
rect 9596 -4777 9609 -4731
rect 9537 -4825 9609 -4777
rect 9537 -4871 9550 -4825
rect 9596 -4871 9609 -4825
rect 9537 -4919 9609 -4871
rect 9537 -4965 9550 -4919
rect 9596 -4965 9609 -4919
rect 9537 -5013 9609 -4965
rect 9537 -5059 9550 -5013
rect 9596 -5059 9609 -5013
rect 9537 -5107 9609 -5059
rect 9537 -5153 9550 -5107
rect 9596 -5153 9609 -5107
rect 9537 -5201 9609 -5153
rect 9537 -5247 9550 -5201
rect 9596 -5247 9609 -5201
rect 9537 -5295 9609 -5247
rect 9537 -5341 9550 -5295
rect 9596 -5341 9609 -5295
rect 9537 -5389 9609 -5341
rect 9537 -5435 9550 -5389
rect 9596 -5435 9609 -5389
rect 9537 -5483 9609 -5435
rect 9537 -5529 9550 -5483
rect 9596 -5529 9609 -5483
rect 9537 -5577 9609 -5529
rect 9537 -5623 9550 -5577
rect 9596 -5623 9609 -5577
rect 9537 -5671 9609 -5623
rect 9537 -5717 9550 -5671
rect 9596 -5717 9609 -5671
rect 9537 -5765 9609 -5717
rect 9537 -5811 9550 -5765
rect 9596 -5811 9609 -5765
rect 9537 -5859 9609 -5811
rect 9537 -5905 9550 -5859
rect 9596 -5905 9609 -5859
rect 9537 -5953 9609 -5905
rect 9537 -5999 9550 -5953
rect 9596 -5999 9609 -5953
rect 9537 -6047 9609 -5999
rect 9537 -6093 9550 -6047
rect 9596 -6093 9609 -6047
rect 6435 -6187 6448 -6141
rect 6494 -6187 6507 -6141
rect 6435 -6235 6507 -6187
rect 6435 -6281 6448 -6235
rect 6494 -6281 6507 -6235
rect 6435 -6316 6507 -6281
rect 9537 -6141 9609 -6093
rect 9537 -6187 9550 -6141
rect 9596 -6187 9609 -6141
rect 9537 -6235 9609 -6187
rect 9537 -6281 9550 -6235
rect 9596 -6281 9609 -6235
rect 5401 -6329 6507 -6316
rect 5401 -6375 5414 -6329
rect 5460 -6375 5508 -6329
rect 5554 -6375 5602 -6329
rect 5648 -6375 5696 -6329
rect 5742 -6375 5790 -6329
rect 5836 -6375 5884 -6329
rect 5930 -6375 5978 -6329
rect 6024 -6375 6072 -6329
rect 6118 -6375 6166 -6329
rect 6212 -6375 6260 -6329
rect 6306 -6375 6354 -6329
rect 6400 -6375 6448 -6329
rect 6494 -6375 6507 -6329
rect 5401 -6388 6507 -6375
rect 9537 -6316 9609 -6281
rect 11515 -4688 17133 -4675
rect 11515 -4734 11528 -4688
rect 11574 -4734 11622 -4688
rect 11668 -4734 11716 -4688
rect 11762 -4734 11810 -4688
rect 11856 -4734 11904 -4688
rect 11950 -4734 11998 -4688
rect 12044 -4734 12092 -4688
rect 12138 -4734 12186 -4688
rect 12232 -4734 12280 -4688
rect 12326 -4734 12374 -4688
rect 12420 -4734 12468 -4688
rect 12514 -4734 12562 -4688
rect 12608 -4734 12656 -4688
rect 12702 -4734 12750 -4688
rect 12796 -4734 12844 -4688
rect 12890 -4734 12938 -4688
rect 12984 -4734 13032 -4688
rect 13078 -4734 13126 -4688
rect 13172 -4734 13220 -4688
rect 13266 -4734 13314 -4688
rect 13360 -4734 13408 -4688
rect 13454 -4734 13502 -4688
rect 13548 -4734 13596 -4688
rect 13642 -4734 13690 -4688
rect 13736 -4734 13784 -4688
rect 13830 -4734 13878 -4688
rect 13924 -4734 13972 -4688
rect 14018 -4734 14066 -4688
rect 14112 -4734 14160 -4688
rect 14206 -4734 14254 -4688
rect 14300 -4734 14348 -4688
rect 14394 -4734 14442 -4688
rect 14488 -4734 14536 -4688
rect 14582 -4734 14630 -4688
rect 14676 -4734 14724 -4688
rect 14770 -4734 14818 -4688
rect 14864 -4734 14912 -4688
rect 14958 -4734 15006 -4688
rect 15052 -4734 15100 -4688
rect 15146 -4734 15194 -4688
rect 15240 -4734 15288 -4688
rect 15334 -4734 15382 -4688
rect 15428 -4734 15476 -4688
rect 15522 -4734 15570 -4688
rect 15616 -4734 15664 -4688
rect 15710 -4734 15758 -4688
rect 15804 -4734 15852 -4688
rect 15898 -4734 15946 -4688
rect 15992 -4734 16040 -4688
rect 16086 -4734 16134 -4688
rect 16180 -4734 16228 -4688
rect 16274 -4734 16322 -4688
rect 16368 -4734 16416 -4688
rect 16462 -4734 16510 -4688
rect 16556 -4734 16604 -4688
rect 16650 -4734 16698 -4688
rect 16744 -4734 16792 -4688
rect 16838 -4734 16886 -4688
rect 16932 -4734 16980 -4688
rect 17026 -4734 17074 -4688
rect 17120 -4734 17133 -4688
rect 11515 -4747 17133 -4734
rect 11515 -4782 11587 -4747
rect 11515 -4828 11528 -4782
rect 11574 -4828 11587 -4782
rect 11515 -4876 11587 -4828
rect 11515 -4922 11528 -4876
rect 11574 -4922 11587 -4876
rect 11515 -4970 11587 -4922
rect 11515 -5016 11528 -4970
rect 11574 -5016 11587 -4970
rect 11515 -5064 11587 -5016
rect 11515 -5110 11528 -5064
rect 11574 -5110 11587 -5064
rect 17061 -4782 17133 -4747
rect 17061 -4828 17074 -4782
rect 17120 -4828 17133 -4782
rect 17061 -4876 17133 -4828
rect 17061 -4922 17074 -4876
rect 17120 -4922 17133 -4876
rect 17061 -4970 17133 -4922
rect 17061 -5016 17074 -4970
rect 17120 -5016 17133 -4970
rect 17061 -5064 17133 -5016
rect 11515 -5158 11587 -5110
rect 11515 -5204 11528 -5158
rect 11574 -5204 11587 -5158
rect 11515 -5252 11587 -5204
rect 11515 -5298 11528 -5252
rect 11574 -5298 11587 -5252
rect 11515 -5346 11587 -5298
rect 11515 -5392 11528 -5346
rect 11574 -5392 11587 -5346
rect 17061 -5110 17074 -5064
rect 17120 -5110 17133 -5064
rect 17061 -5158 17133 -5110
rect 17061 -5204 17074 -5158
rect 17120 -5204 17133 -5158
rect 17061 -5252 17133 -5204
rect 17061 -5298 17074 -5252
rect 17120 -5298 17133 -5252
rect 17061 -5346 17133 -5298
rect 11515 -5440 11587 -5392
rect 11515 -5486 11528 -5440
rect 11574 -5486 11587 -5440
rect 11515 -5534 11587 -5486
rect 11515 -5580 11528 -5534
rect 11574 -5580 11587 -5534
rect 11515 -5628 11587 -5580
rect 11515 -5674 11528 -5628
rect 11574 -5674 11587 -5628
rect 11515 -5722 11587 -5674
rect 11515 -5768 11528 -5722
rect 11574 -5768 11587 -5722
rect 11515 -5816 11587 -5768
rect 17061 -5392 17074 -5346
rect 17120 -5392 17133 -5346
rect 17061 -5440 17133 -5392
rect 17061 -5486 17074 -5440
rect 17120 -5486 17133 -5440
rect 17061 -5534 17133 -5486
rect 17061 -5580 17074 -5534
rect 17120 -5580 17133 -5534
rect 17061 -5628 17133 -5580
rect 17061 -5674 17074 -5628
rect 17120 -5674 17133 -5628
rect 17061 -5722 17133 -5674
rect 17061 -5768 17074 -5722
rect 17120 -5768 17133 -5722
rect 11515 -5862 11528 -5816
rect 11574 -5862 11587 -5816
rect 11515 -5910 11587 -5862
rect 11515 -5956 11528 -5910
rect 11574 -5956 11587 -5910
rect 11515 -6004 11587 -5956
rect 11515 -6050 11528 -6004
rect 11574 -6050 11587 -6004
rect 11515 -6098 11587 -6050
rect 11515 -6144 11528 -6098
rect 11574 -6144 11587 -6098
rect 11515 -6192 11587 -6144
rect 11515 -6238 11528 -6192
rect 11574 -6238 11587 -6192
rect 11515 -6286 11587 -6238
rect 9537 -6329 10643 -6316
rect 9537 -6375 9550 -6329
rect 9596 -6375 9644 -6329
rect 9690 -6375 9738 -6329
rect 9784 -6375 9832 -6329
rect 9878 -6375 9926 -6329
rect 9972 -6375 10020 -6329
rect 10066 -6375 10114 -6329
rect 10160 -6375 10208 -6329
rect 10254 -6375 10302 -6329
rect 10348 -6375 10396 -6329
rect 10442 -6375 10490 -6329
rect 10536 -6375 10584 -6329
rect 10630 -6375 10643 -6329
rect 5401 -6423 5473 -6388
rect 9537 -6388 10643 -6375
rect 10571 -6423 10643 -6388
rect 5401 -6469 5414 -6423
rect 5460 -6469 5473 -6423
rect 5401 -6517 5473 -6469
rect 10571 -6469 10584 -6423
rect 10630 -6469 10643 -6423
rect 5401 -6563 5414 -6517
rect 5460 -6563 5473 -6517
rect 5401 -6611 5473 -6563
rect 5401 -6657 5414 -6611
rect 5460 -6657 5473 -6611
rect 5401 -6705 5473 -6657
rect 5401 -6751 5414 -6705
rect 5460 -6751 5473 -6705
rect 10571 -6517 10643 -6469
rect 10571 -6563 10584 -6517
rect 10630 -6563 10643 -6517
rect 10571 -6611 10643 -6563
rect 10571 -6657 10584 -6611
rect 10630 -6657 10643 -6611
rect 10571 -6705 10643 -6657
rect 5401 -6799 5473 -6751
rect 5401 -6845 5414 -6799
rect 5460 -6845 5473 -6799
rect 5401 -6893 5473 -6845
rect 5401 -6939 5414 -6893
rect 5460 -6939 5473 -6893
rect 10571 -6751 10584 -6705
rect 10630 -6751 10643 -6705
rect 10571 -6799 10643 -6751
rect 10571 -6845 10584 -6799
rect 10630 -6845 10643 -6799
rect 10571 -6893 10643 -6845
rect 5401 -6987 5473 -6939
rect 5401 -7033 5414 -6987
rect 5460 -7033 5473 -6987
rect 5401 -7081 5473 -7033
rect 5401 -7127 5414 -7081
rect 5460 -7127 5473 -7081
rect 10571 -6939 10584 -6893
rect 10630 -6939 10643 -6893
rect 10571 -6987 10643 -6939
rect 10571 -7033 10584 -6987
rect 10630 -7033 10643 -6987
rect 10571 -7081 10643 -7033
rect 5401 -7175 5473 -7127
rect 5401 -7221 5414 -7175
rect 5460 -7221 5473 -7175
rect 10571 -7127 10584 -7081
rect 10630 -7127 10643 -7081
rect 10571 -7175 10643 -7127
rect 5401 -7269 5473 -7221
rect 5401 -7315 5414 -7269
rect 5460 -7315 5473 -7269
rect 5401 -7363 5473 -7315
rect 5401 -7409 5414 -7363
rect 5460 -7409 5473 -7363
rect 10571 -7221 10584 -7175
rect 10630 -7221 10643 -7175
rect 10571 -7269 10643 -7221
rect 10571 -7315 10584 -7269
rect 10630 -7315 10643 -7269
rect 10571 -7363 10643 -7315
rect 5401 -7457 5473 -7409
rect 5401 -7503 5414 -7457
rect 5460 -7503 5473 -7457
rect 5401 -7551 5473 -7503
rect 5401 -7597 5414 -7551
rect 5460 -7597 5473 -7551
rect 5401 -7645 5473 -7597
rect 5401 -7691 5414 -7645
rect 5460 -7691 5473 -7645
rect 5401 -7739 5473 -7691
rect 5401 -7785 5414 -7739
rect 5460 -7785 5473 -7739
rect 5401 -7820 5473 -7785
rect 10571 -7409 10584 -7363
rect 10630 -7409 10643 -7363
rect 10571 -7457 10643 -7409
rect 10571 -7503 10584 -7457
rect 10630 -7503 10643 -7457
rect 10571 -7551 10643 -7503
rect 10571 -7597 10584 -7551
rect 10630 -7597 10643 -7551
rect 10571 -7645 10643 -7597
rect 10571 -7691 10584 -7645
rect 10630 -7691 10643 -7645
rect 10571 -7739 10643 -7691
rect 10571 -7785 10584 -7739
rect 10630 -7785 10643 -7739
rect 10571 -7820 10643 -7785
rect 5401 -7833 10643 -7820
rect 5401 -7879 5414 -7833
rect 5460 -7879 5508 -7833
rect 5554 -7879 5602 -7833
rect 5648 -7879 5696 -7833
rect 5742 -7879 5790 -7833
rect 5836 -7879 5884 -7833
rect 5930 -7879 5978 -7833
rect 6024 -7879 6072 -7833
rect 6118 -7879 6166 -7833
rect 6212 -7879 6260 -7833
rect 6306 -7879 6354 -7833
rect 6400 -7879 6448 -7833
rect 6494 -7879 6542 -7833
rect 6588 -7879 6636 -7833
rect 6682 -7879 6730 -7833
rect 6776 -7879 6824 -7833
rect 6870 -7879 6918 -7833
rect 6964 -7879 7012 -7833
rect 7058 -7879 7106 -7833
rect 7152 -7879 7200 -7833
rect 7246 -7879 7294 -7833
rect 7340 -7879 7388 -7833
rect 7434 -7879 7482 -7833
rect 7528 -7879 7576 -7833
rect 7622 -7879 7670 -7833
rect 7716 -7879 7764 -7833
rect 7810 -7879 7858 -7833
rect 7904 -7879 7952 -7833
rect 7998 -7879 8046 -7833
rect 8092 -7879 8140 -7833
rect 8186 -7879 8234 -7833
rect 8280 -7879 8328 -7833
rect 8374 -7879 8422 -7833
rect 8468 -7879 8516 -7833
rect 8562 -7879 8610 -7833
rect 8656 -7879 8704 -7833
rect 8750 -7879 8798 -7833
rect 8844 -7879 8892 -7833
rect 8938 -7879 8986 -7833
rect 9032 -7879 9080 -7833
rect 9126 -7879 9174 -7833
rect 9220 -7879 9268 -7833
rect 9314 -7879 9362 -7833
rect 9408 -7879 9456 -7833
rect 9502 -7879 9550 -7833
rect 9596 -7879 9644 -7833
rect 9690 -7879 9738 -7833
rect 9784 -7879 9832 -7833
rect 9878 -7879 9926 -7833
rect 9972 -7879 10020 -7833
rect 10066 -7879 10114 -7833
rect 10160 -7879 10208 -7833
rect 10254 -7879 10302 -7833
rect 10348 -7879 10396 -7833
rect 10442 -7879 10490 -7833
rect 10536 -7879 10584 -7833
rect 10630 -7879 10643 -7833
rect 11515 -6332 11528 -6286
rect 11574 -6332 11587 -6286
rect 11515 -6380 11587 -6332
rect 11515 -6426 11528 -6380
rect 11574 -6426 11587 -6380
rect 11515 -6474 11587 -6426
rect 11515 -6520 11528 -6474
rect 11574 -6520 11587 -6474
rect 11515 -6568 11587 -6520
rect 11515 -6614 11528 -6568
rect 11574 -6614 11587 -6568
rect 11515 -6662 11587 -6614
rect 11515 -6708 11528 -6662
rect 11574 -6708 11587 -6662
rect 11515 -6756 11587 -6708
rect 17061 -5816 17133 -5768
rect 17061 -5862 17074 -5816
rect 17120 -5862 17133 -5816
rect 17061 -5910 17133 -5862
rect 17061 -5956 17074 -5910
rect 17120 -5956 17133 -5910
rect 17061 -6004 17133 -5956
rect 17061 -6050 17074 -6004
rect 17120 -6050 17133 -6004
rect 17061 -6098 17133 -6050
rect 17061 -6144 17074 -6098
rect 17120 -6144 17133 -6098
rect 17061 -6192 17133 -6144
rect 17061 -6238 17074 -6192
rect 17120 -6238 17133 -6192
rect 17061 -6286 17133 -6238
rect 17061 -6332 17074 -6286
rect 17120 -6332 17133 -6286
rect 17061 -6380 17133 -6332
rect 17061 -6426 17074 -6380
rect 17120 -6426 17133 -6380
rect 17061 -6474 17133 -6426
rect 17061 -6520 17074 -6474
rect 17120 -6520 17133 -6474
rect 17061 -6568 17133 -6520
rect 17061 -6614 17074 -6568
rect 17120 -6614 17133 -6568
rect 17061 -6662 17133 -6614
rect 17061 -6708 17074 -6662
rect 17120 -6708 17133 -6662
rect 11515 -6802 11528 -6756
rect 11574 -6802 11587 -6756
rect 11515 -6850 11587 -6802
rect 11515 -6896 11528 -6850
rect 11574 -6896 11587 -6850
rect 11515 -6944 11587 -6896
rect 11515 -6990 11528 -6944
rect 11574 -6990 11587 -6944
rect 11515 -7038 11587 -6990
rect 11515 -7084 11528 -7038
rect 11574 -7084 11587 -7038
rect 11515 -7132 11587 -7084
rect 11515 -7178 11528 -7132
rect 11574 -7178 11587 -7132
rect 17061 -6756 17133 -6708
rect 17061 -6802 17074 -6756
rect 17120 -6802 17133 -6756
rect 17061 -6850 17133 -6802
rect 17061 -6896 17074 -6850
rect 17120 -6896 17133 -6850
rect 17061 -6944 17133 -6896
rect 17061 -6990 17074 -6944
rect 17120 -6990 17133 -6944
rect 17061 -7038 17133 -6990
rect 17061 -7084 17074 -7038
rect 17120 -7084 17133 -7038
rect 17061 -7132 17133 -7084
rect 11515 -7226 11587 -7178
rect 11515 -7272 11528 -7226
rect 11574 -7272 11587 -7226
rect 11515 -7320 11587 -7272
rect 11515 -7366 11528 -7320
rect 11574 -7366 11587 -7320
rect 11515 -7414 11587 -7366
rect 11515 -7460 11528 -7414
rect 11574 -7460 11587 -7414
rect 11515 -7508 11587 -7460
rect 11515 -7554 11528 -7508
rect 11574 -7554 11587 -7508
rect 17061 -7178 17074 -7132
rect 17120 -7178 17133 -7132
rect 17061 -7226 17133 -7178
rect 17061 -7272 17074 -7226
rect 17120 -7272 17133 -7226
rect 17061 -7320 17133 -7272
rect 17061 -7366 17074 -7320
rect 17120 -7366 17133 -7320
rect 17061 -7414 17133 -7366
rect 17061 -7460 17074 -7414
rect 17120 -7460 17133 -7414
rect 17061 -7508 17133 -7460
rect 11515 -7602 11587 -7554
rect 11515 -7648 11528 -7602
rect 11574 -7648 11587 -7602
rect 11515 -7696 11587 -7648
rect 11515 -7742 11528 -7696
rect 11574 -7742 11587 -7696
rect 11515 -7777 11587 -7742
rect 17061 -7554 17074 -7508
rect 17120 -7554 17133 -7508
rect 17061 -7602 17133 -7554
rect 17061 -7648 17074 -7602
rect 17120 -7648 17133 -7602
rect 17061 -7696 17133 -7648
rect 17061 -7742 17074 -7696
rect 17120 -7742 17133 -7696
rect 17061 -7777 17133 -7742
rect 11515 -7790 17133 -7777
rect 11515 -7836 11528 -7790
rect 11574 -7836 11622 -7790
rect 11668 -7836 11716 -7790
rect 11762 -7836 11810 -7790
rect 11856 -7836 11904 -7790
rect 11950 -7836 11998 -7790
rect 12044 -7836 12092 -7790
rect 12138 -7836 12186 -7790
rect 12232 -7836 12280 -7790
rect 12326 -7836 12374 -7790
rect 12420 -7836 12468 -7790
rect 12514 -7836 12562 -7790
rect 12608 -7836 12656 -7790
rect 12702 -7836 12750 -7790
rect 12796 -7836 12844 -7790
rect 12890 -7836 12938 -7790
rect 12984 -7836 13032 -7790
rect 13078 -7836 13126 -7790
rect 13172 -7836 13220 -7790
rect 13266 -7836 13314 -7790
rect 13360 -7836 13408 -7790
rect 13454 -7836 13502 -7790
rect 13548 -7836 13596 -7790
rect 13642 -7836 13690 -7790
rect 13736 -7836 13784 -7790
rect 13830 -7836 13878 -7790
rect 13924 -7836 13972 -7790
rect 14018 -7836 14066 -7790
rect 14112 -7836 14160 -7790
rect 14206 -7836 14254 -7790
rect 14300 -7836 14348 -7790
rect 14394 -7836 14442 -7790
rect 14488 -7836 14536 -7790
rect 14582 -7836 14630 -7790
rect 14676 -7836 14724 -7790
rect 14770 -7836 14818 -7790
rect 14864 -7836 14912 -7790
rect 14958 -7836 15006 -7790
rect 15052 -7836 15100 -7790
rect 15146 -7836 15194 -7790
rect 15240 -7836 15288 -7790
rect 15334 -7836 15382 -7790
rect 15428 -7836 15476 -7790
rect 15522 -7836 15570 -7790
rect 15616 -7836 15664 -7790
rect 15710 -7836 15758 -7790
rect 15804 -7836 15852 -7790
rect 15898 -7836 15946 -7790
rect 15992 -7836 16040 -7790
rect 16086 -7836 16134 -7790
rect 16180 -7836 16228 -7790
rect 16274 -7836 16322 -7790
rect 16368 -7836 16416 -7790
rect 16462 -7836 16510 -7790
rect 16556 -7836 16604 -7790
rect 16650 -7836 16698 -7790
rect 16744 -7836 16792 -7790
rect 16838 -7836 16886 -7790
rect 16932 -7836 16980 -7790
rect 17026 -7836 17074 -7790
rect 17120 -7836 17133 -7790
rect 11515 -7849 17133 -7836
rect 5401 -7892 10643 -7879
<< nsubdiff >>
rect 2945 5217 5179 5230
rect 2945 5171 2958 5217
rect 3004 5171 3052 5217
rect 3098 5171 3146 5217
rect 3192 5171 3240 5217
rect 3286 5171 3334 5217
rect 3380 5171 3428 5217
rect 3474 5171 3522 5217
rect 3568 5171 3616 5217
rect 3662 5171 3710 5217
rect 3756 5171 3804 5217
rect 3850 5171 3898 5217
rect 3944 5171 3992 5217
rect 4038 5171 4086 5217
rect 4132 5171 4180 5217
rect 4226 5171 4274 5217
rect 4320 5171 4368 5217
rect 4414 5171 4462 5217
rect 4508 5171 4556 5217
rect 4602 5171 4650 5217
rect 4696 5171 4744 5217
rect 4790 5171 4838 5217
rect 4884 5171 4932 5217
rect 4978 5171 5026 5217
rect 5072 5171 5120 5217
rect 5166 5171 5179 5217
rect 2945 5158 5179 5171
rect 2945 5123 3017 5158
rect 2945 5077 2958 5123
rect 3004 5077 3017 5123
rect 2945 5029 3017 5077
rect 5107 5123 5179 5158
rect 5107 5077 5120 5123
rect 5166 5077 5179 5123
rect 2945 4983 2958 5029
rect 3004 4983 3017 5029
rect 5107 5029 5179 5077
rect 2945 4935 3017 4983
rect 2945 4889 2958 4935
rect 3004 4889 3017 4935
rect 2945 4841 3017 4889
rect 5107 4983 5120 5029
rect 5166 4983 5179 5029
rect 5107 4935 5179 4983
rect 5107 4889 5120 4935
rect 5166 4889 5179 4935
rect 2945 4795 2958 4841
rect 3004 4795 3017 4841
rect 2945 4747 3017 4795
rect 2945 4701 2958 4747
rect 3004 4701 3017 4747
rect 2945 4653 3017 4701
rect 2945 4607 2958 4653
rect 3004 4607 3017 4653
rect 2945 4559 3017 4607
rect 2945 4513 2958 4559
rect 3004 4513 3017 4559
rect 2945 4465 3017 4513
rect 2945 4419 2958 4465
rect 3004 4419 3017 4465
rect 2945 4371 3017 4419
rect 2945 4325 2958 4371
rect 3004 4325 3017 4371
rect 2945 4277 3017 4325
rect 2945 4231 2958 4277
rect 3004 4231 3017 4277
rect 2945 4183 3017 4231
rect 2945 4137 2958 4183
rect 3004 4137 3017 4183
rect 2945 4089 3017 4137
rect 5107 4841 5179 4889
rect 5107 4795 5120 4841
rect 5166 4795 5179 4841
rect 5107 4747 5179 4795
rect 5107 4701 5120 4747
rect 5166 4701 5179 4747
rect 5107 4653 5179 4701
rect 5107 4607 5120 4653
rect 5166 4607 5179 4653
rect 5107 4559 5179 4607
rect 5107 4513 5120 4559
rect 5166 4513 5179 4559
rect 5107 4465 5179 4513
rect 5107 4419 5120 4465
rect 5166 4419 5179 4465
rect 5107 4371 5179 4419
rect 5107 4325 5120 4371
rect 5166 4325 5179 4371
rect 5107 4277 5179 4325
rect 5107 4231 5120 4277
rect 5166 4231 5179 4277
rect 5107 4183 5179 4231
rect 5107 4137 5120 4183
rect 5166 4137 5179 4183
rect 2945 4043 2958 4089
rect 3004 4043 3017 4089
rect 2945 3995 3017 4043
rect 2945 3949 2958 3995
rect 3004 3949 3017 3995
rect 2945 3901 3017 3949
rect 2945 3855 2958 3901
rect 3004 3855 3017 3901
rect 2945 3807 3017 3855
rect 2945 3761 2958 3807
rect 3004 3761 3017 3807
rect 2945 3713 3017 3761
rect 5107 4089 5179 4137
rect 5107 4043 5120 4089
rect 5166 4043 5179 4089
rect 5107 3995 5179 4043
rect 5107 3949 5120 3995
rect 5166 3949 5179 3995
rect 5107 3901 5179 3949
rect 5107 3855 5120 3901
rect 5166 3855 5179 3901
rect 5107 3807 5179 3855
rect 5107 3761 5120 3807
rect 5166 3761 5179 3807
rect 2945 3667 2958 3713
rect 3004 3667 3017 3713
rect 2945 3619 3017 3667
rect 2945 3573 2958 3619
rect 3004 3573 3017 3619
rect 2945 3525 3017 3573
rect 2945 3479 2958 3525
rect 3004 3479 3017 3525
rect 2945 3431 3017 3479
rect 2945 3385 2958 3431
rect 3004 3385 3017 3431
rect 2945 3337 3017 3385
rect 2945 3291 2958 3337
rect 3004 3291 3017 3337
rect 2945 3243 3017 3291
rect 2945 3197 2958 3243
rect 3004 3197 3017 3243
rect 2945 3149 3017 3197
rect 2945 3103 2958 3149
rect 3004 3103 3017 3149
rect 2945 3055 3017 3103
rect 2945 3009 2958 3055
rect 3004 3009 3017 3055
rect 2945 2961 3017 3009
rect 5107 3713 5179 3761
rect 5107 3667 5120 3713
rect 5166 3667 5179 3713
rect 5107 3619 5179 3667
rect 5107 3573 5120 3619
rect 5166 3573 5179 3619
rect 5107 3525 5179 3573
rect 5107 3479 5120 3525
rect 5166 3479 5179 3525
rect 5107 3431 5179 3479
rect 5107 3385 5120 3431
rect 5166 3385 5179 3431
rect 5107 3337 5179 3385
rect 5107 3291 5120 3337
rect 5166 3291 5179 3337
rect 5107 3243 5179 3291
rect 5107 3197 5120 3243
rect 5166 3197 5179 3243
rect 5107 3149 5179 3197
rect 5107 3103 5120 3149
rect 5166 3103 5179 3149
rect 5107 3055 5179 3103
rect 5107 3009 5120 3055
rect 5166 3009 5179 3055
rect 2945 2915 2958 2961
rect 3004 2915 3017 2961
rect 2945 2867 3017 2915
rect 2945 2821 2958 2867
rect 3004 2821 3017 2867
rect 2945 2773 3017 2821
rect 2945 2727 2958 2773
rect 3004 2727 3017 2773
rect 2945 2679 3017 2727
rect 2945 2633 2958 2679
rect 3004 2633 3017 2679
rect 2945 2585 3017 2633
rect 5107 2961 5179 3009
rect 5107 2915 5120 2961
rect 5166 2915 5179 2961
rect 5107 2867 5179 2915
rect 5107 2821 5120 2867
rect 5166 2821 5179 2867
rect 5107 2773 5179 2821
rect 5107 2727 5120 2773
rect 5166 2727 5179 2773
rect 5107 2679 5179 2727
rect 5107 2633 5120 2679
rect 5166 2633 5179 2679
rect 2945 2539 2958 2585
rect 3004 2539 3017 2585
rect 2945 2491 3017 2539
rect 2945 2445 2958 2491
rect 3004 2445 3017 2491
rect 2945 2397 3017 2445
rect 2945 2351 2958 2397
rect 3004 2351 3017 2397
rect 2945 2303 3017 2351
rect 2945 2257 2958 2303
rect 3004 2257 3017 2303
rect 2945 2209 3017 2257
rect 2945 2163 2958 2209
rect 3004 2163 3017 2209
rect 2945 2115 3017 2163
rect 2945 2069 2958 2115
rect 3004 2069 3017 2115
rect 2945 2021 3017 2069
rect 2945 1975 2958 2021
rect 3004 1975 3017 2021
rect 2945 1927 3017 1975
rect 2945 1881 2958 1927
rect 3004 1881 3017 1927
rect 2945 1833 3017 1881
rect 5107 2585 5179 2633
rect 5107 2539 5120 2585
rect 5166 2539 5179 2585
rect 5107 2491 5179 2539
rect 5107 2445 5120 2491
rect 5166 2445 5179 2491
rect 5107 2397 5179 2445
rect 5107 2351 5120 2397
rect 5166 2351 5179 2397
rect 5107 2303 5179 2351
rect 5107 2257 5120 2303
rect 5166 2257 5179 2303
rect 5107 2209 5179 2257
rect 5107 2163 5120 2209
rect 5166 2163 5179 2209
rect 5107 2115 5179 2163
rect 5107 2069 5120 2115
rect 5166 2069 5179 2115
rect 5107 2021 5179 2069
rect 5107 1975 5120 2021
rect 5166 1975 5179 2021
rect 5107 1927 5179 1975
rect 5107 1881 5120 1927
rect 5166 1881 5179 1927
rect 2945 1787 2958 1833
rect 3004 1787 3017 1833
rect 2945 1752 3017 1787
rect 31 1739 3017 1752
rect 31 1693 44 1739
rect 90 1693 138 1739
rect 184 1693 232 1739
rect 278 1693 326 1739
rect 372 1693 420 1739
rect 466 1693 514 1739
rect 560 1693 608 1739
rect 654 1693 702 1739
rect 748 1693 796 1739
rect 842 1693 890 1739
rect 936 1693 984 1739
rect 1030 1693 1078 1739
rect 1124 1693 1172 1739
rect 1218 1693 1266 1739
rect 1312 1693 1360 1739
rect 1406 1693 1454 1739
rect 1500 1693 1548 1739
rect 1594 1693 1642 1739
rect 1688 1693 1736 1739
rect 1782 1693 1830 1739
rect 1876 1693 1924 1739
rect 1970 1693 2018 1739
rect 2064 1693 2112 1739
rect 2158 1693 2206 1739
rect 2252 1693 2300 1739
rect 2346 1693 2394 1739
rect 2440 1693 2488 1739
rect 2534 1693 2582 1739
rect 2628 1693 2676 1739
rect 2722 1693 2770 1739
rect 2816 1693 2864 1739
rect 2910 1693 2958 1739
rect 3004 1693 3017 1739
rect 31 1680 3017 1693
rect 31 1645 103 1680
rect 31 1599 44 1645
rect 90 1599 103 1645
rect 31 1551 103 1599
rect 31 1505 44 1551
rect 90 1505 103 1551
rect 31 1457 103 1505
rect 31 1411 44 1457
rect 90 1411 103 1457
rect 31 1363 103 1411
rect 31 1317 44 1363
rect 90 1317 103 1363
rect 31 1269 103 1317
rect 31 1223 44 1269
rect 90 1223 103 1269
rect 31 1175 103 1223
rect 31 1129 44 1175
rect 90 1129 103 1175
rect 31 1081 103 1129
rect 31 1035 44 1081
rect 90 1035 103 1081
rect 31 987 103 1035
rect 31 941 44 987
rect 90 941 103 987
rect 31 893 103 941
rect 31 847 44 893
rect 90 847 103 893
rect 31 799 103 847
rect 31 753 44 799
rect 90 753 103 799
rect 2945 1645 3017 1680
rect 2945 1599 2958 1645
rect 3004 1599 3017 1645
rect 2945 1551 3017 1599
rect 2945 1505 2958 1551
rect 3004 1505 3017 1551
rect 2945 1457 3017 1505
rect 5107 1833 5179 1881
rect 5107 1787 5120 1833
rect 5166 1787 5179 1833
rect 5107 1739 5179 1787
rect 5107 1693 5120 1739
rect 5166 1693 5179 1739
rect 5107 1645 5179 1693
rect 5107 1599 5120 1645
rect 5166 1599 5179 1645
rect 5107 1551 5179 1599
rect 5107 1505 5120 1551
rect 5166 1505 5179 1551
rect 2945 1411 2958 1457
rect 3004 1411 3017 1457
rect 2945 1363 3017 1411
rect 2945 1317 2958 1363
rect 3004 1317 3017 1363
rect 2945 1269 3017 1317
rect 2945 1223 2958 1269
rect 3004 1223 3017 1269
rect 2945 1175 3017 1223
rect 2945 1129 2958 1175
rect 3004 1129 3017 1175
rect 2945 1081 3017 1129
rect 2945 1035 2958 1081
rect 3004 1035 3017 1081
rect 2945 987 3017 1035
rect 2945 941 2958 987
rect 3004 941 3017 987
rect 2945 893 3017 941
rect 2945 847 2958 893
rect 3004 847 3017 893
rect 2945 799 3017 847
rect 31 705 103 753
rect 31 659 44 705
rect 90 659 103 705
rect 31 611 103 659
rect 2945 753 2958 799
rect 3004 753 3017 799
rect 2945 705 3017 753
rect 5107 1457 5179 1505
rect 5107 1411 5120 1457
rect 5166 1411 5179 1457
rect 5107 1363 5179 1411
rect 5107 1317 5120 1363
rect 5166 1317 5179 1363
rect 5107 1269 5179 1317
rect 5107 1223 5120 1269
rect 5166 1223 5179 1269
rect 5107 1175 5179 1223
rect 5107 1129 5120 1175
rect 5166 1129 5179 1175
rect 5107 1081 5179 1129
rect 5107 1035 5120 1081
rect 5166 1035 5179 1081
rect 5107 987 5179 1035
rect 5107 941 5120 987
rect 5166 941 5179 987
rect 5107 893 5179 941
rect 5107 847 5120 893
rect 5166 847 5179 893
rect 5107 799 5179 847
rect 5107 753 5120 799
rect 5166 753 5179 799
rect 2945 659 2958 705
rect 3004 659 3017 705
rect 31 565 44 611
rect 90 565 103 611
rect 31 517 103 565
rect 31 471 44 517
rect 90 471 103 517
rect 31 423 103 471
rect 31 377 44 423
rect 90 377 103 423
rect 31 329 103 377
rect 31 283 44 329
rect 90 283 103 329
rect 31 235 103 283
rect 31 189 44 235
rect 90 189 103 235
rect 31 141 103 189
rect 31 95 44 141
rect 90 95 103 141
rect 31 47 103 95
rect 31 1 44 47
rect 90 1 103 47
rect 2945 611 3017 659
rect 2945 565 2958 611
rect 3004 565 3017 611
rect 2945 517 3017 565
rect 2945 471 2958 517
rect 3004 471 3017 517
rect 2945 423 3017 471
rect 2945 377 2958 423
rect 3004 377 3017 423
rect 2945 329 3017 377
rect 5107 705 5179 753
rect 5107 659 5120 705
rect 5166 659 5179 705
rect 5107 611 5179 659
rect 5107 565 5120 611
rect 5166 565 5179 611
rect 5107 517 5179 565
rect 5107 471 5120 517
rect 5166 471 5179 517
rect 5107 423 5179 471
rect 5107 377 5120 423
rect 5166 377 5179 423
rect 2945 283 2958 329
rect 3004 283 3017 329
rect 2945 235 3017 283
rect 2945 189 2958 235
rect 3004 189 3017 235
rect 2945 141 3017 189
rect 2945 95 2958 141
rect 3004 95 3017 141
rect 2945 47 3017 95
rect 31 -47 103 1
rect 31 -93 44 -47
rect 90 -93 103 -47
rect 31 -141 103 -93
rect 2945 1 2958 47
rect 3004 1 3017 47
rect 2945 -47 3017 1
rect 2945 -93 2958 -47
rect 3004 -93 3017 -47
rect 31 -187 44 -141
rect 90 -187 103 -141
rect 31 -235 103 -187
rect 31 -281 44 -235
rect 90 -281 103 -235
rect 31 -329 103 -281
rect 31 -375 44 -329
rect 90 -375 103 -329
rect 31 -423 103 -375
rect 31 -469 44 -423
rect 90 -469 103 -423
rect 31 -517 103 -469
rect 31 -563 44 -517
rect 90 -563 103 -517
rect 31 -611 103 -563
rect 31 -657 44 -611
rect 90 -657 103 -611
rect 31 -705 103 -657
rect 31 -751 44 -705
rect 90 -751 103 -705
rect 2945 -141 3017 -93
rect 2945 -187 2958 -141
rect 3004 -187 3017 -141
rect 2945 -235 3017 -187
rect 2945 -281 2958 -235
rect 3004 -281 3017 -235
rect 2945 -329 3017 -281
rect 2945 -375 2958 -329
rect 3004 -375 3017 -329
rect 2945 -423 3017 -375
rect 5107 329 5179 377
rect 5107 283 5120 329
rect 5166 283 5179 329
rect 5107 235 5179 283
rect 5107 189 5120 235
rect 5166 189 5179 235
rect 5107 141 5179 189
rect 5107 95 5120 141
rect 5166 95 5179 141
rect 5107 47 5179 95
rect 5107 1 5120 47
rect 5166 1 5179 47
rect 5107 -47 5179 1
rect 5107 -93 5120 -47
rect 5166 -93 5179 -47
rect 5107 -141 5179 -93
rect 5107 -187 5120 -141
rect 5166 -187 5179 -141
rect 5107 -235 5179 -187
rect 5107 -281 5120 -235
rect 5166 -281 5179 -235
rect 5107 -329 5179 -281
rect 5107 -375 5120 -329
rect 5166 -375 5179 -329
rect 2945 -469 2958 -423
rect 3004 -469 3017 -423
rect 2945 -517 3017 -469
rect 2945 -563 2958 -517
rect 3004 -563 3017 -517
rect 2945 -611 3017 -563
rect 2945 -657 2958 -611
rect 3004 -657 3017 -611
rect 5107 -423 5179 -375
rect 5107 -469 5120 -423
rect 5166 -469 5179 -423
rect 5107 -517 5179 -469
rect 2945 -705 3017 -657
rect 31 -799 103 -751
rect 31 -845 44 -799
rect 90 -845 103 -799
rect 31 -893 103 -845
rect 2945 -751 2958 -705
rect 3004 -751 3017 -705
rect 2945 -799 3017 -751
rect 5107 -563 5120 -517
rect 5166 -563 5179 -517
rect 5107 -611 5179 -563
rect 5107 -657 5120 -611
rect 5166 -657 5179 -611
rect 5107 -705 5179 -657
rect 5107 -751 5120 -705
rect 5166 -751 5179 -705
rect 2945 -845 2958 -799
rect 3004 -845 3017 -799
rect 31 -939 44 -893
rect 90 -939 103 -893
rect 31 -987 103 -939
rect 31 -1033 44 -987
rect 90 -1033 103 -987
rect 31 -1081 103 -1033
rect 31 -1127 44 -1081
rect 90 -1127 103 -1081
rect 31 -1175 103 -1127
rect 31 -1221 44 -1175
rect 90 -1221 103 -1175
rect 31 -1269 103 -1221
rect 31 -1315 44 -1269
rect 90 -1315 103 -1269
rect 31 -1363 103 -1315
rect 31 -1409 44 -1363
rect 90 -1409 103 -1363
rect 31 -1457 103 -1409
rect 31 -1503 44 -1457
rect 90 -1503 103 -1457
rect 31 -1551 103 -1503
rect 2945 -893 3017 -845
rect 2945 -939 2958 -893
rect 3004 -939 3017 -893
rect 2945 -987 3017 -939
rect 2945 -1033 2958 -987
rect 3004 -1033 3017 -987
rect 2945 -1081 3017 -1033
rect 2945 -1127 2958 -1081
rect 3004 -1127 3017 -1081
rect 2945 -1175 3017 -1127
rect 2945 -1221 2958 -1175
rect 3004 -1221 3017 -1175
rect 2945 -1269 3017 -1221
rect 2945 -1315 2958 -1269
rect 3004 -1315 3017 -1269
rect 2945 -1363 3017 -1315
rect 2945 -1409 2958 -1363
rect 3004 -1409 3017 -1363
rect 2945 -1457 3017 -1409
rect 2945 -1503 2958 -1457
rect 3004 -1503 3017 -1457
rect 31 -1597 44 -1551
rect 90 -1597 103 -1551
rect 31 -1645 103 -1597
rect 2945 -1551 3017 -1503
rect 5107 -799 5179 -751
rect 5107 -845 5120 -799
rect 5166 -845 5179 -799
rect 5107 -893 5179 -845
rect 5107 -939 5120 -893
rect 5166 -939 5179 -893
rect 5107 -987 5179 -939
rect 5107 -1033 5120 -987
rect 5166 -1033 5179 -987
rect 5107 -1081 5179 -1033
rect 5107 -1127 5120 -1081
rect 5166 -1127 5179 -1081
rect 5107 -1175 5179 -1127
rect 5107 -1221 5120 -1175
rect 5166 -1221 5179 -1175
rect 5107 -1269 5179 -1221
rect 5107 -1315 5120 -1269
rect 5166 -1315 5179 -1269
rect 5107 -1363 5179 -1315
rect 5107 -1409 5120 -1363
rect 5166 -1409 5179 -1363
rect 5107 -1457 5179 -1409
rect 5107 -1503 5120 -1457
rect 5166 -1503 5179 -1457
rect 2945 -1597 2958 -1551
rect 3004 -1597 3017 -1551
rect 31 -1691 44 -1645
rect 90 -1691 103 -1645
rect 31 -1739 103 -1691
rect 31 -1785 44 -1739
rect 90 -1785 103 -1739
rect 31 -1820 103 -1785
rect 2945 -1645 3017 -1597
rect 2945 -1691 2958 -1645
rect 3004 -1691 3017 -1645
rect 5107 -1551 5179 -1503
rect 5107 -1597 5120 -1551
rect 5166 -1597 5179 -1551
rect 5107 -1645 5179 -1597
rect 2945 -1739 3017 -1691
rect 5107 -1691 5120 -1645
rect 5166 -1691 5179 -1645
rect 2945 -1785 2958 -1739
rect 3004 -1785 3017 -1739
rect 2945 -1820 3017 -1785
rect 5107 -1739 5179 -1691
rect 5107 -1785 5120 -1739
rect 5166 -1785 5179 -1739
rect 5107 -1820 5179 -1785
rect 31 -1833 5179 -1820
rect 31 -1879 44 -1833
rect 90 -1879 138 -1833
rect 184 -1879 232 -1833
rect 278 -1879 326 -1833
rect 372 -1879 420 -1833
rect 466 -1879 514 -1833
rect 560 -1879 608 -1833
rect 654 -1879 702 -1833
rect 748 -1879 796 -1833
rect 842 -1879 890 -1833
rect 936 -1879 984 -1833
rect 1030 -1879 1078 -1833
rect 1124 -1879 1172 -1833
rect 1218 -1879 1266 -1833
rect 1312 -1879 1360 -1833
rect 1406 -1879 1454 -1833
rect 1500 -1879 1548 -1833
rect 1594 -1879 1642 -1833
rect 1688 -1879 1736 -1833
rect 1782 -1879 1830 -1833
rect 1876 -1879 1924 -1833
rect 1970 -1879 2018 -1833
rect 2064 -1879 2112 -1833
rect 2158 -1879 2206 -1833
rect 2252 -1879 2300 -1833
rect 2346 -1879 2394 -1833
rect 2440 -1879 2488 -1833
rect 2534 -1879 2582 -1833
rect 2628 -1879 2676 -1833
rect 2722 -1879 2770 -1833
rect 2816 -1879 2864 -1833
rect 2910 -1879 2958 -1833
rect 3004 -1879 3052 -1833
rect 3098 -1879 3146 -1833
rect 3192 -1879 3240 -1833
rect 3286 -1879 3334 -1833
rect 3380 -1879 3428 -1833
rect 3474 -1879 3522 -1833
rect 3568 -1879 3616 -1833
rect 3662 -1879 3710 -1833
rect 3756 -1879 3804 -1833
rect 3850 -1879 3898 -1833
rect 3944 -1879 3992 -1833
rect 4038 -1879 4086 -1833
rect 4132 -1879 4180 -1833
rect 4226 -1879 4274 -1833
rect 4320 -1879 4368 -1833
rect 4414 -1879 4462 -1833
rect 4508 -1879 4556 -1833
rect 4602 -1879 4650 -1833
rect 4696 -1879 4744 -1833
rect 4790 -1879 4838 -1833
rect 4884 -1879 4932 -1833
rect 4978 -1879 5026 -1833
rect 5072 -1879 5120 -1833
rect 5166 -1879 5179 -1833
rect 31 -1892 5179 -1879
rect 11401 2585 16549 2598
rect 11401 2539 11414 2585
rect 11460 2539 11508 2585
rect 11554 2539 11602 2585
rect 11648 2539 11696 2585
rect 11742 2539 11790 2585
rect 11836 2539 11884 2585
rect 11930 2539 11978 2585
rect 12024 2539 12072 2585
rect 12118 2539 12166 2585
rect 12212 2539 12260 2585
rect 12306 2539 12354 2585
rect 12400 2539 12448 2585
rect 12494 2539 12542 2585
rect 12588 2539 12636 2585
rect 12682 2539 12730 2585
rect 12776 2539 12824 2585
rect 12870 2539 12918 2585
rect 12964 2539 13012 2585
rect 13058 2539 13106 2585
rect 13152 2539 13200 2585
rect 13246 2539 13294 2585
rect 13340 2539 13388 2585
rect 13434 2539 13482 2585
rect 13528 2539 13576 2585
rect 13622 2539 13670 2585
rect 13716 2539 13764 2585
rect 13810 2539 13858 2585
rect 13904 2539 13952 2585
rect 13998 2539 14046 2585
rect 14092 2539 14140 2585
rect 14186 2539 14234 2585
rect 14280 2539 14328 2585
rect 14374 2539 14422 2585
rect 14468 2539 14516 2585
rect 14562 2539 14610 2585
rect 14656 2539 14704 2585
rect 14750 2539 14798 2585
rect 14844 2539 14892 2585
rect 14938 2539 14986 2585
rect 15032 2539 15080 2585
rect 15126 2539 15174 2585
rect 15220 2539 15268 2585
rect 15314 2539 15362 2585
rect 15408 2539 15456 2585
rect 15502 2539 15550 2585
rect 15596 2539 15644 2585
rect 15690 2539 15738 2585
rect 15784 2539 15832 2585
rect 15878 2539 15926 2585
rect 15972 2539 16020 2585
rect 16066 2539 16114 2585
rect 16160 2539 16208 2585
rect 16254 2539 16302 2585
rect 16348 2539 16396 2585
rect 16442 2539 16490 2585
rect 16536 2539 16549 2585
rect 11401 2526 16549 2539
rect 11401 2491 11473 2526
rect 11401 2445 11414 2491
rect 11460 2445 11473 2491
rect 11401 2397 11473 2445
rect 11401 2351 11414 2397
rect 11460 2351 11473 2397
rect 11401 2303 11473 2351
rect 11401 2257 11414 2303
rect 11460 2257 11473 2303
rect 11401 2209 11473 2257
rect 11401 2163 11414 2209
rect 11460 2163 11473 2209
rect 11401 2115 11473 2163
rect 11401 2069 11414 2115
rect 11460 2069 11473 2115
rect 11401 2021 11473 2069
rect 11401 1975 11414 2021
rect 11460 1975 11473 2021
rect 11401 1927 11473 1975
rect 11401 1881 11414 1927
rect 11460 1881 11473 1927
rect 11401 1833 11473 1881
rect 11401 1787 11414 1833
rect 11460 1787 11473 1833
rect 11401 1739 11473 1787
rect 11401 1693 11414 1739
rect 11460 1693 11473 1739
rect 11401 1645 11473 1693
rect 11401 1599 11414 1645
rect 11460 1599 11473 1645
rect 11401 1551 11473 1599
rect 14127 2491 14199 2526
rect 14127 2445 14140 2491
rect 14186 2445 14199 2491
rect 14127 2397 14199 2445
rect 14127 2351 14140 2397
rect 14186 2351 14199 2397
rect 14127 2303 14199 2351
rect 14127 2257 14140 2303
rect 14186 2257 14199 2303
rect 14127 2209 14199 2257
rect 14127 2163 14140 2209
rect 14186 2163 14199 2209
rect 14127 2115 14199 2163
rect 14127 2069 14140 2115
rect 14186 2069 14199 2115
rect 14127 2021 14199 2069
rect 14127 1975 14140 2021
rect 14186 1975 14199 2021
rect 14127 1927 14199 1975
rect 14127 1881 14140 1927
rect 14186 1881 14199 1927
rect 14127 1833 14199 1881
rect 14127 1787 14140 1833
rect 14186 1787 14199 1833
rect 14127 1739 14199 1787
rect 14127 1693 14140 1739
rect 14186 1693 14199 1739
rect 14127 1645 14199 1693
rect 14127 1599 14140 1645
rect 14186 1599 14199 1645
rect 11401 1505 11414 1551
rect 11460 1505 11473 1551
rect 11401 1457 11473 1505
rect 11401 1411 11414 1457
rect 11460 1411 11473 1457
rect 11401 1363 11473 1411
rect 11401 1317 11414 1363
rect 11460 1317 11473 1363
rect 11401 1269 11473 1317
rect 11401 1223 11414 1269
rect 11460 1223 11473 1269
rect 11401 1175 11473 1223
rect 14127 1551 14199 1599
rect 16477 2491 16549 2526
rect 16477 2445 16490 2491
rect 16536 2445 16549 2491
rect 16477 2397 16549 2445
rect 16477 2351 16490 2397
rect 16536 2351 16549 2397
rect 16477 2303 16549 2351
rect 16477 2257 16490 2303
rect 16536 2257 16549 2303
rect 16477 2209 16549 2257
rect 16477 2163 16490 2209
rect 16536 2163 16549 2209
rect 16477 2115 16549 2163
rect 16477 2069 16490 2115
rect 16536 2069 16549 2115
rect 16477 2021 16549 2069
rect 16477 1975 16490 2021
rect 16536 1975 16549 2021
rect 16477 1927 16549 1975
rect 16477 1881 16490 1927
rect 16536 1881 16549 1927
rect 16477 1833 16549 1881
rect 16477 1787 16490 1833
rect 16536 1787 16549 1833
rect 16477 1739 16549 1787
rect 16477 1693 16490 1739
rect 16536 1693 16549 1739
rect 16477 1645 16549 1693
rect 16477 1599 16490 1645
rect 16536 1599 16549 1645
rect 14127 1505 14140 1551
rect 14186 1505 14199 1551
rect 14127 1457 14199 1505
rect 14127 1411 14140 1457
rect 14186 1411 14199 1457
rect 14127 1363 14199 1411
rect 14127 1317 14140 1363
rect 14186 1317 14199 1363
rect 14127 1269 14199 1317
rect 14127 1223 14140 1269
rect 14186 1223 14199 1269
rect 11401 1129 11414 1175
rect 11460 1129 11473 1175
rect 11401 1081 11473 1129
rect 11401 1035 11414 1081
rect 11460 1035 11473 1081
rect 11401 987 11473 1035
rect 11401 941 11414 987
rect 11460 941 11473 987
rect 11401 893 11473 941
rect 11401 847 11414 893
rect 11460 847 11473 893
rect 11401 799 11473 847
rect 11401 753 11414 799
rect 11460 753 11473 799
rect 11401 705 11473 753
rect 11401 659 11414 705
rect 11460 659 11473 705
rect 11401 611 11473 659
rect 11401 565 11414 611
rect 11460 565 11473 611
rect 11401 517 11473 565
rect 14127 1175 14199 1223
rect 16477 1551 16549 1599
rect 16477 1505 16490 1551
rect 16536 1505 16549 1551
rect 16477 1457 16549 1505
rect 16477 1411 16490 1457
rect 16536 1411 16549 1457
rect 16477 1363 16549 1411
rect 16477 1317 16490 1363
rect 16536 1317 16549 1363
rect 16477 1269 16549 1317
rect 16477 1223 16490 1269
rect 16536 1223 16549 1269
rect 14127 1129 14140 1175
rect 14186 1129 14199 1175
rect 14127 1081 14199 1129
rect 14127 1035 14140 1081
rect 14186 1035 14199 1081
rect 14127 987 14199 1035
rect 14127 941 14140 987
rect 14186 941 14199 987
rect 14127 893 14199 941
rect 14127 847 14140 893
rect 14186 847 14199 893
rect 14127 799 14199 847
rect 14127 753 14140 799
rect 14186 753 14199 799
rect 14127 705 14199 753
rect 14127 659 14140 705
rect 14186 659 14199 705
rect 14127 611 14199 659
rect 14127 565 14140 611
rect 14186 565 14199 611
rect 11401 471 11414 517
rect 11460 471 11473 517
rect 11401 423 11473 471
rect 11401 377 11414 423
rect 11460 377 11473 423
rect 11401 329 11473 377
rect 11401 283 11414 329
rect 11460 283 11473 329
rect 11401 235 11473 283
rect 11401 189 11414 235
rect 11460 189 11473 235
rect 11401 141 11473 189
rect 14127 517 14199 565
rect 16477 1175 16549 1223
rect 16477 1129 16490 1175
rect 16536 1129 16549 1175
rect 16477 1081 16549 1129
rect 16477 1035 16490 1081
rect 16536 1035 16549 1081
rect 16477 987 16549 1035
rect 16477 941 16490 987
rect 16536 941 16549 987
rect 16477 893 16549 941
rect 16477 847 16490 893
rect 16536 847 16549 893
rect 16477 799 16549 847
rect 16477 753 16490 799
rect 16536 753 16549 799
rect 16477 705 16549 753
rect 16477 659 16490 705
rect 16536 659 16549 705
rect 16477 611 16549 659
rect 16477 565 16490 611
rect 16536 565 16549 611
rect 14127 471 14140 517
rect 14186 471 14199 517
rect 14127 423 14199 471
rect 14127 377 14140 423
rect 14186 377 14199 423
rect 14127 329 14199 377
rect 14127 283 14140 329
rect 14186 283 14199 329
rect 14127 235 14199 283
rect 14127 189 14140 235
rect 14186 189 14199 235
rect 11401 95 11414 141
rect 11460 95 11473 141
rect 11401 47 11473 95
rect 11401 1 11414 47
rect 11460 1 11473 47
rect 11401 -47 11473 1
rect 11401 -93 11414 -47
rect 11460 -93 11473 -47
rect 11401 -141 11473 -93
rect 11401 -187 11414 -141
rect 11460 -187 11473 -141
rect 11401 -235 11473 -187
rect 11401 -281 11414 -235
rect 11460 -281 11473 -235
rect 11401 -329 11473 -281
rect 11401 -375 11414 -329
rect 11460 -375 11473 -329
rect 11401 -423 11473 -375
rect 11401 -469 11414 -423
rect 11460 -469 11473 -423
rect 11401 -517 11473 -469
rect 14127 141 14199 189
rect 16477 517 16549 565
rect 16477 471 16490 517
rect 16536 471 16549 517
rect 16477 423 16549 471
rect 16477 377 16490 423
rect 16536 377 16549 423
rect 16477 329 16549 377
rect 16477 283 16490 329
rect 16536 283 16549 329
rect 16477 235 16549 283
rect 16477 189 16490 235
rect 16536 189 16549 235
rect 14127 95 14140 141
rect 14186 95 14199 141
rect 14127 47 14199 95
rect 14127 1 14140 47
rect 14186 1 14199 47
rect 14127 -47 14199 1
rect 14127 -93 14140 -47
rect 14186 -93 14199 -47
rect 14127 -141 14199 -93
rect 14127 -187 14140 -141
rect 14186 -187 14199 -141
rect 14127 -235 14199 -187
rect 14127 -281 14140 -235
rect 14186 -281 14199 -235
rect 14127 -329 14199 -281
rect 14127 -375 14140 -329
rect 14186 -375 14199 -329
rect 14127 -423 14199 -375
rect 14127 -469 14140 -423
rect 14186 -469 14199 -423
rect 11401 -563 11414 -517
rect 11460 -563 11473 -517
rect 11401 -611 11473 -563
rect 11401 -657 11414 -611
rect 11460 -657 11473 -611
rect 11401 -705 11473 -657
rect 11401 -751 11414 -705
rect 11460 -751 11473 -705
rect 11401 -799 11473 -751
rect 14127 -517 14199 -469
rect 16477 141 16549 189
rect 16477 95 16490 141
rect 16536 95 16549 141
rect 16477 47 16549 95
rect 16477 1 16490 47
rect 16536 1 16549 47
rect 16477 -47 16549 1
rect 16477 -93 16490 -47
rect 16536 -93 16549 -47
rect 16477 -141 16549 -93
rect 16477 -187 16490 -141
rect 16536 -187 16549 -141
rect 16477 -235 16549 -187
rect 16477 -281 16490 -235
rect 16536 -281 16549 -235
rect 16477 -329 16549 -281
rect 16477 -375 16490 -329
rect 16536 -375 16549 -329
rect 16477 -423 16549 -375
rect 16477 -469 16490 -423
rect 16536 -469 16549 -423
rect 14127 -563 14140 -517
rect 14186 -563 14199 -517
rect 14127 -611 14199 -563
rect 14127 -657 14140 -611
rect 14186 -657 14199 -611
rect 14127 -705 14199 -657
rect 11401 -845 11414 -799
rect 11460 -845 11473 -799
rect 11401 -893 11473 -845
rect 14127 -751 14140 -705
rect 14186 -751 14199 -705
rect 14127 -799 14199 -751
rect 16477 -517 16549 -469
rect 16477 -563 16490 -517
rect 16536 -563 16549 -517
rect 16477 -611 16549 -563
rect 16477 -657 16490 -611
rect 16536 -657 16549 -611
rect 16477 -705 16549 -657
rect 14127 -845 14140 -799
rect 14186 -845 14199 -799
rect 11401 -939 11414 -893
rect 11460 -939 11473 -893
rect 11401 -987 11473 -939
rect 11401 -1033 11414 -987
rect 11460 -1033 11473 -987
rect 11401 -1081 11473 -1033
rect 11401 -1127 11414 -1081
rect 11460 -1127 11473 -1081
rect 11401 -1175 11473 -1127
rect 11401 -1221 11414 -1175
rect 11460 -1221 11473 -1175
rect 11401 -1269 11473 -1221
rect 11401 -1315 11414 -1269
rect 11460 -1315 11473 -1269
rect 11401 -1363 11473 -1315
rect 11401 -1409 11414 -1363
rect 11460 -1409 11473 -1363
rect 11401 -1457 11473 -1409
rect 11401 -1503 11414 -1457
rect 11460 -1503 11473 -1457
rect 11401 -1551 11473 -1503
rect 11401 -1597 11414 -1551
rect 11460 -1597 11473 -1551
rect 11401 -1645 11473 -1597
rect 11401 -1691 11414 -1645
rect 11460 -1691 11473 -1645
rect 11401 -1739 11473 -1691
rect 11401 -1785 11414 -1739
rect 11460 -1785 11473 -1739
rect 11401 -1820 11473 -1785
rect 14127 -893 14199 -845
rect 16477 -751 16490 -705
rect 16536 -751 16549 -705
rect 16477 -799 16549 -751
rect 16477 -845 16490 -799
rect 16536 -845 16549 -799
rect 14127 -939 14140 -893
rect 14186 -939 14199 -893
rect 14127 -987 14199 -939
rect 14127 -1033 14140 -987
rect 14186 -1033 14199 -987
rect 14127 -1081 14199 -1033
rect 14127 -1127 14140 -1081
rect 14186 -1127 14199 -1081
rect 14127 -1175 14199 -1127
rect 14127 -1221 14140 -1175
rect 14186 -1221 14199 -1175
rect 14127 -1269 14199 -1221
rect 14127 -1315 14140 -1269
rect 14186 -1315 14199 -1269
rect 14127 -1363 14199 -1315
rect 14127 -1409 14140 -1363
rect 14186 -1409 14199 -1363
rect 14127 -1457 14199 -1409
rect 14127 -1503 14140 -1457
rect 14186 -1503 14199 -1457
rect 14127 -1551 14199 -1503
rect 14127 -1597 14140 -1551
rect 14186 -1597 14199 -1551
rect 14127 -1645 14199 -1597
rect 14127 -1691 14140 -1645
rect 14186 -1691 14199 -1645
rect 14127 -1739 14199 -1691
rect 14127 -1785 14140 -1739
rect 14186 -1785 14199 -1739
rect 14127 -1820 14199 -1785
rect 16477 -893 16549 -845
rect 16477 -939 16490 -893
rect 16536 -939 16549 -893
rect 16477 -987 16549 -939
rect 16477 -1033 16490 -987
rect 16536 -1033 16549 -987
rect 16477 -1081 16549 -1033
rect 16477 -1127 16490 -1081
rect 16536 -1127 16549 -1081
rect 16477 -1175 16549 -1127
rect 16477 -1221 16490 -1175
rect 16536 -1221 16549 -1175
rect 16477 -1269 16549 -1221
rect 16477 -1315 16490 -1269
rect 16536 -1315 16549 -1269
rect 16477 -1363 16549 -1315
rect 16477 -1409 16490 -1363
rect 16536 -1409 16549 -1363
rect 16477 -1457 16549 -1409
rect 16477 -1503 16490 -1457
rect 16536 -1503 16549 -1457
rect 16477 -1551 16549 -1503
rect 16477 -1597 16490 -1551
rect 16536 -1597 16549 -1551
rect 16477 -1645 16549 -1597
rect 16477 -1691 16490 -1645
rect 16536 -1691 16549 -1645
rect 16477 -1739 16549 -1691
rect 16477 -1785 16490 -1739
rect 16536 -1785 16549 -1739
rect 16477 -1820 16549 -1785
rect 11401 -1833 16549 -1820
rect 11401 -1879 11414 -1833
rect 11460 -1879 11508 -1833
rect 11554 -1879 11602 -1833
rect 11648 -1879 11696 -1833
rect 11742 -1879 11790 -1833
rect 11836 -1879 11884 -1833
rect 11930 -1879 11978 -1833
rect 12024 -1879 12072 -1833
rect 12118 -1879 12166 -1833
rect 12212 -1879 12260 -1833
rect 12306 -1879 12354 -1833
rect 12400 -1879 12448 -1833
rect 12494 -1879 12542 -1833
rect 12588 -1879 12636 -1833
rect 12682 -1879 12730 -1833
rect 12776 -1879 12824 -1833
rect 12870 -1879 12918 -1833
rect 12964 -1879 13012 -1833
rect 13058 -1879 13106 -1833
rect 13152 -1879 13200 -1833
rect 13246 -1879 13294 -1833
rect 13340 -1879 13388 -1833
rect 13434 -1879 13482 -1833
rect 13528 -1879 13576 -1833
rect 13622 -1879 13670 -1833
rect 13716 -1879 13764 -1833
rect 13810 -1879 13858 -1833
rect 13904 -1879 13952 -1833
rect 13998 -1879 14046 -1833
rect 14092 -1879 14140 -1833
rect 14186 -1879 14234 -1833
rect 14280 -1879 14328 -1833
rect 14374 -1879 14422 -1833
rect 14468 -1879 14516 -1833
rect 14562 -1879 14610 -1833
rect 14656 -1879 14704 -1833
rect 14750 -1879 14798 -1833
rect 14844 -1879 14892 -1833
rect 14938 -1879 14986 -1833
rect 15032 -1879 15080 -1833
rect 15126 -1879 15174 -1833
rect 15220 -1879 15268 -1833
rect 15314 -1879 15362 -1833
rect 15408 -1879 15456 -1833
rect 15502 -1879 15550 -1833
rect 15596 -1879 15644 -1833
rect 15690 -1879 15738 -1833
rect 15784 -1879 15832 -1833
rect 15878 -1879 15926 -1833
rect 15972 -1879 16020 -1833
rect 16066 -1879 16114 -1833
rect 16160 -1879 16208 -1833
rect 16254 -1879 16302 -1833
rect 16348 -1879 16396 -1833
rect 16442 -1879 16490 -1833
rect 16536 -1879 16549 -1833
rect 32130 3062 40474 3075
rect 32130 3016 32143 3062
rect 32189 3016 32237 3062
rect 32283 3016 32331 3062
rect 32377 3016 32425 3062
rect 32471 3016 32519 3062
rect 32565 3016 32613 3062
rect 32659 3016 32707 3062
rect 32753 3016 32801 3062
rect 32847 3016 32895 3062
rect 32941 3016 32989 3062
rect 33035 3016 33083 3062
rect 33129 3016 33177 3062
rect 33223 3016 33271 3062
rect 33317 3016 33365 3062
rect 33411 3016 33459 3062
rect 33505 3016 33553 3062
rect 33599 3016 33647 3062
rect 33693 3016 33741 3062
rect 33787 3016 33835 3062
rect 33881 3016 33929 3062
rect 33975 3016 34023 3062
rect 34069 3016 34117 3062
rect 34163 3016 34211 3062
rect 34257 3016 34305 3062
rect 34351 3016 34399 3062
rect 34445 3016 34493 3062
rect 34539 3016 34587 3062
rect 34633 3016 34681 3062
rect 34727 3016 34775 3062
rect 34821 3016 34869 3062
rect 34915 3016 34963 3062
rect 35009 3016 35057 3062
rect 35103 3016 35151 3062
rect 35197 3016 35245 3062
rect 35291 3016 35339 3062
rect 35385 3016 35433 3062
rect 35479 3016 35527 3062
rect 35573 3016 35621 3062
rect 35667 3016 35715 3062
rect 35761 3016 35809 3062
rect 35855 3016 35903 3062
rect 35949 3016 35997 3062
rect 36043 3016 36091 3062
rect 36137 3016 36185 3062
rect 36231 3016 36279 3062
rect 36325 3016 36373 3062
rect 36419 3016 36467 3062
rect 36513 3016 36561 3062
rect 36607 3016 36655 3062
rect 36701 3016 36749 3062
rect 36795 3016 36843 3062
rect 36889 3016 36937 3062
rect 36983 3016 37031 3062
rect 37077 3016 37125 3062
rect 37171 3016 37219 3062
rect 37265 3016 37313 3062
rect 37359 3016 37407 3062
rect 37453 3016 37501 3062
rect 37547 3016 37595 3062
rect 37641 3016 37689 3062
rect 37735 3016 37783 3062
rect 37829 3016 37877 3062
rect 37923 3016 37971 3062
rect 38017 3016 38065 3062
rect 38111 3016 38159 3062
rect 38205 3016 38253 3062
rect 38299 3016 38347 3062
rect 38393 3016 38441 3062
rect 38487 3016 38535 3062
rect 38581 3016 38629 3062
rect 38675 3016 38723 3062
rect 38769 3016 38817 3062
rect 38863 3016 38911 3062
rect 38957 3016 39005 3062
rect 39051 3016 39099 3062
rect 39145 3016 39193 3062
rect 39239 3016 39287 3062
rect 39333 3016 39381 3062
rect 39427 3016 39475 3062
rect 39521 3016 39569 3062
rect 39615 3016 39663 3062
rect 39709 3016 39757 3062
rect 39803 3016 39851 3062
rect 39897 3016 39945 3062
rect 39991 3016 40039 3062
rect 40085 3016 40133 3062
rect 40179 3016 40227 3062
rect 40273 3016 40321 3062
rect 40367 3016 40415 3062
rect 40461 3016 40474 3062
rect 32130 3003 40474 3016
rect 32130 2968 32202 3003
rect 32130 2922 32143 2968
rect 32189 2922 32202 2968
rect 32130 2874 32202 2922
rect 32130 2828 32143 2874
rect 32189 2828 32202 2874
rect 32130 2780 32202 2828
rect 32130 2734 32143 2780
rect 32189 2734 32202 2780
rect 32130 2686 32202 2734
rect 32130 2640 32143 2686
rect 32189 2640 32202 2686
rect 36266 2968 36338 3003
rect 36266 2922 36279 2968
rect 36325 2922 36338 2968
rect 36266 2874 36338 2922
rect 36266 2828 36279 2874
rect 36325 2828 36338 2874
rect 36266 2780 36338 2828
rect 36266 2734 36279 2780
rect 36325 2734 36338 2780
rect 36266 2686 36338 2734
rect 32130 2592 32202 2640
rect 36266 2640 36279 2686
rect 36325 2640 36338 2686
rect 40402 2968 40474 3003
rect 40402 2922 40415 2968
rect 40461 2922 40474 2968
rect 40402 2874 40474 2922
rect 40402 2828 40415 2874
rect 40461 2828 40474 2874
rect 40402 2780 40474 2828
rect 40402 2734 40415 2780
rect 40461 2734 40474 2780
rect 40402 2686 40474 2734
rect 32130 2546 32143 2592
rect 32189 2546 32202 2592
rect 32130 2498 32202 2546
rect 36266 2592 36338 2640
rect 40402 2640 40415 2686
rect 40461 2640 40474 2686
rect 36266 2546 36279 2592
rect 36325 2546 36338 2592
rect 32130 2452 32143 2498
rect 32189 2452 32202 2498
rect 32130 2404 32202 2452
rect 32130 2358 32143 2404
rect 32189 2358 32202 2404
rect 32130 2310 32202 2358
rect 32130 2264 32143 2310
rect 32189 2264 32202 2310
rect 32130 2216 32202 2264
rect 32130 2170 32143 2216
rect 32189 2170 32202 2216
rect 32130 2122 32202 2170
rect 32130 2076 32143 2122
rect 32189 2076 32202 2122
rect 32130 2028 32202 2076
rect 32130 1982 32143 2028
rect 32189 1982 32202 2028
rect 32130 1934 32202 1982
rect 32130 1888 32143 1934
rect 32189 1888 32202 1934
rect 36266 2498 36338 2546
rect 40402 2592 40474 2640
rect 40402 2546 40415 2592
rect 40461 2546 40474 2592
rect 36266 2452 36279 2498
rect 36325 2452 36338 2498
rect 36266 2404 36338 2452
rect 36266 2358 36279 2404
rect 36325 2358 36338 2404
rect 36266 2310 36338 2358
rect 36266 2264 36279 2310
rect 36325 2264 36338 2310
rect 36266 2216 36338 2264
rect 36266 2170 36279 2216
rect 36325 2170 36338 2216
rect 36266 2122 36338 2170
rect 36266 2076 36279 2122
rect 36325 2076 36338 2122
rect 36266 2028 36338 2076
rect 36266 1982 36279 2028
rect 36325 1982 36338 2028
rect 36266 1934 36338 1982
rect 32130 1840 32202 1888
rect 32130 1794 32143 1840
rect 32189 1794 32202 1840
rect 32130 1746 32202 1794
rect 32130 1700 32143 1746
rect 32189 1700 32202 1746
rect 32130 1652 32202 1700
rect 32130 1606 32143 1652
rect 32189 1606 32202 1652
rect 32130 1558 32202 1606
rect 32130 1512 32143 1558
rect 32189 1512 32202 1558
rect 32130 1464 32202 1512
rect 32130 1418 32143 1464
rect 32189 1418 32202 1464
rect 32130 1370 32202 1418
rect 32130 1324 32143 1370
rect 32189 1324 32202 1370
rect 32130 1276 32202 1324
rect 32130 1230 32143 1276
rect 32189 1230 32202 1276
rect 32130 1182 32202 1230
rect 32130 1136 32143 1182
rect 32189 1136 32202 1182
rect 32130 1088 32202 1136
rect 32130 1042 32143 1088
rect 32189 1042 32202 1088
rect 32130 994 32202 1042
rect 32130 948 32143 994
rect 32189 948 32202 994
rect 32130 900 32202 948
rect 32130 854 32143 900
rect 32189 854 32202 900
rect 32130 806 32202 854
rect 32130 760 32143 806
rect 32189 760 32202 806
rect 32130 712 32202 760
rect 32130 666 32143 712
rect 32189 666 32202 712
rect 32130 618 32202 666
rect 32130 572 32143 618
rect 32189 572 32202 618
rect 32130 524 32202 572
rect 32130 478 32143 524
rect 32189 478 32202 524
rect 32130 430 32202 478
rect 32130 384 32143 430
rect 32189 384 32202 430
rect 32130 336 32202 384
rect 32130 290 32143 336
rect 32189 290 32202 336
rect 32130 242 32202 290
rect 32130 196 32143 242
rect 32189 196 32202 242
rect 32130 148 32202 196
rect 32130 102 32143 148
rect 32189 102 32202 148
rect 32130 54 32202 102
rect 32130 8 32143 54
rect 32189 8 32202 54
rect 32130 -40 32202 8
rect 32130 -86 32143 -40
rect 32189 -86 32202 -40
rect 32130 -134 32202 -86
rect 32130 -180 32143 -134
rect 32189 -180 32202 -134
rect 32130 -228 32202 -180
rect 32130 -274 32143 -228
rect 32189 -274 32202 -228
rect 32130 -322 32202 -274
rect 32130 -368 32143 -322
rect 32189 -368 32202 -322
rect 32130 -416 32202 -368
rect 36266 1888 36279 1934
rect 36325 1888 36338 1934
rect 40402 2498 40474 2546
rect 40402 2452 40415 2498
rect 40461 2452 40474 2498
rect 40402 2404 40474 2452
rect 40402 2358 40415 2404
rect 40461 2358 40474 2404
rect 40402 2310 40474 2358
rect 40402 2264 40415 2310
rect 40461 2264 40474 2310
rect 40402 2216 40474 2264
rect 40402 2170 40415 2216
rect 40461 2170 40474 2216
rect 40402 2122 40474 2170
rect 40402 2076 40415 2122
rect 40461 2076 40474 2122
rect 40402 2028 40474 2076
rect 40402 1982 40415 2028
rect 40461 1982 40474 2028
rect 40402 1934 40474 1982
rect 36266 1840 36338 1888
rect 36266 1794 36279 1840
rect 36325 1794 36338 1840
rect 36266 1746 36338 1794
rect 36266 1700 36279 1746
rect 36325 1700 36338 1746
rect 32130 -462 32143 -416
rect 32189 -462 32202 -416
rect 32130 -510 32202 -462
rect 32130 -556 32143 -510
rect 32189 -556 32202 -510
rect 32130 -604 32202 -556
rect 32130 -650 32143 -604
rect 32189 -650 32202 -604
rect 36266 1652 36338 1700
rect 36266 1606 36279 1652
rect 36325 1606 36338 1652
rect 36266 1558 36338 1606
rect 36266 1512 36279 1558
rect 36325 1512 36338 1558
rect 36266 1464 36338 1512
rect 36266 1418 36279 1464
rect 36325 1418 36338 1464
rect 36266 1370 36338 1418
rect 36266 1324 36279 1370
rect 36325 1324 36338 1370
rect 36266 1276 36338 1324
rect 36266 1230 36279 1276
rect 36325 1230 36338 1276
rect 36266 1182 36338 1230
rect 36266 1136 36279 1182
rect 36325 1136 36338 1182
rect 36266 1088 36338 1136
rect 36266 1042 36279 1088
rect 36325 1042 36338 1088
rect 36266 994 36338 1042
rect 36266 948 36279 994
rect 36325 948 36338 994
rect 36266 900 36338 948
rect 36266 854 36279 900
rect 36325 854 36338 900
rect 36266 806 36338 854
rect 36266 760 36279 806
rect 36325 760 36338 806
rect 36266 712 36338 760
rect 36266 666 36279 712
rect 36325 666 36338 712
rect 36266 618 36338 666
rect 36266 572 36279 618
rect 36325 572 36338 618
rect 36266 524 36338 572
rect 36266 478 36279 524
rect 36325 478 36338 524
rect 36266 430 36338 478
rect 36266 384 36279 430
rect 36325 384 36338 430
rect 36266 336 36338 384
rect 36266 290 36279 336
rect 36325 290 36338 336
rect 36266 242 36338 290
rect 36266 196 36279 242
rect 36325 196 36338 242
rect 36266 148 36338 196
rect 36266 102 36279 148
rect 36325 102 36338 148
rect 36266 54 36338 102
rect 36266 8 36279 54
rect 36325 8 36338 54
rect 36266 -40 36338 8
rect 36266 -86 36279 -40
rect 36325 -86 36338 -40
rect 36266 -134 36338 -86
rect 36266 -180 36279 -134
rect 36325 -180 36338 -134
rect 36266 -228 36338 -180
rect 36266 -274 36279 -228
rect 36325 -274 36338 -228
rect 36266 -322 36338 -274
rect 36266 -368 36279 -322
rect 36325 -368 36338 -322
rect 36266 -416 36338 -368
rect 40402 1888 40415 1934
rect 40461 1888 40474 1934
rect 40402 1840 40474 1888
rect 40402 1794 40415 1840
rect 40461 1794 40474 1840
rect 40402 1746 40474 1794
rect 40402 1700 40415 1746
rect 40461 1700 40474 1746
rect 36266 -462 36279 -416
rect 36325 -462 36338 -416
rect 36266 -510 36338 -462
rect 36266 -556 36279 -510
rect 36325 -556 36338 -510
rect 36266 -604 36338 -556
rect 32130 -698 32202 -650
rect 32130 -744 32143 -698
rect 32189 -744 32202 -698
rect 32130 -792 32202 -744
rect 32130 -838 32143 -792
rect 32189 -838 32202 -792
rect 32130 -886 32202 -838
rect 32130 -932 32143 -886
rect 32189 -932 32202 -886
rect 32130 -980 32202 -932
rect 32130 -1026 32143 -980
rect 32189 -1026 32202 -980
rect 32130 -1074 32202 -1026
rect 32130 -1120 32143 -1074
rect 32189 -1120 32202 -1074
rect 32130 -1168 32202 -1120
rect 32130 -1214 32143 -1168
rect 32189 -1214 32202 -1168
rect 32130 -1262 32202 -1214
rect 32130 -1308 32143 -1262
rect 32189 -1308 32202 -1262
rect 32130 -1356 32202 -1308
rect 32130 -1402 32143 -1356
rect 32189 -1402 32202 -1356
rect 32130 -1450 32202 -1402
rect 32130 -1496 32143 -1450
rect 32189 -1496 32202 -1450
rect 32130 -1544 32202 -1496
rect 32130 -1590 32143 -1544
rect 32189 -1590 32202 -1544
rect 32130 -1638 32202 -1590
rect 32130 -1684 32143 -1638
rect 32189 -1684 32202 -1638
rect 32130 -1719 32202 -1684
rect 36266 -650 36279 -604
rect 36325 -650 36338 -604
rect 40402 1652 40474 1700
rect 40402 1606 40415 1652
rect 40461 1606 40474 1652
rect 40402 1558 40474 1606
rect 40402 1512 40415 1558
rect 40461 1512 40474 1558
rect 40402 1464 40474 1512
rect 40402 1418 40415 1464
rect 40461 1418 40474 1464
rect 40402 1370 40474 1418
rect 40402 1324 40415 1370
rect 40461 1324 40474 1370
rect 40402 1276 40474 1324
rect 40402 1230 40415 1276
rect 40461 1230 40474 1276
rect 40402 1182 40474 1230
rect 40402 1136 40415 1182
rect 40461 1136 40474 1182
rect 40402 1088 40474 1136
rect 40402 1042 40415 1088
rect 40461 1042 40474 1088
rect 40402 994 40474 1042
rect 40402 948 40415 994
rect 40461 948 40474 994
rect 40402 900 40474 948
rect 40402 854 40415 900
rect 40461 854 40474 900
rect 40402 806 40474 854
rect 40402 760 40415 806
rect 40461 760 40474 806
rect 40402 712 40474 760
rect 40402 666 40415 712
rect 40461 666 40474 712
rect 40402 618 40474 666
rect 40402 572 40415 618
rect 40461 572 40474 618
rect 40402 524 40474 572
rect 40402 478 40415 524
rect 40461 478 40474 524
rect 40402 430 40474 478
rect 40402 384 40415 430
rect 40461 384 40474 430
rect 40402 336 40474 384
rect 40402 290 40415 336
rect 40461 290 40474 336
rect 40402 242 40474 290
rect 40402 196 40415 242
rect 40461 196 40474 242
rect 40402 148 40474 196
rect 40402 102 40415 148
rect 40461 102 40474 148
rect 40402 54 40474 102
rect 40402 8 40415 54
rect 40461 8 40474 54
rect 40402 -40 40474 8
rect 40402 -86 40415 -40
rect 40461 -86 40474 -40
rect 40402 -134 40474 -86
rect 40402 -180 40415 -134
rect 40461 -180 40474 -134
rect 40402 -228 40474 -180
rect 40402 -274 40415 -228
rect 40461 -274 40474 -228
rect 40402 -322 40474 -274
rect 40402 -368 40415 -322
rect 40461 -368 40474 -322
rect 40402 -416 40474 -368
rect 40402 -462 40415 -416
rect 40461 -462 40474 -416
rect 40402 -510 40474 -462
rect 40402 -556 40415 -510
rect 40461 -556 40474 -510
rect 40402 -604 40474 -556
rect 36266 -698 36338 -650
rect 36266 -744 36279 -698
rect 36325 -744 36338 -698
rect 36266 -792 36338 -744
rect 36266 -838 36279 -792
rect 36325 -838 36338 -792
rect 36266 -886 36338 -838
rect 36266 -932 36279 -886
rect 36325 -932 36338 -886
rect 36266 -980 36338 -932
rect 36266 -1026 36279 -980
rect 36325 -1026 36338 -980
rect 36266 -1074 36338 -1026
rect 36266 -1120 36279 -1074
rect 36325 -1120 36338 -1074
rect 36266 -1168 36338 -1120
rect 36266 -1214 36279 -1168
rect 36325 -1214 36338 -1168
rect 36266 -1262 36338 -1214
rect 36266 -1308 36279 -1262
rect 36325 -1308 36338 -1262
rect 36266 -1356 36338 -1308
rect 36266 -1402 36279 -1356
rect 36325 -1402 36338 -1356
rect 36266 -1450 36338 -1402
rect 36266 -1496 36279 -1450
rect 36325 -1496 36338 -1450
rect 36266 -1544 36338 -1496
rect 36266 -1590 36279 -1544
rect 36325 -1590 36338 -1544
rect 36266 -1638 36338 -1590
rect 36266 -1684 36279 -1638
rect 36325 -1684 36338 -1638
rect 36266 -1719 36338 -1684
rect 40402 -650 40415 -604
rect 40461 -650 40474 -604
rect 40402 -698 40474 -650
rect 40402 -744 40415 -698
rect 40461 -744 40474 -698
rect 40402 -792 40474 -744
rect 40402 -838 40415 -792
rect 40461 -838 40474 -792
rect 40402 -886 40474 -838
rect 40402 -932 40415 -886
rect 40461 -932 40474 -886
rect 40402 -980 40474 -932
rect 40402 -1026 40415 -980
rect 40461 -1026 40474 -980
rect 40402 -1074 40474 -1026
rect 40402 -1120 40415 -1074
rect 40461 -1120 40474 -1074
rect 40402 -1168 40474 -1120
rect 40402 -1214 40415 -1168
rect 40461 -1214 40474 -1168
rect 40402 -1262 40474 -1214
rect 40402 -1308 40415 -1262
rect 40461 -1308 40474 -1262
rect 40402 -1356 40474 -1308
rect 40402 -1402 40415 -1356
rect 40461 -1402 40474 -1356
rect 40402 -1450 40474 -1402
rect 40402 -1496 40415 -1450
rect 40461 -1496 40474 -1450
rect 40402 -1544 40474 -1496
rect 40402 -1590 40415 -1544
rect 40461 -1590 40474 -1544
rect 40402 -1638 40474 -1590
rect 40402 -1684 40415 -1638
rect 40461 -1684 40474 -1638
rect 40402 -1719 40474 -1684
rect 32130 -1732 40474 -1719
rect 32130 -1778 32143 -1732
rect 32189 -1778 32237 -1732
rect 32283 -1778 32331 -1732
rect 32377 -1778 32425 -1732
rect 32471 -1778 32519 -1732
rect 32565 -1778 32613 -1732
rect 32659 -1778 32707 -1732
rect 32753 -1778 32801 -1732
rect 32847 -1778 32895 -1732
rect 32941 -1778 32989 -1732
rect 33035 -1778 33083 -1732
rect 33129 -1778 33177 -1732
rect 33223 -1778 33271 -1732
rect 33317 -1778 33365 -1732
rect 33411 -1778 33459 -1732
rect 33505 -1778 33553 -1732
rect 33599 -1778 33647 -1732
rect 33693 -1778 33741 -1732
rect 33787 -1778 33835 -1732
rect 33881 -1778 33929 -1732
rect 33975 -1778 34023 -1732
rect 34069 -1778 34117 -1732
rect 34163 -1778 34211 -1732
rect 34257 -1778 34305 -1732
rect 34351 -1778 34399 -1732
rect 34445 -1778 34493 -1732
rect 34539 -1778 34587 -1732
rect 34633 -1778 34681 -1732
rect 34727 -1778 34775 -1732
rect 34821 -1778 34869 -1732
rect 34915 -1778 34963 -1732
rect 35009 -1778 35057 -1732
rect 35103 -1778 35151 -1732
rect 35197 -1778 35245 -1732
rect 35291 -1778 35339 -1732
rect 35385 -1778 35433 -1732
rect 35479 -1778 35527 -1732
rect 35573 -1778 35621 -1732
rect 35667 -1778 35715 -1732
rect 35761 -1778 35809 -1732
rect 35855 -1778 35903 -1732
rect 35949 -1778 35997 -1732
rect 36043 -1778 36091 -1732
rect 36137 -1778 36185 -1732
rect 36231 -1778 36279 -1732
rect 36325 -1778 36373 -1732
rect 36419 -1778 36467 -1732
rect 36513 -1778 36561 -1732
rect 36607 -1778 36655 -1732
rect 36701 -1778 36749 -1732
rect 36795 -1778 36843 -1732
rect 36889 -1778 36937 -1732
rect 36983 -1778 37031 -1732
rect 37077 -1778 37125 -1732
rect 37171 -1778 37219 -1732
rect 37265 -1778 37313 -1732
rect 37359 -1778 37407 -1732
rect 37453 -1778 37501 -1732
rect 37547 -1778 37595 -1732
rect 37641 -1778 37689 -1732
rect 37735 -1778 37783 -1732
rect 37829 -1778 37877 -1732
rect 37923 -1778 37971 -1732
rect 38017 -1778 38065 -1732
rect 38111 -1778 38159 -1732
rect 38205 -1778 38253 -1732
rect 38299 -1778 38347 -1732
rect 38393 -1778 38441 -1732
rect 38487 -1778 38535 -1732
rect 38581 -1778 38629 -1732
rect 38675 -1778 38723 -1732
rect 38769 -1778 38817 -1732
rect 38863 -1778 38911 -1732
rect 38957 -1778 39005 -1732
rect 39051 -1778 39099 -1732
rect 39145 -1778 39193 -1732
rect 39239 -1778 39287 -1732
rect 39333 -1778 39381 -1732
rect 39427 -1778 39475 -1732
rect 39521 -1778 39569 -1732
rect 39615 -1778 39663 -1732
rect 39709 -1778 39757 -1732
rect 39803 -1778 39851 -1732
rect 39897 -1778 39945 -1732
rect 39991 -1778 40039 -1732
rect 40085 -1778 40133 -1732
rect 40179 -1778 40227 -1732
rect 40273 -1778 40321 -1732
rect 40367 -1778 40415 -1732
rect 40461 -1778 40474 -1732
rect 32130 -1791 40474 -1778
rect 41826 3062 50170 3075
rect 41826 3016 41839 3062
rect 41885 3016 41933 3062
rect 41979 3016 42027 3062
rect 42073 3016 42121 3062
rect 42167 3016 42215 3062
rect 42261 3016 42309 3062
rect 42355 3016 42403 3062
rect 42449 3016 42497 3062
rect 42543 3016 42591 3062
rect 42637 3016 42685 3062
rect 42731 3016 42779 3062
rect 42825 3016 42873 3062
rect 42919 3016 42967 3062
rect 43013 3016 43061 3062
rect 43107 3016 43155 3062
rect 43201 3016 43249 3062
rect 43295 3016 43343 3062
rect 43389 3016 43437 3062
rect 43483 3016 43531 3062
rect 43577 3016 43625 3062
rect 43671 3016 43719 3062
rect 43765 3016 43813 3062
rect 43859 3016 43907 3062
rect 43953 3016 44001 3062
rect 44047 3016 44095 3062
rect 44141 3016 44189 3062
rect 44235 3016 44283 3062
rect 44329 3016 44377 3062
rect 44423 3016 44471 3062
rect 44517 3016 44565 3062
rect 44611 3016 44659 3062
rect 44705 3016 44753 3062
rect 44799 3016 44847 3062
rect 44893 3016 44941 3062
rect 44987 3016 45035 3062
rect 45081 3016 45129 3062
rect 45175 3016 45223 3062
rect 45269 3016 45317 3062
rect 45363 3016 45411 3062
rect 45457 3016 45505 3062
rect 45551 3016 45599 3062
rect 45645 3016 45693 3062
rect 45739 3016 45787 3062
rect 45833 3016 45881 3062
rect 45927 3016 45975 3062
rect 46021 3016 46069 3062
rect 46115 3016 46163 3062
rect 46209 3016 46257 3062
rect 46303 3016 46351 3062
rect 46397 3016 46445 3062
rect 46491 3016 46539 3062
rect 46585 3016 46633 3062
rect 46679 3016 46727 3062
rect 46773 3016 46821 3062
rect 46867 3016 46915 3062
rect 46961 3016 47009 3062
rect 47055 3016 47103 3062
rect 47149 3016 47197 3062
rect 47243 3016 47291 3062
rect 47337 3016 47385 3062
rect 47431 3016 47479 3062
rect 47525 3016 47573 3062
rect 47619 3016 47667 3062
rect 47713 3016 47761 3062
rect 47807 3016 47855 3062
rect 47901 3016 47949 3062
rect 47995 3016 48043 3062
rect 48089 3016 48137 3062
rect 48183 3016 48231 3062
rect 48277 3016 48325 3062
rect 48371 3016 48419 3062
rect 48465 3016 48513 3062
rect 48559 3016 48607 3062
rect 48653 3016 48701 3062
rect 48747 3016 48795 3062
rect 48841 3016 48889 3062
rect 48935 3016 48983 3062
rect 49029 3016 49077 3062
rect 49123 3016 49171 3062
rect 49217 3016 49265 3062
rect 49311 3016 49359 3062
rect 49405 3016 49453 3062
rect 49499 3016 49547 3062
rect 49593 3016 49641 3062
rect 49687 3016 49735 3062
rect 49781 3016 49829 3062
rect 49875 3016 49923 3062
rect 49969 3016 50017 3062
rect 50063 3016 50111 3062
rect 50157 3016 50170 3062
rect 41826 3003 50170 3016
rect 41826 2968 41898 3003
rect 41826 2922 41839 2968
rect 41885 2922 41898 2968
rect 41826 2874 41898 2922
rect 41826 2828 41839 2874
rect 41885 2828 41898 2874
rect 41826 2780 41898 2828
rect 41826 2734 41839 2780
rect 41885 2734 41898 2780
rect 41826 2686 41898 2734
rect 41826 2640 41839 2686
rect 41885 2640 41898 2686
rect 45962 2968 46034 3003
rect 45962 2922 45975 2968
rect 46021 2922 46034 2968
rect 45962 2874 46034 2922
rect 45962 2828 45975 2874
rect 46021 2828 46034 2874
rect 45962 2780 46034 2828
rect 45962 2734 45975 2780
rect 46021 2734 46034 2780
rect 45962 2686 46034 2734
rect 41826 2592 41898 2640
rect 45962 2640 45975 2686
rect 46021 2640 46034 2686
rect 50098 2968 50170 3003
rect 50098 2922 50111 2968
rect 50157 2922 50170 2968
rect 50098 2874 50170 2922
rect 50098 2828 50111 2874
rect 50157 2828 50170 2874
rect 50098 2780 50170 2828
rect 50098 2734 50111 2780
rect 50157 2734 50170 2780
rect 50098 2686 50170 2734
rect 41826 2546 41839 2592
rect 41885 2546 41898 2592
rect 41826 2498 41898 2546
rect 45962 2592 46034 2640
rect 50098 2640 50111 2686
rect 50157 2640 50170 2686
rect 45962 2546 45975 2592
rect 46021 2546 46034 2592
rect 41826 2452 41839 2498
rect 41885 2452 41898 2498
rect 41826 2404 41898 2452
rect 41826 2358 41839 2404
rect 41885 2358 41898 2404
rect 41826 2310 41898 2358
rect 41826 2264 41839 2310
rect 41885 2264 41898 2310
rect 41826 2216 41898 2264
rect 41826 2170 41839 2216
rect 41885 2170 41898 2216
rect 41826 2122 41898 2170
rect 41826 2076 41839 2122
rect 41885 2076 41898 2122
rect 41826 2028 41898 2076
rect 41826 1982 41839 2028
rect 41885 1982 41898 2028
rect 41826 1934 41898 1982
rect 41826 1888 41839 1934
rect 41885 1888 41898 1934
rect 45962 2498 46034 2546
rect 50098 2592 50170 2640
rect 50098 2546 50111 2592
rect 50157 2546 50170 2592
rect 45962 2452 45975 2498
rect 46021 2452 46034 2498
rect 45962 2404 46034 2452
rect 45962 2358 45975 2404
rect 46021 2358 46034 2404
rect 45962 2310 46034 2358
rect 45962 2264 45975 2310
rect 46021 2264 46034 2310
rect 45962 2216 46034 2264
rect 45962 2170 45975 2216
rect 46021 2170 46034 2216
rect 45962 2122 46034 2170
rect 45962 2076 45975 2122
rect 46021 2076 46034 2122
rect 45962 2028 46034 2076
rect 45962 1982 45975 2028
rect 46021 1982 46034 2028
rect 45962 1934 46034 1982
rect 41826 1840 41898 1888
rect 41826 1794 41839 1840
rect 41885 1794 41898 1840
rect 41826 1746 41898 1794
rect 41826 1700 41839 1746
rect 41885 1700 41898 1746
rect 41826 1652 41898 1700
rect 41826 1606 41839 1652
rect 41885 1606 41898 1652
rect 41826 1558 41898 1606
rect 41826 1512 41839 1558
rect 41885 1512 41898 1558
rect 41826 1464 41898 1512
rect 41826 1418 41839 1464
rect 41885 1418 41898 1464
rect 41826 1370 41898 1418
rect 41826 1324 41839 1370
rect 41885 1324 41898 1370
rect 41826 1276 41898 1324
rect 41826 1230 41839 1276
rect 41885 1230 41898 1276
rect 41826 1182 41898 1230
rect 41826 1136 41839 1182
rect 41885 1136 41898 1182
rect 41826 1088 41898 1136
rect 41826 1042 41839 1088
rect 41885 1042 41898 1088
rect 41826 994 41898 1042
rect 41826 948 41839 994
rect 41885 948 41898 994
rect 41826 900 41898 948
rect 41826 854 41839 900
rect 41885 854 41898 900
rect 41826 806 41898 854
rect 41826 760 41839 806
rect 41885 760 41898 806
rect 41826 712 41898 760
rect 41826 666 41839 712
rect 41885 666 41898 712
rect 41826 618 41898 666
rect 41826 572 41839 618
rect 41885 572 41898 618
rect 41826 524 41898 572
rect 41826 478 41839 524
rect 41885 478 41898 524
rect 41826 430 41898 478
rect 41826 384 41839 430
rect 41885 384 41898 430
rect 41826 336 41898 384
rect 41826 290 41839 336
rect 41885 290 41898 336
rect 41826 242 41898 290
rect 41826 196 41839 242
rect 41885 196 41898 242
rect 41826 148 41898 196
rect 41826 102 41839 148
rect 41885 102 41898 148
rect 41826 54 41898 102
rect 41826 8 41839 54
rect 41885 8 41898 54
rect 41826 -40 41898 8
rect 41826 -86 41839 -40
rect 41885 -86 41898 -40
rect 41826 -134 41898 -86
rect 41826 -180 41839 -134
rect 41885 -180 41898 -134
rect 41826 -228 41898 -180
rect 41826 -274 41839 -228
rect 41885 -274 41898 -228
rect 41826 -322 41898 -274
rect 41826 -368 41839 -322
rect 41885 -368 41898 -322
rect 41826 -416 41898 -368
rect 45962 1888 45975 1934
rect 46021 1888 46034 1934
rect 50098 2498 50170 2546
rect 50098 2452 50111 2498
rect 50157 2452 50170 2498
rect 50098 2404 50170 2452
rect 50098 2358 50111 2404
rect 50157 2358 50170 2404
rect 50098 2310 50170 2358
rect 50098 2264 50111 2310
rect 50157 2264 50170 2310
rect 50098 2216 50170 2264
rect 50098 2170 50111 2216
rect 50157 2170 50170 2216
rect 50098 2122 50170 2170
rect 50098 2076 50111 2122
rect 50157 2076 50170 2122
rect 50098 2028 50170 2076
rect 50098 1982 50111 2028
rect 50157 1982 50170 2028
rect 50098 1934 50170 1982
rect 45962 1840 46034 1888
rect 45962 1794 45975 1840
rect 46021 1794 46034 1840
rect 45962 1746 46034 1794
rect 45962 1700 45975 1746
rect 46021 1700 46034 1746
rect 41826 -462 41839 -416
rect 41885 -462 41898 -416
rect 41826 -510 41898 -462
rect 41826 -556 41839 -510
rect 41885 -556 41898 -510
rect 41826 -604 41898 -556
rect 41826 -650 41839 -604
rect 41885 -650 41898 -604
rect 45962 1652 46034 1700
rect 45962 1606 45975 1652
rect 46021 1606 46034 1652
rect 45962 1558 46034 1606
rect 45962 1512 45975 1558
rect 46021 1512 46034 1558
rect 45962 1464 46034 1512
rect 45962 1418 45975 1464
rect 46021 1418 46034 1464
rect 45962 1370 46034 1418
rect 45962 1324 45975 1370
rect 46021 1324 46034 1370
rect 45962 1276 46034 1324
rect 45962 1230 45975 1276
rect 46021 1230 46034 1276
rect 45962 1182 46034 1230
rect 45962 1136 45975 1182
rect 46021 1136 46034 1182
rect 45962 1088 46034 1136
rect 45962 1042 45975 1088
rect 46021 1042 46034 1088
rect 45962 994 46034 1042
rect 45962 948 45975 994
rect 46021 948 46034 994
rect 45962 900 46034 948
rect 45962 854 45975 900
rect 46021 854 46034 900
rect 45962 806 46034 854
rect 45962 760 45975 806
rect 46021 760 46034 806
rect 45962 712 46034 760
rect 45962 666 45975 712
rect 46021 666 46034 712
rect 45962 618 46034 666
rect 45962 572 45975 618
rect 46021 572 46034 618
rect 45962 524 46034 572
rect 45962 478 45975 524
rect 46021 478 46034 524
rect 45962 430 46034 478
rect 45962 384 45975 430
rect 46021 384 46034 430
rect 45962 336 46034 384
rect 45962 290 45975 336
rect 46021 290 46034 336
rect 45962 242 46034 290
rect 45962 196 45975 242
rect 46021 196 46034 242
rect 45962 148 46034 196
rect 45962 102 45975 148
rect 46021 102 46034 148
rect 45962 54 46034 102
rect 45962 8 45975 54
rect 46021 8 46034 54
rect 45962 -40 46034 8
rect 45962 -86 45975 -40
rect 46021 -86 46034 -40
rect 45962 -134 46034 -86
rect 45962 -180 45975 -134
rect 46021 -180 46034 -134
rect 45962 -228 46034 -180
rect 45962 -274 45975 -228
rect 46021 -274 46034 -228
rect 45962 -322 46034 -274
rect 45962 -368 45975 -322
rect 46021 -368 46034 -322
rect 45962 -416 46034 -368
rect 50098 1888 50111 1934
rect 50157 1888 50170 1934
rect 50098 1840 50170 1888
rect 50098 1794 50111 1840
rect 50157 1794 50170 1840
rect 50098 1746 50170 1794
rect 50098 1700 50111 1746
rect 50157 1700 50170 1746
rect 45962 -462 45975 -416
rect 46021 -462 46034 -416
rect 45962 -510 46034 -462
rect 45962 -556 45975 -510
rect 46021 -556 46034 -510
rect 45962 -604 46034 -556
rect 41826 -698 41898 -650
rect 41826 -744 41839 -698
rect 41885 -744 41898 -698
rect 41826 -792 41898 -744
rect 41826 -838 41839 -792
rect 41885 -838 41898 -792
rect 41826 -886 41898 -838
rect 41826 -932 41839 -886
rect 41885 -932 41898 -886
rect 41826 -980 41898 -932
rect 41826 -1026 41839 -980
rect 41885 -1026 41898 -980
rect 41826 -1074 41898 -1026
rect 41826 -1120 41839 -1074
rect 41885 -1120 41898 -1074
rect 41826 -1168 41898 -1120
rect 41826 -1214 41839 -1168
rect 41885 -1214 41898 -1168
rect 41826 -1262 41898 -1214
rect 41826 -1308 41839 -1262
rect 41885 -1308 41898 -1262
rect 41826 -1356 41898 -1308
rect 41826 -1402 41839 -1356
rect 41885 -1402 41898 -1356
rect 41826 -1450 41898 -1402
rect 41826 -1496 41839 -1450
rect 41885 -1496 41898 -1450
rect 41826 -1544 41898 -1496
rect 41826 -1590 41839 -1544
rect 41885 -1590 41898 -1544
rect 41826 -1638 41898 -1590
rect 41826 -1684 41839 -1638
rect 41885 -1684 41898 -1638
rect 41826 -1719 41898 -1684
rect 45962 -650 45975 -604
rect 46021 -650 46034 -604
rect 50098 1652 50170 1700
rect 50098 1606 50111 1652
rect 50157 1606 50170 1652
rect 50098 1558 50170 1606
rect 50098 1512 50111 1558
rect 50157 1512 50170 1558
rect 50098 1464 50170 1512
rect 50098 1418 50111 1464
rect 50157 1418 50170 1464
rect 50098 1370 50170 1418
rect 50098 1324 50111 1370
rect 50157 1324 50170 1370
rect 50098 1276 50170 1324
rect 50098 1230 50111 1276
rect 50157 1230 50170 1276
rect 50098 1182 50170 1230
rect 50098 1136 50111 1182
rect 50157 1136 50170 1182
rect 50098 1088 50170 1136
rect 50098 1042 50111 1088
rect 50157 1042 50170 1088
rect 50098 994 50170 1042
rect 50098 948 50111 994
rect 50157 948 50170 994
rect 50098 900 50170 948
rect 50098 854 50111 900
rect 50157 854 50170 900
rect 50098 806 50170 854
rect 50098 760 50111 806
rect 50157 760 50170 806
rect 50098 712 50170 760
rect 50098 666 50111 712
rect 50157 666 50170 712
rect 50098 618 50170 666
rect 50098 572 50111 618
rect 50157 572 50170 618
rect 50098 524 50170 572
rect 50098 478 50111 524
rect 50157 478 50170 524
rect 50098 430 50170 478
rect 50098 384 50111 430
rect 50157 384 50170 430
rect 50098 336 50170 384
rect 50098 290 50111 336
rect 50157 290 50170 336
rect 50098 242 50170 290
rect 50098 196 50111 242
rect 50157 196 50170 242
rect 50098 148 50170 196
rect 50098 102 50111 148
rect 50157 102 50170 148
rect 50098 54 50170 102
rect 50098 8 50111 54
rect 50157 8 50170 54
rect 50098 -40 50170 8
rect 50098 -86 50111 -40
rect 50157 -86 50170 -40
rect 50098 -134 50170 -86
rect 50098 -180 50111 -134
rect 50157 -180 50170 -134
rect 50098 -228 50170 -180
rect 50098 -274 50111 -228
rect 50157 -274 50170 -228
rect 50098 -322 50170 -274
rect 50098 -368 50111 -322
rect 50157 -368 50170 -322
rect 50098 -416 50170 -368
rect 50098 -462 50111 -416
rect 50157 -462 50170 -416
rect 50098 -510 50170 -462
rect 50098 -556 50111 -510
rect 50157 -556 50170 -510
rect 50098 -604 50170 -556
rect 45962 -698 46034 -650
rect 45962 -744 45975 -698
rect 46021 -744 46034 -698
rect 45962 -792 46034 -744
rect 45962 -838 45975 -792
rect 46021 -838 46034 -792
rect 45962 -886 46034 -838
rect 45962 -932 45975 -886
rect 46021 -932 46034 -886
rect 45962 -980 46034 -932
rect 45962 -1026 45975 -980
rect 46021 -1026 46034 -980
rect 45962 -1074 46034 -1026
rect 45962 -1120 45975 -1074
rect 46021 -1120 46034 -1074
rect 45962 -1168 46034 -1120
rect 45962 -1214 45975 -1168
rect 46021 -1214 46034 -1168
rect 45962 -1262 46034 -1214
rect 45962 -1308 45975 -1262
rect 46021 -1308 46034 -1262
rect 45962 -1356 46034 -1308
rect 45962 -1402 45975 -1356
rect 46021 -1402 46034 -1356
rect 45962 -1450 46034 -1402
rect 45962 -1496 45975 -1450
rect 46021 -1496 46034 -1450
rect 45962 -1544 46034 -1496
rect 45962 -1590 45975 -1544
rect 46021 -1590 46034 -1544
rect 45962 -1638 46034 -1590
rect 45962 -1684 45975 -1638
rect 46021 -1684 46034 -1638
rect 45962 -1719 46034 -1684
rect 50098 -650 50111 -604
rect 50157 -650 50170 -604
rect 50098 -698 50170 -650
rect 50098 -744 50111 -698
rect 50157 -744 50170 -698
rect 50098 -792 50170 -744
rect 50098 -838 50111 -792
rect 50157 -838 50170 -792
rect 50098 -886 50170 -838
rect 50098 -932 50111 -886
rect 50157 -932 50170 -886
rect 50098 -980 50170 -932
rect 50098 -1026 50111 -980
rect 50157 -1026 50170 -980
rect 50098 -1074 50170 -1026
rect 50098 -1120 50111 -1074
rect 50157 -1120 50170 -1074
rect 50098 -1168 50170 -1120
rect 50098 -1214 50111 -1168
rect 50157 -1214 50170 -1168
rect 50098 -1262 50170 -1214
rect 50098 -1308 50111 -1262
rect 50157 -1308 50170 -1262
rect 50098 -1356 50170 -1308
rect 50098 -1402 50111 -1356
rect 50157 -1402 50170 -1356
rect 50098 -1450 50170 -1402
rect 50098 -1496 50111 -1450
rect 50157 -1496 50170 -1450
rect 50098 -1544 50170 -1496
rect 50098 -1590 50111 -1544
rect 50157 -1590 50170 -1544
rect 50098 -1638 50170 -1590
rect 50098 -1684 50111 -1638
rect 50157 -1684 50170 -1638
rect 50098 -1719 50170 -1684
rect 41826 -1732 50170 -1719
rect 41826 -1778 41839 -1732
rect 41885 -1778 41933 -1732
rect 41979 -1778 42027 -1732
rect 42073 -1778 42121 -1732
rect 42167 -1778 42215 -1732
rect 42261 -1778 42309 -1732
rect 42355 -1778 42403 -1732
rect 42449 -1778 42497 -1732
rect 42543 -1778 42591 -1732
rect 42637 -1778 42685 -1732
rect 42731 -1778 42779 -1732
rect 42825 -1778 42873 -1732
rect 42919 -1778 42967 -1732
rect 43013 -1778 43061 -1732
rect 43107 -1778 43155 -1732
rect 43201 -1778 43249 -1732
rect 43295 -1778 43343 -1732
rect 43389 -1778 43437 -1732
rect 43483 -1778 43531 -1732
rect 43577 -1778 43625 -1732
rect 43671 -1778 43719 -1732
rect 43765 -1778 43813 -1732
rect 43859 -1778 43907 -1732
rect 43953 -1778 44001 -1732
rect 44047 -1778 44095 -1732
rect 44141 -1778 44189 -1732
rect 44235 -1778 44283 -1732
rect 44329 -1778 44377 -1732
rect 44423 -1778 44471 -1732
rect 44517 -1778 44565 -1732
rect 44611 -1778 44659 -1732
rect 44705 -1778 44753 -1732
rect 44799 -1778 44847 -1732
rect 44893 -1778 44941 -1732
rect 44987 -1778 45035 -1732
rect 45081 -1778 45129 -1732
rect 45175 -1778 45223 -1732
rect 45269 -1778 45317 -1732
rect 45363 -1778 45411 -1732
rect 45457 -1778 45505 -1732
rect 45551 -1778 45599 -1732
rect 45645 -1778 45693 -1732
rect 45739 -1778 45787 -1732
rect 45833 -1778 45881 -1732
rect 45927 -1778 45975 -1732
rect 46021 -1778 46069 -1732
rect 46115 -1778 46163 -1732
rect 46209 -1778 46257 -1732
rect 46303 -1778 46351 -1732
rect 46397 -1778 46445 -1732
rect 46491 -1778 46539 -1732
rect 46585 -1778 46633 -1732
rect 46679 -1778 46727 -1732
rect 46773 -1778 46821 -1732
rect 46867 -1778 46915 -1732
rect 46961 -1778 47009 -1732
rect 47055 -1778 47103 -1732
rect 47149 -1778 47197 -1732
rect 47243 -1778 47291 -1732
rect 47337 -1778 47385 -1732
rect 47431 -1778 47479 -1732
rect 47525 -1778 47573 -1732
rect 47619 -1778 47667 -1732
rect 47713 -1778 47761 -1732
rect 47807 -1778 47855 -1732
rect 47901 -1778 47949 -1732
rect 47995 -1778 48043 -1732
rect 48089 -1778 48137 -1732
rect 48183 -1778 48231 -1732
rect 48277 -1778 48325 -1732
rect 48371 -1778 48419 -1732
rect 48465 -1778 48513 -1732
rect 48559 -1778 48607 -1732
rect 48653 -1778 48701 -1732
rect 48747 -1778 48795 -1732
rect 48841 -1778 48889 -1732
rect 48935 -1778 48983 -1732
rect 49029 -1778 49077 -1732
rect 49123 -1778 49171 -1732
rect 49217 -1778 49265 -1732
rect 49311 -1778 49359 -1732
rect 49405 -1778 49453 -1732
rect 49499 -1778 49547 -1732
rect 49593 -1778 49641 -1732
rect 49687 -1778 49735 -1732
rect 49781 -1778 49829 -1732
rect 49875 -1778 49923 -1732
rect 49969 -1778 50017 -1732
rect 50063 -1778 50111 -1732
rect 50157 -1778 50170 -1732
rect 41826 -1791 50170 -1778
rect 51522 3062 59866 3075
rect 51522 3016 51535 3062
rect 51581 3016 51629 3062
rect 51675 3016 51723 3062
rect 51769 3016 51817 3062
rect 51863 3016 51911 3062
rect 51957 3016 52005 3062
rect 52051 3016 52099 3062
rect 52145 3016 52193 3062
rect 52239 3016 52287 3062
rect 52333 3016 52381 3062
rect 52427 3016 52475 3062
rect 52521 3016 52569 3062
rect 52615 3016 52663 3062
rect 52709 3016 52757 3062
rect 52803 3016 52851 3062
rect 52897 3016 52945 3062
rect 52991 3016 53039 3062
rect 53085 3016 53133 3062
rect 53179 3016 53227 3062
rect 53273 3016 53321 3062
rect 53367 3016 53415 3062
rect 53461 3016 53509 3062
rect 53555 3016 53603 3062
rect 53649 3016 53697 3062
rect 53743 3016 53791 3062
rect 53837 3016 53885 3062
rect 53931 3016 53979 3062
rect 54025 3016 54073 3062
rect 54119 3016 54167 3062
rect 54213 3016 54261 3062
rect 54307 3016 54355 3062
rect 54401 3016 54449 3062
rect 54495 3016 54543 3062
rect 54589 3016 54637 3062
rect 54683 3016 54731 3062
rect 54777 3016 54825 3062
rect 54871 3016 54919 3062
rect 54965 3016 55013 3062
rect 55059 3016 55107 3062
rect 55153 3016 55201 3062
rect 55247 3016 55295 3062
rect 55341 3016 55389 3062
rect 55435 3016 55483 3062
rect 55529 3016 55577 3062
rect 55623 3016 55671 3062
rect 55717 3016 55765 3062
rect 55811 3016 55859 3062
rect 55905 3016 55953 3062
rect 55999 3016 56047 3062
rect 56093 3016 56141 3062
rect 56187 3016 56235 3062
rect 56281 3016 56329 3062
rect 56375 3016 56423 3062
rect 56469 3016 56517 3062
rect 56563 3016 56611 3062
rect 56657 3016 56705 3062
rect 56751 3016 56799 3062
rect 56845 3016 56893 3062
rect 56939 3016 56987 3062
rect 57033 3016 57081 3062
rect 57127 3016 57175 3062
rect 57221 3016 57269 3062
rect 57315 3016 57363 3062
rect 57409 3016 57457 3062
rect 57503 3016 57551 3062
rect 57597 3016 57645 3062
rect 57691 3016 57739 3062
rect 57785 3016 57833 3062
rect 57879 3016 57927 3062
rect 57973 3016 58021 3062
rect 58067 3016 58115 3062
rect 58161 3016 58209 3062
rect 58255 3016 58303 3062
rect 58349 3016 58397 3062
rect 58443 3016 58491 3062
rect 58537 3016 58585 3062
rect 58631 3016 58679 3062
rect 58725 3016 58773 3062
rect 58819 3016 58867 3062
rect 58913 3016 58961 3062
rect 59007 3016 59055 3062
rect 59101 3016 59149 3062
rect 59195 3016 59243 3062
rect 59289 3016 59337 3062
rect 59383 3016 59431 3062
rect 59477 3016 59525 3062
rect 59571 3016 59619 3062
rect 59665 3016 59713 3062
rect 59759 3016 59807 3062
rect 59853 3016 59866 3062
rect 51522 3003 59866 3016
rect 51522 2968 51594 3003
rect 51522 2922 51535 2968
rect 51581 2922 51594 2968
rect 51522 2874 51594 2922
rect 51522 2828 51535 2874
rect 51581 2828 51594 2874
rect 51522 2780 51594 2828
rect 51522 2734 51535 2780
rect 51581 2734 51594 2780
rect 51522 2686 51594 2734
rect 51522 2640 51535 2686
rect 51581 2640 51594 2686
rect 55658 2968 55730 3003
rect 55658 2922 55671 2968
rect 55717 2922 55730 2968
rect 55658 2874 55730 2922
rect 55658 2828 55671 2874
rect 55717 2828 55730 2874
rect 55658 2780 55730 2828
rect 55658 2734 55671 2780
rect 55717 2734 55730 2780
rect 55658 2686 55730 2734
rect 51522 2592 51594 2640
rect 55658 2640 55671 2686
rect 55717 2640 55730 2686
rect 59794 2968 59866 3003
rect 59794 2922 59807 2968
rect 59853 2922 59866 2968
rect 59794 2874 59866 2922
rect 59794 2828 59807 2874
rect 59853 2828 59866 2874
rect 59794 2780 59866 2828
rect 59794 2734 59807 2780
rect 59853 2734 59866 2780
rect 59794 2686 59866 2734
rect 51522 2546 51535 2592
rect 51581 2546 51594 2592
rect 51522 2498 51594 2546
rect 55658 2592 55730 2640
rect 59794 2640 59807 2686
rect 59853 2640 59866 2686
rect 55658 2546 55671 2592
rect 55717 2546 55730 2592
rect 51522 2452 51535 2498
rect 51581 2452 51594 2498
rect 51522 2404 51594 2452
rect 51522 2358 51535 2404
rect 51581 2358 51594 2404
rect 51522 2310 51594 2358
rect 51522 2264 51535 2310
rect 51581 2264 51594 2310
rect 51522 2216 51594 2264
rect 51522 2170 51535 2216
rect 51581 2170 51594 2216
rect 51522 2122 51594 2170
rect 51522 2076 51535 2122
rect 51581 2076 51594 2122
rect 51522 2028 51594 2076
rect 51522 1982 51535 2028
rect 51581 1982 51594 2028
rect 51522 1934 51594 1982
rect 51522 1888 51535 1934
rect 51581 1888 51594 1934
rect 55658 2498 55730 2546
rect 59794 2592 59866 2640
rect 59794 2546 59807 2592
rect 59853 2546 59866 2592
rect 55658 2452 55671 2498
rect 55717 2452 55730 2498
rect 55658 2404 55730 2452
rect 55658 2358 55671 2404
rect 55717 2358 55730 2404
rect 55658 2310 55730 2358
rect 55658 2264 55671 2310
rect 55717 2264 55730 2310
rect 55658 2216 55730 2264
rect 55658 2170 55671 2216
rect 55717 2170 55730 2216
rect 55658 2122 55730 2170
rect 55658 2076 55671 2122
rect 55717 2076 55730 2122
rect 55658 2028 55730 2076
rect 55658 1982 55671 2028
rect 55717 1982 55730 2028
rect 55658 1934 55730 1982
rect 51522 1840 51594 1888
rect 51522 1794 51535 1840
rect 51581 1794 51594 1840
rect 51522 1746 51594 1794
rect 51522 1700 51535 1746
rect 51581 1700 51594 1746
rect 51522 1652 51594 1700
rect 51522 1606 51535 1652
rect 51581 1606 51594 1652
rect 51522 1558 51594 1606
rect 51522 1512 51535 1558
rect 51581 1512 51594 1558
rect 51522 1464 51594 1512
rect 51522 1418 51535 1464
rect 51581 1418 51594 1464
rect 51522 1370 51594 1418
rect 51522 1324 51535 1370
rect 51581 1324 51594 1370
rect 51522 1276 51594 1324
rect 51522 1230 51535 1276
rect 51581 1230 51594 1276
rect 51522 1182 51594 1230
rect 51522 1136 51535 1182
rect 51581 1136 51594 1182
rect 51522 1088 51594 1136
rect 51522 1042 51535 1088
rect 51581 1042 51594 1088
rect 51522 994 51594 1042
rect 51522 948 51535 994
rect 51581 948 51594 994
rect 51522 900 51594 948
rect 51522 854 51535 900
rect 51581 854 51594 900
rect 51522 806 51594 854
rect 51522 760 51535 806
rect 51581 760 51594 806
rect 51522 712 51594 760
rect 51522 666 51535 712
rect 51581 666 51594 712
rect 51522 618 51594 666
rect 51522 572 51535 618
rect 51581 572 51594 618
rect 51522 524 51594 572
rect 51522 478 51535 524
rect 51581 478 51594 524
rect 51522 430 51594 478
rect 51522 384 51535 430
rect 51581 384 51594 430
rect 51522 336 51594 384
rect 51522 290 51535 336
rect 51581 290 51594 336
rect 51522 242 51594 290
rect 51522 196 51535 242
rect 51581 196 51594 242
rect 51522 148 51594 196
rect 51522 102 51535 148
rect 51581 102 51594 148
rect 51522 54 51594 102
rect 51522 8 51535 54
rect 51581 8 51594 54
rect 51522 -40 51594 8
rect 51522 -86 51535 -40
rect 51581 -86 51594 -40
rect 51522 -134 51594 -86
rect 51522 -180 51535 -134
rect 51581 -180 51594 -134
rect 51522 -228 51594 -180
rect 51522 -274 51535 -228
rect 51581 -274 51594 -228
rect 51522 -322 51594 -274
rect 51522 -368 51535 -322
rect 51581 -368 51594 -322
rect 51522 -416 51594 -368
rect 55658 1888 55671 1934
rect 55717 1888 55730 1934
rect 59794 2498 59866 2546
rect 59794 2452 59807 2498
rect 59853 2452 59866 2498
rect 59794 2404 59866 2452
rect 59794 2358 59807 2404
rect 59853 2358 59866 2404
rect 59794 2310 59866 2358
rect 59794 2264 59807 2310
rect 59853 2264 59866 2310
rect 59794 2216 59866 2264
rect 59794 2170 59807 2216
rect 59853 2170 59866 2216
rect 59794 2122 59866 2170
rect 59794 2076 59807 2122
rect 59853 2076 59866 2122
rect 59794 2028 59866 2076
rect 59794 1982 59807 2028
rect 59853 1982 59866 2028
rect 59794 1934 59866 1982
rect 55658 1840 55730 1888
rect 55658 1794 55671 1840
rect 55717 1794 55730 1840
rect 55658 1746 55730 1794
rect 55658 1700 55671 1746
rect 55717 1700 55730 1746
rect 51522 -462 51535 -416
rect 51581 -462 51594 -416
rect 51522 -510 51594 -462
rect 51522 -556 51535 -510
rect 51581 -556 51594 -510
rect 51522 -604 51594 -556
rect 51522 -650 51535 -604
rect 51581 -650 51594 -604
rect 55658 1652 55730 1700
rect 55658 1606 55671 1652
rect 55717 1606 55730 1652
rect 55658 1558 55730 1606
rect 55658 1512 55671 1558
rect 55717 1512 55730 1558
rect 55658 1464 55730 1512
rect 55658 1418 55671 1464
rect 55717 1418 55730 1464
rect 55658 1370 55730 1418
rect 55658 1324 55671 1370
rect 55717 1324 55730 1370
rect 55658 1276 55730 1324
rect 55658 1230 55671 1276
rect 55717 1230 55730 1276
rect 55658 1182 55730 1230
rect 55658 1136 55671 1182
rect 55717 1136 55730 1182
rect 55658 1088 55730 1136
rect 55658 1042 55671 1088
rect 55717 1042 55730 1088
rect 55658 994 55730 1042
rect 55658 948 55671 994
rect 55717 948 55730 994
rect 55658 900 55730 948
rect 55658 854 55671 900
rect 55717 854 55730 900
rect 55658 806 55730 854
rect 55658 760 55671 806
rect 55717 760 55730 806
rect 55658 712 55730 760
rect 55658 666 55671 712
rect 55717 666 55730 712
rect 55658 618 55730 666
rect 55658 572 55671 618
rect 55717 572 55730 618
rect 55658 524 55730 572
rect 55658 478 55671 524
rect 55717 478 55730 524
rect 55658 430 55730 478
rect 55658 384 55671 430
rect 55717 384 55730 430
rect 55658 336 55730 384
rect 55658 290 55671 336
rect 55717 290 55730 336
rect 55658 242 55730 290
rect 55658 196 55671 242
rect 55717 196 55730 242
rect 55658 148 55730 196
rect 55658 102 55671 148
rect 55717 102 55730 148
rect 55658 54 55730 102
rect 55658 8 55671 54
rect 55717 8 55730 54
rect 55658 -40 55730 8
rect 55658 -86 55671 -40
rect 55717 -86 55730 -40
rect 55658 -134 55730 -86
rect 55658 -180 55671 -134
rect 55717 -180 55730 -134
rect 55658 -228 55730 -180
rect 55658 -274 55671 -228
rect 55717 -274 55730 -228
rect 55658 -322 55730 -274
rect 55658 -368 55671 -322
rect 55717 -368 55730 -322
rect 55658 -416 55730 -368
rect 59794 1888 59807 1934
rect 59853 1888 59866 1934
rect 59794 1840 59866 1888
rect 59794 1794 59807 1840
rect 59853 1794 59866 1840
rect 59794 1746 59866 1794
rect 59794 1700 59807 1746
rect 59853 1700 59866 1746
rect 55658 -462 55671 -416
rect 55717 -462 55730 -416
rect 55658 -510 55730 -462
rect 55658 -556 55671 -510
rect 55717 -556 55730 -510
rect 55658 -604 55730 -556
rect 51522 -698 51594 -650
rect 51522 -744 51535 -698
rect 51581 -744 51594 -698
rect 51522 -792 51594 -744
rect 51522 -838 51535 -792
rect 51581 -838 51594 -792
rect 51522 -886 51594 -838
rect 51522 -932 51535 -886
rect 51581 -932 51594 -886
rect 51522 -980 51594 -932
rect 51522 -1026 51535 -980
rect 51581 -1026 51594 -980
rect 51522 -1074 51594 -1026
rect 51522 -1120 51535 -1074
rect 51581 -1120 51594 -1074
rect 51522 -1168 51594 -1120
rect 51522 -1214 51535 -1168
rect 51581 -1214 51594 -1168
rect 51522 -1262 51594 -1214
rect 51522 -1308 51535 -1262
rect 51581 -1308 51594 -1262
rect 51522 -1356 51594 -1308
rect 51522 -1402 51535 -1356
rect 51581 -1402 51594 -1356
rect 51522 -1450 51594 -1402
rect 51522 -1496 51535 -1450
rect 51581 -1496 51594 -1450
rect 51522 -1544 51594 -1496
rect 51522 -1590 51535 -1544
rect 51581 -1590 51594 -1544
rect 51522 -1638 51594 -1590
rect 51522 -1684 51535 -1638
rect 51581 -1684 51594 -1638
rect 51522 -1719 51594 -1684
rect 55658 -650 55671 -604
rect 55717 -650 55730 -604
rect 59794 1652 59866 1700
rect 59794 1606 59807 1652
rect 59853 1606 59866 1652
rect 59794 1558 59866 1606
rect 59794 1512 59807 1558
rect 59853 1512 59866 1558
rect 59794 1464 59866 1512
rect 59794 1418 59807 1464
rect 59853 1418 59866 1464
rect 59794 1370 59866 1418
rect 59794 1324 59807 1370
rect 59853 1324 59866 1370
rect 59794 1276 59866 1324
rect 59794 1230 59807 1276
rect 59853 1230 59866 1276
rect 59794 1182 59866 1230
rect 59794 1136 59807 1182
rect 59853 1136 59866 1182
rect 59794 1088 59866 1136
rect 59794 1042 59807 1088
rect 59853 1042 59866 1088
rect 59794 994 59866 1042
rect 59794 948 59807 994
rect 59853 948 59866 994
rect 59794 900 59866 948
rect 59794 854 59807 900
rect 59853 854 59866 900
rect 59794 806 59866 854
rect 59794 760 59807 806
rect 59853 760 59866 806
rect 59794 712 59866 760
rect 59794 666 59807 712
rect 59853 666 59866 712
rect 59794 618 59866 666
rect 59794 572 59807 618
rect 59853 572 59866 618
rect 59794 524 59866 572
rect 59794 478 59807 524
rect 59853 478 59866 524
rect 59794 430 59866 478
rect 59794 384 59807 430
rect 59853 384 59866 430
rect 59794 336 59866 384
rect 59794 290 59807 336
rect 59853 290 59866 336
rect 59794 242 59866 290
rect 59794 196 59807 242
rect 59853 196 59866 242
rect 59794 148 59866 196
rect 59794 102 59807 148
rect 59853 102 59866 148
rect 59794 54 59866 102
rect 59794 8 59807 54
rect 59853 8 59866 54
rect 59794 -40 59866 8
rect 59794 -86 59807 -40
rect 59853 -86 59866 -40
rect 59794 -134 59866 -86
rect 59794 -180 59807 -134
rect 59853 -180 59866 -134
rect 59794 -228 59866 -180
rect 59794 -274 59807 -228
rect 59853 -274 59866 -228
rect 59794 -322 59866 -274
rect 59794 -368 59807 -322
rect 59853 -368 59866 -322
rect 59794 -416 59866 -368
rect 59794 -462 59807 -416
rect 59853 -462 59866 -416
rect 59794 -510 59866 -462
rect 59794 -556 59807 -510
rect 59853 -556 59866 -510
rect 59794 -604 59866 -556
rect 55658 -698 55730 -650
rect 55658 -744 55671 -698
rect 55717 -744 55730 -698
rect 55658 -792 55730 -744
rect 55658 -838 55671 -792
rect 55717 -838 55730 -792
rect 55658 -886 55730 -838
rect 55658 -932 55671 -886
rect 55717 -932 55730 -886
rect 55658 -980 55730 -932
rect 55658 -1026 55671 -980
rect 55717 -1026 55730 -980
rect 55658 -1074 55730 -1026
rect 55658 -1120 55671 -1074
rect 55717 -1120 55730 -1074
rect 55658 -1168 55730 -1120
rect 55658 -1214 55671 -1168
rect 55717 -1214 55730 -1168
rect 55658 -1262 55730 -1214
rect 55658 -1308 55671 -1262
rect 55717 -1308 55730 -1262
rect 55658 -1356 55730 -1308
rect 55658 -1402 55671 -1356
rect 55717 -1402 55730 -1356
rect 55658 -1450 55730 -1402
rect 55658 -1496 55671 -1450
rect 55717 -1496 55730 -1450
rect 55658 -1544 55730 -1496
rect 55658 -1590 55671 -1544
rect 55717 -1590 55730 -1544
rect 55658 -1638 55730 -1590
rect 55658 -1684 55671 -1638
rect 55717 -1684 55730 -1638
rect 55658 -1719 55730 -1684
rect 59794 -650 59807 -604
rect 59853 -650 59866 -604
rect 59794 -698 59866 -650
rect 59794 -744 59807 -698
rect 59853 -744 59866 -698
rect 59794 -792 59866 -744
rect 59794 -838 59807 -792
rect 59853 -838 59866 -792
rect 59794 -886 59866 -838
rect 59794 -932 59807 -886
rect 59853 -932 59866 -886
rect 59794 -980 59866 -932
rect 59794 -1026 59807 -980
rect 59853 -1026 59866 -980
rect 59794 -1074 59866 -1026
rect 59794 -1120 59807 -1074
rect 59853 -1120 59866 -1074
rect 59794 -1168 59866 -1120
rect 59794 -1214 59807 -1168
rect 59853 -1214 59866 -1168
rect 59794 -1262 59866 -1214
rect 59794 -1308 59807 -1262
rect 59853 -1308 59866 -1262
rect 59794 -1356 59866 -1308
rect 59794 -1402 59807 -1356
rect 59853 -1402 59866 -1356
rect 59794 -1450 59866 -1402
rect 59794 -1496 59807 -1450
rect 59853 -1496 59866 -1450
rect 59794 -1544 59866 -1496
rect 59794 -1590 59807 -1544
rect 59853 -1590 59866 -1544
rect 59794 -1638 59866 -1590
rect 59794 -1684 59807 -1638
rect 59853 -1684 59866 -1638
rect 59794 -1719 59866 -1684
rect 51522 -1732 59866 -1719
rect 51522 -1778 51535 -1732
rect 51581 -1778 51629 -1732
rect 51675 -1778 51723 -1732
rect 51769 -1778 51817 -1732
rect 51863 -1778 51911 -1732
rect 51957 -1778 52005 -1732
rect 52051 -1778 52099 -1732
rect 52145 -1778 52193 -1732
rect 52239 -1778 52287 -1732
rect 52333 -1778 52381 -1732
rect 52427 -1778 52475 -1732
rect 52521 -1778 52569 -1732
rect 52615 -1778 52663 -1732
rect 52709 -1778 52757 -1732
rect 52803 -1778 52851 -1732
rect 52897 -1778 52945 -1732
rect 52991 -1778 53039 -1732
rect 53085 -1778 53133 -1732
rect 53179 -1778 53227 -1732
rect 53273 -1778 53321 -1732
rect 53367 -1778 53415 -1732
rect 53461 -1778 53509 -1732
rect 53555 -1778 53603 -1732
rect 53649 -1778 53697 -1732
rect 53743 -1778 53791 -1732
rect 53837 -1778 53885 -1732
rect 53931 -1778 53979 -1732
rect 54025 -1778 54073 -1732
rect 54119 -1778 54167 -1732
rect 54213 -1778 54261 -1732
rect 54307 -1778 54355 -1732
rect 54401 -1778 54449 -1732
rect 54495 -1778 54543 -1732
rect 54589 -1778 54637 -1732
rect 54683 -1778 54731 -1732
rect 54777 -1778 54825 -1732
rect 54871 -1778 54919 -1732
rect 54965 -1778 55013 -1732
rect 55059 -1778 55107 -1732
rect 55153 -1778 55201 -1732
rect 55247 -1778 55295 -1732
rect 55341 -1778 55389 -1732
rect 55435 -1778 55483 -1732
rect 55529 -1778 55577 -1732
rect 55623 -1778 55671 -1732
rect 55717 -1778 55765 -1732
rect 55811 -1778 55859 -1732
rect 55905 -1778 55953 -1732
rect 55999 -1778 56047 -1732
rect 56093 -1778 56141 -1732
rect 56187 -1778 56235 -1732
rect 56281 -1778 56329 -1732
rect 56375 -1778 56423 -1732
rect 56469 -1778 56517 -1732
rect 56563 -1778 56611 -1732
rect 56657 -1778 56705 -1732
rect 56751 -1778 56799 -1732
rect 56845 -1778 56893 -1732
rect 56939 -1778 56987 -1732
rect 57033 -1778 57081 -1732
rect 57127 -1778 57175 -1732
rect 57221 -1778 57269 -1732
rect 57315 -1778 57363 -1732
rect 57409 -1778 57457 -1732
rect 57503 -1778 57551 -1732
rect 57597 -1778 57645 -1732
rect 57691 -1778 57739 -1732
rect 57785 -1778 57833 -1732
rect 57879 -1778 57927 -1732
rect 57973 -1778 58021 -1732
rect 58067 -1778 58115 -1732
rect 58161 -1778 58209 -1732
rect 58255 -1778 58303 -1732
rect 58349 -1778 58397 -1732
rect 58443 -1778 58491 -1732
rect 58537 -1778 58585 -1732
rect 58631 -1778 58679 -1732
rect 58725 -1778 58773 -1732
rect 58819 -1778 58867 -1732
rect 58913 -1778 58961 -1732
rect 59007 -1778 59055 -1732
rect 59101 -1778 59149 -1732
rect 59195 -1778 59243 -1732
rect 59289 -1778 59337 -1732
rect 59383 -1778 59431 -1732
rect 59477 -1778 59525 -1732
rect 59571 -1778 59619 -1732
rect 59665 -1778 59713 -1732
rect 59759 -1778 59807 -1732
rect 59853 -1778 59866 -1732
rect 51522 -1791 59866 -1778
rect 61218 3062 65426 3075
rect 61218 3016 61231 3062
rect 61277 3016 61325 3062
rect 61371 3016 61419 3062
rect 61465 3016 61513 3062
rect 61559 3016 61607 3062
rect 61653 3016 61701 3062
rect 61747 3016 61795 3062
rect 61841 3016 61889 3062
rect 61935 3016 61983 3062
rect 62029 3016 62077 3062
rect 62123 3016 62171 3062
rect 62217 3016 62265 3062
rect 62311 3016 62359 3062
rect 62405 3016 62453 3062
rect 62499 3016 62547 3062
rect 62593 3016 62641 3062
rect 62687 3016 62735 3062
rect 62781 3016 62829 3062
rect 62875 3016 62923 3062
rect 62969 3016 63017 3062
rect 63063 3016 63111 3062
rect 63157 3016 63205 3062
rect 63251 3016 63299 3062
rect 63345 3016 63393 3062
rect 63439 3016 63487 3062
rect 63533 3016 63581 3062
rect 63627 3016 63675 3062
rect 63721 3016 63769 3062
rect 63815 3016 63863 3062
rect 63909 3016 63957 3062
rect 64003 3016 64051 3062
rect 64097 3016 64145 3062
rect 64191 3016 64239 3062
rect 64285 3016 64333 3062
rect 64379 3016 64427 3062
rect 64473 3016 64521 3062
rect 64567 3016 64615 3062
rect 64661 3016 64709 3062
rect 64755 3016 64803 3062
rect 64849 3016 64897 3062
rect 64943 3016 64991 3062
rect 65037 3016 65085 3062
rect 65131 3016 65179 3062
rect 65225 3016 65273 3062
rect 65319 3016 65367 3062
rect 65413 3016 65426 3062
rect 61218 3003 65426 3016
rect 61218 2968 61290 3003
rect 61218 2922 61231 2968
rect 61277 2922 61290 2968
rect 61218 2874 61290 2922
rect 61218 2828 61231 2874
rect 61277 2828 61290 2874
rect 61218 2780 61290 2828
rect 61218 2734 61231 2780
rect 61277 2734 61290 2780
rect 61218 2686 61290 2734
rect 61218 2640 61231 2686
rect 61277 2640 61290 2686
rect 65354 2968 65426 3003
rect 65354 2922 65367 2968
rect 65413 2922 65426 2968
rect 65354 2874 65426 2922
rect 65354 2828 65367 2874
rect 65413 2828 65426 2874
rect 65354 2780 65426 2828
rect 65354 2734 65367 2780
rect 65413 2734 65426 2780
rect 65354 2686 65426 2734
rect 61218 2592 61290 2640
rect 65354 2640 65367 2686
rect 65413 2640 65426 2686
rect 61218 2546 61231 2592
rect 61277 2546 61290 2592
rect 61218 2498 61290 2546
rect 65354 2592 65426 2640
rect 65354 2546 65367 2592
rect 65413 2546 65426 2592
rect 61218 2452 61231 2498
rect 61277 2452 61290 2498
rect 61218 2404 61290 2452
rect 61218 2358 61231 2404
rect 61277 2358 61290 2404
rect 61218 2310 61290 2358
rect 61218 2264 61231 2310
rect 61277 2264 61290 2310
rect 61218 2216 61290 2264
rect 61218 2170 61231 2216
rect 61277 2170 61290 2216
rect 61218 2122 61290 2170
rect 61218 2076 61231 2122
rect 61277 2076 61290 2122
rect 61218 2028 61290 2076
rect 61218 1982 61231 2028
rect 61277 1982 61290 2028
rect 61218 1934 61290 1982
rect 61218 1888 61231 1934
rect 61277 1888 61290 1934
rect 65354 2498 65426 2546
rect 65354 2452 65367 2498
rect 65413 2452 65426 2498
rect 65354 2404 65426 2452
rect 65354 2358 65367 2404
rect 65413 2358 65426 2404
rect 65354 2310 65426 2358
rect 65354 2264 65367 2310
rect 65413 2264 65426 2310
rect 65354 2216 65426 2264
rect 65354 2170 65367 2216
rect 65413 2170 65426 2216
rect 65354 2122 65426 2170
rect 65354 2076 65367 2122
rect 65413 2076 65426 2122
rect 65354 2028 65426 2076
rect 65354 1982 65367 2028
rect 65413 1982 65426 2028
rect 65354 1934 65426 1982
rect 61218 1840 61290 1888
rect 61218 1794 61231 1840
rect 61277 1794 61290 1840
rect 61218 1746 61290 1794
rect 61218 1700 61231 1746
rect 61277 1700 61290 1746
rect 61218 1652 61290 1700
rect 61218 1606 61231 1652
rect 61277 1606 61290 1652
rect 61218 1558 61290 1606
rect 61218 1512 61231 1558
rect 61277 1512 61290 1558
rect 61218 1464 61290 1512
rect 61218 1418 61231 1464
rect 61277 1418 61290 1464
rect 61218 1370 61290 1418
rect 61218 1324 61231 1370
rect 61277 1324 61290 1370
rect 61218 1276 61290 1324
rect 61218 1230 61231 1276
rect 61277 1230 61290 1276
rect 61218 1182 61290 1230
rect 61218 1136 61231 1182
rect 61277 1136 61290 1182
rect 61218 1088 61290 1136
rect 61218 1042 61231 1088
rect 61277 1042 61290 1088
rect 61218 994 61290 1042
rect 61218 948 61231 994
rect 61277 948 61290 994
rect 61218 900 61290 948
rect 61218 854 61231 900
rect 61277 854 61290 900
rect 61218 806 61290 854
rect 61218 760 61231 806
rect 61277 760 61290 806
rect 61218 712 61290 760
rect 61218 666 61231 712
rect 61277 666 61290 712
rect 61218 618 61290 666
rect 61218 572 61231 618
rect 61277 572 61290 618
rect 61218 524 61290 572
rect 61218 478 61231 524
rect 61277 478 61290 524
rect 61218 430 61290 478
rect 61218 384 61231 430
rect 61277 384 61290 430
rect 61218 336 61290 384
rect 61218 290 61231 336
rect 61277 290 61290 336
rect 61218 242 61290 290
rect 61218 196 61231 242
rect 61277 196 61290 242
rect 61218 148 61290 196
rect 61218 102 61231 148
rect 61277 102 61290 148
rect 61218 54 61290 102
rect 61218 8 61231 54
rect 61277 8 61290 54
rect 61218 -40 61290 8
rect 61218 -86 61231 -40
rect 61277 -86 61290 -40
rect 61218 -134 61290 -86
rect 61218 -180 61231 -134
rect 61277 -180 61290 -134
rect 61218 -228 61290 -180
rect 61218 -274 61231 -228
rect 61277 -274 61290 -228
rect 61218 -322 61290 -274
rect 61218 -368 61231 -322
rect 61277 -368 61290 -322
rect 61218 -416 61290 -368
rect 65354 1888 65367 1934
rect 65413 1888 65426 1934
rect 65354 1840 65426 1888
rect 65354 1794 65367 1840
rect 65413 1794 65426 1840
rect 65354 1746 65426 1794
rect 65354 1700 65367 1746
rect 65413 1700 65426 1746
rect 61218 -462 61231 -416
rect 61277 -462 61290 -416
rect 61218 -510 61290 -462
rect 61218 -556 61231 -510
rect 61277 -556 61290 -510
rect 61218 -604 61290 -556
rect 61218 -650 61231 -604
rect 61277 -650 61290 -604
rect 65354 1652 65426 1700
rect 65354 1606 65367 1652
rect 65413 1606 65426 1652
rect 65354 1558 65426 1606
rect 65354 1512 65367 1558
rect 65413 1512 65426 1558
rect 65354 1464 65426 1512
rect 65354 1418 65367 1464
rect 65413 1418 65426 1464
rect 65354 1370 65426 1418
rect 65354 1324 65367 1370
rect 65413 1324 65426 1370
rect 65354 1276 65426 1324
rect 65354 1230 65367 1276
rect 65413 1230 65426 1276
rect 65354 1182 65426 1230
rect 65354 1136 65367 1182
rect 65413 1136 65426 1182
rect 65354 1088 65426 1136
rect 65354 1042 65367 1088
rect 65413 1042 65426 1088
rect 65354 994 65426 1042
rect 65354 948 65367 994
rect 65413 948 65426 994
rect 65354 900 65426 948
rect 65354 854 65367 900
rect 65413 854 65426 900
rect 65354 806 65426 854
rect 65354 760 65367 806
rect 65413 760 65426 806
rect 65354 712 65426 760
rect 65354 666 65367 712
rect 65413 666 65426 712
rect 65354 618 65426 666
rect 65354 572 65367 618
rect 65413 572 65426 618
rect 65354 524 65426 572
rect 65354 478 65367 524
rect 65413 478 65426 524
rect 65354 430 65426 478
rect 65354 384 65367 430
rect 65413 384 65426 430
rect 65354 336 65426 384
rect 65354 290 65367 336
rect 65413 290 65426 336
rect 65354 242 65426 290
rect 65354 196 65367 242
rect 65413 196 65426 242
rect 65354 148 65426 196
rect 65354 102 65367 148
rect 65413 102 65426 148
rect 65354 54 65426 102
rect 65354 8 65367 54
rect 65413 8 65426 54
rect 65354 -40 65426 8
rect 65354 -86 65367 -40
rect 65413 -86 65426 -40
rect 65354 -134 65426 -86
rect 65354 -180 65367 -134
rect 65413 -180 65426 -134
rect 65354 -228 65426 -180
rect 65354 -274 65367 -228
rect 65413 -274 65426 -228
rect 65354 -322 65426 -274
rect 65354 -368 65367 -322
rect 65413 -368 65426 -322
rect 65354 -416 65426 -368
rect 65354 -462 65367 -416
rect 65413 -462 65426 -416
rect 65354 -510 65426 -462
rect 65354 -556 65367 -510
rect 65413 -556 65426 -510
rect 65354 -604 65426 -556
rect 61218 -698 61290 -650
rect 61218 -744 61231 -698
rect 61277 -744 61290 -698
rect 61218 -792 61290 -744
rect 61218 -838 61231 -792
rect 61277 -838 61290 -792
rect 61218 -886 61290 -838
rect 61218 -932 61231 -886
rect 61277 -932 61290 -886
rect 61218 -980 61290 -932
rect 61218 -1026 61231 -980
rect 61277 -1026 61290 -980
rect 61218 -1074 61290 -1026
rect 61218 -1120 61231 -1074
rect 61277 -1120 61290 -1074
rect 61218 -1168 61290 -1120
rect 61218 -1214 61231 -1168
rect 61277 -1214 61290 -1168
rect 61218 -1262 61290 -1214
rect 61218 -1308 61231 -1262
rect 61277 -1308 61290 -1262
rect 61218 -1356 61290 -1308
rect 61218 -1402 61231 -1356
rect 61277 -1402 61290 -1356
rect 61218 -1450 61290 -1402
rect 61218 -1496 61231 -1450
rect 61277 -1496 61290 -1450
rect 61218 -1544 61290 -1496
rect 61218 -1590 61231 -1544
rect 61277 -1590 61290 -1544
rect 61218 -1638 61290 -1590
rect 61218 -1684 61231 -1638
rect 61277 -1684 61290 -1638
rect 61218 -1719 61290 -1684
rect 65354 -650 65367 -604
rect 65413 -650 65426 -604
rect 65354 -698 65426 -650
rect 65354 -744 65367 -698
rect 65413 -744 65426 -698
rect 65354 -792 65426 -744
rect 65354 -838 65367 -792
rect 65413 -838 65426 -792
rect 65354 -886 65426 -838
rect 65354 -932 65367 -886
rect 65413 -932 65426 -886
rect 65354 -980 65426 -932
rect 65354 -1026 65367 -980
rect 65413 -1026 65426 -980
rect 65354 -1074 65426 -1026
rect 65354 -1120 65367 -1074
rect 65413 -1120 65426 -1074
rect 65354 -1168 65426 -1120
rect 65354 -1214 65367 -1168
rect 65413 -1214 65426 -1168
rect 65354 -1262 65426 -1214
rect 65354 -1308 65367 -1262
rect 65413 -1308 65426 -1262
rect 65354 -1356 65426 -1308
rect 65354 -1402 65367 -1356
rect 65413 -1402 65426 -1356
rect 65354 -1450 65426 -1402
rect 65354 -1496 65367 -1450
rect 65413 -1496 65426 -1450
rect 65354 -1544 65426 -1496
rect 65354 -1590 65367 -1544
rect 65413 -1590 65426 -1544
rect 65354 -1638 65426 -1590
rect 65354 -1684 65367 -1638
rect 65413 -1684 65426 -1638
rect 65354 -1719 65426 -1684
rect 61218 -1732 65426 -1719
rect 61218 -1778 61231 -1732
rect 61277 -1778 61325 -1732
rect 61371 -1778 61419 -1732
rect 61465 -1778 61513 -1732
rect 61559 -1778 61607 -1732
rect 61653 -1778 61701 -1732
rect 61747 -1778 61795 -1732
rect 61841 -1778 61889 -1732
rect 61935 -1778 61983 -1732
rect 62029 -1778 62077 -1732
rect 62123 -1778 62171 -1732
rect 62217 -1778 62265 -1732
rect 62311 -1778 62359 -1732
rect 62405 -1778 62453 -1732
rect 62499 -1778 62547 -1732
rect 62593 -1778 62641 -1732
rect 62687 -1778 62735 -1732
rect 62781 -1778 62829 -1732
rect 62875 -1778 62923 -1732
rect 62969 -1778 63017 -1732
rect 63063 -1778 63111 -1732
rect 63157 -1778 63205 -1732
rect 63251 -1778 63299 -1732
rect 63345 -1778 63393 -1732
rect 63439 -1778 63487 -1732
rect 63533 -1778 63581 -1732
rect 63627 -1778 63675 -1732
rect 63721 -1778 63769 -1732
rect 63815 -1778 63863 -1732
rect 63909 -1778 63957 -1732
rect 64003 -1778 64051 -1732
rect 64097 -1778 64145 -1732
rect 64191 -1778 64239 -1732
rect 64285 -1778 64333 -1732
rect 64379 -1778 64427 -1732
rect 64473 -1778 64521 -1732
rect 64567 -1778 64615 -1732
rect 64661 -1778 64709 -1732
rect 64755 -1778 64803 -1732
rect 64849 -1778 64897 -1732
rect 64943 -1778 64991 -1732
rect 65037 -1778 65085 -1732
rect 65131 -1778 65179 -1732
rect 65225 -1778 65273 -1732
rect 65319 -1778 65367 -1732
rect 65413 -1778 65426 -1732
rect 61218 -1791 65426 -1778
rect 11401 -1892 16549 -1879
rect 430 -4365 4544 -4352
rect 430 -4411 443 -4365
rect 489 -4411 537 -4365
rect 583 -4411 631 -4365
rect 677 -4411 725 -4365
rect 771 -4411 819 -4365
rect 865 -4411 913 -4365
rect 959 -4411 1007 -4365
rect 1053 -4411 1101 -4365
rect 1147 -4411 1195 -4365
rect 1241 -4411 1289 -4365
rect 1335 -4411 1383 -4365
rect 1429 -4411 1477 -4365
rect 1523 -4411 1571 -4365
rect 1617 -4411 1665 -4365
rect 1711 -4411 1759 -4365
rect 1805 -4411 1853 -4365
rect 1899 -4411 1947 -4365
rect 1993 -4411 2041 -4365
rect 2087 -4411 2135 -4365
rect 2181 -4411 2229 -4365
rect 2275 -4411 2323 -4365
rect 2369 -4411 2417 -4365
rect 2463 -4411 2511 -4365
rect 2557 -4411 2605 -4365
rect 2651 -4411 2699 -4365
rect 2745 -4411 2793 -4365
rect 2839 -4411 2887 -4365
rect 2933 -4411 2981 -4365
rect 3027 -4411 3075 -4365
rect 3121 -4411 3169 -4365
rect 3215 -4411 3263 -4365
rect 3309 -4411 3357 -4365
rect 3403 -4411 3451 -4365
rect 3497 -4411 3545 -4365
rect 3591 -4411 3639 -4365
rect 3685 -4411 3733 -4365
rect 3779 -4411 3827 -4365
rect 3873 -4411 3921 -4365
rect 3967 -4411 4015 -4365
rect 4061 -4411 4109 -4365
rect 4155 -4411 4203 -4365
rect 4249 -4411 4297 -4365
rect 4343 -4411 4391 -4365
rect 4437 -4411 4485 -4365
rect 4531 -4411 4544 -4365
rect 430 -4424 4544 -4411
rect 430 -4459 502 -4424
rect 430 -4505 443 -4459
rect 489 -4505 502 -4459
rect 430 -4553 502 -4505
rect 430 -4599 443 -4553
rect 489 -4599 502 -4553
rect 4472 -4459 4544 -4424
rect 4472 -4505 4485 -4459
rect 4531 -4505 4544 -4459
rect 4472 -4553 4544 -4505
rect 430 -4647 502 -4599
rect 430 -4693 443 -4647
rect 489 -4693 502 -4647
rect 430 -4741 502 -4693
rect 4472 -4599 4485 -4553
rect 4531 -4599 4544 -4553
rect 4472 -4647 4544 -4599
rect 4472 -4693 4485 -4647
rect 4531 -4693 4544 -4647
rect 430 -4787 443 -4741
rect 489 -4787 502 -4741
rect 430 -4835 502 -4787
rect 430 -4881 443 -4835
rect 489 -4881 502 -4835
rect 430 -4929 502 -4881
rect 430 -4975 443 -4929
rect 489 -4975 502 -4929
rect 430 -5023 502 -4975
rect 430 -5069 443 -5023
rect 489 -5069 502 -5023
rect 430 -5117 502 -5069
rect 430 -5163 443 -5117
rect 489 -5163 502 -5117
rect 430 -5211 502 -5163
rect 430 -5257 443 -5211
rect 489 -5257 502 -5211
rect 430 -5305 502 -5257
rect 430 -5351 443 -5305
rect 489 -5351 502 -5305
rect 430 -5399 502 -5351
rect 430 -5445 443 -5399
rect 489 -5445 502 -5399
rect 430 -5493 502 -5445
rect 430 -5539 443 -5493
rect 489 -5539 502 -5493
rect 4472 -4741 4544 -4693
rect 4472 -4787 4485 -4741
rect 4531 -4787 4544 -4741
rect 4472 -4835 4544 -4787
rect 4472 -4881 4485 -4835
rect 4531 -4881 4544 -4835
rect 4472 -4929 4544 -4881
rect 4472 -4975 4485 -4929
rect 4531 -4975 4544 -4929
rect 4472 -5023 4544 -4975
rect 4472 -5069 4485 -5023
rect 4531 -5069 4544 -5023
rect 4472 -5117 4544 -5069
rect 4472 -5163 4485 -5117
rect 4531 -5163 4544 -5117
rect 4472 -5211 4544 -5163
rect 4472 -5257 4485 -5211
rect 4531 -5257 4544 -5211
rect 4472 -5305 4544 -5257
rect 4472 -5351 4485 -5305
rect 4531 -5351 4544 -5305
rect 4472 -5399 4544 -5351
rect 4472 -5445 4485 -5399
rect 4531 -5445 4544 -5399
rect 4472 -5493 4544 -5445
rect 430 -5587 502 -5539
rect 430 -5633 443 -5587
rect 489 -5633 502 -5587
rect 430 -5681 502 -5633
rect 430 -5727 443 -5681
rect 489 -5727 502 -5681
rect 430 -5775 502 -5727
rect 430 -5821 443 -5775
rect 489 -5821 502 -5775
rect 430 -5869 502 -5821
rect 430 -5915 443 -5869
rect 489 -5915 502 -5869
rect 430 -5963 502 -5915
rect 430 -6009 443 -5963
rect 489 -6009 502 -5963
rect 4472 -5539 4485 -5493
rect 4531 -5539 4544 -5493
rect 4472 -5587 4544 -5539
rect 4472 -5633 4485 -5587
rect 4531 -5633 4544 -5587
rect 4472 -5681 4544 -5633
rect 4472 -5727 4485 -5681
rect 4531 -5727 4544 -5681
rect 4472 -5775 4544 -5727
rect 4472 -5821 4485 -5775
rect 4531 -5821 4544 -5775
rect 4472 -5869 4544 -5821
rect 4472 -5915 4485 -5869
rect 4531 -5915 4544 -5869
rect 4472 -5963 4544 -5915
rect 430 -6057 502 -6009
rect 430 -6103 443 -6057
rect 489 -6103 502 -6057
rect 430 -6151 502 -6103
rect 430 -6197 443 -6151
rect 489 -6197 502 -6151
rect 430 -6245 502 -6197
rect 430 -6291 443 -6245
rect 489 -6291 502 -6245
rect 430 -6339 502 -6291
rect 430 -6385 443 -6339
rect 489 -6385 502 -6339
rect 430 -6433 502 -6385
rect 430 -6479 443 -6433
rect 489 -6479 502 -6433
rect 430 -6527 502 -6479
rect 430 -6573 443 -6527
rect 489 -6573 502 -6527
rect 430 -6621 502 -6573
rect 430 -6667 443 -6621
rect 489 -6667 502 -6621
rect 430 -6715 502 -6667
rect 430 -6761 443 -6715
rect 489 -6761 502 -6715
rect 430 -6809 502 -6761
rect 4472 -6009 4485 -5963
rect 4531 -6009 4544 -5963
rect 4472 -6057 4544 -6009
rect 4472 -6103 4485 -6057
rect 4531 -6103 4544 -6057
rect 4472 -6151 4544 -6103
rect 4472 -6197 4485 -6151
rect 4531 -6197 4544 -6151
rect 4472 -6245 4544 -6197
rect 4472 -6291 4485 -6245
rect 4531 -6291 4544 -6245
rect 4472 -6339 4544 -6291
rect 17707 -3456 31315 -3443
rect 17707 -3502 17720 -3456
rect 17766 -3502 17814 -3456
rect 17860 -3502 17908 -3456
rect 17954 -3502 18002 -3456
rect 18048 -3502 18096 -3456
rect 18142 -3502 18190 -3456
rect 18236 -3502 18284 -3456
rect 18330 -3502 18378 -3456
rect 18424 -3502 18472 -3456
rect 18518 -3502 18566 -3456
rect 18612 -3502 18660 -3456
rect 18706 -3502 18754 -3456
rect 18800 -3502 18848 -3456
rect 18894 -3502 18942 -3456
rect 18988 -3502 19036 -3456
rect 19082 -3502 19130 -3456
rect 19176 -3502 19224 -3456
rect 19270 -3502 19318 -3456
rect 19364 -3502 19412 -3456
rect 19458 -3502 19506 -3456
rect 19552 -3502 19600 -3456
rect 19646 -3502 19694 -3456
rect 19740 -3502 19788 -3456
rect 19834 -3502 19882 -3456
rect 19928 -3502 19976 -3456
rect 20022 -3502 20070 -3456
rect 20116 -3502 20164 -3456
rect 20210 -3502 20258 -3456
rect 20304 -3502 20352 -3456
rect 20398 -3502 20446 -3456
rect 20492 -3502 20540 -3456
rect 20586 -3502 20634 -3456
rect 20680 -3502 20728 -3456
rect 20774 -3502 20822 -3456
rect 20868 -3502 20916 -3456
rect 20962 -3502 21010 -3456
rect 21056 -3502 21104 -3456
rect 21150 -3502 21198 -3456
rect 21244 -3502 21292 -3456
rect 21338 -3502 21386 -3456
rect 21432 -3502 21480 -3456
rect 21526 -3502 21574 -3456
rect 21620 -3502 21668 -3456
rect 21714 -3502 21762 -3456
rect 21808 -3502 21856 -3456
rect 21902 -3502 21950 -3456
rect 21996 -3502 22044 -3456
rect 22090 -3502 22138 -3456
rect 22184 -3502 22232 -3456
rect 22278 -3502 22326 -3456
rect 22372 -3502 22420 -3456
rect 22466 -3502 22514 -3456
rect 22560 -3502 22608 -3456
rect 22654 -3502 22702 -3456
rect 22748 -3502 22796 -3456
rect 22842 -3502 22890 -3456
rect 22936 -3502 22984 -3456
rect 23030 -3502 23078 -3456
rect 23124 -3502 23172 -3456
rect 23218 -3502 23266 -3456
rect 23312 -3502 23360 -3456
rect 23406 -3502 23454 -3456
rect 23500 -3502 23548 -3456
rect 23594 -3502 23642 -3456
rect 23688 -3502 23736 -3456
rect 23782 -3502 23830 -3456
rect 23876 -3502 23924 -3456
rect 23970 -3502 24018 -3456
rect 24064 -3502 24112 -3456
rect 24158 -3502 24206 -3456
rect 24252 -3502 24300 -3456
rect 24346 -3502 24394 -3456
rect 24440 -3502 24488 -3456
rect 24534 -3502 24582 -3456
rect 24628 -3502 24676 -3456
rect 24722 -3502 24770 -3456
rect 24816 -3502 24864 -3456
rect 24910 -3502 24958 -3456
rect 25004 -3502 25052 -3456
rect 25098 -3502 25146 -3456
rect 25192 -3502 25240 -3456
rect 25286 -3502 25334 -3456
rect 25380 -3502 25428 -3456
rect 25474 -3502 25522 -3456
rect 25568 -3502 25616 -3456
rect 25662 -3502 25710 -3456
rect 25756 -3502 25804 -3456
rect 25850 -3502 25898 -3456
rect 25944 -3502 25992 -3456
rect 26038 -3502 26086 -3456
rect 26132 -3502 26180 -3456
rect 26226 -3502 26274 -3456
rect 26320 -3502 26368 -3456
rect 26414 -3502 26462 -3456
rect 26508 -3502 26556 -3456
rect 26602 -3502 26650 -3456
rect 26696 -3502 26744 -3456
rect 26790 -3502 26838 -3456
rect 26884 -3502 26932 -3456
rect 26978 -3502 27026 -3456
rect 27072 -3502 27120 -3456
rect 27166 -3502 27214 -3456
rect 27260 -3502 27308 -3456
rect 27354 -3502 27402 -3456
rect 27448 -3502 27496 -3456
rect 27542 -3502 27590 -3456
rect 27636 -3502 27684 -3456
rect 27730 -3502 27778 -3456
rect 27824 -3502 27872 -3456
rect 27918 -3502 27966 -3456
rect 28012 -3502 28060 -3456
rect 28106 -3502 28154 -3456
rect 28200 -3502 28248 -3456
rect 28294 -3502 28342 -3456
rect 28388 -3502 28436 -3456
rect 28482 -3502 28530 -3456
rect 28576 -3502 28624 -3456
rect 28670 -3502 28718 -3456
rect 28764 -3502 28812 -3456
rect 28858 -3502 28906 -3456
rect 28952 -3502 29000 -3456
rect 29046 -3502 29094 -3456
rect 29140 -3502 29188 -3456
rect 29234 -3502 29282 -3456
rect 29328 -3502 29376 -3456
rect 29422 -3502 29470 -3456
rect 29516 -3502 29564 -3456
rect 29610 -3502 29658 -3456
rect 29704 -3502 29752 -3456
rect 29798 -3502 29846 -3456
rect 29892 -3502 29940 -3456
rect 29986 -3502 30034 -3456
rect 30080 -3502 30128 -3456
rect 30174 -3502 30222 -3456
rect 30268 -3502 30316 -3456
rect 30362 -3502 30410 -3456
rect 30456 -3502 30504 -3456
rect 30550 -3502 30598 -3456
rect 30644 -3502 30692 -3456
rect 30738 -3502 30786 -3456
rect 30832 -3502 30880 -3456
rect 30926 -3502 30974 -3456
rect 31020 -3502 31068 -3456
rect 31114 -3502 31162 -3456
rect 31208 -3502 31256 -3456
rect 31302 -3502 31315 -3456
rect 17707 -3515 31315 -3502
rect 17707 -3550 17779 -3515
rect 17707 -3596 17720 -3550
rect 17766 -3596 17779 -3550
rect 17707 -3644 17779 -3596
rect 17707 -3690 17720 -3644
rect 17766 -3690 17779 -3644
rect 17707 -3738 17779 -3690
rect 17707 -3784 17720 -3738
rect 17766 -3784 17779 -3738
rect 17707 -3832 17779 -3784
rect 17707 -3878 17720 -3832
rect 17766 -3878 17779 -3832
rect 17707 -3926 17779 -3878
rect 17707 -3972 17720 -3926
rect 17766 -3972 17779 -3926
rect 17707 -4020 17779 -3972
rect 17707 -4066 17720 -4020
rect 17766 -4066 17779 -4020
rect 17707 -4114 17779 -4066
rect 17707 -4160 17720 -4114
rect 17766 -4160 17779 -4114
rect 17707 -4208 17779 -4160
rect 17707 -4254 17720 -4208
rect 17766 -4254 17779 -4208
rect 22501 -3550 22573 -3515
rect 22501 -3596 22514 -3550
rect 22560 -3596 22573 -3550
rect 22501 -3644 22573 -3596
rect 22501 -3690 22514 -3644
rect 22560 -3690 22573 -3644
rect 22501 -3738 22573 -3690
rect 22501 -3784 22514 -3738
rect 22560 -3784 22573 -3738
rect 22501 -3832 22573 -3784
rect 22501 -3878 22514 -3832
rect 22560 -3878 22573 -3832
rect 22501 -3926 22573 -3878
rect 22501 -3972 22514 -3926
rect 22560 -3972 22573 -3926
rect 22501 -4020 22573 -3972
rect 22501 -4066 22514 -4020
rect 22560 -4066 22573 -4020
rect 22501 -4114 22573 -4066
rect 22501 -4160 22514 -4114
rect 22560 -4160 22573 -4114
rect 22501 -4208 22573 -4160
rect 17707 -4302 17779 -4254
rect 17707 -4348 17720 -4302
rect 17766 -4348 17779 -4302
rect 17707 -4396 17779 -4348
rect 22501 -4254 22514 -4208
rect 22560 -4254 22573 -4208
rect 22501 -4302 22573 -4254
rect 22501 -4348 22514 -4302
rect 22560 -4348 22573 -4302
rect 17707 -4442 17720 -4396
rect 17766 -4442 17779 -4396
rect 17707 -4490 17779 -4442
rect 17707 -4536 17720 -4490
rect 17766 -4536 17779 -4490
rect 17707 -4584 17779 -4536
rect 17707 -4630 17720 -4584
rect 17766 -4630 17779 -4584
rect 4472 -6385 4485 -6339
rect 4531 -6385 4544 -6339
rect 4472 -6433 4544 -6385
rect 4472 -6479 4485 -6433
rect 4531 -6479 4544 -6433
rect 4472 -6527 4544 -6479
rect 4472 -6573 4485 -6527
rect 4531 -6573 4544 -6527
rect 4472 -6621 4544 -6573
rect 4472 -6667 4485 -6621
rect 4531 -6667 4544 -6621
rect 4472 -6715 4544 -6667
rect 4472 -6761 4485 -6715
rect 4531 -6761 4544 -6715
rect 430 -6855 443 -6809
rect 489 -6855 502 -6809
rect 430 -6903 502 -6855
rect 430 -6949 443 -6903
rect 489 -6949 502 -6903
rect 430 -6997 502 -6949
rect 430 -7043 443 -6997
rect 489 -7043 502 -6997
rect 430 -7091 502 -7043
rect 430 -7137 443 -7091
rect 489 -7137 502 -7091
rect 430 -7185 502 -7137
rect 430 -7231 443 -7185
rect 489 -7231 502 -7185
rect 430 -7279 502 -7231
rect 4472 -6809 4544 -6761
rect 4472 -6855 4485 -6809
rect 4531 -6855 4544 -6809
rect 4472 -6903 4544 -6855
rect 4472 -6949 4485 -6903
rect 4531 -6949 4544 -6903
rect 4472 -6997 4544 -6949
rect 4472 -7043 4485 -6997
rect 4531 -7043 4544 -6997
rect 4472 -7091 4544 -7043
rect 4472 -7137 4485 -7091
rect 4531 -7137 4544 -7091
rect 4472 -7185 4544 -7137
rect 4472 -7231 4485 -7185
rect 4531 -7231 4544 -7185
rect 430 -7325 443 -7279
rect 489 -7325 502 -7279
rect 430 -7373 502 -7325
rect 430 -7419 443 -7373
rect 489 -7419 502 -7373
rect 4472 -7279 4544 -7231
rect 4472 -7325 4485 -7279
rect 4531 -7325 4544 -7279
rect 4472 -7373 4544 -7325
rect 430 -7467 502 -7419
rect 4472 -7419 4485 -7373
rect 4531 -7419 4544 -7373
rect 430 -7513 443 -7467
rect 489 -7513 502 -7467
rect 430 -7561 502 -7513
rect 430 -7607 443 -7561
rect 489 -7607 502 -7561
rect 430 -7642 502 -7607
rect 4472 -7467 4544 -7419
rect 4472 -7513 4485 -7467
rect 4531 -7513 4544 -7467
rect 4472 -7561 4544 -7513
rect 4472 -7607 4485 -7561
rect 4531 -7607 4544 -7561
rect 4472 -7642 4544 -7607
rect 430 -7655 4544 -7642
rect 430 -7701 443 -7655
rect 489 -7701 537 -7655
rect 583 -7701 631 -7655
rect 677 -7701 725 -7655
rect 771 -7701 819 -7655
rect 865 -7701 913 -7655
rect 959 -7701 1007 -7655
rect 1053 -7701 1101 -7655
rect 1147 -7701 1195 -7655
rect 1241 -7701 1289 -7655
rect 1335 -7701 1383 -7655
rect 1429 -7701 1477 -7655
rect 1523 -7701 1571 -7655
rect 1617 -7701 1665 -7655
rect 1711 -7701 1759 -7655
rect 1805 -7701 1853 -7655
rect 1899 -7701 1947 -7655
rect 1993 -7701 2041 -7655
rect 2087 -7701 2135 -7655
rect 2181 -7701 2229 -7655
rect 2275 -7701 2323 -7655
rect 2369 -7701 2417 -7655
rect 2463 -7701 2511 -7655
rect 2557 -7701 2605 -7655
rect 2651 -7701 2699 -7655
rect 2745 -7701 2793 -7655
rect 2839 -7701 2887 -7655
rect 2933 -7701 2981 -7655
rect 3027 -7701 3075 -7655
rect 3121 -7701 3169 -7655
rect 3215 -7701 3263 -7655
rect 3309 -7701 3357 -7655
rect 3403 -7701 3451 -7655
rect 3497 -7701 3545 -7655
rect 3591 -7701 3639 -7655
rect 3685 -7701 3733 -7655
rect 3779 -7701 3827 -7655
rect 3873 -7701 3921 -7655
rect 3967 -7701 4015 -7655
rect 4061 -7701 4109 -7655
rect 4155 -7701 4203 -7655
rect 4249 -7701 4297 -7655
rect 4343 -7701 4391 -7655
rect 4437 -7701 4485 -7655
rect 4531 -7701 4544 -7655
rect 430 -7714 4544 -7701
rect 17707 -4678 17779 -4630
rect 17707 -4724 17720 -4678
rect 17766 -4724 17779 -4678
rect 17707 -4772 17779 -4724
rect 17707 -4818 17720 -4772
rect 17766 -4818 17779 -4772
rect 17707 -4866 17779 -4818
rect 17707 -4912 17720 -4866
rect 17766 -4912 17779 -4866
rect 17707 -4960 17779 -4912
rect 17707 -5006 17720 -4960
rect 17766 -5006 17779 -4960
rect 22501 -4396 22573 -4348
rect 22501 -4442 22514 -4396
rect 22560 -4442 22573 -4396
rect 22501 -4490 22573 -4442
rect 22501 -4536 22514 -4490
rect 22560 -4536 22573 -4490
rect 22501 -4584 22573 -4536
rect 22501 -4630 22514 -4584
rect 22560 -4630 22573 -4584
rect 22501 -4678 22573 -4630
rect 22501 -4724 22514 -4678
rect 22560 -4724 22573 -4678
rect 22501 -4772 22573 -4724
rect 22501 -4818 22514 -4772
rect 22560 -4818 22573 -4772
rect 22501 -4866 22573 -4818
rect 22501 -4912 22514 -4866
rect 22560 -4912 22573 -4866
rect 22501 -4960 22573 -4912
rect 17707 -5054 17779 -5006
rect 17707 -5100 17720 -5054
rect 17766 -5100 17779 -5054
rect 17707 -5148 17779 -5100
rect 17707 -5194 17720 -5148
rect 17766 -5194 17779 -5148
rect 17707 -5242 17779 -5194
rect 17707 -5288 17720 -5242
rect 17766 -5288 17779 -5242
rect 17707 -5336 17779 -5288
rect 17707 -5382 17720 -5336
rect 17766 -5382 17779 -5336
rect 17707 -5430 17779 -5382
rect 17707 -5476 17720 -5430
rect 17766 -5476 17779 -5430
rect 17707 -5524 17779 -5476
rect 17707 -5570 17720 -5524
rect 17766 -5570 17779 -5524
rect 17707 -5618 17779 -5570
rect 17707 -5664 17720 -5618
rect 17766 -5664 17779 -5618
rect 17707 -5712 17779 -5664
rect 17707 -5758 17720 -5712
rect 17766 -5758 17779 -5712
rect 17707 -5806 17779 -5758
rect 17707 -5852 17720 -5806
rect 17766 -5852 17779 -5806
rect 17707 -5900 17779 -5852
rect 17707 -5946 17720 -5900
rect 17766 -5946 17779 -5900
rect 17707 -5994 17779 -5946
rect 17707 -6040 17720 -5994
rect 17766 -6040 17779 -5994
rect 17707 -6088 17779 -6040
rect 17707 -6134 17720 -6088
rect 17766 -6134 17779 -6088
rect 17707 -6182 17779 -6134
rect 17707 -6228 17720 -6182
rect 17766 -6228 17779 -6182
rect 17707 -6276 17779 -6228
rect 17707 -6322 17720 -6276
rect 17766 -6322 17779 -6276
rect 17707 -6370 17779 -6322
rect 17707 -6416 17720 -6370
rect 17766 -6416 17779 -6370
rect 17707 -6464 17779 -6416
rect 17707 -6510 17720 -6464
rect 17766 -6510 17779 -6464
rect 17707 -6558 17779 -6510
rect 17707 -6604 17720 -6558
rect 17766 -6604 17779 -6558
rect 22501 -5006 22514 -4960
rect 22560 -5006 22573 -4960
rect 22501 -5054 22573 -5006
rect 17707 -6652 17779 -6604
rect 17707 -6698 17720 -6652
rect 17766 -6698 17779 -6652
rect 22501 -5100 22514 -5054
rect 22560 -5100 22573 -5054
rect 22501 -5148 22573 -5100
rect 22501 -5194 22514 -5148
rect 22560 -5194 22573 -5148
rect 22501 -5242 22573 -5194
rect 22501 -5288 22514 -5242
rect 22560 -5288 22573 -5242
rect 22501 -5336 22573 -5288
rect 22501 -5382 22514 -5336
rect 22560 -5382 22573 -5336
rect 22501 -5430 22573 -5382
rect 22501 -5476 22514 -5430
rect 22560 -5476 22573 -5430
rect 22501 -5524 22573 -5476
rect 22501 -5570 22514 -5524
rect 22560 -5570 22573 -5524
rect 22501 -5618 22573 -5570
rect 22501 -5664 22514 -5618
rect 22560 -5664 22573 -5618
rect 22501 -5712 22573 -5664
rect 22501 -5758 22514 -5712
rect 22560 -5758 22573 -5712
rect 22501 -5806 22573 -5758
rect 22501 -5852 22514 -5806
rect 22560 -5852 22573 -5806
rect 22501 -5900 22573 -5852
rect 22501 -5946 22514 -5900
rect 22560 -5946 22573 -5900
rect 22501 -5994 22573 -5946
rect 22501 -6040 22514 -5994
rect 22560 -6040 22573 -5994
rect 22501 -6088 22573 -6040
rect 22501 -6134 22514 -6088
rect 22560 -6134 22573 -6088
rect 22501 -6182 22573 -6134
rect 22501 -6228 22514 -6182
rect 22560 -6228 22573 -6182
rect 22501 -6276 22573 -6228
rect 22501 -6322 22514 -6276
rect 22560 -6322 22573 -6276
rect 22501 -6370 22573 -6322
rect 22501 -6416 22514 -6370
rect 22560 -6416 22573 -6370
rect 22501 -6464 22573 -6416
rect 22501 -6510 22514 -6464
rect 22560 -6510 22573 -6464
rect 22501 -6558 22573 -6510
rect 22501 -6604 22514 -6558
rect 22560 -6604 22573 -6558
rect 22501 -6652 22573 -6604
rect 17707 -6746 17779 -6698
rect 17707 -6792 17720 -6746
rect 17766 -6792 17779 -6746
rect 17707 -6840 17779 -6792
rect 17707 -6886 17720 -6840
rect 17766 -6886 17779 -6840
rect 17707 -6934 17779 -6886
rect 17707 -6980 17720 -6934
rect 17766 -6980 17779 -6934
rect 17707 -7028 17779 -6980
rect 17707 -7074 17720 -7028
rect 17766 -7074 17779 -7028
rect 17707 -7122 17779 -7074
rect 17707 -7168 17720 -7122
rect 17766 -7168 17779 -7122
rect 17707 -7216 17779 -7168
rect 22501 -6698 22514 -6652
rect 22560 -6698 22573 -6652
rect 22501 -6746 22573 -6698
rect 22501 -6792 22514 -6746
rect 22560 -6792 22573 -6746
rect 22501 -6840 22573 -6792
rect 22501 -6886 22514 -6840
rect 22560 -6886 22573 -6840
rect 22501 -6934 22573 -6886
rect 22501 -6980 22514 -6934
rect 22560 -6980 22573 -6934
rect 22501 -7028 22573 -6980
rect 22501 -7074 22514 -7028
rect 22560 -7074 22573 -7028
rect 22501 -7122 22573 -7074
rect 22501 -7168 22514 -7122
rect 22560 -7168 22573 -7122
rect 17707 -7262 17720 -7216
rect 17766 -7262 17779 -7216
rect 17707 -7310 17779 -7262
rect 17707 -7356 17720 -7310
rect 17766 -7356 17779 -7310
rect 22501 -7216 22573 -7168
rect 22501 -7262 22514 -7216
rect 22560 -7262 22573 -7216
rect 22501 -7310 22573 -7262
rect 17707 -7404 17779 -7356
rect 17707 -7450 17720 -7404
rect 17766 -7450 17779 -7404
rect 17707 -7498 17779 -7450
rect 17707 -7544 17720 -7498
rect 17766 -7544 17779 -7498
rect 17707 -7592 17779 -7544
rect 17707 -7638 17720 -7592
rect 17766 -7638 17779 -7592
rect 17707 -7686 17779 -7638
rect 17707 -7732 17720 -7686
rect 17766 -7732 17779 -7686
rect 17707 -7780 17779 -7732
rect 17707 -7826 17720 -7780
rect 17766 -7826 17779 -7780
rect 17707 -7874 17779 -7826
rect 17707 -7920 17720 -7874
rect 17766 -7920 17779 -7874
rect 17707 -7968 17779 -7920
rect 17707 -8014 17720 -7968
rect 17766 -8014 17779 -7968
rect 17707 -8049 17779 -8014
rect 22501 -7356 22514 -7310
rect 22560 -7356 22573 -7310
rect 22501 -7404 22573 -7356
rect 22501 -7450 22514 -7404
rect 22560 -7450 22573 -7404
rect 22501 -7498 22573 -7450
rect 22501 -7544 22514 -7498
rect 22560 -7544 22573 -7498
rect 22501 -7592 22573 -7544
rect 22501 -7638 22514 -7592
rect 22560 -7638 22573 -7592
rect 22501 -7686 22573 -7638
rect 22501 -7732 22514 -7686
rect 22560 -7732 22573 -7686
rect 22501 -7780 22573 -7732
rect 22501 -7826 22514 -7780
rect 22560 -7826 22573 -7780
rect 22501 -7874 22573 -7826
rect 22501 -7920 22514 -7874
rect 22560 -7920 22573 -7874
rect 22501 -7968 22573 -7920
rect 22501 -8014 22514 -7968
rect 22560 -8014 22573 -7968
rect 22501 -8049 22573 -8014
rect 28235 -3550 28307 -3515
rect 28235 -3596 28248 -3550
rect 28294 -3596 28307 -3550
rect 28235 -3644 28307 -3596
rect 28235 -3690 28248 -3644
rect 28294 -3690 28307 -3644
rect 28235 -3738 28307 -3690
rect 28235 -3784 28248 -3738
rect 28294 -3784 28307 -3738
rect 28235 -3832 28307 -3784
rect 28235 -3878 28248 -3832
rect 28294 -3878 28307 -3832
rect 28235 -3926 28307 -3878
rect 28235 -3972 28248 -3926
rect 28294 -3972 28307 -3926
rect 28235 -4020 28307 -3972
rect 28235 -4066 28248 -4020
rect 28294 -4066 28307 -4020
rect 28235 -4114 28307 -4066
rect 28235 -4160 28248 -4114
rect 28294 -4160 28307 -4114
rect 28235 -4208 28307 -4160
rect 28235 -4254 28248 -4208
rect 28294 -4254 28307 -4208
rect 28235 -4302 28307 -4254
rect 28235 -4348 28248 -4302
rect 28294 -4348 28307 -4302
rect 28235 -4396 28307 -4348
rect 28235 -4442 28248 -4396
rect 28294 -4442 28307 -4396
rect 28235 -4490 28307 -4442
rect 28235 -4536 28248 -4490
rect 28294 -4536 28307 -4490
rect 28235 -4584 28307 -4536
rect 28235 -4630 28248 -4584
rect 28294 -4630 28307 -4584
rect 28235 -4678 28307 -4630
rect 28235 -4724 28248 -4678
rect 28294 -4724 28307 -4678
rect 28235 -4772 28307 -4724
rect 28235 -4818 28248 -4772
rect 28294 -4818 28307 -4772
rect 28235 -4866 28307 -4818
rect 28235 -4912 28248 -4866
rect 28294 -4912 28307 -4866
rect 28235 -4960 28307 -4912
rect 28235 -5006 28248 -4960
rect 28294 -5006 28307 -4960
rect 28235 -5054 28307 -5006
rect 28235 -5100 28248 -5054
rect 28294 -5100 28307 -5054
rect 28235 -5148 28307 -5100
rect 28235 -5194 28248 -5148
rect 28294 -5194 28307 -5148
rect 28235 -5242 28307 -5194
rect 28235 -5288 28248 -5242
rect 28294 -5288 28307 -5242
rect 28235 -5336 28307 -5288
rect 28235 -5382 28248 -5336
rect 28294 -5382 28307 -5336
rect 28235 -5430 28307 -5382
rect 28235 -5476 28248 -5430
rect 28294 -5476 28307 -5430
rect 28235 -5524 28307 -5476
rect 28235 -5570 28248 -5524
rect 28294 -5570 28307 -5524
rect 28235 -5618 28307 -5570
rect 28235 -5664 28248 -5618
rect 28294 -5664 28307 -5618
rect 28235 -5712 28307 -5664
rect 28235 -5758 28248 -5712
rect 28294 -5758 28307 -5712
rect 28235 -5806 28307 -5758
rect 28235 -5852 28248 -5806
rect 28294 -5852 28307 -5806
rect 28235 -5900 28307 -5852
rect 28235 -5946 28248 -5900
rect 28294 -5946 28307 -5900
rect 28235 -5994 28307 -5946
rect 28235 -6040 28248 -5994
rect 28294 -6040 28307 -5994
rect 28235 -6088 28307 -6040
rect 28235 -6134 28248 -6088
rect 28294 -6134 28307 -6088
rect 28235 -6182 28307 -6134
rect 28235 -6228 28248 -6182
rect 28294 -6228 28307 -6182
rect 28235 -6276 28307 -6228
rect 28235 -6322 28248 -6276
rect 28294 -6322 28307 -6276
rect 28235 -6370 28307 -6322
rect 28235 -6416 28248 -6370
rect 28294 -6416 28307 -6370
rect 28235 -6464 28307 -6416
rect 28235 -6510 28248 -6464
rect 28294 -6510 28307 -6464
rect 28235 -6558 28307 -6510
rect 28235 -6604 28248 -6558
rect 28294 -6604 28307 -6558
rect 28235 -6652 28307 -6604
rect 28235 -6698 28248 -6652
rect 28294 -6698 28307 -6652
rect 28235 -6746 28307 -6698
rect 28235 -6792 28248 -6746
rect 28294 -6792 28307 -6746
rect 28235 -6840 28307 -6792
rect 28235 -6886 28248 -6840
rect 28294 -6886 28307 -6840
rect 28235 -6934 28307 -6886
rect 28235 -6980 28248 -6934
rect 28294 -6980 28307 -6934
rect 28235 -7028 28307 -6980
rect 28235 -7074 28248 -7028
rect 28294 -7074 28307 -7028
rect 28235 -7122 28307 -7074
rect 28235 -7168 28248 -7122
rect 28294 -7168 28307 -7122
rect 28235 -7216 28307 -7168
rect 28235 -7262 28248 -7216
rect 28294 -7262 28307 -7216
rect 28235 -7310 28307 -7262
rect 28235 -7356 28248 -7310
rect 28294 -7356 28307 -7310
rect 28235 -7404 28307 -7356
rect 28235 -7450 28248 -7404
rect 28294 -7450 28307 -7404
rect 28235 -7498 28307 -7450
rect 28235 -7544 28248 -7498
rect 28294 -7544 28307 -7498
rect 28235 -7592 28307 -7544
rect 28235 -7638 28248 -7592
rect 28294 -7638 28307 -7592
rect 28235 -7686 28307 -7638
rect 28235 -7732 28248 -7686
rect 28294 -7732 28307 -7686
rect 28235 -7780 28307 -7732
rect 28235 -7826 28248 -7780
rect 28294 -7826 28307 -7780
rect 28235 -7874 28307 -7826
rect 28235 -7920 28248 -7874
rect 28294 -7920 28307 -7874
rect 28235 -7968 28307 -7920
rect 28235 -8014 28248 -7968
rect 28294 -8014 28307 -7968
rect 28235 -8049 28307 -8014
rect 31243 -3550 31315 -3515
rect 31243 -3596 31256 -3550
rect 31302 -3596 31315 -3550
rect 31243 -3644 31315 -3596
rect 31243 -3690 31256 -3644
rect 31302 -3690 31315 -3644
rect 31243 -3738 31315 -3690
rect 31243 -3784 31256 -3738
rect 31302 -3784 31315 -3738
rect 31243 -3832 31315 -3784
rect 31243 -3878 31256 -3832
rect 31302 -3878 31315 -3832
rect 31243 -3926 31315 -3878
rect 31243 -3972 31256 -3926
rect 31302 -3972 31315 -3926
rect 31243 -4020 31315 -3972
rect 31243 -4066 31256 -4020
rect 31302 -4066 31315 -4020
rect 31243 -4114 31315 -4066
rect 31243 -4160 31256 -4114
rect 31302 -4160 31315 -4114
rect 31243 -4208 31315 -4160
rect 31243 -4254 31256 -4208
rect 31302 -4254 31315 -4208
rect 31243 -4302 31315 -4254
rect 31243 -4348 31256 -4302
rect 31302 -4348 31315 -4302
rect 31243 -4396 31315 -4348
rect 31243 -4442 31256 -4396
rect 31302 -4442 31315 -4396
rect 31243 -4490 31315 -4442
rect 31243 -4536 31256 -4490
rect 31302 -4536 31315 -4490
rect 31243 -4584 31315 -4536
rect 31243 -4630 31256 -4584
rect 31302 -4630 31315 -4584
rect 31243 -4678 31315 -4630
rect 31243 -4724 31256 -4678
rect 31302 -4724 31315 -4678
rect 31243 -4772 31315 -4724
rect 31243 -4818 31256 -4772
rect 31302 -4818 31315 -4772
rect 31243 -4866 31315 -4818
rect 31243 -4912 31256 -4866
rect 31302 -4912 31315 -4866
rect 31243 -4960 31315 -4912
rect 31243 -5006 31256 -4960
rect 31302 -5006 31315 -4960
rect 31243 -5054 31315 -5006
rect 31243 -5100 31256 -5054
rect 31302 -5100 31315 -5054
rect 31243 -5148 31315 -5100
rect 31243 -5194 31256 -5148
rect 31302 -5194 31315 -5148
rect 31243 -5242 31315 -5194
rect 31243 -5288 31256 -5242
rect 31302 -5288 31315 -5242
rect 31243 -5336 31315 -5288
rect 31243 -5382 31256 -5336
rect 31302 -5382 31315 -5336
rect 31243 -5430 31315 -5382
rect 31243 -5476 31256 -5430
rect 31302 -5476 31315 -5430
rect 31243 -5524 31315 -5476
rect 31243 -5570 31256 -5524
rect 31302 -5570 31315 -5524
rect 31243 -5618 31315 -5570
rect 31243 -5664 31256 -5618
rect 31302 -5664 31315 -5618
rect 31243 -5712 31315 -5664
rect 31243 -5758 31256 -5712
rect 31302 -5758 31315 -5712
rect 31243 -5806 31315 -5758
rect 31243 -5852 31256 -5806
rect 31302 -5852 31315 -5806
rect 31243 -5900 31315 -5852
rect 31243 -5946 31256 -5900
rect 31302 -5946 31315 -5900
rect 31243 -5994 31315 -5946
rect 31243 -6040 31256 -5994
rect 31302 -6040 31315 -5994
rect 31243 -6088 31315 -6040
rect 31243 -6134 31256 -6088
rect 31302 -6134 31315 -6088
rect 31243 -6182 31315 -6134
rect 31243 -6228 31256 -6182
rect 31302 -6228 31315 -6182
rect 31243 -6276 31315 -6228
rect 31243 -6322 31256 -6276
rect 31302 -6322 31315 -6276
rect 31243 -6370 31315 -6322
rect 31243 -6416 31256 -6370
rect 31302 -6416 31315 -6370
rect 31243 -6464 31315 -6416
rect 31243 -6510 31256 -6464
rect 31302 -6510 31315 -6464
rect 31243 -6558 31315 -6510
rect 31243 -6604 31256 -6558
rect 31302 -6604 31315 -6558
rect 31243 -6652 31315 -6604
rect 31243 -6698 31256 -6652
rect 31302 -6698 31315 -6652
rect 31243 -6746 31315 -6698
rect 31243 -6792 31256 -6746
rect 31302 -6792 31315 -6746
rect 31243 -6840 31315 -6792
rect 31243 -6886 31256 -6840
rect 31302 -6886 31315 -6840
rect 31243 -6934 31315 -6886
rect 31243 -6980 31256 -6934
rect 31302 -6980 31315 -6934
rect 31243 -7028 31315 -6980
rect 31243 -7074 31256 -7028
rect 31302 -7074 31315 -7028
rect 31243 -7122 31315 -7074
rect 31243 -7168 31256 -7122
rect 31302 -7168 31315 -7122
rect 31243 -7216 31315 -7168
rect 31243 -7262 31256 -7216
rect 31302 -7262 31315 -7216
rect 31243 -7310 31315 -7262
rect 31243 -7356 31256 -7310
rect 31302 -7356 31315 -7310
rect 31243 -7404 31315 -7356
rect 31243 -7450 31256 -7404
rect 31302 -7450 31315 -7404
rect 31243 -7498 31315 -7450
rect 31243 -7544 31256 -7498
rect 31302 -7544 31315 -7498
rect 31243 -7592 31315 -7544
rect 31243 -7638 31256 -7592
rect 31302 -7638 31315 -7592
rect 31243 -7686 31315 -7638
rect 31243 -7732 31256 -7686
rect 31302 -7732 31315 -7686
rect 31243 -7780 31315 -7732
rect 31243 -7826 31256 -7780
rect 31302 -7826 31315 -7780
rect 31243 -7874 31315 -7826
rect 31243 -7920 31256 -7874
rect 31302 -7920 31315 -7874
rect 31243 -7968 31315 -7920
rect 31243 -8014 31256 -7968
rect 31302 -8014 31315 -7968
rect 31243 -8049 31315 -8014
rect 17707 -8062 31315 -8049
rect 17707 -8108 17720 -8062
rect 17766 -8108 17814 -8062
rect 17860 -8108 17908 -8062
rect 17954 -8108 18002 -8062
rect 18048 -8108 18096 -8062
rect 18142 -8108 18190 -8062
rect 18236 -8108 18284 -8062
rect 18330 -8108 18378 -8062
rect 18424 -8108 18472 -8062
rect 18518 -8108 18566 -8062
rect 18612 -8108 18660 -8062
rect 18706 -8108 18754 -8062
rect 18800 -8108 18848 -8062
rect 18894 -8108 18942 -8062
rect 18988 -8108 19036 -8062
rect 19082 -8108 19130 -8062
rect 19176 -8108 19224 -8062
rect 19270 -8108 19318 -8062
rect 19364 -8108 19412 -8062
rect 19458 -8108 19506 -8062
rect 19552 -8108 19600 -8062
rect 19646 -8108 19694 -8062
rect 19740 -8108 19788 -8062
rect 19834 -8108 19882 -8062
rect 19928 -8108 19976 -8062
rect 20022 -8108 20070 -8062
rect 20116 -8108 20164 -8062
rect 20210 -8108 20258 -8062
rect 20304 -8108 20352 -8062
rect 20398 -8108 20446 -8062
rect 20492 -8108 20540 -8062
rect 20586 -8108 20634 -8062
rect 20680 -8108 20728 -8062
rect 20774 -8108 20822 -8062
rect 20868 -8108 20916 -8062
rect 20962 -8108 21010 -8062
rect 21056 -8108 21104 -8062
rect 21150 -8108 21198 -8062
rect 21244 -8108 21292 -8062
rect 21338 -8108 21386 -8062
rect 21432 -8108 21480 -8062
rect 21526 -8108 21574 -8062
rect 21620 -8108 21668 -8062
rect 21714 -8108 21762 -8062
rect 21808 -8108 21856 -8062
rect 21902 -8108 21950 -8062
rect 21996 -8108 22044 -8062
rect 22090 -8108 22138 -8062
rect 22184 -8108 22232 -8062
rect 22278 -8108 22326 -8062
rect 22372 -8108 22420 -8062
rect 22466 -8108 22514 -8062
rect 22560 -8108 22608 -8062
rect 22654 -8108 22702 -8062
rect 22748 -8108 22796 -8062
rect 22842 -8108 22890 -8062
rect 22936 -8108 22984 -8062
rect 23030 -8108 23078 -8062
rect 23124 -8108 23172 -8062
rect 23218 -8108 23266 -8062
rect 23312 -8108 23360 -8062
rect 23406 -8108 23454 -8062
rect 23500 -8108 23548 -8062
rect 23594 -8108 23642 -8062
rect 23688 -8108 23736 -8062
rect 23782 -8108 23830 -8062
rect 23876 -8108 23924 -8062
rect 23970 -8108 24018 -8062
rect 24064 -8108 24112 -8062
rect 24158 -8108 24206 -8062
rect 24252 -8108 24300 -8062
rect 24346 -8108 24394 -8062
rect 24440 -8108 24488 -8062
rect 24534 -8108 24582 -8062
rect 24628 -8108 24676 -8062
rect 24722 -8108 24770 -8062
rect 24816 -8108 24864 -8062
rect 24910 -8108 24958 -8062
rect 25004 -8108 25052 -8062
rect 25098 -8108 25146 -8062
rect 25192 -8108 25240 -8062
rect 25286 -8108 25334 -8062
rect 25380 -8108 25428 -8062
rect 25474 -8108 25522 -8062
rect 25568 -8108 25616 -8062
rect 25662 -8108 25710 -8062
rect 25756 -8108 25804 -8062
rect 25850 -8108 25898 -8062
rect 25944 -8108 25992 -8062
rect 26038 -8108 26086 -8062
rect 26132 -8108 26180 -8062
rect 26226 -8108 26274 -8062
rect 26320 -8108 26368 -8062
rect 26414 -8108 26462 -8062
rect 26508 -8108 26556 -8062
rect 26602 -8108 26650 -8062
rect 26696 -8108 26744 -8062
rect 26790 -8108 26838 -8062
rect 26884 -8108 26932 -8062
rect 26978 -8108 27026 -8062
rect 27072 -8108 27120 -8062
rect 27166 -8108 27214 -8062
rect 27260 -8108 27308 -8062
rect 27354 -8108 27402 -8062
rect 27448 -8108 27496 -8062
rect 27542 -8108 27590 -8062
rect 27636 -8108 27684 -8062
rect 27730 -8108 27778 -8062
rect 27824 -8108 27872 -8062
rect 27918 -8108 27966 -8062
rect 28012 -8108 28060 -8062
rect 28106 -8108 28154 -8062
rect 28200 -8108 28248 -8062
rect 28294 -8108 28342 -8062
rect 28388 -8108 28436 -8062
rect 28482 -8108 28530 -8062
rect 28576 -8108 28624 -8062
rect 28670 -8108 28718 -8062
rect 28764 -8108 28812 -8062
rect 28858 -8108 28906 -8062
rect 28952 -8108 29000 -8062
rect 29046 -8108 29094 -8062
rect 29140 -8108 29188 -8062
rect 29234 -8108 29282 -8062
rect 29328 -8108 29376 -8062
rect 29422 -8108 29470 -8062
rect 29516 -8108 29564 -8062
rect 29610 -8108 29658 -8062
rect 29704 -8108 29752 -8062
rect 29798 -8108 29846 -8062
rect 29892 -8108 29940 -8062
rect 29986 -8108 30034 -8062
rect 30080 -8108 30128 -8062
rect 30174 -8108 30222 -8062
rect 30268 -8108 30316 -8062
rect 30362 -8108 30410 -8062
rect 30456 -8108 30504 -8062
rect 30550 -8108 30598 -8062
rect 30644 -8108 30692 -8062
rect 30738 -8108 30786 -8062
rect 30832 -8108 30880 -8062
rect 30926 -8108 30974 -8062
rect 31020 -8108 31068 -8062
rect 31114 -8108 31162 -8062
rect 31208 -8108 31256 -8062
rect 31302 -8108 31315 -8062
rect 17707 -8121 31315 -8108
<< psubdiffcont >>
rect 5776 5462 5822 5508
rect 5870 5462 5916 5508
rect 5964 5462 6010 5508
rect 6058 5462 6104 5508
rect 6152 5462 6198 5508
rect 6246 5462 6292 5508
rect 6340 5462 6386 5508
rect 6434 5462 6480 5508
rect 6528 5462 6574 5508
rect 6622 5462 6668 5508
rect 6716 5462 6762 5508
rect 6810 5462 6856 5508
rect 6904 5462 6950 5508
rect 6998 5462 7044 5508
rect 7092 5462 7138 5508
rect 7186 5462 7232 5508
rect 7280 5462 7326 5508
rect 7374 5462 7420 5508
rect 7468 5462 7514 5508
rect 7562 5462 7608 5508
rect 7656 5462 7702 5508
rect 7750 5462 7796 5508
rect 7844 5462 7890 5508
rect 7938 5462 7984 5508
rect 8032 5462 8078 5508
rect 5776 5368 5822 5414
rect 5776 5274 5822 5320
rect 5776 5180 5822 5226
rect 5776 5086 5822 5132
rect 5776 4992 5822 5038
rect 5776 4898 5822 4944
rect 5776 4804 5822 4850
rect 5776 4710 5822 4756
rect 5776 4616 5822 4662
rect 5776 4522 5822 4568
rect 8032 5368 8078 5414
rect 8032 5274 8078 5320
rect 8032 5180 8078 5226
rect 8032 5086 8078 5132
rect 8032 4992 8078 5038
rect 8032 4898 8078 4944
rect 8032 4804 8078 4850
rect 8032 4710 8078 4756
rect 8032 4616 8078 4662
rect 5776 4428 5822 4474
rect 5776 4334 5822 4380
rect 5776 4240 5822 4286
rect 8032 4522 8078 4568
rect 8032 4428 8078 4474
rect 8032 4334 8078 4380
rect 5776 4146 5822 4192
rect 5776 4052 5822 4098
rect 5776 3958 5822 4004
rect 5776 3864 5822 3910
rect 5776 3770 5822 3816
rect 5776 3676 5822 3722
rect 8032 4240 8078 4286
rect 8032 4146 8078 4192
rect 8032 4052 8078 4098
rect 8032 3958 8078 4004
rect 8032 3864 8078 3910
rect 8032 3770 8078 3816
rect 5776 3582 5822 3628
rect 5776 3488 5822 3534
rect 5776 3394 5822 3440
rect 8032 3676 8078 3722
rect 8032 3582 8078 3628
rect 8032 3488 8078 3534
rect 5776 3291 5822 3346
rect 5776 3197 5822 3243
rect 5776 3103 5822 3149
rect 5776 3009 5822 3055
rect 5776 2915 5822 2961
rect 5776 2821 5822 2867
rect 8032 3394 8078 3440
rect 8032 3291 8078 3346
rect 8032 3197 8078 3243
rect 8032 3103 8078 3149
rect 8032 3009 8078 3055
rect 8032 2915 8078 2961
rect 8032 2821 8078 2867
rect 5776 2727 5822 2773
rect 5776 2633 5822 2679
rect 5776 2539 5822 2585
rect 8032 2727 8078 2773
rect 8032 2633 8078 2679
rect 17650 4565 17696 4611
rect 17744 4565 17790 4611
rect 17838 4565 17884 4611
rect 17932 4565 17978 4611
rect 18026 4565 18072 4611
rect 18120 4565 18166 4611
rect 18214 4565 18260 4611
rect 18308 4565 18354 4611
rect 18402 4565 18448 4611
rect 18496 4565 18542 4611
rect 18590 4565 18636 4611
rect 18684 4565 18730 4611
rect 18778 4565 18824 4611
rect 18872 4565 18918 4611
rect 18966 4565 19012 4611
rect 19060 4565 19106 4611
rect 19154 4565 19200 4611
rect 19248 4565 19294 4611
rect 19342 4565 19388 4611
rect 19436 4565 19482 4611
rect 19530 4565 19576 4611
rect 19624 4565 19670 4611
rect 19718 4565 19764 4611
rect 19812 4565 19858 4611
rect 19906 4565 19952 4611
rect 20000 4565 20046 4611
rect 20094 4565 20140 4611
rect 20188 4565 20234 4611
rect 20282 4565 20328 4611
rect 20376 4565 20422 4611
rect 20470 4565 20516 4611
rect 20564 4565 20610 4611
rect 20658 4565 20704 4611
rect 17650 4471 17696 4517
rect 17650 4377 17696 4423
rect 17650 4283 17696 4329
rect 20658 4471 20704 4517
rect 20658 4377 20704 4423
rect 20658 4283 20704 4329
rect 17650 4189 17696 4235
rect 20658 4189 20704 4235
rect 17650 4095 17696 4141
rect 17650 4001 17696 4047
rect 20658 4095 20704 4141
rect 17650 3907 17696 3953
rect 17650 3813 17696 3859
rect 17650 3719 17696 3765
rect 17650 3625 17696 3671
rect 17650 3531 17696 3577
rect 17650 3437 17696 3483
rect 20658 4001 20704 4047
rect 20658 3907 20704 3953
rect 20658 3813 20704 3859
rect 20658 3719 20704 3765
rect 20658 3625 20704 3671
rect 20658 3531 20704 3577
rect 20658 3437 20704 3483
rect 17650 3343 17696 3389
rect 17650 3249 17696 3295
rect 20658 3343 20704 3389
rect 17650 3155 17696 3201
rect 17650 3061 17696 3107
rect 17650 2967 17696 3013
rect 17650 2873 17696 2919
rect 17650 2779 17696 2825
rect 17650 2685 17696 2731
rect 8032 2539 8078 2585
rect 5776 2445 5822 2491
rect 5776 2351 5822 2397
rect 5776 2257 5822 2303
rect 5776 2163 5822 2209
rect 5776 2069 5822 2115
rect 5776 1975 5822 2021
rect 8032 2445 8078 2491
rect 8032 2351 8078 2397
rect 8032 2257 8078 2303
rect 8032 2163 8078 2209
rect 8032 2069 8078 2115
rect 8032 1975 8078 2021
rect 8126 1975 8172 2021
rect 8220 1975 8266 2021
rect 8314 1975 8360 2021
rect 8408 1975 8454 2021
rect 8502 1975 8548 2021
rect 8596 1975 8642 2021
rect 8690 1975 8736 2021
rect 8784 1975 8830 2021
rect 8878 1975 8924 2021
rect 8972 1975 9018 2021
rect 9066 1975 9112 2021
rect 9160 1975 9206 2021
rect 9254 1975 9300 2021
rect 9348 1975 9394 2021
rect 9442 1975 9488 2021
rect 9536 1975 9582 2021
rect 9630 1975 9676 2021
rect 9724 1975 9770 2021
rect 9818 1975 9864 2021
rect 9912 1975 9958 2021
rect 10006 1975 10052 2021
rect 10100 1975 10146 2021
rect 10194 1975 10240 2021
rect 10288 1975 10334 2021
rect 10382 1975 10428 2021
rect 10476 1975 10522 2021
rect 10570 1975 10616 2021
rect 10664 1975 10710 2021
rect 10758 1975 10804 2021
rect 5776 1881 5822 1927
rect 5776 1787 5822 1833
rect 5776 1693 5822 1739
rect 8032 1881 8078 1927
rect 8032 1787 8078 1833
rect 8032 1693 8078 1739
rect 5776 1599 5822 1645
rect 5776 1505 5822 1551
rect 5776 1411 5822 1457
rect 5776 1317 5822 1363
rect 5776 1223 5822 1269
rect 5776 1129 5822 1175
rect 8032 1599 8078 1645
rect 8032 1505 8078 1551
rect 8032 1411 8078 1457
rect 8032 1317 8078 1363
rect 8032 1223 8078 1269
rect 8032 1129 8078 1175
rect 5776 1035 5822 1081
rect 5776 941 5822 987
rect 5776 847 5822 893
rect 8032 1035 8078 1081
rect 10758 1881 10804 1927
rect 10758 1787 10804 1833
rect 10758 1693 10804 1739
rect 10758 1599 10804 1645
rect 10758 1505 10804 1551
rect 10758 1411 10804 1457
rect 10758 1317 10804 1363
rect 10758 1223 10804 1269
rect 10758 1129 10804 1175
rect 8032 941 8078 987
rect 8032 847 8078 893
rect 5776 753 5822 799
rect 5776 659 5822 705
rect 5776 565 5822 611
rect 5776 471 5822 517
rect 5776 377 5822 423
rect 5776 283 5822 329
rect 5776 189 5822 235
rect 8032 753 8078 799
rect 10758 1035 10804 1081
rect 10758 941 10804 987
rect 10758 847 10804 893
rect 8032 659 8078 705
rect 8032 565 8078 611
rect 8032 471 8078 517
rect 8032 377 8078 423
rect 8032 283 8078 329
rect 5776 95 5822 141
rect 5776 1 5822 47
rect 5776 -93 5822 -47
rect 8032 189 8078 235
rect 10758 753 10804 799
rect 10758 659 10804 705
rect 10758 565 10804 611
rect 10758 471 10804 517
rect 10758 377 10804 423
rect 10758 283 10804 329
rect 8032 95 8078 141
rect 8032 1 8078 47
rect 5776 -187 5822 -141
rect 5776 -281 5822 -235
rect 5776 -375 5822 -329
rect 5776 -469 5822 -423
rect 5776 -563 5822 -517
rect 5776 -657 5822 -611
rect 8032 -93 8078 -47
rect 10758 189 10804 235
rect 10758 95 10804 141
rect 10758 1 10804 47
rect 8032 -187 8078 -141
rect 8032 -281 8078 -235
rect 8032 -375 8078 -329
rect 8032 -469 8078 -423
rect 8032 -563 8078 -517
rect 5776 -751 5822 -705
rect 5776 -845 5822 -799
rect 8032 -657 8078 -611
rect 10758 -93 10804 -47
rect 10758 -187 10804 -141
rect 10758 -281 10804 -235
rect 10758 -375 10804 -329
rect 10758 -469 10804 -423
rect 10758 -563 10804 -517
rect 5776 -939 5822 -893
rect 8032 -751 8078 -705
rect 8032 -845 8078 -799
rect 10758 -657 10804 -611
rect 10758 -751 10804 -705
rect 5776 -1033 5822 -987
rect 5776 -1127 5822 -1081
rect 5776 -1221 5822 -1175
rect 5776 -1315 5822 -1269
rect 5776 -1409 5822 -1363
rect 5776 -1503 5822 -1457
rect 5776 -1597 5822 -1551
rect 5776 -1691 5822 -1645
rect 5776 -1785 5822 -1739
rect 8032 -939 8078 -893
rect 10758 -845 10804 -799
rect 8032 -1033 8078 -987
rect 8032 -1127 8078 -1081
rect 8032 -1221 8078 -1175
rect 8032 -1315 8078 -1269
rect 8032 -1409 8078 -1363
rect 8032 -1503 8078 -1457
rect 8032 -1597 8078 -1551
rect 8032 -1691 8078 -1645
rect 8032 -1785 8078 -1739
rect 10758 -939 10804 -893
rect 10758 -1033 10804 -987
rect 10758 -1127 10804 -1081
rect 10758 -1221 10804 -1175
rect 10758 -1315 10804 -1269
rect 10758 -1409 10804 -1363
rect 10758 -1503 10804 -1457
rect 10758 -1597 10804 -1551
rect 10758 -1691 10804 -1645
rect 10758 -1785 10804 -1739
rect 5776 -1879 5822 -1833
rect 5870 -1879 5916 -1833
rect 5964 -1879 6010 -1833
rect 6058 -1879 6104 -1833
rect 6152 -1879 6198 -1833
rect 6246 -1879 6292 -1833
rect 6340 -1879 6386 -1833
rect 6434 -1879 6480 -1833
rect 6528 -1879 6574 -1833
rect 6622 -1879 6668 -1833
rect 6716 -1879 6762 -1833
rect 6810 -1879 6856 -1833
rect 6904 -1879 6950 -1833
rect 6998 -1879 7044 -1833
rect 7092 -1879 7138 -1833
rect 7186 -1879 7232 -1833
rect 7280 -1879 7326 -1833
rect 7374 -1879 7420 -1833
rect 7468 -1879 7514 -1833
rect 7562 -1879 7608 -1833
rect 7656 -1879 7702 -1833
rect 7750 -1879 7796 -1833
rect 7844 -1879 7890 -1833
rect 7938 -1879 7984 -1833
rect 8032 -1879 8078 -1833
rect 8126 -1879 8172 -1833
rect 8220 -1879 8266 -1833
rect 8314 -1879 8360 -1833
rect 8408 -1879 8454 -1833
rect 8502 -1879 8548 -1833
rect 8596 -1879 8642 -1833
rect 8690 -1879 8736 -1833
rect 8784 -1879 8830 -1833
rect 8878 -1879 8924 -1833
rect 8972 -1879 9018 -1833
rect 9066 -1879 9112 -1833
rect 9160 -1879 9206 -1833
rect 9254 -1879 9300 -1833
rect 9348 -1879 9394 -1833
rect 9442 -1879 9488 -1833
rect 9536 -1879 9582 -1833
rect 9630 -1879 9676 -1833
rect 9724 -1879 9770 -1833
rect 9818 -1879 9864 -1833
rect 9912 -1879 9958 -1833
rect 10006 -1879 10052 -1833
rect 10100 -1879 10146 -1833
rect 10194 -1879 10240 -1833
rect 10288 -1879 10334 -1833
rect 10382 -1879 10428 -1833
rect 10476 -1879 10522 -1833
rect 10570 -1879 10616 -1833
rect 10664 -1879 10710 -1833
rect 10758 -1879 10804 -1833
rect 17650 2591 17696 2637
rect 17650 2497 17696 2543
rect 17650 2403 17696 2449
rect 17650 2309 17696 2355
rect 17650 2215 17696 2261
rect 17650 2121 17696 2167
rect 17650 2027 17696 2073
rect 17650 1933 17696 1979
rect 17650 1839 17696 1885
rect 17650 1745 17696 1791
rect 17650 1651 17696 1697
rect 17650 1557 17696 1603
rect 17650 1463 17696 1509
rect 17650 1369 17696 1415
rect 17650 1275 17696 1321
rect 17650 1181 17696 1227
rect 17650 1087 17696 1133
rect 17650 993 17696 1039
rect 17650 899 17696 945
rect 17650 805 17696 851
rect 17650 711 17696 757
rect 17650 617 17696 663
rect 17650 523 17696 569
rect 17650 429 17696 475
rect 17650 335 17696 381
rect 17650 241 17696 287
rect 17650 147 17696 193
rect 17650 53 17696 99
rect 17650 -41 17696 5
rect 17650 -135 17696 -89
rect 17650 -229 17696 -183
rect 17650 -323 17696 -277
rect 17650 -417 17696 -371
rect 20658 3249 20704 3295
rect 17650 -511 17696 -465
rect 20658 3155 20704 3201
rect 20658 3061 20704 3107
rect 20658 2967 20704 3013
rect 20658 2873 20704 2919
rect 20658 2779 20704 2825
rect 20658 2685 20704 2731
rect 20658 2591 20704 2637
rect 20658 2497 20704 2543
rect 20658 2403 20704 2449
rect 20658 2309 20704 2355
rect 20658 2215 20704 2261
rect 20658 2121 20704 2167
rect 20658 2027 20704 2073
rect 20658 1933 20704 1979
rect 20658 1839 20704 1885
rect 20658 1745 20704 1791
rect 20658 1651 20704 1697
rect 20658 1557 20704 1603
rect 20658 1463 20704 1509
rect 20658 1369 20704 1415
rect 20658 1275 20704 1321
rect 20658 1181 20704 1227
rect 20658 1087 20704 1133
rect 20658 993 20704 1039
rect 20658 899 20704 945
rect 20658 805 20704 851
rect 20658 711 20704 757
rect 20658 617 20704 663
rect 20658 523 20704 569
rect 20658 429 20704 475
rect 20658 335 20704 381
rect 20658 241 20704 287
rect 20658 147 20704 193
rect 20658 53 20704 99
rect 20658 -41 20704 5
rect 20658 -135 20704 -89
rect 20658 -229 20704 -183
rect 20658 -323 20704 -277
rect 20658 -417 20704 -371
rect 17650 -605 17696 -559
rect 20658 -511 20704 -465
rect 20658 -605 20704 -559
rect 17650 -699 17696 -653
rect 17650 -793 17696 -747
rect 17650 -887 17696 -841
rect 17650 -981 17696 -935
rect 17650 -1075 17696 -1029
rect 17650 -1169 17696 -1123
rect 17650 -1263 17696 -1217
rect 20658 -699 20704 -653
rect 20658 -793 20704 -747
rect 20658 -887 20704 -841
rect 20658 -981 20704 -935
rect 20658 -1075 20704 -1029
rect 20658 -1169 20704 -1123
rect 17650 -1357 17696 -1311
rect 20658 -1263 20704 -1217
rect 20658 -1357 20704 -1311
rect 17650 -1451 17696 -1405
rect 20658 -1451 20704 -1405
rect 17650 -1545 17696 -1499
rect 17650 -1639 17696 -1593
rect 17650 -1733 17696 -1687
rect 20658 -1545 20704 -1499
rect 20658 -1639 20704 -1593
rect 20658 -1733 20704 -1687
rect 17650 -1827 17696 -1781
rect 17744 -1827 17790 -1781
rect 17838 -1827 17884 -1781
rect 17932 -1827 17978 -1781
rect 18026 -1827 18072 -1781
rect 18120 -1827 18166 -1781
rect 18214 -1827 18260 -1781
rect 18308 -1827 18354 -1781
rect 18402 -1827 18448 -1781
rect 18496 -1827 18542 -1781
rect 18590 -1827 18636 -1781
rect 18684 -1827 18730 -1781
rect 18778 -1827 18824 -1781
rect 18872 -1827 18918 -1781
rect 18966 -1827 19012 -1781
rect 19060 -1827 19106 -1781
rect 19154 -1827 19200 -1781
rect 19248 -1827 19294 -1781
rect 19342 -1827 19388 -1781
rect 19436 -1827 19482 -1781
rect 19530 -1827 19576 -1781
rect 19624 -1827 19670 -1781
rect 19718 -1827 19764 -1781
rect 19812 -1827 19858 -1781
rect 19906 -1827 19952 -1781
rect 20000 -1827 20046 -1781
rect 20094 -1827 20140 -1781
rect 20188 -1827 20234 -1781
rect 20282 -1827 20328 -1781
rect 20376 -1827 20422 -1781
rect 20470 -1827 20516 -1781
rect 20564 -1827 20610 -1781
rect 20658 -1827 20704 -1781
rect 22802 4565 22848 4611
rect 22896 4565 22942 4611
rect 22990 4565 23036 4611
rect 23084 4565 23130 4611
rect 23178 4565 23224 4611
rect 23272 4565 23318 4611
rect 23366 4565 23412 4611
rect 23460 4565 23506 4611
rect 23554 4565 23600 4611
rect 23648 4565 23694 4611
rect 23742 4565 23788 4611
rect 23836 4565 23882 4611
rect 23930 4565 23976 4611
rect 24024 4565 24070 4611
rect 24118 4565 24164 4611
rect 24212 4565 24258 4611
rect 24306 4565 24352 4611
rect 24400 4565 24446 4611
rect 24494 4565 24540 4611
rect 24588 4565 24634 4611
rect 24682 4565 24728 4611
rect 24776 4565 24822 4611
rect 24870 4565 24916 4611
rect 24964 4565 25010 4611
rect 25058 4565 25104 4611
rect 25152 4565 25198 4611
rect 25246 4565 25292 4611
rect 25340 4565 25386 4611
rect 25434 4565 25480 4611
rect 25528 4565 25574 4611
rect 25622 4565 25668 4611
rect 25716 4565 25762 4611
rect 25810 4565 25856 4611
rect 22802 4471 22848 4517
rect 22802 4377 22848 4423
rect 22802 4283 22848 4329
rect 25810 4471 25856 4517
rect 25810 4377 25856 4423
rect 25810 4283 25856 4329
rect 22802 4189 22848 4235
rect 25810 4189 25856 4235
rect 22802 4095 22848 4141
rect 22802 4001 22848 4047
rect 25810 4095 25856 4141
rect 22802 3907 22848 3953
rect 22802 3813 22848 3859
rect 22802 3719 22848 3765
rect 22802 3625 22848 3671
rect 22802 3531 22848 3577
rect 22802 3437 22848 3483
rect 25810 4001 25856 4047
rect 25810 3907 25856 3953
rect 25810 3813 25856 3859
rect 25810 3719 25856 3765
rect 25810 3625 25856 3671
rect 25810 3531 25856 3577
rect 25810 3437 25856 3483
rect 22802 3343 22848 3389
rect 22802 3249 22848 3295
rect 25810 3343 25856 3389
rect 22802 3155 22848 3201
rect 22802 3061 22848 3107
rect 22802 2967 22848 3013
rect 22802 2873 22848 2919
rect 22802 2779 22848 2825
rect 22802 2685 22848 2731
rect 22802 2591 22848 2637
rect 22802 2497 22848 2543
rect 22802 2403 22848 2449
rect 22802 2309 22848 2355
rect 22802 2215 22848 2261
rect 22802 2121 22848 2167
rect 22802 2027 22848 2073
rect 22802 1933 22848 1979
rect 22802 1839 22848 1885
rect 22802 1745 22848 1791
rect 22802 1651 22848 1697
rect 22802 1557 22848 1603
rect 22802 1463 22848 1509
rect 22802 1369 22848 1415
rect 22802 1275 22848 1321
rect 22802 1181 22848 1227
rect 22802 1087 22848 1133
rect 22802 993 22848 1039
rect 22802 899 22848 945
rect 22802 805 22848 851
rect 22802 711 22848 757
rect 22802 617 22848 663
rect 22802 523 22848 569
rect 22802 429 22848 475
rect 22802 335 22848 381
rect 22802 241 22848 287
rect 22802 147 22848 193
rect 22802 53 22848 99
rect 22802 -41 22848 5
rect 22802 -135 22848 -89
rect 22802 -229 22848 -183
rect 22802 -323 22848 -277
rect 22802 -417 22848 -371
rect 25810 3249 25856 3295
rect 22802 -511 22848 -465
rect 25810 3155 25856 3201
rect 25810 3061 25856 3107
rect 25810 2967 25856 3013
rect 25810 2873 25856 2919
rect 25810 2779 25856 2825
rect 25810 2685 25856 2731
rect 25810 2591 25856 2637
rect 25810 2497 25856 2543
rect 25810 2403 25856 2449
rect 25810 2309 25856 2355
rect 25810 2215 25856 2261
rect 25810 2121 25856 2167
rect 25810 2027 25856 2073
rect 25810 1933 25856 1979
rect 25810 1839 25856 1885
rect 25810 1745 25856 1791
rect 25810 1651 25856 1697
rect 25810 1557 25856 1603
rect 25810 1463 25856 1509
rect 25810 1369 25856 1415
rect 25810 1275 25856 1321
rect 25810 1181 25856 1227
rect 25810 1087 25856 1133
rect 25810 993 25856 1039
rect 25810 899 25856 945
rect 25810 805 25856 851
rect 25810 711 25856 757
rect 25810 617 25856 663
rect 25810 523 25856 569
rect 25810 429 25856 475
rect 25810 335 25856 381
rect 25810 241 25856 287
rect 25810 147 25856 193
rect 25810 53 25856 99
rect 25810 -41 25856 5
rect 25810 -135 25856 -89
rect 25810 -229 25856 -183
rect 25810 -323 25856 -277
rect 25810 -417 25856 -371
rect 22802 -605 22848 -559
rect 25810 -511 25856 -465
rect 25810 -605 25856 -559
rect 22802 -699 22848 -653
rect 22802 -793 22848 -747
rect 22802 -887 22848 -841
rect 22802 -981 22848 -935
rect 22802 -1075 22848 -1029
rect 22802 -1169 22848 -1123
rect 22802 -1263 22848 -1217
rect 25810 -699 25856 -653
rect 25810 -793 25856 -747
rect 25810 -887 25856 -841
rect 25810 -981 25856 -935
rect 25810 -1075 25856 -1029
rect 25810 -1169 25856 -1123
rect 22802 -1357 22848 -1311
rect 25810 -1263 25856 -1217
rect 25810 -1357 25856 -1311
rect 22802 -1451 22848 -1405
rect 25810 -1451 25856 -1405
rect 22802 -1545 22848 -1499
rect 22802 -1639 22848 -1593
rect 22802 -1733 22848 -1687
rect 25810 -1545 25856 -1499
rect 25810 -1639 25856 -1593
rect 25810 -1733 25856 -1687
rect 22802 -1827 22848 -1781
rect 22896 -1827 22942 -1781
rect 22990 -1827 23036 -1781
rect 23084 -1827 23130 -1781
rect 23178 -1827 23224 -1781
rect 23272 -1827 23318 -1781
rect 23366 -1827 23412 -1781
rect 23460 -1827 23506 -1781
rect 23554 -1827 23600 -1781
rect 23648 -1827 23694 -1781
rect 23742 -1827 23788 -1781
rect 23836 -1827 23882 -1781
rect 23930 -1827 23976 -1781
rect 24024 -1827 24070 -1781
rect 24118 -1827 24164 -1781
rect 24212 -1827 24258 -1781
rect 24306 -1827 24352 -1781
rect 24400 -1827 24446 -1781
rect 24494 -1827 24540 -1781
rect 24588 -1827 24634 -1781
rect 24682 -1827 24728 -1781
rect 24776 -1827 24822 -1781
rect 24870 -1827 24916 -1781
rect 24964 -1827 25010 -1781
rect 25058 -1827 25104 -1781
rect 25152 -1827 25198 -1781
rect 25246 -1827 25292 -1781
rect 25340 -1827 25386 -1781
rect 25434 -1827 25480 -1781
rect 25528 -1827 25574 -1781
rect 25622 -1827 25668 -1781
rect 25716 -1827 25762 -1781
rect 25810 -1827 25856 -1781
rect 26771 4565 26817 4611
rect 26865 4565 26911 4611
rect 26959 4565 27005 4611
rect 27053 4565 27099 4611
rect 27147 4565 27193 4611
rect 27241 4565 27287 4611
rect 27335 4565 27381 4611
rect 27429 4565 27475 4611
rect 27523 4565 27569 4611
rect 27617 4565 27663 4611
rect 27711 4565 27757 4611
rect 27805 4565 27851 4611
rect 27899 4565 27945 4611
rect 27993 4565 28039 4611
rect 28087 4565 28133 4611
rect 28181 4565 28227 4611
rect 28275 4565 28321 4611
rect 28369 4565 28415 4611
rect 28463 4565 28509 4611
rect 28557 4565 28603 4611
rect 28651 4565 28697 4611
rect 28745 4565 28791 4611
rect 28839 4565 28885 4611
rect 28933 4565 28979 4611
rect 29027 4565 29073 4611
rect 29121 4565 29167 4611
rect 29215 4565 29261 4611
rect 29309 4565 29355 4611
rect 29403 4565 29449 4611
rect 29497 4565 29543 4611
rect 29591 4565 29637 4611
rect 29685 4565 29731 4611
rect 29779 4565 29825 4611
rect 26771 4471 26817 4517
rect 26771 4377 26817 4423
rect 26771 4283 26817 4329
rect 29779 4471 29825 4517
rect 29779 4377 29825 4423
rect 29779 4283 29825 4329
rect 26771 4189 26817 4235
rect 29779 4189 29825 4235
rect 26771 4095 26817 4141
rect 26771 4001 26817 4047
rect 29779 4095 29825 4141
rect 26771 3907 26817 3953
rect 26771 3813 26817 3859
rect 26771 3719 26817 3765
rect 26771 3625 26817 3671
rect 26771 3531 26817 3577
rect 26771 3437 26817 3483
rect 29779 4001 29825 4047
rect 29779 3907 29825 3953
rect 29779 3813 29825 3859
rect 29779 3719 29825 3765
rect 29779 3625 29825 3671
rect 29779 3531 29825 3577
rect 29779 3437 29825 3483
rect 26771 3343 26817 3389
rect 26771 3249 26817 3295
rect 29779 3343 29825 3389
rect 26771 3155 26817 3201
rect 26771 3061 26817 3107
rect 26771 2967 26817 3013
rect 26771 2873 26817 2919
rect 26771 2779 26817 2825
rect 26771 2685 26817 2731
rect 26771 2591 26817 2637
rect 26771 2497 26817 2543
rect 26771 2403 26817 2449
rect 26771 2309 26817 2355
rect 26771 2215 26817 2261
rect 26771 2121 26817 2167
rect 26771 2027 26817 2073
rect 26771 1933 26817 1979
rect 26771 1839 26817 1885
rect 26771 1745 26817 1791
rect 26771 1651 26817 1697
rect 26771 1557 26817 1603
rect 26771 1463 26817 1509
rect 26771 1369 26817 1415
rect 26771 1275 26817 1321
rect 26771 1181 26817 1227
rect 26771 1087 26817 1133
rect 26771 993 26817 1039
rect 26771 899 26817 945
rect 26771 805 26817 851
rect 26771 711 26817 757
rect 26771 617 26817 663
rect 26771 523 26817 569
rect 26771 429 26817 475
rect 26771 335 26817 381
rect 26771 241 26817 287
rect 26771 147 26817 193
rect 26771 53 26817 99
rect 26771 -41 26817 5
rect 26771 -135 26817 -89
rect 26771 -229 26817 -183
rect 26771 -323 26817 -277
rect 26771 -417 26817 -371
rect 29779 3249 29825 3295
rect 26771 -511 26817 -465
rect 29779 3155 29825 3201
rect 29779 3061 29825 3107
rect 29779 2967 29825 3013
rect 29779 2873 29825 2919
rect 29779 2779 29825 2825
rect 29779 2685 29825 2731
rect 29779 2591 29825 2637
rect 29779 2497 29825 2543
rect 29779 2403 29825 2449
rect 29779 2309 29825 2355
rect 29779 2215 29825 2261
rect 29779 2121 29825 2167
rect 29779 2027 29825 2073
rect 29779 1933 29825 1979
rect 29779 1839 29825 1885
rect 29779 1745 29825 1791
rect 29779 1651 29825 1697
rect 29779 1557 29825 1603
rect 29779 1463 29825 1509
rect 29779 1369 29825 1415
rect 29779 1275 29825 1321
rect 29779 1181 29825 1227
rect 29779 1087 29825 1133
rect 29779 993 29825 1039
rect 29779 899 29825 945
rect 29779 805 29825 851
rect 29779 711 29825 757
rect 29779 617 29825 663
rect 29779 523 29825 569
rect 29779 429 29825 475
rect 29779 335 29825 381
rect 29779 241 29825 287
rect 29779 147 29825 193
rect 29779 53 29825 99
rect 29779 -41 29825 5
rect 29779 -135 29825 -89
rect 29779 -229 29825 -183
rect 29779 -323 29825 -277
rect 29779 -417 29825 -371
rect 26771 -605 26817 -559
rect 29779 -511 29825 -465
rect 29779 -605 29825 -559
rect 26771 -699 26817 -653
rect 26771 -793 26817 -747
rect 26771 -887 26817 -841
rect 26771 -981 26817 -935
rect 26771 -1075 26817 -1029
rect 26771 -1169 26817 -1123
rect 26771 -1263 26817 -1217
rect 29779 -699 29825 -653
rect 29779 -793 29825 -747
rect 29779 -887 29825 -841
rect 29779 -981 29825 -935
rect 29779 -1075 29825 -1029
rect 29779 -1169 29825 -1123
rect 26771 -1357 26817 -1311
rect 29779 -1263 29825 -1217
rect 29779 -1357 29825 -1311
rect 26771 -1451 26817 -1405
rect 29779 -1451 29825 -1405
rect 26771 -1545 26817 -1499
rect 26771 -1639 26817 -1593
rect 26771 -1733 26817 -1687
rect 29779 -1545 29825 -1499
rect 29779 -1639 29825 -1593
rect 29779 -1733 29825 -1687
rect 26771 -1827 26817 -1781
rect 26865 -1827 26911 -1781
rect 26959 -1827 27005 -1781
rect 27053 -1827 27099 -1781
rect 27147 -1827 27193 -1781
rect 27241 -1827 27287 -1781
rect 27335 -1827 27381 -1781
rect 27429 -1827 27475 -1781
rect 27523 -1827 27569 -1781
rect 27617 -1827 27663 -1781
rect 27711 -1827 27757 -1781
rect 27805 -1827 27851 -1781
rect 27899 -1827 27945 -1781
rect 27993 -1827 28039 -1781
rect 28087 -1827 28133 -1781
rect 28181 -1827 28227 -1781
rect 28275 -1827 28321 -1781
rect 28369 -1827 28415 -1781
rect 28463 -1827 28509 -1781
rect 28557 -1827 28603 -1781
rect 28651 -1827 28697 -1781
rect 28745 -1827 28791 -1781
rect 28839 -1827 28885 -1781
rect 28933 -1827 28979 -1781
rect 29027 -1827 29073 -1781
rect 29121 -1827 29167 -1781
rect 29215 -1827 29261 -1781
rect 29309 -1827 29355 -1781
rect 29403 -1827 29449 -1781
rect 29497 -1827 29543 -1781
rect 29591 -1827 29637 -1781
rect 29685 -1827 29731 -1781
rect 29779 -1827 29825 -1781
rect 6448 -3085 6494 -3039
rect 6542 -3085 6588 -3039
rect 6636 -3085 6682 -3039
rect 6730 -3085 6776 -3039
rect 6824 -3085 6870 -3039
rect 6918 -3085 6964 -3039
rect 7012 -3085 7058 -3039
rect 7106 -3085 7152 -3039
rect 7200 -3085 7246 -3039
rect 7294 -3085 7340 -3039
rect 7388 -3085 7434 -3039
rect 7482 -3085 7528 -3039
rect 7576 -3085 7622 -3039
rect 7670 -3085 7716 -3039
rect 7764 -3085 7810 -3039
rect 7858 -3085 7904 -3039
rect 7952 -3085 7998 -3039
rect 8046 -3085 8092 -3039
rect 8140 -3085 8186 -3039
rect 8234 -3085 8280 -3039
rect 8328 -3085 8374 -3039
rect 8422 -3085 8468 -3039
rect 8516 -3085 8562 -3039
rect 8610 -3085 8656 -3039
rect 8704 -3085 8750 -3039
rect 8798 -3085 8844 -3039
rect 8892 -3085 8938 -3039
rect 8986 -3085 9032 -3039
rect 9080 -3085 9126 -3039
rect 9174 -3085 9220 -3039
rect 9268 -3085 9314 -3039
rect 9362 -3085 9408 -3039
rect 9456 -3085 9502 -3039
rect 9550 -3085 9596 -3039
rect 6448 -3179 6494 -3133
rect 9550 -3179 9596 -3133
rect 6448 -3273 6494 -3227
rect 6448 -3367 6494 -3321
rect 6448 -3461 6494 -3415
rect 9550 -3273 9596 -3227
rect 9550 -3367 9596 -3321
rect 6448 -3555 6494 -3509
rect 6448 -3649 6494 -3603
rect 9550 -3461 9596 -3415
rect 9550 -3555 9596 -3509
rect 6448 -3743 6494 -3697
rect 6448 -3837 6494 -3791
rect 6448 -3931 6494 -3885
rect 6448 -4025 6494 -3979
rect 6448 -4119 6494 -4073
rect 6448 -4213 6494 -4167
rect 6448 -4307 6494 -4261
rect 6448 -4401 6494 -4355
rect 6448 -4495 6494 -4449
rect 6448 -4589 6494 -4543
rect 6448 -4683 6494 -4637
rect 6448 -4777 6494 -4731
rect 6448 -4871 6494 -4825
rect 6448 -4965 6494 -4919
rect 6448 -5059 6494 -5013
rect 6448 -5153 6494 -5107
rect 6448 -5247 6494 -5201
rect 6448 -5341 6494 -5295
rect 6448 -5435 6494 -5389
rect 6448 -5529 6494 -5483
rect 6448 -5623 6494 -5577
rect 6448 -5717 6494 -5671
rect 6448 -5811 6494 -5765
rect 6448 -5905 6494 -5859
rect 6448 -5999 6494 -5953
rect 6448 -6093 6494 -6047
rect 9550 -3649 9596 -3603
rect 9550 -3743 9596 -3697
rect 9550 -3837 9596 -3791
rect 9550 -3931 9596 -3885
rect 9550 -4025 9596 -3979
rect 9550 -4119 9596 -4073
rect 9550 -4213 9596 -4167
rect 9550 -4307 9596 -4261
rect 9550 -4401 9596 -4355
rect 9550 -4495 9596 -4449
rect 9550 -4589 9596 -4543
rect 9550 -4683 9596 -4637
rect 9550 -4777 9596 -4731
rect 9550 -4871 9596 -4825
rect 9550 -4965 9596 -4919
rect 9550 -5059 9596 -5013
rect 9550 -5153 9596 -5107
rect 9550 -5247 9596 -5201
rect 9550 -5341 9596 -5295
rect 9550 -5435 9596 -5389
rect 9550 -5529 9596 -5483
rect 9550 -5623 9596 -5577
rect 9550 -5717 9596 -5671
rect 9550 -5811 9596 -5765
rect 9550 -5905 9596 -5859
rect 9550 -5999 9596 -5953
rect 9550 -6093 9596 -6047
rect 6448 -6187 6494 -6141
rect 6448 -6281 6494 -6235
rect 9550 -6187 9596 -6141
rect 9550 -6281 9596 -6235
rect 5414 -6375 5460 -6329
rect 5508 -6375 5554 -6329
rect 5602 -6375 5648 -6329
rect 5696 -6375 5742 -6329
rect 5790 -6375 5836 -6329
rect 5884 -6375 5930 -6329
rect 5978 -6375 6024 -6329
rect 6072 -6375 6118 -6329
rect 6166 -6375 6212 -6329
rect 6260 -6375 6306 -6329
rect 6354 -6375 6400 -6329
rect 6448 -6375 6494 -6329
rect 11528 -4734 11574 -4688
rect 11622 -4734 11668 -4688
rect 11716 -4734 11762 -4688
rect 11810 -4734 11856 -4688
rect 11904 -4734 11950 -4688
rect 11998 -4734 12044 -4688
rect 12092 -4734 12138 -4688
rect 12186 -4734 12232 -4688
rect 12280 -4734 12326 -4688
rect 12374 -4734 12420 -4688
rect 12468 -4734 12514 -4688
rect 12562 -4734 12608 -4688
rect 12656 -4734 12702 -4688
rect 12750 -4734 12796 -4688
rect 12844 -4734 12890 -4688
rect 12938 -4734 12984 -4688
rect 13032 -4734 13078 -4688
rect 13126 -4734 13172 -4688
rect 13220 -4734 13266 -4688
rect 13314 -4734 13360 -4688
rect 13408 -4734 13454 -4688
rect 13502 -4734 13548 -4688
rect 13596 -4734 13642 -4688
rect 13690 -4734 13736 -4688
rect 13784 -4734 13830 -4688
rect 13878 -4734 13924 -4688
rect 13972 -4734 14018 -4688
rect 14066 -4734 14112 -4688
rect 14160 -4734 14206 -4688
rect 14254 -4734 14300 -4688
rect 14348 -4734 14394 -4688
rect 14442 -4734 14488 -4688
rect 14536 -4734 14582 -4688
rect 14630 -4734 14676 -4688
rect 14724 -4734 14770 -4688
rect 14818 -4734 14864 -4688
rect 14912 -4734 14958 -4688
rect 15006 -4734 15052 -4688
rect 15100 -4734 15146 -4688
rect 15194 -4734 15240 -4688
rect 15288 -4734 15334 -4688
rect 15382 -4734 15428 -4688
rect 15476 -4734 15522 -4688
rect 15570 -4734 15616 -4688
rect 15664 -4734 15710 -4688
rect 15758 -4734 15804 -4688
rect 15852 -4734 15898 -4688
rect 15946 -4734 15992 -4688
rect 16040 -4734 16086 -4688
rect 16134 -4734 16180 -4688
rect 16228 -4734 16274 -4688
rect 16322 -4734 16368 -4688
rect 16416 -4734 16462 -4688
rect 16510 -4734 16556 -4688
rect 16604 -4734 16650 -4688
rect 16698 -4734 16744 -4688
rect 16792 -4734 16838 -4688
rect 16886 -4734 16932 -4688
rect 16980 -4734 17026 -4688
rect 17074 -4734 17120 -4688
rect 11528 -4828 11574 -4782
rect 11528 -4922 11574 -4876
rect 11528 -5016 11574 -4970
rect 11528 -5110 11574 -5064
rect 17074 -4828 17120 -4782
rect 17074 -4922 17120 -4876
rect 17074 -5016 17120 -4970
rect 11528 -5204 11574 -5158
rect 11528 -5298 11574 -5252
rect 11528 -5392 11574 -5346
rect 17074 -5110 17120 -5064
rect 17074 -5204 17120 -5158
rect 17074 -5298 17120 -5252
rect 11528 -5486 11574 -5440
rect 11528 -5580 11574 -5534
rect 11528 -5674 11574 -5628
rect 11528 -5768 11574 -5722
rect 17074 -5392 17120 -5346
rect 17074 -5486 17120 -5440
rect 17074 -5580 17120 -5534
rect 17074 -5674 17120 -5628
rect 17074 -5768 17120 -5722
rect 11528 -5862 11574 -5816
rect 11528 -5956 11574 -5910
rect 11528 -6050 11574 -6004
rect 11528 -6144 11574 -6098
rect 11528 -6238 11574 -6192
rect 9550 -6375 9596 -6329
rect 9644 -6375 9690 -6329
rect 9738 -6375 9784 -6329
rect 9832 -6375 9878 -6329
rect 9926 -6375 9972 -6329
rect 10020 -6375 10066 -6329
rect 10114 -6375 10160 -6329
rect 10208 -6375 10254 -6329
rect 10302 -6375 10348 -6329
rect 10396 -6375 10442 -6329
rect 10490 -6375 10536 -6329
rect 10584 -6375 10630 -6329
rect 5414 -6469 5460 -6423
rect 10584 -6469 10630 -6423
rect 5414 -6563 5460 -6517
rect 5414 -6657 5460 -6611
rect 5414 -6751 5460 -6705
rect 10584 -6563 10630 -6517
rect 10584 -6657 10630 -6611
rect 5414 -6845 5460 -6799
rect 5414 -6939 5460 -6893
rect 10584 -6751 10630 -6705
rect 10584 -6845 10630 -6799
rect 5414 -7033 5460 -6987
rect 5414 -7127 5460 -7081
rect 10584 -6939 10630 -6893
rect 10584 -7033 10630 -6987
rect 5414 -7221 5460 -7175
rect 10584 -7127 10630 -7081
rect 5414 -7315 5460 -7269
rect 5414 -7409 5460 -7363
rect 10584 -7221 10630 -7175
rect 10584 -7315 10630 -7269
rect 5414 -7503 5460 -7457
rect 5414 -7597 5460 -7551
rect 5414 -7691 5460 -7645
rect 5414 -7785 5460 -7739
rect 10584 -7409 10630 -7363
rect 10584 -7503 10630 -7457
rect 10584 -7597 10630 -7551
rect 10584 -7691 10630 -7645
rect 10584 -7785 10630 -7739
rect 5414 -7879 5460 -7833
rect 5508 -7879 5554 -7833
rect 5602 -7879 5648 -7833
rect 5696 -7879 5742 -7833
rect 5790 -7879 5836 -7833
rect 5884 -7879 5930 -7833
rect 5978 -7879 6024 -7833
rect 6072 -7879 6118 -7833
rect 6166 -7879 6212 -7833
rect 6260 -7879 6306 -7833
rect 6354 -7879 6400 -7833
rect 6448 -7879 6494 -7833
rect 6542 -7879 6588 -7833
rect 6636 -7879 6682 -7833
rect 6730 -7879 6776 -7833
rect 6824 -7879 6870 -7833
rect 6918 -7879 6964 -7833
rect 7012 -7879 7058 -7833
rect 7106 -7879 7152 -7833
rect 7200 -7879 7246 -7833
rect 7294 -7879 7340 -7833
rect 7388 -7879 7434 -7833
rect 7482 -7879 7528 -7833
rect 7576 -7879 7622 -7833
rect 7670 -7879 7716 -7833
rect 7764 -7879 7810 -7833
rect 7858 -7879 7904 -7833
rect 7952 -7879 7998 -7833
rect 8046 -7879 8092 -7833
rect 8140 -7879 8186 -7833
rect 8234 -7879 8280 -7833
rect 8328 -7879 8374 -7833
rect 8422 -7879 8468 -7833
rect 8516 -7879 8562 -7833
rect 8610 -7879 8656 -7833
rect 8704 -7879 8750 -7833
rect 8798 -7879 8844 -7833
rect 8892 -7879 8938 -7833
rect 8986 -7879 9032 -7833
rect 9080 -7879 9126 -7833
rect 9174 -7879 9220 -7833
rect 9268 -7879 9314 -7833
rect 9362 -7879 9408 -7833
rect 9456 -7879 9502 -7833
rect 9550 -7879 9596 -7833
rect 9644 -7879 9690 -7833
rect 9738 -7879 9784 -7833
rect 9832 -7879 9878 -7833
rect 9926 -7879 9972 -7833
rect 10020 -7879 10066 -7833
rect 10114 -7879 10160 -7833
rect 10208 -7879 10254 -7833
rect 10302 -7879 10348 -7833
rect 10396 -7879 10442 -7833
rect 10490 -7879 10536 -7833
rect 10584 -7879 10630 -7833
rect 11528 -6332 11574 -6286
rect 11528 -6426 11574 -6380
rect 11528 -6520 11574 -6474
rect 11528 -6614 11574 -6568
rect 11528 -6708 11574 -6662
rect 17074 -5862 17120 -5816
rect 17074 -5956 17120 -5910
rect 17074 -6050 17120 -6004
rect 17074 -6144 17120 -6098
rect 17074 -6238 17120 -6192
rect 17074 -6332 17120 -6286
rect 17074 -6426 17120 -6380
rect 17074 -6520 17120 -6474
rect 17074 -6614 17120 -6568
rect 17074 -6708 17120 -6662
rect 11528 -6802 11574 -6756
rect 11528 -6896 11574 -6850
rect 11528 -6990 11574 -6944
rect 11528 -7084 11574 -7038
rect 11528 -7178 11574 -7132
rect 17074 -6802 17120 -6756
rect 17074 -6896 17120 -6850
rect 17074 -6990 17120 -6944
rect 17074 -7084 17120 -7038
rect 11528 -7272 11574 -7226
rect 11528 -7366 11574 -7320
rect 11528 -7460 11574 -7414
rect 11528 -7554 11574 -7508
rect 17074 -7178 17120 -7132
rect 17074 -7272 17120 -7226
rect 17074 -7366 17120 -7320
rect 17074 -7460 17120 -7414
rect 11528 -7648 11574 -7602
rect 11528 -7742 11574 -7696
rect 17074 -7554 17120 -7508
rect 17074 -7648 17120 -7602
rect 17074 -7742 17120 -7696
rect 11528 -7836 11574 -7790
rect 11622 -7836 11668 -7790
rect 11716 -7836 11762 -7790
rect 11810 -7836 11856 -7790
rect 11904 -7836 11950 -7790
rect 11998 -7836 12044 -7790
rect 12092 -7836 12138 -7790
rect 12186 -7836 12232 -7790
rect 12280 -7836 12326 -7790
rect 12374 -7836 12420 -7790
rect 12468 -7836 12514 -7790
rect 12562 -7836 12608 -7790
rect 12656 -7836 12702 -7790
rect 12750 -7836 12796 -7790
rect 12844 -7836 12890 -7790
rect 12938 -7836 12984 -7790
rect 13032 -7836 13078 -7790
rect 13126 -7836 13172 -7790
rect 13220 -7836 13266 -7790
rect 13314 -7836 13360 -7790
rect 13408 -7836 13454 -7790
rect 13502 -7836 13548 -7790
rect 13596 -7836 13642 -7790
rect 13690 -7836 13736 -7790
rect 13784 -7836 13830 -7790
rect 13878 -7836 13924 -7790
rect 13972 -7836 14018 -7790
rect 14066 -7836 14112 -7790
rect 14160 -7836 14206 -7790
rect 14254 -7836 14300 -7790
rect 14348 -7836 14394 -7790
rect 14442 -7836 14488 -7790
rect 14536 -7836 14582 -7790
rect 14630 -7836 14676 -7790
rect 14724 -7836 14770 -7790
rect 14818 -7836 14864 -7790
rect 14912 -7836 14958 -7790
rect 15006 -7836 15052 -7790
rect 15100 -7836 15146 -7790
rect 15194 -7836 15240 -7790
rect 15288 -7836 15334 -7790
rect 15382 -7836 15428 -7790
rect 15476 -7836 15522 -7790
rect 15570 -7836 15616 -7790
rect 15664 -7836 15710 -7790
rect 15758 -7836 15804 -7790
rect 15852 -7836 15898 -7790
rect 15946 -7836 15992 -7790
rect 16040 -7836 16086 -7790
rect 16134 -7836 16180 -7790
rect 16228 -7836 16274 -7790
rect 16322 -7836 16368 -7790
rect 16416 -7836 16462 -7790
rect 16510 -7836 16556 -7790
rect 16604 -7836 16650 -7790
rect 16698 -7836 16744 -7790
rect 16792 -7836 16838 -7790
rect 16886 -7836 16932 -7790
rect 16980 -7836 17026 -7790
rect 17074 -7836 17120 -7790
<< nsubdiffcont >>
rect 2958 5171 3004 5217
rect 3052 5171 3098 5217
rect 3146 5171 3192 5217
rect 3240 5171 3286 5217
rect 3334 5171 3380 5217
rect 3428 5171 3474 5217
rect 3522 5171 3568 5217
rect 3616 5171 3662 5217
rect 3710 5171 3756 5217
rect 3804 5171 3850 5217
rect 3898 5171 3944 5217
rect 3992 5171 4038 5217
rect 4086 5171 4132 5217
rect 4180 5171 4226 5217
rect 4274 5171 4320 5217
rect 4368 5171 4414 5217
rect 4462 5171 4508 5217
rect 4556 5171 4602 5217
rect 4650 5171 4696 5217
rect 4744 5171 4790 5217
rect 4838 5171 4884 5217
rect 4932 5171 4978 5217
rect 5026 5171 5072 5217
rect 5120 5171 5166 5217
rect 2958 5077 3004 5123
rect 5120 5077 5166 5123
rect 2958 4983 3004 5029
rect 2958 4889 3004 4935
rect 5120 4983 5166 5029
rect 5120 4889 5166 4935
rect 2958 4795 3004 4841
rect 2958 4701 3004 4747
rect 2958 4607 3004 4653
rect 2958 4513 3004 4559
rect 2958 4419 3004 4465
rect 2958 4325 3004 4371
rect 2958 4231 3004 4277
rect 2958 4137 3004 4183
rect 5120 4795 5166 4841
rect 5120 4701 5166 4747
rect 5120 4607 5166 4653
rect 5120 4513 5166 4559
rect 5120 4419 5166 4465
rect 5120 4325 5166 4371
rect 5120 4231 5166 4277
rect 5120 4137 5166 4183
rect 2958 4043 3004 4089
rect 2958 3949 3004 3995
rect 2958 3855 3004 3901
rect 2958 3761 3004 3807
rect 5120 4043 5166 4089
rect 5120 3949 5166 3995
rect 5120 3855 5166 3901
rect 5120 3761 5166 3807
rect 2958 3667 3004 3713
rect 2958 3573 3004 3619
rect 2958 3479 3004 3525
rect 2958 3385 3004 3431
rect 2958 3291 3004 3337
rect 2958 3197 3004 3243
rect 2958 3103 3004 3149
rect 2958 3009 3004 3055
rect 5120 3667 5166 3713
rect 5120 3573 5166 3619
rect 5120 3479 5166 3525
rect 5120 3385 5166 3431
rect 5120 3291 5166 3337
rect 5120 3197 5166 3243
rect 5120 3103 5166 3149
rect 5120 3009 5166 3055
rect 2958 2915 3004 2961
rect 2958 2821 3004 2867
rect 2958 2727 3004 2773
rect 2958 2633 3004 2679
rect 5120 2915 5166 2961
rect 5120 2821 5166 2867
rect 5120 2727 5166 2773
rect 5120 2633 5166 2679
rect 2958 2539 3004 2585
rect 2958 2445 3004 2491
rect 2958 2351 3004 2397
rect 2958 2257 3004 2303
rect 2958 2163 3004 2209
rect 2958 2069 3004 2115
rect 2958 1975 3004 2021
rect 2958 1881 3004 1927
rect 5120 2539 5166 2585
rect 5120 2445 5166 2491
rect 5120 2351 5166 2397
rect 5120 2257 5166 2303
rect 5120 2163 5166 2209
rect 5120 2069 5166 2115
rect 5120 1975 5166 2021
rect 5120 1881 5166 1927
rect 2958 1787 3004 1833
rect 44 1693 90 1739
rect 138 1693 184 1739
rect 232 1693 278 1739
rect 326 1693 372 1739
rect 420 1693 466 1739
rect 514 1693 560 1739
rect 608 1693 654 1739
rect 702 1693 748 1739
rect 796 1693 842 1739
rect 890 1693 936 1739
rect 984 1693 1030 1739
rect 1078 1693 1124 1739
rect 1172 1693 1218 1739
rect 1266 1693 1312 1739
rect 1360 1693 1406 1739
rect 1454 1693 1500 1739
rect 1548 1693 1594 1739
rect 1642 1693 1688 1739
rect 1736 1693 1782 1739
rect 1830 1693 1876 1739
rect 1924 1693 1970 1739
rect 2018 1693 2064 1739
rect 2112 1693 2158 1739
rect 2206 1693 2252 1739
rect 2300 1693 2346 1739
rect 2394 1693 2440 1739
rect 2488 1693 2534 1739
rect 2582 1693 2628 1739
rect 2676 1693 2722 1739
rect 2770 1693 2816 1739
rect 2864 1693 2910 1739
rect 2958 1693 3004 1739
rect 44 1599 90 1645
rect 44 1505 90 1551
rect 44 1411 90 1457
rect 44 1317 90 1363
rect 44 1223 90 1269
rect 44 1129 90 1175
rect 44 1035 90 1081
rect 44 941 90 987
rect 44 847 90 893
rect 44 753 90 799
rect 2958 1599 3004 1645
rect 2958 1505 3004 1551
rect 5120 1787 5166 1833
rect 5120 1693 5166 1739
rect 5120 1599 5166 1645
rect 5120 1505 5166 1551
rect 2958 1411 3004 1457
rect 2958 1317 3004 1363
rect 2958 1223 3004 1269
rect 2958 1129 3004 1175
rect 2958 1035 3004 1081
rect 2958 941 3004 987
rect 2958 847 3004 893
rect 44 659 90 705
rect 2958 753 3004 799
rect 5120 1411 5166 1457
rect 5120 1317 5166 1363
rect 5120 1223 5166 1269
rect 5120 1129 5166 1175
rect 5120 1035 5166 1081
rect 5120 941 5166 987
rect 5120 847 5166 893
rect 5120 753 5166 799
rect 2958 659 3004 705
rect 44 565 90 611
rect 44 471 90 517
rect 44 377 90 423
rect 44 283 90 329
rect 44 189 90 235
rect 44 95 90 141
rect 44 1 90 47
rect 2958 565 3004 611
rect 2958 471 3004 517
rect 2958 377 3004 423
rect 5120 659 5166 705
rect 5120 565 5166 611
rect 5120 471 5166 517
rect 5120 377 5166 423
rect 2958 283 3004 329
rect 2958 189 3004 235
rect 2958 95 3004 141
rect 44 -93 90 -47
rect 2958 1 3004 47
rect 2958 -93 3004 -47
rect 44 -187 90 -141
rect 44 -281 90 -235
rect 44 -375 90 -329
rect 44 -469 90 -423
rect 44 -563 90 -517
rect 44 -657 90 -611
rect 44 -751 90 -705
rect 2958 -187 3004 -141
rect 2958 -281 3004 -235
rect 2958 -375 3004 -329
rect 5120 283 5166 329
rect 5120 189 5166 235
rect 5120 95 5166 141
rect 5120 1 5166 47
rect 5120 -93 5166 -47
rect 5120 -187 5166 -141
rect 5120 -281 5166 -235
rect 5120 -375 5166 -329
rect 2958 -469 3004 -423
rect 2958 -563 3004 -517
rect 2958 -657 3004 -611
rect 5120 -469 5166 -423
rect 44 -845 90 -799
rect 2958 -751 3004 -705
rect 5120 -563 5166 -517
rect 5120 -657 5166 -611
rect 5120 -751 5166 -705
rect 2958 -845 3004 -799
rect 44 -939 90 -893
rect 44 -1033 90 -987
rect 44 -1127 90 -1081
rect 44 -1221 90 -1175
rect 44 -1315 90 -1269
rect 44 -1409 90 -1363
rect 44 -1503 90 -1457
rect 2958 -939 3004 -893
rect 2958 -1033 3004 -987
rect 2958 -1127 3004 -1081
rect 2958 -1221 3004 -1175
rect 2958 -1315 3004 -1269
rect 2958 -1409 3004 -1363
rect 2958 -1503 3004 -1457
rect 44 -1597 90 -1551
rect 5120 -845 5166 -799
rect 5120 -939 5166 -893
rect 5120 -1033 5166 -987
rect 5120 -1127 5166 -1081
rect 5120 -1221 5166 -1175
rect 5120 -1315 5166 -1269
rect 5120 -1409 5166 -1363
rect 5120 -1503 5166 -1457
rect 2958 -1597 3004 -1551
rect 44 -1691 90 -1645
rect 44 -1785 90 -1739
rect 2958 -1691 3004 -1645
rect 5120 -1597 5166 -1551
rect 5120 -1691 5166 -1645
rect 2958 -1785 3004 -1739
rect 5120 -1785 5166 -1739
rect 44 -1879 90 -1833
rect 138 -1879 184 -1833
rect 232 -1879 278 -1833
rect 326 -1879 372 -1833
rect 420 -1879 466 -1833
rect 514 -1879 560 -1833
rect 608 -1879 654 -1833
rect 702 -1879 748 -1833
rect 796 -1879 842 -1833
rect 890 -1879 936 -1833
rect 984 -1879 1030 -1833
rect 1078 -1879 1124 -1833
rect 1172 -1879 1218 -1833
rect 1266 -1879 1312 -1833
rect 1360 -1879 1406 -1833
rect 1454 -1879 1500 -1833
rect 1548 -1879 1594 -1833
rect 1642 -1879 1688 -1833
rect 1736 -1879 1782 -1833
rect 1830 -1879 1876 -1833
rect 1924 -1879 1970 -1833
rect 2018 -1879 2064 -1833
rect 2112 -1879 2158 -1833
rect 2206 -1879 2252 -1833
rect 2300 -1879 2346 -1833
rect 2394 -1879 2440 -1833
rect 2488 -1879 2534 -1833
rect 2582 -1879 2628 -1833
rect 2676 -1879 2722 -1833
rect 2770 -1879 2816 -1833
rect 2864 -1879 2910 -1833
rect 2958 -1879 3004 -1833
rect 3052 -1879 3098 -1833
rect 3146 -1879 3192 -1833
rect 3240 -1879 3286 -1833
rect 3334 -1879 3380 -1833
rect 3428 -1879 3474 -1833
rect 3522 -1879 3568 -1833
rect 3616 -1879 3662 -1833
rect 3710 -1879 3756 -1833
rect 3804 -1879 3850 -1833
rect 3898 -1879 3944 -1833
rect 3992 -1879 4038 -1833
rect 4086 -1879 4132 -1833
rect 4180 -1879 4226 -1833
rect 4274 -1879 4320 -1833
rect 4368 -1879 4414 -1833
rect 4462 -1879 4508 -1833
rect 4556 -1879 4602 -1833
rect 4650 -1879 4696 -1833
rect 4744 -1879 4790 -1833
rect 4838 -1879 4884 -1833
rect 4932 -1879 4978 -1833
rect 5026 -1879 5072 -1833
rect 5120 -1879 5166 -1833
rect 11414 2539 11460 2585
rect 11508 2539 11554 2585
rect 11602 2539 11648 2585
rect 11696 2539 11742 2585
rect 11790 2539 11836 2585
rect 11884 2539 11930 2585
rect 11978 2539 12024 2585
rect 12072 2539 12118 2585
rect 12166 2539 12212 2585
rect 12260 2539 12306 2585
rect 12354 2539 12400 2585
rect 12448 2539 12494 2585
rect 12542 2539 12588 2585
rect 12636 2539 12682 2585
rect 12730 2539 12776 2585
rect 12824 2539 12870 2585
rect 12918 2539 12964 2585
rect 13012 2539 13058 2585
rect 13106 2539 13152 2585
rect 13200 2539 13246 2585
rect 13294 2539 13340 2585
rect 13388 2539 13434 2585
rect 13482 2539 13528 2585
rect 13576 2539 13622 2585
rect 13670 2539 13716 2585
rect 13764 2539 13810 2585
rect 13858 2539 13904 2585
rect 13952 2539 13998 2585
rect 14046 2539 14092 2585
rect 14140 2539 14186 2585
rect 14234 2539 14280 2585
rect 14328 2539 14374 2585
rect 14422 2539 14468 2585
rect 14516 2539 14562 2585
rect 14610 2539 14656 2585
rect 14704 2539 14750 2585
rect 14798 2539 14844 2585
rect 14892 2539 14938 2585
rect 14986 2539 15032 2585
rect 15080 2539 15126 2585
rect 15174 2539 15220 2585
rect 15268 2539 15314 2585
rect 15362 2539 15408 2585
rect 15456 2539 15502 2585
rect 15550 2539 15596 2585
rect 15644 2539 15690 2585
rect 15738 2539 15784 2585
rect 15832 2539 15878 2585
rect 15926 2539 15972 2585
rect 16020 2539 16066 2585
rect 16114 2539 16160 2585
rect 16208 2539 16254 2585
rect 16302 2539 16348 2585
rect 16396 2539 16442 2585
rect 16490 2539 16536 2585
rect 11414 2445 11460 2491
rect 11414 2351 11460 2397
rect 11414 2257 11460 2303
rect 11414 2163 11460 2209
rect 11414 2069 11460 2115
rect 11414 1975 11460 2021
rect 11414 1881 11460 1927
rect 11414 1787 11460 1833
rect 11414 1693 11460 1739
rect 11414 1599 11460 1645
rect 14140 2445 14186 2491
rect 14140 2351 14186 2397
rect 14140 2257 14186 2303
rect 14140 2163 14186 2209
rect 14140 2069 14186 2115
rect 14140 1975 14186 2021
rect 14140 1881 14186 1927
rect 14140 1787 14186 1833
rect 14140 1693 14186 1739
rect 14140 1599 14186 1645
rect 11414 1505 11460 1551
rect 11414 1411 11460 1457
rect 11414 1317 11460 1363
rect 11414 1223 11460 1269
rect 16490 2445 16536 2491
rect 16490 2351 16536 2397
rect 16490 2257 16536 2303
rect 16490 2163 16536 2209
rect 16490 2069 16536 2115
rect 16490 1975 16536 2021
rect 16490 1881 16536 1927
rect 16490 1787 16536 1833
rect 16490 1693 16536 1739
rect 16490 1599 16536 1645
rect 14140 1505 14186 1551
rect 14140 1411 14186 1457
rect 14140 1317 14186 1363
rect 14140 1223 14186 1269
rect 11414 1129 11460 1175
rect 11414 1035 11460 1081
rect 11414 941 11460 987
rect 11414 847 11460 893
rect 11414 753 11460 799
rect 11414 659 11460 705
rect 11414 565 11460 611
rect 16490 1505 16536 1551
rect 16490 1411 16536 1457
rect 16490 1317 16536 1363
rect 16490 1223 16536 1269
rect 14140 1129 14186 1175
rect 14140 1035 14186 1081
rect 14140 941 14186 987
rect 14140 847 14186 893
rect 14140 753 14186 799
rect 14140 659 14186 705
rect 14140 565 14186 611
rect 11414 471 11460 517
rect 11414 377 11460 423
rect 11414 283 11460 329
rect 11414 189 11460 235
rect 16490 1129 16536 1175
rect 16490 1035 16536 1081
rect 16490 941 16536 987
rect 16490 847 16536 893
rect 16490 753 16536 799
rect 16490 659 16536 705
rect 16490 565 16536 611
rect 14140 471 14186 517
rect 14140 377 14186 423
rect 14140 283 14186 329
rect 14140 189 14186 235
rect 11414 95 11460 141
rect 11414 1 11460 47
rect 11414 -93 11460 -47
rect 11414 -187 11460 -141
rect 11414 -281 11460 -235
rect 11414 -375 11460 -329
rect 11414 -469 11460 -423
rect 16490 471 16536 517
rect 16490 377 16536 423
rect 16490 283 16536 329
rect 16490 189 16536 235
rect 14140 95 14186 141
rect 14140 1 14186 47
rect 14140 -93 14186 -47
rect 14140 -187 14186 -141
rect 14140 -281 14186 -235
rect 14140 -375 14186 -329
rect 14140 -469 14186 -423
rect 11414 -563 11460 -517
rect 11414 -657 11460 -611
rect 11414 -751 11460 -705
rect 16490 95 16536 141
rect 16490 1 16536 47
rect 16490 -93 16536 -47
rect 16490 -187 16536 -141
rect 16490 -281 16536 -235
rect 16490 -375 16536 -329
rect 16490 -469 16536 -423
rect 14140 -563 14186 -517
rect 14140 -657 14186 -611
rect 11414 -845 11460 -799
rect 14140 -751 14186 -705
rect 16490 -563 16536 -517
rect 16490 -657 16536 -611
rect 14140 -845 14186 -799
rect 11414 -939 11460 -893
rect 11414 -1033 11460 -987
rect 11414 -1127 11460 -1081
rect 11414 -1221 11460 -1175
rect 11414 -1315 11460 -1269
rect 11414 -1409 11460 -1363
rect 11414 -1503 11460 -1457
rect 11414 -1597 11460 -1551
rect 11414 -1691 11460 -1645
rect 11414 -1785 11460 -1739
rect 16490 -751 16536 -705
rect 16490 -845 16536 -799
rect 14140 -939 14186 -893
rect 14140 -1033 14186 -987
rect 14140 -1127 14186 -1081
rect 14140 -1221 14186 -1175
rect 14140 -1315 14186 -1269
rect 14140 -1409 14186 -1363
rect 14140 -1503 14186 -1457
rect 14140 -1597 14186 -1551
rect 14140 -1691 14186 -1645
rect 14140 -1785 14186 -1739
rect 16490 -939 16536 -893
rect 16490 -1033 16536 -987
rect 16490 -1127 16536 -1081
rect 16490 -1221 16536 -1175
rect 16490 -1315 16536 -1269
rect 16490 -1409 16536 -1363
rect 16490 -1503 16536 -1457
rect 16490 -1597 16536 -1551
rect 16490 -1691 16536 -1645
rect 16490 -1785 16536 -1739
rect 11414 -1879 11460 -1833
rect 11508 -1879 11554 -1833
rect 11602 -1879 11648 -1833
rect 11696 -1879 11742 -1833
rect 11790 -1879 11836 -1833
rect 11884 -1879 11930 -1833
rect 11978 -1879 12024 -1833
rect 12072 -1879 12118 -1833
rect 12166 -1879 12212 -1833
rect 12260 -1879 12306 -1833
rect 12354 -1879 12400 -1833
rect 12448 -1879 12494 -1833
rect 12542 -1879 12588 -1833
rect 12636 -1879 12682 -1833
rect 12730 -1879 12776 -1833
rect 12824 -1879 12870 -1833
rect 12918 -1879 12964 -1833
rect 13012 -1879 13058 -1833
rect 13106 -1879 13152 -1833
rect 13200 -1879 13246 -1833
rect 13294 -1879 13340 -1833
rect 13388 -1879 13434 -1833
rect 13482 -1879 13528 -1833
rect 13576 -1879 13622 -1833
rect 13670 -1879 13716 -1833
rect 13764 -1879 13810 -1833
rect 13858 -1879 13904 -1833
rect 13952 -1879 13998 -1833
rect 14046 -1879 14092 -1833
rect 14140 -1879 14186 -1833
rect 14234 -1879 14280 -1833
rect 14328 -1879 14374 -1833
rect 14422 -1879 14468 -1833
rect 14516 -1879 14562 -1833
rect 14610 -1879 14656 -1833
rect 14704 -1879 14750 -1833
rect 14798 -1879 14844 -1833
rect 14892 -1879 14938 -1833
rect 14986 -1879 15032 -1833
rect 15080 -1879 15126 -1833
rect 15174 -1879 15220 -1833
rect 15268 -1879 15314 -1833
rect 15362 -1879 15408 -1833
rect 15456 -1879 15502 -1833
rect 15550 -1879 15596 -1833
rect 15644 -1879 15690 -1833
rect 15738 -1879 15784 -1833
rect 15832 -1879 15878 -1833
rect 15926 -1879 15972 -1833
rect 16020 -1879 16066 -1833
rect 16114 -1879 16160 -1833
rect 16208 -1879 16254 -1833
rect 16302 -1879 16348 -1833
rect 16396 -1879 16442 -1833
rect 16490 -1879 16536 -1833
rect 32143 3016 32189 3062
rect 32237 3016 32283 3062
rect 32331 3016 32377 3062
rect 32425 3016 32471 3062
rect 32519 3016 32565 3062
rect 32613 3016 32659 3062
rect 32707 3016 32753 3062
rect 32801 3016 32847 3062
rect 32895 3016 32941 3062
rect 32989 3016 33035 3062
rect 33083 3016 33129 3062
rect 33177 3016 33223 3062
rect 33271 3016 33317 3062
rect 33365 3016 33411 3062
rect 33459 3016 33505 3062
rect 33553 3016 33599 3062
rect 33647 3016 33693 3062
rect 33741 3016 33787 3062
rect 33835 3016 33881 3062
rect 33929 3016 33975 3062
rect 34023 3016 34069 3062
rect 34117 3016 34163 3062
rect 34211 3016 34257 3062
rect 34305 3016 34351 3062
rect 34399 3016 34445 3062
rect 34493 3016 34539 3062
rect 34587 3016 34633 3062
rect 34681 3016 34727 3062
rect 34775 3016 34821 3062
rect 34869 3016 34915 3062
rect 34963 3016 35009 3062
rect 35057 3016 35103 3062
rect 35151 3016 35197 3062
rect 35245 3016 35291 3062
rect 35339 3016 35385 3062
rect 35433 3016 35479 3062
rect 35527 3016 35573 3062
rect 35621 3016 35667 3062
rect 35715 3016 35761 3062
rect 35809 3016 35855 3062
rect 35903 3016 35949 3062
rect 35997 3016 36043 3062
rect 36091 3016 36137 3062
rect 36185 3016 36231 3062
rect 36279 3016 36325 3062
rect 36373 3016 36419 3062
rect 36467 3016 36513 3062
rect 36561 3016 36607 3062
rect 36655 3016 36701 3062
rect 36749 3016 36795 3062
rect 36843 3016 36889 3062
rect 36937 3016 36983 3062
rect 37031 3016 37077 3062
rect 37125 3016 37171 3062
rect 37219 3016 37265 3062
rect 37313 3016 37359 3062
rect 37407 3016 37453 3062
rect 37501 3016 37547 3062
rect 37595 3016 37641 3062
rect 37689 3016 37735 3062
rect 37783 3016 37829 3062
rect 37877 3016 37923 3062
rect 37971 3016 38017 3062
rect 38065 3016 38111 3062
rect 38159 3016 38205 3062
rect 38253 3016 38299 3062
rect 38347 3016 38393 3062
rect 38441 3016 38487 3062
rect 38535 3016 38581 3062
rect 38629 3016 38675 3062
rect 38723 3016 38769 3062
rect 38817 3016 38863 3062
rect 38911 3016 38957 3062
rect 39005 3016 39051 3062
rect 39099 3016 39145 3062
rect 39193 3016 39239 3062
rect 39287 3016 39333 3062
rect 39381 3016 39427 3062
rect 39475 3016 39521 3062
rect 39569 3016 39615 3062
rect 39663 3016 39709 3062
rect 39757 3016 39803 3062
rect 39851 3016 39897 3062
rect 39945 3016 39991 3062
rect 40039 3016 40085 3062
rect 40133 3016 40179 3062
rect 40227 3016 40273 3062
rect 40321 3016 40367 3062
rect 40415 3016 40461 3062
rect 32143 2922 32189 2968
rect 32143 2828 32189 2874
rect 32143 2734 32189 2780
rect 32143 2640 32189 2686
rect 36279 2922 36325 2968
rect 36279 2828 36325 2874
rect 36279 2734 36325 2780
rect 36279 2640 36325 2686
rect 40415 2922 40461 2968
rect 40415 2828 40461 2874
rect 40415 2734 40461 2780
rect 32143 2546 32189 2592
rect 40415 2640 40461 2686
rect 36279 2546 36325 2592
rect 32143 2452 32189 2498
rect 32143 2358 32189 2404
rect 32143 2264 32189 2310
rect 32143 2170 32189 2216
rect 32143 2076 32189 2122
rect 32143 1982 32189 2028
rect 32143 1888 32189 1934
rect 40415 2546 40461 2592
rect 36279 2452 36325 2498
rect 36279 2358 36325 2404
rect 36279 2264 36325 2310
rect 36279 2170 36325 2216
rect 36279 2076 36325 2122
rect 36279 1982 36325 2028
rect 32143 1794 32189 1840
rect 32143 1700 32189 1746
rect 32143 1606 32189 1652
rect 32143 1512 32189 1558
rect 32143 1418 32189 1464
rect 32143 1324 32189 1370
rect 32143 1230 32189 1276
rect 32143 1136 32189 1182
rect 32143 1042 32189 1088
rect 32143 948 32189 994
rect 32143 854 32189 900
rect 32143 760 32189 806
rect 32143 666 32189 712
rect 32143 572 32189 618
rect 32143 478 32189 524
rect 32143 384 32189 430
rect 32143 290 32189 336
rect 32143 196 32189 242
rect 32143 102 32189 148
rect 32143 8 32189 54
rect 32143 -86 32189 -40
rect 32143 -180 32189 -134
rect 32143 -274 32189 -228
rect 32143 -368 32189 -322
rect 36279 1888 36325 1934
rect 40415 2452 40461 2498
rect 40415 2358 40461 2404
rect 40415 2264 40461 2310
rect 40415 2170 40461 2216
rect 40415 2076 40461 2122
rect 40415 1982 40461 2028
rect 36279 1794 36325 1840
rect 36279 1700 36325 1746
rect 32143 -462 32189 -416
rect 32143 -556 32189 -510
rect 32143 -650 32189 -604
rect 36279 1606 36325 1652
rect 36279 1512 36325 1558
rect 36279 1418 36325 1464
rect 36279 1324 36325 1370
rect 36279 1230 36325 1276
rect 36279 1136 36325 1182
rect 36279 1042 36325 1088
rect 36279 948 36325 994
rect 36279 854 36325 900
rect 36279 760 36325 806
rect 36279 666 36325 712
rect 36279 572 36325 618
rect 36279 478 36325 524
rect 36279 384 36325 430
rect 36279 290 36325 336
rect 36279 196 36325 242
rect 36279 102 36325 148
rect 36279 8 36325 54
rect 36279 -86 36325 -40
rect 36279 -180 36325 -134
rect 36279 -274 36325 -228
rect 36279 -368 36325 -322
rect 40415 1888 40461 1934
rect 40415 1794 40461 1840
rect 40415 1700 40461 1746
rect 36279 -462 36325 -416
rect 36279 -556 36325 -510
rect 32143 -744 32189 -698
rect 32143 -838 32189 -792
rect 32143 -932 32189 -886
rect 32143 -1026 32189 -980
rect 32143 -1120 32189 -1074
rect 32143 -1214 32189 -1168
rect 32143 -1308 32189 -1262
rect 32143 -1402 32189 -1356
rect 32143 -1496 32189 -1450
rect 32143 -1590 32189 -1544
rect 32143 -1684 32189 -1638
rect 36279 -650 36325 -604
rect 40415 1606 40461 1652
rect 40415 1512 40461 1558
rect 40415 1418 40461 1464
rect 40415 1324 40461 1370
rect 40415 1230 40461 1276
rect 40415 1136 40461 1182
rect 40415 1042 40461 1088
rect 40415 948 40461 994
rect 40415 854 40461 900
rect 40415 760 40461 806
rect 40415 666 40461 712
rect 40415 572 40461 618
rect 40415 478 40461 524
rect 40415 384 40461 430
rect 40415 290 40461 336
rect 40415 196 40461 242
rect 40415 102 40461 148
rect 40415 8 40461 54
rect 40415 -86 40461 -40
rect 40415 -180 40461 -134
rect 40415 -274 40461 -228
rect 40415 -368 40461 -322
rect 40415 -462 40461 -416
rect 40415 -556 40461 -510
rect 36279 -744 36325 -698
rect 36279 -838 36325 -792
rect 36279 -932 36325 -886
rect 36279 -1026 36325 -980
rect 36279 -1120 36325 -1074
rect 36279 -1214 36325 -1168
rect 36279 -1308 36325 -1262
rect 36279 -1402 36325 -1356
rect 36279 -1496 36325 -1450
rect 36279 -1590 36325 -1544
rect 36279 -1684 36325 -1638
rect 40415 -650 40461 -604
rect 40415 -744 40461 -698
rect 40415 -838 40461 -792
rect 40415 -932 40461 -886
rect 40415 -1026 40461 -980
rect 40415 -1120 40461 -1074
rect 40415 -1214 40461 -1168
rect 40415 -1308 40461 -1262
rect 40415 -1402 40461 -1356
rect 40415 -1496 40461 -1450
rect 40415 -1590 40461 -1544
rect 40415 -1684 40461 -1638
rect 32143 -1778 32189 -1732
rect 32237 -1778 32283 -1732
rect 32331 -1778 32377 -1732
rect 32425 -1778 32471 -1732
rect 32519 -1778 32565 -1732
rect 32613 -1778 32659 -1732
rect 32707 -1778 32753 -1732
rect 32801 -1778 32847 -1732
rect 32895 -1778 32941 -1732
rect 32989 -1778 33035 -1732
rect 33083 -1778 33129 -1732
rect 33177 -1778 33223 -1732
rect 33271 -1778 33317 -1732
rect 33365 -1778 33411 -1732
rect 33459 -1778 33505 -1732
rect 33553 -1778 33599 -1732
rect 33647 -1778 33693 -1732
rect 33741 -1778 33787 -1732
rect 33835 -1778 33881 -1732
rect 33929 -1778 33975 -1732
rect 34023 -1778 34069 -1732
rect 34117 -1778 34163 -1732
rect 34211 -1778 34257 -1732
rect 34305 -1778 34351 -1732
rect 34399 -1778 34445 -1732
rect 34493 -1778 34539 -1732
rect 34587 -1778 34633 -1732
rect 34681 -1778 34727 -1732
rect 34775 -1778 34821 -1732
rect 34869 -1778 34915 -1732
rect 34963 -1778 35009 -1732
rect 35057 -1778 35103 -1732
rect 35151 -1778 35197 -1732
rect 35245 -1778 35291 -1732
rect 35339 -1778 35385 -1732
rect 35433 -1778 35479 -1732
rect 35527 -1778 35573 -1732
rect 35621 -1778 35667 -1732
rect 35715 -1778 35761 -1732
rect 35809 -1778 35855 -1732
rect 35903 -1778 35949 -1732
rect 35997 -1778 36043 -1732
rect 36091 -1778 36137 -1732
rect 36185 -1778 36231 -1732
rect 36279 -1778 36325 -1732
rect 36373 -1778 36419 -1732
rect 36467 -1778 36513 -1732
rect 36561 -1778 36607 -1732
rect 36655 -1778 36701 -1732
rect 36749 -1778 36795 -1732
rect 36843 -1778 36889 -1732
rect 36937 -1778 36983 -1732
rect 37031 -1778 37077 -1732
rect 37125 -1778 37171 -1732
rect 37219 -1778 37265 -1732
rect 37313 -1778 37359 -1732
rect 37407 -1778 37453 -1732
rect 37501 -1778 37547 -1732
rect 37595 -1778 37641 -1732
rect 37689 -1778 37735 -1732
rect 37783 -1778 37829 -1732
rect 37877 -1778 37923 -1732
rect 37971 -1778 38017 -1732
rect 38065 -1778 38111 -1732
rect 38159 -1778 38205 -1732
rect 38253 -1778 38299 -1732
rect 38347 -1778 38393 -1732
rect 38441 -1778 38487 -1732
rect 38535 -1778 38581 -1732
rect 38629 -1778 38675 -1732
rect 38723 -1778 38769 -1732
rect 38817 -1778 38863 -1732
rect 38911 -1778 38957 -1732
rect 39005 -1778 39051 -1732
rect 39099 -1778 39145 -1732
rect 39193 -1778 39239 -1732
rect 39287 -1778 39333 -1732
rect 39381 -1778 39427 -1732
rect 39475 -1778 39521 -1732
rect 39569 -1778 39615 -1732
rect 39663 -1778 39709 -1732
rect 39757 -1778 39803 -1732
rect 39851 -1778 39897 -1732
rect 39945 -1778 39991 -1732
rect 40039 -1778 40085 -1732
rect 40133 -1778 40179 -1732
rect 40227 -1778 40273 -1732
rect 40321 -1778 40367 -1732
rect 40415 -1778 40461 -1732
rect 41839 3016 41885 3062
rect 41933 3016 41979 3062
rect 42027 3016 42073 3062
rect 42121 3016 42167 3062
rect 42215 3016 42261 3062
rect 42309 3016 42355 3062
rect 42403 3016 42449 3062
rect 42497 3016 42543 3062
rect 42591 3016 42637 3062
rect 42685 3016 42731 3062
rect 42779 3016 42825 3062
rect 42873 3016 42919 3062
rect 42967 3016 43013 3062
rect 43061 3016 43107 3062
rect 43155 3016 43201 3062
rect 43249 3016 43295 3062
rect 43343 3016 43389 3062
rect 43437 3016 43483 3062
rect 43531 3016 43577 3062
rect 43625 3016 43671 3062
rect 43719 3016 43765 3062
rect 43813 3016 43859 3062
rect 43907 3016 43953 3062
rect 44001 3016 44047 3062
rect 44095 3016 44141 3062
rect 44189 3016 44235 3062
rect 44283 3016 44329 3062
rect 44377 3016 44423 3062
rect 44471 3016 44517 3062
rect 44565 3016 44611 3062
rect 44659 3016 44705 3062
rect 44753 3016 44799 3062
rect 44847 3016 44893 3062
rect 44941 3016 44987 3062
rect 45035 3016 45081 3062
rect 45129 3016 45175 3062
rect 45223 3016 45269 3062
rect 45317 3016 45363 3062
rect 45411 3016 45457 3062
rect 45505 3016 45551 3062
rect 45599 3016 45645 3062
rect 45693 3016 45739 3062
rect 45787 3016 45833 3062
rect 45881 3016 45927 3062
rect 45975 3016 46021 3062
rect 46069 3016 46115 3062
rect 46163 3016 46209 3062
rect 46257 3016 46303 3062
rect 46351 3016 46397 3062
rect 46445 3016 46491 3062
rect 46539 3016 46585 3062
rect 46633 3016 46679 3062
rect 46727 3016 46773 3062
rect 46821 3016 46867 3062
rect 46915 3016 46961 3062
rect 47009 3016 47055 3062
rect 47103 3016 47149 3062
rect 47197 3016 47243 3062
rect 47291 3016 47337 3062
rect 47385 3016 47431 3062
rect 47479 3016 47525 3062
rect 47573 3016 47619 3062
rect 47667 3016 47713 3062
rect 47761 3016 47807 3062
rect 47855 3016 47901 3062
rect 47949 3016 47995 3062
rect 48043 3016 48089 3062
rect 48137 3016 48183 3062
rect 48231 3016 48277 3062
rect 48325 3016 48371 3062
rect 48419 3016 48465 3062
rect 48513 3016 48559 3062
rect 48607 3016 48653 3062
rect 48701 3016 48747 3062
rect 48795 3016 48841 3062
rect 48889 3016 48935 3062
rect 48983 3016 49029 3062
rect 49077 3016 49123 3062
rect 49171 3016 49217 3062
rect 49265 3016 49311 3062
rect 49359 3016 49405 3062
rect 49453 3016 49499 3062
rect 49547 3016 49593 3062
rect 49641 3016 49687 3062
rect 49735 3016 49781 3062
rect 49829 3016 49875 3062
rect 49923 3016 49969 3062
rect 50017 3016 50063 3062
rect 50111 3016 50157 3062
rect 41839 2922 41885 2968
rect 41839 2828 41885 2874
rect 41839 2734 41885 2780
rect 41839 2640 41885 2686
rect 45975 2922 46021 2968
rect 45975 2828 46021 2874
rect 45975 2734 46021 2780
rect 45975 2640 46021 2686
rect 50111 2922 50157 2968
rect 50111 2828 50157 2874
rect 50111 2734 50157 2780
rect 41839 2546 41885 2592
rect 50111 2640 50157 2686
rect 45975 2546 46021 2592
rect 41839 2452 41885 2498
rect 41839 2358 41885 2404
rect 41839 2264 41885 2310
rect 41839 2170 41885 2216
rect 41839 2076 41885 2122
rect 41839 1982 41885 2028
rect 41839 1888 41885 1934
rect 50111 2546 50157 2592
rect 45975 2452 46021 2498
rect 45975 2358 46021 2404
rect 45975 2264 46021 2310
rect 45975 2170 46021 2216
rect 45975 2076 46021 2122
rect 45975 1982 46021 2028
rect 41839 1794 41885 1840
rect 41839 1700 41885 1746
rect 41839 1606 41885 1652
rect 41839 1512 41885 1558
rect 41839 1418 41885 1464
rect 41839 1324 41885 1370
rect 41839 1230 41885 1276
rect 41839 1136 41885 1182
rect 41839 1042 41885 1088
rect 41839 948 41885 994
rect 41839 854 41885 900
rect 41839 760 41885 806
rect 41839 666 41885 712
rect 41839 572 41885 618
rect 41839 478 41885 524
rect 41839 384 41885 430
rect 41839 290 41885 336
rect 41839 196 41885 242
rect 41839 102 41885 148
rect 41839 8 41885 54
rect 41839 -86 41885 -40
rect 41839 -180 41885 -134
rect 41839 -274 41885 -228
rect 41839 -368 41885 -322
rect 45975 1888 46021 1934
rect 50111 2452 50157 2498
rect 50111 2358 50157 2404
rect 50111 2264 50157 2310
rect 50111 2170 50157 2216
rect 50111 2076 50157 2122
rect 50111 1982 50157 2028
rect 45975 1794 46021 1840
rect 45975 1700 46021 1746
rect 41839 -462 41885 -416
rect 41839 -556 41885 -510
rect 41839 -650 41885 -604
rect 45975 1606 46021 1652
rect 45975 1512 46021 1558
rect 45975 1418 46021 1464
rect 45975 1324 46021 1370
rect 45975 1230 46021 1276
rect 45975 1136 46021 1182
rect 45975 1042 46021 1088
rect 45975 948 46021 994
rect 45975 854 46021 900
rect 45975 760 46021 806
rect 45975 666 46021 712
rect 45975 572 46021 618
rect 45975 478 46021 524
rect 45975 384 46021 430
rect 45975 290 46021 336
rect 45975 196 46021 242
rect 45975 102 46021 148
rect 45975 8 46021 54
rect 45975 -86 46021 -40
rect 45975 -180 46021 -134
rect 45975 -274 46021 -228
rect 45975 -368 46021 -322
rect 50111 1888 50157 1934
rect 50111 1794 50157 1840
rect 50111 1700 50157 1746
rect 45975 -462 46021 -416
rect 45975 -556 46021 -510
rect 41839 -744 41885 -698
rect 41839 -838 41885 -792
rect 41839 -932 41885 -886
rect 41839 -1026 41885 -980
rect 41839 -1120 41885 -1074
rect 41839 -1214 41885 -1168
rect 41839 -1308 41885 -1262
rect 41839 -1402 41885 -1356
rect 41839 -1496 41885 -1450
rect 41839 -1590 41885 -1544
rect 41839 -1684 41885 -1638
rect 45975 -650 46021 -604
rect 50111 1606 50157 1652
rect 50111 1512 50157 1558
rect 50111 1418 50157 1464
rect 50111 1324 50157 1370
rect 50111 1230 50157 1276
rect 50111 1136 50157 1182
rect 50111 1042 50157 1088
rect 50111 948 50157 994
rect 50111 854 50157 900
rect 50111 760 50157 806
rect 50111 666 50157 712
rect 50111 572 50157 618
rect 50111 478 50157 524
rect 50111 384 50157 430
rect 50111 290 50157 336
rect 50111 196 50157 242
rect 50111 102 50157 148
rect 50111 8 50157 54
rect 50111 -86 50157 -40
rect 50111 -180 50157 -134
rect 50111 -274 50157 -228
rect 50111 -368 50157 -322
rect 50111 -462 50157 -416
rect 50111 -556 50157 -510
rect 45975 -744 46021 -698
rect 45975 -838 46021 -792
rect 45975 -932 46021 -886
rect 45975 -1026 46021 -980
rect 45975 -1120 46021 -1074
rect 45975 -1214 46021 -1168
rect 45975 -1308 46021 -1262
rect 45975 -1402 46021 -1356
rect 45975 -1496 46021 -1450
rect 45975 -1590 46021 -1544
rect 45975 -1684 46021 -1638
rect 50111 -650 50157 -604
rect 50111 -744 50157 -698
rect 50111 -838 50157 -792
rect 50111 -932 50157 -886
rect 50111 -1026 50157 -980
rect 50111 -1120 50157 -1074
rect 50111 -1214 50157 -1168
rect 50111 -1308 50157 -1262
rect 50111 -1402 50157 -1356
rect 50111 -1496 50157 -1450
rect 50111 -1590 50157 -1544
rect 50111 -1684 50157 -1638
rect 41839 -1778 41885 -1732
rect 41933 -1778 41979 -1732
rect 42027 -1778 42073 -1732
rect 42121 -1778 42167 -1732
rect 42215 -1778 42261 -1732
rect 42309 -1778 42355 -1732
rect 42403 -1778 42449 -1732
rect 42497 -1778 42543 -1732
rect 42591 -1778 42637 -1732
rect 42685 -1778 42731 -1732
rect 42779 -1778 42825 -1732
rect 42873 -1778 42919 -1732
rect 42967 -1778 43013 -1732
rect 43061 -1778 43107 -1732
rect 43155 -1778 43201 -1732
rect 43249 -1778 43295 -1732
rect 43343 -1778 43389 -1732
rect 43437 -1778 43483 -1732
rect 43531 -1778 43577 -1732
rect 43625 -1778 43671 -1732
rect 43719 -1778 43765 -1732
rect 43813 -1778 43859 -1732
rect 43907 -1778 43953 -1732
rect 44001 -1778 44047 -1732
rect 44095 -1778 44141 -1732
rect 44189 -1778 44235 -1732
rect 44283 -1778 44329 -1732
rect 44377 -1778 44423 -1732
rect 44471 -1778 44517 -1732
rect 44565 -1778 44611 -1732
rect 44659 -1778 44705 -1732
rect 44753 -1778 44799 -1732
rect 44847 -1778 44893 -1732
rect 44941 -1778 44987 -1732
rect 45035 -1778 45081 -1732
rect 45129 -1778 45175 -1732
rect 45223 -1778 45269 -1732
rect 45317 -1778 45363 -1732
rect 45411 -1778 45457 -1732
rect 45505 -1778 45551 -1732
rect 45599 -1778 45645 -1732
rect 45693 -1778 45739 -1732
rect 45787 -1778 45833 -1732
rect 45881 -1778 45927 -1732
rect 45975 -1778 46021 -1732
rect 46069 -1778 46115 -1732
rect 46163 -1778 46209 -1732
rect 46257 -1778 46303 -1732
rect 46351 -1778 46397 -1732
rect 46445 -1778 46491 -1732
rect 46539 -1778 46585 -1732
rect 46633 -1778 46679 -1732
rect 46727 -1778 46773 -1732
rect 46821 -1778 46867 -1732
rect 46915 -1778 46961 -1732
rect 47009 -1778 47055 -1732
rect 47103 -1778 47149 -1732
rect 47197 -1778 47243 -1732
rect 47291 -1778 47337 -1732
rect 47385 -1778 47431 -1732
rect 47479 -1778 47525 -1732
rect 47573 -1778 47619 -1732
rect 47667 -1778 47713 -1732
rect 47761 -1778 47807 -1732
rect 47855 -1778 47901 -1732
rect 47949 -1778 47995 -1732
rect 48043 -1778 48089 -1732
rect 48137 -1778 48183 -1732
rect 48231 -1778 48277 -1732
rect 48325 -1778 48371 -1732
rect 48419 -1778 48465 -1732
rect 48513 -1778 48559 -1732
rect 48607 -1778 48653 -1732
rect 48701 -1778 48747 -1732
rect 48795 -1778 48841 -1732
rect 48889 -1778 48935 -1732
rect 48983 -1778 49029 -1732
rect 49077 -1778 49123 -1732
rect 49171 -1778 49217 -1732
rect 49265 -1778 49311 -1732
rect 49359 -1778 49405 -1732
rect 49453 -1778 49499 -1732
rect 49547 -1778 49593 -1732
rect 49641 -1778 49687 -1732
rect 49735 -1778 49781 -1732
rect 49829 -1778 49875 -1732
rect 49923 -1778 49969 -1732
rect 50017 -1778 50063 -1732
rect 50111 -1778 50157 -1732
rect 51535 3016 51581 3062
rect 51629 3016 51675 3062
rect 51723 3016 51769 3062
rect 51817 3016 51863 3062
rect 51911 3016 51957 3062
rect 52005 3016 52051 3062
rect 52099 3016 52145 3062
rect 52193 3016 52239 3062
rect 52287 3016 52333 3062
rect 52381 3016 52427 3062
rect 52475 3016 52521 3062
rect 52569 3016 52615 3062
rect 52663 3016 52709 3062
rect 52757 3016 52803 3062
rect 52851 3016 52897 3062
rect 52945 3016 52991 3062
rect 53039 3016 53085 3062
rect 53133 3016 53179 3062
rect 53227 3016 53273 3062
rect 53321 3016 53367 3062
rect 53415 3016 53461 3062
rect 53509 3016 53555 3062
rect 53603 3016 53649 3062
rect 53697 3016 53743 3062
rect 53791 3016 53837 3062
rect 53885 3016 53931 3062
rect 53979 3016 54025 3062
rect 54073 3016 54119 3062
rect 54167 3016 54213 3062
rect 54261 3016 54307 3062
rect 54355 3016 54401 3062
rect 54449 3016 54495 3062
rect 54543 3016 54589 3062
rect 54637 3016 54683 3062
rect 54731 3016 54777 3062
rect 54825 3016 54871 3062
rect 54919 3016 54965 3062
rect 55013 3016 55059 3062
rect 55107 3016 55153 3062
rect 55201 3016 55247 3062
rect 55295 3016 55341 3062
rect 55389 3016 55435 3062
rect 55483 3016 55529 3062
rect 55577 3016 55623 3062
rect 55671 3016 55717 3062
rect 55765 3016 55811 3062
rect 55859 3016 55905 3062
rect 55953 3016 55999 3062
rect 56047 3016 56093 3062
rect 56141 3016 56187 3062
rect 56235 3016 56281 3062
rect 56329 3016 56375 3062
rect 56423 3016 56469 3062
rect 56517 3016 56563 3062
rect 56611 3016 56657 3062
rect 56705 3016 56751 3062
rect 56799 3016 56845 3062
rect 56893 3016 56939 3062
rect 56987 3016 57033 3062
rect 57081 3016 57127 3062
rect 57175 3016 57221 3062
rect 57269 3016 57315 3062
rect 57363 3016 57409 3062
rect 57457 3016 57503 3062
rect 57551 3016 57597 3062
rect 57645 3016 57691 3062
rect 57739 3016 57785 3062
rect 57833 3016 57879 3062
rect 57927 3016 57973 3062
rect 58021 3016 58067 3062
rect 58115 3016 58161 3062
rect 58209 3016 58255 3062
rect 58303 3016 58349 3062
rect 58397 3016 58443 3062
rect 58491 3016 58537 3062
rect 58585 3016 58631 3062
rect 58679 3016 58725 3062
rect 58773 3016 58819 3062
rect 58867 3016 58913 3062
rect 58961 3016 59007 3062
rect 59055 3016 59101 3062
rect 59149 3016 59195 3062
rect 59243 3016 59289 3062
rect 59337 3016 59383 3062
rect 59431 3016 59477 3062
rect 59525 3016 59571 3062
rect 59619 3016 59665 3062
rect 59713 3016 59759 3062
rect 59807 3016 59853 3062
rect 51535 2922 51581 2968
rect 51535 2828 51581 2874
rect 51535 2734 51581 2780
rect 51535 2640 51581 2686
rect 55671 2922 55717 2968
rect 55671 2828 55717 2874
rect 55671 2734 55717 2780
rect 55671 2640 55717 2686
rect 59807 2922 59853 2968
rect 59807 2828 59853 2874
rect 59807 2734 59853 2780
rect 51535 2546 51581 2592
rect 59807 2640 59853 2686
rect 55671 2546 55717 2592
rect 51535 2452 51581 2498
rect 51535 2358 51581 2404
rect 51535 2264 51581 2310
rect 51535 2170 51581 2216
rect 51535 2076 51581 2122
rect 51535 1982 51581 2028
rect 51535 1888 51581 1934
rect 59807 2546 59853 2592
rect 55671 2452 55717 2498
rect 55671 2358 55717 2404
rect 55671 2264 55717 2310
rect 55671 2170 55717 2216
rect 55671 2076 55717 2122
rect 55671 1982 55717 2028
rect 51535 1794 51581 1840
rect 51535 1700 51581 1746
rect 51535 1606 51581 1652
rect 51535 1512 51581 1558
rect 51535 1418 51581 1464
rect 51535 1324 51581 1370
rect 51535 1230 51581 1276
rect 51535 1136 51581 1182
rect 51535 1042 51581 1088
rect 51535 948 51581 994
rect 51535 854 51581 900
rect 51535 760 51581 806
rect 51535 666 51581 712
rect 51535 572 51581 618
rect 51535 478 51581 524
rect 51535 384 51581 430
rect 51535 290 51581 336
rect 51535 196 51581 242
rect 51535 102 51581 148
rect 51535 8 51581 54
rect 51535 -86 51581 -40
rect 51535 -180 51581 -134
rect 51535 -274 51581 -228
rect 51535 -368 51581 -322
rect 55671 1888 55717 1934
rect 59807 2452 59853 2498
rect 59807 2358 59853 2404
rect 59807 2264 59853 2310
rect 59807 2170 59853 2216
rect 59807 2076 59853 2122
rect 59807 1982 59853 2028
rect 55671 1794 55717 1840
rect 55671 1700 55717 1746
rect 51535 -462 51581 -416
rect 51535 -556 51581 -510
rect 51535 -650 51581 -604
rect 55671 1606 55717 1652
rect 55671 1512 55717 1558
rect 55671 1418 55717 1464
rect 55671 1324 55717 1370
rect 55671 1230 55717 1276
rect 55671 1136 55717 1182
rect 55671 1042 55717 1088
rect 55671 948 55717 994
rect 55671 854 55717 900
rect 55671 760 55717 806
rect 55671 666 55717 712
rect 55671 572 55717 618
rect 55671 478 55717 524
rect 55671 384 55717 430
rect 55671 290 55717 336
rect 55671 196 55717 242
rect 55671 102 55717 148
rect 55671 8 55717 54
rect 55671 -86 55717 -40
rect 55671 -180 55717 -134
rect 55671 -274 55717 -228
rect 55671 -368 55717 -322
rect 59807 1888 59853 1934
rect 59807 1794 59853 1840
rect 59807 1700 59853 1746
rect 55671 -462 55717 -416
rect 55671 -556 55717 -510
rect 51535 -744 51581 -698
rect 51535 -838 51581 -792
rect 51535 -932 51581 -886
rect 51535 -1026 51581 -980
rect 51535 -1120 51581 -1074
rect 51535 -1214 51581 -1168
rect 51535 -1308 51581 -1262
rect 51535 -1402 51581 -1356
rect 51535 -1496 51581 -1450
rect 51535 -1590 51581 -1544
rect 51535 -1684 51581 -1638
rect 55671 -650 55717 -604
rect 59807 1606 59853 1652
rect 59807 1512 59853 1558
rect 59807 1418 59853 1464
rect 59807 1324 59853 1370
rect 59807 1230 59853 1276
rect 59807 1136 59853 1182
rect 59807 1042 59853 1088
rect 59807 948 59853 994
rect 59807 854 59853 900
rect 59807 760 59853 806
rect 59807 666 59853 712
rect 59807 572 59853 618
rect 59807 478 59853 524
rect 59807 384 59853 430
rect 59807 290 59853 336
rect 59807 196 59853 242
rect 59807 102 59853 148
rect 59807 8 59853 54
rect 59807 -86 59853 -40
rect 59807 -180 59853 -134
rect 59807 -274 59853 -228
rect 59807 -368 59853 -322
rect 59807 -462 59853 -416
rect 59807 -556 59853 -510
rect 55671 -744 55717 -698
rect 55671 -838 55717 -792
rect 55671 -932 55717 -886
rect 55671 -1026 55717 -980
rect 55671 -1120 55717 -1074
rect 55671 -1214 55717 -1168
rect 55671 -1308 55717 -1262
rect 55671 -1402 55717 -1356
rect 55671 -1496 55717 -1450
rect 55671 -1590 55717 -1544
rect 55671 -1684 55717 -1638
rect 59807 -650 59853 -604
rect 59807 -744 59853 -698
rect 59807 -838 59853 -792
rect 59807 -932 59853 -886
rect 59807 -1026 59853 -980
rect 59807 -1120 59853 -1074
rect 59807 -1214 59853 -1168
rect 59807 -1308 59853 -1262
rect 59807 -1402 59853 -1356
rect 59807 -1496 59853 -1450
rect 59807 -1590 59853 -1544
rect 59807 -1684 59853 -1638
rect 51535 -1778 51581 -1732
rect 51629 -1778 51675 -1732
rect 51723 -1778 51769 -1732
rect 51817 -1778 51863 -1732
rect 51911 -1778 51957 -1732
rect 52005 -1778 52051 -1732
rect 52099 -1778 52145 -1732
rect 52193 -1778 52239 -1732
rect 52287 -1778 52333 -1732
rect 52381 -1778 52427 -1732
rect 52475 -1778 52521 -1732
rect 52569 -1778 52615 -1732
rect 52663 -1778 52709 -1732
rect 52757 -1778 52803 -1732
rect 52851 -1778 52897 -1732
rect 52945 -1778 52991 -1732
rect 53039 -1778 53085 -1732
rect 53133 -1778 53179 -1732
rect 53227 -1778 53273 -1732
rect 53321 -1778 53367 -1732
rect 53415 -1778 53461 -1732
rect 53509 -1778 53555 -1732
rect 53603 -1778 53649 -1732
rect 53697 -1778 53743 -1732
rect 53791 -1778 53837 -1732
rect 53885 -1778 53931 -1732
rect 53979 -1778 54025 -1732
rect 54073 -1778 54119 -1732
rect 54167 -1778 54213 -1732
rect 54261 -1778 54307 -1732
rect 54355 -1778 54401 -1732
rect 54449 -1778 54495 -1732
rect 54543 -1778 54589 -1732
rect 54637 -1778 54683 -1732
rect 54731 -1778 54777 -1732
rect 54825 -1778 54871 -1732
rect 54919 -1778 54965 -1732
rect 55013 -1778 55059 -1732
rect 55107 -1778 55153 -1732
rect 55201 -1778 55247 -1732
rect 55295 -1778 55341 -1732
rect 55389 -1778 55435 -1732
rect 55483 -1778 55529 -1732
rect 55577 -1778 55623 -1732
rect 55671 -1778 55717 -1732
rect 55765 -1778 55811 -1732
rect 55859 -1778 55905 -1732
rect 55953 -1778 55999 -1732
rect 56047 -1778 56093 -1732
rect 56141 -1778 56187 -1732
rect 56235 -1778 56281 -1732
rect 56329 -1778 56375 -1732
rect 56423 -1778 56469 -1732
rect 56517 -1778 56563 -1732
rect 56611 -1778 56657 -1732
rect 56705 -1778 56751 -1732
rect 56799 -1778 56845 -1732
rect 56893 -1778 56939 -1732
rect 56987 -1778 57033 -1732
rect 57081 -1778 57127 -1732
rect 57175 -1778 57221 -1732
rect 57269 -1778 57315 -1732
rect 57363 -1778 57409 -1732
rect 57457 -1778 57503 -1732
rect 57551 -1778 57597 -1732
rect 57645 -1778 57691 -1732
rect 57739 -1778 57785 -1732
rect 57833 -1778 57879 -1732
rect 57927 -1778 57973 -1732
rect 58021 -1778 58067 -1732
rect 58115 -1778 58161 -1732
rect 58209 -1778 58255 -1732
rect 58303 -1778 58349 -1732
rect 58397 -1778 58443 -1732
rect 58491 -1778 58537 -1732
rect 58585 -1778 58631 -1732
rect 58679 -1778 58725 -1732
rect 58773 -1778 58819 -1732
rect 58867 -1778 58913 -1732
rect 58961 -1778 59007 -1732
rect 59055 -1778 59101 -1732
rect 59149 -1778 59195 -1732
rect 59243 -1778 59289 -1732
rect 59337 -1778 59383 -1732
rect 59431 -1778 59477 -1732
rect 59525 -1778 59571 -1732
rect 59619 -1778 59665 -1732
rect 59713 -1778 59759 -1732
rect 59807 -1778 59853 -1732
rect 61231 3016 61277 3062
rect 61325 3016 61371 3062
rect 61419 3016 61465 3062
rect 61513 3016 61559 3062
rect 61607 3016 61653 3062
rect 61701 3016 61747 3062
rect 61795 3016 61841 3062
rect 61889 3016 61935 3062
rect 61983 3016 62029 3062
rect 62077 3016 62123 3062
rect 62171 3016 62217 3062
rect 62265 3016 62311 3062
rect 62359 3016 62405 3062
rect 62453 3016 62499 3062
rect 62547 3016 62593 3062
rect 62641 3016 62687 3062
rect 62735 3016 62781 3062
rect 62829 3016 62875 3062
rect 62923 3016 62969 3062
rect 63017 3016 63063 3062
rect 63111 3016 63157 3062
rect 63205 3016 63251 3062
rect 63299 3016 63345 3062
rect 63393 3016 63439 3062
rect 63487 3016 63533 3062
rect 63581 3016 63627 3062
rect 63675 3016 63721 3062
rect 63769 3016 63815 3062
rect 63863 3016 63909 3062
rect 63957 3016 64003 3062
rect 64051 3016 64097 3062
rect 64145 3016 64191 3062
rect 64239 3016 64285 3062
rect 64333 3016 64379 3062
rect 64427 3016 64473 3062
rect 64521 3016 64567 3062
rect 64615 3016 64661 3062
rect 64709 3016 64755 3062
rect 64803 3016 64849 3062
rect 64897 3016 64943 3062
rect 64991 3016 65037 3062
rect 65085 3016 65131 3062
rect 65179 3016 65225 3062
rect 65273 3016 65319 3062
rect 65367 3016 65413 3062
rect 61231 2922 61277 2968
rect 61231 2828 61277 2874
rect 61231 2734 61277 2780
rect 61231 2640 61277 2686
rect 65367 2922 65413 2968
rect 65367 2828 65413 2874
rect 65367 2734 65413 2780
rect 65367 2640 65413 2686
rect 61231 2546 61277 2592
rect 65367 2546 65413 2592
rect 61231 2452 61277 2498
rect 61231 2358 61277 2404
rect 61231 2264 61277 2310
rect 61231 2170 61277 2216
rect 61231 2076 61277 2122
rect 61231 1982 61277 2028
rect 61231 1888 61277 1934
rect 65367 2452 65413 2498
rect 65367 2358 65413 2404
rect 65367 2264 65413 2310
rect 65367 2170 65413 2216
rect 65367 2076 65413 2122
rect 65367 1982 65413 2028
rect 61231 1794 61277 1840
rect 61231 1700 61277 1746
rect 61231 1606 61277 1652
rect 61231 1512 61277 1558
rect 61231 1418 61277 1464
rect 61231 1324 61277 1370
rect 61231 1230 61277 1276
rect 61231 1136 61277 1182
rect 61231 1042 61277 1088
rect 61231 948 61277 994
rect 61231 854 61277 900
rect 61231 760 61277 806
rect 61231 666 61277 712
rect 61231 572 61277 618
rect 61231 478 61277 524
rect 61231 384 61277 430
rect 61231 290 61277 336
rect 61231 196 61277 242
rect 61231 102 61277 148
rect 61231 8 61277 54
rect 61231 -86 61277 -40
rect 61231 -180 61277 -134
rect 61231 -274 61277 -228
rect 61231 -368 61277 -322
rect 65367 1888 65413 1934
rect 65367 1794 65413 1840
rect 65367 1700 65413 1746
rect 61231 -462 61277 -416
rect 61231 -556 61277 -510
rect 61231 -650 61277 -604
rect 65367 1606 65413 1652
rect 65367 1512 65413 1558
rect 65367 1418 65413 1464
rect 65367 1324 65413 1370
rect 65367 1230 65413 1276
rect 65367 1136 65413 1182
rect 65367 1042 65413 1088
rect 65367 948 65413 994
rect 65367 854 65413 900
rect 65367 760 65413 806
rect 65367 666 65413 712
rect 65367 572 65413 618
rect 65367 478 65413 524
rect 65367 384 65413 430
rect 65367 290 65413 336
rect 65367 196 65413 242
rect 65367 102 65413 148
rect 65367 8 65413 54
rect 65367 -86 65413 -40
rect 65367 -180 65413 -134
rect 65367 -274 65413 -228
rect 65367 -368 65413 -322
rect 65367 -462 65413 -416
rect 65367 -556 65413 -510
rect 61231 -744 61277 -698
rect 61231 -838 61277 -792
rect 61231 -932 61277 -886
rect 61231 -1026 61277 -980
rect 61231 -1120 61277 -1074
rect 61231 -1214 61277 -1168
rect 61231 -1308 61277 -1262
rect 61231 -1402 61277 -1356
rect 61231 -1496 61277 -1450
rect 61231 -1590 61277 -1544
rect 61231 -1684 61277 -1638
rect 65367 -650 65413 -604
rect 65367 -744 65413 -698
rect 65367 -838 65413 -792
rect 65367 -932 65413 -886
rect 65367 -1026 65413 -980
rect 65367 -1120 65413 -1074
rect 65367 -1214 65413 -1168
rect 65367 -1308 65413 -1262
rect 65367 -1402 65413 -1356
rect 65367 -1496 65413 -1450
rect 65367 -1590 65413 -1544
rect 65367 -1684 65413 -1638
rect 61231 -1778 61277 -1732
rect 61325 -1778 61371 -1732
rect 61419 -1778 61465 -1732
rect 61513 -1778 61559 -1732
rect 61607 -1778 61653 -1732
rect 61701 -1778 61747 -1732
rect 61795 -1778 61841 -1732
rect 61889 -1778 61935 -1732
rect 61983 -1778 62029 -1732
rect 62077 -1778 62123 -1732
rect 62171 -1778 62217 -1732
rect 62265 -1778 62311 -1732
rect 62359 -1778 62405 -1732
rect 62453 -1778 62499 -1732
rect 62547 -1778 62593 -1732
rect 62641 -1778 62687 -1732
rect 62735 -1778 62781 -1732
rect 62829 -1778 62875 -1732
rect 62923 -1778 62969 -1732
rect 63017 -1778 63063 -1732
rect 63111 -1778 63157 -1732
rect 63205 -1778 63251 -1732
rect 63299 -1778 63345 -1732
rect 63393 -1778 63439 -1732
rect 63487 -1778 63533 -1732
rect 63581 -1778 63627 -1732
rect 63675 -1778 63721 -1732
rect 63769 -1778 63815 -1732
rect 63863 -1778 63909 -1732
rect 63957 -1778 64003 -1732
rect 64051 -1778 64097 -1732
rect 64145 -1778 64191 -1732
rect 64239 -1778 64285 -1732
rect 64333 -1778 64379 -1732
rect 64427 -1778 64473 -1732
rect 64521 -1778 64567 -1732
rect 64615 -1778 64661 -1732
rect 64709 -1778 64755 -1732
rect 64803 -1778 64849 -1732
rect 64897 -1778 64943 -1732
rect 64991 -1778 65037 -1732
rect 65085 -1778 65131 -1732
rect 65179 -1778 65225 -1732
rect 65273 -1778 65319 -1732
rect 65367 -1778 65413 -1732
rect 443 -4411 489 -4365
rect 537 -4411 583 -4365
rect 631 -4411 677 -4365
rect 725 -4411 771 -4365
rect 819 -4411 865 -4365
rect 913 -4411 959 -4365
rect 1007 -4411 1053 -4365
rect 1101 -4411 1147 -4365
rect 1195 -4411 1241 -4365
rect 1289 -4411 1335 -4365
rect 1383 -4411 1429 -4365
rect 1477 -4411 1523 -4365
rect 1571 -4411 1617 -4365
rect 1665 -4411 1711 -4365
rect 1759 -4411 1805 -4365
rect 1853 -4411 1899 -4365
rect 1947 -4411 1993 -4365
rect 2041 -4411 2087 -4365
rect 2135 -4411 2181 -4365
rect 2229 -4411 2275 -4365
rect 2323 -4411 2369 -4365
rect 2417 -4411 2463 -4365
rect 2511 -4411 2557 -4365
rect 2605 -4411 2651 -4365
rect 2699 -4411 2745 -4365
rect 2793 -4411 2839 -4365
rect 2887 -4411 2933 -4365
rect 2981 -4411 3027 -4365
rect 3075 -4411 3121 -4365
rect 3169 -4411 3215 -4365
rect 3263 -4411 3309 -4365
rect 3357 -4411 3403 -4365
rect 3451 -4411 3497 -4365
rect 3545 -4411 3591 -4365
rect 3639 -4411 3685 -4365
rect 3733 -4411 3779 -4365
rect 3827 -4411 3873 -4365
rect 3921 -4411 3967 -4365
rect 4015 -4411 4061 -4365
rect 4109 -4411 4155 -4365
rect 4203 -4411 4249 -4365
rect 4297 -4411 4343 -4365
rect 4391 -4411 4437 -4365
rect 4485 -4411 4531 -4365
rect 443 -4505 489 -4459
rect 443 -4599 489 -4553
rect 4485 -4505 4531 -4459
rect 443 -4693 489 -4647
rect 4485 -4599 4531 -4553
rect 4485 -4693 4531 -4647
rect 443 -4787 489 -4741
rect 443 -4881 489 -4835
rect 443 -4975 489 -4929
rect 443 -5069 489 -5023
rect 443 -5163 489 -5117
rect 443 -5257 489 -5211
rect 443 -5351 489 -5305
rect 443 -5445 489 -5399
rect 443 -5539 489 -5493
rect 4485 -4787 4531 -4741
rect 4485 -4881 4531 -4835
rect 4485 -4975 4531 -4929
rect 4485 -5069 4531 -5023
rect 4485 -5163 4531 -5117
rect 4485 -5257 4531 -5211
rect 4485 -5351 4531 -5305
rect 4485 -5445 4531 -5399
rect 443 -5633 489 -5587
rect 443 -5727 489 -5681
rect 443 -5821 489 -5775
rect 443 -5915 489 -5869
rect 443 -6009 489 -5963
rect 4485 -5539 4531 -5493
rect 4485 -5633 4531 -5587
rect 4485 -5727 4531 -5681
rect 4485 -5821 4531 -5775
rect 4485 -5915 4531 -5869
rect 443 -6103 489 -6057
rect 443 -6197 489 -6151
rect 443 -6291 489 -6245
rect 443 -6385 489 -6339
rect 443 -6479 489 -6433
rect 443 -6573 489 -6527
rect 443 -6667 489 -6621
rect 443 -6761 489 -6715
rect 4485 -6009 4531 -5963
rect 4485 -6103 4531 -6057
rect 4485 -6197 4531 -6151
rect 4485 -6291 4531 -6245
rect 17720 -3502 17766 -3456
rect 17814 -3502 17860 -3456
rect 17908 -3502 17954 -3456
rect 18002 -3502 18048 -3456
rect 18096 -3502 18142 -3456
rect 18190 -3502 18236 -3456
rect 18284 -3502 18330 -3456
rect 18378 -3502 18424 -3456
rect 18472 -3502 18518 -3456
rect 18566 -3502 18612 -3456
rect 18660 -3502 18706 -3456
rect 18754 -3502 18800 -3456
rect 18848 -3502 18894 -3456
rect 18942 -3502 18988 -3456
rect 19036 -3502 19082 -3456
rect 19130 -3502 19176 -3456
rect 19224 -3502 19270 -3456
rect 19318 -3502 19364 -3456
rect 19412 -3502 19458 -3456
rect 19506 -3502 19552 -3456
rect 19600 -3502 19646 -3456
rect 19694 -3502 19740 -3456
rect 19788 -3502 19834 -3456
rect 19882 -3502 19928 -3456
rect 19976 -3502 20022 -3456
rect 20070 -3502 20116 -3456
rect 20164 -3502 20210 -3456
rect 20258 -3502 20304 -3456
rect 20352 -3502 20398 -3456
rect 20446 -3502 20492 -3456
rect 20540 -3502 20586 -3456
rect 20634 -3502 20680 -3456
rect 20728 -3502 20774 -3456
rect 20822 -3502 20868 -3456
rect 20916 -3502 20962 -3456
rect 21010 -3502 21056 -3456
rect 21104 -3502 21150 -3456
rect 21198 -3502 21244 -3456
rect 21292 -3502 21338 -3456
rect 21386 -3502 21432 -3456
rect 21480 -3502 21526 -3456
rect 21574 -3502 21620 -3456
rect 21668 -3502 21714 -3456
rect 21762 -3502 21808 -3456
rect 21856 -3502 21902 -3456
rect 21950 -3502 21996 -3456
rect 22044 -3502 22090 -3456
rect 22138 -3502 22184 -3456
rect 22232 -3502 22278 -3456
rect 22326 -3502 22372 -3456
rect 22420 -3502 22466 -3456
rect 22514 -3502 22560 -3456
rect 22608 -3502 22654 -3456
rect 22702 -3502 22748 -3456
rect 22796 -3502 22842 -3456
rect 22890 -3502 22936 -3456
rect 22984 -3502 23030 -3456
rect 23078 -3502 23124 -3456
rect 23172 -3502 23218 -3456
rect 23266 -3502 23312 -3456
rect 23360 -3502 23406 -3456
rect 23454 -3502 23500 -3456
rect 23548 -3502 23594 -3456
rect 23642 -3502 23688 -3456
rect 23736 -3502 23782 -3456
rect 23830 -3502 23876 -3456
rect 23924 -3502 23970 -3456
rect 24018 -3502 24064 -3456
rect 24112 -3502 24158 -3456
rect 24206 -3502 24252 -3456
rect 24300 -3502 24346 -3456
rect 24394 -3502 24440 -3456
rect 24488 -3502 24534 -3456
rect 24582 -3502 24628 -3456
rect 24676 -3502 24722 -3456
rect 24770 -3502 24816 -3456
rect 24864 -3502 24910 -3456
rect 24958 -3502 25004 -3456
rect 25052 -3502 25098 -3456
rect 25146 -3502 25192 -3456
rect 25240 -3502 25286 -3456
rect 25334 -3502 25380 -3456
rect 25428 -3502 25474 -3456
rect 25522 -3502 25568 -3456
rect 25616 -3502 25662 -3456
rect 25710 -3502 25756 -3456
rect 25804 -3502 25850 -3456
rect 25898 -3502 25944 -3456
rect 25992 -3502 26038 -3456
rect 26086 -3502 26132 -3456
rect 26180 -3502 26226 -3456
rect 26274 -3502 26320 -3456
rect 26368 -3502 26414 -3456
rect 26462 -3502 26508 -3456
rect 26556 -3502 26602 -3456
rect 26650 -3502 26696 -3456
rect 26744 -3502 26790 -3456
rect 26838 -3502 26884 -3456
rect 26932 -3502 26978 -3456
rect 27026 -3502 27072 -3456
rect 27120 -3502 27166 -3456
rect 27214 -3502 27260 -3456
rect 27308 -3502 27354 -3456
rect 27402 -3502 27448 -3456
rect 27496 -3502 27542 -3456
rect 27590 -3502 27636 -3456
rect 27684 -3502 27730 -3456
rect 27778 -3502 27824 -3456
rect 27872 -3502 27918 -3456
rect 27966 -3502 28012 -3456
rect 28060 -3502 28106 -3456
rect 28154 -3502 28200 -3456
rect 28248 -3502 28294 -3456
rect 28342 -3502 28388 -3456
rect 28436 -3502 28482 -3456
rect 28530 -3502 28576 -3456
rect 28624 -3502 28670 -3456
rect 28718 -3502 28764 -3456
rect 28812 -3502 28858 -3456
rect 28906 -3502 28952 -3456
rect 29000 -3502 29046 -3456
rect 29094 -3502 29140 -3456
rect 29188 -3502 29234 -3456
rect 29282 -3502 29328 -3456
rect 29376 -3502 29422 -3456
rect 29470 -3502 29516 -3456
rect 29564 -3502 29610 -3456
rect 29658 -3502 29704 -3456
rect 29752 -3502 29798 -3456
rect 29846 -3502 29892 -3456
rect 29940 -3502 29986 -3456
rect 30034 -3502 30080 -3456
rect 30128 -3502 30174 -3456
rect 30222 -3502 30268 -3456
rect 30316 -3502 30362 -3456
rect 30410 -3502 30456 -3456
rect 30504 -3502 30550 -3456
rect 30598 -3502 30644 -3456
rect 30692 -3502 30738 -3456
rect 30786 -3502 30832 -3456
rect 30880 -3502 30926 -3456
rect 30974 -3502 31020 -3456
rect 31068 -3502 31114 -3456
rect 31162 -3502 31208 -3456
rect 31256 -3502 31302 -3456
rect 17720 -3596 17766 -3550
rect 17720 -3690 17766 -3644
rect 17720 -3784 17766 -3738
rect 17720 -3878 17766 -3832
rect 17720 -3972 17766 -3926
rect 17720 -4066 17766 -4020
rect 17720 -4160 17766 -4114
rect 17720 -4254 17766 -4208
rect 22514 -3596 22560 -3550
rect 22514 -3690 22560 -3644
rect 22514 -3784 22560 -3738
rect 22514 -3878 22560 -3832
rect 22514 -3972 22560 -3926
rect 22514 -4066 22560 -4020
rect 22514 -4160 22560 -4114
rect 17720 -4348 17766 -4302
rect 22514 -4254 22560 -4208
rect 22514 -4348 22560 -4302
rect 17720 -4442 17766 -4396
rect 17720 -4536 17766 -4490
rect 17720 -4630 17766 -4584
rect 4485 -6385 4531 -6339
rect 4485 -6479 4531 -6433
rect 4485 -6573 4531 -6527
rect 4485 -6667 4531 -6621
rect 4485 -6761 4531 -6715
rect 443 -6855 489 -6809
rect 443 -6949 489 -6903
rect 443 -7043 489 -6997
rect 443 -7137 489 -7091
rect 443 -7231 489 -7185
rect 4485 -6855 4531 -6809
rect 4485 -6949 4531 -6903
rect 4485 -7043 4531 -6997
rect 4485 -7137 4531 -7091
rect 4485 -7231 4531 -7185
rect 443 -7325 489 -7279
rect 443 -7419 489 -7373
rect 4485 -7325 4531 -7279
rect 4485 -7419 4531 -7373
rect 443 -7513 489 -7467
rect 443 -7607 489 -7561
rect 4485 -7513 4531 -7467
rect 4485 -7607 4531 -7561
rect 443 -7701 489 -7655
rect 537 -7701 583 -7655
rect 631 -7701 677 -7655
rect 725 -7701 771 -7655
rect 819 -7701 865 -7655
rect 913 -7701 959 -7655
rect 1007 -7701 1053 -7655
rect 1101 -7701 1147 -7655
rect 1195 -7701 1241 -7655
rect 1289 -7701 1335 -7655
rect 1383 -7701 1429 -7655
rect 1477 -7701 1523 -7655
rect 1571 -7701 1617 -7655
rect 1665 -7701 1711 -7655
rect 1759 -7701 1805 -7655
rect 1853 -7701 1899 -7655
rect 1947 -7701 1993 -7655
rect 2041 -7701 2087 -7655
rect 2135 -7701 2181 -7655
rect 2229 -7701 2275 -7655
rect 2323 -7701 2369 -7655
rect 2417 -7701 2463 -7655
rect 2511 -7701 2557 -7655
rect 2605 -7701 2651 -7655
rect 2699 -7701 2745 -7655
rect 2793 -7701 2839 -7655
rect 2887 -7701 2933 -7655
rect 2981 -7701 3027 -7655
rect 3075 -7701 3121 -7655
rect 3169 -7701 3215 -7655
rect 3263 -7701 3309 -7655
rect 3357 -7701 3403 -7655
rect 3451 -7701 3497 -7655
rect 3545 -7701 3591 -7655
rect 3639 -7701 3685 -7655
rect 3733 -7701 3779 -7655
rect 3827 -7701 3873 -7655
rect 3921 -7701 3967 -7655
rect 4015 -7701 4061 -7655
rect 4109 -7701 4155 -7655
rect 4203 -7701 4249 -7655
rect 4297 -7701 4343 -7655
rect 4391 -7701 4437 -7655
rect 4485 -7701 4531 -7655
rect 17720 -4724 17766 -4678
rect 17720 -4818 17766 -4772
rect 17720 -4912 17766 -4866
rect 17720 -5006 17766 -4960
rect 22514 -4442 22560 -4396
rect 22514 -4536 22560 -4490
rect 22514 -4630 22560 -4584
rect 22514 -4724 22560 -4678
rect 22514 -4818 22560 -4772
rect 22514 -4912 22560 -4866
rect 17720 -5100 17766 -5054
rect 17720 -5194 17766 -5148
rect 17720 -5288 17766 -5242
rect 17720 -5382 17766 -5336
rect 17720 -5476 17766 -5430
rect 17720 -5570 17766 -5524
rect 17720 -5664 17766 -5618
rect 17720 -5758 17766 -5712
rect 17720 -5852 17766 -5806
rect 17720 -5946 17766 -5900
rect 17720 -6040 17766 -5994
rect 17720 -6134 17766 -6088
rect 17720 -6228 17766 -6182
rect 17720 -6322 17766 -6276
rect 17720 -6416 17766 -6370
rect 17720 -6510 17766 -6464
rect 17720 -6604 17766 -6558
rect 22514 -5006 22560 -4960
rect 17720 -6698 17766 -6652
rect 22514 -5100 22560 -5054
rect 22514 -5194 22560 -5148
rect 22514 -5288 22560 -5242
rect 22514 -5382 22560 -5336
rect 22514 -5476 22560 -5430
rect 22514 -5570 22560 -5524
rect 22514 -5664 22560 -5618
rect 22514 -5758 22560 -5712
rect 22514 -5852 22560 -5806
rect 22514 -5946 22560 -5900
rect 22514 -6040 22560 -5994
rect 22514 -6134 22560 -6088
rect 22514 -6228 22560 -6182
rect 22514 -6322 22560 -6276
rect 22514 -6416 22560 -6370
rect 22514 -6510 22560 -6464
rect 22514 -6604 22560 -6558
rect 17720 -6792 17766 -6746
rect 17720 -6886 17766 -6840
rect 17720 -6980 17766 -6934
rect 17720 -7074 17766 -7028
rect 17720 -7168 17766 -7122
rect 22514 -6698 22560 -6652
rect 22514 -6792 22560 -6746
rect 22514 -6886 22560 -6840
rect 22514 -6980 22560 -6934
rect 22514 -7074 22560 -7028
rect 22514 -7168 22560 -7122
rect 17720 -7262 17766 -7216
rect 17720 -7356 17766 -7310
rect 22514 -7262 22560 -7216
rect 17720 -7450 17766 -7404
rect 17720 -7544 17766 -7498
rect 17720 -7638 17766 -7592
rect 17720 -7732 17766 -7686
rect 17720 -7826 17766 -7780
rect 17720 -7920 17766 -7874
rect 17720 -8014 17766 -7968
rect 22514 -7356 22560 -7310
rect 22514 -7450 22560 -7404
rect 22514 -7544 22560 -7498
rect 22514 -7638 22560 -7592
rect 22514 -7732 22560 -7686
rect 22514 -7826 22560 -7780
rect 22514 -7920 22560 -7874
rect 22514 -8014 22560 -7968
rect 28248 -3596 28294 -3550
rect 28248 -3690 28294 -3644
rect 28248 -3784 28294 -3738
rect 28248 -3878 28294 -3832
rect 28248 -3972 28294 -3926
rect 28248 -4066 28294 -4020
rect 28248 -4160 28294 -4114
rect 28248 -4254 28294 -4208
rect 28248 -4348 28294 -4302
rect 28248 -4442 28294 -4396
rect 28248 -4536 28294 -4490
rect 28248 -4630 28294 -4584
rect 28248 -4724 28294 -4678
rect 28248 -4818 28294 -4772
rect 28248 -4912 28294 -4866
rect 28248 -5006 28294 -4960
rect 28248 -5100 28294 -5054
rect 28248 -5194 28294 -5148
rect 28248 -5288 28294 -5242
rect 28248 -5382 28294 -5336
rect 28248 -5476 28294 -5430
rect 28248 -5570 28294 -5524
rect 28248 -5664 28294 -5618
rect 28248 -5758 28294 -5712
rect 28248 -5852 28294 -5806
rect 28248 -5946 28294 -5900
rect 28248 -6040 28294 -5994
rect 28248 -6134 28294 -6088
rect 28248 -6228 28294 -6182
rect 28248 -6322 28294 -6276
rect 28248 -6416 28294 -6370
rect 28248 -6510 28294 -6464
rect 28248 -6604 28294 -6558
rect 28248 -6698 28294 -6652
rect 28248 -6792 28294 -6746
rect 28248 -6886 28294 -6840
rect 28248 -6980 28294 -6934
rect 28248 -7074 28294 -7028
rect 28248 -7168 28294 -7122
rect 28248 -7262 28294 -7216
rect 28248 -7356 28294 -7310
rect 28248 -7450 28294 -7404
rect 28248 -7544 28294 -7498
rect 28248 -7638 28294 -7592
rect 28248 -7732 28294 -7686
rect 28248 -7826 28294 -7780
rect 28248 -7920 28294 -7874
rect 28248 -8014 28294 -7968
rect 31256 -3596 31302 -3550
rect 31256 -3690 31302 -3644
rect 31256 -3784 31302 -3738
rect 31256 -3878 31302 -3832
rect 31256 -3972 31302 -3926
rect 31256 -4066 31302 -4020
rect 31256 -4160 31302 -4114
rect 31256 -4254 31302 -4208
rect 31256 -4348 31302 -4302
rect 31256 -4442 31302 -4396
rect 31256 -4536 31302 -4490
rect 31256 -4630 31302 -4584
rect 31256 -4724 31302 -4678
rect 31256 -4818 31302 -4772
rect 31256 -4912 31302 -4866
rect 31256 -5006 31302 -4960
rect 31256 -5100 31302 -5054
rect 31256 -5194 31302 -5148
rect 31256 -5288 31302 -5242
rect 31256 -5382 31302 -5336
rect 31256 -5476 31302 -5430
rect 31256 -5570 31302 -5524
rect 31256 -5664 31302 -5618
rect 31256 -5758 31302 -5712
rect 31256 -5852 31302 -5806
rect 31256 -5946 31302 -5900
rect 31256 -6040 31302 -5994
rect 31256 -6134 31302 -6088
rect 31256 -6228 31302 -6182
rect 31256 -6322 31302 -6276
rect 31256 -6416 31302 -6370
rect 31256 -6510 31302 -6464
rect 31256 -6604 31302 -6558
rect 31256 -6698 31302 -6652
rect 31256 -6792 31302 -6746
rect 31256 -6886 31302 -6840
rect 31256 -6980 31302 -6934
rect 31256 -7074 31302 -7028
rect 31256 -7168 31302 -7122
rect 31256 -7262 31302 -7216
rect 31256 -7356 31302 -7310
rect 31256 -7450 31302 -7404
rect 31256 -7544 31302 -7498
rect 31256 -7638 31302 -7592
rect 31256 -7732 31302 -7686
rect 31256 -7826 31302 -7780
rect 31256 -7920 31302 -7874
rect 31256 -8014 31302 -7968
rect 17720 -8108 17766 -8062
rect 17814 -8108 17860 -8062
rect 17908 -8108 17954 -8062
rect 18002 -8108 18048 -8062
rect 18096 -8108 18142 -8062
rect 18190 -8108 18236 -8062
rect 18284 -8108 18330 -8062
rect 18378 -8108 18424 -8062
rect 18472 -8108 18518 -8062
rect 18566 -8108 18612 -8062
rect 18660 -8108 18706 -8062
rect 18754 -8108 18800 -8062
rect 18848 -8108 18894 -8062
rect 18942 -8108 18988 -8062
rect 19036 -8108 19082 -8062
rect 19130 -8108 19176 -8062
rect 19224 -8108 19270 -8062
rect 19318 -8108 19364 -8062
rect 19412 -8108 19458 -8062
rect 19506 -8108 19552 -8062
rect 19600 -8108 19646 -8062
rect 19694 -8108 19740 -8062
rect 19788 -8108 19834 -8062
rect 19882 -8108 19928 -8062
rect 19976 -8108 20022 -8062
rect 20070 -8108 20116 -8062
rect 20164 -8108 20210 -8062
rect 20258 -8108 20304 -8062
rect 20352 -8108 20398 -8062
rect 20446 -8108 20492 -8062
rect 20540 -8108 20586 -8062
rect 20634 -8108 20680 -8062
rect 20728 -8108 20774 -8062
rect 20822 -8108 20868 -8062
rect 20916 -8108 20962 -8062
rect 21010 -8108 21056 -8062
rect 21104 -8108 21150 -8062
rect 21198 -8108 21244 -8062
rect 21292 -8108 21338 -8062
rect 21386 -8108 21432 -8062
rect 21480 -8108 21526 -8062
rect 21574 -8108 21620 -8062
rect 21668 -8108 21714 -8062
rect 21762 -8108 21808 -8062
rect 21856 -8108 21902 -8062
rect 21950 -8108 21996 -8062
rect 22044 -8108 22090 -8062
rect 22138 -8108 22184 -8062
rect 22232 -8108 22278 -8062
rect 22326 -8108 22372 -8062
rect 22420 -8108 22466 -8062
rect 22514 -8108 22560 -8062
rect 22608 -8108 22654 -8062
rect 22702 -8108 22748 -8062
rect 22796 -8108 22842 -8062
rect 22890 -8108 22936 -8062
rect 22984 -8108 23030 -8062
rect 23078 -8108 23124 -8062
rect 23172 -8108 23218 -8062
rect 23266 -8108 23312 -8062
rect 23360 -8108 23406 -8062
rect 23454 -8108 23500 -8062
rect 23548 -8108 23594 -8062
rect 23642 -8108 23688 -8062
rect 23736 -8108 23782 -8062
rect 23830 -8108 23876 -8062
rect 23924 -8108 23970 -8062
rect 24018 -8108 24064 -8062
rect 24112 -8108 24158 -8062
rect 24206 -8108 24252 -8062
rect 24300 -8108 24346 -8062
rect 24394 -8108 24440 -8062
rect 24488 -8108 24534 -8062
rect 24582 -8108 24628 -8062
rect 24676 -8108 24722 -8062
rect 24770 -8108 24816 -8062
rect 24864 -8108 24910 -8062
rect 24958 -8108 25004 -8062
rect 25052 -8108 25098 -8062
rect 25146 -8108 25192 -8062
rect 25240 -8108 25286 -8062
rect 25334 -8108 25380 -8062
rect 25428 -8108 25474 -8062
rect 25522 -8108 25568 -8062
rect 25616 -8108 25662 -8062
rect 25710 -8108 25756 -8062
rect 25804 -8108 25850 -8062
rect 25898 -8108 25944 -8062
rect 25992 -8108 26038 -8062
rect 26086 -8108 26132 -8062
rect 26180 -8108 26226 -8062
rect 26274 -8108 26320 -8062
rect 26368 -8108 26414 -8062
rect 26462 -8108 26508 -8062
rect 26556 -8108 26602 -8062
rect 26650 -8108 26696 -8062
rect 26744 -8108 26790 -8062
rect 26838 -8108 26884 -8062
rect 26932 -8108 26978 -8062
rect 27026 -8108 27072 -8062
rect 27120 -8108 27166 -8062
rect 27214 -8108 27260 -8062
rect 27308 -8108 27354 -8062
rect 27402 -8108 27448 -8062
rect 27496 -8108 27542 -8062
rect 27590 -8108 27636 -8062
rect 27684 -8108 27730 -8062
rect 27778 -8108 27824 -8062
rect 27872 -8108 27918 -8062
rect 27966 -8108 28012 -8062
rect 28060 -8108 28106 -8062
rect 28154 -8108 28200 -8062
rect 28248 -8108 28294 -8062
rect 28342 -8108 28388 -8062
rect 28436 -8108 28482 -8062
rect 28530 -8108 28576 -8062
rect 28624 -8108 28670 -8062
rect 28718 -8108 28764 -8062
rect 28812 -8108 28858 -8062
rect 28906 -8108 28952 -8062
rect 29000 -8108 29046 -8062
rect 29094 -8108 29140 -8062
rect 29188 -8108 29234 -8062
rect 29282 -8108 29328 -8062
rect 29376 -8108 29422 -8062
rect 29470 -8108 29516 -8062
rect 29564 -8108 29610 -8062
rect 29658 -8108 29704 -8062
rect 29752 -8108 29798 -8062
rect 29846 -8108 29892 -8062
rect 29940 -8108 29986 -8062
rect 30034 -8108 30080 -8062
rect 30128 -8108 30174 -8062
rect 30222 -8108 30268 -8062
rect 30316 -8108 30362 -8062
rect 30410 -8108 30456 -8062
rect 30504 -8108 30550 -8062
rect 30598 -8108 30644 -8062
rect 30692 -8108 30738 -8062
rect 30786 -8108 30832 -8062
rect 30880 -8108 30926 -8062
rect 30974 -8108 31020 -8062
rect 31068 -8108 31114 -8062
rect 31162 -8108 31208 -8062
rect 31256 -8108 31302 -8062
<< polysilicon >>
rect 3466 5062 3538 5075
rect 3466 5016 3479 5062
rect 3525 5016 3538 5062
rect 3466 5003 3538 5016
rect 3946 5062 4018 5075
rect 3946 5016 3959 5062
rect 4005 5016 4018 5062
rect 3946 5003 4018 5016
rect 4586 5062 4658 5075
rect 4586 5016 4599 5062
rect 4645 5016 4658 5062
rect 4586 5003 4658 5016
rect 3474 4869 3530 5003
rect 3954 4945 4010 5003
rect 3954 4889 4170 4945
rect 3954 4869 4010 4889
rect 4594 4869 4650 5003
rect 3186 3739 3242 4119
rect 3634 4099 3690 4119
rect 4274 4099 4330 4119
rect 3634 4043 3850 4099
rect 4274 4043 4490 4099
rect 3634 3947 3690 4043
rect 4274 3947 4330 4043
rect 3466 3934 3538 3947
rect 3466 3888 3479 3934
rect 3525 3888 3538 3934
rect 3466 3875 3538 3888
rect 3626 3934 3698 3947
rect 3626 3888 3639 3934
rect 3685 3888 3698 3934
rect 3626 3875 3698 3888
rect 3946 3934 4018 3947
rect 3946 3888 3959 3934
rect 4005 3888 4018 3934
rect 3946 3875 4018 3888
rect 4266 3934 4338 3947
rect 4266 3888 4279 3934
rect 4325 3888 4338 3934
rect 4266 3875 4338 3888
rect 4586 3934 4658 3947
rect 4586 3888 4599 3934
rect 4645 3888 4658 3934
rect 4586 3875 4658 3888
rect 3474 3739 3530 3875
rect 3954 3815 4010 3875
rect 3954 3759 4170 3815
rect 3954 3739 4010 3759
rect 4594 3739 4650 3875
rect 4882 3739 4938 4119
rect 3186 2609 3242 2989
rect 3634 2913 3850 2969
rect 4274 2913 4490 2969
rect 3634 2819 3690 2913
rect 4274 2819 4330 2913
rect 3466 2806 3538 2819
rect 3466 2760 3479 2806
rect 3525 2760 3538 2806
rect 3466 2745 3538 2760
rect 3626 2806 3698 2819
rect 3626 2760 3639 2806
rect 3685 2760 3698 2806
rect 3626 2747 3698 2760
rect 3946 2806 4018 2819
rect 3946 2760 3959 2806
rect 4005 2760 4018 2806
rect 3946 2745 4018 2760
rect 4266 2806 4338 2819
rect 4266 2760 4279 2806
rect 4325 2760 4338 2806
rect 4266 2747 4338 2760
rect 4586 2806 4658 2819
rect 4586 2760 4599 2806
rect 4645 2760 4658 2806
rect 4586 2745 4658 2760
rect 3474 2609 3530 2745
rect 3954 2685 4010 2745
rect 3954 2629 4170 2685
rect 3954 2609 4010 2629
rect 4594 2609 4650 2745
rect 4882 2609 4938 2989
rect 3186 1479 3242 1859
rect 3474 1479 3530 1859
rect 3634 1479 3690 1859
rect 3794 1479 3850 1859
rect 3954 1479 4010 1859
rect 4114 1479 4170 1859
rect 4274 1479 4330 1859
rect 4434 1479 4490 1859
rect 4594 1479 4650 1859
rect 4882 1479 4938 1859
rect 500 639 612 775
rect 716 639 828 775
rect 932 639 1044 775
rect 1148 639 1260 775
rect 1364 639 1476 775
rect 1580 639 1692 775
rect 1796 639 1908 775
rect 2012 639 2124 775
rect 2228 639 2340 775
rect 2444 639 2556 775
rect 3186 349 3242 729
rect 3634 709 3690 729
rect 4274 709 4330 729
rect 3634 653 3850 709
rect 4274 653 4490 709
rect 3634 559 3690 653
rect 4274 559 4330 653
rect 3466 546 3538 559
rect 3466 500 3479 546
rect 3525 500 3538 546
rect 3466 485 3538 500
rect 3626 546 3698 559
rect 3626 500 3639 546
rect 3685 500 3698 546
rect 3626 487 3698 500
rect 3946 546 4018 559
rect 3946 500 3959 546
rect 4005 500 4018 546
rect 3946 485 4018 500
rect 4266 546 4338 559
rect 4266 500 4279 546
rect 4325 500 4338 546
rect 4266 487 4338 500
rect 4586 546 4658 559
rect 4586 500 4599 546
rect 4645 500 4658 546
rect 4586 485 4658 500
rect 3474 349 3530 485
rect 3954 425 4010 485
rect 3954 369 4170 425
rect 3954 349 4010 369
rect 4594 349 4650 485
rect 4882 349 4938 729
rect 500 -123 612 13
rect 716 -123 828 13
rect 932 -123 1044 13
rect 1148 -123 1260 13
rect 1364 -123 1476 13
rect 1580 -123 1692 13
rect 1796 -123 1908 13
rect 2012 -123 2124 13
rect 2228 -123 2340 13
rect 2444 -123 2556 13
rect 3186 -555 3242 -401
rect 3634 -421 3690 -401
rect 4274 -421 4330 -401
rect 4434 -421 4490 -401
rect 3634 -477 3850 -421
rect 4274 -477 4490 -421
rect 3178 -568 3250 -555
rect 3178 -614 3191 -568
rect 3237 -614 3250 -568
rect 3634 -571 3690 -477
rect 4274 -571 4330 -477
rect 4882 -555 4938 -401
rect 4874 -568 4946 -555
rect 3178 -627 3250 -614
rect 3466 -584 3538 -571
rect 500 -794 612 -749
rect 500 -840 533 -794
rect 579 -840 612 -794
rect 500 -885 612 -840
rect 716 -885 828 -749
rect 932 -885 1044 -749
rect 1148 -885 1260 -749
rect 1364 -885 1476 -749
rect 1580 -885 1692 -749
rect 1796 -885 1908 -749
rect 2012 -885 2124 -749
rect 2228 -885 2340 -749
rect 2444 -794 2556 -749
rect 2444 -840 2477 -794
rect 2523 -840 2556 -794
rect 2444 -885 2556 -840
rect 3186 -781 3242 -627
rect 3466 -630 3479 -584
rect 3525 -630 3538 -584
rect 3466 -643 3538 -630
rect 3626 -584 3698 -571
rect 3626 -630 3639 -584
rect 3685 -630 3698 -584
rect 3626 -643 3698 -630
rect 3946 -584 4018 -571
rect 3946 -630 3959 -584
rect 4005 -630 4018 -584
rect 3474 -781 3530 -643
rect 3946 -645 4018 -630
rect 4266 -584 4338 -571
rect 4266 -630 4279 -584
rect 4325 -630 4338 -584
rect 4266 -643 4338 -630
rect 4586 -584 4658 -571
rect 4586 -630 4599 -584
rect 4645 -630 4658 -584
rect 4874 -614 4887 -568
rect 4933 -614 4946 -568
rect 4874 -627 4946 -614
rect 4586 -643 4658 -630
rect 3954 -705 4010 -645
rect 3954 -761 4170 -705
rect 3954 -781 4010 -761
rect 4114 -781 4170 -761
rect 4594 -781 4650 -643
rect 4882 -781 4938 -627
rect 716 -1531 828 -1511
rect 716 -1577 2340 -1531
rect 716 -1623 756 -1577
rect 802 -1623 860 -1577
rect 906 -1623 2340 -1577
rect 716 -1643 2340 -1623
rect 3634 -1551 3690 -1531
rect 4274 -1551 4330 -1531
rect 3634 -1607 3850 -1551
rect 4274 -1607 4490 -1551
rect 3634 -1655 3690 -1607
rect 4274 -1655 4330 -1607
rect 3626 -1668 3698 -1655
rect 3626 -1714 3639 -1668
rect 3685 -1714 3698 -1668
rect 3626 -1727 3698 -1714
rect 4266 -1668 4338 -1655
rect 4266 -1714 4279 -1668
rect 4325 -1714 4338 -1668
rect 4266 -1727 4338 -1714
rect 6051 4257 6107 4543
rect 6339 4484 6395 4543
rect 6499 4484 6555 4543
rect 6659 4484 6715 4543
rect 6819 4484 6875 4543
rect 6979 4484 7035 4543
rect 7139 4484 7195 4543
rect 7299 4484 7355 4543
rect 7459 4484 7515 4543
rect 6339 4364 7515 4484
rect 6339 4257 6395 4364
rect 6499 4257 6555 4364
rect 6659 4257 6715 4364
rect 6819 4321 7515 4364
rect 6819 4257 6875 4321
rect 6979 4257 7035 4321
rect 7139 4257 7195 4321
rect 7299 4257 7355 4321
rect 7459 4257 7515 4321
rect 7747 4257 7803 4543
rect 6051 3395 6107 3681
rect 6339 3620 6395 3681
rect 6499 3620 6555 3681
rect 6659 3620 6715 3681
rect 6819 3620 6875 3681
rect 6979 3620 7035 3681
rect 7139 3620 7195 3681
rect 7299 3620 7355 3681
rect 7459 3620 7515 3681
rect 6339 3500 7515 3620
rect 6339 3395 6395 3500
rect 6499 3395 6555 3500
rect 6659 3395 6715 3500
rect 6819 3395 6875 3500
rect 6979 3395 7035 3500
rect 7139 3395 7195 3500
rect 7299 3395 7355 3500
rect 7459 3395 7515 3500
rect 7747 3395 7803 3681
rect 6051 2533 6107 2819
rect 6339 2750 6395 2819
rect 6499 2750 6555 2819
rect 6659 2750 6715 2819
rect 6819 2750 6875 2819
rect 6979 2750 7035 2819
rect 7139 2750 7195 2819
rect 7299 2750 7355 2819
rect 7459 2750 7515 2819
rect 6339 2630 7515 2750
rect 6339 2533 6395 2630
rect 6499 2533 6555 2630
rect 6659 2533 6715 2630
rect 6819 2533 6875 2630
rect 6979 2533 7035 2630
rect 7139 2533 7195 2630
rect 7299 2533 7355 2630
rect 7459 2533 7515 2630
rect 7747 2533 7803 2819
rect 18581 4245 18653 4258
rect 18581 4199 18594 4245
rect 18640 4199 18653 4245
rect 18581 4186 18653 4199
rect 19061 4245 19133 4258
rect 19061 4199 19074 4245
rect 19120 4199 19133 4245
rect 19061 4186 19133 4199
rect 19701 4245 19773 4258
rect 19701 4199 19714 4245
rect 19760 4199 19773 4245
rect 19701 4186 19773 4199
rect 18589 4032 18645 4186
rect 19069 4108 19125 4186
rect 19069 4052 19285 4108
rect 19069 4032 19125 4052
rect 19709 4032 19765 4186
rect 18301 3300 18357 3432
rect 18749 3412 18805 3432
rect 19389 3412 19445 3432
rect 18749 3356 18965 3412
rect 19389 3356 19605 3412
rect 18293 3287 18365 3300
rect 18749 3292 18805 3356
rect 19389 3292 19445 3356
rect 19997 3300 20053 3432
rect 18293 3241 18306 3287
rect 18352 3241 18365 3287
rect 18293 3228 18365 3241
rect 18581 3279 18653 3292
rect 18581 3233 18594 3279
rect 18640 3233 18653 3279
rect 6051 1671 6107 1957
rect 6339 1876 6395 1957
rect 6499 1876 6555 1957
rect 6659 1876 6715 1957
rect 6819 1876 6875 1957
rect 6979 1876 7035 1957
rect 7139 1876 7195 1957
rect 7299 1876 7355 1957
rect 7459 1876 7515 1957
rect 6339 1756 7515 1876
rect 6339 1671 6395 1756
rect 6499 1671 6555 1756
rect 6659 1671 6715 1756
rect 6819 1671 6875 1756
rect 6979 1671 7035 1756
rect 7139 1671 7195 1756
rect 7299 1671 7355 1756
rect 7459 1671 7515 1756
rect 7747 1671 7803 1957
rect 6051 809 6107 1095
rect 6339 1016 6395 1095
rect 6499 1016 6555 1095
rect 6659 1016 6715 1095
rect 6819 1016 6875 1095
rect 6979 1016 7035 1095
rect 7139 1016 7195 1095
rect 7299 1016 7355 1095
rect 7459 1016 7515 1095
rect 6339 896 7515 1016
rect 6339 809 6395 896
rect 6499 809 6555 896
rect 6659 809 6715 896
rect 6819 809 6875 896
rect 6979 809 7035 896
rect 7139 809 7195 896
rect 7299 809 7355 896
rect 7459 809 7515 896
rect 7747 809 7803 1095
rect 8286 790 8342 1076
rect 8574 978 8630 1076
rect 8862 978 8918 1076
rect 9022 978 9078 1076
rect 9310 978 9366 1076
rect 9470 978 9526 1076
rect 9758 978 9814 1076
rect 9918 978 9974 1076
rect 10206 978 10262 1076
rect 8574 858 10262 978
rect 8574 790 8630 858
rect 8862 790 8918 858
rect 9022 790 9078 858
rect 9310 790 9366 858
rect 9470 790 9526 858
rect 9758 790 9814 858
rect 9918 790 9974 858
rect 10206 790 10262 858
rect 10494 790 10550 1076
rect 6051 -53 6107 233
rect 6339 160 6395 233
rect 6499 160 6555 233
rect 6659 160 6715 233
rect 6819 160 6875 233
rect 6979 160 7035 233
rect 7139 160 7195 233
rect 7299 160 7355 233
rect 7459 160 7515 233
rect 6339 40 7515 160
rect 6339 -53 6395 40
rect 6499 -53 6555 40
rect 6659 -53 6715 40
rect 6819 -53 6875 40
rect 6979 -53 7035 40
rect 7139 -53 7195 40
rect 7299 -53 7355 40
rect 7459 -53 7515 40
rect 7747 -53 7803 233
rect 8286 -72 8342 214
rect 8574 116 8630 214
rect 8862 116 8918 214
rect 9022 116 9078 214
rect 9310 116 9366 214
rect 9470 116 9526 214
rect 9758 116 9814 214
rect 9918 116 9974 214
rect 10206 116 10262 214
rect 8574 -4 10262 116
rect 8574 -72 8630 -4
rect 8862 -72 8918 -4
rect 9022 -72 9078 -4
rect 9310 -72 9366 -4
rect 9470 -72 9526 -4
rect 9758 -72 9814 -4
rect 9918 -72 9974 -4
rect 10206 -72 10262 -4
rect 10494 -72 10550 214
rect 6051 -736 6107 -629
rect 6043 -749 6115 -736
rect 6043 -795 6056 -749
rect 6102 -795 6115 -749
rect 6043 -808 6115 -795
rect 6339 -741 6395 -629
rect 6499 -741 6555 -629
rect 6659 -741 6715 -629
rect 6819 -741 6875 -629
rect 6979 -741 7035 -629
rect 7139 -741 7195 -629
rect 7299 -741 7355 -629
rect 7459 -681 7515 -629
rect 7459 -683 7534 -681
rect 7459 -696 7577 -683
rect 7459 -741 7518 -696
rect 6339 -742 7518 -741
rect 7564 -742 7577 -696
rect 7747 -736 7803 -629
rect 6339 -800 7577 -742
rect 6051 -915 6107 -808
rect 6339 -846 7518 -800
rect 7564 -846 7577 -800
rect 7739 -749 7811 -736
rect 7739 -795 7752 -749
rect 7798 -795 7811 -749
rect 7739 -808 7811 -795
rect 8286 -755 8342 -648
rect 8574 -716 8630 -648
rect 8862 -716 8918 -648
rect 9022 -716 9078 -648
rect 9310 -716 9366 -648
rect 9470 -716 9526 -648
rect 9758 -716 9814 -648
rect 9918 -716 9974 -648
rect 10206 -694 10262 -648
rect 10206 -707 10310 -694
rect 10206 -716 10251 -707
rect 8574 -753 10251 -716
rect 10297 -753 10310 -707
rect 6339 -859 7577 -846
rect 6339 -861 7534 -859
rect 6339 -915 6395 -861
rect 6499 -915 6555 -861
rect 6659 -915 6715 -861
rect 6819 -915 6875 -861
rect 6979 -915 7035 -861
rect 7139 -915 7195 -861
rect 7299 -915 7355 -861
rect 7459 -915 7515 -861
rect 7747 -915 7803 -808
rect 8278 -768 8350 -755
rect 8278 -814 8291 -768
rect 8337 -814 8350 -768
rect 8278 -827 8350 -814
rect 8574 -811 10310 -753
rect 10494 -755 10550 -648
rect 8286 -934 8342 -827
rect 8574 -836 10251 -811
rect 8574 -934 8630 -836
rect 8862 -934 8918 -836
rect 9022 -934 9078 -836
rect 9310 -934 9366 -836
rect 9470 -934 9526 -836
rect 9758 -934 9814 -836
rect 9918 -934 9974 -836
rect 10206 -857 10251 -836
rect 10297 -857 10310 -811
rect 10486 -768 10558 -755
rect 10486 -814 10499 -768
rect 10545 -814 10558 -768
rect 10486 -827 10558 -814
rect 10206 -870 10310 -857
rect 10206 -934 10262 -870
rect 10494 -934 10550 -827
rect 11668 1184 11724 1594
rect 11956 1448 12012 1594
rect 12244 1448 12300 1594
rect 12404 1448 12460 1594
rect 12692 1448 12748 1594
rect 12852 1448 12908 1594
rect 13140 1448 13196 1594
rect 13300 1448 13356 1594
rect 13588 1448 13644 1594
rect 11956 1328 13644 1448
rect 11956 1184 12012 1328
rect 12244 1184 12300 1328
rect 12404 1184 12460 1328
rect 12692 1184 12748 1328
rect 12852 1184 12908 1328
rect 13140 1184 13196 1328
rect 13300 1184 13356 1328
rect 13588 1184 13644 1328
rect 13876 1184 13932 1594
rect 14462 1184 14518 1594
rect 14750 1433 14806 1594
rect 14910 1433 14966 1594
rect 15070 1433 15126 1594
rect 15230 1433 15286 1594
rect 15390 1433 15446 1594
rect 15550 1433 15606 1594
rect 15710 1433 15766 1594
rect 15870 1433 15926 1594
rect 14750 1313 15926 1433
rect 14750 1184 14806 1313
rect 14910 1184 14966 1313
rect 15070 1184 15126 1313
rect 15230 1184 15286 1313
rect 15390 1184 15446 1313
rect 15550 1184 15606 1313
rect 15710 1184 15766 1313
rect 15870 1184 15926 1313
rect 16158 1184 16214 1594
rect 11668 148 11724 558
rect 11956 398 12012 558
rect 12244 398 12300 558
rect 12404 398 12460 558
rect 12692 398 12748 558
rect 12852 398 12908 558
rect 13140 398 13196 558
rect 13300 398 13356 558
rect 13588 398 13644 558
rect 11956 278 13644 398
rect 11956 148 12012 278
rect 12244 148 12300 278
rect 12404 148 12460 278
rect 12692 148 12748 278
rect 12852 148 12908 278
rect 13140 148 13196 278
rect 13300 148 13356 278
rect 13588 148 13644 278
rect 13876 148 13932 558
rect 14462 148 14518 558
rect 14750 406 14806 558
rect 14910 406 14966 558
rect 15070 406 15126 558
rect 15230 406 15286 558
rect 15390 406 15446 558
rect 15550 406 15606 558
rect 15710 406 15766 558
rect 15870 406 15926 558
rect 14750 286 15926 406
rect 14750 148 14806 286
rect 14910 148 14966 286
rect 15070 148 15126 286
rect 15230 148 15286 286
rect 15390 148 15446 286
rect 15550 148 15606 286
rect 15710 148 15766 286
rect 15870 148 15926 286
rect 16158 148 16214 558
rect 11668 -709 11724 -478
rect 11956 -582 12012 -478
rect 11902 -597 12012 -582
rect 11902 -643 11917 -597
rect 11963 -642 12012 -597
rect 12244 -642 12300 -478
rect 12404 -642 12460 -478
rect 12692 -642 12748 -478
rect 12852 -642 12908 -478
rect 13140 -642 13196 -478
rect 13300 -642 13356 -478
rect 13588 -642 13644 -478
rect 11963 -643 13644 -642
rect 11902 -701 13644 -643
rect 11660 -722 11732 -709
rect 11660 -768 11673 -722
rect 11719 -768 11732 -722
rect 11902 -747 11917 -701
rect 11963 -747 13644 -701
rect 13876 -709 13932 -478
rect 11902 -762 13644 -747
rect 11660 -781 11732 -768
rect 11668 -888 11724 -781
rect 11956 -888 12012 -762
rect 12244 -888 12300 -762
rect 12404 -888 12460 -762
rect 12692 -888 12748 -762
rect 12852 -888 12908 -762
rect 13140 -888 13196 -762
rect 13300 -888 13356 -762
rect 13588 -888 13644 -762
rect 13868 -722 13940 -709
rect 13868 -768 13881 -722
rect 13927 -768 13940 -722
rect 13868 -781 13940 -768
rect 14462 -709 14518 -478
rect 14750 -577 14806 -478
rect 14688 -592 14806 -577
rect 14688 -638 14703 -592
rect 14749 -637 14806 -592
rect 14910 -637 14966 -478
rect 15070 -637 15126 -478
rect 15230 -637 15286 -478
rect 15390 -637 15446 -478
rect 15550 -637 15606 -478
rect 15710 -637 15766 -478
rect 15870 -637 15926 -478
rect 14749 -638 15926 -637
rect 14688 -696 15926 -638
rect 13876 -888 13932 -781
rect 14454 -722 14526 -709
rect 14454 -768 14467 -722
rect 14513 -768 14526 -722
rect 14688 -742 14703 -696
rect 14749 -742 15926 -696
rect 16158 -709 16214 -478
rect 14688 -757 15926 -742
rect 14454 -781 14526 -768
rect 14462 -888 14518 -781
rect 14750 -888 14806 -757
rect 14910 -888 14966 -757
rect 15070 -888 15126 -757
rect 15230 -888 15286 -757
rect 15390 -888 15446 -757
rect 15550 -888 15606 -757
rect 15710 -888 15766 -757
rect 15870 -888 15926 -757
rect 16150 -722 16222 -709
rect 16150 -768 16163 -722
rect 16209 -768 16222 -722
rect 16150 -781 16222 -768
rect 16158 -888 16214 -781
rect 18301 -444 18357 3228
rect 18581 3220 18653 3233
rect 18741 3279 18813 3292
rect 18741 3233 18754 3279
rect 18800 3233 18813 3279
rect 18741 3220 18813 3233
rect 19061 3279 19133 3292
rect 19061 3233 19074 3279
rect 19120 3233 19133 3279
rect 19061 3220 19133 3233
rect 19381 3279 19453 3292
rect 19381 3233 19394 3279
rect 19440 3233 19453 3279
rect 19381 3220 19453 3233
rect 19701 3279 19773 3292
rect 19701 3233 19714 3279
rect 19760 3233 19773 3279
rect 19701 3220 19773 3233
rect 19989 3287 20061 3300
rect 19989 3241 20002 3287
rect 20048 3241 20061 3287
rect 19989 3228 20061 3241
rect 18589 3096 18645 3220
rect 19069 3172 19125 3220
rect 19069 3116 19285 3172
rect 19069 3096 19125 3116
rect 19709 3096 19765 3220
rect 18749 2476 18805 2496
rect 19389 2476 19445 2496
rect 18749 2420 18965 2476
rect 19389 2420 19605 2476
rect 18749 2356 18805 2420
rect 19389 2356 19445 2420
rect 18581 2343 18653 2356
rect 18581 2297 18594 2343
rect 18640 2297 18653 2343
rect 18581 2284 18653 2297
rect 18741 2343 18813 2356
rect 18741 2297 18754 2343
rect 18800 2297 18813 2343
rect 18741 2284 18813 2297
rect 19061 2343 19133 2356
rect 19061 2297 19074 2343
rect 19120 2297 19133 2343
rect 19061 2284 19133 2297
rect 19381 2343 19453 2356
rect 19381 2297 19394 2343
rect 19440 2297 19453 2343
rect 19381 2284 19453 2297
rect 19701 2343 19773 2356
rect 19701 2297 19714 2343
rect 19760 2297 19773 2343
rect 19701 2284 19773 2297
rect 18589 2160 18645 2284
rect 19069 2236 19125 2284
rect 19069 2180 19285 2236
rect 19069 2160 19125 2180
rect 19709 2160 19765 2284
rect 18589 1224 18645 1560
rect 18749 1224 18805 1560
rect 18909 1224 18965 1560
rect 19069 1224 19125 1560
rect 19229 1224 19285 1560
rect 19389 1224 19445 1560
rect 19549 1224 19605 1560
rect 19709 1224 19765 1560
rect 18749 604 18805 624
rect 19389 604 19445 624
rect 18749 548 18965 604
rect 19389 548 19605 604
rect 18749 484 18805 548
rect 19389 484 19445 548
rect 18581 471 18653 484
rect 18581 425 18594 471
rect 18640 425 18653 471
rect 18581 412 18653 425
rect 18741 471 18813 484
rect 18741 425 18754 471
rect 18800 425 18813 471
rect 18741 412 18813 425
rect 19061 471 19133 484
rect 19061 425 19074 471
rect 19120 425 19133 471
rect 19061 412 19133 425
rect 19381 471 19453 484
rect 19381 425 19394 471
rect 19440 425 19453 471
rect 19381 412 19453 425
rect 19701 471 19773 484
rect 19701 425 19714 471
rect 19760 425 19773 471
rect 19701 412 19773 425
rect 18589 288 18645 412
rect 19069 364 19125 412
rect 19069 308 19285 364
rect 19069 288 19125 308
rect 19709 288 19765 412
rect 18749 -332 18805 -312
rect 19389 -332 19445 -312
rect 18749 -388 18965 -332
rect 19389 -388 19605 -332
rect 18293 -457 18365 -444
rect 18749 -452 18805 -388
rect 19389 -452 19445 -388
rect 19997 -444 20053 3228
rect 18293 -503 18306 -457
rect 18352 -503 18365 -457
rect 18293 -516 18365 -503
rect 18581 -465 18653 -452
rect 18581 -511 18594 -465
rect 18640 -511 18653 -465
rect 18301 -648 18357 -516
rect 18581 -524 18653 -511
rect 18741 -465 18813 -452
rect 18741 -511 18754 -465
rect 18800 -511 18813 -465
rect 18741 -524 18813 -511
rect 19061 -465 19133 -452
rect 19061 -511 19074 -465
rect 19120 -511 19133 -465
rect 19061 -524 19133 -511
rect 19381 -465 19453 -452
rect 19381 -511 19394 -465
rect 19440 -511 19453 -465
rect 19381 -524 19453 -511
rect 19701 -465 19773 -452
rect 19701 -511 19714 -465
rect 19760 -511 19773 -465
rect 19701 -524 19773 -511
rect 19989 -457 20061 -444
rect 19989 -503 20002 -457
rect 20048 -503 20061 -457
rect 19989 -516 20061 -503
rect 18589 -648 18645 -524
rect 19069 -572 19125 -524
rect 19069 -628 19285 -572
rect 19069 -648 19125 -628
rect 19709 -648 19765 -524
rect 19997 -648 20053 -516
rect 18749 -1268 18805 -1248
rect 19389 -1268 19445 -1248
rect 18749 -1324 18965 -1268
rect 19389 -1324 19605 -1268
rect 18749 -1388 18805 -1324
rect 19389 -1388 19445 -1324
rect 18741 -1401 18813 -1388
rect 18741 -1447 18754 -1401
rect 18800 -1447 18813 -1401
rect 18741 -1460 18813 -1447
rect 19381 -1401 19453 -1388
rect 19381 -1447 19394 -1401
rect 19440 -1447 19453 -1401
rect 19381 -1460 19453 -1447
rect 23733 4245 23805 4258
rect 23733 4199 23746 4245
rect 23792 4199 23805 4245
rect 23733 4186 23805 4199
rect 24373 4245 24445 4258
rect 24373 4199 24386 4245
rect 24432 4199 24445 4245
rect 24373 4186 24445 4199
rect 24853 4245 24925 4258
rect 24853 4199 24866 4245
rect 24912 4199 24925 4245
rect 24853 4186 24925 4199
rect 23741 4032 23797 4186
rect 24381 4108 24437 4186
rect 24221 4052 24437 4108
rect 24381 4032 24437 4052
rect 24861 4032 24917 4186
rect 23453 3300 23509 3432
rect 24061 3412 24117 3432
rect 24701 3412 24757 3432
rect 23901 3356 24117 3412
rect 24541 3356 24757 3412
rect 23445 3287 23517 3300
rect 24061 3292 24117 3356
rect 24701 3292 24757 3356
rect 25149 3300 25205 3432
rect 23445 3241 23458 3287
rect 23504 3241 23517 3287
rect 23445 3228 23517 3241
rect 23733 3279 23805 3292
rect 23733 3233 23746 3279
rect 23792 3233 23805 3279
rect 23453 -444 23509 3228
rect 23733 3220 23805 3233
rect 24053 3279 24125 3292
rect 24053 3233 24066 3279
rect 24112 3233 24125 3279
rect 24053 3220 24125 3233
rect 24373 3279 24445 3292
rect 24373 3233 24386 3279
rect 24432 3233 24445 3279
rect 24373 3220 24445 3233
rect 24693 3279 24765 3292
rect 24693 3233 24706 3279
rect 24752 3233 24765 3279
rect 24693 3220 24765 3233
rect 24853 3279 24925 3292
rect 24853 3233 24866 3279
rect 24912 3233 24925 3279
rect 24853 3220 24925 3233
rect 25141 3287 25213 3300
rect 25141 3241 25154 3287
rect 25200 3241 25213 3287
rect 25141 3228 25213 3241
rect 23741 3096 23797 3220
rect 24381 3172 24437 3220
rect 24221 3116 24437 3172
rect 24381 3096 24437 3116
rect 24861 3096 24917 3220
rect 24061 2476 24117 2496
rect 24701 2476 24757 2496
rect 23901 2420 24117 2476
rect 24541 2420 24757 2476
rect 24061 2356 24117 2420
rect 24701 2356 24757 2420
rect 23733 2343 23805 2356
rect 23733 2297 23746 2343
rect 23792 2297 23805 2343
rect 23733 2284 23805 2297
rect 24053 2343 24125 2356
rect 24053 2297 24066 2343
rect 24112 2297 24125 2343
rect 24053 2284 24125 2297
rect 24373 2343 24445 2356
rect 24373 2297 24386 2343
rect 24432 2297 24445 2343
rect 24373 2284 24445 2297
rect 24693 2343 24765 2356
rect 24693 2297 24706 2343
rect 24752 2297 24765 2343
rect 24693 2284 24765 2297
rect 24853 2343 24925 2356
rect 24853 2297 24866 2343
rect 24912 2297 24925 2343
rect 24853 2284 24925 2297
rect 23741 2160 23797 2284
rect 24381 2236 24437 2284
rect 24221 2180 24437 2236
rect 24381 2160 24437 2180
rect 24861 2160 24917 2284
rect 23741 1224 23797 1560
rect 23901 1224 23957 1560
rect 24061 1224 24117 1560
rect 24221 1224 24277 1560
rect 24381 1224 24437 1560
rect 24541 1224 24597 1560
rect 24701 1224 24757 1560
rect 24861 1224 24917 1560
rect 24061 604 24117 624
rect 24701 604 24757 624
rect 23901 548 24117 604
rect 24541 548 24757 604
rect 24061 484 24117 548
rect 24701 484 24757 548
rect 23733 471 23805 484
rect 23733 425 23746 471
rect 23792 425 23805 471
rect 23733 412 23805 425
rect 24053 471 24125 484
rect 24053 425 24066 471
rect 24112 425 24125 471
rect 24053 412 24125 425
rect 24373 471 24445 484
rect 24373 425 24386 471
rect 24432 425 24445 471
rect 24373 412 24445 425
rect 24693 471 24765 484
rect 24693 425 24706 471
rect 24752 425 24765 471
rect 24693 412 24765 425
rect 24853 471 24925 484
rect 24853 425 24866 471
rect 24912 425 24925 471
rect 24853 412 24925 425
rect 23741 288 23797 412
rect 24381 364 24437 412
rect 24221 308 24437 364
rect 24381 288 24437 308
rect 24861 288 24917 412
rect 24061 -332 24117 -312
rect 24701 -332 24757 -312
rect 23901 -388 24117 -332
rect 24541 -388 24757 -332
rect 23445 -457 23517 -444
rect 24061 -452 24117 -388
rect 24701 -452 24757 -388
rect 25149 -444 25205 3228
rect 23445 -503 23458 -457
rect 23504 -503 23517 -457
rect 23445 -516 23517 -503
rect 23733 -465 23805 -452
rect 23733 -511 23746 -465
rect 23792 -511 23805 -465
rect 23453 -648 23509 -516
rect 23733 -524 23805 -511
rect 24053 -465 24125 -452
rect 24053 -511 24066 -465
rect 24112 -511 24125 -465
rect 24053 -524 24125 -511
rect 24373 -465 24445 -452
rect 24373 -511 24386 -465
rect 24432 -511 24445 -465
rect 24373 -524 24445 -511
rect 24693 -465 24765 -452
rect 24693 -511 24706 -465
rect 24752 -511 24765 -465
rect 24693 -524 24765 -511
rect 24853 -465 24925 -452
rect 24853 -511 24866 -465
rect 24912 -511 24925 -465
rect 24853 -524 24925 -511
rect 25141 -457 25213 -444
rect 25141 -503 25154 -457
rect 25200 -503 25213 -457
rect 25141 -516 25213 -503
rect 23741 -648 23797 -524
rect 24381 -572 24437 -524
rect 24221 -628 24437 -572
rect 24381 -648 24437 -628
rect 24861 -648 24917 -524
rect 25149 -648 25205 -516
rect 24061 -1268 24117 -1248
rect 24701 -1268 24757 -1248
rect 23901 -1324 24117 -1268
rect 24541 -1324 24757 -1268
rect 24061 -1388 24117 -1324
rect 24701 -1388 24757 -1324
rect 24053 -1401 24125 -1388
rect 24053 -1447 24066 -1401
rect 24112 -1447 24125 -1401
rect 24053 -1460 24125 -1447
rect 24693 -1401 24765 -1388
rect 24693 -1447 24706 -1401
rect 24752 -1447 24765 -1401
rect 24693 -1460 24765 -1447
rect 27702 4245 27774 4258
rect 27702 4199 27715 4245
rect 27761 4199 27774 4245
rect 27702 4186 27774 4199
rect 28182 4245 28254 4258
rect 28182 4199 28195 4245
rect 28241 4199 28254 4245
rect 28182 4186 28254 4199
rect 28822 4245 28894 4258
rect 28822 4199 28835 4245
rect 28881 4199 28894 4245
rect 28822 4186 28894 4199
rect 27710 4032 27766 4186
rect 28190 4108 28246 4186
rect 28190 4052 28406 4108
rect 28190 4032 28246 4052
rect 28830 4032 28886 4186
rect 27422 3300 27478 3432
rect 27870 3412 27926 3432
rect 28510 3412 28566 3432
rect 27870 3356 28086 3412
rect 28510 3356 28726 3412
rect 27414 3287 27486 3300
rect 27870 3292 27926 3356
rect 28510 3292 28566 3356
rect 29118 3300 29174 3432
rect 27414 3241 27427 3287
rect 27473 3241 27486 3287
rect 27414 3228 27486 3241
rect 27702 3279 27774 3292
rect 27702 3233 27715 3279
rect 27761 3233 27774 3279
rect 27422 -444 27478 3228
rect 27702 3220 27774 3233
rect 27862 3279 27934 3292
rect 27862 3233 27875 3279
rect 27921 3233 27934 3279
rect 27862 3220 27934 3233
rect 28182 3279 28254 3292
rect 28182 3233 28195 3279
rect 28241 3233 28254 3279
rect 28182 3220 28254 3233
rect 28502 3279 28574 3292
rect 28502 3233 28515 3279
rect 28561 3233 28574 3279
rect 28502 3220 28574 3233
rect 28822 3279 28894 3292
rect 28822 3233 28835 3279
rect 28881 3233 28894 3279
rect 28822 3220 28894 3233
rect 29110 3287 29182 3300
rect 29110 3241 29123 3287
rect 29169 3241 29182 3287
rect 29110 3228 29182 3241
rect 27710 3096 27766 3220
rect 28190 3172 28246 3220
rect 28190 3116 28406 3172
rect 28190 3096 28246 3116
rect 28830 3096 28886 3220
rect 27870 2476 27926 2496
rect 28510 2476 28566 2496
rect 27870 2420 28086 2476
rect 28510 2420 28726 2476
rect 27870 2356 27926 2420
rect 28510 2356 28566 2420
rect 27702 2343 27774 2356
rect 27702 2297 27715 2343
rect 27761 2297 27774 2343
rect 27702 2284 27774 2297
rect 27862 2343 27934 2356
rect 27862 2297 27875 2343
rect 27921 2297 27934 2343
rect 27862 2284 27934 2297
rect 28182 2343 28254 2356
rect 28182 2297 28195 2343
rect 28241 2297 28254 2343
rect 28182 2284 28254 2297
rect 28502 2343 28574 2356
rect 28502 2297 28515 2343
rect 28561 2297 28574 2343
rect 28502 2284 28574 2297
rect 28822 2343 28894 2356
rect 28822 2297 28835 2343
rect 28881 2297 28894 2343
rect 28822 2284 28894 2297
rect 27710 2160 27766 2284
rect 28190 2236 28246 2284
rect 28190 2180 28406 2236
rect 28190 2160 28246 2180
rect 28830 2160 28886 2284
rect 27710 1224 27766 1560
rect 27870 1224 27926 1560
rect 28030 1224 28086 1560
rect 28190 1224 28246 1560
rect 28350 1224 28406 1560
rect 28510 1224 28566 1560
rect 28670 1224 28726 1560
rect 28830 1224 28886 1560
rect 27870 604 27926 624
rect 28510 604 28566 624
rect 27870 548 28086 604
rect 28510 548 28726 604
rect 27870 484 27926 548
rect 28510 484 28566 548
rect 27702 471 27774 484
rect 27702 425 27715 471
rect 27761 425 27774 471
rect 27702 412 27774 425
rect 27862 471 27934 484
rect 27862 425 27875 471
rect 27921 425 27934 471
rect 27862 412 27934 425
rect 28182 471 28254 484
rect 28182 425 28195 471
rect 28241 425 28254 471
rect 28182 412 28254 425
rect 28502 471 28574 484
rect 28502 425 28515 471
rect 28561 425 28574 471
rect 28502 412 28574 425
rect 28822 471 28894 484
rect 28822 425 28835 471
rect 28881 425 28894 471
rect 28822 412 28894 425
rect 27710 288 27766 412
rect 28190 364 28246 412
rect 28190 308 28406 364
rect 28190 288 28246 308
rect 28830 288 28886 412
rect 27870 -332 27926 -312
rect 28510 -332 28566 -312
rect 27870 -388 28086 -332
rect 28510 -388 28726 -332
rect 27414 -457 27486 -444
rect 27870 -452 27926 -388
rect 28510 -452 28566 -388
rect 29118 -444 29174 3228
rect 27414 -503 27427 -457
rect 27473 -503 27486 -457
rect 27414 -516 27486 -503
rect 27702 -465 27774 -452
rect 27702 -511 27715 -465
rect 27761 -511 27774 -465
rect 27422 -648 27478 -516
rect 27702 -524 27774 -511
rect 27862 -465 27934 -452
rect 27862 -511 27875 -465
rect 27921 -511 27934 -465
rect 27862 -524 27934 -511
rect 28182 -465 28254 -452
rect 28182 -511 28195 -465
rect 28241 -511 28254 -465
rect 28182 -524 28254 -511
rect 28502 -465 28574 -452
rect 28502 -511 28515 -465
rect 28561 -511 28574 -465
rect 28502 -524 28574 -511
rect 28822 -465 28894 -452
rect 28822 -511 28835 -465
rect 28881 -511 28894 -465
rect 28822 -524 28894 -511
rect 29110 -457 29182 -444
rect 29110 -503 29123 -457
rect 29169 -503 29182 -457
rect 29110 -516 29182 -503
rect 27710 -648 27766 -524
rect 28190 -572 28246 -524
rect 28190 -628 28406 -572
rect 28190 -648 28246 -628
rect 28830 -648 28886 -524
rect 29118 -648 29174 -516
rect 27870 -1268 27926 -1248
rect 28510 -1268 28566 -1248
rect 27870 -1324 28086 -1268
rect 28510 -1324 28726 -1268
rect 27870 -1388 27926 -1324
rect 28510 -1388 28566 -1324
rect 27862 -1401 27934 -1388
rect 27862 -1447 27875 -1401
rect 27921 -1447 27934 -1401
rect 27862 -1460 27934 -1447
rect 28502 -1401 28574 -1388
rect 28502 -1447 28515 -1401
rect 28561 -1447 28574 -1401
rect 28502 -1460 28574 -1447
rect 34118 2652 34190 2665
rect 34118 2606 34131 2652
rect 34177 2606 34190 2652
rect 34118 2593 34190 2606
rect 34278 2652 34350 2665
rect 34278 2606 34291 2652
rect 34337 2606 34350 2652
rect 34278 2593 34350 2606
rect 34126 2532 34182 2593
rect 34286 2532 34342 2593
rect 38254 2652 38326 2665
rect 38254 2606 38267 2652
rect 38313 2606 38326 2652
rect 38254 2593 38326 2606
rect 38414 2652 38486 2665
rect 38414 2606 38427 2652
rect 38473 2606 38486 2652
rect 38414 2593 38486 2606
rect 38262 2532 38318 2593
rect 38422 2532 38478 2593
rect 32718 1738 32774 1932
rect 32710 1725 32782 1738
rect 32710 1679 32723 1725
rect 32769 1679 32782 1725
rect 32710 1666 32782 1679
rect 32718 -382 32774 1666
rect 33006 1605 33062 1932
rect 33166 1605 33222 1932
rect 33326 1605 33382 1932
rect 33486 1605 33542 1932
rect 33646 1605 33702 1932
rect 33806 1605 33862 1932
rect 33966 1605 34022 1932
rect 34126 1605 34182 1932
rect 34286 1605 34342 1932
rect 34446 1605 34502 1932
rect 34606 1605 34662 1932
rect 34766 1605 34822 1932
rect 34926 1605 34982 1932
rect 35086 1605 35142 1932
rect 35246 1605 35302 1932
rect 35406 1605 35462 1932
rect 35694 1738 35750 1932
rect 35686 1725 35758 1738
rect 35686 1679 35699 1725
rect 35745 1679 35758 1725
rect 35686 1666 35758 1679
rect 36854 1738 36910 1932
rect 33006 1592 35462 1605
rect 33006 1546 34131 1592
rect 34177 1546 34291 1592
rect 34337 1546 35462 1592
rect 33006 1533 35462 1546
rect 33006 545 33062 1533
rect 33166 545 33222 1533
rect 33326 545 33382 1533
rect 33486 545 33542 1533
rect 33646 545 33702 1533
rect 33806 545 33862 1533
rect 33966 545 34022 1533
rect 34126 545 34182 1533
rect 34286 545 34342 1533
rect 34446 545 34502 1533
rect 34606 545 34662 1533
rect 34766 545 34822 1533
rect 34926 545 34982 1533
rect 35086 545 35142 1533
rect 35246 545 35302 1533
rect 35406 545 35462 1533
rect 33006 532 35462 545
rect 33006 486 34131 532
rect 34177 486 34291 532
rect 34337 486 35462 532
rect 33006 473 35462 486
rect 32710 -395 32782 -382
rect 32710 -441 32723 -395
rect 32769 -441 32782 -395
rect 32710 -454 32782 -441
rect 32718 -648 32774 -454
rect 33006 -515 33062 473
rect 33166 -515 33222 473
rect 33326 -515 33382 473
rect 33486 -515 33542 473
rect 33646 -515 33702 473
rect 33806 -515 33862 473
rect 33966 -515 34022 473
rect 34126 -515 34182 473
rect 34286 -515 34342 473
rect 34446 -515 34502 473
rect 34606 -515 34662 473
rect 34766 -515 34822 473
rect 34926 -515 34982 473
rect 35086 -515 35142 473
rect 35246 -515 35302 473
rect 35406 -515 35462 473
rect 35694 -382 35750 1666
rect 36846 1725 36918 1738
rect 36846 1679 36859 1725
rect 36905 1679 36918 1725
rect 36846 1666 36918 1679
rect 35686 -395 35758 -382
rect 35686 -441 35699 -395
rect 35745 -441 35758 -395
rect 35686 -454 35758 -441
rect 36854 -382 36910 1666
rect 37142 1605 37198 1932
rect 37302 1605 37358 1932
rect 37462 1605 37518 1932
rect 37622 1605 37678 1932
rect 37782 1605 37838 1932
rect 37942 1605 37998 1932
rect 38102 1605 38158 1932
rect 38262 1605 38318 1932
rect 38422 1605 38478 1932
rect 38582 1605 38638 1932
rect 38742 1605 38798 1932
rect 38902 1605 38958 1932
rect 39062 1605 39118 1932
rect 39222 1605 39278 1932
rect 39382 1605 39438 1932
rect 39542 1605 39598 1932
rect 39830 1738 39886 1932
rect 39822 1725 39894 1738
rect 39822 1679 39835 1725
rect 39881 1679 39894 1725
rect 39822 1666 39894 1679
rect 37142 1592 39598 1605
rect 37142 1546 38267 1592
rect 38313 1546 38427 1592
rect 38473 1546 39598 1592
rect 37142 1533 39598 1546
rect 37142 545 37198 1533
rect 37302 545 37358 1533
rect 37462 545 37518 1533
rect 37622 545 37678 1533
rect 37782 545 37838 1533
rect 37942 545 37998 1533
rect 38102 545 38158 1533
rect 38262 545 38318 1533
rect 38422 545 38478 1533
rect 38582 545 38638 1533
rect 38742 545 38798 1533
rect 38902 545 38958 1533
rect 39062 545 39118 1533
rect 39222 545 39278 1533
rect 39382 545 39438 1533
rect 39542 545 39598 1533
rect 37142 532 39598 545
rect 37142 486 38267 532
rect 38313 486 38427 532
rect 38473 486 39598 532
rect 37142 473 39598 486
rect 33006 -528 35462 -515
rect 33006 -574 34131 -528
rect 34177 -574 34291 -528
rect 34337 -574 35462 -528
rect 33006 -587 35462 -574
rect 33006 -648 33062 -587
rect 33166 -648 33222 -587
rect 33326 -648 33382 -587
rect 33486 -648 33542 -587
rect 33646 -648 33702 -587
rect 33806 -648 33862 -587
rect 33966 -648 34022 -587
rect 34126 -648 34182 -587
rect 34286 -648 34342 -587
rect 34446 -648 34502 -587
rect 34606 -648 34662 -587
rect 34766 -648 34822 -587
rect 34926 -648 34982 -587
rect 35086 -648 35142 -587
rect 35246 -648 35302 -587
rect 35406 -648 35462 -587
rect 35694 -648 35750 -454
rect 36846 -395 36918 -382
rect 36846 -441 36859 -395
rect 36905 -441 36918 -395
rect 36846 -454 36918 -441
rect 36854 -648 36910 -454
rect 37142 -515 37198 473
rect 37302 -515 37358 473
rect 37462 -515 37518 473
rect 37622 -515 37678 473
rect 37782 -515 37838 473
rect 37942 -515 37998 473
rect 38102 -515 38158 473
rect 38262 -515 38318 473
rect 38422 -515 38478 473
rect 38582 -515 38638 473
rect 38742 -515 38798 473
rect 38902 -515 38958 473
rect 39062 -515 39118 473
rect 39222 -515 39278 473
rect 39382 -515 39438 473
rect 39542 -515 39598 473
rect 39830 -382 39886 1666
rect 39822 -395 39894 -382
rect 39822 -441 39835 -395
rect 39881 -441 39894 -395
rect 39822 -454 39894 -441
rect 37142 -528 39598 -515
rect 37142 -574 38267 -528
rect 38313 -574 38427 -528
rect 38473 -574 39598 -528
rect 37142 -587 39598 -574
rect 37142 -648 37198 -587
rect 37302 -648 37358 -587
rect 37462 -648 37518 -587
rect 37622 -648 37678 -587
rect 37782 -648 37838 -587
rect 37942 -648 37998 -587
rect 38102 -648 38158 -587
rect 38262 -648 38318 -587
rect 38422 -648 38478 -587
rect 38582 -648 38638 -587
rect 38742 -648 38798 -587
rect 38902 -648 38958 -587
rect 39062 -648 39118 -587
rect 39222 -648 39278 -587
rect 39382 -648 39438 -587
rect 39542 -648 39598 -587
rect 39830 -648 39886 -454
rect 43814 2652 43886 2665
rect 43814 2606 43827 2652
rect 43873 2606 43886 2652
rect 43814 2593 43886 2606
rect 43974 2652 44046 2665
rect 43974 2606 43987 2652
rect 44033 2606 44046 2652
rect 43974 2593 44046 2606
rect 43822 2532 43878 2593
rect 43982 2532 44038 2593
rect 47950 2652 48022 2665
rect 47950 2606 47963 2652
rect 48009 2606 48022 2652
rect 47950 2593 48022 2606
rect 48110 2652 48182 2665
rect 48110 2606 48123 2652
rect 48169 2606 48182 2652
rect 48110 2593 48182 2606
rect 47958 2532 48014 2593
rect 48118 2532 48174 2593
rect 42414 1738 42470 1932
rect 42406 1725 42478 1738
rect 42406 1679 42419 1725
rect 42465 1679 42478 1725
rect 42406 1666 42478 1679
rect 42414 -382 42470 1666
rect 42702 1605 42758 1932
rect 42862 1605 42918 1932
rect 43022 1605 43078 1932
rect 43182 1605 43238 1932
rect 43342 1605 43398 1932
rect 43502 1605 43558 1932
rect 43662 1605 43718 1932
rect 43822 1605 43878 1932
rect 43982 1605 44038 1932
rect 44142 1605 44198 1932
rect 44302 1605 44358 1932
rect 44462 1605 44518 1932
rect 44622 1605 44678 1932
rect 44782 1605 44838 1932
rect 44942 1605 44998 1932
rect 45102 1605 45158 1932
rect 45390 1738 45446 1932
rect 45382 1725 45454 1738
rect 45382 1679 45395 1725
rect 45441 1679 45454 1725
rect 45382 1666 45454 1679
rect 46550 1738 46606 1932
rect 42702 1592 45158 1605
rect 42702 1546 43827 1592
rect 43873 1546 43987 1592
rect 44033 1546 45158 1592
rect 42702 1533 45158 1546
rect 42702 545 42758 1533
rect 42862 545 42918 1533
rect 43022 545 43078 1533
rect 43182 545 43238 1533
rect 43342 545 43398 1533
rect 43502 545 43558 1533
rect 43662 545 43718 1533
rect 43822 545 43878 1533
rect 43982 545 44038 1533
rect 44142 545 44198 1533
rect 44302 545 44358 1533
rect 44462 545 44518 1533
rect 44622 545 44678 1533
rect 44782 545 44838 1533
rect 44942 545 44998 1533
rect 45102 545 45158 1533
rect 42702 532 45158 545
rect 42702 486 43827 532
rect 43873 486 43987 532
rect 44033 486 45158 532
rect 42702 473 45158 486
rect 42406 -395 42478 -382
rect 42406 -441 42419 -395
rect 42465 -441 42478 -395
rect 42406 -454 42478 -441
rect 42414 -648 42470 -454
rect 42702 -515 42758 473
rect 42862 -515 42918 473
rect 43022 -515 43078 473
rect 43182 -515 43238 473
rect 43342 -515 43398 473
rect 43502 -515 43558 473
rect 43662 -515 43718 473
rect 43822 -515 43878 473
rect 43982 -515 44038 473
rect 44142 -515 44198 473
rect 44302 -515 44358 473
rect 44462 -515 44518 473
rect 44622 -515 44678 473
rect 44782 -515 44838 473
rect 44942 -515 44998 473
rect 45102 -515 45158 473
rect 45390 -382 45446 1666
rect 46542 1725 46614 1738
rect 46542 1679 46555 1725
rect 46601 1679 46614 1725
rect 46542 1666 46614 1679
rect 45382 -395 45454 -382
rect 45382 -441 45395 -395
rect 45441 -441 45454 -395
rect 45382 -454 45454 -441
rect 46550 -382 46606 1666
rect 46838 1605 46894 1932
rect 46998 1605 47054 1932
rect 47158 1605 47214 1932
rect 47318 1605 47374 1932
rect 47478 1605 47534 1932
rect 47638 1605 47694 1932
rect 47798 1605 47854 1932
rect 47958 1605 48014 1932
rect 48118 1605 48174 1932
rect 48278 1605 48334 1932
rect 48438 1605 48494 1932
rect 48598 1605 48654 1932
rect 48758 1605 48814 1932
rect 48918 1605 48974 1932
rect 49078 1605 49134 1932
rect 49238 1605 49294 1932
rect 49526 1738 49582 1932
rect 49518 1725 49590 1738
rect 49518 1679 49531 1725
rect 49577 1679 49590 1725
rect 49518 1666 49590 1679
rect 46838 1592 49294 1605
rect 46838 1546 47963 1592
rect 48009 1546 48123 1592
rect 48169 1546 49294 1592
rect 46838 1533 49294 1546
rect 46838 545 46894 1533
rect 46998 545 47054 1533
rect 47158 545 47214 1533
rect 47318 545 47374 1533
rect 47478 545 47534 1533
rect 47638 545 47694 1533
rect 47798 545 47854 1533
rect 47958 545 48014 1533
rect 48118 545 48174 1533
rect 48278 545 48334 1533
rect 48438 545 48494 1533
rect 48598 545 48654 1533
rect 48758 545 48814 1533
rect 48918 545 48974 1533
rect 49078 545 49134 1533
rect 49238 545 49294 1533
rect 46838 532 49294 545
rect 46838 486 47963 532
rect 48009 486 48123 532
rect 48169 486 49294 532
rect 46838 473 49294 486
rect 42702 -528 45158 -515
rect 42702 -574 43827 -528
rect 43873 -574 43987 -528
rect 44033 -574 45158 -528
rect 42702 -587 45158 -574
rect 42702 -648 42758 -587
rect 42862 -648 42918 -587
rect 43022 -648 43078 -587
rect 43182 -648 43238 -587
rect 43342 -648 43398 -587
rect 43502 -648 43558 -587
rect 43662 -648 43718 -587
rect 43822 -648 43878 -587
rect 43982 -648 44038 -587
rect 44142 -648 44198 -587
rect 44302 -648 44358 -587
rect 44462 -648 44518 -587
rect 44622 -648 44678 -587
rect 44782 -648 44838 -587
rect 44942 -648 44998 -587
rect 45102 -648 45158 -587
rect 45390 -648 45446 -454
rect 46542 -395 46614 -382
rect 46542 -441 46555 -395
rect 46601 -441 46614 -395
rect 46542 -454 46614 -441
rect 46550 -648 46606 -454
rect 46838 -515 46894 473
rect 46998 -515 47054 473
rect 47158 -515 47214 473
rect 47318 -515 47374 473
rect 47478 -515 47534 473
rect 47638 -515 47694 473
rect 47798 -515 47854 473
rect 47958 -515 48014 473
rect 48118 -515 48174 473
rect 48278 -515 48334 473
rect 48438 -515 48494 473
rect 48598 -515 48654 473
rect 48758 -515 48814 473
rect 48918 -515 48974 473
rect 49078 -515 49134 473
rect 49238 -515 49294 473
rect 49526 -382 49582 1666
rect 49518 -395 49590 -382
rect 49518 -441 49531 -395
rect 49577 -441 49590 -395
rect 49518 -454 49590 -441
rect 46838 -528 49294 -515
rect 46838 -574 47963 -528
rect 48009 -574 48123 -528
rect 48169 -574 49294 -528
rect 46838 -587 49294 -574
rect 46838 -648 46894 -587
rect 46998 -648 47054 -587
rect 47158 -648 47214 -587
rect 47318 -648 47374 -587
rect 47478 -648 47534 -587
rect 47638 -648 47694 -587
rect 47798 -648 47854 -587
rect 47958 -648 48014 -587
rect 48118 -648 48174 -587
rect 48278 -648 48334 -587
rect 48438 -648 48494 -587
rect 48598 -648 48654 -587
rect 48758 -648 48814 -587
rect 48918 -648 48974 -587
rect 49078 -648 49134 -587
rect 49238 -648 49294 -587
rect 49526 -648 49582 -454
rect 53510 2652 53582 2665
rect 53510 2606 53523 2652
rect 53569 2606 53582 2652
rect 53510 2593 53582 2606
rect 53670 2652 53742 2665
rect 53670 2606 53683 2652
rect 53729 2606 53742 2652
rect 53670 2593 53742 2606
rect 53518 2532 53574 2593
rect 53678 2532 53734 2593
rect 57646 2652 57718 2665
rect 57646 2606 57659 2652
rect 57705 2606 57718 2652
rect 57646 2593 57718 2606
rect 57806 2652 57878 2665
rect 57806 2606 57819 2652
rect 57865 2606 57878 2652
rect 57806 2593 57878 2606
rect 57654 2532 57710 2593
rect 57814 2532 57870 2593
rect 52110 1738 52166 1932
rect 52102 1725 52174 1738
rect 52102 1679 52115 1725
rect 52161 1679 52174 1725
rect 52102 1666 52174 1679
rect 52110 -382 52166 1666
rect 52398 1605 52454 1932
rect 52558 1605 52614 1932
rect 52718 1605 52774 1932
rect 52878 1605 52934 1932
rect 53038 1605 53094 1932
rect 53198 1605 53254 1932
rect 53358 1605 53414 1932
rect 53518 1605 53574 1932
rect 53678 1605 53734 1932
rect 53838 1605 53894 1932
rect 53998 1605 54054 1932
rect 54158 1605 54214 1932
rect 54318 1605 54374 1932
rect 54478 1605 54534 1932
rect 54638 1605 54694 1932
rect 54798 1605 54854 1932
rect 55086 1738 55142 1932
rect 55078 1725 55150 1738
rect 55078 1679 55091 1725
rect 55137 1679 55150 1725
rect 55078 1666 55150 1679
rect 56246 1738 56302 1932
rect 52398 1592 54854 1605
rect 52398 1546 53523 1592
rect 53569 1546 53683 1592
rect 53729 1546 54854 1592
rect 52398 1533 54854 1546
rect 52398 545 52454 1533
rect 52558 545 52614 1533
rect 52718 545 52774 1533
rect 52878 545 52934 1533
rect 53038 545 53094 1533
rect 53198 545 53254 1533
rect 53358 545 53414 1533
rect 53518 545 53574 1533
rect 53678 545 53734 1533
rect 53838 545 53894 1533
rect 53998 545 54054 1533
rect 54158 545 54214 1533
rect 54318 545 54374 1533
rect 54478 545 54534 1533
rect 54638 545 54694 1533
rect 54798 545 54854 1533
rect 52398 532 54854 545
rect 52398 486 53523 532
rect 53569 486 53683 532
rect 53729 486 54854 532
rect 52398 473 54854 486
rect 52102 -395 52174 -382
rect 52102 -441 52115 -395
rect 52161 -441 52174 -395
rect 52102 -454 52174 -441
rect 52110 -648 52166 -454
rect 52398 -515 52454 473
rect 52558 -515 52614 473
rect 52718 -515 52774 473
rect 52878 -515 52934 473
rect 53038 -515 53094 473
rect 53198 -515 53254 473
rect 53358 -515 53414 473
rect 53518 -515 53574 473
rect 53678 -515 53734 473
rect 53838 -515 53894 473
rect 53998 -515 54054 473
rect 54158 -515 54214 473
rect 54318 -515 54374 473
rect 54478 -515 54534 473
rect 54638 -515 54694 473
rect 54798 -515 54854 473
rect 55086 -382 55142 1666
rect 56238 1725 56310 1738
rect 56238 1679 56251 1725
rect 56297 1679 56310 1725
rect 56238 1666 56310 1679
rect 55078 -395 55150 -382
rect 55078 -441 55091 -395
rect 55137 -441 55150 -395
rect 55078 -454 55150 -441
rect 56246 -382 56302 1666
rect 56534 1605 56590 1932
rect 56694 1605 56750 1932
rect 56854 1605 56910 1932
rect 57014 1605 57070 1932
rect 57174 1605 57230 1932
rect 57334 1605 57390 1932
rect 57494 1605 57550 1932
rect 57654 1605 57710 1932
rect 57814 1605 57870 1932
rect 57974 1605 58030 1932
rect 58134 1605 58190 1932
rect 58294 1605 58350 1932
rect 58454 1605 58510 1932
rect 58614 1605 58670 1932
rect 58774 1605 58830 1932
rect 58934 1605 58990 1932
rect 59222 1738 59278 1932
rect 59214 1725 59286 1738
rect 59214 1679 59227 1725
rect 59273 1679 59286 1725
rect 59214 1666 59286 1679
rect 56534 1592 58990 1605
rect 56534 1546 57659 1592
rect 57705 1546 57819 1592
rect 57865 1546 58990 1592
rect 56534 1533 58990 1546
rect 56534 545 56590 1533
rect 56694 545 56750 1533
rect 56854 545 56910 1533
rect 57014 545 57070 1533
rect 57174 545 57230 1533
rect 57334 545 57390 1533
rect 57494 545 57550 1533
rect 57654 545 57710 1533
rect 57814 545 57870 1533
rect 57974 545 58030 1533
rect 58134 545 58190 1533
rect 58294 545 58350 1533
rect 58454 545 58510 1533
rect 58614 545 58670 1533
rect 58774 545 58830 1533
rect 58934 545 58990 1533
rect 56534 532 58990 545
rect 56534 486 57659 532
rect 57705 486 57819 532
rect 57865 486 58990 532
rect 56534 473 58990 486
rect 52398 -528 54854 -515
rect 52398 -574 53523 -528
rect 53569 -574 53683 -528
rect 53729 -574 54854 -528
rect 52398 -587 54854 -574
rect 52398 -648 52454 -587
rect 52558 -648 52614 -587
rect 52718 -648 52774 -587
rect 52878 -648 52934 -587
rect 53038 -648 53094 -587
rect 53198 -648 53254 -587
rect 53358 -648 53414 -587
rect 53518 -648 53574 -587
rect 53678 -648 53734 -587
rect 53838 -648 53894 -587
rect 53998 -648 54054 -587
rect 54158 -648 54214 -587
rect 54318 -648 54374 -587
rect 54478 -648 54534 -587
rect 54638 -648 54694 -587
rect 54798 -648 54854 -587
rect 55086 -648 55142 -454
rect 56238 -395 56310 -382
rect 56238 -441 56251 -395
rect 56297 -441 56310 -395
rect 56238 -454 56310 -441
rect 56246 -648 56302 -454
rect 56534 -515 56590 473
rect 56694 -515 56750 473
rect 56854 -515 56910 473
rect 57014 -515 57070 473
rect 57174 -515 57230 473
rect 57334 -515 57390 473
rect 57494 -515 57550 473
rect 57654 -515 57710 473
rect 57814 -515 57870 473
rect 57974 -515 58030 473
rect 58134 -515 58190 473
rect 58294 -515 58350 473
rect 58454 -515 58510 473
rect 58614 -515 58670 473
rect 58774 -515 58830 473
rect 58934 -515 58990 473
rect 59222 -382 59278 1666
rect 59214 -395 59286 -382
rect 59214 -441 59227 -395
rect 59273 -441 59286 -395
rect 59214 -454 59286 -441
rect 56534 -528 58990 -515
rect 56534 -574 57659 -528
rect 57705 -574 57819 -528
rect 57865 -574 58990 -528
rect 56534 -587 58990 -574
rect 56534 -648 56590 -587
rect 56694 -648 56750 -587
rect 56854 -648 56910 -587
rect 57014 -648 57070 -587
rect 57174 -648 57230 -587
rect 57334 -648 57390 -587
rect 57494 -648 57550 -587
rect 57654 -648 57710 -587
rect 57814 -648 57870 -587
rect 57974 -648 58030 -587
rect 58134 -648 58190 -587
rect 58294 -648 58350 -587
rect 58454 -648 58510 -587
rect 58614 -648 58670 -587
rect 58774 -648 58830 -587
rect 58934 -648 58990 -587
rect 59222 -648 59278 -454
rect 63206 2652 63278 2665
rect 63206 2606 63219 2652
rect 63265 2606 63278 2652
rect 63206 2593 63278 2606
rect 63366 2652 63438 2665
rect 63366 2606 63379 2652
rect 63425 2606 63438 2652
rect 63366 2593 63438 2606
rect 63214 2532 63270 2593
rect 63374 2532 63430 2593
rect 61806 1738 61862 1932
rect 61798 1725 61870 1738
rect 61798 1679 61811 1725
rect 61857 1679 61870 1725
rect 61798 1666 61870 1679
rect 61806 -382 61862 1666
rect 62094 1605 62150 1932
rect 62254 1605 62310 1932
rect 62414 1605 62470 1932
rect 62574 1605 62630 1932
rect 62734 1605 62790 1932
rect 62894 1605 62950 1932
rect 63054 1605 63110 1932
rect 63214 1605 63270 1932
rect 63374 1605 63430 1932
rect 63534 1605 63590 1932
rect 63694 1605 63750 1932
rect 63854 1605 63910 1932
rect 64014 1605 64070 1932
rect 64174 1605 64230 1932
rect 64334 1605 64390 1932
rect 64494 1605 64550 1932
rect 64782 1738 64838 1932
rect 64774 1725 64846 1738
rect 64774 1679 64787 1725
rect 64833 1679 64846 1725
rect 64774 1666 64846 1679
rect 62094 1592 64550 1605
rect 62094 1546 63219 1592
rect 63265 1546 63379 1592
rect 63425 1546 64550 1592
rect 62094 1533 64550 1546
rect 62094 545 62150 1533
rect 62254 545 62310 1533
rect 62414 545 62470 1533
rect 62574 545 62630 1533
rect 62734 545 62790 1533
rect 62894 545 62950 1533
rect 63054 545 63110 1533
rect 63214 545 63270 1533
rect 63374 545 63430 1533
rect 63534 545 63590 1533
rect 63694 545 63750 1533
rect 63854 545 63910 1533
rect 64014 545 64070 1533
rect 64174 545 64230 1533
rect 64334 545 64390 1533
rect 64494 545 64550 1533
rect 62094 532 64550 545
rect 62094 486 63219 532
rect 63265 486 63379 532
rect 63425 486 64550 532
rect 62094 473 64550 486
rect 61798 -395 61870 -382
rect 61798 -441 61811 -395
rect 61857 -441 61870 -395
rect 61798 -454 61870 -441
rect 61806 -648 61862 -454
rect 62094 -515 62150 473
rect 62254 -515 62310 473
rect 62414 -515 62470 473
rect 62574 -515 62630 473
rect 62734 -515 62790 473
rect 62894 -515 62950 473
rect 63054 -515 63110 473
rect 63214 -515 63270 473
rect 63374 -515 63430 473
rect 63534 -515 63590 473
rect 63694 -515 63750 473
rect 63854 -515 63910 473
rect 64014 -515 64070 473
rect 64174 -515 64230 473
rect 64334 -515 64390 473
rect 64494 -515 64550 473
rect 64782 -382 64838 1666
rect 64774 -395 64846 -382
rect 64774 -441 64787 -395
rect 64833 -441 64846 -395
rect 64774 -454 64846 -441
rect 62094 -528 64550 -515
rect 62094 -574 63219 -528
rect 63265 -574 63379 -528
rect 63425 -574 64550 -528
rect 62094 -587 64550 -574
rect 62094 -648 62150 -587
rect 62254 -648 62310 -587
rect 62414 -648 62470 -587
rect 62574 -648 62630 -587
rect 62734 -648 62790 -587
rect 62894 -648 62950 -587
rect 63054 -648 63110 -587
rect 63214 -648 63270 -587
rect 63374 -648 63430 -587
rect 63534 -648 63590 -587
rect 63694 -648 63750 -587
rect 63854 -648 63910 -587
rect 64014 -648 64070 -587
rect 64174 -648 64230 -587
rect 64334 -648 64390 -587
rect 64494 -648 64550 -587
rect 64782 -648 64838 -454
rect 7265 -3223 7337 -3209
rect 7265 -3269 7278 -3223
rect 7324 -3269 7337 -3223
rect 7265 -3281 7337 -3269
rect 7745 -3218 7817 -3209
rect 8225 -3218 8297 -3209
rect 7745 -3223 8297 -3218
rect 7745 -3269 7758 -3223
rect 7804 -3269 8238 -3223
rect 8284 -3269 8297 -3223
rect 7745 -3274 8297 -3269
rect 7745 -3281 7817 -3274
rect 7273 -3419 7329 -3281
rect 7753 -3419 7809 -3281
rect 7913 -3419 7969 -3274
rect 8073 -3419 8129 -3274
rect 8225 -3281 8297 -3274
rect 8705 -3222 8777 -3209
rect 8705 -3268 8718 -3222
rect 8764 -3268 8777 -3222
rect 8705 -3281 8777 -3268
rect 8233 -3419 8289 -3281
rect 8713 -3419 8769 -3281
rect 1455 -4604 3727 -4571
rect 1159 -4642 1231 -4629
rect 1159 -4688 1172 -4642
rect 1218 -4688 1231 -4642
rect 1455 -4650 1704 -4604
rect 1750 -4650 1808 -4604
rect 1854 -4650 3727 -4604
rect 1455 -4683 3727 -4650
rect 3823 -4644 3895 -4631
rect 1159 -4701 1231 -4688
rect 3823 -4690 3836 -4644
rect 3882 -4690 3895 -4644
rect 3823 -4703 3895 -4690
rect 3983 -4644 4055 -4631
rect 3983 -4690 3996 -4644
rect 4042 -4690 4055 -4644
rect 3983 -4703 4055 -4690
rect 3831 -4723 3887 -4703
rect 879 -5889 935 -5523
rect 1463 -5816 2439 -5783
rect 1463 -5862 1616 -5816
rect 1662 -5862 1720 -5816
rect 1766 -5862 1824 -5816
rect 1870 -5862 1928 -5816
rect 1974 -5862 2032 -5816
rect 2078 -5862 2136 -5816
rect 2182 -5862 2439 -5816
rect 871 -5902 943 -5889
rect 871 -5948 884 -5902
rect 930 -5948 943 -5902
rect 871 -5961 943 -5948
rect 1167 -5902 1239 -5889
rect 1167 -5948 1180 -5902
rect 1226 -5948 1239 -5902
rect 1167 -5961 1239 -5948
rect 1463 -5895 2439 -5862
rect 879 -5983 935 -5961
rect 1175 -5981 1231 -5961
rect 1463 -5983 1575 -5895
rect 1679 -5983 1791 -5895
rect 1895 -5983 2007 -5895
rect 2111 -5983 2223 -5895
rect 2327 -5982 2439 -5895
rect 3183 -5983 3295 -5523
rect 3735 -5893 3807 -5880
rect 3735 -5939 3748 -5893
rect 3794 -5939 3807 -5893
rect 3735 -5952 3807 -5939
rect 4031 -5893 4103 -5880
rect 4031 -5939 4044 -5893
rect 4090 -5939 4103 -5893
rect 4031 -5952 4103 -5939
rect 3743 -5983 3799 -5952
rect 6985 -5359 7041 -3619
rect 7433 -3653 7489 -3619
rect 8393 -3653 8449 -3633
rect 7433 -3709 7649 -3653
rect 8393 -3709 8609 -3653
rect 7433 -3760 7489 -3709
rect 8393 -3760 8449 -3709
rect 7265 -3773 7337 -3760
rect 7265 -3819 7278 -3773
rect 7324 -3819 7337 -3773
rect 7265 -3832 7337 -3819
rect 7425 -3773 7497 -3760
rect 7425 -3819 7438 -3773
rect 7484 -3819 7497 -3773
rect 7425 -3832 7497 -3819
rect 7745 -3768 7817 -3760
rect 8225 -3768 8297 -3760
rect 7745 -3773 8297 -3768
rect 7745 -3819 7758 -3773
rect 7804 -3819 8238 -3773
rect 8284 -3819 8297 -3773
rect 7745 -3824 8297 -3819
rect 7745 -3832 7817 -3824
rect 7273 -3955 7329 -3832
rect 7753 -3955 7809 -3832
rect 7913 -3955 7969 -3824
rect 8073 -3955 8129 -3824
rect 8225 -3832 8297 -3824
rect 8385 -3773 8457 -3760
rect 8385 -3819 8398 -3773
rect 8444 -3819 8457 -3773
rect 8385 -3832 8457 -3819
rect 8705 -3773 8777 -3760
rect 8705 -3819 8718 -3773
rect 8764 -3819 8777 -3773
rect 8705 -3832 8777 -3819
rect 8233 -3955 8289 -3832
rect 8713 -3955 8769 -3832
rect 7433 -4177 7489 -4155
rect 7433 -4233 7649 -4177
rect 8393 -4233 8609 -4177
rect 7433 -4281 7489 -4233
rect 8393 -4281 8449 -4233
rect 7265 -4294 7337 -4281
rect 7265 -4340 7278 -4294
rect 7324 -4340 7337 -4294
rect 7265 -4353 7337 -4340
rect 7425 -4294 7497 -4281
rect 7425 -4340 7438 -4294
rect 7484 -4340 7497 -4294
rect 7425 -4353 7497 -4340
rect 7745 -4289 7817 -4281
rect 8225 -4289 8297 -4281
rect 7745 -4294 8297 -4289
rect 7745 -4340 7758 -4294
rect 7804 -4340 8238 -4294
rect 8284 -4340 8297 -4294
rect 7745 -4345 7969 -4340
rect 7745 -4353 7817 -4345
rect 7273 -4491 7329 -4353
rect 7753 -4491 7809 -4353
rect 7913 -4491 7969 -4345
rect 8073 -4491 8129 -4340
rect 8225 -4353 8297 -4340
rect 8385 -4294 8457 -4281
rect 8385 -4340 8398 -4294
rect 8444 -4340 8457 -4294
rect 8385 -4353 8457 -4340
rect 8705 -4294 8777 -4281
rect 8705 -4340 8718 -4294
rect 8764 -4340 8777 -4294
rect 8705 -4353 8777 -4340
rect 8233 -4491 8289 -4353
rect 8713 -4491 8769 -4353
rect 7433 -4711 7489 -4691
rect 7433 -4767 7649 -4711
rect 8393 -4767 8609 -4711
rect 7433 -4815 7489 -4767
rect 8393 -4815 8449 -4767
rect 7265 -4828 7337 -4815
rect 7265 -4874 7278 -4828
rect 7324 -4874 7337 -4828
rect 7265 -4887 7337 -4874
rect 7425 -4828 7497 -4815
rect 7425 -4874 7438 -4828
rect 7484 -4874 7497 -4828
rect 7425 -4887 7497 -4874
rect 7745 -4823 7817 -4815
rect 8225 -4823 8297 -4815
rect 7745 -4828 8297 -4823
rect 7745 -4874 7758 -4828
rect 7804 -4874 8238 -4828
rect 8284 -4874 8297 -4828
rect 7745 -4887 7817 -4874
rect 7273 -5027 7329 -4887
rect 7753 -5027 7809 -4887
rect 7913 -5027 7969 -4874
rect 8073 -5027 8129 -4874
rect 8225 -4887 8297 -4874
rect 8385 -4828 8457 -4815
rect 8385 -4874 8398 -4828
rect 8444 -4874 8457 -4828
rect 8385 -4887 8457 -4874
rect 8705 -4828 8777 -4815
rect 8705 -4874 8718 -4828
rect 8764 -4874 8777 -4828
rect 8705 -4887 8777 -4874
rect 8233 -5027 8289 -4887
rect 8713 -5027 8769 -4887
rect 7433 -5247 7489 -5227
rect 8393 -5247 8449 -5227
rect 7433 -5303 7649 -5247
rect 8393 -5303 8609 -5247
rect 7433 -5351 7489 -5303
rect 8393 -5351 8449 -5303
rect 6977 -5372 7049 -5359
rect 6977 -5418 6990 -5372
rect 7036 -5418 7049 -5372
rect 6977 -5431 7049 -5418
rect 7265 -5364 7337 -5351
rect 7265 -5410 7278 -5364
rect 7324 -5410 7337 -5364
rect 7265 -5423 7337 -5410
rect 7425 -5364 7497 -5351
rect 7425 -5410 7438 -5364
rect 7484 -5410 7497 -5364
rect 7425 -5423 7497 -5410
rect 7745 -5359 7817 -5351
rect 8225 -5359 8297 -5351
rect 7745 -5364 8297 -5359
rect 7745 -5410 7758 -5364
rect 7804 -5410 8238 -5364
rect 8284 -5410 8297 -5364
rect 7745 -5423 7817 -5410
rect 6985 -6099 7041 -5431
rect 7273 -5563 7329 -5423
rect 7753 -5563 7809 -5423
rect 7913 -5563 7969 -5410
rect 8073 -5563 8129 -5410
rect 8225 -5423 8297 -5410
rect 8385 -5364 8457 -5351
rect 8385 -5410 8398 -5364
rect 8444 -5410 8457 -5364
rect 8385 -5423 8457 -5410
rect 8705 -5366 8777 -5353
rect 9001 -5359 9057 -3619
rect 18544 -4242 21000 -4229
rect 18544 -4288 20176 -4242
rect 20222 -4288 20280 -4242
rect 20326 -4288 20869 -4242
rect 20915 -4288 21000 -4242
rect 18544 -4301 21000 -4288
rect 18544 -4378 18600 -4301
rect 18704 -4378 18760 -4301
rect 18864 -4378 18920 -4301
rect 19024 -4378 19080 -4301
rect 19184 -4378 19240 -4301
rect 19344 -4378 19400 -4301
rect 19504 -4378 19560 -4301
rect 19664 -4378 19720 -4301
rect 19824 -4378 19880 -4301
rect 19984 -4378 20040 -4301
rect 20144 -4378 20200 -4301
rect 20304 -4378 20360 -4301
rect 20464 -4378 20520 -4301
rect 20624 -4378 20680 -4301
rect 20784 -4378 20840 -4301
rect 20944 -4378 21000 -4301
rect 8705 -5412 8718 -5366
rect 8764 -5412 8777 -5366
rect 8233 -5563 8289 -5423
rect 8705 -5425 8777 -5412
rect 8992 -5372 9065 -5359
rect 8992 -5418 9006 -5372
rect 9052 -5418 9065 -5372
rect 8713 -5563 8769 -5425
rect 8992 -5431 9065 -5418
rect 7433 -5783 7489 -5763
rect 8393 -5783 8449 -5763
rect 7433 -5839 7649 -5783
rect 8393 -5839 8609 -5783
rect 7433 -5887 7489 -5839
rect 8393 -5887 8449 -5839
rect 7265 -5900 7337 -5887
rect 7265 -5946 7278 -5900
rect 7324 -5946 7337 -5900
rect 7265 -5959 7337 -5946
rect 7425 -5900 7497 -5887
rect 7425 -5946 7438 -5900
rect 7484 -5946 7497 -5900
rect 7425 -5959 7497 -5946
rect 7745 -5895 7817 -5887
rect 8225 -5895 8297 -5887
rect 7745 -5900 8297 -5895
rect 7745 -5946 7758 -5900
rect 7804 -5946 8238 -5900
rect 8284 -5946 8297 -5900
rect 7745 -5959 7817 -5946
rect 7273 -6099 7329 -5959
rect 7753 -6099 7809 -5959
rect 7913 -6099 7969 -5946
rect 8073 -6099 8129 -5946
rect 8225 -5959 8297 -5946
rect 8385 -5900 8457 -5887
rect 8385 -5946 8398 -5900
rect 8444 -5946 8457 -5900
rect 8385 -5959 8457 -5946
rect 8705 -5902 8777 -5889
rect 8705 -5948 8718 -5902
rect 8764 -5948 8777 -5902
rect 8233 -6099 8289 -5959
rect 8705 -5961 8777 -5948
rect 8713 -6099 8769 -5961
rect 9001 -6099 9057 -5431
rect 879 -7243 935 -6783
rect 2543 -6805 2599 -6783
rect 2703 -6805 2759 -6783
rect 2543 -6818 2759 -6805
rect 2543 -6864 2628 -6818
rect 2674 -6864 2759 -6818
rect 2543 -6869 2759 -6864
rect 2863 -6805 2919 -6783
rect 3023 -6805 3079 -6783
rect 2863 -6818 3079 -6805
rect 2863 -6864 2948 -6818
rect 2994 -6864 3079 -6818
rect 2863 -6869 3079 -6864
rect 3183 -6803 3295 -6783
rect 3527 -6803 3639 -6783
rect 3183 -6816 3639 -6803
rect 3183 -6862 3216 -6816
rect 3262 -6862 3639 -6816
rect 2615 -6877 2687 -6869
rect 2935 -6877 3007 -6869
rect 3183 -6895 3639 -6862
rect 4039 -7243 4095 -6783
rect 1327 -7382 1399 -7374
rect 1487 -7382 1559 -7374
rect 1967 -7382 2039 -7374
rect 2607 -7382 2679 -7374
rect 1175 -7387 3935 -7382
rect 1175 -7433 1340 -7387
rect 1386 -7433 1500 -7387
rect 1546 -7433 1980 -7387
rect 2026 -7433 2620 -7387
rect 2666 -7433 3935 -7387
rect 1175 -7438 3935 -7433
rect 1327 -7446 1399 -7438
rect 1487 -7446 1559 -7438
rect 1967 -7446 2039 -7438
rect 2607 -7446 2679 -7438
rect 7433 -6319 7489 -6298
rect 7593 -6319 7649 -6299
rect 7433 -6375 7649 -6319
rect 8393 -6319 8449 -6299
rect 8553 -6319 8609 -6299
rect 8393 -6375 8609 -6319
rect 12704 -5156 12904 -5076
rect 12704 -5202 12734 -5156
rect 12780 -5202 12828 -5156
rect 12874 -5202 12904 -5156
rect 12704 -5250 12904 -5202
rect 12704 -5296 12734 -5250
rect 12780 -5296 12828 -5250
rect 12874 -5296 12904 -5250
rect 12704 -5376 12904 -5296
rect 7433 -6423 7489 -6375
rect 8393 -6423 8449 -6375
rect 7425 -6436 7497 -6423
rect 7425 -6482 7438 -6436
rect 7484 -6482 7497 -6436
rect 7425 -6495 7497 -6482
rect 8385 -6436 8457 -6423
rect 8385 -6482 8398 -6436
rect 8444 -6482 8457 -6436
rect 8385 -6495 8457 -6482
rect 9034 -6524 10146 -6508
rect 9034 -6570 9842 -6524
rect 9888 -6570 9946 -6524
rect 9992 -6570 10146 -6524
rect 6178 -6633 6250 -6625
rect 6338 -6633 6410 -6625
rect 6658 -6633 6730 -6625
rect 6818 -6633 6890 -6625
rect 6978 -6633 7050 -6625
rect 7138 -6633 7210 -6625
rect 7298 -6633 7370 -6625
rect 7458 -6633 7530 -6625
rect 7618 -6633 7690 -6625
rect 7778 -6633 7850 -6625
rect 7938 -6633 8010 -6625
rect 8098 -6633 8170 -6625
rect 8258 -6633 8330 -6625
rect 8418 -6633 8490 -6625
rect 8578 -6633 8650 -6625
rect 8738 -6633 8810 -6625
rect 6026 -6638 6562 -6633
rect 6026 -6684 6191 -6638
rect 6237 -6684 6351 -6638
rect 6397 -6684 6562 -6638
rect 6026 -6689 6562 -6684
rect 6658 -6638 8810 -6633
rect 6658 -6684 6671 -6638
rect 6717 -6684 6831 -6638
rect 6877 -6684 6991 -6638
rect 7037 -6684 7151 -6638
rect 7197 -6684 7311 -6638
rect 7357 -6684 7471 -6638
rect 7517 -6684 7631 -6638
rect 7677 -6684 7791 -6638
rect 7837 -6684 7951 -6638
rect 7997 -6684 8111 -6638
rect 8157 -6684 8271 -6638
rect 8317 -6684 8431 -6638
rect 8477 -6684 8591 -6638
rect 8637 -6684 8751 -6638
rect 8797 -6684 8810 -6638
rect 6658 -6689 8810 -6684
rect 6026 -6728 6082 -6689
rect 6178 -6697 6250 -6689
rect 6338 -6697 6410 -6689
rect 6658 -6697 6730 -6689
rect 6818 -6697 6890 -6689
rect 6978 -6697 7050 -6689
rect 7138 -6697 7210 -6689
rect 7298 -6697 7370 -6689
rect 7458 -6697 7530 -6689
rect 7618 -6697 7690 -6689
rect 7778 -6697 7850 -6689
rect 7938 -6697 8010 -6689
rect 8098 -6697 8170 -6689
rect 8258 -6697 8330 -6689
rect 8418 -6697 8490 -6689
rect 8578 -6697 8650 -6689
rect 8738 -6697 8810 -6689
rect 9034 -6628 10146 -6570
rect 9034 -6674 9842 -6628
rect 9888 -6674 9946 -6628
rect 9992 -6674 10146 -6628
rect 9034 -6708 10146 -6674
rect 9034 -6728 9234 -6708
rect 9946 -6727 10146 -6708
rect 5738 -7111 5794 -6928
rect 10250 -7111 10306 -6928
rect 5730 -7124 5802 -7111
rect 5730 -7170 5743 -7124
rect 5789 -7170 5802 -7124
rect 5730 -7183 5802 -7170
rect 10242 -7124 10314 -7111
rect 10242 -7170 10255 -7124
rect 10301 -7170 10314 -7124
rect 10242 -7183 10314 -7170
rect 5738 -7365 5794 -7183
rect 6026 -7250 7866 -7233
rect 6026 -7296 6041 -7250
rect 6087 -7296 6145 -7250
rect 6191 -7266 7866 -7250
rect 6191 -7296 7585 -7266
rect 6026 -7312 7585 -7296
rect 7631 -7312 7679 -7266
rect 7725 -7312 7773 -7266
rect 7819 -7312 7866 -7266
rect 6026 -7345 7866 -7312
rect 7970 -7275 9202 -7233
rect 7970 -7321 8271 -7275
rect 8317 -7321 8431 -7275
rect 8477 -7321 8591 -7275
rect 8637 -7321 8751 -7275
rect 8797 -7321 8911 -7275
rect 8957 -7321 9071 -7275
rect 9117 -7321 9202 -7275
rect 10250 -7289 10306 -7183
rect 7970 -7345 9202 -7321
rect 9450 -7345 10306 -7289
rect 6026 -7365 6138 -7345
rect 6242 -7365 6354 -7345
rect 6458 -7365 6570 -7345
rect 6674 -7365 6786 -7345
rect 6890 -7365 7002 -7345
rect 7106 -7365 7218 -7345
rect 7322 -7365 7434 -7345
rect 7538 -7365 7650 -7345
rect 7754 -7365 7866 -7345
rect 9450 -7365 9506 -7345
rect 10250 -7365 10306 -7345
rect 12272 -6460 12472 -5776
rect 12704 -5912 12904 -5776
rect 13008 -5912 13208 -5776
rect 13312 -5912 13512 -5776
rect 13616 -5912 13816 -5776
rect 13920 -5912 14120 -5776
rect 14224 -5912 14424 -5776
rect 14656 -5912 14856 -5776
rect 14960 -5912 15160 -5776
rect 15264 -5912 15464 -5776
rect 15568 -5912 15768 -5776
rect 15872 -5912 16072 -5776
rect 12272 -6506 12302 -6460
rect 12348 -6506 12396 -6460
rect 12442 -6506 12472 -6460
rect 12272 -6554 12472 -6506
rect 12272 -6600 12302 -6554
rect 12348 -6600 12396 -6554
rect 12442 -6600 12472 -6554
rect 13008 -6372 13208 -6312
rect 13312 -6372 13512 -6312
rect 13616 -6372 13816 -6312
rect 13920 -6372 14120 -6312
rect 14224 -6372 14424 -6312
rect 14656 -6372 14856 -6312
rect 14960 -6372 15160 -6312
rect 15264 -6372 15464 -6312
rect 15568 -6372 15768 -6312
rect 15872 -6372 16072 -6312
rect 13008 -6397 16072 -6372
rect 13008 -6443 15700 -6397
rect 15746 -6443 15804 -6397
rect 15850 -6443 15908 -6397
rect 15954 -6443 16072 -6397
rect 13008 -6449 16072 -6443
rect 13008 -6495 13143 -6449
rect 13189 -6495 13237 -6449
rect 13283 -6495 13331 -6449
rect 13377 -6495 13751 -6449
rect 13797 -6495 13845 -6449
rect 13891 -6495 13939 -6449
rect 13985 -6495 14359 -6449
rect 14405 -6495 14453 -6449
rect 14499 -6495 14547 -6449
rect 14593 -6495 16072 -6449
rect 13008 -6501 16072 -6495
rect 13008 -6547 15700 -6501
rect 15746 -6547 15804 -6501
rect 15850 -6547 15908 -6501
rect 15954 -6547 16072 -6501
rect 13008 -6572 16072 -6547
rect 16176 -6460 16376 -5776
rect 16176 -6506 16206 -6460
rect 16252 -6506 16300 -6460
rect 16346 -6506 16376 -6460
rect 16176 -6554 16376 -6506
rect 12272 -6748 12472 -6600
rect 16176 -6600 16206 -6554
rect 16252 -6600 16300 -6554
rect 16346 -6600 16376 -6554
rect 16176 -6748 16376 -6600
rect 12704 -7345 12904 -7148
rect 12704 -7391 12729 -7345
rect 12775 -7391 12833 -7345
rect 12879 -7391 12904 -7345
rect 12704 -7449 12904 -7391
rect 13008 -7248 13208 -7148
rect 13312 -7248 13512 -7148
rect 13616 -7248 13816 -7148
rect 13920 -7248 14120 -7148
rect 14224 -7248 14424 -7148
rect 14656 -7248 14856 -7148
rect 14960 -7248 15160 -7148
rect 15264 -7248 15464 -7148
rect 15568 -7248 15768 -7148
rect 15872 -7248 16072 -7148
rect 13008 -7325 16072 -7248
rect 13008 -7371 13143 -7325
rect 13189 -7371 13237 -7325
rect 13283 -7371 13331 -7325
rect 13377 -7371 13741 -7325
rect 13787 -7371 13845 -7325
rect 13891 -7371 13949 -7325
rect 13995 -7371 14359 -7325
rect 14405 -7371 14453 -7325
rect 14499 -7371 14547 -7325
rect 14593 -7371 16072 -7325
rect 13008 -7448 16072 -7371
rect 12704 -7495 12729 -7449
rect 12775 -7495 12833 -7449
rect 12879 -7495 12904 -7449
rect 12704 -7520 12904 -7495
rect 18384 -5010 18440 -4978
rect 18376 -5023 18448 -5010
rect 18376 -5069 18389 -5023
rect 18435 -5069 18448 -5023
rect 18376 -5082 18448 -5069
rect 18384 -6482 18440 -5082
rect 18376 -6495 18448 -6482
rect 18376 -6541 18389 -6495
rect 18435 -6541 18448 -6495
rect 18376 -6554 18448 -6541
rect 18384 -6586 18440 -6554
rect 18544 -6586 18600 -4978
rect 18704 -6586 18760 -4978
rect 18864 -6586 18920 -4978
rect 19024 -6586 19080 -4978
rect 19184 -6586 19240 -4978
rect 19344 -6586 19400 -4978
rect 19504 -6586 19560 -4978
rect 19664 -6586 19720 -4978
rect 19824 -6586 19880 -4978
rect 19984 -6586 20040 -4978
rect 20144 -6586 20200 -4978
rect 20304 -6586 20360 -4978
rect 20464 -6586 20520 -4978
rect 20624 -6586 20680 -4978
rect 20784 -6586 20840 -4978
rect 20944 -6586 21000 -4978
rect 21104 -6586 21160 -4978
rect 21264 -6586 21320 -4978
rect 21552 -5010 21608 -4978
rect 21840 -5010 21896 -4978
rect 21544 -5023 21616 -5010
rect 21544 -5069 21557 -5023
rect 21603 -5069 21616 -5023
rect 21544 -5082 21616 -5069
rect 21832 -5023 21904 -5010
rect 21832 -5069 21845 -5023
rect 21891 -5069 21904 -5023
rect 21832 -5082 21904 -5069
rect 21552 -5114 21608 -5082
rect 21552 -6686 21608 -6450
rect 21840 -6482 21896 -5082
rect 21832 -6495 21904 -6482
rect 21832 -6541 21845 -6495
rect 21891 -6541 21904 -6495
rect 21832 -6554 21904 -6541
rect 21840 -6586 21896 -6554
rect 21104 -7243 21160 -7186
rect 21264 -7243 21320 -7186
rect 21552 -7243 21608 -7186
rect 21104 -7256 21608 -7243
rect 21104 -7302 21160 -7256
rect 21206 -7302 21264 -7256
rect 21310 -7302 21368 -7256
rect 21414 -7302 21477 -7256
rect 21523 -7302 21608 -7256
rect 21104 -7315 21608 -7302
<< polycontact >>
rect 3479 5016 3525 5062
rect 3959 5016 4005 5062
rect 4599 5016 4645 5062
rect 3479 3888 3525 3934
rect 3639 3888 3685 3934
rect 3959 3888 4005 3934
rect 4279 3888 4325 3934
rect 4599 3888 4645 3934
rect 3479 2760 3525 2806
rect 3639 2760 3685 2806
rect 3959 2760 4005 2806
rect 4279 2760 4325 2806
rect 4599 2760 4645 2806
rect 3479 500 3525 546
rect 3639 500 3685 546
rect 3959 500 4005 546
rect 4279 500 4325 546
rect 4599 500 4645 546
rect 3191 -614 3237 -568
rect 533 -840 579 -794
rect 2477 -840 2523 -794
rect 3479 -630 3525 -584
rect 3639 -630 3685 -584
rect 3959 -630 4005 -584
rect 4279 -630 4325 -584
rect 4599 -630 4645 -584
rect 4887 -614 4933 -568
rect 756 -1623 802 -1577
rect 860 -1623 906 -1577
rect 3639 -1714 3685 -1668
rect 4279 -1714 4325 -1668
rect 18594 4199 18640 4245
rect 19074 4199 19120 4245
rect 19714 4199 19760 4245
rect 18306 3241 18352 3287
rect 18594 3233 18640 3279
rect 6056 -795 6102 -749
rect 7518 -742 7564 -696
rect 7518 -846 7564 -800
rect 7752 -795 7798 -749
rect 10251 -753 10297 -707
rect 8291 -814 8337 -768
rect 10251 -857 10297 -811
rect 10499 -814 10545 -768
rect 11917 -643 11963 -597
rect 11673 -768 11719 -722
rect 11917 -747 11963 -701
rect 13881 -768 13927 -722
rect 14703 -638 14749 -592
rect 14467 -768 14513 -722
rect 14703 -742 14749 -696
rect 16163 -768 16209 -722
rect 18754 3233 18800 3279
rect 19074 3233 19120 3279
rect 19394 3233 19440 3279
rect 19714 3233 19760 3279
rect 20002 3241 20048 3287
rect 18594 2297 18640 2343
rect 18754 2297 18800 2343
rect 19074 2297 19120 2343
rect 19394 2297 19440 2343
rect 19714 2297 19760 2343
rect 18594 425 18640 471
rect 18754 425 18800 471
rect 19074 425 19120 471
rect 19394 425 19440 471
rect 19714 425 19760 471
rect 18306 -503 18352 -457
rect 18594 -511 18640 -465
rect 18754 -511 18800 -465
rect 19074 -511 19120 -465
rect 19394 -511 19440 -465
rect 19714 -511 19760 -465
rect 20002 -503 20048 -457
rect 18754 -1447 18800 -1401
rect 19394 -1447 19440 -1401
rect 23746 4199 23792 4245
rect 24386 4199 24432 4245
rect 24866 4199 24912 4245
rect 23458 3241 23504 3287
rect 23746 3233 23792 3279
rect 24066 3233 24112 3279
rect 24386 3233 24432 3279
rect 24706 3233 24752 3279
rect 24866 3233 24912 3279
rect 25154 3241 25200 3287
rect 23746 2297 23792 2343
rect 24066 2297 24112 2343
rect 24386 2297 24432 2343
rect 24706 2297 24752 2343
rect 24866 2297 24912 2343
rect 23746 425 23792 471
rect 24066 425 24112 471
rect 24386 425 24432 471
rect 24706 425 24752 471
rect 24866 425 24912 471
rect 23458 -503 23504 -457
rect 23746 -511 23792 -465
rect 24066 -511 24112 -465
rect 24386 -511 24432 -465
rect 24706 -511 24752 -465
rect 24866 -511 24912 -465
rect 25154 -503 25200 -457
rect 24066 -1447 24112 -1401
rect 24706 -1447 24752 -1401
rect 27715 4199 27761 4245
rect 28195 4199 28241 4245
rect 28835 4199 28881 4245
rect 27427 3241 27473 3287
rect 27715 3233 27761 3279
rect 27875 3233 27921 3279
rect 28195 3233 28241 3279
rect 28515 3233 28561 3279
rect 28835 3233 28881 3279
rect 29123 3241 29169 3287
rect 27715 2297 27761 2343
rect 27875 2297 27921 2343
rect 28195 2297 28241 2343
rect 28515 2297 28561 2343
rect 28835 2297 28881 2343
rect 27715 425 27761 471
rect 27875 425 27921 471
rect 28195 425 28241 471
rect 28515 425 28561 471
rect 28835 425 28881 471
rect 27427 -503 27473 -457
rect 27715 -511 27761 -465
rect 27875 -511 27921 -465
rect 28195 -511 28241 -465
rect 28515 -511 28561 -465
rect 28835 -511 28881 -465
rect 29123 -503 29169 -457
rect 27875 -1447 27921 -1401
rect 28515 -1447 28561 -1401
rect 34131 2606 34177 2652
rect 34291 2606 34337 2652
rect 38267 2606 38313 2652
rect 38427 2606 38473 2652
rect 32723 1679 32769 1725
rect 35699 1679 35745 1725
rect 34131 1546 34177 1592
rect 34291 1546 34337 1592
rect 34131 486 34177 532
rect 34291 486 34337 532
rect 32723 -441 32769 -395
rect 36859 1679 36905 1725
rect 35699 -441 35745 -395
rect 39835 1679 39881 1725
rect 38267 1546 38313 1592
rect 38427 1546 38473 1592
rect 38267 486 38313 532
rect 38427 486 38473 532
rect 34131 -574 34177 -528
rect 34291 -574 34337 -528
rect 36859 -441 36905 -395
rect 39835 -441 39881 -395
rect 38267 -574 38313 -528
rect 38427 -574 38473 -528
rect 43827 2606 43873 2652
rect 43987 2606 44033 2652
rect 47963 2606 48009 2652
rect 48123 2606 48169 2652
rect 42419 1679 42465 1725
rect 45395 1679 45441 1725
rect 43827 1546 43873 1592
rect 43987 1546 44033 1592
rect 43827 486 43873 532
rect 43987 486 44033 532
rect 42419 -441 42465 -395
rect 46555 1679 46601 1725
rect 45395 -441 45441 -395
rect 49531 1679 49577 1725
rect 47963 1546 48009 1592
rect 48123 1546 48169 1592
rect 47963 486 48009 532
rect 48123 486 48169 532
rect 43827 -574 43873 -528
rect 43987 -574 44033 -528
rect 46555 -441 46601 -395
rect 49531 -441 49577 -395
rect 47963 -574 48009 -528
rect 48123 -574 48169 -528
rect 53523 2606 53569 2652
rect 53683 2606 53729 2652
rect 57659 2606 57705 2652
rect 57819 2606 57865 2652
rect 52115 1679 52161 1725
rect 55091 1679 55137 1725
rect 53523 1546 53569 1592
rect 53683 1546 53729 1592
rect 53523 486 53569 532
rect 53683 486 53729 532
rect 52115 -441 52161 -395
rect 56251 1679 56297 1725
rect 55091 -441 55137 -395
rect 59227 1679 59273 1725
rect 57659 1546 57705 1592
rect 57819 1546 57865 1592
rect 57659 486 57705 532
rect 57819 486 57865 532
rect 53523 -574 53569 -528
rect 53683 -574 53729 -528
rect 56251 -441 56297 -395
rect 59227 -441 59273 -395
rect 57659 -574 57705 -528
rect 57819 -574 57865 -528
rect 63219 2606 63265 2652
rect 63379 2606 63425 2652
rect 61811 1679 61857 1725
rect 64787 1679 64833 1725
rect 63219 1546 63265 1592
rect 63379 1546 63425 1592
rect 63219 486 63265 532
rect 63379 486 63425 532
rect 61811 -441 61857 -395
rect 64787 -441 64833 -395
rect 63219 -574 63265 -528
rect 63379 -574 63425 -528
rect 7278 -3269 7324 -3223
rect 7758 -3269 7804 -3223
rect 8238 -3269 8284 -3223
rect 8718 -3268 8764 -3222
rect 1172 -4688 1218 -4642
rect 1704 -4650 1750 -4604
rect 1808 -4650 1854 -4604
rect 3836 -4690 3882 -4644
rect 3996 -4690 4042 -4644
rect 1616 -5862 1662 -5816
rect 1720 -5862 1766 -5816
rect 1824 -5862 1870 -5816
rect 1928 -5862 1974 -5816
rect 2032 -5862 2078 -5816
rect 2136 -5862 2182 -5816
rect 884 -5948 930 -5902
rect 1180 -5948 1226 -5902
rect 3748 -5939 3794 -5893
rect 4044 -5939 4090 -5893
rect 7278 -3819 7324 -3773
rect 7438 -3819 7484 -3773
rect 7758 -3819 7804 -3773
rect 8238 -3819 8284 -3773
rect 8398 -3819 8444 -3773
rect 8718 -3819 8764 -3773
rect 7278 -4340 7324 -4294
rect 7438 -4340 7484 -4294
rect 7758 -4340 7804 -4294
rect 8238 -4340 8284 -4294
rect 8398 -4340 8444 -4294
rect 8718 -4340 8764 -4294
rect 7278 -4874 7324 -4828
rect 7438 -4874 7484 -4828
rect 7758 -4874 7804 -4828
rect 8238 -4874 8284 -4828
rect 8398 -4874 8444 -4828
rect 8718 -4874 8764 -4828
rect 6990 -5418 7036 -5372
rect 7278 -5410 7324 -5364
rect 7438 -5410 7484 -5364
rect 7758 -5410 7804 -5364
rect 8238 -5410 8284 -5364
rect 8398 -5410 8444 -5364
rect 20176 -4288 20222 -4242
rect 20280 -4288 20326 -4242
rect 20869 -4288 20915 -4242
rect 8718 -5412 8764 -5366
rect 9006 -5418 9052 -5372
rect 7278 -5946 7324 -5900
rect 7438 -5946 7484 -5900
rect 7758 -5946 7804 -5900
rect 8238 -5946 8284 -5900
rect 8398 -5946 8444 -5900
rect 8718 -5948 8764 -5902
rect 2628 -6864 2674 -6818
rect 2948 -6864 2994 -6818
rect 3216 -6862 3262 -6816
rect 1340 -7433 1386 -7387
rect 1500 -7433 1546 -7387
rect 1980 -7433 2026 -7387
rect 2620 -7433 2666 -7387
rect 12734 -5202 12780 -5156
rect 12828 -5202 12874 -5156
rect 12734 -5296 12780 -5250
rect 12828 -5296 12874 -5250
rect 7438 -6482 7484 -6436
rect 8398 -6482 8444 -6436
rect 9842 -6570 9888 -6524
rect 9946 -6570 9992 -6524
rect 6191 -6684 6237 -6638
rect 6351 -6684 6397 -6638
rect 6671 -6684 6717 -6638
rect 6831 -6684 6877 -6638
rect 6991 -6684 7037 -6638
rect 7151 -6684 7197 -6638
rect 7311 -6684 7357 -6638
rect 7471 -6684 7517 -6638
rect 7631 -6684 7677 -6638
rect 7791 -6684 7837 -6638
rect 7951 -6684 7997 -6638
rect 8111 -6684 8157 -6638
rect 8271 -6684 8317 -6638
rect 8431 -6684 8477 -6638
rect 8591 -6684 8637 -6638
rect 8751 -6684 8797 -6638
rect 9842 -6674 9888 -6628
rect 9946 -6674 9992 -6628
rect 5743 -7170 5789 -7124
rect 10255 -7170 10301 -7124
rect 6041 -7296 6087 -7250
rect 6145 -7296 6191 -7250
rect 7585 -7312 7631 -7266
rect 7679 -7312 7725 -7266
rect 7773 -7312 7819 -7266
rect 8271 -7321 8317 -7275
rect 8431 -7321 8477 -7275
rect 8591 -7321 8637 -7275
rect 8751 -7321 8797 -7275
rect 8911 -7321 8957 -7275
rect 9071 -7321 9117 -7275
rect 12302 -6506 12348 -6460
rect 12396 -6506 12442 -6460
rect 12302 -6600 12348 -6554
rect 12396 -6600 12442 -6554
rect 15700 -6443 15746 -6397
rect 15804 -6443 15850 -6397
rect 15908 -6443 15954 -6397
rect 13143 -6495 13189 -6449
rect 13237 -6495 13283 -6449
rect 13331 -6495 13377 -6449
rect 13751 -6495 13797 -6449
rect 13845 -6495 13891 -6449
rect 13939 -6495 13985 -6449
rect 14359 -6495 14405 -6449
rect 14453 -6495 14499 -6449
rect 14547 -6495 14593 -6449
rect 15700 -6547 15746 -6501
rect 15804 -6547 15850 -6501
rect 15908 -6547 15954 -6501
rect 16206 -6506 16252 -6460
rect 16300 -6506 16346 -6460
rect 16206 -6600 16252 -6554
rect 16300 -6600 16346 -6554
rect 12729 -7391 12775 -7345
rect 12833 -7391 12879 -7345
rect 13143 -7371 13189 -7325
rect 13237 -7371 13283 -7325
rect 13331 -7371 13377 -7325
rect 13741 -7371 13787 -7325
rect 13845 -7371 13891 -7325
rect 13949 -7371 13995 -7325
rect 14359 -7371 14405 -7325
rect 14453 -7371 14499 -7325
rect 14547 -7371 14593 -7325
rect 12729 -7495 12775 -7449
rect 12833 -7495 12879 -7449
rect 18389 -5069 18435 -5023
rect 18389 -6541 18435 -6495
rect 21557 -5069 21603 -5023
rect 21845 -5069 21891 -5023
rect 21845 -6541 21891 -6495
rect 21160 -7302 21206 -7256
rect 21264 -7302 21310 -7256
rect 21368 -7302 21414 -7256
rect 21477 -7302 21523 -7256
<< metal1 >>
rect 30732 6548 31516 6560
rect 30732 6496 30744 6548
rect 30796 6496 30848 6548
rect 30900 6496 30952 6548
rect 31004 6496 31516 6548
rect 30732 6444 31516 6496
rect 30732 6392 30744 6444
rect 30796 6392 30848 6444
rect 30900 6392 30952 6444
rect 31004 6392 31516 6444
rect 30732 6340 31516 6392
rect 30732 6288 30744 6340
rect 30796 6288 30848 6340
rect 30900 6288 30952 6340
rect 31004 6288 31516 6340
rect 30732 6276 31516 6288
rect 31646 5962 32430 5974
rect 31646 5910 31658 5962
rect 31710 5910 31762 5962
rect 31814 5910 31866 5962
rect 31918 5910 32430 5962
rect 31646 5858 32430 5910
rect 31646 5806 31658 5858
rect 31710 5806 31762 5858
rect 31814 5806 31866 5858
rect 31918 5806 32430 5858
rect 31646 5754 32430 5806
rect 31646 5702 31658 5754
rect 31710 5702 31762 5754
rect 31814 5702 31866 5754
rect 31918 5702 32430 5754
rect 31646 5690 32430 5702
rect 5743 5508 29906 5565
rect 5743 5462 5776 5508
rect 5822 5462 5870 5508
rect 5916 5462 5964 5508
rect 6010 5462 6058 5508
rect 6104 5462 6152 5508
rect 6198 5462 6246 5508
rect 6292 5462 6340 5508
rect 6386 5462 6434 5508
rect 6480 5462 6528 5508
rect 6574 5462 6622 5508
rect 6668 5462 6716 5508
rect 6762 5462 6810 5508
rect 6856 5462 6904 5508
rect 6950 5462 6998 5508
rect 7044 5462 7092 5508
rect 7138 5462 7186 5508
rect 7232 5462 7280 5508
rect 7326 5462 7374 5508
rect 7420 5462 7468 5508
rect 7514 5462 7562 5508
rect 7608 5462 7656 5508
rect 7702 5462 7750 5508
rect 7796 5462 7844 5508
rect 7890 5462 7938 5508
rect 7984 5462 8032 5508
rect 8078 5462 29906 5508
rect 5743 5414 29906 5462
rect 5743 5368 5776 5414
rect 5822 5405 8032 5414
rect 5822 5368 5855 5405
rect 5743 5320 5855 5368
rect 2925 5217 5199 5284
rect -1790 5190 -1465 5201
rect -1790 5134 -1781 5190
rect -1725 5134 -1671 5190
rect -1615 5134 -1561 5190
rect -1505 5171 -1465 5190
rect 2675 5171 2855 5181
rect -1505 5169 2855 5171
rect -1505 5134 2687 5169
rect -1790 5117 2687 5134
rect 2739 5117 2791 5169
rect 2843 5117 2855 5169
rect -1790 5080 2855 5117
rect -1790 5024 -1781 5080
rect -1725 5024 -1671 5080
rect -1615 5024 -1561 5080
rect -1505 5065 2855 5080
rect -1505 5024 2687 5065
rect -1790 5013 2687 5024
rect 2739 5013 2791 5065
rect 2843 5013 2855 5065
rect -1790 5011 2855 5013
rect 2675 5001 2855 5011
rect 2925 5171 2958 5217
rect 3004 5171 3052 5217
rect 3098 5171 3146 5217
rect 3192 5171 3240 5217
rect 3286 5171 3334 5217
rect 3380 5171 3428 5217
rect 3474 5171 3522 5217
rect 3568 5171 3616 5217
rect 3662 5171 3710 5217
rect 3756 5171 3804 5217
rect 3850 5171 3898 5217
rect 3944 5171 3992 5217
rect 4038 5171 4086 5217
rect 4132 5171 4180 5217
rect 4226 5171 4274 5217
rect 4320 5171 4368 5217
rect 4414 5171 4462 5217
rect 4508 5171 4556 5217
rect 4602 5171 4650 5217
rect 4696 5171 4744 5217
rect 4790 5171 4838 5217
rect 4884 5171 4932 5217
rect 4978 5171 5026 5217
rect 5072 5171 5120 5217
rect 5166 5171 5199 5217
rect 2925 5124 5199 5171
rect 5255 5127 5415 5317
rect 2925 5123 3037 5124
rect 2925 5077 2958 5123
rect 3004 5077 3037 5123
rect 2925 5029 3037 5077
rect 2925 4983 2958 5029
rect 3004 4983 3037 5029
rect 2925 4935 3037 4983
rect 2925 4889 2958 4935
rect 3004 4889 3037 4935
rect 2925 4841 3037 4889
rect 3111 4856 3157 5124
rect 3271 4856 3317 5124
rect 3464 5065 3540 5077
rect 3464 5013 3476 5065
rect 3528 5062 3540 5065
rect 3528 5016 3959 5062
rect 4005 5016 4599 5062
rect 4645 5016 4656 5062
rect 3528 5013 3540 5016
rect 3464 5001 3540 5013
rect 3559 4913 4565 4959
rect 3559 4856 3605 4913
rect 3879 4856 3925 4913
rect 4199 4856 4245 4913
rect 4519 4856 4565 4913
rect 4807 4856 4853 5124
rect 4967 4856 5013 5124
rect 5087 5123 5199 5124
rect 5087 5077 5120 5123
rect 5166 5077 5199 5123
rect 5087 5029 5199 5077
rect 5087 4983 5120 5029
rect 5166 4983 5199 5029
rect 5087 4935 5199 4983
rect 5245 5115 5425 5127
rect 5245 5063 5257 5115
rect 5309 5063 5361 5115
rect 5413 5063 5425 5115
rect 5245 5011 5425 5063
rect 5245 4959 5257 5011
rect 5309 4959 5361 5011
rect 5413 4959 5425 5011
rect 5245 4947 5425 4959
rect 5087 4889 5120 4935
rect 5166 4889 5199 4935
rect 2034 4822 2214 4832
rect 1852 4820 2214 4822
rect 1852 4768 2046 4820
rect 2098 4768 2150 4820
rect 2202 4768 2214 4820
rect 1852 4716 2214 4768
rect 1852 4664 2046 4716
rect 2098 4664 2150 4716
rect 2202 4664 2214 4716
rect 1852 4662 2214 4664
rect 2034 4652 2214 4662
rect 2925 4795 2958 4841
rect 3004 4795 3037 4841
rect 5087 4841 5199 4889
rect 2925 4747 3037 4795
rect 2925 4701 2958 4747
rect 3004 4701 3037 4747
rect 2925 4653 3037 4701
rect 2925 4607 2958 4653
rect 3004 4607 3037 4653
rect 3544 4820 3620 4832
rect 3544 4768 3556 4820
rect 3608 4768 3620 4820
rect 3544 4716 3620 4768
rect 3544 4664 3556 4716
rect 3608 4664 3620 4716
rect 3544 4652 3620 4664
rect 3704 4820 3780 4832
rect 3704 4768 3716 4820
rect 3768 4768 3780 4820
rect 3704 4716 3780 4768
rect 3704 4664 3716 4716
rect 3768 4664 3780 4716
rect 3704 4652 3780 4664
rect 4345 4820 4421 4832
rect 4345 4768 4357 4820
rect 4409 4768 4421 4820
rect 4345 4716 4421 4768
rect 4345 4664 4357 4716
rect 4409 4664 4421 4716
rect 4345 4652 4421 4664
rect 5087 4795 5120 4841
rect 5166 4795 5199 4841
rect 5527 4832 5687 5307
rect 5743 5274 5776 5320
rect 5822 5274 5855 5320
rect 5743 5226 5855 5274
rect 5743 5180 5776 5226
rect 5822 5180 5855 5226
rect 5743 5132 5855 5180
rect 5743 5086 5776 5132
rect 5822 5086 5855 5132
rect 5976 5106 6022 5405
rect 6136 5106 6182 5405
rect 6249 5115 6325 5127
rect 5743 5038 5855 5086
rect 5743 4992 5776 5038
rect 5822 4992 5855 5038
rect 5743 4944 5855 4992
rect 6249 5063 6261 5115
rect 6313 5063 6325 5115
rect 6424 5106 6470 5405
rect 6744 5106 6790 5405
rect 6889 5115 6965 5127
rect 6249 5011 6325 5063
rect 6249 4959 6261 5011
rect 6313 4959 6325 5011
rect 6249 4947 6325 4959
rect 6889 5063 6901 5115
rect 6953 5063 6965 5115
rect 7064 5106 7110 5405
rect 7384 5106 7430 5405
rect 7529 5115 7605 5127
rect 6889 5011 6965 5063
rect 6889 4959 6901 5011
rect 6953 4959 6965 5011
rect 6889 4947 6965 4959
rect 7529 5063 7541 5115
rect 7593 5063 7605 5115
rect 7672 5106 7718 5405
rect 7832 5106 7878 5405
rect 7999 5368 8032 5405
rect 8078 5368 29906 5414
rect 7999 5320 29906 5368
rect 7999 5274 8032 5320
rect 8078 5274 29906 5320
rect 7999 5245 29906 5274
rect 7999 5226 8159 5245
rect 7999 5180 8032 5226
rect 8078 5180 8159 5226
rect 7999 5132 8159 5180
rect 7529 5011 7605 5063
rect 7529 4959 7541 5011
rect 7593 4959 7605 5011
rect 7529 4947 7605 4959
rect 7999 5086 8032 5132
rect 8078 5086 8159 5132
rect 7999 5038 8159 5086
rect 7999 4992 8032 5038
rect 8078 4992 8159 5038
rect 5743 4898 5776 4944
rect 5822 4898 5855 4944
rect 5743 4850 5855 4898
rect 5087 4747 5199 4795
rect 5087 4701 5120 4747
rect 5166 4701 5199 4747
rect 5087 4653 5199 4701
rect 2925 4559 3037 4607
rect 2925 4513 2958 4559
rect 3004 4513 3037 4559
rect 2925 4465 3037 4513
rect 2925 4419 2958 4465
rect 3004 4419 3037 4465
rect 2925 4371 3037 4419
rect 2925 4325 2958 4371
rect 3004 4325 3037 4371
rect 5087 4607 5120 4653
rect 5166 4607 5199 4653
rect 5517 4820 5697 4832
rect 5517 4768 5529 4820
rect 5581 4768 5633 4820
rect 5685 4768 5697 4820
rect 5517 4716 5697 4768
rect 5517 4664 5529 4716
rect 5581 4664 5633 4716
rect 5685 4664 5697 4716
rect 5517 4652 5697 4664
rect 5743 4804 5776 4850
rect 5822 4804 5855 4850
rect 7999 4944 8159 4992
rect 7999 4898 8032 4944
rect 8078 4898 8159 4944
rect 7999 4850 8159 4898
rect 5743 4756 5855 4804
rect 5743 4710 5776 4756
rect 5822 4710 5855 4756
rect 5743 4662 5855 4710
rect 5087 4559 5199 4607
rect 5087 4513 5120 4559
rect 5166 4513 5199 4559
rect 5087 4465 5199 4513
rect 5087 4419 5120 4465
rect 5166 4419 5199 4465
rect 5087 4371 5199 4419
rect 2925 4277 3037 4325
rect 2925 4231 2958 4277
rect 3004 4231 3037 4277
rect 2925 4183 3037 4231
rect 2925 4137 2958 4183
rect 3004 4137 3037 4183
rect 3384 4324 3460 4336
rect 3384 4272 3396 4324
rect 3448 4272 3460 4324
rect 3384 4220 3460 4272
rect 3384 4168 3396 4220
rect 3448 4168 3460 4220
rect 3384 4156 3460 4168
rect 4024 4324 4100 4336
rect 4024 4272 4036 4324
rect 4088 4272 4100 4324
rect 4024 4220 4100 4272
rect 4024 4168 4036 4220
rect 4088 4168 4100 4220
rect 4024 4156 4100 4168
rect 4664 4324 4740 4336
rect 4664 4272 4676 4324
rect 4728 4272 4740 4324
rect 4664 4220 4740 4272
rect 4664 4168 4676 4220
rect 4728 4168 4740 4220
rect 4664 4156 4740 4168
rect 5087 4325 5120 4371
rect 5166 4325 5199 4371
rect 5087 4277 5199 4325
rect 5087 4231 5120 4277
rect 5166 4231 5199 4277
rect 5087 4183 5199 4231
rect 2925 4089 3037 4137
rect 5087 4137 5120 4183
rect 5166 4137 5199 4183
rect 2395 4043 2575 4053
rect -1117 4041 2575 4043
rect -1117 4032 2407 4041
rect -1117 3976 -1106 4032
rect -1050 3976 -996 4032
rect -940 3976 -886 4032
rect -830 3989 2407 4032
rect 2459 3989 2511 4041
rect 2563 3989 2575 4041
rect -830 3976 2575 3989
rect -1117 3937 2575 3976
rect -1117 3922 2407 3937
rect -1117 3883 -1106 3922
rect -1115 3866 -1106 3883
rect -1050 3866 -996 3922
rect -940 3866 -886 3922
rect -830 3885 2407 3922
rect 2459 3885 2511 3937
rect 2563 3885 2575 3937
rect -830 3883 2575 3885
rect -830 3866 -789 3883
rect 2395 3873 2575 3883
rect 2925 4043 2958 4089
rect 3004 4043 3037 4089
rect 2925 3995 3037 4043
rect 2925 3949 2958 3995
rect 3004 3949 3037 3995
rect 2925 3901 3037 3949
rect -1115 3853 -789 3866
rect 2925 3855 2958 3901
rect 3004 3855 3037 3901
rect 2925 3807 3037 3855
rect 2925 3761 2958 3807
rect 3004 3761 3037 3807
rect 2925 3713 3037 3761
rect 3111 3726 3157 4132
rect 3271 3726 3317 4132
rect 3464 4041 3540 4053
rect 3464 3989 3476 4041
rect 3528 3989 3540 4041
rect 3464 3937 3540 3989
rect 3464 3885 3476 3937
rect 3528 3934 3540 3937
rect 3528 3888 3639 3934
rect 3685 3888 3959 3934
rect 4005 3888 4279 3934
rect 4325 3888 4599 3934
rect 4645 3888 4656 3934
rect 3528 3885 3540 3888
rect 3464 3873 3540 3885
rect 3559 3783 4565 3829
rect 3559 3726 3605 3783
rect 3879 3726 3925 3783
rect 4199 3726 4245 3783
rect 4519 3726 4565 3783
rect 4807 3726 4853 4132
rect 4967 3726 5013 4132
rect 5087 4089 5199 4137
rect 5087 4043 5120 4089
rect 5166 4043 5199 4089
rect 5087 3995 5199 4043
rect 5087 3949 5120 3995
rect 5166 3949 5199 3995
rect 5087 3901 5199 3949
rect 5087 3855 5120 3901
rect 5166 3855 5199 3901
rect 5087 3807 5199 3855
rect 5087 3761 5120 3807
rect 5166 3761 5199 3807
rect 2925 3667 2958 3713
rect 3004 3667 3037 3713
rect 5087 3713 5199 3761
rect 2925 3619 3037 3667
rect 2925 3573 2958 3619
rect 3004 3573 3037 3619
rect 2925 3525 3037 3573
rect 2925 3479 2958 3525
rect 3004 3479 3037 3525
rect 3544 3690 3620 3702
rect 3544 3638 3556 3690
rect 3608 3638 3620 3690
rect 3544 3586 3620 3638
rect 3544 3534 3556 3586
rect 3608 3534 3620 3586
rect 3544 3522 3620 3534
rect 3704 3690 3780 3702
rect 3704 3638 3716 3690
rect 3768 3638 3780 3690
rect 3704 3586 3780 3638
rect 3704 3534 3716 3586
rect 3768 3534 3780 3586
rect 3704 3522 3780 3534
rect 4345 3690 4421 3702
rect 4345 3638 4357 3690
rect 4409 3638 4421 3690
rect 4345 3586 4421 3638
rect 4345 3534 4357 3586
rect 4409 3534 4421 3586
rect 4345 3522 4421 3534
rect 5087 3667 5120 3713
rect 5166 3667 5199 3713
rect 5087 3619 5199 3667
rect 5087 3573 5120 3619
rect 5166 3573 5199 3619
rect 5087 3525 5199 3573
rect 2925 3431 3037 3479
rect 2925 3385 2958 3431
rect 3004 3385 3037 3431
rect 2925 3337 3037 3385
rect 2925 3291 2958 3337
rect 3004 3291 3037 3337
rect 5087 3479 5120 3525
rect 5166 3479 5199 3525
rect 5087 3431 5199 3479
rect 5087 3385 5120 3431
rect 5166 3385 5199 3431
rect 5087 3337 5199 3385
rect 2925 3243 3037 3291
rect 2925 3197 2958 3243
rect 3004 3197 3037 3243
rect 2925 3149 3037 3197
rect 2925 3103 2958 3149
rect 3004 3103 3037 3149
rect 3384 3298 3460 3310
rect 3384 3246 3396 3298
rect 3448 3246 3460 3298
rect 3384 3194 3460 3246
rect 3384 3142 3396 3194
rect 3448 3142 3460 3194
rect 3384 3130 3460 3142
rect 4024 3298 4100 3310
rect 4024 3246 4036 3298
rect 4088 3246 4100 3298
rect 4024 3194 4100 3246
rect 4024 3142 4036 3194
rect 4088 3142 4100 3194
rect 4024 3130 4100 3142
rect 4664 3298 4740 3310
rect 4664 3246 4676 3298
rect 4728 3246 4740 3298
rect 4664 3194 4740 3246
rect 4664 3142 4676 3194
rect 4728 3142 4740 3194
rect 4664 3130 4740 3142
rect 5087 3291 5120 3337
rect 5166 3291 5199 3337
rect 5087 3243 5199 3291
rect 5087 3197 5120 3243
rect 5166 3197 5199 3243
rect 5087 3149 5199 3197
rect 2925 3055 3037 3103
rect 2925 3009 2958 3055
rect 3004 3009 3037 3055
rect 2925 2961 3037 3009
rect 5087 3103 5120 3149
rect 5166 3103 5199 3149
rect 5087 3055 5199 3103
rect 5087 3009 5120 3055
rect 5166 3009 5199 3055
rect 2925 2915 2958 2961
rect 3004 2915 3037 2961
rect 2925 2867 3037 2915
rect 2925 2821 2958 2867
rect 3004 2821 3037 2867
rect 2925 2773 3037 2821
rect 2925 2727 2958 2773
rect 3004 2727 3037 2773
rect 2925 2679 3037 2727
rect 2925 2633 2958 2679
rect 3004 2633 3037 2679
rect 2925 2585 3037 2633
rect 3111 2596 3157 3002
rect 3271 2596 3317 3002
rect 3464 2911 3540 2923
rect 3464 2859 3476 2911
rect 3528 2859 3540 2911
rect 3464 2807 3540 2859
rect 3464 2755 3476 2807
rect 3528 2806 3540 2807
rect 3528 2760 3639 2806
rect 3685 2760 3959 2806
rect 4005 2760 4279 2806
rect 4325 2760 4599 2806
rect 4645 2760 4656 2806
rect 3528 2755 3540 2760
rect 3464 2743 3540 2755
rect 3559 2653 4565 2699
rect 3559 2596 3605 2653
rect 3719 2596 3765 2607
rect 3879 2596 3925 2653
rect 4039 2596 4085 2607
rect 4199 2596 4245 2653
rect 4359 2596 4405 2607
rect 4519 2596 4565 2653
rect 4807 2596 4853 3002
rect 4967 2596 5013 3002
rect 5087 2961 5199 3009
rect 5087 2915 5120 2961
rect 5166 2915 5199 2961
rect 5087 2867 5199 2915
rect 5087 2821 5120 2867
rect 5166 2821 5199 2867
rect 5087 2773 5199 2821
rect 5087 2727 5120 2773
rect 5166 2727 5199 2773
rect 5087 2679 5199 2727
rect 5087 2633 5120 2679
rect 5166 2633 5199 2679
rect 2925 2539 2958 2585
rect 3004 2539 3037 2585
rect 5087 2585 5199 2633
rect 2925 2491 3037 2539
rect 2925 2445 2958 2491
rect 3004 2445 3037 2491
rect 2925 2397 3037 2445
rect 2925 2351 2958 2397
rect 3004 2351 3037 2397
rect 3704 2560 3780 2572
rect 3704 2508 3716 2560
rect 3768 2508 3780 2560
rect 3704 2456 3780 2508
rect 3704 2404 3716 2456
rect 3768 2404 3780 2456
rect 3704 2392 3780 2404
rect 4345 2560 4421 2572
rect 4345 2508 4357 2560
rect 4409 2508 4421 2560
rect 4345 2456 4421 2508
rect 4345 2404 4357 2456
rect 4409 2404 4421 2456
rect 4345 2392 4421 2404
rect 5087 2539 5120 2585
rect 5166 2539 5199 2585
rect 5087 2491 5199 2539
rect 5087 2445 5120 2491
rect 5166 2445 5199 2491
rect 5087 2397 5199 2445
rect 2925 2303 3037 2351
rect 2925 2257 2958 2303
rect 3004 2257 3037 2303
rect 2925 2209 3037 2257
rect 2925 2163 2958 2209
rect 3004 2163 3037 2209
rect 2925 2115 3037 2163
rect 2925 2069 2958 2115
rect 3004 2069 3037 2115
rect 5087 2351 5120 2397
rect 5166 2351 5199 2397
rect 5087 2303 5199 2351
rect 5087 2257 5120 2303
rect 5166 2257 5199 2303
rect 5087 2209 5199 2257
rect 5087 2163 5120 2209
rect 5166 2163 5199 2209
rect 5087 2115 5199 2163
rect 2925 2021 3037 2069
rect 2925 1975 2958 2021
rect 3004 1975 3037 2021
rect 2925 1927 3037 1975
rect 2925 1881 2958 1927
rect 3004 1881 3037 1927
rect 3384 2064 3460 2076
rect 3384 2012 3396 2064
rect 3448 2012 3460 2064
rect 3384 1960 3460 2012
rect 3384 1908 3396 1960
rect 3448 1908 3460 1960
rect 3384 1896 3460 1908
rect 4024 2064 4100 2076
rect 4024 2012 4036 2064
rect 4088 2012 4100 2064
rect 4024 1960 4100 2012
rect 4024 1908 4036 1960
rect 4088 1908 4100 1960
rect 4024 1896 4100 1908
rect 4664 2064 4740 2076
rect 4664 2012 4676 2064
rect 4728 2012 4740 2064
rect 4664 1960 4740 2012
rect 4664 1908 4676 1960
rect 4728 1908 4740 1960
rect 4664 1896 4740 1908
rect 5087 2069 5120 2115
rect 5166 2069 5199 2115
rect 5087 2021 5199 2069
rect 5087 1975 5120 2021
rect 5166 1975 5199 2021
rect 5087 1927 5199 1975
rect 2925 1833 3037 1881
rect 5087 1881 5120 1927
rect 5166 1881 5199 1927
rect 2925 1796 2958 1833
rect 11 1787 2958 1796
rect 3004 1787 3037 1833
rect 11 1739 3037 1787
rect 11 1693 44 1739
rect 90 1693 138 1739
rect 184 1693 232 1739
rect 278 1693 326 1739
rect 372 1693 420 1739
rect 466 1693 514 1739
rect 560 1693 608 1739
rect 654 1693 702 1739
rect 748 1693 796 1739
rect 842 1693 890 1739
rect 936 1693 984 1739
rect 1030 1693 1078 1739
rect 1124 1693 1172 1739
rect 1218 1693 1266 1739
rect 1312 1693 1360 1739
rect 1406 1693 1454 1739
rect 1500 1693 1548 1739
rect 1594 1693 1642 1739
rect 1688 1693 1736 1739
rect 1782 1693 1830 1739
rect 1876 1693 1924 1739
rect 1970 1693 2018 1739
rect 2064 1693 2112 1739
rect 2158 1693 2206 1739
rect 2252 1693 2300 1739
rect 2346 1693 2394 1739
rect 2440 1693 2488 1739
rect 2534 1693 2582 1739
rect 2628 1693 2676 1739
rect 2722 1693 2770 1739
rect 2816 1693 2864 1739
rect 2910 1693 2958 1739
rect 3004 1693 3037 1739
rect 11 1645 3037 1693
rect 11 1599 44 1645
rect 90 1636 2958 1645
rect 90 1599 123 1636
rect 11 1551 123 1599
rect 11 1505 44 1551
rect 90 1505 123 1551
rect 11 1457 123 1505
rect 11 1411 44 1457
rect 90 1411 123 1457
rect 11 1363 123 1411
rect 425 1388 471 1636
rect 641 1388 687 1636
rect 857 1445 2199 1491
rect 857 1388 903 1445
rect 1289 1388 1335 1445
rect 1721 1388 1767 1445
rect 2153 1388 2199 1445
rect 2369 1388 2415 1636
rect 2585 1388 2631 1636
rect 2925 1599 2958 1636
rect 3004 1599 3037 1645
rect 2925 1551 3037 1599
rect 2925 1505 2958 1551
rect 3004 1505 3037 1551
rect 2925 1457 3037 1505
rect 3111 1466 3157 1872
rect 3271 1466 3317 1872
rect 3399 1466 3445 1872
rect 3559 1466 3605 1872
rect 3719 1466 3765 1872
rect 3879 1466 3925 1872
rect 4039 1466 4085 1872
rect 4199 1466 4245 1872
rect 4359 1466 4405 1872
rect 4519 1466 4565 1872
rect 4679 1466 4725 1872
rect 4807 1466 4853 1872
rect 4967 1466 5013 1872
rect 5087 1833 5199 1881
rect 5087 1787 5120 1833
rect 5166 1787 5199 1833
rect 5087 1739 5199 1787
rect 5087 1693 5120 1739
rect 5166 1693 5199 1739
rect 5087 1645 5199 1693
rect 5087 1599 5120 1645
rect 5166 1599 5199 1645
rect 5087 1551 5199 1599
rect 5087 1505 5120 1551
rect 5166 1505 5199 1551
rect 2925 1411 2958 1457
rect 3004 1411 3037 1457
rect 11 1317 44 1363
rect 90 1317 123 1363
rect 11 1269 123 1317
rect 11 1223 44 1269
rect 90 1223 123 1269
rect 11 1175 123 1223
rect 2925 1363 3037 1411
rect 2925 1317 2958 1363
rect 3004 1317 3037 1363
rect 2925 1269 3037 1317
rect 2925 1223 2958 1269
rect 3004 1223 3037 1269
rect 11 1129 44 1175
rect 90 1129 123 1175
rect 11 1081 123 1129
rect 11 1035 44 1081
rect 90 1035 123 1081
rect 11 987 123 1035
rect 2034 1166 2214 1178
rect 2034 1114 2046 1166
rect 2098 1114 2150 1166
rect 2202 1114 2214 1166
rect 2034 1062 2214 1114
rect 2034 1010 2046 1062
rect 2098 1010 2150 1062
rect 2202 1010 2214 1062
rect 2034 998 2214 1010
rect 2925 1175 3037 1223
rect 5087 1457 5199 1505
rect 5087 1411 5120 1457
rect 5166 1411 5199 1457
rect 5087 1363 5199 1411
rect 5087 1317 5120 1363
rect 5166 1317 5199 1363
rect 5087 1269 5199 1317
rect 5087 1223 5120 1269
rect 5166 1223 5199 1269
rect 2925 1129 2958 1175
rect 3004 1129 3037 1175
rect 2925 1081 3037 1129
rect 2925 1035 2958 1081
rect 3004 1035 3037 1081
rect 11 941 44 987
rect 90 941 123 987
rect 11 893 123 941
rect 11 847 44 893
rect 90 847 123 893
rect 11 799 123 847
rect 11 753 44 799
rect 90 753 123 799
rect 2925 987 3037 1035
rect 3544 1166 3620 1178
rect 3544 1114 3556 1166
rect 3608 1114 3620 1166
rect 3544 1062 3620 1114
rect 3544 1010 3556 1062
rect 3608 1010 3620 1062
rect 3544 998 3620 1010
rect 5087 1175 5199 1223
rect 5087 1129 5120 1175
rect 5166 1129 5199 1175
rect 5087 1081 5199 1129
rect 5087 1035 5120 1081
rect 5166 1035 5199 1081
rect 2925 941 2958 987
rect 3004 941 3037 987
rect 2925 893 3037 941
rect 2925 847 2958 893
rect 3004 847 3037 893
rect 2925 799 3037 847
rect 11 705 123 753
rect 11 659 44 705
rect 90 659 123 705
rect 11 611 123 659
rect 425 626 471 788
rect 641 626 687 788
rect 857 626 903 788
rect 1073 626 1119 788
rect 1289 626 1335 788
rect 1505 626 1551 788
rect 1721 626 1767 788
rect 1937 626 1983 788
rect 2153 626 2199 788
rect 2369 626 2415 788
rect 2585 626 2631 788
rect 2925 753 2958 799
rect 3004 753 3037 799
rect 2925 705 3037 753
rect 5087 987 5199 1035
rect 5087 941 5120 987
rect 5166 941 5199 987
rect 5087 893 5199 941
rect 5087 847 5120 893
rect 5166 847 5199 893
rect 5087 799 5199 847
rect 5087 753 5120 799
rect 5166 753 5199 799
rect 2925 659 2958 705
rect 3004 659 3037 705
rect 11 565 44 611
rect 90 565 123 611
rect 11 517 123 565
rect 11 471 44 517
rect 90 471 123 517
rect 11 423 123 471
rect 11 377 44 423
rect 90 377 123 423
rect 11 329 123 377
rect 11 283 44 329
rect 90 283 123 329
rect 2925 611 3037 659
rect 2925 565 2958 611
rect 3004 565 3037 611
rect 2925 517 3037 565
rect 2925 471 2958 517
rect 3004 471 3037 517
rect 2925 423 3037 471
rect 2925 377 2958 423
rect 3004 377 3037 423
rect 2925 329 3037 377
rect 3111 336 3157 742
rect 3271 336 3317 742
rect 3464 653 3540 665
rect 3464 601 3476 653
rect 3528 601 3540 653
rect 3464 549 3540 601
rect 3464 497 3476 549
rect 3528 546 3540 549
rect 3528 500 3639 546
rect 3685 500 3959 546
rect 4005 500 4279 546
rect 4325 500 4599 546
rect 4645 500 4656 546
rect 3528 497 3540 500
rect 3464 483 3540 497
rect 3559 393 4565 439
rect 3559 336 3605 393
rect 3719 336 3765 347
rect 3879 336 3925 393
rect 4039 336 4085 347
rect 4199 336 4245 393
rect 4359 336 4405 347
rect 4519 336 4565 393
rect 4807 336 4853 742
rect 4967 336 5013 742
rect 5087 705 5199 753
rect 5087 659 5120 705
rect 5166 659 5199 705
rect 5087 611 5199 659
rect 5087 565 5120 611
rect 5166 565 5199 611
rect 5087 517 5199 565
rect 5087 471 5120 517
rect 5166 471 5199 517
rect 5087 423 5199 471
rect 5087 377 5120 423
rect 5166 377 5199 423
rect 11 235 123 283
rect 11 189 44 235
rect 90 189 123 235
rect 11 141 123 189
rect 11 95 44 141
rect 90 95 123 141
rect 2138 300 2214 312
rect 2138 248 2150 300
rect 2202 248 2214 300
rect 2138 196 2214 248
rect 2138 144 2150 196
rect 2202 144 2214 196
rect 2138 132 2214 144
rect 2925 283 2958 329
rect 3004 283 3037 329
rect 5087 329 5199 377
rect 2925 235 3037 283
rect 2925 189 2958 235
rect 3004 189 3037 235
rect 2925 141 3037 189
rect 11 47 123 95
rect 11 1 44 47
rect 90 1 123 47
rect 2925 95 2958 141
rect 3004 95 3037 141
rect 3544 300 3620 312
rect 3544 248 3556 300
rect 3608 248 3620 300
rect 3544 196 3620 248
rect 3544 144 3556 196
rect 3608 144 3620 196
rect 3544 132 3620 144
rect 3704 300 3780 312
rect 3704 248 3716 300
rect 3768 248 3780 300
rect 3704 196 3780 248
rect 3704 144 3716 196
rect 3768 144 3780 196
rect 3704 132 3780 144
rect 4345 300 4421 312
rect 4345 248 4357 300
rect 4409 248 4421 300
rect 4345 196 4421 248
rect 4345 144 4357 196
rect 4409 144 4421 196
rect 4345 132 4421 144
rect 5087 283 5120 329
rect 5166 283 5199 329
rect 5087 235 5199 283
rect 5087 189 5120 235
rect 5166 189 5199 235
rect 5087 141 5199 189
rect 2925 47 3037 95
rect 11 -47 123 1
rect 11 -93 44 -47
rect 90 -93 123 -47
rect 11 -141 123 -93
rect 425 -136 471 26
rect 641 -136 687 26
rect 857 -136 903 26
rect 1073 -136 1119 26
rect 1289 -136 1335 26
rect 1505 -136 1551 26
rect 1721 -136 1767 26
rect 1937 -136 1983 26
rect 2153 -136 2199 26
rect 2369 -136 2415 26
rect 2585 -136 2631 26
rect 2925 1 2958 47
rect 3004 1 3037 47
rect 2925 -47 3037 1
rect 2925 -93 2958 -47
rect 3004 -93 3037 -47
rect 11 -187 44 -141
rect 90 -187 123 -141
rect 11 -235 123 -187
rect 11 -281 44 -235
rect 90 -281 123 -235
rect 11 -329 123 -281
rect 11 -375 44 -329
rect 90 -375 123 -329
rect 11 -423 123 -375
rect 11 -469 44 -423
rect 90 -469 123 -423
rect 11 -517 123 -469
rect 11 -563 44 -517
rect 90 -563 123 -517
rect 11 -611 123 -563
rect 11 -657 44 -611
rect 90 -657 123 -611
rect 11 -705 123 -657
rect 11 -751 44 -705
rect 90 -751 123 -705
rect 2925 -141 3037 -93
rect 2925 -187 2958 -141
rect 3004 -187 3037 -141
rect 5087 95 5120 141
rect 5166 95 5199 141
rect 5087 47 5199 95
rect 5087 1 5120 47
rect 5166 1 5199 47
rect 5087 -47 5199 1
rect 5087 -93 5120 -47
rect 5166 -93 5199 -47
rect 5087 -141 5199 -93
rect 2925 -235 3037 -187
rect 2925 -281 2958 -235
rect 3004 -281 3037 -235
rect 2925 -329 3037 -281
rect 2925 -375 2958 -329
rect 3004 -375 3037 -329
rect 3384 -196 3460 -184
rect 3384 -248 3396 -196
rect 3448 -248 3460 -196
rect 3384 -300 3460 -248
rect 3384 -352 3396 -300
rect 3448 -352 3460 -300
rect 3384 -364 3460 -352
rect 4024 -196 4100 -184
rect 4024 -248 4036 -196
rect 4088 -248 4100 -196
rect 4024 -300 4100 -248
rect 4024 -352 4036 -300
rect 4088 -352 4100 -300
rect 4024 -364 4100 -352
rect 4664 -196 4740 -184
rect 4664 -248 4676 -196
rect 4728 -248 4740 -196
rect 4664 -300 4740 -248
rect 4664 -352 4676 -300
rect 4728 -352 4740 -300
rect 4664 -364 4740 -352
rect 5087 -187 5120 -141
rect 5166 -187 5199 -141
rect 5087 -235 5199 -187
rect 5087 -281 5120 -235
rect 5166 -281 5199 -235
rect 5087 -329 5199 -281
rect 2925 -423 3037 -375
rect 5087 -375 5120 -329
rect 5166 -375 5199 -329
rect 2925 -469 2958 -423
rect 3004 -469 3037 -423
rect 2925 -517 3037 -469
rect 2925 -563 2958 -517
rect 3004 -563 3037 -517
rect 2925 -611 3037 -563
rect 2925 -657 2958 -611
rect 3004 -657 3037 -611
rect 2925 -705 3037 -657
rect 11 -799 123 -751
rect 11 -845 44 -799
rect 90 -845 123 -799
rect 11 -893 123 -845
rect 11 -939 44 -893
rect 90 -939 123 -893
rect 425 -794 471 -736
rect 522 -794 590 -783
rect 641 -794 687 -736
rect 425 -840 533 -794
rect 579 -840 687 -794
rect 425 -898 471 -840
rect 522 -851 590 -840
rect 641 -898 687 -840
rect 857 -898 903 -736
rect 1073 -898 1119 -736
rect 1289 -898 1335 -736
rect 1505 -898 1551 -736
rect 1721 -898 1767 -736
rect 1937 -898 1983 -736
rect 2153 -898 2199 -736
rect 2369 -794 2415 -736
rect 2466 -794 2534 -783
rect 2585 -794 2631 -736
rect 2369 -840 2477 -794
rect 2523 -840 2631 -794
rect 2369 -898 2415 -840
rect 2466 -851 2534 -840
rect 2585 -898 2631 -840
rect 2925 -751 2958 -705
rect 3004 -751 3037 -705
rect 2925 -799 3037 -751
rect 3111 -568 3157 -388
rect 3271 -568 3317 -388
rect 3111 -614 3191 -568
rect 3237 -614 3317 -568
rect 3111 -794 3157 -614
rect 3271 -794 3317 -614
rect 3464 -477 3540 -465
rect 3464 -529 3476 -477
rect 3528 -529 3540 -477
rect 3464 -581 3540 -529
rect 3464 -633 3476 -581
rect 3528 -584 3540 -581
rect 4807 -568 4853 -388
rect 4967 -568 5013 -388
rect 3528 -630 3639 -584
rect 3685 -630 3959 -584
rect 4005 -630 4279 -584
rect 4325 -630 4599 -584
rect 4645 -630 4656 -584
rect 4807 -614 4887 -568
rect 4933 -614 5013 -568
rect 3528 -633 3540 -630
rect 3464 -645 3540 -633
rect 3559 -737 4565 -691
rect 3559 -794 3605 -737
rect 3719 -794 3765 -783
rect 3879 -794 3925 -737
rect 4039 -794 4085 -783
rect 4199 -794 4245 -737
rect 4359 -794 4405 -783
rect 4519 -794 4565 -737
rect 4807 -794 4853 -614
rect 4967 -794 5013 -614
rect 5087 -423 5199 -375
rect 5087 -469 5120 -423
rect 5166 -469 5199 -423
rect 5087 -517 5199 -469
rect 5087 -563 5120 -517
rect 5166 -563 5199 -517
rect 5087 -611 5199 -563
rect 5087 -657 5120 -611
rect 5166 -657 5199 -611
rect 5087 -705 5199 -657
rect 5087 -751 5120 -705
rect 5166 -751 5199 -705
rect 2925 -845 2958 -799
rect 3004 -845 3037 -799
rect 5087 -799 5199 -751
rect 2925 -893 3037 -845
rect 11 -987 123 -939
rect 11 -1033 44 -987
rect 90 -1033 123 -987
rect 2925 -939 2958 -893
rect 3004 -939 3037 -893
rect 2925 -987 3037 -939
rect 11 -1081 123 -1033
rect 11 -1127 44 -1081
rect 90 -1127 123 -1081
rect 11 -1175 123 -1127
rect 11 -1221 44 -1175
rect 90 -1221 123 -1175
rect 2138 -1030 2214 -1018
rect 2138 -1082 2150 -1030
rect 2202 -1082 2214 -1030
rect 2138 -1134 2214 -1082
rect 2138 -1186 2150 -1134
rect 2202 -1186 2214 -1134
rect 2138 -1198 2214 -1186
rect 2925 -1033 2958 -987
rect 3004 -1033 3037 -987
rect 3704 -830 3780 -818
rect 3704 -882 3716 -830
rect 3768 -882 3780 -830
rect 3704 -934 3780 -882
rect 3704 -986 3716 -934
rect 3768 -986 3780 -934
rect 3704 -998 3780 -986
rect 4345 -830 4421 -818
rect 4345 -882 4357 -830
rect 4409 -882 4421 -830
rect 4345 -934 4421 -882
rect 4345 -986 4357 -934
rect 4409 -986 4421 -934
rect 4345 -998 4421 -986
rect 5087 -845 5120 -799
rect 5166 -845 5199 -799
rect 5087 -893 5199 -845
rect 5087 -939 5120 -893
rect 5166 -939 5199 -893
rect 5087 -987 5199 -939
rect 2925 -1081 3037 -1033
rect 2925 -1127 2958 -1081
rect 3004 -1127 3037 -1081
rect 2925 -1175 3037 -1127
rect 11 -1269 123 -1221
rect 11 -1315 44 -1269
rect 90 -1315 123 -1269
rect 11 -1363 123 -1315
rect 11 -1409 44 -1363
rect 90 -1409 123 -1363
rect 11 -1457 123 -1409
rect 11 -1503 44 -1457
rect 90 -1503 123 -1457
rect 2925 -1221 2958 -1175
rect 3004 -1221 3037 -1175
rect 3544 -1030 3620 -1018
rect 3544 -1082 3556 -1030
rect 3608 -1082 3620 -1030
rect 3544 -1134 3620 -1082
rect 3544 -1186 3556 -1134
rect 3608 -1186 3620 -1134
rect 3544 -1198 3620 -1186
rect 5087 -1033 5120 -987
rect 5166 -1033 5199 -987
rect 5087 -1081 5199 -1033
rect 5087 -1127 5120 -1081
rect 5166 -1127 5199 -1081
rect 5087 -1175 5199 -1127
rect 2925 -1269 3037 -1221
rect 2925 -1315 2958 -1269
rect 3004 -1315 3037 -1269
rect 5087 -1221 5120 -1175
rect 5166 -1221 5199 -1175
rect 5087 -1269 5199 -1221
rect 2925 -1363 3037 -1315
rect 2925 -1409 2958 -1363
rect 3004 -1409 3037 -1363
rect 2925 -1457 3037 -1409
rect 11 -1551 123 -1503
rect -260 -1572 -80 -1562
rect -486 -1574 -80 -1572
rect -486 -1626 -248 -1574
rect -196 -1626 -144 -1574
rect -92 -1626 -80 -1574
rect -486 -1678 -80 -1626
rect -486 -1730 -248 -1678
rect -196 -1730 -144 -1678
rect -92 -1730 -80 -1678
rect -486 -1732 -80 -1730
rect -260 -1742 -80 -1732
rect 11 -1597 44 -1551
rect 90 -1597 123 -1551
rect 11 -1645 123 -1597
rect 11 -1691 44 -1645
rect 90 -1691 123 -1645
rect 11 -1739 123 -1691
rect 11 -1785 44 -1739
rect 90 -1776 123 -1739
rect 425 -1776 471 -1498
rect 641 -1776 687 -1498
rect 741 -1574 921 -1562
rect 741 -1626 753 -1574
rect 805 -1626 857 -1574
rect 909 -1626 921 -1574
rect 741 -1638 921 -1626
rect 1073 -1776 1119 -1498
rect 1505 -1776 1551 -1498
rect 1937 -1776 1983 -1498
rect 2369 -1776 2415 -1498
rect 2585 -1776 2631 -1498
rect 2925 -1503 2958 -1457
rect 3004 -1503 3037 -1457
rect 3384 -1326 3460 -1314
rect 3384 -1378 3396 -1326
rect 3448 -1378 3460 -1326
rect 3384 -1430 3460 -1378
rect 3384 -1482 3396 -1430
rect 3448 -1482 3460 -1430
rect 3384 -1494 3460 -1482
rect 4024 -1326 4100 -1314
rect 4024 -1378 4036 -1326
rect 4088 -1378 4100 -1326
rect 4024 -1430 4100 -1378
rect 4024 -1482 4036 -1430
rect 4088 -1482 4100 -1430
rect 4024 -1494 4100 -1482
rect 4664 -1326 4740 -1314
rect 4664 -1378 4676 -1326
rect 4728 -1378 4740 -1326
rect 4664 -1430 4740 -1378
rect 4664 -1482 4676 -1430
rect 4728 -1482 4740 -1430
rect 4664 -1494 4740 -1482
rect 5087 -1315 5120 -1269
rect 5166 -1315 5199 -1269
rect 5087 -1363 5199 -1315
rect 5087 -1409 5120 -1363
rect 5166 -1409 5199 -1363
rect 5087 -1457 5199 -1409
rect 2925 -1551 3037 -1503
rect 5087 -1503 5120 -1457
rect 5166 -1503 5199 -1457
rect 2925 -1597 2958 -1551
rect 3004 -1597 3037 -1551
rect 2925 -1645 3037 -1597
rect 2925 -1691 2958 -1645
rect 3004 -1691 3037 -1645
rect 2925 -1739 3037 -1691
rect 2925 -1776 2958 -1739
rect 90 -1785 2958 -1776
rect 3004 -1776 3037 -1739
rect 3111 -1776 3157 -1518
rect 3271 -1776 3317 -1518
rect 3624 -1665 3700 -1653
rect 3624 -1717 3636 -1665
rect 3688 -1668 3700 -1665
rect 3688 -1714 4279 -1668
rect 4325 -1714 4336 -1668
rect 3688 -1717 3700 -1714
rect 3624 -1729 3700 -1717
rect 4807 -1776 4853 -1518
rect 4967 -1776 5013 -1518
rect 5087 -1551 5199 -1503
rect 5087 -1597 5120 -1551
rect 5166 -1597 5199 -1551
rect 5087 -1645 5199 -1597
rect 5087 -1691 5120 -1645
rect 5166 -1691 5199 -1645
rect 5087 -1739 5199 -1691
rect 5087 -1776 5120 -1739
rect 3004 -1785 5120 -1776
rect 5166 -1785 5199 -1739
rect 11 -1833 5199 -1785
rect 11 -1879 44 -1833
rect 90 -1879 138 -1833
rect 184 -1879 232 -1833
rect 278 -1879 326 -1833
rect 372 -1879 420 -1833
rect 466 -1879 514 -1833
rect 560 -1879 608 -1833
rect 654 -1879 702 -1833
rect 748 -1879 796 -1833
rect 842 -1879 890 -1833
rect 936 -1879 984 -1833
rect 1030 -1879 1078 -1833
rect 1124 -1879 1172 -1833
rect 1218 -1879 1266 -1833
rect 1312 -1879 1360 -1833
rect 1406 -1879 1454 -1833
rect 1500 -1879 1548 -1833
rect 1594 -1879 1642 -1833
rect 1688 -1879 1736 -1833
rect 1782 -1879 1830 -1833
rect 1876 -1879 1924 -1833
rect 1970 -1879 2018 -1833
rect 2064 -1879 2112 -1833
rect 2158 -1879 2206 -1833
rect 2252 -1879 2300 -1833
rect 2346 -1879 2394 -1833
rect 2440 -1879 2488 -1833
rect 2534 -1879 2582 -1833
rect 2628 -1879 2676 -1833
rect 2722 -1879 2770 -1833
rect 2816 -1879 2864 -1833
rect 2910 -1879 2958 -1833
rect 3004 -1879 3052 -1833
rect 3098 -1879 3146 -1833
rect 3192 -1879 3240 -1833
rect 3286 -1879 3334 -1833
rect 3380 -1879 3428 -1833
rect 3474 -1879 3522 -1833
rect 3568 -1879 3616 -1833
rect 3662 -1879 3710 -1833
rect 3756 -1879 3804 -1833
rect 3850 -1879 3898 -1833
rect 3944 -1879 3992 -1833
rect 4038 -1879 4086 -1833
rect 4132 -1879 4180 -1833
rect 4226 -1879 4274 -1833
rect 4320 -1879 4368 -1833
rect 4414 -1879 4462 -1833
rect 4508 -1879 4556 -1833
rect 4602 -1879 4650 -1833
rect 4696 -1879 4744 -1833
rect 4790 -1879 4838 -1833
rect 4884 -1879 4932 -1833
rect 4978 -1879 5026 -1833
rect 5072 -1879 5120 -1833
rect 5166 -1879 5199 -1833
rect 11 -1936 5199 -1879
rect 5743 4616 5776 4662
rect 5822 4616 5855 4662
rect 6569 4820 6645 4832
rect 6569 4768 6581 4820
rect 6633 4768 6645 4820
rect 6569 4716 6645 4768
rect 6569 4664 6581 4716
rect 6633 4664 6645 4716
rect 6569 4652 6645 4664
rect 7209 4820 7285 4832
rect 7209 4768 7221 4820
rect 7273 4768 7285 4820
rect 7209 4716 7285 4768
rect 7209 4664 7221 4716
rect 7273 4664 7285 4716
rect 7209 4652 7285 4664
rect 7999 4804 8032 4850
rect 8078 4804 8159 4850
rect 7999 4756 8159 4804
rect 7999 4710 8032 4756
rect 8078 4720 8159 4756
rect 8667 4720 8827 5245
rect 9372 4720 9532 5245
rect 10186 4720 10346 5245
rect 21527 4720 21847 5245
rect 26164 4720 26484 5245
rect 29586 4720 29906 5245
rect 8078 4710 29906 4720
rect 7999 4662 29906 4710
rect 5743 4568 5855 4616
rect 5743 4522 5776 4568
rect 5822 4522 5855 4568
rect 7999 4616 8032 4662
rect 8078 4616 29906 4662
rect 7999 4611 29906 4616
rect 7999 4568 17650 4611
rect 5743 4474 5855 4522
rect 5743 4428 5776 4474
rect 5822 4428 5855 4474
rect 5743 4380 5855 4428
rect 5743 4334 5776 4380
rect 5822 4334 5855 4380
rect 5743 4286 5855 4334
rect 5743 4240 5776 4286
rect 5822 4240 5855 4286
rect 5976 4244 6022 4556
rect 6136 4244 6182 4556
rect 6424 4244 6470 4556
rect 6744 4244 6790 4556
rect 7064 4244 7110 4556
rect 7384 4244 7430 4556
rect 7672 4244 7718 4556
rect 7832 4244 7878 4556
rect 7999 4522 8032 4568
rect 8078 4565 17650 4568
rect 17696 4565 17744 4611
rect 17790 4565 17838 4611
rect 17884 4565 17932 4611
rect 17978 4565 18026 4611
rect 18072 4565 18120 4611
rect 18166 4565 18214 4611
rect 18260 4565 18308 4611
rect 18354 4565 18402 4611
rect 18448 4565 18496 4611
rect 18542 4565 18590 4611
rect 18636 4565 18684 4611
rect 18730 4565 18778 4611
rect 18824 4565 18872 4611
rect 18918 4565 18966 4611
rect 19012 4565 19060 4611
rect 19106 4565 19154 4611
rect 19200 4565 19248 4611
rect 19294 4565 19342 4611
rect 19388 4565 19436 4611
rect 19482 4565 19530 4611
rect 19576 4565 19624 4611
rect 19670 4565 19718 4611
rect 19764 4565 19812 4611
rect 19858 4565 19906 4611
rect 19952 4565 20000 4611
rect 20046 4565 20094 4611
rect 20140 4565 20188 4611
rect 20234 4565 20282 4611
rect 20328 4565 20376 4611
rect 20422 4565 20470 4611
rect 20516 4565 20564 4611
rect 20610 4565 20658 4611
rect 20704 4565 22802 4611
rect 22848 4565 22896 4611
rect 22942 4565 22990 4611
rect 23036 4565 23084 4611
rect 23130 4565 23178 4611
rect 23224 4565 23272 4611
rect 23318 4565 23366 4611
rect 23412 4565 23460 4611
rect 23506 4565 23554 4611
rect 23600 4565 23648 4611
rect 23694 4565 23742 4611
rect 23788 4565 23836 4611
rect 23882 4565 23930 4611
rect 23976 4565 24024 4611
rect 24070 4565 24118 4611
rect 24164 4565 24212 4611
rect 24258 4565 24306 4611
rect 24352 4565 24400 4611
rect 24446 4565 24494 4611
rect 24540 4565 24588 4611
rect 24634 4565 24682 4611
rect 24728 4565 24776 4611
rect 24822 4565 24870 4611
rect 24916 4565 24964 4611
rect 25010 4565 25058 4611
rect 25104 4565 25152 4611
rect 25198 4565 25246 4611
rect 25292 4565 25340 4611
rect 25386 4565 25434 4611
rect 25480 4565 25528 4611
rect 25574 4565 25622 4611
rect 25668 4565 25716 4611
rect 25762 4565 25810 4611
rect 25856 4565 26771 4611
rect 26817 4565 26865 4611
rect 26911 4565 26959 4611
rect 27005 4565 27053 4611
rect 27099 4565 27147 4611
rect 27193 4565 27241 4611
rect 27287 4565 27335 4611
rect 27381 4565 27429 4611
rect 27475 4565 27523 4611
rect 27569 4565 27617 4611
rect 27663 4565 27711 4611
rect 27757 4565 27805 4611
rect 27851 4565 27899 4611
rect 27945 4565 27993 4611
rect 28039 4565 28087 4611
rect 28133 4565 28181 4611
rect 28227 4565 28275 4611
rect 28321 4565 28369 4611
rect 28415 4565 28463 4611
rect 28509 4565 28557 4611
rect 28603 4565 28651 4611
rect 28697 4565 28745 4611
rect 28791 4565 28839 4611
rect 28885 4565 28933 4611
rect 28979 4565 29027 4611
rect 29073 4565 29121 4611
rect 29167 4565 29215 4611
rect 29261 4565 29309 4611
rect 29355 4565 29403 4611
rect 29449 4565 29497 4611
rect 29543 4565 29591 4611
rect 29637 4565 29685 4611
rect 29731 4565 29779 4611
rect 29825 4565 29906 4611
rect 8078 4522 29906 4565
rect 7999 4517 29906 4522
rect 7999 4474 17650 4517
rect 7999 4428 8032 4474
rect 8078 4471 17650 4474
rect 17696 4471 20658 4517
rect 20704 4471 22802 4517
rect 22848 4471 25810 4517
rect 25856 4471 26771 4517
rect 26817 4471 29779 4517
rect 29825 4471 29906 4517
rect 8078 4428 29906 4471
rect 7999 4423 29906 4428
rect 7999 4400 17650 4423
rect 7999 4380 8159 4400
rect 7999 4334 8032 4380
rect 8078 4334 8159 4380
rect 7999 4286 8159 4334
rect 5743 4192 5855 4240
rect 7999 4240 8032 4286
rect 8078 4240 8159 4286
rect 5743 4146 5776 4192
rect 5822 4146 5855 4192
rect 5743 4098 5855 4146
rect 5743 4052 5776 4098
rect 5822 4052 5855 4098
rect 6569 4220 6645 4232
rect 6569 4168 6581 4220
rect 6633 4168 6645 4220
rect 6569 4116 6645 4168
rect 6569 4064 6581 4116
rect 6633 4064 6645 4116
rect 6569 4052 6645 4064
rect 7209 4220 7285 4232
rect 7209 4168 7221 4220
rect 7273 4168 7285 4220
rect 7209 4116 7285 4168
rect 7209 4064 7221 4116
rect 7273 4064 7285 4116
rect 7209 4052 7285 4064
rect 7999 4192 8159 4240
rect 7999 4146 8032 4192
rect 8078 4146 8159 4192
rect 7999 4098 8159 4146
rect 7999 4052 8032 4098
rect 8078 4052 8159 4098
rect 5743 4004 5855 4052
rect 5743 3958 5776 4004
rect 5822 3958 5855 4004
rect 5743 3910 5855 3958
rect 5743 3864 5776 3910
rect 5822 3864 5855 3910
rect 5743 3816 5855 3864
rect 7999 4004 8159 4052
rect 7999 3958 8032 4004
rect 8078 3958 8159 4004
rect 7999 3920 8159 3958
rect 8667 3920 8827 4400
rect 9372 3920 9532 4400
rect 10186 3920 10346 4400
rect 17569 4377 17650 4400
rect 17696 4400 20658 4423
rect 17696 4377 17889 4400
rect 17569 4329 17889 4377
rect 17569 4283 17650 4329
rect 17696 4283 17889 4329
rect 17569 4235 17889 4283
rect 17569 4189 17650 4235
rect 17696 4189 17889 4235
rect 17569 4141 17889 4189
rect 17569 4095 17650 4141
rect 17696 4095 17889 4141
rect 17569 4047 17889 4095
rect 17569 4001 17650 4047
rect 17696 4001 17889 4047
rect 18226 4019 18272 4400
rect 18386 4019 18432 4400
rect 18579 4248 18655 4260
rect 18579 4196 18591 4248
rect 18643 4245 18655 4248
rect 19699 4248 19775 4260
rect 19699 4245 19711 4248
rect 18643 4199 19074 4245
rect 19120 4199 19711 4245
rect 18643 4196 18655 4199
rect 18579 4184 18655 4196
rect 19699 4196 19711 4199
rect 19763 4196 19775 4248
rect 19699 4184 19775 4196
rect 19922 4019 19968 4400
rect 20082 4019 20128 4400
rect 20465 4377 20658 4400
rect 20704 4400 22802 4423
rect 20704 4377 20785 4400
rect 20465 4329 20785 4377
rect 20465 4283 20658 4329
rect 20704 4283 20785 4329
rect 20465 4235 20785 4283
rect 20465 4189 20658 4235
rect 20704 4189 20785 4235
rect 20465 4141 20785 4189
rect 20465 4095 20658 4141
rect 20704 4095 20785 4141
rect 20465 4047 20785 4095
rect 17569 3953 17889 4001
rect 17569 3920 17650 3953
rect 7999 3910 17650 3920
rect 7999 3864 8032 3910
rect 8078 3907 17650 3910
rect 17696 3907 17889 3953
rect 8078 3864 17889 3907
rect 7999 3859 17889 3864
rect 5743 3770 5776 3816
rect 5822 3770 5855 3816
rect 5743 3722 5855 3770
rect 5743 3676 5776 3722
rect 5822 3676 5855 3722
rect 6249 3841 6325 3853
rect 6249 3789 6261 3841
rect 6313 3789 6325 3841
rect 6249 3737 6325 3789
rect 5743 3628 5855 3676
rect 5743 3582 5776 3628
rect 5822 3582 5855 3628
rect 5743 3534 5855 3582
rect 5743 3488 5776 3534
rect 5822 3488 5855 3534
rect 5743 3440 5855 3488
rect 5743 3394 5776 3440
rect 5822 3394 5855 3440
rect 5743 3346 5855 3394
rect 5976 3382 6022 3694
rect 6136 3382 6182 3694
rect 6249 3685 6261 3737
rect 6313 3685 6325 3737
rect 6889 3841 6965 3853
rect 6889 3789 6901 3841
rect 6953 3789 6965 3841
rect 6889 3737 6965 3789
rect 6249 3673 6325 3685
rect 6424 3382 6470 3694
rect 6744 3382 6790 3694
rect 6889 3685 6901 3737
rect 6953 3685 6965 3737
rect 7529 3841 7605 3853
rect 7529 3789 7541 3841
rect 7593 3789 7605 3841
rect 7529 3737 7605 3789
rect 6889 3673 6965 3685
rect 7064 3382 7110 3694
rect 7384 3382 7430 3694
rect 7529 3685 7541 3737
rect 7593 3685 7605 3737
rect 7999 3816 17650 3859
rect 7999 3770 8032 3816
rect 8078 3813 17650 3816
rect 17696 3813 17889 3859
rect 18819 4007 18895 4019
rect 18819 3955 18831 4007
rect 18883 3955 18895 4007
rect 18819 3903 18895 3955
rect 18819 3851 18831 3903
rect 18883 3851 18895 3903
rect 18819 3839 18895 3851
rect 19459 4007 19535 4019
rect 19459 3955 19471 4007
rect 19523 3955 19535 4007
rect 19459 3903 19535 3955
rect 19459 3851 19471 3903
rect 19523 3851 19535 3903
rect 19459 3839 19535 3851
rect 20465 4001 20658 4047
rect 20704 4001 20785 4047
rect 20465 3953 20785 4001
rect 20465 3907 20658 3953
rect 20704 3907 20785 3953
rect 20465 3859 20785 3907
rect 8078 3770 17889 3813
rect 7999 3765 17889 3770
rect 7999 3722 17650 3765
rect 7529 3673 7605 3685
rect 7672 3382 7718 3694
rect 7832 3382 7878 3694
rect 7999 3676 8032 3722
rect 8078 3719 17650 3722
rect 17696 3719 17889 3765
rect 8078 3676 17889 3719
rect 7999 3671 17889 3676
rect 7999 3628 17650 3671
rect 7999 3582 8032 3628
rect 8078 3625 17650 3628
rect 17696 3625 17889 3671
rect 20465 3813 20658 3859
rect 20704 3813 20785 3859
rect 20465 3765 20785 3813
rect 20465 3719 20658 3765
rect 20704 3719 20785 3765
rect 20465 3671 20785 3719
rect 20465 3625 20658 3671
rect 20704 3625 20785 3671
rect 8078 3600 17889 3625
rect 8078 3582 8159 3600
rect 7999 3534 8159 3582
rect 7999 3488 8032 3534
rect 8078 3488 8159 3534
rect 7999 3440 8159 3488
rect 7999 3394 8032 3440
rect 8078 3394 8159 3440
rect 5743 3291 5776 3346
rect 5822 3291 5855 3346
rect 7999 3346 8159 3394
rect 5743 3243 5855 3291
rect 5743 3197 5776 3243
rect 5822 3197 5855 3243
rect 5743 3149 5855 3197
rect 5743 3103 5776 3149
rect 5822 3103 5855 3149
rect 6569 3298 6645 3310
rect 6569 3246 6581 3298
rect 6633 3246 6645 3298
rect 6569 3194 6645 3246
rect 6569 3142 6581 3194
rect 6633 3142 6645 3194
rect 6569 3130 6645 3142
rect 7209 3298 7285 3310
rect 7209 3246 7221 3298
rect 7273 3246 7285 3298
rect 7209 3194 7285 3246
rect 7209 3142 7221 3194
rect 7273 3142 7285 3194
rect 7209 3130 7285 3142
rect 7999 3291 8032 3346
rect 8078 3291 8159 3346
rect 7999 3243 8159 3291
rect 7999 3197 8032 3243
rect 8078 3197 8159 3243
rect 7999 3149 8159 3197
rect 5743 3055 5855 3103
rect 5743 3009 5776 3055
rect 5822 3009 5855 3055
rect 5743 2961 5855 3009
rect 7999 3103 8032 3149
rect 8078 3103 8159 3149
rect 7999 3055 8159 3103
rect 7999 3009 8032 3055
rect 8078 3009 8159 3055
rect 5743 2915 5776 2961
rect 5822 2915 5855 2961
rect 5743 2867 5855 2915
rect 5743 2821 5776 2867
rect 5822 2821 5855 2867
rect 6249 2979 6325 2991
rect 6249 2927 6261 2979
rect 6313 2927 6325 2979
rect 6889 2979 6965 2991
rect 6249 2875 6325 2927
rect 5743 2773 5855 2821
rect 5743 2727 5776 2773
rect 5822 2727 5855 2773
rect 5743 2679 5855 2727
rect 5743 2633 5776 2679
rect 5822 2633 5855 2679
rect 5743 2585 5855 2633
rect 5743 2539 5776 2585
rect 5822 2539 5855 2585
rect 5743 2491 5855 2539
rect 5976 2520 6022 2832
rect 6136 2520 6182 2832
rect 6249 2823 6261 2875
rect 6313 2823 6325 2875
rect 6249 2811 6325 2823
rect 6424 2520 6470 2936
rect 6744 2520 6790 2936
rect 6889 2927 6901 2979
rect 6953 2927 6965 2979
rect 7529 2979 7605 2991
rect 6889 2875 6965 2927
rect 6889 2823 6901 2875
rect 6953 2823 6965 2875
rect 6889 2811 6965 2823
rect 7064 2520 7110 2936
rect 7384 2520 7430 2936
rect 7529 2927 7541 2979
rect 7593 2927 7605 2979
rect 7529 2875 7605 2927
rect 7529 2823 7541 2875
rect 7593 2823 7605 2875
rect 7999 2961 8159 3009
rect 7999 2915 8032 2961
rect 8078 2915 8159 2961
rect 7999 2867 8159 2915
rect 7529 2811 7605 2823
rect 7672 2520 7718 2832
rect 7832 2520 7878 2832
rect 7999 2821 8032 2867
rect 8078 2821 8159 2867
rect 7999 2773 8159 2821
rect 7999 2727 8032 2773
rect 8078 2727 8159 2773
rect 7999 2679 8159 2727
rect 7999 2633 8032 2679
rect 8078 2633 8159 2679
rect 7999 2585 8159 2633
rect 7999 2539 8032 2585
rect 8078 2539 8159 2585
rect 5743 2445 5776 2491
rect 5822 2445 5855 2491
rect 7999 2491 8159 2539
rect 5743 2397 5855 2445
rect 5743 2351 5776 2397
rect 5822 2351 5855 2397
rect 5743 2303 5855 2351
rect 5743 2257 5776 2303
rect 5822 2257 5855 2303
rect 6249 2456 6325 2468
rect 6249 2404 6261 2456
rect 6313 2404 6325 2456
rect 6249 2352 6325 2404
rect 6249 2300 6261 2352
rect 6313 2300 6325 2352
rect 6249 2288 6325 2300
rect 6889 2456 6965 2468
rect 6889 2404 6901 2456
rect 6953 2404 6965 2456
rect 6889 2352 6965 2404
rect 6889 2300 6901 2352
rect 6953 2300 6965 2352
rect 6889 2288 6965 2300
rect 7529 2456 7605 2468
rect 7529 2404 7541 2456
rect 7593 2404 7605 2456
rect 7529 2352 7605 2404
rect 7529 2300 7541 2352
rect 7593 2300 7605 2352
rect 7529 2288 7605 2300
rect 7999 2445 8032 2491
rect 8078 2445 8159 2491
rect 7999 2397 8159 2445
rect 7999 2351 8032 2397
rect 8078 2351 8159 2397
rect 7999 2303 8159 2351
rect 5743 2209 5855 2257
rect 5743 2163 5776 2209
rect 5822 2163 5855 2209
rect 7999 2257 8032 2303
rect 8078 2257 8159 2303
rect 7999 2209 8159 2257
rect 5743 2115 5855 2163
rect 5743 2069 5776 2115
rect 5822 2069 5855 2115
rect 5743 2021 5855 2069
rect 5743 1975 5776 2021
rect 5822 1975 5855 2021
rect 6569 2168 6645 2180
rect 6569 2116 6581 2168
rect 6633 2116 6645 2168
rect 6569 2064 6645 2116
rect 6569 2012 6581 2064
rect 6633 2012 6645 2064
rect 6569 2000 6645 2012
rect 7209 2168 7285 2180
rect 7209 2116 7221 2168
rect 7273 2116 7285 2168
rect 7209 2064 7285 2116
rect 7209 2012 7221 2064
rect 7273 2012 7285 2064
rect 7209 2000 7285 2012
rect 7999 2163 8032 2209
rect 8078 2163 8159 2209
rect 7999 2115 8159 2163
rect 7999 2069 8032 2115
rect 8078 2078 8159 2115
rect 8667 2078 8827 3600
rect 9372 2078 9532 3600
rect 10186 2078 10346 3600
rect 17569 3577 17889 3600
rect 17569 3531 17650 3577
rect 17696 3531 17889 3577
rect 17569 3483 17889 3531
rect 17569 3437 17650 3483
rect 17696 3437 17889 3483
rect 18499 3613 18575 3625
rect 18499 3561 18511 3613
rect 18563 3561 18575 3613
rect 18499 3509 18575 3561
rect 18499 3457 18511 3509
rect 18563 3457 18575 3509
rect 18499 3445 18575 3457
rect 18659 3613 18735 3625
rect 18659 3561 18671 3613
rect 18723 3561 18735 3613
rect 18659 3509 18735 3561
rect 18659 3457 18671 3509
rect 18723 3457 18735 3509
rect 18659 3445 18735 3457
rect 18979 3613 19055 3625
rect 18979 3561 18991 3613
rect 19043 3561 19055 3613
rect 18979 3509 19055 3561
rect 18979 3457 18991 3509
rect 19043 3457 19055 3509
rect 18979 3445 19055 3457
rect 19139 3613 19215 3625
rect 19139 3561 19151 3613
rect 19203 3561 19215 3613
rect 19139 3509 19215 3561
rect 19139 3457 19151 3509
rect 19203 3457 19215 3509
rect 19139 3445 19215 3457
rect 19299 3613 19375 3625
rect 19299 3561 19311 3613
rect 19363 3561 19375 3613
rect 19299 3509 19375 3561
rect 19299 3457 19311 3509
rect 19363 3457 19375 3509
rect 19299 3445 19375 3457
rect 19619 3613 19695 3625
rect 19619 3561 19631 3613
rect 19683 3561 19695 3613
rect 19619 3509 19695 3561
rect 19619 3457 19631 3509
rect 19683 3457 19695 3509
rect 19619 3445 19695 3457
rect 19779 3613 19855 3625
rect 19779 3561 19791 3613
rect 19843 3561 19855 3613
rect 19779 3509 19855 3561
rect 19779 3457 19791 3509
rect 19843 3457 19855 3509
rect 19779 3445 19855 3457
rect 20465 3577 20785 3625
rect 20465 3531 20658 3577
rect 20704 3531 20785 3577
rect 20465 3483 20785 3531
rect 17569 3389 17889 3437
rect 17569 3343 17650 3389
rect 17696 3343 17889 3389
rect 17569 3295 17889 3343
rect 17569 3249 17650 3295
rect 17696 3249 17889 3295
rect 17569 3201 17889 3249
rect 17569 3155 17650 3201
rect 17696 3155 17889 3201
rect 17569 3107 17889 3155
rect 17569 3061 17650 3107
rect 17696 3061 17889 3107
rect 17569 3013 17889 3061
rect 17569 2967 17650 3013
rect 17696 2967 17889 3013
rect 17569 2919 17889 2967
rect 17569 2873 17650 2919
rect 17696 2873 17889 2919
rect 17569 2825 17889 2873
rect 17569 2779 17650 2825
rect 17696 2779 17889 2825
rect 17569 2731 17889 2779
rect 17569 2685 17650 2731
rect 17696 2685 17889 2731
rect 11381 2585 16569 2642
rect 11381 2539 11414 2585
rect 11460 2539 11508 2585
rect 11554 2539 11602 2585
rect 11648 2539 11696 2585
rect 11742 2539 11790 2585
rect 11836 2539 11884 2585
rect 11930 2539 11978 2585
rect 12024 2539 12072 2585
rect 12118 2539 12166 2585
rect 12212 2539 12260 2585
rect 12306 2539 12354 2585
rect 12400 2539 12448 2585
rect 12494 2539 12542 2585
rect 12588 2539 12636 2585
rect 12682 2539 12730 2585
rect 12776 2539 12824 2585
rect 12870 2539 12918 2585
rect 12964 2539 13012 2585
rect 13058 2539 13106 2585
rect 13152 2539 13200 2585
rect 13246 2539 13294 2585
rect 13340 2539 13388 2585
rect 13434 2539 13482 2585
rect 13528 2539 13576 2585
rect 13622 2539 13670 2585
rect 13716 2539 13764 2585
rect 13810 2539 13858 2585
rect 13904 2539 13952 2585
rect 13998 2539 14046 2585
rect 14092 2539 14140 2585
rect 14186 2539 14234 2585
rect 14280 2539 14328 2585
rect 14374 2539 14422 2585
rect 14468 2539 14516 2585
rect 14562 2539 14610 2585
rect 14656 2539 14704 2585
rect 14750 2539 14798 2585
rect 14844 2539 14892 2585
rect 14938 2539 14986 2585
rect 15032 2539 15080 2585
rect 15126 2539 15174 2585
rect 15220 2539 15268 2585
rect 15314 2539 15362 2585
rect 15408 2539 15456 2585
rect 15502 2539 15550 2585
rect 15596 2539 15644 2585
rect 15690 2539 15738 2585
rect 15784 2539 15832 2585
rect 15878 2539 15926 2585
rect 15972 2539 16020 2585
rect 16066 2539 16114 2585
rect 16160 2539 16208 2585
rect 16254 2539 16302 2585
rect 16348 2539 16396 2585
rect 16442 2539 16490 2585
rect 16536 2539 16569 2585
rect 10895 2228 11055 2518
rect 10885 2216 11065 2228
rect 10885 2164 10897 2216
rect 10949 2164 11001 2216
rect 11053 2164 11065 2216
rect 10885 2112 11065 2164
rect 8078 2069 10837 2078
rect 7999 2021 10837 2069
rect 10885 2060 10897 2112
rect 10949 2060 11001 2112
rect 11053 2060 11065 2112
rect 10885 2048 11065 2060
rect 5743 1927 5855 1975
rect 7999 1975 8032 2021
rect 8078 1975 8126 2021
rect 8172 1975 8220 2021
rect 8266 1975 8314 2021
rect 8360 1975 8408 2021
rect 8454 1975 8502 2021
rect 8548 1975 8596 2021
rect 8642 1975 8690 2021
rect 8736 1975 8784 2021
rect 8830 1975 8878 2021
rect 8924 1975 8972 2021
rect 9018 1975 9066 2021
rect 9112 1975 9160 2021
rect 9206 1975 9254 2021
rect 9300 1975 9348 2021
rect 9394 1975 9442 2021
rect 9488 1975 9536 2021
rect 9582 1975 9630 2021
rect 9676 1975 9724 2021
rect 9770 1975 9818 2021
rect 9864 1975 9912 2021
rect 9958 1975 10006 2021
rect 10052 1975 10100 2021
rect 10146 1975 10194 2021
rect 10240 1975 10288 2021
rect 10334 1975 10382 2021
rect 10428 1975 10476 2021
rect 10522 1975 10570 2021
rect 10616 1975 10664 2021
rect 10710 1975 10758 2021
rect 10804 1975 10837 2021
rect 5743 1881 5776 1927
rect 5822 1881 5855 1927
rect 5743 1833 5855 1881
rect 5743 1787 5776 1833
rect 5822 1787 5855 1833
rect 5743 1739 5855 1787
rect 5743 1693 5776 1739
rect 5822 1693 5855 1739
rect 5743 1645 5855 1693
rect 5976 1658 6022 1970
rect 6136 1658 6182 1970
rect 6264 1658 6310 1970
rect 6424 1658 6470 1970
rect 6584 1658 6630 1970
rect 6744 1658 6790 1970
rect 6904 1658 6950 1970
rect 7064 1658 7110 1970
rect 7224 1658 7270 1970
rect 7384 1658 7430 1970
rect 7544 1658 7590 1970
rect 7672 1658 7718 1970
rect 7832 1658 7878 1970
rect 7999 1927 10837 1975
rect 7999 1881 8032 1927
rect 8078 1918 10758 1927
rect 8078 1881 8111 1918
rect 7999 1833 8111 1881
rect 7999 1787 8032 1833
rect 8078 1787 8111 1833
rect 7999 1739 8111 1787
rect 7999 1693 8032 1739
rect 8078 1693 8111 1739
rect 5743 1599 5776 1645
rect 5822 1599 5855 1645
rect 5743 1551 5855 1599
rect 5743 1505 5776 1551
rect 5822 1505 5855 1551
rect 5743 1457 5855 1505
rect 5743 1411 5776 1457
rect 5822 1411 5855 1457
rect 5743 1363 5855 1411
rect 5743 1317 5776 1363
rect 5822 1317 5855 1363
rect 5743 1269 5855 1317
rect 5743 1223 5776 1269
rect 5822 1223 5855 1269
rect 5743 1175 5855 1223
rect 5743 1129 5776 1175
rect 5822 1129 5855 1175
rect 5743 1081 5855 1129
rect 7999 1645 8111 1693
rect 7999 1599 8032 1645
rect 8078 1599 8111 1645
rect 8211 1639 8257 1918
rect 8371 1639 8417 1918
rect 8659 1696 10177 1742
rect 7999 1551 8111 1599
rect 7999 1505 8032 1551
rect 8078 1505 8111 1551
rect 7999 1457 8111 1505
rect 8484 1637 8560 1649
rect 8659 1639 8705 1696
rect 9235 1639 9281 1696
rect 8484 1585 8496 1637
rect 8548 1585 8560 1637
rect 8484 1533 8560 1585
rect 8484 1481 8496 1533
rect 8548 1481 8560 1533
rect 8484 1469 8560 1481
rect 9380 1637 9456 1649
rect 9555 1639 9601 1696
rect 10131 1639 10177 1696
rect 9380 1585 9392 1637
rect 9444 1585 9456 1637
rect 9380 1533 9456 1585
rect 9380 1481 9392 1533
rect 9444 1481 9456 1533
rect 9380 1469 9456 1481
rect 10276 1637 10352 1649
rect 10419 1639 10465 1918
rect 10579 1639 10625 1918
rect 10725 1881 10758 1918
rect 10804 1881 10837 1927
rect 10725 1833 10837 1881
rect 10725 1787 10758 1833
rect 10804 1787 10837 1833
rect 11163 1808 11323 2518
rect 11381 2491 16569 2539
rect 17569 2637 17889 2685
rect 17569 2591 17650 2637
rect 17696 2591 17889 2637
rect 17569 2543 17889 2591
rect 11381 2445 11414 2491
rect 11460 2482 14140 2491
rect 11460 2445 11493 2482
rect 11381 2397 11493 2445
rect 11381 2351 11414 2397
rect 11460 2351 11493 2397
rect 11381 2303 11493 2351
rect 11381 2257 11414 2303
rect 11460 2257 11493 2303
rect 11381 2209 11493 2257
rect 11381 2163 11414 2209
rect 11460 2163 11493 2209
rect 11593 2207 11639 2482
rect 11753 2207 11799 2482
rect 12041 2287 13559 2333
rect 12041 2207 12087 2287
rect 12314 2216 12390 2228
rect 11381 2115 11493 2163
rect 11381 2069 11414 2115
rect 11460 2069 11493 2115
rect 11381 2021 11493 2069
rect 12314 2164 12326 2216
rect 12378 2164 12390 2216
rect 12617 2207 12663 2287
rect 12937 2207 12983 2287
rect 13513 2228 13559 2287
rect 13210 2216 13286 2228
rect 12314 2112 12390 2164
rect 12314 2060 12326 2112
rect 12378 2060 12390 2112
rect 12314 2048 12390 2060
rect 13210 2164 13222 2216
rect 13274 2164 13286 2216
rect 13210 2112 13286 2164
rect 13210 2060 13222 2112
rect 13274 2060 13286 2112
rect 13210 2048 13286 2060
rect 13498 2216 13574 2228
rect 13498 2164 13510 2216
rect 13562 2164 13574 2216
rect 13801 2207 13847 2482
rect 13961 2207 14007 2482
rect 14107 2445 14140 2482
rect 14186 2482 16490 2491
rect 14186 2445 14219 2482
rect 14107 2397 14219 2445
rect 14107 2351 14140 2397
rect 14186 2351 14219 2397
rect 14107 2303 14219 2351
rect 14107 2257 14140 2303
rect 14186 2257 14219 2303
rect 14107 2209 14219 2257
rect 13498 2112 13574 2164
rect 13498 2060 13510 2112
rect 13562 2060 13574 2112
rect 13498 2048 13574 2060
rect 14107 2163 14140 2209
rect 14186 2163 14219 2209
rect 14387 2207 14433 2482
rect 14547 2207 14593 2482
rect 14660 2216 14736 2228
rect 14107 2115 14219 2163
rect 14107 2069 14140 2115
rect 14186 2069 14219 2115
rect 11381 1975 11414 2021
rect 11460 1975 11493 2021
rect 11381 1927 11493 1975
rect 11381 1881 11414 1927
rect 11460 1881 11493 1927
rect 11381 1833 11493 1881
rect 10725 1739 10837 1787
rect 10725 1693 10758 1739
rect 10804 1693 10837 1739
rect 10725 1645 10837 1693
rect 10276 1585 10288 1637
rect 10340 1585 10352 1637
rect 10276 1533 10352 1585
rect 10276 1481 10288 1533
rect 10340 1481 10352 1533
rect 10276 1469 10352 1481
rect 10725 1599 10758 1645
rect 10804 1599 10837 1645
rect 11153 1796 11333 1808
rect 11153 1744 11165 1796
rect 11217 1744 11269 1796
rect 11321 1744 11333 1796
rect 11153 1692 11333 1744
rect 11153 1640 11165 1692
rect 11217 1640 11269 1692
rect 11321 1640 11333 1692
rect 11153 1628 11333 1640
rect 11381 1787 11414 1833
rect 11460 1787 11493 1833
rect 14107 2021 14219 2069
rect 14660 2164 14672 2216
rect 14724 2164 14736 2216
rect 14835 2207 14881 2482
rect 15155 2207 15201 2482
rect 15300 2216 15376 2228
rect 14660 2112 14736 2164
rect 14660 2060 14672 2112
rect 14724 2060 14736 2112
rect 14660 2048 14736 2060
rect 15300 2164 15312 2216
rect 15364 2164 15376 2216
rect 15475 2207 15521 2482
rect 15795 2207 15841 2482
rect 15940 2216 16016 2228
rect 15300 2112 15376 2164
rect 15300 2060 15312 2112
rect 15364 2060 15376 2112
rect 15300 2048 15376 2060
rect 15940 2164 15952 2216
rect 16004 2164 16016 2216
rect 16083 2207 16129 2482
rect 16243 2207 16289 2482
rect 16457 2445 16490 2482
rect 16536 2445 16569 2491
rect 16457 2397 16569 2445
rect 16457 2351 16490 2397
rect 16536 2351 16569 2397
rect 16457 2303 16569 2351
rect 16457 2257 16490 2303
rect 16536 2257 16569 2303
rect 16457 2209 16569 2257
rect 15940 2112 16016 2164
rect 15940 2060 15952 2112
rect 16004 2060 16016 2112
rect 15940 2048 16016 2060
rect 16457 2163 16490 2209
rect 16536 2163 16569 2209
rect 16457 2115 16569 2163
rect 16457 2069 16490 2115
rect 16536 2069 16569 2115
rect 14107 1975 14140 2021
rect 14186 1975 14219 2021
rect 14107 1927 14219 1975
rect 14107 1881 14140 1927
rect 14186 1881 14219 1927
rect 14107 1833 14219 1881
rect 11381 1739 11493 1787
rect 11381 1693 11414 1739
rect 11460 1693 11493 1739
rect 11381 1645 11493 1693
rect 10725 1551 10837 1599
rect 10725 1505 10758 1551
rect 10804 1505 10837 1551
rect 7999 1411 8032 1457
rect 8078 1411 8111 1457
rect 7999 1363 8111 1411
rect 7999 1317 8032 1363
rect 8078 1317 8111 1363
rect 7999 1269 8111 1317
rect 10725 1457 10837 1505
rect 10725 1411 10758 1457
rect 10804 1411 10837 1457
rect 10725 1363 10837 1411
rect 10725 1317 10758 1363
rect 10804 1317 10837 1363
rect 7999 1223 8032 1269
rect 8078 1223 8111 1269
rect 7999 1175 8111 1223
rect 7999 1129 8032 1175
rect 8078 1129 8111 1175
rect 5743 1035 5776 1081
rect 5822 1035 5855 1081
rect 5743 987 5855 1035
rect 5743 941 5776 987
rect 5822 941 5855 987
rect 5743 893 5855 941
rect 5743 847 5776 893
rect 5822 847 5855 893
rect 5743 799 5855 847
rect 5743 753 5776 799
rect 5822 753 5855 799
rect 5976 796 6022 1108
rect 6136 796 6182 1108
rect 6424 796 6470 1108
rect 6569 805 6645 817
rect 5743 705 5855 753
rect 5743 659 5776 705
rect 5822 659 5855 705
rect 5743 611 5855 659
rect 6569 753 6581 805
rect 6633 753 6645 805
rect 6744 796 6790 1108
rect 7064 796 7110 1108
rect 7209 805 7285 817
rect 6569 701 6645 753
rect 6569 649 6581 701
rect 6633 649 6645 701
rect 6569 637 6645 649
rect 7209 753 7221 805
rect 7273 753 7285 805
rect 7384 796 7430 1108
rect 7672 796 7718 1108
rect 7832 796 7878 1108
rect 7999 1081 8111 1129
rect 8932 1266 9008 1278
rect 8932 1214 8944 1266
rect 8996 1214 9008 1266
rect 8932 1162 9008 1214
rect 8932 1110 8944 1162
rect 8996 1110 9008 1162
rect 8932 1098 9008 1110
rect 9828 1266 9904 1278
rect 9828 1214 9840 1266
rect 9892 1214 9904 1266
rect 9828 1162 9904 1214
rect 9828 1110 9840 1162
rect 9892 1110 9904 1162
rect 9828 1098 9904 1110
rect 10116 1266 10192 1278
rect 10116 1214 10128 1266
rect 10180 1214 10192 1266
rect 10116 1162 10192 1214
rect 10116 1110 10128 1162
rect 10180 1110 10192 1162
rect 10116 1098 10192 1110
rect 10725 1269 10837 1317
rect 10725 1223 10758 1269
rect 10804 1223 10837 1269
rect 10725 1175 10837 1223
rect 10725 1129 10758 1175
rect 10804 1129 10837 1175
rect 7999 1035 8032 1081
rect 8078 1035 8111 1081
rect 7999 987 8111 1035
rect 7999 941 8032 987
rect 8078 941 8111 987
rect 7999 893 8111 941
rect 7999 847 8032 893
rect 8078 847 8111 893
rect 7999 799 8111 847
rect 7209 701 7285 753
rect 7209 649 7221 701
rect 7273 649 7285 701
rect 7209 637 7285 649
rect 7999 753 8032 799
rect 8078 753 8111 799
rect 8211 777 8257 1089
rect 8371 777 8417 1089
rect 8787 1032 8833 1089
rect 9107 1032 9153 1089
rect 9683 1032 9729 1089
rect 10003 1032 10049 1089
rect 8787 986 10049 1032
rect 10003 880 10049 986
rect 8659 834 10177 880
rect 8659 777 8705 834
rect 9235 777 9281 834
rect 9555 777 9601 834
rect 10131 777 10177 834
rect 10419 777 10465 1089
rect 10579 777 10625 1089
rect 10725 1081 10837 1129
rect 10725 1035 10758 1081
rect 10804 1035 10837 1081
rect 10725 987 10837 1035
rect 10725 941 10758 987
rect 10804 941 10837 987
rect 10725 893 10837 941
rect 10725 847 10758 893
rect 10804 847 10837 893
rect 10725 799 10837 847
rect 7999 705 8111 753
rect 7999 659 8032 705
rect 8078 659 8111 705
rect 5743 565 5776 611
rect 5822 565 5855 611
rect 5743 517 5855 565
rect 5743 471 5776 517
rect 5822 471 5855 517
rect 5743 423 5855 471
rect 5743 377 5776 423
rect 5822 377 5855 423
rect 7999 611 8111 659
rect 10725 753 10758 799
rect 10804 753 10837 799
rect 10725 705 10837 753
rect 10725 659 10758 705
rect 10804 659 10837 705
rect 7999 565 8032 611
rect 8078 565 8111 611
rect 7999 517 8111 565
rect 7999 471 8032 517
rect 8078 471 8111 517
rect 7999 423 8111 471
rect 10116 604 10192 616
rect 10116 552 10128 604
rect 10180 552 10192 604
rect 10116 500 10192 552
rect 10116 448 10128 500
rect 10180 448 10192 500
rect 10116 436 10192 448
rect 10725 611 10837 659
rect 10725 565 10758 611
rect 10804 565 10837 611
rect 10725 517 10837 565
rect 10725 471 10758 517
rect 10804 471 10837 517
rect 5743 329 5855 377
rect 5743 283 5776 329
rect 5822 283 5855 329
rect 5743 235 5855 283
rect 6249 404 6325 416
rect 6249 352 6261 404
rect 6313 352 6325 404
rect 6249 300 6325 352
rect 6249 248 6261 300
rect 6313 248 6325 300
rect 5743 189 5776 235
rect 5822 189 5855 235
rect 5743 141 5855 189
rect 5743 95 5776 141
rect 5822 95 5855 141
rect 5743 47 5855 95
rect 5743 1 5776 47
rect 5822 1 5855 47
rect 5743 -47 5855 1
rect 5743 -93 5776 -47
rect 5822 -93 5855 -47
rect 5976 -66 6022 246
rect 6136 -66 6182 246
rect 6249 236 6325 248
rect 6889 404 6965 416
rect 6889 352 6901 404
rect 6953 352 6965 404
rect 6889 300 6965 352
rect 6889 248 6901 300
rect 6953 248 6965 300
rect 6424 -66 6470 246
rect 6744 -66 6790 246
rect 6889 236 6965 248
rect 7529 404 7605 416
rect 7529 352 7541 404
rect 7593 352 7605 404
rect 7529 300 7605 352
rect 7529 248 7541 300
rect 7593 248 7605 300
rect 7064 -66 7110 246
rect 7384 -66 7430 246
rect 7529 236 7605 248
rect 7999 377 8032 423
rect 8078 377 8111 423
rect 10725 423 10837 471
rect 7999 329 8111 377
rect 7999 283 8032 329
rect 8078 283 8111 329
rect 7672 -66 7718 246
rect 7832 -66 7878 246
rect 7999 235 8111 283
rect 8932 404 9008 416
rect 8932 352 8944 404
rect 8996 352 9008 404
rect 8932 300 9008 352
rect 8932 248 8944 300
rect 8996 248 9008 300
rect 8932 236 9008 248
rect 9828 404 9904 416
rect 9828 352 9840 404
rect 9892 352 9904 404
rect 9828 300 9904 352
rect 9828 248 9840 300
rect 9892 248 9904 300
rect 9828 236 9904 248
rect 10725 377 10758 423
rect 10804 377 10837 423
rect 10725 329 10837 377
rect 10725 283 10758 329
rect 10804 283 10837 329
rect 7999 189 8032 235
rect 8078 189 8111 235
rect 10725 235 10837 283
rect 7999 141 8111 189
rect 7999 95 8032 141
rect 8078 95 8111 141
rect 7999 47 8111 95
rect 7999 1 8032 47
rect 8078 1 8111 47
rect 7999 -47 8111 1
rect 5743 -141 5855 -93
rect 5743 -187 5776 -141
rect 5822 -187 5855 -141
rect 7999 -93 8032 -47
rect 8078 -93 8111 -47
rect 8211 -85 8257 227
rect 8371 -85 8417 227
rect 8499 -85 8545 227
rect 8659 -85 8705 227
rect 8787 -85 8833 227
rect 8947 -85 8993 227
rect 9107 -85 9153 227
rect 9235 -85 9281 227
rect 9395 -85 9441 227
rect 9555 -85 9601 227
rect 9683 -85 9729 227
rect 9843 -85 9889 227
rect 10003 -85 10049 227
rect 10131 -85 10177 227
rect 10291 -85 10337 227
rect 10419 -85 10465 227
rect 10579 -85 10625 227
rect 10725 189 10758 235
rect 10804 189 10837 235
rect 10725 141 10837 189
rect 10725 95 10758 141
rect 10804 95 10837 141
rect 10725 47 10837 95
rect 10725 1 10758 47
rect 10804 1 10837 47
rect 10725 -47 10837 1
rect 7999 -141 8111 -93
rect 5743 -235 5855 -187
rect 5743 -281 5776 -235
rect 5822 -281 5855 -235
rect 5743 -329 5855 -281
rect 5743 -375 5776 -329
rect 5822 -375 5855 -329
rect 6249 -196 6325 -184
rect 6249 -248 6261 -196
rect 6313 -248 6325 -196
rect 6249 -300 6325 -248
rect 6249 -352 6261 -300
rect 6313 -352 6325 -300
rect 6249 -364 6325 -352
rect 6889 -196 6965 -184
rect 6889 -248 6901 -196
rect 6953 -248 6965 -196
rect 6889 -300 6965 -248
rect 6889 -352 6901 -300
rect 6953 -352 6965 -300
rect 6889 -364 6965 -352
rect 7529 -196 7605 -184
rect 7529 -248 7541 -196
rect 7593 -248 7605 -196
rect 7529 -300 7605 -248
rect 7529 -352 7541 -300
rect 7593 -352 7605 -300
rect 7529 -364 7605 -352
rect 7999 -187 8032 -141
rect 8078 -187 8111 -141
rect 10725 -93 10758 -47
rect 10804 -93 10837 -47
rect 10725 -141 10837 -93
rect 7999 -235 8111 -187
rect 7999 -281 8032 -235
rect 8078 -281 8111 -235
rect 7999 -329 8111 -281
rect 5743 -423 5855 -375
rect 5743 -469 5776 -423
rect 5822 -469 5855 -423
rect 7999 -375 8032 -329
rect 8078 -375 8111 -329
rect 8484 -196 8560 -184
rect 8484 -248 8496 -196
rect 8548 -248 8560 -196
rect 8484 -300 8560 -248
rect 8484 -352 8496 -300
rect 8548 -352 8560 -300
rect 8484 -364 8560 -352
rect 9380 -196 9456 -184
rect 9380 -248 9392 -196
rect 9444 -248 9456 -196
rect 9380 -300 9456 -248
rect 9380 -352 9392 -300
rect 9444 -352 9456 -300
rect 9380 -364 9456 -352
rect 10276 -196 10352 -184
rect 10276 -248 10288 -196
rect 10340 -248 10352 -196
rect 10276 -300 10352 -248
rect 10276 -352 10288 -300
rect 10340 -352 10352 -300
rect 10276 -364 10352 -352
rect 10725 -187 10758 -141
rect 10804 -187 10837 -141
rect 10725 -235 10837 -187
rect 10725 -281 10758 -235
rect 10804 -281 10837 -235
rect 10725 -329 10837 -281
rect 7999 -423 8111 -375
rect 5743 -517 5855 -469
rect 5743 -563 5776 -517
rect 5822 -563 5855 -517
rect 5743 -611 5855 -563
rect 5743 -657 5776 -611
rect 5822 -657 5855 -611
rect 6569 -469 6645 -457
rect 6569 -521 6581 -469
rect 6633 -521 6645 -469
rect 6569 -573 6645 -521
rect 5743 -705 5855 -657
rect 5743 -751 5776 -705
rect 5822 -751 5855 -705
rect 5743 -799 5855 -751
rect 5743 -845 5776 -799
rect 5822 -845 5855 -799
rect 5743 -893 5855 -845
rect 5743 -939 5776 -893
rect 5822 -939 5855 -893
rect 5976 -749 6022 -616
rect 6136 -749 6182 -616
rect 5976 -795 6056 -749
rect 6102 -795 6182 -749
rect 5976 -928 6022 -795
rect 6136 -928 6182 -795
rect 6424 -928 6470 -616
rect 6569 -625 6581 -573
rect 6633 -625 6645 -573
rect 7209 -469 7285 -457
rect 7209 -521 7221 -469
rect 7273 -521 7285 -469
rect 7209 -573 7285 -521
rect 6569 -637 6645 -625
rect 5743 -987 5855 -939
rect 5743 -1033 5776 -987
rect 5822 -1033 5855 -987
rect 5743 -1081 5855 -1033
rect 5743 -1127 5776 -1081
rect 5822 -1127 5855 -1081
rect 6569 -934 6645 -922
rect 6744 -928 6790 -616
rect 7064 -928 7110 -616
rect 7209 -625 7221 -573
rect 7273 -625 7285 -573
rect 7999 -469 8032 -423
rect 8078 -469 8111 -423
rect 10725 -375 10758 -329
rect 10804 -375 10837 -329
rect 10725 -423 10837 -375
rect 7999 -517 8111 -469
rect 7999 -563 8032 -517
rect 8078 -563 8111 -517
rect 7999 -611 8111 -563
rect 7209 -637 7285 -625
rect 6569 -986 6581 -934
rect 6633 -986 6645 -934
rect 6569 -1038 6645 -986
rect 6569 -1090 6581 -1038
rect 6633 -1090 6645 -1038
rect 6569 -1102 6645 -1090
rect 7209 -934 7285 -922
rect 7384 -928 7430 -616
rect 7503 -693 7579 -681
rect 7503 -745 7515 -693
rect 7567 -745 7579 -693
rect 7503 -797 7579 -745
rect 7503 -849 7515 -797
rect 7567 -849 7579 -797
rect 7503 -861 7579 -849
rect 7672 -749 7718 -616
rect 7832 -749 7878 -616
rect 7672 -795 7752 -749
rect 7798 -795 7878 -749
rect 7672 -928 7718 -795
rect 7832 -928 7878 -795
rect 7999 -657 8032 -611
rect 8078 -657 8111 -611
rect 9988 -454 10064 -442
rect 9988 -506 10000 -454
rect 10052 -506 10064 -454
rect 9988 -558 10064 -506
rect 9988 -610 10000 -558
rect 10052 -610 10064 -558
rect 9988 -622 10064 -610
rect 10725 -469 10758 -423
rect 10804 -469 10837 -423
rect 10725 -517 10837 -469
rect 10725 -563 10758 -517
rect 10804 -563 10837 -517
rect 10725 -611 10837 -563
rect 7999 -705 8111 -657
rect 7999 -751 8032 -705
rect 8078 -751 8111 -705
rect 7999 -799 8111 -751
rect 7999 -845 8032 -799
rect 8078 -845 8111 -799
rect 7999 -893 8111 -845
rect 7209 -986 7221 -934
rect 7273 -986 7285 -934
rect 7209 -1038 7285 -986
rect 7209 -1090 7221 -1038
rect 7273 -1090 7285 -1038
rect 7209 -1102 7285 -1090
rect 7999 -939 8032 -893
rect 8078 -939 8111 -893
rect 7999 -987 8111 -939
rect 8211 -768 8257 -635
rect 8371 -768 8417 -635
rect 8787 -692 8833 -635
rect 9107 -692 9153 -635
rect 9683 -692 9729 -635
rect 10003 -692 10049 -635
rect 8787 -738 10049 -692
rect 8211 -814 8291 -768
rect 8337 -814 8417 -768
rect 8211 -947 8257 -814
rect 8371 -947 8417 -814
rect 10003 -830 10049 -738
rect 10236 -704 10312 -692
rect 10236 -756 10248 -704
rect 10300 -756 10312 -704
rect 10236 -808 10312 -756
rect 8659 -876 10177 -830
rect 10236 -860 10248 -808
rect 10300 -860 10312 -808
rect 10236 -872 10312 -860
rect 10419 -768 10465 -635
rect 10579 -768 10625 -635
rect 10419 -814 10499 -768
rect 10545 -814 10625 -768
rect 8659 -947 8705 -876
rect 8932 -934 9008 -922
rect 7999 -1033 8032 -987
rect 8078 -1033 8111 -987
rect 7999 -1081 8111 -1033
rect 5743 -1175 5855 -1127
rect 5743 -1221 5776 -1175
rect 5822 -1221 5855 -1175
rect 5743 -1269 5855 -1221
rect 5743 -1315 5776 -1269
rect 5822 -1315 5855 -1269
rect 7999 -1127 8032 -1081
rect 8078 -1127 8111 -1081
rect 8932 -986 8944 -934
rect 8996 -986 9008 -934
rect 9235 -947 9281 -876
rect 9555 -947 9601 -876
rect 9828 -934 9904 -922
rect 9683 -937 9729 -936
rect 8932 -1038 9008 -986
rect 8932 -1090 8944 -1038
rect 8996 -1090 9008 -1038
rect 8932 -1102 9008 -1090
rect 9828 -986 9840 -934
rect 9892 -986 9904 -934
rect 9828 -1038 9904 -986
rect 9828 -1090 9840 -1038
rect 9892 -1090 9904 -1038
rect 9828 -1102 9904 -1090
rect 9988 -934 10064 -922
rect 9988 -986 10000 -934
rect 10052 -986 10064 -934
rect 10131 -947 10177 -876
rect 10419 -947 10465 -814
rect 10579 -947 10625 -814
rect 10725 -657 10758 -611
rect 10804 -657 10837 -611
rect 10725 -705 10837 -657
rect 10725 -751 10758 -705
rect 10804 -751 10837 -705
rect 10725 -799 10837 -751
rect 10725 -845 10758 -799
rect 10804 -845 10837 -799
rect 10725 -893 10837 -845
rect 10725 -939 10758 -893
rect 10804 -939 10837 -893
rect 9988 -1038 10064 -986
rect 9988 -1090 10000 -1038
rect 10052 -1090 10064 -1038
rect 9988 -1102 10064 -1090
rect 10725 -987 10837 -939
rect 10725 -1033 10758 -987
rect 10804 -1033 10837 -987
rect 10725 -1081 10837 -1033
rect 7999 -1175 8111 -1127
rect 7999 -1221 8032 -1175
rect 8078 -1221 8111 -1175
rect 7999 -1269 8111 -1221
rect 5743 -1363 5855 -1315
rect 5743 -1409 5776 -1363
rect 5822 -1409 5855 -1363
rect 5743 -1457 5855 -1409
rect 5743 -1503 5776 -1457
rect 5822 -1503 5855 -1457
rect 6249 -1326 6325 -1314
rect 6249 -1378 6261 -1326
rect 6313 -1378 6325 -1326
rect 6249 -1430 6325 -1378
rect 5743 -1551 5855 -1503
rect 5743 -1597 5776 -1551
rect 5822 -1597 5855 -1551
rect 5743 -1645 5855 -1597
rect 5743 -1691 5776 -1645
rect 5822 -1691 5855 -1645
rect 5743 -1739 5855 -1691
rect 5743 -1785 5776 -1739
rect 5822 -1776 5855 -1739
rect 5976 -1776 6022 -1478
rect 6136 -1776 6182 -1478
rect 6249 -1482 6261 -1430
rect 6313 -1482 6325 -1430
rect 6889 -1326 6965 -1314
rect 6889 -1378 6901 -1326
rect 6953 -1378 6965 -1326
rect 6889 -1430 6965 -1378
rect 6249 -1494 6325 -1482
rect 6424 -1766 6470 -1478
rect 6381 -1776 6561 -1766
rect 6744 -1776 6790 -1478
rect 6889 -1482 6901 -1430
rect 6953 -1482 6965 -1430
rect 7529 -1326 7605 -1314
rect 7529 -1378 7541 -1326
rect 7593 -1378 7605 -1326
rect 7529 -1430 7605 -1378
rect 6889 -1494 6965 -1482
rect 7064 -1776 7110 -1478
rect 7384 -1776 7430 -1478
rect 7529 -1482 7541 -1430
rect 7593 -1482 7605 -1430
rect 7999 -1315 8032 -1269
rect 8078 -1315 8111 -1269
rect 10725 -1127 10758 -1081
rect 10804 -1127 10837 -1081
rect 10725 -1175 10837 -1127
rect 10725 -1221 10758 -1175
rect 10804 -1221 10837 -1175
rect 10725 -1269 10837 -1221
rect 7999 -1363 8111 -1315
rect 7999 -1409 8032 -1363
rect 8078 -1409 8111 -1363
rect 7999 -1457 8111 -1409
rect 7529 -1494 7605 -1482
rect 7672 -1776 7718 -1478
rect 7832 -1776 7878 -1478
rect 7999 -1503 8032 -1457
rect 8078 -1503 8111 -1457
rect 8484 -1326 8560 -1314
rect 8484 -1378 8496 -1326
rect 8548 -1378 8560 -1326
rect 8484 -1430 8560 -1378
rect 8484 -1482 8496 -1430
rect 8548 -1482 8560 -1430
rect 7999 -1551 8111 -1503
rect 7999 -1597 8032 -1551
rect 8078 -1597 8111 -1551
rect 7999 -1645 8111 -1597
rect 7999 -1691 8032 -1645
rect 8078 -1691 8111 -1645
rect 7999 -1739 8111 -1691
rect 7999 -1776 8032 -1739
rect 5822 -1778 8032 -1776
rect 5822 -1785 6393 -1778
rect 5743 -1830 6393 -1785
rect 6445 -1830 6497 -1778
rect 6549 -1785 8032 -1778
rect 8078 -1776 8111 -1739
rect 8211 -1776 8257 -1484
rect 8371 -1776 8417 -1484
rect 8484 -1494 8560 -1482
rect 9380 -1326 9456 -1314
rect 9380 -1378 9392 -1326
rect 9444 -1378 9456 -1326
rect 9380 -1430 9456 -1378
rect 9380 -1482 9392 -1430
rect 9444 -1482 9456 -1430
rect 9380 -1494 9456 -1482
rect 10276 -1326 10352 -1314
rect 10276 -1378 10288 -1326
rect 10340 -1378 10352 -1326
rect 10276 -1430 10352 -1378
rect 10276 -1482 10288 -1430
rect 10340 -1482 10352 -1430
rect 10276 -1494 10352 -1482
rect 10725 -1315 10758 -1269
rect 10804 -1315 10837 -1269
rect 10725 -1363 10837 -1315
rect 10725 -1409 10758 -1363
rect 10804 -1409 10837 -1363
rect 10725 -1457 10837 -1409
rect 8787 -1554 8833 -1497
rect 9107 -1554 9153 -1497
rect 9683 -1554 9729 -1497
rect 10003 -1554 10049 -1497
rect 8787 -1600 10049 -1554
rect 9483 -1776 9663 -1766
rect 10419 -1776 10465 -1497
rect 10579 -1776 10625 -1497
rect 10725 -1503 10758 -1457
rect 10804 -1503 10837 -1457
rect 10725 -1551 10837 -1503
rect 10725 -1597 10758 -1551
rect 10804 -1597 10837 -1551
rect 10725 -1645 10837 -1597
rect 10725 -1691 10758 -1645
rect 10804 -1691 10837 -1645
rect 10725 -1739 10837 -1691
rect 10725 -1776 10758 -1739
rect 8078 -1778 10758 -1776
rect 8078 -1785 9495 -1778
rect 6549 -1830 9495 -1785
rect 9547 -1830 9599 -1778
rect 9651 -1785 10758 -1778
rect 10804 -1785 10837 -1739
rect 9651 -1830 10837 -1785
rect 5743 -1833 10837 -1830
rect 5743 -1879 5776 -1833
rect 5822 -1879 5870 -1833
rect 5916 -1879 5964 -1833
rect 6010 -1879 6058 -1833
rect 6104 -1879 6152 -1833
rect 6198 -1879 6246 -1833
rect 6292 -1879 6340 -1833
rect 6386 -1879 6434 -1833
rect 6480 -1879 6528 -1833
rect 6574 -1879 6622 -1833
rect 6668 -1879 6716 -1833
rect 6762 -1879 6810 -1833
rect 6856 -1879 6904 -1833
rect 6950 -1879 6998 -1833
rect 7044 -1879 7092 -1833
rect 7138 -1879 7186 -1833
rect 7232 -1879 7280 -1833
rect 7326 -1879 7374 -1833
rect 7420 -1879 7468 -1833
rect 7514 -1879 7562 -1833
rect 7608 -1879 7656 -1833
rect 7702 -1879 7750 -1833
rect 7796 -1879 7844 -1833
rect 7890 -1879 7938 -1833
rect 7984 -1879 8032 -1833
rect 8078 -1879 8126 -1833
rect 8172 -1879 8220 -1833
rect 8266 -1879 8314 -1833
rect 8360 -1879 8408 -1833
rect 8454 -1879 8502 -1833
rect 8548 -1879 8596 -1833
rect 8642 -1879 8690 -1833
rect 8736 -1879 8784 -1833
rect 8830 -1879 8878 -1833
rect 8924 -1879 8972 -1833
rect 9018 -1879 9066 -1833
rect 9112 -1879 9160 -1833
rect 9206 -1879 9254 -1833
rect 9300 -1879 9348 -1833
rect 9394 -1879 9442 -1833
rect 9488 -1879 9536 -1833
rect 9582 -1879 9630 -1833
rect 9676 -1879 9724 -1833
rect 9770 -1879 9818 -1833
rect 9864 -1879 9912 -1833
rect 9958 -1879 10006 -1833
rect 10052 -1879 10100 -1833
rect 10146 -1879 10194 -1833
rect 10240 -1879 10288 -1833
rect 10334 -1879 10382 -1833
rect 10428 -1879 10476 -1833
rect 10522 -1879 10570 -1833
rect 10616 -1879 10664 -1833
rect 10710 -1879 10758 -1833
rect 10804 -1879 10837 -1833
rect 5743 -1882 10837 -1879
rect 5743 -1934 6393 -1882
rect 6445 -1934 6497 -1882
rect 6549 -1934 9495 -1882
rect 9547 -1934 9599 -1882
rect 9651 -1934 10837 -1882
rect 5743 -1936 10837 -1934
rect 11381 1599 11414 1645
rect 11460 1599 11493 1645
rect 11866 1796 11942 1808
rect 11866 1744 11878 1796
rect 11930 1744 11942 1796
rect 11866 1692 11942 1744
rect 11866 1640 11878 1692
rect 11930 1640 11942 1692
rect 11866 1628 11942 1640
rect 12762 1796 12838 1808
rect 12762 1744 12774 1796
rect 12826 1744 12838 1796
rect 12762 1692 12838 1744
rect 12762 1640 12774 1692
rect 12826 1640 12838 1692
rect 12762 1628 12838 1640
rect 13658 1796 13734 1808
rect 13658 1744 13670 1796
rect 13722 1744 13734 1796
rect 13658 1692 13734 1744
rect 13658 1640 13670 1692
rect 13722 1640 13734 1692
rect 13658 1628 13734 1640
rect 14107 1787 14140 1833
rect 14186 1787 14219 1833
rect 16457 2021 16569 2069
rect 16457 1975 16490 2021
rect 16536 1975 16569 2021
rect 16457 1927 16569 1975
rect 16457 1881 16490 1927
rect 16536 1881 16569 1927
rect 16457 1833 16569 1881
rect 14107 1739 14219 1787
rect 14107 1693 14140 1739
rect 14186 1693 14219 1739
rect 14107 1645 14219 1693
rect 11381 1551 11493 1599
rect 11381 1505 11414 1551
rect 11460 1505 11493 1551
rect 11381 1457 11493 1505
rect 11381 1411 11414 1457
rect 11460 1411 11493 1457
rect 11381 1363 11493 1411
rect 11381 1317 11414 1363
rect 11460 1317 11493 1363
rect 11381 1269 11493 1317
rect 11381 1223 11414 1269
rect 11460 1223 11493 1269
rect 11381 1175 11493 1223
rect 11381 1129 11414 1175
rect 11460 1129 11493 1175
rect 11593 1171 11639 1607
rect 11753 1171 11799 1607
rect 12169 1527 12215 1607
rect 12489 1527 12535 1607
rect 13065 1527 13111 1607
rect 13385 1527 13431 1607
rect 12169 1481 13431 1527
rect 13385 1297 13431 1481
rect 12041 1251 13559 1297
rect 12041 1171 12087 1251
rect 12169 1171 12215 1182
rect 11381 1081 11493 1129
rect 11381 1035 11414 1081
rect 11460 1035 11493 1081
rect 11381 987 11493 1035
rect 12314 1162 12390 1174
rect 12489 1171 12535 1182
rect 12617 1171 12663 1251
rect 12777 1171 12823 1182
rect 12937 1171 12983 1251
rect 13065 1171 13111 1182
rect 12314 1110 12326 1162
rect 12378 1110 12390 1162
rect 12314 1058 12390 1110
rect 12314 1006 12326 1058
rect 12378 1006 12390 1058
rect 12314 994 12390 1006
rect 13210 1162 13286 1174
rect 13385 1171 13431 1182
rect 13513 1171 13559 1251
rect 13801 1171 13847 1607
rect 13961 1171 14007 1607
rect 14107 1599 14140 1645
rect 14186 1599 14219 1645
rect 14980 1796 15056 1808
rect 14980 1744 14992 1796
rect 15044 1744 15056 1796
rect 14980 1692 15056 1744
rect 14980 1640 14992 1692
rect 15044 1640 15056 1692
rect 14980 1628 15056 1640
rect 15620 1796 15696 1808
rect 15620 1744 15632 1796
rect 15684 1744 15696 1796
rect 15620 1692 15696 1744
rect 15620 1640 15632 1692
rect 15684 1640 15696 1692
rect 15620 1628 15696 1640
rect 16457 1787 16490 1833
rect 16536 1787 16569 1833
rect 16627 1808 16787 2470
rect 16889 2228 17049 2518
rect 17569 2497 17650 2543
rect 17696 2497 17889 2543
rect 17569 2449 17889 2497
rect 17569 2403 17650 2449
rect 17696 2403 17889 2449
rect 17569 2355 17889 2403
rect 17569 2309 17650 2355
rect 17696 2309 17889 2355
rect 17569 2261 17889 2309
rect 16879 2216 17059 2228
rect 16879 2164 16891 2216
rect 16943 2164 16995 2216
rect 17047 2164 17059 2216
rect 16879 2112 17059 2164
rect 16879 2060 16891 2112
rect 16943 2060 16995 2112
rect 17047 2060 17059 2112
rect 16879 2048 17059 2060
rect 17569 2215 17650 2261
rect 17696 2215 17889 2261
rect 17569 2167 17889 2215
rect 17569 2121 17650 2167
rect 17696 2121 17889 2167
rect 17569 2073 17889 2121
rect 17569 2027 17650 2073
rect 17696 2027 17889 2073
rect 17569 1979 17889 2027
rect 17569 1933 17650 1979
rect 17696 1933 17889 1979
rect 17569 1885 17889 1933
rect 17569 1839 17650 1885
rect 17696 1839 17889 1885
rect 16457 1739 16569 1787
rect 16457 1693 16490 1739
rect 16536 1693 16569 1739
rect 16457 1645 16569 1693
rect 14107 1551 14219 1599
rect 14107 1505 14140 1551
rect 14186 1505 14219 1551
rect 14107 1457 14219 1505
rect 14107 1411 14140 1457
rect 14186 1411 14219 1457
rect 14107 1363 14219 1411
rect 14107 1317 14140 1363
rect 14186 1317 14219 1363
rect 14107 1269 14219 1317
rect 14107 1223 14140 1269
rect 14186 1223 14219 1269
rect 14107 1175 14219 1223
rect 13210 1110 13222 1162
rect 13274 1110 13286 1162
rect 13210 1058 13286 1110
rect 13210 1006 13222 1058
rect 13274 1006 13286 1058
rect 13210 994 13286 1006
rect 13498 1136 13574 1148
rect 13498 1084 13510 1136
rect 13562 1084 13574 1136
rect 13498 1032 13574 1084
rect 11381 941 11414 987
rect 11460 941 11493 987
rect 13498 980 13510 1032
rect 13562 980 13574 1032
rect 13498 968 13574 980
rect 14107 1129 14140 1175
rect 14186 1129 14219 1175
rect 14387 1171 14433 1607
rect 14547 1171 14593 1607
rect 14835 1171 14881 1607
rect 15155 1171 15201 1607
rect 15475 1171 15521 1607
rect 15795 1171 15841 1607
rect 16083 1171 16129 1607
rect 16243 1171 16289 1607
rect 16457 1599 16490 1645
rect 16536 1599 16569 1645
rect 16617 1796 16797 1808
rect 16617 1744 16629 1796
rect 16681 1744 16733 1796
rect 16785 1744 16797 1796
rect 16617 1692 16797 1744
rect 16617 1640 16629 1692
rect 16681 1640 16733 1692
rect 16785 1640 16797 1692
rect 16617 1628 16797 1640
rect 17569 1791 17889 1839
rect 17569 1745 17650 1791
rect 17696 1745 17889 1791
rect 17569 1697 17889 1745
rect 17569 1651 17650 1697
rect 17696 1651 17889 1697
rect 16457 1551 16569 1599
rect 16457 1505 16490 1551
rect 16536 1505 16569 1551
rect 16457 1457 16569 1505
rect 16457 1411 16490 1457
rect 16536 1411 16569 1457
rect 16457 1363 16569 1411
rect 16457 1317 16490 1363
rect 16536 1317 16569 1363
rect 16457 1269 16569 1317
rect 16457 1223 16490 1269
rect 16536 1223 16569 1269
rect 16457 1175 16569 1223
rect 14107 1081 14219 1129
rect 14107 1035 14140 1081
rect 14186 1035 14219 1081
rect 14107 987 14219 1035
rect 11381 893 11493 941
rect 11381 847 11414 893
rect 11460 847 11493 893
rect 11381 799 11493 847
rect 11381 753 11414 799
rect 11460 753 11493 799
rect 11381 705 11493 753
rect 11381 659 11414 705
rect 11460 659 11493 705
rect 11381 611 11493 659
rect 11381 565 11414 611
rect 11460 565 11493 611
rect 14107 941 14140 987
rect 14186 941 14219 987
rect 14660 1136 14736 1148
rect 14660 1084 14672 1136
rect 14724 1084 14736 1136
rect 14660 1032 14736 1084
rect 14660 980 14672 1032
rect 14724 980 14736 1032
rect 14660 968 14736 980
rect 15300 1136 15376 1148
rect 15300 1084 15312 1136
rect 15364 1084 15376 1136
rect 15300 1032 15376 1084
rect 15300 980 15312 1032
rect 15364 980 15376 1032
rect 15300 968 15376 980
rect 15940 1136 16016 1148
rect 15940 1084 15952 1136
rect 16004 1084 16016 1136
rect 15940 1032 16016 1084
rect 15940 980 15952 1032
rect 16004 980 16016 1032
rect 15940 968 16016 980
rect 16457 1129 16490 1175
rect 16536 1129 16569 1175
rect 16457 1081 16569 1129
rect 16457 1035 16490 1081
rect 16536 1035 16569 1081
rect 16457 987 16569 1035
rect 14107 893 14219 941
rect 14107 847 14140 893
rect 14186 847 14219 893
rect 14107 799 14219 847
rect 14107 753 14140 799
rect 14186 753 14219 799
rect 14107 705 14219 753
rect 14107 659 14140 705
rect 14186 659 14219 705
rect 14107 611 14219 659
rect 11381 517 11493 565
rect 11381 471 11414 517
rect 11460 471 11493 517
rect 11381 423 11493 471
rect 11381 377 11414 423
rect 11460 377 11493 423
rect 11381 329 11493 377
rect 11381 283 11414 329
rect 11460 283 11493 329
rect 11381 235 11493 283
rect 11381 189 11414 235
rect 11460 189 11493 235
rect 11381 141 11493 189
rect 11381 95 11414 141
rect 11460 95 11493 141
rect 11593 135 11639 571
rect 11753 135 11799 571
rect 11881 135 11927 571
rect 12041 135 12087 571
rect 12169 135 12215 571
rect 12329 135 12375 571
rect 12489 135 12535 571
rect 12617 135 12663 571
rect 12777 135 12823 571
rect 12937 135 12983 571
rect 13065 135 13111 571
rect 13225 135 13271 571
rect 13385 135 13431 571
rect 13513 135 13559 571
rect 13673 135 13719 571
rect 13801 135 13847 571
rect 13961 135 14007 571
rect 14107 565 14140 611
rect 14186 565 14219 611
rect 16457 941 16490 987
rect 16536 941 16569 987
rect 16457 893 16569 941
rect 16457 847 16490 893
rect 16536 847 16569 893
rect 16457 799 16569 847
rect 16457 753 16490 799
rect 16536 753 16569 799
rect 16457 705 16569 753
rect 16457 659 16490 705
rect 16536 659 16569 705
rect 16457 611 16569 659
rect 14107 517 14219 565
rect 14107 471 14140 517
rect 14186 471 14219 517
rect 14107 423 14219 471
rect 14107 377 14140 423
rect 14186 377 14219 423
rect 14107 329 14219 377
rect 14107 283 14140 329
rect 14186 283 14219 329
rect 14107 235 14219 283
rect 14107 189 14140 235
rect 14186 189 14219 235
rect 14107 141 14219 189
rect 11381 47 11493 95
rect 11381 1 11414 47
rect 11460 1 11493 47
rect 11381 -47 11493 1
rect 11381 -93 11414 -47
rect 11460 -93 11493 -47
rect 11866 116 11942 128
rect 11866 64 11878 116
rect 11930 64 11942 116
rect 11866 12 11942 64
rect 11866 -40 11878 12
rect 11930 -40 11942 12
rect 11866 -52 11942 -40
rect 12762 116 12838 128
rect 12762 64 12774 116
rect 12826 64 12838 116
rect 12762 12 12838 64
rect 12762 -40 12774 12
rect 12826 -40 12838 12
rect 12762 -52 12838 -40
rect 13658 116 13734 128
rect 13658 64 13670 116
rect 13722 64 13734 116
rect 13658 12 13734 64
rect 13658 -40 13670 12
rect 13722 -40 13734 12
rect 13658 -52 13734 -40
rect 14107 95 14140 141
rect 14186 95 14219 141
rect 14387 135 14433 571
rect 14547 135 14593 571
rect 14675 135 14721 571
rect 14835 135 14881 571
rect 14995 135 15041 571
rect 15155 135 15201 571
rect 15315 135 15361 571
rect 15475 135 15521 571
rect 15635 135 15681 571
rect 15795 135 15841 571
rect 15955 135 16001 571
rect 16083 135 16129 571
rect 16243 135 16289 571
rect 16457 565 16490 611
rect 16536 565 16569 611
rect 16457 517 16569 565
rect 16457 471 16490 517
rect 16536 471 16569 517
rect 16457 423 16569 471
rect 16457 377 16490 423
rect 16536 377 16569 423
rect 16457 329 16569 377
rect 16457 283 16490 329
rect 16536 283 16569 329
rect 16457 235 16569 283
rect 16457 189 16490 235
rect 16536 189 16569 235
rect 16457 141 16569 189
rect 14107 47 14219 95
rect 14107 1 14140 47
rect 14186 1 14219 47
rect 14107 -47 14219 1
rect 11381 -141 11493 -93
rect 11381 -187 11414 -141
rect 11460 -187 11493 -141
rect 11381 -235 11493 -187
rect 11381 -281 11414 -235
rect 11460 -281 11493 -235
rect 14107 -93 14140 -47
rect 14186 -93 14219 -47
rect 14107 -141 14219 -93
rect 14107 -187 14140 -141
rect 14186 -187 14219 -141
rect 14107 -235 14219 -187
rect 11381 -329 11493 -281
rect 11381 -375 11414 -329
rect 11460 -375 11493 -329
rect 11381 -423 11493 -375
rect 11381 -469 11414 -423
rect 11460 -469 11493 -423
rect 13370 -284 13446 -272
rect 13370 -336 13382 -284
rect 13434 -336 13446 -284
rect 13370 -388 13446 -336
rect 13370 -440 13382 -388
rect 13434 -440 13446 -388
rect 13370 -452 13446 -440
rect 14107 -281 14140 -235
rect 14186 -281 14219 -235
rect 16457 95 16490 141
rect 16536 95 16569 141
rect 16457 47 16569 95
rect 16457 1 16490 47
rect 16536 1 16569 47
rect 16457 -47 16569 1
rect 16457 -93 16490 -47
rect 16536 -93 16569 -47
rect 16457 -141 16569 -93
rect 16457 -187 16490 -141
rect 16536 -187 16569 -141
rect 16457 -235 16569 -187
rect 14107 -329 14219 -281
rect 14107 -375 14140 -329
rect 14186 -375 14219 -329
rect 14107 -423 14219 -375
rect 11381 -517 11493 -469
rect 11381 -563 11414 -517
rect 11460 -563 11493 -517
rect 11381 -611 11493 -563
rect 11381 -657 11414 -611
rect 11460 -657 11493 -611
rect 11381 -705 11493 -657
rect 11381 -751 11414 -705
rect 11460 -751 11493 -705
rect 11381 -799 11493 -751
rect 11381 -845 11414 -799
rect 11460 -845 11493 -799
rect 11381 -893 11493 -845
rect 11381 -939 11414 -893
rect 11460 -939 11493 -893
rect 11593 -722 11639 -465
rect 11753 -722 11799 -465
rect 12169 -545 12215 -465
rect 12489 -545 12535 -465
rect 13065 -545 13111 -465
rect 13385 -545 13431 -465
rect 11593 -768 11673 -722
rect 11719 -768 11799 -722
rect 11902 -594 11978 -582
rect 12169 -591 13431 -545
rect 11902 -646 11914 -594
rect 11966 -646 11978 -594
rect 11902 -698 11978 -646
rect 11902 -750 11914 -698
rect 11966 -750 11978 -698
rect 11902 -762 11978 -750
rect 11593 -901 11639 -768
rect 11753 -901 11799 -768
rect 13385 -775 13431 -591
rect 13801 -722 13847 -465
rect 13961 -722 14007 -465
rect 13801 -768 13881 -722
rect 13927 -768 14007 -722
rect 12041 -821 13559 -775
rect 12041 -901 12087 -821
rect 12169 -901 12215 -890
rect 12489 -901 12535 -890
rect 12617 -901 12663 -821
rect 12777 -901 12823 -890
rect 12937 -901 12983 -821
rect 13065 -901 13111 -890
rect 13385 -901 13431 -890
rect 13513 -901 13559 -821
rect 13801 -901 13847 -768
rect 13961 -901 14007 -768
rect 14107 -469 14140 -423
rect 14186 -469 14219 -423
rect 14980 -284 15056 -272
rect 14980 -336 14992 -284
rect 15044 -336 15056 -284
rect 14980 -388 15056 -336
rect 14980 -440 14992 -388
rect 15044 -440 15056 -388
rect 14980 -452 15056 -440
rect 15620 -284 15696 -272
rect 15620 -336 15632 -284
rect 15684 -336 15696 -284
rect 15620 -388 15696 -336
rect 15620 -440 15632 -388
rect 15684 -440 15696 -388
rect 15620 -452 15696 -440
rect 16457 -281 16490 -235
rect 16536 -281 16569 -235
rect 16457 -329 16569 -281
rect 16457 -375 16490 -329
rect 16536 -375 16569 -329
rect 16457 -423 16569 -375
rect 14107 -517 14219 -469
rect 14107 -563 14140 -517
rect 14186 -563 14219 -517
rect 14107 -611 14219 -563
rect 14107 -657 14140 -611
rect 14186 -657 14219 -611
rect 14107 -705 14219 -657
rect 14107 -751 14140 -705
rect 14186 -751 14219 -705
rect 14107 -799 14219 -751
rect 14107 -845 14140 -799
rect 14186 -845 14219 -799
rect 14107 -893 14219 -845
rect 11381 -987 11493 -939
rect 11381 -1033 11414 -987
rect 11460 -1033 11493 -987
rect 11381 -1081 11493 -1033
rect 11381 -1127 11414 -1081
rect 11460 -1127 11493 -1081
rect 12314 -934 12390 -922
rect 12314 -986 12326 -934
rect 12378 -986 12390 -934
rect 12314 -1038 12390 -986
rect 12314 -1090 12326 -1038
rect 12378 -1090 12390 -1038
rect 12314 -1102 12390 -1090
rect 13210 -934 13286 -922
rect 13210 -986 13222 -934
rect 13274 -986 13286 -934
rect 13210 -1038 13286 -986
rect 13210 -1090 13222 -1038
rect 13274 -1090 13286 -1038
rect 13210 -1102 13286 -1090
rect 13370 -934 13446 -922
rect 13370 -986 13382 -934
rect 13434 -986 13446 -934
rect 13370 -1038 13446 -986
rect 13370 -1090 13382 -1038
rect 13434 -1090 13446 -1038
rect 13370 -1102 13446 -1090
rect 14107 -939 14140 -893
rect 14186 -939 14219 -893
rect 14387 -722 14433 -465
rect 14547 -722 14593 -465
rect 14387 -768 14467 -722
rect 14513 -768 14593 -722
rect 14688 -589 14764 -577
rect 14688 -641 14700 -589
rect 14752 -641 14764 -589
rect 14688 -693 14764 -641
rect 14688 -745 14700 -693
rect 14752 -745 14764 -693
rect 14688 -757 14764 -745
rect 14387 -901 14433 -768
rect 14547 -901 14593 -768
rect 14835 -901 14881 -465
rect 15155 -901 15201 -465
rect 15475 -901 15521 -465
rect 15795 -901 15841 -465
rect 16083 -722 16129 -465
rect 16243 -722 16289 -465
rect 16083 -768 16163 -722
rect 16209 -768 16289 -722
rect 16083 -901 16129 -768
rect 16243 -901 16289 -768
rect 16457 -469 16490 -423
rect 16536 -469 16569 -423
rect 16457 -517 16569 -469
rect 16457 -563 16490 -517
rect 16536 -563 16569 -517
rect 16457 -611 16569 -563
rect 16457 -657 16490 -611
rect 16536 -657 16569 -611
rect 16457 -705 16569 -657
rect 16457 -751 16490 -705
rect 16536 -751 16569 -705
rect 16457 -799 16569 -751
rect 16457 -845 16490 -799
rect 16536 -845 16569 -799
rect 16457 -893 16569 -845
rect 14107 -987 14219 -939
rect 14107 -1033 14140 -987
rect 14186 -1033 14219 -987
rect 14107 -1081 14219 -1033
rect 11381 -1175 11493 -1127
rect 11381 -1221 11414 -1175
rect 11460 -1221 11493 -1175
rect 11381 -1269 11493 -1221
rect 11381 -1315 11414 -1269
rect 11460 -1315 11493 -1269
rect 11381 -1363 11493 -1315
rect 14107 -1127 14140 -1081
rect 14186 -1127 14219 -1081
rect 14980 -934 15056 -922
rect 14980 -986 14992 -934
rect 15044 -986 15056 -934
rect 14980 -1038 15056 -986
rect 14980 -1090 14992 -1038
rect 15044 -1090 15056 -1038
rect 14980 -1102 15056 -1090
rect 15620 -934 15696 -922
rect 15620 -986 15632 -934
rect 15684 -986 15696 -934
rect 15620 -1038 15696 -986
rect 15620 -1090 15632 -1038
rect 15684 -1090 15696 -1038
rect 15620 -1102 15696 -1090
rect 16457 -939 16490 -893
rect 16536 -939 16569 -893
rect 16457 -987 16569 -939
rect 16457 -1033 16490 -987
rect 16536 -1033 16569 -987
rect 16457 -1081 16569 -1033
rect 14107 -1175 14219 -1127
rect 14107 -1221 14140 -1175
rect 14186 -1221 14219 -1175
rect 14107 -1269 14219 -1221
rect 14107 -1315 14140 -1269
rect 14186 -1315 14219 -1269
rect 16457 -1127 16490 -1081
rect 16536 -1127 16569 -1081
rect 16457 -1175 16569 -1127
rect 16457 -1221 16490 -1175
rect 16536 -1221 16569 -1175
rect 16457 -1269 16569 -1221
rect 11381 -1409 11414 -1363
rect 11460 -1409 11493 -1363
rect 11381 -1457 11493 -1409
rect 11381 -1503 11414 -1457
rect 11460 -1503 11493 -1457
rect 11866 -1334 11942 -1322
rect 11866 -1386 11878 -1334
rect 11930 -1386 11942 -1334
rect 11866 -1438 11942 -1386
rect 11866 -1490 11878 -1438
rect 11930 -1490 11942 -1438
rect 11381 -1551 11493 -1503
rect 11381 -1597 11414 -1551
rect 11460 -1597 11493 -1551
rect 11381 -1645 11493 -1597
rect 11381 -1691 11414 -1645
rect 11460 -1691 11493 -1645
rect 11381 -1739 11493 -1691
rect 11381 -1785 11414 -1739
rect 11460 -1776 11493 -1739
rect 11593 -1776 11639 -1501
rect 11753 -1776 11799 -1501
rect 11866 -1502 11942 -1490
rect 12762 -1334 12838 -1322
rect 12762 -1386 12774 -1334
rect 12826 -1386 12838 -1334
rect 12762 -1438 12838 -1386
rect 12762 -1490 12774 -1438
rect 12826 -1490 12838 -1438
rect 12169 -1581 12215 -1501
rect 12329 -1512 12375 -1501
rect 12489 -1581 12535 -1501
rect 12617 -1512 12663 -1501
rect 12762 -1502 12838 -1490
rect 13658 -1334 13734 -1322
rect 13658 -1386 13670 -1334
rect 13722 -1386 13734 -1334
rect 13658 -1438 13734 -1386
rect 13658 -1490 13670 -1438
rect 13722 -1490 13734 -1438
rect 12777 -1512 12823 -1502
rect 12937 -1512 12983 -1501
rect 13065 -1581 13111 -1501
rect 13225 -1512 13271 -1501
rect 13385 -1581 13431 -1501
rect 13658 -1502 13734 -1490
rect 14107 -1363 14219 -1315
rect 14107 -1409 14140 -1363
rect 14186 -1409 14219 -1363
rect 14107 -1457 14219 -1409
rect 12169 -1627 13431 -1581
rect 13801 -1776 13847 -1501
rect 13961 -1776 14007 -1501
rect 14107 -1503 14140 -1457
rect 14186 -1503 14219 -1457
rect 14660 -1324 14736 -1312
rect 14660 -1376 14672 -1324
rect 14724 -1376 14736 -1324
rect 14660 -1428 14736 -1376
rect 14660 -1480 14672 -1428
rect 14724 -1480 14736 -1428
rect 14660 -1492 14736 -1480
rect 15300 -1324 15376 -1312
rect 15300 -1376 15312 -1324
rect 15364 -1376 15376 -1324
rect 15300 -1428 15376 -1376
rect 15300 -1480 15312 -1428
rect 15364 -1480 15376 -1428
rect 15300 -1492 15376 -1480
rect 15940 -1324 16016 -1312
rect 15940 -1376 15952 -1324
rect 16004 -1376 16016 -1324
rect 15940 -1428 16016 -1376
rect 15940 -1480 15952 -1428
rect 16004 -1480 16016 -1428
rect 15940 -1492 16016 -1480
rect 16457 -1315 16490 -1269
rect 16536 -1315 16569 -1269
rect 16457 -1363 16569 -1315
rect 16457 -1409 16490 -1363
rect 16536 -1409 16569 -1363
rect 16457 -1457 16569 -1409
rect 14107 -1551 14219 -1503
rect 14107 -1597 14140 -1551
rect 14186 -1597 14219 -1551
rect 14107 -1645 14219 -1597
rect 14107 -1691 14140 -1645
rect 14186 -1691 14219 -1645
rect 14107 -1739 14219 -1691
rect 14107 -1776 14140 -1739
rect 11460 -1785 14140 -1776
rect 14186 -1776 14219 -1739
rect 14835 -1776 14881 -1501
rect 15155 -1776 15201 -1501
rect 15475 -1776 15521 -1501
rect 15795 -1776 15841 -1501
rect 16083 -1776 16129 -1501
rect 16243 -1776 16289 -1501
rect 16457 -1503 16490 -1457
rect 16536 -1503 16569 -1457
rect 16457 -1551 16569 -1503
rect 16457 -1597 16490 -1551
rect 16536 -1597 16569 -1551
rect 16457 -1616 16569 -1597
rect 17569 1603 17889 1651
rect 17569 1557 17650 1603
rect 17696 1557 17889 1603
rect 17569 1509 17889 1557
rect 17569 1463 17650 1509
rect 17696 1463 17889 1509
rect 17569 1415 17889 1463
rect 17569 1369 17650 1415
rect 17696 1369 17889 1415
rect 17569 1321 17889 1369
rect 17569 1275 17650 1321
rect 17696 1275 17889 1321
rect 17569 1227 17889 1275
rect 17569 1181 17650 1227
rect 17696 1181 17889 1227
rect 17569 1133 17889 1181
rect 17569 1087 17650 1133
rect 17696 1087 17889 1133
rect 17569 1039 17889 1087
rect 17569 993 17650 1039
rect 17696 993 17889 1039
rect 17569 945 17889 993
rect 17569 899 17650 945
rect 17696 899 17889 945
rect 17569 851 17889 899
rect 17569 805 17650 851
rect 17696 805 17889 851
rect 17569 757 17889 805
rect 17569 711 17650 757
rect 17696 711 17889 757
rect 17569 663 17889 711
rect 17569 617 17650 663
rect 17696 617 17889 663
rect 17569 569 17889 617
rect 17569 523 17650 569
rect 17696 523 17889 569
rect 17569 475 17889 523
rect 17569 429 17650 475
rect 17696 429 17889 475
rect 17569 381 17889 429
rect 17569 335 17650 381
rect 17696 335 17889 381
rect 17569 287 17889 335
rect 17569 241 17650 287
rect 17696 241 17889 287
rect 17569 193 17889 241
rect 17569 147 17650 193
rect 17696 147 17889 193
rect 17569 99 17889 147
rect 17569 53 17650 99
rect 17696 53 17889 99
rect 17569 5 17889 53
rect 17569 -41 17650 5
rect 17696 -41 17889 5
rect 17569 -89 17889 -41
rect 17569 -135 17650 -89
rect 17696 -135 17889 -89
rect 17569 -183 17889 -135
rect 17569 -229 17650 -183
rect 17696 -229 17889 -183
rect 17569 -277 17889 -229
rect 17569 -323 17650 -277
rect 17696 -323 17889 -277
rect 17569 -371 17889 -323
rect 17569 -417 17650 -371
rect 17696 -417 17889 -371
rect 17569 -465 17889 -417
rect 17569 -511 17650 -465
rect 17696 -511 17889 -465
rect 17569 -559 17889 -511
rect 17569 -605 17650 -559
rect 17696 -605 17889 -559
rect 17569 -653 17889 -605
rect 17569 -699 17650 -653
rect 17696 -699 17889 -653
rect 18226 3287 18272 3445
rect 18386 3287 18432 3445
rect 18674 3386 18720 3445
rect 18834 3434 18880 3445
rect 18994 3386 19040 3445
rect 18674 3340 19040 3386
rect 18226 3241 18306 3287
rect 18352 3241 18432 3287
rect 18226 -457 18272 3241
rect 18386 -457 18432 3241
rect 18579 3282 18655 3294
rect 18579 3230 18591 3282
rect 18643 3279 18655 3282
rect 19922 3287 19968 3445
rect 20082 3287 20128 3445
rect 18643 3233 18754 3279
rect 18800 3233 19074 3279
rect 19120 3233 19394 3279
rect 19440 3233 19714 3279
rect 19760 3233 19771 3279
rect 19922 3241 20002 3287
rect 20048 3241 20128 3287
rect 18643 3230 18655 3233
rect 18579 3218 18655 3230
rect 18819 3071 18895 3083
rect 18819 3019 18831 3071
rect 18883 3019 18895 3071
rect 18819 2967 18895 3019
rect 18819 2915 18831 2967
rect 18883 2915 18895 2967
rect 18819 2903 18895 2915
rect 19459 3071 19535 3083
rect 19459 3019 19471 3071
rect 19523 3019 19535 3071
rect 19459 2967 19535 3019
rect 19459 2915 19471 2967
rect 19523 2915 19535 2967
rect 19459 2903 19535 2915
rect 18499 2677 18575 2689
rect 18499 2625 18511 2677
rect 18563 2625 18575 2677
rect 18499 2573 18575 2625
rect 18499 2521 18511 2573
rect 18563 2521 18575 2573
rect 18499 2509 18575 2521
rect 18659 2677 18735 2689
rect 18659 2625 18671 2677
rect 18723 2625 18735 2677
rect 18659 2573 18735 2625
rect 18659 2521 18671 2573
rect 18723 2521 18735 2573
rect 18659 2509 18735 2521
rect 18979 2677 19055 2689
rect 18979 2625 18991 2677
rect 19043 2625 19055 2677
rect 18979 2573 19055 2625
rect 18979 2521 18991 2573
rect 19043 2521 19055 2573
rect 18979 2509 19055 2521
rect 19139 2677 19215 2689
rect 19139 2625 19151 2677
rect 19203 2625 19215 2677
rect 19139 2573 19215 2625
rect 19139 2521 19151 2573
rect 19203 2521 19215 2573
rect 19139 2509 19215 2521
rect 19299 2677 19375 2689
rect 19299 2625 19311 2677
rect 19363 2625 19375 2677
rect 19299 2573 19375 2625
rect 19299 2521 19311 2573
rect 19363 2521 19375 2573
rect 19299 2509 19375 2521
rect 19619 2677 19695 2689
rect 19619 2625 19631 2677
rect 19683 2625 19695 2677
rect 19619 2573 19695 2625
rect 19619 2521 19631 2573
rect 19683 2521 19695 2573
rect 19619 2509 19695 2521
rect 19779 2677 19855 2689
rect 19779 2625 19791 2677
rect 19843 2625 19855 2677
rect 19779 2573 19855 2625
rect 19779 2521 19791 2573
rect 19843 2521 19855 2573
rect 19779 2509 19855 2521
rect 18674 2450 18720 2509
rect 18834 2498 18880 2509
rect 18994 2450 19040 2509
rect 18674 2404 19040 2450
rect 18579 2346 18655 2358
rect 18579 2294 18591 2346
rect 18643 2343 18655 2346
rect 18643 2297 18754 2343
rect 18800 2297 19074 2343
rect 19120 2297 19394 2343
rect 19440 2297 19714 2343
rect 19760 2297 19771 2343
rect 18643 2294 18655 2297
rect 18579 2282 18655 2294
rect 18819 2135 18895 2147
rect 18819 2083 18831 2135
rect 18883 2083 18895 2135
rect 18819 2031 18895 2083
rect 18819 1979 18831 2031
rect 18883 1979 18895 2031
rect 18819 1967 18895 1979
rect 19459 2135 19535 2147
rect 19459 2083 19471 2135
rect 19523 2083 19535 2135
rect 19459 2031 19535 2083
rect 19459 1979 19471 2031
rect 19523 1979 19535 2031
rect 19459 1967 19535 1979
rect 18499 1741 18575 1753
rect 18499 1689 18511 1741
rect 18563 1689 18575 1741
rect 18499 1637 18575 1689
rect 18499 1585 18511 1637
rect 18563 1585 18575 1637
rect 18499 1573 18575 1585
rect 18659 1741 18735 1753
rect 18659 1689 18671 1741
rect 18723 1689 18735 1741
rect 18659 1637 18735 1689
rect 18659 1585 18671 1637
rect 18723 1585 18735 1637
rect 18659 1573 18735 1585
rect 18979 1741 19055 1753
rect 18979 1689 18991 1741
rect 19043 1689 19055 1741
rect 18979 1637 19055 1689
rect 18979 1585 18991 1637
rect 19043 1585 19055 1637
rect 18979 1573 19055 1585
rect 19139 1741 19215 1753
rect 19139 1689 19151 1741
rect 19203 1689 19215 1741
rect 19139 1637 19215 1689
rect 19139 1585 19151 1637
rect 19203 1585 19215 1637
rect 19139 1573 19215 1585
rect 19299 1741 19375 1753
rect 19299 1689 19311 1741
rect 19363 1689 19375 1741
rect 19299 1637 19375 1689
rect 19299 1585 19311 1637
rect 19363 1585 19375 1637
rect 19299 1573 19375 1585
rect 19619 1741 19695 1753
rect 19619 1689 19631 1741
rect 19683 1689 19695 1741
rect 19619 1637 19695 1689
rect 19619 1585 19631 1637
rect 19683 1585 19695 1637
rect 19619 1573 19695 1585
rect 19779 1741 19855 1753
rect 19779 1689 19791 1741
rect 19843 1689 19855 1741
rect 19779 1637 19855 1689
rect 19779 1585 19791 1637
rect 19843 1585 19855 1637
rect 19779 1573 19855 1585
rect 18514 1211 18560 1573
rect 18674 1211 18720 1573
rect 18834 1211 18880 1573
rect 18994 1211 19040 1573
rect 19154 1211 19200 1573
rect 19314 1211 19360 1573
rect 19474 1211 19520 1573
rect 19634 1211 19680 1573
rect 19794 1211 19840 1573
rect 18819 1199 18895 1211
rect 18819 1147 18831 1199
rect 18883 1147 18895 1199
rect 18819 1095 18895 1147
rect 18819 1043 18831 1095
rect 18883 1043 18895 1095
rect 18819 1031 18895 1043
rect 19459 1199 19535 1211
rect 19459 1147 19471 1199
rect 19523 1147 19535 1199
rect 19459 1095 19535 1147
rect 19459 1043 19471 1095
rect 19523 1043 19535 1095
rect 19459 1031 19535 1043
rect 18499 805 18575 817
rect 18499 753 18511 805
rect 18563 753 18575 805
rect 18499 701 18575 753
rect 18499 649 18511 701
rect 18563 649 18575 701
rect 18499 637 18575 649
rect 19139 805 19215 817
rect 19139 753 19151 805
rect 19203 753 19215 805
rect 19139 701 19215 753
rect 19139 649 19151 701
rect 19203 649 19215 701
rect 19139 637 19215 649
rect 19779 805 19855 817
rect 19779 753 19791 805
rect 19843 753 19855 805
rect 19779 701 19855 753
rect 19779 649 19791 701
rect 19843 649 19855 701
rect 19779 637 19855 649
rect 18674 578 18720 637
rect 18834 626 18880 637
rect 18994 578 19040 637
rect 18674 532 19040 578
rect 18579 474 18655 486
rect 18579 422 18591 474
rect 18643 471 18655 474
rect 18643 425 18754 471
rect 18800 425 19074 471
rect 19120 425 19394 471
rect 19440 425 19714 471
rect 19760 425 19771 471
rect 18643 422 18655 425
rect 18579 410 18655 422
rect 18819 263 18895 275
rect 18819 211 18831 263
rect 18883 211 18895 263
rect 18819 159 18895 211
rect 18819 107 18831 159
rect 18883 107 18895 159
rect 18819 95 18895 107
rect 19459 263 19535 275
rect 19459 211 19471 263
rect 19523 211 19535 263
rect 19459 159 19535 211
rect 19459 107 19471 159
rect 19523 107 19535 159
rect 19459 95 19535 107
rect 18499 -131 18575 -119
rect 18499 -183 18511 -131
rect 18563 -183 18575 -131
rect 18499 -235 18575 -183
rect 18499 -287 18511 -235
rect 18563 -287 18575 -235
rect 18499 -299 18575 -287
rect 18659 -131 18735 -119
rect 18659 -183 18671 -131
rect 18723 -183 18735 -131
rect 18659 -235 18735 -183
rect 18659 -287 18671 -235
rect 18723 -287 18735 -235
rect 18659 -299 18735 -287
rect 18979 -131 19055 -119
rect 18979 -183 18991 -131
rect 19043 -183 19055 -131
rect 18979 -235 19055 -183
rect 18979 -287 18991 -235
rect 19043 -287 19055 -235
rect 18979 -299 19055 -287
rect 19139 -131 19215 -119
rect 19139 -183 19151 -131
rect 19203 -183 19215 -131
rect 19139 -235 19215 -183
rect 19139 -287 19151 -235
rect 19203 -287 19215 -235
rect 19139 -299 19215 -287
rect 19299 -131 19375 -119
rect 19299 -183 19311 -131
rect 19363 -183 19375 -131
rect 19299 -235 19375 -183
rect 19299 -287 19311 -235
rect 19363 -287 19375 -235
rect 19299 -299 19375 -287
rect 19619 -131 19695 -119
rect 19619 -183 19631 -131
rect 19683 -183 19695 -131
rect 19619 -235 19695 -183
rect 19619 -287 19631 -235
rect 19683 -287 19695 -235
rect 19619 -299 19695 -287
rect 19779 -131 19855 -119
rect 19779 -183 19791 -131
rect 19843 -183 19855 -131
rect 19779 -235 19855 -183
rect 19779 -287 19791 -235
rect 19843 -287 19855 -235
rect 19779 -299 19855 -287
rect 18674 -358 18720 -299
rect 18834 -310 18880 -299
rect 18994 -358 19040 -299
rect 18674 -404 19040 -358
rect 18226 -503 18306 -457
rect 18352 -503 18432 -457
rect 18226 -661 18272 -503
rect 18386 -661 18432 -503
rect 18579 -462 18655 -450
rect 18579 -514 18591 -462
rect 18643 -465 18655 -462
rect 19922 -457 19968 3241
rect 20082 -457 20128 3241
rect 18643 -511 18754 -465
rect 18800 -511 19074 -465
rect 19120 -511 19394 -465
rect 19440 -511 19714 -465
rect 19760 -511 19771 -465
rect 19922 -503 20002 -457
rect 20048 -503 20128 -457
rect 18643 -514 18655 -511
rect 18579 -526 18655 -514
rect 19922 -661 19968 -503
rect 20082 -661 20128 -503
rect 20465 3437 20658 3483
rect 20704 3437 20785 3483
rect 20465 3389 20785 3437
rect 20465 3343 20658 3389
rect 20704 3343 20785 3389
rect 20465 3295 20785 3343
rect 20465 3249 20658 3295
rect 20704 3249 20785 3295
rect 20465 3201 20785 3249
rect 20465 3155 20658 3201
rect 20704 3155 20785 3201
rect 20465 3107 20785 3155
rect 20465 3061 20658 3107
rect 20704 3061 20785 3107
rect 20465 3013 20785 3061
rect 20465 2967 20658 3013
rect 20704 2967 20785 3013
rect 20465 2919 20785 2967
rect 20465 2873 20658 2919
rect 20704 2873 20785 2919
rect 20465 2825 20785 2873
rect 20465 2779 20658 2825
rect 20704 2779 20785 2825
rect 20465 2731 20785 2779
rect 20465 2685 20658 2731
rect 20704 2685 20785 2731
rect 20465 2637 20785 2685
rect 20465 2591 20658 2637
rect 20704 2591 20785 2637
rect 20465 2543 20785 2591
rect 20465 2497 20658 2543
rect 20704 2497 20785 2543
rect 20465 2449 20785 2497
rect 20465 2403 20658 2449
rect 20704 2403 20785 2449
rect 20465 2355 20785 2403
rect 20465 2309 20658 2355
rect 20704 2309 20785 2355
rect 20465 2261 20785 2309
rect 20465 2215 20658 2261
rect 20704 2215 20785 2261
rect 20465 2167 20785 2215
rect 20465 2121 20658 2167
rect 20704 2121 20785 2167
rect 20465 2073 20785 2121
rect 20465 2027 20658 2073
rect 20704 2027 20785 2073
rect 20465 1979 20785 2027
rect 20465 1933 20658 1979
rect 20704 1933 20785 1979
rect 20465 1885 20785 1933
rect 20465 1839 20658 1885
rect 20704 1839 20785 1885
rect 20465 1791 20785 1839
rect 20465 1745 20658 1791
rect 20704 1745 20785 1791
rect 20465 1697 20785 1745
rect 20465 1651 20658 1697
rect 20704 1651 20785 1697
rect 20465 1603 20785 1651
rect 20465 1557 20658 1603
rect 20704 1557 20785 1603
rect 20465 1509 20785 1557
rect 20465 1463 20658 1509
rect 20704 1463 20785 1509
rect 20465 1415 20785 1463
rect 20465 1369 20658 1415
rect 20704 1369 20785 1415
rect 20465 1321 20785 1369
rect 20465 1275 20658 1321
rect 20704 1275 20785 1321
rect 20465 1227 20785 1275
rect 20465 1181 20658 1227
rect 20704 1181 20785 1227
rect 20465 1133 20785 1181
rect 20465 1087 20658 1133
rect 20704 1087 20785 1133
rect 20465 1039 20785 1087
rect 20465 993 20658 1039
rect 20704 993 20785 1039
rect 20465 945 20785 993
rect 20465 899 20658 945
rect 20704 899 20785 945
rect 20465 851 20785 899
rect 20465 805 20658 851
rect 20704 805 20785 851
rect 20465 757 20785 805
rect 20465 711 20658 757
rect 20704 711 20785 757
rect 20465 663 20785 711
rect 20465 617 20658 663
rect 20704 617 20785 663
rect 20465 569 20785 617
rect 20465 523 20658 569
rect 20704 523 20785 569
rect 20465 475 20785 523
rect 20465 429 20658 475
rect 20704 429 20785 475
rect 20465 381 20785 429
rect 20465 335 20658 381
rect 20704 335 20785 381
rect 20465 287 20785 335
rect 20465 241 20658 287
rect 20704 241 20785 287
rect 20465 193 20785 241
rect 20465 147 20658 193
rect 20704 147 20785 193
rect 20465 99 20785 147
rect 20465 53 20658 99
rect 20704 53 20785 99
rect 20465 5 20785 53
rect 20465 -41 20658 5
rect 20704 -41 20785 5
rect 20465 -89 20785 -41
rect 20465 -135 20658 -89
rect 20704 -135 20785 -89
rect 20465 -183 20785 -135
rect 20465 -229 20658 -183
rect 20704 -229 20785 -183
rect 20465 -277 20785 -229
rect 20465 -323 20658 -277
rect 20704 -323 20785 -277
rect 20465 -371 20785 -323
rect 20465 -417 20658 -371
rect 20704 -417 20785 -371
rect 20465 -465 20785 -417
rect 20465 -511 20658 -465
rect 20704 -511 20785 -465
rect 20465 -559 20785 -511
rect 20465 -605 20658 -559
rect 20704 -605 20785 -559
rect 20465 -653 20785 -605
rect 17569 -747 17889 -699
rect 17569 -793 17650 -747
rect 17696 -793 17889 -747
rect 17569 -841 17889 -793
rect 18819 -673 18895 -661
rect 18819 -725 18831 -673
rect 18883 -725 18895 -673
rect 18819 -777 18895 -725
rect 18819 -829 18831 -777
rect 18883 -829 18895 -777
rect 18819 -841 18895 -829
rect 19459 -673 19535 -661
rect 19459 -725 19471 -673
rect 19523 -725 19535 -673
rect 19459 -777 19535 -725
rect 19459 -829 19471 -777
rect 19523 -829 19535 -777
rect 19459 -841 19535 -829
rect 20465 -699 20658 -653
rect 20704 -699 20785 -653
rect 20465 -747 20785 -699
rect 20465 -793 20658 -747
rect 20704 -793 20785 -747
rect 20465 -841 20785 -793
rect 17569 -887 17650 -841
rect 17696 -887 17889 -841
rect 17569 -935 17889 -887
rect 17569 -981 17650 -935
rect 17696 -981 17889 -935
rect 17569 -1029 17889 -981
rect 17569 -1075 17650 -1029
rect 17696 -1075 17889 -1029
rect 20465 -887 20658 -841
rect 20704 -887 20785 -841
rect 20465 -935 20785 -887
rect 20465 -981 20658 -935
rect 20704 -981 20785 -935
rect 20465 -1029 20785 -981
rect 17569 -1123 17889 -1075
rect 17569 -1169 17650 -1123
rect 17696 -1169 17889 -1123
rect 17569 -1217 17889 -1169
rect 17569 -1263 17650 -1217
rect 17696 -1263 17889 -1217
rect 18499 -1067 18575 -1055
rect 18499 -1119 18511 -1067
rect 18563 -1119 18575 -1067
rect 18499 -1171 18575 -1119
rect 18499 -1223 18511 -1171
rect 18563 -1223 18575 -1171
rect 18499 -1235 18575 -1223
rect 18659 -1067 18735 -1055
rect 18659 -1119 18671 -1067
rect 18723 -1119 18735 -1067
rect 18659 -1171 18735 -1119
rect 18659 -1223 18671 -1171
rect 18723 -1223 18735 -1171
rect 18659 -1235 18735 -1223
rect 18979 -1067 19055 -1055
rect 18979 -1119 18991 -1067
rect 19043 -1119 19055 -1067
rect 18979 -1171 19055 -1119
rect 18979 -1223 18991 -1171
rect 19043 -1223 19055 -1171
rect 18979 -1235 19055 -1223
rect 19139 -1067 19215 -1055
rect 19139 -1119 19151 -1067
rect 19203 -1119 19215 -1067
rect 19139 -1171 19215 -1119
rect 19139 -1223 19151 -1171
rect 19203 -1223 19215 -1171
rect 19139 -1235 19215 -1223
rect 19299 -1067 19375 -1055
rect 19299 -1119 19311 -1067
rect 19363 -1119 19375 -1067
rect 19299 -1171 19375 -1119
rect 19299 -1223 19311 -1171
rect 19363 -1223 19375 -1171
rect 19299 -1235 19375 -1223
rect 19619 -1067 19695 -1055
rect 19619 -1119 19631 -1067
rect 19683 -1119 19695 -1067
rect 19619 -1171 19695 -1119
rect 19619 -1223 19631 -1171
rect 19683 -1223 19695 -1171
rect 19619 -1235 19695 -1223
rect 19779 -1067 19855 -1055
rect 19779 -1119 19791 -1067
rect 19843 -1119 19855 -1067
rect 19779 -1171 19855 -1119
rect 19779 -1223 19791 -1171
rect 19843 -1223 19855 -1171
rect 19779 -1235 19855 -1223
rect 20465 -1075 20658 -1029
rect 20704 -1075 20785 -1029
rect 20465 -1123 20785 -1075
rect 20465 -1169 20658 -1123
rect 20704 -1169 20785 -1123
rect 20465 -1217 20785 -1169
rect 17569 -1311 17889 -1263
rect 17569 -1357 17650 -1311
rect 17696 -1357 17889 -1311
rect 17569 -1405 17889 -1357
rect 17569 -1451 17650 -1405
rect 17696 -1451 17889 -1405
rect 17569 -1499 17889 -1451
rect 17569 -1545 17650 -1499
rect 17696 -1545 17889 -1499
rect 17569 -1593 17889 -1545
rect 16457 -1645 16573 -1616
rect 16457 -1691 16490 -1645
rect 16536 -1691 16573 -1645
rect 16457 -1739 16573 -1691
rect 16457 -1776 16490 -1739
rect 14186 -1785 16490 -1776
rect 16536 -1785 16573 -1739
rect 11381 -1833 16573 -1785
rect 11381 -1879 11414 -1833
rect 11460 -1879 11508 -1833
rect 11554 -1879 11602 -1833
rect 11648 -1879 11696 -1833
rect 11742 -1879 11790 -1833
rect 11836 -1879 11884 -1833
rect 11930 -1879 11978 -1833
rect 12024 -1879 12072 -1833
rect 12118 -1879 12166 -1833
rect 12212 -1879 12260 -1833
rect 12306 -1879 12354 -1833
rect 12400 -1879 12448 -1833
rect 12494 -1879 12542 -1833
rect 12588 -1879 12636 -1833
rect 12682 -1879 12730 -1833
rect 12776 -1879 12824 -1833
rect 12870 -1879 12918 -1833
rect 12964 -1879 13012 -1833
rect 13058 -1879 13106 -1833
rect 13152 -1879 13200 -1833
rect 13246 -1879 13294 -1833
rect 13340 -1879 13388 -1833
rect 13434 -1879 13482 -1833
rect 13528 -1879 13576 -1833
rect 13622 -1879 13670 -1833
rect 13716 -1879 13764 -1833
rect 13810 -1879 13858 -1833
rect 13904 -1879 13952 -1833
rect 13998 -1879 14046 -1833
rect 14092 -1879 14140 -1833
rect 14186 -1879 14234 -1833
rect 14280 -1879 14328 -1833
rect 14374 -1879 14422 -1833
rect 14468 -1879 14516 -1833
rect 14562 -1879 14610 -1833
rect 14656 -1879 14704 -1833
rect 14750 -1879 14798 -1833
rect 14844 -1879 14892 -1833
rect 14938 -1879 14986 -1833
rect 15032 -1879 15080 -1833
rect 15126 -1879 15174 -1833
rect 15220 -1879 15268 -1833
rect 15314 -1879 15362 -1833
rect 15408 -1879 15456 -1833
rect 15502 -1879 15550 -1833
rect 15596 -1879 15644 -1833
rect 15690 -1879 15738 -1833
rect 15784 -1879 15832 -1833
rect 15878 -1879 15926 -1833
rect 15972 -1879 16020 -1833
rect 16066 -1879 16114 -1833
rect 16160 -1879 16208 -1833
rect 16254 -1879 16302 -1833
rect 16348 -1879 16396 -1833
rect 16442 -1879 16490 -1833
rect 16536 -1879 16573 -1833
rect 11381 -1936 16573 -1879
rect 17569 -1639 17650 -1593
rect 17696 -1616 17889 -1593
rect 18226 -1616 18272 -1235
rect 18386 -1616 18432 -1235
rect 18674 -1294 18720 -1235
rect 18994 -1294 19040 -1235
rect 19314 -1294 19360 -1235
rect 19634 -1294 19680 -1235
rect 18674 -1340 19680 -1294
rect 18739 -1398 18815 -1386
rect 18739 -1450 18751 -1398
rect 18803 -1401 18815 -1398
rect 19379 -1398 19455 -1386
rect 19379 -1401 19391 -1398
rect 18803 -1447 19391 -1401
rect 18803 -1450 18815 -1447
rect 18739 -1462 18815 -1450
rect 19379 -1450 19391 -1447
rect 19443 -1450 19455 -1398
rect 19379 -1462 19455 -1450
rect 19634 -1616 19680 -1340
rect 19922 -1616 19968 -1235
rect 20082 -1616 20128 -1235
rect 20465 -1263 20658 -1217
rect 20704 -1263 20785 -1217
rect 20465 -1311 20785 -1263
rect 20465 -1357 20658 -1311
rect 20704 -1357 20785 -1311
rect 20465 -1405 20785 -1357
rect 20465 -1451 20658 -1405
rect 20704 -1451 20785 -1405
rect 20465 -1499 20785 -1451
rect 20465 -1545 20658 -1499
rect 20704 -1545 20785 -1499
rect 20465 -1593 20785 -1545
rect 20465 -1616 20658 -1593
rect 17696 -1639 20658 -1616
rect 20704 -1616 20785 -1593
rect 22721 4377 22802 4400
rect 22848 4400 25810 4423
rect 22848 4377 23041 4400
rect 22721 4329 23041 4377
rect 22721 4283 22802 4329
rect 22848 4283 23041 4329
rect 22721 4235 23041 4283
rect 22721 4189 22802 4235
rect 22848 4189 23041 4235
rect 22721 4141 23041 4189
rect 22721 4095 22802 4141
rect 22848 4095 23041 4141
rect 22721 4047 23041 4095
rect 22721 4001 22802 4047
rect 22848 4001 23041 4047
rect 23378 4019 23424 4400
rect 23538 4019 23584 4400
rect 23731 4248 23807 4260
rect 23731 4196 23743 4248
rect 23795 4245 23807 4248
rect 24851 4248 24927 4260
rect 24851 4245 24863 4248
rect 23795 4199 24386 4245
rect 24432 4199 24863 4245
rect 23795 4196 23807 4199
rect 23731 4184 23807 4196
rect 24851 4196 24863 4199
rect 24915 4196 24927 4248
rect 24851 4184 24927 4196
rect 25074 4019 25120 4400
rect 25234 4019 25280 4400
rect 25617 4377 25810 4400
rect 25856 4400 26771 4423
rect 25856 4377 25937 4400
rect 25617 4329 25937 4377
rect 25617 4283 25810 4329
rect 25856 4283 25937 4329
rect 25617 4235 25937 4283
rect 25617 4189 25810 4235
rect 25856 4189 25937 4235
rect 25617 4141 25937 4189
rect 25617 4095 25810 4141
rect 25856 4095 25937 4141
rect 25617 4047 25937 4095
rect 22721 3953 23041 4001
rect 22721 3907 22802 3953
rect 22848 3907 23041 3953
rect 22721 3859 23041 3907
rect 22721 3813 22802 3859
rect 22848 3813 23041 3859
rect 23971 4007 24047 4019
rect 23971 3955 23983 4007
rect 24035 3955 24047 4007
rect 23971 3903 24047 3955
rect 23971 3851 23983 3903
rect 24035 3851 24047 3903
rect 23971 3839 24047 3851
rect 24611 4007 24687 4019
rect 24611 3955 24623 4007
rect 24675 3955 24687 4007
rect 24611 3903 24687 3955
rect 24611 3851 24623 3903
rect 24675 3851 24687 3903
rect 24611 3839 24687 3851
rect 25617 4001 25810 4047
rect 25856 4001 25937 4047
rect 25617 3953 25937 4001
rect 25617 3907 25810 3953
rect 25856 3907 25937 3953
rect 25617 3859 25937 3907
rect 22721 3765 23041 3813
rect 22721 3719 22802 3765
rect 22848 3719 23041 3765
rect 22721 3671 23041 3719
rect 22721 3625 22802 3671
rect 22848 3625 23041 3671
rect 25617 3813 25810 3859
rect 25856 3813 25937 3859
rect 25617 3765 25937 3813
rect 25617 3719 25810 3765
rect 25856 3719 25937 3765
rect 25617 3671 25937 3719
rect 25617 3625 25810 3671
rect 25856 3625 25937 3671
rect 22721 3577 23041 3625
rect 22721 3531 22802 3577
rect 22848 3531 23041 3577
rect 22721 3483 23041 3531
rect 22721 3437 22802 3483
rect 22848 3437 23041 3483
rect 23651 3613 23727 3625
rect 23651 3561 23663 3613
rect 23715 3561 23727 3613
rect 23651 3509 23727 3561
rect 23651 3457 23663 3509
rect 23715 3457 23727 3509
rect 23651 3445 23727 3457
rect 23811 3613 23887 3625
rect 23811 3561 23823 3613
rect 23875 3561 23887 3613
rect 23811 3509 23887 3561
rect 23811 3457 23823 3509
rect 23875 3457 23887 3509
rect 23811 3445 23887 3457
rect 24131 3613 24207 3625
rect 24131 3561 24143 3613
rect 24195 3561 24207 3613
rect 24131 3509 24207 3561
rect 24131 3457 24143 3509
rect 24195 3457 24207 3509
rect 24131 3445 24207 3457
rect 24291 3613 24367 3625
rect 24291 3561 24303 3613
rect 24355 3561 24367 3613
rect 24291 3509 24367 3561
rect 24291 3457 24303 3509
rect 24355 3457 24367 3509
rect 24291 3445 24367 3457
rect 24451 3613 24527 3625
rect 24451 3561 24463 3613
rect 24515 3561 24527 3613
rect 24451 3509 24527 3561
rect 24451 3457 24463 3509
rect 24515 3457 24527 3509
rect 24451 3445 24527 3457
rect 24771 3613 24847 3625
rect 24771 3561 24783 3613
rect 24835 3561 24847 3613
rect 24771 3509 24847 3561
rect 24771 3457 24783 3509
rect 24835 3457 24847 3509
rect 24771 3445 24847 3457
rect 24931 3613 25007 3625
rect 24931 3561 24943 3613
rect 24995 3561 25007 3613
rect 24931 3509 25007 3561
rect 24931 3457 24943 3509
rect 24995 3457 25007 3509
rect 24931 3445 25007 3457
rect 25617 3577 25937 3625
rect 25617 3531 25810 3577
rect 25856 3531 25937 3577
rect 25617 3483 25937 3531
rect 22721 3389 23041 3437
rect 22721 3343 22802 3389
rect 22848 3343 23041 3389
rect 22721 3295 23041 3343
rect 22721 3249 22802 3295
rect 22848 3249 23041 3295
rect 22721 3201 23041 3249
rect 22721 3155 22802 3201
rect 22848 3155 23041 3201
rect 22721 3107 23041 3155
rect 22721 3061 22802 3107
rect 22848 3061 23041 3107
rect 22721 3013 23041 3061
rect 22721 2967 22802 3013
rect 22848 2967 23041 3013
rect 22721 2919 23041 2967
rect 22721 2873 22802 2919
rect 22848 2873 23041 2919
rect 22721 2825 23041 2873
rect 22721 2779 22802 2825
rect 22848 2779 23041 2825
rect 22721 2731 23041 2779
rect 22721 2685 22802 2731
rect 22848 2685 23041 2731
rect 22721 2637 23041 2685
rect 22721 2591 22802 2637
rect 22848 2591 23041 2637
rect 22721 2543 23041 2591
rect 22721 2497 22802 2543
rect 22848 2497 23041 2543
rect 22721 2449 23041 2497
rect 22721 2403 22802 2449
rect 22848 2403 23041 2449
rect 22721 2355 23041 2403
rect 22721 2309 22802 2355
rect 22848 2309 23041 2355
rect 22721 2261 23041 2309
rect 22721 2215 22802 2261
rect 22848 2215 23041 2261
rect 22721 2167 23041 2215
rect 22721 2121 22802 2167
rect 22848 2121 23041 2167
rect 22721 2073 23041 2121
rect 22721 2027 22802 2073
rect 22848 2027 23041 2073
rect 22721 1979 23041 2027
rect 22721 1933 22802 1979
rect 22848 1933 23041 1979
rect 22721 1885 23041 1933
rect 22721 1839 22802 1885
rect 22848 1839 23041 1885
rect 22721 1791 23041 1839
rect 22721 1745 22802 1791
rect 22848 1745 23041 1791
rect 22721 1697 23041 1745
rect 22721 1651 22802 1697
rect 22848 1651 23041 1697
rect 22721 1603 23041 1651
rect 22721 1557 22802 1603
rect 22848 1557 23041 1603
rect 22721 1509 23041 1557
rect 22721 1463 22802 1509
rect 22848 1463 23041 1509
rect 22721 1415 23041 1463
rect 22721 1369 22802 1415
rect 22848 1369 23041 1415
rect 22721 1321 23041 1369
rect 22721 1275 22802 1321
rect 22848 1275 23041 1321
rect 22721 1227 23041 1275
rect 22721 1181 22802 1227
rect 22848 1181 23041 1227
rect 22721 1133 23041 1181
rect 22721 1087 22802 1133
rect 22848 1087 23041 1133
rect 22721 1039 23041 1087
rect 22721 993 22802 1039
rect 22848 993 23041 1039
rect 22721 945 23041 993
rect 22721 899 22802 945
rect 22848 899 23041 945
rect 22721 851 23041 899
rect 22721 805 22802 851
rect 22848 805 23041 851
rect 22721 757 23041 805
rect 22721 711 22802 757
rect 22848 711 23041 757
rect 22721 663 23041 711
rect 22721 617 22802 663
rect 22848 617 23041 663
rect 22721 569 23041 617
rect 22721 523 22802 569
rect 22848 523 23041 569
rect 22721 475 23041 523
rect 22721 429 22802 475
rect 22848 429 23041 475
rect 22721 381 23041 429
rect 22721 335 22802 381
rect 22848 335 23041 381
rect 22721 287 23041 335
rect 22721 241 22802 287
rect 22848 241 23041 287
rect 22721 193 23041 241
rect 22721 147 22802 193
rect 22848 147 23041 193
rect 22721 99 23041 147
rect 22721 53 22802 99
rect 22848 53 23041 99
rect 22721 5 23041 53
rect 22721 -41 22802 5
rect 22848 -41 23041 5
rect 22721 -89 23041 -41
rect 22721 -135 22802 -89
rect 22848 -135 23041 -89
rect 22721 -183 23041 -135
rect 22721 -229 22802 -183
rect 22848 -229 23041 -183
rect 22721 -277 23041 -229
rect 22721 -323 22802 -277
rect 22848 -323 23041 -277
rect 22721 -371 23041 -323
rect 22721 -417 22802 -371
rect 22848 -417 23041 -371
rect 22721 -465 23041 -417
rect 22721 -511 22802 -465
rect 22848 -511 23041 -465
rect 22721 -559 23041 -511
rect 22721 -605 22802 -559
rect 22848 -605 23041 -559
rect 22721 -653 23041 -605
rect 22721 -699 22802 -653
rect 22848 -699 23041 -653
rect 23378 3287 23424 3445
rect 23538 3287 23584 3445
rect 24466 3386 24512 3445
rect 24626 3434 24672 3445
rect 24786 3386 24832 3445
rect 24466 3340 24832 3386
rect 23378 3241 23458 3287
rect 23504 3241 23584 3287
rect 24851 3282 24927 3294
rect 24851 3279 24863 3282
rect 23378 -457 23424 3241
rect 23538 -457 23584 3241
rect 23735 3233 23746 3279
rect 23792 3233 24066 3279
rect 24112 3233 24386 3279
rect 24432 3233 24706 3279
rect 24752 3233 24863 3279
rect 24851 3230 24863 3233
rect 24915 3230 24927 3282
rect 24851 3218 24927 3230
rect 25074 3287 25120 3445
rect 25234 3287 25280 3445
rect 25074 3241 25154 3287
rect 25200 3241 25280 3287
rect 23971 3071 24047 3083
rect 23971 3019 23983 3071
rect 24035 3019 24047 3071
rect 23971 2967 24047 3019
rect 23971 2915 23983 2967
rect 24035 2915 24047 2967
rect 23971 2903 24047 2915
rect 24611 3071 24687 3083
rect 24611 3019 24623 3071
rect 24675 3019 24687 3071
rect 24611 2967 24687 3019
rect 24611 2915 24623 2967
rect 24675 2915 24687 2967
rect 24611 2903 24687 2915
rect 23651 2677 23727 2689
rect 23651 2625 23663 2677
rect 23715 2625 23727 2677
rect 23651 2573 23727 2625
rect 23651 2521 23663 2573
rect 23715 2521 23727 2573
rect 23651 2509 23727 2521
rect 23811 2677 23887 2689
rect 23811 2625 23823 2677
rect 23875 2625 23887 2677
rect 23811 2573 23887 2625
rect 23811 2521 23823 2573
rect 23875 2521 23887 2573
rect 23811 2509 23887 2521
rect 24131 2677 24207 2689
rect 24131 2625 24143 2677
rect 24195 2625 24207 2677
rect 24131 2573 24207 2625
rect 24131 2521 24143 2573
rect 24195 2521 24207 2573
rect 24131 2509 24207 2521
rect 24291 2677 24367 2689
rect 24291 2625 24303 2677
rect 24355 2625 24367 2677
rect 24291 2573 24367 2625
rect 24291 2521 24303 2573
rect 24355 2521 24367 2573
rect 24291 2509 24367 2521
rect 24451 2677 24527 2689
rect 24451 2625 24463 2677
rect 24515 2625 24527 2677
rect 24451 2573 24527 2625
rect 24451 2521 24463 2573
rect 24515 2521 24527 2573
rect 24451 2509 24527 2521
rect 24771 2677 24847 2689
rect 24771 2625 24783 2677
rect 24835 2625 24847 2677
rect 24771 2573 24847 2625
rect 24771 2521 24783 2573
rect 24835 2521 24847 2573
rect 24771 2509 24847 2521
rect 24931 2677 25007 2689
rect 24931 2625 24943 2677
rect 24995 2625 25007 2677
rect 24931 2573 25007 2625
rect 24931 2521 24943 2573
rect 24995 2521 25007 2573
rect 24931 2509 25007 2521
rect 24466 2450 24512 2509
rect 24626 2498 24672 2509
rect 24786 2450 24832 2509
rect 24466 2404 24832 2450
rect 24851 2346 24927 2358
rect 24851 2343 24863 2346
rect 23735 2297 23746 2343
rect 23792 2297 24066 2343
rect 24112 2297 24386 2343
rect 24432 2297 24706 2343
rect 24752 2297 24863 2343
rect 24851 2294 24863 2297
rect 24915 2294 24927 2346
rect 24851 2282 24927 2294
rect 23971 2135 24047 2147
rect 23971 2083 23983 2135
rect 24035 2083 24047 2135
rect 23971 2031 24047 2083
rect 23971 1979 23983 2031
rect 24035 1979 24047 2031
rect 23971 1967 24047 1979
rect 24611 2135 24687 2147
rect 24611 2083 24623 2135
rect 24675 2083 24687 2135
rect 24611 2031 24687 2083
rect 24611 1979 24623 2031
rect 24675 1979 24687 2031
rect 24611 1967 24687 1979
rect 23651 1741 23727 1753
rect 23651 1689 23663 1741
rect 23715 1689 23727 1741
rect 23651 1637 23727 1689
rect 23651 1585 23663 1637
rect 23715 1585 23727 1637
rect 23651 1573 23727 1585
rect 23811 1741 23887 1753
rect 23811 1689 23823 1741
rect 23875 1689 23887 1741
rect 23811 1637 23887 1689
rect 23811 1585 23823 1637
rect 23875 1585 23887 1637
rect 23811 1573 23887 1585
rect 24131 1741 24207 1753
rect 24131 1689 24143 1741
rect 24195 1689 24207 1741
rect 24131 1637 24207 1689
rect 24131 1585 24143 1637
rect 24195 1585 24207 1637
rect 24131 1573 24207 1585
rect 24291 1741 24367 1753
rect 24291 1689 24303 1741
rect 24355 1689 24367 1741
rect 24291 1637 24367 1689
rect 24291 1585 24303 1637
rect 24355 1585 24367 1637
rect 24291 1573 24367 1585
rect 24451 1741 24527 1753
rect 24451 1689 24463 1741
rect 24515 1689 24527 1741
rect 24451 1637 24527 1689
rect 24451 1585 24463 1637
rect 24515 1585 24527 1637
rect 24451 1573 24527 1585
rect 24771 1741 24847 1753
rect 24771 1689 24783 1741
rect 24835 1689 24847 1741
rect 24771 1637 24847 1689
rect 24771 1585 24783 1637
rect 24835 1585 24847 1637
rect 24771 1573 24847 1585
rect 24931 1741 25007 1753
rect 24931 1689 24943 1741
rect 24995 1689 25007 1741
rect 24931 1637 25007 1689
rect 24931 1585 24943 1637
rect 24995 1585 25007 1637
rect 24931 1573 25007 1585
rect 23666 1211 23712 1573
rect 23826 1211 23872 1573
rect 23986 1211 24032 1573
rect 24146 1211 24192 1573
rect 24306 1211 24352 1573
rect 24466 1211 24512 1573
rect 24626 1211 24672 1573
rect 24786 1211 24832 1573
rect 24946 1211 24992 1573
rect 23971 1199 24047 1211
rect 23971 1147 23983 1199
rect 24035 1147 24047 1199
rect 23971 1095 24047 1147
rect 23971 1043 23983 1095
rect 24035 1043 24047 1095
rect 23971 1031 24047 1043
rect 24611 1199 24687 1211
rect 24611 1147 24623 1199
rect 24675 1147 24687 1199
rect 24611 1095 24687 1147
rect 24611 1043 24623 1095
rect 24675 1043 24687 1095
rect 24611 1031 24687 1043
rect 23651 805 23727 817
rect 23651 753 23663 805
rect 23715 753 23727 805
rect 23651 701 23727 753
rect 23651 649 23663 701
rect 23715 649 23727 701
rect 23651 637 23727 649
rect 24291 805 24367 817
rect 24291 753 24303 805
rect 24355 753 24367 805
rect 24291 701 24367 753
rect 24291 649 24303 701
rect 24355 649 24367 701
rect 24291 637 24367 649
rect 24931 805 25007 817
rect 24931 753 24943 805
rect 24995 753 25007 805
rect 24931 701 25007 753
rect 24931 649 24943 701
rect 24995 649 25007 701
rect 24931 637 25007 649
rect 24466 578 24512 637
rect 24626 626 24672 637
rect 24786 578 24832 637
rect 24466 532 24832 578
rect 24851 474 24927 486
rect 24851 471 24863 474
rect 23735 425 23746 471
rect 23792 425 24066 471
rect 24112 425 24386 471
rect 24432 425 24706 471
rect 24752 425 24863 471
rect 24851 422 24863 425
rect 24915 422 24927 474
rect 24851 410 24927 422
rect 23971 263 24047 275
rect 23971 211 23983 263
rect 24035 211 24047 263
rect 23971 159 24047 211
rect 23971 107 23983 159
rect 24035 107 24047 159
rect 23971 95 24047 107
rect 24611 263 24687 275
rect 24611 211 24623 263
rect 24675 211 24687 263
rect 24611 159 24687 211
rect 24611 107 24623 159
rect 24675 107 24687 159
rect 24611 95 24687 107
rect 23651 -131 23727 -119
rect 23651 -183 23663 -131
rect 23715 -183 23727 -131
rect 23651 -235 23727 -183
rect 23651 -287 23663 -235
rect 23715 -287 23727 -235
rect 23651 -299 23727 -287
rect 23811 -131 23887 -119
rect 23811 -183 23823 -131
rect 23875 -183 23887 -131
rect 23811 -235 23887 -183
rect 23811 -287 23823 -235
rect 23875 -287 23887 -235
rect 23811 -299 23887 -287
rect 24131 -131 24207 -119
rect 24131 -183 24143 -131
rect 24195 -183 24207 -131
rect 24131 -235 24207 -183
rect 24131 -287 24143 -235
rect 24195 -287 24207 -235
rect 24131 -299 24207 -287
rect 24291 -131 24367 -119
rect 24291 -183 24303 -131
rect 24355 -183 24367 -131
rect 24291 -235 24367 -183
rect 24291 -287 24303 -235
rect 24355 -287 24367 -235
rect 24291 -299 24367 -287
rect 24451 -131 24527 -119
rect 24451 -183 24463 -131
rect 24515 -183 24527 -131
rect 24451 -235 24527 -183
rect 24451 -287 24463 -235
rect 24515 -287 24527 -235
rect 24451 -299 24527 -287
rect 24771 -131 24847 -119
rect 24771 -183 24783 -131
rect 24835 -183 24847 -131
rect 24771 -235 24847 -183
rect 24771 -287 24783 -235
rect 24835 -287 24847 -235
rect 24771 -299 24847 -287
rect 24931 -131 25007 -119
rect 24931 -183 24943 -131
rect 24995 -183 25007 -131
rect 24931 -235 25007 -183
rect 24931 -287 24943 -235
rect 24995 -287 25007 -235
rect 24931 -299 25007 -287
rect 24466 -358 24512 -299
rect 24626 -310 24672 -299
rect 24786 -358 24832 -299
rect 24466 -404 24832 -358
rect 23378 -503 23458 -457
rect 23504 -503 23584 -457
rect 24851 -462 24927 -450
rect 24851 -465 24863 -462
rect 23378 -661 23424 -503
rect 23538 -661 23584 -503
rect 23735 -511 23746 -465
rect 23792 -511 24066 -465
rect 24112 -511 24386 -465
rect 24432 -511 24706 -465
rect 24752 -511 24863 -465
rect 24851 -514 24863 -511
rect 24915 -514 24927 -462
rect 24851 -526 24927 -514
rect 25074 -457 25120 3241
rect 25234 -457 25280 3241
rect 25074 -503 25154 -457
rect 25200 -503 25280 -457
rect 25074 -661 25120 -503
rect 25234 -661 25280 -503
rect 25617 3437 25810 3483
rect 25856 3437 25937 3483
rect 25617 3389 25937 3437
rect 25617 3343 25810 3389
rect 25856 3343 25937 3389
rect 25617 3295 25937 3343
rect 25617 3249 25810 3295
rect 25856 3249 25937 3295
rect 25617 3201 25937 3249
rect 25617 3155 25810 3201
rect 25856 3155 25937 3201
rect 25617 3107 25937 3155
rect 25617 3061 25810 3107
rect 25856 3061 25937 3107
rect 25617 3013 25937 3061
rect 25617 2967 25810 3013
rect 25856 2967 25937 3013
rect 25617 2919 25937 2967
rect 25617 2873 25810 2919
rect 25856 2873 25937 2919
rect 25617 2825 25937 2873
rect 25617 2779 25810 2825
rect 25856 2779 25937 2825
rect 25617 2731 25937 2779
rect 25617 2685 25810 2731
rect 25856 2685 25937 2731
rect 25617 2637 25937 2685
rect 25617 2591 25810 2637
rect 25856 2591 25937 2637
rect 25617 2543 25937 2591
rect 25617 2497 25810 2543
rect 25856 2497 25937 2543
rect 25617 2449 25937 2497
rect 25617 2403 25810 2449
rect 25856 2403 25937 2449
rect 25617 2355 25937 2403
rect 25617 2309 25810 2355
rect 25856 2309 25937 2355
rect 25617 2261 25937 2309
rect 25617 2215 25810 2261
rect 25856 2215 25937 2261
rect 25617 2167 25937 2215
rect 25617 2121 25810 2167
rect 25856 2121 25937 2167
rect 25617 2073 25937 2121
rect 25617 2027 25810 2073
rect 25856 2027 25937 2073
rect 25617 1979 25937 2027
rect 25617 1933 25810 1979
rect 25856 1933 25937 1979
rect 25617 1885 25937 1933
rect 25617 1839 25810 1885
rect 25856 1839 25937 1885
rect 25617 1791 25937 1839
rect 25617 1745 25810 1791
rect 25856 1745 25937 1791
rect 25617 1697 25937 1745
rect 25617 1651 25810 1697
rect 25856 1651 25937 1697
rect 25617 1603 25937 1651
rect 25617 1557 25810 1603
rect 25856 1557 25937 1603
rect 25617 1509 25937 1557
rect 25617 1463 25810 1509
rect 25856 1463 25937 1509
rect 25617 1415 25937 1463
rect 25617 1369 25810 1415
rect 25856 1369 25937 1415
rect 25617 1321 25937 1369
rect 25617 1275 25810 1321
rect 25856 1275 25937 1321
rect 25617 1227 25937 1275
rect 25617 1181 25810 1227
rect 25856 1181 25937 1227
rect 25617 1133 25937 1181
rect 25617 1087 25810 1133
rect 25856 1087 25937 1133
rect 25617 1039 25937 1087
rect 25617 993 25810 1039
rect 25856 993 25937 1039
rect 25617 945 25937 993
rect 25617 899 25810 945
rect 25856 899 25937 945
rect 25617 851 25937 899
rect 25617 805 25810 851
rect 25856 805 25937 851
rect 25617 757 25937 805
rect 25617 711 25810 757
rect 25856 711 25937 757
rect 25617 663 25937 711
rect 25617 617 25810 663
rect 25856 617 25937 663
rect 25617 569 25937 617
rect 25617 523 25810 569
rect 25856 523 25937 569
rect 25617 475 25937 523
rect 25617 429 25810 475
rect 25856 429 25937 475
rect 25617 381 25937 429
rect 25617 335 25810 381
rect 25856 335 25937 381
rect 25617 287 25937 335
rect 25617 241 25810 287
rect 25856 241 25937 287
rect 25617 193 25937 241
rect 25617 147 25810 193
rect 25856 147 25937 193
rect 25617 99 25937 147
rect 25617 53 25810 99
rect 25856 53 25937 99
rect 25617 5 25937 53
rect 25617 -41 25810 5
rect 25856 -41 25937 5
rect 25617 -89 25937 -41
rect 25617 -135 25810 -89
rect 25856 -135 25937 -89
rect 25617 -183 25937 -135
rect 25617 -229 25810 -183
rect 25856 -229 25937 -183
rect 25617 -277 25937 -229
rect 25617 -323 25810 -277
rect 25856 -323 25937 -277
rect 25617 -371 25937 -323
rect 25617 -417 25810 -371
rect 25856 -417 25937 -371
rect 25617 -465 25937 -417
rect 25617 -511 25810 -465
rect 25856 -511 25937 -465
rect 25617 -559 25937 -511
rect 25617 -605 25810 -559
rect 25856 -605 25937 -559
rect 25617 -653 25937 -605
rect 22721 -747 23041 -699
rect 22721 -793 22802 -747
rect 22848 -793 23041 -747
rect 22721 -841 23041 -793
rect 23971 -673 24047 -661
rect 23971 -725 23983 -673
rect 24035 -725 24047 -673
rect 23971 -777 24047 -725
rect 23971 -829 23983 -777
rect 24035 -829 24047 -777
rect 23971 -841 24047 -829
rect 24611 -673 24687 -661
rect 24611 -725 24623 -673
rect 24675 -725 24687 -673
rect 24611 -777 24687 -725
rect 24611 -829 24623 -777
rect 24675 -829 24687 -777
rect 24611 -841 24687 -829
rect 25617 -699 25810 -653
rect 25856 -699 25937 -653
rect 25617 -747 25937 -699
rect 25617 -793 25810 -747
rect 25856 -793 25937 -747
rect 25617 -841 25937 -793
rect 22721 -887 22802 -841
rect 22848 -887 23041 -841
rect 22721 -935 23041 -887
rect 22721 -981 22802 -935
rect 22848 -981 23041 -935
rect 22721 -1029 23041 -981
rect 22721 -1075 22802 -1029
rect 22848 -1075 23041 -1029
rect 25617 -887 25810 -841
rect 25856 -887 25937 -841
rect 25617 -935 25937 -887
rect 25617 -981 25810 -935
rect 25856 -981 25937 -935
rect 25617 -1029 25937 -981
rect 22721 -1123 23041 -1075
rect 22721 -1169 22802 -1123
rect 22848 -1169 23041 -1123
rect 22721 -1217 23041 -1169
rect 22721 -1263 22802 -1217
rect 22848 -1263 23041 -1217
rect 23651 -1067 23727 -1055
rect 23651 -1119 23663 -1067
rect 23715 -1119 23727 -1067
rect 23651 -1171 23727 -1119
rect 23651 -1223 23663 -1171
rect 23715 -1223 23727 -1171
rect 23651 -1235 23727 -1223
rect 23811 -1067 23887 -1055
rect 23811 -1119 23823 -1067
rect 23875 -1119 23887 -1067
rect 23811 -1171 23887 -1119
rect 23811 -1223 23823 -1171
rect 23875 -1223 23887 -1171
rect 23811 -1235 23887 -1223
rect 24131 -1067 24207 -1055
rect 24131 -1119 24143 -1067
rect 24195 -1119 24207 -1067
rect 24131 -1171 24207 -1119
rect 24131 -1223 24143 -1171
rect 24195 -1223 24207 -1171
rect 24131 -1235 24207 -1223
rect 24291 -1067 24367 -1055
rect 24291 -1119 24303 -1067
rect 24355 -1119 24367 -1067
rect 24291 -1171 24367 -1119
rect 24291 -1223 24303 -1171
rect 24355 -1223 24367 -1171
rect 24291 -1235 24367 -1223
rect 24451 -1067 24527 -1055
rect 24451 -1119 24463 -1067
rect 24515 -1119 24527 -1067
rect 24451 -1171 24527 -1119
rect 24451 -1223 24463 -1171
rect 24515 -1223 24527 -1171
rect 24451 -1235 24527 -1223
rect 24771 -1067 24847 -1055
rect 24771 -1119 24783 -1067
rect 24835 -1119 24847 -1067
rect 24771 -1171 24847 -1119
rect 24771 -1223 24783 -1171
rect 24835 -1223 24847 -1171
rect 24771 -1235 24847 -1223
rect 24931 -1067 25007 -1055
rect 24931 -1119 24943 -1067
rect 24995 -1119 25007 -1067
rect 24931 -1171 25007 -1119
rect 24931 -1223 24943 -1171
rect 24995 -1223 25007 -1171
rect 24931 -1235 25007 -1223
rect 25617 -1075 25810 -1029
rect 25856 -1075 25937 -1029
rect 25617 -1123 25937 -1075
rect 25617 -1169 25810 -1123
rect 25856 -1169 25937 -1123
rect 25617 -1217 25937 -1169
rect 22721 -1311 23041 -1263
rect 22721 -1357 22802 -1311
rect 22848 -1357 23041 -1311
rect 22721 -1405 23041 -1357
rect 22721 -1451 22802 -1405
rect 22848 -1451 23041 -1405
rect 22721 -1499 23041 -1451
rect 22721 -1545 22802 -1499
rect 22848 -1545 23041 -1499
rect 22721 -1593 23041 -1545
rect 22721 -1616 22802 -1593
rect 20704 -1639 22802 -1616
rect 22848 -1616 23041 -1593
rect 23378 -1616 23424 -1235
rect 23538 -1616 23584 -1235
rect 23826 -1294 23872 -1235
rect 24146 -1294 24192 -1235
rect 24466 -1294 24512 -1235
rect 24786 -1294 24832 -1235
rect 23826 -1340 24832 -1294
rect 23826 -1616 23872 -1340
rect 24051 -1398 24127 -1386
rect 24051 -1450 24063 -1398
rect 24115 -1401 24127 -1398
rect 24691 -1398 24767 -1386
rect 24691 -1401 24703 -1398
rect 24115 -1447 24703 -1401
rect 24115 -1450 24127 -1447
rect 24051 -1462 24127 -1450
rect 24691 -1450 24703 -1447
rect 24755 -1450 24767 -1398
rect 24691 -1462 24767 -1450
rect 25074 -1616 25120 -1235
rect 25234 -1616 25280 -1235
rect 25617 -1263 25810 -1217
rect 25856 -1263 25937 -1217
rect 25617 -1311 25937 -1263
rect 25617 -1357 25810 -1311
rect 25856 -1357 25937 -1311
rect 25617 -1405 25937 -1357
rect 25617 -1451 25810 -1405
rect 25856 -1451 25937 -1405
rect 25617 -1499 25937 -1451
rect 25617 -1545 25810 -1499
rect 25856 -1545 25937 -1499
rect 25617 -1593 25937 -1545
rect 25617 -1616 25810 -1593
rect 22848 -1639 25810 -1616
rect 25856 -1616 25937 -1593
rect 26690 4377 26771 4400
rect 26817 4400 29779 4423
rect 26817 4377 27010 4400
rect 26690 4329 27010 4377
rect 26690 4283 26771 4329
rect 26817 4283 27010 4329
rect 26690 4235 27010 4283
rect 26690 4189 26771 4235
rect 26817 4189 27010 4235
rect 26690 4141 27010 4189
rect 26690 4095 26771 4141
rect 26817 4095 27010 4141
rect 26690 4047 27010 4095
rect 26690 4001 26771 4047
rect 26817 4001 27010 4047
rect 27347 4019 27393 4400
rect 27507 4019 27553 4400
rect 27700 4248 27776 4260
rect 27700 4196 27712 4248
rect 27764 4245 27776 4248
rect 27764 4199 28195 4245
rect 28241 4199 28835 4245
rect 28881 4199 28892 4245
rect 27764 4196 27776 4199
rect 27700 4184 27776 4196
rect 29043 4019 29089 4400
rect 29203 4019 29249 4400
rect 29586 4377 29779 4400
rect 29825 4377 29906 4423
rect 29586 4329 29906 4377
rect 29586 4283 29779 4329
rect 29825 4283 29906 4329
rect 29586 4235 29906 4283
rect 29586 4189 29779 4235
rect 29825 4189 29906 4235
rect 29586 4141 29906 4189
rect 29586 4095 29779 4141
rect 29825 4095 29906 4141
rect 29586 4047 29906 4095
rect 26690 3953 27010 4001
rect 26690 3907 26771 3953
rect 26817 3907 27010 3953
rect 26690 3859 27010 3907
rect 26690 3813 26771 3859
rect 26817 3813 27010 3859
rect 27940 4007 28016 4019
rect 27940 3955 27952 4007
rect 28004 3955 28016 4007
rect 27940 3903 28016 3955
rect 27940 3851 27952 3903
rect 28004 3851 28016 3903
rect 27940 3839 28016 3851
rect 28580 4007 28656 4019
rect 28580 3955 28592 4007
rect 28644 3955 28656 4007
rect 28580 3903 28656 3955
rect 28580 3851 28592 3903
rect 28644 3851 28656 3903
rect 28580 3839 28656 3851
rect 29586 4001 29779 4047
rect 29825 4001 29906 4047
rect 29586 3953 29906 4001
rect 29586 3907 29779 3953
rect 29825 3907 29906 3953
rect 29586 3859 29906 3907
rect 26690 3765 27010 3813
rect 26690 3719 26771 3765
rect 26817 3719 27010 3765
rect 26690 3671 27010 3719
rect 26690 3625 26771 3671
rect 26817 3625 27010 3671
rect 29586 3813 29779 3859
rect 29825 3813 29906 3859
rect 29586 3765 29906 3813
rect 29586 3719 29779 3765
rect 29825 3719 29906 3765
rect 29586 3671 29906 3719
rect 29586 3625 29779 3671
rect 29825 3625 29906 3671
rect 26690 3577 27010 3625
rect 26690 3531 26771 3577
rect 26817 3531 27010 3577
rect 26690 3483 27010 3531
rect 26690 3437 26771 3483
rect 26817 3437 27010 3483
rect 27620 3613 27696 3625
rect 27620 3561 27632 3613
rect 27684 3561 27696 3613
rect 27620 3509 27696 3561
rect 27620 3457 27632 3509
rect 27684 3457 27696 3509
rect 27620 3445 27696 3457
rect 27780 3613 27856 3625
rect 27780 3561 27792 3613
rect 27844 3561 27856 3613
rect 27780 3509 27856 3561
rect 27780 3457 27792 3509
rect 27844 3457 27856 3509
rect 27780 3445 27856 3457
rect 28100 3613 28176 3625
rect 28100 3561 28112 3613
rect 28164 3561 28176 3613
rect 28100 3509 28176 3561
rect 28100 3457 28112 3509
rect 28164 3457 28176 3509
rect 28100 3445 28176 3457
rect 28260 3613 28336 3625
rect 28260 3561 28272 3613
rect 28324 3561 28336 3613
rect 28260 3509 28336 3561
rect 28260 3457 28272 3509
rect 28324 3457 28336 3509
rect 28260 3445 28336 3457
rect 28420 3613 28496 3625
rect 28420 3561 28432 3613
rect 28484 3561 28496 3613
rect 28420 3509 28496 3561
rect 28420 3457 28432 3509
rect 28484 3457 28496 3509
rect 28420 3445 28496 3457
rect 28740 3613 28816 3625
rect 28740 3561 28752 3613
rect 28804 3561 28816 3613
rect 28740 3509 28816 3561
rect 28740 3457 28752 3509
rect 28804 3457 28816 3509
rect 28740 3445 28816 3457
rect 28900 3613 28976 3625
rect 28900 3561 28912 3613
rect 28964 3561 28976 3613
rect 28900 3509 28976 3561
rect 28900 3457 28912 3509
rect 28964 3457 28976 3509
rect 28900 3445 28976 3457
rect 29586 3577 29906 3625
rect 29586 3531 29779 3577
rect 29825 3531 29906 3577
rect 29586 3483 29906 3531
rect 26690 3389 27010 3437
rect 26690 3343 26771 3389
rect 26817 3343 27010 3389
rect 26690 3295 27010 3343
rect 26690 3249 26771 3295
rect 26817 3249 27010 3295
rect 26690 3201 27010 3249
rect 26690 3155 26771 3201
rect 26817 3155 27010 3201
rect 26690 3107 27010 3155
rect 26690 3061 26771 3107
rect 26817 3061 27010 3107
rect 26690 3013 27010 3061
rect 26690 2967 26771 3013
rect 26817 2967 27010 3013
rect 26690 2919 27010 2967
rect 26690 2873 26771 2919
rect 26817 2873 27010 2919
rect 26690 2825 27010 2873
rect 26690 2779 26771 2825
rect 26817 2779 27010 2825
rect 26690 2731 27010 2779
rect 26690 2685 26771 2731
rect 26817 2685 27010 2731
rect 26690 2637 27010 2685
rect 26690 2591 26771 2637
rect 26817 2591 27010 2637
rect 26690 2543 27010 2591
rect 26690 2497 26771 2543
rect 26817 2497 27010 2543
rect 26690 2449 27010 2497
rect 26690 2403 26771 2449
rect 26817 2403 27010 2449
rect 26690 2355 27010 2403
rect 26690 2309 26771 2355
rect 26817 2309 27010 2355
rect 26690 2261 27010 2309
rect 26690 2215 26771 2261
rect 26817 2215 27010 2261
rect 26690 2167 27010 2215
rect 26690 2121 26771 2167
rect 26817 2121 27010 2167
rect 26690 2073 27010 2121
rect 26690 2027 26771 2073
rect 26817 2027 27010 2073
rect 26690 1979 27010 2027
rect 26690 1933 26771 1979
rect 26817 1933 27010 1979
rect 26690 1885 27010 1933
rect 26690 1839 26771 1885
rect 26817 1839 27010 1885
rect 26690 1791 27010 1839
rect 26690 1745 26771 1791
rect 26817 1745 27010 1791
rect 26690 1697 27010 1745
rect 26690 1651 26771 1697
rect 26817 1651 27010 1697
rect 26690 1603 27010 1651
rect 26690 1557 26771 1603
rect 26817 1557 27010 1603
rect 26690 1509 27010 1557
rect 26690 1463 26771 1509
rect 26817 1463 27010 1509
rect 26690 1415 27010 1463
rect 26690 1369 26771 1415
rect 26817 1369 27010 1415
rect 26690 1321 27010 1369
rect 26690 1275 26771 1321
rect 26817 1275 27010 1321
rect 26690 1227 27010 1275
rect 26690 1181 26771 1227
rect 26817 1181 27010 1227
rect 26690 1133 27010 1181
rect 26690 1087 26771 1133
rect 26817 1087 27010 1133
rect 26690 1039 27010 1087
rect 26690 993 26771 1039
rect 26817 993 27010 1039
rect 26690 945 27010 993
rect 26690 899 26771 945
rect 26817 899 27010 945
rect 26690 851 27010 899
rect 26690 805 26771 851
rect 26817 805 27010 851
rect 26690 757 27010 805
rect 26690 711 26771 757
rect 26817 711 27010 757
rect 26690 663 27010 711
rect 26690 617 26771 663
rect 26817 617 27010 663
rect 26690 569 27010 617
rect 26690 523 26771 569
rect 26817 523 27010 569
rect 26690 475 27010 523
rect 26690 429 26771 475
rect 26817 429 27010 475
rect 26690 381 27010 429
rect 26690 335 26771 381
rect 26817 335 27010 381
rect 26690 287 27010 335
rect 26690 241 26771 287
rect 26817 241 27010 287
rect 26690 193 27010 241
rect 26690 147 26771 193
rect 26817 147 27010 193
rect 26690 99 27010 147
rect 26690 53 26771 99
rect 26817 53 27010 99
rect 26690 5 27010 53
rect 26690 -41 26771 5
rect 26817 -41 27010 5
rect 26690 -89 27010 -41
rect 26690 -135 26771 -89
rect 26817 -135 27010 -89
rect 26690 -183 27010 -135
rect 26690 -229 26771 -183
rect 26817 -229 27010 -183
rect 26690 -277 27010 -229
rect 26690 -323 26771 -277
rect 26817 -323 27010 -277
rect 26690 -371 27010 -323
rect 26690 -417 26771 -371
rect 26817 -417 27010 -371
rect 26690 -465 27010 -417
rect 26690 -511 26771 -465
rect 26817 -511 27010 -465
rect 26690 -559 27010 -511
rect 26690 -605 26771 -559
rect 26817 -605 27010 -559
rect 26690 -653 27010 -605
rect 26690 -699 26771 -653
rect 26817 -699 27010 -653
rect 27347 3287 27393 3445
rect 27507 3287 27553 3445
rect 27795 3386 27841 3445
rect 27955 3434 28001 3445
rect 28115 3386 28161 3445
rect 27795 3340 28161 3386
rect 27347 3241 27427 3287
rect 27473 3241 27553 3287
rect 27347 -457 27393 3241
rect 27507 -457 27553 3241
rect 27700 3282 27776 3294
rect 27700 3230 27712 3282
rect 27764 3279 27776 3282
rect 29043 3287 29089 3445
rect 29203 3287 29249 3445
rect 27764 3233 27875 3279
rect 27921 3233 28195 3279
rect 28241 3233 28515 3279
rect 28561 3233 28835 3279
rect 28881 3233 28892 3279
rect 29043 3241 29123 3287
rect 29169 3241 29249 3287
rect 27764 3230 27776 3233
rect 27700 3218 27776 3230
rect 27940 3071 28016 3083
rect 27940 3019 27952 3071
rect 28004 3019 28016 3071
rect 27940 2967 28016 3019
rect 27940 2915 27952 2967
rect 28004 2915 28016 2967
rect 27940 2903 28016 2915
rect 28580 3071 28656 3083
rect 28580 3019 28592 3071
rect 28644 3019 28656 3071
rect 28580 2967 28656 3019
rect 28580 2915 28592 2967
rect 28644 2915 28656 2967
rect 28580 2903 28656 2915
rect 27620 2677 27696 2689
rect 27620 2625 27632 2677
rect 27684 2625 27696 2677
rect 27620 2573 27696 2625
rect 27620 2521 27632 2573
rect 27684 2521 27696 2573
rect 27620 2509 27696 2521
rect 27780 2677 27856 2689
rect 27780 2625 27792 2677
rect 27844 2625 27856 2677
rect 27780 2573 27856 2625
rect 27780 2521 27792 2573
rect 27844 2521 27856 2573
rect 27780 2509 27856 2521
rect 28100 2677 28176 2689
rect 28100 2625 28112 2677
rect 28164 2625 28176 2677
rect 28100 2573 28176 2625
rect 28100 2521 28112 2573
rect 28164 2521 28176 2573
rect 28100 2509 28176 2521
rect 28260 2677 28336 2689
rect 28260 2625 28272 2677
rect 28324 2625 28336 2677
rect 28260 2573 28336 2625
rect 28260 2521 28272 2573
rect 28324 2521 28336 2573
rect 28260 2509 28336 2521
rect 28420 2677 28496 2689
rect 28420 2625 28432 2677
rect 28484 2625 28496 2677
rect 28420 2573 28496 2625
rect 28420 2521 28432 2573
rect 28484 2521 28496 2573
rect 28420 2509 28496 2521
rect 28740 2677 28816 2689
rect 28740 2625 28752 2677
rect 28804 2625 28816 2677
rect 28740 2573 28816 2625
rect 28740 2521 28752 2573
rect 28804 2521 28816 2573
rect 28740 2509 28816 2521
rect 28900 2677 28976 2689
rect 28900 2625 28912 2677
rect 28964 2625 28976 2677
rect 28900 2573 28976 2625
rect 28900 2521 28912 2573
rect 28964 2521 28976 2573
rect 28900 2509 28976 2521
rect 27795 2450 27841 2509
rect 27955 2498 28001 2509
rect 28115 2450 28161 2509
rect 27795 2404 28161 2450
rect 27700 2346 27776 2358
rect 27700 2294 27712 2346
rect 27764 2343 27776 2346
rect 27764 2297 27875 2343
rect 27921 2297 28195 2343
rect 28241 2297 28515 2343
rect 28561 2297 28835 2343
rect 28881 2297 28892 2343
rect 27764 2294 27776 2297
rect 27700 2282 27776 2294
rect 27940 2135 28016 2147
rect 27940 2083 27952 2135
rect 28004 2083 28016 2135
rect 27940 2031 28016 2083
rect 27940 1979 27952 2031
rect 28004 1979 28016 2031
rect 27940 1967 28016 1979
rect 28580 2135 28656 2147
rect 28580 2083 28592 2135
rect 28644 2083 28656 2135
rect 28580 2031 28656 2083
rect 28580 1979 28592 2031
rect 28644 1979 28656 2031
rect 28580 1967 28656 1979
rect 27620 1741 27696 1753
rect 27620 1689 27632 1741
rect 27684 1689 27696 1741
rect 27620 1637 27696 1689
rect 27620 1585 27632 1637
rect 27684 1585 27696 1637
rect 27620 1573 27696 1585
rect 27780 1741 27856 1753
rect 27780 1689 27792 1741
rect 27844 1689 27856 1741
rect 27780 1637 27856 1689
rect 27780 1585 27792 1637
rect 27844 1585 27856 1637
rect 27780 1573 27856 1585
rect 28100 1741 28176 1753
rect 28100 1689 28112 1741
rect 28164 1689 28176 1741
rect 28100 1637 28176 1689
rect 28100 1585 28112 1637
rect 28164 1585 28176 1637
rect 28100 1573 28176 1585
rect 28260 1741 28336 1753
rect 28260 1689 28272 1741
rect 28324 1689 28336 1741
rect 28260 1637 28336 1689
rect 28260 1585 28272 1637
rect 28324 1585 28336 1637
rect 28260 1573 28336 1585
rect 28420 1741 28496 1753
rect 28420 1689 28432 1741
rect 28484 1689 28496 1741
rect 28420 1637 28496 1689
rect 28420 1585 28432 1637
rect 28484 1585 28496 1637
rect 28420 1573 28496 1585
rect 28740 1741 28816 1753
rect 28740 1689 28752 1741
rect 28804 1689 28816 1741
rect 28740 1637 28816 1689
rect 28740 1585 28752 1637
rect 28804 1585 28816 1637
rect 28740 1573 28816 1585
rect 28900 1741 28976 1753
rect 28900 1689 28912 1741
rect 28964 1689 28976 1741
rect 28900 1637 28976 1689
rect 28900 1585 28912 1637
rect 28964 1585 28976 1637
rect 28900 1573 28976 1585
rect 27635 1211 27681 1573
rect 27795 1211 27841 1573
rect 27955 1211 28001 1573
rect 28115 1211 28161 1573
rect 28275 1211 28321 1573
rect 28435 1211 28481 1573
rect 28595 1211 28641 1573
rect 28755 1211 28801 1573
rect 28915 1211 28961 1573
rect 27940 1199 28016 1211
rect 27940 1147 27952 1199
rect 28004 1147 28016 1199
rect 27940 1095 28016 1147
rect 27940 1043 27952 1095
rect 28004 1043 28016 1095
rect 27940 1031 28016 1043
rect 28580 1199 28656 1211
rect 28580 1147 28592 1199
rect 28644 1147 28656 1199
rect 28580 1095 28656 1147
rect 28580 1043 28592 1095
rect 28644 1043 28656 1095
rect 28580 1031 28656 1043
rect 27620 805 27696 817
rect 27620 753 27632 805
rect 27684 753 27696 805
rect 27620 701 27696 753
rect 27620 649 27632 701
rect 27684 649 27696 701
rect 27620 637 27696 649
rect 28260 805 28336 817
rect 28260 753 28272 805
rect 28324 753 28336 805
rect 28260 701 28336 753
rect 28260 649 28272 701
rect 28324 649 28336 701
rect 28260 637 28336 649
rect 28900 805 28976 817
rect 28900 753 28912 805
rect 28964 753 28976 805
rect 28900 701 28976 753
rect 28900 649 28912 701
rect 28964 649 28976 701
rect 28900 637 28976 649
rect 27795 578 27841 637
rect 27955 626 28001 637
rect 28115 578 28161 637
rect 27795 532 28161 578
rect 27700 474 27776 486
rect 27700 422 27712 474
rect 27764 471 27776 474
rect 27764 425 27875 471
rect 27921 425 28195 471
rect 28241 425 28515 471
rect 28561 425 28835 471
rect 28881 425 28892 471
rect 27764 422 27776 425
rect 27700 410 27776 422
rect 27940 263 28016 275
rect 27940 211 27952 263
rect 28004 211 28016 263
rect 27940 159 28016 211
rect 27940 107 27952 159
rect 28004 107 28016 159
rect 27940 95 28016 107
rect 28580 263 28656 275
rect 28580 211 28592 263
rect 28644 211 28656 263
rect 28580 159 28656 211
rect 28580 107 28592 159
rect 28644 107 28656 159
rect 28580 95 28656 107
rect 27620 -131 27696 -119
rect 27620 -183 27632 -131
rect 27684 -183 27696 -131
rect 27620 -235 27696 -183
rect 27620 -287 27632 -235
rect 27684 -287 27696 -235
rect 27620 -299 27696 -287
rect 27780 -131 27856 -119
rect 27780 -183 27792 -131
rect 27844 -183 27856 -131
rect 27780 -235 27856 -183
rect 27780 -287 27792 -235
rect 27844 -287 27856 -235
rect 27780 -299 27856 -287
rect 28100 -131 28176 -119
rect 28100 -183 28112 -131
rect 28164 -183 28176 -131
rect 28100 -235 28176 -183
rect 28100 -287 28112 -235
rect 28164 -287 28176 -235
rect 28100 -299 28176 -287
rect 28260 -131 28336 -119
rect 28260 -183 28272 -131
rect 28324 -183 28336 -131
rect 28260 -235 28336 -183
rect 28260 -287 28272 -235
rect 28324 -287 28336 -235
rect 28260 -299 28336 -287
rect 28420 -131 28496 -119
rect 28420 -183 28432 -131
rect 28484 -183 28496 -131
rect 28420 -235 28496 -183
rect 28420 -287 28432 -235
rect 28484 -287 28496 -235
rect 28420 -299 28496 -287
rect 28740 -131 28816 -119
rect 28740 -183 28752 -131
rect 28804 -183 28816 -131
rect 28740 -235 28816 -183
rect 28740 -287 28752 -235
rect 28804 -287 28816 -235
rect 28740 -299 28816 -287
rect 28900 -131 28976 -119
rect 28900 -183 28912 -131
rect 28964 -183 28976 -131
rect 28900 -235 28976 -183
rect 28900 -287 28912 -235
rect 28964 -287 28976 -235
rect 28900 -299 28976 -287
rect 27795 -358 27841 -299
rect 27955 -310 28001 -299
rect 28115 -358 28161 -299
rect 27795 -404 28161 -358
rect 27347 -503 27427 -457
rect 27473 -503 27553 -457
rect 27347 -661 27393 -503
rect 27507 -661 27553 -503
rect 27700 -462 27776 -450
rect 27700 -514 27712 -462
rect 27764 -465 27776 -462
rect 29043 -457 29089 3241
rect 29203 -457 29249 3241
rect 27764 -511 27875 -465
rect 27921 -511 28195 -465
rect 28241 -511 28515 -465
rect 28561 -511 28835 -465
rect 28881 -511 28892 -465
rect 29043 -503 29123 -457
rect 29169 -503 29249 -457
rect 27764 -514 27776 -511
rect 27700 -526 27776 -514
rect 29043 -661 29089 -503
rect 29203 -661 29249 -503
rect 29586 3437 29779 3483
rect 29825 3437 29906 3483
rect 29586 3389 29906 3437
rect 29586 3343 29779 3389
rect 29825 3343 29906 3389
rect 29586 3295 29906 3343
rect 29586 3249 29779 3295
rect 29825 3249 29906 3295
rect 29586 3201 29906 3249
rect 29586 3155 29779 3201
rect 29825 3155 29906 3201
rect 29586 3107 29906 3155
rect 29586 3061 29779 3107
rect 29825 3061 29906 3107
rect 29586 3013 29906 3061
rect 29586 2967 29779 3013
rect 29825 2967 29906 3013
rect 29586 2919 29906 2967
rect 29586 2873 29779 2919
rect 29825 2873 29906 2919
rect 29586 2825 29906 2873
rect 29586 2779 29779 2825
rect 29825 2779 29906 2825
rect 29586 2731 29906 2779
rect 29586 2685 29779 2731
rect 29825 2685 29906 2731
rect 29586 2637 29906 2685
rect 29586 2591 29779 2637
rect 29825 2591 29906 2637
rect 29586 2543 29906 2591
rect 29586 2497 29779 2543
rect 29825 2497 29906 2543
rect 29586 2449 29906 2497
rect 29586 2403 29779 2449
rect 29825 2403 29906 2449
rect 29586 2355 29906 2403
rect 29586 2309 29779 2355
rect 29825 2309 29906 2355
rect 29586 2261 29906 2309
rect 29586 2215 29779 2261
rect 29825 2215 29906 2261
rect 29586 2167 29906 2215
rect 29586 2121 29779 2167
rect 29825 2121 29906 2167
rect 29586 2073 29906 2121
rect 29586 2027 29779 2073
rect 29825 2027 29906 2073
rect 29586 1979 29906 2027
rect 29586 1933 29779 1979
rect 29825 1933 29906 1979
rect 29586 1885 29906 1933
rect 29586 1839 29779 1885
rect 29825 1839 29906 1885
rect 29586 1791 29906 1839
rect 29586 1745 29779 1791
rect 29825 1745 29906 1791
rect 29586 1697 29906 1745
rect 29586 1651 29779 1697
rect 29825 1651 29906 1697
rect 29586 1603 29906 1651
rect 29586 1557 29779 1603
rect 29825 1557 29906 1603
rect 29586 1509 29906 1557
rect 29586 1463 29779 1509
rect 29825 1463 29906 1509
rect 29586 1415 29906 1463
rect 29586 1369 29779 1415
rect 29825 1369 29906 1415
rect 29586 1321 29906 1369
rect 29586 1275 29779 1321
rect 29825 1275 29906 1321
rect 29586 1227 29906 1275
rect 29586 1181 29779 1227
rect 29825 1181 29906 1227
rect 29586 1133 29906 1181
rect 29586 1087 29779 1133
rect 29825 1087 29906 1133
rect 29586 1039 29906 1087
rect 29586 993 29779 1039
rect 29825 993 29906 1039
rect 29586 945 29906 993
rect 29586 899 29779 945
rect 29825 899 29906 945
rect 29586 851 29906 899
rect 29586 805 29779 851
rect 29825 805 29906 851
rect 29586 757 29906 805
rect 29586 711 29779 757
rect 29825 711 29906 757
rect 29586 663 29906 711
rect 29586 617 29779 663
rect 29825 617 29906 663
rect 29586 569 29906 617
rect 29586 523 29779 569
rect 29825 523 29906 569
rect 29586 475 29906 523
rect 29586 429 29779 475
rect 29825 429 29906 475
rect 29586 381 29906 429
rect 29586 335 29779 381
rect 29825 335 29906 381
rect 29586 287 29906 335
rect 29586 241 29779 287
rect 29825 241 29906 287
rect 29586 193 29906 241
rect 29586 147 29779 193
rect 29825 147 29906 193
rect 29586 99 29906 147
rect 29586 53 29779 99
rect 29825 53 29906 99
rect 29586 5 29906 53
rect 29586 -41 29779 5
rect 29825 -41 29906 5
rect 29586 -89 29906 -41
rect 29586 -135 29779 -89
rect 29825 -135 29906 -89
rect 29586 -183 29906 -135
rect 29586 -229 29779 -183
rect 29825 -229 29906 -183
rect 29586 -277 29906 -229
rect 29586 -323 29779 -277
rect 29825 -323 29906 -277
rect 29586 -371 29906 -323
rect 29586 -417 29779 -371
rect 29825 -417 29906 -371
rect 29586 -465 29906 -417
rect 29586 -511 29779 -465
rect 29825 -511 29906 -465
rect 29586 -559 29906 -511
rect 29586 -605 29779 -559
rect 29825 -605 29906 -559
rect 29586 -653 29906 -605
rect 26690 -747 27010 -699
rect 26690 -793 26771 -747
rect 26817 -793 27010 -747
rect 26690 -841 27010 -793
rect 27940 -673 28016 -661
rect 27940 -725 27952 -673
rect 28004 -725 28016 -673
rect 27940 -777 28016 -725
rect 27940 -829 27952 -777
rect 28004 -829 28016 -777
rect 27940 -841 28016 -829
rect 28580 -673 28656 -661
rect 28580 -725 28592 -673
rect 28644 -725 28656 -673
rect 28580 -777 28656 -725
rect 28580 -829 28592 -777
rect 28644 -829 28656 -777
rect 28580 -841 28656 -829
rect 29586 -699 29779 -653
rect 29825 -699 29906 -653
rect 29586 -747 29906 -699
rect 29586 -793 29779 -747
rect 29825 -793 29906 -747
rect 29586 -841 29906 -793
rect 26690 -887 26771 -841
rect 26817 -887 27010 -841
rect 26690 -935 27010 -887
rect 26690 -981 26771 -935
rect 26817 -981 27010 -935
rect 26690 -1029 27010 -981
rect 26690 -1075 26771 -1029
rect 26817 -1075 27010 -1029
rect 29586 -887 29779 -841
rect 29825 -887 29906 -841
rect 29586 -935 29906 -887
rect 29586 -981 29779 -935
rect 29825 -981 29906 -935
rect 29586 -1029 29906 -981
rect 26690 -1123 27010 -1075
rect 26690 -1169 26771 -1123
rect 26817 -1169 27010 -1123
rect 26690 -1217 27010 -1169
rect 26690 -1263 26771 -1217
rect 26817 -1263 27010 -1217
rect 27620 -1067 27696 -1055
rect 27620 -1119 27632 -1067
rect 27684 -1119 27696 -1067
rect 27620 -1171 27696 -1119
rect 27620 -1223 27632 -1171
rect 27684 -1223 27696 -1171
rect 27620 -1235 27696 -1223
rect 27780 -1067 27856 -1055
rect 27780 -1119 27792 -1067
rect 27844 -1119 27856 -1067
rect 27780 -1171 27856 -1119
rect 27780 -1223 27792 -1171
rect 27844 -1223 27856 -1171
rect 27780 -1235 27856 -1223
rect 28100 -1067 28176 -1055
rect 28100 -1119 28112 -1067
rect 28164 -1119 28176 -1067
rect 28100 -1171 28176 -1119
rect 28100 -1223 28112 -1171
rect 28164 -1223 28176 -1171
rect 28100 -1235 28176 -1223
rect 28260 -1067 28336 -1055
rect 28260 -1119 28272 -1067
rect 28324 -1119 28336 -1067
rect 28260 -1171 28336 -1119
rect 28260 -1223 28272 -1171
rect 28324 -1223 28336 -1171
rect 28260 -1235 28336 -1223
rect 28420 -1067 28496 -1055
rect 28420 -1119 28432 -1067
rect 28484 -1119 28496 -1067
rect 28420 -1171 28496 -1119
rect 28420 -1223 28432 -1171
rect 28484 -1223 28496 -1171
rect 28420 -1235 28496 -1223
rect 28740 -1067 28816 -1055
rect 28740 -1119 28752 -1067
rect 28804 -1119 28816 -1067
rect 28740 -1171 28816 -1119
rect 28740 -1223 28752 -1171
rect 28804 -1223 28816 -1171
rect 28740 -1235 28816 -1223
rect 28900 -1067 28976 -1055
rect 28900 -1119 28912 -1067
rect 28964 -1119 28976 -1067
rect 28900 -1171 28976 -1119
rect 28900 -1223 28912 -1171
rect 28964 -1223 28976 -1171
rect 28900 -1235 28976 -1223
rect 29586 -1075 29779 -1029
rect 29825 -1075 29906 -1029
rect 29586 -1123 29906 -1075
rect 29586 -1169 29779 -1123
rect 29825 -1169 29906 -1123
rect 29586 -1217 29906 -1169
rect 26690 -1311 27010 -1263
rect 26690 -1357 26771 -1311
rect 26817 -1357 27010 -1311
rect 26690 -1405 27010 -1357
rect 26690 -1451 26771 -1405
rect 26817 -1451 27010 -1405
rect 26690 -1499 27010 -1451
rect 26690 -1545 26771 -1499
rect 26817 -1545 27010 -1499
rect 26690 -1593 27010 -1545
rect 26690 -1616 26771 -1593
rect 25856 -1639 26771 -1616
rect 26817 -1616 27010 -1593
rect 27347 -1616 27393 -1235
rect 27507 -1616 27553 -1235
rect 27795 -1294 27841 -1235
rect 28115 -1294 28161 -1235
rect 28435 -1294 28481 -1235
rect 28755 -1294 28801 -1235
rect 27795 -1340 28801 -1294
rect 27860 -1398 27936 -1386
rect 27860 -1450 27872 -1398
rect 27924 -1401 27936 -1398
rect 27924 -1447 28515 -1401
rect 28561 -1447 28572 -1401
rect 27924 -1450 27936 -1447
rect 27860 -1462 27936 -1450
rect 28755 -1616 28801 -1340
rect 29043 -1616 29089 -1235
rect 29203 -1616 29249 -1235
rect 29586 -1263 29779 -1217
rect 29825 -1263 29906 -1217
rect 29586 -1311 29906 -1263
rect 29586 -1357 29779 -1311
rect 29825 -1357 29906 -1311
rect 29586 -1405 29906 -1357
rect 29586 -1451 29779 -1405
rect 29825 -1451 29906 -1405
rect 29586 -1499 29906 -1451
rect 29586 -1545 29779 -1499
rect 29825 -1545 29906 -1499
rect 29586 -1593 29906 -1545
rect 29586 -1616 29779 -1593
rect 26817 -1639 29779 -1616
rect 29825 -1639 29906 -1593
rect 17569 -1687 29906 -1639
rect 17569 -1733 17650 -1687
rect 17696 -1733 20658 -1687
rect 20704 -1733 22802 -1687
rect 22848 -1733 25810 -1687
rect 25856 -1733 26771 -1687
rect 26817 -1733 29779 -1687
rect 29825 -1733 29906 -1687
rect 17569 -1781 29906 -1733
rect 17569 -1827 17650 -1781
rect 17696 -1827 17744 -1781
rect 17790 -1827 17838 -1781
rect 17884 -1827 17932 -1781
rect 17978 -1827 18026 -1781
rect 18072 -1827 18120 -1781
rect 18166 -1827 18214 -1781
rect 18260 -1827 18308 -1781
rect 18354 -1827 18402 -1781
rect 18448 -1827 18496 -1781
rect 18542 -1827 18590 -1781
rect 18636 -1827 18684 -1781
rect 18730 -1827 18778 -1781
rect 18824 -1827 18872 -1781
rect 18918 -1827 18966 -1781
rect 19012 -1827 19060 -1781
rect 19106 -1827 19154 -1781
rect 19200 -1827 19248 -1781
rect 19294 -1827 19342 -1781
rect 19388 -1827 19436 -1781
rect 19482 -1827 19530 -1781
rect 19576 -1827 19624 -1781
rect 19670 -1827 19718 -1781
rect 19764 -1827 19812 -1781
rect 19858 -1827 19906 -1781
rect 19952 -1827 20000 -1781
rect 20046 -1827 20094 -1781
rect 20140 -1827 20188 -1781
rect 20234 -1827 20282 -1781
rect 20328 -1827 20376 -1781
rect 20422 -1827 20470 -1781
rect 20516 -1827 20564 -1781
rect 20610 -1827 20658 -1781
rect 20704 -1827 22802 -1781
rect 22848 -1827 22896 -1781
rect 22942 -1827 22990 -1781
rect 23036 -1827 23084 -1781
rect 23130 -1827 23178 -1781
rect 23224 -1827 23272 -1781
rect 23318 -1827 23366 -1781
rect 23412 -1827 23460 -1781
rect 23506 -1827 23554 -1781
rect 23600 -1827 23648 -1781
rect 23694 -1827 23742 -1781
rect 23788 -1827 23836 -1781
rect 23882 -1827 23930 -1781
rect 23976 -1827 24024 -1781
rect 24070 -1827 24118 -1781
rect 24164 -1827 24212 -1781
rect 24258 -1827 24306 -1781
rect 24352 -1827 24400 -1781
rect 24446 -1827 24494 -1781
rect 24540 -1827 24588 -1781
rect 24634 -1827 24682 -1781
rect 24728 -1827 24776 -1781
rect 24822 -1827 24870 -1781
rect 24916 -1827 24964 -1781
rect 25010 -1827 25058 -1781
rect 25104 -1827 25152 -1781
rect 25198 -1827 25246 -1781
rect 25292 -1827 25340 -1781
rect 25386 -1827 25434 -1781
rect 25480 -1827 25528 -1781
rect 25574 -1827 25622 -1781
rect 25668 -1827 25716 -1781
rect 25762 -1827 25810 -1781
rect 25856 -1827 26771 -1781
rect 26817 -1827 26865 -1781
rect 26911 -1827 26959 -1781
rect 27005 -1827 27053 -1781
rect 27099 -1827 27147 -1781
rect 27193 -1827 27241 -1781
rect 27287 -1827 27335 -1781
rect 27381 -1827 27429 -1781
rect 27475 -1827 27523 -1781
rect 27569 -1827 27617 -1781
rect 27663 -1827 27711 -1781
rect 27757 -1827 27805 -1781
rect 27851 -1827 27899 -1781
rect 27945 -1827 27993 -1781
rect 28039 -1827 28087 -1781
rect 28133 -1827 28181 -1781
rect 28227 -1827 28275 -1781
rect 28321 -1827 28369 -1781
rect 28415 -1827 28463 -1781
rect 28509 -1827 28557 -1781
rect 28603 -1827 28651 -1781
rect 28697 -1827 28745 -1781
rect 28791 -1827 28839 -1781
rect 28885 -1827 28933 -1781
rect 28979 -1827 29027 -1781
rect 29073 -1827 29121 -1781
rect 29167 -1827 29215 -1781
rect 29261 -1827 29309 -1781
rect 29355 -1827 29403 -1781
rect 29449 -1827 29497 -1781
rect 29543 -1827 29591 -1781
rect 29637 -1827 29685 -1781
rect 29731 -1827 29779 -1781
rect 29825 -1827 29906 -1781
rect 17569 -1936 29906 -1827
rect 32024 4760 65532 5080
rect 32024 3182 32344 4760
rect 36160 3182 36480 4760
rect 40260 3182 40580 4760
rect 41720 3182 42040 4760
rect 45856 3182 46176 4760
rect 49956 3182 50276 4760
rect 51452 3182 51772 4760
rect 55552 3182 55872 4760
rect 59652 3182 59972 4760
rect 61112 3182 61432 4760
rect 65212 3182 65532 4760
rect 66428 3891 67202 3903
rect 66428 3839 66440 3891
rect 66492 3839 66544 3891
rect 66596 3839 66648 3891
rect 66700 3839 67202 3891
rect 66428 3787 67202 3839
rect 66428 3735 66440 3787
rect 66492 3735 66544 3787
rect 66596 3735 66648 3787
rect 66700 3735 67202 3787
rect 66428 3683 67202 3735
rect 66428 3631 66440 3683
rect 66492 3631 66544 3683
rect 66596 3631 66648 3683
rect 66700 3631 67202 3683
rect 66428 3619 67202 3631
rect 32024 3062 65532 3182
rect 32024 3016 32143 3062
rect 32189 3016 32237 3062
rect 32283 3016 32331 3062
rect 32377 3016 32425 3062
rect 32471 3016 32519 3062
rect 32565 3016 32613 3062
rect 32659 3016 32707 3062
rect 32753 3016 32801 3062
rect 32847 3016 32895 3062
rect 32941 3016 32989 3062
rect 33035 3016 33083 3062
rect 33129 3016 33177 3062
rect 33223 3016 33271 3062
rect 33317 3016 33365 3062
rect 33411 3016 33459 3062
rect 33505 3016 33553 3062
rect 33599 3016 33647 3062
rect 33693 3016 33741 3062
rect 33787 3016 33835 3062
rect 33881 3016 33929 3062
rect 33975 3016 34023 3062
rect 34069 3016 34117 3062
rect 34163 3016 34211 3062
rect 34257 3016 34305 3062
rect 34351 3016 34399 3062
rect 34445 3016 34493 3062
rect 34539 3016 34587 3062
rect 34633 3016 34681 3062
rect 34727 3016 34775 3062
rect 34821 3016 34869 3062
rect 34915 3016 34963 3062
rect 35009 3016 35057 3062
rect 35103 3016 35151 3062
rect 35197 3016 35245 3062
rect 35291 3016 35339 3062
rect 35385 3016 35433 3062
rect 35479 3016 35527 3062
rect 35573 3016 35621 3062
rect 35667 3016 35715 3062
rect 35761 3016 35809 3062
rect 35855 3016 35903 3062
rect 35949 3016 35997 3062
rect 36043 3016 36091 3062
rect 36137 3016 36185 3062
rect 36231 3016 36279 3062
rect 36325 3016 36373 3062
rect 36419 3016 36467 3062
rect 36513 3016 36561 3062
rect 36607 3016 36655 3062
rect 36701 3016 36749 3062
rect 36795 3016 36843 3062
rect 36889 3016 36937 3062
rect 36983 3016 37031 3062
rect 37077 3016 37125 3062
rect 37171 3016 37219 3062
rect 37265 3016 37313 3062
rect 37359 3016 37407 3062
rect 37453 3016 37501 3062
rect 37547 3016 37595 3062
rect 37641 3016 37689 3062
rect 37735 3016 37783 3062
rect 37829 3016 37877 3062
rect 37923 3016 37971 3062
rect 38017 3016 38065 3062
rect 38111 3016 38159 3062
rect 38205 3016 38253 3062
rect 38299 3016 38347 3062
rect 38393 3016 38441 3062
rect 38487 3016 38535 3062
rect 38581 3016 38629 3062
rect 38675 3016 38723 3062
rect 38769 3016 38817 3062
rect 38863 3016 38911 3062
rect 38957 3016 39005 3062
rect 39051 3016 39099 3062
rect 39145 3016 39193 3062
rect 39239 3016 39287 3062
rect 39333 3016 39381 3062
rect 39427 3016 39475 3062
rect 39521 3016 39569 3062
rect 39615 3016 39663 3062
rect 39709 3016 39757 3062
rect 39803 3016 39851 3062
rect 39897 3016 39945 3062
rect 39991 3016 40039 3062
rect 40085 3016 40133 3062
rect 40179 3016 40227 3062
rect 40273 3016 40321 3062
rect 40367 3016 40415 3062
rect 40461 3016 41839 3062
rect 41885 3016 41933 3062
rect 41979 3016 42027 3062
rect 42073 3016 42121 3062
rect 42167 3016 42215 3062
rect 42261 3016 42309 3062
rect 42355 3016 42403 3062
rect 42449 3016 42497 3062
rect 42543 3016 42591 3062
rect 42637 3016 42685 3062
rect 42731 3016 42779 3062
rect 42825 3016 42873 3062
rect 42919 3016 42967 3062
rect 43013 3016 43061 3062
rect 43107 3016 43155 3062
rect 43201 3016 43249 3062
rect 43295 3016 43343 3062
rect 43389 3016 43437 3062
rect 43483 3016 43531 3062
rect 43577 3016 43625 3062
rect 43671 3016 43719 3062
rect 43765 3016 43813 3062
rect 43859 3016 43907 3062
rect 43953 3016 44001 3062
rect 44047 3016 44095 3062
rect 44141 3016 44189 3062
rect 44235 3016 44283 3062
rect 44329 3016 44377 3062
rect 44423 3016 44471 3062
rect 44517 3016 44565 3062
rect 44611 3016 44659 3062
rect 44705 3016 44753 3062
rect 44799 3016 44847 3062
rect 44893 3016 44941 3062
rect 44987 3016 45035 3062
rect 45081 3016 45129 3062
rect 45175 3016 45223 3062
rect 45269 3016 45317 3062
rect 45363 3016 45411 3062
rect 45457 3016 45505 3062
rect 45551 3016 45599 3062
rect 45645 3016 45693 3062
rect 45739 3016 45787 3062
rect 45833 3016 45881 3062
rect 45927 3016 45975 3062
rect 46021 3016 46069 3062
rect 46115 3016 46163 3062
rect 46209 3016 46257 3062
rect 46303 3016 46351 3062
rect 46397 3016 46445 3062
rect 46491 3016 46539 3062
rect 46585 3016 46633 3062
rect 46679 3016 46727 3062
rect 46773 3016 46821 3062
rect 46867 3016 46915 3062
rect 46961 3016 47009 3062
rect 47055 3016 47103 3062
rect 47149 3016 47197 3062
rect 47243 3016 47291 3062
rect 47337 3016 47385 3062
rect 47431 3016 47479 3062
rect 47525 3016 47573 3062
rect 47619 3016 47667 3062
rect 47713 3016 47761 3062
rect 47807 3016 47855 3062
rect 47901 3016 47949 3062
rect 47995 3016 48043 3062
rect 48089 3016 48137 3062
rect 48183 3016 48231 3062
rect 48277 3016 48325 3062
rect 48371 3016 48419 3062
rect 48465 3016 48513 3062
rect 48559 3016 48607 3062
rect 48653 3016 48701 3062
rect 48747 3016 48795 3062
rect 48841 3016 48889 3062
rect 48935 3016 48983 3062
rect 49029 3016 49077 3062
rect 49123 3016 49171 3062
rect 49217 3016 49265 3062
rect 49311 3016 49359 3062
rect 49405 3016 49453 3062
rect 49499 3016 49547 3062
rect 49593 3016 49641 3062
rect 49687 3016 49735 3062
rect 49781 3016 49829 3062
rect 49875 3016 49923 3062
rect 49969 3016 50017 3062
rect 50063 3016 50111 3062
rect 50157 3016 51535 3062
rect 51581 3016 51629 3062
rect 51675 3016 51723 3062
rect 51769 3016 51817 3062
rect 51863 3016 51911 3062
rect 51957 3016 52005 3062
rect 52051 3016 52099 3062
rect 52145 3016 52193 3062
rect 52239 3016 52287 3062
rect 52333 3016 52381 3062
rect 52427 3016 52475 3062
rect 52521 3016 52569 3062
rect 52615 3016 52663 3062
rect 52709 3016 52757 3062
rect 52803 3016 52851 3062
rect 52897 3016 52945 3062
rect 52991 3016 53039 3062
rect 53085 3016 53133 3062
rect 53179 3016 53227 3062
rect 53273 3016 53321 3062
rect 53367 3016 53415 3062
rect 53461 3016 53509 3062
rect 53555 3016 53603 3062
rect 53649 3016 53697 3062
rect 53743 3016 53791 3062
rect 53837 3016 53885 3062
rect 53931 3016 53979 3062
rect 54025 3016 54073 3062
rect 54119 3016 54167 3062
rect 54213 3016 54261 3062
rect 54307 3016 54355 3062
rect 54401 3016 54449 3062
rect 54495 3016 54543 3062
rect 54589 3016 54637 3062
rect 54683 3016 54731 3062
rect 54777 3016 54825 3062
rect 54871 3016 54919 3062
rect 54965 3016 55013 3062
rect 55059 3016 55107 3062
rect 55153 3016 55201 3062
rect 55247 3016 55295 3062
rect 55341 3016 55389 3062
rect 55435 3016 55483 3062
rect 55529 3016 55577 3062
rect 55623 3016 55671 3062
rect 55717 3016 55765 3062
rect 55811 3016 55859 3062
rect 55905 3016 55953 3062
rect 55999 3016 56047 3062
rect 56093 3016 56141 3062
rect 56187 3016 56235 3062
rect 56281 3016 56329 3062
rect 56375 3016 56423 3062
rect 56469 3016 56517 3062
rect 56563 3016 56611 3062
rect 56657 3016 56705 3062
rect 56751 3016 56799 3062
rect 56845 3016 56893 3062
rect 56939 3016 56987 3062
rect 57033 3016 57081 3062
rect 57127 3016 57175 3062
rect 57221 3016 57269 3062
rect 57315 3016 57363 3062
rect 57409 3016 57457 3062
rect 57503 3016 57551 3062
rect 57597 3016 57645 3062
rect 57691 3016 57739 3062
rect 57785 3016 57833 3062
rect 57879 3016 57927 3062
rect 57973 3016 58021 3062
rect 58067 3016 58115 3062
rect 58161 3016 58209 3062
rect 58255 3016 58303 3062
rect 58349 3016 58397 3062
rect 58443 3016 58491 3062
rect 58537 3016 58585 3062
rect 58631 3016 58679 3062
rect 58725 3016 58773 3062
rect 58819 3016 58867 3062
rect 58913 3016 58961 3062
rect 59007 3016 59055 3062
rect 59101 3016 59149 3062
rect 59195 3016 59243 3062
rect 59289 3016 59337 3062
rect 59383 3016 59431 3062
rect 59477 3016 59525 3062
rect 59571 3016 59619 3062
rect 59665 3016 59713 3062
rect 59759 3016 59807 3062
rect 59853 3016 61231 3062
rect 61277 3016 61325 3062
rect 61371 3016 61419 3062
rect 61465 3016 61513 3062
rect 61559 3016 61607 3062
rect 61653 3016 61701 3062
rect 61747 3016 61795 3062
rect 61841 3016 61889 3062
rect 61935 3016 61983 3062
rect 62029 3016 62077 3062
rect 62123 3016 62171 3062
rect 62217 3016 62265 3062
rect 62311 3016 62359 3062
rect 62405 3016 62453 3062
rect 62499 3016 62547 3062
rect 62593 3016 62641 3062
rect 62687 3016 62735 3062
rect 62781 3016 62829 3062
rect 62875 3016 62923 3062
rect 62969 3016 63017 3062
rect 63063 3016 63111 3062
rect 63157 3016 63205 3062
rect 63251 3016 63299 3062
rect 63345 3016 63393 3062
rect 63439 3016 63487 3062
rect 63533 3016 63581 3062
rect 63627 3016 63675 3062
rect 63721 3016 63769 3062
rect 63815 3016 63863 3062
rect 63909 3016 63957 3062
rect 64003 3016 64051 3062
rect 64097 3016 64145 3062
rect 64191 3016 64239 3062
rect 64285 3016 64333 3062
rect 64379 3016 64427 3062
rect 64473 3016 64521 3062
rect 64567 3016 64615 3062
rect 64661 3016 64709 3062
rect 64755 3016 64803 3062
rect 64849 3016 64897 3062
rect 64943 3016 64991 3062
rect 65037 3016 65085 3062
rect 65131 3016 65179 3062
rect 65225 3016 65273 3062
rect 65319 3016 65367 3062
rect 65413 3016 65532 3062
rect 32024 2968 65532 3016
rect 32024 2922 32143 2968
rect 32189 2922 36279 2968
rect 36325 2922 40415 2968
rect 40461 2922 41839 2968
rect 41885 2922 45975 2968
rect 46021 2922 50111 2968
rect 50157 2922 51535 2968
rect 51581 2922 55671 2968
rect 55717 2922 59807 2968
rect 59853 2922 61231 2968
rect 61277 2922 65367 2968
rect 65413 2922 65532 2968
rect 32024 2874 65532 2922
rect 32024 2828 32143 2874
rect 32189 2862 36279 2874
rect 32189 2828 32344 2862
rect 32024 2780 32344 2828
rect 32024 2734 32143 2780
rect 32189 2734 32344 2780
rect 32024 2686 32344 2734
rect 32024 2640 32143 2686
rect 32189 2640 32344 2686
rect 32024 2592 32344 2640
rect 32024 2546 32143 2592
rect 32189 2546 32344 2592
rect 32024 2498 32344 2546
rect 32643 2519 32689 2862
rect 32803 2519 32849 2862
rect 32024 2452 32143 2498
rect 32189 2452 32344 2498
rect 32024 2404 32344 2452
rect 32024 2358 32143 2404
rect 32189 2358 32344 2404
rect 32024 2310 32344 2358
rect 32024 2264 32143 2310
rect 32189 2264 32344 2310
rect 32024 2216 32344 2264
rect 32024 2170 32143 2216
rect 32189 2170 32344 2216
rect 32024 2122 32344 2170
rect 32024 2076 32143 2122
rect 32189 2076 32344 2122
rect 32024 2028 32344 2076
rect 32024 1982 32143 2028
rect 32189 1982 32344 2028
rect 32024 1934 32344 1982
rect 32916 2113 32992 2125
rect 32916 2061 32928 2113
rect 32980 2061 32992 2113
rect 32916 2009 32992 2061
rect 32916 1957 32928 2009
rect 32980 1957 32992 2009
rect 32916 1945 32992 1957
rect 32024 1888 32143 1934
rect 32189 1888 32344 1934
rect 32024 1840 32344 1888
rect 32024 1794 32143 1840
rect 32189 1794 32344 1840
rect 32024 1746 32344 1794
rect 32024 1700 32143 1746
rect 32189 1700 32344 1746
rect 32024 1652 32344 1700
rect 32024 1606 32143 1652
rect 32189 1606 32344 1652
rect 32024 1558 32344 1606
rect 32024 1512 32143 1558
rect 32189 1512 32344 1558
rect 32024 1464 32344 1512
rect 32024 1418 32143 1464
rect 32189 1418 32344 1464
rect 32024 1370 32344 1418
rect 32024 1324 32143 1370
rect 32189 1324 32344 1370
rect 32024 1276 32344 1324
rect 32024 1230 32143 1276
rect 32189 1230 32344 1276
rect 32024 1182 32344 1230
rect 32024 1136 32143 1182
rect 32189 1136 32344 1182
rect 32024 1088 32344 1136
rect 32024 1042 32143 1088
rect 32189 1042 32344 1088
rect 32024 994 32344 1042
rect 32024 948 32143 994
rect 32189 948 32344 994
rect 32024 900 32344 948
rect 32024 854 32143 900
rect 32189 854 32344 900
rect 32024 806 32344 854
rect 32024 760 32143 806
rect 32189 760 32344 806
rect 32024 712 32344 760
rect 32024 666 32143 712
rect 32189 666 32344 712
rect 32024 618 32344 666
rect 32024 572 32143 618
rect 32189 572 32344 618
rect 32024 524 32344 572
rect 32024 478 32143 524
rect 32189 478 32344 524
rect 32024 430 32344 478
rect 32024 384 32143 430
rect 32189 384 32344 430
rect 32024 336 32344 384
rect 32024 290 32143 336
rect 32189 290 32344 336
rect 32024 242 32344 290
rect 32024 196 32143 242
rect 32189 196 32344 242
rect 32024 148 32344 196
rect 32024 102 32143 148
rect 32189 102 32344 148
rect 32024 54 32344 102
rect 32024 8 32143 54
rect 32189 8 32344 54
rect 32024 -40 32344 8
rect 32024 -86 32143 -40
rect 32189 -86 32344 -40
rect 32024 -134 32344 -86
rect 32024 -180 32143 -134
rect 32189 -180 32344 -134
rect 32024 -228 32344 -180
rect 32024 -274 32143 -228
rect 32189 -274 32344 -228
rect 32024 -322 32344 -274
rect 32024 -368 32143 -322
rect 32189 -368 32344 -322
rect 32024 -416 32344 -368
rect 32024 -462 32143 -416
rect 32189 -462 32344 -416
rect 32024 -510 32344 -462
rect 32024 -556 32143 -510
rect 32189 -556 32344 -510
rect 32024 -604 32344 -556
rect 32024 -650 32143 -604
rect 32189 -650 32344 -604
rect 32024 -698 32344 -650
rect 32024 -744 32143 -698
rect 32189 -744 32344 -698
rect 32024 -792 32344 -744
rect 32024 -838 32143 -792
rect 32189 -838 32344 -792
rect 32024 -886 32344 -838
rect 32024 -932 32143 -886
rect 32189 -932 32344 -886
rect 32024 -980 32344 -932
rect 32024 -1026 32143 -980
rect 32189 -1026 32344 -980
rect 32024 -1074 32344 -1026
rect 32024 -1120 32143 -1074
rect 32189 -1120 32344 -1074
rect 32024 -1168 32344 -1120
rect 32024 -1214 32143 -1168
rect 32189 -1214 32344 -1168
rect 32024 -1262 32344 -1214
rect 32024 -1308 32143 -1262
rect 32189 -1308 32344 -1262
rect 32024 -1356 32344 -1308
rect 32024 -1402 32143 -1356
rect 32189 -1402 32344 -1356
rect 32024 -1450 32344 -1402
rect 32024 -1496 32143 -1450
rect 32189 -1496 32344 -1450
rect 32024 -1544 32344 -1496
rect 32024 -1590 32143 -1544
rect 32189 -1578 32344 -1544
rect 32643 1725 32689 1945
rect 32803 1725 32849 1945
rect 32643 1679 32723 1725
rect 32769 1679 32849 1725
rect 32643 -395 32689 1679
rect 32803 -395 32849 1679
rect 32916 1053 32992 1065
rect 32916 1001 32928 1053
rect 32980 1001 32992 1053
rect 32916 949 32992 1001
rect 32916 897 32928 949
rect 32980 897 32992 949
rect 32916 885 32992 897
rect 32916 -7 32992 5
rect 32916 -59 32928 -7
rect 32980 -59 32992 -7
rect 32916 -111 32992 -59
rect 32916 -163 32928 -111
rect 32980 -163 32992 -111
rect 32916 -175 32992 -163
rect 32643 -441 32723 -395
rect 32769 -441 32849 -395
rect 32643 -1578 32689 -441
rect 32803 -1578 32849 -441
rect 32916 -1067 32992 -1055
rect 32916 -1119 32928 -1067
rect 32980 -1119 32992 -1067
rect 32916 -1171 32992 -1119
rect 32916 -1223 32928 -1171
rect 32980 -1223 32992 -1171
rect 32916 -1235 32992 -1223
rect 33091 -1578 33137 2862
rect 33237 2507 33313 2519
rect 33237 2455 33249 2507
rect 33301 2455 33313 2507
rect 33237 2403 33313 2455
rect 33237 2351 33249 2403
rect 33301 2351 33313 2403
rect 33237 2339 33313 2351
rect 33237 1447 33313 1459
rect 33237 1395 33249 1447
rect 33301 1395 33313 1447
rect 33237 1343 33313 1395
rect 33237 1291 33249 1343
rect 33301 1291 33313 1343
rect 33237 1279 33313 1291
rect 33237 387 33313 399
rect 33237 335 33249 387
rect 33301 335 33313 387
rect 33237 283 33313 335
rect 33237 231 33249 283
rect 33301 231 33313 283
rect 33237 219 33313 231
rect 33237 -673 33313 -661
rect 33237 -725 33249 -673
rect 33301 -725 33313 -673
rect 33237 -777 33313 -725
rect 33237 -829 33249 -777
rect 33301 -829 33313 -777
rect 33237 -841 33313 -829
rect 33411 -1578 33457 2862
rect 33556 2113 33632 2125
rect 33556 2061 33568 2113
rect 33620 2061 33632 2113
rect 33556 2009 33632 2061
rect 33556 1957 33568 2009
rect 33620 1957 33632 2009
rect 33556 1945 33632 1957
rect 33731 1888 33777 2862
rect 34116 2655 34192 2667
rect 34116 2603 34128 2655
rect 34180 2652 34192 2655
rect 34276 2655 34352 2667
rect 34276 2652 34288 2655
rect 34180 2603 34288 2652
rect 34340 2603 34352 2655
rect 34116 2591 34352 2603
rect 34211 2519 34257 2591
rect 33877 2507 33953 2519
rect 33877 2455 33889 2507
rect 33941 2455 33953 2507
rect 33877 2403 33953 2455
rect 33877 2351 33889 2403
rect 33941 2351 33953 2403
rect 33877 2339 33953 2351
rect 34517 2507 34593 2519
rect 34517 2455 34529 2507
rect 34581 2455 34593 2507
rect 34517 2403 34593 2455
rect 34517 2351 34529 2403
rect 34581 2351 34593 2403
rect 34517 2339 34593 2351
rect 34051 1888 34097 1945
rect 34371 1888 34417 1945
rect 33731 1842 34417 1888
rect 33556 1053 33632 1065
rect 33556 1001 33568 1053
rect 33620 1001 33632 1053
rect 33556 949 33632 1001
rect 33556 897 33568 949
rect 33620 897 33632 949
rect 33556 885 33632 897
rect 33731 828 33777 1842
rect 34116 1595 34192 1607
rect 34116 1543 34128 1595
rect 34180 1592 34192 1595
rect 34276 1595 34352 1607
rect 34276 1592 34288 1595
rect 34180 1543 34288 1592
rect 34340 1543 34352 1595
rect 34116 1531 34352 1543
rect 34211 1459 34257 1531
rect 33877 1447 33953 1459
rect 33877 1395 33889 1447
rect 33941 1395 33953 1447
rect 33877 1343 33953 1395
rect 33877 1291 33889 1343
rect 33941 1291 33953 1343
rect 33877 1279 33953 1291
rect 34517 1447 34593 1459
rect 34517 1395 34529 1447
rect 34581 1395 34593 1447
rect 34517 1343 34593 1395
rect 34517 1291 34529 1343
rect 34581 1291 34593 1343
rect 34517 1279 34593 1291
rect 34051 828 34097 885
rect 34371 828 34417 885
rect 33731 782 34417 828
rect 33556 -7 33632 5
rect 33556 -59 33568 -7
rect 33620 -59 33632 -7
rect 33556 -111 33632 -59
rect 33556 -163 33568 -111
rect 33620 -163 33632 -111
rect 33556 -175 33632 -163
rect 33731 -232 33777 782
rect 34116 535 34192 547
rect 34116 483 34128 535
rect 34180 532 34192 535
rect 34276 535 34352 547
rect 34276 532 34288 535
rect 34180 483 34288 532
rect 34340 483 34352 535
rect 34116 471 34352 483
rect 34211 399 34257 471
rect 33877 387 33953 399
rect 33877 335 33889 387
rect 33941 335 33953 387
rect 33877 283 33953 335
rect 33877 231 33889 283
rect 33941 231 33953 283
rect 33877 219 33953 231
rect 34517 387 34593 399
rect 34517 335 34529 387
rect 34581 335 34593 387
rect 34517 283 34593 335
rect 34517 231 34529 283
rect 34581 231 34593 283
rect 34517 219 34593 231
rect 34051 -232 34097 -175
rect 34371 -232 34417 -175
rect 33731 -278 34417 -232
rect 33556 -1067 33632 -1055
rect 33556 -1119 33568 -1067
rect 33620 -1119 33632 -1067
rect 33556 -1171 33632 -1119
rect 33556 -1223 33568 -1171
rect 33620 -1223 33632 -1171
rect 33556 -1235 33632 -1223
rect 33731 -1578 33777 -278
rect 34116 -525 34192 -513
rect 34116 -577 34128 -525
rect 34180 -528 34192 -525
rect 34276 -525 34352 -513
rect 34276 -528 34288 -525
rect 34180 -577 34288 -528
rect 34340 -577 34352 -525
rect 34116 -589 34352 -577
rect 34211 -661 34257 -589
rect 33877 -673 33953 -661
rect 33877 -725 33889 -673
rect 33941 -725 33953 -673
rect 33877 -777 33953 -725
rect 33877 -829 33889 -777
rect 33941 -829 33953 -777
rect 33877 -841 33953 -829
rect 34517 -673 34593 -661
rect 34517 -725 34529 -673
rect 34581 -725 34593 -673
rect 34517 -777 34593 -725
rect 34517 -829 34529 -777
rect 34581 -829 34593 -777
rect 34517 -841 34593 -829
rect 34051 -1578 34097 -1235
rect 34371 -1578 34417 -1235
rect 34691 -1578 34737 2862
rect 34836 2113 34912 2125
rect 34836 2061 34848 2113
rect 34900 2061 34912 2113
rect 34836 2009 34912 2061
rect 34836 1957 34848 2009
rect 34900 1957 34912 2009
rect 34836 1945 34912 1957
rect 34836 1053 34912 1065
rect 34836 1001 34848 1053
rect 34900 1001 34912 1053
rect 34836 949 34912 1001
rect 34836 897 34848 949
rect 34900 897 34912 949
rect 34836 885 34912 897
rect 34836 -7 34912 5
rect 34836 -59 34848 -7
rect 34900 -59 34912 -7
rect 34836 -111 34912 -59
rect 34836 -163 34848 -111
rect 34900 -163 34912 -111
rect 34836 -175 34912 -163
rect 34836 -1067 34912 -1055
rect 34836 -1119 34848 -1067
rect 34900 -1119 34912 -1067
rect 34836 -1171 34912 -1119
rect 34836 -1223 34848 -1171
rect 34900 -1223 34912 -1171
rect 34836 -1235 34912 -1223
rect 35011 -1578 35057 2862
rect 35157 2507 35233 2519
rect 35157 2455 35169 2507
rect 35221 2455 35233 2507
rect 35157 2403 35233 2455
rect 35157 2351 35169 2403
rect 35221 2351 35233 2403
rect 35157 2339 35233 2351
rect 35157 1447 35233 1459
rect 35157 1395 35169 1447
rect 35221 1395 35233 1447
rect 35157 1343 35233 1395
rect 35157 1291 35169 1343
rect 35221 1291 35233 1343
rect 35157 1279 35233 1291
rect 35157 387 35233 399
rect 35157 335 35169 387
rect 35221 335 35233 387
rect 35157 283 35233 335
rect 35157 231 35169 283
rect 35221 231 35233 283
rect 35157 219 35233 231
rect 35157 -673 35233 -661
rect 35157 -725 35169 -673
rect 35221 -725 35233 -673
rect 35157 -777 35233 -725
rect 35157 -829 35169 -777
rect 35221 -829 35233 -777
rect 35157 -841 35233 -829
rect 35331 -1578 35377 2862
rect 35619 2519 35665 2862
rect 35779 2519 35825 2862
rect 36124 2828 36279 2862
rect 36325 2862 40415 2874
rect 36325 2828 36480 2862
rect 36124 2780 36480 2828
rect 36124 2734 36279 2780
rect 36325 2734 36480 2780
rect 36124 2686 36480 2734
rect 36124 2640 36279 2686
rect 36325 2640 36480 2686
rect 36124 2592 36480 2640
rect 36124 2546 36279 2592
rect 36325 2546 36480 2592
rect 36124 2498 36480 2546
rect 36779 2519 36825 2862
rect 36939 2519 36985 2862
rect 36124 2452 36279 2498
rect 36325 2452 36480 2498
rect 36124 2404 36480 2452
rect 36124 2358 36279 2404
rect 36325 2358 36480 2404
rect 36124 2310 36480 2358
rect 36124 2264 36279 2310
rect 36325 2264 36480 2310
rect 36124 2216 36480 2264
rect 36124 2170 36279 2216
rect 36325 2170 36480 2216
rect 35476 2113 35552 2125
rect 35476 2061 35488 2113
rect 35540 2061 35552 2113
rect 35476 2009 35552 2061
rect 35476 1957 35488 2009
rect 35540 1957 35552 2009
rect 35476 1945 35552 1957
rect 36124 2122 36480 2170
rect 36124 2076 36279 2122
rect 36325 2076 36480 2122
rect 36124 2028 36480 2076
rect 36124 1982 36279 2028
rect 36325 1982 36480 2028
rect 35619 1725 35665 1945
rect 35779 1725 35825 1945
rect 35619 1679 35699 1725
rect 35745 1679 35825 1725
rect 35476 1053 35552 1065
rect 35476 1001 35488 1053
rect 35540 1001 35552 1053
rect 35476 949 35552 1001
rect 35476 897 35488 949
rect 35540 897 35552 949
rect 35476 885 35552 897
rect 35476 -7 35552 5
rect 35476 -59 35488 -7
rect 35540 -59 35552 -7
rect 35476 -111 35552 -59
rect 35476 -163 35488 -111
rect 35540 -163 35552 -111
rect 35476 -175 35552 -163
rect 35619 -395 35665 1679
rect 35779 -395 35825 1679
rect 35619 -441 35699 -395
rect 35745 -441 35825 -395
rect 35476 -1067 35552 -1055
rect 35476 -1119 35488 -1067
rect 35540 -1119 35552 -1067
rect 35476 -1171 35552 -1119
rect 35476 -1223 35488 -1171
rect 35540 -1223 35552 -1171
rect 35476 -1235 35552 -1223
rect 35619 -1578 35665 -441
rect 35779 -1578 35825 -441
rect 36124 1934 36480 1982
rect 37052 2113 37128 2125
rect 37052 2061 37064 2113
rect 37116 2061 37128 2113
rect 37052 2009 37128 2061
rect 37052 1957 37064 2009
rect 37116 1957 37128 2009
rect 37052 1945 37128 1957
rect 36124 1888 36279 1934
rect 36325 1888 36480 1934
rect 36124 1840 36480 1888
rect 36124 1794 36279 1840
rect 36325 1794 36480 1840
rect 36124 1746 36480 1794
rect 36124 1700 36279 1746
rect 36325 1700 36480 1746
rect 36124 1652 36480 1700
rect 36124 1606 36279 1652
rect 36325 1606 36480 1652
rect 36124 1558 36480 1606
rect 36124 1512 36279 1558
rect 36325 1512 36480 1558
rect 36124 1464 36480 1512
rect 36124 1418 36279 1464
rect 36325 1418 36480 1464
rect 36124 1370 36480 1418
rect 36124 1324 36279 1370
rect 36325 1324 36480 1370
rect 36124 1276 36480 1324
rect 36124 1230 36279 1276
rect 36325 1230 36480 1276
rect 36124 1182 36480 1230
rect 36124 1136 36279 1182
rect 36325 1136 36480 1182
rect 36124 1088 36480 1136
rect 36124 1042 36279 1088
rect 36325 1042 36480 1088
rect 36124 994 36480 1042
rect 36124 948 36279 994
rect 36325 948 36480 994
rect 36124 900 36480 948
rect 36124 854 36279 900
rect 36325 854 36480 900
rect 36124 806 36480 854
rect 36124 760 36279 806
rect 36325 760 36480 806
rect 36124 712 36480 760
rect 36124 666 36279 712
rect 36325 666 36480 712
rect 36124 618 36480 666
rect 36124 572 36279 618
rect 36325 572 36480 618
rect 36124 524 36480 572
rect 36124 478 36279 524
rect 36325 478 36480 524
rect 36124 430 36480 478
rect 36124 384 36279 430
rect 36325 384 36480 430
rect 36124 336 36480 384
rect 36124 290 36279 336
rect 36325 290 36480 336
rect 36124 242 36480 290
rect 36124 196 36279 242
rect 36325 196 36480 242
rect 36124 148 36480 196
rect 36124 102 36279 148
rect 36325 102 36480 148
rect 36124 54 36480 102
rect 36124 8 36279 54
rect 36325 8 36480 54
rect 36124 -40 36480 8
rect 36124 -86 36279 -40
rect 36325 -86 36480 -40
rect 36124 -134 36480 -86
rect 36124 -180 36279 -134
rect 36325 -180 36480 -134
rect 36124 -228 36480 -180
rect 36124 -274 36279 -228
rect 36325 -274 36480 -228
rect 36124 -322 36480 -274
rect 36124 -368 36279 -322
rect 36325 -368 36480 -322
rect 36124 -416 36480 -368
rect 36124 -462 36279 -416
rect 36325 -462 36480 -416
rect 36124 -510 36480 -462
rect 36124 -556 36279 -510
rect 36325 -556 36480 -510
rect 36124 -604 36480 -556
rect 36124 -650 36279 -604
rect 36325 -650 36480 -604
rect 36124 -698 36480 -650
rect 36124 -744 36279 -698
rect 36325 -744 36480 -698
rect 36124 -792 36480 -744
rect 36124 -838 36279 -792
rect 36325 -838 36480 -792
rect 36124 -886 36480 -838
rect 36124 -932 36279 -886
rect 36325 -932 36480 -886
rect 36124 -980 36480 -932
rect 36124 -1026 36279 -980
rect 36325 -1026 36480 -980
rect 36124 -1074 36480 -1026
rect 36124 -1120 36279 -1074
rect 36325 -1120 36480 -1074
rect 36124 -1168 36480 -1120
rect 36124 -1214 36279 -1168
rect 36325 -1214 36480 -1168
rect 36124 -1262 36480 -1214
rect 36124 -1308 36279 -1262
rect 36325 -1308 36480 -1262
rect 36124 -1356 36480 -1308
rect 36124 -1402 36279 -1356
rect 36325 -1402 36480 -1356
rect 36124 -1450 36480 -1402
rect 36124 -1496 36279 -1450
rect 36325 -1496 36480 -1450
rect 36124 -1544 36480 -1496
rect 36124 -1578 36279 -1544
rect 32189 -1590 36279 -1578
rect 36325 -1578 36480 -1544
rect 36779 1725 36825 1945
rect 36939 1725 36985 1945
rect 36779 1679 36859 1725
rect 36905 1679 36985 1725
rect 36779 -395 36825 1679
rect 36939 -395 36985 1679
rect 37052 1053 37128 1065
rect 37052 1001 37064 1053
rect 37116 1001 37128 1053
rect 37052 949 37128 1001
rect 37052 897 37064 949
rect 37116 897 37128 949
rect 37052 885 37128 897
rect 37052 -7 37128 5
rect 37052 -59 37064 -7
rect 37116 -59 37128 -7
rect 37052 -111 37128 -59
rect 37052 -163 37064 -111
rect 37116 -163 37128 -111
rect 37052 -175 37128 -163
rect 36779 -441 36859 -395
rect 36905 -441 36985 -395
rect 36779 -1578 36825 -441
rect 36939 -1578 36985 -441
rect 37052 -1067 37128 -1055
rect 37052 -1119 37064 -1067
rect 37116 -1119 37128 -1067
rect 37052 -1171 37128 -1119
rect 37052 -1223 37064 -1171
rect 37116 -1223 37128 -1171
rect 37052 -1235 37128 -1223
rect 37227 -1578 37273 2862
rect 37371 2507 37447 2519
rect 37371 2455 37383 2507
rect 37435 2455 37447 2507
rect 37371 2403 37447 2455
rect 37371 2351 37383 2403
rect 37435 2351 37447 2403
rect 37371 2339 37447 2351
rect 37371 1447 37447 1459
rect 37371 1395 37383 1447
rect 37435 1395 37447 1447
rect 37371 1343 37447 1395
rect 37371 1291 37383 1343
rect 37435 1291 37447 1343
rect 37371 1279 37447 1291
rect 37371 387 37447 399
rect 37371 335 37383 387
rect 37435 335 37447 387
rect 37371 283 37447 335
rect 37371 231 37383 283
rect 37435 231 37447 283
rect 37371 219 37447 231
rect 37371 -673 37447 -661
rect 37371 -725 37383 -673
rect 37435 -725 37447 -673
rect 37371 -777 37447 -725
rect 37371 -829 37383 -777
rect 37435 -829 37447 -777
rect 37371 -841 37447 -829
rect 37547 -1578 37593 2862
rect 37692 2113 37768 2125
rect 37692 2061 37704 2113
rect 37756 2061 37768 2113
rect 37692 2009 37768 2061
rect 37692 1957 37704 2009
rect 37756 1957 37768 2009
rect 37692 1945 37768 1957
rect 37692 1053 37768 1065
rect 37692 1001 37704 1053
rect 37756 1001 37768 1053
rect 37692 949 37768 1001
rect 37692 897 37704 949
rect 37756 897 37768 949
rect 37692 885 37768 897
rect 37692 -7 37768 5
rect 37692 -59 37704 -7
rect 37756 -59 37768 -7
rect 37692 -111 37768 -59
rect 37692 -163 37704 -111
rect 37756 -163 37768 -111
rect 37692 -175 37768 -163
rect 37692 -1067 37768 -1055
rect 37692 -1119 37704 -1067
rect 37756 -1119 37768 -1067
rect 37692 -1171 37768 -1119
rect 37692 -1223 37704 -1171
rect 37756 -1223 37768 -1171
rect 37692 -1235 37768 -1223
rect 37867 -1578 37913 2862
rect 38252 2655 38328 2667
rect 38252 2603 38264 2655
rect 38316 2652 38328 2655
rect 38412 2655 38488 2667
rect 38412 2652 38424 2655
rect 38316 2603 38424 2652
rect 38476 2603 38488 2655
rect 38252 2591 38488 2603
rect 38347 2519 38393 2591
rect 38011 2507 38087 2519
rect 38011 2455 38023 2507
rect 38075 2455 38087 2507
rect 38011 2403 38087 2455
rect 38011 2351 38023 2403
rect 38075 2351 38087 2403
rect 38011 2339 38087 2351
rect 38651 2507 38727 2519
rect 38651 2455 38663 2507
rect 38715 2455 38727 2507
rect 38651 2403 38727 2455
rect 38651 2351 38663 2403
rect 38715 2351 38727 2403
rect 38651 2339 38727 2351
rect 38187 1888 38233 1945
rect 38507 1888 38553 1945
rect 38827 1888 38873 2862
rect 38972 2113 39048 2125
rect 38972 2061 38984 2113
rect 39036 2061 39048 2113
rect 38972 2009 39048 2061
rect 38972 1957 38984 2009
rect 39036 1957 39048 2009
rect 38972 1945 39048 1957
rect 38187 1842 38873 1888
rect 38252 1595 38328 1607
rect 38252 1543 38264 1595
rect 38316 1592 38328 1595
rect 38412 1595 38488 1607
rect 38412 1592 38424 1595
rect 38316 1543 38424 1592
rect 38476 1543 38488 1595
rect 38252 1531 38488 1543
rect 38347 1459 38393 1531
rect 38011 1447 38087 1459
rect 38011 1395 38023 1447
rect 38075 1395 38087 1447
rect 38011 1343 38087 1395
rect 38011 1291 38023 1343
rect 38075 1291 38087 1343
rect 38011 1279 38087 1291
rect 38651 1447 38727 1459
rect 38651 1395 38663 1447
rect 38715 1395 38727 1447
rect 38651 1343 38727 1395
rect 38651 1291 38663 1343
rect 38715 1291 38727 1343
rect 38651 1279 38727 1291
rect 38187 828 38233 885
rect 38507 828 38553 885
rect 38827 828 38873 1842
rect 38972 1053 39048 1065
rect 38972 1001 38984 1053
rect 39036 1001 39048 1053
rect 38972 949 39048 1001
rect 38972 897 38984 949
rect 39036 897 39048 949
rect 38972 885 39048 897
rect 38187 782 38873 828
rect 38252 535 38328 547
rect 38252 483 38264 535
rect 38316 532 38328 535
rect 38412 535 38488 547
rect 38412 532 38424 535
rect 38316 483 38424 532
rect 38476 483 38488 535
rect 38252 471 38488 483
rect 38347 399 38393 471
rect 38011 387 38087 399
rect 38011 335 38023 387
rect 38075 335 38087 387
rect 38011 283 38087 335
rect 38011 231 38023 283
rect 38075 231 38087 283
rect 38011 219 38087 231
rect 38651 387 38727 399
rect 38651 335 38663 387
rect 38715 335 38727 387
rect 38651 283 38727 335
rect 38651 231 38663 283
rect 38715 231 38727 283
rect 38651 219 38727 231
rect 38187 -232 38233 -175
rect 38507 -232 38553 -175
rect 38827 -232 38873 782
rect 38972 -7 39048 5
rect 38972 -59 38984 -7
rect 39036 -59 39048 -7
rect 38972 -111 39048 -59
rect 38972 -163 38984 -111
rect 39036 -163 39048 -111
rect 38972 -175 39048 -163
rect 38187 -278 38873 -232
rect 38252 -525 38328 -513
rect 38252 -577 38264 -525
rect 38316 -528 38328 -525
rect 38412 -525 38488 -513
rect 38412 -528 38424 -525
rect 38316 -577 38424 -528
rect 38476 -577 38488 -525
rect 38252 -589 38488 -577
rect 38347 -661 38393 -589
rect 38011 -673 38087 -661
rect 38011 -725 38023 -673
rect 38075 -725 38087 -673
rect 38011 -777 38087 -725
rect 38011 -829 38023 -777
rect 38075 -829 38087 -777
rect 38011 -841 38087 -829
rect 38651 -673 38727 -661
rect 38651 -725 38663 -673
rect 38715 -725 38727 -673
rect 38651 -777 38727 -725
rect 38651 -829 38663 -777
rect 38715 -829 38727 -777
rect 38651 -841 38727 -829
rect 38187 -1578 38233 -1235
rect 38507 -1578 38553 -1235
rect 38827 -1578 38873 -278
rect 38972 -1067 39048 -1055
rect 38972 -1119 38984 -1067
rect 39036 -1119 39048 -1067
rect 38972 -1171 39048 -1119
rect 38972 -1223 38984 -1171
rect 39036 -1223 39048 -1171
rect 38972 -1235 39048 -1223
rect 39147 -1578 39193 2862
rect 39291 2507 39367 2519
rect 39291 2455 39303 2507
rect 39355 2455 39367 2507
rect 39291 2403 39367 2455
rect 39291 2351 39303 2403
rect 39355 2351 39367 2403
rect 39291 2339 39367 2351
rect 39291 1447 39367 1459
rect 39291 1395 39303 1447
rect 39355 1395 39367 1447
rect 39291 1343 39367 1395
rect 39291 1291 39303 1343
rect 39355 1291 39367 1343
rect 39291 1279 39367 1291
rect 39291 387 39367 399
rect 39291 335 39303 387
rect 39355 335 39367 387
rect 39291 283 39367 335
rect 39291 231 39303 283
rect 39355 231 39367 283
rect 39291 219 39367 231
rect 39291 -673 39367 -661
rect 39291 -725 39303 -673
rect 39355 -725 39367 -673
rect 39291 -777 39367 -725
rect 39291 -829 39303 -777
rect 39355 -829 39367 -777
rect 39291 -841 39367 -829
rect 39467 -1578 39513 2862
rect 39755 2519 39801 2862
rect 39915 2519 39961 2862
rect 40260 2828 40415 2862
rect 40461 2862 41839 2874
rect 40461 2828 40580 2862
rect 40260 2780 40580 2828
rect 40260 2734 40415 2780
rect 40461 2734 40580 2780
rect 40260 2686 40580 2734
rect 40260 2640 40415 2686
rect 40461 2640 40580 2686
rect 40260 2592 40580 2640
rect 40260 2546 40415 2592
rect 40461 2546 40580 2592
rect 40260 2498 40580 2546
rect 40260 2452 40415 2498
rect 40461 2452 40580 2498
rect 40260 2404 40580 2452
rect 40260 2358 40415 2404
rect 40461 2358 40580 2404
rect 40260 2310 40580 2358
rect 40260 2264 40415 2310
rect 40461 2264 40580 2310
rect 40260 2216 40580 2264
rect 40260 2170 40415 2216
rect 40461 2170 40580 2216
rect 39612 2113 39688 2125
rect 39612 2061 39624 2113
rect 39676 2061 39688 2113
rect 39612 2009 39688 2061
rect 39612 1957 39624 2009
rect 39676 1957 39688 2009
rect 39612 1945 39688 1957
rect 40260 2122 40580 2170
rect 40260 2076 40415 2122
rect 40461 2076 40580 2122
rect 40260 2028 40580 2076
rect 40260 1982 40415 2028
rect 40461 1982 40580 2028
rect 39755 1725 39801 1945
rect 39915 1725 39961 1945
rect 39755 1679 39835 1725
rect 39881 1679 39961 1725
rect 39612 1053 39688 1065
rect 39612 1001 39624 1053
rect 39676 1001 39688 1053
rect 39612 949 39688 1001
rect 39612 897 39624 949
rect 39676 897 39688 949
rect 39612 885 39688 897
rect 39612 -7 39688 5
rect 39612 -59 39624 -7
rect 39676 -59 39688 -7
rect 39612 -111 39688 -59
rect 39612 -163 39624 -111
rect 39676 -163 39688 -111
rect 39612 -175 39688 -163
rect 39755 -395 39801 1679
rect 39915 -395 39961 1679
rect 39755 -441 39835 -395
rect 39881 -441 39961 -395
rect 39612 -1067 39688 -1055
rect 39612 -1119 39624 -1067
rect 39676 -1119 39688 -1067
rect 39612 -1171 39688 -1119
rect 39612 -1223 39624 -1171
rect 39676 -1223 39688 -1171
rect 39612 -1235 39688 -1223
rect 39755 -1578 39801 -441
rect 39915 -1578 39961 -441
rect 40260 1934 40580 1982
rect 40260 1888 40415 1934
rect 40461 1888 40580 1934
rect 40260 1840 40580 1888
rect 40260 1794 40415 1840
rect 40461 1794 40580 1840
rect 40260 1746 40580 1794
rect 40260 1700 40415 1746
rect 40461 1700 40580 1746
rect 40260 1652 40580 1700
rect 40260 1606 40415 1652
rect 40461 1606 40580 1652
rect 40260 1558 40580 1606
rect 40260 1512 40415 1558
rect 40461 1512 40580 1558
rect 40260 1464 40580 1512
rect 40260 1418 40415 1464
rect 40461 1418 40580 1464
rect 40260 1370 40580 1418
rect 40260 1324 40415 1370
rect 40461 1324 40580 1370
rect 40260 1276 40580 1324
rect 40260 1230 40415 1276
rect 40461 1230 40580 1276
rect 40260 1182 40580 1230
rect 40260 1136 40415 1182
rect 40461 1136 40580 1182
rect 40260 1088 40580 1136
rect 40260 1042 40415 1088
rect 40461 1042 40580 1088
rect 40260 994 40580 1042
rect 40260 948 40415 994
rect 40461 948 40580 994
rect 40260 900 40580 948
rect 40260 854 40415 900
rect 40461 854 40580 900
rect 40260 806 40580 854
rect 40260 760 40415 806
rect 40461 760 40580 806
rect 40260 712 40580 760
rect 40260 666 40415 712
rect 40461 666 40580 712
rect 40260 618 40580 666
rect 40260 572 40415 618
rect 40461 572 40580 618
rect 40260 524 40580 572
rect 40260 478 40415 524
rect 40461 478 40580 524
rect 40260 430 40580 478
rect 40260 384 40415 430
rect 40461 384 40580 430
rect 40260 336 40580 384
rect 40260 290 40415 336
rect 40461 290 40580 336
rect 40260 242 40580 290
rect 40260 196 40415 242
rect 40461 196 40580 242
rect 40260 148 40580 196
rect 40260 102 40415 148
rect 40461 102 40580 148
rect 40260 54 40580 102
rect 40260 8 40415 54
rect 40461 8 40580 54
rect 40260 -40 40580 8
rect 40260 -86 40415 -40
rect 40461 -86 40580 -40
rect 40260 -134 40580 -86
rect 40260 -180 40415 -134
rect 40461 -180 40580 -134
rect 40260 -228 40580 -180
rect 40260 -274 40415 -228
rect 40461 -274 40580 -228
rect 40260 -322 40580 -274
rect 40260 -368 40415 -322
rect 40461 -368 40580 -322
rect 40260 -416 40580 -368
rect 40260 -462 40415 -416
rect 40461 -462 40580 -416
rect 40260 -510 40580 -462
rect 40260 -556 40415 -510
rect 40461 -556 40580 -510
rect 40260 -604 40580 -556
rect 40260 -650 40415 -604
rect 40461 -650 40580 -604
rect 40260 -698 40580 -650
rect 40260 -744 40415 -698
rect 40461 -744 40580 -698
rect 40260 -792 40580 -744
rect 40260 -838 40415 -792
rect 40461 -838 40580 -792
rect 40260 -886 40580 -838
rect 40260 -932 40415 -886
rect 40461 -932 40580 -886
rect 40260 -980 40580 -932
rect 40260 -1026 40415 -980
rect 40461 -1026 40580 -980
rect 40260 -1074 40580 -1026
rect 40260 -1120 40415 -1074
rect 40461 -1120 40580 -1074
rect 40260 -1168 40580 -1120
rect 40260 -1214 40415 -1168
rect 40461 -1214 40580 -1168
rect 40260 -1262 40580 -1214
rect 40260 -1308 40415 -1262
rect 40461 -1308 40580 -1262
rect 40260 -1356 40580 -1308
rect 40260 -1402 40415 -1356
rect 40461 -1402 40580 -1356
rect 40260 -1450 40580 -1402
rect 40260 -1496 40415 -1450
rect 40461 -1496 40580 -1450
rect 40260 -1544 40580 -1496
rect 40260 -1578 40415 -1544
rect 36325 -1590 40415 -1578
rect 40461 -1578 40580 -1544
rect 41720 2828 41839 2862
rect 41885 2862 45975 2874
rect 41885 2828 42040 2862
rect 41720 2780 42040 2828
rect 41720 2734 41839 2780
rect 41885 2734 42040 2780
rect 41720 2686 42040 2734
rect 41720 2640 41839 2686
rect 41885 2640 42040 2686
rect 41720 2592 42040 2640
rect 41720 2546 41839 2592
rect 41885 2546 42040 2592
rect 41720 2498 42040 2546
rect 42339 2519 42385 2862
rect 42499 2519 42545 2862
rect 41720 2452 41839 2498
rect 41885 2452 42040 2498
rect 41720 2404 42040 2452
rect 41720 2358 41839 2404
rect 41885 2358 42040 2404
rect 41720 2310 42040 2358
rect 41720 2264 41839 2310
rect 41885 2264 42040 2310
rect 41720 2216 42040 2264
rect 41720 2170 41839 2216
rect 41885 2170 42040 2216
rect 41720 2122 42040 2170
rect 41720 2076 41839 2122
rect 41885 2076 42040 2122
rect 41720 2028 42040 2076
rect 41720 1982 41839 2028
rect 41885 1982 42040 2028
rect 41720 1934 42040 1982
rect 42612 2113 42688 2125
rect 42612 2061 42624 2113
rect 42676 2061 42688 2113
rect 42612 2009 42688 2061
rect 42612 1957 42624 2009
rect 42676 1957 42688 2009
rect 42612 1945 42688 1957
rect 41720 1888 41839 1934
rect 41885 1888 42040 1934
rect 41720 1840 42040 1888
rect 41720 1794 41839 1840
rect 41885 1794 42040 1840
rect 41720 1746 42040 1794
rect 41720 1700 41839 1746
rect 41885 1700 42040 1746
rect 41720 1652 42040 1700
rect 41720 1606 41839 1652
rect 41885 1606 42040 1652
rect 41720 1558 42040 1606
rect 41720 1512 41839 1558
rect 41885 1512 42040 1558
rect 41720 1464 42040 1512
rect 41720 1418 41839 1464
rect 41885 1418 42040 1464
rect 41720 1370 42040 1418
rect 41720 1324 41839 1370
rect 41885 1324 42040 1370
rect 41720 1276 42040 1324
rect 41720 1230 41839 1276
rect 41885 1230 42040 1276
rect 41720 1182 42040 1230
rect 41720 1136 41839 1182
rect 41885 1136 42040 1182
rect 41720 1088 42040 1136
rect 41720 1042 41839 1088
rect 41885 1042 42040 1088
rect 41720 994 42040 1042
rect 41720 948 41839 994
rect 41885 948 42040 994
rect 41720 900 42040 948
rect 41720 854 41839 900
rect 41885 854 42040 900
rect 41720 806 42040 854
rect 41720 760 41839 806
rect 41885 760 42040 806
rect 41720 712 42040 760
rect 41720 666 41839 712
rect 41885 666 42040 712
rect 41720 618 42040 666
rect 41720 572 41839 618
rect 41885 572 42040 618
rect 41720 524 42040 572
rect 41720 478 41839 524
rect 41885 478 42040 524
rect 41720 430 42040 478
rect 41720 384 41839 430
rect 41885 384 42040 430
rect 41720 336 42040 384
rect 41720 290 41839 336
rect 41885 290 42040 336
rect 41720 242 42040 290
rect 41720 196 41839 242
rect 41885 196 42040 242
rect 41720 148 42040 196
rect 41720 102 41839 148
rect 41885 102 42040 148
rect 41720 54 42040 102
rect 41720 8 41839 54
rect 41885 8 42040 54
rect 41720 -40 42040 8
rect 41720 -86 41839 -40
rect 41885 -86 42040 -40
rect 41720 -134 42040 -86
rect 41720 -180 41839 -134
rect 41885 -180 42040 -134
rect 41720 -228 42040 -180
rect 41720 -274 41839 -228
rect 41885 -274 42040 -228
rect 41720 -322 42040 -274
rect 41720 -368 41839 -322
rect 41885 -368 42040 -322
rect 41720 -416 42040 -368
rect 41720 -462 41839 -416
rect 41885 -462 42040 -416
rect 41720 -510 42040 -462
rect 41720 -556 41839 -510
rect 41885 -556 42040 -510
rect 41720 -604 42040 -556
rect 41720 -650 41839 -604
rect 41885 -650 42040 -604
rect 41720 -698 42040 -650
rect 41720 -744 41839 -698
rect 41885 -744 42040 -698
rect 41720 -792 42040 -744
rect 41720 -838 41839 -792
rect 41885 -838 42040 -792
rect 41720 -886 42040 -838
rect 41720 -932 41839 -886
rect 41885 -932 42040 -886
rect 41720 -980 42040 -932
rect 41720 -1026 41839 -980
rect 41885 -1026 42040 -980
rect 41720 -1074 42040 -1026
rect 41720 -1120 41839 -1074
rect 41885 -1120 42040 -1074
rect 41720 -1168 42040 -1120
rect 41720 -1214 41839 -1168
rect 41885 -1214 42040 -1168
rect 41720 -1262 42040 -1214
rect 41720 -1308 41839 -1262
rect 41885 -1308 42040 -1262
rect 41720 -1356 42040 -1308
rect 41720 -1402 41839 -1356
rect 41885 -1402 42040 -1356
rect 41720 -1450 42040 -1402
rect 41720 -1496 41839 -1450
rect 41885 -1496 42040 -1450
rect 41720 -1544 42040 -1496
rect 41720 -1578 41839 -1544
rect 40461 -1590 41839 -1578
rect 41885 -1578 42040 -1544
rect 42339 1725 42385 1945
rect 42499 1725 42545 1945
rect 42339 1679 42419 1725
rect 42465 1679 42545 1725
rect 42339 -395 42385 1679
rect 42499 -395 42545 1679
rect 42612 1053 42688 1065
rect 42612 1001 42624 1053
rect 42676 1001 42688 1053
rect 42612 949 42688 1001
rect 42612 897 42624 949
rect 42676 897 42688 949
rect 42612 885 42688 897
rect 42612 -7 42688 5
rect 42612 -59 42624 -7
rect 42676 -59 42688 -7
rect 42612 -111 42688 -59
rect 42612 -163 42624 -111
rect 42676 -163 42688 -111
rect 42612 -175 42688 -163
rect 42339 -441 42419 -395
rect 42465 -441 42545 -395
rect 42339 -1578 42385 -441
rect 42499 -1578 42545 -441
rect 42612 -1067 42688 -1055
rect 42612 -1119 42624 -1067
rect 42676 -1119 42688 -1067
rect 42612 -1171 42688 -1119
rect 42612 -1223 42624 -1171
rect 42676 -1223 42688 -1171
rect 42612 -1235 42688 -1223
rect 42787 -1578 42833 2862
rect 42933 2507 43009 2519
rect 42933 2455 42945 2507
rect 42997 2455 43009 2507
rect 42933 2403 43009 2455
rect 42933 2351 42945 2403
rect 42997 2351 43009 2403
rect 42933 2339 43009 2351
rect 42933 1447 43009 1459
rect 42933 1395 42945 1447
rect 42997 1395 43009 1447
rect 42933 1343 43009 1395
rect 42933 1291 42945 1343
rect 42997 1291 43009 1343
rect 42933 1279 43009 1291
rect 42933 387 43009 399
rect 42933 335 42945 387
rect 42997 335 43009 387
rect 42933 283 43009 335
rect 42933 231 42945 283
rect 42997 231 43009 283
rect 42933 219 43009 231
rect 42933 -673 43009 -661
rect 42933 -725 42945 -673
rect 42997 -725 43009 -673
rect 42933 -777 43009 -725
rect 42933 -829 42945 -777
rect 42997 -829 43009 -777
rect 42933 -841 43009 -829
rect 43107 -1578 43153 2862
rect 43252 2113 43328 2125
rect 43252 2061 43264 2113
rect 43316 2061 43328 2113
rect 43252 2009 43328 2061
rect 43252 1957 43264 2009
rect 43316 1957 43328 2009
rect 43252 1945 43328 1957
rect 43427 1888 43473 2862
rect 43812 2655 43888 2667
rect 43812 2603 43824 2655
rect 43876 2652 43888 2655
rect 43972 2655 44048 2667
rect 43972 2652 43984 2655
rect 43876 2603 43984 2652
rect 44036 2603 44048 2655
rect 43812 2591 44048 2603
rect 43907 2519 43953 2591
rect 43573 2507 43649 2519
rect 43573 2455 43585 2507
rect 43637 2455 43649 2507
rect 43573 2403 43649 2455
rect 43573 2351 43585 2403
rect 43637 2351 43649 2403
rect 43573 2339 43649 2351
rect 44213 2507 44289 2519
rect 44213 2455 44225 2507
rect 44277 2455 44289 2507
rect 44213 2403 44289 2455
rect 44213 2351 44225 2403
rect 44277 2351 44289 2403
rect 44213 2339 44289 2351
rect 43747 1888 43793 1945
rect 44067 1888 44113 1945
rect 43427 1842 44113 1888
rect 43252 1053 43328 1065
rect 43252 1001 43264 1053
rect 43316 1001 43328 1053
rect 43252 949 43328 1001
rect 43252 897 43264 949
rect 43316 897 43328 949
rect 43252 885 43328 897
rect 43427 828 43473 1842
rect 43812 1595 43888 1607
rect 43812 1543 43824 1595
rect 43876 1592 43888 1595
rect 43972 1595 44048 1607
rect 43972 1592 43984 1595
rect 43876 1543 43984 1592
rect 44036 1543 44048 1595
rect 43812 1531 44048 1543
rect 43907 1459 43953 1531
rect 43573 1447 43649 1459
rect 43573 1395 43585 1447
rect 43637 1395 43649 1447
rect 43573 1343 43649 1395
rect 43573 1291 43585 1343
rect 43637 1291 43649 1343
rect 43573 1279 43649 1291
rect 44213 1447 44289 1459
rect 44213 1395 44225 1447
rect 44277 1395 44289 1447
rect 44213 1343 44289 1395
rect 44213 1291 44225 1343
rect 44277 1291 44289 1343
rect 44213 1279 44289 1291
rect 43747 828 43793 885
rect 44067 828 44113 885
rect 43427 782 44113 828
rect 43252 -7 43328 5
rect 43252 -59 43264 -7
rect 43316 -59 43328 -7
rect 43252 -111 43328 -59
rect 43252 -163 43264 -111
rect 43316 -163 43328 -111
rect 43252 -175 43328 -163
rect 43427 -232 43473 782
rect 43812 535 43888 547
rect 43812 483 43824 535
rect 43876 532 43888 535
rect 43972 535 44048 547
rect 43972 532 43984 535
rect 43876 483 43984 532
rect 44036 483 44048 535
rect 43812 471 44048 483
rect 43907 399 43953 471
rect 43573 387 43649 399
rect 43573 335 43585 387
rect 43637 335 43649 387
rect 43573 283 43649 335
rect 43573 231 43585 283
rect 43637 231 43649 283
rect 43573 219 43649 231
rect 44213 387 44289 399
rect 44213 335 44225 387
rect 44277 335 44289 387
rect 44213 283 44289 335
rect 44213 231 44225 283
rect 44277 231 44289 283
rect 44213 219 44289 231
rect 43747 -232 43793 -175
rect 44067 -232 44113 -175
rect 43427 -278 44113 -232
rect 43252 -1067 43328 -1055
rect 43252 -1119 43264 -1067
rect 43316 -1119 43328 -1067
rect 43252 -1171 43328 -1119
rect 43252 -1223 43264 -1171
rect 43316 -1223 43328 -1171
rect 43252 -1235 43328 -1223
rect 43427 -1578 43473 -278
rect 43812 -525 43888 -513
rect 43812 -577 43824 -525
rect 43876 -528 43888 -525
rect 43972 -525 44048 -513
rect 43972 -528 43984 -525
rect 43876 -577 43984 -528
rect 44036 -577 44048 -525
rect 43812 -589 44048 -577
rect 43907 -661 43953 -589
rect 43573 -673 43649 -661
rect 43573 -725 43585 -673
rect 43637 -725 43649 -673
rect 43573 -777 43649 -725
rect 43573 -829 43585 -777
rect 43637 -829 43649 -777
rect 43573 -841 43649 -829
rect 44213 -673 44289 -661
rect 44213 -725 44225 -673
rect 44277 -725 44289 -673
rect 44213 -777 44289 -725
rect 44213 -829 44225 -777
rect 44277 -829 44289 -777
rect 44213 -841 44289 -829
rect 43747 -1578 43793 -1235
rect 44067 -1578 44113 -1235
rect 44387 -1578 44433 2862
rect 44532 2113 44608 2125
rect 44532 2061 44544 2113
rect 44596 2061 44608 2113
rect 44532 2009 44608 2061
rect 44532 1957 44544 2009
rect 44596 1957 44608 2009
rect 44532 1945 44608 1957
rect 44532 1053 44608 1065
rect 44532 1001 44544 1053
rect 44596 1001 44608 1053
rect 44532 949 44608 1001
rect 44532 897 44544 949
rect 44596 897 44608 949
rect 44532 885 44608 897
rect 44532 -7 44608 5
rect 44532 -59 44544 -7
rect 44596 -59 44608 -7
rect 44532 -111 44608 -59
rect 44532 -163 44544 -111
rect 44596 -163 44608 -111
rect 44532 -175 44608 -163
rect 44532 -1067 44608 -1055
rect 44532 -1119 44544 -1067
rect 44596 -1119 44608 -1067
rect 44532 -1171 44608 -1119
rect 44532 -1223 44544 -1171
rect 44596 -1223 44608 -1171
rect 44532 -1235 44608 -1223
rect 44707 -1578 44753 2862
rect 44853 2507 44929 2519
rect 44853 2455 44865 2507
rect 44917 2455 44929 2507
rect 44853 2403 44929 2455
rect 44853 2351 44865 2403
rect 44917 2351 44929 2403
rect 44853 2339 44929 2351
rect 44853 1447 44929 1459
rect 44853 1395 44865 1447
rect 44917 1395 44929 1447
rect 44853 1343 44929 1395
rect 44853 1291 44865 1343
rect 44917 1291 44929 1343
rect 44853 1279 44929 1291
rect 44853 387 44929 399
rect 44853 335 44865 387
rect 44917 335 44929 387
rect 44853 283 44929 335
rect 44853 231 44865 283
rect 44917 231 44929 283
rect 44853 219 44929 231
rect 44853 -673 44929 -661
rect 44853 -725 44865 -673
rect 44917 -725 44929 -673
rect 44853 -777 44929 -725
rect 44853 -829 44865 -777
rect 44917 -829 44929 -777
rect 44853 -841 44929 -829
rect 45027 -1578 45073 2862
rect 45315 2519 45361 2862
rect 45475 2519 45521 2862
rect 45820 2828 45975 2862
rect 46021 2862 50111 2874
rect 46021 2828 46176 2862
rect 45820 2780 46176 2828
rect 45820 2734 45975 2780
rect 46021 2734 46176 2780
rect 45820 2686 46176 2734
rect 45820 2640 45975 2686
rect 46021 2640 46176 2686
rect 45820 2592 46176 2640
rect 45820 2546 45975 2592
rect 46021 2546 46176 2592
rect 45820 2498 46176 2546
rect 46475 2519 46521 2862
rect 46635 2519 46681 2862
rect 45820 2452 45975 2498
rect 46021 2452 46176 2498
rect 45820 2404 46176 2452
rect 45820 2358 45975 2404
rect 46021 2358 46176 2404
rect 45820 2310 46176 2358
rect 45820 2264 45975 2310
rect 46021 2264 46176 2310
rect 45820 2216 46176 2264
rect 45820 2170 45975 2216
rect 46021 2170 46176 2216
rect 45172 2113 45248 2125
rect 45172 2061 45184 2113
rect 45236 2061 45248 2113
rect 45172 2009 45248 2061
rect 45172 1957 45184 2009
rect 45236 1957 45248 2009
rect 45172 1945 45248 1957
rect 45820 2122 46176 2170
rect 45820 2076 45975 2122
rect 46021 2076 46176 2122
rect 45820 2028 46176 2076
rect 45820 1982 45975 2028
rect 46021 1982 46176 2028
rect 45315 1725 45361 1945
rect 45475 1725 45521 1945
rect 45315 1679 45395 1725
rect 45441 1679 45521 1725
rect 45172 1053 45248 1065
rect 45172 1001 45184 1053
rect 45236 1001 45248 1053
rect 45172 949 45248 1001
rect 45172 897 45184 949
rect 45236 897 45248 949
rect 45172 885 45248 897
rect 45172 -7 45248 5
rect 45172 -59 45184 -7
rect 45236 -59 45248 -7
rect 45172 -111 45248 -59
rect 45172 -163 45184 -111
rect 45236 -163 45248 -111
rect 45172 -175 45248 -163
rect 45315 -395 45361 1679
rect 45475 -395 45521 1679
rect 45315 -441 45395 -395
rect 45441 -441 45521 -395
rect 45172 -1067 45248 -1055
rect 45172 -1119 45184 -1067
rect 45236 -1119 45248 -1067
rect 45172 -1171 45248 -1119
rect 45172 -1223 45184 -1171
rect 45236 -1223 45248 -1171
rect 45172 -1235 45248 -1223
rect 45315 -1578 45361 -441
rect 45475 -1578 45521 -441
rect 45820 1934 46176 1982
rect 46748 2113 46824 2125
rect 46748 2061 46760 2113
rect 46812 2061 46824 2113
rect 46748 2009 46824 2061
rect 46748 1957 46760 2009
rect 46812 1957 46824 2009
rect 46748 1945 46824 1957
rect 45820 1888 45975 1934
rect 46021 1888 46176 1934
rect 45820 1840 46176 1888
rect 45820 1794 45975 1840
rect 46021 1794 46176 1840
rect 45820 1746 46176 1794
rect 45820 1700 45975 1746
rect 46021 1700 46176 1746
rect 45820 1652 46176 1700
rect 45820 1606 45975 1652
rect 46021 1606 46176 1652
rect 45820 1558 46176 1606
rect 45820 1512 45975 1558
rect 46021 1512 46176 1558
rect 45820 1464 46176 1512
rect 45820 1418 45975 1464
rect 46021 1418 46176 1464
rect 45820 1370 46176 1418
rect 45820 1324 45975 1370
rect 46021 1324 46176 1370
rect 45820 1276 46176 1324
rect 45820 1230 45975 1276
rect 46021 1230 46176 1276
rect 45820 1182 46176 1230
rect 45820 1136 45975 1182
rect 46021 1136 46176 1182
rect 45820 1088 46176 1136
rect 45820 1042 45975 1088
rect 46021 1042 46176 1088
rect 45820 994 46176 1042
rect 45820 948 45975 994
rect 46021 948 46176 994
rect 45820 900 46176 948
rect 45820 854 45975 900
rect 46021 854 46176 900
rect 45820 806 46176 854
rect 45820 760 45975 806
rect 46021 760 46176 806
rect 45820 712 46176 760
rect 45820 666 45975 712
rect 46021 666 46176 712
rect 45820 618 46176 666
rect 45820 572 45975 618
rect 46021 572 46176 618
rect 45820 524 46176 572
rect 45820 478 45975 524
rect 46021 478 46176 524
rect 45820 430 46176 478
rect 45820 384 45975 430
rect 46021 384 46176 430
rect 45820 336 46176 384
rect 45820 290 45975 336
rect 46021 290 46176 336
rect 45820 242 46176 290
rect 45820 196 45975 242
rect 46021 196 46176 242
rect 45820 148 46176 196
rect 45820 102 45975 148
rect 46021 102 46176 148
rect 45820 54 46176 102
rect 45820 8 45975 54
rect 46021 8 46176 54
rect 45820 -40 46176 8
rect 45820 -86 45975 -40
rect 46021 -86 46176 -40
rect 45820 -134 46176 -86
rect 45820 -180 45975 -134
rect 46021 -180 46176 -134
rect 45820 -228 46176 -180
rect 45820 -274 45975 -228
rect 46021 -274 46176 -228
rect 45820 -322 46176 -274
rect 45820 -368 45975 -322
rect 46021 -368 46176 -322
rect 45820 -416 46176 -368
rect 45820 -462 45975 -416
rect 46021 -462 46176 -416
rect 45820 -510 46176 -462
rect 45820 -556 45975 -510
rect 46021 -556 46176 -510
rect 45820 -604 46176 -556
rect 45820 -650 45975 -604
rect 46021 -650 46176 -604
rect 45820 -698 46176 -650
rect 45820 -744 45975 -698
rect 46021 -744 46176 -698
rect 45820 -792 46176 -744
rect 45820 -838 45975 -792
rect 46021 -838 46176 -792
rect 45820 -886 46176 -838
rect 45820 -932 45975 -886
rect 46021 -932 46176 -886
rect 45820 -980 46176 -932
rect 45820 -1026 45975 -980
rect 46021 -1026 46176 -980
rect 45820 -1074 46176 -1026
rect 45820 -1120 45975 -1074
rect 46021 -1120 46176 -1074
rect 45820 -1168 46176 -1120
rect 45820 -1214 45975 -1168
rect 46021 -1214 46176 -1168
rect 45820 -1262 46176 -1214
rect 45820 -1308 45975 -1262
rect 46021 -1308 46176 -1262
rect 45820 -1356 46176 -1308
rect 45820 -1402 45975 -1356
rect 46021 -1402 46176 -1356
rect 45820 -1450 46176 -1402
rect 45820 -1496 45975 -1450
rect 46021 -1496 46176 -1450
rect 45820 -1544 46176 -1496
rect 45820 -1578 45975 -1544
rect 41885 -1590 45975 -1578
rect 46021 -1578 46176 -1544
rect 46475 1725 46521 1945
rect 46635 1725 46681 1945
rect 46475 1679 46555 1725
rect 46601 1679 46681 1725
rect 46475 -395 46521 1679
rect 46635 -395 46681 1679
rect 46748 1053 46824 1065
rect 46748 1001 46760 1053
rect 46812 1001 46824 1053
rect 46748 949 46824 1001
rect 46748 897 46760 949
rect 46812 897 46824 949
rect 46748 885 46824 897
rect 46748 -7 46824 5
rect 46748 -59 46760 -7
rect 46812 -59 46824 -7
rect 46748 -111 46824 -59
rect 46748 -163 46760 -111
rect 46812 -163 46824 -111
rect 46748 -175 46824 -163
rect 46475 -441 46555 -395
rect 46601 -441 46681 -395
rect 46475 -1578 46521 -441
rect 46635 -1578 46681 -441
rect 46748 -1067 46824 -1055
rect 46748 -1119 46760 -1067
rect 46812 -1119 46824 -1067
rect 46748 -1171 46824 -1119
rect 46748 -1223 46760 -1171
rect 46812 -1223 46824 -1171
rect 46748 -1235 46824 -1223
rect 46923 -1578 46969 2862
rect 47067 2507 47143 2519
rect 47067 2455 47079 2507
rect 47131 2455 47143 2507
rect 47067 2403 47143 2455
rect 47067 2351 47079 2403
rect 47131 2351 47143 2403
rect 47067 2339 47143 2351
rect 47067 1447 47143 1459
rect 47067 1395 47079 1447
rect 47131 1395 47143 1447
rect 47067 1343 47143 1395
rect 47067 1291 47079 1343
rect 47131 1291 47143 1343
rect 47067 1279 47143 1291
rect 47067 387 47143 399
rect 47067 335 47079 387
rect 47131 335 47143 387
rect 47067 283 47143 335
rect 47067 231 47079 283
rect 47131 231 47143 283
rect 47067 219 47143 231
rect 47067 -673 47143 -661
rect 47067 -725 47079 -673
rect 47131 -725 47143 -673
rect 47067 -777 47143 -725
rect 47067 -829 47079 -777
rect 47131 -829 47143 -777
rect 47067 -841 47143 -829
rect 47243 -1578 47289 2862
rect 47388 2113 47464 2125
rect 47388 2061 47400 2113
rect 47452 2061 47464 2113
rect 47388 2009 47464 2061
rect 47388 1957 47400 2009
rect 47452 1957 47464 2009
rect 47388 1945 47464 1957
rect 47388 1053 47464 1065
rect 47388 1001 47400 1053
rect 47452 1001 47464 1053
rect 47388 949 47464 1001
rect 47388 897 47400 949
rect 47452 897 47464 949
rect 47388 885 47464 897
rect 47388 -7 47464 5
rect 47388 -59 47400 -7
rect 47452 -59 47464 -7
rect 47388 -111 47464 -59
rect 47388 -163 47400 -111
rect 47452 -163 47464 -111
rect 47388 -175 47464 -163
rect 47388 -1067 47464 -1055
rect 47388 -1119 47400 -1067
rect 47452 -1119 47464 -1067
rect 47388 -1171 47464 -1119
rect 47388 -1223 47400 -1171
rect 47452 -1223 47464 -1171
rect 47388 -1235 47464 -1223
rect 47563 -1578 47609 2862
rect 47948 2655 48024 2667
rect 47948 2603 47960 2655
rect 48012 2652 48024 2655
rect 48108 2655 48184 2667
rect 48108 2652 48120 2655
rect 48012 2603 48120 2652
rect 48172 2603 48184 2655
rect 47948 2591 48184 2603
rect 48043 2519 48089 2591
rect 47707 2507 47783 2519
rect 47707 2455 47719 2507
rect 47771 2455 47783 2507
rect 47707 2403 47783 2455
rect 47707 2351 47719 2403
rect 47771 2351 47783 2403
rect 47707 2339 47783 2351
rect 48347 2507 48423 2519
rect 48347 2455 48359 2507
rect 48411 2455 48423 2507
rect 48347 2403 48423 2455
rect 48347 2351 48359 2403
rect 48411 2351 48423 2403
rect 48347 2339 48423 2351
rect 47883 1888 47929 1945
rect 48203 1888 48249 1945
rect 48523 1888 48569 2862
rect 48668 2113 48744 2125
rect 48668 2061 48680 2113
rect 48732 2061 48744 2113
rect 48668 2009 48744 2061
rect 48668 1957 48680 2009
rect 48732 1957 48744 2009
rect 48668 1945 48744 1957
rect 47883 1842 48569 1888
rect 47948 1595 48024 1607
rect 47948 1543 47960 1595
rect 48012 1592 48024 1595
rect 48108 1595 48184 1607
rect 48108 1592 48120 1595
rect 48012 1543 48120 1592
rect 48172 1543 48184 1595
rect 47948 1531 48184 1543
rect 48043 1459 48089 1531
rect 47707 1447 47783 1459
rect 47707 1395 47719 1447
rect 47771 1395 47783 1447
rect 47707 1343 47783 1395
rect 47707 1291 47719 1343
rect 47771 1291 47783 1343
rect 47707 1279 47783 1291
rect 48347 1447 48423 1459
rect 48347 1395 48359 1447
rect 48411 1395 48423 1447
rect 48347 1343 48423 1395
rect 48347 1291 48359 1343
rect 48411 1291 48423 1343
rect 48347 1279 48423 1291
rect 47883 828 47929 885
rect 48203 828 48249 885
rect 48523 828 48569 1842
rect 48668 1053 48744 1065
rect 48668 1001 48680 1053
rect 48732 1001 48744 1053
rect 48668 949 48744 1001
rect 48668 897 48680 949
rect 48732 897 48744 949
rect 48668 885 48744 897
rect 47883 782 48569 828
rect 47948 535 48024 547
rect 47948 483 47960 535
rect 48012 532 48024 535
rect 48108 535 48184 547
rect 48108 532 48120 535
rect 48012 483 48120 532
rect 48172 483 48184 535
rect 47948 471 48184 483
rect 48043 399 48089 471
rect 47707 387 47783 399
rect 47707 335 47719 387
rect 47771 335 47783 387
rect 47707 283 47783 335
rect 47707 231 47719 283
rect 47771 231 47783 283
rect 47707 219 47783 231
rect 48347 387 48423 399
rect 48347 335 48359 387
rect 48411 335 48423 387
rect 48347 283 48423 335
rect 48347 231 48359 283
rect 48411 231 48423 283
rect 48347 219 48423 231
rect 47883 -232 47929 -175
rect 48203 -232 48249 -175
rect 48523 -232 48569 782
rect 48668 -7 48744 5
rect 48668 -59 48680 -7
rect 48732 -59 48744 -7
rect 48668 -111 48744 -59
rect 48668 -163 48680 -111
rect 48732 -163 48744 -111
rect 48668 -175 48744 -163
rect 47883 -278 48569 -232
rect 47948 -525 48024 -513
rect 47948 -577 47960 -525
rect 48012 -528 48024 -525
rect 48108 -525 48184 -513
rect 48108 -528 48120 -525
rect 48012 -577 48120 -528
rect 48172 -577 48184 -525
rect 47948 -589 48184 -577
rect 48043 -661 48089 -589
rect 47707 -673 47783 -661
rect 47707 -725 47719 -673
rect 47771 -725 47783 -673
rect 47707 -777 47783 -725
rect 47707 -829 47719 -777
rect 47771 -829 47783 -777
rect 47707 -841 47783 -829
rect 48347 -673 48423 -661
rect 48347 -725 48359 -673
rect 48411 -725 48423 -673
rect 48347 -777 48423 -725
rect 48347 -829 48359 -777
rect 48411 -829 48423 -777
rect 48347 -841 48423 -829
rect 47883 -1578 47929 -1235
rect 48203 -1578 48249 -1235
rect 48523 -1578 48569 -278
rect 48668 -1067 48744 -1055
rect 48668 -1119 48680 -1067
rect 48732 -1119 48744 -1067
rect 48668 -1171 48744 -1119
rect 48668 -1223 48680 -1171
rect 48732 -1223 48744 -1171
rect 48668 -1235 48744 -1223
rect 48843 -1578 48889 2862
rect 48987 2507 49063 2519
rect 48987 2455 48999 2507
rect 49051 2455 49063 2507
rect 48987 2403 49063 2455
rect 48987 2351 48999 2403
rect 49051 2351 49063 2403
rect 48987 2339 49063 2351
rect 48987 1447 49063 1459
rect 48987 1395 48999 1447
rect 49051 1395 49063 1447
rect 48987 1343 49063 1395
rect 48987 1291 48999 1343
rect 49051 1291 49063 1343
rect 48987 1279 49063 1291
rect 48987 387 49063 399
rect 48987 335 48999 387
rect 49051 335 49063 387
rect 48987 283 49063 335
rect 48987 231 48999 283
rect 49051 231 49063 283
rect 48987 219 49063 231
rect 48987 -673 49063 -661
rect 48987 -725 48999 -673
rect 49051 -725 49063 -673
rect 48987 -777 49063 -725
rect 48987 -829 48999 -777
rect 49051 -829 49063 -777
rect 48987 -841 49063 -829
rect 49163 -1578 49209 2862
rect 49451 2519 49497 2862
rect 49611 2519 49657 2862
rect 49956 2828 50111 2862
rect 50157 2862 51535 2874
rect 50157 2828 50276 2862
rect 49956 2780 50276 2828
rect 49956 2734 50111 2780
rect 50157 2734 50276 2780
rect 49956 2686 50276 2734
rect 49956 2640 50111 2686
rect 50157 2640 50276 2686
rect 49956 2592 50276 2640
rect 49956 2546 50111 2592
rect 50157 2546 50276 2592
rect 49956 2498 50276 2546
rect 49956 2452 50111 2498
rect 50157 2452 50276 2498
rect 49956 2404 50276 2452
rect 49956 2358 50111 2404
rect 50157 2358 50276 2404
rect 49956 2310 50276 2358
rect 49956 2264 50111 2310
rect 50157 2264 50276 2310
rect 49956 2216 50276 2264
rect 49956 2170 50111 2216
rect 50157 2170 50276 2216
rect 49308 2113 49384 2125
rect 49308 2061 49320 2113
rect 49372 2061 49384 2113
rect 49308 2009 49384 2061
rect 49308 1957 49320 2009
rect 49372 1957 49384 2009
rect 49308 1945 49384 1957
rect 49956 2122 50276 2170
rect 49956 2076 50111 2122
rect 50157 2076 50276 2122
rect 49956 2028 50276 2076
rect 49956 1982 50111 2028
rect 50157 1982 50276 2028
rect 49451 1725 49497 1945
rect 49611 1725 49657 1945
rect 49451 1679 49531 1725
rect 49577 1679 49657 1725
rect 49308 1053 49384 1065
rect 49308 1001 49320 1053
rect 49372 1001 49384 1053
rect 49308 949 49384 1001
rect 49308 897 49320 949
rect 49372 897 49384 949
rect 49308 885 49384 897
rect 49308 -7 49384 5
rect 49308 -59 49320 -7
rect 49372 -59 49384 -7
rect 49308 -111 49384 -59
rect 49308 -163 49320 -111
rect 49372 -163 49384 -111
rect 49308 -175 49384 -163
rect 49451 -395 49497 1679
rect 49611 -395 49657 1679
rect 49451 -441 49531 -395
rect 49577 -441 49657 -395
rect 49308 -1067 49384 -1055
rect 49308 -1119 49320 -1067
rect 49372 -1119 49384 -1067
rect 49308 -1171 49384 -1119
rect 49308 -1223 49320 -1171
rect 49372 -1223 49384 -1171
rect 49308 -1235 49384 -1223
rect 49451 -1578 49497 -441
rect 49611 -1578 49657 -441
rect 49956 1934 50276 1982
rect 49956 1888 50111 1934
rect 50157 1888 50276 1934
rect 49956 1840 50276 1888
rect 49956 1794 50111 1840
rect 50157 1794 50276 1840
rect 49956 1746 50276 1794
rect 49956 1700 50111 1746
rect 50157 1700 50276 1746
rect 49956 1652 50276 1700
rect 49956 1606 50111 1652
rect 50157 1606 50276 1652
rect 49956 1558 50276 1606
rect 49956 1512 50111 1558
rect 50157 1512 50276 1558
rect 49956 1464 50276 1512
rect 49956 1418 50111 1464
rect 50157 1418 50276 1464
rect 49956 1370 50276 1418
rect 49956 1324 50111 1370
rect 50157 1324 50276 1370
rect 49956 1276 50276 1324
rect 49956 1230 50111 1276
rect 50157 1230 50276 1276
rect 49956 1182 50276 1230
rect 49956 1136 50111 1182
rect 50157 1136 50276 1182
rect 49956 1088 50276 1136
rect 49956 1042 50111 1088
rect 50157 1042 50276 1088
rect 49956 994 50276 1042
rect 49956 948 50111 994
rect 50157 948 50276 994
rect 49956 900 50276 948
rect 49956 854 50111 900
rect 50157 854 50276 900
rect 49956 806 50276 854
rect 49956 760 50111 806
rect 50157 760 50276 806
rect 49956 712 50276 760
rect 49956 666 50111 712
rect 50157 666 50276 712
rect 49956 618 50276 666
rect 49956 572 50111 618
rect 50157 572 50276 618
rect 49956 524 50276 572
rect 49956 478 50111 524
rect 50157 478 50276 524
rect 49956 430 50276 478
rect 49956 384 50111 430
rect 50157 384 50276 430
rect 49956 336 50276 384
rect 49956 290 50111 336
rect 50157 290 50276 336
rect 49956 242 50276 290
rect 49956 196 50111 242
rect 50157 196 50276 242
rect 49956 148 50276 196
rect 49956 102 50111 148
rect 50157 102 50276 148
rect 49956 54 50276 102
rect 49956 8 50111 54
rect 50157 8 50276 54
rect 49956 -40 50276 8
rect 49956 -86 50111 -40
rect 50157 -86 50276 -40
rect 49956 -134 50276 -86
rect 49956 -180 50111 -134
rect 50157 -180 50276 -134
rect 49956 -228 50276 -180
rect 49956 -274 50111 -228
rect 50157 -274 50276 -228
rect 49956 -322 50276 -274
rect 49956 -368 50111 -322
rect 50157 -368 50276 -322
rect 49956 -416 50276 -368
rect 49956 -462 50111 -416
rect 50157 -462 50276 -416
rect 49956 -510 50276 -462
rect 49956 -556 50111 -510
rect 50157 -556 50276 -510
rect 49956 -604 50276 -556
rect 49956 -650 50111 -604
rect 50157 -650 50276 -604
rect 49956 -698 50276 -650
rect 49956 -744 50111 -698
rect 50157 -744 50276 -698
rect 49956 -792 50276 -744
rect 49956 -838 50111 -792
rect 50157 -838 50276 -792
rect 49956 -886 50276 -838
rect 49956 -932 50111 -886
rect 50157 -932 50276 -886
rect 49956 -980 50276 -932
rect 49956 -1026 50111 -980
rect 50157 -1026 50276 -980
rect 49956 -1074 50276 -1026
rect 49956 -1120 50111 -1074
rect 50157 -1120 50276 -1074
rect 49956 -1168 50276 -1120
rect 49956 -1214 50111 -1168
rect 50157 -1214 50276 -1168
rect 49956 -1262 50276 -1214
rect 49956 -1308 50111 -1262
rect 50157 -1308 50276 -1262
rect 49956 -1356 50276 -1308
rect 49956 -1402 50111 -1356
rect 50157 -1402 50276 -1356
rect 49956 -1450 50276 -1402
rect 49956 -1496 50111 -1450
rect 50157 -1496 50276 -1450
rect 49956 -1544 50276 -1496
rect 49956 -1578 50111 -1544
rect 46021 -1590 50111 -1578
rect 50157 -1578 50276 -1544
rect 51416 2828 51535 2862
rect 51581 2862 55671 2874
rect 51581 2828 51736 2862
rect 51416 2780 51736 2828
rect 51416 2734 51535 2780
rect 51581 2734 51736 2780
rect 51416 2686 51736 2734
rect 51416 2640 51535 2686
rect 51581 2640 51736 2686
rect 51416 2592 51736 2640
rect 51416 2546 51535 2592
rect 51581 2546 51736 2592
rect 51416 2498 51736 2546
rect 52035 2519 52081 2862
rect 52195 2519 52241 2862
rect 51416 2452 51535 2498
rect 51581 2452 51736 2498
rect 51416 2404 51736 2452
rect 51416 2358 51535 2404
rect 51581 2358 51736 2404
rect 51416 2310 51736 2358
rect 51416 2264 51535 2310
rect 51581 2264 51736 2310
rect 51416 2216 51736 2264
rect 51416 2170 51535 2216
rect 51581 2170 51736 2216
rect 51416 2122 51736 2170
rect 51416 2076 51535 2122
rect 51581 2076 51736 2122
rect 51416 2028 51736 2076
rect 51416 1982 51535 2028
rect 51581 1982 51736 2028
rect 51416 1934 51736 1982
rect 52308 2113 52384 2125
rect 52308 2061 52320 2113
rect 52372 2061 52384 2113
rect 52308 2009 52384 2061
rect 52308 1957 52320 2009
rect 52372 1957 52384 2009
rect 52308 1945 52384 1957
rect 51416 1888 51535 1934
rect 51581 1888 51736 1934
rect 51416 1840 51736 1888
rect 51416 1794 51535 1840
rect 51581 1794 51736 1840
rect 51416 1746 51736 1794
rect 51416 1700 51535 1746
rect 51581 1700 51736 1746
rect 51416 1652 51736 1700
rect 51416 1606 51535 1652
rect 51581 1606 51736 1652
rect 51416 1558 51736 1606
rect 51416 1512 51535 1558
rect 51581 1512 51736 1558
rect 51416 1464 51736 1512
rect 51416 1418 51535 1464
rect 51581 1418 51736 1464
rect 51416 1370 51736 1418
rect 51416 1324 51535 1370
rect 51581 1324 51736 1370
rect 51416 1276 51736 1324
rect 51416 1230 51535 1276
rect 51581 1230 51736 1276
rect 51416 1182 51736 1230
rect 51416 1136 51535 1182
rect 51581 1136 51736 1182
rect 51416 1088 51736 1136
rect 51416 1042 51535 1088
rect 51581 1042 51736 1088
rect 51416 994 51736 1042
rect 51416 948 51535 994
rect 51581 948 51736 994
rect 51416 900 51736 948
rect 51416 854 51535 900
rect 51581 854 51736 900
rect 51416 806 51736 854
rect 51416 760 51535 806
rect 51581 760 51736 806
rect 51416 712 51736 760
rect 51416 666 51535 712
rect 51581 666 51736 712
rect 51416 618 51736 666
rect 51416 572 51535 618
rect 51581 572 51736 618
rect 51416 524 51736 572
rect 51416 478 51535 524
rect 51581 478 51736 524
rect 51416 430 51736 478
rect 51416 384 51535 430
rect 51581 384 51736 430
rect 51416 336 51736 384
rect 51416 290 51535 336
rect 51581 290 51736 336
rect 51416 242 51736 290
rect 51416 196 51535 242
rect 51581 196 51736 242
rect 51416 148 51736 196
rect 51416 102 51535 148
rect 51581 102 51736 148
rect 51416 54 51736 102
rect 51416 8 51535 54
rect 51581 8 51736 54
rect 51416 -40 51736 8
rect 51416 -86 51535 -40
rect 51581 -86 51736 -40
rect 51416 -134 51736 -86
rect 51416 -180 51535 -134
rect 51581 -180 51736 -134
rect 51416 -228 51736 -180
rect 51416 -274 51535 -228
rect 51581 -274 51736 -228
rect 51416 -322 51736 -274
rect 51416 -368 51535 -322
rect 51581 -368 51736 -322
rect 51416 -416 51736 -368
rect 51416 -462 51535 -416
rect 51581 -462 51736 -416
rect 51416 -510 51736 -462
rect 51416 -556 51535 -510
rect 51581 -556 51736 -510
rect 51416 -604 51736 -556
rect 51416 -650 51535 -604
rect 51581 -650 51736 -604
rect 51416 -698 51736 -650
rect 51416 -744 51535 -698
rect 51581 -744 51736 -698
rect 51416 -792 51736 -744
rect 51416 -838 51535 -792
rect 51581 -838 51736 -792
rect 51416 -886 51736 -838
rect 51416 -932 51535 -886
rect 51581 -932 51736 -886
rect 51416 -980 51736 -932
rect 51416 -1026 51535 -980
rect 51581 -1026 51736 -980
rect 51416 -1074 51736 -1026
rect 51416 -1120 51535 -1074
rect 51581 -1120 51736 -1074
rect 51416 -1168 51736 -1120
rect 51416 -1214 51535 -1168
rect 51581 -1214 51736 -1168
rect 51416 -1262 51736 -1214
rect 51416 -1308 51535 -1262
rect 51581 -1308 51736 -1262
rect 51416 -1356 51736 -1308
rect 51416 -1402 51535 -1356
rect 51581 -1402 51736 -1356
rect 51416 -1450 51736 -1402
rect 51416 -1496 51535 -1450
rect 51581 -1496 51736 -1450
rect 51416 -1544 51736 -1496
rect 51416 -1578 51535 -1544
rect 50157 -1590 51535 -1578
rect 51581 -1578 51736 -1544
rect 52035 1725 52081 1945
rect 52195 1725 52241 1945
rect 52035 1679 52115 1725
rect 52161 1679 52241 1725
rect 52035 -395 52081 1679
rect 52195 -395 52241 1679
rect 52308 1053 52384 1065
rect 52308 1001 52320 1053
rect 52372 1001 52384 1053
rect 52308 949 52384 1001
rect 52308 897 52320 949
rect 52372 897 52384 949
rect 52308 885 52384 897
rect 52308 -7 52384 5
rect 52308 -59 52320 -7
rect 52372 -59 52384 -7
rect 52308 -111 52384 -59
rect 52308 -163 52320 -111
rect 52372 -163 52384 -111
rect 52308 -175 52384 -163
rect 52035 -441 52115 -395
rect 52161 -441 52241 -395
rect 52035 -1578 52081 -441
rect 52195 -1578 52241 -441
rect 52308 -1067 52384 -1055
rect 52308 -1119 52320 -1067
rect 52372 -1119 52384 -1067
rect 52308 -1171 52384 -1119
rect 52308 -1223 52320 -1171
rect 52372 -1223 52384 -1171
rect 52308 -1235 52384 -1223
rect 52483 -1578 52529 2862
rect 52629 2507 52705 2519
rect 52629 2455 52641 2507
rect 52693 2455 52705 2507
rect 52629 2403 52705 2455
rect 52629 2351 52641 2403
rect 52693 2351 52705 2403
rect 52629 2339 52705 2351
rect 52629 1447 52705 1459
rect 52629 1395 52641 1447
rect 52693 1395 52705 1447
rect 52629 1343 52705 1395
rect 52629 1291 52641 1343
rect 52693 1291 52705 1343
rect 52629 1279 52705 1291
rect 52629 387 52705 399
rect 52629 335 52641 387
rect 52693 335 52705 387
rect 52629 283 52705 335
rect 52629 231 52641 283
rect 52693 231 52705 283
rect 52629 219 52705 231
rect 52629 -673 52705 -661
rect 52629 -725 52641 -673
rect 52693 -725 52705 -673
rect 52629 -777 52705 -725
rect 52629 -829 52641 -777
rect 52693 -829 52705 -777
rect 52629 -841 52705 -829
rect 52803 -1578 52849 2862
rect 52948 2113 53024 2125
rect 52948 2061 52960 2113
rect 53012 2061 53024 2113
rect 52948 2009 53024 2061
rect 52948 1957 52960 2009
rect 53012 1957 53024 2009
rect 52948 1945 53024 1957
rect 53123 1888 53169 2862
rect 53508 2655 53584 2667
rect 53508 2603 53520 2655
rect 53572 2652 53584 2655
rect 53668 2655 53744 2667
rect 53668 2652 53680 2655
rect 53572 2603 53680 2652
rect 53732 2603 53744 2655
rect 53508 2591 53744 2603
rect 53603 2519 53649 2591
rect 53269 2507 53345 2519
rect 53269 2455 53281 2507
rect 53333 2455 53345 2507
rect 53269 2403 53345 2455
rect 53269 2351 53281 2403
rect 53333 2351 53345 2403
rect 53269 2339 53345 2351
rect 53909 2507 53985 2519
rect 53909 2455 53921 2507
rect 53973 2455 53985 2507
rect 53909 2403 53985 2455
rect 53909 2351 53921 2403
rect 53973 2351 53985 2403
rect 53909 2339 53985 2351
rect 53443 1888 53489 1945
rect 53763 1888 53809 1945
rect 53123 1842 53809 1888
rect 52948 1053 53024 1065
rect 52948 1001 52960 1053
rect 53012 1001 53024 1053
rect 52948 949 53024 1001
rect 52948 897 52960 949
rect 53012 897 53024 949
rect 52948 885 53024 897
rect 53123 828 53169 1842
rect 53508 1595 53584 1607
rect 53508 1543 53520 1595
rect 53572 1592 53584 1595
rect 53668 1595 53744 1607
rect 53668 1592 53680 1595
rect 53572 1543 53680 1592
rect 53732 1543 53744 1595
rect 53508 1531 53744 1543
rect 53603 1459 53649 1531
rect 53269 1447 53345 1459
rect 53269 1395 53281 1447
rect 53333 1395 53345 1447
rect 53269 1343 53345 1395
rect 53269 1291 53281 1343
rect 53333 1291 53345 1343
rect 53269 1279 53345 1291
rect 53909 1447 53985 1459
rect 53909 1395 53921 1447
rect 53973 1395 53985 1447
rect 53909 1343 53985 1395
rect 53909 1291 53921 1343
rect 53973 1291 53985 1343
rect 53909 1279 53985 1291
rect 53443 828 53489 885
rect 53763 828 53809 885
rect 53123 782 53809 828
rect 52948 -7 53024 5
rect 52948 -59 52960 -7
rect 53012 -59 53024 -7
rect 52948 -111 53024 -59
rect 52948 -163 52960 -111
rect 53012 -163 53024 -111
rect 52948 -175 53024 -163
rect 53123 -232 53169 782
rect 53508 535 53584 547
rect 53508 483 53520 535
rect 53572 532 53584 535
rect 53668 535 53744 547
rect 53668 532 53680 535
rect 53572 483 53680 532
rect 53732 483 53744 535
rect 53508 471 53744 483
rect 53603 399 53649 471
rect 53269 387 53345 399
rect 53269 335 53281 387
rect 53333 335 53345 387
rect 53269 283 53345 335
rect 53269 231 53281 283
rect 53333 231 53345 283
rect 53269 219 53345 231
rect 53909 387 53985 399
rect 53909 335 53921 387
rect 53973 335 53985 387
rect 53909 283 53985 335
rect 53909 231 53921 283
rect 53973 231 53985 283
rect 53909 219 53985 231
rect 53443 -232 53489 -175
rect 53763 -232 53809 -175
rect 53123 -278 53809 -232
rect 52948 -1067 53024 -1055
rect 52948 -1119 52960 -1067
rect 53012 -1119 53024 -1067
rect 52948 -1171 53024 -1119
rect 52948 -1223 52960 -1171
rect 53012 -1223 53024 -1171
rect 52948 -1235 53024 -1223
rect 53123 -1578 53169 -278
rect 53508 -525 53584 -513
rect 53508 -577 53520 -525
rect 53572 -528 53584 -525
rect 53668 -525 53744 -513
rect 53668 -528 53680 -525
rect 53572 -577 53680 -528
rect 53732 -577 53744 -525
rect 53508 -589 53744 -577
rect 53603 -661 53649 -589
rect 53269 -673 53345 -661
rect 53269 -725 53281 -673
rect 53333 -725 53345 -673
rect 53269 -777 53345 -725
rect 53269 -829 53281 -777
rect 53333 -829 53345 -777
rect 53269 -841 53345 -829
rect 53909 -673 53985 -661
rect 53909 -725 53921 -673
rect 53973 -725 53985 -673
rect 53909 -777 53985 -725
rect 53909 -829 53921 -777
rect 53973 -829 53985 -777
rect 53909 -841 53985 -829
rect 53443 -1578 53489 -1235
rect 53763 -1578 53809 -1235
rect 54083 -1578 54129 2862
rect 54228 2113 54304 2125
rect 54228 2061 54240 2113
rect 54292 2061 54304 2113
rect 54228 2009 54304 2061
rect 54228 1957 54240 2009
rect 54292 1957 54304 2009
rect 54228 1945 54304 1957
rect 54228 1053 54304 1065
rect 54228 1001 54240 1053
rect 54292 1001 54304 1053
rect 54228 949 54304 1001
rect 54228 897 54240 949
rect 54292 897 54304 949
rect 54228 885 54304 897
rect 54228 -7 54304 5
rect 54228 -59 54240 -7
rect 54292 -59 54304 -7
rect 54228 -111 54304 -59
rect 54228 -163 54240 -111
rect 54292 -163 54304 -111
rect 54228 -175 54304 -163
rect 54228 -1067 54304 -1055
rect 54228 -1119 54240 -1067
rect 54292 -1119 54304 -1067
rect 54228 -1171 54304 -1119
rect 54228 -1223 54240 -1171
rect 54292 -1223 54304 -1171
rect 54228 -1235 54304 -1223
rect 54403 -1578 54449 2862
rect 54549 2507 54625 2519
rect 54549 2455 54561 2507
rect 54613 2455 54625 2507
rect 54549 2403 54625 2455
rect 54549 2351 54561 2403
rect 54613 2351 54625 2403
rect 54549 2339 54625 2351
rect 54549 1447 54625 1459
rect 54549 1395 54561 1447
rect 54613 1395 54625 1447
rect 54549 1343 54625 1395
rect 54549 1291 54561 1343
rect 54613 1291 54625 1343
rect 54549 1279 54625 1291
rect 54549 387 54625 399
rect 54549 335 54561 387
rect 54613 335 54625 387
rect 54549 283 54625 335
rect 54549 231 54561 283
rect 54613 231 54625 283
rect 54549 219 54625 231
rect 54549 -673 54625 -661
rect 54549 -725 54561 -673
rect 54613 -725 54625 -673
rect 54549 -777 54625 -725
rect 54549 -829 54561 -777
rect 54613 -829 54625 -777
rect 54549 -841 54625 -829
rect 54723 -1578 54769 2862
rect 55011 2519 55057 2862
rect 55171 2519 55217 2862
rect 55516 2828 55671 2862
rect 55717 2862 59807 2874
rect 55717 2828 55872 2862
rect 55516 2780 55872 2828
rect 55516 2734 55671 2780
rect 55717 2734 55872 2780
rect 55516 2686 55872 2734
rect 55516 2640 55671 2686
rect 55717 2640 55872 2686
rect 55516 2592 55872 2640
rect 55516 2546 55671 2592
rect 55717 2546 55872 2592
rect 55516 2498 55872 2546
rect 56171 2519 56217 2862
rect 56331 2519 56377 2862
rect 55516 2452 55671 2498
rect 55717 2452 55872 2498
rect 55516 2404 55872 2452
rect 55516 2358 55671 2404
rect 55717 2358 55872 2404
rect 55516 2310 55872 2358
rect 55516 2264 55671 2310
rect 55717 2264 55872 2310
rect 55516 2216 55872 2264
rect 55516 2170 55671 2216
rect 55717 2170 55872 2216
rect 54868 2113 54944 2125
rect 54868 2061 54880 2113
rect 54932 2061 54944 2113
rect 54868 2009 54944 2061
rect 54868 1957 54880 2009
rect 54932 1957 54944 2009
rect 54868 1945 54944 1957
rect 55516 2122 55872 2170
rect 55516 2076 55671 2122
rect 55717 2076 55872 2122
rect 55516 2028 55872 2076
rect 55516 1982 55671 2028
rect 55717 1982 55872 2028
rect 55011 1725 55057 1945
rect 55171 1725 55217 1945
rect 55011 1679 55091 1725
rect 55137 1679 55217 1725
rect 54868 1053 54944 1065
rect 54868 1001 54880 1053
rect 54932 1001 54944 1053
rect 54868 949 54944 1001
rect 54868 897 54880 949
rect 54932 897 54944 949
rect 54868 885 54944 897
rect 54868 -7 54944 5
rect 54868 -59 54880 -7
rect 54932 -59 54944 -7
rect 54868 -111 54944 -59
rect 54868 -163 54880 -111
rect 54932 -163 54944 -111
rect 54868 -175 54944 -163
rect 55011 -395 55057 1679
rect 55171 -395 55217 1679
rect 55011 -441 55091 -395
rect 55137 -441 55217 -395
rect 54868 -1067 54944 -1055
rect 54868 -1119 54880 -1067
rect 54932 -1119 54944 -1067
rect 54868 -1171 54944 -1119
rect 54868 -1223 54880 -1171
rect 54932 -1223 54944 -1171
rect 54868 -1235 54944 -1223
rect 55011 -1578 55057 -441
rect 55171 -1578 55217 -441
rect 55516 1934 55872 1982
rect 56444 2113 56520 2125
rect 56444 2061 56456 2113
rect 56508 2061 56520 2113
rect 56444 2009 56520 2061
rect 56444 1957 56456 2009
rect 56508 1957 56520 2009
rect 56444 1945 56520 1957
rect 55516 1888 55671 1934
rect 55717 1888 55872 1934
rect 55516 1840 55872 1888
rect 55516 1794 55671 1840
rect 55717 1794 55872 1840
rect 55516 1746 55872 1794
rect 55516 1700 55671 1746
rect 55717 1700 55872 1746
rect 55516 1652 55872 1700
rect 55516 1606 55671 1652
rect 55717 1606 55872 1652
rect 55516 1558 55872 1606
rect 55516 1512 55671 1558
rect 55717 1512 55872 1558
rect 55516 1464 55872 1512
rect 55516 1418 55671 1464
rect 55717 1418 55872 1464
rect 55516 1370 55872 1418
rect 55516 1324 55671 1370
rect 55717 1324 55872 1370
rect 55516 1276 55872 1324
rect 55516 1230 55671 1276
rect 55717 1230 55872 1276
rect 55516 1182 55872 1230
rect 55516 1136 55671 1182
rect 55717 1136 55872 1182
rect 55516 1088 55872 1136
rect 55516 1042 55671 1088
rect 55717 1042 55872 1088
rect 55516 994 55872 1042
rect 55516 948 55671 994
rect 55717 948 55872 994
rect 55516 900 55872 948
rect 55516 854 55671 900
rect 55717 854 55872 900
rect 55516 806 55872 854
rect 55516 760 55671 806
rect 55717 760 55872 806
rect 55516 712 55872 760
rect 55516 666 55671 712
rect 55717 666 55872 712
rect 55516 618 55872 666
rect 55516 572 55671 618
rect 55717 572 55872 618
rect 55516 524 55872 572
rect 55516 478 55671 524
rect 55717 478 55872 524
rect 55516 430 55872 478
rect 55516 384 55671 430
rect 55717 384 55872 430
rect 55516 336 55872 384
rect 55516 290 55671 336
rect 55717 290 55872 336
rect 55516 242 55872 290
rect 55516 196 55671 242
rect 55717 196 55872 242
rect 55516 148 55872 196
rect 55516 102 55671 148
rect 55717 102 55872 148
rect 55516 54 55872 102
rect 55516 8 55671 54
rect 55717 8 55872 54
rect 55516 -40 55872 8
rect 55516 -86 55671 -40
rect 55717 -86 55872 -40
rect 55516 -134 55872 -86
rect 55516 -180 55671 -134
rect 55717 -180 55872 -134
rect 55516 -228 55872 -180
rect 55516 -274 55671 -228
rect 55717 -274 55872 -228
rect 55516 -322 55872 -274
rect 55516 -368 55671 -322
rect 55717 -368 55872 -322
rect 55516 -416 55872 -368
rect 55516 -462 55671 -416
rect 55717 -462 55872 -416
rect 55516 -510 55872 -462
rect 55516 -556 55671 -510
rect 55717 -556 55872 -510
rect 55516 -604 55872 -556
rect 55516 -650 55671 -604
rect 55717 -650 55872 -604
rect 55516 -698 55872 -650
rect 55516 -744 55671 -698
rect 55717 -744 55872 -698
rect 55516 -792 55872 -744
rect 55516 -838 55671 -792
rect 55717 -838 55872 -792
rect 55516 -886 55872 -838
rect 55516 -932 55671 -886
rect 55717 -932 55872 -886
rect 55516 -980 55872 -932
rect 55516 -1026 55671 -980
rect 55717 -1026 55872 -980
rect 55516 -1074 55872 -1026
rect 55516 -1120 55671 -1074
rect 55717 -1120 55872 -1074
rect 55516 -1168 55872 -1120
rect 55516 -1214 55671 -1168
rect 55717 -1214 55872 -1168
rect 55516 -1262 55872 -1214
rect 55516 -1308 55671 -1262
rect 55717 -1308 55872 -1262
rect 55516 -1356 55872 -1308
rect 55516 -1402 55671 -1356
rect 55717 -1402 55872 -1356
rect 55516 -1450 55872 -1402
rect 55516 -1496 55671 -1450
rect 55717 -1496 55872 -1450
rect 55516 -1544 55872 -1496
rect 55516 -1578 55671 -1544
rect 51581 -1590 55671 -1578
rect 55717 -1578 55872 -1544
rect 56171 1725 56217 1945
rect 56331 1725 56377 1945
rect 56171 1679 56251 1725
rect 56297 1679 56377 1725
rect 56171 -395 56217 1679
rect 56331 -395 56377 1679
rect 56444 1053 56520 1065
rect 56444 1001 56456 1053
rect 56508 1001 56520 1053
rect 56444 949 56520 1001
rect 56444 897 56456 949
rect 56508 897 56520 949
rect 56444 885 56520 897
rect 56444 -7 56520 5
rect 56444 -59 56456 -7
rect 56508 -59 56520 -7
rect 56444 -111 56520 -59
rect 56444 -163 56456 -111
rect 56508 -163 56520 -111
rect 56444 -175 56520 -163
rect 56171 -441 56251 -395
rect 56297 -441 56377 -395
rect 56171 -1578 56217 -441
rect 56331 -1578 56377 -441
rect 56444 -1067 56520 -1055
rect 56444 -1119 56456 -1067
rect 56508 -1119 56520 -1067
rect 56444 -1171 56520 -1119
rect 56444 -1223 56456 -1171
rect 56508 -1223 56520 -1171
rect 56444 -1235 56520 -1223
rect 56619 -1578 56665 2862
rect 56763 2507 56839 2519
rect 56763 2455 56775 2507
rect 56827 2455 56839 2507
rect 56763 2403 56839 2455
rect 56763 2351 56775 2403
rect 56827 2351 56839 2403
rect 56763 2339 56839 2351
rect 56763 1447 56839 1459
rect 56763 1395 56775 1447
rect 56827 1395 56839 1447
rect 56763 1343 56839 1395
rect 56763 1291 56775 1343
rect 56827 1291 56839 1343
rect 56763 1279 56839 1291
rect 56763 387 56839 399
rect 56763 335 56775 387
rect 56827 335 56839 387
rect 56763 283 56839 335
rect 56763 231 56775 283
rect 56827 231 56839 283
rect 56763 219 56839 231
rect 56763 -673 56839 -661
rect 56763 -725 56775 -673
rect 56827 -725 56839 -673
rect 56763 -777 56839 -725
rect 56763 -829 56775 -777
rect 56827 -829 56839 -777
rect 56763 -841 56839 -829
rect 56939 -1578 56985 2862
rect 57084 2113 57160 2125
rect 57084 2061 57096 2113
rect 57148 2061 57160 2113
rect 57084 2009 57160 2061
rect 57084 1957 57096 2009
rect 57148 1957 57160 2009
rect 57084 1945 57160 1957
rect 57084 1053 57160 1065
rect 57084 1001 57096 1053
rect 57148 1001 57160 1053
rect 57084 949 57160 1001
rect 57084 897 57096 949
rect 57148 897 57160 949
rect 57084 885 57160 897
rect 57084 -7 57160 5
rect 57084 -59 57096 -7
rect 57148 -59 57160 -7
rect 57084 -111 57160 -59
rect 57084 -163 57096 -111
rect 57148 -163 57160 -111
rect 57084 -175 57160 -163
rect 57084 -1067 57160 -1055
rect 57084 -1119 57096 -1067
rect 57148 -1119 57160 -1067
rect 57084 -1171 57160 -1119
rect 57084 -1223 57096 -1171
rect 57148 -1223 57160 -1171
rect 57084 -1235 57160 -1223
rect 57259 -1578 57305 2862
rect 57644 2655 57720 2667
rect 57644 2603 57656 2655
rect 57708 2652 57720 2655
rect 57804 2655 57880 2667
rect 57804 2652 57816 2655
rect 57708 2603 57816 2652
rect 57868 2603 57880 2655
rect 57644 2591 57880 2603
rect 57739 2519 57785 2591
rect 57403 2507 57479 2519
rect 57403 2455 57415 2507
rect 57467 2455 57479 2507
rect 57403 2403 57479 2455
rect 57403 2351 57415 2403
rect 57467 2351 57479 2403
rect 57403 2339 57479 2351
rect 58043 2507 58119 2519
rect 58043 2455 58055 2507
rect 58107 2455 58119 2507
rect 58043 2403 58119 2455
rect 58043 2351 58055 2403
rect 58107 2351 58119 2403
rect 58043 2339 58119 2351
rect 57579 1888 57625 1945
rect 57899 1888 57945 1945
rect 58219 1888 58265 2862
rect 58364 2113 58440 2125
rect 58364 2061 58376 2113
rect 58428 2061 58440 2113
rect 58364 2009 58440 2061
rect 58364 1957 58376 2009
rect 58428 1957 58440 2009
rect 58364 1945 58440 1957
rect 57579 1842 58265 1888
rect 57644 1595 57720 1607
rect 57644 1543 57656 1595
rect 57708 1592 57720 1595
rect 57804 1595 57880 1607
rect 57804 1592 57816 1595
rect 57708 1543 57816 1592
rect 57868 1543 57880 1595
rect 57644 1531 57880 1543
rect 57739 1459 57785 1531
rect 57403 1447 57479 1459
rect 57403 1395 57415 1447
rect 57467 1395 57479 1447
rect 57403 1343 57479 1395
rect 57403 1291 57415 1343
rect 57467 1291 57479 1343
rect 57403 1279 57479 1291
rect 58043 1447 58119 1459
rect 58043 1395 58055 1447
rect 58107 1395 58119 1447
rect 58043 1343 58119 1395
rect 58043 1291 58055 1343
rect 58107 1291 58119 1343
rect 58043 1279 58119 1291
rect 57579 828 57625 885
rect 57899 828 57945 885
rect 58219 828 58265 1842
rect 58364 1053 58440 1065
rect 58364 1001 58376 1053
rect 58428 1001 58440 1053
rect 58364 949 58440 1001
rect 58364 897 58376 949
rect 58428 897 58440 949
rect 58364 885 58440 897
rect 57579 782 58265 828
rect 57644 535 57720 547
rect 57644 483 57656 535
rect 57708 532 57720 535
rect 57804 535 57880 547
rect 57804 532 57816 535
rect 57708 483 57816 532
rect 57868 483 57880 535
rect 57644 471 57880 483
rect 57739 399 57785 471
rect 57403 387 57479 399
rect 57403 335 57415 387
rect 57467 335 57479 387
rect 57403 283 57479 335
rect 57403 231 57415 283
rect 57467 231 57479 283
rect 57403 219 57479 231
rect 58043 387 58119 399
rect 58043 335 58055 387
rect 58107 335 58119 387
rect 58043 283 58119 335
rect 58043 231 58055 283
rect 58107 231 58119 283
rect 58043 219 58119 231
rect 57579 -232 57625 -175
rect 57899 -232 57945 -175
rect 58219 -232 58265 782
rect 58364 -7 58440 5
rect 58364 -59 58376 -7
rect 58428 -59 58440 -7
rect 58364 -111 58440 -59
rect 58364 -163 58376 -111
rect 58428 -163 58440 -111
rect 58364 -175 58440 -163
rect 57579 -278 58265 -232
rect 57644 -525 57720 -513
rect 57644 -577 57656 -525
rect 57708 -528 57720 -525
rect 57804 -525 57880 -513
rect 57804 -528 57816 -525
rect 57708 -577 57816 -528
rect 57868 -577 57880 -525
rect 57644 -589 57880 -577
rect 57739 -661 57785 -589
rect 57403 -673 57479 -661
rect 57403 -725 57415 -673
rect 57467 -725 57479 -673
rect 57403 -777 57479 -725
rect 57403 -829 57415 -777
rect 57467 -829 57479 -777
rect 57403 -841 57479 -829
rect 58043 -673 58119 -661
rect 58043 -725 58055 -673
rect 58107 -725 58119 -673
rect 58043 -777 58119 -725
rect 58043 -829 58055 -777
rect 58107 -829 58119 -777
rect 58043 -841 58119 -829
rect 57579 -1578 57625 -1235
rect 57899 -1578 57945 -1235
rect 58219 -1578 58265 -278
rect 58364 -1067 58440 -1055
rect 58364 -1119 58376 -1067
rect 58428 -1119 58440 -1067
rect 58364 -1171 58440 -1119
rect 58364 -1223 58376 -1171
rect 58428 -1223 58440 -1171
rect 58364 -1235 58440 -1223
rect 58539 -1578 58585 2862
rect 58683 2507 58759 2519
rect 58683 2455 58695 2507
rect 58747 2455 58759 2507
rect 58683 2403 58759 2455
rect 58683 2351 58695 2403
rect 58747 2351 58759 2403
rect 58683 2339 58759 2351
rect 58683 1447 58759 1459
rect 58683 1395 58695 1447
rect 58747 1395 58759 1447
rect 58683 1343 58759 1395
rect 58683 1291 58695 1343
rect 58747 1291 58759 1343
rect 58683 1279 58759 1291
rect 58683 387 58759 399
rect 58683 335 58695 387
rect 58747 335 58759 387
rect 58683 283 58759 335
rect 58683 231 58695 283
rect 58747 231 58759 283
rect 58683 219 58759 231
rect 58683 -673 58759 -661
rect 58683 -725 58695 -673
rect 58747 -725 58759 -673
rect 58683 -777 58759 -725
rect 58683 -829 58695 -777
rect 58747 -829 58759 -777
rect 58683 -841 58759 -829
rect 58859 -1578 58905 2862
rect 59147 2519 59193 2862
rect 59307 2519 59353 2862
rect 59652 2828 59807 2862
rect 59853 2862 61231 2874
rect 59853 2828 59972 2862
rect 59652 2780 59972 2828
rect 59652 2734 59807 2780
rect 59853 2734 59972 2780
rect 59652 2686 59972 2734
rect 59652 2640 59807 2686
rect 59853 2640 59972 2686
rect 59652 2592 59972 2640
rect 59652 2546 59807 2592
rect 59853 2546 59972 2592
rect 59652 2498 59972 2546
rect 59652 2452 59807 2498
rect 59853 2452 59972 2498
rect 59652 2404 59972 2452
rect 59652 2358 59807 2404
rect 59853 2358 59972 2404
rect 59652 2310 59972 2358
rect 59652 2264 59807 2310
rect 59853 2264 59972 2310
rect 59652 2216 59972 2264
rect 59652 2170 59807 2216
rect 59853 2170 59972 2216
rect 59004 2113 59080 2125
rect 59004 2061 59016 2113
rect 59068 2061 59080 2113
rect 59004 2009 59080 2061
rect 59004 1957 59016 2009
rect 59068 1957 59080 2009
rect 59004 1945 59080 1957
rect 59652 2122 59972 2170
rect 59652 2076 59807 2122
rect 59853 2076 59972 2122
rect 59652 2028 59972 2076
rect 59652 1982 59807 2028
rect 59853 1982 59972 2028
rect 59147 1725 59193 1945
rect 59307 1725 59353 1945
rect 59147 1679 59227 1725
rect 59273 1679 59353 1725
rect 59004 1053 59080 1065
rect 59004 1001 59016 1053
rect 59068 1001 59080 1053
rect 59004 949 59080 1001
rect 59004 897 59016 949
rect 59068 897 59080 949
rect 59004 885 59080 897
rect 59004 -7 59080 5
rect 59004 -59 59016 -7
rect 59068 -59 59080 -7
rect 59004 -111 59080 -59
rect 59004 -163 59016 -111
rect 59068 -163 59080 -111
rect 59004 -175 59080 -163
rect 59147 -395 59193 1679
rect 59307 -395 59353 1679
rect 59147 -441 59227 -395
rect 59273 -441 59353 -395
rect 59004 -1067 59080 -1055
rect 59004 -1119 59016 -1067
rect 59068 -1119 59080 -1067
rect 59004 -1171 59080 -1119
rect 59004 -1223 59016 -1171
rect 59068 -1223 59080 -1171
rect 59004 -1235 59080 -1223
rect 59147 -1578 59193 -441
rect 59307 -1578 59353 -441
rect 59652 1934 59972 1982
rect 59652 1888 59807 1934
rect 59853 1888 59972 1934
rect 59652 1840 59972 1888
rect 59652 1794 59807 1840
rect 59853 1794 59972 1840
rect 59652 1746 59972 1794
rect 59652 1700 59807 1746
rect 59853 1700 59972 1746
rect 59652 1652 59972 1700
rect 59652 1606 59807 1652
rect 59853 1606 59972 1652
rect 59652 1558 59972 1606
rect 59652 1512 59807 1558
rect 59853 1512 59972 1558
rect 59652 1464 59972 1512
rect 59652 1418 59807 1464
rect 59853 1418 59972 1464
rect 59652 1370 59972 1418
rect 59652 1324 59807 1370
rect 59853 1324 59972 1370
rect 59652 1276 59972 1324
rect 59652 1230 59807 1276
rect 59853 1230 59972 1276
rect 59652 1182 59972 1230
rect 59652 1136 59807 1182
rect 59853 1136 59972 1182
rect 59652 1088 59972 1136
rect 59652 1042 59807 1088
rect 59853 1042 59972 1088
rect 59652 994 59972 1042
rect 59652 948 59807 994
rect 59853 948 59972 994
rect 59652 900 59972 948
rect 59652 854 59807 900
rect 59853 854 59972 900
rect 59652 806 59972 854
rect 59652 760 59807 806
rect 59853 760 59972 806
rect 59652 712 59972 760
rect 59652 666 59807 712
rect 59853 666 59972 712
rect 59652 618 59972 666
rect 59652 572 59807 618
rect 59853 572 59972 618
rect 59652 524 59972 572
rect 59652 478 59807 524
rect 59853 478 59972 524
rect 59652 430 59972 478
rect 59652 384 59807 430
rect 59853 384 59972 430
rect 59652 336 59972 384
rect 59652 290 59807 336
rect 59853 290 59972 336
rect 59652 242 59972 290
rect 59652 196 59807 242
rect 59853 196 59972 242
rect 59652 148 59972 196
rect 59652 102 59807 148
rect 59853 102 59972 148
rect 59652 54 59972 102
rect 59652 8 59807 54
rect 59853 8 59972 54
rect 59652 -40 59972 8
rect 59652 -86 59807 -40
rect 59853 -86 59972 -40
rect 59652 -134 59972 -86
rect 59652 -180 59807 -134
rect 59853 -180 59972 -134
rect 59652 -228 59972 -180
rect 59652 -274 59807 -228
rect 59853 -274 59972 -228
rect 59652 -322 59972 -274
rect 59652 -368 59807 -322
rect 59853 -368 59972 -322
rect 59652 -416 59972 -368
rect 59652 -462 59807 -416
rect 59853 -462 59972 -416
rect 59652 -510 59972 -462
rect 59652 -556 59807 -510
rect 59853 -556 59972 -510
rect 59652 -604 59972 -556
rect 59652 -650 59807 -604
rect 59853 -650 59972 -604
rect 59652 -698 59972 -650
rect 59652 -744 59807 -698
rect 59853 -744 59972 -698
rect 59652 -792 59972 -744
rect 59652 -838 59807 -792
rect 59853 -838 59972 -792
rect 59652 -886 59972 -838
rect 59652 -932 59807 -886
rect 59853 -932 59972 -886
rect 59652 -980 59972 -932
rect 59652 -1026 59807 -980
rect 59853 -1026 59972 -980
rect 59652 -1074 59972 -1026
rect 59652 -1120 59807 -1074
rect 59853 -1120 59972 -1074
rect 59652 -1168 59972 -1120
rect 59652 -1214 59807 -1168
rect 59853 -1214 59972 -1168
rect 59652 -1262 59972 -1214
rect 59652 -1308 59807 -1262
rect 59853 -1308 59972 -1262
rect 59652 -1356 59972 -1308
rect 59652 -1402 59807 -1356
rect 59853 -1402 59972 -1356
rect 59652 -1450 59972 -1402
rect 59652 -1496 59807 -1450
rect 59853 -1496 59972 -1450
rect 59652 -1544 59972 -1496
rect 59652 -1578 59807 -1544
rect 55717 -1590 59807 -1578
rect 59853 -1578 59972 -1544
rect 61112 2828 61231 2862
rect 61277 2862 65367 2874
rect 61277 2828 61432 2862
rect 61112 2780 61432 2828
rect 61112 2734 61231 2780
rect 61277 2734 61432 2780
rect 61112 2686 61432 2734
rect 61112 2640 61231 2686
rect 61277 2640 61432 2686
rect 61112 2592 61432 2640
rect 61112 2546 61231 2592
rect 61277 2546 61432 2592
rect 61112 2498 61432 2546
rect 61731 2519 61777 2862
rect 61891 2519 61937 2862
rect 61112 2452 61231 2498
rect 61277 2452 61432 2498
rect 61112 2404 61432 2452
rect 61112 2358 61231 2404
rect 61277 2358 61432 2404
rect 61112 2310 61432 2358
rect 61112 2264 61231 2310
rect 61277 2264 61432 2310
rect 61112 2216 61432 2264
rect 61112 2170 61231 2216
rect 61277 2170 61432 2216
rect 61112 2122 61432 2170
rect 61112 2076 61231 2122
rect 61277 2076 61432 2122
rect 61112 2028 61432 2076
rect 61112 1982 61231 2028
rect 61277 1982 61432 2028
rect 61112 1934 61432 1982
rect 62004 2113 62080 2125
rect 62004 2061 62016 2113
rect 62068 2061 62080 2113
rect 62004 2009 62080 2061
rect 62004 1957 62016 2009
rect 62068 1957 62080 2009
rect 62004 1945 62080 1957
rect 61112 1888 61231 1934
rect 61277 1888 61432 1934
rect 61112 1840 61432 1888
rect 61112 1794 61231 1840
rect 61277 1794 61432 1840
rect 61112 1746 61432 1794
rect 61112 1700 61231 1746
rect 61277 1700 61432 1746
rect 61112 1652 61432 1700
rect 61112 1606 61231 1652
rect 61277 1606 61432 1652
rect 61112 1558 61432 1606
rect 61112 1512 61231 1558
rect 61277 1512 61432 1558
rect 61112 1464 61432 1512
rect 61112 1418 61231 1464
rect 61277 1418 61432 1464
rect 61112 1370 61432 1418
rect 61112 1324 61231 1370
rect 61277 1324 61432 1370
rect 61112 1276 61432 1324
rect 61112 1230 61231 1276
rect 61277 1230 61432 1276
rect 61112 1182 61432 1230
rect 61112 1136 61231 1182
rect 61277 1136 61432 1182
rect 61112 1088 61432 1136
rect 61112 1042 61231 1088
rect 61277 1042 61432 1088
rect 61112 994 61432 1042
rect 61112 948 61231 994
rect 61277 948 61432 994
rect 61112 900 61432 948
rect 61112 854 61231 900
rect 61277 854 61432 900
rect 61112 806 61432 854
rect 61112 760 61231 806
rect 61277 760 61432 806
rect 61112 712 61432 760
rect 61112 666 61231 712
rect 61277 666 61432 712
rect 61112 618 61432 666
rect 61112 572 61231 618
rect 61277 572 61432 618
rect 61112 524 61432 572
rect 61112 478 61231 524
rect 61277 478 61432 524
rect 61112 430 61432 478
rect 61112 384 61231 430
rect 61277 384 61432 430
rect 61112 336 61432 384
rect 61112 290 61231 336
rect 61277 290 61432 336
rect 61112 242 61432 290
rect 61112 196 61231 242
rect 61277 196 61432 242
rect 61112 148 61432 196
rect 61112 102 61231 148
rect 61277 102 61432 148
rect 61112 54 61432 102
rect 61112 8 61231 54
rect 61277 8 61432 54
rect 61112 -40 61432 8
rect 61112 -86 61231 -40
rect 61277 -86 61432 -40
rect 61112 -134 61432 -86
rect 61112 -180 61231 -134
rect 61277 -180 61432 -134
rect 61112 -228 61432 -180
rect 61112 -274 61231 -228
rect 61277 -274 61432 -228
rect 61112 -322 61432 -274
rect 61112 -368 61231 -322
rect 61277 -368 61432 -322
rect 61112 -416 61432 -368
rect 61112 -462 61231 -416
rect 61277 -462 61432 -416
rect 61112 -510 61432 -462
rect 61112 -556 61231 -510
rect 61277 -556 61432 -510
rect 61112 -604 61432 -556
rect 61112 -650 61231 -604
rect 61277 -650 61432 -604
rect 61112 -698 61432 -650
rect 61112 -744 61231 -698
rect 61277 -744 61432 -698
rect 61112 -792 61432 -744
rect 61112 -838 61231 -792
rect 61277 -838 61432 -792
rect 61112 -886 61432 -838
rect 61112 -932 61231 -886
rect 61277 -932 61432 -886
rect 61112 -980 61432 -932
rect 61112 -1026 61231 -980
rect 61277 -1026 61432 -980
rect 61112 -1074 61432 -1026
rect 61112 -1120 61231 -1074
rect 61277 -1120 61432 -1074
rect 61112 -1168 61432 -1120
rect 61112 -1214 61231 -1168
rect 61277 -1214 61432 -1168
rect 61112 -1262 61432 -1214
rect 61112 -1308 61231 -1262
rect 61277 -1308 61432 -1262
rect 61112 -1356 61432 -1308
rect 61112 -1402 61231 -1356
rect 61277 -1402 61432 -1356
rect 61112 -1450 61432 -1402
rect 61112 -1496 61231 -1450
rect 61277 -1496 61432 -1450
rect 61112 -1544 61432 -1496
rect 61112 -1578 61231 -1544
rect 59853 -1590 61231 -1578
rect 61277 -1578 61432 -1544
rect 61731 1725 61777 1945
rect 61891 1725 61937 1945
rect 61731 1679 61811 1725
rect 61857 1679 61937 1725
rect 61731 -395 61777 1679
rect 61891 -395 61937 1679
rect 62004 1053 62080 1065
rect 62004 1001 62016 1053
rect 62068 1001 62080 1053
rect 62004 949 62080 1001
rect 62004 897 62016 949
rect 62068 897 62080 949
rect 62004 885 62080 897
rect 62004 -7 62080 5
rect 62004 -59 62016 -7
rect 62068 -59 62080 -7
rect 62004 -111 62080 -59
rect 62004 -163 62016 -111
rect 62068 -163 62080 -111
rect 62004 -175 62080 -163
rect 61731 -441 61811 -395
rect 61857 -441 61937 -395
rect 61731 -1578 61777 -441
rect 61891 -1578 61937 -441
rect 62004 -1067 62080 -1055
rect 62004 -1119 62016 -1067
rect 62068 -1119 62080 -1067
rect 62004 -1171 62080 -1119
rect 62004 -1223 62016 -1171
rect 62068 -1223 62080 -1171
rect 62004 -1235 62080 -1223
rect 62179 -1578 62225 2862
rect 62325 2507 62401 2519
rect 62325 2455 62337 2507
rect 62389 2455 62401 2507
rect 62325 2403 62401 2455
rect 62325 2351 62337 2403
rect 62389 2351 62401 2403
rect 62325 2339 62401 2351
rect 62325 1447 62401 1459
rect 62325 1395 62337 1447
rect 62389 1395 62401 1447
rect 62325 1343 62401 1395
rect 62325 1291 62337 1343
rect 62389 1291 62401 1343
rect 62325 1279 62401 1291
rect 62325 387 62401 399
rect 62325 335 62337 387
rect 62389 335 62401 387
rect 62325 283 62401 335
rect 62325 231 62337 283
rect 62389 231 62401 283
rect 62325 219 62401 231
rect 62325 -673 62401 -661
rect 62325 -725 62337 -673
rect 62389 -725 62401 -673
rect 62325 -777 62401 -725
rect 62325 -829 62337 -777
rect 62389 -829 62401 -777
rect 62325 -841 62401 -829
rect 62499 -1578 62545 2862
rect 62644 2113 62720 2125
rect 62644 2061 62656 2113
rect 62708 2061 62720 2113
rect 62644 2009 62720 2061
rect 62644 1957 62656 2009
rect 62708 1957 62720 2009
rect 62644 1945 62720 1957
rect 62819 1888 62865 2862
rect 63204 2655 63280 2667
rect 63204 2603 63216 2655
rect 63268 2652 63280 2655
rect 63364 2655 63440 2667
rect 63364 2652 63376 2655
rect 63268 2603 63376 2652
rect 63428 2603 63440 2655
rect 63204 2591 63440 2603
rect 63299 2519 63345 2591
rect 62965 2507 63041 2519
rect 62965 2455 62977 2507
rect 63029 2455 63041 2507
rect 62965 2403 63041 2455
rect 62965 2351 62977 2403
rect 63029 2351 63041 2403
rect 62965 2339 63041 2351
rect 63605 2507 63681 2519
rect 63605 2455 63617 2507
rect 63669 2455 63681 2507
rect 63605 2403 63681 2455
rect 63605 2351 63617 2403
rect 63669 2351 63681 2403
rect 63605 2339 63681 2351
rect 63139 1888 63185 1945
rect 63459 1888 63505 1945
rect 62819 1842 63505 1888
rect 62644 1053 62720 1065
rect 62644 1001 62656 1053
rect 62708 1001 62720 1053
rect 62644 949 62720 1001
rect 62644 897 62656 949
rect 62708 897 62720 949
rect 62644 885 62720 897
rect 62819 828 62865 1842
rect 63204 1595 63280 1607
rect 63204 1543 63216 1595
rect 63268 1592 63280 1595
rect 63364 1595 63440 1607
rect 63364 1592 63376 1595
rect 63268 1543 63376 1592
rect 63428 1543 63440 1595
rect 63204 1531 63440 1543
rect 63299 1459 63345 1531
rect 62965 1447 63041 1459
rect 62965 1395 62977 1447
rect 63029 1395 63041 1447
rect 62965 1343 63041 1395
rect 62965 1291 62977 1343
rect 63029 1291 63041 1343
rect 62965 1279 63041 1291
rect 63605 1447 63681 1459
rect 63605 1395 63617 1447
rect 63669 1395 63681 1447
rect 63605 1343 63681 1395
rect 63605 1291 63617 1343
rect 63669 1291 63681 1343
rect 63605 1279 63681 1291
rect 63139 828 63185 885
rect 63459 828 63505 885
rect 62819 782 63505 828
rect 62644 -7 62720 5
rect 62644 -59 62656 -7
rect 62708 -59 62720 -7
rect 62644 -111 62720 -59
rect 62644 -163 62656 -111
rect 62708 -163 62720 -111
rect 62644 -175 62720 -163
rect 62819 -232 62865 782
rect 63204 535 63280 547
rect 63204 483 63216 535
rect 63268 532 63280 535
rect 63364 535 63440 547
rect 63364 532 63376 535
rect 63268 483 63376 532
rect 63428 483 63440 535
rect 63204 471 63440 483
rect 63299 399 63345 471
rect 62965 387 63041 399
rect 62965 335 62977 387
rect 63029 335 63041 387
rect 62965 283 63041 335
rect 62965 231 62977 283
rect 63029 231 63041 283
rect 62965 219 63041 231
rect 63605 387 63681 399
rect 63605 335 63617 387
rect 63669 335 63681 387
rect 63605 283 63681 335
rect 63605 231 63617 283
rect 63669 231 63681 283
rect 63605 219 63681 231
rect 63139 -232 63185 -175
rect 63459 -232 63505 -175
rect 62819 -278 63505 -232
rect 62644 -1067 62720 -1055
rect 62644 -1119 62656 -1067
rect 62708 -1119 62720 -1067
rect 62644 -1171 62720 -1119
rect 62644 -1223 62656 -1171
rect 62708 -1223 62720 -1171
rect 62644 -1235 62720 -1223
rect 62819 -1578 62865 -278
rect 63204 -525 63280 -513
rect 63204 -577 63216 -525
rect 63268 -528 63280 -525
rect 63364 -525 63440 -513
rect 63364 -528 63376 -525
rect 63268 -577 63376 -528
rect 63428 -577 63440 -525
rect 63204 -589 63440 -577
rect 63299 -661 63345 -589
rect 62965 -673 63041 -661
rect 62965 -725 62977 -673
rect 63029 -725 63041 -673
rect 62965 -777 63041 -725
rect 62965 -829 62977 -777
rect 63029 -829 63041 -777
rect 62965 -841 63041 -829
rect 63605 -673 63681 -661
rect 63605 -725 63617 -673
rect 63669 -725 63681 -673
rect 63605 -777 63681 -725
rect 63605 -829 63617 -777
rect 63669 -829 63681 -777
rect 63605 -841 63681 -829
rect 63139 -1578 63185 -1235
rect 63459 -1578 63505 -1235
rect 63779 -1578 63825 2862
rect 63924 2113 64000 2125
rect 63924 2061 63936 2113
rect 63988 2061 64000 2113
rect 63924 2009 64000 2061
rect 63924 1957 63936 2009
rect 63988 1957 64000 2009
rect 63924 1945 64000 1957
rect 63924 1053 64000 1065
rect 63924 1001 63936 1053
rect 63988 1001 64000 1053
rect 63924 949 64000 1001
rect 63924 897 63936 949
rect 63988 897 64000 949
rect 63924 885 64000 897
rect 63924 -7 64000 5
rect 63924 -59 63936 -7
rect 63988 -59 64000 -7
rect 63924 -111 64000 -59
rect 63924 -163 63936 -111
rect 63988 -163 64000 -111
rect 63924 -175 64000 -163
rect 63924 -1067 64000 -1055
rect 63924 -1119 63936 -1067
rect 63988 -1119 64000 -1067
rect 63924 -1171 64000 -1119
rect 63924 -1223 63936 -1171
rect 63988 -1223 64000 -1171
rect 63924 -1235 64000 -1223
rect 64099 -1578 64145 2862
rect 64245 2507 64321 2519
rect 64245 2455 64257 2507
rect 64309 2455 64321 2507
rect 64245 2403 64321 2455
rect 64245 2351 64257 2403
rect 64309 2351 64321 2403
rect 64245 2339 64321 2351
rect 64245 1447 64321 1459
rect 64245 1395 64257 1447
rect 64309 1395 64321 1447
rect 64245 1343 64321 1395
rect 64245 1291 64257 1343
rect 64309 1291 64321 1343
rect 64245 1279 64321 1291
rect 64245 387 64321 399
rect 64245 335 64257 387
rect 64309 335 64321 387
rect 64245 283 64321 335
rect 64245 231 64257 283
rect 64309 231 64321 283
rect 64245 219 64321 231
rect 64245 -673 64321 -661
rect 64245 -725 64257 -673
rect 64309 -725 64321 -673
rect 64245 -777 64321 -725
rect 64245 -829 64257 -777
rect 64309 -829 64321 -777
rect 64245 -841 64321 -829
rect 64419 -1578 64465 2862
rect 64707 2519 64753 2862
rect 64867 2519 64913 2862
rect 65212 2828 65367 2862
rect 65413 2828 65532 2874
rect 65212 2780 65532 2828
rect 65212 2734 65367 2780
rect 65413 2734 65532 2780
rect 65212 2686 65532 2734
rect 65212 2640 65367 2686
rect 65413 2640 65532 2686
rect 65212 2592 65532 2640
rect 65212 2546 65367 2592
rect 65413 2546 65532 2592
rect 65212 2498 65532 2546
rect 65212 2452 65367 2498
rect 65413 2452 65532 2498
rect 65212 2404 65532 2452
rect 65212 2358 65367 2404
rect 65413 2358 65532 2404
rect 65212 2310 65532 2358
rect 65212 2264 65367 2310
rect 65413 2264 65532 2310
rect 65212 2216 65532 2264
rect 65212 2170 65367 2216
rect 65413 2170 65532 2216
rect 64564 2113 64640 2125
rect 64564 2061 64576 2113
rect 64628 2061 64640 2113
rect 64564 2009 64640 2061
rect 64564 1957 64576 2009
rect 64628 1957 64640 2009
rect 64564 1945 64640 1957
rect 65212 2122 65532 2170
rect 65212 2076 65367 2122
rect 65413 2076 65532 2122
rect 65212 2028 65532 2076
rect 65212 1982 65367 2028
rect 65413 1982 65532 2028
rect 64707 1725 64753 1945
rect 64867 1725 64913 1945
rect 64707 1679 64787 1725
rect 64833 1679 64913 1725
rect 64564 1053 64640 1065
rect 64564 1001 64576 1053
rect 64628 1001 64640 1053
rect 64564 949 64640 1001
rect 64564 897 64576 949
rect 64628 897 64640 949
rect 64564 885 64640 897
rect 64564 -7 64640 5
rect 64564 -59 64576 -7
rect 64628 -59 64640 -7
rect 64564 -111 64640 -59
rect 64564 -163 64576 -111
rect 64628 -163 64640 -111
rect 64564 -175 64640 -163
rect 64707 -395 64753 1679
rect 64867 -395 64913 1679
rect 64707 -441 64787 -395
rect 64833 -441 64913 -395
rect 64564 -1067 64640 -1055
rect 64564 -1119 64576 -1067
rect 64628 -1119 64640 -1067
rect 64564 -1171 64640 -1119
rect 64564 -1223 64576 -1171
rect 64628 -1223 64640 -1171
rect 64564 -1235 64640 -1223
rect 64707 -1578 64753 -441
rect 64867 -1578 64913 -441
rect 65212 1934 65532 1982
rect 65212 1888 65367 1934
rect 65413 1888 65532 1934
rect 65212 1840 65532 1888
rect 65212 1794 65367 1840
rect 65413 1794 65532 1840
rect 65212 1746 65532 1794
rect 65212 1700 65367 1746
rect 65413 1700 65532 1746
rect 65212 1652 65532 1700
rect 65212 1606 65367 1652
rect 65413 1606 65532 1652
rect 65212 1558 65532 1606
rect 65212 1512 65367 1558
rect 65413 1512 65532 1558
rect 65212 1464 65532 1512
rect 65212 1418 65367 1464
rect 65413 1418 65532 1464
rect 65212 1370 65532 1418
rect 65212 1324 65367 1370
rect 65413 1324 65532 1370
rect 65212 1276 65532 1324
rect 65212 1230 65367 1276
rect 65413 1230 65532 1276
rect 65212 1182 65532 1230
rect 65212 1136 65367 1182
rect 65413 1136 65532 1182
rect 65212 1088 65532 1136
rect 65212 1042 65367 1088
rect 65413 1042 65532 1088
rect 65212 994 65532 1042
rect 65212 948 65367 994
rect 65413 948 65532 994
rect 65212 900 65532 948
rect 65212 854 65367 900
rect 65413 854 65532 900
rect 65212 806 65532 854
rect 65212 760 65367 806
rect 65413 760 65532 806
rect 65212 712 65532 760
rect 65212 666 65367 712
rect 65413 666 65532 712
rect 65212 618 65532 666
rect 65212 572 65367 618
rect 65413 572 65532 618
rect 65212 524 65532 572
rect 65212 478 65367 524
rect 65413 478 65532 524
rect 65212 430 65532 478
rect 65212 384 65367 430
rect 65413 384 65532 430
rect 65212 336 65532 384
rect 65212 290 65367 336
rect 65413 290 65532 336
rect 65212 242 65532 290
rect 65212 196 65367 242
rect 65413 196 65532 242
rect 65212 148 65532 196
rect 65212 102 65367 148
rect 65413 102 65532 148
rect 65212 54 65532 102
rect 65212 8 65367 54
rect 65413 8 65532 54
rect 65212 -40 65532 8
rect 65212 -86 65367 -40
rect 65413 -86 65532 -40
rect 65212 -134 65532 -86
rect 65212 -180 65367 -134
rect 65413 -180 65532 -134
rect 65212 -228 65532 -180
rect 65212 -274 65367 -228
rect 65413 -274 65532 -228
rect 65212 -322 65532 -274
rect 65212 -368 65367 -322
rect 65413 -368 65532 -322
rect 65212 -416 65532 -368
rect 65212 -462 65367 -416
rect 65413 -462 65532 -416
rect 65212 -510 65532 -462
rect 65212 -556 65367 -510
rect 65413 -556 65532 -510
rect 65212 -604 65532 -556
rect 65212 -650 65367 -604
rect 65413 -650 65532 -604
rect 65212 -698 65532 -650
rect 65212 -744 65367 -698
rect 65413 -744 65532 -698
rect 65212 -792 65532 -744
rect 65212 -838 65367 -792
rect 65413 -838 65532 -792
rect 65212 -886 65532 -838
rect 65212 -932 65367 -886
rect 65413 -932 65532 -886
rect 65212 -980 65532 -932
rect 65212 -1026 65367 -980
rect 65413 -1026 65532 -980
rect 65212 -1074 65532 -1026
rect 65212 -1120 65367 -1074
rect 65413 -1120 65532 -1074
rect 65212 -1168 65532 -1120
rect 65212 -1214 65367 -1168
rect 65413 -1214 65532 -1168
rect 65212 -1262 65532 -1214
rect 65212 -1308 65367 -1262
rect 65413 -1308 65532 -1262
rect 65212 -1356 65532 -1308
rect 65212 -1402 65367 -1356
rect 65413 -1402 65532 -1356
rect 65212 -1450 65532 -1402
rect 65212 -1496 65367 -1450
rect 65413 -1496 65532 -1450
rect 65212 -1544 65532 -1496
rect 65212 -1578 65367 -1544
rect 61277 -1590 65367 -1578
rect 65413 -1590 65532 -1544
rect 32024 -1638 65532 -1590
rect 32024 -1684 32143 -1638
rect 32189 -1684 36279 -1638
rect 36325 -1684 40415 -1638
rect 40461 -1684 41839 -1638
rect 41885 -1684 45975 -1638
rect 46021 -1684 50111 -1638
rect 50157 -1684 51535 -1638
rect 51581 -1684 55671 -1638
rect 55717 -1684 59807 -1638
rect 59853 -1684 61231 -1638
rect 61277 -1684 65367 -1638
rect 65413 -1684 65532 -1638
rect 32024 -1732 65532 -1684
rect 32024 -1778 32143 -1732
rect 32189 -1778 32237 -1732
rect 32283 -1778 32331 -1732
rect 32377 -1778 32425 -1732
rect 32471 -1778 32519 -1732
rect 32565 -1778 32613 -1732
rect 32659 -1778 32707 -1732
rect 32753 -1778 32801 -1732
rect 32847 -1778 32895 -1732
rect 32941 -1778 32989 -1732
rect 33035 -1778 33083 -1732
rect 33129 -1778 33177 -1732
rect 33223 -1778 33271 -1732
rect 33317 -1778 33365 -1732
rect 33411 -1778 33459 -1732
rect 33505 -1778 33553 -1732
rect 33599 -1778 33647 -1732
rect 33693 -1778 33741 -1732
rect 33787 -1778 33835 -1732
rect 33881 -1778 33929 -1732
rect 33975 -1778 34023 -1732
rect 34069 -1778 34117 -1732
rect 34163 -1778 34211 -1732
rect 34257 -1778 34305 -1732
rect 34351 -1778 34399 -1732
rect 34445 -1778 34493 -1732
rect 34539 -1778 34587 -1732
rect 34633 -1778 34681 -1732
rect 34727 -1778 34775 -1732
rect 34821 -1778 34869 -1732
rect 34915 -1778 34963 -1732
rect 35009 -1778 35057 -1732
rect 35103 -1778 35151 -1732
rect 35197 -1778 35245 -1732
rect 35291 -1778 35339 -1732
rect 35385 -1778 35433 -1732
rect 35479 -1778 35527 -1732
rect 35573 -1778 35621 -1732
rect 35667 -1778 35715 -1732
rect 35761 -1778 35809 -1732
rect 35855 -1778 35903 -1732
rect 35949 -1778 35997 -1732
rect 36043 -1778 36091 -1732
rect 36137 -1778 36185 -1732
rect 36231 -1778 36279 -1732
rect 36325 -1778 36373 -1732
rect 36419 -1778 36467 -1732
rect 36513 -1778 36561 -1732
rect 36607 -1778 36655 -1732
rect 36701 -1778 36749 -1732
rect 36795 -1778 36843 -1732
rect 36889 -1778 36937 -1732
rect 36983 -1778 37031 -1732
rect 37077 -1778 37125 -1732
rect 37171 -1778 37219 -1732
rect 37265 -1778 37313 -1732
rect 37359 -1778 37407 -1732
rect 37453 -1778 37501 -1732
rect 37547 -1778 37595 -1732
rect 37641 -1778 37689 -1732
rect 37735 -1778 37783 -1732
rect 37829 -1778 37877 -1732
rect 37923 -1778 37971 -1732
rect 38017 -1778 38065 -1732
rect 38111 -1778 38159 -1732
rect 38205 -1778 38253 -1732
rect 38299 -1778 38347 -1732
rect 38393 -1778 38441 -1732
rect 38487 -1778 38535 -1732
rect 38581 -1778 38629 -1732
rect 38675 -1778 38723 -1732
rect 38769 -1778 38817 -1732
rect 38863 -1778 38911 -1732
rect 38957 -1778 39005 -1732
rect 39051 -1778 39099 -1732
rect 39145 -1778 39193 -1732
rect 39239 -1778 39287 -1732
rect 39333 -1778 39381 -1732
rect 39427 -1778 39475 -1732
rect 39521 -1778 39569 -1732
rect 39615 -1778 39663 -1732
rect 39709 -1778 39757 -1732
rect 39803 -1778 39851 -1732
rect 39897 -1778 39945 -1732
rect 39991 -1778 40039 -1732
rect 40085 -1778 40133 -1732
rect 40179 -1778 40227 -1732
rect 40273 -1778 40321 -1732
rect 40367 -1778 40415 -1732
rect 40461 -1778 41839 -1732
rect 41885 -1778 41933 -1732
rect 41979 -1778 42027 -1732
rect 42073 -1778 42121 -1732
rect 42167 -1778 42215 -1732
rect 42261 -1778 42309 -1732
rect 42355 -1778 42403 -1732
rect 42449 -1778 42497 -1732
rect 42543 -1778 42591 -1732
rect 42637 -1778 42685 -1732
rect 42731 -1778 42779 -1732
rect 42825 -1778 42873 -1732
rect 42919 -1778 42967 -1732
rect 43013 -1778 43061 -1732
rect 43107 -1778 43155 -1732
rect 43201 -1778 43249 -1732
rect 43295 -1778 43343 -1732
rect 43389 -1778 43437 -1732
rect 43483 -1778 43531 -1732
rect 43577 -1778 43625 -1732
rect 43671 -1778 43719 -1732
rect 43765 -1778 43813 -1732
rect 43859 -1778 43907 -1732
rect 43953 -1778 44001 -1732
rect 44047 -1778 44095 -1732
rect 44141 -1778 44189 -1732
rect 44235 -1778 44283 -1732
rect 44329 -1778 44377 -1732
rect 44423 -1778 44471 -1732
rect 44517 -1778 44565 -1732
rect 44611 -1778 44659 -1732
rect 44705 -1778 44753 -1732
rect 44799 -1778 44847 -1732
rect 44893 -1778 44941 -1732
rect 44987 -1778 45035 -1732
rect 45081 -1778 45129 -1732
rect 45175 -1778 45223 -1732
rect 45269 -1778 45317 -1732
rect 45363 -1778 45411 -1732
rect 45457 -1778 45505 -1732
rect 45551 -1778 45599 -1732
rect 45645 -1778 45693 -1732
rect 45739 -1778 45787 -1732
rect 45833 -1778 45881 -1732
rect 45927 -1778 45975 -1732
rect 46021 -1778 46069 -1732
rect 46115 -1778 46163 -1732
rect 46209 -1778 46257 -1732
rect 46303 -1778 46351 -1732
rect 46397 -1778 46445 -1732
rect 46491 -1778 46539 -1732
rect 46585 -1778 46633 -1732
rect 46679 -1778 46727 -1732
rect 46773 -1778 46821 -1732
rect 46867 -1778 46915 -1732
rect 46961 -1778 47009 -1732
rect 47055 -1778 47103 -1732
rect 47149 -1778 47197 -1732
rect 47243 -1778 47291 -1732
rect 47337 -1778 47385 -1732
rect 47431 -1778 47479 -1732
rect 47525 -1778 47573 -1732
rect 47619 -1778 47667 -1732
rect 47713 -1778 47761 -1732
rect 47807 -1778 47855 -1732
rect 47901 -1778 47949 -1732
rect 47995 -1778 48043 -1732
rect 48089 -1778 48137 -1732
rect 48183 -1778 48231 -1732
rect 48277 -1778 48325 -1732
rect 48371 -1778 48419 -1732
rect 48465 -1778 48513 -1732
rect 48559 -1778 48607 -1732
rect 48653 -1778 48701 -1732
rect 48747 -1778 48795 -1732
rect 48841 -1778 48889 -1732
rect 48935 -1778 48983 -1732
rect 49029 -1778 49077 -1732
rect 49123 -1778 49171 -1732
rect 49217 -1778 49265 -1732
rect 49311 -1778 49359 -1732
rect 49405 -1778 49453 -1732
rect 49499 -1778 49547 -1732
rect 49593 -1778 49641 -1732
rect 49687 -1778 49735 -1732
rect 49781 -1778 49829 -1732
rect 49875 -1778 49923 -1732
rect 49969 -1778 50017 -1732
rect 50063 -1778 50111 -1732
rect 50157 -1778 51535 -1732
rect 51581 -1778 51629 -1732
rect 51675 -1778 51723 -1732
rect 51769 -1778 51817 -1732
rect 51863 -1778 51911 -1732
rect 51957 -1778 52005 -1732
rect 52051 -1778 52099 -1732
rect 52145 -1778 52193 -1732
rect 52239 -1778 52287 -1732
rect 52333 -1778 52381 -1732
rect 52427 -1778 52475 -1732
rect 52521 -1778 52569 -1732
rect 52615 -1778 52663 -1732
rect 52709 -1778 52757 -1732
rect 52803 -1778 52851 -1732
rect 52897 -1778 52945 -1732
rect 52991 -1778 53039 -1732
rect 53085 -1778 53133 -1732
rect 53179 -1778 53227 -1732
rect 53273 -1778 53321 -1732
rect 53367 -1778 53415 -1732
rect 53461 -1778 53509 -1732
rect 53555 -1778 53603 -1732
rect 53649 -1778 53697 -1732
rect 53743 -1778 53791 -1732
rect 53837 -1778 53885 -1732
rect 53931 -1778 53979 -1732
rect 54025 -1778 54073 -1732
rect 54119 -1778 54167 -1732
rect 54213 -1778 54261 -1732
rect 54307 -1778 54355 -1732
rect 54401 -1778 54449 -1732
rect 54495 -1778 54543 -1732
rect 54589 -1778 54637 -1732
rect 54683 -1778 54731 -1732
rect 54777 -1778 54825 -1732
rect 54871 -1778 54919 -1732
rect 54965 -1778 55013 -1732
rect 55059 -1778 55107 -1732
rect 55153 -1778 55201 -1732
rect 55247 -1778 55295 -1732
rect 55341 -1778 55389 -1732
rect 55435 -1778 55483 -1732
rect 55529 -1778 55577 -1732
rect 55623 -1778 55671 -1732
rect 55717 -1778 55765 -1732
rect 55811 -1778 55859 -1732
rect 55905 -1778 55953 -1732
rect 55999 -1778 56047 -1732
rect 56093 -1778 56141 -1732
rect 56187 -1778 56235 -1732
rect 56281 -1778 56329 -1732
rect 56375 -1778 56423 -1732
rect 56469 -1778 56517 -1732
rect 56563 -1778 56611 -1732
rect 56657 -1778 56705 -1732
rect 56751 -1778 56799 -1732
rect 56845 -1778 56893 -1732
rect 56939 -1778 56987 -1732
rect 57033 -1778 57081 -1732
rect 57127 -1778 57175 -1732
rect 57221 -1778 57269 -1732
rect 57315 -1778 57363 -1732
rect 57409 -1778 57457 -1732
rect 57503 -1778 57551 -1732
rect 57597 -1778 57645 -1732
rect 57691 -1778 57739 -1732
rect 57785 -1778 57833 -1732
rect 57879 -1778 57927 -1732
rect 57973 -1778 58021 -1732
rect 58067 -1778 58115 -1732
rect 58161 -1778 58209 -1732
rect 58255 -1778 58303 -1732
rect 58349 -1778 58397 -1732
rect 58443 -1778 58491 -1732
rect 58537 -1778 58585 -1732
rect 58631 -1778 58679 -1732
rect 58725 -1778 58773 -1732
rect 58819 -1778 58867 -1732
rect 58913 -1778 58961 -1732
rect 59007 -1778 59055 -1732
rect 59101 -1778 59149 -1732
rect 59195 -1778 59243 -1732
rect 59289 -1778 59337 -1732
rect 59383 -1778 59431 -1732
rect 59477 -1778 59525 -1732
rect 59571 -1778 59619 -1732
rect 59665 -1778 59713 -1732
rect 59759 -1778 59807 -1732
rect 59853 -1778 61231 -1732
rect 61277 -1778 61325 -1732
rect 61371 -1778 61419 -1732
rect 61465 -1778 61513 -1732
rect 61559 -1778 61607 -1732
rect 61653 -1778 61701 -1732
rect 61747 -1778 61795 -1732
rect 61841 -1778 61889 -1732
rect 61935 -1778 61983 -1732
rect 62029 -1778 62077 -1732
rect 62123 -1778 62171 -1732
rect 62217 -1778 62265 -1732
rect 62311 -1778 62359 -1732
rect 62405 -1778 62453 -1732
rect 62499 -1778 62547 -1732
rect 62593 -1778 62641 -1732
rect 62687 -1778 62735 -1732
rect 62781 -1778 62829 -1732
rect 62875 -1778 62923 -1732
rect 62969 -1778 63017 -1732
rect 63063 -1778 63111 -1732
rect 63157 -1778 63205 -1732
rect 63251 -1778 63299 -1732
rect 63345 -1778 63393 -1732
rect 63439 -1778 63487 -1732
rect 63533 -1778 63581 -1732
rect 63627 -1778 63675 -1732
rect 63721 -1778 63769 -1732
rect 63815 -1778 63863 -1732
rect 63909 -1778 63957 -1732
rect 64003 -1778 64051 -1732
rect 64097 -1778 64145 -1732
rect 64191 -1778 64239 -1732
rect 64285 -1778 64333 -1732
rect 64379 -1778 64427 -1732
rect 64473 -1778 64521 -1732
rect 64567 -1778 64615 -1732
rect 64661 -1778 64709 -1732
rect 64755 -1778 64803 -1732
rect 64849 -1778 64897 -1732
rect 64943 -1778 64991 -1732
rect 65037 -1778 65085 -1732
rect 65131 -1778 65179 -1732
rect 65225 -1778 65273 -1732
rect 65319 -1778 65367 -1732
rect 65413 -1778 65532 -1732
rect 32024 -1898 65532 -1778
rect 1137 -4308 1297 -1936
rect 1689 -3845 1869 -3837
rect 1689 -3849 2157 -3845
rect 1689 -3901 1701 -3849
rect 1753 -3901 1805 -3849
rect 1857 -3901 2157 -3849
rect 1689 -3953 2157 -3901
rect 1689 -4005 1701 -3953
rect 1753 -4005 1805 -3953
rect 1857 -4005 2157 -3953
rect 2571 -3972 2731 -3682
rect 2561 -3984 2741 -3972
rect 1689 -4017 1869 -4005
rect 2561 -4036 2573 -3984
rect 2625 -4036 2677 -3984
rect 2729 -4036 2741 -3984
rect 2561 -4088 2741 -4036
rect 2561 -4140 2573 -4088
rect 2625 -4140 2677 -4088
rect 2729 -4140 2741 -4088
rect 2561 -4152 2741 -4140
rect 3439 -4308 3599 -1936
rect 4428 -2297 4588 -1936
rect 5039 -2153 5199 -1936
rect 6381 -1946 6448 -1936
rect 6494 -1946 6561 -1936
rect 9483 -1946 9663 -1936
rect 11381 -2153 11541 -1936
rect 5039 -2297 11541 -2153
rect 4428 -2331 11541 -2297
rect 11781 -2331 11941 -1936
rect 16413 -2331 16573 -1936
rect 32024 -2331 32344 -1898
rect 36124 -2331 36444 -1898
rect 40224 -2331 40544 -1898
rect 41684 -2331 42004 -1898
rect 45784 -2331 46104 -1898
rect 49884 -2331 50204 -1898
rect 51344 -2331 51664 -1898
rect 55444 -2331 55764 -1898
rect 59544 -2331 59864 -1898
rect 61004 -2331 61324 -1898
rect 65212 -2331 65532 -1898
rect 4428 -2651 65532 -2331
rect 4428 -4308 4588 -2651
rect 10885 -2721 16917 -2709
rect 7789 -2746 7969 -2736
rect 7789 -2748 8259 -2746
rect 7789 -2800 7801 -2748
rect 7853 -2800 7905 -2748
rect 7957 -2800 8259 -2748
rect 7789 -2852 8259 -2800
rect 7789 -2904 7801 -2852
rect 7853 -2904 7905 -2852
rect 7957 -2904 8259 -2852
rect 7789 -2906 8259 -2904
rect 10885 -2773 10897 -2721
rect 10949 -2773 11001 -2721
rect 11053 -2773 16645 -2721
rect 16697 -2773 16749 -2721
rect 16801 -2773 16853 -2721
rect 16905 -2773 16917 -2721
rect 10885 -2825 16917 -2773
rect 10885 -2877 10897 -2825
rect 10949 -2877 11001 -2825
rect 11053 -2877 16645 -2825
rect 16697 -2877 16749 -2825
rect 16801 -2877 16853 -2825
rect 16905 -2877 16917 -2825
rect 7789 -2916 7969 -2906
rect 10885 -2929 16917 -2877
rect 6381 -2982 6561 -2972
rect 9483 -2982 9663 -2972
rect 6381 -2984 9663 -2982
rect 6381 -3036 6393 -2984
rect 6445 -3036 6497 -2984
rect 6549 -3036 9495 -2984
rect 9547 -3036 9599 -2984
rect 9651 -3036 9663 -2984
rect 10885 -2981 10897 -2929
rect 10949 -2981 11001 -2929
rect 11053 -2981 16645 -2929
rect 16697 -2981 16749 -2929
rect 16801 -2981 16853 -2929
rect 16905 -2981 16917 -2929
rect 10885 -2993 16917 -2981
rect 6381 -3039 9663 -3036
rect 6391 -3085 6448 -3039
rect 6494 -3085 6542 -3039
rect 6588 -3085 6636 -3039
rect 6682 -3085 6730 -3039
rect 6776 -3085 6824 -3039
rect 6870 -3085 6918 -3039
rect 6964 -3085 7012 -3039
rect 7058 -3085 7106 -3039
rect 7152 -3085 7200 -3039
rect 7246 -3085 7294 -3039
rect 7340 -3085 7388 -3039
rect 7434 -3085 7482 -3039
rect 7528 -3085 7576 -3039
rect 7622 -3085 7670 -3039
rect 7716 -3085 7764 -3039
rect 7810 -3085 7858 -3039
rect 7904 -3085 7952 -3039
rect 7998 -3085 8046 -3039
rect 8092 -3085 8140 -3039
rect 8186 -3085 8234 -3039
rect 8280 -3085 8328 -3039
rect 8374 -3085 8422 -3039
rect 8468 -3085 8516 -3039
rect 8562 -3085 8610 -3039
rect 8656 -3085 8704 -3039
rect 8750 -3085 8798 -3039
rect 8844 -3085 8892 -3039
rect 8938 -3085 8986 -3039
rect 9032 -3085 9080 -3039
rect 9126 -3085 9174 -3039
rect 9220 -3085 9268 -3039
rect 9314 -3085 9362 -3039
rect 9408 -3085 9456 -3039
rect 9502 -3085 9550 -3039
rect 9596 -3085 9663 -3039
rect 6381 -3088 9663 -3085
rect 6381 -3140 6393 -3088
rect 6445 -3133 6497 -3088
rect 6445 -3140 6448 -3133
rect 6381 -3152 6448 -3140
rect 6391 -3179 6448 -3152
rect 6494 -3140 6497 -3133
rect 6549 -3140 9495 -3088
rect 9547 -3133 9599 -3088
rect 9547 -3140 9550 -3133
rect 6494 -3142 9550 -3140
rect 6494 -3152 6561 -3142
rect 6494 -3179 6551 -3152
rect 6391 -3227 6551 -3179
rect 6391 -3273 6448 -3227
rect 6494 -3273 6551 -3227
rect 6391 -3321 6551 -3273
rect 6391 -3367 6448 -3321
rect 6494 -3367 6551 -3321
rect 6391 -3415 6551 -3367
rect 6391 -3461 6448 -3415
rect 6494 -3461 6551 -3415
rect 6391 -3509 6551 -3461
rect 6391 -3555 6448 -3509
rect 6494 -3555 6551 -3509
rect 6391 -3603 6551 -3555
rect 6391 -3649 6448 -3603
rect 6494 -3649 6551 -3603
rect 4658 -3694 4838 -3686
rect 4658 -3698 5138 -3694
rect 4658 -3750 4670 -3698
rect 4722 -3750 4774 -3698
rect 4826 -3750 5138 -3698
rect 4658 -3802 5138 -3750
rect 4658 -3854 4670 -3802
rect 4722 -3854 4774 -3802
rect 4826 -3854 5138 -3802
rect 6391 -3697 6551 -3649
rect 6391 -3743 6448 -3697
rect 6494 -3743 6551 -3697
rect 6391 -3791 6551 -3743
rect 6391 -3837 6448 -3791
rect 6494 -3837 6551 -3791
rect 4658 -3866 4838 -3854
rect 386 -4365 4588 -4308
rect 386 -4411 443 -4365
rect 489 -4411 537 -4365
rect 583 -4411 631 -4365
rect 677 -4411 725 -4365
rect 771 -4411 819 -4365
rect 865 -4411 913 -4365
rect 959 -4411 1007 -4365
rect 1053 -4411 1101 -4365
rect 1147 -4411 1195 -4365
rect 1241 -4411 1289 -4365
rect 1335 -4411 1383 -4365
rect 1429 -4411 1477 -4365
rect 1523 -4411 1571 -4365
rect 1617 -4411 1665 -4365
rect 1711 -4411 1759 -4365
rect 1805 -4411 1853 -4365
rect 1899 -4411 1947 -4365
rect 1993 -4411 2041 -4365
rect 2087 -4411 2135 -4365
rect 2181 -4411 2229 -4365
rect 2275 -4411 2323 -4365
rect 2369 -4411 2417 -4365
rect 2463 -4411 2511 -4365
rect 2557 -4411 2605 -4365
rect 2651 -4411 2699 -4365
rect 2745 -4411 2793 -4365
rect 2839 -4411 2887 -4365
rect 2933 -4411 2981 -4365
rect 3027 -4411 3075 -4365
rect 3121 -4411 3169 -4365
rect 3215 -4411 3263 -4365
rect 3309 -4411 3357 -4365
rect 3403 -4411 3451 -4365
rect 3497 -4411 3545 -4365
rect 3591 -4411 3639 -4365
rect 3685 -4411 3733 -4365
rect 3779 -4411 3827 -4365
rect 3873 -4411 3921 -4365
rect 3967 -4411 4015 -4365
rect 4061 -4411 4109 -4365
rect 4155 -4411 4203 -4365
rect 4249 -4411 4297 -4365
rect 4343 -4411 4391 -4365
rect 4437 -4411 4485 -4365
rect 4531 -4411 4588 -4365
rect 386 -4459 4588 -4411
rect 386 -4505 443 -4459
rect 489 -4468 4485 -4459
rect 489 -4505 546 -4468
rect 386 -4553 546 -4505
rect 386 -4599 443 -4553
rect 489 -4599 546 -4553
rect 386 -4647 546 -4599
rect 386 -4693 443 -4647
rect 489 -4693 546 -4647
rect 386 -4741 546 -4693
rect 804 -4642 850 -4468
rect 964 -4642 1010 -4468
rect 1092 -4642 1138 -4468
rect 1252 -4642 1298 -4468
rect 804 -4688 1172 -4642
rect 1218 -4688 1298 -4642
rect 804 -4736 850 -4688
rect 964 -4736 1010 -4688
rect 1092 -4734 1138 -4688
rect 1252 -4734 1298 -4688
rect 1596 -4736 1642 -4468
rect 1689 -4601 1869 -4589
rect 1689 -4653 1701 -4601
rect 1753 -4653 1805 -4601
rect 1857 -4653 1869 -4601
rect 1689 -4665 1869 -4653
rect 2028 -4736 2074 -4468
rect 386 -4787 443 -4741
rect 489 -4787 546 -4741
rect 386 -4835 546 -4787
rect 386 -4881 443 -4835
rect 489 -4881 546 -4835
rect 386 -4929 546 -4881
rect 2229 -4738 2305 -4726
rect 2460 -4736 2506 -4468
rect 2892 -4736 2938 -4468
rect 3324 -4736 3370 -4468
rect 3756 -4644 3802 -4468
rect 3916 -4644 3962 -4468
rect 4076 -4644 4122 -4468
rect 3756 -4690 3836 -4644
rect 3882 -4690 3996 -4644
rect 4042 -4690 4122 -4644
rect 3756 -4736 3802 -4690
rect 3916 -4736 3962 -4690
rect 4076 -4736 4122 -4690
rect 4428 -4505 4485 -4468
rect 4531 -4505 4588 -4459
rect 4428 -4553 4588 -4505
rect 4428 -4599 4485 -4553
rect 4531 -4599 4588 -4553
rect 4428 -4647 4588 -4599
rect 4428 -4693 4485 -4647
rect 4531 -4693 4588 -4647
rect 2229 -4790 2241 -4738
rect 2293 -4790 2305 -4738
rect 2229 -4842 2305 -4790
rect 2229 -4894 2241 -4842
rect 2293 -4894 2305 -4842
rect 2229 -4906 2305 -4894
rect 4428 -4741 4588 -4693
rect 4428 -4787 4485 -4741
rect 4531 -4787 4588 -4741
rect 6391 -3885 6551 -3837
rect 6391 -3931 6448 -3885
rect 6494 -3931 6551 -3885
rect 6391 -3979 6551 -3931
rect 6391 -4025 6448 -3979
rect 6494 -4025 6551 -3979
rect 6391 -4073 6551 -4025
rect 6391 -4119 6448 -4073
rect 6494 -4119 6551 -4073
rect 6391 -4167 6551 -4119
rect 6391 -4213 6448 -4167
rect 6494 -4213 6551 -4167
rect 6391 -4261 6551 -4213
rect 6391 -4307 6448 -4261
rect 6494 -4307 6551 -4261
rect 6391 -4355 6551 -4307
rect 6391 -4401 6448 -4355
rect 6494 -4401 6551 -4355
rect 6391 -4449 6551 -4401
rect 6391 -4495 6448 -4449
rect 6494 -4495 6551 -4449
rect 6391 -4543 6551 -4495
rect 6391 -4589 6448 -4543
rect 6494 -4589 6551 -4543
rect 6391 -4637 6551 -4589
rect 6391 -4683 6448 -4637
rect 6494 -4683 6551 -4637
rect 6391 -4731 6551 -4683
rect 4428 -4835 4588 -4787
rect 4428 -4881 4485 -4835
rect 4531 -4881 4588 -4835
rect 386 -4975 443 -4929
rect 489 -4975 546 -4929
rect 386 -5023 546 -4975
rect 4428 -4929 4588 -4881
rect 4428 -4975 4485 -4929
rect 4531 -4975 4588 -4929
rect 386 -5069 443 -5023
rect 489 -5069 546 -5023
rect 386 -5117 546 -5069
rect 386 -5163 443 -5117
rect 489 -5163 546 -5117
rect 386 -5211 546 -5163
rect 3525 -5028 3601 -5016
rect 3525 -5080 3537 -5028
rect 3589 -5080 3601 -5028
rect 3525 -5132 3601 -5080
rect 3525 -5184 3537 -5132
rect 3589 -5184 3601 -5132
rect 3525 -5196 3601 -5184
rect 4428 -5023 4588 -4975
rect 4428 -5069 4485 -5023
rect 4531 -5069 4588 -5023
rect 6068 -5044 6228 -4754
rect 6391 -4777 6448 -4731
rect 6494 -4777 6551 -4731
rect 6391 -4825 6551 -4777
rect 6391 -4871 6448 -4825
rect 6494 -4871 6551 -4825
rect 6391 -4919 6551 -4871
rect 6391 -4965 6448 -4919
rect 6494 -4965 6551 -4919
rect 6391 -5013 6551 -4965
rect 4428 -5117 4588 -5069
rect 4428 -5163 4485 -5117
rect 4531 -5163 4588 -5117
rect 386 -5257 443 -5211
rect 489 -5257 546 -5211
rect 386 -5305 546 -5257
rect 386 -5351 443 -5305
rect 489 -5351 546 -5305
rect 4428 -5211 4588 -5163
rect 4428 -5257 4485 -5211
rect 4531 -5257 4588 -5211
rect 6058 -5056 6238 -5044
rect 6058 -5108 6070 -5056
rect 6122 -5108 6174 -5056
rect 6226 -5108 6238 -5056
rect 6058 -5160 6238 -5108
rect 6058 -5212 6070 -5160
rect 6122 -5212 6174 -5160
rect 6226 -5212 6238 -5160
rect 6058 -5224 6238 -5212
rect 6391 -5059 6448 -5013
rect 6494 -5059 6551 -5013
rect 6391 -5107 6551 -5059
rect 6391 -5153 6448 -5107
rect 6494 -5153 6551 -5107
rect 6391 -5201 6551 -5153
rect 4428 -5305 4588 -5257
rect 386 -5399 546 -5351
rect 386 -5445 443 -5399
rect 489 -5445 546 -5399
rect 386 -5493 546 -5445
rect 386 -5539 443 -5493
rect 489 -5539 546 -5493
rect 3093 -5352 3169 -5340
rect 3093 -5404 3105 -5352
rect 3157 -5404 3169 -5352
rect 3093 -5456 3169 -5404
rect 3093 -5508 3105 -5456
rect 3157 -5508 3169 -5456
rect 386 -5587 546 -5539
rect 386 -5633 443 -5587
rect 489 -5633 546 -5587
rect 386 -5681 546 -5633
rect 386 -5727 443 -5681
rect 489 -5727 546 -5681
rect 386 -5775 546 -5727
rect 386 -5821 443 -5775
rect 489 -5821 546 -5775
rect 386 -5869 546 -5821
rect 386 -5915 443 -5869
rect 489 -5915 546 -5869
rect 386 -5963 546 -5915
rect 386 -6009 443 -5963
rect 489 -6009 546 -5963
rect 804 -5902 850 -5510
rect 964 -5902 1010 -5510
rect 1380 -5567 1426 -5510
rect 1812 -5567 1858 -5510
rect 2244 -5567 2290 -5511
rect 1380 -5613 2290 -5567
rect 2676 -5567 2722 -5510
rect 3093 -5520 3169 -5508
rect 4428 -5351 4485 -5305
rect 4531 -5351 4588 -5305
rect 4428 -5399 4588 -5351
rect 4428 -5445 4485 -5399
rect 4531 -5445 4588 -5399
rect 4428 -5493 4588 -5445
rect 3108 -5567 3154 -5520
rect 2676 -5613 3154 -5567
rect 4428 -5539 4485 -5493
rect 4531 -5539 4588 -5493
rect 4428 -5587 4588 -5539
rect 4428 -5633 4485 -5587
rect 4531 -5633 4588 -5587
rect 4428 -5681 4588 -5633
rect 4428 -5727 4485 -5681
rect 4531 -5727 4588 -5681
rect 4428 -5775 4588 -5727
rect 1388 -5862 1616 -5816
rect 1662 -5862 1720 -5816
rect 1766 -5862 1824 -5816
rect 1870 -5862 1928 -5816
rect 1974 -5862 2032 -5816
rect 2078 -5862 2136 -5816
rect 2182 -5862 2298 -5816
rect 804 -5948 884 -5902
rect 930 -5948 1180 -5902
rect 1226 -5948 1306 -5902
rect 804 -5996 850 -5948
rect 964 -5996 1010 -5948
rect 1100 -5994 1146 -5948
rect 1260 -5994 1306 -5948
rect 1388 -5996 1434 -5862
rect 1820 -5996 1866 -5862
rect 2252 -5986 2298 -5862
rect 4428 -5821 4485 -5775
rect 4531 -5821 4588 -5775
rect 4428 -5869 4588 -5821
rect 2788 -5939 3748 -5893
rect 3794 -5939 4044 -5893
rect 4090 -5939 4170 -5893
rect 386 -6057 546 -6009
rect 386 -6103 443 -6057
rect 489 -6103 546 -6057
rect 386 -6151 546 -6103
rect 386 -6197 443 -6151
rect 489 -6197 546 -6151
rect 2239 -5998 2315 -5986
rect 2239 -6050 2251 -5998
rect 2303 -6050 2315 -5998
rect 2239 -6102 2315 -6050
rect 2239 -6154 2251 -6102
rect 2303 -6154 2315 -6102
rect 2239 -6166 2315 -6154
rect 2613 -5998 2689 -5986
rect 2788 -5996 2834 -5939
rect 2613 -6050 2625 -5998
rect 2677 -6050 2689 -5998
rect 2613 -6102 2689 -6050
rect 2613 -6154 2625 -6102
rect 2677 -6154 2689 -6102
rect 2613 -6166 2689 -6154
rect 2933 -5998 3009 -5986
rect 3108 -5996 3154 -5939
rect 3668 -5996 3714 -5939
rect 3828 -5996 3874 -5939
rect 3964 -5996 4010 -5939
rect 4124 -5996 4170 -5939
rect 4428 -5915 4485 -5869
rect 4531 -5915 4588 -5869
rect 4428 -5963 4588 -5915
rect 2933 -6050 2945 -5998
rect 2997 -6050 3009 -5998
rect 2933 -6102 3009 -6050
rect 2933 -6154 2945 -6102
rect 2997 -6154 3009 -6102
rect 2933 -6166 3009 -6154
rect 4428 -6009 4485 -5963
rect 4531 -6009 4588 -5963
rect 4428 -6057 4588 -6009
rect 4428 -6103 4485 -6057
rect 4531 -6103 4588 -6057
rect 4428 -6151 4588 -6103
rect 386 -6245 546 -6197
rect 386 -6291 443 -6245
rect 489 -6291 546 -6245
rect 386 -6339 546 -6291
rect 386 -6385 443 -6339
rect 489 -6385 546 -6339
rect 386 -6433 546 -6385
rect 386 -6479 443 -6433
rect 489 -6479 546 -6433
rect 386 -6527 546 -6479
rect 386 -6573 443 -6527
rect 489 -6573 546 -6527
rect 386 -6621 546 -6573
rect 4428 -6197 4485 -6151
rect 4531 -6197 4588 -6151
rect 4428 -6245 4588 -6197
rect 4428 -6291 4485 -6245
rect 4531 -6291 4588 -6245
rect 6391 -5247 6448 -5201
rect 6494 -5247 6551 -5201
rect 6391 -5295 6551 -5247
rect 6391 -5341 6448 -5295
rect 6494 -5341 6551 -5295
rect 6391 -5389 6551 -5341
rect 6391 -5435 6448 -5389
rect 6494 -5435 6551 -5389
rect 6391 -5483 6551 -5435
rect 6391 -5529 6448 -5483
rect 6494 -5529 6551 -5483
rect 6391 -5577 6551 -5529
rect 6391 -5623 6448 -5577
rect 6494 -5623 6551 -5577
rect 6391 -5671 6551 -5623
rect 6391 -5717 6448 -5671
rect 6494 -5717 6551 -5671
rect 6391 -5765 6551 -5717
rect 6391 -5811 6448 -5765
rect 6494 -5811 6551 -5765
rect 6391 -5859 6551 -5811
rect 6391 -5905 6448 -5859
rect 6494 -5905 6551 -5859
rect 6391 -5953 6551 -5905
rect 6391 -5999 6448 -5953
rect 6494 -5999 6551 -5953
rect 6391 -6047 6551 -5999
rect 6391 -6093 6448 -6047
rect 6494 -6093 6551 -6047
rect 6391 -6141 6551 -6093
rect 6910 -5372 6956 -3142
rect 7070 -5372 7116 -3142
rect 8703 -3219 8779 -3207
rect 8703 -3222 8715 -3219
rect 7267 -3223 7815 -3222
rect 7267 -3269 7278 -3223
rect 7324 -3269 7758 -3223
rect 7804 -3269 7815 -3223
rect 8227 -3223 8715 -3222
rect 8227 -3269 8238 -3223
rect 8284 -3269 8715 -3223
rect 8767 -3271 8779 -3219
rect 8715 -3283 8779 -3271
rect 7198 -3375 8844 -3329
rect 7198 -3432 7244 -3375
rect 7838 -3432 7884 -3375
rect 8158 -3432 8204 -3375
rect 8798 -3432 8844 -3375
rect 7183 -3448 7259 -3436
rect 7183 -3500 7195 -3448
rect 7247 -3500 7259 -3448
rect 7183 -3552 7259 -3500
rect 7183 -3604 7195 -3552
rect 7247 -3604 7259 -3552
rect 7183 -3616 7259 -3604
rect 7343 -3448 7419 -3436
rect 7343 -3500 7355 -3448
rect 7407 -3500 7419 -3448
rect 7343 -3552 7419 -3500
rect 7343 -3604 7355 -3552
rect 7407 -3604 7419 -3552
rect 7343 -3616 7358 -3604
rect 7404 -3616 7419 -3604
rect 7663 -3448 7739 -3436
rect 7663 -3500 7675 -3448
rect 7727 -3500 7739 -3448
rect 7663 -3552 7739 -3500
rect 7663 -3604 7675 -3552
rect 7727 -3604 7739 -3552
rect 7518 -3663 7564 -3606
rect 7663 -3616 7678 -3604
rect 7724 -3616 7739 -3604
rect 7983 -3448 8059 -3436
rect 7983 -3500 7995 -3448
rect 8047 -3500 8059 -3448
rect 7983 -3552 8059 -3500
rect 7983 -3604 7995 -3552
rect 8047 -3604 8059 -3552
rect 7983 -3616 7998 -3604
rect 8044 -3616 8059 -3604
rect 8303 -3448 8379 -3436
rect 8303 -3500 8315 -3448
rect 8367 -3500 8379 -3448
rect 8303 -3552 8379 -3500
rect 8303 -3604 8315 -3552
rect 8367 -3604 8379 -3552
rect 8303 -3616 8318 -3604
rect 8364 -3616 8379 -3604
rect 8463 -3448 8539 -3437
rect 8463 -3500 8475 -3448
rect 8527 -3500 8539 -3448
rect 8463 -3552 8539 -3500
rect 8463 -3604 8475 -3552
rect 8527 -3604 8539 -3552
rect 8463 -3617 8539 -3604
rect 8623 -3448 8699 -3436
rect 8623 -3500 8635 -3448
rect 8687 -3500 8699 -3448
rect 8623 -3552 8699 -3500
rect 8623 -3604 8635 -3552
rect 8687 -3604 8699 -3552
rect 8623 -3616 8638 -3604
rect 8684 -3616 8699 -3604
rect 8478 -3663 8524 -3617
rect 7518 -3709 8524 -3663
rect 7267 -3819 7278 -3773
rect 7324 -3819 7438 -3773
rect 7484 -3819 7758 -3773
rect 7804 -3819 7815 -3773
rect 8010 -3865 8056 -3709
rect 8782 -3755 8858 -3743
rect 8782 -3773 8794 -3755
rect 8227 -3819 8238 -3773
rect 8284 -3819 8398 -3773
rect 8444 -3819 8718 -3773
rect 8764 -3807 8794 -3773
rect 8846 -3807 8858 -3755
rect 8764 -3819 8858 -3807
rect 7198 -3911 8844 -3865
rect 7198 -3968 7244 -3911
rect 7838 -3968 7884 -3911
rect 8158 -3968 8204 -3911
rect 8798 -3968 8844 -3911
rect 7343 -3984 7419 -3972
rect 7343 -4036 7355 -3984
rect 7407 -4036 7419 -3984
rect 7343 -4088 7419 -4036
rect 7343 -4140 7355 -4088
rect 7407 -4140 7419 -4088
rect 7343 -4142 7358 -4140
rect 7404 -4142 7419 -4140
rect 7343 -4152 7419 -4142
rect 7503 -3984 7579 -3973
rect 7503 -4036 7515 -3984
rect 7567 -4036 7579 -3984
rect 7503 -4088 7579 -4036
rect 7503 -4140 7515 -4088
rect 7567 -4140 7579 -4088
rect 7503 -4153 7579 -4140
rect 7663 -3984 7739 -3972
rect 7663 -4036 7675 -3984
rect 7727 -4036 7739 -3984
rect 7663 -4088 7739 -4036
rect 7663 -4140 7675 -4088
rect 7727 -4140 7739 -4088
rect 7663 -4142 7678 -4140
rect 7724 -4142 7739 -4140
rect 7663 -4152 7739 -4142
rect 7983 -3984 8059 -3972
rect 7983 -4036 7995 -3984
rect 8047 -4036 8059 -3984
rect 7983 -4088 8059 -4036
rect 7983 -4140 7995 -4088
rect 8047 -4140 8059 -4088
rect 7983 -4142 7998 -4140
rect 8044 -4142 8059 -4140
rect 7983 -4152 8059 -4142
rect 8303 -3984 8379 -3972
rect 8303 -4036 8315 -3984
rect 8367 -4036 8379 -3984
rect 8303 -4088 8379 -4036
rect 8303 -4140 8315 -4088
rect 8367 -4140 8379 -4088
rect 8303 -4142 8318 -4140
rect 8364 -4142 8379 -4140
rect 8623 -3984 8699 -3972
rect 8623 -4036 8635 -3984
rect 8687 -4036 8699 -3984
rect 8623 -4088 8699 -4036
rect 8623 -4140 8635 -4088
rect 8687 -4140 8699 -4088
rect 8623 -4142 8638 -4140
rect 8684 -4142 8699 -4140
rect 8303 -4152 8379 -4142
rect 7518 -4199 7564 -4153
rect 8478 -4199 8524 -4142
rect 8623 -4152 8699 -4142
rect 7518 -4245 8524 -4199
rect 7267 -4340 7278 -4294
rect 7324 -4340 7438 -4294
rect 7484 -4340 7758 -4294
rect 7804 -4340 7815 -4294
rect 7993 -4401 8039 -4245
rect 8585 -4291 8661 -4279
rect 8585 -4294 8597 -4291
rect 8227 -4340 8238 -4294
rect 8284 -4340 8398 -4294
rect 8444 -4340 8597 -4294
rect 8585 -4343 8597 -4340
rect 8649 -4294 8661 -4291
rect 8649 -4340 8718 -4294
rect 8764 -4340 8775 -4294
rect 8649 -4343 8661 -4340
rect 8585 -4355 8661 -4343
rect 7198 -4447 8844 -4401
rect 7198 -4504 7244 -4447
rect 7838 -4504 7884 -4447
rect 8158 -4504 8204 -4447
rect 8798 -4504 8844 -4447
rect 7183 -4520 7259 -4508
rect 7183 -4572 7195 -4520
rect 7247 -4572 7259 -4520
rect 7183 -4624 7259 -4572
rect 7183 -4676 7195 -4624
rect 7247 -4676 7259 -4624
rect 7183 -4688 7259 -4676
rect 7343 -4520 7419 -4508
rect 7343 -4572 7355 -4520
rect 7407 -4572 7419 -4520
rect 7343 -4624 7419 -4572
rect 7343 -4676 7355 -4624
rect 7407 -4676 7419 -4624
rect 7343 -4688 7358 -4676
rect 7404 -4688 7419 -4676
rect 7663 -4520 7739 -4508
rect 7663 -4572 7675 -4520
rect 7727 -4572 7739 -4520
rect 7663 -4624 7739 -4572
rect 7663 -4676 7675 -4624
rect 7727 -4676 7739 -4624
rect 7663 -4678 7678 -4676
rect 7724 -4678 7739 -4676
rect 7518 -4735 7564 -4678
rect 7663 -4688 7739 -4678
rect 7983 -4520 8059 -4508
rect 7983 -4572 7995 -4520
rect 8047 -4572 8059 -4520
rect 7983 -4624 8059 -4572
rect 7983 -4676 7995 -4624
rect 8047 -4676 8059 -4624
rect 7983 -4678 7998 -4676
rect 8044 -4678 8059 -4676
rect 7983 -4688 8059 -4678
rect 8303 -4520 8379 -4508
rect 8303 -4572 8315 -4520
rect 8367 -4572 8379 -4520
rect 8303 -4624 8379 -4572
rect 8303 -4676 8315 -4624
rect 8367 -4676 8379 -4624
rect 8303 -4678 8318 -4676
rect 8364 -4678 8379 -4676
rect 8303 -4688 8379 -4678
rect 8463 -4520 8539 -4508
rect 8463 -4572 8475 -4520
rect 8527 -4572 8539 -4520
rect 8463 -4624 8539 -4572
rect 8463 -4676 8475 -4624
rect 8527 -4676 8539 -4624
rect 8463 -4689 8539 -4676
rect 8623 -4520 8699 -4508
rect 8623 -4572 8635 -4520
rect 8687 -4572 8699 -4520
rect 8623 -4624 8699 -4572
rect 8623 -4676 8635 -4624
rect 8687 -4676 8699 -4624
rect 8623 -4678 8638 -4676
rect 8684 -4678 8699 -4676
rect 8623 -4688 8699 -4678
rect 8478 -4735 8524 -4689
rect 7518 -4781 8524 -4735
rect 7267 -4874 7278 -4828
rect 7324 -4874 7438 -4828
rect 7484 -4874 7758 -4828
rect 7804 -4874 7815 -4828
rect 7993 -4937 8039 -4781
rect 8703 -4825 8779 -4813
rect 8703 -4828 8715 -4825
rect 8227 -4874 8238 -4828
rect 8284 -4874 8398 -4828
rect 8444 -4874 8715 -4828
rect 8703 -4877 8715 -4874
rect 8767 -4877 8779 -4825
rect 8703 -4889 8779 -4877
rect 7198 -4983 8844 -4937
rect 7198 -5040 7244 -4983
rect 7838 -5040 7884 -4983
rect 8158 -5040 8204 -4983
rect 8798 -5040 8844 -4983
rect 7343 -5056 7419 -5044
rect 7343 -5108 7355 -5056
rect 7407 -5108 7419 -5056
rect 7343 -5160 7419 -5108
rect 7343 -5212 7355 -5160
rect 7407 -5212 7419 -5160
rect 7343 -5224 7358 -5212
rect 7404 -5224 7419 -5212
rect 7503 -5056 7579 -5045
rect 7503 -5108 7515 -5056
rect 7567 -5108 7579 -5056
rect 7503 -5160 7579 -5108
rect 7503 -5212 7515 -5160
rect 7567 -5212 7579 -5160
rect 7503 -5225 7579 -5212
rect 7663 -5056 7739 -5044
rect 7663 -5108 7675 -5056
rect 7727 -5108 7739 -5056
rect 7663 -5160 7739 -5108
rect 7663 -5212 7675 -5160
rect 7727 -5212 7739 -5160
rect 7663 -5224 7678 -5212
rect 7724 -5224 7739 -5212
rect 7983 -5056 8059 -5044
rect 7983 -5108 7995 -5056
rect 8047 -5108 8059 -5056
rect 7983 -5160 8059 -5108
rect 7983 -5212 7995 -5160
rect 8047 -5212 8059 -5160
rect 7983 -5224 7998 -5212
rect 8044 -5224 8059 -5212
rect 8303 -5056 8379 -5044
rect 8303 -5108 8315 -5056
rect 8367 -5108 8379 -5056
rect 8303 -5160 8379 -5108
rect 8303 -5212 8315 -5160
rect 8367 -5212 8379 -5160
rect 8623 -5056 8699 -5044
rect 8623 -5108 8635 -5056
rect 8687 -5108 8699 -5056
rect 8623 -5160 8699 -5108
rect 8623 -5212 8635 -5160
rect 8687 -5212 8699 -5160
rect 8303 -5224 8318 -5212
rect 8364 -5224 8379 -5212
rect 7518 -5271 7564 -5225
rect 8478 -5271 8524 -5212
rect 8623 -5224 8638 -5212
rect 8684 -5224 8699 -5212
rect 7518 -5317 8524 -5271
rect 6910 -5418 6990 -5372
rect 7036 -5418 7116 -5372
rect 7267 -5410 7278 -5364
rect 7324 -5410 7438 -5364
rect 7484 -5410 7758 -5364
rect 7804 -5410 7815 -5364
rect 6910 -6112 6956 -5418
rect 7070 -6112 7116 -5418
rect 7993 -5473 8039 -5317
rect 8782 -5361 8858 -5349
rect 8782 -5364 8794 -5361
rect 8227 -5410 8238 -5364
rect 8284 -5410 8398 -5364
rect 8444 -5366 8794 -5364
rect 8444 -5410 8718 -5366
rect 8705 -5412 8718 -5410
rect 8764 -5412 8794 -5366
rect 8782 -5413 8794 -5412
rect 8846 -5413 8858 -5361
rect 8782 -5425 8858 -5413
rect 8926 -5372 8972 -3142
rect 9086 -5372 9132 -3142
rect 9483 -3152 9550 -3142
rect 8926 -5418 9006 -5372
rect 9052 -5418 9132 -5372
rect 7198 -5519 8844 -5473
rect 7198 -5576 7244 -5519
rect 7343 -5584 7358 -5572
rect 7404 -5584 7419 -5572
rect 7343 -5636 7355 -5584
rect 7407 -5636 7419 -5584
rect 7343 -5688 7419 -5636
rect 7343 -5740 7355 -5688
rect 7407 -5740 7419 -5688
rect 7343 -5752 7419 -5740
rect 7663 -5584 7678 -5572
rect 7724 -5584 7739 -5572
rect 7838 -5576 7884 -5519
rect 7663 -5636 7675 -5584
rect 7727 -5636 7739 -5584
rect 7663 -5688 7739 -5636
rect 7663 -5740 7675 -5688
rect 7727 -5740 7739 -5688
rect 7518 -5807 7564 -5748
rect 7663 -5752 7678 -5740
rect 7724 -5752 7739 -5740
rect 7983 -5584 7998 -5572
rect 8044 -5584 8059 -5572
rect 8158 -5576 8204 -5519
rect 7983 -5636 7995 -5584
rect 8047 -5636 8059 -5584
rect 7983 -5688 8059 -5636
rect 7983 -5740 7995 -5688
rect 8047 -5740 8059 -5688
rect 7983 -5752 7998 -5740
rect 8044 -5752 8059 -5740
rect 8303 -5584 8318 -5572
rect 8364 -5584 8379 -5572
rect 8303 -5636 8315 -5584
rect 8367 -5636 8379 -5584
rect 8303 -5688 8379 -5636
rect 8303 -5740 8315 -5688
rect 8367 -5740 8379 -5688
rect 8303 -5752 8318 -5740
rect 8364 -5752 8379 -5740
rect 8463 -5592 8539 -5580
rect 8463 -5644 8475 -5592
rect 8527 -5644 8539 -5592
rect 8463 -5696 8539 -5644
rect 8463 -5748 8475 -5696
rect 8527 -5748 8539 -5696
rect 8463 -5761 8539 -5748
rect 8623 -5584 8638 -5572
rect 8684 -5584 8699 -5572
rect 8798 -5576 8844 -5519
rect 8623 -5636 8635 -5584
rect 8687 -5636 8699 -5584
rect 8623 -5688 8699 -5636
rect 8623 -5740 8635 -5688
rect 8687 -5740 8699 -5688
rect 8623 -5752 8638 -5740
rect 8684 -5752 8699 -5740
rect 8478 -5807 8524 -5761
rect 7518 -5853 8524 -5807
rect 7267 -5946 7278 -5900
rect 7324 -5946 7438 -5900
rect 7484 -5946 7758 -5900
rect 7804 -5946 7815 -5900
rect 7993 -6009 8039 -5853
rect 8782 -5876 8858 -5864
rect 8782 -5900 8794 -5876
rect 8227 -5946 8238 -5900
rect 8284 -5946 8398 -5900
rect 8444 -5902 8794 -5900
rect 8444 -5946 8718 -5902
rect 8707 -5948 8718 -5946
rect 8764 -5928 8794 -5902
rect 8846 -5928 8858 -5876
rect 8764 -5946 8858 -5928
rect 8764 -5948 8775 -5946
rect 7198 -6055 8844 -6009
rect 7198 -6112 7244 -6055
rect 6391 -6187 6448 -6141
rect 6494 -6187 6551 -6141
rect 6391 -6235 6551 -6187
rect 6391 -6272 6448 -6235
rect 4428 -6339 4588 -6291
rect 4428 -6385 4485 -6339
rect 4531 -6385 4588 -6339
rect 4428 -6433 4588 -6385
rect 4428 -6479 4485 -6433
rect 4531 -6479 4588 -6433
rect 4428 -6527 4588 -6479
rect 4428 -6573 4485 -6527
rect 4531 -6573 4588 -6527
rect 386 -6667 443 -6621
rect 489 -6667 546 -6621
rect 386 -6715 546 -6667
rect 386 -6761 443 -6715
rect 489 -6761 546 -6715
rect 386 -6809 546 -6761
rect 3437 -6614 3513 -6602
rect 3437 -6666 3449 -6614
rect 3501 -6666 3513 -6614
rect 3437 -6718 3513 -6666
rect 3437 -6770 3449 -6718
rect 3501 -6770 3513 -6718
rect 4428 -6621 4588 -6573
rect 4428 -6667 4485 -6621
rect 4531 -6667 4588 -6621
rect 4428 -6715 4588 -6667
rect 4428 -6761 4485 -6715
rect 4531 -6761 4588 -6715
rect 386 -6855 443 -6809
rect 489 -6855 546 -6809
rect 386 -6903 546 -6855
rect 386 -6949 443 -6903
rect 489 -6949 546 -6903
rect 386 -6997 546 -6949
rect 386 -7043 443 -6997
rect 489 -7043 546 -6997
rect 386 -7091 546 -7043
rect 386 -7137 443 -7091
rect 489 -7137 546 -7091
rect 386 -7185 546 -7137
rect 386 -7231 443 -7185
rect 489 -7231 546 -7185
rect 386 -7279 546 -7231
rect 386 -7325 443 -7279
rect 489 -7325 546 -7279
rect 386 -7373 546 -7325
rect 386 -7419 443 -7373
rect 489 -7419 546 -7373
rect 386 -7467 546 -7419
rect 386 -7513 443 -7467
rect 489 -7513 546 -7467
rect 386 -7561 546 -7513
rect 386 -7607 443 -7561
rect 489 -7598 546 -7561
rect 804 -7598 850 -6770
rect 964 -7598 1010 -6770
rect 1260 -6827 1306 -6770
rect 1604 -6827 1650 -6770
rect 2036 -6827 2082 -6770
rect 2468 -6827 2514 -6770
rect 2628 -6807 2674 -6770
rect 2948 -6807 2994 -6770
rect 1260 -6873 2514 -6827
rect 2617 -6818 2685 -6807
rect 2617 -6864 2628 -6818
rect 2674 -6864 2685 -6818
rect 2617 -6875 2685 -6864
rect 2937 -6818 3005 -6807
rect 2937 -6864 2948 -6818
rect 2994 -6864 3005 -6818
rect 2937 -6875 3005 -6864
rect 3205 -6816 3273 -6805
rect 3324 -6816 3370 -6770
rect 3437 -6782 3513 -6770
rect 3205 -6862 3216 -6816
rect 3262 -6862 3370 -6816
rect 3205 -6873 3273 -6862
rect 1100 -7199 3706 -7153
rect 1100 -7256 1146 -7199
rect 1420 -7256 1466 -7199
rect 1740 -7256 1786 -7199
rect 2060 -7256 2106 -7199
rect 2380 -7256 2426 -7199
rect 2700 -7256 2746 -7199
rect 3020 -7256 3066 -7199
rect 3340 -7256 3386 -7199
rect 3660 -7256 3706 -7199
rect 1260 -7387 1306 -7330
rect 1580 -7387 1626 -7329
rect 1900 -7387 1946 -7330
rect 2220 -7387 2266 -7330
rect 2540 -7387 2586 -7330
rect 2860 -7387 2906 -7331
rect 3180 -7387 3226 -7330
rect 3500 -7372 3546 -7330
rect 3485 -7384 3561 -7372
rect 3485 -7387 3497 -7384
rect 1260 -7433 1340 -7387
rect 1386 -7433 1500 -7387
rect 1546 -7433 1980 -7387
rect 2026 -7433 2620 -7387
rect 2666 -7433 3497 -7387
rect 2860 -7434 2906 -7433
rect 3485 -7436 3497 -7433
rect 3549 -7436 3561 -7384
rect 3485 -7488 3561 -7436
rect 3485 -7540 3497 -7488
rect 3549 -7540 3561 -7488
rect 3485 -7552 3561 -7540
rect 3964 -7598 4010 -6770
rect 4124 -7598 4170 -6770
rect 4428 -6809 4588 -6761
rect 4428 -6855 4485 -6809
rect 4531 -6855 4588 -6809
rect 4428 -6903 4588 -6855
rect 4428 -6949 4485 -6903
rect 4531 -6949 4588 -6903
rect 4428 -6997 4588 -6949
rect 4428 -7043 4485 -6997
rect 4531 -7043 4588 -6997
rect 4428 -7091 4588 -7043
rect 4428 -7137 4485 -7091
rect 4531 -7137 4588 -7091
rect 4428 -7185 4588 -7137
rect 4428 -7231 4485 -7185
rect 4531 -7231 4588 -7185
rect 4428 -7279 4588 -7231
rect 4428 -7325 4485 -7279
rect 4531 -7325 4588 -7279
rect 4428 -7373 4588 -7325
rect 4428 -7419 4485 -7373
rect 4531 -7419 4588 -7373
rect 4428 -7467 4588 -7419
rect 4428 -7513 4485 -7467
rect 4531 -7513 4588 -7467
rect 4428 -7561 4588 -7513
rect 4428 -7598 4485 -7561
rect 489 -7607 4485 -7598
rect 4531 -7607 4588 -7561
rect 386 -7655 4588 -7607
rect 386 -7701 443 -7655
rect 489 -7701 537 -7655
rect 583 -7701 631 -7655
rect 677 -7701 725 -7655
rect 771 -7701 819 -7655
rect 865 -7701 913 -7655
rect 959 -7701 1007 -7655
rect 1053 -7701 1101 -7655
rect 1147 -7701 1195 -7655
rect 1241 -7701 1289 -7655
rect 1335 -7701 1383 -7655
rect 1429 -7701 1477 -7655
rect 1523 -7701 1571 -7655
rect 1617 -7701 1665 -7655
rect 1711 -7701 1759 -7655
rect 1805 -7701 1853 -7655
rect 1899 -7701 1947 -7655
rect 1993 -7701 2041 -7655
rect 2087 -7701 2135 -7655
rect 2181 -7701 2229 -7655
rect 2275 -7701 2323 -7655
rect 2369 -7701 2417 -7655
rect 2463 -7701 2511 -7655
rect 2557 -7701 2605 -7655
rect 2651 -7701 2699 -7655
rect 2745 -7701 2793 -7655
rect 2839 -7701 2887 -7655
rect 2933 -7701 2981 -7655
rect 3027 -7701 3075 -7655
rect 3121 -7701 3169 -7655
rect 3215 -7701 3263 -7655
rect 3309 -7701 3357 -7655
rect 3403 -7701 3451 -7655
rect 3497 -7701 3545 -7655
rect 3591 -7701 3639 -7655
rect 3685 -7701 3733 -7655
rect 3779 -7701 3827 -7655
rect 3873 -7701 3921 -7655
rect 3967 -7701 4015 -7655
rect 4061 -7701 4109 -7655
rect 4155 -7701 4203 -7655
rect 4249 -7701 4297 -7655
rect 4343 -7701 4391 -7655
rect 4437 -7701 4485 -7655
rect 4531 -7701 4588 -7655
rect 386 -7758 4588 -7701
rect 5357 -6281 6448 -6272
rect 6494 -6281 6551 -6235
rect 5357 -6329 6551 -6281
rect 7343 -6120 7419 -6108
rect 7343 -6172 7355 -6120
rect 7407 -6172 7419 -6120
rect 7343 -6224 7419 -6172
rect 7343 -6276 7355 -6224
rect 7407 -6276 7419 -6224
rect 7343 -6288 7419 -6276
rect 7503 -6128 7579 -6117
rect 7503 -6180 7515 -6128
rect 7567 -6180 7579 -6128
rect 7503 -6232 7579 -6180
rect 7503 -6284 7515 -6232
rect 7567 -6284 7579 -6232
rect 7503 -6297 7579 -6284
rect 7663 -6120 7678 -6108
rect 7724 -6120 7739 -6108
rect 7838 -6112 7884 -6055
rect 7663 -6172 7675 -6120
rect 7727 -6172 7739 -6120
rect 7663 -6224 7739 -6172
rect 7663 -6276 7675 -6224
rect 7727 -6276 7739 -6224
rect 7663 -6288 7739 -6276
rect 7983 -6120 7998 -6108
rect 8044 -6120 8059 -6108
rect 8158 -6112 8204 -6055
rect 7983 -6172 7995 -6120
rect 8047 -6172 8059 -6120
rect 7983 -6224 8059 -6172
rect 7983 -6276 7995 -6224
rect 8047 -6276 8059 -6224
rect 7983 -6288 8059 -6276
rect 8303 -6120 8318 -6108
rect 8364 -6120 8379 -6108
rect 8303 -6172 8315 -6120
rect 8367 -6172 8379 -6120
rect 8303 -6224 8379 -6172
rect 8303 -6276 8315 -6224
rect 8367 -6276 8379 -6224
rect 8303 -6288 8379 -6276
rect 8623 -6120 8638 -6108
rect 8684 -6120 8699 -6108
rect 8798 -6112 8844 -6055
rect 8926 -6112 8972 -5418
rect 9086 -6112 9132 -5418
rect 9493 -3179 9550 -3152
rect 9596 -3140 9599 -3133
rect 9651 -3140 9663 -3088
rect 11153 -3063 17354 -3051
rect 9596 -3152 9663 -3140
rect 9792 -3113 9972 -3103
rect 9792 -3115 10262 -3113
rect 9596 -3179 9653 -3152
rect 9493 -3227 9653 -3179
rect 9493 -3273 9550 -3227
rect 9596 -3273 9653 -3227
rect 9493 -3321 9653 -3273
rect 9792 -3167 9804 -3115
rect 9856 -3167 9908 -3115
rect 9960 -3167 10262 -3115
rect 9792 -3219 10262 -3167
rect 9792 -3271 9804 -3219
rect 9856 -3271 9908 -3219
rect 9960 -3271 10262 -3219
rect 9792 -3273 10262 -3271
rect 11153 -3115 11165 -3063
rect 11217 -3115 11269 -3063
rect 11321 -3115 17082 -3063
rect 17134 -3115 17186 -3063
rect 17238 -3115 17290 -3063
rect 17342 -3115 17354 -3063
rect 11153 -3167 17354 -3115
rect 11153 -3219 11165 -3167
rect 11217 -3219 11269 -3167
rect 11321 -3219 17082 -3167
rect 17134 -3219 17186 -3167
rect 17238 -3219 17290 -3167
rect 17342 -3219 17354 -3167
rect 11153 -3271 17354 -3219
rect 9792 -3283 9972 -3273
rect 9493 -3367 9550 -3321
rect 9596 -3367 9653 -3321
rect 11153 -3323 11165 -3271
rect 11217 -3323 11269 -3271
rect 11321 -3323 17082 -3271
rect 17134 -3323 17186 -3271
rect 17238 -3323 17290 -3271
rect 17342 -3323 17354 -3271
rect 11153 -3335 17354 -3323
rect 9493 -3415 9653 -3367
rect 9493 -3461 9550 -3415
rect 9596 -3461 9653 -3415
rect 17590 -3346 17910 -2651
rect 18090 -3346 18410 -2651
rect 18590 -3346 18910 -2651
rect 19090 -3346 19410 -2651
rect 19590 -3346 19910 -2651
rect 20090 -3346 20410 -2651
rect 20590 -3346 20910 -2651
rect 21090 -3346 21410 -2651
rect 21590 -3346 21910 -2651
rect 22370 -3346 22690 -2651
rect 28104 -3346 28424 -2651
rect 31112 -3346 31432 -2651
rect 57013 -3096 58818 -2651
rect 9493 -3509 9653 -3461
rect 9493 -3555 9550 -3509
rect 9596 -3555 9653 -3509
rect 9493 -3603 9653 -3555
rect 9493 -3649 9550 -3603
rect 9596 -3649 9653 -3603
rect 14200 -3444 14380 -3436
rect 14200 -3448 14668 -3444
rect 14200 -3500 14212 -3448
rect 14264 -3500 14316 -3448
rect 14368 -3500 14668 -3448
rect 14200 -3552 14668 -3500
rect 14200 -3604 14212 -3552
rect 14264 -3604 14316 -3552
rect 14368 -3604 14668 -3552
rect 17590 -3456 31432 -3346
rect 17590 -3502 17720 -3456
rect 17766 -3502 17814 -3456
rect 17860 -3502 17908 -3456
rect 17954 -3502 18002 -3456
rect 18048 -3502 18096 -3456
rect 18142 -3502 18190 -3456
rect 18236 -3502 18284 -3456
rect 18330 -3502 18378 -3456
rect 18424 -3502 18472 -3456
rect 18518 -3502 18566 -3456
rect 18612 -3502 18660 -3456
rect 18706 -3502 18754 -3456
rect 18800 -3502 18848 -3456
rect 18894 -3502 18942 -3456
rect 18988 -3502 19036 -3456
rect 19082 -3502 19130 -3456
rect 19176 -3502 19224 -3456
rect 19270 -3502 19318 -3456
rect 19364 -3502 19412 -3456
rect 19458 -3502 19506 -3456
rect 19552 -3502 19600 -3456
rect 19646 -3502 19694 -3456
rect 19740 -3502 19788 -3456
rect 19834 -3502 19882 -3456
rect 19928 -3502 19976 -3456
rect 20022 -3502 20070 -3456
rect 20116 -3502 20164 -3456
rect 20210 -3502 20258 -3456
rect 20304 -3502 20352 -3456
rect 20398 -3502 20446 -3456
rect 20492 -3502 20540 -3456
rect 20586 -3502 20634 -3456
rect 20680 -3502 20728 -3456
rect 20774 -3502 20822 -3456
rect 20868 -3502 20916 -3456
rect 20962 -3502 21010 -3456
rect 21056 -3502 21104 -3456
rect 21150 -3502 21198 -3456
rect 21244 -3502 21292 -3456
rect 21338 -3502 21386 -3456
rect 21432 -3502 21480 -3456
rect 21526 -3502 21574 -3456
rect 21620 -3502 21668 -3456
rect 21714 -3502 21762 -3456
rect 21808 -3502 21856 -3456
rect 21902 -3502 21950 -3456
rect 21996 -3502 22044 -3456
rect 22090 -3502 22138 -3456
rect 22184 -3502 22232 -3456
rect 22278 -3502 22326 -3456
rect 22372 -3502 22420 -3456
rect 22466 -3502 22514 -3456
rect 22560 -3502 22608 -3456
rect 22654 -3502 22702 -3456
rect 22748 -3502 22796 -3456
rect 22842 -3502 22890 -3456
rect 22936 -3502 22984 -3456
rect 23030 -3502 23078 -3456
rect 23124 -3502 23172 -3456
rect 23218 -3502 23266 -3456
rect 23312 -3502 23360 -3456
rect 23406 -3502 23454 -3456
rect 23500 -3502 23548 -3456
rect 23594 -3502 23642 -3456
rect 23688 -3502 23736 -3456
rect 23782 -3502 23830 -3456
rect 23876 -3502 23924 -3456
rect 23970 -3502 24018 -3456
rect 24064 -3502 24112 -3456
rect 24158 -3502 24206 -3456
rect 24252 -3502 24300 -3456
rect 24346 -3502 24394 -3456
rect 24440 -3502 24488 -3456
rect 24534 -3502 24582 -3456
rect 24628 -3502 24676 -3456
rect 24722 -3502 24770 -3456
rect 24816 -3502 24864 -3456
rect 24910 -3502 24958 -3456
rect 25004 -3502 25052 -3456
rect 25098 -3502 25146 -3456
rect 25192 -3502 25240 -3456
rect 25286 -3502 25334 -3456
rect 25380 -3502 25428 -3456
rect 25474 -3502 25522 -3456
rect 25568 -3502 25616 -3456
rect 25662 -3502 25710 -3456
rect 25756 -3502 25804 -3456
rect 25850 -3502 25898 -3456
rect 25944 -3502 25992 -3456
rect 26038 -3502 26086 -3456
rect 26132 -3502 26180 -3456
rect 26226 -3502 26274 -3456
rect 26320 -3502 26368 -3456
rect 26414 -3502 26462 -3456
rect 26508 -3502 26556 -3456
rect 26602 -3502 26650 -3456
rect 26696 -3502 26744 -3456
rect 26790 -3502 26838 -3456
rect 26884 -3502 26932 -3456
rect 26978 -3502 27026 -3456
rect 27072 -3502 27120 -3456
rect 27166 -3502 27214 -3456
rect 27260 -3502 27308 -3456
rect 27354 -3502 27402 -3456
rect 27448 -3502 27496 -3456
rect 27542 -3502 27590 -3456
rect 27636 -3502 27684 -3456
rect 27730 -3502 27778 -3456
rect 27824 -3502 27872 -3456
rect 27918 -3502 27966 -3456
rect 28012 -3502 28060 -3456
rect 28106 -3502 28154 -3456
rect 28200 -3502 28248 -3456
rect 28294 -3502 28342 -3456
rect 28388 -3502 28436 -3456
rect 28482 -3502 28530 -3456
rect 28576 -3502 28624 -3456
rect 28670 -3502 28718 -3456
rect 28764 -3502 28812 -3456
rect 28858 -3502 28906 -3456
rect 28952 -3502 29000 -3456
rect 29046 -3502 29094 -3456
rect 29140 -3502 29188 -3456
rect 29234 -3502 29282 -3456
rect 29328 -3502 29376 -3456
rect 29422 -3502 29470 -3456
rect 29516 -3502 29564 -3456
rect 29610 -3502 29658 -3456
rect 29704 -3502 29752 -3456
rect 29798 -3502 29846 -3456
rect 29892 -3502 29940 -3456
rect 29986 -3502 30034 -3456
rect 30080 -3502 30128 -3456
rect 30174 -3502 30222 -3456
rect 30268 -3502 30316 -3456
rect 30362 -3502 30410 -3456
rect 30456 -3502 30504 -3456
rect 30550 -3502 30598 -3456
rect 30644 -3502 30692 -3456
rect 30738 -3502 30786 -3456
rect 30832 -3502 30880 -3456
rect 30926 -3502 30974 -3456
rect 31020 -3502 31068 -3456
rect 31114 -3502 31162 -3456
rect 31208 -3502 31256 -3456
rect 31302 -3502 31432 -3456
rect 17590 -3550 31432 -3502
rect 17590 -3596 17720 -3550
rect 17766 -3596 22514 -3550
rect 22560 -3596 28248 -3550
rect 28294 -3596 31256 -3550
rect 31302 -3596 31432 -3550
rect 14200 -3616 14380 -3604
rect 9493 -3697 9653 -3649
rect 9493 -3743 9550 -3697
rect 9596 -3743 9653 -3697
rect 17590 -3644 31432 -3596
rect 54292 -3569 54491 -3556
rect 54292 -3625 54309 -3569
rect 54365 -3625 54419 -3569
rect 54475 -3579 54491 -3569
rect 54475 -3625 56701 -3579
rect 54292 -3642 54491 -3625
rect 17590 -3690 17720 -3644
rect 17766 -3666 22514 -3644
rect 17766 -3690 17910 -3666
rect 9493 -3791 9653 -3743
rect 9493 -3837 9550 -3791
rect 9596 -3837 9653 -3791
rect 9493 -3885 9653 -3837
rect 10058 -3711 10238 -3701
rect 16848 -3711 17028 -3701
rect 10058 -3713 17028 -3711
rect 10058 -3765 10070 -3713
rect 10122 -3765 10174 -3713
rect 10226 -3765 16860 -3713
rect 16912 -3765 16964 -3713
rect 17016 -3765 17028 -3713
rect 10058 -3817 17028 -3765
rect 10058 -3869 10070 -3817
rect 10122 -3869 10174 -3817
rect 10226 -3869 16860 -3817
rect 16912 -3869 16964 -3817
rect 17016 -3869 17028 -3817
rect 10058 -3871 17028 -3869
rect 10058 -3881 10238 -3871
rect 16848 -3881 17028 -3871
rect 17590 -3738 17910 -3690
rect 17590 -3784 17720 -3738
rect 17766 -3784 17910 -3738
rect 17590 -3832 17910 -3784
rect 17590 -3878 17720 -3832
rect 17766 -3878 17910 -3832
rect 9493 -3931 9550 -3885
rect 9596 -3931 9653 -3885
rect 9493 -3979 9653 -3931
rect 9493 -4025 9550 -3979
rect 9596 -4025 9653 -3979
rect 9493 -4073 9653 -4025
rect 9493 -4119 9550 -4073
rect 9596 -4119 9653 -4073
rect 9493 -4167 9653 -4119
rect 9493 -4213 9550 -4167
rect 9596 -4213 9653 -4167
rect 9493 -4261 9653 -4213
rect 9493 -4307 9550 -4261
rect 9596 -4307 9653 -4261
rect 9493 -4355 9653 -4307
rect 9493 -4401 9550 -4355
rect 9596 -4401 9653 -4355
rect 9493 -4449 9653 -4401
rect 9493 -4495 9550 -4449
rect 9596 -4495 9653 -4449
rect 9493 -4543 9653 -4495
rect 9493 -4589 9550 -4543
rect 9596 -4588 9653 -4543
rect 17590 -3926 17910 -3878
rect 17590 -3972 17720 -3926
rect 17766 -3972 17910 -3926
rect 17590 -4020 17910 -3972
rect 17590 -4066 17720 -4020
rect 17766 -4066 17910 -4020
rect 17590 -4114 17910 -4066
rect 17590 -4160 17720 -4114
rect 17766 -4160 17910 -4114
rect 17590 -4208 17910 -4160
rect 17590 -4254 17720 -4208
rect 17766 -4254 17910 -4208
rect 17590 -4302 17910 -4254
rect 17590 -4348 17720 -4302
rect 17766 -4348 17910 -4302
rect 17590 -4396 17910 -4348
rect 17590 -4442 17720 -4396
rect 17766 -4442 17910 -4396
rect 17590 -4490 17910 -4442
rect 17590 -4536 17720 -4490
rect 17766 -4536 17910 -4490
rect 17590 -4584 17910 -4536
rect 9596 -4589 17208 -4588
rect 9493 -4637 17208 -4589
rect 9493 -4683 9550 -4637
rect 9596 -4683 17208 -4637
rect 9493 -4688 17208 -4683
rect 9493 -4731 11528 -4688
rect 9493 -4777 9550 -4731
rect 9596 -4734 11528 -4731
rect 11574 -4734 11622 -4688
rect 11668 -4734 11716 -4688
rect 11762 -4734 11810 -4688
rect 11856 -4734 11904 -4688
rect 11950 -4734 11998 -4688
rect 12044 -4734 12092 -4688
rect 12138 -4734 12186 -4688
rect 12232 -4734 12280 -4688
rect 12326 -4734 12374 -4688
rect 12420 -4734 12468 -4688
rect 12514 -4734 12562 -4688
rect 12608 -4734 12656 -4688
rect 12702 -4734 12750 -4688
rect 12796 -4734 12844 -4688
rect 12890 -4734 12938 -4688
rect 12984 -4734 13032 -4688
rect 13078 -4734 13126 -4688
rect 13172 -4734 13220 -4688
rect 13266 -4734 13314 -4688
rect 13360 -4734 13408 -4688
rect 13454 -4734 13502 -4688
rect 13548 -4734 13596 -4688
rect 13642 -4734 13690 -4688
rect 13736 -4734 13784 -4688
rect 13830 -4734 13878 -4688
rect 13924 -4734 13972 -4688
rect 14018 -4734 14066 -4688
rect 14112 -4734 14160 -4688
rect 14206 -4734 14254 -4688
rect 14300 -4734 14348 -4688
rect 14394 -4734 14442 -4688
rect 14488 -4734 14536 -4688
rect 14582 -4734 14630 -4688
rect 14676 -4734 14724 -4688
rect 14770 -4734 14818 -4688
rect 14864 -4734 14912 -4688
rect 14958 -4734 15006 -4688
rect 15052 -4734 15100 -4688
rect 15146 -4734 15194 -4688
rect 15240 -4734 15288 -4688
rect 15334 -4734 15382 -4688
rect 15428 -4734 15476 -4688
rect 15522 -4734 15570 -4688
rect 15616 -4734 15664 -4688
rect 15710 -4734 15758 -4688
rect 15804 -4734 15852 -4688
rect 15898 -4734 15946 -4688
rect 15992 -4734 16040 -4688
rect 16086 -4734 16134 -4688
rect 16180 -4734 16228 -4688
rect 16274 -4734 16322 -4688
rect 16368 -4734 16416 -4688
rect 16462 -4734 16510 -4688
rect 16556 -4734 16604 -4688
rect 16650 -4734 16698 -4688
rect 16744 -4734 16792 -4688
rect 16838 -4734 16886 -4688
rect 16932 -4734 16980 -4688
rect 17026 -4734 17074 -4688
rect 17120 -4734 17208 -4688
rect 9596 -4777 17208 -4734
rect 9493 -4782 17208 -4777
rect 9493 -4825 11528 -4782
rect 9493 -4871 9550 -4825
rect 9596 -4828 11528 -4825
rect 11574 -4828 17074 -4782
rect 17120 -4828 17208 -4782
rect 9596 -4871 17208 -4828
rect 9493 -4876 17208 -4871
rect 9493 -4908 11528 -4876
rect 9493 -4919 9653 -4908
rect 9493 -4965 9550 -4919
rect 9596 -4965 9653 -4919
rect 9493 -5013 9653 -4965
rect 9493 -5059 9550 -5013
rect 9596 -5059 9653 -5013
rect 9493 -5107 9653 -5059
rect 9493 -5153 9550 -5107
rect 9596 -5153 9653 -5107
rect 9493 -5201 9653 -5153
rect 9493 -5247 9550 -5201
rect 9596 -5247 9653 -5201
rect 9493 -5295 9653 -5247
rect 9493 -5341 9550 -5295
rect 9596 -5341 9653 -5295
rect 9493 -5389 9653 -5341
rect 9493 -5435 9550 -5389
rect 9596 -5435 9653 -5389
rect 9493 -5483 9653 -5435
rect 9493 -5529 9550 -5483
rect 9596 -5529 9653 -5483
rect 9493 -5577 9653 -5529
rect 9493 -5623 9550 -5577
rect 9596 -5616 9653 -5577
rect 11440 -4922 11528 -4908
rect 11574 -4908 17074 -4876
rect 11574 -4922 11760 -4908
rect 11440 -4970 11760 -4922
rect 11440 -5016 11528 -4970
rect 11574 -5016 11760 -4970
rect 11440 -5064 11760 -5016
rect 11440 -5110 11528 -5064
rect 11574 -5110 11760 -5064
rect 11440 -5158 11760 -5110
rect 11440 -5204 11528 -5158
rect 11574 -5204 11760 -5158
rect 11440 -5252 11760 -5204
rect 11440 -5298 11528 -5252
rect 11574 -5298 11760 -5252
rect 11440 -5346 11760 -5298
rect 11440 -5392 11528 -5346
rect 11574 -5392 11760 -5346
rect 11440 -5440 11760 -5392
rect 11440 -5486 11528 -5440
rect 11574 -5486 11760 -5440
rect 11440 -5534 11760 -5486
rect 11440 -5580 11528 -5534
rect 11574 -5580 11760 -5534
rect 11440 -5616 11760 -5580
rect 9596 -5623 11760 -5616
rect 9493 -5628 11760 -5623
rect 9493 -5671 11528 -5628
rect 9493 -5717 9550 -5671
rect 9596 -5674 11528 -5671
rect 11574 -5674 11760 -5628
rect 9596 -5717 11760 -5674
rect 9493 -5722 11760 -5717
rect 9493 -5765 11528 -5722
rect 9493 -5811 9550 -5765
rect 9596 -5768 11528 -5765
rect 11574 -5768 11760 -5722
rect 9596 -5811 11760 -5768
rect 9493 -5816 11760 -5811
rect 9493 -5859 11528 -5816
rect 9493 -5905 9550 -5859
rect 9596 -5862 11528 -5859
rect 11574 -5862 11760 -5816
rect 9596 -5905 11760 -5862
rect 9493 -5910 11760 -5905
rect 9493 -5936 11528 -5910
rect 9493 -5953 9653 -5936
rect 9493 -5999 9550 -5953
rect 9596 -5999 9653 -5953
rect 9493 -6047 9653 -5999
rect 9493 -6093 9550 -6047
rect 9596 -6093 9653 -6047
rect 8623 -6172 8635 -6120
rect 8687 -6172 8699 -6120
rect 8623 -6224 8699 -6172
rect 8623 -6276 8635 -6224
rect 8687 -6276 8699 -6224
rect 5357 -6375 5414 -6329
rect 5460 -6375 5508 -6329
rect 5554 -6375 5602 -6329
rect 5648 -6375 5696 -6329
rect 5742 -6375 5790 -6329
rect 5836 -6375 5884 -6329
rect 5930 -6375 5978 -6329
rect 6024 -6375 6072 -6329
rect 6118 -6375 6166 -6329
rect 6212 -6375 6260 -6329
rect 6306 -6375 6354 -6329
rect 6400 -6375 6448 -6329
rect 6494 -6375 6551 -6329
rect 5357 -6423 6551 -6375
rect 7518 -6343 7564 -6297
rect 8478 -6343 8524 -6286
rect 8623 -6288 8699 -6276
rect 9493 -6141 9653 -6093
rect 9493 -6187 9550 -6141
rect 9596 -6187 9653 -6141
rect 9493 -6235 9653 -6187
rect 9493 -6281 9550 -6235
rect 9596 -6272 9653 -6235
rect 11440 -5956 11528 -5936
rect 11574 -5956 11760 -5910
rect 11440 -6004 11760 -5956
rect 11440 -6050 11528 -6004
rect 11574 -6050 11760 -6004
rect 11440 -6098 11760 -6050
rect 11440 -6144 11528 -6098
rect 11574 -6144 11760 -6098
rect 11440 -6192 11760 -6144
rect 11440 -6238 11528 -6192
rect 11574 -6238 11760 -6192
rect 11440 -6272 11760 -6238
rect 9596 -6281 11760 -6272
rect 9493 -6286 11760 -6281
rect 7518 -6389 8524 -6343
rect 9493 -6329 11528 -6286
rect 9493 -6375 9550 -6329
rect 9596 -6375 9644 -6329
rect 9690 -6375 9738 -6329
rect 9784 -6375 9832 -6329
rect 9878 -6375 9926 -6329
rect 9972 -6375 10020 -6329
rect 10066 -6375 10114 -6329
rect 10160 -6375 10208 -6329
rect 10254 -6375 10302 -6329
rect 10348 -6375 10396 -6329
rect 10442 -6375 10490 -6329
rect 10536 -6375 10584 -6329
rect 10630 -6332 11528 -6329
rect 11574 -6332 11760 -6286
rect 10630 -6375 11760 -6332
rect 9493 -6380 11760 -6375
rect 5357 -6469 5414 -6423
rect 5460 -6432 6551 -6423
rect 9493 -6423 11528 -6380
rect 9493 -6432 10584 -6423
rect 5460 -6469 5517 -6432
rect 5357 -6517 5517 -6469
rect 5357 -6563 5414 -6517
rect 5460 -6563 5517 -6517
rect 5357 -6611 5517 -6563
rect 5357 -6657 5414 -6611
rect 5460 -6657 5517 -6611
rect 5357 -6705 5517 -6657
rect 5357 -6751 5414 -6705
rect 5460 -6751 5517 -6705
rect 5357 -6799 5517 -6751
rect 5357 -6845 5414 -6799
rect 5460 -6845 5517 -6799
rect 5357 -6893 5517 -6845
rect 5357 -6939 5414 -6893
rect 5460 -6939 5517 -6893
rect 5357 -6987 5517 -6939
rect 5357 -7033 5414 -6987
rect 5460 -7033 5517 -6987
rect 5357 -7081 5517 -7033
rect 5357 -7127 5414 -7081
rect 5460 -7127 5517 -7081
rect 5357 -7175 5517 -7127
rect 5357 -7221 5414 -7175
rect 5460 -7221 5517 -7175
rect 5357 -7269 5517 -7221
rect 5357 -7315 5414 -7269
rect 5460 -7315 5517 -7269
rect 5357 -7363 5517 -7315
rect 5357 -7409 5414 -7363
rect 5460 -7409 5517 -7363
rect 5357 -7457 5517 -7409
rect 5357 -7503 5414 -7457
rect 5460 -7503 5517 -7457
rect 5357 -7551 5517 -7503
rect 5357 -7597 5414 -7551
rect 5460 -7597 5517 -7551
rect 5357 -7645 5517 -7597
rect 5357 -7691 5414 -7645
rect 5460 -7691 5517 -7645
rect 5357 -7739 5517 -7691
rect 3250 -14035 3847 -7758
rect 5357 -7785 5414 -7739
rect 5460 -7776 5517 -7739
rect 5663 -7124 5709 -6432
rect 5823 -7124 5869 -6432
rect 7427 -6482 7438 -6436
rect 7484 -6448 8398 -6436
rect 8444 -6448 8459 -6436
rect 7484 -6482 8395 -6448
rect 8383 -6500 8395 -6482
rect 8447 -6500 8459 -6448
rect 6898 -6518 7078 -6504
rect 8383 -6512 8459 -6500
rect 6898 -6570 6908 -6518
rect 6960 -6570 7012 -6518
rect 7064 -6570 7078 -6518
rect 6898 -6622 7078 -6570
rect 6898 -6638 6908 -6622
rect 6111 -6684 6191 -6638
rect 6237 -6684 6351 -6638
rect 6397 -6684 6477 -6638
rect 6111 -6741 6157 -6684
rect 6431 -6741 6477 -6684
rect 6591 -6684 6671 -6638
rect 6717 -6684 6831 -6638
rect 6877 -6674 6908 -6638
rect 6960 -6638 7012 -6622
rect 7064 -6638 7078 -6622
rect 9827 -6521 10007 -6509
rect 9827 -6573 9839 -6521
rect 9891 -6573 9943 -6521
rect 9995 -6573 10007 -6521
rect 9827 -6625 10007 -6573
rect 6960 -6674 6991 -6638
rect 7064 -6674 7151 -6638
rect 6877 -6684 6991 -6674
rect 7037 -6684 7151 -6674
rect 7197 -6684 7311 -6638
rect 7357 -6684 7471 -6638
rect 7517 -6684 7631 -6638
rect 7677 -6684 7791 -6638
rect 7837 -6684 7951 -6638
rect 7997 -6684 8111 -6638
rect 8157 -6684 8271 -6638
rect 8317 -6684 8431 -6638
rect 8477 -6684 8591 -6638
rect 8637 -6684 8751 -6638
rect 8797 -6684 8877 -6638
rect 6591 -6741 6637 -6684
rect 6911 -6741 6957 -6684
rect 7231 -6741 7277 -6684
rect 7551 -6741 7597 -6684
rect 7871 -6741 7917 -6684
rect 8191 -6741 8237 -6684
rect 8511 -6741 8557 -6684
rect 8831 -6741 8877 -6684
rect 9827 -6677 9839 -6625
rect 9891 -6677 9943 -6625
rect 9995 -6677 10007 -6625
rect 9827 -6689 10007 -6677
rect 9871 -6741 9917 -6689
rect 6096 -6757 6172 -6745
rect 6096 -6809 6108 -6757
rect 6160 -6809 6172 -6757
rect 6096 -6861 6172 -6809
rect 6096 -6913 6108 -6861
rect 6160 -6913 6172 -6861
rect 6096 -6925 6172 -6913
rect 9251 -6753 9431 -6741
rect 9251 -6805 9263 -6753
rect 9315 -6805 9367 -6753
rect 9419 -6805 9431 -6753
rect 9251 -6857 9431 -6805
rect 9251 -6909 9263 -6857
rect 9315 -6909 9367 -6857
rect 9419 -6909 9431 -6857
rect 5951 -6972 5997 -6925
rect 6271 -6972 6317 -6915
rect 6591 -6972 6637 -6915
rect 5951 -7018 6637 -6972
rect 6751 -6972 6797 -6915
rect 7071 -6972 7117 -6915
rect 7391 -6972 7437 -6915
rect 7711 -6972 7757 -6915
rect 8031 -6972 8077 -6915
rect 8351 -6972 8397 -6915
rect 8671 -6972 8717 -6915
rect 8959 -6972 9005 -6915
rect 9251 -6921 9431 -6909
rect 9567 -6972 9613 -6915
rect 10175 -6972 10221 -6432
rect 6751 -7018 10221 -6972
rect 5663 -7170 5743 -7124
rect 5789 -7170 5869 -7124
rect 10175 -7124 10221 -7018
rect 10335 -7124 10381 -6432
rect 5663 -7776 5709 -7170
rect 5823 -7776 5869 -7170
rect 8910 -7153 9090 -7141
rect 8910 -7205 8922 -7153
rect 8974 -7205 9026 -7153
rect 9078 -7205 9090 -7153
rect 6026 -7247 6206 -7233
rect 6026 -7299 6038 -7247
rect 6090 -7299 6142 -7247
rect 6194 -7299 6206 -7247
rect 8910 -7257 9090 -7205
rect 8910 -7264 8922 -7257
rect 6026 -7311 6206 -7299
rect 6383 -7321 7293 -7275
rect 7574 -7312 7585 -7266
rect 7631 -7312 7679 -7266
rect 7725 -7312 7773 -7266
rect 7819 -7312 7830 -7266
rect 8271 -7275 8922 -7264
rect 5936 -7386 6012 -7374
rect 6383 -7378 6429 -7321
rect 6815 -7378 6861 -7321
rect 7247 -7378 7293 -7321
rect 7679 -7378 7725 -7312
rect 8317 -7321 8431 -7275
rect 8477 -7321 8591 -7275
rect 8637 -7321 8751 -7275
rect 8797 -7321 8911 -7275
rect 8974 -7309 9026 -7257
rect 9078 -7264 9090 -7257
rect 10175 -7170 10255 -7124
rect 10301 -7170 10381 -7124
rect 9078 -7275 9277 -7264
rect 8957 -7321 9071 -7309
rect 9117 -7321 9277 -7275
rect 8271 -7378 8317 -7321
rect 8591 -7378 8637 -7321
rect 8911 -7378 8957 -7321
rect 9231 -7378 9277 -7321
rect 5936 -7438 5948 -7386
rect 6000 -7438 6012 -7386
rect 5936 -7490 6012 -7438
rect 5936 -7542 5948 -7490
rect 6000 -7542 6012 -7490
rect 5936 -7554 6012 -7542
rect 6368 -7392 6444 -7380
rect 6368 -7444 6380 -7392
rect 6432 -7444 6444 -7392
rect 6368 -7496 6444 -7444
rect 6368 -7548 6380 -7496
rect 6432 -7548 6444 -7496
rect 6167 -7776 6213 -7552
rect 6368 -7560 6444 -7548
rect 6599 -7776 6645 -7552
rect 7031 -7776 7077 -7552
rect 7463 -7776 7509 -7552
rect 7895 -7776 7941 -7552
rect 8111 -7609 8157 -7552
rect 8431 -7609 8477 -7552
rect 8751 -7609 8797 -7552
rect 9071 -7609 9117 -7552
rect 8111 -7655 9117 -7609
rect 9375 -7776 9421 -7552
rect 9535 -7776 9581 -7552
rect 9695 -7776 9741 -7552
rect 9855 -7776 9901 -7552
rect 10015 -7776 10061 -7552
rect 10175 -7776 10221 -7170
rect 10335 -7776 10381 -7170
rect 10527 -6469 10584 -6432
rect 10630 -6426 11528 -6423
rect 11574 -6426 11760 -6380
rect 10630 -6469 11760 -6426
rect 10527 -6474 11760 -6469
rect 10527 -6517 11528 -6474
rect 10527 -6563 10584 -6517
rect 10630 -6520 11528 -6517
rect 11574 -6520 11760 -6474
rect 10630 -6563 11760 -6520
rect 10527 -6568 11760 -6563
rect 10527 -6592 11528 -6568
rect 10527 -6611 10687 -6592
rect 10527 -6657 10584 -6611
rect 10630 -6657 10687 -6611
rect 10527 -6705 10687 -6657
rect 10527 -6751 10584 -6705
rect 10630 -6751 10687 -6705
rect 10527 -6799 10687 -6751
rect 10527 -6845 10584 -6799
rect 10630 -6845 10687 -6799
rect 10527 -6893 10687 -6845
rect 10527 -6939 10584 -6893
rect 10630 -6939 10687 -6893
rect 10527 -6987 10687 -6939
rect 10527 -7033 10584 -6987
rect 10630 -7033 10687 -6987
rect 10527 -7081 10687 -7033
rect 10527 -7127 10584 -7081
rect 10630 -7127 10687 -7081
rect 10527 -7175 10687 -7127
rect 11440 -6614 11528 -6592
rect 11574 -6614 11760 -6568
rect 11440 -6662 11760 -6614
rect 11440 -6708 11528 -6662
rect 11574 -6708 11760 -6662
rect 11440 -6756 11760 -6708
rect 11440 -6802 11528 -6756
rect 11574 -6802 11760 -6756
rect 11440 -6850 11760 -6802
rect 11440 -6896 11528 -6850
rect 11574 -6896 11760 -6850
rect 11440 -6944 11760 -6896
rect 11440 -6990 11528 -6944
rect 11574 -6990 11760 -6944
rect 11440 -7038 11760 -6990
rect 11440 -7084 11528 -7038
rect 11574 -7084 11760 -7038
rect 11440 -7132 11760 -7084
rect 10527 -7221 10584 -7175
rect 10630 -7221 10687 -7175
rect 10527 -7269 10687 -7221
rect 10527 -7315 10584 -7269
rect 10630 -7315 10687 -7269
rect 10527 -7363 10687 -7315
rect 10819 -7151 10999 -7141
rect 10819 -7153 11291 -7151
rect 10819 -7205 10831 -7153
rect 10883 -7205 10935 -7153
rect 10987 -7205 11291 -7153
rect 10819 -7257 11291 -7205
rect 10819 -7309 10831 -7257
rect 10883 -7309 10935 -7257
rect 10987 -7309 11291 -7257
rect 10819 -7311 11291 -7309
rect 11440 -7178 11528 -7132
rect 11574 -7178 11760 -7132
rect 11440 -7226 11760 -7178
rect 11440 -7272 11528 -7226
rect 11574 -7272 11760 -7226
rect 10819 -7321 10999 -7311
rect 11440 -7320 11760 -7272
rect 10527 -7409 10584 -7363
rect 10630 -7409 10687 -7363
rect 10527 -7457 10687 -7409
rect 10527 -7503 10584 -7457
rect 10630 -7503 10687 -7457
rect 10527 -7551 10687 -7503
rect 10527 -7597 10584 -7551
rect 10630 -7597 10687 -7551
rect 10527 -7616 10687 -7597
rect 11440 -7366 11528 -7320
rect 11574 -7366 11760 -7320
rect 11440 -7414 11760 -7366
rect 11440 -7460 11528 -7414
rect 11574 -7460 11760 -7414
rect 11440 -7508 11760 -7460
rect 11440 -7554 11528 -7508
rect 11574 -7554 11760 -7508
rect 11440 -7602 11760 -7554
rect 11440 -7616 11528 -7602
rect 10527 -7645 11528 -7616
rect 10527 -7691 10584 -7645
rect 10630 -7648 11528 -7645
rect 11574 -7616 11760 -7602
rect 12197 -6460 12243 -4908
rect 12501 -6460 12547 -4908
rect 12629 -5925 12675 -4908
rect 12723 -5156 12885 -4908
rect 12723 -5202 12734 -5156
rect 12780 -5202 12828 -5156
rect 12874 -5202 12885 -5156
rect 12723 -5250 12885 -5202
rect 12723 -5296 12734 -5250
rect 12780 -5296 12828 -5250
rect 12874 -5296 12885 -5250
rect 12723 -5307 12885 -5296
rect 12197 -6506 12302 -6460
rect 12348 -6506 12396 -6460
rect 12442 -6506 12547 -6460
rect 12197 -6554 12547 -6506
rect 12197 -6600 12302 -6554
rect 12348 -6600 12396 -6554
rect 12442 -6600 12547 -6554
rect 12197 -7616 12243 -6600
rect 12501 -7616 12547 -6600
rect 12933 -6761 12979 -4908
rect 13237 -6449 13283 -5763
rect 13132 -6495 13143 -6449
rect 13189 -6495 13237 -6449
rect 13283 -6495 13331 -6449
rect 13377 -6495 13388 -6449
rect 12614 -6863 12690 -6851
rect 12614 -6915 12626 -6863
rect 12678 -6915 12690 -6863
rect 12614 -6967 12690 -6915
rect 12614 -7019 12626 -6967
rect 12678 -7019 12690 -6967
rect 12614 -7071 12690 -7019
rect 12614 -7123 12626 -7071
rect 12678 -7123 12690 -7071
rect 12614 -7135 12690 -7123
rect 13237 -7325 13283 -7135
rect 12714 -7342 12894 -7330
rect 12714 -7394 12726 -7342
rect 12778 -7394 12830 -7342
rect 12882 -7394 12894 -7342
rect 13132 -7371 13143 -7325
rect 13189 -7371 13237 -7325
rect 13283 -7371 13331 -7325
rect 13377 -7371 13388 -7325
rect 12714 -7446 12894 -7394
rect 12714 -7498 12726 -7446
rect 12778 -7498 12830 -7446
rect 12882 -7498 12894 -7446
rect 12714 -7510 12894 -7498
rect 13541 -7616 13587 -4908
rect 13845 -6449 13891 -5763
rect 13740 -6495 13751 -6449
rect 13797 -6495 13845 -6449
rect 13891 -6495 13939 -6449
rect 13985 -6495 13996 -6449
rect 13845 -7310 13891 -7135
rect 13726 -7322 14010 -7310
rect 13726 -7374 13738 -7322
rect 13790 -7374 13842 -7322
rect 13894 -7374 13946 -7322
rect 13998 -7374 14010 -7322
rect 13726 -7386 14010 -7374
rect 14149 -7616 14195 -4908
rect 14566 -5595 14642 -5583
rect 14566 -5647 14578 -5595
rect 14630 -5647 14642 -5595
rect 14566 -5699 14642 -5647
rect 14566 -5751 14578 -5699
rect 14630 -5751 14642 -5699
rect 14566 -5763 14642 -5751
rect 14453 -6449 14499 -5763
rect 14581 -5925 14627 -5763
rect 14885 -6299 14931 -4908
rect 15174 -5595 15250 -5583
rect 15174 -5647 15186 -5595
rect 15238 -5647 15250 -5595
rect 15174 -5699 15250 -5647
rect 15174 -5751 15186 -5699
rect 15238 -5751 15250 -5699
rect 15174 -5763 15250 -5751
rect 15189 -5925 15235 -5763
rect 15493 -6299 15539 -4908
rect 15782 -5595 15858 -5583
rect 15782 -5647 15794 -5595
rect 15846 -5647 15858 -5595
rect 15782 -5699 15858 -5647
rect 15782 -5751 15794 -5699
rect 15846 -5751 15858 -5699
rect 15782 -5763 15858 -5751
rect 15797 -5925 15843 -5763
rect 15685 -6394 15969 -6372
rect 15685 -6446 15697 -6394
rect 15749 -6446 15801 -6394
rect 15853 -6446 15905 -6394
rect 15957 -6446 15969 -6394
rect 14348 -6495 14359 -6449
rect 14405 -6495 14453 -6449
rect 14499 -6495 14547 -6449
rect 14593 -6495 14604 -6449
rect 15685 -6498 15969 -6446
rect 15685 -6550 15697 -6498
rect 15749 -6550 15801 -6498
rect 15853 -6550 15905 -6498
rect 15957 -6550 15969 -6498
rect 15685 -6572 15969 -6550
rect 16101 -6460 16147 -4908
rect 16405 -6460 16451 -4908
rect 16101 -6506 16206 -6460
rect 16252 -6506 16300 -6460
rect 16346 -6506 16451 -6460
rect 16101 -6554 16451 -6506
rect 16101 -6600 16206 -6554
rect 16252 -6600 16300 -6554
rect 16346 -6600 16451 -6554
rect 14581 -6704 15843 -6658
rect 14581 -6761 14627 -6704
rect 15189 -6761 15235 -6704
rect 15797 -6761 15843 -6704
rect 14453 -7325 14499 -7135
rect 14348 -7371 14359 -7325
rect 14405 -7371 14453 -7325
rect 14499 -7371 14547 -7325
rect 14593 -7371 14604 -7325
rect 14885 -7616 14931 -6761
rect 15174 -6863 15250 -6851
rect 15174 -6915 15186 -6863
rect 15238 -6915 15250 -6863
rect 15174 -6967 15250 -6915
rect 15174 -7019 15186 -6967
rect 15238 -7019 15250 -6967
rect 15174 -7071 15250 -7019
rect 15174 -7123 15186 -7071
rect 15238 -7123 15250 -7071
rect 15174 -7135 15250 -7123
rect 15493 -7616 15539 -6761
rect 16101 -7616 16147 -6600
rect 16405 -7616 16451 -6600
rect 16888 -4922 17074 -4908
rect 17120 -4922 17208 -4876
rect 16888 -4970 17208 -4922
rect 16888 -5016 17074 -4970
rect 17120 -5016 17208 -4970
rect 16888 -5064 17208 -5016
rect 16888 -5110 17074 -5064
rect 17120 -5110 17208 -5064
rect 16888 -5158 17208 -5110
rect 16888 -5204 17074 -5158
rect 17120 -5204 17208 -5158
rect 16888 -5252 17208 -5204
rect 16888 -5298 17074 -5252
rect 17120 -5298 17208 -5252
rect 16888 -5346 17208 -5298
rect 16888 -5392 17074 -5346
rect 17120 -5392 17208 -5346
rect 16888 -5440 17208 -5392
rect 16888 -5486 17074 -5440
rect 17120 -5486 17208 -5440
rect 16888 -5534 17208 -5486
rect 16888 -5580 17074 -5534
rect 17120 -5580 17208 -5534
rect 16888 -5628 17208 -5580
rect 16888 -5674 17074 -5628
rect 17120 -5674 17208 -5628
rect 16888 -5722 17208 -5674
rect 16888 -5768 17074 -5722
rect 17120 -5768 17208 -5722
rect 16888 -5816 17208 -5768
rect 16888 -5862 17074 -5816
rect 17120 -5862 17208 -5816
rect 16888 -5910 17208 -5862
rect 16888 -5956 17074 -5910
rect 17120 -5956 17208 -5910
rect 16888 -6004 17208 -5956
rect 16888 -6050 17074 -6004
rect 17120 -6050 17208 -6004
rect 16888 -6098 17208 -6050
rect 16888 -6144 17074 -6098
rect 17120 -6144 17208 -6098
rect 16888 -6192 17208 -6144
rect 16888 -6238 17074 -6192
rect 17120 -6238 17208 -6192
rect 16888 -6286 17208 -6238
rect 16888 -6332 17074 -6286
rect 17120 -6332 17208 -6286
rect 16888 -6380 17208 -6332
rect 16888 -6426 17074 -6380
rect 17120 -6426 17208 -6380
rect 16888 -6474 17208 -6426
rect 16888 -6520 17074 -6474
rect 17120 -6520 17208 -6474
rect 16888 -6568 17208 -6520
rect 16888 -6614 17074 -6568
rect 17120 -6614 17208 -6568
rect 16888 -6662 17208 -6614
rect 16888 -6708 17074 -6662
rect 17120 -6708 17208 -6662
rect 16888 -6756 17208 -6708
rect 16888 -6802 17074 -6756
rect 17120 -6802 17208 -6756
rect 16888 -6850 17208 -6802
rect 16888 -6896 17074 -6850
rect 17120 -6896 17208 -6850
rect 16888 -6944 17208 -6896
rect 16888 -6990 17074 -6944
rect 17120 -6990 17208 -6944
rect 16888 -7038 17208 -6990
rect 16888 -7084 17074 -7038
rect 17120 -7084 17208 -7038
rect 16888 -7132 17208 -7084
rect 16888 -7178 17074 -7132
rect 17120 -7178 17208 -7132
rect 16888 -7226 17208 -7178
rect 16888 -7272 17074 -7226
rect 17120 -7272 17208 -7226
rect 16888 -7320 17208 -7272
rect 16888 -7366 17074 -7320
rect 17120 -7366 17208 -7320
rect 16888 -7414 17208 -7366
rect 16888 -7460 17074 -7414
rect 17120 -7460 17208 -7414
rect 16888 -7508 17208 -7460
rect 16888 -7554 17074 -7508
rect 17120 -7554 17208 -7508
rect 16888 -7602 17208 -7554
rect 16888 -7616 17074 -7602
rect 11574 -7648 17074 -7616
rect 17120 -7648 17208 -7602
rect 10630 -7691 17208 -7648
rect 10527 -7696 17208 -7691
rect 10527 -7739 11528 -7696
rect 10527 -7776 10584 -7739
rect 5460 -7785 10584 -7776
rect 10630 -7742 11528 -7739
rect 11574 -7742 17074 -7696
rect 17120 -7742 17208 -7696
rect 10630 -7785 17208 -7742
rect 5357 -7790 17208 -7785
rect 5357 -7833 11528 -7790
rect 5357 -7879 5414 -7833
rect 5460 -7879 5508 -7833
rect 5554 -7879 5602 -7833
rect 5648 -7879 5696 -7833
rect 5742 -7879 5790 -7833
rect 5836 -7879 5884 -7833
rect 5930 -7879 5978 -7833
rect 6024 -7879 6072 -7833
rect 6118 -7879 6166 -7833
rect 6212 -7879 6260 -7833
rect 6306 -7879 6354 -7833
rect 6400 -7879 6448 -7833
rect 6494 -7879 6542 -7833
rect 6588 -7879 6636 -7833
rect 6682 -7879 6730 -7833
rect 6776 -7879 6824 -7833
rect 6870 -7879 6918 -7833
rect 6964 -7879 7012 -7833
rect 7058 -7879 7106 -7833
rect 7152 -7879 7200 -7833
rect 7246 -7879 7294 -7833
rect 7340 -7879 7388 -7833
rect 7434 -7879 7482 -7833
rect 7528 -7879 7576 -7833
rect 7622 -7879 7670 -7833
rect 7716 -7879 7764 -7833
rect 7810 -7879 7858 -7833
rect 7904 -7879 7952 -7833
rect 7998 -7879 8046 -7833
rect 8092 -7879 8140 -7833
rect 8186 -7879 8234 -7833
rect 8280 -7879 8328 -7833
rect 8374 -7879 8422 -7833
rect 8468 -7879 8516 -7833
rect 8562 -7879 8610 -7833
rect 8656 -7879 8704 -7833
rect 8750 -7879 8798 -7833
rect 8844 -7879 8892 -7833
rect 8938 -7879 8986 -7833
rect 9032 -7879 9080 -7833
rect 9126 -7879 9174 -7833
rect 9220 -7879 9268 -7833
rect 9314 -7879 9362 -7833
rect 9408 -7879 9456 -7833
rect 9502 -7879 9550 -7833
rect 9596 -7879 9644 -7833
rect 9690 -7879 9738 -7833
rect 9784 -7879 9832 -7833
rect 9878 -7879 9926 -7833
rect 9972 -7879 10020 -7833
rect 10066 -7879 10114 -7833
rect 10160 -7879 10208 -7833
rect 10254 -7879 10302 -7833
rect 10348 -7879 10396 -7833
rect 10442 -7879 10490 -7833
rect 10536 -7879 10584 -7833
rect 10630 -7836 11528 -7833
rect 11574 -7836 11622 -7790
rect 11668 -7836 11716 -7790
rect 11762 -7836 11810 -7790
rect 11856 -7836 11904 -7790
rect 11950 -7836 11998 -7790
rect 12044 -7836 12092 -7790
rect 12138 -7836 12186 -7790
rect 12232 -7836 12280 -7790
rect 12326 -7836 12374 -7790
rect 12420 -7836 12468 -7790
rect 12514 -7836 12562 -7790
rect 12608 -7836 12656 -7790
rect 12702 -7836 12750 -7790
rect 12796 -7836 12844 -7790
rect 12890 -7836 12938 -7790
rect 12984 -7836 13032 -7790
rect 13078 -7836 13126 -7790
rect 13172 -7836 13220 -7790
rect 13266 -7836 13314 -7790
rect 13360 -7836 13408 -7790
rect 13454 -7836 13502 -7790
rect 13548 -7836 13596 -7790
rect 13642 -7836 13690 -7790
rect 13736 -7836 13784 -7790
rect 13830 -7836 13878 -7790
rect 13924 -7836 13972 -7790
rect 14018 -7836 14066 -7790
rect 14112 -7836 14160 -7790
rect 14206 -7836 14254 -7790
rect 14300 -7836 14348 -7790
rect 14394 -7836 14442 -7790
rect 14488 -7836 14536 -7790
rect 14582 -7836 14630 -7790
rect 14676 -7836 14724 -7790
rect 14770 -7836 14818 -7790
rect 14864 -7836 14912 -7790
rect 14958 -7836 15006 -7790
rect 15052 -7836 15100 -7790
rect 15146 -7836 15194 -7790
rect 15240 -7836 15288 -7790
rect 15334 -7836 15382 -7790
rect 15428 -7836 15476 -7790
rect 15522 -7836 15570 -7790
rect 15616 -7836 15664 -7790
rect 15710 -7836 15758 -7790
rect 15804 -7836 15852 -7790
rect 15898 -7836 15946 -7790
rect 15992 -7836 16040 -7790
rect 16086 -7836 16134 -7790
rect 16180 -7836 16228 -7790
rect 16274 -7836 16322 -7790
rect 16368 -7836 16416 -7790
rect 16462 -7836 16510 -7790
rect 16556 -7836 16604 -7790
rect 16650 -7836 16698 -7790
rect 16744 -7836 16792 -7790
rect 16838 -7836 16886 -7790
rect 16932 -7836 16980 -7790
rect 17026 -7836 17074 -7790
rect 17120 -7836 17208 -7790
rect 10630 -7879 17208 -7836
rect 5357 -7936 17208 -7879
rect 17590 -4630 17720 -4584
rect 17766 -4630 17910 -4584
rect 17590 -4678 17910 -4630
rect 17590 -4724 17720 -4678
rect 17766 -4724 17910 -4678
rect 17590 -4772 17910 -4724
rect 17590 -4818 17720 -4772
rect 17766 -4818 17910 -4772
rect 17590 -4866 17910 -4818
rect 17590 -4912 17720 -4866
rect 17766 -4912 17910 -4866
rect 17590 -4960 17910 -4912
rect 17590 -5006 17720 -4960
rect 17766 -5006 17910 -4960
rect 17590 -5054 17910 -5006
rect 17590 -5100 17720 -5054
rect 17766 -5100 17910 -5054
rect 17590 -5148 17910 -5100
rect 17590 -5194 17720 -5148
rect 17766 -5194 17910 -5148
rect 17590 -5242 17910 -5194
rect 17590 -5288 17720 -5242
rect 17766 -5288 17910 -5242
rect 17590 -5336 17910 -5288
rect 17590 -5382 17720 -5336
rect 17766 -5382 17910 -5336
rect 17590 -5430 17910 -5382
rect 17590 -5476 17720 -5430
rect 17766 -5476 17910 -5430
rect 17590 -5524 17910 -5476
rect 17590 -5570 17720 -5524
rect 17766 -5570 17910 -5524
rect 17590 -5618 17910 -5570
rect 17590 -5664 17720 -5618
rect 17766 -5664 17910 -5618
rect 17590 -5712 17910 -5664
rect 17590 -5758 17720 -5712
rect 17766 -5758 17910 -5712
rect 17590 -5806 17910 -5758
rect 17590 -5852 17720 -5806
rect 17766 -5852 17910 -5806
rect 17590 -5900 17910 -5852
rect 17590 -5946 17720 -5900
rect 17766 -5946 17910 -5900
rect 17590 -5994 17910 -5946
rect 17590 -6040 17720 -5994
rect 17766 -6040 17910 -5994
rect 17590 -6088 17910 -6040
rect 17590 -6134 17720 -6088
rect 17766 -6134 17910 -6088
rect 17590 -6182 17910 -6134
rect 17590 -6228 17720 -6182
rect 17766 -6228 17910 -6182
rect 17590 -6276 17910 -6228
rect 17590 -6322 17720 -6276
rect 17766 -6322 17910 -6276
rect 17590 -6370 17910 -6322
rect 17590 -6416 17720 -6370
rect 17766 -6416 17910 -6370
rect 17590 -6464 17910 -6416
rect 17590 -6510 17720 -6464
rect 17766 -6510 17910 -6464
rect 17590 -6558 17910 -6510
rect 17590 -6604 17720 -6558
rect 17766 -6604 17910 -6558
rect 17590 -6652 17910 -6604
rect 17590 -6698 17720 -6652
rect 17766 -6698 17910 -6652
rect 17590 -6746 17910 -6698
rect 17590 -6792 17720 -6746
rect 17766 -6792 17910 -6746
rect 17590 -6840 17910 -6792
rect 17590 -6886 17720 -6840
rect 17766 -6886 17910 -6840
rect 17590 -6934 17910 -6886
rect 17590 -6980 17720 -6934
rect 17766 -6980 17910 -6934
rect 17590 -7028 17910 -6980
rect 17590 -7074 17720 -7028
rect 17766 -7074 17910 -7028
rect 17590 -7122 17910 -7074
rect 17590 -7168 17720 -7122
rect 17766 -7168 17910 -7122
rect 17590 -7216 17910 -7168
rect 17590 -7262 17720 -7216
rect 17766 -7262 17910 -7216
rect 17590 -7310 17910 -7262
rect 17590 -7356 17720 -7310
rect 17766 -7356 17910 -7310
rect 17590 -7404 17910 -7356
rect 17590 -7450 17720 -7404
rect 17766 -7450 17910 -7404
rect 17590 -7498 17910 -7450
rect 17590 -7544 17720 -7498
rect 17766 -7544 17910 -7498
rect 17590 -7592 17910 -7544
rect 17590 -7638 17720 -7592
rect 17766 -7638 17910 -7592
rect 17590 -7686 17910 -7638
rect 17590 -7732 17720 -7686
rect 17766 -7732 17910 -7686
rect 17590 -7780 17910 -7732
rect 17590 -7826 17720 -7780
rect 17766 -7826 17910 -7780
rect 17590 -7874 17910 -7826
rect 17590 -7920 17720 -7874
rect 17766 -7898 17910 -7874
rect 18309 -5023 18355 -3666
rect 18469 -5023 18515 -3666
rect 18309 -5069 18389 -5023
rect 18435 -5069 18515 -5023
rect 18309 -6495 18355 -5069
rect 18469 -6495 18515 -5069
rect 18309 -6541 18389 -6495
rect 18435 -6541 18515 -6495
rect 18309 -7898 18355 -6541
rect 18469 -7898 18515 -6541
rect 18629 -6599 18675 -4965
rect 18789 -6599 18835 -3666
rect 18949 -6599 18995 -4965
rect 19109 -6599 19155 -3666
rect 19269 -6599 19315 -4965
rect 19429 -6599 19475 -3666
rect 19589 -6599 19635 -4965
rect 19749 -6599 19795 -3666
rect 19909 -6599 19955 -4965
rect 20069 -6599 20115 -3666
rect 20161 -4239 20341 -4227
rect 20161 -4291 20173 -4239
rect 20225 -4291 20277 -4239
rect 20329 -4291 20341 -4239
rect 20161 -4303 20341 -4291
rect 20229 -6599 20275 -4965
rect 20389 -6599 20435 -3666
rect 20549 -6599 20595 -4965
rect 18614 -6901 18690 -6889
rect 18614 -6953 18626 -6901
rect 18678 -6953 18690 -6901
rect 18614 -7005 18690 -6953
rect 18614 -7057 18626 -7005
rect 18678 -7057 18690 -7005
rect 18614 -7109 18690 -7057
rect 18614 -7161 18626 -7109
rect 18678 -7161 18690 -7109
rect 18614 -7173 18690 -7161
rect 18934 -6901 19010 -6889
rect 18934 -6953 18946 -6901
rect 18998 -6953 19010 -6901
rect 18934 -7005 19010 -6953
rect 18934 -7057 18946 -7005
rect 18998 -7057 19010 -7005
rect 18934 -7109 19010 -7057
rect 18934 -7161 18946 -7109
rect 18998 -7161 19010 -7109
rect 18934 -7173 19010 -7161
rect 19254 -6901 19330 -6889
rect 19254 -6953 19266 -6901
rect 19318 -6953 19330 -6901
rect 19254 -7005 19330 -6953
rect 19254 -7057 19266 -7005
rect 19318 -7057 19330 -7005
rect 19254 -7109 19330 -7057
rect 19254 -7161 19266 -7109
rect 19318 -7161 19330 -7109
rect 19254 -7173 19330 -7161
rect 19574 -6901 19650 -6889
rect 19574 -6953 19586 -6901
rect 19638 -6953 19650 -6901
rect 19574 -7005 19650 -6953
rect 19574 -7057 19586 -7005
rect 19638 -7057 19650 -7005
rect 19574 -7109 19650 -7057
rect 19574 -7161 19586 -7109
rect 19638 -7161 19650 -7109
rect 19574 -7173 19650 -7161
rect 19894 -6901 19970 -6889
rect 19894 -6953 19906 -6901
rect 19958 -6953 19970 -6901
rect 19894 -7005 19970 -6953
rect 19894 -7057 19906 -7005
rect 19958 -7057 19970 -7005
rect 19894 -7109 19970 -7057
rect 19894 -7161 19906 -7109
rect 19958 -7161 19970 -7109
rect 19894 -7173 19970 -7161
rect 20214 -6901 20290 -6889
rect 20214 -6953 20226 -6901
rect 20278 -6953 20290 -6901
rect 20214 -7005 20290 -6953
rect 20214 -7057 20226 -7005
rect 20278 -7057 20290 -7005
rect 20214 -7109 20290 -7057
rect 20214 -7161 20226 -7109
rect 20278 -7161 20290 -7109
rect 20214 -7173 20290 -7161
rect 20534 -6901 20610 -6889
rect 20534 -6953 20546 -6901
rect 20598 -6953 20610 -6901
rect 20534 -7005 20610 -6953
rect 20534 -7057 20546 -7005
rect 20598 -7057 20610 -7005
rect 20534 -7109 20610 -7057
rect 20534 -7161 20546 -7109
rect 20598 -7161 20610 -7109
rect 20534 -7173 20610 -7161
rect 18629 -7260 18675 -7173
rect 18949 -7260 18995 -7173
rect 19269 -7260 19315 -7173
rect 19589 -7260 19635 -7173
rect 19909 -7260 19955 -7173
rect 20229 -7260 20275 -7173
rect 20549 -7260 20595 -7173
rect 18629 -7306 20595 -7260
rect 20709 -7898 20755 -3666
rect 20869 -4242 20915 -4231
rect 20869 -4391 20915 -4288
rect 20869 -6599 20915 -4965
rect 21029 -7898 21075 -3666
rect 21174 -4693 21250 -4681
rect 21174 -4745 21186 -4693
rect 21238 -4745 21250 -4693
rect 21174 -4797 21250 -4745
rect 21174 -4849 21186 -4797
rect 21238 -4849 21250 -4797
rect 21174 -4901 21250 -4849
rect 21174 -4953 21186 -4901
rect 21238 -4953 21250 -4901
rect 21174 -4965 21250 -4953
rect 21189 -6599 21235 -4965
rect 21349 -6599 21395 -3666
rect 21477 -5023 21523 -3666
rect 21637 -5023 21683 -3666
rect 21477 -5069 21557 -5023
rect 21603 -5069 21683 -5023
rect 21477 -5127 21523 -5069
rect 21477 -6699 21523 -6437
rect 21145 -7253 21429 -7241
rect 21145 -7305 21157 -7253
rect 21209 -7305 21261 -7253
rect 21313 -7305 21365 -7253
rect 21417 -7305 21429 -7253
rect 21145 -7315 21429 -7305
rect 21477 -7256 21523 -7173
rect 21477 -7313 21523 -7302
rect 21637 -7898 21683 -5069
rect 21765 -5023 21811 -3666
rect 21925 -5023 21971 -3666
rect 21765 -5069 21845 -5023
rect 21891 -5069 21971 -5023
rect 21765 -6495 21811 -5069
rect 21925 -6495 21971 -5069
rect 21765 -6541 21845 -6495
rect 21891 -6541 21971 -6495
rect 21765 -7898 21811 -6541
rect 21925 -7898 21971 -6541
rect 22370 -3690 22514 -3666
rect 22560 -3666 28248 -3644
rect 22560 -3690 22690 -3666
rect 22370 -3738 22690 -3690
rect 22370 -3784 22514 -3738
rect 22560 -3784 22690 -3738
rect 22370 -3832 22690 -3784
rect 22370 -3878 22514 -3832
rect 22560 -3878 22690 -3832
rect 22370 -3926 22690 -3878
rect 22370 -3972 22514 -3926
rect 22560 -3972 22690 -3926
rect 22370 -4020 22690 -3972
rect 22370 -4066 22514 -4020
rect 22560 -4066 22690 -4020
rect 22370 -4114 22690 -4066
rect 22370 -4160 22514 -4114
rect 22560 -4160 22690 -4114
rect 22370 -4208 22690 -4160
rect 22370 -4254 22514 -4208
rect 22560 -4254 22690 -4208
rect 22370 -4302 22690 -4254
rect 22370 -4348 22514 -4302
rect 22560 -4348 22690 -4302
rect 22370 -4396 22690 -4348
rect 22370 -4442 22514 -4396
rect 22560 -4442 22690 -4396
rect 22370 -4490 22690 -4442
rect 22370 -4536 22514 -4490
rect 22560 -4536 22690 -4490
rect 22370 -4584 22690 -4536
rect 22370 -4630 22514 -4584
rect 22560 -4630 22690 -4584
rect 22370 -4678 22690 -4630
rect 22370 -4724 22514 -4678
rect 22560 -4724 22690 -4678
rect 22370 -4772 22690 -4724
rect 22370 -4818 22514 -4772
rect 22560 -4818 22690 -4772
rect 22370 -4866 22690 -4818
rect 22370 -4912 22514 -4866
rect 22560 -4912 22690 -4866
rect 22370 -4960 22690 -4912
rect 22370 -5006 22514 -4960
rect 22560 -5006 22690 -4960
rect 22370 -5054 22690 -5006
rect 22370 -5100 22514 -5054
rect 22560 -5100 22690 -5054
rect 22370 -5148 22690 -5100
rect 22370 -5194 22514 -5148
rect 22560 -5194 22690 -5148
rect 22370 -5242 22690 -5194
rect 22370 -5288 22514 -5242
rect 22560 -5288 22690 -5242
rect 22370 -5336 22690 -5288
rect 22370 -5382 22514 -5336
rect 22560 -5382 22690 -5336
rect 22370 -5430 22690 -5382
rect 22370 -5476 22514 -5430
rect 22560 -5476 22690 -5430
rect 22370 -5524 22690 -5476
rect 22370 -5570 22514 -5524
rect 22560 -5570 22690 -5524
rect 22370 -5618 22690 -5570
rect 22370 -5664 22514 -5618
rect 22560 -5664 22690 -5618
rect 22370 -5712 22690 -5664
rect 22370 -5758 22514 -5712
rect 22560 -5758 22690 -5712
rect 22370 -5806 22690 -5758
rect 22370 -5852 22514 -5806
rect 22560 -5852 22690 -5806
rect 22370 -5900 22690 -5852
rect 22370 -5946 22514 -5900
rect 22560 -5946 22690 -5900
rect 22370 -5994 22690 -5946
rect 22370 -6040 22514 -5994
rect 22560 -6040 22690 -5994
rect 22370 -6088 22690 -6040
rect 22370 -6134 22514 -6088
rect 22560 -6134 22690 -6088
rect 22370 -6182 22690 -6134
rect 22370 -6228 22514 -6182
rect 22560 -6228 22690 -6182
rect 22370 -6276 22690 -6228
rect 22370 -6322 22514 -6276
rect 22560 -6322 22690 -6276
rect 22370 -6370 22690 -6322
rect 22370 -6416 22514 -6370
rect 22560 -6416 22690 -6370
rect 22370 -6464 22690 -6416
rect 22370 -6510 22514 -6464
rect 22560 -6510 22690 -6464
rect 22370 -6558 22690 -6510
rect 22370 -6604 22514 -6558
rect 22560 -6604 22690 -6558
rect 22370 -6652 22690 -6604
rect 22370 -6698 22514 -6652
rect 22560 -6698 22690 -6652
rect 22370 -6746 22690 -6698
rect 22370 -6792 22514 -6746
rect 22560 -6792 22690 -6746
rect 22370 -6840 22690 -6792
rect 22370 -6886 22514 -6840
rect 22560 -6886 22690 -6840
rect 22370 -6934 22690 -6886
rect 22370 -6980 22514 -6934
rect 22560 -6980 22690 -6934
rect 22370 -7028 22690 -6980
rect 22370 -7074 22514 -7028
rect 22560 -7074 22690 -7028
rect 22370 -7122 22690 -7074
rect 22370 -7168 22514 -7122
rect 22560 -7168 22690 -7122
rect 22370 -7216 22690 -7168
rect 22370 -7262 22514 -7216
rect 22560 -7262 22690 -7216
rect 22370 -7310 22690 -7262
rect 22370 -7356 22514 -7310
rect 22560 -7356 22690 -7310
rect 22370 -7404 22690 -7356
rect 22370 -7450 22514 -7404
rect 22560 -7450 22690 -7404
rect 22370 -7498 22690 -7450
rect 22370 -7544 22514 -7498
rect 22560 -7544 22690 -7498
rect 22370 -7592 22690 -7544
rect 22370 -7638 22514 -7592
rect 22560 -7638 22690 -7592
rect 22370 -7686 22690 -7638
rect 22370 -7732 22514 -7686
rect 22560 -7732 22690 -7686
rect 22370 -7780 22690 -7732
rect 22370 -7826 22514 -7780
rect 22560 -7826 22690 -7780
rect 22370 -7874 22690 -7826
rect 22370 -7898 22514 -7874
rect 17766 -7920 22514 -7898
rect 22560 -7898 22690 -7874
rect 23176 -7898 23372 -3666
rect 23632 -4144 23812 -4132
rect 23632 -4196 23644 -4144
rect 23696 -4196 23748 -4144
rect 23800 -4196 23812 -4144
rect 23632 -4248 23812 -4196
rect 23632 -4300 23644 -4248
rect 23696 -4300 23748 -4248
rect 23800 -4300 23812 -4248
rect 24352 -4160 25724 -3964
rect 23820 -4297 24268 -4251
rect 24352 -4297 24548 -4160
rect 24800 -4297 25276 -4251
rect 25528 -4297 25724 -4160
rect 25808 -4160 27180 -3964
rect 25808 -4297 26004 -4160
rect 26256 -4297 26732 -4251
rect 26984 -4297 27180 -4160
rect 23632 -4312 23812 -4300
rect 26994 -4852 27174 -4840
rect 26556 -4904 27006 -4852
rect 27058 -4904 27110 -4852
rect 27162 -4904 27174 -4852
rect 26556 -4956 27174 -4904
rect 26556 -5008 27006 -4956
rect 27058 -5008 27110 -4956
rect 27162 -5008 27174 -4956
rect 26556 -5383 26716 -5008
rect 26994 -5020 27174 -5008
rect 23624 -5520 23820 -5383
rect 24072 -5429 24548 -5383
rect 24800 -5520 24996 -5383
rect 23624 -5716 24996 -5520
rect 25080 -5520 25276 -5383
rect 25528 -5429 26004 -5383
rect 26256 -5520 26452 -5383
rect 26536 -5429 26732 -5383
rect 25080 -5716 26452 -5520
rect 26984 -5736 27180 -5383
rect 26536 -5932 27180 -5736
rect 23624 -6132 24996 -5936
rect 23624 -6269 23820 -6132
rect 24072 -6269 24548 -6223
rect 24800 -6269 24996 -6132
rect 25080 -6132 26452 -5936
rect 25080 -6269 25276 -6132
rect 25528 -6269 26004 -6223
rect 26256 -6269 26452 -6132
rect 26536 -6269 26732 -5932
rect 26992 -6220 27172 -6208
rect 26992 -6272 27004 -6220
rect 27056 -6272 27108 -6220
rect 27160 -6272 27172 -6220
rect 26992 -6324 27172 -6272
rect 26992 -6376 27004 -6324
rect 27056 -6376 27108 -6324
rect 27160 -6376 27172 -6324
rect 26992 -6388 27172 -6376
rect 23632 -7352 23812 -7340
rect 23632 -7404 23644 -7352
rect 23696 -7404 23748 -7352
rect 23800 -7404 23812 -7352
rect 23632 -7456 23812 -7404
rect 23632 -7508 23644 -7456
rect 23696 -7508 23748 -7456
rect 23800 -7508 23812 -7456
rect 23632 -7520 23812 -7508
rect 24082 -7352 24262 -7338
rect 24082 -7404 24092 -7352
rect 24144 -7404 24196 -7352
rect 24248 -7404 24262 -7352
rect 24082 -7456 24262 -7404
rect 24082 -7508 24092 -7456
rect 24144 -7508 24196 -7456
rect 24248 -7508 24262 -7456
rect 24082 -7518 24262 -7508
rect 24352 -7492 24548 -7355
rect 24800 -7401 25276 -7355
rect 25528 -7492 25724 -7355
rect 24352 -7688 25724 -7492
rect 25808 -7492 26004 -7355
rect 26256 -7401 26732 -7355
rect 26984 -7492 27180 -7355
rect 25808 -7688 27180 -7492
rect 27456 -7898 27652 -3666
rect 28104 -3690 28248 -3666
rect 28294 -3666 31256 -3644
rect 28294 -3690 28424 -3666
rect 28104 -3738 28424 -3690
rect 28104 -3784 28248 -3738
rect 28294 -3784 28424 -3738
rect 28104 -3832 28424 -3784
rect 28104 -3878 28248 -3832
rect 28294 -3878 28424 -3832
rect 28104 -3926 28424 -3878
rect 28104 -3972 28248 -3926
rect 28294 -3972 28424 -3926
rect 28104 -4020 28424 -3972
rect 28104 -4066 28248 -4020
rect 28294 -4066 28424 -4020
rect 28104 -4114 28424 -4066
rect 28104 -4160 28248 -4114
rect 28294 -4160 28424 -4114
rect 28104 -4208 28424 -4160
rect 28104 -4254 28248 -4208
rect 28294 -4254 28424 -4208
rect 28104 -4302 28424 -4254
rect 28104 -4348 28248 -4302
rect 28294 -4348 28424 -4302
rect 28104 -4396 28424 -4348
rect 28104 -4442 28248 -4396
rect 28294 -4442 28424 -4396
rect 28104 -4490 28424 -4442
rect 28104 -4536 28248 -4490
rect 28294 -4536 28424 -4490
rect 28104 -4584 28424 -4536
rect 28104 -4630 28248 -4584
rect 28294 -4630 28424 -4584
rect 28104 -4678 28424 -4630
rect 28104 -4724 28248 -4678
rect 28294 -4724 28424 -4678
rect 28104 -4772 28424 -4724
rect 28104 -4818 28248 -4772
rect 28294 -4818 28424 -4772
rect 28104 -4866 28424 -4818
rect 28104 -4912 28248 -4866
rect 28294 -4912 28424 -4866
rect 28104 -4960 28424 -4912
rect 28104 -5006 28248 -4960
rect 28294 -5006 28424 -4960
rect 28104 -5054 28424 -5006
rect 28104 -5100 28248 -5054
rect 28294 -5100 28424 -5054
rect 28104 -5148 28424 -5100
rect 28104 -5194 28248 -5148
rect 28294 -5194 28424 -5148
rect 28104 -5242 28424 -5194
rect 28104 -5288 28248 -5242
rect 28294 -5288 28424 -5242
rect 28104 -5336 28424 -5288
rect 28104 -5382 28248 -5336
rect 28294 -5382 28424 -5336
rect 28104 -5430 28424 -5382
rect 28104 -5476 28248 -5430
rect 28294 -5476 28424 -5430
rect 28104 -5524 28424 -5476
rect 28802 -5485 28998 -3666
rect 29250 -4064 30294 -4052
rect 29250 -4116 29814 -4064
rect 29866 -4116 29918 -4064
rect 29970 -4116 30022 -4064
rect 30074 -4116 30126 -4064
rect 30178 -4116 30230 -4064
rect 30282 -4116 30294 -4064
rect 29250 -4168 30294 -4116
rect 29250 -4220 29814 -4168
rect 29866 -4220 29918 -4168
rect 29970 -4220 30022 -4168
rect 30074 -4220 30126 -4168
rect 30178 -4220 30230 -4168
rect 30282 -4220 30294 -4168
rect 29250 -4272 30294 -4220
rect 29250 -4324 29814 -4272
rect 29866 -4324 29918 -4272
rect 29970 -4324 30022 -4272
rect 30074 -4324 30126 -4272
rect 30178 -4324 30230 -4272
rect 30282 -4324 30294 -4272
rect 29250 -4336 30294 -4324
rect 29250 -5020 30294 -5008
rect 29250 -5072 29814 -5020
rect 29866 -5072 29918 -5020
rect 29970 -5072 30022 -5020
rect 30074 -5072 30126 -5020
rect 30178 -5072 30230 -5020
rect 30282 -5072 30294 -5020
rect 29250 -5124 30294 -5072
rect 29250 -5176 29814 -5124
rect 29866 -5176 29918 -5124
rect 29970 -5176 30022 -5124
rect 30074 -5176 30126 -5124
rect 30178 -5176 30230 -5124
rect 30282 -5176 30294 -5124
rect 29250 -5228 30294 -5176
rect 29250 -5280 29814 -5228
rect 29866 -5280 29918 -5228
rect 29970 -5280 30022 -5228
rect 30074 -5280 30126 -5228
rect 30178 -5280 30230 -5228
rect 30282 -5280 30294 -5228
rect 29250 -5332 30294 -5280
rect 29250 -5384 29814 -5332
rect 29866 -5384 29918 -5332
rect 29970 -5384 30022 -5332
rect 30074 -5384 30126 -5332
rect 30178 -5384 30230 -5332
rect 30282 -5384 30294 -5332
rect 29250 -5436 30294 -5384
rect 29250 -5488 29814 -5436
rect 29866 -5488 29918 -5436
rect 29970 -5488 30022 -5436
rect 30074 -5488 30126 -5436
rect 30178 -5488 30230 -5436
rect 30282 -5488 30294 -5436
rect 30538 -5485 30734 -3666
rect 31112 -3690 31256 -3666
rect 31302 -3690 31432 -3644
rect 31112 -3738 31432 -3690
rect 31112 -3784 31256 -3738
rect 31302 -3784 31432 -3738
rect 31112 -3832 31432 -3784
rect 31112 -3878 31256 -3832
rect 31302 -3878 31432 -3832
rect 31112 -3926 31432 -3878
rect 31112 -3972 31256 -3926
rect 31302 -3972 31432 -3926
rect 31112 -4020 31432 -3972
rect 31112 -4066 31256 -4020
rect 31302 -4066 31432 -4020
rect 31112 -4114 31432 -4066
rect 31112 -4160 31256 -4114
rect 31302 -4160 31432 -4114
rect 31112 -4208 31432 -4160
rect 31112 -4254 31256 -4208
rect 31302 -4254 31432 -4208
rect 31112 -4302 31432 -4254
rect 31112 -4348 31256 -4302
rect 31302 -4348 31432 -4302
rect 31112 -4396 31432 -4348
rect 31112 -4442 31256 -4396
rect 31302 -4442 31432 -4396
rect 31112 -4490 31432 -4442
rect 31112 -4536 31256 -4490
rect 31302 -4536 31432 -4490
rect 54527 -4444 54726 -4431
rect 54527 -4500 54544 -4444
rect 54600 -4500 54654 -4444
rect 54710 -4450 54726 -4444
rect 54710 -4496 56719 -4450
rect 54710 -4500 54726 -4496
rect 54527 -4517 54726 -4500
rect 31112 -4584 31432 -4536
rect 31112 -4630 31256 -4584
rect 31302 -4630 31432 -4584
rect 31112 -4678 31432 -4630
rect 31112 -4724 31256 -4678
rect 31302 -4724 31432 -4678
rect 31112 -4772 31432 -4724
rect 31112 -4818 31256 -4772
rect 31302 -4818 31432 -4772
rect 31112 -4866 31432 -4818
rect 31112 -4912 31256 -4866
rect 31302 -4912 31432 -4866
rect 31112 -4960 31432 -4912
rect 31112 -5006 31256 -4960
rect 31302 -5006 31432 -4960
rect 31112 -5054 31432 -5006
rect 31112 -5100 31256 -5054
rect 31302 -5100 31432 -5054
rect 31112 -5148 31432 -5100
rect 31112 -5194 31256 -5148
rect 31302 -5194 31432 -5148
rect 31112 -5242 31432 -5194
rect 31112 -5288 31256 -5242
rect 31302 -5288 31432 -5242
rect 31112 -5336 31432 -5288
rect 31112 -5382 31256 -5336
rect 31302 -5382 31432 -5336
rect 31112 -5430 31432 -5382
rect 31112 -5476 31256 -5430
rect 31302 -5476 31432 -5430
rect 29250 -5500 30294 -5488
rect 28104 -5570 28248 -5524
rect 28294 -5570 28424 -5524
rect 28104 -5618 28424 -5570
rect 28104 -5664 28248 -5618
rect 28294 -5664 28424 -5618
rect 28104 -5712 28424 -5664
rect 28104 -5758 28248 -5712
rect 28294 -5758 28424 -5712
rect 28104 -5806 28424 -5758
rect 28104 -5852 28248 -5806
rect 28294 -5852 28424 -5806
rect 28104 -5900 28424 -5852
rect 28104 -5946 28248 -5900
rect 28294 -5946 28424 -5900
rect 28104 -5994 28424 -5946
rect 28104 -6040 28248 -5994
rect 28294 -6040 28424 -5994
rect 28104 -6088 28424 -6040
rect 31112 -5524 31432 -5476
rect 31112 -5570 31256 -5524
rect 31302 -5570 31432 -5524
rect 54800 -5481 54999 -5468
rect 54800 -5537 54817 -5481
rect 54873 -5537 54927 -5481
rect 54983 -5493 54999 -5481
rect 54983 -5537 56707 -5493
rect 54800 -5539 56707 -5537
rect 54800 -5554 54999 -5539
rect 31112 -5618 31432 -5570
rect 31112 -5664 31256 -5618
rect 31302 -5664 31432 -5618
rect 31112 -5712 31432 -5664
rect 31112 -5758 31256 -5712
rect 31302 -5758 31432 -5712
rect 31112 -5806 31432 -5758
rect 31112 -5852 31256 -5806
rect 31302 -5852 31432 -5806
rect 31112 -5900 31432 -5852
rect 31112 -5946 31256 -5900
rect 31302 -5946 31432 -5900
rect 31112 -5994 31432 -5946
rect 31112 -6040 31256 -5994
rect 31302 -6040 31432 -5994
rect 29242 -6076 30286 -6064
rect 28104 -6134 28248 -6088
rect 28294 -6134 28424 -6088
rect 28104 -6182 28424 -6134
rect 28104 -6228 28248 -6182
rect 28294 -6228 28424 -6182
rect 28104 -6276 28424 -6228
rect 28104 -6322 28248 -6276
rect 28294 -6322 28424 -6276
rect 28104 -6370 28424 -6322
rect 28104 -6416 28248 -6370
rect 28294 -6416 28424 -6370
rect 28104 -6464 28424 -6416
rect 28104 -6510 28248 -6464
rect 28294 -6510 28424 -6464
rect 28104 -6558 28424 -6510
rect 28104 -6604 28248 -6558
rect 28294 -6604 28424 -6558
rect 28104 -6652 28424 -6604
rect 28104 -6698 28248 -6652
rect 28294 -6698 28424 -6652
rect 28104 -6746 28424 -6698
rect 28104 -6792 28248 -6746
rect 28294 -6792 28424 -6746
rect 28104 -6840 28424 -6792
rect 28104 -6886 28248 -6840
rect 28294 -6886 28424 -6840
rect 28104 -6934 28424 -6886
rect 28104 -6980 28248 -6934
rect 28294 -6980 28424 -6934
rect 28104 -7028 28424 -6980
rect 28104 -7074 28248 -7028
rect 28294 -7074 28424 -7028
rect 28104 -7122 28424 -7074
rect 28104 -7168 28248 -7122
rect 28294 -7168 28424 -7122
rect 28104 -7216 28424 -7168
rect 28104 -7262 28248 -7216
rect 28294 -7262 28424 -7216
rect 28104 -7310 28424 -7262
rect 28104 -7356 28248 -7310
rect 28294 -7356 28424 -7310
rect 28104 -7404 28424 -7356
rect 28104 -7450 28248 -7404
rect 28294 -7450 28424 -7404
rect 28104 -7498 28424 -7450
rect 28104 -7544 28248 -7498
rect 28294 -7544 28424 -7498
rect 28104 -7592 28424 -7544
rect 28104 -7638 28248 -7592
rect 28294 -7638 28424 -7592
rect 28104 -7686 28424 -7638
rect 28104 -7732 28248 -7686
rect 28294 -7732 28424 -7686
rect 28104 -7780 28424 -7732
rect 28104 -7826 28248 -7780
rect 28294 -7826 28424 -7780
rect 28104 -7874 28424 -7826
rect 28104 -7898 28248 -7874
rect 22560 -7920 28248 -7898
rect 28294 -7898 28424 -7874
rect 28802 -7898 28998 -6079
rect 29242 -6128 29254 -6076
rect 29306 -6128 29358 -6076
rect 29410 -6128 29462 -6076
rect 29514 -6128 29566 -6076
rect 29618 -6128 29670 -6076
rect 29722 -6128 30286 -6076
rect 29242 -6180 30286 -6128
rect 29242 -6232 29254 -6180
rect 29306 -6232 29358 -6180
rect 29410 -6232 29462 -6180
rect 29514 -6232 29566 -6180
rect 29618 -6232 29670 -6180
rect 29722 -6232 30286 -6180
rect 29242 -6284 30286 -6232
rect 29242 -6336 29254 -6284
rect 29306 -6336 29358 -6284
rect 29410 -6336 29462 -6284
rect 29514 -6336 29566 -6284
rect 29618 -6336 29670 -6284
rect 29722 -6336 30286 -6284
rect 29242 -6348 30286 -6336
rect 29250 -7032 30294 -7020
rect 29250 -7084 29814 -7032
rect 29866 -7084 29918 -7032
rect 29970 -7084 30022 -7032
rect 30074 -7084 30126 -7032
rect 30178 -7084 30230 -7032
rect 30282 -7084 30294 -7032
rect 29250 -7136 30294 -7084
rect 29250 -7188 29814 -7136
rect 29866 -7188 29918 -7136
rect 29970 -7188 30022 -7136
rect 30074 -7188 30126 -7136
rect 30178 -7188 30230 -7136
rect 30282 -7188 30294 -7136
rect 29250 -7240 30294 -7188
rect 29250 -7292 29814 -7240
rect 29866 -7292 29918 -7240
rect 29970 -7292 30022 -7240
rect 30074 -7292 30126 -7240
rect 30178 -7292 30230 -7240
rect 30282 -7292 30294 -7240
rect 29250 -7344 30294 -7292
rect 29250 -7396 29814 -7344
rect 29866 -7396 29918 -7344
rect 29970 -7396 30022 -7344
rect 30074 -7396 30126 -7344
rect 30178 -7396 30230 -7344
rect 30282 -7396 30294 -7344
rect 29250 -7448 30294 -7396
rect 29250 -7500 29814 -7448
rect 29866 -7500 29918 -7448
rect 29970 -7500 30022 -7448
rect 30074 -7500 30126 -7448
rect 30178 -7500 30230 -7448
rect 30282 -7500 30294 -7448
rect 29250 -7512 30294 -7500
rect 30538 -7898 30734 -6079
rect 31112 -6088 31432 -6040
rect 31112 -6134 31256 -6088
rect 31302 -6134 31432 -6088
rect 31112 -6182 31432 -6134
rect 31112 -6228 31256 -6182
rect 31302 -6228 31432 -6182
rect 31112 -6276 31432 -6228
rect 31112 -6322 31256 -6276
rect 31302 -6322 31432 -6276
rect 31112 -6370 31432 -6322
rect 31112 -6416 31256 -6370
rect 31302 -6416 31432 -6370
rect 31112 -6464 31432 -6416
rect 55049 -6355 55248 -6342
rect 55049 -6411 55066 -6355
rect 55122 -6411 55176 -6355
rect 55232 -6364 55248 -6355
rect 55232 -6410 56911 -6364
rect 55232 -6411 55248 -6410
rect 55049 -6428 55248 -6411
rect 31112 -6510 31256 -6464
rect 31302 -6510 31432 -6464
rect 31112 -6558 31432 -6510
rect 31112 -6604 31256 -6558
rect 31302 -6604 31432 -6558
rect 31112 -6652 31432 -6604
rect 31112 -6698 31256 -6652
rect 31302 -6698 31432 -6652
rect 31112 -6746 31432 -6698
rect 31112 -6792 31256 -6746
rect 31302 -6792 31432 -6746
rect 31112 -6840 31432 -6792
rect 31112 -6886 31256 -6840
rect 31302 -6886 31432 -6840
rect 31112 -6934 31432 -6886
rect 31112 -6980 31256 -6934
rect 31302 -6980 31432 -6934
rect 31112 -7028 31432 -6980
rect 31112 -7074 31256 -7028
rect 31302 -7074 31432 -7028
rect 31112 -7122 31432 -7074
rect 31112 -7168 31256 -7122
rect 31302 -7168 31432 -7122
rect 31112 -7216 31432 -7168
rect 31112 -7262 31256 -7216
rect 31302 -7262 31432 -7216
rect 31112 -7310 31432 -7262
rect 31112 -7356 31256 -7310
rect 31302 -7356 31432 -7310
rect 31112 -7404 31432 -7356
rect 31112 -7450 31256 -7404
rect 31302 -7450 31432 -7404
rect 31112 -7498 31432 -7450
rect 55298 -7404 55497 -7391
rect 55298 -7460 55315 -7404
rect 55371 -7460 55425 -7404
rect 55481 -7407 55497 -7404
rect 55481 -7453 56718 -7407
rect 55481 -7460 55497 -7453
rect 55298 -7477 55497 -7460
rect 31112 -7544 31256 -7498
rect 31302 -7544 31432 -7498
rect 31112 -7592 31432 -7544
rect 31112 -7638 31256 -7592
rect 31302 -7638 31432 -7592
rect 31112 -7686 31432 -7638
rect 31112 -7732 31256 -7686
rect 31302 -7732 31432 -7686
rect 31112 -7780 31432 -7732
rect 31112 -7826 31256 -7780
rect 31302 -7826 31432 -7780
rect 31112 -7874 31432 -7826
rect 31112 -7898 31256 -7874
rect 28294 -7920 31256 -7898
rect 31302 -7920 31432 -7874
rect 6168 -12783 6682 -7936
rect 17590 -7968 31432 -7920
rect 17590 -8014 17720 -7968
rect 17766 -8014 22514 -7968
rect 22560 -8014 28248 -7968
rect 28294 -8014 31256 -7968
rect 31302 -8014 31432 -7968
rect 11532 -8026 11712 -8018
rect 11532 -8030 12000 -8026
rect 11532 -8082 11544 -8030
rect 11596 -8082 11648 -8030
rect 11700 -8082 12000 -8030
rect 11532 -8134 12000 -8082
rect 11532 -8186 11544 -8134
rect 11596 -8186 11648 -8134
rect 11700 -8186 12000 -8134
rect 17590 -8062 31432 -8014
rect 44536 -7956 50146 -7944
rect 44536 -8008 44548 -7956
rect 44600 -8008 44652 -7956
rect 44704 -8008 44756 -7956
rect 44808 -8008 44860 -7956
rect 44912 -8008 44964 -7956
rect 45016 -8008 48988 -7956
rect 49040 -8008 49092 -7956
rect 49144 -8008 49196 -7956
rect 49248 -8008 49300 -7956
rect 49352 -8008 49404 -7956
rect 49456 -8008 50146 -7956
rect 17590 -8108 17720 -8062
rect 17766 -8108 17814 -8062
rect 17860 -8108 17908 -8062
rect 17954 -8108 18002 -8062
rect 18048 -8108 18096 -8062
rect 18142 -8108 18190 -8062
rect 18236 -8108 18284 -8062
rect 18330 -8108 18378 -8062
rect 18424 -8108 18472 -8062
rect 18518 -8108 18566 -8062
rect 18612 -8108 18660 -8062
rect 18706 -8108 18754 -8062
rect 18800 -8108 18848 -8062
rect 18894 -8108 18942 -8062
rect 18988 -8108 19036 -8062
rect 19082 -8108 19130 -8062
rect 19176 -8108 19224 -8062
rect 19270 -8108 19318 -8062
rect 19364 -8108 19412 -8062
rect 19458 -8108 19506 -8062
rect 19552 -8108 19600 -8062
rect 19646 -8108 19694 -8062
rect 19740 -8108 19788 -8062
rect 19834 -8108 19882 -8062
rect 19928 -8108 19976 -8062
rect 20022 -8108 20070 -8062
rect 20116 -8108 20164 -8062
rect 20210 -8108 20258 -8062
rect 20304 -8108 20352 -8062
rect 20398 -8108 20446 -8062
rect 20492 -8108 20540 -8062
rect 20586 -8108 20634 -8062
rect 20680 -8108 20728 -8062
rect 20774 -8108 20822 -8062
rect 20868 -8108 20916 -8062
rect 20962 -8108 21010 -8062
rect 21056 -8108 21104 -8062
rect 21150 -8108 21198 -8062
rect 21244 -8108 21292 -8062
rect 21338 -8108 21386 -8062
rect 21432 -8108 21480 -8062
rect 21526 -8108 21574 -8062
rect 21620 -8108 21668 -8062
rect 21714 -8108 21762 -8062
rect 21808 -8108 21856 -8062
rect 21902 -8108 21950 -8062
rect 21996 -8108 22044 -8062
rect 22090 -8108 22138 -8062
rect 22184 -8108 22232 -8062
rect 22278 -8108 22326 -8062
rect 22372 -8108 22420 -8062
rect 22466 -8108 22514 -8062
rect 22560 -8108 22608 -8062
rect 22654 -8108 22702 -8062
rect 22748 -8108 22796 -8062
rect 22842 -8108 22890 -8062
rect 22936 -8108 22984 -8062
rect 23030 -8108 23078 -8062
rect 23124 -8108 23172 -8062
rect 23218 -8108 23266 -8062
rect 23312 -8108 23360 -8062
rect 23406 -8108 23454 -8062
rect 23500 -8108 23548 -8062
rect 23594 -8108 23642 -8062
rect 23688 -8108 23736 -8062
rect 23782 -8108 23830 -8062
rect 23876 -8108 23924 -8062
rect 23970 -8108 24018 -8062
rect 24064 -8108 24112 -8062
rect 24158 -8108 24206 -8062
rect 24252 -8108 24300 -8062
rect 24346 -8108 24394 -8062
rect 24440 -8108 24488 -8062
rect 24534 -8108 24582 -8062
rect 24628 -8108 24676 -8062
rect 24722 -8108 24770 -8062
rect 24816 -8108 24864 -8062
rect 24910 -8108 24958 -8062
rect 25004 -8108 25052 -8062
rect 25098 -8108 25146 -8062
rect 25192 -8108 25240 -8062
rect 25286 -8108 25334 -8062
rect 25380 -8108 25428 -8062
rect 25474 -8108 25522 -8062
rect 25568 -8108 25616 -8062
rect 25662 -8108 25710 -8062
rect 25756 -8108 25804 -8062
rect 25850 -8108 25898 -8062
rect 25944 -8108 25992 -8062
rect 26038 -8108 26086 -8062
rect 26132 -8108 26180 -8062
rect 26226 -8108 26274 -8062
rect 26320 -8108 26368 -8062
rect 26414 -8108 26462 -8062
rect 26508 -8108 26556 -8062
rect 26602 -8108 26650 -8062
rect 26696 -8108 26744 -8062
rect 26790 -8108 26838 -8062
rect 26884 -8108 26932 -8062
rect 26978 -8108 27026 -8062
rect 27072 -8108 27120 -8062
rect 27166 -8108 27214 -8062
rect 27260 -8108 27308 -8062
rect 27354 -8108 27402 -8062
rect 27448 -8108 27496 -8062
rect 27542 -8108 27590 -8062
rect 27636 -8108 27684 -8062
rect 27730 -8108 27778 -8062
rect 27824 -8108 27872 -8062
rect 27918 -8108 27966 -8062
rect 28012 -8108 28060 -8062
rect 28106 -8108 28154 -8062
rect 28200 -8108 28248 -8062
rect 28294 -8108 28342 -8062
rect 28388 -8108 28436 -8062
rect 28482 -8108 28530 -8062
rect 28576 -8108 28624 -8062
rect 28670 -8108 28718 -8062
rect 28764 -8108 28812 -8062
rect 28858 -8108 28906 -8062
rect 28952 -8108 29000 -8062
rect 29046 -8108 29094 -8062
rect 29140 -8108 29188 -8062
rect 29234 -8108 29282 -8062
rect 29328 -8108 29376 -8062
rect 29422 -8108 29470 -8062
rect 29516 -8108 29564 -8062
rect 29610 -8108 29658 -8062
rect 29704 -8108 29752 -8062
rect 29798 -8108 29846 -8062
rect 29892 -8108 29940 -8062
rect 29986 -8108 30034 -8062
rect 30080 -8108 30128 -8062
rect 30174 -8108 30222 -8062
rect 30268 -8108 30316 -8062
rect 30362 -8108 30410 -8062
rect 30456 -8108 30504 -8062
rect 30550 -8108 30598 -8062
rect 30644 -8108 30692 -8062
rect 30738 -8108 30786 -8062
rect 30832 -8108 30880 -8062
rect 30926 -8108 30974 -8062
rect 31020 -8108 31068 -8062
rect 31114 -8108 31162 -8062
rect 31208 -8108 31256 -8062
rect 31302 -8108 31432 -8062
rect 11532 -8198 11712 -8186
rect 17590 -8218 31432 -8108
rect 34706 -8056 40316 -8044
rect 34706 -8108 34718 -8056
rect 34770 -8108 34822 -8056
rect 34874 -8108 34926 -8056
rect 34978 -8108 35030 -8056
rect 35082 -8108 35134 -8056
rect 35186 -8108 39158 -8056
rect 39210 -8108 39262 -8056
rect 39314 -8108 39366 -8056
rect 39418 -8108 39470 -8056
rect 39522 -8108 39574 -8056
rect 39626 -8108 40316 -8056
rect 34706 -8160 40316 -8108
rect 34706 -8212 34718 -8160
rect 34770 -8212 34822 -8160
rect 34874 -8212 34926 -8160
rect 34978 -8212 35030 -8160
rect 35082 -8212 35134 -8160
rect 35186 -8212 39158 -8160
rect 39210 -8212 39262 -8160
rect 39314 -8212 39366 -8160
rect 39418 -8212 39470 -8160
rect 39522 -8212 39574 -8160
rect 39626 -8212 40316 -8160
rect 15070 -8885 15854 -8873
rect 15070 -8937 15082 -8885
rect 15134 -8937 15186 -8885
rect 15238 -8937 15290 -8885
rect 15342 -8937 15854 -8885
rect 15070 -8989 15854 -8937
rect 15070 -9041 15082 -8989
rect 15134 -9041 15186 -8989
rect 15238 -9041 15290 -8989
rect 15342 -9041 15854 -8989
rect 15070 -9093 15854 -9041
rect 15070 -9145 15082 -9093
rect 15134 -9145 15186 -9093
rect 15238 -9145 15290 -9093
rect 15342 -9145 15854 -9093
rect 15070 -9157 15854 -9145
rect 17671 -11721 18384 -8218
rect 21145 -8385 21989 -8373
rect 21145 -8437 21157 -8385
rect 21209 -8437 21261 -8385
rect 21313 -8437 21365 -8385
rect 21417 -8437 21989 -8385
rect 21145 -8489 21989 -8437
rect 21145 -8541 21157 -8489
rect 21209 -8541 21261 -8489
rect 21313 -8541 21365 -8489
rect 21417 -8541 21989 -8489
rect 21145 -8593 21989 -8541
rect 21145 -8645 21157 -8593
rect 21209 -8645 21261 -8593
rect 21313 -8645 21365 -8593
rect 21417 -8645 21989 -8593
rect 21145 -8657 21989 -8645
rect 26397 -11714 27285 -8218
rect 34706 -8264 40316 -8212
rect 34706 -8316 34718 -8264
rect 34770 -8316 34822 -8264
rect 34874 -8316 34926 -8264
rect 34978 -8316 35030 -8264
rect 35082 -8316 35134 -8264
rect 35186 -8316 39158 -8264
rect 39210 -8316 39262 -8264
rect 39314 -8316 39366 -8264
rect 39418 -8316 39470 -8264
rect 39522 -8316 39574 -8264
rect 39626 -8316 40316 -8264
rect 34706 -8368 40316 -8316
rect 34706 -8420 34718 -8368
rect 34770 -8420 34822 -8368
rect 34874 -8420 34926 -8368
rect 34978 -8420 35030 -8368
rect 35082 -8420 35134 -8368
rect 35186 -8420 39158 -8368
rect 39210 -8420 39262 -8368
rect 39314 -8420 39366 -8368
rect 39418 -8420 39470 -8368
rect 39522 -8420 39574 -8368
rect 39626 -8420 40316 -8368
rect 34706 -8472 40316 -8420
rect 44536 -8060 50146 -8008
rect 44536 -8112 44548 -8060
rect 44600 -8112 44652 -8060
rect 44704 -8112 44756 -8060
rect 44808 -8112 44860 -8060
rect 44912 -8112 44964 -8060
rect 45016 -8112 48988 -8060
rect 49040 -8112 49092 -8060
rect 49144 -8112 49196 -8060
rect 49248 -8112 49300 -8060
rect 49352 -8112 49404 -8060
rect 49456 -8112 50146 -8060
rect 44536 -8164 50146 -8112
rect 44536 -8216 44548 -8164
rect 44600 -8216 44652 -8164
rect 44704 -8216 44756 -8164
rect 44808 -8216 44860 -8164
rect 44912 -8216 44964 -8164
rect 45016 -8216 48988 -8164
rect 49040 -8216 49092 -8164
rect 49144 -8216 49196 -8164
rect 49248 -8216 49300 -8164
rect 49352 -8216 49404 -8164
rect 49456 -8216 50146 -8164
rect 44536 -8268 50146 -8216
rect 44536 -8320 44548 -8268
rect 44600 -8320 44652 -8268
rect 44704 -8320 44756 -8268
rect 44808 -8320 44860 -8268
rect 44912 -8320 44964 -8268
rect 45016 -8320 48988 -8268
rect 49040 -8320 49092 -8268
rect 49144 -8320 49196 -8268
rect 49248 -8320 49300 -8268
rect 49352 -8320 49404 -8268
rect 49456 -8320 50146 -8268
rect 44536 -8372 50146 -8320
rect 44536 -8424 44548 -8372
rect 44600 -8424 44652 -8372
rect 44704 -8424 44756 -8372
rect 44808 -8424 44860 -8372
rect 44912 -8424 44964 -8372
rect 45016 -8424 48988 -8372
rect 49040 -8424 49092 -8372
rect 49144 -8424 49196 -8372
rect 49248 -8424 49300 -8372
rect 49352 -8424 49404 -8372
rect 49456 -8424 50146 -8372
rect 44536 -8436 50146 -8424
rect 34706 -8524 34718 -8472
rect 34770 -8524 34822 -8472
rect 34874 -8524 34926 -8472
rect 34978 -8524 35030 -8472
rect 35082 -8524 35134 -8472
rect 35186 -8524 39158 -8472
rect 39210 -8524 39262 -8472
rect 39314 -8524 39366 -8472
rect 39418 -8524 39470 -8472
rect 39522 -8524 39574 -8472
rect 39626 -8524 40316 -8472
rect 34706 -8536 40316 -8524
rect 55644 -8742 55843 -8729
rect 55644 -8798 55661 -8742
rect 55717 -8798 55771 -8742
rect 55827 -8743 55843 -8742
rect 55827 -8790 56693 -8743
rect 55827 -8798 55843 -8790
rect 55644 -8815 55843 -8798
rect 56523 -10479 57347 -10312
rect 7380 -11849 18417 -11721
rect 24371 -11842 35408 -11714
rect 8450 -12287 8649 -12274
rect 8450 -12314 8467 -12287
rect 8342 -12343 8467 -12314
rect 8523 -12343 8577 -12287
rect 8633 -12343 8649 -12287
rect 10443 -12287 10642 -12274
rect 10443 -12314 10460 -12287
rect 6865 -12363 7064 -12350
rect 8342 -12360 8649 -12343
rect 10356 -12343 10460 -12314
rect 10516 -12343 10570 -12287
rect 10626 -12343 10642 -12287
rect 12472 -12287 12671 -12274
rect 12472 -12314 12489 -12287
rect 8866 -12360 9065 -12347
rect 10356 -12360 10642 -12343
rect 12365 -12343 12489 -12314
rect 12545 -12343 12599 -12287
rect 12655 -12343 12671 -12287
rect 14475 -12287 14674 -12274
rect 14475 -12314 14492 -12287
rect 6865 -12419 6882 -12363
rect 6938 -12419 6992 -12363
rect 7048 -12366 7064 -12363
rect 7048 -12419 7396 -12366
rect 6865 -12420 7396 -12419
rect 8866 -12416 8883 -12360
rect 8939 -12416 8993 -12360
rect 9049 -12366 9065 -12360
rect 10891 -12363 11090 -12350
rect 12365 -12360 12671 -12343
rect 14365 -12343 14492 -12314
rect 14548 -12343 14602 -12287
rect 14658 -12343 14674 -12287
rect 16490 -12288 16689 -12275
rect 16490 -12314 16507 -12288
rect 9049 -12416 9383 -12366
rect 8866 -12420 9383 -12416
rect 10891 -12419 10908 -12363
rect 10964 -12419 11018 -12363
rect 11074 -12366 11090 -12363
rect 12900 -12362 13099 -12349
rect 14365 -12360 14674 -12343
rect 16365 -12344 16507 -12314
rect 16563 -12344 16617 -12288
rect 16673 -12344 16689 -12288
rect 18511 -12287 18710 -12274
rect 18511 -12314 18528 -12287
rect 11074 -12419 11409 -12366
rect 10891 -12420 11409 -12419
rect 12900 -12418 12917 -12362
rect 12973 -12418 13027 -12362
rect 13083 -12366 13099 -12362
rect 14870 -12362 15069 -12349
rect 16365 -12360 16689 -12344
rect 18365 -12343 18528 -12314
rect 18584 -12343 18638 -12287
rect 18694 -12343 18710 -12287
rect 25450 -12287 25649 -12274
rect 25450 -12314 25467 -12287
rect 16490 -12361 16689 -12360
rect 16905 -12358 17104 -12345
rect 13083 -12418 13391 -12366
rect 12900 -12420 13391 -12418
rect 14870 -12418 14887 -12362
rect 14943 -12418 14997 -12362
rect 15053 -12366 15069 -12362
rect 15053 -12418 15406 -12366
rect 14870 -12420 15406 -12418
rect 16905 -12414 16922 -12358
rect 16978 -12414 17032 -12358
rect 17088 -12366 17104 -12358
rect 18365 -12360 18710 -12343
rect 25342 -12343 25467 -12314
rect 25523 -12343 25577 -12287
rect 25633 -12343 25649 -12287
rect 27443 -12287 27642 -12274
rect 27443 -12314 27460 -12287
rect 23865 -12363 24064 -12350
rect 25342 -12360 25649 -12343
rect 27356 -12343 27460 -12314
rect 27516 -12343 27570 -12287
rect 27626 -12343 27642 -12287
rect 29472 -12287 29671 -12274
rect 29472 -12314 29489 -12287
rect 25866 -12360 26065 -12347
rect 27356 -12360 27642 -12343
rect 29365 -12343 29489 -12314
rect 29545 -12343 29599 -12287
rect 29655 -12343 29671 -12287
rect 31475 -12287 31674 -12274
rect 31475 -12314 31492 -12287
rect 17088 -12414 17409 -12366
rect 16905 -12420 17409 -12414
rect 23865 -12419 23882 -12363
rect 23938 -12419 23992 -12363
rect 24048 -12366 24064 -12363
rect 24048 -12419 24396 -12366
rect 23865 -12420 24396 -12419
rect 25866 -12416 25883 -12360
rect 25939 -12416 25993 -12360
rect 26049 -12366 26065 -12360
rect 27891 -12363 28090 -12350
rect 29365 -12360 29671 -12343
rect 31365 -12343 31492 -12314
rect 31548 -12343 31602 -12287
rect 31658 -12343 31674 -12287
rect 33490 -12288 33689 -12275
rect 33490 -12314 33507 -12288
rect 26049 -12416 26383 -12366
rect 25866 -12420 26383 -12416
rect 27891 -12419 27908 -12363
rect 27964 -12419 28018 -12363
rect 28074 -12366 28090 -12363
rect 29900 -12362 30099 -12349
rect 31365 -12360 31674 -12343
rect 33365 -12344 33507 -12314
rect 33563 -12344 33617 -12288
rect 33673 -12344 33689 -12288
rect 35511 -12287 35710 -12274
rect 35511 -12314 35528 -12287
rect 28074 -12419 28409 -12366
rect 27891 -12420 28409 -12419
rect 29900 -12418 29917 -12362
rect 29973 -12418 30027 -12362
rect 30083 -12366 30099 -12362
rect 31870 -12362 32069 -12349
rect 33365 -12360 33689 -12344
rect 35365 -12343 35528 -12314
rect 35584 -12343 35638 -12287
rect 35694 -12343 35710 -12287
rect 33490 -12361 33689 -12360
rect 33905 -12358 34104 -12345
rect 30083 -12418 30391 -12366
rect 29900 -12420 30391 -12418
rect 31870 -12418 31887 -12362
rect 31943 -12418 31997 -12362
rect 32053 -12366 32069 -12362
rect 32053 -12418 32406 -12366
rect 31870 -12420 32406 -12418
rect 33905 -12414 33922 -12358
rect 33978 -12414 34032 -12358
rect 34088 -12366 34104 -12358
rect 35365 -12360 35710 -12343
rect 35883 -12314 36082 -12301
rect 34088 -12414 34409 -12366
rect 35883 -12370 35900 -12314
rect 35956 -12370 36010 -12314
rect 36066 -12370 36082 -12314
rect 35883 -12387 36082 -12370
rect 33905 -12420 34409 -12414
rect 6865 -12436 7064 -12420
rect 8866 -12433 9065 -12420
rect 10891 -12436 11090 -12420
rect 12900 -12435 13099 -12420
rect 14870 -12435 15069 -12420
rect 16905 -12431 17104 -12420
rect 23865 -12436 24064 -12420
rect 25866 -12433 26065 -12420
rect 27891 -12436 28090 -12420
rect 29900 -12435 30099 -12420
rect 31870 -12435 32069 -12420
rect 33905 -12431 34104 -12420
rect 56530 -12783 56785 -10479
rect 6168 -12838 56787 -12783
rect 6166 -13182 56787 -12838
rect 3250 -14632 7285 -14035
rect 17267 -14730 24286 -14038
rect 34747 -16138 39578 -16035
rect 17744 -16201 19290 -16175
rect 17744 -16257 18977 -16201
rect 19033 -16257 19087 -16201
rect 19143 -16257 19197 -16201
rect 19253 -16257 19290 -16201
rect 17744 -16311 19290 -16257
rect 17744 -16367 18977 -16311
rect 19033 -16367 19087 -16311
rect 19143 -16367 19197 -16311
rect 19253 -16367 19290 -16311
rect 17744 -16421 19290 -16367
rect 17744 -16477 18977 -16421
rect 19033 -16477 19087 -16421
rect 19143 -16477 19197 -16421
rect 19253 -16477 19290 -16421
rect 34747 -16194 39211 -16138
rect 39267 -16194 39321 -16138
rect 39377 -16194 39431 -16138
rect 39487 -16194 39578 -16138
rect 34747 -16248 39578 -16194
rect 34747 -16304 39211 -16248
rect 39267 -16304 39321 -16248
rect 39377 -16304 39431 -16248
rect 39487 -16304 39578 -16248
rect 34747 -16358 39578 -16304
rect 34747 -16414 39211 -16358
rect 39267 -16414 39321 -16358
rect 39377 -16414 39431 -16358
rect 39487 -16414 39578 -16358
rect 34747 -16439 39578 -16414
rect 17744 -16486 19290 -16477
rect 6909 -17853 6972 -16834
rect 5115 -18387 6972 -17853
rect 23909 -17964 23972 -16982
rect 6909 -18418 6972 -18387
rect 22058 -18615 23972 -17964
rect 23909 -18646 23972 -18615
<< via1 >>
rect 30744 6496 30796 6548
rect 30848 6496 30900 6548
rect 30952 6496 31004 6548
rect 30744 6392 30796 6444
rect 30848 6392 30900 6444
rect 30952 6392 31004 6444
rect 30744 6288 30796 6340
rect 30848 6288 30900 6340
rect 30952 6288 31004 6340
rect 31658 5910 31710 5962
rect 31762 5910 31814 5962
rect 31866 5910 31918 5962
rect 31658 5806 31710 5858
rect 31762 5806 31814 5858
rect 31866 5806 31918 5858
rect 31658 5702 31710 5754
rect 31762 5702 31814 5754
rect 31866 5702 31918 5754
rect -1781 5134 -1725 5190
rect -1671 5134 -1615 5190
rect -1561 5134 -1505 5190
rect 2687 5117 2739 5169
rect 2791 5117 2843 5169
rect -1781 5024 -1725 5080
rect -1671 5024 -1615 5080
rect -1561 5024 -1505 5080
rect 2687 5013 2739 5065
rect 2791 5013 2843 5065
rect 3476 5062 3528 5065
rect 3476 5016 3479 5062
rect 3479 5016 3525 5062
rect 3525 5016 3528 5062
rect 3476 5013 3528 5016
rect 5257 5063 5309 5115
rect 5361 5063 5413 5115
rect 5257 4959 5309 5011
rect 5361 4959 5413 5011
rect 2046 4768 2098 4820
rect 2150 4768 2202 4820
rect 2046 4664 2098 4716
rect 2150 4664 2202 4716
rect 3556 4768 3608 4820
rect 3556 4664 3608 4716
rect 3716 4768 3768 4820
rect 3716 4664 3768 4716
rect 4357 4768 4409 4820
rect 4357 4664 4409 4716
rect 6261 5063 6313 5115
rect 6261 4959 6313 5011
rect 6901 5063 6953 5115
rect 6901 4959 6953 5011
rect 7541 5063 7593 5115
rect 7541 4959 7593 5011
rect 5529 4768 5581 4820
rect 5633 4768 5685 4820
rect 5529 4664 5581 4716
rect 5633 4664 5685 4716
rect 3396 4272 3448 4324
rect 3396 4168 3448 4220
rect 4036 4272 4088 4324
rect 4036 4168 4088 4220
rect 4676 4272 4728 4324
rect 4676 4168 4728 4220
rect -1106 3976 -1050 4032
rect -996 3976 -940 4032
rect -886 3976 -830 4032
rect 2407 3989 2459 4041
rect 2511 3989 2563 4041
rect -1106 3866 -1050 3922
rect -996 3866 -940 3922
rect -886 3866 -830 3922
rect 2407 3885 2459 3937
rect 2511 3885 2563 3937
rect 3476 3989 3528 4041
rect 3476 3934 3528 3937
rect 3476 3888 3479 3934
rect 3479 3888 3525 3934
rect 3525 3888 3528 3934
rect 3476 3885 3528 3888
rect 3556 3638 3608 3690
rect 3556 3534 3608 3586
rect 3716 3638 3768 3690
rect 3716 3534 3768 3586
rect 4357 3638 4409 3690
rect 4357 3534 4409 3586
rect 3396 3246 3448 3298
rect 3396 3142 3448 3194
rect 4036 3246 4088 3298
rect 4036 3142 4088 3194
rect 4676 3246 4728 3298
rect 4676 3142 4728 3194
rect 3476 2859 3528 2911
rect 3476 2806 3528 2807
rect 3476 2760 3479 2806
rect 3479 2760 3525 2806
rect 3525 2760 3528 2806
rect 3476 2755 3528 2760
rect 3716 2508 3768 2560
rect 3716 2404 3768 2456
rect 4357 2508 4409 2560
rect 4357 2404 4409 2456
rect 3396 2012 3448 2064
rect 3396 1908 3448 1960
rect 4036 2012 4088 2064
rect 4036 1908 4088 1960
rect 4676 2012 4728 2064
rect 4676 1908 4728 1960
rect 2046 1114 2098 1166
rect 2150 1114 2202 1166
rect 2046 1010 2098 1062
rect 2150 1010 2202 1062
rect 3556 1114 3608 1166
rect 3556 1010 3608 1062
rect 3476 601 3528 653
rect 3476 546 3528 549
rect 3476 500 3479 546
rect 3479 500 3525 546
rect 3525 500 3528 546
rect 3476 497 3528 500
rect 2150 248 2202 300
rect 2150 144 2202 196
rect 3556 248 3608 300
rect 3556 144 3608 196
rect 3716 248 3768 300
rect 3716 144 3768 196
rect 4357 248 4409 300
rect 4357 144 4409 196
rect 3396 -248 3448 -196
rect 3396 -352 3448 -300
rect 4036 -248 4088 -196
rect 4036 -352 4088 -300
rect 4676 -248 4728 -196
rect 4676 -352 4728 -300
rect 3476 -529 3528 -477
rect 3476 -584 3528 -581
rect 3476 -630 3479 -584
rect 3479 -630 3525 -584
rect 3525 -630 3528 -584
rect 3476 -633 3528 -630
rect 2150 -1082 2202 -1030
rect 2150 -1186 2202 -1134
rect 3716 -882 3768 -830
rect 3716 -986 3768 -934
rect 4357 -882 4409 -830
rect 4357 -986 4409 -934
rect 3556 -1082 3608 -1030
rect 3556 -1186 3608 -1134
rect -248 -1626 -196 -1574
rect -144 -1626 -92 -1574
rect -248 -1730 -196 -1678
rect -144 -1730 -92 -1678
rect 753 -1577 805 -1574
rect 753 -1623 756 -1577
rect 756 -1623 802 -1577
rect 802 -1623 805 -1577
rect 753 -1626 805 -1623
rect 857 -1577 909 -1574
rect 857 -1623 860 -1577
rect 860 -1623 906 -1577
rect 906 -1623 909 -1577
rect 857 -1626 909 -1623
rect 3396 -1378 3448 -1326
rect 3396 -1482 3448 -1430
rect 4036 -1378 4088 -1326
rect 4036 -1482 4088 -1430
rect 4676 -1378 4728 -1326
rect 4676 -1482 4728 -1430
rect 3636 -1668 3688 -1665
rect 3636 -1714 3639 -1668
rect 3639 -1714 3685 -1668
rect 3685 -1714 3688 -1668
rect 3636 -1717 3688 -1714
rect 6581 4768 6633 4820
rect 6581 4664 6633 4716
rect 7221 4768 7273 4820
rect 7221 4664 7273 4716
rect 6581 4168 6633 4220
rect 6581 4064 6633 4116
rect 7221 4168 7273 4220
rect 7221 4064 7273 4116
rect 18591 4245 18643 4248
rect 19711 4245 19763 4248
rect 18591 4199 18594 4245
rect 18594 4199 18640 4245
rect 18640 4199 18643 4245
rect 19711 4199 19714 4245
rect 19714 4199 19760 4245
rect 19760 4199 19763 4245
rect 18591 4196 18643 4199
rect 19711 4196 19763 4199
rect 6261 3789 6313 3841
rect 6261 3685 6313 3737
rect 6901 3789 6953 3841
rect 6901 3685 6953 3737
rect 7541 3789 7593 3841
rect 7541 3685 7593 3737
rect 18831 3955 18883 4007
rect 18831 3851 18883 3903
rect 19471 3955 19523 4007
rect 19471 3851 19523 3903
rect 6581 3246 6633 3298
rect 6581 3142 6633 3194
rect 7221 3246 7273 3298
rect 7221 3142 7273 3194
rect 6261 2927 6313 2979
rect 6261 2823 6313 2875
rect 6901 2927 6953 2979
rect 6901 2823 6953 2875
rect 7541 2927 7593 2979
rect 7541 2823 7593 2875
rect 6261 2404 6313 2456
rect 6261 2300 6313 2352
rect 6901 2404 6953 2456
rect 6901 2300 6953 2352
rect 7541 2404 7593 2456
rect 7541 2300 7593 2352
rect 6581 2116 6633 2168
rect 6581 2012 6633 2064
rect 7221 2116 7273 2168
rect 7221 2012 7273 2064
rect 18511 3561 18563 3613
rect 18511 3457 18563 3509
rect 18671 3561 18723 3613
rect 18671 3457 18723 3509
rect 18991 3561 19043 3613
rect 18991 3457 19043 3509
rect 19151 3561 19203 3613
rect 19151 3457 19203 3509
rect 19311 3561 19363 3613
rect 19311 3457 19363 3509
rect 19631 3561 19683 3613
rect 19631 3457 19683 3509
rect 19791 3561 19843 3613
rect 19791 3457 19843 3509
rect 10897 2164 10949 2216
rect 11001 2164 11053 2216
rect 10897 2060 10949 2112
rect 11001 2060 11053 2112
rect 8496 1585 8548 1637
rect 8496 1481 8548 1533
rect 9392 1585 9444 1637
rect 9392 1481 9444 1533
rect 12326 2164 12378 2216
rect 12326 2060 12378 2112
rect 13222 2164 13274 2216
rect 13222 2060 13274 2112
rect 13510 2164 13562 2216
rect 13510 2060 13562 2112
rect 10288 1585 10340 1637
rect 10288 1481 10340 1533
rect 11165 1744 11217 1796
rect 11269 1744 11321 1796
rect 11165 1640 11217 1692
rect 11269 1640 11321 1692
rect 14672 2164 14724 2216
rect 14672 2060 14724 2112
rect 15312 2164 15364 2216
rect 15312 2060 15364 2112
rect 15952 2164 16004 2216
rect 15952 2060 16004 2112
rect 6581 753 6633 805
rect 6581 649 6633 701
rect 7221 753 7273 805
rect 8944 1214 8996 1266
rect 8944 1110 8996 1162
rect 9840 1214 9892 1266
rect 9840 1110 9892 1162
rect 10128 1214 10180 1266
rect 10128 1110 10180 1162
rect 7221 649 7273 701
rect 10128 552 10180 604
rect 10128 448 10180 500
rect 6261 352 6313 404
rect 6261 248 6313 300
rect 6901 352 6953 404
rect 6901 248 6953 300
rect 7541 352 7593 404
rect 7541 248 7593 300
rect 8944 352 8996 404
rect 8944 248 8996 300
rect 9840 352 9892 404
rect 9840 248 9892 300
rect 6261 -248 6313 -196
rect 6261 -352 6313 -300
rect 6901 -248 6953 -196
rect 6901 -352 6953 -300
rect 7541 -248 7593 -196
rect 7541 -352 7593 -300
rect 8496 -248 8548 -196
rect 8496 -352 8548 -300
rect 9392 -248 9444 -196
rect 9392 -352 9444 -300
rect 10288 -248 10340 -196
rect 10288 -352 10340 -300
rect 6581 -521 6633 -469
rect 6581 -625 6633 -573
rect 7221 -521 7273 -469
rect 7221 -625 7273 -573
rect 6581 -986 6633 -934
rect 6581 -1090 6633 -1038
rect 7515 -696 7567 -693
rect 7515 -742 7518 -696
rect 7518 -742 7564 -696
rect 7564 -742 7567 -696
rect 7515 -745 7567 -742
rect 7515 -800 7567 -797
rect 7515 -846 7518 -800
rect 7518 -846 7564 -800
rect 7564 -846 7567 -800
rect 7515 -849 7567 -846
rect 10000 -506 10052 -454
rect 10000 -610 10052 -558
rect 7221 -986 7273 -934
rect 7221 -1090 7273 -1038
rect 10248 -707 10300 -704
rect 10248 -753 10251 -707
rect 10251 -753 10297 -707
rect 10297 -753 10300 -707
rect 10248 -756 10300 -753
rect 10248 -811 10300 -808
rect 10248 -857 10251 -811
rect 10251 -857 10297 -811
rect 10297 -857 10300 -811
rect 10248 -860 10300 -857
rect 8944 -986 8996 -934
rect 8944 -1090 8996 -1038
rect 9840 -986 9892 -934
rect 9840 -1090 9892 -1038
rect 10000 -986 10052 -934
rect 10000 -1090 10052 -1038
rect 6261 -1378 6313 -1326
rect 6261 -1482 6313 -1430
rect 6901 -1378 6953 -1326
rect 6901 -1482 6953 -1430
rect 7541 -1378 7593 -1326
rect 7541 -1482 7593 -1430
rect 8496 -1378 8548 -1326
rect 8496 -1482 8548 -1430
rect 6393 -1830 6445 -1778
rect 6497 -1830 6549 -1778
rect 9392 -1378 9444 -1326
rect 9392 -1482 9444 -1430
rect 10288 -1378 10340 -1326
rect 10288 -1482 10340 -1430
rect 9495 -1830 9547 -1778
rect 9599 -1830 9651 -1778
rect 6393 -1934 6445 -1882
rect 6497 -1934 6549 -1882
rect 9495 -1934 9547 -1882
rect 9599 -1934 9651 -1882
rect 11878 1744 11930 1796
rect 11878 1640 11930 1692
rect 12774 1744 12826 1796
rect 12774 1640 12826 1692
rect 13670 1744 13722 1796
rect 13670 1640 13722 1692
rect 12326 1110 12378 1162
rect 12326 1006 12378 1058
rect 14992 1744 15044 1796
rect 14992 1640 15044 1692
rect 15632 1744 15684 1796
rect 15632 1640 15684 1692
rect 16891 2164 16943 2216
rect 16995 2164 17047 2216
rect 16891 2060 16943 2112
rect 16995 2060 17047 2112
rect 13222 1110 13274 1162
rect 13222 1006 13274 1058
rect 13510 1084 13562 1136
rect 13510 980 13562 1032
rect 16629 1744 16681 1796
rect 16733 1744 16785 1796
rect 16629 1640 16681 1692
rect 16733 1640 16785 1692
rect 14672 1084 14724 1136
rect 14672 980 14724 1032
rect 15312 1084 15364 1136
rect 15312 980 15364 1032
rect 15952 1084 16004 1136
rect 15952 980 16004 1032
rect 11878 64 11930 116
rect 11878 -40 11930 12
rect 12774 64 12826 116
rect 12774 -40 12826 12
rect 13670 64 13722 116
rect 13670 -40 13722 12
rect 13382 -336 13434 -284
rect 13382 -440 13434 -388
rect 11914 -597 11966 -594
rect 11914 -643 11917 -597
rect 11917 -643 11963 -597
rect 11963 -643 11966 -597
rect 11914 -646 11966 -643
rect 11914 -701 11966 -698
rect 11914 -747 11917 -701
rect 11917 -747 11963 -701
rect 11963 -747 11966 -701
rect 11914 -750 11966 -747
rect 14992 -336 15044 -284
rect 14992 -440 15044 -388
rect 15632 -336 15684 -284
rect 15632 -440 15684 -388
rect 12326 -986 12378 -934
rect 12326 -1090 12378 -1038
rect 13222 -986 13274 -934
rect 13222 -1090 13274 -1038
rect 13382 -986 13434 -934
rect 13382 -1090 13434 -1038
rect 14700 -592 14752 -589
rect 14700 -638 14703 -592
rect 14703 -638 14749 -592
rect 14749 -638 14752 -592
rect 14700 -641 14752 -638
rect 14700 -696 14752 -693
rect 14700 -742 14703 -696
rect 14703 -742 14749 -696
rect 14749 -742 14752 -696
rect 14700 -745 14752 -742
rect 14992 -986 15044 -934
rect 14992 -1090 15044 -1038
rect 15632 -986 15684 -934
rect 15632 -1090 15684 -1038
rect 11878 -1386 11930 -1334
rect 11878 -1490 11930 -1438
rect 12774 -1386 12826 -1334
rect 12774 -1490 12826 -1438
rect 13670 -1386 13722 -1334
rect 13670 -1490 13722 -1438
rect 14672 -1376 14724 -1324
rect 14672 -1480 14724 -1428
rect 15312 -1376 15364 -1324
rect 15312 -1480 15364 -1428
rect 15952 -1376 16004 -1324
rect 15952 -1480 16004 -1428
rect 18591 3279 18643 3282
rect 18591 3233 18594 3279
rect 18594 3233 18640 3279
rect 18640 3233 18643 3279
rect 18591 3230 18643 3233
rect 18831 3019 18883 3071
rect 18831 2915 18883 2967
rect 19471 3019 19523 3071
rect 19471 2915 19523 2967
rect 18511 2625 18563 2677
rect 18511 2521 18563 2573
rect 18671 2625 18723 2677
rect 18671 2521 18723 2573
rect 18991 2625 19043 2677
rect 18991 2521 19043 2573
rect 19151 2625 19203 2677
rect 19151 2521 19203 2573
rect 19311 2625 19363 2677
rect 19311 2521 19363 2573
rect 19631 2625 19683 2677
rect 19631 2521 19683 2573
rect 19791 2625 19843 2677
rect 19791 2521 19843 2573
rect 18591 2343 18643 2346
rect 18591 2297 18594 2343
rect 18594 2297 18640 2343
rect 18640 2297 18643 2343
rect 18591 2294 18643 2297
rect 18831 2083 18883 2135
rect 18831 1979 18883 2031
rect 19471 2083 19523 2135
rect 19471 1979 19523 2031
rect 18511 1689 18563 1741
rect 18511 1585 18563 1637
rect 18671 1689 18723 1741
rect 18671 1585 18723 1637
rect 18991 1689 19043 1741
rect 18991 1585 19043 1637
rect 19151 1689 19203 1741
rect 19151 1585 19203 1637
rect 19311 1689 19363 1741
rect 19311 1585 19363 1637
rect 19631 1689 19683 1741
rect 19631 1585 19683 1637
rect 19791 1689 19843 1741
rect 19791 1585 19843 1637
rect 18831 1147 18883 1199
rect 18831 1043 18883 1095
rect 19471 1147 19523 1199
rect 19471 1043 19523 1095
rect 18511 753 18563 805
rect 18511 649 18563 701
rect 19151 753 19203 805
rect 19151 649 19203 701
rect 19791 753 19843 805
rect 19791 649 19843 701
rect 18591 471 18643 474
rect 18591 425 18594 471
rect 18594 425 18640 471
rect 18640 425 18643 471
rect 18591 422 18643 425
rect 18831 211 18883 263
rect 18831 107 18883 159
rect 19471 211 19523 263
rect 19471 107 19523 159
rect 18511 -183 18563 -131
rect 18511 -287 18563 -235
rect 18671 -183 18723 -131
rect 18671 -287 18723 -235
rect 18991 -183 19043 -131
rect 18991 -287 19043 -235
rect 19151 -183 19203 -131
rect 19151 -287 19203 -235
rect 19311 -183 19363 -131
rect 19311 -287 19363 -235
rect 19631 -183 19683 -131
rect 19631 -287 19683 -235
rect 19791 -183 19843 -131
rect 19791 -287 19843 -235
rect 18591 -465 18643 -462
rect 18591 -511 18594 -465
rect 18594 -511 18640 -465
rect 18640 -511 18643 -465
rect 18591 -514 18643 -511
rect 18831 -725 18883 -673
rect 18831 -829 18883 -777
rect 19471 -725 19523 -673
rect 19471 -829 19523 -777
rect 18511 -1119 18563 -1067
rect 18511 -1223 18563 -1171
rect 18671 -1119 18723 -1067
rect 18671 -1223 18723 -1171
rect 18991 -1119 19043 -1067
rect 18991 -1223 19043 -1171
rect 19151 -1119 19203 -1067
rect 19151 -1223 19203 -1171
rect 19311 -1119 19363 -1067
rect 19311 -1223 19363 -1171
rect 19631 -1119 19683 -1067
rect 19631 -1223 19683 -1171
rect 19791 -1119 19843 -1067
rect 19791 -1223 19843 -1171
rect 18751 -1401 18803 -1398
rect 19391 -1401 19443 -1398
rect 18751 -1447 18754 -1401
rect 18754 -1447 18800 -1401
rect 18800 -1447 18803 -1401
rect 19391 -1447 19394 -1401
rect 19394 -1447 19440 -1401
rect 19440 -1447 19443 -1401
rect 18751 -1450 18803 -1447
rect 19391 -1450 19443 -1447
rect 23743 4245 23795 4248
rect 24863 4245 24915 4248
rect 23743 4199 23746 4245
rect 23746 4199 23792 4245
rect 23792 4199 23795 4245
rect 24863 4199 24866 4245
rect 24866 4199 24912 4245
rect 24912 4199 24915 4245
rect 23743 4196 23795 4199
rect 24863 4196 24915 4199
rect 23983 3955 24035 4007
rect 23983 3851 24035 3903
rect 24623 3955 24675 4007
rect 24623 3851 24675 3903
rect 23663 3561 23715 3613
rect 23663 3457 23715 3509
rect 23823 3561 23875 3613
rect 23823 3457 23875 3509
rect 24143 3561 24195 3613
rect 24143 3457 24195 3509
rect 24303 3561 24355 3613
rect 24303 3457 24355 3509
rect 24463 3561 24515 3613
rect 24463 3457 24515 3509
rect 24783 3561 24835 3613
rect 24783 3457 24835 3509
rect 24943 3561 24995 3613
rect 24943 3457 24995 3509
rect 24863 3279 24915 3282
rect 24863 3233 24866 3279
rect 24866 3233 24912 3279
rect 24912 3233 24915 3279
rect 24863 3230 24915 3233
rect 23983 3019 24035 3071
rect 23983 2915 24035 2967
rect 24623 3019 24675 3071
rect 24623 2915 24675 2967
rect 23663 2625 23715 2677
rect 23663 2521 23715 2573
rect 23823 2625 23875 2677
rect 23823 2521 23875 2573
rect 24143 2625 24195 2677
rect 24143 2521 24195 2573
rect 24303 2625 24355 2677
rect 24303 2521 24355 2573
rect 24463 2625 24515 2677
rect 24463 2521 24515 2573
rect 24783 2625 24835 2677
rect 24783 2521 24835 2573
rect 24943 2625 24995 2677
rect 24943 2521 24995 2573
rect 24863 2343 24915 2346
rect 24863 2297 24866 2343
rect 24866 2297 24912 2343
rect 24912 2297 24915 2343
rect 24863 2294 24915 2297
rect 23983 2083 24035 2135
rect 23983 1979 24035 2031
rect 24623 2083 24675 2135
rect 24623 1979 24675 2031
rect 23663 1689 23715 1741
rect 23663 1585 23715 1637
rect 23823 1689 23875 1741
rect 23823 1585 23875 1637
rect 24143 1689 24195 1741
rect 24143 1585 24195 1637
rect 24303 1689 24355 1741
rect 24303 1585 24355 1637
rect 24463 1689 24515 1741
rect 24463 1585 24515 1637
rect 24783 1689 24835 1741
rect 24783 1585 24835 1637
rect 24943 1689 24995 1741
rect 24943 1585 24995 1637
rect 23983 1147 24035 1199
rect 23983 1043 24035 1095
rect 24623 1147 24675 1199
rect 24623 1043 24675 1095
rect 23663 753 23715 805
rect 23663 649 23715 701
rect 24303 753 24355 805
rect 24303 649 24355 701
rect 24943 753 24995 805
rect 24943 649 24995 701
rect 24863 471 24915 474
rect 24863 425 24866 471
rect 24866 425 24912 471
rect 24912 425 24915 471
rect 24863 422 24915 425
rect 23983 211 24035 263
rect 23983 107 24035 159
rect 24623 211 24675 263
rect 24623 107 24675 159
rect 23663 -183 23715 -131
rect 23663 -287 23715 -235
rect 23823 -183 23875 -131
rect 23823 -287 23875 -235
rect 24143 -183 24195 -131
rect 24143 -287 24195 -235
rect 24303 -183 24355 -131
rect 24303 -287 24355 -235
rect 24463 -183 24515 -131
rect 24463 -287 24515 -235
rect 24783 -183 24835 -131
rect 24783 -287 24835 -235
rect 24943 -183 24995 -131
rect 24943 -287 24995 -235
rect 24863 -465 24915 -462
rect 24863 -511 24866 -465
rect 24866 -511 24912 -465
rect 24912 -511 24915 -465
rect 24863 -514 24915 -511
rect 23983 -725 24035 -673
rect 23983 -829 24035 -777
rect 24623 -725 24675 -673
rect 24623 -829 24675 -777
rect 23663 -1119 23715 -1067
rect 23663 -1223 23715 -1171
rect 23823 -1119 23875 -1067
rect 23823 -1223 23875 -1171
rect 24143 -1119 24195 -1067
rect 24143 -1223 24195 -1171
rect 24303 -1119 24355 -1067
rect 24303 -1223 24355 -1171
rect 24463 -1119 24515 -1067
rect 24463 -1223 24515 -1171
rect 24783 -1119 24835 -1067
rect 24783 -1223 24835 -1171
rect 24943 -1119 24995 -1067
rect 24943 -1223 24995 -1171
rect 24063 -1401 24115 -1398
rect 24703 -1401 24755 -1398
rect 24063 -1447 24066 -1401
rect 24066 -1447 24112 -1401
rect 24112 -1447 24115 -1401
rect 24703 -1447 24706 -1401
rect 24706 -1447 24752 -1401
rect 24752 -1447 24755 -1401
rect 24063 -1450 24115 -1447
rect 24703 -1450 24755 -1447
rect 27712 4245 27764 4248
rect 27712 4199 27715 4245
rect 27715 4199 27761 4245
rect 27761 4199 27764 4245
rect 27712 4196 27764 4199
rect 27952 3955 28004 4007
rect 27952 3851 28004 3903
rect 28592 3955 28644 4007
rect 28592 3851 28644 3903
rect 27632 3561 27684 3613
rect 27632 3457 27684 3509
rect 27792 3561 27844 3613
rect 27792 3457 27844 3509
rect 28112 3561 28164 3613
rect 28112 3457 28164 3509
rect 28272 3561 28324 3613
rect 28272 3457 28324 3509
rect 28432 3561 28484 3613
rect 28432 3457 28484 3509
rect 28752 3561 28804 3613
rect 28752 3457 28804 3509
rect 28912 3561 28964 3613
rect 28912 3457 28964 3509
rect 27712 3279 27764 3282
rect 27712 3233 27715 3279
rect 27715 3233 27761 3279
rect 27761 3233 27764 3279
rect 27712 3230 27764 3233
rect 27952 3019 28004 3071
rect 27952 2915 28004 2967
rect 28592 3019 28644 3071
rect 28592 2915 28644 2967
rect 27632 2625 27684 2677
rect 27632 2521 27684 2573
rect 27792 2625 27844 2677
rect 27792 2521 27844 2573
rect 28112 2625 28164 2677
rect 28112 2521 28164 2573
rect 28272 2625 28324 2677
rect 28272 2521 28324 2573
rect 28432 2625 28484 2677
rect 28432 2521 28484 2573
rect 28752 2625 28804 2677
rect 28752 2521 28804 2573
rect 28912 2625 28964 2677
rect 28912 2521 28964 2573
rect 27712 2343 27764 2346
rect 27712 2297 27715 2343
rect 27715 2297 27761 2343
rect 27761 2297 27764 2343
rect 27712 2294 27764 2297
rect 27952 2083 28004 2135
rect 27952 1979 28004 2031
rect 28592 2083 28644 2135
rect 28592 1979 28644 2031
rect 27632 1689 27684 1741
rect 27632 1585 27684 1637
rect 27792 1689 27844 1741
rect 27792 1585 27844 1637
rect 28112 1689 28164 1741
rect 28112 1585 28164 1637
rect 28272 1689 28324 1741
rect 28272 1585 28324 1637
rect 28432 1689 28484 1741
rect 28432 1585 28484 1637
rect 28752 1689 28804 1741
rect 28752 1585 28804 1637
rect 28912 1689 28964 1741
rect 28912 1585 28964 1637
rect 27952 1147 28004 1199
rect 27952 1043 28004 1095
rect 28592 1147 28644 1199
rect 28592 1043 28644 1095
rect 27632 753 27684 805
rect 27632 649 27684 701
rect 28272 753 28324 805
rect 28272 649 28324 701
rect 28912 753 28964 805
rect 28912 649 28964 701
rect 27712 471 27764 474
rect 27712 425 27715 471
rect 27715 425 27761 471
rect 27761 425 27764 471
rect 27712 422 27764 425
rect 27952 211 28004 263
rect 27952 107 28004 159
rect 28592 211 28644 263
rect 28592 107 28644 159
rect 27632 -183 27684 -131
rect 27632 -287 27684 -235
rect 27792 -183 27844 -131
rect 27792 -287 27844 -235
rect 28112 -183 28164 -131
rect 28112 -287 28164 -235
rect 28272 -183 28324 -131
rect 28272 -287 28324 -235
rect 28432 -183 28484 -131
rect 28432 -287 28484 -235
rect 28752 -183 28804 -131
rect 28752 -287 28804 -235
rect 28912 -183 28964 -131
rect 28912 -287 28964 -235
rect 27712 -465 27764 -462
rect 27712 -511 27715 -465
rect 27715 -511 27761 -465
rect 27761 -511 27764 -465
rect 27712 -514 27764 -511
rect 27952 -725 28004 -673
rect 27952 -829 28004 -777
rect 28592 -725 28644 -673
rect 28592 -829 28644 -777
rect 27632 -1119 27684 -1067
rect 27632 -1223 27684 -1171
rect 27792 -1119 27844 -1067
rect 27792 -1223 27844 -1171
rect 28112 -1119 28164 -1067
rect 28112 -1223 28164 -1171
rect 28272 -1119 28324 -1067
rect 28272 -1223 28324 -1171
rect 28432 -1119 28484 -1067
rect 28432 -1223 28484 -1171
rect 28752 -1119 28804 -1067
rect 28752 -1223 28804 -1171
rect 28912 -1119 28964 -1067
rect 28912 -1223 28964 -1171
rect 27872 -1401 27924 -1398
rect 27872 -1447 27875 -1401
rect 27875 -1447 27921 -1401
rect 27921 -1447 27924 -1401
rect 27872 -1450 27924 -1447
rect 66440 3839 66492 3891
rect 66544 3839 66596 3891
rect 66648 3839 66700 3891
rect 66440 3735 66492 3787
rect 66544 3735 66596 3787
rect 66648 3735 66700 3787
rect 66440 3631 66492 3683
rect 66544 3631 66596 3683
rect 66648 3631 66700 3683
rect 32928 2061 32980 2113
rect 32928 1957 32980 2009
rect 32928 1001 32980 1053
rect 32928 897 32980 949
rect 32928 -59 32980 -7
rect 32928 -163 32980 -111
rect 32928 -1119 32980 -1067
rect 32928 -1223 32980 -1171
rect 33249 2455 33301 2507
rect 33249 2351 33301 2403
rect 33249 1395 33301 1447
rect 33249 1291 33301 1343
rect 33249 335 33301 387
rect 33249 231 33301 283
rect 33249 -725 33301 -673
rect 33249 -829 33301 -777
rect 33568 2061 33620 2113
rect 33568 1957 33620 2009
rect 34128 2652 34180 2655
rect 34288 2652 34340 2655
rect 34128 2606 34131 2652
rect 34131 2606 34177 2652
rect 34177 2606 34180 2652
rect 34128 2603 34180 2606
rect 34288 2606 34291 2652
rect 34291 2606 34337 2652
rect 34337 2606 34340 2652
rect 34288 2603 34340 2606
rect 33889 2455 33941 2507
rect 33889 2351 33941 2403
rect 34529 2455 34581 2507
rect 34529 2351 34581 2403
rect 33568 1001 33620 1053
rect 33568 897 33620 949
rect 34128 1592 34180 1595
rect 34288 1592 34340 1595
rect 34128 1546 34131 1592
rect 34131 1546 34177 1592
rect 34177 1546 34180 1592
rect 34128 1543 34180 1546
rect 34288 1546 34291 1592
rect 34291 1546 34337 1592
rect 34337 1546 34340 1592
rect 34288 1543 34340 1546
rect 33889 1395 33941 1447
rect 33889 1291 33941 1343
rect 34529 1395 34581 1447
rect 34529 1291 34581 1343
rect 33568 -59 33620 -7
rect 33568 -163 33620 -111
rect 34128 532 34180 535
rect 34288 532 34340 535
rect 34128 486 34131 532
rect 34131 486 34177 532
rect 34177 486 34180 532
rect 34128 483 34180 486
rect 34288 486 34291 532
rect 34291 486 34337 532
rect 34337 486 34340 532
rect 34288 483 34340 486
rect 33889 335 33941 387
rect 33889 231 33941 283
rect 34529 335 34581 387
rect 34529 231 34581 283
rect 33568 -1119 33620 -1067
rect 33568 -1223 33620 -1171
rect 34128 -528 34180 -525
rect 34288 -528 34340 -525
rect 34128 -574 34131 -528
rect 34131 -574 34177 -528
rect 34177 -574 34180 -528
rect 34128 -577 34180 -574
rect 34288 -574 34291 -528
rect 34291 -574 34337 -528
rect 34337 -574 34340 -528
rect 34288 -577 34340 -574
rect 33889 -725 33941 -673
rect 33889 -829 33941 -777
rect 34529 -725 34581 -673
rect 34529 -829 34581 -777
rect 34848 2061 34900 2113
rect 34848 1957 34900 2009
rect 34848 1001 34900 1053
rect 34848 897 34900 949
rect 34848 -59 34900 -7
rect 34848 -163 34900 -111
rect 34848 -1119 34900 -1067
rect 34848 -1223 34900 -1171
rect 35169 2455 35221 2507
rect 35169 2351 35221 2403
rect 35169 1395 35221 1447
rect 35169 1291 35221 1343
rect 35169 335 35221 387
rect 35169 231 35221 283
rect 35169 -725 35221 -673
rect 35169 -829 35221 -777
rect 35488 2061 35540 2113
rect 35488 1957 35540 2009
rect 35488 1001 35540 1053
rect 35488 897 35540 949
rect 35488 -59 35540 -7
rect 35488 -163 35540 -111
rect 35488 -1119 35540 -1067
rect 35488 -1223 35540 -1171
rect 37064 2061 37116 2113
rect 37064 1957 37116 2009
rect 37064 1001 37116 1053
rect 37064 897 37116 949
rect 37064 -59 37116 -7
rect 37064 -163 37116 -111
rect 37064 -1119 37116 -1067
rect 37064 -1223 37116 -1171
rect 37383 2455 37435 2507
rect 37383 2351 37435 2403
rect 37383 1395 37435 1447
rect 37383 1291 37435 1343
rect 37383 335 37435 387
rect 37383 231 37435 283
rect 37383 -725 37435 -673
rect 37383 -829 37435 -777
rect 37704 2061 37756 2113
rect 37704 1957 37756 2009
rect 37704 1001 37756 1053
rect 37704 897 37756 949
rect 37704 -59 37756 -7
rect 37704 -163 37756 -111
rect 37704 -1119 37756 -1067
rect 37704 -1223 37756 -1171
rect 38264 2652 38316 2655
rect 38424 2652 38476 2655
rect 38264 2606 38267 2652
rect 38267 2606 38313 2652
rect 38313 2606 38316 2652
rect 38264 2603 38316 2606
rect 38424 2606 38427 2652
rect 38427 2606 38473 2652
rect 38473 2606 38476 2652
rect 38424 2603 38476 2606
rect 38023 2455 38075 2507
rect 38023 2351 38075 2403
rect 38663 2455 38715 2507
rect 38663 2351 38715 2403
rect 38984 2061 39036 2113
rect 38984 1957 39036 2009
rect 38264 1592 38316 1595
rect 38424 1592 38476 1595
rect 38264 1546 38267 1592
rect 38267 1546 38313 1592
rect 38313 1546 38316 1592
rect 38264 1543 38316 1546
rect 38424 1546 38427 1592
rect 38427 1546 38473 1592
rect 38473 1546 38476 1592
rect 38424 1543 38476 1546
rect 38023 1395 38075 1447
rect 38023 1291 38075 1343
rect 38663 1395 38715 1447
rect 38663 1291 38715 1343
rect 38984 1001 39036 1053
rect 38984 897 39036 949
rect 38264 532 38316 535
rect 38424 532 38476 535
rect 38264 486 38267 532
rect 38267 486 38313 532
rect 38313 486 38316 532
rect 38264 483 38316 486
rect 38424 486 38427 532
rect 38427 486 38473 532
rect 38473 486 38476 532
rect 38424 483 38476 486
rect 38023 335 38075 387
rect 38023 231 38075 283
rect 38663 335 38715 387
rect 38663 231 38715 283
rect 38984 -59 39036 -7
rect 38984 -163 39036 -111
rect 38264 -528 38316 -525
rect 38424 -528 38476 -525
rect 38264 -574 38267 -528
rect 38267 -574 38313 -528
rect 38313 -574 38316 -528
rect 38264 -577 38316 -574
rect 38424 -574 38427 -528
rect 38427 -574 38473 -528
rect 38473 -574 38476 -528
rect 38424 -577 38476 -574
rect 38023 -725 38075 -673
rect 38023 -829 38075 -777
rect 38663 -725 38715 -673
rect 38663 -829 38715 -777
rect 38984 -1119 39036 -1067
rect 38984 -1223 39036 -1171
rect 39303 2455 39355 2507
rect 39303 2351 39355 2403
rect 39303 1395 39355 1447
rect 39303 1291 39355 1343
rect 39303 335 39355 387
rect 39303 231 39355 283
rect 39303 -725 39355 -673
rect 39303 -829 39355 -777
rect 39624 2061 39676 2113
rect 39624 1957 39676 2009
rect 39624 1001 39676 1053
rect 39624 897 39676 949
rect 39624 -59 39676 -7
rect 39624 -163 39676 -111
rect 39624 -1119 39676 -1067
rect 39624 -1223 39676 -1171
rect 42624 2061 42676 2113
rect 42624 1957 42676 2009
rect 42624 1001 42676 1053
rect 42624 897 42676 949
rect 42624 -59 42676 -7
rect 42624 -163 42676 -111
rect 42624 -1119 42676 -1067
rect 42624 -1223 42676 -1171
rect 42945 2455 42997 2507
rect 42945 2351 42997 2403
rect 42945 1395 42997 1447
rect 42945 1291 42997 1343
rect 42945 335 42997 387
rect 42945 231 42997 283
rect 42945 -725 42997 -673
rect 42945 -829 42997 -777
rect 43264 2061 43316 2113
rect 43264 1957 43316 2009
rect 43824 2652 43876 2655
rect 43984 2652 44036 2655
rect 43824 2606 43827 2652
rect 43827 2606 43873 2652
rect 43873 2606 43876 2652
rect 43824 2603 43876 2606
rect 43984 2606 43987 2652
rect 43987 2606 44033 2652
rect 44033 2606 44036 2652
rect 43984 2603 44036 2606
rect 43585 2455 43637 2507
rect 43585 2351 43637 2403
rect 44225 2455 44277 2507
rect 44225 2351 44277 2403
rect 43264 1001 43316 1053
rect 43264 897 43316 949
rect 43824 1592 43876 1595
rect 43984 1592 44036 1595
rect 43824 1546 43827 1592
rect 43827 1546 43873 1592
rect 43873 1546 43876 1592
rect 43824 1543 43876 1546
rect 43984 1546 43987 1592
rect 43987 1546 44033 1592
rect 44033 1546 44036 1592
rect 43984 1543 44036 1546
rect 43585 1395 43637 1447
rect 43585 1291 43637 1343
rect 44225 1395 44277 1447
rect 44225 1291 44277 1343
rect 43264 -59 43316 -7
rect 43264 -163 43316 -111
rect 43824 532 43876 535
rect 43984 532 44036 535
rect 43824 486 43827 532
rect 43827 486 43873 532
rect 43873 486 43876 532
rect 43824 483 43876 486
rect 43984 486 43987 532
rect 43987 486 44033 532
rect 44033 486 44036 532
rect 43984 483 44036 486
rect 43585 335 43637 387
rect 43585 231 43637 283
rect 44225 335 44277 387
rect 44225 231 44277 283
rect 43264 -1119 43316 -1067
rect 43264 -1223 43316 -1171
rect 43824 -528 43876 -525
rect 43984 -528 44036 -525
rect 43824 -574 43827 -528
rect 43827 -574 43873 -528
rect 43873 -574 43876 -528
rect 43824 -577 43876 -574
rect 43984 -574 43987 -528
rect 43987 -574 44033 -528
rect 44033 -574 44036 -528
rect 43984 -577 44036 -574
rect 43585 -725 43637 -673
rect 43585 -829 43637 -777
rect 44225 -725 44277 -673
rect 44225 -829 44277 -777
rect 44544 2061 44596 2113
rect 44544 1957 44596 2009
rect 44544 1001 44596 1053
rect 44544 897 44596 949
rect 44544 -59 44596 -7
rect 44544 -163 44596 -111
rect 44544 -1119 44596 -1067
rect 44544 -1223 44596 -1171
rect 44865 2455 44917 2507
rect 44865 2351 44917 2403
rect 44865 1395 44917 1447
rect 44865 1291 44917 1343
rect 44865 335 44917 387
rect 44865 231 44917 283
rect 44865 -725 44917 -673
rect 44865 -829 44917 -777
rect 45184 2061 45236 2113
rect 45184 1957 45236 2009
rect 45184 1001 45236 1053
rect 45184 897 45236 949
rect 45184 -59 45236 -7
rect 45184 -163 45236 -111
rect 45184 -1119 45236 -1067
rect 45184 -1223 45236 -1171
rect 46760 2061 46812 2113
rect 46760 1957 46812 2009
rect 46760 1001 46812 1053
rect 46760 897 46812 949
rect 46760 -59 46812 -7
rect 46760 -163 46812 -111
rect 46760 -1119 46812 -1067
rect 46760 -1223 46812 -1171
rect 47079 2455 47131 2507
rect 47079 2351 47131 2403
rect 47079 1395 47131 1447
rect 47079 1291 47131 1343
rect 47079 335 47131 387
rect 47079 231 47131 283
rect 47079 -725 47131 -673
rect 47079 -829 47131 -777
rect 47400 2061 47452 2113
rect 47400 1957 47452 2009
rect 47400 1001 47452 1053
rect 47400 897 47452 949
rect 47400 -59 47452 -7
rect 47400 -163 47452 -111
rect 47400 -1119 47452 -1067
rect 47400 -1223 47452 -1171
rect 47960 2652 48012 2655
rect 48120 2652 48172 2655
rect 47960 2606 47963 2652
rect 47963 2606 48009 2652
rect 48009 2606 48012 2652
rect 47960 2603 48012 2606
rect 48120 2606 48123 2652
rect 48123 2606 48169 2652
rect 48169 2606 48172 2652
rect 48120 2603 48172 2606
rect 47719 2455 47771 2507
rect 47719 2351 47771 2403
rect 48359 2455 48411 2507
rect 48359 2351 48411 2403
rect 48680 2061 48732 2113
rect 48680 1957 48732 2009
rect 47960 1592 48012 1595
rect 48120 1592 48172 1595
rect 47960 1546 47963 1592
rect 47963 1546 48009 1592
rect 48009 1546 48012 1592
rect 47960 1543 48012 1546
rect 48120 1546 48123 1592
rect 48123 1546 48169 1592
rect 48169 1546 48172 1592
rect 48120 1543 48172 1546
rect 47719 1395 47771 1447
rect 47719 1291 47771 1343
rect 48359 1395 48411 1447
rect 48359 1291 48411 1343
rect 48680 1001 48732 1053
rect 48680 897 48732 949
rect 47960 532 48012 535
rect 48120 532 48172 535
rect 47960 486 47963 532
rect 47963 486 48009 532
rect 48009 486 48012 532
rect 47960 483 48012 486
rect 48120 486 48123 532
rect 48123 486 48169 532
rect 48169 486 48172 532
rect 48120 483 48172 486
rect 47719 335 47771 387
rect 47719 231 47771 283
rect 48359 335 48411 387
rect 48359 231 48411 283
rect 48680 -59 48732 -7
rect 48680 -163 48732 -111
rect 47960 -528 48012 -525
rect 48120 -528 48172 -525
rect 47960 -574 47963 -528
rect 47963 -574 48009 -528
rect 48009 -574 48012 -528
rect 47960 -577 48012 -574
rect 48120 -574 48123 -528
rect 48123 -574 48169 -528
rect 48169 -574 48172 -528
rect 48120 -577 48172 -574
rect 47719 -725 47771 -673
rect 47719 -829 47771 -777
rect 48359 -725 48411 -673
rect 48359 -829 48411 -777
rect 48680 -1119 48732 -1067
rect 48680 -1223 48732 -1171
rect 48999 2455 49051 2507
rect 48999 2351 49051 2403
rect 48999 1395 49051 1447
rect 48999 1291 49051 1343
rect 48999 335 49051 387
rect 48999 231 49051 283
rect 48999 -725 49051 -673
rect 48999 -829 49051 -777
rect 49320 2061 49372 2113
rect 49320 1957 49372 2009
rect 49320 1001 49372 1053
rect 49320 897 49372 949
rect 49320 -59 49372 -7
rect 49320 -163 49372 -111
rect 49320 -1119 49372 -1067
rect 49320 -1223 49372 -1171
rect 52320 2061 52372 2113
rect 52320 1957 52372 2009
rect 52320 1001 52372 1053
rect 52320 897 52372 949
rect 52320 -59 52372 -7
rect 52320 -163 52372 -111
rect 52320 -1119 52372 -1067
rect 52320 -1223 52372 -1171
rect 52641 2455 52693 2507
rect 52641 2351 52693 2403
rect 52641 1395 52693 1447
rect 52641 1291 52693 1343
rect 52641 335 52693 387
rect 52641 231 52693 283
rect 52641 -725 52693 -673
rect 52641 -829 52693 -777
rect 52960 2061 53012 2113
rect 52960 1957 53012 2009
rect 53520 2652 53572 2655
rect 53680 2652 53732 2655
rect 53520 2606 53523 2652
rect 53523 2606 53569 2652
rect 53569 2606 53572 2652
rect 53520 2603 53572 2606
rect 53680 2606 53683 2652
rect 53683 2606 53729 2652
rect 53729 2606 53732 2652
rect 53680 2603 53732 2606
rect 53281 2455 53333 2507
rect 53281 2351 53333 2403
rect 53921 2455 53973 2507
rect 53921 2351 53973 2403
rect 52960 1001 53012 1053
rect 52960 897 53012 949
rect 53520 1592 53572 1595
rect 53680 1592 53732 1595
rect 53520 1546 53523 1592
rect 53523 1546 53569 1592
rect 53569 1546 53572 1592
rect 53520 1543 53572 1546
rect 53680 1546 53683 1592
rect 53683 1546 53729 1592
rect 53729 1546 53732 1592
rect 53680 1543 53732 1546
rect 53281 1395 53333 1447
rect 53281 1291 53333 1343
rect 53921 1395 53973 1447
rect 53921 1291 53973 1343
rect 52960 -59 53012 -7
rect 52960 -163 53012 -111
rect 53520 532 53572 535
rect 53680 532 53732 535
rect 53520 486 53523 532
rect 53523 486 53569 532
rect 53569 486 53572 532
rect 53520 483 53572 486
rect 53680 486 53683 532
rect 53683 486 53729 532
rect 53729 486 53732 532
rect 53680 483 53732 486
rect 53281 335 53333 387
rect 53281 231 53333 283
rect 53921 335 53973 387
rect 53921 231 53973 283
rect 52960 -1119 53012 -1067
rect 52960 -1223 53012 -1171
rect 53520 -528 53572 -525
rect 53680 -528 53732 -525
rect 53520 -574 53523 -528
rect 53523 -574 53569 -528
rect 53569 -574 53572 -528
rect 53520 -577 53572 -574
rect 53680 -574 53683 -528
rect 53683 -574 53729 -528
rect 53729 -574 53732 -528
rect 53680 -577 53732 -574
rect 53281 -725 53333 -673
rect 53281 -829 53333 -777
rect 53921 -725 53973 -673
rect 53921 -829 53973 -777
rect 54240 2061 54292 2113
rect 54240 1957 54292 2009
rect 54240 1001 54292 1053
rect 54240 897 54292 949
rect 54240 -59 54292 -7
rect 54240 -163 54292 -111
rect 54240 -1119 54292 -1067
rect 54240 -1223 54292 -1171
rect 54561 2455 54613 2507
rect 54561 2351 54613 2403
rect 54561 1395 54613 1447
rect 54561 1291 54613 1343
rect 54561 335 54613 387
rect 54561 231 54613 283
rect 54561 -725 54613 -673
rect 54561 -829 54613 -777
rect 54880 2061 54932 2113
rect 54880 1957 54932 2009
rect 54880 1001 54932 1053
rect 54880 897 54932 949
rect 54880 -59 54932 -7
rect 54880 -163 54932 -111
rect 54880 -1119 54932 -1067
rect 54880 -1223 54932 -1171
rect 56456 2061 56508 2113
rect 56456 1957 56508 2009
rect 56456 1001 56508 1053
rect 56456 897 56508 949
rect 56456 -59 56508 -7
rect 56456 -163 56508 -111
rect 56456 -1119 56508 -1067
rect 56456 -1223 56508 -1171
rect 56775 2455 56827 2507
rect 56775 2351 56827 2403
rect 56775 1395 56827 1447
rect 56775 1291 56827 1343
rect 56775 335 56827 387
rect 56775 231 56827 283
rect 56775 -725 56827 -673
rect 56775 -829 56827 -777
rect 57096 2061 57148 2113
rect 57096 1957 57148 2009
rect 57096 1001 57148 1053
rect 57096 897 57148 949
rect 57096 -59 57148 -7
rect 57096 -163 57148 -111
rect 57096 -1119 57148 -1067
rect 57096 -1223 57148 -1171
rect 57656 2652 57708 2655
rect 57816 2652 57868 2655
rect 57656 2606 57659 2652
rect 57659 2606 57705 2652
rect 57705 2606 57708 2652
rect 57656 2603 57708 2606
rect 57816 2606 57819 2652
rect 57819 2606 57865 2652
rect 57865 2606 57868 2652
rect 57816 2603 57868 2606
rect 57415 2455 57467 2507
rect 57415 2351 57467 2403
rect 58055 2455 58107 2507
rect 58055 2351 58107 2403
rect 58376 2061 58428 2113
rect 58376 1957 58428 2009
rect 57656 1592 57708 1595
rect 57816 1592 57868 1595
rect 57656 1546 57659 1592
rect 57659 1546 57705 1592
rect 57705 1546 57708 1592
rect 57656 1543 57708 1546
rect 57816 1546 57819 1592
rect 57819 1546 57865 1592
rect 57865 1546 57868 1592
rect 57816 1543 57868 1546
rect 57415 1395 57467 1447
rect 57415 1291 57467 1343
rect 58055 1395 58107 1447
rect 58055 1291 58107 1343
rect 58376 1001 58428 1053
rect 58376 897 58428 949
rect 57656 532 57708 535
rect 57816 532 57868 535
rect 57656 486 57659 532
rect 57659 486 57705 532
rect 57705 486 57708 532
rect 57656 483 57708 486
rect 57816 486 57819 532
rect 57819 486 57865 532
rect 57865 486 57868 532
rect 57816 483 57868 486
rect 57415 335 57467 387
rect 57415 231 57467 283
rect 58055 335 58107 387
rect 58055 231 58107 283
rect 58376 -59 58428 -7
rect 58376 -163 58428 -111
rect 57656 -528 57708 -525
rect 57816 -528 57868 -525
rect 57656 -574 57659 -528
rect 57659 -574 57705 -528
rect 57705 -574 57708 -528
rect 57656 -577 57708 -574
rect 57816 -574 57819 -528
rect 57819 -574 57865 -528
rect 57865 -574 57868 -528
rect 57816 -577 57868 -574
rect 57415 -725 57467 -673
rect 57415 -829 57467 -777
rect 58055 -725 58107 -673
rect 58055 -829 58107 -777
rect 58376 -1119 58428 -1067
rect 58376 -1223 58428 -1171
rect 58695 2455 58747 2507
rect 58695 2351 58747 2403
rect 58695 1395 58747 1447
rect 58695 1291 58747 1343
rect 58695 335 58747 387
rect 58695 231 58747 283
rect 58695 -725 58747 -673
rect 58695 -829 58747 -777
rect 59016 2061 59068 2113
rect 59016 1957 59068 2009
rect 59016 1001 59068 1053
rect 59016 897 59068 949
rect 59016 -59 59068 -7
rect 59016 -163 59068 -111
rect 59016 -1119 59068 -1067
rect 59016 -1223 59068 -1171
rect 62016 2061 62068 2113
rect 62016 1957 62068 2009
rect 62016 1001 62068 1053
rect 62016 897 62068 949
rect 62016 -59 62068 -7
rect 62016 -163 62068 -111
rect 62016 -1119 62068 -1067
rect 62016 -1223 62068 -1171
rect 62337 2455 62389 2507
rect 62337 2351 62389 2403
rect 62337 1395 62389 1447
rect 62337 1291 62389 1343
rect 62337 335 62389 387
rect 62337 231 62389 283
rect 62337 -725 62389 -673
rect 62337 -829 62389 -777
rect 62656 2061 62708 2113
rect 62656 1957 62708 2009
rect 63216 2652 63268 2655
rect 63376 2652 63428 2655
rect 63216 2606 63219 2652
rect 63219 2606 63265 2652
rect 63265 2606 63268 2652
rect 63216 2603 63268 2606
rect 63376 2606 63379 2652
rect 63379 2606 63425 2652
rect 63425 2606 63428 2652
rect 63376 2603 63428 2606
rect 62977 2455 63029 2507
rect 62977 2351 63029 2403
rect 63617 2455 63669 2507
rect 63617 2351 63669 2403
rect 62656 1001 62708 1053
rect 62656 897 62708 949
rect 63216 1592 63268 1595
rect 63376 1592 63428 1595
rect 63216 1546 63219 1592
rect 63219 1546 63265 1592
rect 63265 1546 63268 1592
rect 63216 1543 63268 1546
rect 63376 1546 63379 1592
rect 63379 1546 63425 1592
rect 63425 1546 63428 1592
rect 63376 1543 63428 1546
rect 62977 1395 63029 1447
rect 62977 1291 63029 1343
rect 63617 1395 63669 1447
rect 63617 1291 63669 1343
rect 62656 -59 62708 -7
rect 62656 -163 62708 -111
rect 63216 532 63268 535
rect 63376 532 63428 535
rect 63216 486 63219 532
rect 63219 486 63265 532
rect 63265 486 63268 532
rect 63216 483 63268 486
rect 63376 486 63379 532
rect 63379 486 63425 532
rect 63425 486 63428 532
rect 63376 483 63428 486
rect 62977 335 63029 387
rect 62977 231 63029 283
rect 63617 335 63669 387
rect 63617 231 63669 283
rect 62656 -1119 62708 -1067
rect 62656 -1223 62708 -1171
rect 63216 -528 63268 -525
rect 63376 -528 63428 -525
rect 63216 -574 63219 -528
rect 63219 -574 63265 -528
rect 63265 -574 63268 -528
rect 63216 -577 63268 -574
rect 63376 -574 63379 -528
rect 63379 -574 63425 -528
rect 63425 -574 63428 -528
rect 63376 -577 63428 -574
rect 62977 -725 63029 -673
rect 62977 -829 63029 -777
rect 63617 -725 63669 -673
rect 63617 -829 63669 -777
rect 63936 2061 63988 2113
rect 63936 1957 63988 2009
rect 63936 1001 63988 1053
rect 63936 897 63988 949
rect 63936 -59 63988 -7
rect 63936 -163 63988 -111
rect 63936 -1119 63988 -1067
rect 63936 -1223 63988 -1171
rect 64257 2455 64309 2507
rect 64257 2351 64309 2403
rect 64257 1395 64309 1447
rect 64257 1291 64309 1343
rect 64257 335 64309 387
rect 64257 231 64309 283
rect 64257 -725 64309 -673
rect 64257 -829 64309 -777
rect 64576 2061 64628 2113
rect 64576 1957 64628 2009
rect 64576 1001 64628 1053
rect 64576 897 64628 949
rect 64576 -59 64628 -7
rect 64576 -163 64628 -111
rect 64576 -1119 64628 -1067
rect 64576 -1223 64628 -1171
rect 1701 -3901 1753 -3849
rect 1805 -3901 1857 -3849
rect 1701 -4005 1753 -3953
rect 1805 -4005 1857 -3953
rect 2573 -4036 2625 -3984
rect 2677 -4036 2729 -3984
rect 2573 -4140 2625 -4088
rect 2677 -4140 2729 -4088
rect 7801 -2800 7853 -2748
rect 7905 -2800 7957 -2748
rect 7801 -2904 7853 -2852
rect 7905 -2904 7957 -2852
rect 10897 -2773 10949 -2721
rect 11001 -2773 11053 -2721
rect 16645 -2773 16697 -2721
rect 16749 -2773 16801 -2721
rect 16853 -2773 16905 -2721
rect 10897 -2877 10949 -2825
rect 11001 -2877 11053 -2825
rect 16645 -2877 16697 -2825
rect 16749 -2877 16801 -2825
rect 16853 -2877 16905 -2825
rect 6393 -3036 6445 -2984
rect 6497 -3036 6549 -2984
rect 9495 -3036 9547 -2984
rect 9599 -3036 9651 -2984
rect 10897 -2981 10949 -2929
rect 11001 -2981 11053 -2929
rect 16645 -2981 16697 -2929
rect 16749 -2981 16801 -2929
rect 16853 -2981 16905 -2929
rect 6393 -3140 6445 -3088
rect 6497 -3140 6549 -3088
rect 9495 -3140 9547 -3088
rect 4670 -3750 4722 -3698
rect 4774 -3750 4826 -3698
rect 4670 -3854 4722 -3802
rect 4774 -3854 4826 -3802
rect 1701 -4604 1753 -4601
rect 1701 -4650 1704 -4604
rect 1704 -4650 1750 -4604
rect 1750 -4650 1753 -4604
rect 1701 -4653 1753 -4650
rect 1805 -4604 1857 -4601
rect 1805 -4650 1808 -4604
rect 1808 -4650 1854 -4604
rect 1854 -4650 1857 -4604
rect 1805 -4653 1857 -4650
rect 2241 -4790 2293 -4738
rect 2241 -4894 2293 -4842
rect 3537 -5080 3589 -5028
rect 3537 -5184 3589 -5132
rect 6070 -5108 6122 -5056
rect 6174 -5108 6226 -5056
rect 6070 -5212 6122 -5160
rect 6174 -5212 6226 -5160
rect 3105 -5404 3157 -5352
rect 3105 -5508 3157 -5456
rect 2251 -6050 2303 -5998
rect 2251 -6154 2303 -6102
rect 2625 -6050 2677 -5998
rect 2625 -6154 2677 -6102
rect 2945 -6050 2997 -5998
rect 2945 -6154 2997 -6102
rect 8715 -3222 8767 -3219
rect 8715 -3268 8718 -3222
rect 8718 -3268 8764 -3222
rect 8764 -3268 8767 -3222
rect 8715 -3271 8767 -3268
rect 7195 -3500 7247 -3448
rect 7195 -3604 7247 -3552
rect 7355 -3500 7407 -3448
rect 7355 -3604 7407 -3552
rect 7675 -3500 7727 -3448
rect 7675 -3604 7727 -3552
rect 7995 -3500 8047 -3448
rect 7995 -3604 8047 -3552
rect 8315 -3500 8367 -3448
rect 8315 -3604 8367 -3552
rect 8475 -3500 8527 -3448
rect 8475 -3604 8527 -3552
rect 8635 -3500 8687 -3448
rect 8635 -3604 8687 -3552
rect 8794 -3807 8846 -3755
rect 7355 -4036 7407 -3984
rect 7355 -4140 7407 -4088
rect 7515 -4036 7567 -3984
rect 7515 -4140 7567 -4088
rect 7675 -4036 7727 -3984
rect 7675 -4140 7727 -4088
rect 7995 -4036 8047 -3984
rect 7995 -4140 8047 -4088
rect 8315 -4036 8367 -3984
rect 8315 -4140 8367 -4088
rect 8635 -4036 8687 -3984
rect 8635 -4140 8687 -4088
rect 8597 -4343 8649 -4291
rect 7195 -4572 7247 -4520
rect 7195 -4676 7247 -4624
rect 7355 -4572 7407 -4520
rect 7355 -4676 7407 -4624
rect 7675 -4572 7727 -4520
rect 7675 -4676 7727 -4624
rect 7995 -4572 8047 -4520
rect 7995 -4676 8047 -4624
rect 8315 -4572 8367 -4520
rect 8315 -4676 8367 -4624
rect 8475 -4572 8527 -4520
rect 8475 -4676 8527 -4624
rect 8635 -4572 8687 -4520
rect 8635 -4676 8687 -4624
rect 8715 -4828 8767 -4825
rect 8715 -4874 8718 -4828
rect 8718 -4874 8764 -4828
rect 8764 -4874 8767 -4828
rect 8715 -4877 8767 -4874
rect 7355 -5108 7407 -5056
rect 7355 -5212 7407 -5160
rect 7515 -5108 7567 -5056
rect 7515 -5212 7567 -5160
rect 7675 -5108 7727 -5056
rect 7675 -5212 7727 -5160
rect 7995 -5108 8047 -5056
rect 7995 -5212 8047 -5160
rect 8315 -5108 8367 -5056
rect 8315 -5212 8367 -5160
rect 8635 -5108 8687 -5056
rect 8635 -5212 8687 -5160
rect 8794 -5413 8846 -5361
rect 7355 -5636 7407 -5584
rect 7355 -5740 7407 -5688
rect 7675 -5636 7727 -5584
rect 7675 -5740 7727 -5688
rect 7995 -5636 8047 -5584
rect 7995 -5740 8047 -5688
rect 8315 -5636 8367 -5584
rect 8315 -5740 8367 -5688
rect 8475 -5644 8527 -5592
rect 8475 -5748 8527 -5696
rect 8635 -5636 8687 -5584
rect 8635 -5740 8687 -5688
rect 8794 -5928 8846 -5876
rect 3449 -6666 3501 -6614
rect 3449 -6770 3501 -6718
rect 3497 -7436 3549 -7384
rect 3497 -7540 3549 -7488
rect 7355 -6172 7407 -6120
rect 7355 -6276 7407 -6224
rect 7515 -6180 7567 -6128
rect 7515 -6284 7567 -6232
rect 7675 -6172 7727 -6120
rect 7675 -6276 7727 -6224
rect 7995 -6172 8047 -6120
rect 7995 -6276 8047 -6224
rect 8315 -6172 8367 -6120
rect 8315 -6276 8367 -6224
rect 9599 -3140 9651 -3088
rect 9804 -3167 9856 -3115
rect 9908 -3167 9960 -3115
rect 9804 -3271 9856 -3219
rect 9908 -3271 9960 -3219
rect 11165 -3115 11217 -3063
rect 11269 -3115 11321 -3063
rect 17082 -3115 17134 -3063
rect 17186 -3115 17238 -3063
rect 17290 -3115 17342 -3063
rect 11165 -3219 11217 -3167
rect 11269 -3219 11321 -3167
rect 17082 -3219 17134 -3167
rect 17186 -3219 17238 -3167
rect 17290 -3219 17342 -3167
rect 11165 -3323 11217 -3271
rect 11269 -3323 11321 -3271
rect 17082 -3323 17134 -3271
rect 17186 -3323 17238 -3271
rect 17290 -3323 17342 -3271
rect 14212 -3500 14264 -3448
rect 14316 -3500 14368 -3448
rect 14212 -3604 14264 -3552
rect 14316 -3604 14368 -3552
rect 54309 -3625 54365 -3569
rect 54419 -3625 54475 -3569
rect 10070 -3765 10122 -3713
rect 10174 -3765 10226 -3713
rect 16860 -3765 16912 -3713
rect 16964 -3765 17016 -3713
rect 10070 -3869 10122 -3817
rect 10174 -3869 10226 -3817
rect 16860 -3869 16912 -3817
rect 16964 -3869 17016 -3817
rect 8635 -6172 8687 -6120
rect 8635 -6276 8687 -6224
rect 8395 -6482 8398 -6448
rect 8398 -6482 8444 -6448
rect 8444 -6482 8447 -6448
rect 8395 -6500 8447 -6482
rect 6908 -6570 6960 -6518
rect 7012 -6570 7064 -6518
rect 6908 -6674 6960 -6622
rect 7012 -6638 7064 -6622
rect 9839 -6524 9891 -6521
rect 9839 -6570 9842 -6524
rect 9842 -6570 9888 -6524
rect 9888 -6570 9891 -6524
rect 9839 -6573 9891 -6570
rect 9943 -6524 9995 -6521
rect 9943 -6570 9946 -6524
rect 9946 -6570 9992 -6524
rect 9992 -6570 9995 -6524
rect 9943 -6573 9995 -6570
rect 7012 -6674 7037 -6638
rect 7037 -6674 7064 -6638
rect 9839 -6628 9891 -6625
rect 9839 -6674 9842 -6628
rect 9842 -6674 9888 -6628
rect 9888 -6674 9891 -6628
rect 9839 -6677 9891 -6674
rect 9943 -6628 9995 -6625
rect 9943 -6674 9946 -6628
rect 9946 -6674 9992 -6628
rect 9992 -6674 9995 -6628
rect 9943 -6677 9995 -6674
rect 6108 -6809 6160 -6757
rect 6108 -6913 6160 -6861
rect 9263 -6805 9315 -6753
rect 9367 -6805 9419 -6753
rect 9263 -6909 9315 -6857
rect 9367 -6909 9419 -6857
rect 8922 -7205 8974 -7153
rect 9026 -7205 9078 -7153
rect 6038 -7250 6090 -7247
rect 6038 -7296 6041 -7250
rect 6041 -7296 6087 -7250
rect 6087 -7296 6090 -7250
rect 6038 -7299 6090 -7296
rect 6142 -7250 6194 -7247
rect 6142 -7296 6145 -7250
rect 6145 -7296 6191 -7250
rect 6191 -7296 6194 -7250
rect 6142 -7299 6194 -7296
rect 8922 -7275 8974 -7257
rect 8922 -7309 8957 -7275
rect 8957 -7309 8974 -7275
rect 9026 -7275 9078 -7257
rect 9026 -7309 9071 -7275
rect 9071 -7309 9078 -7275
rect 5948 -7438 6000 -7386
rect 5948 -7542 6000 -7490
rect 6380 -7444 6432 -7392
rect 6380 -7548 6432 -7496
rect 10831 -7205 10883 -7153
rect 10935 -7205 10987 -7153
rect 10831 -7309 10883 -7257
rect 10935 -7309 10987 -7257
rect 12626 -6915 12678 -6863
rect 12626 -7019 12678 -6967
rect 12626 -7123 12678 -7071
rect 12726 -7345 12778 -7342
rect 12726 -7391 12729 -7345
rect 12729 -7391 12775 -7345
rect 12775 -7391 12778 -7345
rect 12726 -7394 12778 -7391
rect 12830 -7345 12882 -7342
rect 12830 -7391 12833 -7345
rect 12833 -7391 12879 -7345
rect 12879 -7391 12882 -7345
rect 12830 -7394 12882 -7391
rect 12726 -7449 12778 -7446
rect 12726 -7495 12729 -7449
rect 12729 -7495 12775 -7449
rect 12775 -7495 12778 -7449
rect 12726 -7498 12778 -7495
rect 12830 -7449 12882 -7446
rect 12830 -7495 12833 -7449
rect 12833 -7495 12879 -7449
rect 12879 -7495 12882 -7449
rect 12830 -7498 12882 -7495
rect 13738 -7325 13790 -7322
rect 13738 -7371 13741 -7325
rect 13741 -7371 13787 -7325
rect 13787 -7371 13790 -7325
rect 13738 -7374 13790 -7371
rect 13842 -7325 13894 -7322
rect 13842 -7371 13845 -7325
rect 13845 -7371 13891 -7325
rect 13891 -7371 13894 -7325
rect 13842 -7374 13894 -7371
rect 13946 -7325 13998 -7322
rect 13946 -7371 13949 -7325
rect 13949 -7371 13995 -7325
rect 13995 -7371 13998 -7325
rect 13946 -7374 13998 -7371
rect 14578 -5647 14630 -5595
rect 14578 -5751 14630 -5699
rect 15186 -5647 15238 -5595
rect 15186 -5751 15238 -5699
rect 15794 -5647 15846 -5595
rect 15794 -5751 15846 -5699
rect 15697 -6397 15749 -6394
rect 15697 -6443 15700 -6397
rect 15700 -6443 15746 -6397
rect 15746 -6443 15749 -6397
rect 15697 -6446 15749 -6443
rect 15801 -6397 15853 -6394
rect 15801 -6443 15804 -6397
rect 15804 -6443 15850 -6397
rect 15850 -6443 15853 -6397
rect 15801 -6446 15853 -6443
rect 15905 -6397 15957 -6394
rect 15905 -6443 15908 -6397
rect 15908 -6443 15954 -6397
rect 15954 -6443 15957 -6397
rect 15905 -6446 15957 -6443
rect 15697 -6501 15749 -6498
rect 15697 -6547 15700 -6501
rect 15700 -6547 15746 -6501
rect 15746 -6547 15749 -6501
rect 15697 -6550 15749 -6547
rect 15801 -6501 15853 -6498
rect 15801 -6547 15804 -6501
rect 15804 -6547 15850 -6501
rect 15850 -6547 15853 -6501
rect 15801 -6550 15853 -6547
rect 15905 -6501 15957 -6498
rect 15905 -6547 15908 -6501
rect 15908 -6547 15954 -6501
rect 15954 -6547 15957 -6501
rect 15905 -6550 15957 -6547
rect 15186 -6915 15238 -6863
rect 15186 -7019 15238 -6967
rect 15186 -7123 15238 -7071
rect 20173 -4242 20225 -4239
rect 20173 -4288 20176 -4242
rect 20176 -4288 20222 -4242
rect 20222 -4288 20225 -4242
rect 20173 -4291 20225 -4288
rect 20277 -4242 20329 -4239
rect 20277 -4288 20280 -4242
rect 20280 -4288 20326 -4242
rect 20326 -4288 20329 -4242
rect 20277 -4291 20329 -4288
rect 18626 -6953 18678 -6901
rect 18626 -7057 18678 -7005
rect 18626 -7161 18678 -7109
rect 18946 -6953 18998 -6901
rect 18946 -7057 18998 -7005
rect 18946 -7161 18998 -7109
rect 19266 -6953 19318 -6901
rect 19266 -7057 19318 -7005
rect 19266 -7161 19318 -7109
rect 19586 -6953 19638 -6901
rect 19586 -7057 19638 -7005
rect 19586 -7161 19638 -7109
rect 19906 -6953 19958 -6901
rect 19906 -7057 19958 -7005
rect 19906 -7161 19958 -7109
rect 20226 -6953 20278 -6901
rect 20226 -7057 20278 -7005
rect 20226 -7161 20278 -7109
rect 20546 -6953 20598 -6901
rect 20546 -7057 20598 -7005
rect 20546 -7161 20598 -7109
rect 21186 -4745 21238 -4693
rect 21186 -4849 21238 -4797
rect 21186 -4953 21238 -4901
rect 21157 -7256 21209 -7253
rect 21157 -7302 21160 -7256
rect 21160 -7302 21206 -7256
rect 21206 -7302 21209 -7256
rect 21157 -7305 21209 -7302
rect 21261 -7256 21313 -7253
rect 21261 -7302 21264 -7256
rect 21264 -7302 21310 -7256
rect 21310 -7302 21313 -7256
rect 21261 -7305 21313 -7302
rect 21365 -7256 21417 -7253
rect 21365 -7302 21368 -7256
rect 21368 -7302 21414 -7256
rect 21414 -7302 21417 -7256
rect 21365 -7305 21417 -7302
rect 23644 -4196 23696 -4144
rect 23748 -4196 23800 -4144
rect 23644 -4300 23696 -4248
rect 23748 -4300 23800 -4248
rect 27006 -4904 27058 -4852
rect 27110 -4904 27162 -4852
rect 27006 -5008 27058 -4956
rect 27110 -5008 27162 -4956
rect 27004 -6272 27056 -6220
rect 27108 -6272 27160 -6220
rect 27004 -6376 27056 -6324
rect 27108 -6376 27160 -6324
rect 23644 -7404 23696 -7352
rect 23748 -7404 23800 -7352
rect 23644 -7508 23696 -7456
rect 23748 -7508 23800 -7456
rect 24092 -7404 24144 -7352
rect 24196 -7404 24248 -7352
rect 24092 -7508 24144 -7456
rect 24196 -7508 24248 -7456
rect 29814 -4116 29866 -4064
rect 29918 -4116 29970 -4064
rect 30022 -4116 30074 -4064
rect 30126 -4116 30178 -4064
rect 30230 -4116 30282 -4064
rect 29814 -4220 29866 -4168
rect 29918 -4220 29970 -4168
rect 30022 -4220 30074 -4168
rect 30126 -4220 30178 -4168
rect 30230 -4220 30282 -4168
rect 29814 -4324 29866 -4272
rect 29918 -4324 29970 -4272
rect 30022 -4324 30074 -4272
rect 30126 -4324 30178 -4272
rect 30230 -4324 30282 -4272
rect 29814 -5072 29866 -5020
rect 29918 -5072 29970 -5020
rect 30022 -5072 30074 -5020
rect 30126 -5072 30178 -5020
rect 30230 -5072 30282 -5020
rect 29814 -5176 29866 -5124
rect 29918 -5176 29970 -5124
rect 30022 -5176 30074 -5124
rect 30126 -5176 30178 -5124
rect 30230 -5176 30282 -5124
rect 29814 -5280 29866 -5228
rect 29918 -5280 29970 -5228
rect 30022 -5280 30074 -5228
rect 30126 -5280 30178 -5228
rect 30230 -5280 30282 -5228
rect 29814 -5384 29866 -5332
rect 29918 -5384 29970 -5332
rect 30022 -5384 30074 -5332
rect 30126 -5384 30178 -5332
rect 30230 -5384 30282 -5332
rect 29814 -5488 29866 -5436
rect 29918 -5488 29970 -5436
rect 30022 -5488 30074 -5436
rect 30126 -5488 30178 -5436
rect 30230 -5488 30282 -5436
rect 54544 -4500 54600 -4444
rect 54654 -4500 54710 -4444
rect 54817 -5537 54873 -5481
rect 54927 -5537 54983 -5481
rect 29254 -6128 29306 -6076
rect 29358 -6128 29410 -6076
rect 29462 -6128 29514 -6076
rect 29566 -6128 29618 -6076
rect 29670 -6128 29722 -6076
rect 29254 -6232 29306 -6180
rect 29358 -6232 29410 -6180
rect 29462 -6232 29514 -6180
rect 29566 -6232 29618 -6180
rect 29670 -6232 29722 -6180
rect 29254 -6336 29306 -6284
rect 29358 -6336 29410 -6284
rect 29462 -6336 29514 -6284
rect 29566 -6336 29618 -6284
rect 29670 -6336 29722 -6284
rect 29814 -7084 29866 -7032
rect 29918 -7084 29970 -7032
rect 30022 -7084 30074 -7032
rect 30126 -7084 30178 -7032
rect 30230 -7084 30282 -7032
rect 29814 -7188 29866 -7136
rect 29918 -7188 29970 -7136
rect 30022 -7188 30074 -7136
rect 30126 -7188 30178 -7136
rect 30230 -7188 30282 -7136
rect 29814 -7292 29866 -7240
rect 29918 -7292 29970 -7240
rect 30022 -7292 30074 -7240
rect 30126 -7292 30178 -7240
rect 30230 -7292 30282 -7240
rect 29814 -7396 29866 -7344
rect 29918 -7396 29970 -7344
rect 30022 -7396 30074 -7344
rect 30126 -7396 30178 -7344
rect 30230 -7396 30282 -7344
rect 29814 -7500 29866 -7448
rect 29918 -7500 29970 -7448
rect 30022 -7500 30074 -7448
rect 30126 -7500 30178 -7448
rect 30230 -7500 30282 -7448
rect 55066 -6411 55122 -6355
rect 55176 -6411 55232 -6355
rect 55315 -7460 55371 -7404
rect 55425 -7460 55481 -7404
rect 11544 -8082 11596 -8030
rect 11648 -8082 11700 -8030
rect 11544 -8186 11596 -8134
rect 11648 -8186 11700 -8134
rect 44548 -8008 44600 -7956
rect 44652 -8008 44704 -7956
rect 44756 -8008 44808 -7956
rect 44860 -8008 44912 -7956
rect 44964 -8008 45016 -7956
rect 48988 -8008 49040 -7956
rect 49092 -8008 49144 -7956
rect 49196 -8008 49248 -7956
rect 49300 -8008 49352 -7956
rect 49404 -8008 49456 -7956
rect 34718 -8108 34770 -8056
rect 34822 -8108 34874 -8056
rect 34926 -8108 34978 -8056
rect 35030 -8108 35082 -8056
rect 35134 -8108 35186 -8056
rect 39158 -8108 39210 -8056
rect 39262 -8108 39314 -8056
rect 39366 -8108 39418 -8056
rect 39470 -8108 39522 -8056
rect 39574 -8108 39626 -8056
rect 34718 -8212 34770 -8160
rect 34822 -8212 34874 -8160
rect 34926 -8212 34978 -8160
rect 35030 -8212 35082 -8160
rect 35134 -8212 35186 -8160
rect 39158 -8212 39210 -8160
rect 39262 -8212 39314 -8160
rect 39366 -8212 39418 -8160
rect 39470 -8212 39522 -8160
rect 39574 -8212 39626 -8160
rect 15082 -8937 15134 -8885
rect 15186 -8937 15238 -8885
rect 15290 -8937 15342 -8885
rect 15082 -9041 15134 -8989
rect 15186 -9041 15238 -8989
rect 15290 -9041 15342 -8989
rect 15082 -9145 15134 -9093
rect 15186 -9145 15238 -9093
rect 15290 -9145 15342 -9093
rect 21157 -8437 21209 -8385
rect 21261 -8437 21313 -8385
rect 21365 -8437 21417 -8385
rect 21157 -8541 21209 -8489
rect 21261 -8541 21313 -8489
rect 21365 -8541 21417 -8489
rect 21157 -8645 21209 -8593
rect 21261 -8645 21313 -8593
rect 21365 -8645 21417 -8593
rect 34718 -8316 34770 -8264
rect 34822 -8316 34874 -8264
rect 34926 -8316 34978 -8264
rect 35030 -8316 35082 -8264
rect 35134 -8316 35186 -8264
rect 39158 -8316 39210 -8264
rect 39262 -8316 39314 -8264
rect 39366 -8316 39418 -8264
rect 39470 -8316 39522 -8264
rect 39574 -8316 39626 -8264
rect 34718 -8420 34770 -8368
rect 34822 -8420 34874 -8368
rect 34926 -8420 34978 -8368
rect 35030 -8420 35082 -8368
rect 35134 -8420 35186 -8368
rect 39158 -8420 39210 -8368
rect 39262 -8420 39314 -8368
rect 39366 -8420 39418 -8368
rect 39470 -8420 39522 -8368
rect 39574 -8420 39626 -8368
rect 44548 -8112 44600 -8060
rect 44652 -8112 44704 -8060
rect 44756 -8112 44808 -8060
rect 44860 -8112 44912 -8060
rect 44964 -8112 45016 -8060
rect 48988 -8112 49040 -8060
rect 49092 -8112 49144 -8060
rect 49196 -8112 49248 -8060
rect 49300 -8112 49352 -8060
rect 49404 -8112 49456 -8060
rect 44548 -8216 44600 -8164
rect 44652 -8216 44704 -8164
rect 44756 -8216 44808 -8164
rect 44860 -8216 44912 -8164
rect 44964 -8216 45016 -8164
rect 48988 -8216 49040 -8164
rect 49092 -8216 49144 -8164
rect 49196 -8216 49248 -8164
rect 49300 -8216 49352 -8164
rect 49404 -8216 49456 -8164
rect 44548 -8320 44600 -8268
rect 44652 -8320 44704 -8268
rect 44756 -8320 44808 -8268
rect 44860 -8320 44912 -8268
rect 44964 -8320 45016 -8268
rect 48988 -8320 49040 -8268
rect 49092 -8320 49144 -8268
rect 49196 -8320 49248 -8268
rect 49300 -8320 49352 -8268
rect 49404 -8320 49456 -8268
rect 44548 -8424 44600 -8372
rect 44652 -8424 44704 -8372
rect 44756 -8424 44808 -8372
rect 44860 -8424 44912 -8372
rect 44964 -8424 45016 -8372
rect 48988 -8424 49040 -8372
rect 49092 -8424 49144 -8372
rect 49196 -8424 49248 -8372
rect 49300 -8424 49352 -8372
rect 49404 -8424 49456 -8372
rect 34718 -8524 34770 -8472
rect 34822 -8524 34874 -8472
rect 34926 -8524 34978 -8472
rect 35030 -8524 35082 -8472
rect 35134 -8524 35186 -8472
rect 39158 -8524 39210 -8472
rect 39262 -8524 39314 -8472
rect 39366 -8524 39418 -8472
rect 39470 -8524 39522 -8472
rect 39574 -8524 39626 -8472
rect 55661 -8798 55717 -8742
rect 55771 -8798 55827 -8742
rect 8467 -12343 8523 -12287
rect 8577 -12343 8633 -12287
rect 10460 -12343 10516 -12287
rect 10570 -12343 10626 -12287
rect 12489 -12343 12545 -12287
rect 12599 -12343 12655 -12287
rect 6882 -12419 6938 -12363
rect 6992 -12419 7048 -12363
rect 8883 -12416 8939 -12360
rect 8993 -12416 9049 -12360
rect 14492 -12343 14548 -12287
rect 14602 -12343 14658 -12287
rect 10908 -12419 10964 -12363
rect 11018 -12419 11074 -12363
rect 16507 -12344 16563 -12288
rect 16617 -12344 16673 -12288
rect 12917 -12418 12973 -12362
rect 13027 -12418 13083 -12362
rect 18528 -12343 18584 -12287
rect 18638 -12343 18694 -12287
rect 14887 -12418 14943 -12362
rect 14997 -12418 15053 -12362
rect 16922 -12414 16978 -12358
rect 17032 -12414 17088 -12358
rect 25467 -12343 25523 -12287
rect 25577 -12343 25633 -12287
rect 27460 -12343 27516 -12287
rect 27570 -12343 27626 -12287
rect 29489 -12343 29545 -12287
rect 29599 -12343 29655 -12287
rect 23882 -12419 23938 -12363
rect 23992 -12419 24048 -12363
rect 25883 -12416 25939 -12360
rect 25993 -12416 26049 -12360
rect 31492 -12343 31548 -12287
rect 31602 -12343 31658 -12287
rect 27908 -12419 27964 -12363
rect 28018 -12419 28074 -12363
rect 33507 -12344 33563 -12288
rect 33617 -12344 33673 -12288
rect 29917 -12418 29973 -12362
rect 30027 -12418 30083 -12362
rect 35528 -12343 35584 -12287
rect 35638 -12343 35694 -12287
rect 31887 -12418 31943 -12362
rect 31997 -12418 32053 -12362
rect 33922 -12414 33978 -12358
rect 34032 -12414 34088 -12358
rect 35900 -12370 35956 -12314
rect 36010 -12370 36066 -12314
rect 18977 -16257 19033 -16201
rect 19087 -16257 19143 -16201
rect 19197 -16257 19253 -16201
rect 18977 -16367 19033 -16311
rect 19087 -16367 19143 -16311
rect 19197 -16367 19253 -16311
rect 18977 -16477 19033 -16421
rect 19087 -16477 19143 -16421
rect 19197 -16477 19253 -16421
rect 39211 -16194 39267 -16138
rect 39321 -16194 39377 -16138
rect 39431 -16194 39487 -16138
rect 39211 -16304 39267 -16248
rect 39321 -16304 39377 -16248
rect 39431 -16304 39487 -16248
rect 39211 -16414 39267 -16358
rect 39321 -16414 39377 -16358
rect 39431 -16414 39487 -16358
<< metal2 >>
rect 30732 6548 31016 6560
rect 30732 6496 30744 6548
rect 30796 6496 30848 6548
rect 30900 6496 30952 6548
rect 31004 6496 31016 6548
rect 30732 6444 31016 6496
rect 30732 6392 30744 6444
rect 30796 6392 30848 6444
rect 30900 6392 30952 6444
rect 31004 6392 31016 6444
rect 30732 6340 31016 6392
rect 30732 6288 30744 6340
rect 30796 6288 30848 6340
rect 30900 6288 30952 6340
rect 31004 6288 31016 6340
rect -1790 5190 -1465 5201
rect -1790 5134 -1781 5190
rect -1725 5134 -1671 5190
rect -1615 5134 -1561 5190
rect -1505 5134 -1465 5190
rect -1790 5080 -1465 5134
rect -1790 5024 -1781 5080
rect -1725 5024 -1671 5080
rect -1615 5024 -1561 5080
rect -1505 5024 -1465 5080
rect -1790 -10864 -1465 5024
rect 2675 5171 2855 5181
rect 2675 5115 2685 5171
rect 2741 5115 2789 5171
rect 2845 5115 2855 5171
rect 2675 5067 2855 5115
rect 2675 5011 2685 5067
rect 2741 5011 2789 5067
rect 2845 5011 2855 5067
rect 2675 5001 2855 5011
rect 3464 5171 3540 5181
rect 3464 5115 3474 5171
rect 3530 5115 3540 5171
rect 3464 5067 3540 5115
rect 3464 5011 3474 5067
rect 3530 5011 3540 5067
rect 3464 5001 3540 5011
rect 5245 5117 5425 5127
rect 5245 5061 5255 5117
rect 5311 5061 5359 5117
rect 5415 5061 5425 5117
rect 5245 5013 5425 5061
rect 2034 4822 2214 4832
rect 2034 4766 2044 4822
rect 2100 4766 2148 4822
rect 2204 4766 2214 4822
rect 2034 4718 2214 4766
rect 2034 4662 2044 4718
rect 2100 4662 2148 4718
rect 2204 4662 2214 4718
rect 2034 4652 2214 4662
rect -1115 4032 -790 4045
rect -1115 3976 -1106 4032
rect -1050 3976 -996 4032
rect -940 3976 -886 4032
rect -830 3976 -790 4032
rect -1115 3922 -790 3976
rect -1115 3866 -1106 3922
rect -1050 3866 -996 3922
rect -940 3866 -886 3922
rect -830 3910 -790 3922
rect -830 3866 -789 3910
rect -1115 3853 -789 3866
rect -1790 -11017 -1314 -10864
rect -1790 -11018 -1524 -11017
rect -1790 -11074 -1761 -11018
rect -1705 -11074 -1651 -11018
rect -1595 -11073 -1524 -11018
rect -1468 -11073 -1414 -11017
rect -1358 -11073 -1314 -11017
rect -1595 -11074 -1314 -11073
rect -1790 -11127 -1314 -11074
rect -1790 -11128 -1524 -11127
rect -1790 -11184 -1761 -11128
rect -1705 -11184 -1651 -11128
rect -1595 -11183 -1524 -11128
rect -1468 -11183 -1414 -11127
rect -1358 -11183 -1314 -11127
rect -1595 -11184 -1314 -11183
rect -1790 -11188 -1314 -11184
rect -1790 -11189 -1465 -11188
rect -1115 -11433 -790 3853
rect 2044 3702 2204 4652
rect 2395 4043 2575 4053
rect 2395 3987 2405 4043
rect 2461 3987 2509 4043
rect 2565 3987 2575 4043
rect 2395 3939 2575 3987
rect 2395 3883 2405 3939
rect 2461 3883 2509 3939
rect 2565 3883 2575 3939
rect 2395 3873 2575 3883
rect 2034 3692 2214 3702
rect 2034 3636 2044 3692
rect 2100 3636 2148 3692
rect 2204 3636 2214 3692
rect 2034 3588 2214 3636
rect 2034 3532 2044 3588
rect 2100 3532 2148 3588
rect 2204 3532 2214 3588
rect 2034 3522 2214 3532
rect 2044 1178 2204 3522
rect 2034 1168 2214 1178
rect 2034 1112 2044 1168
rect 2100 1112 2148 1168
rect 2204 1112 2214 1168
rect 2034 1064 2214 1112
rect 2034 1008 2044 1064
rect 2100 1008 2148 1064
rect 2204 1008 2214 1064
rect 2034 998 2214 1008
rect 2405 665 2565 3873
rect 2685 2923 2845 5001
rect 5245 4957 5255 5013
rect 5311 4957 5359 5013
rect 5415 4957 5425 5013
rect 5245 4947 5425 4957
rect 6249 5117 6325 5127
rect 6249 5061 6259 5117
rect 6315 5061 6325 5117
rect 6249 5013 6325 5061
rect 6249 4957 6259 5013
rect 6315 4957 6325 5013
rect 6249 4947 6325 4957
rect 6889 5117 6965 5127
rect 6889 5061 6899 5117
rect 6955 5061 6965 5117
rect 6889 5013 6965 5061
rect 6889 4957 6899 5013
rect 6955 4957 6965 5013
rect 6889 4947 6965 4957
rect 7529 5117 7605 5127
rect 7529 5061 7539 5117
rect 7595 5061 7605 5117
rect 7529 5013 7605 5061
rect 7529 4957 7539 5013
rect 7595 4957 7605 5013
rect 7529 4947 7605 4957
rect 3544 4822 3620 4832
rect 3544 4766 3554 4822
rect 3610 4766 3620 4822
rect 3544 4718 3620 4766
rect 3544 4662 3554 4718
rect 3610 4662 3620 4718
rect 3544 4652 3620 4662
rect 3704 4822 3780 4832
rect 3704 4766 3714 4822
rect 3770 4766 3780 4822
rect 3704 4718 3780 4766
rect 3704 4662 3714 4718
rect 3770 4662 3780 4718
rect 3704 4652 3780 4662
rect 4345 4822 4421 4832
rect 4345 4766 4355 4822
rect 4411 4766 4421 4822
rect 4345 4718 4421 4766
rect 4345 4662 4355 4718
rect 4411 4662 4421 4718
rect 4345 4652 4421 4662
rect 5255 4336 5415 4947
rect 5517 4822 5697 4832
rect 5517 4766 5527 4822
rect 5583 4766 5631 4822
rect 5687 4766 5697 4822
rect 5517 4718 5697 4766
rect 5517 4662 5527 4718
rect 5583 4662 5631 4718
rect 5687 4662 5697 4718
rect 5517 4652 5697 4662
rect 6569 4822 6645 4832
rect 6569 4766 6579 4822
rect 6635 4766 6645 4822
rect 6569 4718 6645 4766
rect 6569 4662 6579 4718
rect 6635 4662 6645 4718
rect 6569 4652 6645 4662
rect 7209 4822 7285 4832
rect 7209 4766 7219 4822
rect 7275 4766 7285 4822
rect 7209 4718 7285 4766
rect 7209 4662 7219 4718
rect 7275 4662 7285 4718
rect 7209 4652 7285 4662
rect 3384 4326 3460 4336
rect 3384 4270 3394 4326
rect 3450 4270 3460 4326
rect 3384 4222 3460 4270
rect 3384 4166 3394 4222
rect 3450 4166 3460 4222
rect 3384 4156 3460 4166
rect 4024 4326 4100 4336
rect 4024 4270 4034 4326
rect 4090 4270 4100 4326
rect 4024 4222 4100 4270
rect 4024 4166 4034 4222
rect 4090 4166 4100 4222
rect 4024 4156 4100 4166
rect 4664 4326 4740 4336
rect 4664 4270 4674 4326
rect 4730 4270 4740 4326
rect 4664 4222 4740 4270
rect 4664 4166 4674 4222
rect 4730 4166 4740 4222
rect 4664 4156 4740 4166
rect 5245 4326 5425 4336
rect 5245 4270 5255 4326
rect 5311 4270 5359 4326
rect 5415 4270 5425 4326
rect 5245 4222 5425 4270
rect 5245 4166 5255 4222
rect 5311 4166 5359 4222
rect 5415 4166 5425 4222
rect 5245 4118 5425 4166
rect 5245 4062 5255 4118
rect 5311 4062 5359 4118
rect 5415 4062 5425 4118
rect 3464 4043 3540 4053
rect 5245 4052 5425 4062
rect 3464 3987 3474 4043
rect 3530 3987 3540 4043
rect 3464 3939 3540 3987
rect 3464 3883 3474 3939
rect 3530 3883 3540 3939
rect 3464 3873 3540 3883
rect 5255 3702 5415 4052
rect 5527 3853 5687 4652
rect 11153 4302 11333 4312
rect 11153 4246 11163 4302
rect 11219 4246 11267 4302
rect 11323 4246 11333 4302
rect 6569 4222 6645 4232
rect 6569 4166 6579 4222
rect 6635 4166 6645 4222
rect 6569 4118 6645 4166
rect 6569 4062 6579 4118
rect 6635 4062 6645 4118
rect 6569 4052 6645 4062
rect 7209 4222 7285 4232
rect 7209 4166 7219 4222
rect 7275 4166 7285 4222
rect 7209 4118 7285 4166
rect 11153 4198 11333 4246
rect 11153 4142 11163 4198
rect 11219 4142 11267 4198
rect 11323 4142 11333 4198
rect 11153 4132 11333 4142
rect 17155 4250 17230 4260
rect 17155 4194 17165 4250
rect 17221 4194 17230 4250
rect 7209 4062 7219 4118
rect 7275 4062 7285 4118
rect 7209 4052 7285 4062
rect 5517 3843 5697 3853
rect 5517 3787 5527 3843
rect 5583 3787 5631 3843
rect 5687 3787 5697 3843
rect 5517 3739 5697 3787
rect 3544 3692 3620 3702
rect 3544 3636 3554 3692
rect 3610 3636 3620 3692
rect 3544 3588 3620 3636
rect 3544 3532 3554 3588
rect 3610 3532 3620 3588
rect 3544 3522 3620 3532
rect 3704 3692 3780 3702
rect 3704 3636 3714 3692
rect 3770 3636 3780 3692
rect 3704 3588 3780 3636
rect 3704 3532 3714 3588
rect 3770 3532 3780 3588
rect 3704 3522 3780 3532
rect 4345 3692 4421 3702
rect 4345 3636 4355 3692
rect 4411 3636 4421 3692
rect 4345 3588 4421 3636
rect 4345 3532 4355 3588
rect 4411 3532 4421 3588
rect 4345 3522 4421 3532
rect 5245 3692 5425 3702
rect 5245 3636 5255 3692
rect 5311 3636 5359 3692
rect 5415 3636 5425 3692
rect 5517 3683 5527 3739
rect 5583 3683 5631 3739
rect 5687 3683 5697 3739
rect 5517 3673 5697 3683
rect 6249 3843 6325 3853
rect 6249 3787 6259 3843
rect 6315 3787 6325 3843
rect 6249 3739 6325 3787
rect 6249 3683 6259 3739
rect 6315 3683 6325 3739
rect 6249 3673 6325 3683
rect 6889 3843 6965 3853
rect 6889 3787 6899 3843
rect 6955 3787 6965 3843
rect 6889 3739 6965 3787
rect 6889 3683 6899 3739
rect 6955 3683 6965 3739
rect 6889 3673 6965 3683
rect 7529 3843 7605 3853
rect 7529 3787 7539 3843
rect 7595 3787 7605 3843
rect 7529 3739 7605 3787
rect 7529 3683 7539 3739
rect 7595 3683 7605 3739
rect 7529 3673 7605 3683
rect 5245 3588 5425 3636
rect 5245 3532 5255 3588
rect 5311 3532 5359 3588
rect 5415 3532 5425 3588
rect 5245 3522 5425 3532
rect 3384 3300 3460 3310
rect 3384 3244 3394 3300
rect 3450 3244 3460 3300
rect 3384 3196 3460 3244
rect 3384 3140 3394 3196
rect 3450 3140 3460 3196
rect 3384 3130 3460 3140
rect 4024 3300 4100 3310
rect 4024 3244 4034 3300
rect 4090 3244 4100 3300
rect 4024 3196 4100 3244
rect 4024 3140 4034 3196
rect 4090 3140 4100 3196
rect 4024 3130 4100 3140
rect 4664 3300 4740 3310
rect 4664 3244 4674 3300
rect 4730 3244 4740 3300
rect 4664 3196 4740 3244
rect 4664 3140 4674 3196
rect 4730 3140 4740 3196
rect 4664 3130 4740 3140
rect 5255 2991 5415 3522
rect 5527 3310 5687 3673
rect 10885 3336 11065 3346
rect 5517 3300 5697 3310
rect 5517 3244 5527 3300
rect 5583 3244 5631 3300
rect 5687 3244 5697 3300
rect 5517 3196 5697 3244
rect 5517 3140 5527 3196
rect 5583 3140 5631 3196
rect 5687 3140 5697 3196
rect 5517 3130 5697 3140
rect 6569 3300 6645 3310
rect 6569 3244 6579 3300
rect 6635 3244 6645 3300
rect 6569 3196 6645 3244
rect 6569 3140 6579 3196
rect 6635 3140 6645 3196
rect 6569 3130 6645 3140
rect 7209 3300 7285 3310
rect 7209 3244 7219 3300
rect 7275 3244 7285 3300
rect 7209 3196 7285 3244
rect 7209 3140 7219 3196
rect 7275 3140 7285 3196
rect 10885 3280 10895 3336
rect 10951 3280 10999 3336
rect 11055 3280 11065 3336
rect 10885 3232 11065 3280
rect 10885 3176 10895 3232
rect 10951 3176 10999 3232
rect 11055 3176 11065 3232
rect 10885 3166 11065 3176
rect 7209 3130 7285 3140
rect 5245 2981 5425 2991
rect 5245 2925 5255 2981
rect 5311 2925 5359 2981
rect 5415 2925 5425 2981
rect 2675 2913 2855 2923
rect 2675 2857 2685 2913
rect 2741 2857 2789 2913
rect 2845 2857 2855 2913
rect 2675 2809 2855 2857
rect 2675 2753 2685 2809
rect 2741 2753 2789 2809
rect 2845 2753 2855 2809
rect 2675 2743 2855 2753
rect 3464 2913 3540 2923
rect 3464 2857 3474 2913
rect 3530 2857 3540 2913
rect 3464 2809 3540 2857
rect 5245 2877 5425 2925
rect 5245 2821 5255 2877
rect 5311 2821 5359 2877
rect 5415 2821 5425 2877
rect 5245 2811 5425 2821
rect 3464 2753 3474 2809
rect 3530 2753 3540 2809
rect 3464 2743 3540 2753
rect 2395 655 2575 665
rect 2395 599 2405 655
rect 2461 599 2509 655
rect 2565 599 2575 655
rect 2395 551 2575 599
rect 2395 495 2405 551
rect 2461 495 2509 551
rect 2565 495 2575 551
rect 2395 485 2575 495
rect 2138 302 2214 312
rect 2138 246 2148 302
rect 2204 246 2214 302
rect 2138 198 2214 246
rect 2138 142 2148 198
rect 2204 142 2214 198
rect 2138 132 2214 142
rect 2138 -1028 2214 -1018
rect 2138 -1084 2148 -1028
rect 2204 -1084 2214 -1028
rect 2138 -1132 2214 -1084
rect 2138 -1188 2148 -1132
rect 2204 -1188 2214 -1132
rect 2138 -1198 2214 -1188
rect -260 -1572 -80 -1562
rect -260 -1628 -250 -1572
rect -194 -1628 -146 -1572
rect -90 -1628 -80 -1572
rect -260 -1676 -80 -1628
rect -260 -1732 -250 -1676
rect -194 -1732 -146 -1676
rect -90 -1732 -80 -1676
rect -260 -1742 -80 -1732
rect 741 -1572 921 -1562
rect 741 -1628 751 -1572
rect 807 -1628 855 -1572
rect 911 -1628 921 -1572
rect 741 -1676 921 -1628
rect 2405 -1653 2565 485
rect 2685 -465 2845 2743
rect 3704 2562 3780 2572
rect 3704 2506 3714 2562
rect 3770 2506 3780 2562
rect 3704 2458 3780 2506
rect 3704 2402 3714 2458
rect 3770 2402 3780 2458
rect 3704 2392 3780 2402
rect 4345 2562 4421 2572
rect 4345 2506 4355 2562
rect 4411 2506 4421 2562
rect 4345 2458 4421 2506
rect 4345 2402 4355 2458
rect 4411 2402 4421 2458
rect 4345 2392 4421 2402
rect 5255 2180 5415 2811
rect 5527 2572 5687 3130
rect 6249 2981 6325 2991
rect 6249 2925 6259 2981
rect 6315 2925 6325 2981
rect 6249 2877 6325 2925
rect 6249 2821 6259 2877
rect 6315 2821 6325 2877
rect 6249 2811 6325 2821
rect 6889 2981 6965 2991
rect 6889 2925 6899 2981
rect 6955 2925 6965 2981
rect 6889 2877 6965 2925
rect 6889 2821 6899 2877
rect 6955 2821 6965 2877
rect 6889 2811 6965 2821
rect 7529 2981 7605 2991
rect 7529 2925 7539 2981
rect 7595 2925 7605 2981
rect 7529 2877 7605 2925
rect 7529 2821 7539 2877
rect 7595 2821 7605 2877
rect 7529 2811 7605 2821
rect 5517 2562 5697 2572
rect 5517 2506 5527 2562
rect 5583 2506 5631 2562
rect 5687 2506 5697 2562
rect 5517 2458 5697 2506
rect 5517 2402 5527 2458
rect 5583 2402 5631 2458
rect 5687 2402 5697 2458
rect 5517 2354 5697 2402
rect 5517 2298 5527 2354
rect 5583 2298 5631 2354
rect 5687 2298 5697 2354
rect 5517 2288 5697 2298
rect 6249 2458 6325 2468
rect 6249 2402 6259 2458
rect 6315 2402 6325 2458
rect 6249 2354 6325 2402
rect 6249 2298 6259 2354
rect 6315 2298 6325 2354
rect 6249 2288 6325 2298
rect 6889 2458 6965 2468
rect 6889 2402 6899 2458
rect 6955 2402 6965 2458
rect 6889 2354 6965 2402
rect 6889 2298 6899 2354
rect 6955 2298 6965 2354
rect 6889 2288 6965 2298
rect 7529 2458 7605 2468
rect 7529 2402 7539 2458
rect 7595 2402 7605 2458
rect 7529 2354 7605 2402
rect 7529 2298 7539 2354
rect 7595 2298 7605 2354
rect 7529 2288 7605 2298
rect 5245 2170 5425 2180
rect 5245 2114 5255 2170
rect 5311 2114 5359 2170
rect 5415 2114 5425 2170
rect 3384 2066 3460 2076
rect 3384 2010 3394 2066
rect 3450 2010 3460 2066
rect 3384 1962 3460 2010
rect 3384 1906 3394 1962
rect 3450 1906 3460 1962
rect 3384 1896 3460 1906
rect 4024 2066 4100 2076
rect 4024 2010 4034 2066
rect 4090 2010 4100 2066
rect 4024 1962 4100 2010
rect 4024 1906 4034 1962
rect 4090 1906 4100 1962
rect 4024 1896 4100 1906
rect 4664 2066 4740 2076
rect 4664 2010 4674 2066
rect 4730 2010 4740 2066
rect 4664 1962 4740 2010
rect 4664 1906 4674 1962
rect 4730 1906 4740 1962
rect 4664 1896 4740 1906
rect 5245 2066 5425 2114
rect 5245 2010 5255 2066
rect 5311 2010 5359 2066
rect 5415 2010 5425 2066
rect 5245 1962 5425 2010
rect 5245 1906 5255 1962
rect 5311 1906 5359 1962
rect 5415 1906 5425 1962
rect 5245 1896 5425 1906
rect 5255 1649 5415 1896
rect 5245 1639 5425 1649
rect 5245 1583 5255 1639
rect 5311 1583 5359 1639
rect 5415 1583 5425 1639
rect 5245 1535 5425 1583
rect 5245 1479 5255 1535
rect 5311 1479 5359 1535
rect 5415 1479 5425 1535
rect 5245 1469 5425 1479
rect 3544 1168 3620 1178
rect 3544 1112 3554 1168
rect 3610 1112 3620 1168
rect 3544 1064 3620 1112
rect 3544 1008 3554 1064
rect 3610 1008 3620 1064
rect 3544 998 3620 1008
rect 3464 655 3540 665
rect 3464 599 3474 655
rect 3530 599 3540 655
rect 3464 551 3540 599
rect 3464 495 3474 551
rect 3530 495 3540 551
rect 3464 483 3540 495
rect 5255 416 5415 1469
rect 5527 1278 5687 2288
rect 10895 2228 11055 3166
rect 10885 2218 11065 2228
rect 6569 2170 6645 2180
rect 6569 2114 6579 2170
rect 6635 2114 6645 2170
rect 6569 2066 6645 2114
rect 6569 2010 6579 2066
rect 6635 2010 6645 2066
rect 6569 2000 6645 2010
rect 7209 2170 7285 2180
rect 7209 2114 7219 2170
rect 7275 2114 7285 2170
rect 7209 2066 7285 2114
rect 7209 2010 7219 2066
rect 7275 2010 7285 2066
rect 10885 2162 10895 2218
rect 10951 2162 10999 2218
rect 11055 2162 11065 2218
rect 10885 2114 11065 2162
rect 10885 2058 10895 2114
rect 10951 2058 10999 2114
rect 11055 2058 11065 2114
rect 10885 2048 11065 2058
rect 7209 2000 7285 2010
rect 8484 1639 8560 1649
rect 8484 1583 8494 1639
rect 8550 1583 8560 1639
rect 8484 1535 8560 1583
rect 8484 1479 8494 1535
rect 8550 1479 8560 1535
rect 8484 1469 8560 1479
rect 9380 1639 9456 1649
rect 9380 1583 9390 1639
rect 9446 1583 9456 1639
rect 9380 1535 9456 1583
rect 9380 1479 9390 1535
rect 9446 1479 9456 1535
rect 9380 1469 9456 1479
rect 10276 1639 10352 1649
rect 10276 1583 10286 1639
rect 10342 1583 10352 1639
rect 10276 1535 10352 1583
rect 10276 1479 10286 1535
rect 10342 1479 10352 1535
rect 10276 1469 10352 1479
rect 5517 1268 5697 1278
rect 5517 1212 5527 1268
rect 5583 1212 5631 1268
rect 5687 1212 5697 1268
rect 5517 1164 5697 1212
rect 5517 1108 5527 1164
rect 5583 1108 5631 1164
rect 5687 1108 5697 1164
rect 5517 1098 5697 1108
rect 8932 1268 9008 1278
rect 8932 1212 8942 1268
rect 8998 1212 9008 1268
rect 8932 1164 9008 1212
rect 8932 1108 8942 1164
rect 8998 1108 9008 1164
rect 8932 1098 9008 1108
rect 9828 1268 9904 1278
rect 9828 1212 9838 1268
rect 9894 1212 9904 1268
rect 9828 1164 9904 1212
rect 9828 1108 9838 1164
rect 9894 1108 9904 1164
rect 9828 1098 9904 1108
rect 10116 1268 10192 1278
rect 10116 1212 10126 1268
rect 10182 1212 10192 1268
rect 10116 1164 10192 1212
rect 10116 1108 10126 1164
rect 10182 1108 10192 1164
rect 10116 1098 10192 1108
rect 5527 817 5687 1098
rect 5517 807 5697 817
rect 5517 751 5527 807
rect 5583 751 5631 807
rect 5687 751 5697 807
rect 5517 703 5697 751
rect 5517 647 5527 703
rect 5583 647 5631 703
rect 5687 647 5697 703
rect 5517 637 5697 647
rect 6569 807 6645 817
rect 6569 751 6579 807
rect 6635 751 6645 807
rect 6569 703 6645 751
rect 6569 647 6579 703
rect 6635 647 6645 703
rect 6569 637 6645 647
rect 7209 807 7285 817
rect 7209 751 7219 807
rect 7275 751 7285 807
rect 7209 703 7285 751
rect 7209 647 7219 703
rect 7275 647 7285 703
rect 7209 637 7285 647
rect 5245 406 5425 416
rect 5245 350 5255 406
rect 5311 350 5359 406
rect 5415 350 5425 406
rect 3544 302 3620 312
rect 3544 246 3554 302
rect 3610 246 3620 302
rect 3544 198 3620 246
rect 3544 142 3554 198
rect 3610 142 3620 198
rect 3544 132 3620 142
rect 3704 302 3780 312
rect 3704 246 3714 302
rect 3770 246 3780 302
rect 3704 198 3780 246
rect 3704 142 3714 198
rect 3770 142 3780 198
rect 3704 132 3780 142
rect 4345 302 4421 312
rect 4345 246 4355 302
rect 4411 246 4421 302
rect 4345 198 4421 246
rect 4345 142 4355 198
rect 4411 142 4421 198
rect 4345 132 4421 142
rect 5245 302 5425 350
rect 5245 246 5255 302
rect 5311 246 5359 302
rect 5415 246 5425 302
rect 5245 198 5425 246
rect 5245 142 5255 198
rect 5311 142 5359 198
rect 5415 142 5425 198
rect 5245 132 5425 142
rect 3384 -194 3460 -184
rect 3384 -250 3394 -194
rect 3450 -250 3460 -194
rect 3384 -298 3460 -250
rect 3384 -354 3394 -298
rect 3450 -354 3460 -298
rect 3384 -364 3460 -354
rect 4024 -194 4100 -184
rect 4024 -250 4034 -194
rect 4090 -250 4100 -194
rect 4024 -298 4100 -250
rect 4024 -354 4034 -298
rect 4090 -354 4100 -298
rect 4024 -364 4100 -354
rect 4664 -194 4740 -184
rect 4664 -250 4674 -194
rect 4730 -250 4740 -194
rect 4664 -298 4740 -250
rect 4664 -354 4674 -298
rect 4730 -354 4740 -298
rect 4664 -364 4740 -354
rect 5255 -457 5415 132
rect 5527 -184 5687 637
rect 10895 616 11055 2048
rect 11163 1808 11323 4132
rect 17155 2348 17230 4194
rect 18579 4250 18655 4260
rect 18579 4194 18589 4250
rect 18645 4194 18655 4250
rect 18579 4184 18655 4194
rect 19699 4250 19775 4260
rect 19699 4194 19709 4250
rect 19765 4194 19775 4250
rect 19699 4184 19775 4194
rect 23731 4250 23807 4260
rect 23731 4194 23741 4250
rect 23797 4194 23807 4250
rect 23731 4184 23807 4194
rect 24851 4250 24927 4260
rect 24851 4194 24861 4250
rect 24917 4194 24927 4250
rect 24851 4184 24927 4194
rect 26276 4250 26351 4260
rect 26276 4194 26285 4250
rect 26342 4194 26351 4250
rect 21611 4113 21895 4123
rect 21611 4057 21621 4113
rect 21677 4057 21725 4113
rect 21781 4057 21829 4113
rect 21885 4057 21895 4113
rect 18819 4009 18895 4019
rect 18819 3953 18829 4009
rect 18885 3953 18895 4009
rect 18819 3905 18895 3953
rect 18819 3849 18829 3905
rect 18885 3849 18895 3905
rect 18819 3839 18895 3849
rect 19459 4009 19535 4019
rect 19459 3953 19469 4009
rect 19525 3953 19535 4009
rect 19459 3905 19535 3953
rect 19459 3849 19469 3905
rect 19525 3849 19535 3905
rect 19459 3839 19535 3849
rect 21611 4009 21895 4057
rect 21611 3953 21621 4009
rect 21677 3953 21725 4009
rect 21781 3953 21829 4009
rect 21885 3953 21895 4009
rect 21611 3905 21895 3953
rect 21611 3849 21621 3905
rect 21677 3849 21725 3905
rect 21781 3849 21829 3905
rect 21885 3849 21895 3905
rect 20962 3719 21246 3729
rect 20962 3663 20972 3719
rect 21028 3663 21076 3719
rect 21132 3663 21180 3719
rect 21236 3663 21246 3719
rect 18499 3615 18575 3625
rect 18499 3559 18509 3615
rect 18565 3559 18575 3615
rect 18499 3511 18575 3559
rect 18499 3455 18509 3511
rect 18565 3455 18575 3511
rect 18499 3445 18575 3455
rect 18659 3613 18735 3625
rect 18659 3561 18671 3613
rect 18723 3561 18735 3613
rect 18659 3509 18735 3561
rect 18659 3457 18671 3509
rect 18723 3457 18735 3509
rect 18659 3445 18735 3457
rect 18979 3613 19055 3625
rect 18979 3561 18991 3613
rect 19043 3561 19055 3613
rect 18979 3509 19055 3561
rect 18979 3457 18991 3509
rect 19043 3457 19055 3509
rect 18979 3445 19055 3457
rect 19139 3615 19215 3625
rect 19139 3559 19149 3615
rect 19205 3559 19215 3615
rect 19139 3511 19215 3559
rect 19139 3455 19149 3511
rect 19205 3455 19215 3511
rect 19139 3445 19215 3455
rect 19299 3613 19375 3625
rect 19299 3561 19311 3613
rect 19363 3561 19375 3613
rect 19299 3509 19375 3561
rect 19299 3457 19311 3509
rect 19363 3457 19375 3509
rect 19299 3445 19375 3457
rect 19619 3613 19695 3625
rect 19619 3561 19631 3613
rect 19683 3561 19695 3613
rect 19619 3509 19695 3561
rect 19619 3457 19631 3509
rect 19683 3457 19695 3509
rect 19619 3445 19695 3457
rect 19779 3615 19855 3625
rect 19779 3559 19789 3615
rect 19845 3559 19855 3615
rect 19779 3511 19855 3559
rect 19779 3455 19789 3511
rect 19845 3455 19855 3511
rect 19779 3445 19855 3455
rect 20962 3615 21246 3663
rect 20962 3559 20972 3615
rect 21028 3559 21076 3615
rect 21132 3559 21180 3615
rect 21236 3559 21246 3615
rect 20962 3511 21246 3559
rect 20962 3455 20972 3511
rect 21028 3455 21076 3511
rect 21132 3455 21180 3511
rect 21236 3455 21246 3511
rect 17155 2292 17165 2348
rect 17221 2292 17230 2348
rect 12314 2218 12390 2228
rect 12314 2162 12324 2218
rect 12380 2162 12390 2218
rect 12314 2114 12390 2162
rect 12314 2058 12324 2114
rect 12380 2058 12390 2114
rect 12314 2048 12390 2058
rect 13210 2218 13286 2228
rect 13210 2162 13220 2218
rect 13276 2162 13286 2218
rect 13210 2114 13286 2162
rect 13210 2058 13220 2114
rect 13276 2058 13286 2114
rect 13210 2048 13286 2058
rect 13498 2218 13574 2228
rect 13498 2162 13508 2218
rect 13564 2162 13574 2218
rect 13498 2114 13574 2162
rect 13498 2058 13508 2114
rect 13564 2058 13574 2114
rect 13498 2048 13574 2058
rect 14660 2218 14736 2228
rect 14660 2162 14670 2218
rect 14726 2162 14736 2218
rect 14660 2114 14736 2162
rect 14660 2058 14670 2114
rect 14726 2058 14736 2114
rect 14660 2048 14736 2058
rect 15300 2218 15376 2228
rect 15300 2162 15310 2218
rect 15366 2162 15376 2218
rect 15300 2114 15376 2162
rect 15300 2058 15310 2114
rect 15366 2058 15376 2114
rect 15300 2048 15376 2058
rect 15940 2218 16016 2228
rect 15940 2162 15950 2218
rect 16006 2162 16016 2218
rect 15940 2114 16016 2162
rect 15940 2058 15950 2114
rect 16006 2058 16016 2114
rect 15940 2048 16016 2058
rect 16879 2218 17059 2228
rect 16879 2162 16889 2218
rect 16945 2162 16993 2218
rect 17049 2162 17059 2218
rect 16879 2114 17059 2162
rect 16879 2058 16889 2114
rect 16945 2058 16993 2114
rect 17049 2058 17059 2114
rect 16879 2048 17059 2058
rect 11153 1798 11333 1808
rect 11153 1742 11163 1798
rect 11219 1742 11267 1798
rect 11323 1742 11333 1798
rect 11153 1694 11333 1742
rect 11153 1638 11163 1694
rect 11219 1638 11267 1694
rect 11323 1638 11333 1694
rect 11153 1628 11333 1638
rect 11866 1798 11942 1808
rect 11866 1742 11876 1798
rect 11932 1742 11942 1798
rect 11866 1694 11942 1742
rect 11866 1638 11876 1694
rect 11932 1638 11942 1694
rect 11866 1628 11942 1638
rect 12762 1798 12838 1808
rect 12762 1742 12772 1798
rect 12828 1742 12838 1798
rect 12762 1694 12838 1742
rect 12762 1638 12772 1694
rect 12828 1638 12838 1694
rect 12762 1628 12838 1638
rect 13658 1798 13734 1808
rect 13658 1742 13668 1798
rect 13724 1742 13734 1798
rect 13658 1694 13734 1742
rect 13658 1638 13668 1694
rect 13724 1638 13734 1694
rect 13658 1628 13734 1638
rect 14980 1798 15056 1808
rect 14980 1742 14990 1798
rect 15046 1742 15056 1798
rect 14980 1694 15056 1742
rect 14980 1638 14990 1694
rect 15046 1638 15056 1694
rect 14980 1628 15056 1638
rect 15620 1798 15696 1808
rect 15620 1742 15630 1798
rect 15686 1742 15696 1798
rect 15620 1694 15696 1742
rect 15620 1638 15630 1694
rect 15686 1638 15696 1694
rect 15620 1628 15696 1638
rect 16617 1798 16797 1808
rect 16617 1742 16627 1798
rect 16683 1742 16731 1798
rect 16787 1742 16797 1798
rect 16617 1694 16797 1742
rect 16617 1638 16627 1694
rect 16683 1638 16731 1694
rect 16787 1638 16797 1694
rect 16617 1628 16797 1638
rect 11163 1278 11323 1628
rect 11153 1268 11333 1278
rect 11153 1212 11163 1268
rect 11219 1212 11267 1268
rect 11323 1212 11333 1268
rect 11153 1164 11333 1212
rect 11153 1108 11163 1164
rect 11219 1108 11267 1164
rect 11323 1108 11333 1164
rect 11153 1060 11333 1108
rect 11153 1004 11163 1060
rect 11219 1004 11267 1060
rect 11323 1004 11333 1060
rect 11153 994 11333 1004
rect 12314 1164 12390 1174
rect 12314 1108 12324 1164
rect 12380 1108 12390 1164
rect 12314 1060 12390 1108
rect 12314 1004 12324 1060
rect 12380 1004 12390 1060
rect 12314 994 12390 1004
rect 13210 1164 13286 1174
rect 13210 1108 13220 1164
rect 13276 1108 13286 1164
rect 16627 1148 16787 1628
rect 13210 1060 13286 1108
rect 13210 1004 13220 1060
rect 13276 1004 13286 1060
rect 13210 994 13286 1004
rect 13498 1138 13574 1148
rect 13498 1082 13508 1138
rect 13564 1082 13574 1138
rect 13498 1034 13574 1082
rect 10116 606 10192 616
rect 10116 550 10126 606
rect 10182 550 10192 606
rect 10116 502 10192 550
rect 10116 446 10126 502
rect 10182 446 10192 502
rect 10116 436 10192 446
rect 10885 606 11065 616
rect 10885 550 10895 606
rect 10951 550 10999 606
rect 11055 550 11065 606
rect 10885 502 11065 550
rect 10885 446 10895 502
rect 10951 446 10999 502
rect 11055 446 11065 502
rect 10885 436 11065 446
rect 6249 406 6325 416
rect 6249 350 6259 406
rect 6315 350 6325 406
rect 6249 302 6325 350
rect 6249 246 6259 302
rect 6315 246 6325 302
rect 6249 236 6325 246
rect 6889 406 6965 416
rect 6889 350 6899 406
rect 6955 350 6965 406
rect 6889 302 6965 350
rect 6889 246 6899 302
rect 6955 246 6965 302
rect 6889 236 6965 246
rect 7529 406 7605 416
rect 7529 350 7539 406
rect 7595 350 7605 406
rect 7529 302 7605 350
rect 7529 246 7539 302
rect 7595 246 7605 302
rect 7529 236 7605 246
rect 8932 406 9008 416
rect 8932 350 8942 406
rect 8998 350 9008 406
rect 8932 302 9008 350
rect 8932 246 8942 302
rect 8998 246 9008 302
rect 8932 236 9008 246
rect 9828 406 9904 416
rect 9828 350 9838 406
rect 9894 350 9904 406
rect 9828 302 9904 350
rect 9828 246 9838 302
rect 9894 246 9904 302
rect 9828 236 9904 246
rect 10895 128 11055 436
rect 10885 118 11065 128
rect 10885 62 10895 118
rect 10951 62 10999 118
rect 11055 62 11065 118
rect 10885 14 11065 62
rect 10885 -42 10895 14
rect 10951 -42 10999 14
rect 11055 -42 11065 14
rect 10885 -52 11065 -42
rect 5517 -194 5697 -184
rect 5517 -250 5527 -194
rect 5583 -250 5631 -194
rect 5687 -250 5697 -194
rect 5517 -298 5697 -250
rect 5517 -354 5527 -298
rect 5583 -354 5631 -298
rect 5687 -354 5697 -298
rect 5517 -364 5697 -354
rect 6249 -194 6325 -184
rect 6249 -250 6259 -194
rect 6315 -250 6325 -194
rect 6249 -298 6325 -250
rect 6249 -354 6259 -298
rect 6315 -354 6325 -298
rect 6249 -364 6325 -354
rect 6889 -194 6965 -184
rect 6889 -250 6899 -194
rect 6955 -250 6965 -194
rect 6889 -298 6965 -250
rect 6889 -354 6899 -298
rect 6955 -354 6965 -298
rect 6889 -364 6965 -354
rect 7529 -194 7605 -184
rect 7529 -250 7539 -194
rect 7595 -250 7605 -194
rect 7529 -298 7605 -250
rect 7529 -354 7539 -298
rect 7595 -354 7605 -298
rect 7529 -364 7605 -354
rect 8484 -194 8560 -184
rect 8484 -250 8494 -194
rect 8550 -250 8560 -194
rect 8484 -298 8560 -250
rect 8484 -354 8494 -298
rect 8550 -354 8560 -298
rect 8484 -364 8560 -354
rect 9380 -194 9456 -184
rect 9380 -250 9390 -194
rect 9446 -250 9456 -194
rect 9380 -298 9456 -250
rect 9380 -354 9390 -298
rect 9446 -354 9456 -298
rect 9380 -364 9456 -354
rect 10276 -194 10352 -184
rect 10276 -250 10286 -194
rect 10342 -250 10352 -194
rect 10276 -298 10352 -250
rect 10276 -354 10286 -298
rect 10342 -354 10352 -298
rect 10276 -364 10352 -354
rect 2675 -475 2855 -465
rect 2675 -531 2685 -475
rect 2741 -531 2789 -475
rect 2845 -531 2855 -475
rect 2675 -579 2855 -531
rect 2675 -635 2685 -579
rect 2741 -635 2789 -579
rect 2845 -635 2855 -579
rect 2675 -645 2855 -635
rect 3464 -475 3540 -465
rect 3464 -531 3474 -475
rect 3530 -531 3540 -475
rect 3464 -579 3540 -531
rect 3464 -635 3474 -579
rect 3530 -635 3540 -579
rect 3464 -645 3540 -635
rect 5245 -467 5425 -457
rect 5245 -523 5255 -467
rect 5311 -523 5359 -467
rect 5415 -523 5425 -467
rect 5245 -571 5425 -523
rect 5245 -627 5255 -571
rect 5311 -627 5359 -571
rect 5415 -627 5425 -571
rect 5245 -637 5425 -627
rect 3704 -828 3780 -818
rect 3704 -884 3714 -828
rect 3770 -884 3780 -828
rect 3704 -932 3780 -884
rect 3704 -988 3714 -932
rect 3770 -988 3780 -932
rect 3704 -998 3780 -988
rect 4345 -828 4421 -818
rect 4345 -884 4355 -828
rect 4411 -884 4421 -828
rect 4345 -932 4421 -884
rect 4345 -988 4355 -932
rect 4411 -988 4421 -932
rect 4345 -998 4421 -988
rect 3544 -1028 3620 -1018
rect 3544 -1084 3554 -1028
rect 3610 -1084 3620 -1028
rect 3544 -1132 3620 -1084
rect 3544 -1188 3554 -1132
rect 3610 -1188 3620 -1132
rect 3544 -1198 3620 -1188
rect 5255 -1314 5415 -637
rect 5527 -818 5687 -364
rect 9988 -452 10064 -442
rect 6569 -467 6645 -457
rect 6569 -523 6579 -467
rect 6635 -523 6645 -467
rect 6569 -571 6645 -523
rect 6569 -627 6579 -571
rect 6635 -627 6645 -571
rect 6569 -637 6645 -627
rect 7209 -467 7285 -457
rect 7209 -523 7219 -467
rect 7275 -523 7285 -467
rect 7209 -571 7285 -523
rect 7209 -627 7219 -571
rect 7275 -627 7285 -571
rect 9988 -508 9998 -452
rect 10054 -508 10064 -452
rect 9988 -556 10064 -508
rect 9988 -612 9998 -556
rect 10054 -612 10064 -556
rect 9988 -622 10064 -612
rect 7209 -637 7285 -627
rect 7503 -691 7579 -681
rect 7503 -747 7513 -691
rect 7569 -747 7579 -691
rect 7503 -795 7579 -747
rect 5517 -828 5697 -818
rect 5517 -884 5527 -828
rect 5583 -884 5631 -828
rect 5687 -884 5697 -828
rect 7503 -851 7513 -795
rect 7569 -851 7579 -795
rect 7503 -861 7579 -851
rect 7789 -691 7969 -681
rect 7789 -747 7799 -691
rect 7855 -747 7903 -691
rect 7959 -747 7969 -691
rect 7789 -795 7969 -747
rect 7789 -851 7799 -795
rect 7855 -851 7903 -795
rect 7959 -851 7969 -795
rect 7789 -861 7969 -851
rect 10236 -702 10312 -692
rect 10236 -758 10246 -702
rect 10302 -758 10312 -702
rect 10236 -806 10312 -758
rect 5517 -932 5697 -884
rect 5517 -988 5527 -932
rect 5583 -988 5631 -932
rect 5687 -988 5697 -932
rect 5517 -1036 5697 -988
rect 5517 -1092 5527 -1036
rect 5583 -1092 5631 -1036
rect 5687 -1092 5697 -1036
rect 5517 -1102 5697 -1092
rect 6569 -932 6645 -922
rect 6569 -988 6579 -932
rect 6635 -988 6645 -932
rect 6569 -1036 6645 -988
rect 6569 -1092 6579 -1036
rect 6635 -1092 6645 -1036
rect 6569 -1102 6645 -1092
rect 7209 -932 7285 -922
rect 7209 -988 7219 -932
rect 7275 -988 7285 -932
rect 7209 -1036 7285 -988
rect 7209 -1092 7219 -1036
rect 7275 -1092 7285 -1036
rect 7209 -1102 7285 -1092
rect 3384 -1324 3460 -1314
rect 3384 -1380 3394 -1324
rect 3450 -1380 3460 -1324
rect 3384 -1428 3460 -1380
rect 3384 -1484 3394 -1428
rect 3450 -1484 3460 -1428
rect 3384 -1494 3460 -1484
rect 4024 -1324 4100 -1314
rect 4024 -1380 4034 -1324
rect 4090 -1380 4100 -1324
rect 4024 -1428 4100 -1380
rect 4024 -1484 4034 -1428
rect 4090 -1484 4100 -1428
rect 4024 -1494 4100 -1484
rect 4664 -1324 4740 -1314
rect 4664 -1380 4674 -1324
rect 4730 -1380 4740 -1324
rect 4664 -1428 4740 -1380
rect 4664 -1484 4674 -1428
rect 4730 -1484 4740 -1428
rect 4664 -1494 4740 -1484
rect 5245 -1324 5425 -1314
rect 5245 -1380 5255 -1324
rect 5311 -1380 5359 -1324
rect 5415 -1380 5425 -1324
rect 5245 -1428 5425 -1380
rect 5245 -1484 5255 -1428
rect 5311 -1484 5359 -1428
rect 5415 -1484 5425 -1428
rect 5245 -1494 5425 -1484
rect 6249 -1324 6325 -1314
rect 6249 -1380 6259 -1324
rect 6315 -1380 6325 -1324
rect 6249 -1428 6325 -1380
rect 6249 -1484 6259 -1428
rect 6315 -1484 6325 -1428
rect 6249 -1494 6325 -1484
rect 6889 -1324 6965 -1314
rect 6889 -1380 6899 -1324
rect 6955 -1380 6965 -1324
rect 6889 -1428 6965 -1380
rect 6889 -1484 6899 -1428
rect 6955 -1484 6965 -1428
rect 6889 -1494 6965 -1484
rect 7529 -1324 7605 -1314
rect 7529 -1380 7539 -1324
rect 7595 -1380 7605 -1324
rect 7529 -1428 7605 -1380
rect 7529 -1484 7539 -1428
rect 7595 -1484 7605 -1428
rect 7529 -1494 7605 -1484
rect 741 -1732 751 -1676
rect 807 -1732 855 -1676
rect 911 -1732 921 -1676
rect 741 -1742 921 -1732
rect 2395 -1663 2575 -1653
rect 2395 -1719 2405 -1663
rect 2461 -1719 2509 -1663
rect 2565 -1719 2575 -1663
rect 751 -5986 911 -1742
rect 2395 -1767 2575 -1719
rect 2395 -1823 2405 -1767
rect 2461 -1823 2509 -1767
rect 2565 -1823 2575 -1767
rect 2395 -1833 2575 -1823
rect 3624 -1663 3700 -1653
rect 3624 -1719 3634 -1663
rect 3690 -1719 3700 -1663
rect 3624 -1767 3700 -1719
rect 3624 -1823 3634 -1767
rect 3690 -1823 3700 -1767
rect 3624 -1833 3700 -1823
rect 6381 -1778 6561 -1766
rect 6381 -1830 6393 -1778
rect 6445 -1830 6497 -1778
rect 6549 -1830 6561 -1778
rect 6381 -1882 6561 -1830
rect 6381 -1934 6393 -1882
rect 6445 -1934 6497 -1882
rect 6549 -1934 6561 -1882
rect 6381 -1946 6561 -1934
rect 6393 -2972 6553 -1946
rect 7799 -2736 7959 -861
rect 10236 -862 10246 -806
rect 10302 -862 10312 -806
rect 10236 -872 10312 -862
rect 10432 -702 10612 -692
rect 10432 -758 10442 -702
rect 10498 -758 10546 -702
rect 10602 -758 10612 -702
rect 10432 -806 10612 -758
rect 10432 -862 10442 -806
rect 10498 -862 10546 -806
rect 10602 -862 10612 -806
rect 10432 -872 10612 -862
rect 8932 -932 9008 -922
rect 8932 -988 8942 -932
rect 8998 -988 9008 -932
rect 8932 -1036 9008 -988
rect 8932 -1092 8942 -1036
rect 8998 -1092 9008 -1036
rect 8932 -1102 9008 -1092
rect 9828 -932 9904 -922
rect 9828 -988 9838 -932
rect 9894 -988 9904 -932
rect 9828 -1036 9904 -988
rect 9828 -1092 9838 -1036
rect 9894 -1092 9904 -1036
rect 9828 -1102 9904 -1092
rect 9988 -932 10064 -922
rect 9988 -988 9998 -932
rect 10054 -988 10064 -932
rect 9988 -1036 10064 -988
rect 9988 -1092 9998 -1036
rect 10054 -1092 10064 -1036
rect 9988 -1102 10064 -1092
rect 8484 -1324 8560 -1314
rect 8484 -1380 8494 -1324
rect 8550 -1380 8560 -1324
rect 8484 -1428 8560 -1380
rect 8484 -1484 8494 -1428
rect 8550 -1484 8560 -1428
rect 8484 -1494 8560 -1484
rect 9380 -1324 9456 -1314
rect 9380 -1380 9390 -1324
rect 9446 -1380 9456 -1324
rect 9380 -1428 9456 -1380
rect 9380 -1484 9390 -1428
rect 9446 -1484 9456 -1428
rect 9380 -1494 9456 -1484
rect 10276 -1324 10352 -1314
rect 10276 -1380 10286 -1324
rect 10342 -1380 10352 -1324
rect 10276 -1428 10352 -1380
rect 10276 -1484 10286 -1428
rect 10342 -1484 10352 -1428
rect 10276 -1494 10352 -1484
rect 9483 -1778 9663 -1766
rect 9483 -1830 9495 -1778
rect 9547 -1830 9599 -1778
rect 9651 -1830 9663 -1778
rect 9483 -1882 9663 -1830
rect 9483 -1934 9495 -1882
rect 9547 -1934 9599 -1882
rect 9651 -1934 9663 -1882
rect 9483 -1946 9663 -1934
rect 6896 -2746 7076 -2736
rect 6896 -2802 6906 -2746
rect 6962 -2802 7010 -2746
rect 7066 -2802 7076 -2746
rect 6896 -2850 7076 -2802
rect 6896 -2906 6906 -2850
rect 6962 -2906 7010 -2850
rect 7066 -2906 7076 -2850
rect 6896 -2916 7076 -2906
rect 7789 -2746 7969 -2736
rect 7789 -2802 7799 -2746
rect 7855 -2802 7903 -2746
rect 7959 -2802 7969 -2746
rect 7789 -2850 7969 -2802
rect 7789 -2906 7799 -2850
rect 7855 -2906 7903 -2850
rect 7959 -2906 7969 -2850
rect 7789 -2916 7969 -2906
rect 6381 -2984 6561 -2972
rect 6381 -3036 6393 -2984
rect 6445 -3036 6497 -2984
rect 6549 -3036 6561 -2984
rect 6381 -3088 6561 -3036
rect 6381 -3140 6393 -3088
rect 6445 -3140 6497 -3088
rect 6549 -3140 6561 -3088
rect 6381 -3152 6561 -3140
rect 4658 -3698 4838 -3686
rect 4658 -3750 4670 -3698
rect 4722 -3750 4774 -3698
rect 4826 -3750 4838 -3698
rect 4658 -3802 4838 -3750
rect 1689 -3849 1869 -3837
rect 1689 -3901 1701 -3849
rect 1753 -3901 1805 -3849
rect 1857 -3901 1869 -3849
rect 4658 -3854 4670 -3802
rect 4722 -3854 4774 -3802
rect 4826 -3854 4838 -3802
rect 4658 -3866 4838 -3854
rect 1689 -3953 1869 -3901
rect 1689 -4005 1701 -3953
rect 1753 -4005 1805 -3953
rect 1857 -4005 1869 -3953
rect 1689 -4017 1869 -4005
rect 2561 -3982 2741 -3972
rect 1699 -4589 1859 -4017
rect 2561 -4038 2571 -3982
rect 2627 -4038 2675 -3982
rect 2731 -4038 2741 -3982
rect 2561 -4086 2741 -4038
rect 2561 -4142 2571 -4086
rect 2627 -4142 2675 -4086
rect 2731 -4142 2741 -4086
rect 2561 -4152 2741 -4142
rect 1689 -4601 1869 -4589
rect 1689 -4653 1701 -4601
rect 1753 -4653 1805 -4601
rect 1857 -4653 1869 -4601
rect 1689 -4665 1869 -4653
rect 2229 -4736 2305 -4726
rect 2229 -4792 2239 -4736
rect 2295 -4792 2305 -4736
rect 2229 -4840 2305 -4792
rect 2229 -4896 2239 -4840
rect 2295 -4896 2305 -4840
rect 2229 -4906 2305 -4896
rect 2623 -5986 2679 -4152
rect 3525 -5026 3601 -5016
rect 3525 -5082 3535 -5026
rect 3591 -5082 3601 -5026
rect 3525 -5130 3601 -5082
rect 3525 -5186 3535 -5130
rect 3591 -5186 3601 -5130
rect 3525 -5196 3601 -5186
rect 3093 -5350 3169 -5340
rect 3093 -5406 3103 -5350
rect 3159 -5406 3169 -5350
rect 3093 -5454 3169 -5406
rect 3093 -5510 3103 -5454
rect 3159 -5510 3169 -5454
rect 3093 -5520 3169 -5510
rect 2933 -5752 3113 -5742
rect 2933 -5808 2943 -5752
rect 2999 -5808 3047 -5752
rect 3103 -5808 3113 -5752
rect 2933 -5856 3113 -5808
rect 2933 -5912 2943 -5856
rect 2999 -5912 3047 -5856
rect 3103 -5912 3113 -5856
rect 2933 -5922 3113 -5912
rect 2943 -5986 2999 -5922
rect 741 -5996 921 -5986
rect 741 -6052 751 -5996
rect 807 -6052 855 -5996
rect 911 -6052 921 -5996
rect 741 -6100 921 -6052
rect 741 -6156 751 -6100
rect 807 -6156 855 -6100
rect 911 -6156 921 -6100
rect 741 -6166 921 -6156
rect 2239 -5996 2315 -5986
rect 2239 -6052 2249 -5996
rect 2305 -6052 2315 -5996
rect 2239 -6100 2315 -6052
rect 2239 -6156 2249 -6100
rect 2305 -6156 2315 -6100
rect 2239 -6166 2315 -6156
rect 2613 -5998 2689 -5986
rect 2613 -6050 2625 -5998
rect 2677 -6050 2689 -5998
rect 2613 -6102 2689 -6050
rect 2613 -6154 2625 -6102
rect 2677 -6154 2689 -6102
rect 2613 -6166 2689 -6154
rect 2933 -5998 3009 -5986
rect 2933 -6050 2945 -5998
rect 2997 -6050 3009 -5998
rect 2933 -6102 3009 -6050
rect 2933 -6154 2945 -6102
rect 2997 -6154 3009 -6102
rect 2933 -6166 3009 -6154
rect 4668 -6602 4828 -3866
rect 5134 -4736 5314 -4726
rect 5134 -4792 5144 -4736
rect 5200 -4792 5248 -4736
rect 5304 -4792 5314 -4736
rect 5134 -4840 5314 -4792
rect 5134 -4896 5144 -4840
rect 5200 -4896 5248 -4840
rect 5304 -4896 5314 -4840
rect 5134 -4906 5314 -4896
rect 4898 -5350 5078 -5340
rect 4898 -5406 4908 -5350
rect 4964 -5406 5012 -5350
rect 5068 -5406 5078 -5350
rect 4898 -5454 5078 -5406
rect 4898 -5510 4908 -5454
rect 4964 -5510 5012 -5454
rect 5068 -5510 5078 -5454
rect 4898 -5520 5078 -5510
rect 3437 -6612 3513 -6602
rect 3437 -6668 3447 -6612
rect 3503 -6668 3513 -6612
rect 3437 -6716 3513 -6668
rect 3437 -6772 3447 -6716
rect 3503 -6772 3513 -6716
rect 3437 -6782 3513 -6772
rect 4658 -6612 4838 -6602
rect 4658 -6668 4668 -6612
rect 4724 -6668 4772 -6612
rect 4828 -6668 4838 -6612
rect 4658 -6716 4838 -6668
rect 4658 -6772 4668 -6716
rect 4724 -6772 4772 -6716
rect 4828 -6772 4838 -6716
rect 4908 -6745 5068 -5520
rect 4658 -6782 4838 -6772
rect 4898 -6755 5078 -6745
rect 4668 -7131 4828 -6782
rect 4898 -6811 4908 -6755
rect 4964 -6811 5012 -6755
rect 5068 -6811 5078 -6755
rect 4898 -6859 5078 -6811
rect 4898 -6915 4908 -6859
rect 4964 -6915 5012 -6859
rect 5068 -6915 5078 -6859
rect 4898 -6925 5078 -6915
rect 4658 -7141 4838 -7131
rect 4658 -7197 4668 -7141
rect 4724 -7197 4772 -7141
rect 4828 -7197 4838 -7141
rect 4658 -7245 4838 -7197
rect 4658 -7301 4668 -7245
rect 4724 -7301 4772 -7245
rect 4828 -7301 4838 -7245
rect 4658 -7311 4838 -7301
rect 3485 -7382 3561 -7372
rect 3485 -7438 3495 -7382
rect 3551 -7438 3561 -7382
rect 3485 -7486 3561 -7438
rect 3485 -7542 3495 -7486
rect 3551 -7542 3561 -7486
rect 3485 -7552 3561 -7542
rect 4668 -8590 4828 -7311
rect 5144 -8270 5304 -4906
rect 5607 -5026 5787 -5016
rect 5607 -5082 5617 -5026
rect 5673 -5082 5721 -5026
rect 5777 -5082 5787 -5026
rect 5607 -5130 5787 -5082
rect 5607 -5186 5617 -5130
rect 5673 -5186 5721 -5130
rect 5777 -5186 5787 -5130
rect 5607 -5196 5787 -5186
rect 6058 -5054 6238 -5044
rect 6058 -5110 6068 -5054
rect 6124 -5110 6172 -5054
rect 6228 -5110 6238 -5054
rect 6058 -5158 6238 -5110
rect 5365 -5544 5545 -5534
rect 5365 -5600 5375 -5544
rect 5431 -5600 5479 -5544
rect 5535 -5600 5545 -5544
rect 5365 -5648 5545 -5600
rect 5365 -5704 5375 -5648
rect 5431 -5704 5479 -5648
rect 5535 -5704 5545 -5648
rect 5365 -5752 5545 -5704
rect 5365 -5808 5375 -5752
rect 5431 -5808 5479 -5752
rect 5535 -5808 5545 -5752
rect 5365 -5856 5545 -5808
rect 5365 -5912 5375 -5856
rect 5431 -5912 5479 -5856
rect 5535 -5912 5545 -5856
rect 5365 -5922 5545 -5912
rect 5617 -6258 5777 -5196
rect 6058 -5214 6068 -5158
rect 6124 -5214 6172 -5158
rect 6228 -5214 6238 -5158
rect 6058 -5224 6238 -5214
rect 6368 -5054 6548 -5044
rect 6368 -5110 6378 -5054
rect 6434 -5110 6482 -5054
rect 6538 -5110 6548 -5054
rect 6368 -5158 6548 -5110
rect 6368 -5214 6378 -5158
rect 6434 -5214 6482 -5158
rect 6538 -5214 6548 -5158
rect 6368 -5224 6548 -5214
rect 5607 -6268 5787 -6258
rect 5607 -6324 5617 -6268
rect 5673 -6324 5721 -6268
rect 5777 -6324 5787 -6268
rect 5607 -6372 5787 -6324
rect 5607 -6428 5617 -6372
rect 5673 -6428 5721 -6372
rect 5777 -6428 5787 -6372
rect 5607 -6438 5787 -6428
rect 6096 -6755 6172 -6745
rect 6096 -6811 6106 -6755
rect 6162 -6811 6172 -6755
rect 6096 -6859 6172 -6811
rect 6096 -6915 6106 -6859
rect 6162 -6915 6172 -6859
rect 6096 -6925 6172 -6915
rect 6026 -7141 6206 -7131
rect 6026 -7197 6036 -7141
rect 6092 -7197 6140 -7141
rect 6196 -7197 6206 -7141
rect 6026 -7245 6206 -7197
rect 6026 -7301 6036 -7245
rect 6092 -7301 6140 -7245
rect 6196 -7301 6206 -7245
rect 6026 -7311 6206 -7301
rect 5936 -7384 6012 -7374
rect 6378 -7380 6538 -5224
rect 6632 -6268 6812 -6258
rect 6632 -6324 6642 -6268
rect 6698 -6324 6746 -6268
rect 6802 -6324 6812 -6268
rect 6632 -6372 6812 -6324
rect 6632 -6428 6642 -6372
rect 6698 -6428 6746 -6372
rect 6802 -6428 6812 -6372
rect 6632 -6438 6812 -6428
rect 6642 -7141 6802 -6438
rect 6906 -6504 7066 -2916
rect 9493 -2972 9653 -1946
rect 9483 -2984 9663 -2972
rect 9483 -3036 9495 -2984
rect 9547 -3036 9599 -2984
rect 9651 -3036 9663 -2984
rect 9483 -3088 9663 -3036
rect 8703 -3113 8779 -3103
rect 8703 -3169 8713 -3113
rect 8769 -3169 8779 -3113
rect 9483 -3140 9495 -3088
rect 9547 -3140 9599 -3088
rect 9651 -3140 9663 -3088
rect 9483 -3152 9663 -3140
rect 9792 -3113 9972 -3103
rect 8703 -3217 8779 -3169
rect 8703 -3273 8713 -3217
rect 8769 -3273 8779 -3217
rect 8703 -3283 8779 -3273
rect 9792 -3169 9802 -3113
rect 9858 -3169 9906 -3113
rect 9962 -3169 9972 -3113
rect 9792 -3217 9972 -3169
rect 9792 -3273 9802 -3217
rect 9858 -3273 9906 -3217
rect 9962 -3273 9972 -3217
rect 9792 -3283 9972 -3273
rect 7183 -3448 7259 -3436
rect 7183 -3500 7195 -3448
rect 7247 -3500 7259 -3448
rect 7183 -3552 7259 -3500
rect 7183 -3604 7195 -3552
rect 7247 -3604 7259 -3552
rect 7183 -3616 7259 -3604
rect 7343 -3446 7419 -3436
rect 7343 -3502 7353 -3446
rect 7409 -3502 7419 -3446
rect 7343 -3550 7419 -3502
rect 7343 -3606 7353 -3550
rect 7409 -3606 7419 -3550
rect 7343 -3616 7419 -3606
rect 7663 -3446 7739 -3436
rect 7663 -3502 7673 -3446
rect 7729 -3502 7739 -3446
rect 7663 -3550 7739 -3502
rect 7663 -3606 7673 -3550
rect 7729 -3606 7739 -3550
rect 7663 -3616 7739 -3606
rect 7983 -3446 8059 -3436
rect 7983 -3502 7993 -3446
rect 8049 -3502 8059 -3446
rect 7983 -3550 8059 -3502
rect 7983 -3606 7993 -3550
rect 8049 -3606 8059 -3550
rect 7983 -3616 8059 -3606
rect 8303 -3446 8379 -3436
rect 8303 -3502 8313 -3446
rect 8369 -3502 8379 -3446
rect 8303 -3550 8379 -3502
rect 8303 -3606 8313 -3550
rect 8369 -3606 8379 -3550
rect 8303 -3616 8379 -3606
rect 8463 -3446 8539 -3437
rect 8463 -3502 8473 -3446
rect 8529 -3502 8539 -3446
rect 8463 -3550 8539 -3502
rect 8463 -3606 8473 -3550
rect 8529 -3606 8539 -3550
rect 7193 -4508 7249 -3616
rect 7353 -3972 7409 -3616
rect 8463 -3617 8539 -3606
rect 8623 -3448 8699 -3436
rect 8623 -3500 8635 -3448
rect 8687 -3500 8699 -3448
rect 8623 -3552 8699 -3500
rect 8623 -3604 8635 -3552
rect 8687 -3604 8699 -3552
rect 8623 -3616 8699 -3604
rect 7343 -3984 7419 -3972
rect 7343 -4036 7355 -3984
rect 7407 -4036 7419 -3984
rect 7343 -4088 7419 -4036
rect 7343 -4140 7355 -4088
rect 7407 -4140 7419 -4088
rect 7343 -4152 7419 -4140
rect 7503 -3982 7579 -3973
rect 7503 -4038 7513 -3982
rect 7569 -4038 7579 -3982
rect 7503 -4086 7579 -4038
rect 7503 -4142 7513 -4086
rect 7569 -4142 7579 -4086
rect 7353 -4508 7409 -4152
rect 7503 -4153 7579 -4142
rect 7663 -3982 7739 -3972
rect 7663 -4038 7673 -3982
rect 7729 -4038 7739 -3982
rect 7663 -4086 7739 -4038
rect 7663 -4142 7673 -4086
rect 7729 -4142 7739 -4086
rect 7663 -4152 7739 -4142
rect 7983 -3982 8059 -3972
rect 7983 -4038 7993 -3982
rect 8049 -4038 8059 -3982
rect 7983 -4086 8059 -4038
rect 7983 -4142 7993 -4086
rect 8049 -4142 8059 -4086
rect 7983 -4152 8059 -4142
rect 8303 -3982 8379 -3972
rect 8303 -4038 8313 -3982
rect 8369 -4038 8379 -3982
rect 8303 -4086 8379 -4038
rect 8303 -4142 8313 -4086
rect 8369 -4142 8379 -4086
rect 8303 -4152 8379 -4142
rect 7183 -4520 7259 -4508
rect 7183 -4572 7195 -4520
rect 7247 -4572 7259 -4520
rect 7183 -4624 7259 -4572
rect 7183 -4676 7195 -4624
rect 7247 -4676 7259 -4624
rect 7183 -4688 7259 -4676
rect 7343 -4518 7419 -4508
rect 7343 -4574 7353 -4518
rect 7409 -4574 7419 -4518
rect 7343 -4622 7419 -4574
rect 7343 -4678 7353 -4622
rect 7409 -4678 7419 -4622
rect 7343 -4688 7419 -4678
rect 7353 -5044 7409 -4688
rect 7343 -5054 7419 -5044
rect 7513 -5045 7569 -4153
rect 7673 -4508 7729 -4152
rect 8473 -4508 8529 -3617
rect 8633 -3972 8689 -3616
rect 8782 -3753 8858 -3743
rect 8782 -3809 8792 -3753
rect 8848 -3809 8858 -3753
rect 8782 -3819 8858 -3809
rect 8623 -3982 8699 -3972
rect 8623 -4038 8633 -3982
rect 8689 -4038 8699 -3982
rect 8623 -4086 8699 -4038
rect 8623 -4142 8633 -4086
rect 8689 -4142 8699 -4086
rect 8623 -4152 8699 -4142
rect 9802 -4227 9962 -3283
rect 10058 -3711 10238 -3701
rect 10058 -3767 10068 -3711
rect 10124 -3767 10172 -3711
rect 10228 -3767 10238 -3711
rect 10058 -3815 10238 -3767
rect 10058 -3871 10068 -3815
rect 10124 -3871 10172 -3815
rect 10228 -3871 10238 -3815
rect 10058 -3881 10238 -3871
rect 9792 -4237 9972 -4227
rect 8585 -4289 8661 -4279
rect 8585 -4345 8595 -4289
rect 8651 -4345 8661 -4289
rect 8585 -4355 8661 -4345
rect 9792 -4293 9802 -4237
rect 9858 -4293 9906 -4237
rect 9962 -4293 9972 -4237
rect 9792 -4341 9972 -4293
rect 9792 -4397 9802 -4341
rect 9858 -4397 9906 -4341
rect 9962 -4397 9972 -4341
rect 9792 -4407 9972 -4397
rect 7663 -4518 7739 -4508
rect 7663 -4574 7673 -4518
rect 7729 -4574 7739 -4518
rect 7663 -4622 7739 -4574
rect 7663 -4678 7673 -4622
rect 7729 -4678 7739 -4622
rect 7663 -4688 7739 -4678
rect 7983 -4518 8059 -4508
rect 7983 -4574 7993 -4518
rect 8049 -4574 8059 -4518
rect 7983 -4622 8059 -4574
rect 7983 -4678 7993 -4622
rect 8049 -4678 8059 -4622
rect 7983 -4688 8059 -4678
rect 8303 -4518 8379 -4508
rect 8303 -4574 8313 -4518
rect 8369 -4574 8379 -4518
rect 8303 -4622 8379 -4574
rect 8303 -4678 8313 -4622
rect 8369 -4678 8379 -4622
rect 8303 -4688 8379 -4678
rect 8463 -4520 8539 -4508
rect 8463 -4572 8475 -4520
rect 8527 -4572 8539 -4520
rect 8463 -4624 8539 -4572
rect 8463 -4676 8475 -4624
rect 8527 -4676 8539 -4624
rect 8463 -4689 8539 -4676
rect 8623 -4518 8699 -4508
rect 8623 -4574 8633 -4518
rect 8689 -4574 8699 -4518
rect 8623 -4622 8699 -4574
rect 8623 -4678 8633 -4622
rect 8689 -4678 8699 -4622
rect 8623 -4688 8699 -4678
rect 7343 -5110 7353 -5054
rect 7409 -5110 7419 -5054
rect 7343 -5158 7419 -5110
rect 7343 -5214 7353 -5158
rect 7409 -5214 7419 -5158
rect 7343 -5224 7419 -5214
rect 7503 -5056 7579 -5045
rect 7503 -5108 7515 -5056
rect 7567 -5108 7579 -5056
rect 7503 -5160 7579 -5108
rect 7503 -5212 7515 -5160
rect 7567 -5212 7579 -5160
rect 7353 -5572 7409 -5224
rect 7503 -5225 7579 -5212
rect 7663 -5054 7739 -5044
rect 7663 -5110 7673 -5054
rect 7729 -5110 7739 -5054
rect 7663 -5158 7739 -5110
rect 7663 -5214 7673 -5158
rect 7729 -5214 7739 -5158
rect 7663 -5224 7739 -5214
rect 7983 -5054 8059 -5044
rect 7983 -5110 7993 -5054
rect 8049 -5110 8059 -5054
rect 7983 -5158 8059 -5110
rect 7983 -5214 7993 -5158
rect 8049 -5214 8059 -5158
rect 7983 -5224 8059 -5214
rect 8303 -5054 8379 -5044
rect 8303 -5110 8313 -5054
rect 8369 -5110 8379 -5054
rect 8303 -5158 8379 -5110
rect 8303 -5214 8313 -5158
rect 8369 -5214 8379 -5158
rect 8303 -5224 8379 -5214
rect 7343 -5584 7419 -5572
rect 7343 -5636 7355 -5584
rect 7407 -5636 7419 -5584
rect 7343 -5688 7419 -5636
rect 7343 -5740 7355 -5688
rect 7407 -5740 7419 -5688
rect 7343 -5752 7419 -5740
rect 7353 -6108 7409 -5752
rect 7343 -6120 7419 -6108
rect 7513 -6117 7569 -5225
rect 7673 -5572 7729 -5224
rect 7993 -5572 8049 -5224
rect 8313 -5572 8369 -5224
rect 7663 -5584 7739 -5572
rect 7663 -5636 7675 -5584
rect 7727 -5636 7739 -5584
rect 7663 -5688 7739 -5636
rect 7663 -5740 7675 -5688
rect 7727 -5740 7739 -5688
rect 7663 -5752 7739 -5740
rect 7983 -5584 8059 -5572
rect 7983 -5636 7995 -5584
rect 8047 -5636 8059 -5584
rect 7983 -5688 8059 -5636
rect 7983 -5740 7995 -5688
rect 8047 -5740 8059 -5688
rect 7983 -5752 8059 -5740
rect 8303 -5584 8379 -5572
rect 8473 -5580 8529 -4689
rect 8703 -4823 8779 -4813
rect 8703 -4879 8713 -4823
rect 8769 -4879 8779 -4823
rect 8703 -4889 8779 -4879
rect 8623 -5054 8699 -5044
rect 8623 -5110 8633 -5054
rect 8689 -5110 8699 -5054
rect 8623 -5158 8699 -5110
rect 8623 -5214 8633 -5158
rect 8689 -5214 8699 -5158
rect 8623 -5224 8699 -5214
rect 8633 -5572 8689 -5224
rect 8782 -5255 8858 -5245
rect 8782 -5311 8792 -5255
rect 8848 -5311 8858 -5255
rect 8782 -5359 8858 -5311
rect 8782 -5415 8792 -5359
rect 8848 -5415 8858 -5359
rect 8782 -5425 8858 -5415
rect 9520 -5255 9700 -5245
rect 9802 -5247 9962 -4407
rect 10068 -4761 10228 -3881
rect 10058 -4771 10238 -4761
rect 10058 -4827 10068 -4771
rect 10124 -4827 10172 -4771
rect 10228 -4827 10238 -4771
rect 10058 -4875 10238 -4827
rect 10058 -4931 10068 -4875
rect 10124 -4931 10172 -4875
rect 10228 -4931 10238 -4875
rect 10058 -4941 10238 -4931
rect 9520 -5311 9530 -5255
rect 9586 -5311 9634 -5255
rect 9690 -5311 9700 -5255
rect 9520 -5359 9700 -5311
rect 9520 -5415 9530 -5359
rect 9586 -5415 9634 -5359
rect 9690 -5415 9700 -5359
rect 9520 -5425 9700 -5415
rect 9792 -5257 9972 -5247
rect 9792 -5313 9802 -5257
rect 9858 -5313 9906 -5257
rect 9962 -5313 9972 -5257
rect 9792 -5361 9972 -5313
rect 9792 -5417 9802 -5361
rect 9858 -5417 9906 -5361
rect 9962 -5417 9972 -5361
rect 8303 -5636 8315 -5584
rect 8367 -5636 8379 -5584
rect 8303 -5688 8379 -5636
rect 8303 -5740 8315 -5688
rect 8367 -5740 8379 -5688
rect 8303 -5752 8379 -5740
rect 8463 -5590 8539 -5580
rect 8463 -5646 8473 -5590
rect 8529 -5646 8539 -5590
rect 8463 -5694 8539 -5646
rect 8463 -5750 8473 -5694
rect 8529 -5750 8539 -5694
rect 7673 -6108 7729 -5752
rect 7993 -6108 8049 -5752
rect 8313 -6108 8369 -5752
rect 8463 -5761 8539 -5750
rect 8623 -5584 8699 -5572
rect 8623 -5636 8635 -5584
rect 8687 -5636 8699 -5584
rect 8623 -5688 8699 -5636
rect 8623 -5740 8635 -5688
rect 8687 -5740 8699 -5688
rect 8623 -5752 8699 -5740
rect 8633 -6108 8689 -5752
rect 8782 -5770 8858 -5760
rect 8782 -5826 8792 -5770
rect 8848 -5826 8858 -5770
rect 8782 -5874 8858 -5826
rect 8782 -5930 8792 -5874
rect 8848 -5930 8858 -5874
rect 8782 -5940 8858 -5930
rect 9253 -5996 9433 -5986
rect 9253 -6052 9263 -5996
rect 9319 -6052 9367 -5996
rect 9423 -6052 9433 -5996
rect 9253 -6100 9433 -6052
rect 7343 -6172 7355 -6120
rect 7407 -6172 7419 -6120
rect 7343 -6224 7419 -6172
rect 7343 -6276 7355 -6224
rect 7407 -6276 7419 -6224
rect 7343 -6288 7419 -6276
rect 7503 -6128 7579 -6117
rect 7503 -6180 7515 -6128
rect 7567 -6180 7579 -6128
rect 7503 -6232 7579 -6180
rect 7503 -6284 7515 -6232
rect 7567 -6284 7579 -6232
rect 7503 -6297 7579 -6284
rect 7663 -6120 7739 -6108
rect 7663 -6172 7675 -6120
rect 7727 -6172 7739 -6120
rect 7663 -6224 7739 -6172
rect 7663 -6276 7675 -6224
rect 7727 -6276 7739 -6224
rect 7663 -6288 7739 -6276
rect 7983 -6120 8059 -6108
rect 7983 -6172 7995 -6120
rect 8047 -6172 8059 -6120
rect 7983 -6224 8059 -6172
rect 7983 -6276 7995 -6224
rect 8047 -6276 8059 -6224
rect 7983 -6288 8059 -6276
rect 8303 -6120 8379 -6108
rect 8303 -6172 8315 -6120
rect 8367 -6172 8379 -6120
rect 8303 -6224 8379 -6172
rect 8303 -6276 8315 -6224
rect 8367 -6276 8379 -6224
rect 8303 -6288 8379 -6276
rect 8623 -6120 8699 -6108
rect 8623 -6172 8635 -6120
rect 8687 -6172 8699 -6120
rect 9253 -6156 9263 -6100
rect 9319 -6156 9367 -6100
rect 9423 -6156 9433 -6100
rect 9253 -6166 9433 -6156
rect 8623 -6224 8699 -6172
rect 8623 -6276 8635 -6224
rect 8687 -6276 8699 -6224
rect 8623 -6288 8699 -6276
rect 8383 -6446 8459 -6436
rect 8383 -6502 8393 -6446
rect 8449 -6502 8459 -6446
rect 6898 -6518 7078 -6504
rect 6898 -6570 6908 -6518
rect 6960 -6570 7012 -6518
rect 7064 -6570 7078 -6518
rect 6898 -6622 7078 -6570
rect 8383 -6550 8459 -6502
rect 8383 -6606 8393 -6550
rect 8449 -6606 8459 -6550
rect 8383 -6616 8459 -6606
rect 6898 -6674 6908 -6622
rect 6960 -6674 7012 -6622
rect 7064 -6674 7078 -6622
rect 6898 -6684 7078 -6674
rect 9263 -6741 9423 -6166
rect 9530 -6436 9690 -5425
rect 9792 -5427 9972 -5417
rect 10068 -5760 10228 -4941
rect 10058 -5770 10238 -5760
rect 10058 -5826 10068 -5770
rect 10124 -5826 10172 -5770
rect 10228 -5826 10238 -5770
rect 10058 -5874 10238 -5826
rect 10058 -5930 10068 -5874
rect 10124 -5930 10172 -5874
rect 10228 -5930 10238 -5874
rect 10058 -5940 10238 -5930
rect 9520 -6446 9700 -6436
rect 9520 -6502 9530 -6446
rect 9586 -6502 9634 -6446
rect 9690 -6502 9700 -6446
rect 9520 -6550 9700 -6502
rect 9520 -6606 9530 -6550
rect 9586 -6606 9634 -6550
rect 9690 -6606 9700 -6550
rect 9520 -6616 9700 -6606
rect 9827 -6521 10007 -6509
rect 9827 -6573 9839 -6521
rect 9891 -6573 9943 -6521
rect 9995 -6573 10007 -6521
rect 9827 -6625 10007 -6573
rect 9827 -6677 9839 -6625
rect 9891 -6677 9943 -6625
rect 9995 -6677 10007 -6625
rect 9827 -6689 10007 -6677
rect 9251 -6753 9431 -6741
rect 9251 -6805 9263 -6753
rect 9315 -6805 9367 -6753
rect 9419 -6805 9431 -6753
rect 9251 -6857 9431 -6805
rect 9251 -6909 9263 -6857
rect 9315 -6909 9367 -6857
rect 9419 -6909 9431 -6857
rect 9251 -6921 9431 -6909
rect 6632 -7151 6812 -7141
rect 6632 -7207 6642 -7151
rect 6698 -7207 6746 -7151
rect 6802 -7207 6812 -7151
rect 6632 -7255 6812 -7207
rect 6632 -7311 6642 -7255
rect 6698 -7311 6746 -7255
rect 6802 -7311 6812 -7255
rect 6632 -7321 6812 -7311
rect 8910 -7151 9090 -7141
rect 8910 -7207 8920 -7151
rect 8976 -7207 9024 -7151
rect 9080 -7207 9090 -7151
rect 8910 -7255 9090 -7207
rect 8910 -7311 8920 -7255
rect 8976 -7311 9024 -7255
rect 9080 -7311 9090 -7255
rect 8910 -7321 9090 -7311
rect 5936 -7440 5946 -7384
rect 6002 -7440 6012 -7384
rect 5936 -7488 6012 -7440
rect 5936 -7544 5946 -7488
rect 6002 -7544 6012 -7488
rect 5936 -7554 6012 -7544
rect 6368 -7390 6548 -7380
rect 6368 -7446 6378 -7390
rect 6434 -7446 6482 -7390
rect 6538 -7446 6548 -7390
rect 6368 -7494 6548 -7446
rect 6368 -7550 6378 -7494
rect 6434 -7550 6482 -7494
rect 6538 -7550 6548 -7494
rect 5946 -8018 6002 -7554
rect 6368 -7560 6548 -7550
rect 5884 -8028 6064 -8018
rect 5884 -8084 5894 -8028
rect 5950 -8084 5998 -8028
rect 6054 -8084 6064 -8028
rect 5884 -8132 6064 -8084
rect 5884 -8188 5894 -8132
rect 5950 -8188 5998 -8132
rect 6054 -8188 6064 -8132
rect 5884 -8198 6064 -8188
rect 9837 -8270 9997 -6689
rect 10442 -7141 10602 -872
rect 10895 -922 11055 -52
rect 11163 -442 11323 994
rect 13498 978 13508 1034
rect 13564 978 13574 1034
rect 13498 968 13574 978
rect 14660 1138 14736 1148
rect 14660 1082 14670 1138
rect 14726 1082 14736 1138
rect 14660 1034 14736 1082
rect 14660 978 14670 1034
rect 14726 978 14736 1034
rect 14660 968 14736 978
rect 15300 1138 15376 1148
rect 15300 1082 15310 1138
rect 15366 1082 15376 1138
rect 15300 1034 15376 1082
rect 15300 978 15310 1034
rect 15366 978 15376 1034
rect 15300 968 15376 978
rect 15940 1138 16016 1148
rect 15940 1082 15950 1138
rect 16006 1082 16016 1138
rect 15940 1034 16016 1082
rect 15940 978 15950 1034
rect 16006 978 16016 1034
rect 15940 968 16016 978
rect 16617 1138 16797 1148
rect 16617 1082 16627 1138
rect 16683 1082 16731 1138
rect 16787 1082 16797 1138
rect 16617 1034 16797 1082
rect 16617 978 16627 1034
rect 16683 978 16731 1034
rect 16787 978 16797 1034
rect 16617 968 16797 978
rect 11866 118 11942 128
rect 11866 62 11876 118
rect 11932 62 11942 118
rect 11866 14 11942 62
rect 11866 -42 11876 14
rect 11932 -42 11942 14
rect 11866 -52 11942 -42
rect 12762 118 12838 128
rect 12762 62 12772 118
rect 12828 62 12838 118
rect 12762 14 12838 62
rect 12762 -42 12772 14
rect 12828 -42 12838 14
rect 12762 -52 12838 -42
rect 13658 118 13734 128
rect 13658 62 13668 118
rect 13724 62 13734 118
rect 13658 14 13734 62
rect 13658 -42 13668 14
rect 13724 -42 13734 14
rect 13658 -52 13734 -42
rect 13370 -282 13446 -272
rect 13370 -338 13380 -282
rect 13436 -338 13446 -282
rect 13370 -386 13446 -338
rect 13370 -442 13380 -386
rect 13436 -442 13446 -386
rect 11153 -452 11333 -442
rect 13370 -452 13446 -442
rect 14980 -282 15056 -272
rect 14980 -338 14990 -282
rect 15046 -338 15056 -282
rect 14980 -386 15056 -338
rect 14980 -442 14990 -386
rect 15046 -442 15056 -386
rect 14980 -452 15056 -442
rect 15620 -282 15696 -272
rect 15620 -338 15630 -282
rect 15686 -338 15696 -282
rect 15620 -386 15696 -338
rect 15620 -442 15630 -386
rect 15686 -442 15696 -386
rect 15620 -452 15696 -442
rect 11153 -508 11163 -452
rect 11219 -508 11267 -452
rect 11323 -508 11333 -452
rect 11153 -556 11333 -508
rect 11153 -612 11163 -556
rect 11219 -612 11267 -556
rect 11323 -612 11333 -556
rect 11153 -622 11333 -612
rect 11532 -592 11712 -582
rect 10885 -932 11065 -922
rect 10885 -988 10895 -932
rect 10951 -988 10999 -932
rect 11055 -988 11065 -932
rect 10885 -1036 11065 -988
rect 10885 -1092 10895 -1036
rect 10951 -1092 10999 -1036
rect 11055 -1092 11065 -1036
rect 10885 -1102 11065 -1092
rect 10895 -2709 11055 -1102
rect 11163 -1322 11323 -622
rect 11532 -648 11542 -592
rect 11598 -648 11646 -592
rect 11702 -648 11712 -592
rect 11532 -696 11712 -648
rect 11532 -752 11542 -696
rect 11598 -752 11646 -696
rect 11702 -752 11712 -696
rect 11532 -762 11712 -752
rect 11902 -592 11978 -582
rect 11902 -648 11912 -592
rect 11968 -648 11978 -592
rect 11902 -696 11978 -648
rect 11902 -752 11912 -696
rect 11968 -752 11978 -696
rect 11902 -762 11978 -752
rect 14200 -587 14380 -577
rect 14200 -643 14210 -587
rect 14266 -643 14314 -587
rect 14370 -643 14380 -587
rect 14200 -691 14380 -643
rect 14200 -747 14210 -691
rect 14266 -747 14314 -691
rect 14370 -747 14380 -691
rect 14200 -757 14380 -747
rect 14688 -587 14764 -577
rect 14688 -643 14698 -587
rect 14754 -643 14764 -587
rect 14688 -691 14764 -643
rect 14688 -747 14698 -691
rect 14754 -747 14764 -691
rect 14688 -757 14764 -747
rect 11153 -1332 11333 -1322
rect 11153 -1388 11163 -1332
rect 11219 -1388 11267 -1332
rect 11323 -1388 11333 -1332
rect 11153 -1436 11333 -1388
rect 11153 -1492 11163 -1436
rect 11219 -1492 11267 -1436
rect 11323 -1492 11333 -1436
rect 11153 -1502 11333 -1492
rect 10885 -2721 11065 -2709
rect 10885 -2773 10897 -2721
rect 10949 -2773 11001 -2721
rect 11053 -2773 11065 -2721
rect 10885 -2825 11065 -2773
rect 10885 -2877 10897 -2825
rect 10949 -2877 11001 -2825
rect 11053 -2877 11065 -2825
rect 10885 -2929 11065 -2877
rect 10885 -2981 10897 -2929
rect 10949 -2981 11001 -2929
rect 11053 -2981 11065 -2929
rect 10885 -2993 11065 -2981
rect 11163 -3051 11323 -1502
rect 11153 -3063 11333 -3051
rect 11153 -3115 11165 -3063
rect 11217 -3115 11269 -3063
rect 11321 -3115 11333 -3063
rect 11153 -3167 11333 -3115
rect 11153 -3219 11165 -3167
rect 11217 -3219 11269 -3167
rect 11321 -3219 11333 -3167
rect 11153 -3271 11333 -3219
rect 11153 -3323 11165 -3271
rect 11217 -3323 11269 -3271
rect 11321 -3323 11333 -3271
rect 11153 -3335 11333 -3323
rect 10432 -7151 10612 -7141
rect 10432 -7207 10442 -7151
rect 10498 -7207 10546 -7151
rect 10602 -7207 10612 -7151
rect 10432 -7255 10612 -7207
rect 10432 -7311 10442 -7255
rect 10498 -7311 10546 -7255
rect 10602 -7311 10612 -7255
rect 10432 -7321 10612 -7311
rect 10819 -7151 10999 -7141
rect 10819 -7207 10829 -7151
rect 10885 -7207 10933 -7151
rect 10989 -7207 10999 -7151
rect 10819 -7255 10999 -7207
rect 10819 -7311 10829 -7255
rect 10885 -7311 10933 -7255
rect 10989 -7311 10999 -7255
rect 10819 -7321 10999 -7311
rect 11542 -8018 11702 -762
rect 12314 -932 12390 -922
rect 12314 -988 12324 -932
rect 12380 -988 12390 -932
rect 12314 -1036 12390 -988
rect 12314 -1092 12324 -1036
rect 12380 -1092 12390 -1036
rect 12314 -1102 12390 -1092
rect 13210 -932 13286 -922
rect 13210 -988 13220 -932
rect 13276 -988 13286 -932
rect 13210 -1036 13286 -988
rect 13210 -1092 13220 -1036
rect 13276 -1092 13286 -1036
rect 13210 -1102 13286 -1092
rect 13370 -932 13446 -922
rect 13370 -988 13380 -932
rect 13436 -988 13446 -932
rect 13370 -1036 13446 -988
rect 13370 -1092 13380 -1036
rect 13436 -1092 13446 -1036
rect 13370 -1102 13446 -1092
rect 11866 -1332 11942 -1322
rect 11866 -1388 11876 -1332
rect 11932 -1388 11942 -1332
rect 11866 -1436 11942 -1388
rect 11866 -1492 11876 -1436
rect 11932 -1492 11942 -1436
rect 11866 -1502 11942 -1492
rect 12762 -1332 12838 -1322
rect 12762 -1388 12772 -1332
rect 12828 -1388 12838 -1332
rect 12762 -1436 12838 -1388
rect 12762 -1492 12772 -1436
rect 12828 -1492 12838 -1436
rect 12762 -1502 12838 -1492
rect 13658 -1332 13734 -1322
rect 13658 -1388 13668 -1332
rect 13724 -1388 13734 -1332
rect 13658 -1436 13734 -1388
rect 13658 -1492 13668 -1436
rect 13724 -1492 13734 -1436
rect 13658 -1502 13734 -1492
rect 14210 -3436 14370 -757
rect 16627 -922 16787 968
rect 16889 -272 17049 2048
rect 16879 -282 17059 -272
rect 16879 -338 16889 -282
rect 16945 -338 16993 -282
rect 17049 -338 17059 -282
rect 16879 -386 17059 -338
rect 16879 -442 16889 -386
rect 16945 -442 16993 -386
rect 17049 -442 17059 -386
rect 16879 -452 17059 -442
rect 14980 -932 15056 -922
rect 14980 -988 14990 -932
rect 15046 -988 15056 -932
rect 14980 -1036 15056 -988
rect 14980 -1092 14990 -1036
rect 15046 -1092 15056 -1036
rect 14980 -1102 15056 -1092
rect 15620 -932 15696 -922
rect 15620 -988 15630 -932
rect 15686 -988 15696 -932
rect 15620 -1036 15696 -988
rect 15620 -1092 15630 -1036
rect 15686 -1092 15696 -1036
rect 15620 -1102 15696 -1092
rect 16617 -932 16797 -922
rect 16617 -988 16627 -932
rect 16683 -988 16731 -932
rect 16787 -988 16797 -932
rect 16617 -1036 16797 -988
rect 16617 -1092 16627 -1036
rect 16683 -1092 16731 -1036
rect 16787 -1092 16797 -1036
rect 16617 -1102 16797 -1092
rect 16889 -1312 17049 -452
rect 17155 -460 17230 2292
rect 17155 -516 17165 -460
rect 17221 -516 17230 -460
rect 17155 -526 17230 -516
rect 17355 3284 17431 3294
rect 17355 3228 17365 3284
rect 17421 3228 17431 3284
rect 17355 476 17431 3228
rect 18579 3284 18655 3294
rect 18579 3228 18589 3284
rect 18645 3228 18655 3284
rect 18579 3218 18655 3228
rect 18819 3073 18895 3083
rect 18819 3017 18829 3073
rect 18885 3017 18895 3073
rect 18819 2969 18895 3017
rect 18819 2913 18829 2969
rect 18885 2913 18895 2969
rect 18819 2903 18895 2913
rect 18989 2689 19045 3445
rect 19309 2689 19365 3445
rect 19459 3073 19535 3083
rect 19459 3017 19469 3073
rect 19525 3017 19535 3073
rect 19459 2969 19535 3017
rect 19459 2913 19469 2969
rect 19525 2913 19535 2969
rect 19459 2903 19535 2913
rect 19629 2689 19685 3445
rect 20962 3177 21246 3455
rect 20962 3121 20972 3177
rect 21028 3121 21076 3177
rect 21132 3121 21180 3177
rect 21236 3121 21246 3177
rect 20962 3073 21246 3121
rect 20962 3017 20972 3073
rect 21028 3017 21076 3073
rect 21132 3017 21180 3073
rect 21236 3017 21246 3073
rect 20962 2969 21246 3017
rect 20962 2913 20972 2969
rect 21028 2913 21076 2969
rect 21132 2913 21180 2969
rect 21236 2913 21246 2969
rect 18499 2679 18575 2689
rect 18499 2623 18509 2679
rect 18565 2623 18575 2679
rect 18499 2575 18575 2623
rect 18499 2519 18509 2575
rect 18565 2519 18575 2575
rect 18499 2509 18575 2519
rect 18659 2677 18735 2689
rect 18659 2625 18671 2677
rect 18723 2625 18735 2677
rect 18659 2573 18735 2625
rect 18659 2521 18671 2573
rect 18723 2521 18735 2573
rect 18659 2509 18735 2521
rect 18979 2677 19055 2689
rect 18979 2625 18991 2677
rect 19043 2625 19055 2677
rect 18979 2573 19055 2625
rect 18979 2521 18991 2573
rect 19043 2521 19055 2573
rect 18979 2509 19055 2521
rect 19139 2679 19215 2689
rect 19139 2623 19149 2679
rect 19205 2623 19215 2679
rect 19139 2575 19215 2623
rect 19139 2519 19149 2575
rect 19205 2519 19215 2575
rect 19139 2509 19215 2519
rect 19299 2677 19375 2689
rect 19299 2625 19311 2677
rect 19363 2625 19375 2677
rect 19299 2573 19375 2625
rect 19299 2521 19311 2573
rect 19363 2521 19375 2573
rect 19299 2509 19375 2521
rect 19619 2677 19695 2689
rect 19619 2625 19631 2677
rect 19683 2625 19695 2677
rect 19619 2573 19695 2625
rect 19619 2521 19631 2573
rect 19683 2521 19695 2573
rect 19619 2509 19695 2521
rect 19779 2679 19855 2689
rect 19779 2623 19789 2679
rect 19845 2623 19855 2679
rect 19779 2575 19855 2623
rect 19779 2519 19789 2575
rect 19845 2519 19855 2575
rect 19779 2509 19855 2519
rect 18579 2348 18655 2358
rect 18579 2292 18589 2348
rect 18645 2292 18655 2348
rect 18579 2282 18655 2292
rect 18819 2137 18895 2147
rect 18819 2081 18829 2137
rect 18885 2081 18895 2137
rect 18819 2033 18895 2081
rect 18819 1977 18829 2033
rect 18885 1977 18895 2033
rect 18819 1967 18895 1977
rect 18989 1753 19045 2509
rect 19309 1753 19365 2509
rect 19459 2137 19535 2147
rect 19459 2081 19469 2137
rect 19525 2081 19535 2137
rect 19459 2033 19535 2081
rect 19459 1977 19469 2033
rect 19525 1977 19535 2033
rect 19459 1967 19535 1977
rect 19629 1753 19685 2509
rect 20962 1847 21246 2913
rect 20962 1791 20972 1847
rect 21028 1791 21076 1847
rect 21132 1791 21180 1847
rect 21236 1791 21246 1847
rect 18499 1743 18575 1753
rect 18499 1687 18509 1743
rect 18565 1687 18575 1743
rect 18499 1639 18575 1687
rect 18499 1583 18509 1639
rect 18565 1583 18575 1639
rect 18499 1573 18575 1583
rect 18659 1741 18735 1753
rect 18659 1689 18671 1741
rect 18723 1689 18735 1741
rect 18659 1637 18735 1689
rect 18659 1585 18671 1637
rect 18723 1585 18735 1637
rect 18659 1573 18735 1585
rect 18979 1741 19055 1753
rect 18979 1689 18991 1741
rect 19043 1689 19055 1741
rect 18979 1637 19055 1689
rect 18979 1585 18991 1637
rect 19043 1585 19055 1637
rect 18979 1573 19055 1585
rect 19139 1743 19215 1753
rect 19139 1687 19149 1743
rect 19205 1687 19215 1743
rect 19139 1639 19215 1687
rect 19139 1583 19149 1639
rect 19205 1583 19215 1639
rect 19139 1573 19215 1583
rect 19299 1741 19375 1753
rect 19299 1689 19311 1741
rect 19363 1689 19375 1741
rect 19299 1637 19375 1689
rect 19299 1585 19311 1637
rect 19363 1585 19375 1637
rect 19299 1573 19375 1585
rect 19619 1741 19695 1753
rect 19619 1689 19631 1741
rect 19683 1689 19695 1741
rect 19619 1637 19695 1689
rect 19619 1585 19631 1637
rect 19683 1585 19695 1637
rect 19619 1573 19695 1585
rect 19779 1743 19855 1753
rect 19779 1687 19789 1743
rect 19845 1687 19855 1743
rect 19779 1639 19855 1687
rect 19779 1583 19789 1639
rect 19845 1583 19855 1639
rect 19779 1573 19855 1583
rect 20962 1743 21246 1791
rect 20962 1687 20972 1743
rect 21028 1687 21076 1743
rect 21132 1687 21180 1743
rect 21236 1687 21246 1743
rect 20962 1639 21246 1687
rect 20962 1583 20972 1639
rect 21028 1583 21076 1639
rect 21132 1583 21180 1639
rect 21236 1583 21246 1639
rect 18819 1201 18895 1211
rect 18819 1145 18829 1201
rect 18885 1145 18895 1201
rect 18819 1097 18895 1145
rect 18819 1041 18829 1097
rect 18885 1041 18895 1097
rect 18819 1031 18895 1041
rect 18499 807 18575 817
rect 18499 751 18509 807
rect 18565 751 18575 807
rect 18499 703 18575 751
rect 18499 647 18509 703
rect 18565 647 18575 703
rect 18499 637 18575 647
rect 17355 420 17365 476
rect 17421 420 17431 476
rect 14660 -1322 14736 -1312
rect 14660 -1378 14670 -1322
rect 14726 -1378 14736 -1322
rect 14660 -1426 14736 -1378
rect 14660 -1482 14670 -1426
rect 14726 -1482 14736 -1426
rect 14660 -1492 14736 -1482
rect 15300 -1322 15376 -1312
rect 15300 -1378 15310 -1322
rect 15366 -1378 15376 -1322
rect 15300 -1426 15376 -1378
rect 15300 -1482 15310 -1426
rect 15366 -1482 15376 -1426
rect 15300 -1492 15376 -1482
rect 15940 -1322 16016 -1312
rect 15940 -1378 15950 -1322
rect 16006 -1378 16016 -1322
rect 15940 -1426 16016 -1378
rect 15940 -1482 15950 -1426
rect 16006 -1482 16016 -1426
rect 15940 -1492 16016 -1482
rect 16879 -1322 17059 -1312
rect 16879 -1378 16889 -1322
rect 16945 -1378 16993 -1322
rect 17049 -1378 17059 -1322
rect 16879 -1426 17059 -1378
rect 16879 -1482 16889 -1426
rect 16945 -1482 16993 -1426
rect 17049 -1482 17059 -1426
rect 17355 -1396 17431 420
rect 18579 476 18655 486
rect 18579 420 18589 476
rect 18645 420 18655 476
rect 18579 410 18655 420
rect 18819 265 18895 275
rect 18819 209 18829 265
rect 18885 209 18895 265
rect 18819 161 18895 209
rect 18819 105 18829 161
rect 18885 105 18895 161
rect 18819 95 18895 105
rect 18989 -119 19045 1573
rect 19139 807 19215 817
rect 19139 751 19149 807
rect 19205 751 19215 807
rect 19139 703 19215 751
rect 19139 647 19149 703
rect 19205 647 19215 703
rect 19139 637 19215 647
rect 19309 -119 19365 1573
rect 19459 1201 19535 1211
rect 19459 1145 19469 1201
rect 19525 1145 19535 1201
rect 19459 1097 19535 1145
rect 19459 1041 19469 1097
rect 19525 1041 19535 1097
rect 19459 1031 19535 1041
rect 19459 265 19535 275
rect 19459 209 19469 265
rect 19525 209 19535 265
rect 19459 161 19535 209
rect 19459 105 19469 161
rect 19525 105 19535 161
rect 19459 95 19535 105
rect 19629 -119 19685 1573
rect 20962 911 21246 1583
rect 20962 855 20972 911
rect 21028 855 21076 911
rect 21132 855 21180 911
rect 21236 855 21246 911
rect 19779 807 19855 817
rect 19779 751 19789 807
rect 19845 751 19855 807
rect 19779 703 19855 751
rect 19779 647 19789 703
rect 19845 647 19855 703
rect 19779 637 19855 647
rect 20962 807 21246 855
rect 20962 751 20972 807
rect 21028 751 21076 807
rect 21132 751 21180 807
rect 21236 751 21246 807
rect 20962 703 21246 751
rect 20962 647 20972 703
rect 21028 647 21076 703
rect 21132 647 21180 703
rect 21236 647 21246 703
rect 20962 369 21246 647
rect 20962 313 20972 369
rect 21028 313 21076 369
rect 21132 313 21180 369
rect 21236 313 21246 369
rect 20962 265 21246 313
rect 20962 209 20972 265
rect 21028 209 21076 265
rect 21132 209 21180 265
rect 21236 209 21246 265
rect 20962 161 21246 209
rect 20962 105 20972 161
rect 21028 105 21076 161
rect 21132 105 21180 161
rect 21236 105 21246 161
rect 18499 -129 18575 -119
rect 18499 -185 18509 -129
rect 18565 -185 18575 -129
rect 18499 -233 18575 -185
rect 18499 -289 18509 -233
rect 18565 -289 18575 -233
rect 18499 -299 18575 -289
rect 18659 -131 18735 -119
rect 18659 -183 18671 -131
rect 18723 -183 18735 -131
rect 18659 -235 18735 -183
rect 18659 -287 18671 -235
rect 18723 -287 18735 -235
rect 18659 -299 18735 -287
rect 18979 -131 19055 -119
rect 18979 -183 18991 -131
rect 19043 -183 19055 -131
rect 18979 -235 19055 -183
rect 18979 -287 18991 -235
rect 19043 -287 19055 -235
rect 18979 -299 19055 -287
rect 19139 -129 19215 -119
rect 19139 -185 19149 -129
rect 19205 -185 19215 -129
rect 19139 -233 19215 -185
rect 19139 -289 19149 -233
rect 19205 -289 19215 -233
rect 19139 -299 19215 -289
rect 19299 -131 19375 -119
rect 19299 -183 19311 -131
rect 19363 -183 19375 -131
rect 19299 -235 19375 -183
rect 19299 -287 19311 -235
rect 19363 -287 19375 -235
rect 19299 -299 19375 -287
rect 19619 -131 19695 -119
rect 19619 -183 19631 -131
rect 19683 -183 19695 -131
rect 19619 -235 19695 -183
rect 19619 -287 19631 -235
rect 19683 -287 19695 -235
rect 19619 -299 19695 -287
rect 19779 -129 19855 -119
rect 19779 -185 19789 -129
rect 19845 -185 19855 -129
rect 19779 -233 19855 -185
rect 19779 -289 19789 -233
rect 19845 -289 19855 -233
rect 19779 -299 19855 -289
rect 18579 -460 18655 -450
rect 18579 -516 18589 -460
rect 18645 -516 18655 -460
rect 18579 -526 18655 -516
rect 18819 -671 18895 -661
rect 18819 -727 18829 -671
rect 18885 -727 18895 -671
rect 18819 -775 18895 -727
rect 18819 -831 18829 -775
rect 18885 -831 18895 -775
rect 18819 -841 18895 -831
rect 18989 -1055 19045 -299
rect 19309 -1055 19365 -299
rect 19459 -671 19535 -661
rect 19459 -727 19469 -671
rect 19525 -727 19535 -671
rect 19459 -775 19535 -727
rect 19459 -831 19469 -775
rect 19525 -831 19535 -775
rect 19459 -841 19535 -831
rect 19629 -1055 19685 -299
rect 20962 -961 21246 105
rect 21611 2783 21895 3849
rect 23971 4009 24047 4019
rect 23971 3953 23981 4009
rect 24037 3953 24047 4009
rect 23971 3905 24047 3953
rect 23971 3849 23981 3905
rect 24037 3849 24047 3905
rect 23971 3839 24047 3849
rect 24611 4009 24687 4019
rect 24611 3953 24621 4009
rect 24677 3953 24687 4009
rect 24611 3905 24687 3953
rect 24611 3849 24621 3905
rect 24677 3849 24687 3905
rect 24611 3839 24687 3849
rect 21611 2727 21621 2783
rect 21677 2727 21725 2783
rect 21781 2727 21829 2783
rect 21885 2727 21895 2783
rect 21611 2679 21895 2727
rect 21611 2623 21621 2679
rect 21677 2623 21725 2679
rect 21781 2623 21829 2679
rect 21885 2623 21895 2679
rect 21611 2575 21895 2623
rect 21611 2519 21621 2575
rect 21677 2519 21725 2575
rect 21781 2519 21829 2575
rect 21885 2519 21895 2575
rect 21611 2241 21895 2519
rect 21611 2185 21621 2241
rect 21677 2185 21725 2241
rect 21781 2185 21829 2241
rect 21885 2185 21895 2241
rect 21611 2137 21895 2185
rect 21611 2081 21621 2137
rect 21677 2081 21725 2137
rect 21781 2081 21829 2137
rect 21885 2081 21895 2137
rect 21611 2033 21895 2081
rect 21611 1977 21621 2033
rect 21677 1977 21725 2033
rect 21781 1977 21829 2033
rect 21885 1977 21895 2033
rect 21611 1305 21895 1977
rect 21611 1249 21621 1305
rect 21677 1249 21725 1305
rect 21781 1249 21829 1305
rect 21885 1249 21895 1305
rect 21611 1201 21895 1249
rect 21611 1145 21621 1201
rect 21677 1145 21725 1201
rect 21781 1145 21829 1201
rect 21885 1145 21895 1201
rect 21611 1097 21895 1145
rect 21611 1041 21621 1097
rect 21677 1041 21725 1097
rect 21781 1041 21829 1097
rect 21885 1041 21895 1097
rect 21611 -25 21895 1041
rect 21611 -81 21621 -25
rect 21677 -81 21725 -25
rect 21781 -81 21829 -25
rect 21885 -81 21895 -25
rect 21611 -129 21895 -81
rect 21611 -185 21621 -129
rect 21677 -185 21725 -129
rect 21781 -185 21829 -129
rect 21885 -185 21895 -129
rect 21611 -233 21895 -185
rect 21611 -289 21621 -233
rect 21677 -289 21725 -233
rect 21781 -289 21829 -233
rect 21885 -289 21895 -233
rect 21611 -567 21895 -289
rect 21611 -623 21621 -567
rect 21677 -623 21725 -567
rect 21781 -623 21829 -567
rect 21885 -623 21895 -567
rect 21611 -671 21895 -623
rect 21611 -727 21621 -671
rect 21677 -727 21725 -671
rect 21781 -727 21829 -671
rect 21885 -727 21895 -671
rect 21611 -775 21895 -727
rect 21611 -831 21621 -775
rect 21677 -831 21725 -775
rect 21781 -831 21829 -775
rect 21885 -831 21895 -775
rect 21611 -841 21895 -831
rect 22260 3719 22544 3729
rect 22260 3663 22270 3719
rect 22326 3663 22374 3719
rect 22430 3663 22478 3719
rect 22534 3663 22544 3719
rect 22260 3615 22544 3663
rect 22260 3559 22270 3615
rect 22326 3559 22374 3615
rect 22430 3559 22478 3615
rect 22534 3559 22544 3615
rect 22260 3511 22544 3559
rect 22260 3455 22270 3511
rect 22326 3455 22374 3511
rect 22430 3455 22478 3511
rect 22534 3455 22544 3511
rect 22260 3177 22544 3455
rect 23651 3615 23727 3625
rect 23651 3559 23661 3615
rect 23717 3559 23727 3615
rect 23651 3511 23727 3559
rect 23651 3455 23661 3511
rect 23717 3455 23727 3511
rect 23651 3445 23727 3455
rect 23811 3613 23887 3625
rect 23811 3561 23823 3613
rect 23875 3561 23887 3613
rect 23811 3509 23887 3561
rect 23811 3457 23823 3509
rect 23875 3457 23887 3509
rect 23811 3445 23887 3457
rect 24131 3613 24207 3625
rect 24131 3561 24143 3613
rect 24195 3561 24207 3613
rect 24131 3509 24207 3561
rect 24131 3457 24143 3509
rect 24195 3457 24207 3509
rect 24131 3445 24207 3457
rect 24291 3615 24367 3625
rect 24291 3559 24301 3615
rect 24357 3559 24367 3615
rect 24291 3511 24367 3559
rect 24291 3455 24301 3511
rect 24357 3455 24367 3511
rect 24291 3445 24367 3455
rect 24451 3613 24527 3625
rect 24451 3561 24463 3613
rect 24515 3561 24527 3613
rect 24451 3509 24527 3561
rect 24451 3457 24463 3509
rect 24515 3457 24527 3509
rect 24451 3445 24527 3457
rect 24771 3613 24847 3625
rect 24771 3561 24783 3613
rect 24835 3561 24847 3613
rect 24771 3509 24847 3561
rect 24771 3457 24783 3509
rect 24835 3457 24847 3509
rect 24771 3445 24847 3457
rect 24931 3615 25007 3625
rect 24931 3559 24941 3615
rect 24997 3559 25007 3615
rect 24931 3511 25007 3559
rect 24931 3455 24941 3511
rect 24997 3455 25007 3511
rect 24931 3445 25007 3455
rect 22260 3121 22270 3177
rect 22326 3121 22374 3177
rect 22430 3121 22478 3177
rect 22534 3121 22544 3177
rect 22260 3073 22544 3121
rect 22260 3017 22270 3073
rect 22326 3017 22374 3073
rect 22430 3017 22478 3073
rect 22534 3017 22544 3073
rect 22260 2969 22544 3017
rect 22260 2913 22270 2969
rect 22326 2913 22374 2969
rect 22430 2913 22478 2969
rect 22534 2913 22544 2969
rect 22260 1847 22544 2913
rect 23821 2689 23877 3445
rect 23971 3073 24047 3083
rect 23971 3017 23981 3073
rect 24037 3017 24047 3073
rect 23971 2969 24047 3017
rect 23971 2913 23981 2969
rect 24037 2913 24047 2969
rect 23971 2903 24047 2913
rect 24141 2689 24197 3445
rect 24461 2689 24517 3445
rect 24851 3284 24927 3294
rect 24851 3228 24861 3284
rect 24917 3228 24927 3284
rect 24851 3218 24927 3228
rect 26075 3284 26151 3294
rect 26075 3228 26085 3284
rect 26141 3228 26151 3284
rect 24611 3073 24687 3083
rect 24611 3017 24621 3073
rect 24677 3017 24687 3073
rect 24611 2969 24687 3017
rect 24611 2913 24621 2969
rect 24677 2913 24687 2969
rect 24611 2903 24687 2913
rect 23651 2679 23727 2689
rect 23651 2623 23661 2679
rect 23717 2623 23727 2679
rect 23651 2575 23727 2623
rect 23651 2519 23661 2575
rect 23717 2519 23727 2575
rect 23651 2509 23727 2519
rect 23811 2677 23887 2689
rect 23811 2625 23823 2677
rect 23875 2625 23887 2677
rect 23811 2573 23887 2625
rect 23811 2521 23823 2573
rect 23875 2521 23887 2573
rect 23811 2509 23887 2521
rect 24131 2677 24207 2689
rect 24131 2625 24143 2677
rect 24195 2625 24207 2677
rect 24131 2573 24207 2625
rect 24131 2521 24143 2573
rect 24195 2521 24207 2573
rect 24131 2509 24207 2521
rect 24291 2679 24367 2689
rect 24291 2623 24301 2679
rect 24357 2623 24367 2679
rect 24291 2575 24367 2623
rect 24291 2519 24301 2575
rect 24357 2519 24367 2575
rect 24291 2509 24367 2519
rect 24451 2677 24527 2689
rect 24451 2625 24463 2677
rect 24515 2625 24527 2677
rect 24451 2573 24527 2625
rect 24451 2521 24463 2573
rect 24515 2521 24527 2573
rect 24451 2509 24527 2521
rect 24771 2677 24847 2689
rect 24771 2625 24783 2677
rect 24835 2625 24847 2677
rect 24771 2573 24847 2625
rect 24771 2521 24783 2573
rect 24835 2521 24847 2573
rect 24771 2509 24847 2521
rect 24931 2679 25007 2689
rect 24931 2623 24941 2679
rect 24997 2623 25007 2679
rect 24931 2575 25007 2623
rect 24931 2519 24941 2575
rect 24997 2519 25007 2575
rect 24931 2509 25007 2519
rect 22260 1791 22270 1847
rect 22326 1791 22374 1847
rect 22430 1791 22478 1847
rect 22534 1791 22544 1847
rect 22260 1743 22544 1791
rect 23821 1753 23877 2509
rect 23971 2137 24047 2147
rect 23971 2081 23981 2137
rect 24037 2081 24047 2137
rect 23971 2033 24047 2081
rect 23971 1977 23981 2033
rect 24037 1977 24047 2033
rect 23971 1967 24047 1977
rect 24141 1753 24197 2509
rect 24461 1753 24517 2509
rect 24851 2348 24927 2358
rect 24851 2292 24861 2348
rect 24917 2292 24927 2348
rect 24851 2282 24927 2292
rect 24611 2137 24687 2147
rect 24611 2081 24621 2137
rect 24677 2081 24687 2137
rect 24611 2033 24687 2081
rect 24611 1977 24621 2033
rect 24677 1977 24687 2033
rect 24611 1967 24687 1977
rect 22260 1687 22270 1743
rect 22326 1687 22374 1743
rect 22430 1687 22478 1743
rect 22534 1687 22544 1743
rect 22260 1639 22544 1687
rect 22260 1583 22270 1639
rect 22326 1583 22374 1639
rect 22430 1583 22478 1639
rect 22534 1583 22544 1639
rect 22260 911 22544 1583
rect 23651 1743 23727 1753
rect 23651 1687 23661 1743
rect 23717 1687 23727 1743
rect 23651 1639 23727 1687
rect 23651 1583 23661 1639
rect 23717 1583 23727 1639
rect 23651 1573 23727 1583
rect 23811 1741 23887 1753
rect 23811 1689 23823 1741
rect 23875 1689 23887 1741
rect 23811 1637 23887 1689
rect 23811 1585 23823 1637
rect 23875 1585 23887 1637
rect 23811 1573 23887 1585
rect 24131 1741 24207 1753
rect 24131 1689 24143 1741
rect 24195 1689 24207 1741
rect 24131 1637 24207 1689
rect 24131 1585 24143 1637
rect 24195 1585 24207 1637
rect 24131 1573 24207 1585
rect 24291 1743 24367 1753
rect 24291 1687 24301 1743
rect 24357 1687 24367 1743
rect 24291 1639 24367 1687
rect 24291 1583 24301 1639
rect 24357 1583 24367 1639
rect 24291 1573 24367 1583
rect 24451 1741 24527 1753
rect 24451 1689 24463 1741
rect 24515 1689 24527 1741
rect 24451 1637 24527 1689
rect 24451 1585 24463 1637
rect 24515 1585 24527 1637
rect 24451 1573 24527 1585
rect 24771 1741 24847 1753
rect 24771 1689 24783 1741
rect 24835 1689 24847 1741
rect 24771 1637 24847 1689
rect 24771 1585 24783 1637
rect 24835 1585 24847 1637
rect 24771 1573 24847 1585
rect 24931 1743 25007 1753
rect 24931 1687 24941 1743
rect 24997 1687 25007 1743
rect 24931 1639 25007 1687
rect 24931 1583 24941 1639
rect 24997 1583 25007 1639
rect 24931 1573 25007 1583
rect 22260 855 22270 911
rect 22326 855 22374 911
rect 22430 855 22478 911
rect 22534 855 22544 911
rect 22260 807 22544 855
rect 22260 751 22270 807
rect 22326 751 22374 807
rect 22430 751 22478 807
rect 22534 751 22544 807
rect 22260 703 22544 751
rect 22260 647 22270 703
rect 22326 647 22374 703
rect 22430 647 22478 703
rect 22534 647 22544 703
rect 22260 369 22544 647
rect 23651 807 23727 817
rect 23651 751 23661 807
rect 23717 751 23727 807
rect 23651 703 23727 751
rect 23651 647 23661 703
rect 23717 647 23727 703
rect 23651 637 23727 647
rect 22260 313 22270 369
rect 22326 313 22374 369
rect 22430 313 22478 369
rect 22534 313 22544 369
rect 22260 265 22544 313
rect 22260 209 22270 265
rect 22326 209 22374 265
rect 22430 209 22478 265
rect 22534 209 22544 265
rect 22260 161 22544 209
rect 22260 105 22270 161
rect 22326 105 22374 161
rect 22430 105 22478 161
rect 22534 105 22544 161
rect 20962 -1017 20972 -961
rect 21028 -1017 21076 -961
rect 21132 -1017 21180 -961
rect 21236 -1017 21246 -961
rect 18499 -1065 18575 -1055
rect 18499 -1121 18509 -1065
rect 18565 -1121 18575 -1065
rect 18499 -1169 18575 -1121
rect 18499 -1225 18509 -1169
rect 18565 -1225 18575 -1169
rect 18499 -1235 18575 -1225
rect 18659 -1067 18735 -1055
rect 18659 -1119 18671 -1067
rect 18723 -1119 18735 -1067
rect 18659 -1171 18735 -1119
rect 18659 -1223 18671 -1171
rect 18723 -1223 18735 -1171
rect 18659 -1235 18735 -1223
rect 18979 -1067 19055 -1055
rect 18979 -1119 18991 -1067
rect 19043 -1119 19055 -1067
rect 18979 -1171 19055 -1119
rect 18979 -1223 18991 -1171
rect 19043 -1223 19055 -1171
rect 18979 -1235 19055 -1223
rect 19139 -1065 19215 -1055
rect 19139 -1121 19149 -1065
rect 19205 -1121 19215 -1065
rect 19139 -1169 19215 -1121
rect 19139 -1225 19149 -1169
rect 19205 -1225 19215 -1169
rect 19139 -1235 19215 -1225
rect 19299 -1067 19375 -1055
rect 19299 -1119 19311 -1067
rect 19363 -1119 19375 -1067
rect 19299 -1171 19375 -1119
rect 19299 -1223 19311 -1171
rect 19363 -1223 19375 -1171
rect 19299 -1235 19375 -1223
rect 19619 -1067 19695 -1055
rect 19619 -1119 19631 -1067
rect 19683 -1119 19695 -1067
rect 19619 -1171 19695 -1119
rect 19619 -1223 19631 -1171
rect 19683 -1223 19695 -1171
rect 19619 -1235 19695 -1223
rect 19779 -1065 19855 -1055
rect 19779 -1121 19789 -1065
rect 19845 -1121 19855 -1065
rect 19779 -1169 19855 -1121
rect 19779 -1225 19789 -1169
rect 19845 -1225 19855 -1169
rect 19779 -1235 19855 -1225
rect 20962 -1065 21246 -1017
rect 20962 -1121 20972 -1065
rect 21028 -1121 21076 -1065
rect 21132 -1121 21180 -1065
rect 21236 -1121 21246 -1065
rect 20962 -1169 21246 -1121
rect 20962 -1225 20972 -1169
rect 21028 -1225 21076 -1169
rect 21132 -1225 21180 -1169
rect 21236 -1225 21246 -1169
rect 20962 -1235 21246 -1225
rect 22260 -961 22544 105
rect 23821 -119 23877 1573
rect 23971 1201 24047 1211
rect 23971 1145 23981 1201
rect 24037 1145 24047 1201
rect 23971 1097 24047 1145
rect 23971 1041 23981 1097
rect 24037 1041 24047 1097
rect 23971 1031 24047 1041
rect 23971 265 24047 275
rect 23971 209 23981 265
rect 24037 209 24047 265
rect 23971 161 24047 209
rect 23971 105 23981 161
rect 24037 105 24047 161
rect 23971 95 24047 105
rect 24141 -119 24197 1573
rect 24291 807 24367 817
rect 24291 751 24301 807
rect 24357 751 24367 807
rect 24291 703 24367 751
rect 24291 647 24301 703
rect 24357 647 24367 703
rect 24291 637 24367 647
rect 24461 -119 24517 1573
rect 24611 1201 24687 1211
rect 24611 1145 24621 1201
rect 24677 1145 24687 1201
rect 24611 1097 24687 1145
rect 24611 1041 24621 1097
rect 24677 1041 24687 1097
rect 24611 1031 24687 1041
rect 24931 807 25007 817
rect 24931 751 24941 807
rect 24997 751 25007 807
rect 24931 703 25007 751
rect 24931 647 24941 703
rect 24997 647 25007 703
rect 24931 637 25007 647
rect 24851 476 24927 486
rect 24851 420 24861 476
rect 24917 420 24927 476
rect 24851 410 24927 420
rect 26075 476 26151 3228
rect 26075 420 26085 476
rect 26141 420 26151 476
rect 24611 265 24687 275
rect 24611 209 24621 265
rect 24677 209 24687 265
rect 24611 161 24687 209
rect 24611 105 24621 161
rect 24677 105 24687 161
rect 24611 95 24687 105
rect 23651 -129 23727 -119
rect 23651 -185 23661 -129
rect 23717 -185 23727 -129
rect 23651 -233 23727 -185
rect 23651 -289 23661 -233
rect 23717 -289 23727 -233
rect 23651 -299 23727 -289
rect 23811 -131 23887 -119
rect 23811 -183 23823 -131
rect 23875 -183 23887 -131
rect 23811 -235 23887 -183
rect 23811 -287 23823 -235
rect 23875 -287 23887 -235
rect 23811 -299 23887 -287
rect 24131 -131 24207 -119
rect 24131 -183 24143 -131
rect 24195 -183 24207 -131
rect 24131 -235 24207 -183
rect 24131 -287 24143 -235
rect 24195 -287 24207 -235
rect 24131 -299 24207 -287
rect 24291 -129 24367 -119
rect 24291 -185 24301 -129
rect 24357 -185 24367 -129
rect 24291 -233 24367 -185
rect 24291 -289 24301 -233
rect 24357 -289 24367 -233
rect 24291 -299 24367 -289
rect 24451 -131 24527 -119
rect 24451 -183 24463 -131
rect 24515 -183 24527 -131
rect 24451 -235 24527 -183
rect 24451 -287 24463 -235
rect 24515 -287 24527 -235
rect 24451 -299 24527 -287
rect 24771 -131 24847 -119
rect 24771 -183 24783 -131
rect 24835 -183 24847 -131
rect 24771 -235 24847 -183
rect 24771 -287 24783 -235
rect 24835 -287 24847 -235
rect 24771 -299 24847 -287
rect 24931 -129 25007 -119
rect 24931 -185 24941 -129
rect 24997 -185 25007 -129
rect 24931 -233 25007 -185
rect 24931 -289 24941 -233
rect 24997 -289 25007 -233
rect 24931 -299 25007 -289
rect 22260 -1017 22270 -961
rect 22326 -1017 22374 -961
rect 22430 -1017 22478 -961
rect 22534 -1017 22544 -961
rect 22260 -1065 22544 -1017
rect 23821 -1055 23877 -299
rect 23971 -671 24047 -661
rect 23971 -727 23981 -671
rect 24037 -727 24047 -671
rect 23971 -775 24047 -727
rect 23971 -831 23981 -775
rect 24037 -831 24047 -775
rect 23971 -841 24047 -831
rect 24141 -1055 24197 -299
rect 24461 -1055 24517 -299
rect 24851 -460 24927 -450
rect 24851 -516 24861 -460
rect 24917 -516 24927 -460
rect 24851 -526 24927 -516
rect 24611 -671 24687 -661
rect 24611 -727 24621 -671
rect 24677 -727 24687 -671
rect 24611 -775 24687 -727
rect 24611 -831 24621 -775
rect 24677 -831 24687 -775
rect 24611 -841 24687 -831
rect 22260 -1121 22270 -1065
rect 22326 -1121 22374 -1065
rect 22430 -1121 22478 -1065
rect 22534 -1121 22544 -1065
rect 22260 -1169 22544 -1121
rect 22260 -1225 22270 -1169
rect 22326 -1225 22374 -1169
rect 22430 -1225 22478 -1169
rect 22534 -1225 22544 -1169
rect 22260 -1235 22544 -1225
rect 23651 -1065 23727 -1055
rect 23651 -1121 23661 -1065
rect 23717 -1121 23727 -1065
rect 23651 -1169 23727 -1121
rect 23651 -1225 23661 -1169
rect 23717 -1225 23727 -1169
rect 23651 -1235 23727 -1225
rect 23811 -1067 23887 -1055
rect 23811 -1119 23823 -1067
rect 23875 -1119 23887 -1067
rect 23811 -1171 23887 -1119
rect 23811 -1223 23823 -1171
rect 23875 -1223 23887 -1171
rect 23811 -1235 23887 -1223
rect 24131 -1067 24207 -1055
rect 24131 -1119 24143 -1067
rect 24195 -1119 24207 -1067
rect 24131 -1171 24207 -1119
rect 24131 -1223 24143 -1171
rect 24195 -1223 24207 -1171
rect 24131 -1235 24207 -1223
rect 24291 -1065 24367 -1055
rect 24291 -1121 24301 -1065
rect 24357 -1121 24367 -1065
rect 24291 -1169 24367 -1121
rect 24291 -1225 24301 -1169
rect 24357 -1225 24367 -1169
rect 24291 -1235 24367 -1225
rect 24451 -1067 24527 -1055
rect 24451 -1119 24463 -1067
rect 24515 -1119 24527 -1067
rect 24451 -1171 24527 -1119
rect 24451 -1223 24463 -1171
rect 24515 -1223 24527 -1171
rect 24451 -1235 24527 -1223
rect 24771 -1067 24847 -1055
rect 24771 -1119 24783 -1067
rect 24835 -1119 24847 -1067
rect 24771 -1171 24847 -1119
rect 24771 -1223 24783 -1171
rect 24835 -1223 24847 -1171
rect 24771 -1235 24847 -1223
rect 24931 -1065 25007 -1055
rect 24931 -1121 24941 -1065
rect 24997 -1121 25007 -1065
rect 24931 -1169 25007 -1121
rect 24931 -1225 24941 -1169
rect 24997 -1225 25007 -1169
rect 24931 -1235 25007 -1225
rect 17355 -1452 17365 -1396
rect 17421 -1452 17431 -1396
rect 17355 -1462 17431 -1452
rect 18739 -1396 18815 -1386
rect 18739 -1452 18749 -1396
rect 18805 -1452 18815 -1396
rect 18739 -1462 18815 -1452
rect 19379 -1396 19455 -1386
rect 19379 -1452 19389 -1396
rect 19445 -1452 19455 -1396
rect 19379 -1462 19455 -1452
rect 24051 -1396 24127 -1386
rect 24051 -1452 24061 -1396
rect 24117 -1452 24127 -1396
rect 24051 -1462 24127 -1452
rect 24691 -1396 24767 -1386
rect 24691 -1452 24701 -1396
rect 24757 -1452 24767 -1396
rect 24691 -1462 24767 -1452
rect 26075 -1396 26151 420
rect 26276 2348 26351 4194
rect 27700 4250 27776 4260
rect 27700 4194 27710 4250
rect 27766 4194 27776 4250
rect 27700 4184 27776 4194
rect 30732 4113 31016 6288
rect 30732 4057 30742 4113
rect 30798 4057 30846 4113
rect 30902 4057 30950 4113
rect 31006 4057 31016 4113
rect 27940 4009 28016 4019
rect 27940 3953 27950 4009
rect 28006 3953 28016 4009
rect 27940 3905 28016 3953
rect 27940 3849 27950 3905
rect 28006 3849 28016 3905
rect 27940 3839 28016 3849
rect 28580 4009 28656 4019
rect 28580 3953 28590 4009
rect 28646 3953 28656 4009
rect 28580 3905 28656 3953
rect 28580 3849 28590 3905
rect 28646 3849 28656 3905
rect 28580 3839 28656 3849
rect 30732 4009 31016 4057
rect 30732 3953 30742 4009
rect 30798 3953 30846 4009
rect 30902 3953 30950 4009
rect 31006 3953 31016 4009
rect 30732 3905 31016 3953
rect 30732 3849 30742 3905
rect 30798 3849 30846 3905
rect 30902 3849 30950 3905
rect 31006 3849 31016 3905
rect 30083 3719 30367 3729
rect 30083 3663 30093 3719
rect 30149 3663 30197 3719
rect 30253 3663 30301 3719
rect 30357 3663 30367 3719
rect 27620 3615 27696 3625
rect 27620 3559 27630 3615
rect 27686 3559 27696 3615
rect 27620 3511 27696 3559
rect 27620 3455 27630 3511
rect 27686 3455 27696 3511
rect 27620 3445 27696 3455
rect 27780 3613 27856 3625
rect 27780 3561 27792 3613
rect 27844 3561 27856 3613
rect 27780 3509 27856 3561
rect 27780 3457 27792 3509
rect 27844 3457 27856 3509
rect 27780 3445 27856 3457
rect 28100 3613 28176 3625
rect 28100 3561 28112 3613
rect 28164 3561 28176 3613
rect 28100 3509 28176 3561
rect 28100 3457 28112 3509
rect 28164 3457 28176 3509
rect 28100 3445 28176 3457
rect 28260 3615 28336 3625
rect 28260 3559 28270 3615
rect 28326 3559 28336 3615
rect 28260 3511 28336 3559
rect 28260 3455 28270 3511
rect 28326 3455 28336 3511
rect 28260 3445 28336 3455
rect 28420 3613 28496 3625
rect 28420 3561 28432 3613
rect 28484 3561 28496 3613
rect 28420 3509 28496 3561
rect 28420 3457 28432 3509
rect 28484 3457 28496 3509
rect 28420 3445 28496 3457
rect 28740 3613 28816 3625
rect 28740 3561 28752 3613
rect 28804 3561 28816 3613
rect 28740 3509 28816 3561
rect 28740 3457 28752 3509
rect 28804 3457 28816 3509
rect 28740 3445 28816 3457
rect 28900 3615 28976 3625
rect 28900 3559 28910 3615
rect 28966 3559 28976 3615
rect 28900 3511 28976 3559
rect 28900 3455 28910 3511
rect 28966 3455 28976 3511
rect 28900 3445 28976 3455
rect 30083 3615 30367 3663
rect 30083 3559 30093 3615
rect 30149 3559 30197 3615
rect 30253 3559 30301 3615
rect 30357 3559 30367 3615
rect 30083 3511 30367 3559
rect 30083 3455 30093 3511
rect 30149 3455 30197 3511
rect 30253 3455 30301 3511
rect 30357 3455 30367 3511
rect 26276 2292 26285 2348
rect 26342 2292 26351 2348
rect 26276 -460 26351 2292
rect 26276 -516 26285 -460
rect 26342 -516 26351 -460
rect 26276 -526 26351 -516
rect 26476 3284 26552 3294
rect 26476 3228 26486 3284
rect 26542 3228 26552 3284
rect 26476 476 26552 3228
rect 27700 3284 27776 3294
rect 27700 3228 27710 3284
rect 27766 3228 27776 3284
rect 27700 3218 27776 3228
rect 27940 3073 28016 3083
rect 27940 3017 27950 3073
rect 28006 3017 28016 3073
rect 27940 2969 28016 3017
rect 27940 2913 27950 2969
rect 28006 2913 28016 2969
rect 27940 2903 28016 2913
rect 28110 2689 28166 3445
rect 28430 2689 28486 3445
rect 28580 3073 28656 3083
rect 28580 3017 28590 3073
rect 28646 3017 28656 3073
rect 28580 2969 28656 3017
rect 28580 2913 28590 2969
rect 28646 2913 28656 2969
rect 28580 2903 28656 2913
rect 28750 2689 28806 3445
rect 30083 3177 30367 3455
rect 30083 3121 30093 3177
rect 30149 3121 30197 3177
rect 30253 3121 30301 3177
rect 30357 3121 30367 3177
rect 30083 3073 30367 3121
rect 30083 3017 30093 3073
rect 30149 3017 30197 3073
rect 30253 3017 30301 3073
rect 30357 3017 30367 3073
rect 30083 2969 30367 3017
rect 30083 2913 30093 2969
rect 30149 2913 30197 2969
rect 30253 2913 30301 2969
rect 30357 2913 30367 2969
rect 27620 2679 27696 2689
rect 27620 2623 27630 2679
rect 27686 2623 27696 2679
rect 27620 2575 27696 2623
rect 27620 2519 27630 2575
rect 27686 2519 27696 2575
rect 27620 2509 27696 2519
rect 27780 2677 27856 2689
rect 27780 2625 27792 2677
rect 27844 2625 27856 2677
rect 27780 2573 27856 2625
rect 27780 2521 27792 2573
rect 27844 2521 27856 2573
rect 27780 2509 27856 2521
rect 28100 2677 28176 2689
rect 28100 2625 28112 2677
rect 28164 2625 28176 2677
rect 28100 2573 28176 2625
rect 28100 2521 28112 2573
rect 28164 2521 28176 2573
rect 28100 2509 28176 2521
rect 28260 2679 28336 2689
rect 28260 2623 28270 2679
rect 28326 2623 28336 2679
rect 28260 2575 28336 2623
rect 28260 2519 28270 2575
rect 28326 2519 28336 2575
rect 28260 2509 28336 2519
rect 28420 2677 28496 2689
rect 28420 2625 28432 2677
rect 28484 2625 28496 2677
rect 28420 2573 28496 2625
rect 28420 2521 28432 2573
rect 28484 2521 28496 2573
rect 28420 2509 28496 2521
rect 28740 2677 28816 2689
rect 28740 2625 28752 2677
rect 28804 2625 28816 2677
rect 28740 2573 28816 2625
rect 28740 2521 28752 2573
rect 28804 2521 28816 2573
rect 28740 2509 28816 2521
rect 28900 2679 28976 2689
rect 28900 2623 28910 2679
rect 28966 2623 28976 2679
rect 28900 2575 28976 2623
rect 28900 2519 28910 2575
rect 28966 2519 28976 2575
rect 28900 2509 28976 2519
rect 27700 2348 27776 2358
rect 27700 2292 27710 2348
rect 27766 2292 27776 2348
rect 27700 2282 27776 2292
rect 27940 2137 28016 2147
rect 27940 2081 27950 2137
rect 28006 2081 28016 2137
rect 27940 2033 28016 2081
rect 27940 1977 27950 2033
rect 28006 1977 28016 2033
rect 27940 1967 28016 1977
rect 28110 1753 28166 2509
rect 28430 1753 28486 2509
rect 28580 2137 28656 2147
rect 28580 2081 28590 2137
rect 28646 2081 28656 2137
rect 28580 2033 28656 2081
rect 28580 1977 28590 2033
rect 28646 1977 28656 2033
rect 28580 1967 28656 1977
rect 28750 1753 28806 2509
rect 30083 1847 30367 2913
rect 30083 1791 30093 1847
rect 30149 1791 30197 1847
rect 30253 1791 30301 1847
rect 30357 1791 30367 1847
rect 27620 1743 27696 1753
rect 27620 1687 27630 1743
rect 27686 1687 27696 1743
rect 27620 1639 27696 1687
rect 27620 1583 27630 1639
rect 27686 1583 27696 1639
rect 27620 1573 27696 1583
rect 27780 1741 27856 1753
rect 27780 1689 27792 1741
rect 27844 1689 27856 1741
rect 27780 1637 27856 1689
rect 27780 1585 27792 1637
rect 27844 1585 27856 1637
rect 27780 1573 27856 1585
rect 28100 1741 28176 1753
rect 28100 1689 28112 1741
rect 28164 1689 28176 1741
rect 28100 1637 28176 1689
rect 28100 1585 28112 1637
rect 28164 1585 28176 1637
rect 28100 1573 28176 1585
rect 28260 1743 28336 1753
rect 28260 1687 28270 1743
rect 28326 1687 28336 1743
rect 28260 1639 28336 1687
rect 28260 1583 28270 1639
rect 28326 1583 28336 1639
rect 28260 1573 28336 1583
rect 28420 1741 28496 1753
rect 28420 1689 28432 1741
rect 28484 1689 28496 1741
rect 28420 1637 28496 1689
rect 28420 1585 28432 1637
rect 28484 1585 28496 1637
rect 28420 1573 28496 1585
rect 28740 1741 28816 1753
rect 28740 1689 28752 1741
rect 28804 1689 28816 1741
rect 28740 1637 28816 1689
rect 28740 1585 28752 1637
rect 28804 1585 28816 1637
rect 28740 1573 28816 1585
rect 28900 1743 28976 1753
rect 28900 1687 28910 1743
rect 28966 1687 28976 1743
rect 28900 1639 28976 1687
rect 28900 1583 28910 1639
rect 28966 1583 28976 1639
rect 28900 1573 28976 1583
rect 30083 1743 30367 1791
rect 30083 1687 30093 1743
rect 30149 1687 30197 1743
rect 30253 1687 30301 1743
rect 30357 1687 30367 1743
rect 30083 1639 30367 1687
rect 30083 1583 30093 1639
rect 30149 1583 30197 1639
rect 30253 1583 30301 1639
rect 30357 1583 30367 1639
rect 27940 1201 28016 1211
rect 27940 1145 27950 1201
rect 28006 1145 28016 1201
rect 27940 1097 28016 1145
rect 27940 1041 27950 1097
rect 28006 1041 28016 1097
rect 27940 1031 28016 1041
rect 27620 807 27696 817
rect 27620 751 27630 807
rect 27686 751 27696 807
rect 27620 703 27696 751
rect 27620 647 27630 703
rect 27686 647 27696 703
rect 27620 637 27696 647
rect 26476 420 26486 476
rect 26542 420 26552 476
rect 26075 -1452 26085 -1396
rect 26141 -1452 26151 -1396
rect 26075 -1462 26151 -1452
rect 26476 -1396 26552 420
rect 27700 476 27776 486
rect 27700 420 27710 476
rect 27766 420 27776 476
rect 27700 410 27776 420
rect 27940 265 28016 275
rect 27940 209 27950 265
rect 28006 209 28016 265
rect 27940 161 28016 209
rect 27940 105 27950 161
rect 28006 105 28016 161
rect 27940 95 28016 105
rect 28110 -119 28166 1573
rect 28260 807 28336 817
rect 28260 751 28270 807
rect 28326 751 28336 807
rect 28260 703 28336 751
rect 28260 647 28270 703
rect 28326 647 28336 703
rect 28260 637 28336 647
rect 28430 -119 28486 1573
rect 28580 1201 28656 1211
rect 28580 1145 28590 1201
rect 28646 1145 28656 1201
rect 28580 1097 28656 1145
rect 28580 1041 28590 1097
rect 28646 1041 28656 1097
rect 28580 1031 28656 1041
rect 28580 265 28656 275
rect 28580 209 28590 265
rect 28646 209 28656 265
rect 28580 161 28656 209
rect 28580 105 28590 161
rect 28646 105 28656 161
rect 28580 95 28656 105
rect 28750 -119 28806 1573
rect 30083 911 30367 1583
rect 30083 855 30093 911
rect 30149 855 30197 911
rect 30253 855 30301 911
rect 30357 855 30367 911
rect 28900 807 28976 817
rect 28900 751 28910 807
rect 28966 751 28976 807
rect 28900 703 28976 751
rect 28900 647 28910 703
rect 28966 647 28976 703
rect 28900 637 28976 647
rect 30083 807 30367 855
rect 30083 751 30093 807
rect 30149 751 30197 807
rect 30253 751 30301 807
rect 30357 751 30367 807
rect 30083 703 30367 751
rect 30083 647 30093 703
rect 30149 647 30197 703
rect 30253 647 30301 703
rect 30357 647 30367 703
rect 30083 369 30367 647
rect 30083 313 30093 369
rect 30149 313 30197 369
rect 30253 313 30301 369
rect 30357 313 30367 369
rect 30083 265 30367 313
rect 30083 209 30093 265
rect 30149 209 30197 265
rect 30253 209 30301 265
rect 30357 209 30367 265
rect 30083 161 30367 209
rect 30083 105 30093 161
rect 30149 105 30197 161
rect 30253 105 30301 161
rect 30357 105 30367 161
rect 27620 -129 27696 -119
rect 27620 -185 27630 -129
rect 27686 -185 27696 -129
rect 27620 -233 27696 -185
rect 27620 -289 27630 -233
rect 27686 -289 27696 -233
rect 27620 -299 27696 -289
rect 27780 -131 27856 -119
rect 27780 -183 27792 -131
rect 27844 -183 27856 -131
rect 27780 -235 27856 -183
rect 27780 -287 27792 -235
rect 27844 -287 27856 -235
rect 27780 -299 27856 -287
rect 28100 -131 28176 -119
rect 28100 -183 28112 -131
rect 28164 -183 28176 -131
rect 28100 -235 28176 -183
rect 28100 -287 28112 -235
rect 28164 -287 28176 -235
rect 28100 -299 28176 -287
rect 28260 -129 28336 -119
rect 28260 -185 28270 -129
rect 28326 -185 28336 -129
rect 28260 -233 28336 -185
rect 28260 -289 28270 -233
rect 28326 -289 28336 -233
rect 28260 -299 28336 -289
rect 28420 -131 28496 -119
rect 28420 -183 28432 -131
rect 28484 -183 28496 -131
rect 28420 -235 28496 -183
rect 28420 -287 28432 -235
rect 28484 -287 28496 -235
rect 28420 -299 28496 -287
rect 28740 -131 28816 -119
rect 28740 -183 28752 -131
rect 28804 -183 28816 -131
rect 28740 -235 28816 -183
rect 28740 -287 28752 -235
rect 28804 -287 28816 -235
rect 28740 -299 28816 -287
rect 28900 -129 28976 -119
rect 28900 -185 28910 -129
rect 28966 -185 28976 -129
rect 28900 -233 28976 -185
rect 28900 -289 28910 -233
rect 28966 -289 28976 -233
rect 28900 -299 28976 -289
rect 27700 -460 27776 -450
rect 27700 -516 27710 -460
rect 27766 -516 27776 -460
rect 27700 -526 27776 -516
rect 27940 -671 28016 -661
rect 27940 -727 27950 -671
rect 28006 -727 28016 -671
rect 27940 -775 28016 -727
rect 27940 -831 27950 -775
rect 28006 -831 28016 -775
rect 27940 -841 28016 -831
rect 28110 -1055 28166 -299
rect 28430 -1055 28486 -299
rect 28580 -671 28656 -661
rect 28580 -727 28590 -671
rect 28646 -727 28656 -671
rect 28580 -775 28656 -727
rect 28580 -831 28590 -775
rect 28646 -831 28656 -775
rect 28580 -841 28656 -831
rect 28750 -1055 28806 -299
rect 30083 -961 30367 105
rect 30083 -1017 30093 -961
rect 30149 -1017 30197 -961
rect 30253 -1017 30301 -961
rect 30357 -1017 30367 -961
rect 27620 -1065 27696 -1055
rect 27620 -1121 27630 -1065
rect 27686 -1121 27696 -1065
rect 27620 -1169 27696 -1121
rect 27620 -1225 27630 -1169
rect 27686 -1225 27696 -1169
rect 27620 -1235 27696 -1225
rect 27780 -1067 27856 -1055
rect 27780 -1119 27792 -1067
rect 27844 -1119 27856 -1067
rect 27780 -1171 27856 -1119
rect 27780 -1223 27792 -1171
rect 27844 -1223 27856 -1171
rect 27780 -1235 27856 -1223
rect 28100 -1067 28176 -1055
rect 28100 -1119 28112 -1067
rect 28164 -1119 28176 -1067
rect 28100 -1171 28176 -1119
rect 28100 -1223 28112 -1171
rect 28164 -1223 28176 -1171
rect 28100 -1235 28176 -1223
rect 28260 -1065 28336 -1055
rect 28260 -1121 28270 -1065
rect 28326 -1121 28336 -1065
rect 28260 -1169 28336 -1121
rect 28260 -1225 28270 -1169
rect 28326 -1225 28336 -1169
rect 28260 -1235 28336 -1225
rect 28420 -1067 28496 -1055
rect 28420 -1119 28432 -1067
rect 28484 -1119 28496 -1067
rect 28420 -1171 28496 -1119
rect 28420 -1223 28432 -1171
rect 28484 -1223 28496 -1171
rect 28420 -1235 28496 -1223
rect 28740 -1067 28816 -1055
rect 28740 -1119 28752 -1067
rect 28804 -1119 28816 -1067
rect 28740 -1171 28816 -1119
rect 28740 -1223 28752 -1171
rect 28804 -1223 28816 -1171
rect 28740 -1235 28816 -1223
rect 28900 -1065 28976 -1055
rect 28900 -1121 28910 -1065
rect 28966 -1121 28976 -1065
rect 28900 -1169 28976 -1121
rect 28900 -1225 28910 -1169
rect 28966 -1225 28976 -1169
rect 28900 -1235 28976 -1225
rect 30083 -1065 30367 -1017
rect 30083 -1121 30093 -1065
rect 30149 -1121 30197 -1065
rect 30253 -1121 30301 -1065
rect 30357 -1121 30367 -1065
rect 30083 -1169 30367 -1121
rect 30083 -1225 30093 -1169
rect 30149 -1225 30197 -1169
rect 30253 -1225 30301 -1169
rect 30357 -1225 30367 -1169
rect 30083 -1235 30367 -1225
rect 30732 2783 31016 3849
rect 31646 5962 31930 5974
rect 31646 5910 31658 5962
rect 31710 5910 31762 5962
rect 31814 5910 31866 5962
rect 31918 5910 31930 5962
rect 31646 5858 31930 5910
rect 31646 5806 31658 5858
rect 31710 5806 31762 5858
rect 31814 5806 31866 5858
rect 31918 5806 31930 5858
rect 31646 5754 31930 5806
rect 31646 5702 31658 5754
rect 31710 5702 31762 5754
rect 31814 5702 31866 5754
rect 31918 5702 31930 5754
rect 31646 5690 31930 5702
rect 31646 3729 31924 5690
rect 30732 2727 30742 2783
rect 30798 2727 30846 2783
rect 30902 2727 30950 2783
rect 31006 2727 31016 2783
rect 30732 2679 31016 2727
rect 30732 2623 30742 2679
rect 30798 2623 30846 2679
rect 30902 2623 30950 2679
rect 31006 2623 31016 2679
rect 31640 3719 31924 3729
rect 31640 3663 31650 3719
rect 31706 3663 31754 3719
rect 31810 3663 31858 3719
rect 31914 3663 31924 3719
rect 31640 3615 31924 3663
rect 34092 3893 34376 3903
rect 34092 3837 34102 3893
rect 34158 3837 34206 3893
rect 34262 3837 34310 3893
rect 34366 3837 34376 3893
rect 34092 3789 34376 3837
rect 34092 3733 34102 3789
rect 34158 3733 34206 3789
rect 34262 3733 34310 3789
rect 34366 3733 34376 3789
rect 34092 3685 34376 3733
rect 34092 3629 34102 3685
rect 34158 3629 34206 3685
rect 34262 3629 34310 3685
rect 34366 3629 34376 3685
rect 34092 3619 34376 3629
rect 38228 3893 38512 3903
rect 38228 3837 38238 3893
rect 38294 3837 38342 3893
rect 38398 3837 38446 3893
rect 38502 3837 38512 3893
rect 38228 3789 38512 3837
rect 38228 3733 38238 3789
rect 38294 3733 38342 3789
rect 38398 3733 38446 3789
rect 38502 3733 38512 3789
rect 38228 3685 38512 3733
rect 38228 3629 38238 3685
rect 38294 3629 38342 3685
rect 38398 3629 38446 3685
rect 38502 3629 38512 3685
rect 38228 3619 38512 3629
rect 43788 3893 44072 3903
rect 43788 3837 43798 3893
rect 43854 3837 43902 3893
rect 43958 3837 44006 3893
rect 44062 3837 44072 3893
rect 43788 3789 44072 3837
rect 43788 3733 43798 3789
rect 43854 3733 43902 3789
rect 43958 3733 44006 3789
rect 44062 3733 44072 3789
rect 43788 3685 44072 3733
rect 43788 3629 43798 3685
rect 43854 3629 43902 3685
rect 43958 3629 44006 3685
rect 44062 3629 44072 3685
rect 43788 3619 44072 3629
rect 47924 3893 48208 3903
rect 47924 3837 47934 3893
rect 47990 3837 48038 3893
rect 48094 3837 48142 3893
rect 48198 3837 48208 3893
rect 47924 3789 48208 3837
rect 47924 3733 47934 3789
rect 47990 3733 48038 3789
rect 48094 3733 48142 3789
rect 48198 3733 48208 3789
rect 47924 3685 48208 3733
rect 47924 3629 47934 3685
rect 47990 3629 48038 3685
rect 48094 3629 48142 3685
rect 48198 3629 48208 3685
rect 47924 3619 48208 3629
rect 53484 3893 53768 3903
rect 53484 3837 53494 3893
rect 53550 3837 53598 3893
rect 53654 3837 53702 3893
rect 53758 3837 53768 3893
rect 53484 3789 53768 3837
rect 53484 3733 53494 3789
rect 53550 3733 53598 3789
rect 53654 3733 53702 3789
rect 53758 3733 53768 3789
rect 53484 3685 53768 3733
rect 53484 3629 53494 3685
rect 53550 3629 53598 3685
rect 53654 3629 53702 3685
rect 53758 3629 53768 3685
rect 53484 3619 53768 3629
rect 57620 3893 57904 3903
rect 57620 3837 57630 3893
rect 57686 3837 57734 3893
rect 57790 3837 57838 3893
rect 57894 3837 57904 3893
rect 57620 3789 57904 3837
rect 57620 3733 57630 3789
rect 57686 3733 57734 3789
rect 57790 3733 57838 3789
rect 57894 3733 57904 3789
rect 57620 3685 57904 3733
rect 57620 3629 57630 3685
rect 57686 3629 57734 3685
rect 57790 3629 57838 3685
rect 57894 3629 57904 3685
rect 57620 3619 57904 3629
rect 63180 3893 63464 3903
rect 63180 3837 63190 3893
rect 63246 3837 63294 3893
rect 63350 3837 63398 3893
rect 63454 3837 63464 3893
rect 63180 3789 63464 3837
rect 63180 3733 63190 3789
rect 63246 3733 63294 3789
rect 63350 3733 63398 3789
rect 63454 3733 63464 3789
rect 63180 3685 63464 3733
rect 63180 3629 63190 3685
rect 63246 3629 63294 3685
rect 63350 3629 63398 3685
rect 63454 3629 63464 3685
rect 63180 3619 63464 3629
rect 66428 3893 66712 3903
rect 66428 3837 66438 3893
rect 66494 3837 66542 3893
rect 66598 3837 66646 3893
rect 66702 3837 66712 3893
rect 66428 3789 66712 3837
rect 66428 3733 66438 3789
rect 66494 3733 66542 3789
rect 66598 3733 66646 3789
rect 66702 3733 66712 3789
rect 66428 3685 66712 3733
rect 66428 3629 66438 3685
rect 66494 3629 66542 3685
rect 66598 3629 66646 3685
rect 66702 3629 66712 3685
rect 66428 3619 66712 3629
rect 31640 3559 31650 3615
rect 31706 3559 31754 3615
rect 31810 3559 31858 3615
rect 31914 3559 31924 3615
rect 31640 3511 31924 3559
rect 31640 3455 31650 3511
rect 31706 3455 31754 3511
rect 31810 3455 31858 3511
rect 31914 3455 31924 3511
rect 31640 3177 31924 3455
rect 31640 3121 31650 3177
rect 31706 3121 31754 3177
rect 31810 3121 31858 3177
rect 31914 3121 31924 3177
rect 31640 3073 31924 3121
rect 31640 3017 31650 3073
rect 31706 3017 31754 3073
rect 31810 3017 31858 3073
rect 31914 3017 31924 3073
rect 31640 2969 31924 3017
rect 31640 2913 31650 2969
rect 31706 2913 31754 2969
rect 31810 2913 31858 2969
rect 31914 2913 31924 2969
rect 30732 2575 31016 2623
rect 30732 2519 30742 2575
rect 30798 2519 30846 2575
rect 30902 2519 30950 2575
rect 31006 2519 31016 2575
rect 30732 2241 31016 2519
rect 30732 2185 30742 2241
rect 30798 2185 30846 2241
rect 30902 2185 30950 2241
rect 31006 2185 31016 2241
rect 30732 2137 31016 2185
rect 30732 2081 30742 2137
rect 30798 2081 30846 2137
rect 30902 2081 30950 2137
rect 31006 2081 31016 2137
rect 30732 2033 31016 2081
rect 30732 1977 30742 2033
rect 30798 1977 30846 2033
rect 30902 1977 30950 2033
rect 31006 1977 31016 2033
rect 30732 1305 31016 1977
rect 30732 1249 30742 1305
rect 30798 1249 30846 1305
rect 30902 1249 30950 1305
rect 31006 1249 31016 1305
rect 30732 1201 31016 1249
rect 30732 1145 30742 1201
rect 30798 1145 30846 1201
rect 30902 1145 30950 1201
rect 31006 1145 31016 1201
rect 30732 1097 31016 1145
rect 30732 1041 30742 1097
rect 30798 1041 30846 1097
rect 30902 1041 30950 1097
rect 31006 1041 31016 1097
rect 30732 -25 31016 1041
rect 30732 -81 30742 -25
rect 30798 -81 30846 -25
rect 30902 -81 30950 -25
rect 31006 -81 31016 -25
rect 30732 -129 31016 -81
rect 30732 -185 30742 -129
rect 30798 -185 30846 -129
rect 30902 -185 30950 -129
rect 31006 -185 31016 -129
rect 30732 -233 31016 -185
rect 30732 -289 30742 -233
rect 30798 -289 30846 -233
rect 30902 -289 30950 -233
rect 31006 -289 31016 -233
rect 30732 -567 31016 -289
rect 30732 -623 30742 -567
rect 30798 -623 30846 -567
rect 30902 -623 30950 -567
rect 31006 -623 31016 -567
rect 30732 -671 31016 -623
rect 30732 -727 30742 -671
rect 30798 -727 30846 -671
rect 30902 -727 30950 -671
rect 31006 -727 31016 -671
rect 30732 -775 31016 -727
rect 30732 -831 30742 -775
rect 30798 -831 30846 -775
rect 30902 -831 30950 -775
rect 31006 -831 31016 -775
rect 26476 -1452 26486 -1396
rect 26542 -1452 26552 -1396
rect 26476 -1462 26552 -1452
rect 27860 -1396 27936 -1386
rect 27860 -1452 27870 -1396
rect 27926 -1452 27936 -1396
rect 27860 -1462 27936 -1452
rect 16879 -1492 17059 -1482
rect 16633 -2719 16917 -2709
rect 16633 -2775 16643 -2719
rect 16699 -2775 16747 -2719
rect 16803 -2775 16851 -2719
rect 16907 -2775 16917 -2719
rect 16633 -2823 16917 -2775
rect 16633 -2879 16643 -2823
rect 16699 -2879 16747 -2823
rect 16803 -2879 16851 -2823
rect 16907 -2879 16917 -2823
rect 16633 -2927 16917 -2879
rect 16633 -2983 16643 -2927
rect 16699 -2983 16747 -2927
rect 16803 -2983 16851 -2927
rect 16907 -2983 16917 -2927
rect 16633 -2993 16917 -2983
rect 29802 -2719 30294 -2709
rect 29802 -2775 29812 -2719
rect 29868 -2775 29916 -2719
rect 29972 -2775 30020 -2719
rect 30076 -2775 30124 -2719
rect 30180 -2775 30228 -2719
rect 30284 -2775 30294 -2719
rect 29802 -2823 30294 -2775
rect 29802 -2879 29812 -2823
rect 29868 -2879 29916 -2823
rect 29972 -2879 30020 -2823
rect 30076 -2879 30124 -2823
rect 30180 -2879 30228 -2823
rect 30284 -2879 30294 -2823
rect 29802 -2927 30294 -2879
rect 29802 -2983 29812 -2927
rect 29868 -2983 29916 -2927
rect 29972 -2983 30020 -2927
rect 30076 -2983 30124 -2927
rect 30180 -2983 30228 -2927
rect 30284 -2983 30294 -2927
rect 17070 -3061 17354 -3051
rect 17070 -3117 17080 -3061
rect 17136 -3117 17184 -3061
rect 17240 -3117 17288 -3061
rect 17344 -3117 17354 -3061
rect 17070 -3165 17354 -3117
rect 17070 -3221 17080 -3165
rect 17136 -3221 17184 -3165
rect 17240 -3221 17288 -3165
rect 17344 -3221 17354 -3165
rect 17070 -3269 17354 -3221
rect 17070 -3325 17080 -3269
rect 17136 -3325 17184 -3269
rect 17240 -3325 17288 -3269
rect 17344 -3325 17354 -3269
rect 17070 -3335 17354 -3325
rect 29242 -3061 29734 -3051
rect 29242 -3117 29252 -3061
rect 29308 -3117 29356 -3061
rect 29412 -3117 29460 -3061
rect 29516 -3117 29564 -3061
rect 29620 -3117 29668 -3061
rect 29724 -3117 29734 -3061
rect 29242 -3165 29734 -3117
rect 29242 -3221 29252 -3165
rect 29308 -3221 29356 -3165
rect 29412 -3221 29460 -3165
rect 29516 -3221 29564 -3165
rect 29620 -3221 29668 -3165
rect 29724 -3221 29734 -3165
rect 29242 -3269 29734 -3221
rect 29242 -3325 29252 -3269
rect 29308 -3325 29356 -3269
rect 29412 -3325 29460 -3269
rect 29516 -3325 29564 -3269
rect 29620 -3325 29668 -3269
rect 29724 -3325 29734 -3269
rect 14200 -3446 14380 -3436
rect 14200 -3502 14210 -3446
rect 14266 -3502 14314 -3446
rect 14370 -3502 14380 -3446
rect 14200 -3550 14380 -3502
rect 14200 -3606 14210 -3550
rect 14266 -3606 14314 -3550
rect 14370 -3606 14380 -3550
rect 14200 -3616 14380 -3606
rect 16848 -3711 17028 -3701
rect 16848 -3767 16858 -3711
rect 16914 -3767 16962 -3711
rect 17018 -3767 17028 -3711
rect 16848 -3815 17028 -3767
rect 16848 -3871 16858 -3815
rect 16914 -3871 16962 -3815
rect 17018 -3871 17028 -3815
rect 16848 -3881 17028 -3871
rect 23634 -3711 23814 -3701
rect 23634 -3767 23644 -3711
rect 23700 -3767 23748 -3711
rect 23804 -3767 23814 -3711
rect 23634 -3815 23814 -3767
rect 23634 -3871 23644 -3815
rect 23700 -3871 23748 -3815
rect 23804 -3871 23814 -3815
rect 23634 -3881 23814 -3871
rect 23644 -4132 23804 -3881
rect 23632 -4144 23812 -4132
rect 23632 -4196 23644 -4144
rect 23696 -4196 23748 -4144
rect 23800 -4196 23812 -4144
rect 20084 -4239 20368 -4227
rect 20084 -4291 20173 -4239
rect 20225 -4291 20277 -4239
rect 20329 -4291 20368 -4239
rect 13726 -4691 14010 -4681
rect 13726 -4747 13736 -4691
rect 13792 -4747 13840 -4691
rect 13896 -4747 13944 -4691
rect 14000 -4747 14010 -4691
rect 13726 -4795 14010 -4747
rect 13726 -4851 13736 -4795
rect 13792 -4851 13840 -4795
rect 13896 -4851 13944 -4795
rect 14000 -4851 14010 -4795
rect 13726 -4899 14010 -4851
rect 13726 -4955 13736 -4899
rect 13792 -4955 13840 -4899
rect 13896 -4955 13944 -4899
rect 14000 -4955 14010 -4899
rect 12614 -6861 12690 -6851
rect 12614 -6917 12624 -6861
rect 12680 -6917 12690 -6861
rect 12614 -6965 12690 -6917
rect 12614 -7021 12624 -6965
rect 12680 -7021 12690 -6965
rect 12614 -7069 12690 -7021
rect 12614 -7125 12624 -7069
rect 12680 -7125 12690 -7069
rect 12614 -7135 12690 -7125
rect 13726 -7322 14010 -4955
rect 14566 -5593 14642 -5583
rect 14566 -5649 14576 -5593
rect 14632 -5649 14642 -5593
rect 14566 -5697 14642 -5649
rect 14566 -5753 14576 -5697
rect 14632 -5753 14642 -5697
rect 14566 -5763 14642 -5753
rect 15174 -5593 15250 -5583
rect 15174 -5649 15184 -5593
rect 15240 -5649 15250 -5593
rect 15174 -5697 15250 -5649
rect 15174 -5753 15184 -5697
rect 15240 -5753 15250 -5697
rect 15174 -5763 15250 -5753
rect 15782 -5593 15858 -5583
rect 15782 -5649 15792 -5593
rect 15848 -5649 15858 -5593
rect 15782 -5697 15858 -5649
rect 15782 -5753 15792 -5697
rect 15848 -5753 15858 -5697
rect 15782 -5763 15858 -5753
rect 15070 -5993 15354 -5983
rect 15070 -6049 15080 -5993
rect 15136 -6049 15184 -5993
rect 15240 -6049 15288 -5993
rect 15344 -6049 15354 -5993
rect 15070 -6097 15354 -6049
rect 15070 -6153 15080 -6097
rect 15136 -6153 15184 -6097
rect 15240 -6153 15288 -6097
rect 15344 -6153 15354 -6097
rect 15070 -6201 15354 -6153
rect 15070 -6257 15080 -6201
rect 15136 -6257 15184 -6201
rect 15240 -6257 15288 -6201
rect 15344 -6257 15354 -6201
rect 12714 -7342 12894 -7330
rect 12714 -7394 12726 -7342
rect 12778 -7394 12830 -7342
rect 12882 -7394 12894 -7342
rect 13726 -7374 13738 -7322
rect 13790 -7374 13842 -7322
rect 13894 -7374 13946 -7322
rect 13998 -7374 14010 -7322
rect 13726 -7386 14010 -7374
rect 14403 -6861 14687 -6851
rect 14403 -6917 14413 -6861
rect 14469 -6917 14517 -6861
rect 14573 -6917 14621 -6861
rect 14677 -6917 14687 -6861
rect 14403 -6965 14687 -6917
rect 14403 -7021 14413 -6965
rect 14469 -7021 14517 -6965
rect 14573 -7021 14621 -6965
rect 14677 -7021 14687 -6965
rect 14403 -7069 14687 -7021
rect 14403 -7125 14413 -7069
rect 14469 -7125 14517 -7069
rect 14573 -7125 14621 -7069
rect 14677 -7125 14687 -7069
rect 12714 -7446 12894 -7394
rect 12714 -7498 12726 -7446
rect 12778 -7498 12830 -7446
rect 12882 -7498 12894 -7446
rect 11532 -8028 11712 -8018
rect 11532 -8084 11542 -8028
rect 11598 -8084 11646 -8028
rect 11702 -8084 11712 -8028
rect 11532 -8132 11712 -8084
rect 11532 -8188 11542 -8132
rect 11598 -8188 11646 -8132
rect 11702 -8188 11712 -8132
rect 11532 -8198 11712 -8188
rect 5134 -8280 5314 -8270
rect 5134 -8336 5144 -8280
rect 5200 -8336 5248 -8280
rect 5304 -8336 5314 -8280
rect 5134 -8384 5314 -8336
rect 5134 -8440 5144 -8384
rect 5200 -8440 5248 -8384
rect 5304 -8440 5314 -8384
rect 5134 -8450 5314 -8440
rect 9827 -8280 10007 -8270
rect 9827 -8336 9837 -8280
rect 9893 -8336 9941 -8280
rect 9997 -8336 10007 -8280
rect 9827 -8384 10007 -8336
rect 9827 -8440 9837 -8384
rect 9893 -8440 9941 -8384
rect 9997 -8440 10007 -8384
rect 9827 -8450 10007 -8440
rect 4658 -8600 4838 -8590
rect 4658 -8656 4668 -8600
rect 4724 -8656 4772 -8600
rect 4828 -8656 4838 -8600
rect 4658 -8704 4838 -8656
rect 4658 -8760 4668 -8704
rect 4724 -8760 4772 -8704
rect 4828 -8760 4838 -8704
rect 4658 -8770 4838 -8760
rect 12714 -8600 12894 -7498
rect 12714 -8656 12724 -8600
rect 12780 -8656 12828 -8600
rect 12884 -8656 12894 -8600
rect 12714 -8704 12894 -8656
rect 14403 -8383 14687 -7125
rect 14403 -8439 14413 -8383
rect 14469 -8439 14517 -8383
rect 14573 -8439 14621 -8383
rect 14677 -8439 14687 -8383
rect 14403 -8487 14687 -8439
rect 14403 -8543 14413 -8487
rect 14469 -8543 14517 -8487
rect 14573 -8543 14621 -8487
rect 14677 -8543 14687 -8487
rect 14403 -8591 14687 -8543
rect 14403 -8647 14413 -8591
rect 14469 -8647 14517 -8591
rect 14573 -8647 14621 -8591
rect 14677 -8647 14687 -8591
rect 14403 -8657 14687 -8647
rect 15070 -6861 15354 -6257
rect 20084 -5993 20368 -4291
rect 23632 -4248 23812 -4196
rect 23632 -4300 23644 -4248
rect 23696 -4300 23748 -4248
rect 23800 -4300 23812 -4248
rect 23632 -4312 23812 -4300
rect 21174 -4691 21250 -4681
rect 21174 -4747 21184 -4691
rect 21240 -4747 21250 -4691
rect 21174 -4795 21250 -4747
rect 21174 -4851 21184 -4795
rect 21240 -4851 21250 -4795
rect 21174 -4899 21250 -4851
rect 21174 -4955 21184 -4899
rect 21240 -4955 21250 -4899
rect 21174 -4965 21250 -4955
rect 26994 -4852 27174 -4840
rect 26994 -4904 27006 -4852
rect 27058 -4904 27110 -4852
rect 27162 -4904 27174 -4852
rect 26994 -4956 27174 -4904
rect 26994 -5008 27006 -4956
rect 27058 -5008 27110 -4956
rect 27162 -5008 27174 -4956
rect 20084 -6049 20094 -5993
rect 20150 -6049 20198 -5993
rect 20254 -6049 20302 -5993
rect 20358 -6049 20368 -5993
rect 20084 -6097 20368 -6049
rect 20084 -6153 20094 -6097
rect 20150 -6153 20198 -6097
rect 20254 -6153 20302 -6097
rect 20358 -6153 20368 -6097
rect 20084 -6201 20368 -6153
rect 20084 -6257 20094 -6201
rect 20150 -6257 20198 -6201
rect 20254 -6257 20302 -6201
rect 20358 -6257 20368 -6201
rect 20084 -6267 20368 -6257
rect 26992 -6220 27174 -5008
rect 26992 -6272 27004 -6220
rect 27056 -6272 27108 -6220
rect 27160 -6222 27174 -6220
rect 29242 -6076 29734 -3325
rect 29802 -4064 30294 -2983
rect 29802 -4116 29814 -4064
rect 29866 -4116 29918 -4064
rect 29970 -4116 30022 -4064
rect 30074 -4116 30126 -4064
rect 30178 -4116 30230 -4064
rect 30282 -4116 30294 -4064
rect 29802 -4168 30294 -4116
rect 29802 -4220 29814 -4168
rect 29866 -4220 29918 -4168
rect 29970 -4220 30022 -4168
rect 30074 -4220 30126 -4168
rect 30178 -4220 30230 -4168
rect 30282 -4220 30294 -4168
rect 29802 -4272 30294 -4220
rect 29802 -4324 29814 -4272
rect 29866 -4324 29918 -4272
rect 29970 -4324 30022 -4272
rect 30074 -4324 30126 -4272
rect 30178 -4324 30230 -4272
rect 30282 -4324 30294 -4272
rect 29802 -4336 30294 -4324
rect 29802 -5018 30294 -5008
rect 29802 -5074 29812 -5018
rect 29868 -5074 29916 -5018
rect 29972 -5074 30020 -5018
rect 30076 -5074 30124 -5018
rect 30180 -5074 30228 -5018
rect 30284 -5074 30294 -5018
rect 29802 -5122 30294 -5074
rect 29802 -5178 29812 -5122
rect 29868 -5178 29916 -5122
rect 29972 -5178 30020 -5122
rect 30076 -5178 30124 -5122
rect 30180 -5178 30228 -5122
rect 30284 -5178 30294 -5122
rect 29802 -5226 30294 -5178
rect 29802 -5282 29812 -5226
rect 29868 -5282 29916 -5226
rect 29972 -5282 30020 -5226
rect 30076 -5282 30124 -5226
rect 30180 -5282 30228 -5226
rect 30284 -5282 30294 -5226
rect 29802 -5330 30294 -5282
rect 29802 -5386 29812 -5330
rect 29868 -5386 29916 -5330
rect 29972 -5386 30020 -5330
rect 30076 -5386 30124 -5330
rect 30180 -5386 30228 -5330
rect 30284 -5386 30294 -5330
rect 29802 -5434 30294 -5386
rect 29802 -5490 29812 -5434
rect 29868 -5490 29916 -5434
rect 29972 -5490 30020 -5434
rect 30076 -5490 30124 -5434
rect 30180 -5490 30228 -5434
rect 30284 -5490 30294 -5434
rect 29802 -5500 30294 -5490
rect 29242 -6128 29254 -6076
rect 29306 -6128 29358 -6076
rect 29410 -6128 29462 -6076
rect 29514 -6128 29566 -6076
rect 29618 -6128 29670 -6076
rect 29722 -6128 29734 -6076
rect 29242 -6180 29734 -6128
rect 27160 -6272 27172 -6222
rect 26992 -6324 27172 -6272
rect 15070 -6917 15080 -6861
rect 15136 -6917 15184 -6861
rect 15240 -6917 15288 -6861
rect 15344 -6917 15354 -6861
rect 15070 -6965 15354 -6917
rect 15070 -7021 15080 -6965
rect 15136 -7021 15184 -6965
rect 15240 -7021 15288 -6965
rect 15344 -7021 15354 -6965
rect 15070 -7069 15354 -7021
rect 15070 -7125 15080 -7069
rect 15136 -7125 15184 -7069
rect 15240 -7125 15288 -7069
rect 15344 -7125 15354 -7069
rect 12714 -8760 12724 -8704
rect 12780 -8760 12828 -8704
rect 12884 -8760 12894 -8704
rect 12714 -8770 12894 -8760
rect 15070 -8885 15354 -7125
rect 15685 -6394 15969 -6372
rect 26992 -6376 27004 -6324
rect 27056 -6376 27108 -6324
rect 27160 -6376 27172 -6324
rect 29242 -6232 29254 -6180
rect 29306 -6232 29358 -6180
rect 29410 -6232 29462 -6180
rect 29514 -6232 29566 -6180
rect 29618 -6232 29670 -6180
rect 29722 -6232 29734 -6180
rect 29242 -6284 29734 -6232
rect 29242 -6336 29254 -6284
rect 29306 -6336 29358 -6284
rect 29410 -6336 29462 -6284
rect 29514 -6336 29566 -6284
rect 29618 -6336 29670 -6284
rect 29722 -6336 29734 -6284
rect 29242 -6348 29734 -6336
rect 26992 -6388 27172 -6376
rect 15685 -6446 15697 -6394
rect 15749 -6446 15801 -6394
rect 15853 -6446 15905 -6394
rect 15957 -6446 15969 -6394
rect 15685 -6498 15969 -6446
rect 15685 -6550 15697 -6498
rect 15749 -6550 15801 -6498
rect 15853 -6550 15905 -6498
rect 15957 -6550 15969 -6498
rect 15685 -6899 15969 -6550
rect 15685 -6955 15695 -6899
rect 15751 -6955 15799 -6899
rect 15855 -6955 15903 -6899
rect 15959 -6955 15969 -6899
rect 15685 -7003 15969 -6955
rect 15685 -7059 15695 -7003
rect 15751 -7059 15799 -7003
rect 15855 -7059 15903 -7003
rect 15959 -7059 15969 -7003
rect 15685 -7107 15969 -7059
rect 15685 -7163 15695 -7107
rect 15751 -7163 15799 -7107
rect 15855 -7163 15903 -7107
rect 15959 -7163 15969 -7107
rect 15685 -7173 15969 -7163
rect 18614 -6899 18690 -6889
rect 18614 -6955 18624 -6899
rect 18680 -6955 18690 -6899
rect 18614 -7003 18690 -6955
rect 18614 -7059 18624 -7003
rect 18680 -7059 18690 -7003
rect 18614 -7107 18690 -7059
rect 18614 -7163 18624 -7107
rect 18680 -7163 18690 -7107
rect 18614 -7173 18690 -7163
rect 18934 -6899 19010 -6889
rect 18934 -6955 18944 -6899
rect 19000 -6955 19010 -6899
rect 18934 -7003 19010 -6955
rect 18934 -7059 18944 -7003
rect 19000 -7059 19010 -7003
rect 18934 -7107 19010 -7059
rect 18934 -7163 18944 -7107
rect 19000 -7163 19010 -7107
rect 18934 -7173 19010 -7163
rect 19254 -6899 19330 -6889
rect 19254 -6955 19264 -6899
rect 19320 -6955 19330 -6899
rect 19254 -7003 19330 -6955
rect 19254 -7059 19264 -7003
rect 19320 -7059 19330 -7003
rect 19254 -7107 19330 -7059
rect 19254 -7163 19264 -7107
rect 19320 -7163 19330 -7107
rect 19254 -7173 19330 -7163
rect 19574 -6899 19650 -6889
rect 19574 -6955 19584 -6899
rect 19640 -6955 19650 -6899
rect 19574 -7003 19650 -6955
rect 19574 -7059 19584 -7003
rect 19640 -7059 19650 -7003
rect 19574 -7107 19650 -7059
rect 19574 -7163 19584 -7107
rect 19640 -7163 19650 -7107
rect 19574 -7173 19650 -7163
rect 19894 -6899 19970 -6889
rect 19894 -6955 19904 -6899
rect 19960 -6955 19970 -6899
rect 19894 -7003 19970 -6955
rect 19894 -7059 19904 -7003
rect 19960 -7059 19970 -7003
rect 19894 -7107 19970 -7059
rect 19894 -7163 19904 -7107
rect 19960 -7163 19970 -7107
rect 19894 -7173 19970 -7163
rect 20214 -6899 20290 -6889
rect 20214 -6955 20224 -6899
rect 20280 -6955 20290 -6899
rect 20214 -7003 20290 -6955
rect 20214 -7059 20224 -7003
rect 20280 -7059 20290 -7003
rect 20214 -7107 20290 -7059
rect 20214 -7163 20224 -7107
rect 20280 -7163 20290 -7107
rect 20214 -7173 20290 -7163
rect 20534 -6899 20610 -6889
rect 20534 -6955 20544 -6899
rect 20600 -6955 20610 -6899
rect 20534 -7003 20610 -6955
rect 20534 -7059 20544 -7003
rect 20600 -7059 20610 -7003
rect 20534 -7107 20610 -7059
rect 20534 -7163 20544 -7107
rect 20600 -7163 20610 -7107
rect 20534 -7173 20610 -7163
rect 29802 -7030 30294 -7020
rect 29802 -7086 29812 -7030
rect 29868 -7086 29916 -7030
rect 29972 -7086 30020 -7030
rect 30076 -7086 30124 -7030
rect 30180 -7086 30228 -7030
rect 30284 -7086 30294 -7030
rect 29802 -7134 30294 -7086
rect 29802 -7190 29812 -7134
rect 29868 -7190 29916 -7134
rect 29972 -7190 30020 -7134
rect 30076 -7190 30124 -7134
rect 30180 -7190 30228 -7134
rect 30284 -7190 30294 -7134
rect 29802 -7238 30294 -7190
rect 21145 -7253 21429 -7241
rect 21145 -7305 21157 -7253
rect 21209 -7305 21261 -7253
rect 21313 -7305 21365 -7253
rect 21417 -7305 21429 -7253
rect 21145 -8383 21429 -7305
rect 29802 -7294 29812 -7238
rect 29868 -7294 29916 -7238
rect 29972 -7294 30020 -7238
rect 30076 -7294 30124 -7238
rect 30180 -7294 30228 -7238
rect 30284 -7294 30294 -7238
rect 21145 -8439 21155 -8383
rect 21211 -8439 21259 -8383
rect 21315 -8439 21363 -8383
rect 21419 -8439 21429 -8383
rect 21145 -8487 21429 -8439
rect 21145 -8543 21155 -8487
rect 21211 -8543 21259 -8487
rect 21315 -8543 21363 -8487
rect 21419 -8543 21429 -8487
rect 21145 -8591 21429 -8543
rect 21145 -8647 21155 -8591
rect 21211 -8647 21259 -8591
rect 21315 -8647 21363 -8591
rect 21419 -8647 21429 -8591
rect 23632 -7352 23812 -7340
rect 23632 -7404 23644 -7352
rect 23696 -7404 23748 -7352
rect 23800 -7404 23812 -7352
rect 23632 -7456 23812 -7404
rect 23632 -7508 23644 -7456
rect 23696 -7508 23748 -7456
rect 23800 -7508 23812 -7456
rect 23632 -8370 23812 -7508
rect 23632 -8426 23642 -8370
rect 23698 -8426 23746 -8370
rect 23802 -8426 23812 -8370
rect 23632 -8474 23812 -8426
rect 23632 -8530 23642 -8474
rect 23698 -8530 23746 -8474
rect 23802 -8530 23812 -8474
rect 23632 -8578 23812 -8530
rect 23632 -8634 23642 -8578
rect 23698 -8634 23746 -8578
rect 23802 -8634 23812 -8578
rect 23632 -8644 23812 -8634
rect 24082 -7352 24262 -7338
rect 24082 -7404 24092 -7352
rect 24144 -7404 24196 -7352
rect 24248 -7404 24262 -7352
rect 24082 -7456 24262 -7404
rect 24082 -7508 24092 -7456
rect 24144 -7508 24196 -7456
rect 24248 -7508 24262 -7456
rect 21145 -8657 21429 -8647
rect 18953 -8771 19258 -8761
rect 18953 -8795 18963 -8771
rect 15070 -8937 15082 -8885
rect 15134 -8937 15186 -8885
rect 15238 -8937 15290 -8885
rect 15342 -8937 15354 -8885
rect 15070 -8989 15354 -8937
rect 15070 -9041 15082 -8989
rect 15134 -9041 15186 -8989
rect 15238 -9041 15290 -8989
rect 15342 -9041 15354 -8989
rect 15070 -9093 15354 -9041
rect 15070 -9145 15082 -9093
rect 15134 -9145 15186 -9093
rect 15238 -9145 15290 -9093
rect 15342 -9145 15354 -9093
rect 15070 -9157 15354 -9145
rect 18952 -8827 18963 -8795
rect 19019 -8827 19067 -8771
rect 19123 -8827 19190 -8771
rect 19246 -8827 19258 -8771
rect 18952 -8875 19258 -8827
rect 18952 -8931 18963 -8875
rect 19019 -8931 19067 -8875
rect 19123 -8931 19190 -8875
rect 19246 -8931 19258 -8875
rect 18952 -8979 19258 -8931
rect 18952 -9035 18963 -8979
rect 19019 -9035 19067 -8979
rect 19123 -9035 19190 -8979
rect 19246 -9035 19258 -8979
rect 18952 -9045 19258 -9035
rect 24082 -8771 24262 -7508
rect 29802 -7342 30294 -7294
rect 29802 -7398 29812 -7342
rect 29868 -7398 29916 -7342
rect 29972 -7398 30020 -7342
rect 30076 -7398 30124 -7342
rect 30180 -7398 30228 -7342
rect 30284 -7398 30294 -7342
rect 29802 -7446 30294 -7398
rect 29802 -7502 29812 -7446
rect 29868 -7502 29916 -7446
rect 29972 -7502 30020 -7446
rect 30076 -7502 30124 -7446
rect 30180 -7502 30228 -7446
rect 30284 -7502 30294 -7446
rect 29802 -7512 30294 -7502
rect 30732 -8370 31016 -831
rect 31260 2613 31544 2623
rect 31260 2557 31270 2613
rect 31326 2557 31374 2613
rect 31430 2557 31478 2613
rect 31534 2557 31544 2613
rect 31260 2509 31544 2557
rect 31260 2453 31270 2509
rect 31326 2453 31374 2509
rect 31430 2453 31478 2509
rect 31534 2453 31544 2509
rect 31260 2405 31544 2453
rect 31260 2349 31270 2405
rect 31326 2349 31374 2405
rect 31430 2349 31478 2405
rect 31534 2349 31544 2405
rect 31260 1159 31544 2349
rect 31260 1103 31270 1159
rect 31326 1103 31374 1159
rect 31430 1103 31478 1159
rect 31534 1103 31544 1159
rect 31260 1055 31544 1103
rect 31260 999 31270 1055
rect 31326 999 31374 1055
rect 31430 999 31478 1055
rect 31534 999 31544 1055
rect 31260 951 31544 999
rect 31260 895 31270 951
rect 31326 895 31374 951
rect 31430 895 31478 951
rect 31534 895 31544 951
rect 31260 99 31544 895
rect 31260 43 31270 99
rect 31326 43 31374 99
rect 31430 43 31478 99
rect 31534 43 31544 99
rect 31260 -5 31544 43
rect 31260 -61 31270 -5
rect 31326 -61 31374 -5
rect 31430 -61 31478 -5
rect 31534 -61 31544 -5
rect 31260 -109 31544 -61
rect 31260 -165 31270 -109
rect 31326 -165 31374 -109
rect 31430 -165 31478 -109
rect 31534 -165 31544 -109
rect 31260 -567 31544 -165
rect 31260 -623 31270 -567
rect 31326 -623 31374 -567
rect 31430 -623 31478 -567
rect 31534 -623 31544 -567
rect 31260 -671 31544 -623
rect 31260 -727 31270 -671
rect 31326 -727 31374 -671
rect 31430 -727 31478 -671
rect 31534 -727 31544 -671
rect 31260 -775 31544 -727
rect 31260 -831 31270 -775
rect 31326 -831 31374 -775
rect 31430 -831 31478 -775
rect 31534 -831 31544 -775
rect 31260 -841 31544 -831
rect 31640 2219 31924 2913
rect 34116 2655 34352 3619
rect 34116 2603 34128 2655
rect 34180 2603 34288 2655
rect 34340 2603 34352 2655
rect 33237 2509 33313 2519
rect 33237 2453 33247 2509
rect 33303 2453 33313 2509
rect 33237 2405 33313 2453
rect 33237 2349 33247 2405
rect 33303 2349 33313 2405
rect 33237 2339 33313 2349
rect 33877 2509 33953 2519
rect 33877 2453 33887 2509
rect 33943 2453 33953 2509
rect 33877 2405 33953 2453
rect 33877 2349 33887 2405
rect 33943 2349 33953 2405
rect 33877 2339 33953 2349
rect 31640 2163 31650 2219
rect 31706 2163 31754 2219
rect 31810 2163 31858 2219
rect 31914 2163 31924 2219
rect 31640 2115 31924 2163
rect 31640 2059 31650 2115
rect 31706 2059 31754 2115
rect 31810 2059 31858 2115
rect 31914 2059 31924 2115
rect 31640 2011 31924 2059
rect 31640 1955 31650 2011
rect 31706 1955 31754 2011
rect 31810 1955 31858 2011
rect 31914 1955 31924 2011
rect 31640 1553 31924 1955
rect 32916 2115 32992 2125
rect 32916 2059 32926 2115
rect 32982 2059 32992 2115
rect 32916 2011 32992 2059
rect 32916 1955 32926 2011
rect 32982 1955 32992 2011
rect 32916 1945 32992 1955
rect 33556 2115 33632 2125
rect 33556 2059 33566 2115
rect 33622 2059 33632 2115
rect 33556 2011 33632 2059
rect 33556 1955 33566 2011
rect 33622 1955 33632 2011
rect 33556 1945 33632 1955
rect 31640 1497 31650 1553
rect 31706 1497 31754 1553
rect 31810 1497 31858 1553
rect 31914 1497 31924 1553
rect 31640 1449 31924 1497
rect 34116 1595 34352 2603
rect 38252 2655 38488 3619
rect 38252 2603 38264 2655
rect 38316 2603 38424 2655
rect 38476 2603 38488 2655
rect 43812 2655 44048 3619
rect 34517 2509 34593 2519
rect 34517 2453 34527 2509
rect 34583 2453 34593 2509
rect 34517 2405 34593 2453
rect 34517 2349 34527 2405
rect 34583 2349 34593 2405
rect 34517 2339 34593 2349
rect 35157 2509 35233 2519
rect 35157 2453 35167 2509
rect 35223 2453 35233 2509
rect 35157 2405 35233 2453
rect 35157 2349 35167 2405
rect 35223 2349 35233 2405
rect 35157 2339 35233 2349
rect 37371 2509 37447 2519
rect 37371 2453 37381 2509
rect 37437 2453 37447 2509
rect 37371 2405 37447 2453
rect 37371 2349 37381 2405
rect 37437 2349 37447 2405
rect 37371 2339 37447 2349
rect 38011 2509 38087 2519
rect 38011 2453 38021 2509
rect 38077 2453 38087 2509
rect 38011 2405 38087 2453
rect 38011 2349 38021 2405
rect 38077 2349 38087 2405
rect 38011 2339 38087 2349
rect 34836 2115 34912 2125
rect 34836 2059 34846 2115
rect 34902 2059 34912 2115
rect 34836 2011 34912 2059
rect 34836 1955 34846 2011
rect 34902 1955 34912 2011
rect 34836 1945 34912 1955
rect 35476 2115 35552 2125
rect 35476 2059 35486 2115
rect 35542 2059 35552 2115
rect 35476 2011 35552 2059
rect 35476 1955 35486 2011
rect 35542 1955 35552 2011
rect 35476 1945 35552 1955
rect 37052 2115 37128 2125
rect 37052 2059 37062 2115
rect 37118 2059 37128 2115
rect 37052 2011 37128 2059
rect 37052 1955 37062 2011
rect 37118 1955 37128 2011
rect 37052 1945 37128 1955
rect 37692 2115 37768 2125
rect 37692 2059 37702 2115
rect 37758 2059 37768 2115
rect 37692 2011 37768 2059
rect 37692 1955 37702 2011
rect 37758 1955 37768 2011
rect 37692 1945 37768 1955
rect 34116 1543 34128 1595
rect 34180 1543 34288 1595
rect 34340 1543 34352 1595
rect 31640 1393 31650 1449
rect 31706 1393 31754 1449
rect 31810 1393 31858 1449
rect 31914 1393 31924 1449
rect 31640 1345 31924 1393
rect 31640 1289 31650 1345
rect 31706 1289 31754 1345
rect 31810 1289 31858 1345
rect 31914 1289 31924 1345
rect 31640 493 31924 1289
rect 33237 1449 33313 1459
rect 33237 1393 33247 1449
rect 33303 1393 33313 1449
rect 33237 1345 33313 1393
rect 33237 1289 33247 1345
rect 33303 1289 33313 1345
rect 33237 1279 33313 1289
rect 33877 1449 33953 1459
rect 33877 1393 33887 1449
rect 33943 1393 33953 1449
rect 33877 1345 33953 1393
rect 33877 1289 33887 1345
rect 33943 1289 33953 1345
rect 33877 1279 33953 1289
rect 32916 1055 32992 1065
rect 32916 999 32926 1055
rect 32982 999 32992 1055
rect 32916 951 32992 999
rect 32916 895 32926 951
rect 32982 895 32992 951
rect 32916 885 32992 895
rect 33556 1055 33632 1065
rect 33556 999 33566 1055
rect 33622 999 33632 1055
rect 33556 951 33632 999
rect 33556 895 33566 951
rect 33622 895 33632 951
rect 33556 885 33632 895
rect 31640 437 31650 493
rect 31706 437 31754 493
rect 31810 437 31858 493
rect 31914 437 31924 493
rect 31640 389 31924 437
rect 34116 535 34352 1543
rect 38252 1595 38488 2603
rect 40987 2613 41271 2623
rect 40987 2557 40997 2613
rect 41053 2557 41101 2613
rect 41157 2557 41205 2613
rect 41261 2557 41271 2613
rect 38651 2509 38727 2519
rect 38651 2453 38661 2509
rect 38717 2453 38727 2509
rect 38651 2405 38727 2453
rect 38651 2349 38661 2405
rect 38717 2349 38727 2405
rect 38651 2339 38727 2349
rect 39291 2509 39367 2519
rect 39291 2453 39301 2509
rect 39357 2453 39367 2509
rect 39291 2405 39367 2453
rect 39291 2349 39301 2405
rect 39357 2349 39367 2405
rect 39291 2339 39367 2349
rect 40987 2509 41271 2557
rect 43812 2603 43824 2655
rect 43876 2603 43984 2655
rect 44036 2603 44048 2655
rect 40987 2453 40997 2509
rect 41053 2453 41101 2509
rect 41157 2453 41205 2509
rect 41261 2453 41271 2509
rect 40987 2405 41271 2453
rect 40987 2349 40997 2405
rect 41053 2349 41101 2405
rect 41157 2349 41205 2405
rect 41261 2349 41271 2405
rect 40626 2219 40910 2229
rect 40626 2163 40636 2219
rect 40692 2163 40740 2219
rect 40796 2163 40844 2219
rect 40900 2163 40910 2219
rect 38972 2115 39048 2125
rect 38972 2059 38982 2115
rect 39038 2059 39048 2115
rect 38972 2011 39048 2059
rect 38972 1955 38982 2011
rect 39038 1955 39048 2011
rect 38972 1945 39048 1955
rect 39612 2115 39688 2125
rect 39612 2059 39622 2115
rect 39678 2059 39688 2115
rect 39612 2011 39688 2059
rect 39612 1955 39622 2011
rect 39678 1955 39688 2011
rect 39612 1945 39688 1955
rect 40626 2115 40910 2163
rect 40626 2059 40636 2115
rect 40692 2059 40740 2115
rect 40796 2059 40844 2115
rect 40900 2059 40910 2115
rect 40626 2011 40910 2059
rect 40626 1955 40636 2011
rect 40692 1955 40740 2011
rect 40796 1955 40844 2011
rect 40900 1955 40910 2011
rect 38252 1543 38264 1595
rect 38316 1543 38424 1595
rect 38476 1543 38488 1595
rect 34517 1449 34593 1459
rect 34517 1393 34527 1449
rect 34583 1393 34593 1449
rect 34517 1345 34593 1393
rect 34517 1289 34527 1345
rect 34583 1289 34593 1345
rect 34517 1279 34593 1289
rect 35157 1449 35233 1459
rect 35157 1393 35167 1449
rect 35223 1393 35233 1449
rect 35157 1345 35233 1393
rect 35157 1289 35167 1345
rect 35223 1289 35233 1345
rect 35157 1279 35233 1289
rect 37371 1449 37447 1459
rect 37371 1393 37381 1449
rect 37437 1393 37447 1449
rect 37371 1345 37447 1393
rect 37371 1289 37381 1345
rect 37437 1289 37447 1345
rect 37371 1279 37447 1289
rect 38011 1449 38087 1459
rect 38011 1393 38021 1449
rect 38077 1393 38087 1449
rect 38011 1345 38087 1393
rect 38011 1289 38021 1345
rect 38077 1289 38087 1345
rect 38011 1279 38087 1289
rect 34836 1055 34912 1065
rect 34836 999 34846 1055
rect 34902 999 34912 1055
rect 34836 951 34912 999
rect 34836 895 34846 951
rect 34902 895 34912 951
rect 34836 885 34912 895
rect 35476 1055 35552 1065
rect 35476 999 35486 1055
rect 35542 999 35552 1055
rect 35476 951 35552 999
rect 35476 895 35486 951
rect 35542 895 35552 951
rect 35476 885 35552 895
rect 37052 1055 37128 1065
rect 37052 999 37062 1055
rect 37118 999 37128 1055
rect 37052 951 37128 999
rect 37052 895 37062 951
rect 37118 895 37128 951
rect 37052 885 37128 895
rect 37692 1055 37768 1065
rect 37692 999 37702 1055
rect 37758 999 37768 1055
rect 37692 951 37768 999
rect 37692 895 37702 951
rect 37758 895 37768 951
rect 37692 885 37768 895
rect 34116 483 34128 535
rect 34180 483 34288 535
rect 34340 483 34352 535
rect 31640 333 31650 389
rect 31706 333 31754 389
rect 31810 333 31858 389
rect 31914 333 31924 389
rect 31640 285 31924 333
rect 31640 229 31650 285
rect 31706 229 31754 285
rect 31810 229 31858 285
rect 31914 229 31924 285
rect 30732 -8426 30742 -8370
rect 30798 -8426 30846 -8370
rect 30902 -8426 30950 -8370
rect 31006 -8426 31016 -8370
rect 30732 -8474 31016 -8426
rect 30732 -8530 30742 -8474
rect 30798 -8530 30846 -8474
rect 30902 -8530 30950 -8474
rect 31006 -8530 31016 -8474
rect 30732 -8578 31016 -8530
rect 30732 -8634 30742 -8578
rect 30798 -8634 30846 -8578
rect 30902 -8634 30950 -8578
rect 31006 -8634 31016 -8578
rect 30732 -8644 31016 -8634
rect 31640 -961 31924 229
rect 33237 389 33313 399
rect 33237 333 33247 389
rect 33303 333 33313 389
rect 33237 285 33313 333
rect 33237 229 33247 285
rect 33303 229 33313 285
rect 33237 219 33313 229
rect 33877 389 33953 399
rect 33877 333 33887 389
rect 33943 333 33953 389
rect 33877 285 33953 333
rect 33877 229 33887 285
rect 33943 229 33953 285
rect 33877 219 33953 229
rect 32916 -5 32992 5
rect 32916 -61 32926 -5
rect 32982 -61 32992 -5
rect 32916 -109 32992 -61
rect 32916 -165 32926 -109
rect 32982 -165 32992 -109
rect 32916 -175 32992 -165
rect 33556 -5 33632 5
rect 33556 -61 33566 -5
rect 33622 -61 33632 -5
rect 33556 -109 33632 -61
rect 33556 -165 33566 -109
rect 33622 -165 33632 -109
rect 33556 -175 33632 -165
rect 34116 -525 34352 483
rect 38252 535 38488 1543
rect 40626 1553 40910 1955
rect 40626 1497 40636 1553
rect 40692 1497 40740 1553
rect 40796 1497 40844 1553
rect 40900 1497 40910 1553
rect 38651 1449 38727 1459
rect 38651 1393 38661 1449
rect 38717 1393 38727 1449
rect 38651 1345 38727 1393
rect 38651 1289 38661 1345
rect 38717 1289 38727 1345
rect 38651 1279 38727 1289
rect 39291 1449 39367 1459
rect 39291 1393 39301 1449
rect 39357 1393 39367 1449
rect 39291 1345 39367 1393
rect 39291 1289 39301 1345
rect 39357 1289 39367 1345
rect 39291 1279 39367 1289
rect 40626 1449 40910 1497
rect 40626 1393 40636 1449
rect 40692 1393 40740 1449
rect 40796 1393 40844 1449
rect 40900 1393 40910 1449
rect 40626 1345 40910 1393
rect 40626 1289 40636 1345
rect 40692 1289 40740 1345
rect 40796 1289 40844 1345
rect 40900 1289 40910 1345
rect 38972 1055 39048 1065
rect 38972 999 38982 1055
rect 39038 999 39048 1055
rect 38972 951 39048 999
rect 38972 895 38982 951
rect 39038 895 39048 951
rect 38972 885 39048 895
rect 39612 1055 39688 1065
rect 39612 999 39622 1055
rect 39678 999 39688 1055
rect 39612 951 39688 999
rect 39612 895 39622 951
rect 39678 895 39688 951
rect 39612 885 39688 895
rect 38252 483 38264 535
rect 38316 483 38424 535
rect 38476 483 38488 535
rect 34517 389 34593 399
rect 34517 333 34527 389
rect 34583 333 34593 389
rect 34517 285 34593 333
rect 34517 229 34527 285
rect 34583 229 34593 285
rect 34517 219 34593 229
rect 35157 389 35233 399
rect 35157 333 35167 389
rect 35223 333 35233 389
rect 35157 285 35233 333
rect 35157 229 35167 285
rect 35223 229 35233 285
rect 35157 219 35233 229
rect 37371 389 37447 399
rect 37371 333 37381 389
rect 37437 333 37447 389
rect 37371 285 37447 333
rect 37371 229 37381 285
rect 37437 229 37447 285
rect 37371 219 37447 229
rect 38011 389 38087 399
rect 38011 333 38021 389
rect 38077 333 38087 389
rect 38011 285 38087 333
rect 38011 229 38021 285
rect 38077 229 38087 285
rect 38011 219 38087 229
rect 34836 -5 34912 5
rect 34836 -61 34846 -5
rect 34902 -61 34912 -5
rect 34836 -109 34912 -61
rect 34836 -165 34846 -109
rect 34902 -165 34912 -109
rect 34836 -175 34912 -165
rect 35476 -5 35552 5
rect 35476 -61 35486 -5
rect 35542 -61 35552 -5
rect 35476 -109 35552 -61
rect 35476 -165 35486 -109
rect 35542 -165 35552 -109
rect 35476 -175 35552 -165
rect 37052 -5 37128 5
rect 37052 -61 37062 -5
rect 37118 -61 37128 -5
rect 37052 -109 37128 -61
rect 37052 -165 37062 -109
rect 37118 -165 37128 -109
rect 37052 -175 37128 -165
rect 37692 -5 37768 5
rect 37692 -61 37702 -5
rect 37758 -61 37768 -5
rect 37692 -109 37768 -61
rect 37692 -165 37702 -109
rect 37758 -165 37768 -109
rect 37692 -175 37768 -165
rect 34116 -577 34128 -525
rect 34180 -577 34288 -525
rect 34340 -577 34352 -525
rect 33237 -671 33313 -661
rect 33237 -727 33247 -671
rect 33303 -727 33313 -671
rect 33237 -775 33313 -727
rect 33237 -831 33247 -775
rect 33303 -831 33313 -775
rect 33237 -841 33313 -831
rect 33877 -671 33953 -661
rect 33877 -727 33887 -671
rect 33943 -727 33953 -671
rect 33877 -775 33953 -727
rect 33877 -831 33887 -775
rect 33943 -831 33953 -775
rect 33877 -841 33953 -831
rect 31640 -1017 31650 -961
rect 31706 -1017 31754 -961
rect 31810 -1017 31858 -961
rect 31914 -1017 31924 -961
rect 31640 -1065 31924 -1017
rect 31640 -1121 31650 -1065
rect 31706 -1121 31754 -1065
rect 31810 -1121 31858 -1065
rect 31914 -1121 31924 -1065
rect 31640 -1169 31924 -1121
rect 31640 -1225 31650 -1169
rect 31706 -1225 31754 -1169
rect 31810 -1225 31858 -1169
rect 31914 -1225 31924 -1169
rect 24082 -8827 24092 -8771
rect 24148 -8827 24196 -8771
rect 24252 -8827 24262 -8771
rect 24082 -8875 24262 -8827
rect 24082 -8931 24092 -8875
rect 24148 -8931 24196 -8875
rect 24252 -8931 24262 -8875
rect 24082 -8979 24262 -8931
rect 24082 -9035 24092 -8979
rect 24148 -9035 24196 -8979
rect 24252 -9035 24262 -8979
rect 24082 -9045 24262 -9035
rect 31640 -8771 31924 -1225
rect 32916 -1065 32992 -1055
rect 32916 -1121 32926 -1065
rect 32982 -1121 32992 -1065
rect 32916 -1169 32992 -1121
rect 32916 -1225 32926 -1169
rect 32982 -1225 32992 -1169
rect 32916 -1235 32992 -1225
rect 33556 -1065 33632 -1055
rect 33556 -1121 33566 -1065
rect 33622 -1121 33632 -1065
rect 33556 -1169 33632 -1121
rect 33556 -1225 33566 -1169
rect 33622 -1225 33632 -1169
rect 33556 -1235 33632 -1225
rect 34116 -5593 34352 -577
rect 38252 -525 38488 483
rect 40626 493 40910 1289
rect 40626 437 40636 493
rect 40692 437 40740 493
rect 40796 437 40844 493
rect 40900 437 40910 493
rect 38651 389 38727 399
rect 38651 333 38661 389
rect 38717 333 38727 389
rect 38651 285 38727 333
rect 38651 229 38661 285
rect 38717 229 38727 285
rect 38651 219 38727 229
rect 39291 389 39367 399
rect 39291 333 39301 389
rect 39357 333 39367 389
rect 39291 285 39367 333
rect 39291 229 39301 285
rect 39357 229 39367 285
rect 39291 219 39367 229
rect 40626 389 40910 437
rect 40626 333 40636 389
rect 40692 333 40740 389
rect 40796 333 40844 389
rect 40900 333 40910 389
rect 40626 285 40910 333
rect 40626 229 40636 285
rect 40692 229 40740 285
rect 40796 229 40844 285
rect 40900 229 40910 285
rect 38972 -5 39048 5
rect 38972 -61 38982 -5
rect 39038 -61 39048 -5
rect 38972 -109 39048 -61
rect 38972 -165 38982 -109
rect 39038 -165 39048 -109
rect 38972 -175 39048 -165
rect 39612 -5 39688 5
rect 39612 -61 39622 -5
rect 39678 -61 39688 -5
rect 39612 -109 39688 -61
rect 39612 -165 39622 -109
rect 39678 -165 39688 -109
rect 39612 -175 39688 -165
rect 38252 -577 38264 -525
rect 38316 -577 38424 -525
rect 38476 -577 38488 -525
rect 38252 -589 38488 -577
rect 34517 -671 34593 -661
rect 34517 -727 34527 -671
rect 34583 -727 34593 -671
rect 34517 -775 34593 -727
rect 34517 -831 34527 -775
rect 34583 -831 34593 -775
rect 34517 -841 34593 -831
rect 35157 -671 35233 -661
rect 35157 -727 35167 -671
rect 35223 -727 35233 -671
rect 35157 -775 35233 -727
rect 35157 -831 35167 -775
rect 35223 -831 35233 -775
rect 35157 -841 35233 -831
rect 37371 -671 37447 -661
rect 37371 -727 37381 -671
rect 37437 -727 37447 -671
rect 37371 -775 37447 -727
rect 37371 -831 37381 -775
rect 37437 -831 37447 -775
rect 37371 -841 37447 -831
rect 38011 -671 38087 -661
rect 38011 -727 38021 -671
rect 38077 -727 38087 -671
rect 38011 -775 38087 -727
rect 38011 -831 38021 -775
rect 38077 -831 38087 -775
rect 38011 -841 38087 -831
rect 38651 -671 38727 -661
rect 38651 -727 38661 -671
rect 38717 -727 38727 -671
rect 38651 -775 38727 -727
rect 38651 -831 38661 -775
rect 38717 -831 38727 -775
rect 38651 -841 38727 -831
rect 39291 -671 39367 -661
rect 39291 -727 39301 -671
rect 39357 -727 39367 -671
rect 39291 -775 39367 -727
rect 39291 -831 39301 -775
rect 39357 -831 39367 -775
rect 39291 -841 39367 -831
rect 40626 -961 40910 229
rect 40987 1159 41271 2349
rect 42933 2509 43009 2519
rect 42933 2453 42943 2509
rect 42999 2453 43009 2509
rect 42933 2405 43009 2453
rect 42933 2349 42943 2405
rect 42999 2349 43009 2405
rect 42933 2339 43009 2349
rect 43573 2509 43649 2519
rect 43573 2453 43583 2509
rect 43639 2453 43649 2509
rect 43573 2405 43649 2453
rect 43573 2349 43583 2405
rect 43639 2349 43649 2405
rect 43573 2339 43649 2349
rect 40987 1103 40997 1159
rect 41053 1103 41101 1159
rect 41157 1103 41205 1159
rect 41261 1103 41271 1159
rect 40987 1055 41271 1103
rect 40987 999 40997 1055
rect 41053 999 41101 1055
rect 41157 999 41205 1055
rect 41261 999 41271 1055
rect 40987 951 41271 999
rect 40987 895 40997 951
rect 41053 895 41101 951
rect 41157 895 41205 951
rect 41261 895 41271 951
rect 40987 99 41271 895
rect 40987 43 40997 99
rect 41053 43 41101 99
rect 41157 43 41205 99
rect 41261 43 41271 99
rect 40987 -5 41271 43
rect 40987 -61 40997 -5
rect 41053 -61 41101 -5
rect 41157 -61 41205 -5
rect 41261 -61 41271 -5
rect 40987 -109 41271 -61
rect 40987 -165 40997 -109
rect 41053 -165 41101 -109
rect 41157 -165 41205 -109
rect 41261 -165 41271 -109
rect 40987 -567 41271 -165
rect 40987 -623 40997 -567
rect 41053 -623 41101 -567
rect 41157 -623 41205 -567
rect 41261 -623 41271 -567
rect 40987 -671 41271 -623
rect 40987 -727 40997 -671
rect 41053 -727 41101 -671
rect 41157 -727 41205 -671
rect 41261 -727 41271 -671
rect 40987 -775 41271 -727
rect 40987 -831 40997 -775
rect 41053 -831 41101 -775
rect 41157 -831 41205 -775
rect 41261 -831 41271 -775
rect 40987 -841 41271 -831
rect 41346 2219 41630 2229
rect 41346 2163 41356 2219
rect 41412 2163 41460 2219
rect 41516 2163 41564 2219
rect 41620 2163 41630 2219
rect 41346 2115 41630 2163
rect 41346 2059 41356 2115
rect 41412 2059 41460 2115
rect 41516 2059 41564 2115
rect 41620 2059 41630 2115
rect 41346 2011 41630 2059
rect 41346 1955 41356 2011
rect 41412 1955 41460 2011
rect 41516 1955 41564 2011
rect 41620 1955 41630 2011
rect 41346 1553 41630 1955
rect 42612 2115 42688 2125
rect 42612 2059 42622 2115
rect 42678 2059 42688 2115
rect 42612 2011 42688 2059
rect 42612 1955 42622 2011
rect 42678 1955 42688 2011
rect 42612 1945 42688 1955
rect 43252 2115 43328 2125
rect 43252 2059 43262 2115
rect 43318 2059 43328 2115
rect 43252 2011 43328 2059
rect 43252 1955 43262 2011
rect 43318 1955 43328 2011
rect 43252 1945 43328 1955
rect 41346 1497 41356 1553
rect 41412 1497 41460 1553
rect 41516 1497 41564 1553
rect 41620 1497 41630 1553
rect 41346 1449 41630 1497
rect 43812 1595 44048 2603
rect 47948 2655 48184 3619
rect 47948 2603 47960 2655
rect 48012 2603 48120 2655
rect 48172 2603 48184 2655
rect 53508 2655 53744 3619
rect 44213 2509 44289 2519
rect 44213 2453 44223 2509
rect 44279 2453 44289 2509
rect 44213 2405 44289 2453
rect 44213 2349 44223 2405
rect 44279 2349 44289 2405
rect 44213 2339 44289 2349
rect 44853 2509 44929 2519
rect 44853 2453 44863 2509
rect 44919 2453 44929 2509
rect 44853 2405 44929 2453
rect 44853 2349 44863 2405
rect 44919 2349 44929 2405
rect 44853 2339 44929 2349
rect 47067 2509 47143 2519
rect 47067 2453 47077 2509
rect 47133 2453 47143 2509
rect 47067 2405 47143 2453
rect 47067 2349 47077 2405
rect 47133 2349 47143 2405
rect 47067 2339 47143 2349
rect 47707 2509 47783 2519
rect 47707 2453 47717 2509
rect 47773 2453 47783 2509
rect 47707 2405 47783 2453
rect 47707 2349 47717 2405
rect 47773 2349 47783 2405
rect 47707 2339 47783 2349
rect 44532 2115 44608 2125
rect 44532 2059 44542 2115
rect 44598 2059 44608 2115
rect 44532 2011 44608 2059
rect 44532 1955 44542 2011
rect 44598 1955 44608 2011
rect 44532 1945 44608 1955
rect 45172 2115 45248 2125
rect 45172 2059 45182 2115
rect 45238 2059 45248 2115
rect 45172 2011 45248 2059
rect 45172 1955 45182 2011
rect 45238 1955 45248 2011
rect 45172 1945 45248 1955
rect 46748 2115 46824 2125
rect 46748 2059 46758 2115
rect 46814 2059 46824 2115
rect 46748 2011 46824 2059
rect 46748 1955 46758 2011
rect 46814 1955 46824 2011
rect 46748 1945 46824 1955
rect 47388 2115 47464 2125
rect 47388 2059 47398 2115
rect 47454 2059 47464 2115
rect 47388 2011 47464 2059
rect 47388 1955 47398 2011
rect 47454 1955 47464 2011
rect 47388 1945 47464 1955
rect 43812 1543 43824 1595
rect 43876 1543 43984 1595
rect 44036 1543 44048 1595
rect 41346 1393 41356 1449
rect 41412 1393 41460 1449
rect 41516 1393 41564 1449
rect 41620 1393 41630 1449
rect 41346 1345 41630 1393
rect 41346 1289 41356 1345
rect 41412 1289 41460 1345
rect 41516 1289 41564 1345
rect 41620 1289 41630 1345
rect 41346 493 41630 1289
rect 42933 1449 43009 1459
rect 42933 1393 42943 1449
rect 42999 1393 43009 1449
rect 42933 1345 43009 1393
rect 42933 1289 42943 1345
rect 42999 1289 43009 1345
rect 42933 1279 43009 1289
rect 43573 1449 43649 1459
rect 43573 1393 43583 1449
rect 43639 1393 43649 1449
rect 43573 1345 43649 1393
rect 43573 1289 43583 1345
rect 43639 1289 43649 1345
rect 43573 1279 43649 1289
rect 42612 1055 42688 1065
rect 42612 999 42622 1055
rect 42678 999 42688 1055
rect 42612 951 42688 999
rect 42612 895 42622 951
rect 42678 895 42688 951
rect 42612 885 42688 895
rect 43252 1055 43328 1065
rect 43252 999 43262 1055
rect 43318 999 43328 1055
rect 43252 951 43328 999
rect 43252 895 43262 951
rect 43318 895 43328 951
rect 43252 885 43328 895
rect 41346 437 41356 493
rect 41412 437 41460 493
rect 41516 437 41564 493
rect 41620 437 41630 493
rect 41346 389 41630 437
rect 43812 535 44048 1543
rect 47948 1595 48184 2603
rect 50642 2613 50926 2623
rect 50642 2557 50652 2613
rect 50708 2557 50756 2613
rect 50812 2557 50860 2613
rect 50916 2557 50926 2613
rect 48347 2509 48423 2519
rect 48347 2453 48357 2509
rect 48413 2453 48423 2509
rect 48347 2405 48423 2453
rect 48347 2349 48357 2405
rect 48413 2349 48423 2405
rect 48347 2339 48423 2349
rect 48987 2509 49063 2519
rect 48987 2453 48997 2509
rect 49053 2453 49063 2509
rect 48987 2405 49063 2453
rect 48987 2349 48997 2405
rect 49053 2349 49063 2405
rect 48987 2339 49063 2349
rect 50642 2509 50926 2557
rect 53508 2603 53520 2655
rect 53572 2603 53680 2655
rect 53732 2603 53744 2655
rect 50642 2453 50652 2509
rect 50708 2453 50756 2509
rect 50812 2453 50860 2509
rect 50916 2453 50926 2509
rect 50642 2405 50926 2453
rect 50642 2349 50652 2405
rect 50708 2349 50756 2405
rect 50812 2349 50860 2405
rect 50916 2349 50926 2405
rect 50302 2219 50586 2229
rect 50302 2163 50312 2219
rect 50368 2163 50416 2219
rect 50472 2163 50520 2219
rect 50576 2163 50586 2219
rect 48668 2115 48744 2125
rect 48668 2059 48678 2115
rect 48734 2059 48744 2115
rect 48668 2011 48744 2059
rect 48668 1955 48678 2011
rect 48734 1955 48744 2011
rect 48668 1945 48744 1955
rect 49308 2115 49384 2125
rect 49308 2059 49318 2115
rect 49374 2059 49384 2115
rect 49308 2011 49384 2059
rect 49308 1955 49318 2011
rect 49374 1955 49384 2011
rect 49308 1945 49384 1955
rect 50302 2115 50586 2163
rect 50302 2059 50312 2115
rect 50368 2059 50416 2115
rect 50472 2059 50520 2115
rect 50576 2059 50586 2115
rect 50302 2011 50586 2059
rect 50302 1955 50312 2011
rect 50368 1955 50416 2011
rect 50472 1955 50520 2011
rect 50576 1955 50586 2011
rect 47948 1543 47960 1595
rect 48012 1543 48120 1595
rect 48172 1543 48184 1595
rect 44213 1449 44289 1459
rect 44213 1393 44223 1449
rect 44279 1393 44289 1449
rect 44213 1345 44289 1393
rect 44213 1289 44223 1345
rect 44279 1289 44289 1345
rect 44213 1279 44289 1289
rect 44853 1449 44929 1459
rect 44853 1393 44863 1449
rect 44919 1393 44929 1449
rect 44853 1345 44929 1393
rect 44853 1289 44863 1345
rect 44919 1289 44929 1345
rect 44853 1279 44929 1289
rect 47067 1449 47143 1459
rect 47067 1393 47077 1449
rect 47133 1393 47143 1449
rect 47067 1345 47143 1393
rect 47067 1289 47077 1345
rect 47133 1289 47143 1345
rect 47067 1279 47143 1289
rect 47707 1449 47783 1459
rect 47707 1393 47717 1449
rect 47773 1393 47783 1449
rect 47707 1345 47783 1393
rect 47707 1289 47717 1345
rect 47773 1289 47783 1345
rect 47707 1279 47783 1289
rect 44532 1055 44608 1065
rect 44532 999 44542 1055
rect 44598 999 44608 1055
rect 44532 951 44608 999
rect 44532 895 44542 951
rect 44598 895 44608 951
rect 44532 885 44608 895
rect 45172 1055 45248 1065
rect 45172 999 45182 1055
rect 45238 999 45248 1055
rect 45172 951 45248 999
rect 45172 895 45182 951
rect 45238 895 45248 951
rect 45172 885 45248 895
rect 46748 1055 46824 1065
rect 46748 999 46758 1055
rect 46814 999 46824 1055
rect 46748 951 46824 999
rect 46748 895 46758 951
rect 46814 895 46824 951
rect 46748 885 46824 895
rect 47388 1055 47464 1065
rect 47388 999 47398 1055
rect 47454 999 47464 1055
rect 47388 951 47464 999
rect 47388 895 47398 951
rect 47454 895 47464 951
rect 47388 885 47464 895
rect 43812 483 43824 535
rect 43876 483 43984 535
rect 44036 483 44048 535
rect 41346 333 41356 389
rect 41412 333 41460 389
rect 41516 333 41564 389
rect 41620 333 41630 389
rect 41346 285 41630 333
rect 41346 229 41356 285
rect 41412 229 41460 285
rect 41516 229 41564 285
rect 41620 229 41630 285
rect 40626 -1017 40636 -961
rect 40692 -1017 40740 -961
rect 40796 -1017 40844 -961
rect 40900 -1017 40910 -961
rect 34836 -1065 34912 -1055
rect 34836 -1121 34846 -1065
rect 34902 -1121 34912 -1065
rect 34836 -1169 34912 -1121
rect 34836 -1225 34846 -1169
rect 34902 -1225 34912 -1169
rect 34836 -1235 34912 -1225
rect 35476 -1065 35552 -1055
rect 35476 -1121 35486 -1065
rect 35542 -1121 35552 -1065
rect 35476 -1169 35552 -1121
rect 35476 -1225 35486 -1169
rect 35542 -1225 35552 -1169
rect 35476 -1235 35552 -1225
rect 37052 -1065 37128 -1055
rect 37052 -1121 37062 -1065
rect 37118 -1121 37128 -1065
rect 37052 -1169 37128 -1121
rect 37052 -1225 37062 -1169
rect 37118 -1225 37128 -1169
rect 37052 -1235 37128 -1225
rect 37692 -1065 37768 -1055
rect 37692 -1121 37702 -1065
rect 37758 -1121 37768 -1065
rect 37692 -1169 37768 -1121
rect 37692 -1225 37702 -1169
rect 37758 -1225 37768 -1169
rect 37692 -1235 37768 -1225
rect 38972 -1065 39048 -1055
rect 38972 -1121 38982 -1065
rect 39038 -1121 39048 -1065
rect 38972 -1169 39048 -1121
rect 38972 -1225 38982 -1169
rect 39038 -1225 39048 -1169
rect 38972 -1235 39048 -1225
rect 39612 -1065 39688 -1055
rect 39612 -1121 39622 -1065
rect 39678 -1121 39688 -1065
rect 39612 -1169 39688 -1121
rect 39612 -1225 39622 -1169
rect 39678 -1225 39688 -1169
rect 39612 -1235 39688 -1225
rect 40626 -1065 40910 -1017
rect 40626 -1121 40636 -1065
rect 40692 -1121 40740 -1065
rect 40796 -1121 40844 -1065
rect 40900 -1121 40910 -1065
rect 40626 -1169 40910 -1121
rect 40626 -1225 40636 -1169
rect 40692 -1225 40740 -1169
rect 40796 -1225 40844 -1169
rect 40900 -1225 40910 -1169
rect 40626 -1235 40910 -1225
rect 41346 -961 41630 229
rect 42933 389 43009 399
rect 42933 333 42943 389
rect 42999 333 43009 389
rect 42933 285 43009 333
rect 42933 229 42943 285
rect 42999 229 43009 285
rect 42933 219 43009 229
rect 43573 389 43649 399
rect 43573 333 43583 389
rect 43639 333 43649 389
rect 43573 285 43649 333
rect 43573 229 43583 285
rect 43639 229 43649 285
rect 43573 219 43649 229
rect 42612 -5 42688 5
rect 42612 -61 42622 -5
rect 42678 -61 42688 -5
rect 42612 -109 42688 -61
rect 42612 -165 42622 -109
rect 42678 -165 42688 -109
rect 42612 -175 42688 -165
rect 43252 -5 43328 5
rect 43252 -61 43262 -5
rect 43318 -61 43328 -5
rect 43252 -109 43328 -61
rect 43252 -165 43262 -109
rect 43318 -165 43328 -109
rect 43252 -175 43328 -165
rect 43812 -525 44048 483
rect 47948 535 48184 1543
rect 50302 1553 50586 1955
rect 50302 1497 50312 1553
rect 50368 1497 50416 1553
rect 50472 1497 50520 1553
rect 50576 1497 50586 1553
rect 48347 1449 48423 1459
rect 48347 1393 48357 1449
rect 48413 1393 48423 1449
rect 48347 1345 48423 1393
rect 48347 1289 48357 1345
rect 48413 1289 48423 1345
rect 48347 1279 48423 1289
rect 48987 1449 49063 1459
rect 48987 1393 48997 1449
rect 49053 1393 49063 1449
rect 48987 1345 49063 1393
rect 48987 1289 48997 1345
rect 49053 1289 49063 1345
rect 48987 1279 49063 1289
rect 50302 1449 50586 1497
rect 50302 1393 50312 1449
rect 50368 1393 50416 1449
rect 50472 1393 50520 1449
rect 50576 1393 50586 1449
rect 50302 1345 50586 1393
rect 50302 1289 50312 1345
rect 50368 1289 50416 1345
rect 50472 1289 50520 1345
rect 50576 1289 50586 1345
rect 48668 1055 48744 1065
rect 48668 999 48678 1055
rect 48734 999 48744 1055
rect 48668 951 48744 999
rect 48668 895 48678 951
rect 48734 895 48744 951
rect 48668 885 48744 895
rect 49308 1055 49384 1065
rect 49308 999 49318 1055
rect 49374 999 49384 1055
rect 49308 951 49384 999
rect 49308 895 49318 951
rect 49374 895 49384 951
rect 49308 885 49384 895
rect 47948 483 47960 535
rect 48012 483 48120 535
rect 48172 483 48184 535
rect 44213 389 44289 399
rect 44213 333 44223 389
rect 44279 333 44289 389
rect 44213 285 44289 333
rect 44213 229 44223 285
rect 44279 229 44289 285
rect 44213 219 44289 229
rect 44853 389 44929 399
rect 44853 333 44863 389
rect 44919 333 44929 389
rect 44853 285 44929 333
rect 44853 229 44863 285
rect 44919 229 44929 285
rect 44853 219 44929 229
rect 47067 389 47143 399
rect 47067 333 47077 389
rect 47133 333 47143 389
rect 47067 285 47143 333
rect 47067 229 47077 285
rect 47133 229 47143 285
rect 47067 219 47143 229
rect 47707 389 47783 399
rect 47707 333 47717 389
rect 47773 333 47783 389
rect 47707 285 47783 333
rect 47707 229 47717 285
rect 47773 229 47783 285
rect 47707 219 47783 229
rect 44532 -5 44608 5
rect 44532 -61 44542 -5
rect 44598 -61 44608 -5
rect 44532 -109 44608 -61
rect 44532 -165 44542 -109
rect 44598 -165 44608 -109
rect 44532 -175 44608 -165
rect 45172 -5 45248 5
rect 45172 -61 45182 -5
rect 45238 -61 45248 -5
rect 45172 -109 45248 -61
rect 45172 -165 45182 -109
rect 45238 -165 45248 -109
rect 45172 -175 45248 -165
rect 46748 -5 46824 5
rect 46748 -61 46758 -5
rect 46814 -61 46824 -5
rect 46748 -109 46824 -61
rect 46748 -165 46758 -109
rect 46814 -165 46824 -109
rect 46748 -175 46824 -165
rect 47388 -5 47464 5
rect 47388 -61 47398 -5
rect 47454 -61 47464 -5
rect 47388 -109 47464 -61
rect 47388 -165 47398 -109
rect 47454 -165 47464 -109
rect 47388 -175 47464 -165
rect 43812 -577 43824 -525
rect 43876 -577 43984 -525
rect 44036 -577 44048 -525
rect 43812 -589 44048 -577
rect 47948 -525 48184 483
rect 50302 493 50586 1289
rect 50302 437 50312 493
rect 50368 437 50416 493
rect 50472 437 50520 493
rect 50576 437 50586 493
rect 48347 389 48423 399
rect 48347 333 48357 389
rect 48413 333 48423 389
rect 48347 285 48423 333
rect 48347 229 48357 285
rect 48413 229 48423 285
rect 48347 219 48423 229
rect 48987 389 49063 399
rect 48987 333 48997 389
rect 49053 333 49063 389
rect 48987 285 49063 333
rect 48987 229 48997 285
rect 49053 229 49063 285
rect 48987 219 49063 229
rect 50302 389 50586 437
rect 50302 333 50312 389
rect 50368 333 50416 389
rect 50472 333 50520 389
rect 50576 333 50586 389
rect 50302 285 50586 333
rect 50302 229 50312 285
rect 50368 229 50416 285
rect 50472 229 50520 285
rect 50576 229 50586 285
rect 48668 -5 48744 5
rect 48668 -61 48678 -5
rect 48734 -61 48744 -5
rect 48668 -109 48744 -61
rect 48668 -165 48678 -109
rect 48734 -165 48744 -109
rect 48668 -175 48744 -165
rect 49308 -5 49384 5
rect 49308 -61 49318 -5
rect 49374 -61 49384 -5
rect 49308 -109 49384 -61
rect 49308 -165 49318 -109
rect 49374 -165 49384 -109
rect 49308 -175 49384 -165
rect 47948 -577 47960 -525
rect 48012 -577 48120 -525
rect 48172 -577 48184 -525
rect 47948 -589 48184 -577
rect 42933 -671 43009 -661
rect 42933 -727 42943 -671
rect 42999 -727 43009 -671
rect 42933 -775 43009 -727
rect 42933 -831 42943 -775
rect 42999 -831 43009 -775
rect 42933 -841 43009 -831
rect 43573 -671 43649 -661
rect 43573 -727 43583 -671
rect 43639 -727 43649 -671
rect 43573 -775 43649 -727
rect 43573 -831 43583 -775
rect 43639 -831 43649 -775
rect 43573 -841 43649 -831
rect 44213 -671 44289 -661
rect 44213 -727 44223 -671
rect 44279 -727 44289 -671
rect 44213 -775 44289 -727
rect 44213 -831 44223 -775
rect 44279 -831 44289 -775
rect 44213 -841 44289 -831
rect 44853 -671 44929 -661
rect 44853 -727 44863 -671
rect 44919 -727 44929 -671
rect 44853 -775 44929 -727
rect 44853 -831 44863 -775
rect 44919 -831 44929 -775
rect 44853 -841 44929 -831
rect 47067 -671 47143 -661
rect 47067 -727 47077 -671
rect 47133 -727 47143 -671
rect 47067 -775 47143 -727
rect 47067 -831 47077 -775
rect 47133 -831 47143 -775
rect 47067 -841 47143 -831
rect 47707 -671 47783 -661
rect 47707 -727 47717 -671
rect 47773 -727 47783 -671
rect 47707 -775 47783 -727
rect 47707 -831 47717 -775
rect 47773 -831 47783 -775
rect 47707 -841 47783 -831
rect 48347 -671 48423 -661
rect 48347 -727 48357 -671
rect 48413 -727 48423 -671
rect 48347 -775 48423 -727
rect 48347 -831 48357 -775
rect 48413 -831 48423 -775
rect 48347 -841 48423 -831
rect 48987 -671 49063 -661
rect 48987 -727 48997 -671
rect 49053 -727 49063 -671
rect 48987 -775 49063 -727
rect 48987 -831 48997 -775
rect 49053 -831 49063 -775
rect 48987 -841 49063 -831
rect 41346 -1017 41356 -961
rect 41412 -1017 41460 -961
rect 41516 -1017 41564 -961
rect 41620 -1017 41630 -961
rect 41346 -1065 41630 -1017
rect 50302 -961 50586 229
rect 50642 1159 50926 2349
rect 52629 2509 52705 2519
rect 52629 2453 52639 2509
rect 52695 2453 52705 2509
rect 52629 2405 52705 2453
rect 52629 2349 52639 2405
rect 52695 2349 52705 2405
rect 52629 2339 52705 2349
rect 53269 2509 53345 2519
rect 53269 2453 53279 2509
rect 53335 2453 53345 2509
rect 53269 2405 53345 2453
rect 53269 2349 53279 2405
rect 53335 2349 53345 2405
rect 53269 2339 53345 2349
rect 50642 1103 50652 1159
rect 50708 1103 50756 1159
rect 50812 1103 50860 1159
rect 50916 1103 50926 1159
rect 50642 1055 50926 1103
rect 50642 999 50652 1055
rect 50708 999 50756 1055
rect 50812 999 50860 1055
rect 50916 999 50926 1055
rect 50642 951 50926 999
rect 50642 895 50652 951
rect 50708 895 50756 951
rect 50812 895 50860 951
rect 50916 895 50926 951
rect 50642 99 50926 895
rect 50642 43 50652 99
rect 50708 43 50756 99
rect 50812 43 50860 99
rect 50916 43 50926 99
rect 50642 -5 50926 43
rect 50642 -61 50652 -5
rect 50708 -61 50756 -5
rect 50812 -61 50860 -5
rect 50916 -61 50926 -5
rect 50642 -109 50926 -61
rect 50642 -165 50652 -109
rect 50708 -165 50756 -109
rect 50812 -165 50860 -109
rect 50916 -165 50926 -109
rect 50642 -567 50926 -165
rect 50642 -623 50652 -567
rect 50708 -623 50756 -567
rect 50812 -623 50860 -567
rect 50916 -623 50926 -567
rect 50642 -671 50926 -623
rect 50642 -727 50652 -671
rect 50708 -727 50756 -671
rect 50812 -727 50860 -671
rect 50916 -727 50926 -671
rect 50642 -775 50926 -727
rect 50642 -831 50652 -775
rect 50708 -831 50756 -775
rect 50812 -831 50860 -775
rect 50916 -831 50926 -775
rect 50642 -841 50926 -831
rect 51034 2219 51318 2229
rect 51034 2163 51044 2219
rect 51100 2163 51148 2219
rect 51204 2163 51252 2219
rect 51308 2163 51318 2219
rect 51034 2115 51318 2163
rect 51034 2059 51044 2115
rect 51100 2059 51148 2115
rect 51204 2059 51252 2115
rect 51308 2059 51318 2115
rect 51034 2011 51318 2059
rect 51034 1955 51044 2011
rect 51100 1955 51148 2011
rect 51204 1955 51252 2011
rect 51308 1955 51318 2011
rect 51034 1553 51318 1955
rect 52308 2115 52384 2125
rect 52308 2059 52318 2115
rect 52374 2059 52384 2115
rect 52308 2011 52384 2059
rect 52308 1955 52318 2011
rect 52374 1955 52384 2011
rect 52308 1945 52384 1955
rect 52948 2115 53024 2125
rect 52948 2059 52958 2115
rect 53014 2059 53024 2115
rect 52948 2011 53024 2059
rect 52948 1955 52958 2011
rect 53014 1955 53024 2011
rect 52948 1945 53024 1955
rect 51034 1497 51044 1553
rect 51100 1497 51148 1553
rect 51204 1497 51252 1553
rect 51308 1497 51318 1553
rect 51034 1449 51318 1497
rect 53508 1595 53744 2603
rect 57644 2655 57880 3619
rect 57644 2603 57656 2655
rect 57708 2603 57816 2655
rect 57868 2603 57880 2655
rect 63204 2655 63440 3619
rect 53909 2509 53985 2519
rect 53909 2453 53919 2509
rect 53975 2453 53985 2509
rect 53909 2405 53985 2453
rect 53909 2349 53919 2405
rect 53975 2349 53985 2405
rect 53909 2339 53985 2349
rect 54549 2509 54625 2519
rect 54549 2453 54559 2509
rect 54615 2453 54625 2509
rect 54549 2405 54625 2453
rect 54549 2349 54559 2405
rect 54615 2349 54625 2405
rect 54549 2339 54625 2349
rect 56763 2509 56839 2519
rect 56763 2453 56773 2509
rect 56829 2453 56839 2509
rect 56763 2405 56839 2453
rect 56763 2349 56773 2405
rect 56829 2349 56839 2405
rect 56763 2339 56839 2349
rect 57403 2509 57479 2519
rect 57403 2453 57413 2509
rect 57469 2453 57479 2509
rect 57403 2405 57479 2453
rect 57403 2349 57413 2405
rect 57469 2349 57479 2405
rect 57403 2339 57479 2349
rect 54228 2115 54304 2125
rect 54228 2059 54238 2115
rect 54294 2059 54304 2115
rect 54228 2011 54304 2059
rect 54228 1955 54238 2011
rect 54294 1955 54304 2011
rect 54228 1945 54304 1955
rect 54868 2115 54944 2125
rect 54868 2059 54878 2115
rect 54934 2059 54944 2115
rect 54868 2011 54944 2059
rect 54868 1955 54878 2011
rect 54934 1955 54944 2011
rect 54868 1945 54944 1955
rect 56444 2115 56520 2125
rect 56444 2059 56454 2115
rect 56510 2059 56520 2115
rect 56444 2011 56520 2059
rect 56444 1955 56454 2011
rect 56510 1955 56520 2011
rect 56444 1945 56520 1955
rect 57084 2115 57160 2125
rect 57084 2059 57094 2115
rect 57150 2059 57160 2115
rect 57084 2011 57160 2059
rect 57084 1955 57094 2011
rect 57150 1955 57160 2011
rect 57084 1945 57160 1955
rect 53508 1543 53520 1595
rect 53572 1543 53680 1595
rect 53732 1543 53744 1595
rect 51034 1393 51044 1449
rect 51100 1393 51148 1449
rect 51204 1393 51252 1449
rect 51308 1393 51318 1449
rect 51034 1345 51318 1393
rect 51034 1289 51044 1345
rect 51100 1289 51148 1345
rect 51204 1289 51252 1345
rect 51308 1289 51318 1345
rect 51034 493 51318 1289
rect 52629 1449 52705 1459
rect 52629 1393 52639 1449
rect 52695 1393 52705 1449
rect 52629 1345 52705 1393
rect 52629 1289 52639 1345
rect 52695 1289 52705 1345
rect 52629 1279 52705 1289
rect 53269 1449 53345 1459
rect 53269 1393 53279 1449
rect 53335 1393 53345 1449
rect 53269 1345 53345 1393
rect 53269 1289 53279 1345
rect 53335 1289 53345 1345
rect 53269 1279 53345 1289
rect 52308 1055 52384 1065
rect 52308 999 52318 1055
rect 52374 999 52384 1055
rect 52308 951 52384 999
rect 52308 895 52318 951
rect 52374 895 52384 951
rect 52308 885 52384 895
rect 52948 1055 53024 1065
rect 52948 999 52958 1055
rect 53014 999 53024 1055
rect 52948 951 53024 999
rect 52948 895 52958 951
rect 53014 895 53024 951
rect 52948 885 53024 895
rect 51034 437 51044 493
rect 51100 437 51148 493
rect 51204 437 51252 493
rect 51308 437 51318 493
rect 51034 389 51318 437
rect 53508 535 53744 1543
rect 57644 1595 57880 2603
rect 60423 2613 60707 2623
rect 60423 2557 60433 2613
rect 60489 2557 60537 2613
rect 60593 2557 60641 2613
rect 60697 2557 60707 2613
rect 58043 2509 58119 2519
rect 58043 2453 58053 2509
rect 58109 2453 58119 2509
rect 58043 2405 58119 2453
rect 58043 2349 58053 2405
rect 58109 2349 58119 2405
rect 58043 2339 58119 2349
rect 58683 2509 58759 2519
rect 58683 2453 58693 2509
rect 58749 2453 58759 2509
rect 58683 2405 58759 2453
rect 58683 2349 58693 2405
rect 58749 2349 58759 2405
rect 58683 2339 58759 2349
rect 60423 2509 60707 2557
rect 63204 2603 63216 2655
rect 63268 2603 63376 2655
rect 63428 2603 63440 2655
rect 60423 2453 60433 2509
rect 60489 2453 60537 2509
rect 60593 2453 60641 2509
rect 60697 2453 60707 2509
rect 60423 2405 60707 2453
rect 60423 2349 60433 2405
rect 60489 2349 60537 2405
rect 60593 2349 60641 2405
rect 60697 2349 60707 2405
rect 60018 2219 60302 2229
rect 60018 2163 60028 2219
rect 60084 2163 60132 2219
rect 60188 2163 60236 2219
rect 60292 2163 60302 2219
rect 58364 2115 58440 2125
rect 58364 2059 58374 2115
rect 58430 2059 58440 2115
rect 58364 2011 58440 2059
rect 58364 1955 58374 2011
rect 58430 1955 58440 2011
rect 58364 1945 58440 1955
rect 59004 2115 59080 2125
rect 59004 2059 59014 2115
rect 59070 2059 59080 2115
rect 59004 2011 59080 2059
rect 59004 1955 59014 2011
rect 59070 1955 59080 2011
rect 59004 1945 59080 1955
rect 60018 2115 60302 2163
rect 60018 2059 60028 2115
rect 60084 2059 60132 2115
rect 60188 2059 60236 2115
rect 60292 2059 60302 2115
rect 60018 2011 60302 2059
rect 60018 1955 60028 2011
rect 60084 1955 60132 2011
rect 60188 1955 60236 2011
rect 60292 1955 60302 2011
rect 57644 1543 57656 1595
rect 57708 1543 57816 1595
rect 57868 1543 57880 1595
rect 53909 1449 53985 1459
rect 53909 1393 53919 1449
rect 53975 1393 53985 1449
rect 53909 1345 53985 1393
rect 53909 1289 53919 1345
rect 53975 1289 53985 1345
rect 53909 1279 53985 1289
rect 54549 1449 54625 1459
rect 54549 1393 54559 1449
rect 54615 1393 54625 1449
rect 54549 1345 54625 1393
rect 54549 1289 54559 1345
rect 54615 1289 54625 1345
rect 54549 1279 54625 1289
rect 56763 1449 56839 1459
rect 56763 1393 56773 1449
rect 56829 1393 56839 1449
rect 56763 1345 56839 1393
rect 56763 1289 56773 1345
rect 56829 1289 56839 1345
rect 56763 1279 56839 1289
rect 57403 1449 57479 1459
rect 57403 1393 57413 1449
rect 57469 1393 57479 1449
rect 57403 1345 57479 1393
rect 57403 1289 57413 1345
rect 57469 1289 57479 1345
rect 57403 1279 57479 1289
rect 54228 1055 54304 1065
rect 54228 999 54238 1055
rect 54294 999 54304 1055
rect 54228 951 54304 999
rect 54228 895 54238 951
rect 54294 895 54304 951
rect 54228 885 54304 895
rect 54868 1055 54944 1065
rect 54868 999 54878 1055
rect 54934 999 54944 1055
rect 54868 951 54944 999
rect 54868 895 54878 951
rect 54934 895 54944 951
rect 54868 885 54944 895
rect 56444 1055 56520 1065
rect 56444 999 56454 1055
rect 56510 999 56520 1055
rect 56444 951 56520 999
rect 56444 895 56454 951
rect 56510 895 56520 951
rect 56444 885 56520 895
rect 57084 1055 57160 1065
rect 57084 999 57094 1055
rect 57150 999 57160 1055
rect 57084 951 57160 999
rect 57084 895 57094 951
rect 57150 895 57160 951
rect 57084 885 57160 895
rect 53508 483 53520 535
rect 53572 483 53680 535
rect 53732 483 53744 535
rect 51034 333 51044 389
rect 51100 333 51148 389
rect 51204 333 51252 389
rect 51308 333 51318 389
rect 51034 285 51318 333
rect 51034 229 51044 285
rect 51100 229 51148 285
rect 51204 229 51252 285
rect 51308 229 51318 285
rect 50302 -1017 50312 -961
rect 50368 -1017 50416 -961
rect 50472 -1017 50520 -961
rect 50576 -1017 50586 -961
rect 41346 -1121 41356 -1065
rect 41412 -1121 41460 -1065
rect 41516 -1121 41564 -1065
rect 41620 -1121 41630 -1065
rect 41346 -1169 41630 -1121
rect 41346 -1225 41356 -1169
rect 41412 -1225 41460 -1169
rect 41516 -1225 41564 -1169
rect 41620 -1225 41630 -1169
rect 41346 -1235 41630 -1225
rect 42612 -1065 42688 -1055
rect 42612 -1121 42622 -1065
rect 42678 -1121 42688 -1065
rect 42612 -1169 42688 -1121
rect 42612 -1225 42622 -1169
rect 42678 -1225 42688 -1169
rect 42612 -1235 42688 -1225
rect 43252 -1065 43328 -1055
rect 43252 -1121 43262 -1065
rect 43318 -1121 43328 -1065
rect 43252 -1169 43328 -1121
rect 43252 -1225 43262 -1169
rect 43318 -1225 43328 -1169
rect 43252 -1235 43328 -1225
rect 44532 -1065 44608 -1055
rect 44532 -1121 44542 -1065
rect 44598 -1121 44608 -1065
rect 44532 -1169 44608 -1121
rect 44532 -1225 44542 -1169
rect 44598 -1225 44608 -1169
rect 44532 -1235 44608 -1225
rect 45172 -1065 45248 -1055
rect 45172 -1121 45182 -1065
rect 45238 -1121 45248 -1065
rect 45172 -1169 45248 -1121
rect 45172 -1225 45182 -1169
rect 45238 -1225 45248 -1169
rect 45172 -1235 45248 -1225
rect 46748 -1065 46824 -1055
rect 46748 -1121 46758 -1065
rect 46814 -1121 46824 -1065
rect 46748 -1169 46824 -1121
rect 46748 -1225 46758 -1169
rect 46814 -1225 46824 -1169
rect 46748 -1235 46824 -1225
rect 47388 -1065 47464 -1055
rect 47388 -1121 47398 -1065
rect 47454 -1121 47464 -1065
rect 47388 -1169 47464 -1121
rect 47388 -1225 47398 -1169
rect 47454 -1225 47464 -1169
rect 47388 -1235 47464 -1225
rect 48668 -1065 48744 -1055
rect 48668 -1121 48678 -1065
rect 48734 -1121 48744 -1065
rect 48668 -1169 48744 -1121
rect 48668 -1225 48678 -1169
rect 48734 -1225 48744 -1169
rect 48668 -1235 48744 -1225
rect 49308 -1065 49384 -1055
rect 49308 -1121 49318 -1065
rect 49374 -1121 49384 -1065
rect 49308 -1169 49384 -1121
rect 49308 -1225 49318 -1169
rect 49374 -1225 49384 -1169
rect 49308 -1235 49384 -1225
rect 50302 -1065 50586 -1017
rect 50302 -1121 50312 -1065
rect 50368 -1121 50416 -1065
rect 50472 -1121 50520 -1065
rect 50576 -1121 50586 -1065
rect 50302 -1169 50586 -1121
rect 50302 -1225 50312 -1169
rect 50368 -1225 50416 -1169
rect 50472 -1225 50520 -1169
rect 50576 -1225 50586 -1169
rect 50302 -1235 50586 -1225
rect 51034 -961 51318 229
rect 52629 389 52705 399
rect 52629 333 52639 389
rect 52695 333 52705 389
rect 52629 285 52705 333
rect 52629 229 52639 285
rect 52695 229 52705 285
rect 52629 219 52705 229
rect 53269 389 53345 399
rect 53269 333 53279 389
rect 53335 333 53345 389
rect 53269 285 53345 333
rect 53269 229 53279 285
rect 53335 229 53345 285
rect 53269 219 53345 229
rect 52308 -5 52384 5
rect 52308 -61 52318 -5
rect 52374 -61 52384 -5
rect 52308 -109 52384 -61
rect 52308 -165 52318 -109
rect 52374 -165 52384 -109
rect 52308 -175 52384 -165
rect 52948 -5 53024 5
rect 52948 -61 52958 -5
rect 53014 -61 53024 -5
rect 52948 -109 53024 -61
rect 52948 -165 52958 -109
rect 53014 -165 53024 -109
rect 52948 -175 53024 -165
rect 53508 -525 53744 483
rect 57644 535 57880 1543
rect 60018 1553 60302 1955
rect 60018 1497 60028 1553
rect 60084 1497 60132 1553
rect 60188 1497 60236 1553
rect 60292 1497 60302 1553
rect 58043 1449 58119 1459
rect 58043 1393 58053 1449
rect 58109 1393 58119 1449
rect 58043 1345 58119 1393
rect 58043 1289 58053 1345
rect 58109 1289 58119 1345
rect 58043 1279 58119 1289
rect 58683 1449 58759 1459
rect 58683 1393 58693 1449
rect 58749 1393 58759 1449
rect 58683 1345 58759 1393
rect 58683 1289 58693 1345
rect 58749 1289 58759 1345
rect 58683 1279 58759 1289
rect 60018 1449 60302 1497
rect 60018 1393 60028 1449
rect 60084 1393 60132 1449
rect 60188 1393 60236 1449
rect 60292 1393 60302 1449
rect 60018 1345 60302 1393
rect 60018 1289 60028 1345
rect 60084 1289 60132 1345
rect 60188 1289 60236 1345
rect 60292 1289 60302 1345
rect 58364 1055 58440 1065
rect 58364 999 58374 1055
rect 58430 999 58440 1055
rect 58364 951 58440 999
rect 58364 895 58374 951
rect 58430 895 58440 951
rect 58364 885 58440 895
rect 59004 1055 59080 1065
rect 59004 999 59014 1055
rect 59070 999 59080 1055
rect 59004 951 59080 999
rect 59004 895 59014 951
rect 59070 895 59080 951
rect 59004 885 59080 895
rect 57644 483 57656 535
rect 57708 483 57816 535
rect 57868 483 57880 535
rect 53909 389 53985 399
rect 53909 333 53919 389
rect 53975 333 53985 389
rect 53909 285 53985 333
rect 53909 229 53919 285
rect 53975 229 53985 285
rect 53909 219 53985 229
rect 54549 389 54625 399
rect 54549 333 54559 389
rect 54615 333 54625 389
rect 54549 285 54625 333
rect 54549 229 54559 285
rect 54615 229 54625 285
rect 54549 219 54625 229
rect 56763 389 56839 399
rect 56763 333 56773 389
rect 56829 333 56839 389
rect 56763 285 56839 333
rect 56763 229 56773 285
rect 56829 229 56839 285
rect 56763 219 56839 229
rect 57403 389 57479 399
rect 57403 333 57413 389
rect 57469 333 57479 389
rect 57403 285 57479 333
rect 57403 229 57413 285
rect 57469 229 57479 285
rect 57403 219 57479 229
rect 54228 -5 54304 5
rect 54228 -61 54238 -5
rect 54294 -61 54304 -5
rect 54228 -109 54304 -61
rect 54228 -165 54238 -109
rect 54294 -165 54304 -109
rect 54228 -175 54304 -165
rect 54868 -5 54944 5
rect 54868 -61 54878 -5
rect 54934 -61 54944 -5
rect 54868 -109 54944 -61
rect 54868 -165 54878 -109
rect 54934 -165 54944 -109
rect 54868 -175 54944 -165
rect 56444 -5 56520 5
rect 56444 -61 56454 -5
rect 56510 -61 56520 -5
rect 56444 -109 56520 -61
rect 56444 -165 56454 -109
rect 56510 -165 56520 -109
rect 56444 -175 56520 -165
rect 57084 -5 57160 5
rect 57084 -61 57094 -5
rect 57150 -61 57160 -5
rect 57084 -109 57160 -61
rect 57084 -165 57094 -109
rect 57150 -165 57160 -109
rect 57084 -175 57160 -165
rect 53508 -577 53520 -525
rect 53572 -577 53680 -525
rect 53732 -577 53744 -525
rect 53508 -589 53744 -577
rect 57644 -525 57880 483
rect 60018 493 60302 1289
rect 60018 437 60028 493
rect 60084 437 60132 493
rect 60188 437 60236 493
rect 60292 437 60302 493
rect 58043 389 58119 399
rect 58043 333 58053 389
rect 58109 333 58119 389
rect 58043 285 58119 333
rect 58043 229 58053 285
rect 58109 229 58119 285
rect 58043 219 58119 229
rect 58683 389 58759 399
rect 58683 333 58693 389
rect 58749 333 58759 389
rect 58683 285 58759 333
rect 58683 229 58693 285
rect 58749 229 58759 285
rect 58683 219 58759 229
rect 60018 389 60302 437
rect 60018 333 60028 389
rect 60084 333 60132 389
rect 60188 333 60236 389
rect 60292 333 60302 389
rect 60018 285 60302 333
rect 60018 229 60028 285
rect 60084 229 60132 285
rect 60188 229 60236 285
rect 60292 229 60302 285
rect 58364 -5 58440 5
rect 58364 -61 58374 -5
rect 58430 -61 58440 -5
rect 58364 -109 58440 -61
rect 58364 -165 58374 -109
rect 58430 -165 58440 -109
rect 58364 -175 58440 -165
rect 59004 -5 59080 5
rect 59004 -61 59014 -5
rect 59070 -61 59080 -5
rect 59004 -109 59080 -61
rect 59004 -165 59014 -109
rect 59070 -165 59080 -109
rect 59004 -175 59080 -165
rect 57644 -577 57656 -525
rect 57708 -577 57816 -525
rect 57868 -577 57880 -525
rect 57644 -589 57880 -577
rect 52629 -671 52705 -661
rect 52629 -727 52639 -671
rect 52695 -727 52705 -671
rect 52629 -775 52705 -727
rect 52629 -831 52639 -775
rect 52695 -831 52705 -775
rect 52629 -841 52705 -831
rect 53269 -671 53345 -661
rect 53269 -727 53279 -671
rect 53335 -727 53345 -671
rect 53269 -775 53345 -727
rect 53269 -831 53279 -775
rect 53335 -831 53345 -775
rect 53269 -841 53345 -831
rect 53909 -671 53985 -661
rect 53909 -727 53919 -671
rect 53975 -727 53985 -671
rect 53909 -775 53985 -727
rect 53909 -831 53919 -775
rect 53975 -831 53985 -775
rect 53909 -841 53985 -831
rect 54549 -671 54625 -661
rect 54549 -727 54559 -671
rect 54615 -727 54625 -671
rect 54549 -775 54625 -727
rect 54549 -831 54559 -775
rect 54615 -831 54625 -775
rect 54549 -841 54625 -831
rect 56763 -671 56839 -661
rect 56763 -727 56773 -671
rect 56829 -727 56839 -671
rect 56763 -775 56839 -727
rect 56763 -831 56773 -775
rect 56829 -831 56839 -775
rect 56763 -841 56839 -831
rect 57403 -671 57479 -661
rect 57403 -727 57413 -671
rect 57469 -727 57479 -671
rect 57403 -775 57479 -727
rect 57403 -831 57413 -775
rect 57469 -831 57479 -775
rect 57403 -841 57479 -831
rect 58043 -671 58119 -661
rect 58043 -727 58053 -671
rect 58109 -727 58119 -671
rect 58043 -775 58119 -727
rect 58043 -831 58053 -775
rect 58109 -831 58119 -775
rect 58043 -841 58119 -831
rect 58683 -671 58759 -661
rect 58683 -727 58693 -671
rect 58749 -727 58759 -671
rect 58683 -775 58759 -727
rect 58683 -831 58693 -775
rect 58749 -831 58759 -775
rect 58683 -841 58759 -831
rect 51034 -1017 51044 -961
rect 51100 -1017 51148 -961
rect 51204 -1017 51252 -961
rect 51308 -1017 51318 -961
rect 51034 -1065 51318 -1017
rect 60018 -961 60302 229
rect 60423 1159 60707 2349
rect 62325 2509 62401 2519
rect 62325 2453 62335 2509
rect 62391 2453 62401 2509
rect 62325 2405 62401 2453
rect 62325 2349 62335 2405
rect 62391 2349 62401 2405
rect 62325 2339 62401 2349
rect 62965 2509 63041 2519
rect 62965 2453 62975 2509
rect 63031 2453 63041 2509
rect 62965 2405 63041 2453
rect 62965 2349 62975 2405
rect 63031 2349 63041 2405
rect 62965 2339 63041 2349
rect 60423 1103 60433 1159
rect 60489 1103 60537 1159
rect 60593 1103 60641 1159
rect 60697 1103 60707 1159
rect 60423 1055 60707 1103
rect 60423 999 60433 1055
rect 60489 999 60537 1055
rect 60593 999 60641 1055
rect 60697 999 60707 1055
rect 60423 951 60707 999
rect 60423 895 60433 951
rect 60489 895 60537 951
rect 60593 895 60641 951
rect 60697 895 60707 951
rect 60423 99 60707 895
rect 60423 43 60433 99
rect 60489 43 60537 99
rect 60593 43 60641 99
rect 60697 43 60707 99
rect 60423 -5 60707 43
rect 60423 -61 60433 -5
rect 60489 -61 60537 -5
rect 60593 -61 60641 -5
rect 60697 -61 60707 -5
rect 60423 -109 60707 -61
rect 60423 -165 60433 -109
rect 60489 -165 60537 -109
rect 60593 -165 60641 -109
rect 60697 -165 60707 -109
rect 60423 -567 60707 -165
rect 60423 -623 60433 -567
rect 60489 -623 60537 -567
rect 60593 -623 60641 -567
rect 60697 -623 60707 -567
rect 60423 -671 60707 -623
rect 60423 -727 60433 -671
rect 60489 -727 60537 -671
rect 60593 -727 60641 -671
rect 60697 -727 60707 -671
rect 60423 -775 60707 -727
rect 60423 -831 60433 -775
rect 60489 -831 60537 -775
rect 60593 -831 60641 -775
rect 60697 -831 60707 -775
rect 60423 -841 60707 -831
rect 60782 2219 61066 2229
rect 60782 2163 60792 2219
rect 60848 2163 60896 2219
rect 60952 2163 61000 2219
rect 61056 2163 61066 2219
rect 60782 2115 61066 2163
rect 60782 2059 60792 2115
rect 60848 2059 60896 2115
rect 60952 2059 61000 2115
rect 61056 2059 61066 2115
rect 60782 2011 61066 2059
rect 60782 1955 60792 2011
rect 60848 1955 60896 2011
rect 60952 1955 61000 2011
rect 61056 1955 61066 2011
rect 60782 1553 61066 1955
rect 62004 2115 62080 2125
rect 62004 2059 62014 2115
rect 62070 2059 62080 2115
rect 62004 2011 62080 2059
rect 62004 1955 62014 2011
rect 62070 1955 62080 2011
rect 62004 1945 62080 1955
rect 62644 2115 62720 2125
rect 62644 2059 62654 2115
rect 62710 2059 62720 2115
rect 62644 2011 62720 2059
rect 62644 1955 62654 2011
rect 62710 1955 62720 2011
rect 62644 1945 62720 1955
rect 60782 1497 60792 1553
rect 60848 1497 60896 1553
rect 60952 1497 61000 1553
rect 61056 1497 61066 1553
rect 60782 1449 61066 1497
rect 63204 1595 63440 2603
rect 63605 2509 63681 2519
rect 63605 2453 63615 2509
rect 63671 2453 63681 2509
rect 63605 2405 63681 2453
rect 63605 2349 63615 2405
rect 63671 2349 63681 2405
rect 63605 2339 63681 2349
rect 64245 2509 64321 2519
rect 64245 2453 64255 2509
rect 64311 2453 64321 2509
rect 64245 2405 64321 2453
rect 64245 2349 64255 2405
rect 64311 2349 64321 2405
rect 64245 2339 64321 2349
rect 63924 2115 64000 2125
rect 63924 2059 63934 2115
rect 63990 2059 64000 2115
rect 63924 2011 64000 2059
rect 63924 1955 63934 2011
rect 63990 1955 64000 2011
rect 63924 1945 64000 1955
rect 64564 2115 64640 2125
rect 64564 2059 64574 2115
rect 64630 2059 64640 2115
rect 64564 2011 64640 2059
rect 64564 1955 64574 2011
rect 64630 1955 64640 2011
rect 64564 1945 64640 1955
rect 63204 1543 63216 1595
rect 63268 1543 63376 1595
rect 63428 1543 63440 1595
rect 60782 1393 60792 1449
rect 60848 1393 60896 1449
rect 60952 1393 61000 1449
rect 61056 1393 61066 1449
rect 60782 1345 61066 1393
rect 60782 1289 60792 1345
rect 60848 1289 60896 1345
rect 60952 1289 61000 1345
rect 61056 1289 61066 1345
rect 60782 493 61066 1289
rect 62325 1449 62401 1459
rect 62325 1393 62335 1449
rect 62391 1393 62401 1449
rect 62325 1345 62401 1393
rect 62325 1289 62335 1345
rect 62391 1289 62401 1345
rect 62325 1279 62401 1289
rect 62965 1449 63041 1459
rect 62965 1393 62975 1449
rect 63031 1393 63041 1449
rect 62965 1345 63041 1393
rect 62965 1289 62975 1345
rect 63031 1289 63041 1345
rect 62965 1279 63041 1289
rect 62004 1055 62080 1065
rect 62004 999 62014 1055
rect 62070 999 62080 1055
rect 62004 951 62080 999
rect 62004 895 62014 951
rect 62070 895 62080 951
rect 62004 885 62080 895
rect 62644 1055 62720 1065
rect 62644 999 62654 1055
rect 62710 999 62720 1055
rect 62644 951 62720 999
rect 62644 895 62654 951
rect 62710 895 62720 951
rect 62644 885 62720 895
rect 60782 437 60792 493
rect 60848 437 60896 493
rect 60952 437 61000 493
rect 61056 437 61066 493
rect 60782 389 61066 437
rect 63204 535 63440 1543
rect 63605 1449 63681 1459
rect 63605 1393 63615 1449
rect 63671 1393 63681 1449
rect 63605 1345 63681 1393
rect 63605 1289 63615 1345
rect 63671 1289 63681 1345
rect 63605 1279 63681 1289
rect 64245 1449 64321 1459
rect 64245 1393 64255 1449
rect 64311 1393 64321 1449
rect 64245 1345 64321 1393
rect 64245 1289 64255 1345
rect 64311 1289 64321 1345
rect 64245 1279 64321 1289
rect 63924 1055 64000 1065
rect 63924 999 63934 1055
rect 63990 999 64000 1055
rect 63924 951 64000 999
rect 63924 895 63934 951
rect 63990 895 64000 951
rect 63924 885 64000 895
rect 64564 1055 64640 1065
rect 64564 999 64574 1055
rect 64630 999 64640 1055
rect 64564 951 64640 999
rect 64564 895 64574 951
rect 64630 895 64640 951
rect 64564 885 64640 895
rect 63204 483 63216 535
rect 63268 483 63376 535
rect 63428 483 63440 535
rect 60782 333 60792 389
rect 60848 333 60896 389
rect 60952 333 61000 389
rect 61056 333 61066 389
rect 60782 285 61066 333
rect 60782 229 60792 285
rect 60848 229 60896 285
rect 60952 229 61000 285
rect 61056 229 61066 285
rect 60018 -1017 60028 -961
rect 60084 -1017 60132 -961
rect 60188 -1017 60236 -961
rect 60292 -1017 60302 -961
rect 51034 -1121 51044 -1065
rect 51100 -1121 51148 -1065
rect 51204 -1121 51252 -1065
rect 51308 -1121 51318 -1065
rect 51034 -1169 51318 -1121
rect 51034 -1225 51044 -1169
rect 51100 -1225 51148 -1169
rect 51204 -1225 51252 -1169
rect 51308 -1225 51318 -1169
rect 51034 -1235 51318 -1225
rect 52308 -1065 52384 -1055
rect 52308 -1121 52318 -1065
rect 52374 -1121 52384 -1065
rect 52308 -1169 52384 -1121
rect 52308 -1225 52318 -1169
rect 52374 -1225 52384 -1169
rect 52308 -1235 52384 -1225
rect 52948 -1065 53024 -1055
rect 52948 -1121 52958 -1065
rect 53014 -1121 53024 -1065
rect 52948 -1169 53024 -1121
rect 52948 -1225 52958 -1169
rect 53014 -1225 53024 -1169
rect 52948 -1235 53024 -1225
rect 54228 -1065 54304 -1055
rect 54228 -1121 54238 -1065
rect 54294 -1121 54304 -1065
rect 54228 -1169 54304 -1121
rect 54228 -1225 54238 -1169
rect 54294 -1225 54304 -1169
rect 54228 -1235 54304 -1225
rect 54868 -1065 54944 -1055
rect 54868 -1121 54878 -1065
rect 54934 -1121 54944 -1065
rect 54868 -1169 54944 -1121
rect 54868 -1225 54878 -1169
rect 54934 -1225 54944 -1169
rect 54868 -1235 54944 -1225
rect 56444 -1065 56520 -1055
rect 56444 -1121 56454 -1065
rect 56510 -1121 56520 -1065
rect 56444 -1169 56520 -1121
rect 56444 -1225 56454 -1169
rect 56510 -1225 56520 -1169
rect 56444 -1235 56520 -1225
rect 57084 -1065 57160 -1055
rect 57084 -1121 57094 -1065
rect 57150 -1121 57160 -1065
rect 57084 -1169 57160 -1121
rect 57084 -1225 57094 -1169
rect 57150 -1225 57160 -1169
rect 57084 -1235 57160 -1225
rect 58364 -1065 58440 -1055
rect 58364 -1121 58374 -1065
rect 58430 -1121 58440 -1065
rect 58364 -1169 58440 -1121
rect 58364 -1225 58374 -1169
rect 58430 -1225 58440 -1169
rect 58364 -1235 58440 -1225
rect 59004 -1065 59080 -1055
rect 59004 -1121 59014 -1065
rect 59070 -1121 59080 -1065
rect 59004 -1169 59080 -1121
rect 59004 -1225 59014 -1169
rect 59070 -1225 59080 -1169
rect 59004 -1235 59080 -1225
rect 60018 -1065 60302 -1017
rect 60018 -1121 60028 -1065
rect 60084 -1121 60132 -1065
rect 60188 -1121 60236 -1065
rect 60292 -1121 60302 -1065
rect 60018 -1169 60302 -1121
rect 60018 -1225 60028 -1169
rect 60084 -1225 60132 -1169
rect 60188 -1225 60236 -1169
rect 60292 -1225 60302 -1169
rect 60018 -1235 60302 -1225
rect 60782 -961 61066 229
rect 62325 389 62401 399
rect 62325 333 62335 389
rect 62391 333 62401 389
rect 62325 285 62401 333
rect 62325 229 62335 285
rect 62391 229 62401 285
rect 62325 219 62401 229
rect 62965 389 63041 399
rect 62965 333 62975 389
rect 63031 333 63041 389
rect 62965 285 63041 333
rect 62965 229 62975 285
rect 63031 229 63041 285
rect 62965 219 63041 229
rect 62004 -5 62080 5
rect 62004 -61 62014 -5
rect 62070 -61 62080 -5
rect 62004 -109 62080 -61
rect 62004 -165 62014 -109
rect 62070 -165 62080 -109
rect 62004 -175 62080 -165
rect 62644 -5 62720 5
rect 62644 -61 62654 -5
rect 62710 -61 62720 -5
rect 62644 -109 62720 -61
rect 62644 -165 62654 -109
rect 62710 -165 62720 -109
rect 62644 -175 62720 -165
rect 63204 -525 63440 483
rect 63605 389 63681 399
rect 63605 333 63615 389
rect 63671 333 63681 389
rect 63605 285 63681 333
rect 63605 229 63615 285
rect 63671 229 63681 285
rect 63605 219 63681 229
rect 64245 389 64321 399
rect 64245 333 64255 389
rect 64311 333 64321 389
rect 64245 285 64321 333
rect 64245 229 64255 285
rect 64311 229 64321 285
rect 64245 219 64321 229
rect 63924 -5 64000 5
rect 63924 -61 63934 -5
rect 63990 -61 64000 -5
rect 63924 -109 64000 -61
rect 63924 -165 63934 -109
rect 63990 -165 64000 -109
rect 63924 -175 64000 -165
rect 64564 -5 64640 5
rect 64564 -61 64574 -5
rect 64630 -61 64640 -5
rect 64564 -109 64640 -61
rect 64564 -165 64574 -109
rect 64630 -165 64640 -109
rect 64564 -175 64640 -165
rect 63204 -577 63216 -525
rect 63268 -577 63376 -525
rect 63428 -577 63440 -525
rect 63204 -589 63440 -577
rect 62325 -671 62401 -661
rect 62325 -727 62335 -671
rect 62391 -727 62401 -671
rect 62325 -775 62401 -727
rect 62325 -831 62335 -775
rect 62391 -831 62401 -775
rect 62325 -841 62401 -831
rect 62965 -671 63041 -661
rect 62965 -727 62975 -671
rect 63031 -727 63041 -671
rect 62965 -775 63041 -727
rect 62965 -831 62975 -775
rect 63031 -831 63041 -775
rect 62965 -841 63041 -831
rect 63605 -671 63681 -661
rect 63605 -727 63615 -671
rect 63671 -727 63681 -671
rect 63605 -775 63681 -727
rect 63605 -831 63615 -775
rect 63671 -831 63681 -775
rect 63605 -841 63681 -831
rect 64245 -671 64321 -661
rect 64245 -727 64255 -671
rect 64311 -727 64321 -671
rect 64245 -775 64321 -727
rect 64245 -831 64255 -775
rect 64311 -831 64321 -775
rect 64245 -841 64321 -831
rect 60782 -1017 60792 -961
rect 60848 -1017 60896 -961
rect 60952 -1017 61000 -961
rect 61056 -1017 61066 -961
rect 60782 -1065 61066 -1017
rect 60782 -1121 60792 -1065
rect 60848 -1121 60896 -1065
rect 60952 -1121 61000 -1065
rect 61056 -1121 61066 -1065
rect 60782 -1169 61066 -1121
rect 60782 -1225 60792 -1169
rect 60848 -1225 60896 -1169
rect 60952 -1225 61000 -1169
rect 61056 -1225 61066 -1169
rect 60782 -1235 61066 -1225
rect 62004 -1065 62080 -1055
rect 62004 -1121 62014 -1065
rect 62070 -1121 62080 -1065
rect 62004 -1169 62080 -1121
rect 62004 -1225 62014 -1169
rect 62070 -1225 62080 -1169
rect 62004 -1235 62080 -1225
rect 62644 -1065 62720 -1055
rect 62644 -1121 62654 -1065
rect 62710 -1121 62720 -1065
rect 62644 -1169 62720 -1121
rect 62644 -1225 62654 -1169
rect 62710 -1225 62720 -1169
rect 62644 -1235 62720 -1225
rect 63924 -1065 64000 -1055
rect 63924 -1121 63934 -1065
rect 63990 -1121 64000 -1065
rect 63924 -1169 64000 -1121
rect 63924 -1225 63934 -1169
rect 63990 -1225 64000 -1169
rect 63924 -1235 64000 -1225
rect 64564 -1065 64640 -1055
rect 64564 -1121 64574 -1065
rect 64630 -1121 64640 -1065
rect 64564 -1169 64640 -1121
rect 64564 -1225 64574 -1169
rect 64630 -1225 64640 -1169
rect 64564 -1235 64640 -1225
rect 54292 -3569 54491 -3556
rect 54292 -3625 54309 -3569
rect 54365 -3625 54419 -3569
rect 54475 -3625 54491 -3569
rect 54292 -3642 54491 -3625
rect 34116 -5649 34154 -5593
rect 34210 -5649 34258 -5593
rect 34314 -5649 34352 -5593
rect 34116 -5697 34352 -5649
rect 34116 -5753 34154 -5697
rect 34210 -5753 34258 -5697
rect 34314 -5753 34352 -5697
rect 34116 -5763 34352 -5753
rect 44536 -7954 45028 -7944
rect 44536 -8010 44546 -7954
rect 44602 -8010 44650 -7954
rect 44706 -8010 44754 -7954
rect 44810 -8010 44858 -7954
rect 44914 -8010 44962 -7954
rect 45018 -8010 45028 -7954
rect 34706 -8054 35198 -8044
rect 34706 -8110 34716 -8054
rect 34772 -8110 34820 -8054
rect 34876 -8110 34924 -8054
rect 34980 -8110 35028 -8054
rect 35084 -8110 35132 -8054
rect 35188 -8110 35198 -8054
rect 34706 -8158 35198 -8110
rect 34706 -8214 34716 -8158
rect 34772 -8214 34820 -8158
rect 34876 -8214 34924 -8158
rect 34980 -8214 35028 -8158
rect 35084 -8214 35132 -8158
rect 35188 -8214 35198 -8158
rect 34706 -8262 35198 -8214
rect 34706 -8318 34716 -8262
rect 34772 -8318 34820 -8262
rect 34876 -8318 34924 -8262
rect 34980 -8318 35028 -8262
rect 35084 -8318 35132 -8262
rect 35188 -8318 35198 -8262
rect 34706 -8366 35198 -8318
rect 34706 -8422 34716 -8366
rect 34772 -8422 34820 -8366
rect 34876 -8422 34924 -8366
rect 34980 -8422 35028 -8366
rect 35084 -8422 35132 -8366
rect 35188 -8422 35198 -8366
rect 34706 -8470 35198 -8422
rect 34706 -8526 34716 -8470
rect 34772 -8526 34820 -8470
rect 34876 -8526 34924 -8470
rect 34980 -8526 35028 -8470
rect 35084 -8526 35132 -8470
rect 35188 -8526 35198 -8470
rect 34706 -8536 35198 -8526
rect 39146 -8054 39638 -8044
rect 39146 -8110 39156 -8054
rect 39212 -8110 39260 -8054
rect 39316 -8110 39364 -8054
rect 39420 -8110 39468 -8054
rect 39524 -8110 39572 -8054
rect 39628 -8110 39638 -8054
rect 39146 -8158 39638 -8110
rect 39146 -8214 39156 -8158
rect 39212 -8214 39260 -8158
rect 39316 -8214 39364 -8158
rect 39420 -8214 39468 -8158
rect 39524 -8214 39572 -8158
rect 39628 -8214 39638 -8158
rect 39146 -8262 39638 -8214
rect 39146 -8318 39156 -8262
rect 39212 -8318 39260 -8262
rect 39316 -8318 39364 -8262
rect 39420 -8318 39468 -8262
rect 39524 -8318 39572 -8262
rect 39628 -8318 39638 -8262
rect 39146 -8366 39638 -8318
rect 39146 -8422 39156 -8366
rect 39212 -8422 39260 -8366
rect 39316 -8422 39364 -8366
rect 39420 -8422 39468 -8366
rect 39524 -8422 39572 -8366
rect 39628 -8422 39638 -8366
rect 39146 -8470 39638 -8422
rect 44536 -8058 45028 -8010
rect 44536 -8114 44546 -8058
rect 44602 -8114 44650 -8058
rect 44706 -8114 44754 -8058
rect 44810 -8114 44858 -8058
rect 44914 -8114 44962 -8058
rect 45018 -8114 45028 -8058
rect 44536 -8162 45028 -8114
rect 44536 -8218 44546 -8162
rect 44602 -8218 44650 -8162
rect 44706 -8218 44754 -8162
rect 44810 -8218 44858 -8162
rect 44914 -8218 44962 -8162
rect 45018 -8218 45028 -8162
rect 44536 -8266 45028 -8218
rect 44536 -8322 44546 -8266
rect 44602 -8322 44650 -8266
rect 44706 -8322 44754 -8266
rect 44810 -8322 44858 -8266
rect 44914 -8322 44962 -8266
rect 45018 -8322 45028 -8266
rect 44536 -8370 45028 -8322
rect 44536 -8426 44546 -8370
rect 44602 -8426 44650 -8370
rect 44706 -8426 44754 -8370
rect 44810 -8426 44858 -8370
rect 44914 -8426 44962 -8370
rect 45018 -8426 45028 -8370
rect 44536 -8436 45028 -8426
rect 48976 -7954 49468 -7944
rect 48976 -8010 48986 -7954
rect 49042 -8010 49090 -7954
rect 49146 -8010 49194 -7954
rect 49250 -8010 49298 -7954
rect 49354 -8010 49402 -7954
rect 49458 -8010 49468 -7954
rect 48976 -8058 49468 -8010
rect 48976 -8114 48986 -8058
rect 49042 -8114 49090 -8058
rect 49146 -8114 49194 -8058
rect 49250 -8114 49298 -8058
rect 49354 -8114 49402 -8058
rect 49458 -8114 49468 -8058
rect 48976 -8162 49468 -8114
rect 48976 -8218 48986 -8162
rect 49042 -8218 49090 -8162
rect 49146 -8218 49194 -8162
rect 49250 -8218 49298 -8162
rect 49354 -8218 49402 -8162
rect 49458 -8218 49468 -8162
rect 48976 -8266 49468 -8218
rect 48976 -8322 48986 -8266
rect 49042 -8322 49090 -8266
rect 49146 -8322 49194 -8266
rect 49250 -8322 49298 -8266
rect 49354 -8322 49402 -8266
rect 49458 -8322 49468 -8266
rect 48976 -8370 49468 -8322
rect 48976 -8426 48986 -8370
rect 49042 -8426 49090 -8370
rect 49146 -8426 49194 -8370
rect 49250 -8426 49298 -8370
rect 49354 -8426 49402 -8370
rect 49458 -8426 49468 -8370
rect 48976 -8436 49468 -8426
rect 39146 -8526 39156 -8470
rect 39212 -8526 39260 -8470
rect 39316 -8526 39364 -8470
rect 39420 -8526 39468 -8470
rect 39524 -8526 39572 -8470
rect 39628 -8526 39638 -8470
rect 39146 -8536 39638 -8526
rect 31640 -8827 31650 -8771
rect 31706 -8827 31754 -8771
rect 31810 -8827 31858 -8771
rect 31914 -8827 31924 -8771
rect 31640 -8875 31924 -8827
rect 31640 -8931 31650 -8875
rect 31706 -8931 31754 -8875
rect 31810 -8931 31858 -8875
rect 31914 -8931 31924 -8875
rect 31640 -8979 31924 -8931
rect 31640 -9035 31650 -8979
rect 31706 -9035 31754 -8979
rect 31810 -9035 31858 -8979
rect 31914 -9035 31924 -8979
rect 31640 -9045 31924 -9035
rect 16938 -9391 17159 -9382
rect 16938 -9447 16967 -9391
rect 17023 -9447 17077 -9391
rect 17133 -9447 17159 -9391
rect 16938 -9501 17159 -9447
rect 16938 -9557 16967 -9501
rect 17023 -9557 17077 -9501
rect 17133 -9557 17159 -9501
rect 16938 -9562 17159 -9557
rect 14917 -9633 15138 -9624
rect 14917 -9689 14946 -9633
rect 15002 -9689 15056 -9633
rect 15112 -9689 15138 -9633
rect 14917 -9743 15138 -9689
rect 14917 -9799 14946 -9743
rect 15002 -9799 15056 -9743
rect 15112 -9799 15138 -9743
rect 14917 -9804 15138 -9799
rect 12954 -9875 13175 -9866
rect 12954 -9931 12983 -9875
rect 13039 -9931 13093 -9875
rect 13149 -9931 13175 -9875
rect 12954 -9985 13175 -9931
rect 12954 -10041 12983 -9985
rect 13039 -10041 13093 -9985
rect 13149 -10041 13175 -9985
rect 12954 -10046 13175 -10041
rect 10947 -10120 11168 -10111
rect 10947 -10176 10976 -10120
rect 11032 -10176 11086 -10120
rect 11142 -10176 11168 -10120
rect 10947 -10230 11168 -10176
rect 10947 -10286 10976 -10230
rect 11032 -10286 11086 -10230
rect 11142 -10286 11168 -10230
rect 10947 -10291 11168 -10286
rect 8912 -10356 9133 -10347
rect 8912 -10412 8941 -10356
rect 8997 -10412 9051 -10356
rect 9107 -10412 9133 -10356
rect 8912 -10466 9133 -10412
rect 8912 -10522 8941 -10466
rect 8997 -10522 9051 -10466
rect 9107 -10522 9133 -10466
rect 8912 -10527 9133 -10522
rect 6825 -10598 7046 -10589
rect 6825 -10654 6854 -10598
rect 6910 -10654 6964 -10598
rect 7020 -10654 7046 -10598
rect 6825 -10708 7046 -10654
rect 6825 -10764 6854 -10708
rect 6910 -10764 6964 -10708
rect 7020 -10764 7046 -10708
rect 6825 -10769 7046 -10764
rect -1115 -11442 -667 -11433
rect -1115 -11498 -1086 -11442
rect -1030 -11498 -976 -11442
rect -920 -11498 -858 -11442
rect -802 -11498 -748 -11442
rect -692 -11498 -667 -11442
rect -1115 -11552 -667 -11498
rect -1115 -11608 -1086 -11552
rect -1030 -11608 -976 -11552
rect -920 -11608 -858 -11552
rect -802 -11608 -748 -11552
rect -692 -11608 -667 -11552
rect -1115 -11613 -667 -11608
rect 6933 -12350 7037 -10769
rect 8372 -11425 8592 -11416
rect 8372 -11481 8401 -11425
rect 8457 -11481 8511 -11425
rect 8567 -11481 8592 -11425
rect 8372 -11535 8592 -11481
rect 8372 -11591 8401 -11535
rect 8457 -11591 8511 -11535
rect 8567 -11591 8592 -11535
rect 8372 -11596 8592 -11591
rect 7129 -12111 7399 -12086
rect 7128 -12160 7399 -12111
rect 6865 -12363 7064 -12350
rect 6865 -12419 6882 -12363
rect 6938 -12419 6992 -12363
rect 7048 -12419 7064 -12363
rect 6865 -12436 7064 -12419
rect 7128 -12943 7232 -12160
rect 8458 -12274 8562 -11596
rect 8450 -12287 8649 -12274
rect 8450 -12343 8467 -12287
rect 8523 -12343 8577 -12287
rect 8633 -12343 8649 -12287
rect 8450 -12360 8649 -12343
rect 8912 -12347 9016 -10527
rect 10375 -11401 10595 -11392
rect 10375 -11457 10404 -11401
rect 10460 -11457 10514 -11401
rect 10570 -11457 10595 -11401
rect 10375 -11511 10595 -11457
rect 10375 -11567 10404 -11511
rect 10460 -11567 10514 -11511
rect 10570 -11567 10595 -11511
rect 10375 -11572 10595 -11567
rect 9150 -12160 9394 -12086
rect 8866 -12360 9065 -12347
rect 8866 -12416 8883 -12360
rect 8939 -12416 8993 -12360
rect 9049 -12416 9065 -12360
rect 8866 -12433 9065 -12416
rect 7127 -12960 7318 -12943
rect 7127 -13016 7132 -12960
rect 7188 -13016 7242 -12960
rect 7298 -13016 7318 -12960
rect 7127 -13037 7318 -13016
rect 9151 -13093 9255 -12160
rect 10443 -12274 10547 -11572
rect 10443 -12287 10642 -12274
rect 10443 -12343 10460 -12287
rect 10516 -12343 10570 -12287
rect 10626 -12343 10642 -12287
rect 10443 -12360 10642 -12343
rect 10947 -12350 11051 -10291
rect 12399 -11397 12619 -11388
rect 12399 -11453 12428 -11397
rect 12484 -11453 12538 -11397
rect 12594 -11453 12619 -11397
rect 12399 -11507 12619 -11453
rect 12399 -11563 12428 -11507
rect 12484 -11563 12538 -11507
rect 12594 -11563 12619 -11507
rect 12399 -11568 12619 -11563
rect 11172 -12109 11394 -12086
rect 11171 -12160 11394 -12109
rect 10443 -12368 10547 -12360
rect 10891 -12363 11090 -12350
rect 10891 -12419 10908 -12363
rect 10964 -12419 11018 -12363
rect 11074 -12419 11090 -12363
rect 10891 -12436 11090 -12419
rect 10947 -12438 11051 -12436
rect 7083 -13110 7274 -13093
rect 7083 -13166 7088 -13110
rect 7144 -13166 7198 -13110
rect 7254 -13166 7274 -13110
rect 7083 -13187 7274 -13166
rect 9151 -13110 9342 -13093
rect 9151 -13166 9156 -13110
rect 9212 -13166 9266 -13110
rect 9322 -13166 9342 -13110
rect 9151 -13187 9342 -13166
rect 6699 -13410 6890 -13393
rect 6699 -13466 6704 -13410
rect 6760 -13466 6814 -13410
rect 6870 -13466 6890 -13410
rect 6699 -13487 6890 -13466
rect 6459 -13710 6650 -13693
rect 6459 -13766 6464 -13710
rect 6520 -13766 6574 -13710
rect 6630 -13766 6650 -13710
rect 6459 -13787 6650 -13766
rect 6518 -15925 6613 -13787
rect 6712 -15358 6804 -13487
rect 7093 -14849 7159 -13187
rect 11171 -13243 11275 -12160
rect 12472 -12274 12576 -11568
rect 12472 -12287 12671 -12274
rect 12472 -12343 12489 -12287
rect 12545 -12343 12599 -12287
rect 12655 -12343 12671 -12287
rect 12472 -12360 12671 -12343
rect 12954 -12349 13058 -10046
rect 14433 -11388 14653 -11379
rect 14433 -11444 14462 -11388
rect 14518 -11444 14572 -11388
rect 14628 -11444 14653 -11388
rect 14433 -11498 14653 -11444
rect 14433 -11554 14462 -11498
rect 14518 -11554 14572 -11498
rect 14628 -11554 14653 -11498
rect 14433 -11559 14653 -11554
rect 13161 -12160 13394 -12086
rect 12472 -12364 12576 -12360
rect 12900 -12362 13099 -12349
rect 12900 -12418 12917 -12362
rect 12973 -12418 13027 -12362
rect 13083 -12418 13099 -12362
rect 12900 -12435 13099 -12418
rect 12954 -12443 13058 -12435
rect 11171 -13260 11362 -13243
rect 11171 -13316 11176 -13260
rect 11232 -13316 11286 -13260
rect 11342 -13316 11362 -13260
rect 11171 -13337 11362 -13316
rect 13161 -13393 13265 -12160
rect 14475 -12274 14579 -11559
rect 14475 -12287 14674 -12274
rect 14475 -12343 14492 -12287
rect 14548 -12343 14602 -12287
rect 14658 -12343 14674 -12287
rect 14475 -12360 14674 -12343
rect 14917 -12349 15021 -9804
rect 16429 -11387 16649 -11378
rect 16429 -11443 16458 -11387
rect 16514 -11443 16568 -11387
rect 16624 -11443 16649 -11387
rect 16429 -11497 16649 -11443
rect 16429 -11553 16458 -11497
rect 16514 -11553 16568 -11497
rect 16624 -11553 16649 -11497
rect 16429 -11558 16649 -11553
rect 15186 -12160 15401 -12086
rect 14475 -12363 14579 -12360
rect 14870 -12362 15069 -12349
rect 14870 -12418 14887 -12362
rect 14943 -12418 14997 -12362
rect 15053 -12418 15069 -12362
rect 14870 -12435 15069 -12418
rect 14917 -12440 15021 -12435
rect 13161 -13410 13352 -13393
rect 13161 -13466 13166 -13410
rect 13222 -13466 13276 -13410
rect 13332 -13466 13352 -13410
rect 13161 -13487 13352 -13466
rect 15188 -13543 15292 -12160
rect 16502 -12275 16606 -11558
rect 16490 -12288 16689 -12275
rect 16490 -12344 16507 -12288
rect 16563 -12344 16617 -12288
rect 16673 -12344 16689 -12288
rect 16490 -12361 16689 -12344
rect 16938 -12345 17042 -9562
rect 18419 -11384 18639 -11375
rect 18419 -11440 18448 -11384
rect 18504 -11440 18558 -11384
rect 18614 -11440 18639 -11384
rect 18419 -11494 18639 -11440
rect 18419 -11550 18448 -11494
rect 18504 -11550 18558 -11494
rect 18614 -11550 18639 -11494
rect 18419 -11555 18639 -11550
rect 17165 -12106 17394 -12086
rect 17164 -12160 17394 -12106
rect 16905 -12358 17104 -12345
rect 16502 -12365 16606 -12361
rect 16905 -12414 16922 -12358
rect 16978 -12414 17032 -12358
rect 17088 -12414 17104 -12358
rect 16905 -12431 17104 -12414
rect 15188 -13560 15379 -13543
rect 15188 -13616 15193 -13560
rect 15249 -13616 15303 -13560
rect 15359 -13616 15379 -13560
rect 15188 -13637 15379 -13616
rect 17164 -13693 17268 -12160
rect 18532 -12274 18636 -11555
rect 18511 -12287 18710 -12274
rect 18511 -12343 18528 -12287
rect 18584 -12343 18638 -12287
rect 18694 -12343 18710 -12287
rect 18511 -12360 18710 -12343
rect 18532 -12363 18636 -12360
rect 17440 -12960 17631 -12943
rect 17440 -13016 17445 -12960
rect 17501 -13016 17555 -12960
rect 17611 -13016 17631 -12960
rect 17440 -13037 17631 -13016
rect 17117 -13710 17308 -13693
rect 17117 -13766 17122 -13710
rect 17178 -13766 17232 -13710
rect 17288 -13766 17308 -13710
rect 17117 -13787 17308 -13766
rect 7042 -15058 7159 -14849
rect 7093 -15103 7159 -15058
rect 17440 -15103 17506 -13037
rect 17623 -13260 17808 -13243
rect 17623 -13316 17628 -13260
rect 17684 -13316 17738 -13260
rect 17794 -13316 17808 -13260
rect 17623 -13337 17808 -13316
rect 6712 -15450 6829 -15358
rect 17623 -15527 17689 -13337
rect 17780 -13553 17971 -13543
rect 17486 -15676 17689 -15527
rect 17779 -13560 17971 -13553
rect 17779 -13616 17785 -13560
rect 17841 -13616 17895 -13560
rect 17951 -13616 17971 -13560
rect 17779 -13637 17971 -13616
rect 17779 -15752 17874 -13637
rect 17663 -15847 17874 -15752
rect 6518 -15928 6674 -15925
rect 6518 -16023 6678 -15928
rect 18952 -16201 19286 -9045
rect 33938 -9391 34159 -9382
rect 33938 -9447 33967 -9391
rect 34023 -9447 34077 -9391
rect 34133 -9447 34159 -9391
rect 33938 -9501 34159 -9447
rect 33938 -9557 33967 -9501
rect 34023 -9557 34077 -9501
rect 34133 -9557 34159 -9501
rect 33938 -9562 34159 -9557
rect 31917 -9633 32138 -9624
rect 31917 -9689 31946 -9633
rect 32002 -9689 32056 -9633
rect 32112 -9689 32138 -9633
rect 31917 -9743 32138 -9689
rect 31917 -9799 31946 -9743
rect 32002 -9799 32056 -9743
rect 32112 -9799 32138 -9743
rect 31917 -9804 32138 -9799
rect 29954 -9875 30175 -9866
rect 29954 -9931 29983 -9875
rect 30039 -9931 30093 -9875
rect 30149 -9931 30175 -9875
rect 29954 -9985 30175 -9931
rect 29954 -10041 29983 -9985
rect 30039 -10041 30093 -9985
rect 30149 -10041 30175 -9985
rect 29954 -10046 30175 -10041
rect 27947 -10120 28168 -10111
rect 27947 -10176 27976 -10120
rect 28032 -10176 28086 -10120
rect 28142 -10176 28168 -10120
rect 27947 -10230 28168 -10176
rect 27947 -10286 27976 -10230
rect 28032 -10286 28086 -10230
rect 28142 -10286 28168 -10230
rect 27947 -10291 28168 -10286
rect 25912 -10356 26133 -10347
rect 25912 -10412 25941 -10356
rect 25997 -10412 26051 -10356
rect 26107 -10412 26133 -10356
rect 25912 -10466 26133 -10412
rect 25912 -10522 25941 -10466
rect 25997 -10522 26051 -10466
rect 26107 -10522 26133 -10466
rect 25912 -10527 26133 -10522
rect 23825 -10598 24046 -10589
rect 23825 -10654 23854 -10598
rect 23910 -10654 23964 -10598
rect 24020 -10654 24046 -10598
rect 23825 -10708 24046 -10654
rect 23825 -10764 23854 -10708
rect 23910 -10764 23964 -10708
rect 24020 -10764 24046 -10708
rect 23825 -10769 24046 -10764
rect 23933 -12350 24037 -10769
rect 25366 -10977 25587 -10968
rect 25366 -11033 25395 -10977
rect 25451 -11033 25505 -10977
rect 25561 -11033 25587 -10977
rect 25366 -11087 25587 -11033
rect 25366 -11143 25395 -11087
rect 25451 -11143 25505 -11087
rect 25561 -11143 25587 -11087
rect 25366 -11148 25587 -11143
rect 24129 -12111 24399 -12086
rect 24128 -12160 24399 -12111
rect 23865 -12363 24064 -12350
rect 23865 -12419 23882 -12363
rect 23938 -12419 23992 -12363
rect 24048 -12419 24064 -12363
rect 23865 -12436 24064 -12419
rect 24128 -12943 24232 -12160
rect 25458 -12274 25562 -11148
rect 25450 -12287 25649 -12274
rect 25450 -12343 25467 -12287
rect 25523 -12343 25577 -12287
rect 25633 -12343 25649 -12287
rect 25450 -12360 25649 -12343
rect 25912 -12347 26016 -10527
rect 27368 -10947 27589 -10938
rect 27368 -11003 27397 -10947
rect 27453 -11003 27507 -10947
rect 27563 -11003 27589 -10947
rect 27368 -11057 27589 -11003
rect 27368 -11113 27397 -11057
rect 27453 -11113 27507 -11057
rect 27563 -11113 27589 -11057
rect 27368 -11118 27589 -11113
rect 26150 -12160 26394 -12086
rect 25866 -12360 26065 -12347
rect 25866 -12416 25883 -12360
rect 25939 -12416 25993 -12360
rect 26049 -12416 26065 -12360
rect 25866 -12433 26065 -12416
rect 24127 -12960 24318 -12943
rect 24127 -13016 24132 -12960
rect 24188 -13016 24242 -12960
rect 24298 -13016 24318 -12960
rect 24127 -13037 24318 -13016
rect 26151 -13093 26255 -12160
rect 27443 -12274 27547 -11118
rect 27443 -12287 27642 -12274
rect 27443 -12343 27460 -12287
rect 27516 -12343 27570 -12287
rect 27626 -12343 27642 -12287
rect 27443 -12360 27642 -12343
rect 27947 -12350 28051 -10291
rect 29421 -10937 29642 -10928
rect 29421 -10993 29450 -10937
rect 29506 -10993 29560 -10937
rect 29616 -10993 29642 -10937
rect 29421 -11047 29642 -10993
rect 29421 -11103 29450 -11047
rect 29506 -11103 29560 -11047
rect 29616 -11103 29642 -11047
rect 29421 -11108 29642 -11103
rect 28172 -12109 28394 -12086
rect 28171 -12160 28394 -12109
rect 27443 -12368 27547 -12360
rect 27891 -12363 28090 -12350
rect 27891 -12419 27908 -12363
rect 27964 -12419 28018 -12363
rect 28074 -12419 28090 -12363
rect 27891 -12436 28090 -12419
rect 27947 -12438 28051 -12436
rect 24083 -13110 24274 -13093
rect 24083 -13166 24088 -13110
rect 24144 -13166 24198 -13110
rect 24254 -13166 24274 -13110
rect 24083 -13187 24274 -13166
rect 26151 -13110 26342 -13093
rect 26151 -13166 26156 -13110
rect 26212 -13166 26266 -13110
rect 26322 -13166 26342 -13110
rect 26151 -13187 26342 -13166
rect 23699 -13410 23890 -13393
rect 23699 -13466 23704 -13410
rect 23760 -13466 23814 -13410
rect 23870 -13466 23890 -13410
rect 23699 -13487 23890 -13466
rect 23459 -13710 23650 -13693
rect 23459 -13766 23464 -13710
rect 23520 -13766 23574 -13710
rect 23630 -13766 23650 -13710
rect 23459 -13787 23650 -13766
rect 23518 -15925 23613 -13787
rect 23712 -15358 23804 -13487
rect 24093 -14849 24159 -13187
rect 28171 -13243 28275 -12160
rect 29472 -12274 29576 -11108
rect 29472 -12287 29671 -12274
rect 29472 -12343 29489 -12287
rect 29545 -12343 29599 -12287
rect 29655 -12343 29671 -12287
rect 29472 -12360 29671 -12343
rect 29954 -12349 30058 -10046
rect 31424 -10933 31645 -10924
rect 31424 -10989 31453 -10933
rect 31509 -10989 31563 -10933
rect 31619 -10989 31645 -10933
rect 31424 -11043 31645 -10989
rect 31424 -11099 31453 -11043
rect 31509 -11099 31563 -11043
rect 31619 -11099 31645 -11043
rect 31424 -11104 31645 -11099
rect 30161 -12160 30394 -12086
rect 29472 -12364 29576 -12360
rect 29900 -12362 30099 -12349
rect 29900 -12418 29917 -12362
rect 29973 -12418 30027 -12362
rect 30083 -12418 30099 -12362
rect 29900 -12435 30099 -12418
rect 29954 -12443 30058 -12435
rect 28171 -13260 28362 -13243
rect 28171 -13316 28176 -13260
rect 28232 -13316 28286 -13260
rect 28342 -13316 28362 -13260
rect 28171 -13337 28362 -13316
rect 30161 -13393 30265 -12160
rect 31475 -12274 31579 -11104
rect 31475 -12287 31674 -12274
rect 31475 -12343 31492 -12287
rect 31548 -12343 31602 -12287
rect 31658 -12343 31674 -12287
rect 31475 -12360 31674 -12343
rect 31917 -12349 32021 -9804
rect 33477 -10933 33698 -10924
rect 33477 -10989 33506 -10933
rect 33562 -10989 33616 -10933
rect 33672 -10989 33698 -10933
rect 33477 -11043 33698 -10989
rect 33477 -11099 33506 -11043
rect 33562 -11099 33616 -11043
rect 33672 -11099 33698 -11043
rect 33477 -11104 33698 -11099
rect 32186 -12160 32401 -12086
rect 31475 -12363 31579 -12360
rect 31870 -12362 32069 -12349
rect 31870 -12418 31887 -12362
rect 31943 -12418 31997 -12362
rect 32053 -12418 32069 -12362
rect 31870 -12435 32069 -12418
rect 31917 -12440 32021 -12435
rect 30161 -13410 30352 -13393
rect 30161 -13466 30166 -13410
rect 30222 -13466 30276 -13410
rect 30332 -13466 30352 -13410
rect 30161 -13487 30352 -13466
rect 32188 -13543 32292 -12160
rect 33502 -12275 33606 -11104
rect 33490 -12288 33689 -12275
rect 33490 -12344 33507 -12288
rect 33563 -12344 33617 -12288
rect 33673 -12344 33689 -12288
rect 33490 -12361 33689 -12344
rect 33938 -12345 34042 -9562
rect 35528 -10933 35749 -10924
rect 35528 -10989 35557 -10933
rect 35613 -10989 35667 -10933
rect 35723 -10989 35749 -10933
rect 35528 -11043 35749 -10989
rect 35528 -11099 35557 -11043
rect 35613 -11099 35667 -11043
rect 35723 -11099 35749 -11043
rect 35528 -11104 35749 -11099
rect 34165 -12106 34394 -12086
rect 34164 -12160 34394 -12106
rect 33905 -12358 34104 -12345
rect 33502 -12365 33606 -12361
rect 33905 -12414 33922 -12358
rect 33978 -12414 34032 -12358
rect 34088 -12414 34104 -12358
rect 33905 -12431 34104 -12414
rect 32188 -13560 32379 -13543
rect 32188 -13616 32193 -13560
rect 32249 -13616 32303 -13560
rect 32359 -13616 32379 -13560
rect 32188 -13637 32379 -13616
rect 34164 -13693 34268 -12160
rect 35532 -12274 35636 -11104
rect 35511 -12287 35710 -12274
rect 35511 -12343 35528 -12287
rect 35584 -12343 35638 -12287
rect 35694 -12343 35710 -12287
rect 35511 -12360 35710 -12343
rect 35883 -12314 36082 -12301
rect 35532 -12363 35636 -12360
rect 35883 -12370 35900 -12314
rect 35956 -12370 36010 -12314
rect 36066 -12370 36082 -12314
rect 35883 -12387 36082 -12370
rect 34440 -12960 34631 -12943
rect 34440 -13016 34445 -12960
rect 34501 -13016 34555 -12960
rect 34611 -13016 34631 -12960
rect 34440 -13037 34631 -13016
rect 34117 -13710 34308 -13693
rect 34117 -13766 34122 -13710
rect 34178 -13766 34232 -13710
rect 34288 -13766 34308 -13710
rect 34117 -13787 34308 -13766
rect 24042 -15058 24159 -14849
rect 24093 -15103 24159 -15058
rect 34440 -15103 34506 -13037
rect 34623 -13260 34808 -13243
rect 34623 -13316 34628 -13260
rect 34684 -13316 34738 -13260
rect 34794 -13316 34808 -13260
rect 34623 -13337 34808 -13316
rect 23712 -15450 23829 -15358
rect 34623 -15527 34689 -13337
rect 34780 -13553 34971 -13543
rect 34486 -15676 34689 -15527
rect 34779 -13560 34971 -13553
rect 34779 -13616 34785 -13560
rect 34841 -13616 34895 -13560
rect 34951 -13616 34971 -13560
rect 34779 -13637 34971 -13616
rect 34779 -15752 34874 -13637
rect 34663 -15847 34874 -15752
rect 23518 -15928 23674 -15925
rect 23518 -16023 23678 -15928
rect 18952 -16257 18977 -16201
rect 19033 -16257 19087 -16201
rect 19143 -16257 19197 -16201
rect 19253 -16257 19286 -16201
rect 18952 -16311 19286 -16257
rect 18952 -16367 18977 -16311
rect 19033 -16367 19087 -16311
rect 19143 -16367 19197 -16311
rect 19253 -16367 19286 -16311
rect 18952 -16421 19286 -16367
rect 18952 -16477 18977 -16421
rect 19033 -16477 19087 -16421
rect 19143 -16477 19197 -16421
rect 19253 -16477 19286 -16421
rect 39179 -16138 39576 -8536
rect 54314 -9382 54424 -3642
rect 54527 -4444 54726 -4431
rect 54527 -4500 54544 -4444
rect 54600 -4500 54654 -4444
rect 54710 -4500 54726 -4444
rect 54527 -4517 54726 -4500
rect 54204 -9391 54425 -9382
rect 54204 -9447 54233 -9391
rect 54289 -9447 54343 -9391
rect 54399 -9447 54425 -9391
rect 54204 -9501 54425 -9447
rect 54204 -9557 54233 -9501
rect 54289 -9557 54343 -9501
rect 54399 -9557 54425 -9501
rect 54204 -9562 54425 -9557
rect 54527 -9624 54644 -4517
rect 54800 -5481 54999 -5468
rect 54800 -5537 54817 -5481
rect 54873 -5537 54927 -5481
rect 54983 -5537 54999 -5481
rect 54800 -5554 54999 -5537
rect 54423 -9633 54644 -9624
rect 54423 -9689 54452 -9633
rect 54508 -9689 54562 -9633
rect 54618 -9689 54644 -9633
rect 54423 -9743 54644 -9689
rect 54423 -9799 54452 -9743
rect 54508 -9799 54562 -9743
rect 54618 -9799 54644 -9743
rect 54423 -9804 54644 -9799
rect 54828 -9866 54910 -5554
rect 55049 -6355 55248 -6342
rect 55049 -6411 55066 -6355
rect 55122 -6411 55176 -6355
rect 55232 -6411 55248 -6355
rect 55049 -6428 55248 -6411
rect 54725 -9875 54946 -9866
rect 54725 -9931 54754 -9875
rect 54810 -9931 54864 -9875
rect 54920 -9931 54946 -9875
rect 54725 -9985 54946 -9931
rect 54725 -10041 54754 -9985
rect 54810 -10041 54864 -9985
rect 54920 -10041 54946 -9985
rect 54725 -10046 54946 -10041
rect 55090 -10111 55184 -6428
rect 55298 -7404 55497 -7391
rect 55298 -7460 55315 -7404
rect 55371 -7460 55425 -7404
rect 55481 -7460 55497 -7404
rect 55298 -7477 55497 -7460
rect 54961 -10120 55184 -10111
rect 54961 -10176 54990 -10120
rect 55046 -10176 55100 -10120
rect 55156 -10176 55184 -10120
rect 54961 -10230 55184 -10176
rect 54961 -10286 54990 -10230
rect 55046 -10286 55100 -10230
rect 55156 -10286 55184 -10230
rect 54961 -10290 55184 -10286
rect 54961 -10291 55182 -10290
rect 55321 -10347 55415 -7477
rect 55644 -8742 55843 -8729
rect 55644 -8798 55661 -8742
rect 55717 -8798 55771 -8742
rect 55827 -8798 55843 -8742
rect 55644 -8815 55843 -8798
rect 55222 -10356 55443 -10347
rect 55222 -10412 55251 -10356
rect 55307 -10412 55361 -10356
rect 55417 -10412 55443 -10356
rect 55222 -10466 55443 -10412
rect 55222 -10522 55251 -10466
rect 55307 -10522 55361 -10466
rect 55417 -10522 55443 -10466
rect 55222 -10527 55443 -10522
rect 55654 -10588 55748 -8815
rect 55539 -10597 55760 -10588
rect 55539 -10653 55568 -10597
rect 55624 -10653 55678 -10597
rect 55734 -10653 55760 -10597
rect 55539 -10707 55760 -10653
rect 55539 -10763 55568 -10707
rect 55624 -10763 55678 -10707
rect 55734 -10763 55760 -10707
rect 55539 -10768 55760 -10763
rect 59300 -11865 59356 -10203
rect 59564 -11544 59620 -10258
rect 59818 -11140 59874 -10134
rect 39179 -16194 39211 -16138
rect 39267 -16194 39321 -16138
rect 39377 -16194 39431 -16138
rect 39487 -16194 39576 -16138
rect 39179 -16248 39576 -16194
rect 39179 -16304 39211 -16248
rect 39267 -16304 39321 -16248
rect 39377 -16304 39431 -16248
rect 39487 -16304 39576 -16248
rect 39179 -16358 39576 -16304
rect 39179 -16414 39211 -16358
rect 39267 -16414 39321 -16358
rect 39377 -16414 39431 -16358
rect 39487 -16414 39576 -16358
rect 39179 -16430 39576 -16414
rect 18952 -16485 19286 -16477
<< via2 >>
rect 2685 5169 2741 5171
rect 2685 5117 2687 5169
rect 2687 5117 2739 5169
rect 2739 5117 2741 5169
rect 2685 5115 2741 5117
rect 2789 5169 2845 5171
rect 2789 5117 2791 5169
rect 2791 5117 2843 5169
rect 2843 5117 2845 5169
rect 2789 5115 2845 5117
rect 2685 5065 2741 5067
rect 2685 5013 2687 5065
rect 2687 5013 2739 5065
rect 2739 5013 2741 5065
rect 2685 5011 2741 5013
rect 2789 5065 2845 5067
rect 2789 5013 2791 5065
rect 2791 5013 2843 5065
rect 2843 5013 2845 5065
rect 2789 5011 2845 5013
rect 3474 5115 3530 5171
rect 3474 5065 3530 5067
rect 3474 5013 3476 5065
rect 3476 5013 3528 5065
rect 3528 5013 3530 5065
rect 3474 5011 3530 5013
rect 5255 5115 5311 5117
rect 5255 5063 5257 5115
rect 5257 5063 5309 5115
rect 5309 5063 5311 5115
rect 5255 5061 5311 5063
rect 5359 5115 5415 5117
rect 5359 5063 5361 5115
rect 5361 5063 5413 5115
rect 5413 5063 5415 5115
rect 5359 5061 5415 5063
rect 2044 4820 2100 4822
rect 2044 4768 2046 4820
rect 2046 4768 2098 4820
rect 2098 4768 2100 4820
rect 2044 4766 2100 4768
rect 2148 4820 2204 4822
rect 2148 4768 2150 4820
rect 2150 4768 2202 4820
rect 2202 4768 2204 4820
rect 2148 4766 2204 4768
rect 2044 4716 2100 4718
rect 2044 4664 2046 4716
rect 2046 4664 2098 4716
rect 2098 4664 2100 4716
rect 2044 4662 2100 4664
rect 2148 4716 2204 4718
rect 2148 4664 2150 4716
rect 2150 4664 2202 4716
rect 2202 4664 2204 4716
rect 2148 4662 2204 4664
rect -1761 -11074 -1705 -11018
rect -1651 -11074 -1595 -11018
rect -1524 -11073 -1468 -11017
rect -1414 -11073 -1358 -11017
rect -1761 -11184 -1705 -11128
rect -1651 -11184 -1595 -11128
rect -1524 -11183 -1468 -11127
rect -1414 -11183 -1358 -11127
rect 2405 4041 2461 4043
rect 2405 3989 2407 4041
rect 2407 3989 2459 4041
rect 2459 3989 2461 4041
rect 2405 3987 2461 3989
rect 2509 4041 2565 4043
rect 2509 3989 2511 4041
rect 2511 3989 2563 4041
rect 2563 3989 2565 4041
rect 2509 3987 2565 3989
rect 2405 3937 2461 3939
rect 2405 3885 2407 3937
rect 2407 3885 2459 3937
rect 2459 3885 2461 3937
rect 2405 3883 2461 3885
rect 2509 3937 2565 3939
rect 2509 3885 2511 3937
rect 2511 3885 2563 3937
rect 2563 3885 2565 3937
rect 2509 3883 2565 3885
rect 2044 3636 2100 3692
rect 2148 3636 2204 3692
rect 2044 3532 2100 3588
rect 2148 3532 2204 3588
rect 2044 1166 2100 1168
rect 2044 1114 2046 1166
rect 2046 1114 2098 1166
rect 2098 1114 2100 1166
rect 2044 1112 2100 1114
rect 2148 1166 2204 1168
rect 2148 1114 2150 1166
rect 2150 1114 2202 1166
rect 2202 1114 2204 1166
rect 2148 1112 2204 1114
rect 2044 1062 2100 1064
rect 2044 1010 2046 1062
rect 2046 1010 2098 1062
rect 2098 1010 2100 1062
rect 2044 1008 2100 1010
rect 2148 1062 2204 1064
rect 2148 1010 2150 1062
rect 2150 1010 2202 1062
rect 2202 1010 2204 1062
rect 2148 1008 2204 1010
rect 5255 5011 5311 5013
rect 5255 4959 5257 5011
rect 5257 4959 5309 5011
rect 5309 4959 5311 5011
rect 5255 4957 5311 4959
rect 5359 5011 5415 5013
rect 5359 4959 5361 5011
rect 5361 4959 5413 5011
rect 5413 4959 5415 5011
rect 5359 4957 5415 4959
rect 6259 5115 6315 5117
rect 6259 5063 6261 5115
rect 6261 5063 6313 5115
rect 6313 5063 6315 5115
rect 6259 5061 6315 5063
rect 6259 5011 6315 5013
rect 6259 4959 6261 5011
rect 6261 4959 6313 5011
rect 6313 4959 6315 5011
rect 6259 4957 6315 4959
rect 6899 5115 6955 5117
rect 6899 5063 6901 5115
rect 6901 5063 6953 5115
rect 6953 5063 6955 5115
rect 6899 5061 6955 5063
rect 6899 5011 6955 5013
rect 6899 4959 6901 5011
rect 6901 4959 6953 5011
rect 6953 4959 6955 5011
rect 6899 4957 6955 4959
rect 7539 5115 7595 5117
rect 7539 5063 7541 5115
rect 7541 5063 7593 5115
rect 7593 5063 7595 5115
rect 7539 5061 7595 5063
rect 7539 5011 7595 5013
rect 7539 4959 7541 5011
rect 7541 4959 7593 5011
rect 7593 4959 7595 5011
rect 7539 4957 7595 4959
rect 3554 4820 3610 4822
rect 3554 4768 3556 4820
rect 3556 4768 3608 4820
rect 3608 4768 3610 4820
rect 3554 4766 3610 4768
rect 3554 4716 3610 4718
rect 3554 4664 3556 4716
rect 3556 4664 3608 4716
rect 3608 4664 3610 4716
rect 3554 4662 3610 4664
rect 3714 4820 3770 4822
rect 3714 4768 3716 4820
rect 3716 4768 3768 4820
rect 3768 4768 3770 4820
rect 3714 4766 3770 4768
rect 3714 4716 3770 4718
rect 3714 4664 3716 4716
rect 3716 4664 3768 4716
rect 3768 4664 3770 4716
rect 3714 4662 3770 4664
rect 4355 4820 4411 4822
rect 4355 4768 4357 4820
rect 4357 4768 4409 4820
rect 4409 4768 4411 4820
rect 4355 4766 4411 4768
rect 4355 4716 4411 4718
rect 4355 4664 4357 4716
rect 4357 4664 4409 4716
rect 4409 4664 4411 4716
rect 4355 4662 4411 4664
rect 5527 4820 5583 4822
rect 5527 4768 5529 4820
rect 5529 4768 5581 4820
rect 5581 4768 5583 4820
rect 5527 4766 5583 4768
rect 5631 4820 5687 4822
rect 5631 4768 5633 4820
rect 5633 4768 5685 4820
rect 5685 4768 5687 4820
rect 5631 4766 5687 4768
rect 5527 4716 5583 4718
rect 5527 4664 5529 4716
rect 5529 4664 5581 4716
rect 5581 4664 5583 4716
rect 5527 4662 5583 4664
rect 5631 4716 5687 4718
rect 5631 4664 5633 4716
rect 5633 4664 5685 4716
rect 5685 4664 5687 4716
rect 5631 4662 5687 4664
rect 6579 4820 6635 4822
rect 6579 4768 6581 4820
rect 6581 4768 6633 4820
rect 6633 4768 6635 4820
rect 6579 4766 6635 4768
rect 6579 4716 6635 4718
rect 6579 4664 6581 4716
rect 6581 4664 6633 4716
rect 6633 4664 6635 4716
rect 6579 4662 6635 4664
rect 7219 4820 7275 4822
rect 7219 4768 7221 4820
rect 7221 4768 7273 4820
rect 7273 4768 7275 4820
rect 7219 4766 7275 4768
rect 7219 4716 7275 4718
rect 7219 4664 7221 4716
rect 7221 4664 7273 4716
rect 7273 4664 7275 4716
rect 7219 4662 7275 4664
rect 3394 4324 3450 4326
rect 3394 4272 3396 4324
rect 3396 4272 3448 4324
rect 3448 4272 3450 4324
rect 3394 4270 3450 4272
rect 3394 4220 3450 4222
rect 3394 4168 3396 4220
rect 3396 4168 3448 4220
rect 3448 4168 3450 4220
rect 3394 4166 3450 4168
rect 4034 4324 4090 4326
rect 4034 4272 4036 4324
rect 4036 4272 4088 4324
rect 4088 4272 4090 4324
rect 4034 4270 4090 4272
rect 4034 4220 4090 4222
rect 4034 4168 4036 4220
rect 4036 4168 4088 4220
rect 4088 4168 4090 4220
rect 4034 4166 4090 4168
rect 4674 4324 4730 4326
rect 4674 4272 4676 4324
rect 4676 4272 4728 4324
rect 4728 4272 4730 4324
rect 4674 4270 4730 4272
rect 4674 4220 4730 4222
rect 4674 4168 4676 4220
rect 4676 4168 4728 4220
rect 4728 4168 4730 4220
rect 4674 4166 4730 4168
rect 5255 4270 5311 4326
rect 5359 4270 5415 4326
rect 5255 4166 5311 4222
rect 5359 4166 5415 4222
rect 5255 4062 5311 4118
rect 5359 4062 5415 4118
rect 3474 4041 3530 4043
rect 3474 3989 3476 4041
rect 3476 3989 3528 4041
rect 3528 3989 3530 4041
rect 3474 3987 3530 3989
rect 3474 3937 3530 3939
rect 3474 3885 3476 3937
rect 3476 3885 3528 3937
rect 3528 3885 3530 3937
rect 3474 3883 3530 3885
rect 11163 4246 11219 4302
rect 11267 4246 11323 4302
rect 6579 4220 6635 4222
rect 6579 4168 6581 4220
rect 6581 4168 6633 4220
rect 6633 4168 6635 4220
rect 6579 4166 6635 4168
rect 6579 4116 6635 4118
rect 6579 4064 6581 4116
rect 6581 4064 6633 4116
rect 6633 4064 6635 4116
rect 6579 4062 6635 4064
rect 7219 4220 7275 4222
rect 7219 4168 7221 4220
rect 7221 4168 7273 4220
rect 7273 4168 7275 4220
rect 7219 4166 7275 4168
rect 11163 4142 11219 4198
rect 11267 4142 11323 4198
rect 17165 4194 17221 4250
rect 7219 4116 7275 4118
rect 7219 4064 7221 4116
rect 7221 4064 7273 4116
rect 7273 4064 7275 4116
rect 7219 4062 7275 4064
rect 5527 3787 5583 3843
rect 5631 3787 5687 3843
rect 3554 3690 3610 3692
rect 3554 3638 3556 3690
rect 3556 3638 3608 3690
rect 3608 3638 3610 3690
rect 3554 3636 3610 3638
rect 3554 3586 3610 3588
rect 3554 3534 3556 3586
rect 3556 3534 3608 3586
rect 3608 3534 3610 3586
rect 3554 3532 3610 3534
rect 3714 3690 3770 3692
rect 3714 3638 3716 3690
rect 3716 3638 3768 3690
rect 3768 3638 3770 3690
rect 3714 3636 3770 3638
rect 3714 3586 3770 3588
rect 3714 3534 3716 3586
rect 3716 3534 3768 3586
rect 3768 3534 3770 3586
rect 3714 3532 3770 3534
rect 4355 3690 4411 3692
rect 4355 3638 4357 3690
rect 4357 3638 4409 3690
rect 4409 3638 4411 3690
rect 4355 3636 4411 3638
rect 4355 3586 4411 3588
rect 4355 3534 4357 3586
rect 4357 3534 4409 3586
rect 4409 3534 4411 3586
rect 4355 3532 4411 3534
rect 5255 3636 5311 3692
rect 5359 3636 5415 3692
rect 5527 3683 5583 3739
rect 5631 3683 5687 3739
rect 6259 3841 6315 3843
rect 6259 3789 6261 3841
rect 6261 3789 6313 3841
rect 6313 3789 6315 3841
rect 6259 3787 6315 3789
rect 6259 3737 6315 3739
rect 6259 3685 6261 3737
rect 6261 3685 6313 3737
rect 6313 3685 6315 3737
rect 6259 3683 6315 3685
rect 6899 3841 6955 3843
rect 6899 3789 6901 3841
rect 6901 3789 6953 3841
rect 6953 3789 6955 3841
rect 6899 3787 6955 3789
rect 6899 3737 6955 3739
rect 6899 3685 6901 3737
rect 6901 3685 6953 3737
rect 6953 3685 6955 3737
rect 6899 3683 6955 3685
rect 7539 3841 7595 3843
rect 7539 3789 7541 3841
rect 7541 3789 7593 3841
rect 7593 3789 7595 3841
rect 7539 3787 7595 3789
rect 7539 3737 7595 3739
rect 7539 3685 7541 3737
rect 7541 3685 7593 3737
rect 7593 3685 7595 3737
rect 7539 3683 7595 3685
rect 5255 3532 5311 3588
rect 5359 3532 5415 3588
rect 3394 3298 3450 3300
rect 3394 3246 3396 3298
rect 3396 3246 3448 3298
rect 3448 3246 3450 3298
rect 3394 3244 3450 3246
rect 3394 3194 3450 3196
rect 3394 3142 3396 3194
rect 3396 3142 3448 3194
rect 3448 3142 3450 3194
rect 3394 3140 3450 3142
rect 4034 3298 4090 3300
rect 4034 3246 4036 3298
rect 4036 3246 4088 3298
rect 4088 3246 4090 3298
rect 4034 3244 4090 3246
rect 4034 3194 4090 3196
rect 4034 3142 4036 3194
rect 4036 3142 4088 3194
rect 4088 3142 4090 3194
rect 4034 3140 4090 3142
rect 4674 3298 4730 3300
rect 4674 3246 4676 3298
rect 4676 3246 4728 3298
rect 4728 3246 4730 3298
rect 4674 3244 4730 3246
rect 4674 3194 4730 3196
rect 4674 3142 4676 3194
rect 4676 3142 4728 3194
rect 4728 3142 4730 3194
rect 4674 3140 4730 3142
rect 5527 3244 5583 3300
rect 5631 3244 5687 3300
rect 5527 3140 5583 3196
rect 5631 3140 5687 3196
rect 6579 3298 6635 3300
rect 6579 3246 6581 3298
rect 6581 3246 6633 3298
rect 6633 3246 6635 3298
rect 6579 3244 6635 3246
rect 6579 3194 6635 3196
rect 6579 3142 6581 3194
rect 6581 3142 6633 3194
rect 6633 3142 6635 3194
rect 6579 3140 6635 3142
rect 7219 3298 7275 3300
rect 7219 3246 7221 3298
rect 7221 3246 7273 3298
rect 7273 3246 7275 3298
rect 7219 3244 7275 3246
rect 7219 3194 7275 3196
rect 7219 3142 7221 3194
rect 7221 3142 7273 3194
rect 7273 3142 7275 3194
rect 7219 3140 7275 3142
rect 10895 3280 10951 3336
rect 10999 3280 11055 3336
rect 10895 3176 10951 3232
rect 10999 3176 11055 3232
rect 5255 2925 5311 2981
rect 5359 2925 5415 2981
rect 2685 2857 2741 2913
rect 2789 2857 2845 2913
rect 2685 2753 2741 2809
rect 2789 2753 2845 2809
rect 3474 2911 3530 2913
rect 3474 2859 3476 2911
rect 3476 2859 3528 2911
rect 3528 2859 3530 2911
rect 3474 2857 3530 2859
rect 5255 2821 5311 2877
rect 5359 2821 5415 2877
rect 3474 2807 3530 2809
rect 3474 2755 3476 2807
rect 3476 2755 3528 2807
rect 3528 2755 3530 2807
rect 3474 2753 3530 2755
rect 2405 599 2461 655
rect 2509 599 2565 655
rect 2405 495 2461 551
rect 2509 495 2565 551
rect 2148 300 2204 302
rect 2148 248 2150 300
rect 2150 248 2202 300
rect 2202 248 2204 300
rect 2148 246 2204 248
rect 2148 196 2204 198
rect 2148 144 2150 196
rect 2150 144 2202 196
rect 2202 144 2204 196
rect 2148 142 2204 144
rect 2148 -1030 2204 -1028
rect 2148 -1082 2150 -1030
rect 2150 -1082 2202 -1030
rect 2202 -1082 2204 -1030
rect 2148 -1084 2204 -1082
rect 2148 -1134 2204 -1132
rect 2148 -1186 2150 -1134
rect 2150 -1186 2202 -1134
rect 2202 -1186 2204 -1134
rect 2148 -1188 2204 -1186
rect -250 -1574 -194 -1572
rect -250 -1626 -248 -1574
rect -248 -1626 -196 -1574
rect -196 -1626 -194 -1574
rect -250 -1628 -194 -1626
rect -146 -1574 -90 -1572
rect -146 -1626 -144 -1574
rect -144 -1626 -92 -1574
rect -92 -1626 -90 -1574
rect -146 -1628 -90 -1626
rect -250 -1678 -194 -1676
rect -250 -1730 -248 -1678
rect -248 -1730 -196 -1678
rect -196 -1730 -194 -1678
rect -250 -1732 -194 -1730
rect -146 -1678 -90 -1676
rect -146 -1730 -144 -1678
rect -144 -1730 -92 -1678
rect -92 -1730 -90 -1678
rect -146 -1732 -90 -1730
rect 751 -1574 807 -1572
rect 751 -1626 753 -1574
rect 753 -1626 805 -1574
rect 805 -1626 807 -1574
rect 751 -1628 807 -1626
rect 855 -1574 911 -1572
rect 855 -1626 857 -1574
rect 857 -1626 909 -1574
rect 909 -1626 911 -1574
rect 855 -1628 911 -1626
rect 3714 2560 3770 2562
rect 3714 2508 3716 2560
rect 3716 2508 3768 2560
rect 3768 2508 3770 2560
rect 3714 2506 3770 2508
rect 3714 2456 3770 2458
rect 3714 2404 3716 2456
rect 3716 2404 3768 2456
rect 3768 2404 3770 2456
rect 3714 2402 3770 2404
rect 4355 2560 4411 2562
rect 4355 2508 4357 2560
rect 4357 2508 4409 2560
rect 4409 2508 4411 2560
rect 4355 2506 4411 2508
rect 4355 2456 4411 2458
rect 4355 2404 4357 2456
rect 4357 2404 4409 2456
rect 4409 2404 4411 2456
rect 4355 2402 4411 2404
rect 6259 2979 6315 2981
rect 6259 2927 6261 2979
rect 6261 2927 6313 2979
rect 6313 2927 6315 2979
rect 6259 2925 6315 2927
rect 6259 2875 6315 2877
rect 6259 2823 6261 2875
rect 6261 2823 6313 2875
rect 6313 2823 6315 2875
rect 6259 2821 6315 2823
rect 6899 2979 6955 2981
rect 6899 2927 6901 2979
rect 6901 2927 6953 2979
rect 6953 2927 6955 2979
rect 6899 2925 6955 2927
rect 6899 2875 6955 2877
rect 6899 2823 6901 2875
rect 6901 2823 6953 2875
rect 6953 2823 6955 2875
rect 6899 2821 6955 2823
rect 7539 2979 7595 2981
rect 7539 2927 7541 2979
rect 7541 2927 7593 2979
rect 7593 2927 7595 2979
rect 7539 2925 7595 2927
rect 7539 2875 7595 2877
rect 7539 2823 7541 2875
rect 7541 2823 7593 2875
rect 7593 2823 7595 2875
rect 7539 2821 7595 2823
rect 5527 2506 5583 2562
rect 5631 2506 5687 2562
rect 5527 2402 5583 2458
rect 5631 2402 5687 2458
rect 5527 2298 5583 2354
rect 5631 2298 5687 2354
rect 6259 2456 6315 2458
rect 6259 2404 6261 2456
rect 6261 2404 6313 2456
rect 6313 2404 6315 2456
rect 6259 2402 6315 2404
rect 6259 2352 6315 2354
rect 6259 2300 6261 2352
rect 6261 2300 6313 2352
rect 6313 2300 6315 2352
rect 6259 2298 6315 2300
rect 6899 2456 6955 2458
rect 6899 2404 6901 2456
rect 6901 2404 6953 2456
rect 6953 2404 6955 2456
rect 6899 2402 6955 2404
rect 6899 2352 6955 2354
rect 6899 2300 6901 2352
rect 6901 2300 6953 2352
rect 6953 2300 6955 2352
rect 6899 2298 6955 2300
rect 7539 2456 7595 2458
rect 7539 2404 7541 2456
rect 7541 2404 7593 2456
rect 7593 2404 7595 2456
rect 7539 2402 7595 2404
rect 7539 2352 7595 2354
rect 7539 2300 7541 2352
rect 7541 2300 7593 2352
rect 7593 2300 7595 2352
rect 7539 2298 7595 2300
rect 5255 2114 5311 2170
rect 5359 2114 5415 2170
rect 3394 2064 3450 2066
rect 3394 2012 3396 2064
rect 3396 2012 3448 2064
rect 3448 2012 3450 2064
rect 3394 2010 3450 2012
rect 3394 1960 3450 1962
rect 3394 1908 3396 1960
rect 3396 1908 3448 1960
rect 3448 1908 3450 1960
rect 3394 1906 3450 1908
rect 4034 2064 4090 2066
rect 4034 2012 4036 2064
rect 4036 2012 4088 2064
rect 4088 2012 4090 2064
rect 4034 2010 4090 2012
rect 4034 1960 4090 1962
rect 4034 1908 4036 1960
rect 4036 1908 4088 1960
rect 4088 1908 4090 1960
rect 4034 1906 4090 1908
rect 4674 2064 4730 2066
rect 4674 2012 4676 2064
rect 4676 2012 4728 2064
rect 4728 2012 4730 2064
rect 4674 2010 4730 2012
rect 4674 1960 4730 1962
rect 4674 1908 4676 1960
rect 4676 1908 4728 1960
rect 4728 1908 4730 1960
rect 4674 1906 4730 1908
rect 5255 2010 5311 2066
rect 5359 2010 5415 2066
rect 5255 1906 5311 1962
rect 5359 1906 5415 1962
rect 5255 1583 5311 1639
rect 5359 1583 5415 1639
rect 5255 1479 5311 1535
rect 5359 1479 5415 1535
rect 3554 1166 3610 1168
rect 3554 1114 3556 1166
rect 3556 1114 3608 1166
rect 3608 1114 3610 1166
rect 3554 1112 3610 1114
rect 3554 1062 3610 1064
rect 3554 1010 3556 1062
rect 3556 1010 3608 1062
rect 3608 1010 3610 1062
rect 3554 1008 3610 1010
rect 3474 653 3530 655
rect 3474 601 3476 653
rect 3476 601 3528 653
rect 3528 601 3530 653
rect 3474 599 3530 601
rect 3474 549 3530 551
rect 3474 497 3476 549
rect 3476 497 3528 549
rect 3528 497 3530 549
rect 3474 495 3530 497
rect 6579 2168 6635 2170
rect 6579 2116 6581 2168
rect 6581 2116 6633 2168
rect 6633 2116 6635 2168
rect 6579 2114 6635 2116
rect 6579 2064 6635 2066
rect 6579 2012 6581 2064
rect 6581 2012 6633 2064
rect 6633 2012 6635 2064
rect 6579 2010 6635 2012
rect 7219 2168 7275 2170
rect 7219 2116 7221 2168
rect 7221 2116 7273 2168
rect 7273 2116 7275 2168
rect 7219 2114 7275 2116
rect 7219 2064 7275 2066
rect 7219 2012 7221 2064
rect 7221 2012 7273 2064
rect 7273 2012 7275 2064
rect 7219 2010 7275 2012
rect 10895 2216 10951 2218
rect 10895 2164 10897 2216
rect 10897 2164 10949 2216
rect 10949 2164 10951 2216
rect 10895 2162 10951 2164
rect 10999 2216 11055 2218
rect 10999 2164 11001 2216
rect 11001 2164 11053 2216
rect 11053 2164 11055 2216
rect 10999 2162 11055 2164
rect 10895 2112 10951 2114
rect 10895 2060 10897 2112
rect 10897 2060 10949 2112
rect 10949 2060 10951 2112
rect 10895 2058 10951 2060
rect 10999 2112 11055 2114
rect 10999 2060 11001 2112
rect 11001 2060 11053 2112
rect 11053 2060 11055 2112
rect 10999 2058 11055 2060
rect 8494 1637 8550 1639
rect 8494 1585 8496 1637
rect 8496 1585 8548 1637
rect 8548 1585 8550 1637
rect 8494 1583 8550 1585
rect 8494 1533 8550 1535
rect 8494 1481 8496 1533
rect 8496 1481 8548 1533
rect 8548 1481 8550 1533
rect 8494 1479 8550 1481
rect 9390 1637 9446 1639
rect 9390 1585 9392 1637
rect 9392 1585 9444 1637
rect 9444 1585 9446 1637
rect 9390 1583 9446 1585
rect 9390 1533 9446 1535
rect 9390 1481 9392 1533
rect 9392 1481 9444 1533
rect 9444 1481 9446 1533
rect 9390 1479 9446 1481
rect 10286 1637 10342 1639
rect 10286 1585 10288 1637
rect 10288 1585 10340 1637
rect 10340 1585 10342 1637
rect 10286 1583 10342 1585
rect 10286 1533 10342 1535
rect 10286 1481 10288 1533
rect 10288 1481 10340 1533
rect 10340 1481 10342 1533
rect 10286 1479 10342 1481
rect 5527 1212 5583 1268
rect 5631 1212 5687 1268
rect 5527 1108 5583 1164
rect 5631 1108 5687 1164
rect 8942 1266 8998 1268
rect 8942 1214 8944 1266
rect 8944 1214 8996 1266
rect 8996 1214 8998 1266
rect 8942 1212 8998 1214
rect 8942 1162 8998 1164
rect 8942 1110 8944 1162
rect 8944 1110 8996 1162
rect 8996 1110 8998 1162
rect 8942 1108 8998 1110
rect 9838 1266 9894 1268
rect 9838 1214 9840 1266
rect 9840 1214 9892 1266
rect 9892 1214 9894 1266
rect 9838 1212 9894 1214
rect 9838 1162 9894 1164
rect 9838 1110 9840 1162
rect 9840 1110 9892 1162
rect 9892 1110 9894 1162
rect 9838 1108 9894 1110
rect 10126 1266 10182 1268
rect 10126 1214 10128 1266
rect 10128 1214 10180 1266
rect 10180 1214 10182 1266
rect 10126 1212 10182 1214
rect 10126 1162 10182 1164
rect 10126 1110 10128 1162
rect 10128 1110 10180 1162
rect 10180 1110 10182 1162
rect 10126 1108 10182 1110
rect 5527 751 5583 807
rect 5631 751 5687 807
rect 5527 647 5583 703
rect 5631 647 5687 703
rect 6579 805 6635 807
rect 6579 753 6581 805
rect 6581 753 6633 805
rect 6633 753 6635 805
rect 6579 751 6635 753
rect 6579 701 6635 703
rect 6579 649 6581 701
rect 6581 649 6633 701
rect 6633 649 6635 701
rect 6579 647 6635 649
rect 7219 805 7275 807
rect 7219 753 7221 805
rect 7221 753 7273 805
rect 7273 753 7275 805
rect 7219 751 7275 753
rect 7219 701 7275 703
rect 7219 649 7221 701
rect 7221 649 7273 701
rect 7273 649 7275 701
rect 7219 647 7275 649
rect 5255 350 5311 406
rect 5359 350 5415 406
rect 3554 300 3610 302
rect 3554 248 3556 300
rect 3556 248 3608 300
rect 3608 248 3610 300
rect 3554 246 3610 248
rect 3554 196 3610 198
rect 3554 144 3556 196
rect 3556 144 3608 196
rect 3608 144 3610 196
rect 3554 142 3610 144
rect 3714 300 3770 302
rect 3714 248 3716 300
rect 3716 248 3768 300
rect 3768 248 3770 300
rect 3714 246 3770 248
rect 3714 196 3770 198
rect 3714 144 3716 196
rect 3716 144 3768 196
rect 3768 144 3770 196
rect 3714 142 3770 144
rect 4355 300 4411 302
rect 4355 248 4357 300
rect 4357 248 4409 300
rect 4409 248 4411 300
rect 4355 246 4411 248
rect 4355 196 4411 198
rect 4355 144 4357 196
rect 4357 144 4409 196
rect 4409 144 4411 196
rect 4355 142 4411 144
rect 5255 246 5311 302
rect 5359 246 5415 302
rect 5255 142 5311 198
rect 5359 142 5415 198
rect 3394 -196 3450 -194
rect 3394 -248 3396 -196
rect 3396 -248 3448 -196
rect 3448 -248 3450 -196
rect 3394 -250 3450 -248
rect 3394 -300 3450 -298
rect 3394 -352 3396 -300
rect 3396 -352 3448 -300
rect 3448 -352 3450 -300
rect 3394 -354 3450 -352
rect 4034 -196 4090 -194
rect 4034 -248 4036 -196
rect 4036 -248 4088 -196
rect 4088 -248 4090 -196
rect 4034 -250 4090 -248
rect 4034 -300 4090 -298
rect 4034 -352 4036 -300
rect 4036 -352 4088 -300
rect 4088 -352 4090 -300
rect 4034 -354 4090 -352
rect 4674 -196 4730 -194
rect 4674 -248 4676 -196
rect 4676 -248 4728 -196
rect 4728 -248 4730 -196
rect 4674 -250 4730 -248
rect 4674 -300 4730 -298
rect 4674 -352 4676 -300
rect 4676 -352 4728 -300
rect 4728 -352 4730 -300
rect 4674 -354 4730 -352
rect 18589 4248 18645 4250
rect 18589 4196 18591 4248
rect 18591 4196 18643 4248
rect 18643 4196 18645 4248
rect 18589 4194 18645 4196
rect 19709 4248 19765 4250
rect 19709 4196 19711 4248
rect 19711 4196 19763 4248
rect 19763 4196 19765 4248
rect 19709 4194 19765 4196
rect 23741 4248 23797 4250
rect 23741 4196 23743 4248
rect 23743 4196 23795 4248
rect 23795 4196 23797 4248
rect 23741 4194 23797 4196
rect 24861 4248 24917 4250
rect 24861 4196 24863 4248
rect 24863 4196 24915 4248
rect 24915 4196 24917 4248
rect 24861 4194 24917 4196
rect 26285 4194 26342 4250
rect 21621 4057 21677 4113
rect 21725 4057 21781 4113
rect 21829 4057 21885 4113
rect 18829 4007 18885 4009
rect 18829 3955 18831 4007
rect 18831 3955 18883 4007
rect 18883 3955 18885 4007
rect 18829 3953 18885 3955
rect 18829 3903 18885 3905
rect 18829 3851 18831 3903
rect 18831 3851 18883 3903
rect 18883 3851 18885 3903
rect 18829 3849 18885 3851
rect 19469 4007 19525 4009
rect 19469 3955 19471 4007
rect 19471 3955 19523 4007
rect 19523 3955 19525 4007
rect 19469 3953 19525 3955
rect 19469 3903 19525 3905
rect 19469 3851 19471 3903
rect 19471 3851 19523 3903
rect 19523 3851 19525 3903
rect 19469 3849 19525 3851
rect 21621 3953 21677 4009
rect 21725 3953 21781 4009
rect 21829 3953 21885 4009
rect 21621 3849 21677 3905
rect 21725 3849 21781 3905
rect 21829 3849 21885 3905
rect 20972 3663 21028 3719
rect 21076 3663 21132 3719
rect 21180 3663 21236 3719
rect 18509 3613 18565 3615
rect 18509 3561 18511 3613
rect 18511 3561 18563 3613
rect 18563 3561 18565 3613
rect 18509 3559 18565 3561
rect 18509 3509 18565 3511
rect 18509 3457 18511 3509
rect 18511 3457 18563 3509
rect 18563 3457 18565 3509
rect 18509 3455 18565 3457
rect 19149 3613 19205 3615
rect 19149 3561 19151 3613
rect 19151 3561 19203 3613
rect 19203 3561 19205 3613
rect 19149 3559 19205 3561
rect 19149 3509 19205 3511
rect 19149 3457 19151 3509
rect 19151 3457 19203 3509
rect 19203 3457 19205 3509
rect 19149 3455 19205 3457
rect 19789 3613 19845 3615
rect 19789 3561 19791 3613
rect 19791 3561 19843 3613
rect 19843 3561 19845 3613
rect 19789 3559 19845 3561
rect 19789 3509 19845 3511
rect 19789 3457 19791 3509
rect 19791 3457 19843 3509
rect 19843 3457 19845 3509
rect 19789 3455 19845 3457
rect 20972 3559 21028 3615
rect 21076 3559 21132 3615
rect 21180 3559 21236 3615
rect 20972 3455 21028 3511
rect 21076 3455 21132 3511
rect 21180 3455 21236 3511
rect 17165 2292 17221 2348
rect 12324 2216 12380 2218
rect 12324 2164 12326 2216
rect 12326 2164 12378 2216
rect 12378 2164 12380 2216
rect 12324 2162 12380 2164
rect 12324 2112 12380 2114
rect 12324 2060 12326 2112
rect 12326 2060 12378 2112
rect 12378 2060 12380 2112
rect 12324 2058 12380 2060
rect 13220 2216 13276 2218
rect 13220 2164 13222 2216
rect 13222 2164 13274 2216
rect 13274 2164 13276 2216
rect 13220 2162 13276 2164
rect 13220 2112 13276 2114
rect 13220 2060 13222 2112
rect 13222 2060 13274 2112
rect 13274 2060 13276 2112
rect 13220 2058 13276 2060
rect 13508 2216 13564 2218
rect 13508 2164 13510 2216
rect 13510 2164 13562 2216
rect 13562 2164 13564 2216
rect 13508 2162 13564 2164
rect 13508 2112 13564 2114
rect 13508 2060 13510 2112
rect 13510 2060 13562 2112
rect 13562 2060 13564 2112
rect 13508 2058 13564 2060
rect 14670 2216 14726 2218
rect 14670 2164 14672 2216
rect 14672 2164 14724 2216
rect 14724 2164 14726 2216
rect 14670 2162 14726 2164
rect 14670 2112 14726 2114
rect 14670 2060 14672 2112
rect 14672 2060 14724 2112
rect 14724 2060 14726 2112
rect 14670 2058 14726 2060
rect 15310 2216 15366 2218
rect 15310 2164 15312 2216
rect 15312 2164 15364 2216
rect 15364 2164 15366 2216
rect 15310 2162 15366 2164
rect 15310 2112 15366 2114
rect 15310 2060 15312 2112
rect 15312 2060 15364 2112
rect 15364 2060 15366 2112
rect 15310 2058 15366 2060
rect 15950 2216 16006 2218
rect 15950 2164 15952 2216
rect 15952 2164 16004 2216
rect 16004 2164 16006 2216
rect 15950 2162 16006 2164
rect 15950 2112 16006 2114
rect 15950 2060 15952 2112
rect 15952 2060 16004 2112
rect 16004 2060 16006 2112
rect 15950 2058 16006 2060
rect 16889 2216 16945 2218
rect 16889 2164 16891 2216
rect 16891 2164 16943 2216
rect 16943 2164 16945 2216
rect 16889 2162 16945 2164
rect 16993 2216 17049 2218
rect 16993 2164 16995 2216
rect 16995 2164 17047 2216
rect 17047 2164 17049 2216
rect 16993 2162 17049 2164
rect 16889 2112 16945 2114
rect 16889 2060 16891 2112
rect 16891 2060 16943 2112
rect 16943 2060 16945 2112
rect 16889 2058 16945 2060
rect 16993 2112 17049 2114
rect 16993 2060 16995 2112
rect 16995 2060 17047 2112
rect 17047 2060 17049 2112
rect 16993 2058 17049 2060
rect 11163 1796 11219 1798
rect 11163 1744 11165 1796
rect 11165 1744 11217 1796
rect 11217 1744 11219 1796
rect 11163 1742 11219 1744
rect 11267 1796 11323 1798
rect 11267 1744 11269 1796
rect 11269 1744 11321 1796
rect 11321 1744 11323 1796
rect 11267 1742 11323 1744
rect 11163 1692 11219 1694
rect 11163 1640 11165 1692
rect 11165 1640 11217 1692
rect 11217 1640 11219 1692
rect 11163 1638 11219 1640
rect 11267 1692 11323 1694
rect 11267 1640 11269 1692
rect 11269 1640 11321 1692
rect 11321 1640 11323 1692
rect 11267 1638 11323 1640
rect 11876 1796 11932 1798
rect 11876 1744 11878 1796
rect 11878 1744 11930 1796
rect 11930 1744 11932 1796
rect 11876 1742 11932 1744
rect 11876 1692 11932 1694
rect 11876 1640 11878 1692
rect 11878 1640 11930 1692
rect 11930 1640 11932 1692
rect 11876 1638 11932 1640
rect 12772 1796 12828 1798
rect 12772 1744 12774 1796
rect 12774 1744 12826 1796
rect 12826 1744 12828 1796
rect 12772 1742 12828 1744
rect 12772 1692 12828 1694
rect 12772 1640 12774 1692
rect 12774 1640 12826 1692
rect 12826 1640 12828 1692
rect 12772 1638 12828 1640
rect 13668 1796 13724 1798
rect 13668 1744 13670 1796
rect 13670 1744 13722 1796
rect 13722 1744 13724 1796
rect 13668 1742 13724 1744
rect 13668 1692 13724 1694
rect 13668 1640 13670 1692
rect 13670 1640 13722 1692
rect 13722 1640 13724 1692
rect 13668 1638 13724 1640
rect 14990 1796 15046 1798
rect 14990 1744 14992 1796
rect 14992 1744 15044 1796
rect 15044 1744 15046 1796
rect 14990 1742 15046 1744
rect 14990 1692 15046 1694
rect 14990 1640 14992 1692
rect 14992 1640 15044 1692
rect 15044 1640 15046 1692
rect 14990 1638 15046 1640
rect 15630 1796 15686 1798
rect 15630 1744 15632 1796
rect 15632 1744 15684 1796
rect 15684 1744 15686 1796
rect 15630 1742 15686 1744
rect 15630 1692 15686 1694
rect 15630 1640 15632 1692
rect 15632 1640 15684 1692
rect 15684 1640 15686 1692
rect 15630 1638 15686 1640
rect 16627 1796 16683 1798
rect 16627 1744 16629 1796
rect 16629 1744 16681 1796
rect 16681 1744 16683 1796
rect 16627 1742 16683 1744
rect 16731 1796 16787 1798
rect 16731 1744 16733 1796
rect 16733 1744 16785 1796
rect 16785 1744 16787 1796
rect 16731 1742 16787 1744
rect 16627 1692 16683 1694
rect 16627 1640 16629 1692
rect 16629 1640 16681 1692
rect 16681 1640 16683 1692
rect 16627 1638 16683 1640
rect 16731 1692 16787 1694
rect 16731 1640 16733 1692
rect 16733 1640 16785 1692
rect 16785 1640 16787 1692
rect 16731 1638 16787 1640
rect 11163 1212 11219 1268
rect 11267 1212 11323 1268
rect 11163 1108 11219 1164
rect 11267 1108 11323 1164
rect 11163 1004 11219 1060
rect 11267 1004 11323 1060
rect 12324 1162 12380 1164
rect 12324 1110 12326 1162
rect 12326 1110 12378 1162
rect 12378 1110 12380 1162
rect 12324 1108 12380 1110
rect 12324 1058 12380 1060
rect 12324 1006 12326 1058
rect 12326 1006 12378 1058
rect 12378 1006 12380 1058
rect 12324 1004 12380 1006
rect 13220 1162 13276 1164
rect 13220 1110 13222 1162
rect 13222 1110 13274 1162
rect 13274 1110 13276 1162
rect 13220 1108 13276 1110
rect 13220 1058 13276 1060
rect 13220 1006 13222 1058
rect 13222 1006 13274 1058
rect 13274 1006 13276 1058
rect 13220 1004 13276 1006
rect 13508 1136 13564 1138
rect 13508 1084 13510 1136
rect 13510 1084 13562 1136
rect 13562 1084 13564 1136
rect 13508 1082 13564 1084
rect 10126 604 10182 606
rect 10126 552 10128 604
rect 10128 552 10180 604
rect 10180 552 10182 604
rect 10126 550 10182 552
rect 10126 500 10182 502
rect 10126 448 10128 500
rect 10128 448 10180 500
rect 10180 448 10182 500
rect 10126 446 10182 448
rect 10895 550 10951 606
rect 10999 550 11055 606
rect 10895 446 10951 502
rect 10999 446 11055 502
rect 6259 404 6315 406
rect 6259 352 6261 404
rect 6261 352 6313 404
rect 6313 352 6315 404
rect 6259 350 6315 352
rect 6259 300 6315 302
rect 6259 248 6261 300
rect 6261 248 6313 300
rect 6313 248 6315 300
rect 6259 246 6315 248
rect 6899 404 6955 406
rect 6899 352 6901 404
rect 6901 352 6953 404
rect 6953 352 6955 404
rect 6899 350 6955 352
rect 6899 300 6955 302
rect 6899 248 6901 300
rect 6901 248 6953 300
rect 6953 248 6955 300
rect 6899 246 6955 248
rect 7539 404 7595 406
rect 7539 352 7541 404
rect 7541 352 7593 404
rect 7593 352 7595 404
rect 7539 350 7595 352
rect 7539 300 7595 302
rect 7539 248 7541 300
rect 7541 248 7593 300
rect 7593 248 7595 300
rect 7539 246 7595 248
rect 8942 404 8998 406
rect 8942 352 8944 404
rect 8944 352 8996 404
rect 8996 352 8998 404
rect 8942 350 8998 352
rect 8942 300 8998 302
rect 8942 248 8944 300
rect 8944 248 8996 300
rect 8996 248 8998 300
rect 8942 246 8998 248
rect 9838 404 9894 406
rect 9838 352 9840 404
rect 9840 352 9892 404
rect 9892 352 9894 404
rect 9838 350 9894 352
rect 9838 300 9894 302
rect 9838 248 9840 300
rect 9840 248 9892 300
rect 9892 248 9894 300
rect 9838 246 9894 248
rect 10895 62 10951 118
rect 10999 62 11055 118
rect 10895 -42 10951 14
rect 10999 -42 11055 14
rect 5527 -250 5583 -194
rect 5631 -250 5687 -194
rect 5527 -354 5583 -298
rect 5631 -354 5687 -298
rect 6259 -196 6315 -194
rect 6259 -248 6261 -196
rect 6261 -248 6313 -196
rect 6313 -248 6315 -196
rect 6259 -250 6315 -248
rect 6259 -300 6315 -298
rect 6259 -352 6261 -300
rect 6261 -352 6313 -300
rect 6313 -352 6315 -300
rect 6259 -354 6315 -352
rect 6899 -196 6955 -194
rect 6899 -248 6901 -196
rect 6901 -248 6953 -196
rect 6953 -248 6955 -196
rect 6899 -250 6955 -248
rect 6899 -300 6955 -298
rect 6899 -352 6901 -300
rect 6901 -352 6953 -300
rect 6953 -352 6955 -300
rect 6899 -354 6955 -352
rect 7539 -196 7595 -194
rect 7539 -248 7541 -196
rect 7541 -248 7593 -196
rect 7593 -248 7595 -196
rect 7539 -250 7595 -248
rect 7539 -300 7595 -298
rect 7539 -352 7541 -300
rect 7541 -352 7593 -300
rect 7593 -352 7595 -300
rect 7539 -354 7595 -352
rect 8494 -196 8550 -194
rect 8494 -248 8496 -196
rect 8496 -248 8548 -196
rect 8548 -248 8550 -196
rect 8494 -250 8550 -248
rect 8494 -300 8550 -298
rect 8494 -352 8496 -300
rect 8496 -352 8548 -300
rect 8548 -352 8550 -300
rect 8494 -354 8550 -352
rect 9390 -196 9446 -194
rect 9390 -248 9392 -196
rect 9392 -248 9444 -196
rect 9444 -248 9446 -196
rect 9390 -250 9446 -248
rect 9390 -300 9446 -298
rect 9390 -352 9392 -300
rect 9392 -352 9444 -300
rect 9444 -352 9446 -300
rect 9390 -354 9446 -352
rect 10286 -196 10342 -194
rect 10286 -248 10288 -196
rect 10288 -248 10340 -196
rect 10340 -248 10342 -196
rect 10286 -250 10342 -248
rect 10286 -300 10342 -298
rect 10286 -352 10288 -300
rect 10288 -352 10340 -300
rect 10340 -352 10342 -300
rect 10286 -354 10342 -352
rect 2685 -531 2741 -475
rect 2789 -531 2845 -475
rect 2685 -635 2741 -579
rect 2789 -635 2845 -579
rect 3474 -477 3530 -475
rect 3474 -529 3476 -477
rect 3476 -529 3528 -477
rect 3528 -529 3530 -477
rect 3474 -531 3530 -529
rect 3474 -581 3530 -579
rect 3474 -633 3476 -581
rect 3476 -633 3528 -581
rect 3528 -633 3530 -581
rect 3474 -635 3530 -633
rect 5255 -523 5311 -467
rect 5359 -523 5415 -467
rect 5255 -627 5311 -571
rect 5359 -627 5415 -571
rect 3714 -830 3770 -828
rect 3714 -882 3716 -830
rect 3716 -882 3768 -830
rect 3768 -882 3770 -830
rect 3714 -884 3770 -882
rect 3714 -934 3770 -932
rect 3714 -986 3716 -934
rect 3716 -986 3768 -934
rect 3768 -986 3770 -934
rect 3714 -988 3770 -986
rect 4355 -830 4411 -828
rect 4355 -882 4357 -830
rect 4357 -882 4409 -830
rect 4409 -882 4411 -830
rect 4355 -884 4411 -882
rect 4355 -934 4411 -932
rect 4355 -986 4357 -934
rect 4357 -986 4409 -934
rect 4409 -986 4411 -934
rect 4355 -988 4411 -986
rect 3554 -1030 3610 -1028
rect 3554 -1082 3556 -1030
rect 3556 -1082 3608 -1030
rect 3608 -1082 3610 -1030
rect 3554 -1084 3610 -1082
rect 3554 -1134 3610 -1132
rect 3554 -1186 3556 -1134
rect 3556 -1186 3608 -1134
rect 3608 -1186 3610 -1134
rect 3554 -1188 3610 -1186
rect 6579 -469 6635 -467
rect 6579 -521 6581 -469
rect 6581 -521 6633 -469
rect 6633 -521 6635 -469
rect 6579 -523 6635 -521
rect 6579 -573 6635 -571
rect 6579 -625 6581 -573
rect 6581 -625 6633 -573
rect 6633 -625 6635 -573
rect 6579 -627 6635 -625
rect 7219 -469 7275 -467
rect 7219 -521 7221 -469
rect 7221 -521 7273 -469
rect 7273 -521 7275 -469
rect 7219 -523 7275 -521
rect 7219 -573 7275 -571
rect 7219 -625 7221 -573
rect 7221 -625 7273 -573
rect 7273 -625 7275 -573
rect 7219 -627 7275 -625
rect 9998 -454 10054 -452
rect 9998 -506 10000 -454
rect 10000 -506 10052 -454
rect 10052 -506 10054 -454
rect 9998 -508 10054 -506
rect 9998 -558 10054 -556
rect 9998 -610 10000 -558
rect 10000 -610 10052 -558
rect 10052 -610 10054 -558
rect 9998 -612 10054 -610
rect 7513 -693 7569 -691
rect 7513 -745 7515 -693
rect 7515 -745 7567 -693
rect 7567 -745 7569 -693
rect 7513 -747 7569 -745
rect 5527 -884 5583 -828
rect 5631 -884 5687 -828
rect 7513 -797 7569 -795
rect 7513 -849 7515 -797
rect 7515 -849 7567 -797
rect 7567 -849 7569 -797
rect 7513 -851 7569 -849
rect 7799 -747 7855 -691
rect 7903 -747 7959 -691
rect 7799 -851 7855 -795
rect 7903 -851 7959 -795
rect 10246 -704 10302 -702
rect 10246 -756 10248 -704
rect 10248 -756 10300 -704
rect 10300 -756 10302 -704
rect 10246 -758 10302 -756
rect 5527 -988 5583 -932
rect 5631 -988 5687 -932
rect 5527 -1092 5583 -1036
rect 5631 -1092 5687 -1036
rect 6579 -934 6635 -932
rect 6579 -986 6581 -934
rect 6581 -986 6633 -934
rect 6633 -986 6635 -934
rect 6579 -988 6635 -986
rect 6579 -1038 6635 -1036
rect 6579 -1090 6581 -1038
rect 6581 -1090 6633 -1038
rect 6633 -1090 6635 -1038
rect 6579 -1092 6635 -1090
rect 7219 -934 7275 -932
rect 7219 -986 7221 -934
rect 7221 -986 7273 -934
rect 7273 -986 7275 -934
rect 7219 -988 7275 -986
rect 7219 -1038 7275 -1036
rect 7219 -1090 7221 -1038
rect 7221 -1090 7273 -1038
rect 7273 -1090 7275 -1038
rect 7219 -1092 7275 -1090
rect 3394 -1326 3450 -1324
rect 3394 -1378 3396 -1326
rect 3396 -1378 3448 -1326
rect 3448 -1378 3450 -1326
rect 3394 -1380 3450 -1378
rect 3394 -1430 3450 -1428
rect 3394 -1482 3396 -1430
rect 3396 -1482 3448 -1430
rect 3448 -1482 3450 -1430
rect 3394 -1484 3450 -1482
rect 4034 -1326 4090 -1324
rect 4034 -1378 4036 -1326
rect 4036 -1378 4088 -1326
rect 4088 -1378 4090 -1326
rect 4034 -1380 4090 -1378
rect 4034 -1430 4090 -1428
rect 4034 -1482 4036 -1430
rect 4036 -1482 4088 -1430
rect 4088 -1482 4090 -1430
rect 4034 -1484 4090 -1482
rect 4674 -1326 4730 -1324
rect 4674 -1378 4676 -1326
rect 4676 -1378 4728 -1326
rect 4728 -1378 4730 -1326
rect 4674 -1380 4730 -1378
rect 4674 -1430 4730 -1428
rect 4674 -1482 4676 -1430
rect 4676 -1482 4728 -1430
rect 4728 -1482 4730 -1430
rect 4674 -1484 4730 -1482
rect 5255 -1380 5311 -1324
rect 5359 -1380 5415 -1324
rect 5255 -1484 5311 -1428
rect 5359 -1484 5415 -1428
rect 6259 -1326 6315 -1324
rect 6259 -1378 6261 -1326
rect 6261 -1378 6313 -1326
rect 6313 -1378 6315 -1326
rect 6259 -1380 6315 -1378
rect 6259 -1430 6315 -1428
rect 6259 -1482 6261 -1430
rect 6261 -1482 6313 -1430
rect 6313 -1482 6315 -1430
rect 6259 -1484 6315 -1482
rect 6899 -1326 6955 -1324
rect 6899 -1378 6901 -1326
rect 6901 -1378 6953 -1326
rect 6953 -1378 6955 -1326
rect 6899 -1380 6955 -1378
rect 6899 -1430 6955 -1428
rect 6899 -1482 6901 -1430
rect 6901 -1482 6953 -1430
rect 6953 -1482 6955 -1430
rect 6899 -1484 6955 -1482
rect 7539 -1326 7595 -1324
rect 7539 -1378 7541 -1326
rect 7541 -1378 7593 -1326
rect 7593 -1378 7595 -1326
rect 7539 -1380 7595 -1378
rect 7539 -1430 7595 -1428
rect 7539 -1482 7541 -1430
rect 7541 -1482 7593 -1430
rect 7593 -1482 7595 -1430
rect 7539 -1484 7595 -1482
rect 751 -1732 807 -1676
rect 855 -1732 911 -1676
rect 2405 -1719 2461 -1663
rect 2509 -1719 2565 -1663
rect 2405 -1823 2461 -1767
rect 2509 -1823 2565 -1767
rect 3634 -1665 3690 -1663
rect 3634 -1717 3636 -1665
rect 3636 -1717 3688 -1665
rect 3688 -1717 3690 -1665
rect 3634 -1719 3690 -1717
rect 3634 -1823 3690 -1767
rect 10246 -808 10302 -806
rect 10246 -860 10248 -808
rect 10248 -860 10300 -808
rect 10300 -860 10302 -808
rect 10246 -862 10302 -860
rect 10442 -758 10498 -702
rect 10546 -758 10602 -702
rect 10442 -862 10498 -806
rect 10546 -862 10602 -806
rect 8942 -934 8998 -932
rect 8942 -986 8944 -934
rect 8944 -986 8996 -934
rect 8996 -986 8998 -934
rect 8942 -988 8998 -986
rect 8942 -1038 8998 -1036
rect 8942 -1090 8944 -1038
rect 8944 -1090 8996 -1038
rect 8996 -1090 8998 -1038
rect 8942 -1092 8998 -1090
rect 9838 -934 9894 -932
rect 9838 -986 9840 -934
rect 9840 -986 9892 -934
rect 9892 -986 9894 -934
rect 9838 -988 9894 -986
rect 9838 -1038 9894 -1036
rect 9838 -1090 9840 -1038
rect 9840 -1090 9892 -1038
rect 9892 -1090 9894 -1038
rect 9838 -1092 9894 -1090
rect 9998 -934 10054 -932
rect 9998 -986 10000 -934
rect 10000 -986 10052 -934
rect 10052 -986 10054 -934
rect 9998 -988 10054 -986
rect 9998 -1038 10054 -1036
rect 9998 -1090 10000 -1038
rect 10000 -1090 10052 -1038
rect 10052 -1090 10054 -1038
rect 9998 -1092 10054 -1090
rect 8494 -1326 8550 -1324
rect 8494 -1378 8496 -1326
rect 8496 -1378 8548 -1326
rect 8548 -1378 8550 -1326
rect 8494 -1380 8550 -1378
rect 8494 -1430 8550 -1428
rect 8494 -1482 8496 -1430
rect 8496 -1482 8548 -1430
rect 8548 -1482 8550 -1430
rect 8494 -1484 8550 -1482
rect 9390 -1326 9446 -1324
rect 9390 -1378 9392 -1326
rect 9392 -1378 9444 -1326
rect 9444 -1378 9446 -1326
rect 9390 -1380 9446 -1378
rect 9390 -1430 9446 -1428
rect 9390 -1482 9392 -1430
rect 9392 -1482 9444 -1430
rect 9444 -1482 9446 -1430
rect 9390 -1484 9446 -1482
rect 10286 -1326 10342 -1324
rect 10286 -1378 10288 -1326
rect 10288 -1378 10340 -1326
rect 10340 -1378 10342 -1326
rect 10286 -1380 10342 -1378
rect 10286 -1430 10342 -1428
rect 10286 -1482 10288 -1430
rect 10288 -1482 10340 -1430
rect 10340 -1482 10342 -1430
rect 10286 -1484 10342 -1482
rect 6906 -2802 6962 -2746
rect 7010 -2802 7066 -2746
rect 6906 -2906 6962 -2850
rect 7010 -2906 7066 -2850
rect 7799 -2748 7855 -2746
rect 7799 -2800 7801 -2748
rect 7801 -2800 7853 -2748
rect 7853 -2800 7855 -2748
rect 7799 -2802 7855 -2800
rect 7903 -2748 7959 -2746
rect 7903 -2800 7905 -2748
rect 7905 -2800 7957 -2748
rect 7957 -2800 7959 -2748
rect 7903 -2802 7959 -2800
rect 7799 -2852 7855 -2850
rect 7799 -2904 7801 -2852
rect 7801 -2904 7853 -2852
rect 7853 -2904 7855 -2852
rect 7799 -2906 7855 -2904
rect 7903 -2852 7959 -2850
rect 7903 -2904 7905 -2852
rect 7905 -2904 7957 -2852
rect 7957 -2904 7959 -2852
rect 7903 -2906 7959 -2904
rect 2571 -3984 2627 -3982
rect 2571 -4036 2573 -3984
rect 2573 -4036 2625 -3984
rect 2625 -4036 2627 -3984
rect 2571 -4038 2627 -4036
rect 2675 -3984 2731 -3982
rect 2675 -4036 2677 -3984
rect 2677 -4036 2729 -3984
rect 2729 -4036 2731 -3984
rect 2675 -4038 2731 -4036
rect 2571 -4088 2627 -4086
rect 2571 -4140 2573 -4088
rect 2573 -4140 2625 -4088
rect 2625 -4140 2627 -4088
rect 2571 -4142 2627 -4140
rect 2675 -4088 2731 -4086
rect 2675 -4140 2677 -4088
rect 2677 -4140 2729 -4088
rect 2729 -4140 2731 -4088
rect 2675 -4142 2731 -4140
rect 2239 -4738 2295 -4736
rect 2239 -4790 2241 -4738
rect 2241 -4790 2293 -4738
rect 2293 -4790 2295 -4738
rect 2239 -4792 2295 -4790
rect 2239 -4842 2295 -4840
rect 2239 -4894 2241 -4842
rect 2241 -4894 2293 -4842
rect 2293 -4894 2295 -4842
rect 2239 -4896 2295 -4894
rect 3535 -5028 3591 -5026
rect 3535 -5080 3537 -5028
rect 3537 -5080 3589 -5028
rect 3589 -5080 3591 -5028
rect 3535 -5082 3591 -5080
rect 3535 -5132 3591 -5130
rect 3535 -5184 3537 -5132
rect 3537 -5184 3589 -5132
rect 3589 -5184 3591 -5132
rect 3535 -5186 3591 -5184
rect 3103 -5352 3159 -5350
rect 3103 -5404 3105 -5352
rect 3105 -5404 3157 -5352
rect 3157 -5404 3159 -5352
rect 3103 -5406 3159 -5404
rect 3103 -5456 3159 -5454
rect 3103 -5508 3105 -5456
rect 3105 -5508 3157 -5456
rect 3157 -5508 3159 -5456
rect 3103 -5510 3159 -5508
rect 2943 -5808 2999 -5752
rect 3047 -5808 3103 -5752
rect 2943 -5912 2999 -5856
rect 3047 -5912 3103 -5856
rect 751 -6052 807 -5996
rect 855 -6052 911 -5996
rect 751 -6156 807 -6100
rect 855 -6156 911 -6100
rect 2249 -5998 2305 -5996
rect 2249 -6050 2251 -5998
rect 2251 -6050 2303 -5998
rect 2303 -6050 2305 -5998
rect 2249 -6052 2305 -6050
rect 2249 -6102 2305 -6100
rect 2249 -6154 2251 -6102
rect 2251 -6154 2303 -6102
rect 2303 -6154 2305 -6102
rect 2249 -6156 2305 -6154
rect 5144 -4792 5200 -4736
rect 5248 -4792 5304 -4736
rect 5144 -4896 5200 -4840
rect 5248 -4896 5304 -4840
rect 4908 -5406 4964 -5350
rect 5012 -5406 5068 -5350
rect 4908 -5510 4964 -5454
rect 5012 -5510 5068 -5454
rect 3447 -6614 3503 -6612
rect 3447 -6666 3449 -6614
rect 3449 -6666 3501 -6614
rect 3501 -6666 3503 -6614
rect 3447 -6668 3503 -6666
rect 3447 -6718 3503 -6716
rect 3447 -6770 3449 -6718
rect 3449 -6770 3501 -6718
rect 3501 -6770 3503 -6718
rect 3447 -6772 3503 -6770
rect 4668 -6668 4724 -6612
rect 4772 -6668 4828 -6612
rect 4668 -6772 4724 -6716
rect 4772 -6772 4828 -6716
rect 4908 -6811 4964 -6755
rect 5012 -6811 5068 -6755
rect 4908 -6915 4964 -6859
rect 5012 -6915 5068 -6859
rect 4668 -7197 4724 -7141
rect 4772 -7197 4828 -7141
rect 4668 -7301 4724 -7245
rect 4772 -7301 4828 -7245
rect 3495 -7384 3551 -7382
rect 3495 -7436 3497 -7384
rect 3497 -7436 3549 -7384
rect 3549 -7436 3551 -7384
rect 3495 -7438 3551 -7436
rect 3495 -7488 3551 -7486
rect 3495 -7540 3497 -7488
rect 3497 -7540 3549 -7488
rect 3549 -7540 3551 -7488
rect 3495 -7542 3551 -7540
rect 5617 -5082 5673 -5026
rect 5721 -5082 5777 -5026
rect 5617 -5186 5673 -5130
rect 5721 -5186 5777 -5130
rect 6068 -5056 6124 -5054
rect 6068 -5108 6070 -5056
rect 6070 -5108 6122 -5056
rect 6122 -5108 6124 -5056
rect 6068 -5110 6124 -5108
rect 6172 -5056 6228 -5054
rect 6172 -5108 6174 -5056
rect 6174 -5108 6226 -5056
rect 6226 -5108 6228 -5056
rect 6172 -5110 6228 -5108
rect 5375 -5600 5431 -5544
rect 5479 -5600 5535 -5544
rect 5375 -5704 5431 -5648
rect 5479 -5704 5535 -5648
rect 5375 -5808 5431 -5752
rect 5479 -5808 5535 -5752
rect 5375 -5912 5431 -5856
rect 5479 -5912 5535 -5856
rect 6068 -5160 6124 -5158
rect 6068 -5212 6070 -5160
rect 6070 -5212 6122 -5160
rect 6122 -5212 6124 -5160
rect 6068 -5214 6124 -5212
rect 6172 -5160 6228 -5158
rect 6172 -5212 6174 -5160
rect 6174 -5212 6226 -5160
rect 6226 -5212 6228 -5160
rect 6172 -5214 6228 -5212
rect 6378 -5110 6434 -5054
rect 6482 -5110 6538 -5054
rect 6378 -5214 6434 -5158
rect 6482 -5214 6538 -5158
rect 5617 -6324 5673 -6268
rect 5721 -6324 5777 -6268
rect 5617 -6428 5673 -6372
rect 5721 -6428 5777 -6372
rect 6106 -6757 6162 -6755
rect 6106 -6809 6108 -6757
rect 6108 -6809 6160 -6757
rect 6160 -6809 6162 -6757
rect 6106 -6811 6162 -6809
rect 6106 -6861 6162 -6859
rect 6106 -6913 6108 -6861
rect 6108 -6913 6160 -6861
rect 6160 -6913 6162 -6861
rect 6106 -6915 6162 -6913
rect 6036 -7197 6092 -7141
rect 6140 -7197 6196 -7141
rect 6036 -7247 6092 -7245
rect 6036 -7299 6038 -7247
rect 6038 -7299 6090 -7247
rect 6090 -7299 6092 -7247
rect 6036 -7301 6092 -7299
rect 6140 -7247 6196 -7245
rect 6140 -7299 6142 -7247
rect 6142 -7299 6194 -7247
rect 6194 -7299 6196 -7247
rect 6140 -7301 6196 -7299
rect 6642 -6324 6698 -6268
rect 6746 -6324 6802 -6268
rect 6642 -6428 6698 -6372
rect 6746 -6428 6802 -6372
rect 8713 -3169 8769 -3113
rect 8713 -3219 8769 -3217
rect 8713 -3271 8715 -3219
rect 8715 -3271 8767 -3219
rect 8767 -3271 8769 -3219
rect 8713 -3273 8769 -3271
rect 9802 -3115 9858 -3113
rect 9802 -3167 9804 -3115
rect 9804 -3167 9856 -3115
rect 9856 -3167 9858 -3115
rect 9802 -3169 9858 -3167
rect 9906 -3115 9962 -3113
rect 9906 -3167 9908 -3115
rect 9908 -3167 9960 -3115
rect 9960 -3167 9962 -3115
rect 9906 -3169 9962 -3167
rect 9802 -3219 9858 -3217
rect 9802 -3271 9804 -3219
rect 9804 -3271 9856 -3219
rect 9856 -3271 9858 -3219
rect 9802 -3273 9858 -3271
rect 9906 -3219 9962 -3217
rect 9906 -3271 9908 -3219
rect 9908 -3271 9960 -3219
rect 9960 -3271 9962 -3219
rect 9906 -3273 9962 -3271
rect 7353 -3448 7409 -3446
rect 7353 -3500 7355 -3448
rect 7355 -3500 7407 -3448
rect 7407 -3500 7409 -3448
rect 7353 -3502 7409 -3500
rect 7353 -3552 7409 -3550
rect 7353 -3604 7355 -3552
rect 7355 -3604 7407 -3552
rect 7407 -3604 7409 -3552
rect 7353 -3606 7409 -3604
rect 7673 -3448 7729 -3446
rect 7673 -3500 7675 -3448
rect 7675 -3500 7727 -3448
rect 7727 -3500 7729 -3448
rect 7673 -3502 7729 -3500
rect 7673 -3552 7729 -3550
rect 7673 -3604 7675 -3552
rect 7675 -3604 7727 -3552
rect 7727 -3604 7729 -3552
rect 7673 -3606 7729 -3604
rect 7993 -3448 8049 -3446
rect 7993 -3500 7995 -3448
rect 7995 -3500 8047 -3448
rect 8047 -3500 8049 -3448
rect 7993 -3502 8049 -3500
rect 7993 -3552 8049 -3550
rect 7993 -3604 7995 -3552
rect 7995 -3604 8047 -3552
rect 8047 -3604 8049 -3552
rect 7993 -3606 8049 -3604
rect 8313 -3448 8369 -3446
rect 8313 -3500 8315 -3448
rect 8315 -3500 8367 -3448
rect 8367 -3500 8369 -3448
rect 8313 -3502 8369 -3500
rect 8313 -3552 8369 -3550
rect 8313 -3604 8315 -3552
rect 8315 -3604 8367 -3552
rect 8367 -3604 8369 -3552
rect 8313 -3606 8369 -3604
rect 8473 -3448 8529 -3446
rect 8473 -3500 8475 -3448
rect 8475 -3500 8527 -3448
rect 8527 -3500 8529 -3448
rect 8473 -3502 8529 -3500
rect 8473 -3552 8529 -3550
rect 8473 -3604 8475 -3552
rect 8475 -3604 8527 -3552
rect 8527 -3604 8529 -3552
rect 8473 -3606 8529 -3604
rect 7513 -3984 7569 -3982
rect 7513 -4036 7515 -3984
rect 7515 -4036 7567 -3984
rect 7567 -4036 7569 -3984
rect 7513 -4038 7569 -4036
rect 7513 -4088 7569 -4086
rect 7513 -4140 7515 -4088
rect 7515 -4140 7567 -4088
rect 7567 -4140 7569 -4088
rect 7513 -4142 7569 -4140
rect 7673 -3984 7729 -3982
rect 7673 -4036 7675 -3984
rect 7675 -4036 7727 -3984
rect 7727 -4036 7729 -3984
rect 7673 -4038 7729 -4036
rect 7673 -4088 7729 -4086
rect 7673 -4140 7675 -4088
rect 7675 -4140 7727 -4088
rect 7727 -4140 7729 -4088
rect 7673 -4142 7729 -4140
rect 7993 -3984 8049 -3982
rect 7993 -4036 7995 -3984
rect 7995 -4036 8047 -3984
rect 8047 -4036 8049 -3984
rect 7993 -4038 8049 -4036
rect 7993 -4088 8049 -4086
rect 7993 -4140 7995 -4088
rect 7995 -4140 8047 -4088
rect 8047 -4140 8049 -4088
rect 7993 -4142 8049 -4140
rect 8313 -3984 8369 -3982
rect 8313 -4036 8315 -3984
rect 8315 -4036 8367 -3984
rect 8367 -4036 8369 -3984
rect 8313 -4038 8369 -4036
rect 8313 -4088 8369 -4086
rect 8313 -4140 8315 -4088
rect 8315 -4140 8367 -4088
rect 8367 -4140 8369 -4088
rect 8313 -4142 8369 -4140
rect 7353 -4520 7409 -4518
rect 7353 -4572 7355 -4520
rect 7355 -4572 7407 -4520
rect 7407 -4572 7409 -4520
rect 7353 -4574 7409 -4572
rect 7353 -4624 7409 -4622
rect 7353 -4676 7355 -4624
rect 7355 -4676 7407 -4624
rect 7407 -4676 7409 -4624
rect 7353 -4678 7409 -4676
rect 8792 -3755 8848 -3753
rect 8792 -3807 8794 -3755
rect 8794 -3807 8846 -3755
rect 8846 -3807 8848 -3755
rect 8792 -3809 8848 -3807
rect 8633 -3984 8689 -3982
rect 8633 -4036 8635 -3984
rect 8635 -4036 8687 -3984
rect 8687 -4036 8689 -3984
rect 8633 -4038 8689 -4036
rect 8633 -4088 8689 -4086
rect 8633 -4140 8635 -4088
rect 8635 -4140 8687 -4088
rect 8687 -4140 8689 -4088
rect 8633 -4142 8689 -4140
rect 10068 -3713 10124 -3711
rect 10068 -3765 10070 -3713
rect 10070 -3765 10122 -3713
rect 10122 -3765 10124 -3713
rect 10068 -3767 10124 -3765
rect 10172 -3713 10228 -3711
rect 10172 -3765 10174 -3713
rect 10174 -3765 10226 -3713
rect 10226 -3765 10228 -3713
rect 10172 -3767 10228 -3765
rect 10068 -3817 10124 -3815
rect 10068 -3869 10070 -3817
rect 10070 -3869 10122 -3817
rect 10122 -3869 10124 -3817
rect 10068 -3871 10124 -3869
rect 10172 -3817 10228 -3815
rect 10172 -3869 10174 -3817
rect 10174 -3869 10226 -3817
rect 10226 -3869 10228 -3817
rect 10172 -3871 10228 -3869
rect 8595 -4291 8651 -4289
rect 8595 -4343 8597 -4291
rect 8597 -4343 8649 -4291
rect 8649 -4343 8651 -4291
rect 8595 -4345 8651 -4343
rect 9802 -4293 9858 -4237
rect 9906 -4293 9962 -4237
rect 9802 -4397 9858 -4341
rect 9906 -4397 9962 -4341
rect 7673 -4520 7729 -4518
rect 7673 -4572 7675 -4520
rect 7675 -4572 7727 -4520
rect 7727 -4572 7729 -4520
rect 7673 -4574 7729 -4572
rect 7673 -4624 7729 -4622
rect 7673 -4676 7675 -4624
rect 7675 -4676 7727 -4624
rect 7727 -4676 7729 -4624
rect 7673 -4678 7729 -4676
rect 7993 -4520 8049 -4518
rect 7993 -4572 7995 -4520
rect 7995 -4572 8047 -4520
rect 8047 -4572 8049 -4520
rect 7993 -4574 8049 -4572
rect 7993 -4624 8049 -4622
rect 7993 -4676 7995 -4624
rect 7995 -4676 8047 -4624
rect 8047 -4676 8049 -4624
rect 7993 -4678 8049 -4676
rect 8313 -4520 8369 -4518
rect 8313 -4572 8315 -4520
rect 8315 -4572 8367 -4520
rect 8367 -4572 8369 -4520
rect 8313 -4574 8369 -4572
rect 8313 -4624 8369 -4622
rect 8313 -4676 8315 -4624
rect 8315 -4676 8367 -4624
rect 8367 -4676 8369 -4624
rect 8313 -4678 8369 -4676
rect 8633 -4520 8689 -4518
rect 8633 -4572 8635 -4520
rect 8635 -4572 8687 -4520
rect 8687 -4572 8689 -4520
rect 8633 -4574 8689 -4572
rect 8633 -4624 8689 -4622
rect 8633 -4676 8635 -4624
rect 8635 -4676 8687 -4624
rect 8687 -4676 8689 -4624
rect 8633 -4678 8689 -4676
rect 7353 -5056 7409 -5054
rect 7353 -5108 7355 -5056
rect 7355 -5108 7407 -5056
rect 7407 -5108 7409 -5056
rect 7353 -5110 7409 -5108
rect 7353 -5160 7409 -5158
rect 7353 -5212 7355 -5160
rect 7355 -5212 7407 -5160
rect 7407 -5212 7409 -5160
rect 7353 -5214 7409 -5212
rect 7673 -5056 7729 -5054
rect 7673 -5108 7675 -5056
rect 7675 -5108 7727 -5056
rect 7727 -5108 7729 -5056
rect 7673 -5110 7729 -5108
rect 7673 -5160 7729 -5158
rect 7673 -5212 7675 -5160
rect 7675 -5212 7727 -5160
rect 7727 -5212 7729 -5160
rect 7673 -5214 7729 -5212
rect 7993 -5056 8049 -5054
rect 7993 -5108 7995 -5056
rect 7995 -5108 8047 -5056
rect 8047 -5108 8049 -5056
rect 7993 -5110 8049 -5108
rect 7993 -5160 8049 -5158
rect 7993 -5212 7995 -5160
rect 7995 -5212 8047 -5160
rect 8047 -5212 8049 -5160
rect 7993 -5214 8049 -5212
rect 8313 -5056 8369 -5054
rect 8313 -5108 8315 -5056
rect 8315 -5108 8367 -5056
rect 8367 -5108 8369 -5056
rect 8313 -5110 8369 -5108
rect 8313 -5160 8369 -5158
rect 8313 -5212 8315 -5160
rect 8315 -5212 8367 -5160
rect 8367 -5212 8369 -5160
rect 8313 -5214 8369 -5212
rect 8713 -4825 8769 -4823
rect 8713 -4877 8715 -4825
rect 8715 -4877 8767 -4825
rect 8767 -4877 8769 -4825
rect 8713 -4879 8769 -4877
rect 8633 -5056 8689 -5054
rect 8633 -5108 8635 -5056
rect 8635 -5108 8687 -5056
rect 8687 -5108 8689 -5056
rect 8633 -5110 8689 -5108
rect 8633 -5160 8689 -5158
rect 8633 -5212 8635 -5160
rect 8635 -5212 8687 -5160
rect 8687 -5212 8689 -5160
rect 8633 -5214 8689 -5212
rect 8792 -5311 8848 -5255
rect 8792 -5361 8848 -5359
rect 8792 -5413 8794 -5361
rect 8794 -5413 8846 -5361
rect 8846 -5413 8848 -5361
rect 8792 -5415 8848 -5413
rect 10068 -4827 10124 -4771
rect 10172 -4827 10228 -4771
rect 10068 -4931 10124 -4875
rect 10172 -4931 10228 -4875
rect 9530 -5311 9586 -5255
rect 9634 -5311 9690 -5255
rect 9530 -5415 9586 -5359
rect 9634 -5415 9690 -5359
rect 9802 -5313 9858 -5257
rect 9906 -5313 9962 -5257
rect 9802 -5417 9858 -5361
rect 9906 -5417 9962 -5361
rect 8473 -5592 8529 -5590
rect 8473 -5644 8475 -5592
rect 8475 -5644 8527 -5592
rect 8527 -5644 8529 -5592
rect 8473 -5646 8529 -5644
rect 8473 -5696 8529 -5694
rect 8473 -5748 8475 -5696
rect 8475 -5748 8527 -5696
rect 8527 -5748 8529 -5696
rect 8473 -5750 8529 -5748
rect 8792 -5826 8848 -5770
rect 8792 -5876 8848 -5874
rect 8792 -5928 8794 -5876
rect 8794 -5928 8846 -5876
rect 8846 -5928 8848 -5876
rect 8792 -5930 8848 -5928
rect 9263 -6052 9319 -5996
rect 9367 -6052 9423 -5996
rect 9263 -6156 9319 -6100
rect 9367 -6156 9423 -6100
rect 8393 -6448 8449 -6446
rect 8393 -6500 8395 -6448
rect 8395 -6500 8447 -6448
rect 8447 -6500 8449 -6448
rect 8393 -6502 8449 -6500
rect 8393 -6606 8449 -6550
rect 10068 -5826 10124 -5770
rect 10172 -5826 10228 -5770
rect 10068 -5930 10124 -5874
rect 10172 -5930 10228 -5874
rect 9530 -6502 9586 -6446
rect 9634 -6502 9690 -6446
rect 9530 -6606 9586 -6550
rect 9634 -6606 9690 -6550
rect 6642 -7207 6698 -7151
rect 6746 -7207 6802 -7151
rect 6642 -7311 6698 -7255
rect 6746 -7311 6802 -7255
rect 8920 -7153 8976 -7151
rect 8920 -7205 8922 -7153
rect 8922 -7205 8974 -7153
rect 8974 -7205 8976 -7153
rect 8920 -7207 8976 -7205
rect 9024 -7153 9080 -7151
rect 9024 -7205 9026 -7153
rect 9026 -7205 9078 -7153
rect 9078 -7205 9080 -7153
rect 9024 -7207 9080 -7205
rect 8920 -7257 8976 -7255
rect 8920 -7309 8922 -7257
rect 8922 -7309 8974 -7257
rect 8974 -7309 8976 -7257
rect 8920 -7311 8976 -7309
rect 9024 -7257 9080 -7255
rect 9024 -7309 9026 -7257
rect 9026 -7309 9078 -7257
rect 9078 -7309 9080 -7257
rect 9024 -7311 9080 -7309
rect 5946 -7386 6002 -7384
rect 5946 -7438 5948 -7386
rect 5948 -7438 6000 -7386
rect 6000 -7438 6002 -7386
rect 5946 -7440 6002 -7438
rect 5946 -7490 6002 -7488
rect 5946 -7542 5948 -7490
rect 5948 -7542 6000 -7490
rect 6000 -7542 6002 -7490
rect 5946 -7544 6002 -7542
rect 6378 -7392 6434 -7390
rect 6378 -7444 6380 -7392
rect 6380 -7444 6432 -7392
rect 6432 -7444 6434 -7392
rect 6378 -7446 6434 -7444
rect 6482 -7446 6538 -7390
rect 6378 -7496 6434 -7494
rect 6378 -7548 6380 -7496
rect 6380 -7548 6432 -7496
rect 6432 -7548 6434 -7496
rect 6378 -7550 6434 -7548
rect 6482 -7550 6538 -7494
rect 5894 -8084 5950 -8028
rect 5998 -8084 6054 -8028
rect 5894 -8188 5950 -8132
rect 5998 -8188 6054 -8132
rect 13508 1032 13564 1034
rect 13508 980 13510 1032
rect 13510 980 13562 1032
rect 13562 980 13564 1032
rect 13508 978 13564 980
rect 14670 1136 14726 1138
rect 14670 1084 14672 1136
rect 14672 1084 14724 1136
rect 14724 1084 14726 1136
rect 14670 1082 14726 1084
rect 14670 1032 14726 1034
rect 14670 980 14672 1032
rect 14672 980 14724 1032
rect 14724 980 14726 1032
rect 14670 978 14726 980
rect 15310 1136 15366 1138
rect 15310 1084 15312 1136
rect 15312 1084 15364 1136
rect 15364 1084 15366 1136
rect 15310 1082 15366 1084
rect 15310 1032 15366 1034
rect 15310 980 15312 1032
rect 15312 980 15364 1032
rect 15364 980 15366 1032
rect 15310 978 15366 980
rect 15950 1136 16006 1138
rect 15950 1084 15952 1136
rect 15952 1084 16004 1136
rect 16004 1084 16006 1136
rect 15950 1082 16006 1084
rect 15950 1032 16006 1034
rect 15950 980 15952 1032
rect 15952 980 16004 1032
rect 16004 980 16006 1032
rect 15950 978 16006 980
rect 16627 1082 16683 1138
rect 16731 1082 16787 1138
rect 16627 978 16683 1034
rect 16731 978 16787 1034
rect 11876 116 11932 118
rect 11876 64 11878 116
rect 11878 64 11930 116
rect 11930 64 11932 116
rect 11876 62 11932 64
rect 11876 12 11932 14
rect 11876 -40 11878 12
rect 11878 -40 11930 12
rect 11930 -40 11932 12
rect 11876 -42 11932 -40
rect 12772 116 12828 118
rect 12772 64 12774 116
rect 12774 64 12826 116
rect 12826 64 12828 116
rect 12772 62 12828 64
rect 12772 12 12828 14
rect 12772 -40 12774 12
rect 12774 -40 12826 12
rect 12826 -40 12828 12
rect 12772 -42 12828 -40
rect 13668 116 13724 118
rect 13668 64 13670 116
rect 13670 64 13722 116
rect 13722 64 13724 116
rect 13668 62 13724 64
rect 13668 12 13724 14
rect 13668 -40 13670 12
rect 13670 -40 13722 12
rect 13722 -40 13724 12
rect 13668 -42 13724 -40
rect 13380 -284 13436 -282
rect 13380 -336 13382 -284
rect 13382 -336 13434 -284
rect 13434 -336 13436 -284
rect 13380 -338 13436 -336
rect 13380 -388 13436 -386
rect 13380 -440 13382 -388
rect 13382 -440 13434 -388
rect 13434 -440 13436 -388
rect 13380 -442 13436 -440
rect 14990 -284 15046 -282
rect 14990 -336 14992 -284
rect 14992 -336 15044 -284
rect 15044 -336 15046 -284
rect 14990 -338 15046 -336
rect 14990 -388 15046 -386
rect 14990 -440 14992 -388
rect 14992 -440 15044 -388
rect 15044 -440 15046 -388
rect 14990 -442 15046 -440
rect 15630 -284 15686 -282
rect 15630 -336 15632 -284
rect 15632 -336 15684 -284
rect 15684 -336 15686 -284
rect 15630 -338 15686 -336
rect 15630 -388 15686 -386
rect 15630 -440 15632 -388
rect 15632 -440 15684 -388
rect 15684 -440 15686 -388
rect 15630 -442 15686 -440
rect 11163 -508 11219 -452
rect 11267 -508 11323 -452
rect 11163 -612 11219 -556
rect 11267 -612 11323 -556
rect 10895 -988 10951 -932
rect 10999 -988 11055 -932
rect 10895 -1092 10951 -1036
rect 10999 -1092 11055 -1036
rect 11542 -648 11598 -592
rect 11646 -648 11702 -592
rect 11542 -752 11598 -696
rect 11646 -752 11702 -696
rect 11912 -594 11968 -592
rect 11912 -646 11914 -594
rect 11914 -646 11966 -594
rect 11966 -646 11968 -594
rect 11912 -648 11968 -646
rect 11912 -698 11968 -696
rect 11912 -750 11914 -698
rect 11914 -750 11966 -698
rect 11966 -750 11968 -698
rect 11912 -752 11968 -750
rect 14210 -643 14266 -587
rect 14314 -643 14370 -587
rect 14210 -747 14266 -691
rect 14314 -747 14370 -691
rect 14698 -589 14754 -587
rect 14698 -641 14700 -589
rect 14700 -641 14752 -589
rect 14752 -641 14754 -589
rect 14698 -643 14754 -641
rect 14698 -693 14754 -691
rect 14698 -745 14700 -693
rect 14700 -745 14752 -693
rect 14752 -745 14754 -693
rect 14698 -747 14754 -745
rect 11163 -1388 11219 -1332
rect 11267 -1388 11323 -1332
rect 11163 -1492 11219 -1436
rect 11267 -1492 11323 -1436
rect 10442 -7207 10498 -7151
rect 10546 -7207 10602 -7151
rect 10442 -7311 10498 -7255
rect 10546 -7311 10602 -7255
rect 10829 -7153 10885 -7151
rect 10829 -7205 10831 -7153
rect 10831 -7205 10883 -7153
rect 10883 -7205 10885 -7153
rect 10829 -7207 10885 -7205
rect 10933 -7153 10989 -7151
rect 10933 -7205 10935 -7153
rect 10935 -7205 10987 -7153
rect 10987 -7205 10989 -7153
rect 10933 -7207 10989 -7205
rect 10829 -7257 10885 -7255
rect 10829 -7309 10831 -7257
rect 10831 -7309 10883 -7257
rect 10883 -7309 10885 -7257
rect 10829 -7311 10885 -7309
rect 10933 -7257 10989 -7255
rect 10933 -7309 10935 -7257
rect 10935 -7309 10987 -7257
rect 10987 -7309 10989 -7257
rect 10933 -7311 10989 -7309
rect 12324 -934 12380 -932
rect 12324 -986 12326 -934
rect 12326 -986 12378 -934
rect 12378 -986 12380 -934
rect 12324 -988 12380 -986
rect 12324 -1038 12380 -1036
rect 12324 -1090 12326 -1038
rect 12326 -1090 12378 -1038
rect 12378 -1090 12380 -1038
rect 12324 -1092 12380 -1090
rect 13220 -934 13276 -932
rect 13220 -986 13222 -934
rect 13222 -986 13274 -934
rect 13274 -986 13276 -934
rect 13220 -988 13276 -986
rect 13220 -1038 13276 -1036
rect 13220 -1090 13222 -1038
rect 13222 -1090 13274 -1038
rect 13274 -1090 13276 -1038
rect 13220 -1092 13276 -1090
rect 13380 -934 13436 -932
rect 13380 -986 13382 -934
rect 13382 -986 13434 -934
rect 13434 -986 13436 -934
rect 13380 -988 13436 -986
rect 13380 -1038 13436 -1036
rect 13380 -1090 13382 -1038
rect 13382 -1090 13434 -1038
rect 13434 -1090 13436 -1038
rect 13380 -1092 13436 -1090
rect 11876 -1334 11932 -1332
rect 11876 -1386 11878 -1334
rect 11878 -1386 11930 -1334
rect 11930 -1386 11932 -1334
rect 11876 -1388 11932 -1386
rect 11876 -1438 11932 -1436
rect 11876 -1490 11878 -1438
rect 11878 -1490 11930 -1438
rect 11930 -1490 11932 -1438
rect 11876 -1492 11932 -1490
rect 12772 -1334 12828 -1332
rect 12772 -1386 12774 -1334
rect 12774 -1386 12826 -1334
rect 12826 -1386 12828 -1334
rect 12772 -1388 12828 -1386
rect 12772 -1438 12828 -1436
rect 12772 -1490 12774 -1438
rect 12774 -1490 12826 -1438
rect 12826 -1490 12828 -1438
rect 12772 -1492 12828 -1490
rect 13668 -1334 13724 -1332
rect 13668 -1386 13670 -1334
rect 13670 -1386 13722 -1334
rect 13722 -1386 13724 -1334
rect 13668 -1388 13724 -1386
rect 13668 -1438 13724 -1436
rect 13668 -1490 13670 -1438
rect 13670 -1490 13722 -1438
rect 13722 -1490 13724 -1438
rect 13668 -1492 13724 -1490
rect 16889 -338 16945 -282
rect 16993 -338 17049 -282
rect 16889 -442 16945 -386
rect 16993 -442 17049 -386
rect 14990 -934 15046 -932
rect 14990 -986 14992 -934
rect 14992 -986 15044 -934
rect 15044 -986 15046 -934
rect 14990 -988 15046 -986
rect 14990 -1038 15046 -1036
rect 14990 -1090 14992 -1038
rect 14992 -1090 15044 -1038
rect 15044 -1090 15046 -1038
rect 14990 -1092 15046 -1090
rect 15630 -934 15686 -932
rect 15630 -986 15632 -934
rect 15632 -986 15684 -934
rect 15684 -986 15686 -934
rect 15630 -988 15686 -986
rect 15630 -1038 15686 -1036
rect 15630 -1090 15632 -1038
rect 15632 -1090 15684 -1038
rect 15684 -1090 15686 -1038
rect 15630 -1092 15686 -1090
rect 16627 -988 16683 -932
rect 16731 -988 16787 -932
rect 16627 -1092 16683 -1036
rect 16731 -1092 16787 -1036
rect 17165 -516 17221 -460
rect 17365 3228 17421 3284
rect 18589 3282 18645 3284
rect 18589 3230 18591 3282
rect 18591 3230 18643 3282
rect 18643 3230 18645 3282
rect 18589 3228 18645 3230
rect 18829 3071 18885 3073
rect 18829 3019 18831 3071
rect 18831 3019 18883 3071
rect 18883 3019 18885 3071
rect 18829 3017 18885 3019
rect 18829 2967 18885 2969
rect 18829 2915 18831 2967
rect 18831 2915 18883 2967
rect 18883 2915 18885 2967
rect 18829 2913 18885 2915
rect 19469 3071 19525 3073
rect 19469 3019 19471 3071
rect 19471 3019 19523 3071
rect 19523 3019 19525 3071
rect 19469 3017 19525 3019
rect 19469 2967 19525 2969
rect 19469 2915 19471 2967
rect 19471 2915 19523 2967
rect 19523 2915 19525 2967
rect 19469 2913 19525 2915
rect 20972 3121 21028 3177
rect 21076 3121 21132 3177
rect 21180 3121 21236 3177
rect 20972 3017 21028 3073
rect 21076 3017 21132 3073
rect 21180 3017 21236 3073
rect 20972 2913 21028 2969
rect 21076 2913 21132 2969
rect 21180 2913 21236 2969
rect 18509 2677 18565 2679
rect 18509 2625 18511 2677
rect 18511 2625 18563 2677
rect 18563 2625 18565 2677
rect 18509 2623 18565 2625
rect 18509 2573 18565 2575
rect 18509 2521 18511 2573
rect 18511 2521 18563 2573
rect 18563 2521 18565 2573
rect 18509 2519 18565 2521
rect 19149 2677 19205 2679
rect 19149 2625 19151 2677
rect 19151 2625 19203 2677
rect 19203 2625 19205 2677
rect 19149 2623 19205 2625
rect 19149 2573 19205 2575
rect 19149 2521 19151 2573
rect 19151 2521 19203 2573
rect 19203 2521 19205 2573
rect 19149 2519 19205 2521
rect 19789 2677 19845 2679
rect 19789 2625 19791 2677
rect 19791 2625 19843 2677
rect 19843 2625 19845 2677
rect 19789 2623 19845 2625
rect 19789 2573 19845 2575
rect 19789 2521 19791 2573
rect 19791 2521 19843 2573
rect 19843 2521 19845 2573
rect 19789 2519 19845 2521
rect 18589 2346 18645 2348
rect 18589 2294 18591 2346
rect 18591 2294 18643 2346
rect 18643 2294 18645 2346
rect 18589 2292 18645 2294
rect 18829 2135 18885 2137
rect 18829 2083 18831 2135
rect 18831 2083 18883 2135
rect 18883 2083 18885 2135
rect 18829 2081 18885 2083
rect 18829 2031 18885 2033
rect 18829 1979 18831 2031
rect 18831 1979 18883 2031
rect 18883 1979 18885 2031
rect 18829 1977 18885 1979
rect 19469 2135 19525 2137
rect 19469 2083 19471 2135
rect 19471 2083 19523 2135
rect 19523 2083 19525 2135
rect 19469 2081 19525 2083
rect 19469 2031 19525 2033
rect 19469 1979 19471 2031
rect 19471 1979 19523 2031
rect 19523 1979 19525 2031
rect 19469 1977 19525 1979
rect 20972 1791 21028 1847
rect 21076 1791 21132 1847
rect 21180 1791 21236 1847
rect 18509 1741 18565 1743
rect 18509 1689 18511 1741
rect 18511 1689 18563 1741
rect 18563 1689 18565 1741
rect 18509 1687 18565 1689
rect 18509 1637 18565 1639
rect 18509 1585 18511 1637
rect 18511 1585 18563 1637
rect 18563 1585 18565 1637
rect 18509 1583 18565 1585
rect 19149 1741 19205 1743
rect 19149 1689 19151 1741
rect 19151 1689 19203 1741
rect 19203 1689 19205 1741
rect 19149 1687 19205 1689
rect 19149 1637 19205 1639
rect 19149 1585 19151 1637
rect 19151 1585 19203 1637
rect 19203 1585 19205 1637
rect 19149 1583 19205 1585
rect 19789 1741 19845 1743
rect 19789 1689 19791 1741
rect 19791 1689 19843 1741
rect 19843 1689 19845 1741
rect 19789 1687 19845 1689
rect 19789 1637 19845 1639
rect 19789 1585 19791 1637
rect 19791 1585 19843 1637
rect 19843 1585 19845 1637
rect 19789 1583 19845 1585
rect 20972 1687 21028 1743
rect 21076 1687 21132 1743
rect 21180 1687 21236 1743
rect 20972 1583 21028 1639
rect 21076 1583 21132 1639
rect 21180 1583 21236 1639
rect 18829 1199 18885 1201
rect 18829 1147 18831 1199
rect 18831 1147 18883 1199
rect 18883 1147 18885 1199
rect 18829 1145 18885 1147
rect 18829 1095 18885 1097
rect 18829 1043 18831 1095
rect 18831 1043 18883 1095
rect 18883 1043 18885 1095
rect 18829 1041 18885 1043
rect 18509 805 18565 807
rect 18509 753 18511 805
rect 18511 753 18563 805
rect 18563 753 18565 805
rect 18509 751 18565 753
rect 18509 701 18565 703
rect 18509 649 18511 701
rect 18511 649 18563 701
rect 18563 649 18565 701
rect 18509 647 18565 649
rect 17365 420 17421 476
rect 14670 -1324 14726 -1322
rect 14670 -1376 14672 -1324
rect 14672 -1376 14724 -1324
rect 14724 -1376 14726 -1324
rect 14670 -1378 14726 -1376
rect 14670 -1428 14726 -1426
rect 14670 -1480 14672 -1428
rect 14672 -1480 14724 -1428
rect 14724 -1480 14726 -1428
rect 14670 -1482 14726 -1480
rect 15310 -1324 15366 -1322
rect 15310 -1376 15312 -1324
rect 15312 -1376 15364 -1324
rect 15364 -1376 15366 -1324
rect 15310 -1378 15366 -1376
rect 15310 -1428 15366 -1426
rect 15310 -1480 15312 -1428
rect 15312 -1480 15364 -1428
rect 15364 -1480 15366 -1428
rect 15310 -1482 15366 -1480
rect 15950 -1324 16006 -1322
rect 15950 -1376 15952 -1324
rect 15952 -1376 16004 -1324
rect 16004 -1376 16006 -1324
rect 15950 -1378 16006 -1376
rect 15950 -1428 16006 -1426
rect 15950 -1480 15952 -1428
rect 15952 -1480 16004 -1428
rect 16004 -1480 16006 -1428
rect 15950 -1482 16006 -1480
rect 16889 -1378 16945 -1322
rect 16993 -1378 17049 -1322
rect 16889 -1482 16945 -1426
rect 16993 -1482 17049 -1426
rect 18589 474 18645 476
rect 18589 422 18591 474
rect 18591 422 18643 474
rect 18643 422 18645 474
rect 18589 420 18645 422
rect 18829 263 18885 265
rect 18829 211 18831 263
rect 18831 211 18883 263
rect 18883 211 18885 263
rect 18829 209 18885 211
rect 18829 159 18885 161
rect 18829 107 18831 159
rect 18831 107 18883 159
rect 18883 107 18885 159
rect 18829 105 18885 107
rect 19149 805 19205 807
rect 19149 753 19151 805
rect 19151 753 19203 805
rect 19203 753 19205 805
rect 19149 751 19205 753
rect 19149 701 19205 703
rect 19149 649 19151 701
rect 19151 649 19203 701
rect 19203 649 19205 701
rect 19149 647 19205 649
rect 19469 1199 19525 1201
rect 19469 1147 19471 1199
rect 19471 1147 19523 1199
rect 19523 1147 19525 1199
rect 19469 1145 19525 1147
rect 19469 1095 19525 1097
rect 19469 1043 19471 1095
rect 19471 1043 19523 1095
rect 19523 1043 19525 1095
rect 19469 1041 19525 1043
rect 19469 263 19525 265
rect 19469 211 19471 263
rect 19471 211 19523 263
rect 19523 211 19525 263
rect 19469 209 19525 211
rect 19469 159 19525 161
rect 19469 107 19471 159
rect 19471 107 19523 159
rect 19523 107 19525 159
rect 19469 105 19525 107
rect 20972 855 21028 911
rect 21076 855 21132 911
rect 21180 855 21236 911
rect 19789 805 19845 807
rect 19789 753 19791 805
rect 19791 753 19843 805
rect 19843 753 19845 805
rect 19789 751 19845 753
rect 19789 701 19845 703
rect 19789 649 19791 701
rect 19791 649 19843 701
rect 19843 649 19845 701
rect 19789 647 19845 649
rect 20972 751 21028 807
rect 21076 751 21132 807
rect 21180 751 21236 807
rect 20972 647 21028 703
rect 21076 647 21132 703
rect 21180 647 21236 703
rect 20972 313 21028 369
rect 21076 313 21132 369
rect 21180 313 21236 369
rect 20972 209 21028 265
rect 21076 209 21132 265
rect 21180 209 21236 265
rect 20972 105 21028 161
rect 21076 105 21132 161
rect 21180 105 21236 161
rect 18509 -131 18565 -129
rect 18509 -183 18511 -131
rect 18511 -183 18563 -131
rect 18563 -183 18565 -131
rect 18509 -185 18565 -183
rect 18509 -235 18565 -233
rect 18509 -287 18511 -235
rect 18511 -287 18563 -235
rect 18563 -287 18565 -235
rect 18509 -289 18565 -287
rect 19149 -131 19205 -129
rect 19149 -183 19151 -131
rect 19151 -183 19203 -131
rect 19203 -183 19205 -131
rect 19149 -185 19205 -183
rect 19149 -235 19205 -233
rect 19149 -287 19151 -235
rect 19151 -287 19203 -235
rect 19203 -287 19205 -235
rect 19149 -289 19205 -287
rect 19789 -131 19845 -129
rect 19789 -183 19791 -131
rect 19791 -183 19843 -131
rect 19843 -183 19845 -131
rect 19789 -185 19845 -183
rect 19789 -235 19845 -233
rect 19789 -287 19791 -235
rect 19791 -287 19843 -235
rect 19843 -287 19845 -235
rect 19789 -289 19845 -287
rect 18589 -462 18645 -460
rect 18589 -514 18591 -462
rect 18591 -514 18643 -462
rect 18643 -514 18645 -462
rect 18589 -516 18645 -514
rect 18829 -673 18885 -671
rect 18829 -725 18831 -673
rect 18831 -725 18883 -673
rect 18883 -725 18885 -673
rect 18829 -727 18885 -725
rect 18829 -777 18885 -775
rect 18829 -829 18831 -777
rect 18831 -829 18883 -777
rect 18883 -829 18885 -777
rect 18829 -831 18885 -829
rect 19469 -673 19525 -671
rect 19469 -725 19471 -673
rect 19471 -725 19523 -673
rect 19523 -725 19525 -673
rect 19469 -727 19525 -725
rect 19469 -777 19525 -775
rect 19469 -829 19471 -777
rect 19471 -829 19523 -777
rect 19523 -829 19525 -777
rect 19469 -831 19525 -829
rect 23981 4007 24037 4009
rect 23981 3955 23983 4007
rect 23983 3955 24035 4007
rect 24035 3955 24037 4007
rect 23981 3953 24037 3955
rect 23981 3903 24037 3905
rect 23981 3851 23983 3903
rect 23983 3851 24035 3903
rect 24035 3851 24037 3903
rect 23981 3849 24037 3851
rect 24621 4007 24677 4009
rect 24621 3955 24623 4007
rect 24623 3955 24675 4007
rect 24675 3955 24677 4007
rect 24621 3953 24677 3955
rect 24621 3903 24677 3905
rect 24621 3851 24623 3903
rect 24623 3851 24675 3903
rect 24675 3851 24677 3903
rect 24621 3849 24677 3851
rect 21621 2727 21677 2783
rect 21725 2727 21781 2783
rect 21829 2727 21885 2783
rect 21621 2623 21677 2679
rect 21725 2623 21781 2679
rect 21829 2623 21885 2679
rect 21621 2519 21677 2575
rect 21725 2519 21781 2575
rect 21829 2519 21885 2575
rect 21621 2185 21677 2241
rect 21725 2185 21781 2241
rect 21829 2185 21885 2241
rect 21621 2081 21677 2137
rect 21725 2081 21781 2137
rect 21829 2081 21885 2137
rect 21621 1977 21677 2033
rect 21725 1977 21781 2033
rect 21829 1977 21885 2033
rect 21621 1249 21677 1305
rect 21725 1249 21781 1305
rect 21829 1249 21885 1305
rect 21621 1145 21677 1201
rect 21725 1145 21781 1201
rect 21829 1145 21885 1201
rect 21621 1041 21677 1097
rect 21725 1041 21781 1097
rect 21829 1041 21885 1097
rect 21621 -81 21677 -25
rect 21725 -81 21781 -25
rect 21829 -81 21885 -25
rect 21621 -185 21677 -129
rect 21725 -185 21781 -129
rect 21829 -185 21885 -129
rect 21621 -289 21677 -233
rect 21725 -289 21781 -233
rect 21829 -289 21885 -233
rect 21621 -623 21677 -567
rect 21725 -623 21781 -567
rect 21829 -623 21885 -567
rect 21621 -727 21677 -671
rect 21725 -727 21781 -671
rect 21829 -727 21885 -671
rect 21621 -831 21677 -775
rect 21725 -831 21781 -775
rect 21829 -831 21885 -775
rect 22270 3663 22326 3719
rect 22374 3663 22430 3719
rect 22478 3663 22534 3719
rect 22270 3559 22326 3615
rect 22374 3559 22430 3615
rect 22478 3559 22534 3615
rect 22270 3455 22326 3511
rect 22374 3455 22430 3511
rect 22478 3455 22534 3511
rect 23661 3613 23717 3615
rect 23661 3561 23663 3613
rect 23663 3561 23715 3613
rect 23715 3561 23717 3613
rect 23661 3559 23717 3561
rect 23661 3509 23717 3511
rect 23661 3457 23663 3509
rect 23663 3457 23715 3509
rect 23715 3457 23717 3509
rect 23661 3455 23717 3457
rect 24301 3613 24357 3615
rect 24301 3561 24303 3613
rect 24303 3561 24355 3613
rect 24355 3561 24357 3613
rect 24301 3559 24357 3561
rect 24301 3509 24357 3511
rect 24301 3457 24303 3509
rect 24303 3457 24355 3509
rect 24355 3457 24357 3509
rect 24301 3455 24357 3457
rect 24941 3613 24997 3615
rect 24941 3561 24943 3613
rect 24943 3561 24995 3613
rect 24995 3561 24997 3613
rect 24941 3559 24997 3561
rect 24941 3509 24997 3511
rect 24941 3457 24943 3509
rect 24943 3457 24995 3509
rect 24995 3457 24997 3509
rect 24941 3455 24997 3457
rect 22270 3121 22326 3177
rect 22374 3121 22430 3177
rect 22478 3121 22534 3177
rect 22270 3017 22326 3073
rect 22374 3017 22430 3073
rect 22478 3017 22534 3073
rect 22270 2913 22326 2969
rect 22374 2913 22430 2969
rect 22478 2913 22534 2969
rect 23981 3071 24037 3073
rect 23981 3019 23983 3071
rect 23983 3019 24035 3071
rect 24035 3019 24037 3071
rect 23981 3017 24037 3019
rect 23981 2967 24037 2969
rect 23981 2915 23983 2967
rect 23983 2915 24035 2967
rect 24035 2915 24037 2967
rect 23981 2913 24037 2915
rect 24861 3282 24917 3284
rect 24861 3230 24863 3282
rect 24863 3230 24915 3282
rect 24915 3230 24917 3282
rect 24861 3228 24917 3230
rect 26085 3228 26141 3284
rect 24621 3071 24677 3073
rect 24621 3019 24623 3071
rect 24623 3019 24675 3071
rect 24675 3019 24677 3071
rect 24621 3017 24677 3019
rect 24621 2967 24677 2969
rect 24621 2915 24623 2967
rect 24623 2915 24675 2967
rect 24675 2915 24677 2967
rect 24621 2913 24677 2915
rect 23661 2677 23717 2679
rect 23661 2625 23663 2677
rect 23663 2625 23715 2677
rect 23715 2625 23717 2677
rect 23661 2623 23717 2625
rect 23661 2573 23717 2575
rect 23661 2521 23663 2573
rect 23663 2521 23715 2573
rect 23715 2521 23717 2573
rect 23661 2519 23717 2521
rect 24301 2677 24357 2679
rect 24301 2625 24303 2677
rect 24303 2625 24355 2677
rect 24355 2625 24357 2677
rect 24301 2623 24357 2625
rect 24301 2573 24357 2575
rect 24301 2521 24303 2573
rect 24303 2521 24355 2573
rect 24355 2521 24357 2573
rect 24301 2519 24357 2521
rect 24941 2677 24997 2679
rect 24941 2625 24943 2677
rect 24943 2625 24995 2677
rect 24995 2625 24997 2677
rect 24941 2623 24997 2625
rect 24941 2573 24997 2575
rect 24941 2521 24943 2573
rect 24943 2521 24995 2573
rect 24995 2521 24997 2573
rect 24941 2519 24997 2521
rect 22270 1791 22326 1847
rect 22374 1791 22430 1847
rect 22478 1791 22534 1847
rect 23981 2135 24037 2137
rect 23981 2083 23983 2135
rect 23983 2083 24035 2135
rect 24035 2083 24037 2135
rect 23981 2081 24037 2083
rect 23981 2031 24037 2033
rect 23981 1979 23983 2031
rect 23983 1979 24035 2031
rect 24035 1979 24037 2031
rect 23981 1977 24037 1979
rect 24861 2346 24917 2348
rect 24861 2294 24863 2346
rect 24863 2294 24915 2346
rect 24915 2294 24917 2346
rect 24861 2292 24917 2294
rect 24621 2135 24677 2137
rect 24621 2083 24623 2135
rect 24623 2083 24675 2135
rect 24675 2083 24677 2135
rect 24621 2081 24677 2083
rect 24621 2031 24677 2033
rect 24621 1979 24623 2031
rect 24623 1979 24675 2031
rect 24675 1979 24677 2031
rect 24621 1977 24677 1979
rect 22270 1687 22326 1743
rect 22374 1687 22430 1743
rect 22478 1687 22534 1743
rect 22270 1583 22326 1639
rect 22374 1583 22430 1639
rect 22478 1583 22534 1639
rect 23661 1741 23717 1743
rect 23661 1689 23663 1741
rect 23663 1689 23715 1741
rect 23715 1689 23717 1741
rect 23661 1687 23717 1689
rect 23661 1637 23717 1639
rect 23661 1585 23663 1637
rect 23663 1585 23715 1637
rect 23715 1585 23717 1637
rect 23661 1583 23717 1585
rect 24301 1741 24357 1743
rect 24301 1689 24303 1741
rect 24303 1689 24355 1741
rect 24355 1689 24357 1741
rect 24301 1687 24357 1689
rect 24301 1637 24357 1639
rect 24301 1585 24303 1637
rect 24303 1585 24355 1637
rect 24355 1585 24357 1637
rect 24301 1583 24357 1585
rect 24941 1741 24997 1743
rect 24941 1689 24943 1741
rect 24943 1689 24995 1741
rect 24995 1689 24997 1741
rect 24941 1687 24997 1689
rect 24941 1637 24997 1639
rect 24941 1585 24943 1637
rect 24943 1585 24995 1637
rect 24995 1585 24997 1637
rect 24941 1583 24997 1585
rect 22270 855 22326 911
rect 22374 855 22430 911
rect 22478 855 22534 911
rect 22270 751 22326 807
rect 22374 751 22430 807
rect 22478 751 22534 807
rect 22270 647 22326 703
rect 22374 647 22430 703
rect 22478 647 22534 703
rect 23661 805 23717 807
rect 23661 753 23663 805
rect 23663 753 23715 805
rect 23715 753 23717 805
rect 23661 751 23717 753
rect 23661 701 23717 703
rect 23661 649 23663 701
rect 23663 649 23715 701
rect 23715 649 23717 701
rect 23661 647 23717 649
rect 22270 313 22326 369
rect 22374 313 22430 369
rect 22478 313 22534 369
rect 22270 209 22326 265
rect 22374 209 22430 265
rect 22478 209 22534 265
rect 22270 105 22326 161
rect 22374 105 22430 161
rect 22478 105 22534 161
rect 20972 -1017 21028 -961
rect 21076 -1017 21132 -961
rect 21180 -1017 21236 -961
rect 18509 -1067 18565 -1065
rect 18509 -1119 18511 -1067
rect 18511 -1119 18563 -1067
rect 18563 -1119 18565 -1067
rect 18509 -1121 18565 -1119
rect 18509 -1171 18565 -1169
rect 18509 -1223 18511 -1171
rect 18511 -1223 18563 -1171
rect 18563 -1223 18565 -1171
rect 18509 -1225 18565 -1223
rect 19149 -1067 19205 -1065
rect 19149 -1119 19151 -1067
rect 19151 -1119 19203 -1067
rect 19203 -1119 19205 -1067
rect 19149 -1121 19205 -1119
rect 19149 -1171 19205 -1169
rect 19149 -1223 19151 -1171
rect 19151 -1223 19203 -1171
rect 19203 -1223 19205 -1171
rect 19149 -1225 19205 -1223
rect 19789 -1067 19845 -1065
rect 19789 -1119 19791 -1067
rect 19791 -1119 19843 -1067
rect 19843 -1119 19845 -1067
rect 19789 -1121 19845 -1119
rect 19789 -1171 19845 -1169
rect 19789 -1223 19791 -1171
rect 19791 -1223 19843 -1171
rect 19843 -1223 19845 -1171
rect 19789 -1225 19845 -1223
rect 20972 -1121 21028 -1065
rect 21076 -1121 21132 -1065
rect 21180 -1121 21236 -1065
rect 20972 -1225 21028 -1169
rect 21076 -1225 21132 -1169
rect 21180 -1225 21236 -1169
rect 23981 1199 24037 1201
rect 23981 1147 23983 1199
rect 23983 1147 24035 1199
rect 24035 1147 24037 1199
rect 23981 1145 24037 1147
rect 23981 1095 24037 1097
rect 23981 1043 23983 1095
rect 23983 1043 24035 1095
rect 24035 1043 24037 1095
rect 23981 1041 24037 1043
rect 23981 263 24037 265
rect 23981 211 23983 263
rect 23983 211 24035 263
rect 24035 211 24037 263
rect 23981 209 24037 211
rect 23981 159 24037 161
rect 23981 107 23983 159
rect 23983 107 24035 159
rect 24035 107 24037 159
rect 23981 105 24037 107
rect 24301 805 24357 807
rect 24301 753 24303 805
rect 24303 753 24355 805
rect 24355 753 24357 805
rect 24301 751 24357 753
rect 24301 701 24357 703
rect 24301 649 24303 701
rect 24303 649 24355 701
rect 24355 649 24357 701
rect 24301 647 24357 649
rect 24621 1199 24677 1201
rect 24621 1147 24623 1199
rect 24623 1147 24675 1199
rect 24675 1147 24677 1199
rect 24621 1145 24677 1147
rect 24621 1095 24677 1097
rect 24621 1043 24623 1095
rect 24623 1043 24675 1095
rect 24675 1043 24677 1095
rect 24621 1041 24677 1043
rect 24941 805 24997 807
rect 24941 753 24943 805
rect 24943 753 24995 805
rect 24995 753 24997 805
rect 24941 751 24997 753
rect 24941 701 24997 703
rect 24941 649 24943 701
rect 24943 649 24995 701
rect 24995 649 24997 701
rect 24941 647 24997 649
rect 24861 474 24917 476
rect 24861 422 24863 474
rect 24863 422 24915 474
rect 24915 422 24917 474
rect 24861 420 24917 422
rect 26085 420 26141 476
rect 24621 263 24677 265
rect 24621 211 24623 263
rect 24623 211 24675 263
rect 24675 211 24677 263
rect 24621 209 24677 211
rect 24621 159 24677 161
rect 24621 107 24623 159
rect 24623 107 24675 159
rect 24675 107 24677 159
rect 24621 105 24677 107
rect 23661 -131 23717 -129
rect 23661 -183 23663 -131
rect 23663 -183 23715 -131
rect 23715 -183 23717 -131
rect 23661 -185 23717 -183
rect 23661 -235 23717 -233
rect 23661 -287 23663 -235
rect 23663 -287 23715 -235
rect 23715 -287 23717 -235
rect 23661 -289 23717 -287
rect 24301 -131 24357 -129
rect 24301 -183 24303 -131
rect 24303 -183 24355 -131
rect 24355 -183 24357 -131
rect 24301 -185 24357 -183
rect 24301 -235 24357 -233
rect 24301 -287 24303 -235
rect 24303 -287 24355 -235
rect 24355 -287 24357 -235
rect 24301 -289 24357 -287
rect 24941 -131 24997 -129
rect 24941 -183 24943 -131
rect 24943 -183 24995 -131
rect 24995 -183 24997 -131
rect 24941 -185 24997 -183
rect 24941 -235 24997 -233
rect 24941 -287 24943 -235
rect 24943 -287 24995 -235
rect 24995 -287 24997 -235
rect 24941 -289 24997 -287
rect 22270 -1017 22326 -961
rect 22374 -1017 22430 -961
rect 22478 -1017 22534 -961
rect 23981 -673 24037 -671
rect 23981 -725 23983 -673
rect 23983 -725 24035 -673
rect 24035 -725 24037 -673
rect 23981 -727 24037 -725
rect 23981 -777 24037 -775
rect 23981 -829 23983 -777
rect 23983 -829 24035 -777
rect 24035 -829 24037 -777
rect 23981 -831 24037 -829
rect 24861 -462 24917 -460
rect 24861 -514 24863 -462
rect 24863 -514 24915 -462
rect 24915 -514 24917 -462
rect 24861 -516 24917 -514
rect 24621 -673 24677 -671
rect 24621 -725 24623 -673
rect 24623 -725 24675 -673
rect 24675 -725 24677 -673
rect 24621 -727 24677 -725
rect 24621 -777 24677 -775
rect 24621 -829 24623 -777
rect 24623 -829 24675 -777
rect 24675 -829 24677 -777
rect 24621 -831 24677 -829
rect 22270 -1121 22326 -1065
rect 22374 -1121 22430 -1065
rect 22478 -1121 22534 -1065
rect 22270 -1225 22326 -1169
rect 22374 -1225 22430 -1169
rect 22478 -1225 22534 -1169
rect 23661 -1067 23717 -1065
rect 23661 -1119 23663 -1067
rect 23663 -1119 23715 -1067
rect 23715 -1119 23717 -1067
rect 23661 -1121 23717 -1119
rect 23661 -1171 23717 -1169
rect 23661 -1223 23663 -1171
rect 23663 -1223 23715 -1171
rect 23715 -1223 23717 -1171
rect 23661 -1225 23717 -1223
rect 24301 -1067 24357 -1065
rect 24301 -1119 24303 -1067
rect 24303 -1119 24355 -1067
rect 24355 -1119 24357 -1067
rect 24301 -1121 24357 -1119
rect 24301 -1171 24357 -1169
rect 24301 -1223 24303 -1171
rect 24303 -1223 24355 -1171
rect 24355 -1223 24357 -1171
rect 24301 -1225 24357 -1223
rect 24941 -1067 24997 -1065
rect 24941 -1119 24943 -1067
rect 24943 -1119 24995 -1067
rect 24995 -1119 24997 -1067
rect 24941 -1121 24997 -1119
rect 24941 -1171 24997 -1169
rect 24941 -1223 24943 -1171
rect 24943 -1223 24995 -1171
rect 24995 -1223 24997 -1171
rect 24941 -1225 24997 -1223
rect 17365 -1452 17421 -1396
rect 18749 -1398 18805 -1396
rect 18749 -1450 18751 -1398
rect 18751 -1450 18803 -1398
rect 18803 -1450 18805 -1398
rect 18749 -1452 18805 -1450
rect 19389 -1398 19445 -1396
rect 19389 -1450 19391 -1398
rect 19391 -1450 19443 -1398
rect 19443 -1450 19445 -1398
rect 19389 -1452 19445 -1450
rect 24061 -1398 24117 -1396
rect 24061 -1450 24063 -1398
rect 24063 -1450 24115 -1398
rect 24115 -1450 24117 -1398
rect 24061 -1452 24117 -1450
rect 24701 -1398 24757 -1396
rect 24701 -1450 24703 -1398
rect 24703 -1450 24755 -1398
rect 24755 -1450 24757 -1398
rect 24701 -1452 24757 -1450
rect 27710 4248 27766 4250
rect 27710 4196 27712 4248
rect 27712 4196 27764 4248
rect 27764 4196 27766 4248
rect 27710 4194 27766 4196
rect 30742 4057 30798 4113
rect 30846 4057 30902 4113
rect 30950 4057 31006 4113
rect 27950 4007 28006 4009
rect 27950 3955 27952 4007
rect 27952 3955 28004 4007
rect 28004 3955 28006 4007
rect 27950 3953 28006 3955
rect 27950 3903 28006 3905
rect 27950 3851 27952 3903
rect 27952 3851 28004 3903
rect 28004 3851 28006 3903
rect 27950 3849 28006 3851
rect 28590 4007 28646 4009
rect 28590 3955 28592 4007
rect 28592 3955 28644 4007
rect 28644 3955 28646 4007
rect 28590 3953 28646 3955
rect 28590 3903 28646 3905
rect 28590 3851 28592 3903
rect 28592 3851 28644 3903
rect 28644 3851 28646 3903
rect 28590 3849 28646 3851
rect 30742 3953 30798 4009
rect 30846 3953 30902 4009
rect 30950 3953 31006 4009
rect 30742 3849 30798 3905
rect 30846 3849 30902 3905
rect 30950 3849 31006 3905
rect 30093 3663 30149 3719
rect 30197 3663 30253 3719
rect 30301 3663 30357 3719
rect 27630 3613 27686 3615
rect 27630 3561 27632 3613
rect 27632 3561 27684 3613
rect 27684 3561 27686 3613
rect 27630 3559 27686 3561
rect 27630 3509 27686 3511
rect 27630 3457 27632 3509
rect 27632 3457 27684 3509
rect 27684 3457 27686 3509
rect 27630 3455 27686 3457
rect 28270 3613 28326 3615
rect 28270 3561 28272 3613
rect 28272 3561 28324 3613
rect 28324 3561 28326 3613
rect 28270 3559 28326 3561
rect 28270 3509 28326 3511
rect 28270 3457 28272 3509
rect 28272 3457 28324 3509
rect 28324 3457 28326 3509
rect 28270 3455 28326 3457
rect 28910 3613 28966 3615
rect 28910 3561 28912 3613
rect 28912 3561 28964 3613
rect 28964 3561 28966 3613
rect 28910 3559 28966 3561
rect 28910 3509 28966 3511
rect 28910 3457 28912 3509
rect 28912 3457 28964 3509
rect 28964 3457 28966 3509
rect 28910 3455 28966 3457
rect 30093 3559 30149 3615
rect 30197 3559 30253 3615
rect 30301 3559 30357 3615
rect 30093 3455 30149 3511
rect 30197 3455 30253 3511
rect 30301 3455 30357 3511
rect 26285 2292 26342 2348
rect 26285 -516 26342 -460
rect 26486 3228 26542 3284
rect 27710 3282 27766 3284
rect 27710 3230 27712 3282
rect 27712 3230 27764 3282
rect 27764 3230 27766 3282
rect 27710 3228 27766 3230
rect 27950 3071 28006 3073
rect 27950 3019 27952 3071
rect 27952 3019 28004 3071
rect 28004 3019 28006 3071
rect 27950 3017 28006 3019
rect 27950 2967 28006 2969
rect 27950 2915 27952 2967
rect 27952 2915 28004 2967
rect 28004 2915 28006 2967
rect 27950 2913 28006 2915
rect 28590 3071 28646 3073
rect 28590 3019 28592 3071
rect 28592 3019 28644 3071
rect 28644 3019 28646 3071
rect 28590 3017 28646 3019
rect 28590 2967 28646 2969
rect 28590 2915 28592 2967
rect 28592 2915 28644 2967
rect 28644 2915 28646 2967
rect 28590 2913 28646 2915
rect 30093 3121 30149 3177
rect 30197 3121 30253 3177
rect 30301 3121 30357 3177
rect 30093 3017 30149 3073
rect 30197 3017 30253 3073
rect 30301 3017 30357 3073
rect 30093 2913 30149 2969
rect 30197 2913 30253 2969
rect 30301 2913 30357 2969
rect 27630 2677 27686 2679
rect 27630 2625 27632 2677
rect 27632 2625 27684 2677
rect 27684 2625 27686 2677
rect 27630 2623 27686 2625
rect 27630 2573 27686 2575
rect 27630 2521 27632 2573
rect 27632 2521 27684 2573
rect 27684 2521 27686 2573
rect 27630 2519 27686 2521
rect 28270 2677 28326 2679
rect 28270 2625 28272 2677
rect 28272 2625 28324 2677
rect 28324 2625 28326 2677
rect 28270 2623 28326 2625
rect 28270 2573 28326 2575
rect 28270 2521 28272 2573
rect 28272 2521 28324 2573
rect 28324 2521 28326 2573
rect 28270 2519 28326 2521
rect 28910 2677 28966 2679
rect 28910 2625 28912 2677
rect 28912 2625 28964 2677
rect 28964 2625 28966 2677
rect 28910 2623 28966 2625
rect 28910 2573 28966 2575
rect 28910 2521 28912 2573
rect 28912 2521 28964 2573
rect 28964 2521 28966 2573
rect 28910 2519 28966 2521
rect 27710 2346 27766 2348
rect 27710 2294 27712 2346
rect 27712 2294 27764 2346
rect 27764 2294 27766 2346
rect 27710 2292 27766 2294
rect 27950 2135 28006 2137
rect 27950 2083 27952 2135
rect 27952 2083 28004 2135
rect 28004 2083 28006 2135
rect 27950 2081 28006 2083
rect 27950 2031 28006 2033
rect 27950 1979 27952 2031
rect 27952 1979 28004 2031
rect 28004 1979 28006 2031
rect 27950 1977 28006 1979
rect 28590 2135 28646 2137
rect 28590 2083 28592 2135
rect 28592 2083 28644 2135
rect 28644 2083 28646 2135
rect 28590 2081 28646 2083
rect 28590 2031 28646 2033
rect 28590 1979 28592 2031
rect 28592 1979 28644 2031
rect 28644 1979 28646 2031
rect 28590 1977 28646 1979
rect 30093 1791 30149 1847
rect 30197 1791 30253 1847
rect 30301 1791 30357 1847
rect 27630 1741 27686 1743
rect 27630 1689 27632 1741
rect 27632 1689 27684 1741
rect 27684 1689 27686 1741
rect 27630 1687 27686 1689
rect 27630 1637 27686 1639
rect 27630 1585 27632 1637
rect 27632 1585 27684 1637
rect 27684 1585 27686 1637
rect 27630 1583 27686 1585
rect 28270 1741 28326 1743
rect 28270 1689 28272 1741
rect 28272 1689 28324 1741
rect 28324 1689 28326 1741
rect 28270 1687 28326 1689
rect 28270 1637 28326 1639
rect 28270 1585 28272 1637
rect 28272 1585 28324 1637
rect 28324 1585 28326 1637
rect 28270 1583 28326 1585
rect 28910 1741 28966 1743
rect 28910 1689 28912 1741
rect 28912 1689 28964 1741
rect 28964 1689 28966 1741
rect 28910 1687 28966 1689
rect 28910 1637 28966 1639
rect 28910 1585 28912 1637
rect 28912 1585 28964 1637
rect 28964 1585 28966 1637
rect 28910 1583 28966 1585
rect 30093 1687 30149 1743
rect 30197 1687 30253 1743
rect 30301 1687 30357 1743
rect 30093 1583 30149 1639
rect 30197 1583 30253 1639
rect 30301 1583 30357 1639
rect 27950 1199 28006 1201
rect 27950 1147 27952 1199
rect 27952 1147 28004 1199
rect 28004 1147 28006 1199
rect 27950 1145 28006 1147
rect 27950 1095 28006 1097
rect 27950 1043 27952 1095
rect 27952 1043 28004 1095
rect 28004 1043 28006 1095
rect 27950 1041 28006 1043
rect 27630 805 27686 807
rect 27630 753 27632 805
rect 27632 753 27684 805
rect 27684 753 27686 805
rect 27630 751 27686 753
rect 27630 701 27686 703
rect 27630 649 27632 701
rect 27632 649 27684 701
rect 27684 649 27686 701
rect 27630 647 27686 649
rect 26486 420 26542 476
rect 26085 -1452 26141 -1396
rect 27710 474 27766 476
rect 27710 422 27712 474
rect 27712 422 27764 474
rect 27764 422 27766 474
rect 27710 420 27766 422
rect 27950 263 28006 265
rect 27950 211 27952 263
rect 27952 211 28004 263
rect 28004 211 28006 263
rect 27950 209 28006 211
rect 27950 159 28006 161
rect 27950 107 27952 159
rect 27952 107 28004 159
rect 28004 107 28006 159
rect 27950 105 28006 107
rect 28270 805 28326 807
rect 28270 753 28272 805
rect 28272 753 28324 805
rect 28324 753 28326 805
rect 28270 751 28326 753
rect 28270 701 28326 703
rect 28270 649 28272 701
rect 28272 649 28324 701
rect 28324 649 28326 701
rect 28270 647 28326 649
rect 28590 1199 28646 1201
rect 28590 1147 28592 1199
rect 28592 1147 28644 1199
rect 28644 1147 28646 1199
rect 28590 1145 28646 1147
rect 28590 1095 28646 1097
rect 28590 1043 28592 1095
rect 28592 1043 28644 1095
rect 28644 1043 28646 1095
rect 28590 1041 28646 1043
rect 28590 263 28646 265
rect 28590 211 28592 263
rect 28592 211 28644 263
rect 28644 211 28646 263
rect 28590 209 28646 211
rect 28590 159 28646 161
rect 28590 107 28592 159
rect 28592 107 28644 159
rect 28644 107 28646 159
rect 28590 105 28646 107
rect 30093 855 30149 911
rect 30197 855 30253 911
rect 30301 855 30357 911
rect 28910 805 28966 807
rect 28910 753 28912 805
rect 28912 753 28964 805
rect 28964 753 28966 805
rect 28910 751 28966 753
rect 28910 701 28966 703
rect 28910 649 28912 701
rect 28912 649 28964 701
rect 28964 649 28966 701
rect 28910 647 28966 649
rect 30093 751 30149 807
rect 30197 751 30253 807
rect 30301 751 30357 807
rect 30093 647 30149 703
rect 30197 647 30253 703
rect 30301 647 30357 703
rect 30093 313 30149 369
rect 30197 313 30253 369
rect 30301 313 30357 369
rect 30093 209 30149 265
rect 30197 209 30253 265
rect 30301 209 30357 265
rect 30093 105 30149 161
rect 30197 105 30253 161
rect 30301 105 30357 161
rect 27630 -131 27686 -129
rect 27630 -183 27632 -131
rect 27632 -183 27684 -131
rect 27684 -183 27686 -131
rect 27630 -185 27686 -183
rect 27630 -235 27686 -233
rect 27630 -287 27632 -235
rect 27632 -287 27684 -235
rect 27684 -287 27686 -235
rect 27630 -289 27686 -287
rect 28270 -131 28326 -129
rect 28270 -183 28272 -131
rect 28272 -183 28324 -131
rect 28324 -183 28326 -131
rect 28270 -185 28326 -183
rect 28270 -235 28326 -233
rect 28270 -287 28272 -235
rect 28272 -287 28324 -235
rect 28324 -287 28326 -235
rect 28270 -289 28326 -287
rect 28910 -131 28966 -129
rect 28910 -183 28912 -131
rect 28912 -183 28964 -131
rect 28964 -183 28966 -131
rect 28910 -185 28966 -183
rect 28910 -235 28966 -233
rect 28910 -287 28912 -235
rect 28912 -287 28964 -235
rect 28964 -287 28966 -235
rect 28910 -289 28966 -287
rect 27710 -462 27766 -460
rect 27710 -514 27712 -462
rect 27712 -514 27764 -462
rect 27764 -514 27766 -462
rect 27710 -516 27766 -514
rect 27950 -673 28006 -671
rect 27950 -725 27952 -673
rect 27952 -725 28004 -673
rect 28004 -725 28006 -673
rect 27950 -727 28006 -725
rect 27950 -777 28006 -775
rect 27950 -829 27952 -777
rect 27952 -829 28004 -777
rect 28004 -829 28006 -777
rect 27950 -831 28006 -829
rect 28590 -673 28646 -671
rect 28590 -725 28592 -673
rect 28592 -725 28644 -673
rect 28644 -725 28646 -673
rect 28590 -727 28646 -725
rect 28590 -777 28646 -775
rect 28590 -829 28592 -777
rect 28592 -829 28644 -777
rect 28644 -829 28646 -777
rect 28590 -831 28646 -829
rect 30093 -1017 30149 -961
rect 30197 -1017 30253 -961
rect 30301 -1017 30357 -961
rect 27630 -1067 27686 -1065
rect 27630 -1119 27632 -1067
rect 27632 -1119 27684 -1067
rect 27684 -1119 27686 -1067
rect 27630 -1121 27686 -1119
rect 27630 -1171 27686 -1169
rect 27630 -1223 27632 -1171
rect 27632 -1223 27684 -1171
rect 27684 -1223 27686 -1171
rect 27630 -1225 27686 -1223
rect 28270 -1067 28326 -1065
rect 28270 -1119 28272 -1067
rect 28272 -1119 28324 -1067
rect 28324 -1119 28326 -1067
rect 28270 -1121 28326 -1119
rect 28270 -1171 28326 -1169
rect 28270 -1223 28272 -1171
rect 28272 -1223 28324 -1171
rect 28324 -1223 28326 -1171
rect 28270 -1225 28326 -1223
rect 28910 -1067 28966 -1065
rect 28910 -1119 28912 -1067
rect 28912 -1119 28964 -1067
rect 28964 -1119 28966 -1067
rect 28910 -1121 28966 -1119
rect 28910 -1171 28966 -1169
rect 28910 -1223 28912 -1171
rect 28912 -1223 28964 -1171
rect 28964 -1223 28966 -1171
rect 28910 -1225 28966 -1223
rect 30093 -1121 30149 -1065
rect 30197 -1121 30253 -1065
rect 30301 -1121 30357 -1065
rect 30093 -1225 30149 -1169
rect 30197 -1225 30253 -1169
rect 30301 -1225 30357 -1169
rect 30742 2727 30798 2783
rect 30846 2727 30902 2783
rect 30950 2727 31006 2783
rect 30742 2623 30798 2679
rect 30846 2623 30902 2679
rect 30950 2623 31006 2679
rect 31650 3663 31706 3719
rect 31754 3663 31810 3719
rect 31858 3663 31914 3719
rect 34102 3837 34158 3893
rect 34206 3837 34262 3893
rect 34310 3837 34366 3893
rect 34102 3733 34158 3789
rect 34206 3733 34262 3789
rect 34310 3733 34366 3789
rect 34102 3629 34158 3685
rect 34206 3629 34262 3685
rect 34310 3629 34366 3685
rect 38238 3837 38294 3893
rect 38342 3837 38398 3893
rect 38446 3837 38502 3893
rect 38238 3733 38294 3789
rect 38342 3733 38398 3789
rect 38446 3733 38502 3789
rect 38238 3629 38294 3685
rect 38342 3629 38398 3685
rect 38446 3629 38502 3685
rect 43798 3837 43854 3893
rect 43902 3837 43958 3893
rect 44006 3837 44062 3893
rect 43798 3733 43854 3789
rect 43902 3733 43958 3789
rect 44006 3733 44062 3789
rect 43798 3629 43854 3685
rect 43902 3629 43958 3685
rect 44006 3629 44062 3685
rect 47934 3837 47990 3893
rect 48038 3837 48094 3893
rect 48142 3837 48198 3893
rect 47934 3733 47990 3789
rect 48038 3733 48094 3789
rect 48142 3733 48198 3789
rect 47934 3629 47990 3685
rect 48038 3629 48094 3685
rect 48142 3629 48198 3685
rect 53494 3837 53550 3893
rect 53598 3837 53654 3893
rect 53702 3837 53758 3893
rect 53494 3733 53550 3789
rect 53598 3733 53654 3789
rect 53702 3733 53758 3789
rect 53494 3629 53550 3685
rect 53598 3629 53654 3685
rect 53702 3629 53758 3685
rect 57630 3837 57686 3893
rect 57734 3837 57790 3893
rect 57838 3837 57894 3893
rect 57630 3733 57686 3789
rect 57734 3733 57790 3789
rect 57838 3733 57894 3789
rect 57630 3629 57686 3685
rect 57734 3629 57790 3685
rect 57838 3629 57894 3685
rect 63190 3837 63246 3893
rect 63294 3837 63350 3893
rect 63398 3837 63454 3893
rect 63190 3733 63246 3789
rect 63294 3733 63350 3789
rect 63398 3733 63454 3789
rect 63190 3629 63246 3685
rect 63294 3629 63350 3685
rect 63398 3629 63454 3685
rect 66438 3891 66494 3893
rect 66438 3839 66440 3891
rect 66440 3839 66492 3891
rect 66492 3839 66494 3891
rect 66438 3837 66494 3839
rect 66542 3891 66598 3893
rect 66542 3839 66544 3891
rect 66544 3839 66596 3891
rect 66596 3839 66598 3891
rect 66542 3837 66598 3839
rect 66646 3891 66702 3893
rect 66646 3839 66648 3891
rect 66648 3839 66700 3891
rect 66700 3839 66702 3891
rect 66646 3837 66702 3839
rect 66438 3787 66494 3789
rect 66438 3735 66440 3787
rect 66440 3735 66492 3787
rect 66492 3735 66494 3787
rect 66438 3733 66494 3735
rect 66542 3787 66598 3789
rect 66542 3735 66544 3787
rect 66544 3735 66596 3787
rect 66596 3735 66598 3787
rect 66542 3733 66598 3735
rect 66646 3787 66702 3789
rect 66646 3735 66648 3787
rect 66648 3735 66700 3787
rect 66700 3735 66702 3787
rect 66646 3733 66702 3735
rect 66438 3683 66494 3685
rect 66438 3631 66440 3683
rect 66440 3631 66492 3683
rect 66492 3631 66494 3683
rect 66438 3629 66494 3631
rect 66542 3683 66598 3685
rect 66542 3631 66544 3683
rect 66544 3631 66596 3683
rect 66596 3631 66598 3683
rect 66542 3629 66598 3631
rect 66646 3683 66702 3685
rect 66646 3631 66648 3683
rect 66648 3631 66700 3683
rect 66700 3631 66702 3683
rect 66646 3629 66702 3631
rect 31650 3559 31706 3615
rect 31754 3559 31810 3615
rect 31858 3559 31914 3615
rect 31650 3455 31706 3511
rect 31754 3455 31810 3511
rect 31858 3455 31914 3511
rect 31650 3121 31706 3177
rect 31754 3121 31810 3177
rect 31858 3121 31914 3177
rect 31650 3017 31706 3073
rect 31754 3017 31810 3073
rect 31858 3017 31914 3073
rect 31650 2913 31706 2969
rect 31754 2913 31810 2969
rect 31858 2913 31914 2969
rect 30742 2519 30798 2575
rect 30846 2519 30902 2575
rect 30950 2519 31006 2575
rect 30742 2185 30798 2241
rect 30846 2185 30902 2241
rect 30950 2185 31006 2241
rect 30742 2081 30798 2137
rect 30846 2081 30902 2137
rect 30950 2081 31006 2137
rect 30742 1977 30798 2033
rect 30846 1977 30902 2033
rect 30950 1977 31006 2033
rect 30742 1249 30798 1305
rect 30846 1249 30902 1305
rect 30950 1249 31006 1305
rect 30742 1145 30798 1201
rect 30846 1145 30902 1201
rect 30950 1145 31006 1201
rect 30742 1041 30798 1097
rect 30846 1041 30902 1097
rect 30950 1041 31006 1097
rect 30742 -81 30798 -25
rect 30846 -81 30902 -25
rect 30950 -81 31006 -25
rect 30742 -185 30798 -129
rect 30846 -185 30902 -129
rect 30950 -185 31006 -129
rect 30742 -289 30798 -233
rect 30846 -289 30902 -233
rect 30950 -289 31006 -233
rect 30742 -623 30798 -567
rect 30846 -623 30902 -567
rect 30950 -623 31006 -567
rect 30742 -727 30798 -671
rect 30846 -727 30902 -671
rect 30950 -727 31006 -671
rect 30742 -831 30798 -775
rect 30846 -831 30902 -775
rect 30950 -831 31006 -775
rect 26486 -1452 26542 -1396
rect 27870 -1398 27926 -1396
rect 27870 -1450 27872 -1398
rect 27872 -1450 27924 -1398
rect 27924 -1450 27926 -1398
rect 27870 -1452 27926 -1450
rect 16643 -2721 16699 -2719
rect 16643 -2773 16645 -2721
rect 16645 -2773 16697 -2721
rect 16697 -2773 16699 -2721
rect 16643 -2775 16699 -2773
rect 16747 -2721 16803 -2719
rect 16747 -2773 16749 -2721
rect 16749 -2773 16801 -2721
rect 16801 -2773 16803 -2721
rect 16747 -2775 16803 -2773
rect 16851 -2721 16907 -2719
rect 16851 -2773 16853 -2721
rect 16853 -2773 16905 -2721
rect 16905 -2773 16907 -2721
rect 16851 -2775 16907 -2773
rect 16643 -2825 16699 -2823
rect 16643 -2877 16645 -2825
rect 16645 -2877 16697 -2825
rect 16697 -2877 16699 -2825
rect 16643 -2879 16699 -2877
rect 16747 -2825 16803 -2823
rect 16747 -2877 16749 -2825
rect 16749 -2877 16801 -2825
rect 16801 -2877 16803 -2825
rect 16747 -2879 16803 -2877
rect 16851 -2825 16907 -2823
rect 16851 -2877 16853 -2825
rect 16853 -2877 16905 -2825
rect 16905 -2877 16907 -2825
rect 16851 -2879 16907 -2877
rect 16643 -2929 16699 -2927
rect 16643 -2981 16645 -2929
rect 16645 -2981 16697 -2929
rect 16697 -2981 16699 -2929
rect 16643 -2983 16699 -2981
rect 16747 -2929 16803 -2927
rect 16747 -2981 16749 -2929
rect 16749 -2981 16801 -2929
rect 16801 -2981 16803 -2929
rect 16747 -2983 16803 -2981
rect 16851 -2929 16907 -2927
rect 16851 -2981 16853 -2929
rect 16853 -2981 16905 -2929
rect 16905 -2981 16907 -2929
rect 16851 -2983 16907 -2981
rect 29812 -2775 29868 -2719
rect 29916 -2775 29972 -2719
rect 30020 -2775 30076 -2719
rect 30124 -2775 30180 -2719
rect 30228 -2775 30284 -2719
rect 29812 -2879 29868 -2823
rect 29916 -2879 29972 -2823
rect 30020 -2879 30076 -2823
rect 30124 -2879 30180 -2823
rect 30228 -2879 30284 -2823
rect 29812 -2983 29868 -2927
rect 29916 -2983 29972 -2927
rect 30020 -2983 30076 -2927
rect 30124 -2983 30180 -2927
rect 30228 -2983 30284 -2927
rect 17080 -3063 17136 -3061
rect 17080 -3115 17082 -3063
rect 17082 -3115 17134 -3063
rect 17134 -3115 17136 -3063
rect 17080 -3117 17136 -3115
rect 17184 -3063 17240 -3061
rect 17184 -3115 17186 -3063
rect 17186 -3115 17238 -3063
rect 17238 -3115 17240 -3063
rect 17184 -3117 17240 -3115
rect 17288 -3063 17344 -3061
rect 17288 -3115 17290 -3063
rect 17290 -3115 17342 -3063
rect 17342 -3115 17344 -3063
rect 17288 -3117 17344 -3115
rect 17080 -3167 17136 -3165
rect 17080 -3219 17082 -3167
rect 17082 -3219 17134 -3167
rect 17134 -3219 17136 -3167
rect 17080 -3221 17136 -3219
rect 17184 -3167 17240 -3165
rect 17184 -3219 17186 -3167
rect 17186 -3219 17238 -3167
rect 17238 -3219 17240 -3167
rect 17184 -3221 17240 -3219
rect 17288 -3167 17344 -3165
rect 17288 -3219 17290 -3167
rect 17290 -3219 17342 -3167
rect 17342 -3219 17344 -3167
rect 17288 -3221 17344 -3219
rect 17080 -3271 17136 -3269
rect 17080 -3323 17082 -3271
rect 17082 -3323 17134 -3271
rect 17134 -3323 17136 -3271
rect 17080 -3325 17136 -3323
rect 17184 -3271 17240 -3269
rect 17184 -3323 17186 -3271
rect 17186 -3323 17238 -3271
rect 17238 -3323 17240 -3271
rect 17184 -3325 17240 -3323
rect 17288 -3271 17344 -3269
rect 17288 -3323 17290 -3271
rect 17290 -3323 17342 -3271
rect 17342 -3323 17344 -3271
rect 17288 -3325 17344 -3323
rect 29252 -3117 29308 -3061
rect 29356 -3117 29412 -3061
rect 29460 -3117 29516 -3061
rect 29564 -3117 29620 -3061
rect 29668 -3117 29724 -3061
rect 29252 -3221 29308 -3165
rect 29356 -3221 29412 -3165
rect 29460 -3221 29516 -3165
rect 29564 -3221 29620 -3165
rect 29668 -3221 29724 -3165
rect 29252 -3325 29308 -3269
rect 29356 -3325 29412 -3269
rect 29460 -3325 29516 -3269
rect 29564 -3325 29620 -3269
rect 29668 -3325 29724 -3269
rect 14210 -3448 14266 -3446
rect 14210 -3500 14212 -3448
rect 14212 -3500 14264 -3448
rect 14264 -3500 14266 -3448
rect 14210 -3502 14266 -3500
rect 14314 -3448 14370 -3446
rect 14314 -3500 14316 -3448
rect 14316 -3500 14368 -3448
rect 14368 -3500 14370 -3448
rect 14314 -3502 14370 -3500
rect 14210 -3552 14266 -3550
rect 14210 -3604 14212 -3552
rect 14212 -3604 14264 -3552
rect 14264 -3604 14266 -3552
rect 14210 -3606 14266 -3604
rect 14314 -3552 14370 -3550
rect 14314 -3604 14316 -3552
rect 14316 -3604 14368 -3552
rect 14368 -3604 14370 -3552
rect 14314 -3606 14370 -3604
rect 16858 -3713 16914 -3711
rect 16858 -3765 16860 -3713
rect 16860 -3765 16912 -3713
rect 16912 -3765 16914 -3713
rect 16858 -3767 16914 -3765
rect 16962 -3713 17018 -3711
rect 16962 -3765 16964 -3713
rect 16964 -3765 17016 -3713
rect 17016 -3765 17018 -3713
rect 16962 -3767 17018 -3765
rect 16858 -3817 16914 -3815
rect 16858 -3869 16860 -3817
rect 16860 -3869 16912 -3817
rect 16912 -3869 16914 -3817
rect 16858 -3871 16914 -3869
rect 16962 -3817 17018 -3815
rect 16962 -3869 16964 -3817
rect 16964 -3869 17016 -3817
rect 17016 -3869 17018 -3817
rect 16962 -3871 17018 -3869
rect 23644 -3767 23700 -3711
rect 23748 -3767 23804 -3711
rect 23644 -3871 23700 -3815
rect 23748 -3871 23804 -3815
rect 13736 -4747 13792 -4691
rect 13840 -4747 13896 -4691
rect 13944 -4747 14000 -4691
rect 13736 -4851 13792 -4795
rect 13840 -4851 13896 -4795
rect 13944 -4851 14000 -4795
rect 13736 -4955 13792 -4899
rect 13840 -4955 13896 -4899
rect 13944 -4955 14000 -4899
rect 12624 -6863 12680 -6861
rect 12624 -6915 12626 -6863
rect 12626 -6915 12678 -6863
rect 12678 -6915 12680 -6863
rect 12624 -6917 12680 -6915
rect 12624 -6967 12680 -6965
rect 12624 -7019 12626 -6967
rect 12626 -7019 12678 -6967
rect 12678 -7019 12680 -6967
rect 12624 -7021 12680 -7019
rect 12624 -7071 12680 -7069
rect 12624 -7123 12626 -7071
rect 12626 -7123 12678 -7071
rect 12678 -7123 12680 -7071
rect 12624 -7125 12680 -7123
rect 14576 -5595 14632 -5593
rect 14576 -5647 14578 -5595
rect 14578 -5647 14630 -5595
rect 14630 -5647 14632 -5595
rect 14576 -5649 14632 -5647
rect 14576 -5699 14632 -5697
rect 14576 -5751 14578 -5699
rect 14578 -5751 14630 -5699
rect 14630 -5751 14632 -5699
rect 14576 -5753 14632 -5751
rect 15184 -5595 15240 -5593
rect 15184 -5647 15186 -5595
rect 15186 -5647 15238 -5595
rect 15238 -5647 15240 -5595
rect 15184 -5649 15240 -5647
rect 15184 -5699 15240 -5697
rect 15184 -5751 15186 -5699
rect 15186 -5751 15238 -5699
rect 15238 -5751 15240 -5699
rect 15184 -5753 15240 -5751
rect 15792 -5595 15848 -5593
rect 15792 -5647 15794 -5595
rect 15794 -5647 15846 -5595
rect 15846 -5647 15848 -5595
rect 15792 -5649 15848 -5647
rect 15792 -5699 15848 -5697
rect 15792 -5751 15794 -5699
rect 15794 -5751 15846 -5699
rect 15846 -5751 15848 -5699
rect 15792 -5753 15848 -5751
rect 15080 -6049 15136 -5993
rect 15184 -6049 15240 -5993
rect 15288 -6049 15344 -5993
rect 15080 -6153 15136 -6097
rect 15184 -6153 15240 -6097
rect 15288 -6153 15344 -6097
rect 15080 -6257 15136 -6201
rect 15184 -6257 15240 -6201
rect 15288 -6257 15344 -6201
rect 14413 -6917 14469 -6861
rect 14517 -6917 14573 -6861
rect 14621 -6917 14677 -6861
rect 14413 -7021 14469 -6965
rect 14517 -7021 14573 -6965
rect 14621 -7021 14677 -6965
rect 14413 -7125 14469 -7069
rect 14517 -7125 14573 -7069
rect 14621 -7125 14677 -7069
rect 11542 -8030 11598 -8028
rect 11542 -8082 11544 -8030
rect 11544 -8082 11596 -8030
rect 11596 -8082 11598 -8030
rect 11542 -8084 11598 -8082
rect 11646 -8030 11702 -8028
rect 11646 -8082 11648 -8030
rect 11648 -8082 11700 -8030
rect 11700 -8082 11702 -8030
rect 11646 -8084 11702 -8082
rect 11542 -8134 11598 -8132
rect 11542 -8186 11544 -8134
rect 11544 -8186 11596 -8134
rect 11596 -8186 11598 -8134
rect 11542 -8188 11598 -8186
rect 11646 -8134 11702 -8132
rect 11646 -8186 11648 -8134
rect 11648 -8186 11700 -8134
rect 11700 -8186 11702 -8134
rect 11646 -8188 11702 -8186
rect 5144 -8336 5200 -8280
rect 5248 -8336 5304 -8280
rect 5144 -8440 5200 -8384
rect 5248 -8440 5304 -8384
rect 9837 -8336 9893 -8280
rect 9941 -8336 9997 -8280
rect 9837 -8440 9893 -8384
rect 9941 -8440 9997 -8384
rect 4668 -8656 4724 -8600
rect 4772 -8656 4828 -8600
rect 4668 -8760 4724 -8704
rect 4772 -8760 4828 -8704
rect 12724 -8656 12780 -8600
rect 12828 -8656 12884 -8600
rect 14413 -8439 14469 -8383
rect 14517 -8439 14573 -8383
rect 14621 -8439 14677 -8383
rect 14413 -8543 14469 -8487
rect 14517 -8543 14573 -8487
rect 14621 -8543 14677 -8487
rect 14413 -8647 14469 -8591
rect 14517 -8647 14573 -8591
rect 14621 -8647 14677 -8591
rect 21184 -4693 21240 -4691
rect 21184 -4745 21186 -4693
rect 21186 -4745 21238 -4693
rect 21238 -4745 21240 -4693
rect 21184 -4747 21240 -4745
rect 21184 -4797 21240 -4795
rect 21184 -4849 21186 -4797
rect 21186 -4849 21238 -4797
rect 21238 -4849 21240 -4797
rect 21184 -4851 21240 -4849
rect 21184 -4901 21240 -4899
rect 21184 -4953 21186 -4901
rect 21186 -4953 21238 -4901
rect 21238 -4953 21240 -4901
rect 21184 -4955 21240 -4953
rect 20094 -6049 20150 -5993
rect 20198 -6049 20254 -5993
rect 20302 -6049 20358 -5993
rect 20094 -6153 20150 -6097
rect 20198 -6153 20254 -6097
rect 20302 -6153 20358 -6097
rect 20094 -6257 20150 -6201
rect 20198 -6257 20254 -6201
rect 20302 -6257 20358 -6201
rect 29812 -5020 29868 -5018
rect 29812 -5072 29814 -5020
rect 29814 -5072 29866 -5020
rect 29866 -5072 29868 -5020
rect 29812 -5074 29868 -5072
rect 29916 -5020 29972 -5018
rect 29916 -5072 29918 -5020
rect 29918 -5072 29970 -5020
rect 29970 -5072 29972 -5020
rect 29916 -5074 29972 -5072
rect 30020 -5020 30076 -5018
rect 30020 -5072 30022 -5020
rect 30022 -5072 30074 -5020
rect 30074 -5072 30076 -5020
rect 30020 -5074 30076 -5072
rect 30124 -5020 30180 -5018
rect 30124 -5072 30126 -5020
rect 30126 -5072 30178 -5020
rect 30178 -5072 30180 -5020
rect 30124 -5074 30180 -5072
rect 30228 -5020 30284 -5018
rect 30228 -5072 30230 -5020
rect 30230 -5072 30282 -5020
rect 30282 -5072 30284 -5020
rect 30228 -5074 30284 -5072
rect 29812 -5124 29868 -5122
rect 29812 -5176 29814 -5124
rect 29814 -5176 29866 -5124
rect 29866 -5176 29868 -5124
rect 29812 -5178 29868 -5176
rect 29916 -5124 29972 -5122
rect 29916 -5176 29918 -5124
rect 29918 -5176 29970 -5124
rect 29970 -5176 29972 -5124
rect 29916 -5178 29972 -5176
rect 30020 -5124 30076 -5122
rect 30020 -5176 30022 -5124
rect 30022 -5176 30074 -5124
rect 30074 -5176 30076 -5124
rect 30020 -5178 30076 -5176
rect 30124 -5124 30180 -5122
rect 30124 -5176 30126 -5124
rect 30126 -5176 30178 -5124
rect 30178 -5176 30180 -5124
rect 30124 -5178 30180 -5176
rect 30228 -5124 30284 -5122
rect 30228 -5176 30230 -5124
rect 30230 -5176 30282 -5124
rect 30282 -5176 30284 -5124
rect 30228 -5178 30284 -5176
rect 29812 -5228 29868 -5226
rect 29812 -5280 29814 -5228
rect 29814 -5280 29866 -5228
rect 29866 -5280 29868 -5228
rect 29812 -5282 29868 -5280
rect 29916 -5228 29972 -5226
rect 29916 -5280 29918 -5228
rect 29918 -5280 29970 -5228
rect 29970 -5280 29972 -5228
rect 29916 -5282 29972 -5280
rect 30020 -5228 30076 -5226
rect 30020 -5280 30022 -5228
rect 30022 -5280 30074 -5228
rect 30074 -5280 30076 -5228
rect 30020 -5282 30076 -5280
rect 30124 -5228 30180 -5226
rect 30124 -5280 30126 -5228
rect 30126 -5280 30178 -5228
rect 30178 -5280 30180 -5228
rect 30124 -5282 30180 -5280
rect 30228 -5228 30284 -5226
rect 30228 -5280 30230 -5228
rect 30230 -5280 30282 -5228
rect 30282 -5280 30284 -5228
rect 30228 -5282 30284 -5280
rect 29812 -5332 29868 -5330
rect 29812 -5384 29814 -5332
rect 29814 -5384 29866 -5332
rect 29866 -5384 29868 -5332
rect 29812 -5386 29868 -5384
rect 29916 -5332 29972 -5330
rect 29916 -5384 29918 -5332
rect 29918 -5384 29970 -5332
rect 29970 -5384 29972 -5332
rect 29916 -5386 29972 -5384
rect 30020 -5332 30076 -5330
rect 30020 -5384 30022 -5332
rect 30022 -5384 30074 -5332
rect 30074 -5384 30076 -5332
rect 30020 -5386 30076 -5384
rect 30124 -5332 30180 -5330
rect 30124 -5384 30126 -5332
rect 30126 -5384 30178 -5332
rect 30178 -5384 30180 -5332
rect 30124 -5386 30180 -5384
rect 30228 -5332 30284 -5330
rect 30228 -5384 30230 -5332
rect 30230 -5384 30282 -5332
rect 30282 -5384 30284 -5332
rect 30228 -5386 30284 -5384
rect 29812 -5436 29868 -5434
rect 29812 -5488 29814 -5436
rect 29814 -5488 29866 -5436
rect 29866 -5488 29868 -5436
rect 29812 -5490 29868 -5488
rect 29916 -5436 29972 -5434
rect 29916 -5488 29918 -5436
rect 29918 -5488 29970 -5436
rect 29970 -5488 29972 -5436
rect 29916 -5490 29972 -5488
rect 30020 -5436 30076 -5434
rect 30020 -5488 30022 -5436
rect 30022 -5488 30074 -5436
rect 30074 -5488 30076 -5436
rect 30020 -5490 30076 -5488
rect 30124 -5436 30180 -5434
rect 30124 -5488 30126 -5436
rect 30126 -5488 30178 -5436
rect 30178 -5488 30180 -5436
rect 30124 -5490 30180 -5488
rect 30228 -5436 30284 -5434
rect 30228 -5488 30230 -5436
rect 30230 -5488 30282 -5436
rect 30282 -5488 30284 -5436
rect 30228 -5490 30284 -5488
rect 15080 -6917 15136 -6861
rect 15184 -6863 15240 -6861
rect 15184 -6915 15186 -6863
rect 15186 -6915 15238 -6863
rect 15238 -6915 15240 -6863
rect 15184 -6917 15240 -6915
rect 15288 -6917 15344 -6861
rect 15080 -7021 15136 -6965
rect 15184 -6967 15240 -6965
rect 15184 -7019 15186 -6967
rect 15186 -7019 15238 -6967
rect 15238 -7019 15240 -6967
rect 15184 -7021 15240 -7019
rect 15288 -7021 15344 -6965
rect 15080 -7125 15136 -7069
rect 15184 -7071 15240 -7069
rect 15184 -7123 15186 -7071
rect 15186 -7123 15238 -7071
rect 15238 -7123 15240 -7071
rect 15184 -7125 15240 -7123
rect 15288 -7125 15344 -7069
rect 12724 -8760 12780 -8704
rect 12828 -8760 12884 -8704
rect 15695 -6955 15751 -6899
rect 15799 -6955 15855 -6899
rect 15903 -6955 15959 -6899
rect 15695 -7059 15751 -7003
rect 15799 -7059 15855 -7003
rect 15903 -7059 15959 -7003
rect 15695 -7163 15751 -7107
rect 15799 -7163 15855 -7107
rect 15903 -7163 15959 -7107
rect 18624 -6901 18680 -6899
rect 18624 -6953 18626 -6901
rect 18626 -6953 18678 -6901
rect 18678 -6953 18680 -6901
rect 18624 -6955 18680 -6953
rect 18624 -7005 18680 -7003
rect 18624 -7057 18626 -7005
rect 18626 -7057 18678 -7005
rect 18678 -7057 18680 -7005
rect 18624 -7059 18680 -7057
rect 18624 -7109 18680 -7107
rect 18624 -7161 18626 -7109
rect 18626 -7161 18678 -7109
rect 18678 -7161 18680 -7109
rect 18624 -7163 18680 -7161
rect 18944 -6901 19000 -6899
rect 18944 -6953 18946 -6901
rect 18946 -6953 18998 -6901
rect 18998 -6953 19000 -6901
rect 18944 -6955 19000 -6953
rect 18944 -7005 19000 -7003
rect 18944 -7057 18946 -7005
rect 18946 -7057 18998 -7005
rect 18998 -7057 19000 -7005
rect 18944 -7059 19000 -7057
rect 18944 -7109 19000 -7107
rect 18944 -7161 18946 -7109
rect 18946 -7161 18998 -7109
rect 18998 -7161 19000 -7109
rect 18944 -7163 19000 -7161
rect 19264 -6901 19320 -6899
rect 19264 -6953 19266 -6901
rect 19266 -6953 19318 -6901
rect 19318 -6953 19320 -6901
rect 19264 -6955 19320 -6953
rect 19264 -7005 19320 -7003
rect 19264 -7057 19266 -7005
rect 19266 -7057 19318 -7005
rect 19318 -7057 19320 -7005
rect 19264 -7059 19320 -7057
rect 19264 -7109 19320 -7107
rect 19264 -7161 19266 -7109
rect 19266 -7161 19318 -7109
rect 19318 -7161 19320 -7109
rect 19264 -7163 19320 -7161
rect 19584 -6901 19640 -6899
rect 19584 -6953 19586 -6901
rect 19586 -6953 19638 -6901
rect 19638 -6953 19640 -6901
rect 19584 -6955 19640 -6953
rect 19584 -7005 19640 -7003
rect 19584 -7057 19586 -7005
rect 19586 -7057 19638 -7005
rect 19638 -7057 19640 -7005
rect 19584 -7059 19640 -7057
rect 19584 -7109 19640 -7107
rect 19584 -7161 19586 -7109
rect 19586 -7161 19638 -7109
rect 19638 -7161 19640 -7109
rect 19584 -7163 19640 -7161
rect 19904 -6901 19960 -6899
rect 19904 -6953 19906 -6901
rect 19906 -6953 19958 -6901
rect 19958 -6953 19960 -6901
rect 19904 -6955 19960 -6953
rect 19904 -7005 19960 -7003
rect 19904 -7057 19906 -7005
rect 19906 -7057 19958 -7005
rect 19958 -7057 19960 -7005
rect 19904 -7059 19960 -7057
rect 19904 -7109 19960 -7107
rect 19904 -7161 19906 -7109
rect 19906 -7161 19958 -7109
rect 19958 -7161 19960 -7109
rect 19904 -7163 19960 -7161
rect 20224 -6901 20280 -6899
rect 20224 -6953 20226 -6901
rect 20226 -6953 20278 -6901
rect 20278 -6953 20280 -6901
rect 20224 -6955 20280 -6953
rect 20224 -7005 20280 -7003
rect 20224 -7057 20226 -7005
rect 20226 -7057 20278 -7005
rect 20278 -7057 20280 -7005
rect 20224 -7059 20280 -7057
rect 20224 -7109 20280 -7107
rect 20224 -7161 20226 -7109
rect 20226 -7161 20278 -7109
rect 20278 -7161 20280 -7109
rect 20224 -7163 20280 -7161
rect 20544 -6901 20600 -6899
rect 20544 -6953 20546 -6901
rect 20546 -6953 20598 -6901
rect 20598 -6953 20600 -6901
rect 20544 -6955 20600 -6953
rect 20544 -7005 20600 -7003
rect 20544 -7057 20546 -7005
rect 20546 -7057 20598 -7005
rect 20598 -7057 20600 -7005
rect 20544 -7059 20600 -7057
rect 20544 -7109 20600 -7107
rect 20544 -7161 20546 -7109
rect 20546 -7161 20598 -7109
rect 20598 -7161 20600 -7109
rect 20544 -7163 20600 -7161
rect 29812 -7032 29868 -7030
rect 29812 -7084 29814 -7032
rect 29814 -7084 29866 -7032
rect 29866 -7084 29868 -7032
rect 29812 -7086 29868 -7084
rect 29916 -7032 29972 -7030
rect 29916 -7084 29918 -7032
rect 29918 -7084 29970 -7032
rect 29970 -7084 29972 -7032
rect 29916 -7086 29972 -7084
rect 30020 -7032 30076 -7030
rect 30020 -7084 30022 -7032
rect 30022 -7084 30074 -7032
rect 30074 -7084 30076 -7032
rect 30020 -7086 30076 -7084
rect 30124 -7032 30180 -7030
rect 30124 -7084 30126 -7032
rect 30126 -7084 30178 -7032
rect 30178 -7084 30180 -7032
rect 30124 -7086 30180 -7084
rect 30228 -7032 30284 -7030
rect 30228 -7084 30230 -7032
rect 30230 -7084 30282 -7032
rect 30282 -7084 30284 -7032
rect 30228 -7086 30284 -7084
rect 29812 -7136 29868 -7134
rect 29812 -7188 29814 -7136
rect 29814 -7188 29866 -7136
rect 29866 -7188 29868 -7136
rect 29812 -7190 29868 -7188
rect 29916 -7136 29972 -7134
rect 29916 -7188 29918 -7136
rect 29918 -7188 29970 -7136
rect 29970 -7188 29972 -7136
rect 29916 -7190 29972 -7188
rect 30020 -7136 30076 -7134
rect 30020 -7188 30022 -7136
rect 30022 -7188 30074 -7136
rect 30074 -7188 30076 -7136
rect 30020 -7190 30076 -7188
rect 30124 -7136 30180 -7134
rect 30124 -7188 30126 -7136
rect 30126 -7188 30178 -7136
rect 30178 -7188 30180 -7136
rect 30124 -7190 30180 -7188
rect 30228 -7136 30284 -7134
rect 30228 -7188 30230 -7136
rect 30230 -7188 30282 -7136
rect 30282 -7188 30284 -7136
rect 30228 -7190 30284 -7188
rect 29812 -7240 29868 -7238
rect 29812 -7292 29814 -7240
rect 29814 -7292 29866 -7240
rect 29866 -7292 29868 -7240
rect 29812 -7294 29868 -7292
rect 29916 -7240 29972 -7238
rect 29916 -7292 29918 -7240
rect 29918 -7292 29970 -7240
rect 29970 -7292 29972 -7240
rect 29916 -7294 29972 -7292
rect 30020 -7240 30076 -7238
rect 30020 -7292 30022 -7240
rect 30022 -7292 30074 -7240
rect 30074 -7292 30076 -7240
rect 30020 -7294 30076 -7292
rect 30124 -7240 30180 -7238
rect 30124 -7292 30126 -7240
rect 30126 -7292 30178 -7240
rect 30178 -7292 30180 -7240
rect 30124 -7294 30180 -7292
rect 30228 -7240 30284 -7238
rect 30228 -7292 30230 -7240
rect 30230 -7292 30282 -7240
rect 30282 -7292 30284 -7240
rect 30228 -7294 30284 -7292
rect 21155 -8385 21211 -8383
rect 21155 -8437 21157 -8385
rect 21157 -8437 21209 -8385
rect 21209 -8437 21211 -8385
rect 21155 -8439 21211 -8437
rect 21259 -8385 21315 -8383
rect 21259 -8437 21261 -8385
rect 21261 -8437 21313 -8385
rect 21313 -8437 21315 -8385
rect 21259 -8439 21315 -8437
rect 21363 -8385 21419 -8383
rect 21363 -8437 21365 -8385
rect 21365 -8437 21417 -8385
rect 21417 -8437 21419 -8385
rect 21363 -8439 21419 -8437
rect 21155 -8489 21211 -8487
rect 21155 -8541 21157 -8489
rect 21157 -8541 21209 -8489
rect 21209 -8541 21211 -8489
rect 21155 -8543 21211 -8541
rect 21259 -8489 21315 -8487
rect 21259 -8541 21261 -8489
rect 21261 -8541 21313 -8489
rect 21313 -8541 21315 -8489
rect 21259 -8543 21315 -8541
rect 21363 -8489 21419 -8487
rect 21363 -8541 21365 -8489
rect 21365 -8541 21417 -8489
rect 21417 -8541 21419 -8489
rect 21363 -8543 21419 -8541
rect 21155 -8593 21211 -8591
rect 21155 -8645 21157 -8593
rect 21157 -8645 21209 -8593
rect 21209 -8645 21211 -8593
rect 21155 -8647 21211 -8645
rect 21259 -8593 21315 -8591
rect 21259 -8645 21261 -8593
rect 21261 -8645 21313 -8593
rect 21313 -8645 21315 -8593
rect 21259 -8647 21315 -8645
rect 21363 -8593 21419 -8591
rect 21363 -8645 21365 -8593
rect 21365 -8645 21417 -8593
rect 21417 -8645 21419 -8593
rect 21363 -8647 21419 -8645
rect 23642 -8426 23698 -8370
rect 23746 -8426 23802 -8370
rect 23642 -8530 23698 -8474
rect 23746 -8530 23802 -8474
rect 23642 -8634 23698 -8578
rect 23746 -8634 23802 -8578
rect 18963 -8827 19019 -8771
rect 19067 -8827 19123 -8771
rect 19190 -8827 19246 -8771
rect 18963 -8931 19019 -8875
rect 19067 -8931 19123 -8875
rect 19190 -8931 19246 -8875
rect 18963 -9035 19019 -8979
rect 19067 -9035 19123 -8979
rect 19190 -9035 19246 -8979
rect 29812 -7344 29868 -7342
rect 29812 -7396 29814 -7344
rect 29814 -7396 29866 -7344
rect 29866 -7396 29868 -7344
rect 29812 -7398 29868 -7396
rect 29916 -7344 29972 -7342
rect 29916 -7396 29918 -7344
rect 29918 -7396 29970 -7344
rect 29970 -7396 29972 -7344
rect 29916 -7398 29972 -7396
rect 30020 -7344 30076 -7342
rect 30020 -7396 30022 -7344
rect 30022 -7396 30074 -7344
rect 30074 -7396 30076 -7344
rect 30020 -7398 30076 -7396
rect 30124 -7344 30180 -7342
rect 30124 -7396 30126 -7344
rect 30126 -7396 30178 -7344
rect 30178 -7396 30180 -7344
rect 30124 -7398 30180 -7396
rect 30228 -7344 30284 -7342
rect 30228 -7396 30230 -7344
rect 30230 -7396 30282 -7344
rect 30282 -7396 30284 -7344
rect 30228 -7398 30284 -7396
rect 29812 -7448 29868 -7446
rect 29812 -7500 29814 -7448
rect 29814 -7500 29866 -7448
rect 29866 -7500 29868 -7448
rect 29812 -7502 29868 -7500
rect 29916 -7448 29972 -7446
rect 29916 -7500 29918 -7448
rect 29918 -7500 29970 -7448
rect 29970 -7500 29972 -7448
rect 29916 -7502 29972 -7500
rect 30020 -7448 30076 -7446
rect 30020 -7500 30022 -7448
rect 30022 -7500 30074 -7448
rect 30074 -7500 30076 -7448
rect 30020 -7502 30076 -7500
rect 30124 -7448 30180 -7446
rect 30124 -7500 30126 -7448
rect 30126 -7500 30178 -7448
rect 30178 -7500 30180 -7448
rect 30124 -7502 30180 -7500
rect 30228 -7448 30284 -7446
rect 30228 -7500 30230 -7448
rect 30230 -7500 30282 -7448
rect 30282 -7500 30284 -7448
rect 30228 -7502 30284 -7500
rect 31270 2557 31326 2613
rect 31374 2557 31430 2613
rect 31478 2557 31534 2613
rect 31270 2453 31326 2509
rect 31374 2453 31430 2509
rect 31478 2453 31534 2509
rect 31270 2349 31326 2405
rect 31374 2349 31430 2405
rect 31478 2349 31534 2405
rect 31270 1103 31326 1159
rect 31374 1103 31430 1159
rect 31478 1103 31534 1159
rect 31270 999 31326 1055
rect 31374 999 31430 1055
rect 31478 999 31534 1055
rect 31270 895 31326 951
rect 31374 895 31430 951
rect 31478 895 31534 951
rect 31270 43 31326 99
rect 31374 43 31430 99
rect 31478 43 31534 99
rect 31270 -61 31326 -5
rect 31374 -61 31430 -5
rect 31478 -61 31534 -5
rect 31270 -165 31326 -109
rect 31374 -165 31430 -109
rect 31478 -165 31534 -109
rect 31270 -623 31326 -567
rect 31374 -623 31430 -567
rect 31478 -623 31534 -567
rect 31270 -727 31326 -671
rect 31374 -727 31430 -671
rect 31478 -727 31534 -671
rect 31270 -831 31326 -775
rect 31374 -831 31430 -775
rect 31478 -831 31534 -775
rect 33247 2507 33303 2509
rect 33247 2455 33249 2507
rect 33249 2455 33301 2507
rect 33301 2455 33303 2507
rect 33247 2453 33303 2455
rect 33247 2403 33303 2405
rect 33247 2351 33249 2403
rect 33249 2351 33301 2403
rect 33301 2351 33303 2403
rect 33247 2349 33303 2351
rect 33887 2507 33943 2509
rect 33887 2455 33889 2507
rect 33889 2455 33941 2507
rect 33941 2455 33943 2507
rect 33887 2453 33943 2455
rect 33887 2403 33943 2405
rect 33887 2351 33889 2403
rect 33889 2351 33941 2403
rect 33941 2351 33943 2403
rect 33887 2349 33943 2351
rect 31650 2163 31706 2219
rect 31754 2163 31810 2219
rect 31858 2163 31914 2219
rect 31650 2059 31706 2115
rect 31754 2059 31810 2115
rect 31858 2059 31914 2115
rect 31650 1955 31706 2011
rect 31754 1955 31810 2011
rect 31858 1955 31914 2011
rect 32926 2113 32982 2115
rect 32926 2061 32928 2113
rect 32928 2061 32980 2113
rect 32980 2061 32982 2113
rect 32926 2059 32982 2061
rect 32926 2009 32982 2011
rect 32926 1957 32928 2009
rect 32928 1957 32980 2009
rect 32980 1957 32982 2009
rect 32926 1955 32982 1957
rect 33566 2113 33622 2115
rect 33566 2061 33568 2113
rect 33568 2061 33620 2113
rect 33620 2061 33622 2113
rect 33566 2059 33622 2061
rect 33566 2009 33622 2011
rect 33566 1957 33568 2009
rect 33568 1957 33620 2009
rect 33620 1957 33622 2009
rect 33566 1955 33622 1957
rect 31650 1497 31706 1553
rect 31754 1497 31810 1553
rect 31858 1497 31914 1553
rect 34527 2507 34583 2509
rect 34527 2455 34529 2507
rect 34529 2455 34581 2507
rect 34581 2455 34583 2507
rect 34527 2453 34583 2455
rect 34527 2403 34583 2405
rect 34527 2351 34529 2403
rect 34529 2351 34581 2403
rect 34581 2351 34583 2403
rect 34527 2349 34583 2351
rect 35167 2507 35223 2509
rect 35167 2455 35169 2507
rect 35169 2455 35221 2507
rect 35221 2455 35223 2507
rect 35167 2453 35223 2455
rect 35167 2403 35223 2405
rect 35167 2351 35169 2403
rect 35169 2351 35221 2403
rect 35221 2351 35223 2403
rect 35167 2349 35223 2351
rect 37381 2507 37437 2509
rect 37381 2455 37383 2507
rect 37383 2455 37435 2507
rect 37435 2455 37437 2507
rect 37381 2453 37437 2455
rect 37381 2403 37437 2405
rect 37381 2351 37383 2403
rect 37383 2351 37435 2403
rect 37435 2351 37437 2403
rect 37381 2349 37437 2351
rect 38021 2507 38077 2509
rect 38021 2455 38023 2507
rect 38023 2455 38075 2507
rect 38075 2455 38077 2507
rect 38021 2453 38077 2455
rect 38021 2403 38077 2405
rect 38021 2351 38023 2403
rect 38023 2351 38075 2403
rect 38075 2351 38077 2403
rect 38021 2349 38077 2351
rect 34846 2113 34902 2115
rect 34846 2061 34848 2113
rect 34848 2061 34900 2113
rect 34900 2061 34902 2113
rect 34846 2059 34902 2061
rect 34846 2009 34902 2011
rect 34846 1957 34848 2009
rect 34848 1957 34900 2009
rect 34900 1957 34902 2009
rect 34846 1955 34902 1957
rect 35486 2113 35542 2115
rect 35486 2061 35488 2113
rect 35488 2061 35540 2113
rect 35540 2061 35542 2113
rect 35486 2059 35542 2061
rect 35486 2009 35542 2011
rect 35486 1957 35488 2009
rect 35488 1957 35540 2009
rect 35540 1957 35542 2009
rect 35486 1955 35542 1957
rect 37062 2113 37118 2115
rect 37062 2061 37064 2113
rect 37064 2061 37116 2113
rect 37116 2061 37118 2113
rect 37062 2059 37118 2061
rect 37062 2009 37118 2011
rect 37062 1957 37064 2009
rect 37064 1957 37116 2009
rect 37116 1957 37118 2009
rect 37062 1955 37118 1957
rect 37702 2113 37758 2115
rect 37702 2061 37704 2113
rect 37704 2061 37756 2113
rect 37756 2061 37758 2113
rect 37702 2059 37758 2061
rect 37702 2009 37758 2011
rect 37702 1957 37704 2009
rect 37704 1957 37756 2009
rect 37756 1957 37758 2009
rect 37702 1955 37758 1957
rect 31650 1393 31706 1449
rect 31754 1393 31810 1449
rect 31858 1393 31914 1449
rect 31650 1289 31706 1345
rect 31754 1289 31810 1345
rect 31858 1289 31914 1345
rect 33247 1447 33303 1449
rect 33247 1395 33249 1447
rect 33249 1395 33301 1447
rect 33301 1395 33303 1447
rect 33247 1393 33303 1395
rect 33247 1343 33303 1345
rect 33247 1291 33249 1343
rect 33249 1291 33301 1343
rect 33301 1291 33303 1343
rect 33247 1289 33303 1291
rect 33887 1447 33943 1449
rect 33887 1395 33889 1447
rect 33889 1395 33941 1447
rect 33941 1395 33943 1447
rect 33887 1393 33943 1395
rect 33887 1343 33943 1345
rect 33887 1291 33889 1343
rect 33889 1291 33941 1343
rect 33941 1291 33943 1343
rect 33887 1289 33943 1291
rect 32926 1053 32982 1055
rect 32926 1001 32928 1053
rect 32928 1001 32980 1053
rect 32980 1001 32982 1053
rect 32926 999 32982 1001
rect 32926 949 32982 951
rect 32926 897 32928 949
rect 32928 897 32980 949
rect 32980 897 32982 949
rect 32926 895 32982 897
rect 33566 1053 33622 1055
rect 33566 1001 33568 1053
rect 33568 1001 33620 1053
rect 33620 1001 33622 1053
rect 33566 999 33622 1001
rect 33566 949 33622 951
rect 33566 897 33568 949
rect 33568 897 33620 949
rect 33620 897 33622 949
rect 33566 895 33622 897
rect 31650 437 31706 493
rect 31754 437 31810 493
rect 31858 437 31914 493
rect 40997 2557 41053 2613
rect 41101 2557 41157 2613
rect 41205 2557 41261 2613
rect 38661 2507 38717 2509
rect 38661 2455 38663 2507
rect 38663 2455 38715 2507
rect 38715 2455 38717 2507
rect 38661 2453 38717 2455
rect 38661 2403 38717 2405
rect 38661 2351 38663 2403
rect 38663 2351 38715 2403
rect 38715 2351 38717 2403
rect 38661 2349 38717 2351
rect 39301 2507 39357 2509
rect 39301 2455 39303 2507
rect 39303 2455 39355 2507
rect 39355 2455 39357 2507
rect 39301 2453 39357 2455
rect 39301 2403 39357 2405
rect 39301 2351 39303 2403
rect 39303 2351 39355 2403
rect 39355 2351 39357 2403
rect 39301 2349 39357 2351
rect 40997 2453 41053 2509
rect 41101 2453 41157 2509
rect 41205 2453 41261 2509
rect 40997 2349 41053 2405
rect 41101 2349 41157 2405
rect 41205 2349 41261 2405
rect 40636 2163 40692 2219
rect 40740 2163 40796 2219
rect 40844 2163 40900 2219
rect 38982 2113 39038 2115
rect 38982 2061 38984 2113
rect 38984 2061 39036 2113
rect 39036 2061 39038 2113
rect 38982 2059 39038 2061
rect 38982 2009 39038 2011
rect 38982 1957 38984 2009
rect 38984 1957 39036 2009
rect 39036 1957 39038 2009
rect 38982 1955 39038 1957
rect 39622 2113 39678 2115
rect 39622 2061 39624 2113
rect 39624 2061 39676 2113
rect 39676 2061 39678 2113
rect 39622 2059 39678 2061
rect 39622 2009 39678 2011
rect 39622 1957 39624 2009
rect 39624 1957 39676 2009
rect 39676 1957 39678 2009
rect 39622 1955 39678 1957
rect 40636 2059 40692 2115
rect 40740 2059 40796 2115
rect 40844 2059 40900 2115
rect 40636 1955 40692 2011
rect 40740 1955 40796 2011
rect 40844 1955 40900 2011
rect 34527 1447 34583 1449
rect 34527 1395 34529 1447
rect 34529 1395 34581 1447
rect 34581 1395 34583 1447
rect 34527 1393 34583 1395
rect 34527 1343 34583 1345
rect 34527 1291 34529 1343
rect 34529 1291 34581 1343
rect 34581 1291 34583 1343
rect 34527 1289 34583 1291
rect 35167 1447 35223 1449
rect 35167 1395 35169 1447
rect 35169 1395 35221 1447
rect 35221 1395 35223 1447
rect 35167 1393 35223 1395
rect 35167 1343 35223 1345
rect 35167 1291 35169 1343
rect 35169 1291 35221 1343
rect 35221 1291 35223 1343
rect 35167 1289 35223 1291
rect 37381 1447 37437 1449
rect 37381 1395 37383 1447
rect 37383 1395 37435 1447
rect 37435 1395 37437 1447
rect 37381 1393 37437 1395
rect 37381 1343 37437 1345
rect 37381 1291 37383 1343
rect 37383 1291 37435 1343
rect 37435 1291 37437 1343
rect 37381 1289 37437 1291
rect 38021 1447 38077 1449
rect 38021 1395 38023 1447
rect 38023 1395 38075 1447
rect 38075 1395 38077 1447
rect 38021 1393 38077 1395
rect 38021 1343 38077 1345
rect 38021 1291 38023 1343
rect 38023 1291 38075 1343
rect 38075 1291 38077 1343
rect 38021 1289 38077 1291
rect 34846 1053 34902 1055
rect 34846 1001 34848 1053
rect 34848 1001 34900 1053
rect 34900 1001 34902 1053
rect 34846 999 34902 1001
rect 34846 949 34902 951
rect 34846 897 34848 949
rect 34848 897 34900 949
rect 34900 897 34902 949
rect 34846 895 34902 897
rect 35486 1053 35542 1055
rect 35486 1001 35488 1053
rect 35488 1001 35540 1053
rect 35540 1001 35542 1053
rect 35486 999 35542 1001
rect 35486 949 35542 951
rect 35486 897 35488 949
rect 35488 897 35540 949
rect 35540 897 35542 949
rect 35486 895 35542 897
rect 37062 1053 37118 1055
rect 37062 1001 37064 1053
rect 37064 1001 37116 1053
rect 37116 1001 37118 1053
rect 37062 999 37118 1001
rect 37062 949 37118 951
rect 37062 897 37064 949
rect 37064 897 37116 949
rect 37116 897 37118 949
rect 37062 895 37118 897
rect 37702 1053 37758 1055
rect 37702 1001 37704 1053
rect 37704 1001 37756 1053
rect 37756 1001 37758 1053
rect 37702 999 37758 1001
rect 37702 949 37758 951
rect 37702 897 37704 949
rect 37704 897 37756 949
rect 37756 897 37758 949
rect 37702 895 37758 897
rect 31650 333 31706 389
rect 31754 333 31810 389
rect 31858 333 31914 389
rect 31650 229 31706 285
rect 31754 229 31810 285
rect 31858 229 31914 285
rect 30742 -8426 30798 -8370
rect 30846 -8426 30902 -8370
rect 30950 -8426 31006 -8370
rect 30742 -8530 30798 -8474
rect 30846 -8530 30902 -8474
rect 30950 -8530 31006 -8474
rect 30742 -8634 30798 -8578
rect 30846 -8634 30902 -8578
rect 30950 -8634 31006 -8578
rect 33247 387 33303 389
rect 33247 335 33249 387
rect 33249 335 33301 387
rect 33301 335 33303 387
rect 33247 333 33303 335
rect 33247 283 33303 285
rect 33247 231 33249 283
rect 33249 231 33301 283
rect 33301 231 33303 283
rect 33247 229 33303 231
rect 33887 387 33943 389
rect 33887 335 33889 387
rect 33889 335 33941 387
rect 33941 335 33943 387
rect 33887 333 33943 335
rect 33887 283 33943 285
rect 33887 231 33889 283
rect 33889 231 33941 283
rect 33941 231 33943 283
rect 33887 229 33943 231
rect 32926 -7 32982 -5
rect 32926 -59 32928 -7
rect 32928 -59 32980 -7
rect 32980 -59 32982 -7
rect 32926 -61 32982 -59
rect 32926 -111 32982 -109
rect 32926 -163 32928 -111
rect 32928 -163 32980 -111
rect 32980 -163 32982 -111
rect 32926 -165 32982 -163
rect 33566 -7 33622 -5
rect 33566 -59 33568 -7
rect 33568 -59 33620 -7
rect 33620 -59 33622 -7
rect 33566 -61 33622 -59
rect 33566 -111 33622 -109
rect 33566 -163 33568 -111
rect 33568 -163 33620 -111
rect 33620 -163 33622 -111
rect 33566 -165 33622 -163
rect 40636 1497 40692 1553
rect 40740 1497 40796 1553
rect 40844 1497 40900 1553
rect 38661 1447 38717 1449
rect 38661 1395 38663 1447
rect 38663 1395 38715 1447
rect 38715 1395 38717 1447
rect 38661 1393 38717 1395
rect 38661 1343 38717 1345
rect 38661 1291 38663 1343
rect 38663 1291 38715 1343
rect 38715 1291 38717 1343
rect 38661 1289 38717 1291
rect 39301 1447 39357 1449
rect 39301 1395 39303 1447
rect 39303 1395 39355 1447
rect 39355 1395 39357 1447
rect 39301 1393 39357 1395
rect 39301 1343 39357 1345
rect 39301 1291 39303 1343
rect 39303 1291 39355 1343
rect 39355 1291 39357 1343
rect 39301 1289 39357 1291
rect 40636 1393 40692 1449
rect 40740 1393 40796 1449
rect 40844 1393 40900 1449
rect 40636 1289 40692 1345
rect 40740 1289 40796 1345
rect 40844 1289 40900 1345
rect 38982 1053 39038 1055
rect 38982 1001 38984 1053
rect 38984 1001 39036 1053
rect 39036 1001 39038 1053
rect 38982 999 39038 1001
rect 38982 949 39038 951
rect 38982 897 38984 949
rect 38984 897 39036 949
rect 39036 897 39038 949
rect 38982 895 39038 897
rect 39622 1053 39678 1055
rect 39622 1001 39624 1053
rect 39624 1001 39676 1053
rect 39676 1001 39678 1053
rect 39622 999 39678 1001
rect 39622 949 39678 951
rect 39622 897 39624 949
rect 39624 897 39676 949
rect 39676 897 39678 949
rect 39622 895 39678 897
rect 34527 387 34583 389
rect 34527 335 34529 387
rect 34529 335 34581 387
rect 34581 335 34583 387
rect 34527 333 34583 335
rect 34527 283 34583 285
rect 34527 231 34529 283
rect 34529 231 34581 283
rect 34581 231 34583 283
rect 34527 229 34583 231
rect 35167 387 35223 389
rect 35167 335 35169 387
rect 35169 335 35221 387
rect 35221 335 35223 387
rect 35167 333 35223 335
rect 35167 283 35223 285
rect 35167 231 35169 283
rect 35169 231 35221 283
rect 35221 231 35223 283
rect 35167 229 35223 231
rect 37381 387 37437 389
rect 37381 335 37383 387
rect 37383 335 37435 387
rect 37435 335 37437 387
rect 37381 333 37437 335
rect 37381 283 37437 285
rect 37381 231 37383 283
rect 37383 231 37435 283
rect 37435 231 37437 283
rect 37381 229 37437 231
rect 38021 387 38077 389
rect 38021 335 38023 387
rect 38023 335 38075 387
rect 38075 335 38077 387
rect 38021 333 38077 335
rect 38021 283 38077 285
rect 38021 231 38023 283
rect 38023 231 38075 283
rect 38075 231 38077 283
rect 38021 229 38077 231
rect 34846 -7 34902 -5
rect 34846 -59 34848 -7
rect 34848 -59 34900 -7
rect 34900 -59 34902 -7
rect 34846 -61 34902 -59
rect 34846 -111 34902 -109
rect 34846 -163 34848 -111
rect 34848 -163 34900 -111
rect 34900 -163 34902 -111
rect 34846 -165 34902 -163
rect 35486 -7 35542 -5
rect 35486 -59 35488 -7
rect 35488 -59 35540 -7
rect 35540 -59 35542 -7
rect 35486 -61 35542 -59
rect 35486 -111 35542 -109
rect 35486 -163 35488 -111
rect 35488 -163 35540 -111
rect 35540 -163 35542 -111
rect 35486 -165 35542 -163
rect 37062 -7 37118 -5
rect 37062 -59 37064 -7
rect 37064 -59 37116 -7
rect 37116 -59 37118 -7
rect 37062 -61 37118 -59
rect 37062 -111 37118 -109
rect 37062 -163 37064 -111
rect 37064 -163 37116 -111
rect 37116 -163 37118 -111
rect 37062 -165 37118 -163
rect 37702 -7 37758 -5
rect 37702 -59 37704 -7
rect 37704 -59 37756 -7
rect 37756 -59 37758 -7
rect 37702 -61 37758 -59
rect 37702 -111 37758 -109
rect 37702 -163 37704 -111
rect 37704 -163 37756 -111
rect 37756 -163 37758 -111
rect 37702 -165 37758 -163
rect 33247 -673 33303 -671
rect 33247 -725 33249 -673
rect 33249 -725 33301 -673
rect 33301 -725 33303 -673
rect 33247 -727 33303 -725
rect 33247 -777 33303 -775
rect 33247 -829 33249 -777
rect 33249 -829 33301 -777
rect 33301 -829 33303 -777
rect 33247 -831 33303 -829
rect 33887 -673 33943 -671
rect 33887 -725 33889 -673
rect 33889 -725 33941 -673
rect 33941 -725 33943 -673
rect 33887 -727 33943 -725
rect 33887 -777 33943 -775
rect 33887 -829 33889 -777
rect 33889 -829 33941 -777
rect 33941 -829 33943 -777
rect 33887 -831 33943 -829
rect 31650 -1017 31706 -961
rect 31754 -1017 31810 -961
rect 31858 -1017 31914 -961
rect 31650 -1121 31706 -1065
rect 31754 -1121 31810 -1065
rect 31858 -1121 31914 -1065
rect 31650 -1225 31706 -1169
rect 31754 -1225 31810 -1169
rect 31858 -1225 31914 -1169
rect 24092 -8827 24148 -8771
rect 24196 -8827 24252 -8771
rect 24092 -8931 24148 -8875
rect 24196 -8931 24252 -8875
rect 24092 -9035 24148 -8979
rect 24196 -9035 24252 -8979
rect 32926 -1067 32982 -1065
rect 32926 -1119 32928 -1067
rect 32928 -1119 32980 -1067
rect 32980 -1119 32982 -1067
rect 32926 -1121 32982 -1119
rect 32926 -1171 32982 -1169
rect 32926 -1223 32928 -1171
rect 32928 -1223 32980 -1171
rect 32980 -1223 32982 -1171
rect 32926 -1225 32982 -1223
rect 33566 -1067 33622 -1065
rect 33566 -1119 33568 -1067
rect 33568 -1119 33620 -1067
rect 33620 -1119 33622 -1067
rect 33566 -1121 33622 -1119
rect 33566 -1171 33622 -1169
rect 33566 -1223 33568 -1171
rect 33568 -1223 33620 -1171
rect 33620 -1223 33622 -1171
rect 33566 -1225 33622 -1223
rect 40636 437 40692 493
rect 40740 437 40796 493
rect 40844 437 40900 493
rect 38661 387 38717 389
rect 38661 335 38663 387
rect 38663 335 38715 387
rect 38715 335 38717 387
rect 38661 333 38717 335
rect 38661 283 38717 285
rect 38661 231 38663 283
rect 38663 231 38715 283
rect 38715 231 38717 283
rect 38661 229 38717 231
rect 39301 387 39357 389
rect 39301 335 39303 387
rect 39303 335 39355 387
rect 39355 335 39357 387
rect 39301 333 39357 335
rect 39301 283 39357 285
rect 39301 231 39303 283
rect 39303 231 39355 283
rect 39355 231 39357 283
rect 39301 229 39357 231
rect 40636 333 40692 389
rect 40740 333 40796 389
rect 40844 333 40900 389
rect 40636 229 40692 285
rect 40740 229 40796 285
rect 40844 229 40900 285
rect 38982 -7 39038 -5
rect 38982 -59 38984 -7
rect 38984 -59 39036 -7
rect 39036 -59 39038 -7
rect 38982 -61 39038 -59
rect 38982 -111 39038 -109
rect 38982 -163 38984 -111
rect 38984 -163 39036 -111
rect 39036 -163 39038 -111
rect 38982 -165 39038 -163
rect 39622 -7 39678 -5
rect 39622 -59 39624 -7
rect 39624 -59 39676 -7
rect 39676 -59 39678 -7
rect 39622 -61 39678 -59
rect 39622 -111 39678 -109
rect 39622 -163 39624 -111
rect 39624 -163 39676 -111
rect 39676 -163 39678 -111
rect 39622 -165 39678 -163
rect 34527 -673 34583 -671
rect 34527 -725 34529 -673
rect 34529 -725 34581 -673
rect 34581 -725 34583 -673
rect 34527 -727 34583 -725
rect 34527 -777 34583 -775
rect 34527 -829 34529 -777
rect 34529 -829 34581 -777
rect 34581 -829 34583 -777
rect 34527 -831 34583 -829
rect 35167 -673 35223 -671
rect 35167 -725 35169 -673
rect 35169 -725 35221 -673
rect 35221 -725 35223 -673
rect 35167 -727 35223 -725
rect 35167 -777 35223 -775
rect 35167 -829 35169 -777
rect 35169 -829 35221 -777
rect 35221 -829 35223 -777
rect 35167 -831 35223 -829
rect 37381 -673 37437 -671
rect 37381 -725 37383 -673
rect 37383 -725 37435 -673
rect 37435 -725 37437 -673
rect 37381 -727 37437 -725
rect 37381 -777 37437 -775
rect 37381 -829 37383 -777
rect 37383 -829 37435 -777
rect 37435 -829 37437 -777
rect 37381 -831 37437 -829
rect 38021 -673 38077 -671
rect 38021 -725 38023 -673
rect 38023 -725 38075 -673
rect 38075 -725 38077 -673
rect 38021 -727 38077 -725
rect 38021 -777 38077 -775
rect 38021 -829 38023 -777
rect 38023 -829 38075 -777
rect 38075 -829 38077 -777
rect 38021 -831 38077 -829
rect 38661 -673 38717 -671
rect 38661 -725 38663 -673
rect 38663 -725 38715 -673
rect 38715 -725 38717 -673
rect 38661 -727 38717 -725
rect 38661 -777 38717 -775
rect 38661 -829 38663 -777
rect 38663 -829 38715 -777
rect 38715 -829 38717 -777
rect 38661 -831 38717 -829
rect 39301 -673 39357 -671
rect 39301 -725 39303 -673
rect 39303 -725 39355 -673
rect 39355 -725 39357 -673
rect 39301 -727 39357 -725
rect 39301 -777 39357 -775
rect 39301 -829 39303 -777
rect 39303 -829 39355 -777
rect 39355 -829 39357 -777
rect 39301 -831 39357 -829
rect 42943 2507 42999 2509
rect 42943 2455 42945 2507
rect 42945 2455 42997 2507
rect 42997 2455 42999 2507
rect 42943 2453 42999 2455
rect 42943 2403 42999 2405
rect 42943 2351 42945 2403
rect 42945 2351 42997 2403
rect 42997 2351 42999 2403
rect 42943 2349 42999 2351
rect 43583 2507 43639 2509
rect 43583 2455 43585 2507
rect 43585 2455 43637 2507
rect 43637 2455 43639 2507
rect 43583 2453 43639 2455
rect 43583 2403 43639 2405
rect 43583 2351 43585 2403
rect 43585 2351 43637 2403
rect 43637 2351 43639 2403
rect 43583 2349 43639 2351
rect 40997 1103 41053 1159
rect 41101 1103 41157 1159
rect 41205 1103 41261 1159
rect 40997 999 41053 1055
rect 41101 999 41157 1055
rect 41205 999 41261 1055
rect 40997 895 41053 951
rect 41101 895 41157 951
rect 41205 895 41261 951
rect 40997 43 41053 99
rect 41101 43 41157 99
rect 41205 43 41261 99
rect 40997 -61 41053 -5
rect 41101 -61 41157 -5
rect 41205 -61 41261 -5
rect 40997 -165 41053 -109
rect 41101 -165 41157 -109
rect 41205 -165 41261 -109
rect 40997 -623 41053 -567
rect 41101 -623 41157 -567
rect 41205 -623 41261 -567
rect 40997 -727 41053 -671
rect 41101 -727 41157 -671
rect 41205 -727 41261 -671
rect 40997 -831 41053 -775
rect 41101 -831 41157 -775
rect 41205 -831 41261 -775
rect 41356 2163 41412 2219
rect 41460 2163 41516 2219
rect 41564 2163 41620 2219
rect 41356 2059 41412 2115
rect 41460 2059 41516 2115
rect 41564 2059 41620 2115
rect 41356 1955 41412 2011
rect 41460 1955 41516 2011
rect 41564 1955 41620 2011
rect 42622 2113 42678 2115
rect 42622 2061 42624 2113
rect 42624 2061 42676 2113
rect 42676 2061 42678 2113
rect 42622 2059 42678 2061
rect 42622 2009 42678 2011
rect 42622 1957 42624 2009
rect 42624 1957 42676 2009
rect 42676 1957 42678 2009
rect 42622 1955 42678 1957
rect 43262 2113 43318 2115
rect 43262 2061 43264 2113
rect 43264 2061 43316 2113
rect 43316 2061 43318 2113
rect 43262 2059 43318 2061
rect 43262 2009 43318 2011
rect 43262 1957 43264 2009
rect 43264 1957 43316 2009
rect 43316 1957 43318 2009
rect 43262 1955 43318 1957
rect 41356 1497 41412 1553
rect 41460 1497 41516 1553
rect 41564 1497 41620 1553
rect 44223 2507 44279 2509
rect 44223 2455 44225 2507
rect 44225 2455 44277 2507
rect 44277 2455 44279 2507
rect 44223 2453 44279 2455
rect 44223 2403 44279 2405
rect 44223 2351 44225 2403
rect 44225 2351 44277 2403
rect 44277 2351 44279 2403
rect 44223 2349 44279 2351
rect 44863 2507 44919 2509
rect 44863 2455 44865 2507
rect 44865 2455 44917 2507
rect 44917 2455 44919 2507
rect 44863 2453 44919 2455
rect 44863 2403 44919 2405
rect 44863 2351 44865 2403
rect 44865 2351 44917 2403
rect 44917 2351 44919 2403
rect 44863 2349 44919 2351
rect 47077 2507 47133 2509
rect 47077 2455 47079 2507
rect 47079 2455 47131 2507
rect 47131 2455 47133 2507
rect 47077 2453 47133 2455
rect 47077 2403 47133 2405
rect 47077 2351 47079 2403
rect 47079 2351 47131 2403
rect 47131 2351 47133 2403
rect 47077 2349 47133 2351
rect 47717 2507 47773 2509
rect 47717 2455 47719 2507
rect 47719 2455 47771 2507
rect 47771 2455 47773 2507
rect 47717 2453 47773 2455
rect 47717 2403 47773 2405
rect 47717 2351 47719 2403
rect 47719 2351 47771 2403
rect 47771 2351 47773 2403
rect 47717 2349 47773 2351
rect 44542 2113 44598 2115
rect 44542 2061 44544 2113
rect 44544 2061 44596 2113
rect 44596 2061 44598 2113
rect 44542 2059 44598 2061
rect 44542 2009 44598 2011
rect 44542 1957 44544 2009
rect 44544 1957 44596 2009
rect 44596 1957 44598 2009
rect 44542 1955 44598 1957
rect 45182 2113 45238 2115
rect 45182 2061 45184 2113
rect 45184 2061 45236 2113
rect 45236 2061 45238 2113
rect 45182 2059 45238 2061
rect 45182 2009 45238 2011
rect 45182 1957 45184 2009
rect 45184 1957 45236 2009
rect 45236 1957 45238 2009
rect 45182 1955 45238 1957
rect 46758 2113 46814 2115
rect 46758 2061 46760 2113
rect 46760 2061 46812 2113
rect 46812 2061 46814 2113
rect 46758 2059 46814 2061
rect 46758 2009 46814 2011
rect 46758 1957 46760 2009
rect 46760 1957 46812 2009
rect 46812 1957 46814 2009
rect 46758 1955 46814 1957
rect 47398 2113 47454 2115
rect 47398 2061 47400 2113
rect 47400 2061 47452 2113
rect 47452 2061 47454 2113
rect 47398 2059 47454 2061
rect 47398 2009 47454 2011
rect 47398 1957 47400 2009
rect 47400 1957 47452 2009
rect 47452 1957 47454 2009
rect 47398 1955 47454 1957
rect 41356 1393 41412 1449
rect 41460 1393 41516 1449
rect 41564 1393 41620 1449
rect 41356 1289 41412 1345
rect 41460 1289 41516 1345
rect 41564 1289 41620 1345
rect 42943 1447 42999 1449
rect 42943 1395 42945 1447
rect 42945 1395 42997 1447
rect 42997 1395 42999 1447
rect 42943 1393 42999 1395
rect 42943 1343 42999 1345
rect 42943 1291 42945 1343
rect 42945 1291 42997 1343
rect 42997 1291 42999 1343
rect 42943 1289 42999 1291
rect 43583 1447 43639 1449
rect 43583 1395 43585 1447
rect 43585 1395 43637 1447
rect 43637 1395 43639 1447
rect 43583 1393 43639 1395
rect 43583 1343 43639 1345
rect 43583 1291 43585 1343
rect 43585 1291 43637 1343
rect 43637 1291 43639 1343
rect 43583 1289 43639 1291
rect 42622 1053 42678 1055
rect 42622 1001 42624 1053
rect 42624 1001 42676 1053
rect 42676 1001 42678 1053
rect 42622 999 42678 1001
rect 42622 949 42678 951
rect 42622 897 42624 949
rect 42624 897 42676 949
rect 42676 897 42678 949
rect 42622 895 42678 897
rect 43262 1053 43318 1055
rect 43262 1001 43264 1053
rect 43264 1001 43316 1053
rect 43316 1001 43318 1053
rect 43262 999 43318 1001
rect 43262 949 43318 951
rect 43262 897 43264 949
rect 43264 897 43316 949
rect 43316 897 43318 949
rect 43262 895 43318 897
rect 41356 437 41412 493
rect 41460 437 41516 493
rect 41564 437 41620 493
rect 50652 2557 50708 2613
rect 50756 2557 50812 2613
rect 50860 2557 50916 2613
rect 48357 2507 48413 2509
rect 48357 2455 48359 2507
rect 48359 2455 48411 2507
rect 48411 2455 48413 2507
rect 48357 2453 48413 2455
rect 48357 2403 48413 2405
rect 48357 2351 48359 2403
rect 48359 2351 48411 2403
rect 48411 2351 48413 2403
rect 48357 2349 48413 2351
rect 48997 2507 49053 2509
rect 48997 2455 48999 2507
rect 48999 2455 49051 2507
rect 49051 2455 49053 2507
rect 48997 2453 49053 2455
rect 48997 2403 49053 2405
rect 48997 2351 48999 2403
rect 48999 2351 49051 2403
rect 49051 2351 49053 2403
rect 48997 2349 49053 2351
rect 50652 2453 50708 2509
rect 50756 2453 50812 2509
rect 50860 2453 50916 2509
rect 50652 2349 50708 2405
rect 50756 2349 50812 2405
rect 50860 2349 50916 2405
rect 50312 2163 50368 2219
rect 50416 2163 50472 2219
rect 50520 2163 50576 2219
rect 48678 2113 48734 2115
rect 48678 2061 48680 2113
rect 48680 2061 48732 2113
rect 48732 2061 48734 2113
rect 48678 2059 48734 2061
rect 48678 2009 48734 2011
rect 48678 1957 48680 2009
rect 48680 1957 48732 2009
rect 48732 1957 48734 2009
rect 48678 1955 48734 1957
rect 49318 2113 49374 2115
rect 49318 2061 49320 2113
rect 49320 2061 49372 2113
rect 49372 2061 49374 2113
rect 49318 2059 49374 2061
rect 49318 2009 49374 2011
rect 49318 1957 49320 2009
rect 49320 1957 49372 2009
rect 49372 1957 49374 2009
rect 49318 1955 49374 1957
rect 50312 2059 50368 2115
rect 50416 2059 50472 2115
rect 50520 2059 50576 2115
rect 50312 1955 50368 2011
rect 50416 1955 50472 2011
rect 50520 1955 50576 2011
rect 44223 1447 44279 1449
rect 44223 1395 44225 1447
rect 44225 1395 44277 1447
rect 44277 1395 44279 1447
rect 44223 1393 44279 1395
rect 44223 1343 44279 1345
rect 44223 1291 44225 1343
rect 44225 1291 44277 1343
rect 44277 1291 44279 1343
rect 44223 1289 44279 1291
rect 44863 1447 44919 1449
rect 44863 1395 44865 1447
rect 44865 1395 44917 1447
rect 44917 1395 44919 1447
rect 44863 1393 44919 1395
rect 44863 1343 44919 1345
rect 44863 1291 44865 1343
rect 44865 1291 44917 1343
rect 44917 1291 44919 1343
rect 44863 1289 44919 1291
rect 47077 1447 47133 1449
rect 47077 1395 47079 1447
rect 47079 1395 47131 1447
rect 47131 1395 47133 1447
rect 47077 1393 47133 1395
rect 47077 1343 47133 1345
rect 47077 1291 47079 1343
rect 47079 1291 47131 1343
rect 47131 1291 47133 1343
rect 47077 1289 47133 1291
rect 47717 1447 47773 1449
rect 47717 1395 47719 1447
rect 47719 1395 47771 1447
rect 47771 1395 47773 1447
rect 47717 1393 47773 1395
rect 47717 1343 47773 1345
rect 47717 1291 47719 1343
rect 47719 1291 47771 1343
rect 47771 1291 47773 1343
rect 47717 1289 47773 1291
rect 44542 1053 44598 1055
rect 44542 1001 44544 1053
rect 44544 1001 44596 1053
rect 44596 1001 44598 1053
rect 44542 999 44598 1001
rect 44542 949 44598 951
rect 44542 897 44544 949
rect 44544 897 44596 949
rect 44596 897 44598 949
rect 44542 895 44598 897
rect 45182 1053 45238 1055
rect 45182 1001 45184 1053
rect 45184 1001 45236 1053
rect 45236 1001 45238 1053
rect 45182 999 45238 1001
rect 45182 949 45238 951
rect 45182 897 45184 949
rect 45184 897 45236 949
rect 45236 897 45238 949
rect 45182 895 45238 897
rect 46758 1053 46814 1055
rect 46758 1001 46760 1053
rect 46760 1001 46812 1053
rect 46812 1001 46814 1053
rect 46758 999 46814 1001
rect 46758 949 46814 951
rect 46758 897 46760 949
rect 46760 897 46812 949
rect 46812 897 46814 949
rect 46758 895 46814 897
rect 47398 1053 47454 1055
rect 47398 1001 47400 1053
rect 47400 1001 47452 1053
rect 47452 1001 47454 1053
rect 47398 999 47454 1001
rect 47398 949 47454 951
rect 47398 897 47400 949
rect 47400 897 47452 949
rect 47452 897 47454 949
rect 47398 895 47454 897
rect 41356 333 41412 389
rect 41460 333 41516 389
rect 41564 333 41620 389
rect 41356 229 41412 285
rect 41460 229 41516 285
rect 41564 229 41620 285
rect 40636 -1017 40692 -961
rect 40740 -1017 40796 -961
rect 40844 -1017 40900 -961
rect 34846 -1067 34902 -1065
rect 34846 -1119 34848 -1067
rect 34848 -1119 34900 -1067
rect 34900 -1119 34902 -1067
rect 34846 -1121 34902 -1119
rect 34846 -1171 34902 -1169
rect 34846 -1223 34848 -1171
rect 34848 -1223 34900 -1171
rect 34900 -1223 34902 -1171
rect 34846 -1225 34902 -1223
rect 35486 -1067 35542 -1065
rect 35486 -1119 35488 -1067
rect 35488 -1119 35540 -1067
rect 35540 -1119 35542 -1067
rect 35486 -1121 35542 -1119
rect 35486 -1171 35542 -1169
rect 35486 -1223 35488 -1171
rect 35488 -1223 35540 -1171
rect 35540 -1223 35542 -1171
rect 35486 -1225 35542 -1223
rect 37062 -1067 37118 -1065
rect 37062 -1119 37064 -1067
rect 37064 -1119 37116 -1067
rect 37116 -1119 37118 -1067
rect 37062 -1121 37118 -1119
rect 37062 -1171 37118 -1169
rect 37062 -1223 37064 -1171
rect 37064 -1223 37116 -1171
rect 37116 -1223 37118 -1171
rect 37062 -1225 37118 -1223
rect 37702 -1067 37758 -1065
rect 37702 -1119 37704 -1067
rect 37704 -1119 37756 -1067
rect 37756 -1119 37758 -1067
rect 37702 -1121 37758 -1119
rect 37702 -1171 37758 -1169
rect 37702 -1223 37704 -1171
rect 37704 -1223 37756 -1171
rect 37756 -1223 37758 -1171
rect 37702 -1225 37758 -1223
rect 38982 -1067 39038 -1065
rect 38982 -1119 38984 -1067
rect 38984 -1119 39036 -1067
rect 39036 -1119 39038 -1067
rect 38982 -1121 39038 -1119
rect 38982 -1171 39038 -1169
rect 38982 -1223 38984 -1171
rect 38984 -1223 39036 -1171
rect 39036 -1223 39038 -1171
rect 38982 -1225 39038 -1223
rect 39622 -1067 39678 -1065
rect 39622 -1119 39624 -1067
rect 39624 -1119 39676 -1067
rect 39676 -1119 39678 -1067
rect 39622 -1121 39678 -1119
rect 39622 -1171 39678 -1169
rect 39622 -1223 39624 -1171
rect 39624 -1223 39676 -1171
rect 39676 -1223 39678 -1171
rect 39622 -1225 39678 -1223
rect 40636 -1121 40692 -1065
rect 40740 -1121 40796 -1065
rect 40844 -1121 40900 -1065
rect 40636 -1225 40692 -1169
rect 40740 -1225 40796 -1169
rect 40844 -1225 40900 -1169
rect 42943 387 42999 389
rect 42943 335 42945 387
rect 42945 335 42997 387
rect 42997 335 42999 387
rect 42943 333 42999 335
rect 42943 283 42999 285
rect 42943 231 42945 283
rect 42945 231 42997 283
rect 42997 231 42999 283
rect 42943 229 42999 231
rect 43583 387 43639 389
rect 43583 335 43585 387
rect 43585 335 43637 387
rect 43637 335 43639 387
rect 43583 333 43639 335
rect 43583 283 43639 285
rect 43583 231 43585 283
rect 43585 231 43637 283
rect 43637 231 43639 283
rect 43583 229 43639 231
rect 42622 -7 42678 -5
rect 42622 -59 42624 -7
rect 42624 -59 42676 -7
rect 42676 -59 42678 -7
rect 42622 -61 42678 -59
rect 42622 -111 42678 -109
rect 42622 -163 42624 -111
rect 42624 -163 42676 -111
rect 42676 -163 42678 -111
rect 42622 -165 42678 -163
rect 43262 -7 43318 -5
rect 43262 -59 43264 -7
rect 43264 -59 43316 -7
rect 43316 -59 43318 -7
rect 43262 -61 43318 -59
rect 43262 -111 43318 -109
rect 43262 -163 43264 -111
rect 43264 -163 43316 -111
rect 43316 -163 43318 -111
rect 43262 -165 43318 -163
rect 50312 1497 50368 1553
rect 50416 1497 50472 1553
rect 50520 1497 50576 1553
rect 48357 1447 48413 1449
rect 48357 1395 48359 1447
rect 48359 1395 48411 1447
rect 48411 1395 48413 1447
rect 48357 1393 48413 1395
rect 48357 1343 48413 1345
rect 48357 1291 48359 1343
rect 48359 1291 48411 1343
rect 48411 1291 48413 1343
rect 48357 1289 48413 1291
rect 48997 1447 49053 1449
rect 48997 1395 48999 1447
rect 48999 1395 49051 1447
rect 49051 1395 49053 1447
rect 48997 1393 49053 1395
rect 48997 1343 49053 1345
rect 48997 1291 48999 1343
rect 48999 1291 49051 1343
rect 49051 1291 49053 1343
rect 48997 1289 49053 1291
rect 50312 1393 50368 1449
rect 50416 1393 50472 1449
rect 50520 1393 50576 1449
rect 50312 1289 50368 1345
rect 50416 1289 50472 1345
rect 50520 1289 50576 1345
rect 48678 1053 48734 1055
rect 48678 1001 48680 1053
rect 48680 1001 48732 1053
rect 48732 1001 48734 1053
rect 48678 999 48734 1001
rect 48678 949 48734 951
rect 48678 897 48680 949
rect 48680 897 48732 949
rect 48732 897 48734 949
rect 48678 895 48734 897
rect 49318 1053 49374 1055
rect 49318 1001 49320 1053
rect 49320 1001 49372 1053
rect 49372 1001 49374 1053
rect 49318 999 49374 1001
rect 49318 949 49374 951
rect 49318 897 49320 949
rect 49320 897 49372 949
rect 49372 897 49374 949
rect 49318 895 49374 897
rect 44223 387 44279 389
rect 44223 335 44225 387
rect 44225 335 44277 387
rect 44277 335 44279 387
rect 44223 333 44279 335
rect 44223 283 44279 285
rect 44223 231 44225 283
rect 44225 231 44277 283
rect 44277 231 44279 283
rect 44223 229 44279 231
rect 44863 387 44919 389
rect 44863 335 44865 387
rect 44865 335 44917 387
rect 44917 335 44919 387
rect 44863 333 44919 335
rect 44863 283 44919 285
rect 44863 231 44865 283
rect 44865 231 44917 283
rect 44917 231 44919 283
rect 44863 229 44919 231
rect 47077 387 47133 389
rect 47077 335 47079 387
rect 47079 335 47131 387
rect 47131 335 47133 387
rect 47077 333 47133 335
rect 47077 283 47133 285
rect 47077 231 47079 283
rect 47079 231 47131 283
rect 47131 231 47133 283
rect 47077 229 47133 231
rect 47717 387 47773 389
rect 47717 335 47719 387
rect 47719 335 47771 387
rect 47771 335 47773 387
rect 47717 333 47773 335
rect 47717 283 47773 285
rect 47717 231 47719 283
rect 47719 231 47771 283
rect 47771 231 47773 283
rect 47717 229 47773 231
rect 44542 -7 44598 -5
rect 44542 -59 44544 -7
rect 44544 -59 44596 -7
rect 44596 -59 44598 -7
rect 44542 -61 44598 -59
rect 44542 -111 44598 -109
rect 44542 -163 44544 -111
rect 44544 -163 44596 -111
rect 44596 -163 44598 -111
rect 44542 -165 44598 -163
rect 45182 -7 45238 -5
rect 45182 -59 45184 -7
rect 45184 -59 45236 -7
rect 45236 -59 45238 -7
rect 45182 -61 45238 -59
rect 45182 -111 45238 -109
rect 45182 -163 45184 -111
rect 45184 -163 45236 -111
rect 45236 -163 45238 -111
rect 45182 -165 45238 -163
rect 46758 -7 46814 -5
rect 46758 -59 46760 -7
rect 46760 -59 46812 -7
rect 46812 -59 46814 -7
rect 46758 -61 46814 -59
rect 46758 -111 46814 -109
rect 46758 -163 46760 -111
rect 46760 -163 46812 -111
rect 46812 -163 46814 -111
rect 46758 -165 46814 -163
rect 47398 -7 47454 -5
rect 47398 -59 47400 -7
rect 47400 -59 47452 -7
rect 47452 -59 47454 -7
rect 47398 -61 47454 -59
rect 47398 -111 47454 -109
rect 47398 -163 47400 -111
rect 47400 -163 47452 -111
rect 47452 -163 47454 -111
rect 47398 -165 47454 -163
rect 50312 437 50368 493
rect 50416 437 50472 493
rect 50520 437 50576 493
rect 48357 387 48413 389
rect 48357 335 48359 387
rect 48359 335 48411 387
rect 48411 335 48413 387
rect 48357 333 48413 335
rect 48357 283 48413 285
rect 48357 231 48359 283
rect 48359 231 48411 283
rect 48411 231 48413 283
rect 48357 229 48413 231
rect 48997 387 49053 389
rect 48997 335 48999 387
rect 48999 335 49051 387
rect 49051 335 49053 387
rect 48997 333 49053 335
rect 48997 283 49053 285
rect 48997 231 48999 283
rect 48999 231 49051 283
rect 49051 231 49053 283
rect 48997 229 49053 231
rect 50312 333 50368 389
rect 50416 333 50472 389
rect 50520 333 50576 389
rect 50312 229 50368 285
rect 50416 229 50472 285
rect 50520 229 50576 285
rect 48678 -7 48734 -5
rect 48678 -59 48680 -7
rect 48680 -59 48732 -7
rect 48732 -59 48734 -7
rect 48678 -61 48734 -59
rect 48678 -111 48734 -109
rect 48678 -163 48680 -111
rect 48680 -163 48732 -111
rect 48732 -163 48734 -111
rect 48678 -165 48734 -163
rect 49318 -7 49374 -5
rect 49318 -59 49320 -7
rect 49320 -59 49372 -7
rect 49372 -59 49374 -7
rect 49318 -61 49374 -59
rect 49318 -111 49374 -109
rect 49318 -163 49320 -111
rect 49320 -163 49372 -111
rect 49372 -163 49374 -111
rect 49318 -165 49374 -163
rect 42943 -673 42999 -671
rect 42943 -725 42945 -673
rect 42945 -725 42997 -673
rect 42997 -725 42999 -673
rect 42943 -727 42999 -725
rect 42943 -777 42999 -775
rect 42943 -829 42945 -777
rect 42945 -829 42997 -777
rect 42997 -829 42999 -777
rect 42943 -831 42999 -829
rect 43583 -673 43639 -671
rect 43583 -725 43585 -673
rect 43585 -725 43637 -673
rect 43637 -725 43639 -673
rect 43583 -727 43639 -725
rect 43583 -777 43639 -775
rect 43583 -829 43585 -777
rect 43585 -829 43637 -777
rect 43637 -829 43639 -777
rect 43583 -831 43639 -829
rect 44223 -673 44279 -671
rect 44223 -725 44225 -673
rect 44225 -725 44277 -673
rect 44277 -725 44279 -673
rect 44223 -727 44279 -725
rect 44223 -777 44279 -775
rect 44223 -829 44225 -777
rect 44225 -829 44277 -777
rect 44277 -829 44279 -777
rect 44223 -831 44279 -829
rect 44863 -673 44919 -671
rect 44863 -725 44865 -673
rect 44865 -725 44917 -673
rect 44917 -725 44919 -673
rect 44863 -727 44919 -725
rect 44863 -777 44919 -775
rect 44863 -829 44865 -777
rect 44865 -829 44917 -777
rect 44917 -829 44919 -777
rect 44863 -831 44919 -829
rect 47077 -673 47133 -671
rect 47077 -725 47079 -673
rect 47079 -725 47131 -673
rect 47131 -725 47133 -673
rect 47077 -727 47133 -725
rect 47077 -777 47133 -775
rect 47077 -829 47079 -777
rect 47079 -829 47131 -777
rect 47131 -829 47133 -777
rect 47077 -831 47133 -829
rect 47717 -673 47773 -671
rect 47717 -725 47719 -673
rect 47719 -725 47771 -673
rect 47771 -725 47773 -673
rect 47717 -727 47773 -725
rect 47717 -777 47773 -775
rect 47717 -829 47719 -777
rect 47719 -829 47771 -777
rect 47771 -829 47773 -777
rect 47717 -831 47773 -829
rect 48357 -673 48413 -671
rect 48357 -725 48359 -673
rect 48359 -725 48411 -673
rect 48411 -725 48413 -673
rect 48357 -727 48413 -725
rect 48357 -777 48413 -775
rect 48357 -829 48359 -777
rect 48359 -829 48411 -777
rect 48411 -829 48413 -777
rect 48357 -831 48413 -829
rect 48997 -673 49053 -671
rect 48997 -725 48999 -673
rect 48999 -725 49051 -673
rect 49051 -725 49053 -673
rect 48997 -727 49053 -725
rect 48997 -777 49053 -775
rect 48997 -829 48999 -777
rect 48999 -829 49051 -777
rect 49051 -829 49053 -777
rect 48997 -831 49053 -829
rect 41356 -1017 41412 -961
rect 41460 -1017 41516 -961
rect 41564 -1017 41620 -961
rect 52639 2507 52695 2509
rect 52639 2455 52641 2507
rect 52641 2455 52693 2507
rect 52693 2455 52695 2507
rect 52639 2453 52695 2455
rect 52639 2403 52695 2405
rect 52639 2351 52641 2403
rect 52641 2351 52693 2403
rect 52693 2351 52695 2403
rect 52639 2349 52695 2351
rect 53279 2507 53335 2509
rect 53279 2455 53281 2507
rect 53281 2455 53333 2507
rect 53333 2455 53335 2507
rect 53279 2453 53335 2455
rect 53279 2403 53335 2405
rect 53279 2351 53281 2403
rect 53281 2351 53333 2403
rect 53333 2351 53335 2403
rect 53279 2349 53335 2351
rect 50652 1103 50708 1159
rect 50756 1103 50812 1159
rect 50860 1103 50916 1159
rect 50652 999 50708 1055
rect 50756 999 50812 1055
rect 50860 999 50916 1055
rect 50652 895 50708 951
rect 50756 895 50812 951
rect 50860 895 50916 951
rect 50652 43 50708 99
rect 50756 43 50812 99
rect 50860 43 50916 99
rect 50652 -61 50708 -5
rect 50756 -61 50812 -5
rect 50860 -61 50916 -5
rect 50652 -165 50708 -109
rect 50756 -165 50812 -109
rect 50860 -165 50916 -109
rect 50652 -623 50708 -567
rect 50756 -623 50812 -567
rect 50860 -623 50916 -567
rect 50652 -727 50708 -671
rect 50756 -727 50812 -671
rect 50860 -727 50916 -671
rect 50652 -831 50708 -775
rect 50756 -831 50812 -775
rect 50860 -831 50916 -775
rect 51044 2163 51100 2219
rect 51148 2163 51204 2219
rect 51252 2163 51308 2219
rect 51044 2059 51100 2115
rect 51148 2059 51204 2115
rect 51252 2059 51308 2115
rect 51044 1955 51100 2011
rect 51148 1955 51204 2011
rect 51252 1955 51308 2011
rect 52318 2113 52374 2115
rect 52318 2061 52320 2113
rect 52320 2061 52372 2113
rect 52372 2061 52374 2113
rect 52318 2059 52374 2061
rect 52318 2009 52374 2011
rect 52318 1957 52320 2009
rect 52320 1957 52372 2009
rect 52372 1957 52374 2009
rect 52318 1955 52374 1957
rect 52958 2113 53014 2115
rect 52958 2061 52960 2113
rect 52960 2061 53012 2113
rect 53012 2061 53014 2113
rect 52958 2059 53014 2061
rect 52958 2009 53014 2011
rect 52958 1957 52960 2009
rect 52960 1957 53012 2009
rect 53012 1957 53014 2009
rect 52958 1955 53014 1957
rect 51044 1497 51100 1553
rect 51148 1497 51204 1553
rect 51252 1497 51308 1553
rect 53919 2507 53975 2509
rect 53919 2455 53921 2507
rect 53921 2455 53973 2507
rect 53973 2455 53975 2507
rect 53919 2453 53975 2455
rect 53919 2403 53975 2405
rect 53919 2351 53921 2403
rect 53921 2351 53973 2403
rect 53973 2351 53975 2403
rect 53919 2349 53975 2351
rect 54559 2507 54615 2509
rect 54559 2455 54561 2507
rect 54561 2455 54613 2507
rect 54613 2455 54615 2507
rect 54559 2453 54615 2455
rect 54559 2403 54615 2405
rect 54559 2351 54561 2403
rect 54561 2351 54613 2403
rect 54613 2351 54615 2403
rect 54559 2349 54615 2351
rect 56773 2507 56829 2509
rect 56773 2455 56775 2507
rect 56775 2455 56827 2507
rect 56827 2455 56829 2507
rect 56773 2453 56829 2455
rect 56773 2403 56829 2405
rect 56773 2351 56775 2403
rect 56775 2351 56827 2403
rect 56827 2351 56829 2403
rect 56773 2349 56829 2351
rect 57413 2507 57469 2509
rect 57413 2455 57415 2507
rect 57415 2455 57467 2507
rect 57467 2455 57469 2507
rect 57413 2453 57469 2455
rect 57413 2403 57469 2405
rect 57413 2351 57415 2403
rect 57415 2351 57467 2403
rect 57467 2351 57469 2403
rect 57413 2349 57469 2351
rect 54238 2113 54294 2115
rect 54238 2061 54240 2113
rect 54240 2061 54292 2113
rect 54292 2061 54294 2113
rect 54238 2059 54294 2061
rect 54238 2009 54294 2011
rect 54238 1957 54240 2009
rect 54240 1957 54292 2009
rect 54292 1957 54294 2009
rect 54238 1955 54294 1957
rect 54878 2113 54934 2115
rect 54878 2061 54880 2113
rect 54880 2061 54932 2113
rect 54932 2061 54934 2113
rect 54878 2059 54934 2061
rect 54878 2009 54934 2011
rect 54878 1957 54880 2009
rect 54880 1957 54932 2009
rect 54932 1957 54934 2009
rect 54878 1955 54934 1957
rect 56454 2113 56510 2115
rect 56454 2061 56456 2113
rect 56456 2061 56508 2113
rect 56508 2061 56510 2113
rect 56454 2059 56510 2061
rect 56454 2009 56510 2011
rect 56454 1957 56456 2009
rect 56456 1957 56508 2009
rect 56508 1957 56510 2009
rect 56454 1955 56510 1957
rect 57094 2113 57150 2115
rect 57094 2061 57096 2113
rect 57096 2061 57148 2113
rect 57148 2061 57150 2113
rect 57094 2059 57150 2061
rect 57094 2009 57150 2011
rect 57094 1957 57096 2009
rect 57096 1957 57148 2009
rect 57148 1957 57150 2009
rect 57094 1955 57150 1957
rect 51044 1393 51100 1449
rect 51148 1393 51204 1449
rect 51252 1393 51308 1449
rect 51044 1289 51100 1345
rect 51148 1289 51204 1345
rect 51252 1289 51308 1345
rect 52639 1447 52695 1449
rect 52639 1395 52641 1447
rect 52641 1395 52693 1447
rect 52693 1395 52695 1447
rect 52639 1393 52695 1395
rect 52639 1343 52695 1345
rect 52639 1291 52641 1343
rect 52641 1291 52693 1343
rect 52693 1291 52695 1343
rect 52639 1289 52695 1291
rect 53279 1447 53335 1449
rect 53279 1395 53281 1447
rect 53281 1395 53333 1447
rect 53333 1395 53335 1447
rect 53279 1393 53335 1395
rect 53279 1343 53335 1345
rect 53279 1291 53281 1343
rect 53281 1291 53333 1343
rect 53333 1291 53335 1343
rect 53279 1289 53335 1291
rect 52318 1053 52374 1055
rect 52318 1001 52320 1053
rect 52320 1001 52372 1053
rect 52372 1001 52374 1053
rect 52318 999 52374 1001
rect 52318 949 52374 951
rect 52318 897 52320 949
rect 52320 897 52372 949
rect 52372 897 52374 949
rect 52318 895 52374 897
rect 52958 1053 53014 1055
rect 52958 1001 52960 1053
rect 52960 1001 53012 1053
rect 53012 1001 53014 1053
rect 52958 999 53014 1001
rect 52958 949 53014 951
rect 52958 897 52960 949
rect 52960 897 53012 949
rect 53012 897 53014 949
rect 52958 895 53014 897
rect 51044 437 51100 493
rect 51148 437 51204 493
rect 51252 437 51308 493
rect 60433 2557 60489 2613
rect 60537 2557 60593 2613
rect 60641 2557 60697 2613
rect 58053 2507 58109 2509
rect 58053 2455 58055 2507
rect 58055 2455 58107 2507
rect 58107 2455 58109 2507
rect 58053 2453 58109 2455
rect 58053 2403 58109 2405
rect 58053 2351 58055 2403
rect 58055 2351 58107 2403
rect 58107 2351 58109 2403
rect 58053 2349 58109 2351
rect 58693 2507 58749 2509
rect 58693 2455 58695 2507
rect 58695 2455 58747 2507
rect 58747 2455 58749 2507
rect 58693 2453 58749 2455
rect 58693 2403 58749 2405
rect 58693 2351 58695 2403
rect 58695 2351 58747 2403
rect 58747 2351 58749 2403
rect 58693 2349 58749 2351
rect 60433 2453 60489 2509
rect 60537 2453 60593 2509
rect 60641 2453 60697 2509
rect 60433 2349 60489 2405
rect 60537 2349 60593 2405
rect 60641 2349 60697 2405
rect 60028 2163 60084 2219
rect 60132 2163 60188 2219
rect 60236 2163 60292 2219
rect 58374 2113 58430 2115
rect 58374 2061 58376 2113
rect 58376 2061 58428 2113
rect 58428 2061 58430 2113
rect 58374 2059 58430 2061
rect 58374 2009 58430 2011
rect 58374 1957 58376 2009
rect 58376 1957 58428 2009
rect 58428 1957 58430 2009
rect 58374 1955 58430 1957
rect 59014 2113 59070 2115
rect 59014 2061 59016 2113
rect 59016 2061 59068 2113
rect 59068 2061 59070 2113
rect 59014 2059 59070 2061
rect 59014 2009 59070 2011
rect 59014 1957 59016 2009
rect 59016 1957 59068 2009
rect 59068 1957 59070 2009
rect 59014 1955 59070 1957
rect 60028 2059 60084 2115
rect 60132 2059 60188 2115
rect 60236 2059 60292 2115
rect 60028 1955 60084 2011
rect 60132 1955 60188 2011
rect 60236 1955 60292 2011
rect 53919 1447 53975 1449
rect 53919 1395 53921 1447
rect 53921 1395 53973 1447
rect 53973 1395 53975 1447
rect 53919 1393 53975 1395
rect 53919 1343 53975 1345
rect 53919 1291 53921 1343
rect 53921 1291 53973 1343
rect 53973 1291 53975 1343
rect 53919 1289 53975 1291
rect 54559 1447 54615 1449
rect 54559 1395 54561 1447
rect 54561 1395 54613 1447
rect 54613 1395 54615 1447
rect 54559 1393 54615 1395
rect 54559 1343 54615 1345
rect 54559 1291 54561 1343
rect 54561 1291 54613 1343
rect 54613 1291 54615 1343
rect 54559 1289 54615 1291
rect 56773 1447 56829 1449
rect 56773 1395 56775 1447
rect 56775 1395 56827 1447
rect 56827 1395 56829 1447
rect 56773 1393 56829 1395
rect 56773 1343 56829 1345
rect 56773 1291 56775 1343
rect 56775 1291 56827 1343
rect 56827 1291 56829 1343
rect 56773 1289 56829 1291
rect 57413 1447 57469 1449
rect 57413 1395 57415 1447
rect 57415 1395 57467 1447
rect 57467 1395 57469 1447
rect 57413 1393 57469 1395
rect 57413 1343 57469 1345
rect 57413 1291 57415 1343
rect 57415 1291 57467 1343
rect 57467 1291 57469 1343
rect 57413 1289 57469 1291
rect 54238 1053 54294 1055
rect 54238 1001 54240 1053
rect 54240 1001 54292 1053
rect 54292 1001 54294 1053
rect 54238 999 54294 1001
rect 54238 949 54294 951
rect 54238 897 54240 949
rect 54240 897 54292 949
rect 54292 897 54294 949
rect 54238 895 54294 897
rect 54878 1053 54934 1055
rect 54878 1001 54880 1053
rect 54880 1001 54932 1053
rect 54932 1001 54934 1053
rect 54878 999 54934 1001
rect 54878 949 54934 951
rect 54878 897 54880 949
rect 54880 897 54932 949
rect 54932 897 54934 949
rect 54878 895 54934 897
rect 56454 1053 56510 1055
rect 56454 1001 56456 1053
rect 56456 1001 56508 1053
rect 56508 1001 56510 1053
rect 56454 999 56510 1001
rect 56454 949 56510 951
rect 56454 897 56456 949
rect 56456 897 56508 949
rect 56508 897 56510 949
rect 56454 895 56510 897
rect 57094 1053 57150 1055
rect 57094 1001 57096 1053
rect 57096 1001 57148 1053
rect 57148 1001 57150 1053
rect 57094 999 57150 1001
rect 57094 949 57150 951
rect 57094 897 57096 949
rect 57096 897 57148 949
rect 57148 897 57150 949
rect 57094 895 57150 897
rect 51044 333 51100 389
rect 51148 333 51204 389
rect 51252 333 51308 389
rect 51044 229 51100 285
rect 51148 229 51204 285
rect 51252 229 51308 285
rect 50312 -1017 50368 -961
rect 50416 -1017 50472 -961
rect 50520 -1017 50576 -961
rect 41356 -1121 41412 -1065
rect 41460 -1121 41516 -1065
rect 41564 -1121 41620 -1065
rect 41356 -1225 41412 -1169
rect 41460 -1225 41516 -1169
rect 41564 -1225 41620 -1169
rect 42622 -1067 42678 -1065
rect 42622 -1119 42624 -1067
rect 42624 -1119 42676 -1067
rect 42676 -1119 42678 -1067
rect 42622 -1121 42678 -1119
rect 42622 -1171 42678 -1169
rect 42622 -1223 42624 -1171
rect 42624 -1223 42676 -1171
rect 42676 -1223 42678 -1171
rect 42622 -1225 42678 -1223
rect 43262 -1067 43318 -1065
rect 43262 -1119 43264 -1067
rect 43264 -1119 43316 -1067
rect 43316 -1119 43318 -1067
rect 43262 -1121 43318 -1119
rect 43262 -1171 43318 -1169
rect 43262 -1223 43264 -1171
rect 43264 -1223 43316 -1171
rect 43316 -1223 43318 -1171
rect 43262 -1225 43318 -1223
rect 44542 -1067 44598 -1065
rect 44542 -1119 44544 -1067
rect 44544 -1119 44596 -1067
rect 44596 -1119 44598 -1067
rect 44542 -1121 44598 -1119
rect 44542 -1171 44598 -1169
rect 44542 -1223 44544 -1171
rect 44544 -1223 44596 -1171
rect 44596 -1223 44598 -1171
rect 44542 -1225 44598 -1223
rect 45182 -1067 45238 -1065
rect 45182 -1119 45184 -1067
rect 45184 -1119 45236 -1067
rect 45236 -1119 45238 -1067
rect 45182 -1121 45238 -1119
rect 45182 -1171 45238 -1169
rect 45182 -1223 45184 -1171
rect 45184 -1223 45236 -1171
rect 45236 -1223 45238 -1171
rect 45182 -1225 45238 -1223
rect 46758 -1067 46814 -1065
rect 46758 -1119 46760 -1067
rect 46760 -1119 46812 -1067
rect 46812 -1119 46814 -1067
rect 46758 -1121 46814 -1119
rect 46758 -1171 46814 -1169
rect 46758 -1223 46760 -1171
rect 46760 -1223 46812 -1171
rect 46812 -1223 46814 -1171
rect 46758 -1225 46814 -1223
rect 47398 -1067 47454 -1065
rect 47398 -1119 47400 -1067
rect 47400 -1119 47452 -1067
rect 47452 -1119 47454 -1067
rect 47398 -1121 47454 -1119
rect 47398 -1171 47454 -1169
rect 47398 -1223 47400 -1171
rect 47400 -1223 47452 -1171
rect 47452 -1223 47454 -1171
rect 47398 -1225 47454 -1223
rect 48678 -1067 48734 -1065
rect 48678 -1119 48680 -1067
rect 48680 -1119 48732 -1067
rect 48732 -1119 48734 -1067
rect 48678 -1121 48734 -1119
rect 48678 -1171 48734 -1169
rect 48678 -1223 48680 -1171
rect 48680 -1223 48732 -1171
rect 48732 -1223 48734 -1171
rect 48678 -1225 48734 -1223
rect 49318 -1067 49374 -1065
rect 49318 -1119 49320 -1067
rect 49320 -1119 49372 -1067
rect 49372 -1119 49374 -1067
rect 49318 -1121 49374 -1119
rect 49318 -1171 49374 -1169
rect 49318 -1223 49320 -1171
rect 49320 -1223 49372 -1171
rect 49372 -1223 49374 -1171
rect 49318 -1225 49374 -1223
rect 50312 -1121 50368 -1065
rect 50416 -1121 50472 -1065
rect 50520 -1121 50576 -1065
rect 50312 -1225 50368 -1169
rect 50416 -1225 50472 -1169
rect 50520 -1225 50576 -1169
rect 52639 387 52695 389
rect 52639 335 52641 387
rect 52641 335 52693 387
rect 52693 335 52695 387
rect 52639 333 52695 335
rect 52639 283 52695 285
rect 52639 231 52641 283
rect 52641 231 52693 283
rect 52693 231 52695 283
rect 52639 229 52695 231
rect 53279 387 53335 389
rect 53279 335 53281 387
rect 53281 335 53333 387
rect 53333 335 53335 387
rect 53279 333 53335 335
rect 53279 283 53335 285
rect 53279 231 53281 283
rect 53281 231 53333 283
rect 53333 231 53335 283
rect 53279 229 53335 231
rect 52318 -7 52374 -5
rect 52318 -59 52320 -7
rect 52320 -59 52372 -7
rect 52372 -59 52374 -7
rect 52318 -61 52374 -59
rect 52318 -111 52374 -109
rect 52318 -163 52320 -111
rect 52320 -163 52372 -111
rect 52372 -163 52374 -111
rect 52318 -165 52374 -163
rect 52958 -7 53014 -5
rect 52958 -59 52960 -7
rect 52960 -59 53012 -7
rect 53012 -59 53014 -7
rect 52958 -61 53014 -59
rect 52958 -111 53014 -109
rect 52958 -163 52960 -111
rect 52960 -163 53012 -111
rect 53012 -163 53014 -111
rect 52958 -165 53014 -163
rect 60028 1497 60084 1553
rect 60132 1497 60188 1553
rect 60236 1497 60292 1553
rect 58053 1447 58109 1449
rect 58053 1395 58055 1447
rect 58055 1395 58107 1447
rect 58107 1395 58109 1447
rect 58053 1393 58109 1395
rect 58053 1343 58109 1345
rect 58053 1291 58055 1343
rect 58055 1291 58107 1343
rect 58107 1291 58109 1343
rect 58053 1289 58109 1291
rect 58693 1447 58749 1449
rect 58693 1395 58695 1447
rect 58695 1395 58747 1447
rect 58747 1395 58749 1447
rect 58693 1393 58749 1395
rect 58693 1343 58749 1345
rect 58693 1291 58695 1343
rect 58695 1291 58747 1343
rect 58747 1291 58749 1343
rect 58693 1289 58749 1291
rect 60028 1393 60084 1449
rect 60132 1393 60188 1449
rect 60236 1393 60292 1449
rect 60028 1289 60084 1345
rect 60132 1289 60188 1345
rect 60236 1289 60292 1345
rect 58374 1053 58430 1055
rect 58374 1001 58376 1053
rect 58376 1001 58428 1053
rect 58428 1001 58430 1053
rect 58374 999 58430 1001
rect 58374 949 58430 951
rect 58374 897 58376 949
rect 58376 897 58428 949
rect 58428 897 58430 949
rect 58374 895 58430 897
rect 59014 1053 59070 1055
rect 59014 1001 59016 1053
rect 59016 1001 59068 1053
rect 59068 1001 59070 1053
rect 59014 999 59070 1001
rect 59014 949 59070 951
rect 59014 897 59016 949
rect 59016 897 59068 949
rect 59068 897 59070 949
rect 59014 895 59070 897
rect 53919 387 53975 389
rect 53919 335 53921 387
rect 53921 335 53973 387
rect 53973 335 53975 387
rect 53919 333 53975 335
rect 53919 283 53975 285
rect 53919 231 53921 283
rect 53921 231 53973 283
rect 53973 231 53975 283
rect 53919 229 53975 231
rect 54559 387 54615 389
rect 54559 335 54561 387
rect 54561 335 54613 387
rect 54613 335 54615 387
rect 54559 333 54615 335
rect 54559 283 54615 285
rect 54559 231 54561 283
rect 54561 231 54613 283
rect 54613 231 54615 283
rect 54559 229 54615 231
rect 56773 387 56829 389
rect 56773 335 56775 387
rect 56775 335 56827 387
rect 56827 335 56829 387
rect 56773 333 56829 335
rect 56773 283 56829 285
rect 56773 231 56775 283
rect 56775 231 56827 283
rect 56827 231 56829 283
rect 56773 229 56829 231
rect 57413 387 57469 389
rect 57413 335 57415 387
rect 57415 335 57467 387
rect 57467 335 57469 387
rect 57413 333 57469 335
rect 57413 283 57469 285
rect 57413 231 57415 283
rect 57415 231 57467 283
rect 57467 231 57469 283
rect 57413 229 57469 231
rect 54238 -7 54294 -5
rect 54238 -59 54240 -7
rect 54240 -59 54292 -7
rect 54292 -59 54294 -7
rect 54238 -61 54294 -59
rect 54238 -111 54294 -109
rect 54238 -163 54240 -111
rect 54240 -163 54292 -111
rect 54292 -163 54294 -111
rect 54238 -165 54294 -163
rect 54878 -7 54934 -5
rect 54878 -59 54880 -7
rect 54880 -59 54932 -7
rect 54932 -59 54934 -7
rect 54878 -61 54934 -59
rect 54878 -111 54934 -109
rect 54878 -163 54880 -111
rect 54880 -163 54932 -111
rect 54932 -163 54934 -111
rect 54878 -165 54934 -163
rect 56454 -7 56510 -5
rect 56454 -59 56456 -7
rect 56456 -59 56508 -7
rect 56508 -59 56510 -7
rect 56454 -61 56510 -59
rect 56454 -111 56510 -109
rect 56454 -163 56456 -111
rect 56456 -163 56508 -111
rect 56508 -163 56510 -111
rect 56454 -165 56510 -163
rect 57094 -7 57150 -5
rect 57094 -59 57096 -7
rect 57096 -59 57148 -7
rect 57148 -59 57150 -7
rect 57094 -61 57150 -59
rect 57094 -111 57150 -109
rect 57094 -163 57096 -111
rect 57096 -163 57148 -111
rect 57148 -163 57150 -111
rect 57094 -165 57150 -163
rect 60028 437 60084 493
rect 60132 437 60188 493
rect 60236 437 60292 493
rect 58053 387 58109 389
rect 58053 335 58055 387
rect 58055 335 58107 387
rect 58107 335 58109 387
rect 58053 333 58109 335
rect 58053 283 58109 285
rect 58053 231 58055 283
rect 58055 231 58107 283
rect 58107 231 58109 283
rect 58053 229 58109 231
rect 58693 387 58749 389
rect 58693 335 58695 387
rect 58695 335 58747 387
rect 58747 335 58749 387
rect 58693 333 58749 335
rect 58693 283 58749 285
rect 58693 231 58695 283
rect 58695 231 58747 283
rect 58747 231 58749 283
rect 58693 229 58749 231
rect 60028 333 60084 389
rect 60132 333 60188 389
rect 60236 333 60292 389
rect 60028 229 60084 285
rect 60132 229 60188 285
rect 60236 229 60292 285
rect 58374 -7 58430 -5
rect 58374 -59 58376 -7
rect 58376 -59 58428 -7
rect 58428 -59 58430 -7
rect 58374 -61 58430 -59
rect 58374 -111 58430 -109
rect 58374 -163 58376 -111
rect 58376 -163 58428 -111
rect 58428 -163 58430 -111
rect 58374 -165 58430 -163
rect 59014 -7 59070 -5
rect 59014 -59 59016 -7
rect 59016 -59 59068 -7
rect 59068 -59 59070 -7
rect 59014 -61 59070 -59
rect 59014 -111 59070 -109
rect 59014 -163 59016 -111
rect 59016 -163 59068 -111
rect 59068 -163 59070 -111
rect 59014 -165 59070 -163
rect 52639 -673 52695 -671
rect 52639 -725 52641 -673
rect 52641 -725 52693 -673
rect 52693 -725 52695 -673
rect 52639 -727 52695 -725
rect 52639 -777 52695 -775
rect 52639 -829 52641 -777
rect 52641 -829 52693 -777
rect 52693 -829 52695 -777
rect 52639 -831 52695 -829
rect 53279 -673 53335 -671
rect 53279 -725 53281 -673
rect 53281 -725 53333 -673
rect 53333 -725 53335 -673
rect 53279 -727 53335 -725
rect 53279 -777 53335 -775
rect 53279 -829 53281 -777
rect 53281 -829 53333 -777
rect 53333 -829 53335 -777
rect 53279 -831 53335 -829
rect 53919 -673 53975 -671
rect 53919 -725 53921 -673
rect 53921 -725 53973 -673
rect 53973 -725 53975 -673
rect 53919 -727 53975 -725
rect 53919 -777 53975 -775
rect 53919 -829 53921 -777
rect 53921 -829 53973 -777
rect 53973 -829 53975 -777
rect 53919 -831 53975 -829
rect 54559 -673 54615 -671
rect 54559 -725 54561 -673
rect 54561 -725 54613 -673
rect 54613 -725 54615 -673
rect 54559 -727 54615 -725
rect 54559 -777 54615 -775
rect 54559 -829 54561 -777
rect 54561 -829 54613 -777
rect 54613 -829 54615 -777
rect 54559 -831 54615 -829
rect 56773 -673 56829 -671
rect 56773 -725 56775 -673
rect 56775 -725 56827 -673
rect 56827 -725 56829 -673
rect 56773 -727 56829 -725
rect 56773 -777 56829 -775
rect 56773 -829 56775 -777
rect 56775 -829 56827 -777
rect 56827 -829 56829 -777
rect 56773 -831 56829 -829
rect 57413 -673 57469 -671
rect 57413 -725 57415 -673
rect 57415 -725 57467 -673
rect 57467 -725 57469 -673
rect 57413 -727 57469 -725
rect 57413 -777 57469 -775
rect 57413 -829 57415 -777
rect 57415 -829 57467 -777
rect 57467 -829 57469 -777
rect 57413 -831 57469 -829
rect 58053 -673 58109 -671
rect 58053 -725 58055 -673
rect 58055 -725 58107 -673
rect 58107 -725 58109 -673
rect 58053 -727 58109 -725
rect 58053 -777 58109 -775
rect 58053 -829 58055 -777
rect 58055 -829 58107 -777
rect 58107 -829 58109 -777
rect 58053 -831 58109 -829
rect 58693 -673 58749 -671
rect 58693 -725 58695 -673
rect 58695 -725 58747 -673
rect 58747 -725 58749 -673
rect 58693 -727 58749 -725
rect 58693 -777 58749 -775
rect 58693 -829 58695 -777
rect 58695 -829 58747 -777
rect 58747 -829 58749 -777
rect 58693 -831 58749 -829
rect 51044 -1017 51100 -961
rect 51148 -1017 51204 -961
rect 51252 -1017 51308 -961
rect 62335 2507 62391 2509
rect 62335 2455 62337 2507
rect 62337 2455 62389 2507
rect 62389 2455 62391 2507
rect 62335 2453 62391 2455
rect 62335 2403 62391 2405
rect 62335 2351 62337 2403
rect 62337 2351 62389 2403
rect 62389 2351 62391 2403
rect 62335 2349 62391 2351
rect 62975 2507 63031 2509
rect 62975 2455 62977 2507
rect 62977 2455 63029 2507
rect 63029 2455 63031 2507
rect 62975 2453 63031 2455
rect 62975 2403 63031 2405
rect 62975 2351 62977 2403
rect 62977 2351 63029 2403
rect 63029 2351 63031 2403
rect 62975 2349 63031 2351
rect 60433 1103 60489 1159
rect 60537 1103 60593 1159
rect 60641 1103 60697 1159
rect 60433 999 60489 1055
rect 60537 999 60593 1055
rect 60641 999 60697 1055
rect 60433 895 60489 951
rect 60537 895 60593 951
rect 60641 895 60697 951
rect 60433 43 60489 99
rect 60537 43 60593 99
rect 60641 43 60697 99
rect 60433 -61 60489 -5
rect 60537 -61 60593 -5
rect 60641 -61 60697 -5
rect 60433 -165 60489 -109
rect 60537 -165 60593 -109
rect 60641 -165 60697 -109
rect 60433 -623 60489 -567
rect 60537 -623 60593 -567
rect 60641 -623 60697 -567
rect 60433 -727 60489 -671
rect 60537 -727 60593 -671
rect 60641 -727 60697 -671
rect 60433 -831 60489 -775
rect 60537 -831 60593 -775
rect 60641 -831 60697 -775
rect 60792 2163 60848 2219
rect 60896 2163 60952 2219
rect 61000 2163 61056 2219
rect 60792 2059 60848 2115
rect 60896 2059 60952 2115
rect 61000 2059 61056 2115
rect 60792 1955 60848 2011
rect 60896 1955 60952 2011
rect 61000 1955 61056 2011
rect 62014 2113 62070 2115
rect 62014 2061 62016 2113
rect 62016 2061 62068 2113
rect 62068 2061 62070 2113
rect 62014 2059 62070 2061
rect 62014 2009 62070 2011
rect 62014 1957 62016 2009
rect 62016 1957 62068 2009
rect 62068 1957 62070 2009
rect 62014 1955 62070 1957
rect 62654 2113 62710 2115
rect 62654 2061 62656 2113
rect 62656 2061 62708 2113
rect 62708 2061 62710 2113
rect 62654 2059 62710 2061
rect 62654 2009 62710 2011
rect 62654 1957 62656 2009
rect 62656 1957 62708 2009
rect 62708 1957 62710 2009
rect 62654 1955 62710 1957
rect 60792 1497 60848 1553
rect 60896 1497 60952 1553
rect 61000 1497 61056 1553
rect 63615 2507 63671 2509
rect 63615 2455 63617 2507
rect 63617 2455 63669 2507
rect 63669 2455 63671 2507
rect 63615 2453 63671 2455
rect 63615 2403 63671 2405
rect 63615 2351 63617 2403
rect 63617 2351 63669 2403
rect 63669 2351 63671 2403
rect 63615 2349 63671 2351
rect 64255 2507 64311 2509
rect 64255 2455 64257 2507
rect 64257 2455 64309 2507
rect 64309 2455 64311 2507
rect 64255 2453 64311 2455
rect 64255 2403 64311 2405
rect 64255 2351 64257 2403
rect 64257 2351 64309 2403
rect 64309 2351 64311 2403
rect 64255 2349 64311 2351
rect 63934 2113 63990 2115
rect 63934 2061 63936 2113
rect 63936 2061 63988 2113
rect 63988 2061 63990 2113
rect 63934 2059 63990 2061
rect 63934 2009 63990 2011
rect 63934 1957 63936 2009
rect 63936 1957 63988 2009
rect 63988 1957 63990 2009
rect 63934 1955 63990 1957
rect 64574 2113 64630 2115
rect 64574 2061 64576 2113
rect 64576 2061 64628 2113
rect 64628 2061 64630 2113
rect 64574 2059 64630 2061
rect 64574 2009 64630 2011
rect 64574 1957 64576 2009
rect 64576 1957 64628 2009
rect 64628 1957 64630 2009
rect 64574 1955 64630 1957
rect 60792 1393 60848 1449
rect 60896 1393 60952 1449
rect 61000 1393 61056 1449
rect 60792 1289 60848 1345
rect 60896 1289 60952 1345
rect 61000 1289 61056 1345
rect 62335 1447 62391 1449
rect 62335 1395 62337 1447
rect 62337 1395 62389 1447
rect 62389 1395 62391 1447
rect 62335 1393 62391 1395
rect 62335 1343 62391 1345
rect 62335 1291 62337 1343
rect 62337 1291 62389 1343
rect 62389 1291 62391 1343
rect 62335 1289 62391 1291
rect 62975 1447 63031 1449
rect 62975 1395 62977 1447
rect 62977 1395 63029 1447
rect 63029 1395 63031 1447
rect 62975 1393 63031 1395
rect 62975 1343 63031 1345
rect 62975 1291 62977 1343
rect 62977 1291 63029 1343
rect 63029 1291 63031 1343
rect 62975 1289 63031 1291
rect 62014 1053 62070 1055
rect 62014 1001 62016 1053
rect 62016 1001 62068 1053
rect 62068 1001 62070 1053
rect 62014 999 62070 1001
rect 62014 949 62070 951
rect 62014 897 62016 949
rect 62016 897 62068 949
rect 62068 897 62070 949
rect 62014 895 62070 897
rect 62654 1053 62710 1055
rect 62654 1001 62656 1053
rect 62656 1001 62708 1053
rect 62708 1001 62710 1053
rect 62654 999 62710 1001
rect 62654 949 62710 951
rect 62654 897 62656 949
rect 62656 897 62708 949
rect 62708 897 62710 949
rect 62654 895 62710 897
rect 60792 437 60848 493
rect 60896 437 60952 493
rect 61000 437 61056 493
rect 63615 1447 63671 1449
rect 63615 1395 63617 1447
rect 63617 1395 63669 1447
rect 63669 1395 63671 1447
rect 63615 1393 63671 1395
rect 63615 1343 63671 1345
rect 63615 1291 63617 1343
rect 63617 1291 63669 1343
rect 63669 1291 63671 1343
rect 63615 1289 63671 1291
rect 64255 1447 64311 1449
rect 64255 1395 64257 1447
rect 64257 1395 64309 1447
rect 64309 1395 64311 1447
rect 64255 1393 64311 1395
rect 64255 1343 64311 1345
rect 64255 1291 64257 1343
rect 64257 1291 64309 1343
rect 64309 1291 64311 1343
rect 64255 1289 64311 1291
rect 63934 1053 63990 1055
rect 63934 1001 63936 1053
rect 63936 1001 63988 1053
rect 63988 1001 63990 1053
rect 63934 999 63990 1001
rect 63934 949 63990 951
rect 63934 897 63936 949
rect 63936 897 63988 949
rect 63988 897 63990 949
rect 63934 895 63990 897
rect 64574 1053 64630 1055
rect 64574 1001 64576 1053
rect 64576 1001 64628 1053
rect 64628 1001 64630 1053
rect 64574 999 64630 1001
rect 64574 949 64630 951
rect 64574 897 64576 949
rect 64576 897 64628 949
rect 64628 897 64630 949
rect 64574 895 64630 897
rect 60792 333 60848 389
rect 60896 333 60952 389
rect 61000 333 61056 389
rect 60792 229 60848 285
rect 60896 229 60952 285
rect 61000 229 61056 285
rect 60028 -1017 60084 -961
rect 60132 -1017 60188 -961
rect 60236 -1017 60292 -961
rect 51044 -1121 51100 -1065
rect 51148 -1121 51204 -1065
rect 51252 -1121 51308 -1065
rect 51044 -1225 51100 -1169
rect 51148 -1225 51204 -1169
rect 51252 -1225 51308 -1169
rect 52318 -1067 52374 -1065
rect 52318 -1119 52320 -1067
rect 52320 -1119 52372 -1067
rect 52372 -1119 52374 -1067
rect 52318 -1121 52374 -1119
rect 52318 -1171 52374 -1169
rect 52318 -1223 52320 -1171
rect 52320 -1223 52372 -1171
rect 52372 -1223 52374 -1171
rect 52318 -1225 52374 -1223
rect 52958 -1067 53014 -1065
rect 52958 -1119 52960 -1067
rect 52960 -1119 53012 -1067
rect 53012 -1119 53014 -1067
rect 52958 -1121 53014 -1119
rect 52958 -1171 53014 -1169
rect 52958 -1223 52960 -1171
rect 52960 -1223 53012 -1171
rect 53012 -1223 53014 -1171
rect 52958 -1225 53014 -1223
rect 54238 -1067 54294 -1065
rect 54238 -1119 54240 -1067
rect 54240 -1119 54292 -1067
rect 54292 -1119 54294 -1067
rect 54238 -1121 54294 -1119
rect 54238 -1171 54294 -1169
rect 54238 -1223 54240 -1171
rect 54240 -1223 54292 -1171
rect 54292 -1223 54294 -1171
rect 54238 -1225 54294 -1223
rect 54878 -1067 54934 -1065
rect 54878 -1119 54880 -1067
rect 54880 -1119 54932 -1067
rect 54932 -1119 54934 -1067
rect 54878 -1121 54934 -1119
rect 54878 -1171 54934 -1169
rect 54878 -1223 54880 -1171
rect 54880 -1223 54932 -1171
rect 54932 -1223 54934 -1171
rect 54878 -1225 54934 -1223
rect 56454 -1067 56510 -1065
rect 56454 -1119 56456 -1067
rect 56456 -1119 56508 -1067
rect 56508 -1119 56510 -1067
rect 56454 -1121 56510 -1119
rect 56454 -1171 56510 -1169
rect 56454 -1223 56456 -1171
rect 56456 -1223 56508 -1171
rect 56508 -1223 56510 -1171
rect 56454 -1225 56510 -1223
rect 57094 -1067 57150 -1065
rect 57094 -1119 57096 -1067
rect 57096 -1119 57148 -1067
rect 57148 -1119 57150 -1067
rect 57094 -1121 57150 -1119
rect 57094 -1171 57150 -1169
rect 57094 -1223 57096 -1171
rect 57096 -1223 57148 -1171
rect 57148 -1223 57150 -1171
rect 57094 -1225 57150 -1223
rect 58374 -1067 58430 -1065
rect 58374 -1119 58376 -1067
rect 58376 -1119 58428 -1067
rect 58428 -1119 58430 -1067
rect 58374 -1121 58430 -1119
rect 58374 -1171 58430 -1169
rect 58374 -1223 58376 -1171
rect 58376 -1223 58428 -1171
rect 58428 -1223 58430 -1171
rect 58374 -1225 58430 -1223
rect 59014 -1067 59070 -1065
rect 59014 -1119 59016 -1067
rect 59016 -1119 59068 -1067
rect 59068 -1119 59070 -1067
rect 59014 -1121 59070 -1119
rect 59014 -1171 59070 -1169
rect 59014 -1223 59016 -1171
rect 59016 -1223 59068 -1171
rect 59068 -1223 59070 -1171
rect 59014 -1225 59070 -1223
rect 60028 -1121 60084 -1065
rect 60132 -1121 60188 -1065
rect 60236 -1121 60292 -1065
rect 60028 -1225 60084 -1169
rect 60132 -1225 60188 -1169
rect 60236 -1225 60292 -1169
rect 62335 387 62391 389
rect 62335 335 62337 387
rect 62337 335 62389 387
rect 62389 335 62391 387
rect 62335 333 62391 335
rect 62335 283 62391 285
rect 62335 231 62337 283
rect 62337 231 62389 283
rect 62389 231 62391 283
rect 62335 229 62391 231
rect 62975 387 63031 389
rect 62975 335 62977 387
rect 62977 335 63029 387
rect 63029 335 63031 387
rect 62975 333 63031 335
rect 62975 283 63031 285
rect 62975 231 62977 283
rect 62977 231 63029 283
rect 63029 231 63031 283
rect 62975 229 63031 231
rect 62014 -7 62070 -5
rect 62014 -59 62016 -7
rect 62016 -59 62068 -7
rect 62068 -59 62070 -7
rect 62014 -61 62070 -59
rect 62014 -111 62070 -109
rect 62014 -163 62016 -111
rect 62016 -163 62068 -111
rect 62068 -163 62070 -111
rect 62014 -165 62070 -163
rect 62654 -7 62710 -5
rect 62654 -59 62656 -7
rect 62656 -59 62708 -7
rect 62708 -59 62710 -7
rect 62654 -61 62710 -59
rect 62654 -111 62710 -109
rect 62654 -163 62656 -111
rect 62656 -163 62708 -111
rect 62708 -163 62710 -111
rect 62654 -165 62710 -163
rect 63615 387 63671 389
rect 63615 335 63617 387
rect 63617 335 63669 387
rect 63669 335 63671 387
rect 63615 333 63671 335
rect 63615 283 63671 285
rect 63615 231 63617 283
rect 63617 231 63669 283
rect 63669 231 63671 283
rect 63615 229 63671 231
rect 64255 387 64311 389
rect 64255 335 64257 387
rect 64257 335 64309 387
rect 64309 335 64311 387
rect 64255 333 64311 335
rect 64255 283 64311 285
rect 64255 231 64257 283
rect 64257 231 64309 283
rect 64309 231 64311 283
rect 64255 229 64311 231
rect 63934 -7 63990 -5
rect 63934 -59 63936 -7
rect 63936 -59 63988 -7
rect 63988 -59 63990 -7
rect 63934 -61 63990 -59
rect 63934 -111 63990 -109
rect 63934 -163 63936 -111
rect 63936 -163 63988 -111
rect 63988 -163 63990 -111
rect 63934 -165 63990 -163
rect 64574 -7 64630 -5
rect 64574 -59 64576 -7
rect 64576 -59 64628 -7
rect 64628 -59 64630 -7
rect 64574 -61 64630 -59
rect 64574 -111 64630 -109
rect 64574 -163 64576 -111
rect 64576 -163 64628 -111
rect 64628 -163 64630 -111
rect 64574 -165 64630 -163
rect 62335 -673 62391 -671
rect 62335 -725 62337 -673
rect 62337 -725 62389 -673
rect 62389 -725 62391 -673
rect 62335 -727 62391 -725
rect 62335 -777 62391 -775
rect 62335 -829 62337 -777
rect 62337 -829 62389 -777
rect 62389 -829 62391 -777
rect 62335 -831 62391 -829
rect 62975 -673 63031 -671
rect 62975 -725 62977 -673
rect 62977 -725 63029 -673
rect 63029 -725 63031 -673
rect 62975 -727 63031 -725
rect 62975 -777 63031 -775
rect 62975 -829 62977 -777
rect 62977 -829 63029 -777
rect 63029 -829 63031 -777
rect 62975 -831 63031 -829
rect 63615 -673 63671 -671
rect 63615 -725 63617 -673
rect 63617 -725 63669 -673
rect 63669 -725 63671 -673
rect 63615 -727 63671 -725
rect 63615 -777 63671 -775
rect 63615 -829 63617 -777
rect 63617 -829 63669 -777
rect 63669 -829 63671 -777
rect 63615 -831 63671 -829
rect 64255 -673 64311 -671
rect 64255 -725 64257 -673
rect 64257 -725 64309 -673
rect 64309 -725 64311 -673
rect 64255 -727 64311 -725
rect 64255 -777 64311 -775
rect 64255 -829 64257 -777
rect 64257 -829 64309 -777
rect 64309 -829 64311 -777
rect 64255 -831 64311 -829
rect 60792 -1017 60848 -961
rect 60896 -1017 60952 -961
rect 61000 -1017 61056 -961
rect 60792 -1121 60848 -1065
rect 60896 -1121 60952 -1065
rect 61000 -1121 61056 -1065
rect 60792 -1225 60848 -1169
rect 60896 -1225 60952 -1169
rect 61000 -1225 61056 -1169
rect 62014 -1067 62070 -1065
rect 62014 -1119 62016 -1067
rect 62016 -1119 62068 -1067
rect 62068 -1119 62070 -1067
rect 62014 -1121 62070 -1119
rect 62014 -1171 62070 -1169
rect 62014 -1223 62016 -1171
rect 62016 -1223 62068 -1171
rect 62068 -1223 62070 -1171
rect 62014 -1225 62070 -1223
rect 62654 -1067 62710 -1065
rect 62654 -1119 62656 -1067
rect 62656 -1119 62708 -1067
rect 62708 -1119 62710 -1067
rect 62654 -1121 62710 -1119
rect 62654 -1171 62710 -1169
rect 62654 -1223 62656 -1171
rect 62656 -1223 62708 -1171
rect 62708 -1223 62710 -1171
rect 62654 -1225 62710 -1223
rect 63934 -1067 63990 -1065
rect 63934 -1119 63936 -1067
rect 63936 -1119 63988 -1067
rect 63988 -1119 63990 -1067
rect 63934 -1121 63990 -1119
rect 63934 -1171 63990 -1169
rect 63934 -1223 63936 -1171
rect 63936 -1223 63988 -1171
rect 63988 -1223 63990 -1171
rect 63934 -1225 63990 -1223
rect 64574 -1067 64630 -1065
rect 64574 -1119 64576 -1067
rect 64576 -1119 64628 -1067
rect 64628 -1119 64630 -1067
rect 64574 -1121 64630 -1119
rect 64574 -1171 64630 -1169
rect 64574 -1223 64576 -1171
rect 64576 -1223 64628 -1171
rect 64628 -1223 64630 -1171
rect 64574 -1225 64630 -1223
rect 34154 -5649 34210 -5593
rect 34258 -5649 34314 -5593
rect 34154 -5753 34210 -5697
rect 34258 -5753 34314 -5697
rect 44546 -7956 44602 -7954
rect 44546 -8008 44548 -7956
rect 44548 -8008 44600 -7956
rect 44600 -8008 44602 -7956
rect 44546 -8010 44602 -8008
rect 44650 -7956 44706 -7954
rect 44650 -8008 44652 -7956
rect 44652 -8008 44704 -7956
rect 44704 -8008 44706 -7956
rect 44650 -8010 44706 -8008
rect 44754 -7956 44810 -7954
rect 44754 -8008 44756 -7956
rect 44756 -8008 44808 -7956
rect 44808 -8008 44810 -7956
rect 44754 -8010 44810 -8008
rect 44858 -7956 44914 -7954
rect 44858 -8008 44860 -7956
rect 44860 -8008 44912 -7956
rect 44912 -8008 44914 -7956
rect 44858 -8010 44914 -8008
rect 44962 -7956 45018 -7954
rect 44962 -8008 44964 -7956
rect 44964 -8008 45016 -7956
rect 45016 -8008 45018 -7956
rect 44962 -8010 45018 -8008
rect 34716 -8056 34772 -8054
rect 34716 -8108 34718 -8056
rect 34718 -8108 34770 -8056
rect 34770 -8108 34772 -8056
rect 34716 -8110 34772 -8108
rect 34820 -8056 34876 -8054
rect 34820 -8108 34822 -8056
rect 34822 -8108 34874 -8056
rect 34874 -8108 34876 -8056
rect 34820 -8110 34876 -8108
rect 34924 -8056 34980 -8054
rect 34924 -8108 34926 -8056
rect 34926 -8108 34978 -8056
rect 34978 -8108 34980 -8056
rect 34924 -8110 34980 -8108
rect 35028 -8056 35084 -8054
rect 35028 -8108 35030 -8056
rect 35030 -8108 35082 -8056
rect 35082 -8108 35084 -8056
rect 35028 -8110 35084 -8108
rect 35132 -8056 35188 -8054
rect 35132 -8108 35134 -8056
rect 35134 -8108 35186 -8056
rect 35186 -8108 35188 -8056
rect 35132 -8110 35188 -8108
rect 34716 -8160 34772 -8158
rect 34716 -8212 34718 -8160
rect 34718 -8212 34770 -8160
rect 34770 -8212 34772 -8160
rect 34716 -8214 34772 -8212
rect 34820 -8160 34876 -8158
rect 34820 -8212 34822 -8160
rect 34822 -8212 34874 -8160
rect 34874 -8212 34876 -8160
rect 34820 -8214 34876 -8212
rect 34924 -8160 34980 -8158
rect 34924 -8212 34926 -8160
rect 34926 -8212 34978 -8160
rect 34978 -8212 34980 -8160
rect 34924 -8214 34980 -8212
rect 35028 -8160 35084 -8158
rect 35028 -8212 35030 -8160
rect 35030 -8212 35082 -8160
rect 35082 -8212 35084 -8160
rect 35028 -8214 35084 -8212
rect 35132 -8160 35188 -8158
rect 35132 -8212 35134 -8160
rect 35134 -8212 35186 -8160
rect 35186 -8212 35188 -8160
rect 35132 -8214 35188 -8212
rect 34716 -8264 34772 -8262
rect 34716 -8316 34718 -8264
rect 34718 -8316 34770 -8264
rect 34770 -8316 34772 -8264
rect 34716 -8318 34772 -8316
rect 34820 -8264 34876 -8262
rect 34820 -8316 34822 -8264
rect 34822 -8316 34874 -8264
rect 34874 -8316 34876 -8264
rect 34820 -8318 34876 -8316
rect 34924 -8264 34980 -8262
rect 34924 -8316 34926 -8264
rect 34926 -8316 34978 -8264
rect 34978 -8316 34980 -8264
rect 34924 -8318 34980 -8316
rect 35028 -8264 35084 -8262
rect 35028 -8316 35030 -8264
rect 35030 -8316 35082 -8264
rect 35082 -8316 35084 -8264
rect 35028 -8318 35084 -8316
rect 35132 -8264 35188 -8262
rect 35132 -8316 35134 -8264
rect 35134 -8316 35186 -8264
rect 35186 -8316 35188 -8264
rect 35132 -8318 35188 -8316
rect 34716 -8368 34772 -8366
rect 34716 -8420 34718 -8368
rect 34718 -8420 34770 -8368
rect 34770 -8420 34772 -8368
rect 34716 -8422 34772 -8420
rect 34820 -8368 34876 -8366
rect 34820 -8420 34822 -8368
rect 34822 -8420 34874 -8368
rect 34874 -8420 34876 -8368
rect 34820 -8422 34876 -8420
rect 34924 -8368 34980 -8366
rect 34924 -8420 34926 -8368
rect 34926 -8420 34978 -8368
rect 34978 -8420 34980 -8368
rect 34924 -8422 34980 -8420
rect 35028 -8368 35084 -8366
rect 35028 -8420 35030 -8368
rect 35030 -8420 35082 -8368
rect 35082 -8420 35084 -8368
rect 35028 -8422 35084 -8420
rect 35132 -8368 35188 -8366
rect 35132 -8420 35134 -8368
rect 35134 -8420 35186 -8368
rect 35186 -8420 35188 -8368
rect 35132 -8422 35188 -8420
rect 34716 -8472 34772 -8470
rect 34716 -8524 34718 -8472
rect 34718 -8524 34770 -8472
rect 34770 -8524 34772 -8472
rect 34716 -8526 34772 -8524
rect 34820 -8472 34876 -8470
rect 34820 -8524 34822 -8472
rect 34822 -8524 34874 -8472
rect 34874 -8524 34876 -8472
rect 34820 -8526 34876 -8524
rect 34924 -8472 34980 -8470
rect 34924 -8524 34926 -8472
rect 34926 -8524 34978 -8472
rect 34978 -8524 34980 -8472
rect 34924 -8526 34980 -8524
rect 35028 -8472 35084 -8470
rect 35028 -8524 35030 -8472
rect 35030 -8524 35082 -8472
rect 35082 -8524 35084 -8472
rect 35028 -8526 35084 -8524
rect 35132 -8472 35188 -8470
rect 35132 -8524 35134 -8472
rect 35134 -8524 35186 -8472
rect 35186 -8524 35188 -8472
rect 35132 -8526 35188 -8524
rect 39156 -8056 39212 -8054
rect 39156 -8108 39158 -8056
rect 39158 -8108 39210 -8056
rect 39210 -8108 39212 -8056
rect 39156 -8110 39212 -8108
rect 39260 -8056 39316 -8054
rect 39260 -8108 39262 -8056
rect 39262 -8108 39314 -8056
rect 39314 -8108 39316 -8056
rect 39260 -8110 39316 -8108
rect 39364 -8056 39420 -8054
rect 39364 -8108 39366 -8056
rect 39366 -8108 39418 -8056
rect 39418 -8108 39420 -8056
rect 39364 -8110 39420 -8108
rect 39468 -8056 39524 -8054
rect 39468 -8108 39470 -8056
rect 39470 -8108 39522 -8056
rect 39522 -8108 39524 -8056
rect 39468 -8110 39524 -8108
rect 39572 -8056 39628 -8054
rect 39572 -8108 39574 -8056
rect 39574 -8108 39626 -8056
rect 39626 -8108 39628 -8056
rect 39572 -8110 39628 -8108
rect 39156 -8160 39212 -8158
rect 39156 -8212 39158 -8160
rect 39158 -8212 39210 -8160
rect 39210 -8212 39212 -8160
rect 39156 -8214 39212 -8212
rect 39260 -8160 39316 -8158
rect 39260 -8212 39262 -8160
rect 39262 -8212 39314 -8160
rect 39314 -8212 39316 -8160
rect 39260 -8214 39316 -8212
rect 39364 -8160 39420 -8158
rect 39364 -8212 39366 -8160
rect 39366 -8212 39418 -8160
rect 39418 -8212 39420 -8160
rect 39364 -8214 39420 -8212
rect 39468 -8160 39524 -8158
rect 39468 -8212 39470 -8160
rect 39470 -8212 39522 -8160
rect 39522 -8212 39524 -8160
rect 39468 -8214 39524 -8212
rect 39572 -8160 39628 -8158
rect 39572 -8212 39574 -8160
rect 39574 -8212 39626 -8160
rect 39626 -8212 39628 -8160
rect 39572 -8214 39628 -8212
rect 39156 -8264 39212 -8262
rect 39156 -8316 39158 -8264
rect 39158 -8316 39210 -8264
rect 39210 -8316 39212 -8264
rect 39156 -8318 39212 -8316
rect 39260 -8264 39316 -8262
rect 39260 -8316 39262 -8264
rect 39262 -8316 39314 -8264
rect 39314 -8316 39316 -8264
rect 39260 -8318 39316 -8316
rect 39364 -8264 39420 -8262
rect 39364 -8316 39366 -8264
rect 39366 -8316 39418 -8264
rect 39418 -8316 39420 -8264
rect 39364 -8318 39420 -8316
rect 39468 -8264 39524 -8262
rect 39468 -8316 39470 -8264
rect 39470 -8316 39522 -8264
rect 39522 -8316 39524 -8264
rect 39468 -8318 39524 -8316
rect 39572 -8264 39628 -8262
rect 39572 -8316 39574 -8264
rect 39574 -8316 39626 -8264
rect 39626 -8316 39628 -8264
rect 39572 -8318 39628 -8316
rect 39156 -8368 39212 -8366
rect 39156 -8420 39158 -8368
rect 39158 -8420 39210 -8368
rect 39210 -8420 39212 -8368
rect 39156 -8422 39212 -8420
rect 39260 -8368 39316 -8366
rect 39260 -8420 39262 -8368
rect 39262 -8420 39314 -8368
rect 39314 -8420 39316 -8368
rect 39260 -8422 39316 -8420
rect 39364 -8368 39420 -8366
rect 39364 -8420 39366 -8368
rect 39366 -8420 39418 -8368
rect 39418 -8420 39420 -8368
rect 39364 -8422 39420 -8420
rect 39468 -8368 39524 -8366
rect 39468 -8420 39470 -8368
rect 39470 -8420 39522 -8368
rect 39522 -8420 39524 -8368
rect 39468 -8422 39524 -8420
rect 39572 -8368 39628 -8366
rect 39572 -8420 39574 -8368
rect 39574 -8420 39626 -8368
rect 39626 -8420 39628 -8368
rect 39572 -8422 39628 -8420
rect 44546 -8060 44602 -8058
rect 44546 -8112 44548 -8060
rect 44548 -8112 44600 -8060
rect 44600 -8112 44602 -8060
rect 44546 -8114 44602 -8112
rect 44650 -8060 44706 -8058
rect 44650 -8112 44652 -8060
rect 44652 -8112 44704 -8060
rect 44704 -8112 44706 -8060
rect 44650 -8114 44706 -8112
rect 44754 -8060 44810 -8058
rect 44754 -8112 44756 -8060
rect 44756 -8112 44808 -8060
rect 44808 -8112 44810 -8060
rect 44754 -8114 44810 -8112
rect 44858 -8060 44914 -8058
rect 44858 -8112 44860 -8060
rect 44860 -8112 44912 -8060
rect 44912 -8112 44914 -8060
rect 44858 -8114 44914 -8112
rect 44962 -8060 45018 -8058
rect 44962 -8112 44964 -8060
rect 44964 -8112 45016 -8060
rect 45016 -8112 45018 -8060
rect 44962 -8114 45018 -8112
rect 44546 -8164 44602 -8162
rect 44546 -8216 44548 -8164
rect 44548 -8216 44600 -8164
rect 44600 -8216 44602 -8164
rect 44546 -8218 44602 -8216
rect 44650 -8164 44706 -8162
rect 44650 -8216 44652 -8164
rect 44652 -8216 44704 -8164
rect 44704 -8216 44706 -8164
rect 44650 -8218 44706 -8216
rect 44754 -8164 44810 -8162
rect 44754 -8216 44756 -8164
rect 44756 -8216 44808 -8164
rect 44808 -8216 44810 -8164
rect 44754 -8218 44810 -8216
rect 44858 -8164 44914 -8162
rect 44858 -8216 44860 -8164
rect 44860 -8216 44912 -8164
rect 44912 -8216 44914 -8164
rect 44858 -8218 44914 -8216
rect 44962 -8164 45018 -8162
rect 44962 -8216 44964 -8164
rect 44964 -8216 45016 -8164
rect 45016 -8216 45018 -8164
rect 44962 -8218 45018 -8216
rect 44546 -8268 44602 -8266
rect 44546 -8320 44548 -8268
rect 44548 -8320 44600 -8268
rect 44600 -8320 44602 -8268
rect 44546 -8322 44602 -8320
rect 44650 -8268 44706 -8266
rect 44650 -8320 44652 -8268
rect 44652 -8320 44704 -8268
rect 44704 -8320 44706 -8268
rect 44650 -8322 44706 -8320
rect 44754 -8268 44810 -8266
rect 44754 -8320 44756 -8268
rect 44756 -8320 44808 -8268
rect 44808 -8320 44810 -8268
rect 44754 -8322 44810 -8320
rect 44858 -8268 44914 -8266
rect 44858 -8320 44860 -8268
rect 44860 -8320 44912 -8268
rect 44912 -8320 44914 -8268
rect 44858 -8322 44914 -8320
rect 44962 -8268 45018 -8266
rect 44962 -8320 44964 -8268
rect 44964 -8320 45016 -8268
rect 45016 -8320 45018 -8268
rect 44962 -8322 45018 -8320
rect 44546 -8372 44602 -8370
rect 44546 -8424 44548 -8372
rect 44548 -8424 44600 -8372
rect 44600 -8424 44602 -8372
rect 44546 -8426 44602 -8424
rect 44650 -8372 44706 -8370
rect 44650 -8424 44652 -8372
rect 44652 -8424 44704 -8372
rect 44704 -8424 44706 -8372
rect 44650 -8426 44706 -8424
rect 44754 -8372 44810 -8370
rect 44754 -8424 44756 -8372
rect 44756 -8424 44808 -8372
rect 44808 -8424 44810 -8372
rect 44754 -8426 44810 -8424
rect 44858 -8372 44914 -8370
rect 44858 -8424 44860 -8372
rect 44860 -8424 44912 -8372
rect 44912 -8424 44914 -8372
rect 44858 -8426 44914 -8424
rect 44962 -8372 45018 -8370
rect 44962 -8424 44964 -8372
rect 44964 -8424 45016 -8372
rect 45016 -8424 45018 -8372
rect 44962 -8426 45018 -8424
rect 48986 -7956 49042 -7954
rect 48986 -8008 48988 -7956
rect 48988 -8008 49040 -7956
rect 49040 -8008 49042 -7956
rect 48986 -8010 49042 -8008
rect 49090 -7956 49146 -7954
rect 49090 -8008 49092 -7956
rect 49092 -8008 49144 -7956
rect 49144 -8008 49146 -7956
rect 49090 -8010 49146 -8008
rect 49194 -7956 49250 -7954
rect 49194 -8008 49196 -7956
rect 49196 -8008 49248 -7956
rect 49248 -8008 49250 -7956
rect 49194 -8010 49250 -8008
rect 49298 -7956 49354 -7954
rect 49298 -8008 49300 -7956
rect 49300 -8008 49352 -7956
rect 49352 -8008 49354 -7956
rect 49298 -8010 49354 -8008
rect 49402 -7956 49458 -7954
rect 49402 -8008 49404 -7956
rect 49404 -8008 49456 -7956
rect 49456 -8008 49458 -7956
rect 49402 -8010 49458 -8008
rect 48986 -8060 49042 -8058
rect 48986 -8112 48988 -8060
rect 48988 -8112 49040 -8060
rect 49040 -8112 49042 -8060
rect 48986 -8114 49042 -8112
rect 49090 -8060 49146 -8058
rect 49090 -8112 49092 -8060
rect 49092 -8112 49144 -8060
rect 49144 -8112 49146 -8060
rect 49090 -8114 49146 -8112
rect 49194 -8060 49250 -8058
rect 49194 -8112 49196 -8060
rect 49196 -8112 49248 -8060
rect 49248 -8112 49250 -8060
rect 49194 -8114 49250 -8112
rect 49298 -8060 49354 -8058
rect 49298 -8112 49300 -8060
rect 49300 -8112 49352 -8060
rect 49352 -8112 49354 -8060
rect 49298 -8114 49354 -8112
rect 49402 -8060 49458 -8058
rect 49402 -8112 49404 -8060
rect 49404 -8112 49456 -8060
rect 49456 -8112 49458 -8060
rect 49402 -8114 49458 -8112
rect 48986 -8164 49042 -8162
rect 48986 -8216 48988 -8164
rect 48988 -8216 49040 -8164
rect 49040 -8216 49042 -8164
rect 48986 -8218 49042 -8216
rect 49090 -8164 49146 -8162
rect 49090 -8216 49092 -8164
rect 49092 -8216 49144 -8164
rect 49144 -8216 49146 -8164
rect 49090 -8218 49146 -8216
rect 49194 -8164 49250 -8162
rect 49194 -8216 49196 -8164
rect 49196 -8216 49248 -8164
rect 49248 -8216 49250 -8164
rect 49194 -8218 49250 -8216
rect 49298 -8164 49354 -8162
rect 49298 -8216 49300 -8164
rect 49300 -8216 49352 -8164
rect 49352 -8216 49354 -8164
rect 49298 -8218 49354 -8216
rect 49402 -8164 49458 -8162
rect 49402 -8216 49404 -8164
rect 49404 -8216 49456 -8164
rect 49456 -8216 49458 -8164
rect 49402 -8218 49458 -8216
rect 48986 -8268 49042 -8266
rect 48986 -8320 48988 -8268
rect 48988 -8320 49040 -8268
rect 49040 -8320 49042 -8268
rect 48986 -8322 49042 -8320
rect 49090 -8268 49146 -8266
rect 49090 -8320 49092 -8268
rect 49092 -8320 49144 -8268
rect 49144 -8320 49146 -8268
rect 49090 -8322 49146 -8320
rect 49194 -8268 49250 -8266
rect 49194 -8320 49196 -8268
rect 49196 -8320 49248 -8268
rect 49248 -8320 49250 -8268
rect 49194 -8322 49250 -8320
rect 49298 -8268 49354 -8266
rect 49298 -8320 49300 -8268
rect 49300 -8320 49352 -8268
rect 49352 -8320 49354 -8268
rect 49298 -8322 49354 -8320
rect 49402 -8268 49458 -8266
rect 49402 -8320 49404 -8268
rect 49404 -8320 49456 -8268
rect 49456 -8320 49458 -8268
rect 49402 -8322 49458 -8320
rect 48986 -8372 49042 -8370
rect 48986 -8424 48988 -8372
rect 48988 -8424 49040 -8372
rect 49040 -8424 49042 -8372
rect 48986 -8426 49042 -8424
rect 49090 -8372 49146 -8370
rect 49090 -8424 49092 -8372
rect 49092 -8424 49144 -8372
rect 49144 -8424 49146 -8372
rect 49090 -8426 49146 -8424
rect 49194 -8372 49250 -8370
rect 49194 -8424 49196 -8372
rect 49196 -8424 49248 -8372
rect 49248 -8424 49250 -8372
rect 49194 -8426 49250 -8424
rect 49298 -8372 49354 -8370
rect 49298 -8424 49300 -8372
rect 49300 -8424 49352 -8372
rect 49352 -8424 49354 -8372
rect 49298 -8426 49354 -8424
rect 49402 -8372 49458 -8370
rect 49402 -8424 49404 -8372
rect 49404 -8424 49456 -8372
rect 49456 -8424 49458 -8372
rect 49402 -8426 49458 -8424
rect 39156 -8472 39212 -8470
rect 39156 -8524 39158 -8472
rect 39158 -8524 39210 -8472
rect 39210 -8524 39212 -8472
rect 39156 -8526 39212 -8524
rect 39260 -8472 39316 -8470
rect 39260 -8524 39262 -8472
rect 39262 -8524 39314 -8472
rect 39314 -8524 39316 -8472
rect 39260 -8526 39316 -8524
rect 39364 -8472 39420 -8470
rect 39364 -8524 39366 -8472
rect 39366 -8524 39418 -8472
rect 39418 -8524 39420 -8472
rect 39364 -8526 39420 -8524
rect 39468 -8472 39524 -8470
rect 39468 -8524 39470 -8472
rect 39470 -8524 39522 -8472
rect 39522 -8524 39524 -8472
rect 39468 -8526 39524 -8524
rect 39572 -8472 39628 -8470
rect 39572 -8524 39574 -8472
rect 39574 -8524 39626 -8472
rect 39626 -8524 39628 -8472
rect 39572 -8526 39628 -8524
rect 31650 -8827 31706 -8771
rect 31754 -8827 31810 -8771
rect 31858 -8827 31914 -8771
rect 31650 -8931 31706 -8875
rect 31754 -8931 31810 -8875
rect 31858 -8931 31914 -8875
rect 31650 -9035 31706 -8979
rect 31754 -9035 31810 -8979
rect 31858 -9035 31914 -8979
rect 16967 -9447 17023 -9391
rect 17077 -9447 17133 -9391
rect 16967 -9557 17023 -9501
rect 17077 -9557 17133 -9501
rect 14946 -9689 15002 -9633
rect 15056 -9689 15112 -9633
rect 14946 -9799 15002 -9743
rect 15056 -9799 15112 -9743
rect 12983 -9931 13039 -9875
rect 13093 -9931 13149 -9875
rect 12983 -10041 13039 -9985
rect 13093 -10041 13149 -9985
rect 10976 -10176 11032 -10120
rect 11086 -10176 11142 -10120
rect 10976 -10286 11032 -10230
rect 11086 -10286 11142 -10230
rect 8941 -10412 8997 -10356
rect 9051 -10412 9107 -10356
rect 8941 -10522 8997 -10466
rect 9051 -10522 9107 -10466
rect 6854 -10654 6910 -10598
rect 6964 -10654 7020 -10598
rect 6854 -10764 6910 -10708
rect 6964 -10764 7020 -10708
rect -1086 -11498 -1030 -11442
rect -976 -11498 -920 -11442
rect -858 -11498 -802 -11442
rect -748 -11498 -692 -11442
rect -1086 -11608 -1030 -11552
rect -976 -11608 -920 -11552
rect -858 -11608 -802 -11552
rect -748 -11608 -692 -11552
rect 8401 -11481 8457 -11425
rect 8511 -11481 8567 -11425
rect 8401 -11591 8457 -11535
rect 8511 -11591 8567 -11535
rect 10404 -11457 10460 -11401
rect 10514 -11457 10570 -11401
rect 10404 -11567 10460 -11511
rect 10514 -11567 10570 -11511
rect 7132 -13016 7188 -12960
rect 7242 -13016 7298 -12960
rect 12428 -11453 12484 -11397
rect 12538 -11453 12594 -11397
rect 12428 -11563 12484 -11507
rect 12538 -11563 12594 -11507
rect 7088 -13166 7144 -13110
rect 7198 -13166 7254 -13110
rect 9156 -13166 9212 -13110
rect 9266 -13166 9322 -13110
rect 6704 -13466 6760 -13410
rect 6814 -13466 6870 -13410
rect 6464 -13766 6520 -13710
rect 6574 -13766 6630 -13710
rect 14462 -11444 14518 -11388
rect 14572 -11444 14628 -11388
rect 14462 -11554 14518 -11498
rect 14572 -11554 14628 -11498
rect 11176 -13316 11232 -13260
rect 11286 -13316 11342 -13260
rect 16458 -11443 16514 -11387
rect 16568 -11443 16624 -11387
rect 16458 -11553 16514 -11497
rect 16568 -11553 16624 -11497
rect 13166 -13466 13222 -13410
rect 13276 -13466 13332 -13410
rect 18448 -11440 18504 -11384
rect 18558 -11440 18614 -11384
rect 18448 -11550 18504 -11494
rect 18558 -11550 18614 -11494
rect 15193 -13616 15249 -13560
rect 15303 -13616 15359 -13560
rect 17445 -13016 17501 -12960
rect 17555 -13016 17611 -12960
rect 17122 -13766 17178 -13710
rect 17232 -13766 17288 -13710
rect 17628 -13316 17684 -13260
rect 17738 -13316 17794 -13260
rect 17785 -13616 17841 -13560
rect 17895 -13616 17951 -13560
rect 33967 -9447 34023 -9391
rect 34077 -9447 34133 -9391
rect 33967 -9557 34023 -9501
rect 34077 -9557 34133 -9501
rect 31946 -9689 32002 -9633
rect 32056 -9689 32112 -9633
rect 31946 -9799 32002 -9743
rect 32056 -9799 32112 -9743
rect 29983 -9931 30039 -9875
rect 30093 -9931 30149 -9875
rect 29983 -10041 30039 -9985
rect 30093 -10041 30149 -9985
rect 27976 -10176 28032 -10120
rect 28086 -10176 28142 -10120
rect 27976 -10286 28032 -10230
rect 28086 -10286 28142 -10230
rect 25941 -10412 25997 -10356
rect 26051 -10412 26107 -10356
rect 25941 -10522 25997 -10466
rect 26051 -10522 26107 -10466
rect 23854 -10654 23910 -10598
rect 23964 -10654 24020 -10598
rect 23854 -10764 23910 -10708
rect 23964 -10764 24020 -10708
rect 25395 -11033 25451 -10977
rect 25505 -11033 25561 -10977
rect 25395 -11143 25451 -11087
rect 25505 -11143 25561 -11087
rect 27397 -11003 27453 -10947
rect 27507 -11003 27563 -10947
rect 27397 -11113 27453 -11057
rect 27507 -11113 27563 -11057
rect 24132 -13016 24188 -12960
rect 24242 -13016 24298 -12960
rect 29450 -10993 29506 -10937
rect 29560 -10993 29616 -10937
rect 29450 -11103 29506 -11047
rect 29560 -11103 29616 -11047
rect 24088 -13166 24144 -13110
rect 24198 -13166 24254 -13110
rect 26156 -13166 26212 -13110
rect 26266 -13166 26322 -13110
rect 23704 -13466 23760 -13410
rect 23814 -13466 23870 -13410
rect 23464 -13766 23520 -13710
rect 23574 -13766 23630 -13710
rect 31453 -10989 31509 -10933
rect 31563 -10989 31619 -10933
rect 31453 -11099 31509 -11043
rect 31563 -11099 31619 -11043
rect 28176 -13316 28232 -13260
rect 28286 -13316 28342 -13260
rect 33506 -10989 33562 -10933
rect 33616 -10989 33672 -10933
rect 33506 -11099 33562 -11043
rect 33616 -11099 33672 -11043
rect 30166 -13466 30222 -13410
rect 30276 -13466 30332 -13410
rect 35557 -10989 35613 -10933
rect 35667 -10989 35723 -10933
rect 35557 -11099 35613 -11043
rect 35667 -11099 35723 -11043
rect 32193 -13616 32249 -13560
rect 32303 -13616 32359 -13560
rect 34445 -13016 34501 -12960
rect 34555 -13016 34611 -12960
rect 34122 -13766 34178 -13710
rect 34232 -13766 34288 -13710
rect 34628 -13316 34684 -13260
rect 34738 -13316 34794 -13260
rect 34785 -13616 34841 -13560
rect 34895 -13616 34951 -13560
rect 54233 -9447 54289 -9391
rect 54343 -9447 54399 -9391
rect 54233 -9557 54289 -9501
rect 54343 -9557 54399 -9501
rect 54452 -9689 54508 -9633
rect 54562 -9689 54618 -9633
rect 54452 -9799 54508 -9743
rect 54562 -9799 54618 -9743
rect 54754 -9931 54810 -9875
rect 54864 -9931 54920 -9875
rect 54754 -10041 54810 -9985
rect 54864 -10041 54920 -9985
rect 54990 -10176 55046 -10120
rect 55100 -10176 55156 -10120
rect 54990 -10286 55046 -10230
rect 55100 -10286 55156 -10230
rect 55251 -10412 55307 -10356
rect 55361 -10412 55417 -10356
rect 55251 -10522 55307 -10466
rect 55361 -10522 55417 -10466
rect 55568 -10653 55624 -10597
rect 55678 -10653 55734 -10597
rect 55568 -10763 55624 -10707
rect 55678 -10763 55734 -10707
<< metal3 >>
rect 2675 5171 2855 5181
rect 3464 5171 3540 5181
rect 2675 5115 2685 5171
rect 2741 5115 2789 5171
rect 2845 5115 3474 5171
rect 3530 5115 3540 5171
rect 2675 5067 3540 5115
rect 2675 5011 2685 5067
rect 2741 5011 2789 5067
rect 2845 5011 3474 5067
rect 3530 5011 3540 5067
rect 2675 5001 2855 5011
rect 3464 5001 3540 5011
rect 5245 5117 5425 5127
rect 6249 5117 6325 5127
rect 6889 5117 6965 5127
rect 7529 5117 7605 5127
rect 5245 5061 5255 5117
rect 5311 5061 5359 5117
rect 5415 5061 6259 5117
rect 6315 5061 6899 5117
rect 6955 5061 7539 5117
rect 7595 5061 7605 5117
rect 5245 5013 7605 5061
rect 5245 4957 5255 5013
rect 5311 4957 5359 5013
rect 5415 4957 6259 5013
rect 6315 4957 6899 5013
rect 6955 4957 7539 5013
rect 7595 4957 7605 5013
rect 5245 4947 5425 4957
rect 6249 4947 6325 4957
rect 6889 4947 6965 4957
rect 7529 4947 7605 4957
rect 2034 4822 2214 4832
rect 3544 4822 3620 4832
rect 2034 4766 2044 4822
rect 2100 4766 2148 4822
rect 2204 4766 3554 4822
rect 3610 4766 3620 4822
rect 2034 4718 3620 4766
rect 2034 4662 2044 4718
rect 2100 4662 2148 4718
rect 2204 4662 3554 4718
rect 3610 4662 3620 4718
rect 2034 4652 2214 4662
rect 3544 4652 3620 4662
rect 3704 4822 3780 4832
rect 4345 4822 4421 4832
rect 5517 4822 5697 4832
rect 6569 4822 6645 4832
rect 7209 4822 7285 4832
rect 3704 4766 3714 4822
rect 3770 4766 4355 4822
rect 4411 4766 5527 4822
rect 5583 4766 5631 4822
rect 5687 4766 6579 4822
rect 6635 4766 7219 4822
rect 7275 4766 7285 4822
rect 3704 4718 7285 4766
rect 3704 4662 3714 4718
rect 3770 4662 4355 4718
rect 4411 4662 5527 4718
rect 5583 4662 5631 4718
rect 5687 4662 6579 4718
rect 6635 4662 7219 4718
rect 7275 4662 7285 4718
rect 3704 4652 3780 4662
rect 4345 4652 4421 4662
rect 5517 4652 5697 4662
rect 6569 4652 6645 4662
rect 7209 4652 7285 4662
rect 3384 4326 3460 4336
rect 4024 4326 4100 4336
rect 4664 4326 4740 4336
rect 5245 4326 5425 4336
rect 3384 4270 3394 4326
rect 3450 4270 4034 4326
rect 4090 4270 4674 4326
rect 4730 4270 5255 4326
rect 5311 4270 5359 4326
rect 5415 4270 5425 4326
rect 3384 4222 5425 4270
rect 11153 4302 11333 4312
rect 11153 4246 11163 4302
rect 11219 4246 11267 4302
rect 11323 4260 11333 4302
rect 11323 4250 18655 4260
rect 11323 4246 17165 4250
rect 6569 4222 6645 4232
rect 7209 4222 7285 4232
rect 3384 4166 3394 4222
rect 3450 4166 4034 4222
rect 4090 4166 4674 4222
rect 4730 4166 5255 4222
rect 5311 4166 5359 4222
rect 5415 4166 6579 4222
rect 6635 4166 7219 4222
rect 7275 4166 7285 4222
rect 3384 4156 3460 4166
rect 4024 4156 4100 4166
rect 4664 4156 4740 4166
rect 5245 4118 7285 4166
rect 11153 4198 17165 4246
rect 11153 4142 11163 4198
rect 11219 4142 11267 4198
rect 11323 4194 17165 4198
rect 17221 4194 18589 4250
rect 18645 4194 18655 4250
rect 11323 4184 18655 4194
rect 19699 4250 23807 4260
rect 19699 4194 19709 4250
rect 19765 4194 23741 4250
rect 23797 4194 23807 4250
rect 19699 4184 23807 4194
rect 24851 4250 27776 4260
rect 24851 4194 24861 4250
rect 24917 4194 26285 4250
rect 26342 4194 27710 4250
rect 27766 4194 27776 4250
rect 24851 4184 27776 4194
rect 11323 4142 11333 4184
rect 11153 4132 11333 4142
rect 5245 4062 5255 4118
rect 5311 4062 5359 4118
rect 5415 4062 6579 4118
rect 6635 4062 7219 4118
rect 7275 4062 7285 4118
rect 2395 4043 2575 4053
rect 3464 4043 3540 4053
rect 5245 4052 5425 4062
rect 6569 4052 6645 4062
rect 7209 4052 7285 4062
rect 18819 4113 24687 4123
rect 18819 4057 21621 4113
rect 21677 4057 21725 4113
rect 21781 4057 21829 4113
rect 21885 4057 24687 4113
rect 2395 3987 2405 4043
rect 2461 3987 2509 4043
rect 2565 3987 3474 4043
rect 3530 3987 3540 4043
rect 2395 3939 3540 3987
rect 2395 3883 2405 3939
rect 2461 3883 2509 3939
rect 2565 3883 3474 3939
rect 3530 3883 3540 3939
rect 2395 3873 2575 3883
rect 3464 3873 3540 3883
rect 18819 4009 24687 4057
rect 18819 3953 18829 4009
rect 18885 3953 19469 4009
rect 19525 3953 21621 4009
rect 21677 3953 21725 4009
rect 21781 3953 21829 4009
rect 21885 3953 23981 4009
rect 24037 3953 24621 4009
rect 24677 3953 24687 4009
rect 18819 3905 24687 3953
rect 5517 3843 5697 3853
rect 6249 3843 6325 3853
rect 6889 3843 6965 3853
rect 7529 3843 7605 3853
rect 5517 3787 5527 3843
rect 5583 3787 5631 3843
rect 5687 3787 6259 3843
rect 6315 3787 6899 3843
rect 6955 3787 7539 3843
rect 7595 3787 7605 3843
rect 18819 3849 18829 3905
rect 18885 3849 19469 3905
rect 19525 3849 21621 3905
rect 21677 3849 21725 3905
rect 21781 3849 21829 3905
rect 21885 3849 23981 3905
rect 24037 3849 24621 3905
rect 24677 3849 24687 3905
rect 18819 3839 24687 3849
rect 27940 4113 31016 4123
rect 27940 4057 30742 4113
rect 30798 4057 30846 4113
rect 30902 4057 30950 4113
rect 31006 4057 31016 4113
rect 27940 4009 31016 4057
rect 27940 3953 27950 4009
rect 28006 3953 28590 4009
rect 28646 3953 30742 4009
rect 30798 3953 30846 4009
rect 30902 3953 30950 4009
rect 31006 3953 31016 4009
rect 27940 3905 31016 3953
rect 27940 3849 27950 3905
rect 28006 3849 28590 3905
rect 28646 3849 30742 3905
rect 30798 3849 30846 3905
rect 30902 3849 30950 3905
rect 31006 3849 31016 3905
rect 27940 3839 31016 3849
rect 34092 3893 66712 3903
rect 5517 3739 7605 3787
rect 2034 3692 2214 3702
rect 3544 3692 3620 3702
rect 2034 3636 2044 3692
rect 2100 3636 2148 3692
rect 2204 3636 3554 3692
rect 3610 3636 3620 3692
rect 2034 3588 3620 3636
rect 2034 3532 2044 3588
rect 2100 3532 2148 3588
rect 2204 3532 3554 3588
rect 3610 3532 3620 3588
rect 2034 3522 2214 3532
rect 3544 3522 3620 3532
rect 3704 3692 3780 3702
rect 4345 3692 4421 3702
rect 5245 3692 5425 3702
rect 3704 3636 3714 3692
rect 3770 3636 4355 3692
rect 4411 3636 5255 3692
rect 5311 3636 5359 3692
rect 5415 3636 5425 3692
rect 5517 3683 5527 3739
rect 5583 3683 5631 3739
rect 5687 3683 6259 3739
rect 6315 3683 6899 3739
rect 6955 3683 7539 3739
rect 7595 3683 7605 3739
rect 34092 3837 34102 3893
rect 34158 3837 34206 3893
rect 34262 3837 34310 3893
rect 34366 3837 38238 3893
rect 38294 3837 38342 3893
rect 38398 3837 38446 3893
rect 38502 3837 43798 3893
rect 43854 3837 43902 3893
rect 43958 3837 44006 3893
rect 44062 3837 47934 3893
rect 47990 3837 48038 3893
rect 48094 3837 48142 3893
rect 48198 3837 53494 3893
rect 53550 3837 53598 3893
rect 53654 3837 53702 3893
rect 53758 3837 57630 3893
rect 57686 3837 57734 3893
rect 57790 3837 57838 3893
rect 57894 3837 63190 3893
rect 63246 3837 63294 3893
rect 63350 3837 63398 3893
rect 63454 3837 66438 3893
rect 66494 3837 66542 3893
rect 66598 3837 66646 3893
rect 66702 3837 66712 3893
rect 34092 3789 66712 3837
rect 34092 3733 34102 3789
rect 34158 3733 34206 3789
rect 34262 3733 34310 3789
rect 34366 3733 38238 3789
rect 38294 3733 38342 3789
rect 38398 3733 38446 3789
rect 38502 3733 43798 3789
rect 43854 3733 43902 3789
rect 43958 3733 44006 3789
rect 44062 3733 47934 3789
rect 47990 3733 48038 3789
rect 48094 3733 48142 3789
rect 48198 3733 53494 3789
rect 53550 3733 53598 3789
rect 53654 3733 53702 3789
rect 53758 3733 57630 3789
rect 57686 3733 57734 3789
rect 57790 3733 57838 3789
rect 57894 3733 63190 3789
rect 63246 3733 63294 3789
rect 63350 3733 63398 3789
rect 63454 3733 66438 3789
rect 66494 3733 66542 3789
rect 66598 3733 66646 3789
rect 66702 3733 66712 3789
rect 5517 3673 5697 3683
rect 6249 3673 6325 3683
rect 6889 3673 6965 3683
rect 7529 3673 7605 3683
rect 18499 3719 31924 3729
rect 3704 3588 5425 3636
rect 3704 3532 3714 3588
rect 3770 3532 4355 3588
rect 4411 3532 5255 3588
rect 5311 3532 5359 3588
rect 5415 3532 5425 3588
rect 3704 3522 3780 3532
rect 4345 3522 4421 3532
rect 5245 3522 5425 3532
rect 18499 3663 20972 3719
rect 21028 3663 21076 3719
rect 21132 3663 21180 3719
rect 21236 3663 22270 3719
rect 22326 3663 22374 3719
rect 22430 3663 22478 3719
rect 22534 3663 30093 3719
rect 30149 3663 30197 3719
rect 30253 3663 30301 3719
rect 30357 3663 31650 3719
rect 31706 3663 31754 3719
rect 31810 3663 31858 3719
rect 31914 3663 31924 3719
rect 18499 3615 31924 3663
rect 34092 3685 66712 3733
rect 34092 3629 34102 3685
rect 34158 3629 34206 3685
rect 34262 3629 34310 3685
rect 34366 3629 38238 3685
rect 38294 3629 38342 3685
rect 38398 3629 38446 3685
rect 38502 3629 43798 3685
rect 43854 3629 43902 3685
rect 43958 3629 44006 3685
rect 44062 3629 47934 3685
rect 47990 3629 48038 3685
rect 48094 3629 48142 3685
rect 48198 3629 53494 3685
rect 53550 3629 53598 3685
rect 53654 3629 53702 3685
rect 53758 3629 57630 3685
rect 57686 3629 57734 3685
rect 57790 3629 57838 3685
rect 57894 3629 63190 3685
rect 63246 3629 63294 3685
rect 63350 3629 63398 3685
rect 63454 3629 66438 3685
rect 66494 3629 66542 3685
rect 66598 3629 66646 3685
rect 66702 3629 66712 3685
rect 34092 3619 66712 3629
rect 18499 3559 18509 3615
rect 18565 3559 19149 3615
rect 19205 3559 19789 3615
rect 19845 3559 20972 3615
rect 21028 3559 21076 3615
rect 21132 3559 21180 3615
rect 21236 3559 22270 3615
rect 22326 3559 22374 3615
rect 22430 3559 22478 3615
rect 22534 3559 23661 3615
rect 23717 3559 24301 3615
rect 24357 3559 24941 3615
rect 24997 3559 27630 3615
rect 27686 3559 28270 3615
rect 28326 3559 28910 3615
rect 28966 3559 30093 3615
rect 30149 3559 30197 3615
rect 30253 3559 30301 3615
rect 30357 3559 31650 3615
rect 31706 3559 31754 3615
rect 31810 3559 31858 3615
rect 31914 3559 31924 3615
rect 18499 3511 31924 3559
rect 18499 3455 18509 3511
rect 18565 3455 19149 3511
rect 19205 3455 19789 3511
rect 19845 3455 20972 3511
rect 21028 3455 21076 3511
rect 21132 3455 21180 3511
rect 21236 3455 22270 3511
rect 22326 3455 22374 3511
rect 22430 3455 22478 3511
rect 22534 3455 23661 3511
rect 23717 3455 24301 3511
rect 24357 3455 24941 3511
rect 24997 3455 27630 3511
rect 27686 3455 28270 3511
rect 28326 3455 28910 3511
rect 28966 3455 30093 3511
rect 30149 3455 30197 3511
rect 30253 3455 30301 3511
rect 30357 3455 31650 3511
rect 31706 3455 31754 3511
rect 31810 3455 31858 3511
rect 31914 3455 31924 3511
rect 18499 3445 31924 3455
rect 10885 3336 11065 3346
rect 3384 3300 3460 3310
rect 4024 3300 4100 3310
rect 4664 3300 4740 3310
rect 5517 3300 5697 3310
rect 6569 3300 6645 3310
rect 7209 3300 7285 3310
rect 3384 3244 3394 3300
rect 3450 3244 4034 3300
rect 4090 3244 4674 3300
rect 4730 3244 5527 3300
rect 5583 3244 5631 3300
rect 5687 3244 6579 3300
rect 6635 3244 7219 3300
rect 7275 3244 7285 3300
rect 3384 3196 7285 3244
rect 3384 3140 3394 3196
rect 3450 3140 4034 3196
rect 4090 3140 4674 3196
rect 4730 3140 5527 3196
rect 5583 3140 5631 3196
rect 5687 3140 6579 3196
rect 6635 3140 7219 3196
rect 7275 3140 7285 3196
rect 10885 3280 10895 3336
rect 10951 3280 10999 3336
rect 11055 3294 11065 3336
rect 11055 3284 18655 3294
rect 11055 3280 17365 3284
rect 10885 3232 17365 3280
rect 10885 3176 10895 3232
rect 10951 3176 10999 3232
rect 11055 3228 17365 3232
rect 17421 3228 18589 3284
rect 18645 3228 18655 3284
rect 11055 3218 18655 3228
rect 24851 3284 27776 3294
rect 24851 3228 24861 3284
rect 24917 3228 26085 3284
rect 26141 3228 26486 3284
rect 26542 3228 27710 3284
rect 27766 3228 27776 3284
rect 24851 3218 27776 3228
rect 11055 3176 11065 3218
rect 10885 3166 11065 3176
rect 18819 3177 24687 3187
rect 3384 3130 3460 3140
rect 4024 3130 4100 3140
rect 4664 3130 4740 3140
rect 5517 3130 5697 3140
rect 6569 3130 6645 3140
rect 7209 3130 7285 3140
rect 18819 3121 20972 3177
rect 21028 3121 21076 3177
rect 21132 3121 21180 3177
rect 21236 3121 22270 3177
rect 22326 3121 22374 3177
rect 22430 3121 22478 3177
rect 22534 3121 24687 3177
rect 18819 3073 24687 3121
rect 18819 3017 18829 3073
rect 18885 3017 19469 3073
rect 19525 3017 20972 3073
rect 21028 3017 21076 3073
rect 21132 3017 21180 3073
rect 21236 3017 22270 3073
rect 22326 3017 22374 3073
rect 22430 3017 22478 3073
rect 22534 3017 23981 3073
rect 24037 3017 24621 3073
rect 24677 3017 24687 3073
rect 5245 2981 5425 2991
rect 6249 2981 6325 2991
rect 6889 2981 6965 2991
rect 7529 2981 7605 2991
rect 5245 2925 5255 2981
rect 5311 2925 5359 2981
rect 5415 2925 6259 2981
rect 6315 2925 6899 2981
rect 6955 2925 7539 2981
rect 7595 2925 7605 2981
rect 2675 2913 2855 2923
rect 3464 2913 3540 2923
rect 2675 2857 2685 2913
rect 2741 2857 2789 2913
rect 2845 2857 3474 2913
rect 3530 2857 3540 2913
rect 2675 2809 3540 2857
rect 5245 2877 7605 2925
rect 18819 2969 24687 3017
rect 18819 2913 18829 2969
rect 18885 2913 19469 2969
rect 19525 2913 20972 2969
rect 21028 2913 21076 2969
rect 21132 2913 21180 2969
rect 21236 2913 22270 2969
rect 22326 2913 22374 2969
rect 22430 2913 22478 2969
rect 22534 2913 23981 2969
rect 24037 2913 24621 2969
rect 24677 2913 24687 2969
rect 18819 2903 24687 2913
rect 27940 3177 31924 3187
rect 27940 3121 30093 3177
rect 30149 3121 30197 3177
rect 30253 3121 30301 3177
rect 30357 3121 31650 3177
rect 31706 3121 31754 3177
rect 31810 3121 31858 3177
rect 31914 3121 31924 3177
rect 27940 3073 31924 3121
rect 27940 3017 27950 3073
rect 28006 3017 28590 3073
rect 28646 3017 30093 3073
rect 30149 3017 30197 3073
rect 30253 3017 30301 3073
rect 30357 3017 31650 3073
rect 31706 3017 31754 3073
rect 31810 3017 31858 3073
rect 31914 3017 31924 3073
rect 27940 2969 31924 3017
rect 27940 2913 27950 2969
rect 28006 2913 28590 2969
rect 28646 2913 30093 2969
rect 30149 2913 30197 2969
rect 30253 2913 30301 2969
rect 30357 2913 31650 2969
rect 31706 2913 31754 2969
rect 31810 2913 31858 2969
rect 31914 2913 31924 2969
rect 27940 2903 31924 2913
rect 5245 2821 5255 2877
rect 5311 2821 5359 2877
rect 5415 2821 6259 2877
rect 6315 2821 6899 2877
rect 6955 2821 7539 2877
rect 7595 2821 7605 2877
rect 5245 2811 5425 2821
rect 6249 2811 6325 2821
rect 6889 2811 6965 2821
rect 7529 2811 7605 2821
rect 2675 2753 2685 2809
rect 2741 2753 2789 2809
rect 2845 2753 3474 2809
rect 3530 2753 3540 2809
rect 2675 2743 2855 2753
rect 3464 2743 3540 2753
rect 18499 2783 31544 2793
rect 18499 2727 21621 2783
rect 21677 2727 21725 2783
rect 21781 2727 21829 2783
rect 21885 2727 30742 2783
rect 30798 2727 30846 2783
rect 30902 2727 30950 2783
rect 31006 2727 31544 2783
rect 18499 2679 31544 2727
rect 18499 2623 18509 2679
rect 18565 2623 19149 2679
rect 19205 2623 19789 2679
rect 19845 2623 21621 2679
rect 21677 2623 21725 2679
rect 21781 2623 21829 2679
rect 21885 2623 23661 2679
rect 23717 2623 24301 2679
rect 24357 2623 24941 2679
rect 24997 2623 27630 2679
rect 27686 2623 28270 2679
rect 28326 2623 28910 2679
rect 28966 2623 30742 2679
rect 30798 2623 30846 2679
rect 30902 2623 30950 2679
rect 31006 2623 31544 2679
rect 18499 2613 64321 2623
rect 18499 2575 31270 2613
rect 3704 2562 3780 2572
rect 4345 2562 4421 2572
rect 5517 2562 5697 2572
rect 3704 2506 3714 2562
rect 3770 2506 4355 2562
rect 4411 2506 5527 2562
rect 5583 2506 5631 2562
rect 5687 2506 5697 2562
rect 18499 2519 18509 2575
rect 18565 2519 19149 2575
rect 19205 2519 19789 2575
rect 19845 2519 21621 2575
rect 21677 2519 21725 2575
rect 21781 2519 21829 2575
rect 21885 2519 23661 2575
rect 23717 2519 24301 2575
rect 24357 2519 24941 2575
rect 24997 2519 27630 2575
rect 27686 2519 28270 2575
rect 28326 2519 28910 2575
rect 28966 2519 30742 2575
rect 30798 2519 30846 2575
rect 30902 2519 30950 2575
rect 31006 2557 31270 2575
rect 31326 2557 31374 2613
rect 31430 2557 31478 2613
rect 31534 2557 40997 2613
rect 41053 2557 41101 2613
rect 41157 2557 41205 2613
rect 41261 2557 50652 2613
rect 50708 2557 50756 2613
rect 50812 2557 50860 2613
rect 50916 2557 60433 2613
rect 60489 2557 60537 2613
rect 60593 2557 60641 2613
rect 60697 2557 64321 2613
rect 31006 2519 64321 2557
rect 18499 2509 64321 2519
rect 3704 2458 5697 2506
rect 6249 2458 6325 2468
rect 6889 2458 6965 2468
rect 7529 2458 7605 2468
rect 3704 2402 3714 2458
rect 3770 2402 4355 2458
rect 4411 2402 5527 2458
rect 5583 2402 5631 2458
rect 5687 2402 6259 2458
rect 6315 2402 6899 2458
rect 6955 2402 7539 2458
rect 7595 2402 7605 2458
rect 3704 2392 3780 2402
rect 4345 2392 4421 2402
rect 5517 2354 7605 2402
rect 31260 2453 31270 2509
rect 31326 2453 31374 2509
rect 31430 2453 31478 2509
rect 31534 2453 33247 2509
rect 33303 2453 33887 2509
rect 33943 2453 34527 2509
rect 34583 2453 35167 2509
rect 35223 2453 37381 2509
rect 37437 2453 38021 2509
rect 38077 2453 38661 2509
rect 38717 2453 39301 2509
rect 39357 2453 40997 2509
rect 41053 2453 41101 2509
rect 41157 2453 41205 2509
rect 41261 2453 42943 2509
rect 42999 2453 43583 2509
rect 43639 2453 44223 2509
rect 44279 2453 44863 2509
rect 44919 2453 47077 2509
rect 47133 2453 47717 2509
rect 47773 2453 48357 2509
rect 48413 2453 48997 2509
rect 49053 2453 50652 2509
rect 50708 2453 50756 2509
rect 50812 2453 50860 2509
rect 50916 2453 52639 2509
rect 52695 2453 53279 2509
rect 53335 2453 53919 2509
rect 53975 2453 54559 2509
rect 54615 2453 56773 2509
rect 56829 2453 57413 2509
rect 57469 2453 58053 2509
rect 58109 2453 58693 2509
rect 58749 2453 60433 2509
rect 60489 2453 60537 2509
rect 60593 2453 60641 2509
rect 60697 2453 62335 2509
rect 62391 2453 62975 2509
rect 63031 2453 63615 2509
rect 63671 2453 64255 2509
rect 64311 2453 64321 2509
rect 31260 2405 64321 2453
rect 5517 2298 5527 2354
rect 5583 2298 5631 2354
rect 5687 2298 6259 2354
rect 6315 2298 6899 2354
rect 6955 2298 7539 2354
rect 7595 2298 7605 2354
rect 5517 2288 5697 2298
rect 6249 2288 6325 2298
rect 6889 2288 6965 2298
rect 7529 2288 7605 2298
rect 17155 2348 18655 2358
rect 17155 2292 17165 2348
rect 17221 2292 18589 2348
rect 18645 2292 18655 2348
rect 17155 2282 18655 2292
rect 24851 2348 27776 2358
rect 24851 2292 24861 2348
rect 24917 2292 26285 2348
rect 26342 2292 27710 2348
rect 27766 2292 27776 2348
rect 31260 2349 31270 2405
rect 31326 2349 31374 2405
rect 31430 2349 31478 2405
rect 31534 2349 33247 2405
rect 33303 2349 33887 2405
rect 33943 2349 34527 2405
rect 34583 2349 35167 2405
rect 35223 2349 37381 2405
rect 37437 2349 38021 2405
rect 38077 2349 38661 2405
rect 38717 2349 39301 2405
rect 39357 2349 40997 2405
rect 41053 2349 41101 2405
rect 41157 2349 41205 2405
rect 41261 2349 42943 2405
rect 42999 2349 43583 2405
rect 43639 2349 44223 2405
rect 44279 2349 44863 2405
rect 44919 2349 47077 2405
rect 47133 2349 47717 2405
rect 47773 2349 48357 2405
rect 48413 2349 48997 2405
rect 49053 2349 50652 2405
rect 50708 2349 50756 2405
rect 50812 2349 50860 2405
rect 50916 2349 52639 2405
rect 52695 2349 53279 2405
rect 53335 2349 53919 2405
rect 53975 2349 54559 2405
rect 54615 2349 56773 2405
rect 56829 2349 57413 2405
rect 57469 2349 58053 2405
rect 58109 2349 58693 2405
rect 58749 2349 60433 2405
rect 60489 2349 60537 2405
rect 60593 2349 60641 2405
rect 60697 2349 62335 2405
rect 62391 2349 62975 2405
rect 63031 2349 63615 2405
rect 63671 2349 64255 2405
rect 64311 2349 64321 2405
rect 31260 2339 64321 2349
rect 24851 2282 27776 2292
rect 18819 2241 24687 2251
rect 10885 2218 11065 2228
rect 12314 2218 12390 2228
rect 13210 2218 13286 2228
rect 5245 2170 5425 2180
rect 6569 2170 6645 2180
rect 7209 2170 7285 2180
rect 5245 2114 5255 2170
rect 5311 2114 5359 2170
rect 5415 2114 6579 2170
rect 6635 2114 7219 2170
rect 7275 2114 7285 2170
rect 3384 2066 3460 2076
rect 4024 2066 4100 2076
rect 4664 2066 4740 2076
rect 5245 2066 7285 2114
rect 3384 2010 3394 2066
rect 3450 2010 4034 2066
rect 4090 2010 4674 2066
rect 4730 2010 5255 2066
rect 5311 2010 5359 2066
rect 5415 2010 6579 2066
rect 6635 2010 7219 2066
rect 7275 2010 7285 2066
rect 10885 2162 10895 2218
rect 10951 2162 10999 2218
rect 11055 2162 12324 2218
rect 12380 2162 13220 2218
rect 13276 2162 13286 2218
rect 10885 2114 13286 2162
rect 10885 2058 10895 2114
rect 10951 2058 10999 2114
rect 11055 2058 12324 2114
rect 12380 2058 13220 2114
rect 13276 2058 13286 2114
rect 10885 2048 11065 2058
rect 12314 2048 12390 2058
rect 13210 2048 13286 2058
rect 13498 2218 13574 2228
rect 14660 2218 14736 2228
rect 15300 2218 15376 2228
rect 15940 2218 16016 2228
rect 16879 2218 17059 2228
rect 13498 2162 13508 2218
rect 13564 2162 14670 2218
rect 14726 2162 15310 2218
rect 15366 2162 15950 2218
rect 16006 2162 16889 2218
rect 16945 2162 16993 2218
rect 17049 2162 17059 2218
rect 13498 2114 17059 2162
rect 13498 2058 13508 2114
rect 13564 2058 14670 2114
rect 14726 2058 15310 2114
rect 15366 2058 15950 2114
rect 16006 2058 16889 2114
rect 16945 2058 16993 2114
rect 17049 2058 17059 2114
rect 13498 2048 13574 2058
rect 14660 2048 14736 2058
rect 15300 2048 15376 2058
rect 15940 2048 16016 2058
rect 16879 2048 17059 2058
rect 18819 2185 21621 2241
rect 21677 2185 21725 2241
rect 21781 2185 21829 2241
rect 21885 2185 24687 2241
rect 18819 2137 24687 2185
rect 18819 2081 18829 2137
rect 18885 2081 19469 2137
rect 19525 2081 21621 2137
rect 21677 2081 21725 2137
rect 21781 2081 21829 2137
rect 21885 2081 23981 2137
rect 24037 2081 24621 2137
rect 24677 2081 24687 2137
rect 3384 1962 5425 2010
rect 6569 2000 6645 2010
rect 7209 2000 7285 2010
rect 18819 2033 24687 2081
rect 18819 1977 18829 2033
rect 18885 1977 19469 2033
rect 19525 1977 21621 2033
rect 21677 1977 21725 2033
rect 21781 1977 21829 2033
rect 21885 1977 23981 2033
rect 24037 1977 24621 2033
rect 24677 1977 24687 2033
rect 18819 1967 24687 1977
rect 27940 2241 31016 2251
rect 27940 2185 30742 2241
rect 30798 2185 30846 2241
rect 30902 2185 30950 2241
rect 31006 2185 31016 2241
rect 27940 2137 31016 2185
rect 27940 2081 27950 2137
rect 28006 2081 28590 2137
rect 28646 2081 30742 2137
rect 30798 2081 30846 2137
rect 30902 2081 30950 2137
rect 31006 2081 31016 2137
rect 27940 2033 31016 2081
rect 27940 1977 27950 2033
rect 28006 1977 28590 2033
rect 28646 1977 30742 2033
rect 30798 1977 30846 2033
rect 30902 1977 30950 2033
rect 31006 1977 31016 2033
rect 27940 1967 31016 1977
rect 31640 2219 64640 2229
rect 31640 2163 31650 2219
rect 31706 2163 31754 2219
rect 31810 2163 31858 2219
rect 31914 2163 40636 2219
rect 40692 2163 40740 2219
rect 40796 2163 40844 2219
rect 40900 2163 41356 2219
rect 41412 2163 41460 2219
rect 41516 2163 41564 2219
rect 41620 2163 50312 2219
rect 50368 2163 50416 2219
rect 50472 2163 50520 2219
rect 50576 2163 51044 2219
rect 51100 2163 51148 2219
rect 51204 2163 51252 2219
rect 51308 2163 60028 2219
rect 60084 2163 60132 2219
rect 60188 2163 60236 2219
rect 60292 2163 60792 2219
rect 60848 2163 60896 2219
rect 60952 2163 61000 2219
rect 61056 2163 64640 2219
rect 31640 2115 64640 2163
rect 31640 2059 31650 2115
rect 31706 2059 31754 2115
rect 31810 2059 31858 2115
rect 31914 2059 32926 2115
rect 32982 2059 33566 2115
rect 33622 2059 34846 2115
rect 34902 2059 35486 2115
rect 35542 2059 37062 2115
rect 37118 2059 37702 2115
rect 37758 2059 38982 2115
rect 39038 2059 39622 2115
rect 39678 2059 40636 2115
rect 40692 2059 40740 2115
rect 40796 2059 40844 2115
rect 40900 2059 41356 2115
rect 41412 2059 41460 2115
rect 41516 2059 41564 2115
rect 41620 2059 42622 2115
rect 42678 2059 43262 2115
rect 43318 2059 44542 2115
rect 44598 2059 45182 2115
rect 45238 2059 46758 2115
rect 46814 2059 47398 2115
rect 47454 2059 48678 2115
rect 48734 2059 49318 2115
rect 49374 2059 50312 2115
rect 50368 2059 50416 2115
rect 50472 2059 50520 2115
rect 50576 2059 51044 2115
rect 51100 2059 51148 2115
rect 51204 2059 51252 2115
rect 51308 2059 52318 2115
rect 52374 2059 52958 2115
rect 53014 2059 54238 2115
rect 54294 2059 54878 2115
rect 54934 2059 56454 2115
rect 56510 2059 57094 2115
rect 57150 2059 58374 2115
rect 58430 2059 59014 2115
rect 59070 2059 60028 2115
rect 60084 2059 60132 2115
rect 60188 2059 60236 2115
rect 60292 2059 60792 2115
rect 60848 2059 60896 2115
rect 60952 2059 61000 2115
rect 61056 2059 62014 2115
rect 62070 2059 62654 2115
rect 62710 2059 63934 2115
rect 63990 2059 64574 2115
rect 64630 2059 64640 2115
rect 31640 2011 64640 2059
rect 3384 1906 3394 1962
rect 3450 1906 4034 1962
rect 4090 1906 4674 1962
rect 4730 1906 5255 1962
rect 5311 1906 5359 1962
rect 5415 1906 5425 1962
rect 31640 1955 31650 2011
rect 31706 1955 31754 2011
rect 31810 1955 31858 2011
rect 31914 1955 32926 2011
rect 32982 1955 33566 2011
rect 33622 1955 34846 2011
rect 34902 1955 35486 2011
rect 35542 1955 37062 2011
rect 37118 1955 37702 2011
rect 37758 1955 38982 2011
rect 39038 1955 39622 2011
rect 39678 1955 40636 2011
rect 40692 1955 40740 2011
rect 40796 1955 40844 2011
rect 40900 1955 41356 2011
rect 41412 1955 41460 2011
rect 41516 1955 41564 2011
rect 41620 1955 42622 2011
rect 42678 1955 43262 2011
rect 43318 1955 44542 2011
rect 44598 1955 45182 2011
rect 45238 1955 46758 2011
rect 46814 1955 47398 2011
rect 47454 1955 48678 2011
rect 48734 1955 49318 2011
rect 49374 1955 50312 2011
rect 50368 1955 50416 2011
rect 50472 1955 50520 2011
rect 50576 1955 51044 2011
rect 51100 1955 51148 2011
rect 51204 1955 51252 2011
rect 51308 1955 52318 2011
rect 52374 1955 52958 2011
rect 53014 1955 54238 2011
rect 54294 1955 54878 2011
rect 54934 1955 56454 2011
rect 56510 1955 57094 2011
rect 57150 1955 58374 2011
rect 58430 1955 59014 2011
rect 59070 1955 60028 2011
rect 60084 1955 60132 2011
rect 60188 1955 60236 2011
rect 60292 1955 60792 2011
rect 60848 1955 60896 2011
rect 60952 1955 61000 2011
rect 61056 1955 62014 2011
rect 62070 1955 62654 2011
rect 62710 1955 63934 2011
rect 63990 1955 64574 2011
rect 64630 1955 64640 2011
rect 31640 1945 64640 1955
rect 3384 1896 3460 1906
rect 4024 1896 4100 1906
rect 4664 1896 4740 1906
rect 5245 1896 5425 1906
rect 18499 1847 25007 1857
rect 11153 1798 11333 1808
rect 11866 1798 11942 1808
rect 12762 1798 12838 1808
rect 13658 1798 13734 1808
rect 11153 1742 11163 1798
rect 11219 1742 11267 1798
rect 11323 1742 11876 1798
rect 11932 1742 12772 1798
rect 12828 1742 13668 1798
rect 13724 1742 13734 1798
rect 11153 1694 13734 1742
rect 5245 1639 5425 1649
rect 8484 1639 8560 1649
rect 9380 1639 9456 1649
rect 10276 1639 10352 1649
rect 5245 1583 5255 1639
rect 5311 1583 5359 1639
rect 5415 1583 8494 1639
rect 8550 1583 9390 1639
rect 9446 1583 10286 1639
rect 10342 1583 10352 1639
rect 11153 1638 11163 1694
rect 11219 1638 11267 1694
rect 11323 1638 11876 1694
rect 11932 1638 12772 1694
rect 12828 1638 13668 1694
rect 13724 1638 13734 1694
rect 11153 1628 11333 1638
rect 11866 1628 11942 1638
rect 12762 1628 12838 1638
rect 13658 1628 13734 1638
rect 14980 1798 15056 1808
rect 15620 1798 15696 1808
rect 16617 1798 16797 1808
rect 14980 1742 14990 1798
rect 15046 1742 15630 1798
rect 15686 1742 16627 1798
rect 16683 1742 16731 1798
rect 16787 1742 16797 1798
rect 14980 1694 16797 1742
rect 14980 1638 14990 1694
rect 15046 1638 15630 1694
rect 15686 1638 16627 1694
rect 16683 1638 16731 1694
rect 16787 1638 16797 1694
rect 14980 1628 15056 1638
rect 15620 1628 15696 1638
rect 16617 1628 16797 1638
rect 18499 1791 20972 1847
rect 21028 1791 21076 1847
rect 21132 1791 21180 1847
rect 21236 1791 22270 1847
rect 22326 1791 22374 1847
rect 22430 1791 22478 1847
rect 22534 1791 25007 1847
rect 18499 1743 25007 1791
rect 18499 1687 18509 1743
rect 18565 1687 19149 1743
rect 19205 1687 19789 1743
rect 19845 1687 20972 1743
rect 21028 1687 21076 1743
rect 21132 1687 21180 1743
rect 21236 1687 22270 1743
rect 22326 1687 22374 1743
rect 22430 1687 22478 1743
rect 22534 1687 23661 1743
rect 23717 1687 24301 1743
rect 24357 1687 24941 1743
rect 24997 1687 25007 1743
rect 18499 1639 25007 1687
rect 5245 1535 10352 1583
rect 18499 1583 18509 1639
rect 18565 1583 19149 1639
rect 19205 1583 19789 1639
rect 19845 1583 20972 1639
rect 21028 1583 21076 1639
rect 21132 1583 21180 1639
rect 21236 1583 22270 1639
rect 22326 1583 22374 1639
rect 22430 1583 22478 1639
rect 22534 1583 23661 1639
rect 23717 1583 24301 1639
rect 24357 1583 24941 1639
rect 24997 1583 25007 1639
rect 18499 1573 25007 1583
rect 27620 1847 30367 1857
rect 27620 1791 30093 1847
rect 30149 1791 30197 1847
rect 30253 1791 30301 1847
rect 30357 1791 30367 1847
rect 27620 1743 30367 1791
rect 27620 1687 27630 1743
rect 27686 1687 28270 1743
rect 28326 1687 28910 1743
rect 28966 1687 30093 1743
rect 30149 1687 30197 1743
rect 30253 1687 30301 1743
rect 30357 1687 30367 1743
rect 27620 1639 30367 1687
rect 27620 1583 27630 1639
rect 27686 1583 28270 1639
rect 28326 1583 28910 1639
rect 28966 1583 30093 1639
rect 30149 1583 30197 1639
rect 30253 1583 30301 1639
rect 30357 1583 30367 1639
rect 27620 1573 30367 1583
rect 5245 1479 5255 1535
rect 5311 1479 5359 1535
rect 5415 1479 8494 1535
rect 8550 1479 9390 1535
rect 9446 1479 10286 1535
rect 10342 1479 10352 1535
rect 5245 1469 5425 1479
rect 8484 1469 8560 1479
rect 9380 1469 9456 1479
rect 10276 1469 10352 1479
rect 31640 1553 64321 1563
rect 31640 1497 31650 1553
rect 31706 1497 31754 1553
rect 31810 1497 31858 1553
rect 31914 1497 40636 1553
rect 40692 1497 40740 1553
rect 40796 1497 40844 1553
rect 40900 1497 41356 1553
rect 41412 1497 41460 1553
rect 41516 1497 41564 1553
rect 41620 1497 50312 1553
rect 50368 1497 50416 1553
rect 50472 1497 50520 1553
rect 50576 1497 51044 1553
rect 51100 1497 51148 1553
rect 51204 1497 51252 1553
rect 51308 1497 60028 1553
rect 60084 1497 60132 1553
rect 60188 1497 60236 1553
rect 60292 1497 60792 1553
rect 60848 1497 60896 1553
rect 60952 1497 61000 1553
rect 61056 1497 64321 1553
rect 31640 1449 64321 1497
rect 31640 1393 31650 1449
rect 31706 1393 31754 1449
rect 31810 1393 31858 1449
rect 31914 1393 33247 1449
rect 33303 1393 33887 1449
rect 33943 1393 34527 1449
rect 34583 1393 35167 1449
rect 35223 1393 37381 1449
rect 37437 1393 38021 1449
rect 38077 1393 38661 1449
rect 38717 1393 39301 1449
rect 39357 1393 40636 1449
rect 40692 1393 40740 1449
rect 40796 1393 40844 1449
rect 40900 1393 41356 1449
rect 41412 1393 41460 1449
rect 41516 1393 41564 1449
rect 41620 1393 42943 1449
rect 42999 1393 43583 1449
rect 43639 1393 44223 1449
rect 44279 1393 44863 1449
rect 44919 1393 47077 1449
rect 47133 1393 47717 1449
rect 47773 1393 48357 1449
rect 48413 1393 48997 1449
rect 49053 1393 50312 1449
rect 50368 1393 50416 1449
rect 50472 1393 50520 1449
rect 50576 1393 51044 1449
rect 51100 1393 51148 1449
rect 51204 1393 51252 1449
rect 51308 1393 52639 1449
rect 52695 1393 53279 1449
rect 53335 1393 53919 1449
rect 53975 1393 54559 1449
rect 54615 1393 56773 1449
rect 56829 1393 57413 1449
rect 57469 1393 58053 1449
rect 58109 1393 58693 1449
rect 58749 1393 60028 1449
rect 60084 1393 60132 1449
rect 60188 1393 60236 1449
rect 60292 1393 60792 1449
rect 60848 1393 60896 1449
rect 60952 1393 61000 1449
rect 61056 1393 62335 1449
rect 62391 1393 62975 1449
rect 63031 1393 63615 1449
rect 63671 1393 64255 1449
rect 64311 1393 64321 1449
rect 31640 1345 64321 1393
rect 18819 1305 31544 1315
rect 5517 1268 5697 1278
rect 8932 1268 9008 1278
rect 9828 1268 9904 1278
rect 5517 1212 5527 1268
rect 5583 1212 5631 1268
rect 5687 1212 8942 1268
rect 8998 1212 9838 1268
rect 9894 1212 9904 1268
rect 2034 1168 2214 1178
rect 3544 1168 3620 1178
rect 2034 1112 2044 1168
rect 2100 1112 2148 1168
rect 2204 1112 3554 1168
rect 3610 1112 3620 1168
rect 2034 1064 3620 1112
rect 5517 1164 9904 1212
rect 5517 1108 5527 1164
rect 5583 1108 5631 1164
rect 5687 1108 8942 1164
rect 8998 1108 9838 1164
rect 9894 1108 9904 1164
rect 5517 1098 5697 1108
rect 8932 1098 9008 1108
rect 9828 1098 9904 1108
rect 10116 1268 10192 1278
rect 11153 1268 11333 1278
rect 10116 1212 10126 1268
rect 10182 1212 11163 1268
rect 11219 1212 11267 1268
rect 11323 1212 11333 1268
rect 10116 1164 11333 1212
rect 18819 1249 21621 1305
rect 21677 1249 21725 1305
rect 21781 1249 21829 1305
rect 21885 1249 30742 1305
rect 30798 1249 30846 1305
rect 30902 1249 30950 1305
rect 31006 1249 31544 1305
rect 31640 1289 31650 1345
rect 31706 1289 31754 1345
rect 31810 1289 31858 1345
rect 31914 1289 33247 1345
rect 33303 1289 33887 1345
rect 33943 1289 34527 1345
rect 34583 1289 35167 1345
rect 35223 1289 37381 1345
rect 37437 1289 38021 1345
rect 38077 1289 38661 1345
rect 38717 1289 39301 1345
rect 39357 1289 40636 1345
rect 40692 1289 40740 1345
rect 40796 1289 40844 1345
rect 40900 1289 41356 1345
rect 41412 1289 41460 1345
rect 41516 1289 41564 1345
rect 41620 1289 42943 1345
rect 42999 1289 43583 1345
rect 43639 1289 44223 1345
rect 44279 1289 44863 1345
rect 44919 1289 47077 1345
rect 47133 1289 47717 1345
rect 47773 1289 48357 1345
rect 48413 1289 48997 1345
rect 49053 1289 50312 1345
rect 50368 1289 50416 1345
rect 50472 1289 50520 1345
rect 50576 1289 51044 1345
rect 51100 1289 51148 1345
rect 51204 1289 51252 1345
rect 51308 1289 52639 1345
rect 52695 1289 53279 1345
rect 53335 1289 53919 1345
rect 53975 1289 54559 1345
rect 54615 1289 56773 1345
rect 56829 1289 57413 1345
rect 57469 1289 58053 1345
rect 58109 1289 58693 1345
rect 58749 1289 60028 1345
rect 60084 1289 60132 1345
rect 60188 1289 60236 1345
rect 60292 1289 60792 1345
rect 60848 1289 60896 1345
rect 60952 1289 61000 1345
rect 61056 1289 62335 1345
rect 62391 1289 62975 1345
rect 63031 1289 63615 1345
rect 63671 1289 64255 1345
rect 64311 1289 64321 1345
rect 31640 1279 64321 1289
rect 18819 1201 31544 1249
rect 12314 1164 12390 1174
rect 13210 1164 13286 1174
rect 10116 1108 10126 1164
rect 10182 1108 11163 1164
rect 11219 1108 11267 1164
rect 11323 1108 12324 1164
rect 12380 1108 13220 1164
rect 13276 1108 13286 1164
rect 10116 1098 10192 1108
rect 2034 1008 2044 1064
rect 2100 1008 2148 1064
rect 2204 1008 3554 1064
rect 3610 1008 3620 1064
rect 2034 998 2214 1008
rect 3544 998 3620 1008
rect 11153 1060 13286 1108
rect 11153 1004 11163 1060
rect 11219 1004 11267 1060
rect 11323 1004 12324 1060
rect 12380 1004 13220 1060
rect 13276 1004 13286 1060
rect 11153 994 11333 1004
rect 12314 994 12390 1004
rect 13210 994 13286 1004
rect 13498 1138 13574 1148
rect 14660 1138 14736 1148
rect 15300 1138 15376 1148
rect 15940 1138 16016 1148
rect 16617 1138 16797 1148
rect 13498 1082 13508 1138
rect 13564 1082 14670 1138
rect 14726 1082 15310 1138
rect 15366 1082 15950 1138
rect 16006 1082 16627 1138
rect 16683 1082 16731 1138
rect 16787 1082 16797 1138
rect 13498 1034 16797 1082
rect 13498 978 13508 1034
rect 13564 978 14670 1034
rect 14726 978 15310 1034
rect 15366 978 15950 1034
rect 16006 978 16627 1034
rect 16683 978 16731 1034
rect 16787 978 16797 1034
rect 18819 1145 18829 1201
rect 18885 1145 19469 1201
rect 19525 1145 21621 1201
rect 21677 1145 21725 1201
rect 21781 1145 21829 1201
rect 21885 1145 23981 1201
rect 24037 1145 24621 1201
rect 24677 1145 27950 1201
rect 28006 1145 28590 1201
rect 28646 1145 30742 1201
rect 30798 1145 30846 1201
rect 30902 1145 30950 1201
rect 31006 1169 31544 1201
rect 31006 1159 64640 1169
rect 31006 1145 31270 1159
rect 18819 1103 31270 1145
rect 31326 1103 31374 1159
rect 31430 1103 31478 1159
rect 31534 1103 40997 1159
rect 41053 1103 41101 1159
rect 41157 1103 41205 1159
rect 41261 1103 50652 1159
rect 50708 1103 50756 1159
rect 50812 1103 50860 1159
rect 50916 1103 60433 1159
rect 60489 1103 60537 1159
rect 60593 1103 60641 1159
rect 60697 1103 64640 1159
rect 18819 1097 64640 1103
rect 18819 1041 18829 1097
rect 18885 1041 19469 1097
rect 19525 1041 21621 1097
rect 21677 1041 21725 1097
rect 21781 1041 21829 1097
rect 21885 1041 23981 1097
rect 24037 1041 24621 1097
rect 24677 1041 27950 1097
rect 28006 1041 28590 1097
rect 28646 1041 30742 1097
rect 30798 1041 30846 1097
rect 30902 1041 30950 1097
rect 31006 1055 64640 1097
rect 31006 1041 31270 1055
rect 18819 1031 31270 1041
rect 13498 968 13574 978
rect 14660 968 14736 978
rect 15300 968 15376 978
rect 15940 968 16016 978
rect 16617 968 16797 978
rect 31260 999 31270 1031
rect 31326 999 31374 1055
rect 31430 999 31478 1055
rect 31534 999 32926 1055
rect 32982 999 33566 1055
rect 33622 999 34846 1055
rect 34902 999 35486 1055
rect 35542 999 37062 1055
rect 37118 999 37702 1055
rect 37758 999 38982 1055
rect 39038 999 39622 1055
rect 39678 999 40997 1055
rect 41053 999 41101 1055
rect 41157 999 41205 1055
rect 41261 999 42622 1055
rect 42678 999 43262 1055
rect 43318 999 44542 1055
rect 44598 999 45182 1055
rect 45238 999 46758 1055
rect 46814 999 47398 1055
rect 47454 999 48678 1055
rect 48734 999 49318 1055
rect 49374 999 50652 1055
rect 50708 999 50756 1055
rect 50812 999 50860 1055
rect 50916 999 52318 1055
rect 52374 999 52958 1055
rect 53014 999 54238 1055
rect 54294 999 54878 1055
rect 54934 999 56454 1055
rect 56510 999 57094 1055
rect 57150 999 58374 1055
rect 58430 999 59014 1055
rect 59070 999 60433 1055
rect 60489 999 60537 1055
rect 60593 999 60641 1055
rect 60697 999 62014 1055
rect 62070 999 62654 1055
rect 62710 999 63934 1055
rect 63990 999 64574 1055
rect 64630 999 64640 1055
rect 31260 951 64640 999
rect 18499 911 25007 921
rect 18499 855 20972 911
rect 21028 855 21076 911
rect 21132 855 21180 911
rect 21236 855 22270 911
rect 22326 855 22374 911
rect 22430 855 22478 911
rect 22534 855 25007 911
rect 5517 807 5697 817
rect 6569 807 6645 817
rect 7209 807 7285 817
rect 5517 751 5527 807
rect 5583 751 5631 807
rect 5687 751 6579 807
rect 6635 751 7219 807
rect 7275 751 7285 807
rect 5517 703 7285 751
rect 2395 655 2575 665
rect 3464 655 3540 665
rect 2395 599 2405 655
rect 2461 599 2509 655
rect 2565 599 3474 655
rect 3530 599 3540 655
rect 5517 647 5527 703
rect 5583 647 5631 703
rect 5687 647 6579 703
rect 6635 647 7219 703
rect 7275 647 7285 703
rect 5517 637 5697 647
rect 6569 637 6645 647
rect 7209 637 7285 647
rect 18499 807 25007 855
rect 18499 751 18509 807
rect 18565 751 19149 807
rect 19205 751 19789 807
rect 19845 751 20972 807
rect 21028 751 21076 807
rect 21132 751 21180 807
rect 21236 751 22270 807
rect 22326 751 22374 807
rect 22430 751 22478 807
rect 22534 751 23661 807
rect 23717 751 24301 807
rect 24357 751 24941 807
rect 24997 751 25007 807
rect 18499 703 25007 751
rect 18499 647 18509 703
rect 18565 647 19149 703
rect 19205 647 19789 703
rect 19845 647 20972 703
rect 21028 647 21076 703
rect 21132 647 21180 703
rect 21236 647 22270 703
rect 22326 647 22374 703
rect 22430 647 22478 703
rect 22534 647 23661 703
rect 23717 647 24301 703
rect 24357 647 24941 703
rect 24997 647 25007 703
rect 18499 637 25007 647
rect 27620 911 30367 921
rect 27620 855 30093 911
rect 30149 855 30197 911
rect 30253 855 30301 911
rect 30357 855 30367 911
rect 31260 895 31270 951
rect 31326 895 31374 951
rect 31430 895 31478 951
rect 31534 895 32926 951
rect 32982 895 33566 951
rect 33622 895 34846 951
rect 34902 895 35486 951
rect 35542 895 37062 951
rect 37118 895 37702 951
rect 37758 895 38982 951
rect 39038 895 39622 951
rect 39678 895 40997 951
rect 41053 895 41101 951
rect 41157 895 41205 951
rect 41261 895 42622 951
rect 42678 895 43262 951
rect 43318 895 44542 951
rect 44598 895 45182 951
rect 45238 895 46758 951
rect 46814 895 47398 951
rect 47454 895 48678 951
rect 48734 895 49318 951
rect 49374 895 50652 951
rect 50708 895 50756 951
rect 50812 895 50860 951
rect 50916 895 52318 951
rect 52374 895 52958 951
rect 53014 895 54238 951
rect 54294 895 54878 951
rect 54934 895 56454 951
rect 56510 895 57094 951
rect 57150 895 58374 951
rect 58430 895 59014 951
rect 59070 895 60433 951
rect 60489 895 60537 951
rect 60593 895 60641 951
rect 60697 895 62014 951
rect 62070 895 62654 951
rect 62710 895 63934 951
rect 63990 895 64574 951
rect 64630 895 64640 951
rect 31260 885 64640 895
rect 27620 807 30367 855
rect 27620 751 27630 807
rect 27686 751 28270 807
rect 28326 751 28910 807
rect 28966 751 30093 807
rect 30149 751 30197 807
rect 30253 751 30301 807
rect 30357 751 30367 807
rect 27620 703 30367 751
rect 27620 647 27630 703
rect 27686 647 28270 703
rect 28326 647 28910 703
rect 28966 647 30093 703
rect 30149 647 30197 703
rect 30253 647 30301 703
rect 30357 647 30367 703
rect 27620 637 30367 647
rect 2395 551 3540 599
rect 2395 495 2405 551
rect 2461 495 2509 551
rect 2565 495 3474 551
rect 3530 495 3540 551
rect 2395 485 2575 495
rect 3464 483 3540 495
rect 10116 606 10192 616
rect 10885 606 11065 616
rect 10116 550 10126 606
rect 10182 550 10895 606
rect 10951 550 10999 606
rect 11055 550 11065 606
rect 10116 502 11065 550
rect 10116 446 10126 502
rect 10182 446 10895 502
rect 10951 446 10999 502
rect 11055 446 11065 502
rect 31640 493 64321 503
rect 10116 436 10192 446
rect 10885 436 11065 446
rect 17355 476 18655 486
rect 17355 420 17365 476
rect 17421 420 18589 476
rect 18645 420 18655 476
rect 5245 406 5425 416
rect 6249 406 6325 416
rect 6889 406 6965 416
rect 7529 406 7605 416
rect 8932 406 9008 416
rect 9828 406 9904 416
rect 17355 410 18655 420
rect 24851 476 27776 486
rect 24851 420 24861 476
rect 24917 420 26085 476
rect 26141 420 26486 476
rect 26542 420 27710 476
rect 27766 420 27776 476
rect 24851 410 27776 420
rect 31640 437 31650 493
rect 31706 437 31754 493
rect 31810 437 31858 493
rect 31914 437 40636 493
rect 40692 437 40740 493
rect 40796 437 40844 493
rect 40900 437 41356 493
rect 41412 437 41460 493
rect 41516 437 41564 493
rect 41620 437 50312 493
rect 50368 437 50416 493
rect 50472 437 50520 493
rect 50576 437 51044 493
rect 51100 437 51148 493
rect 51204 437 51252 493
rect 51308 437 60028 493
rect 60084 437 60132 493
rect 60188 437 60236 493
rect 60292 437 60792 493
rect 60848 437 60896 493
rect 60952 437 61000 493
rect 61056 437 64321 493
rect 5245 350 5255 406
rect 5311 350 5359 406
rect 5415 350 6259 406
rect 6315 350 6899 406
rect 6955 350 7539 406
rect 7595 350 8942 406
rect 8998 350 9838 406
rect 9894 350 9904 406
rect 31640 389 64321 437
rect 2138 302 2214 312
rect 3544 302 3620 312
rect 2138 246 2148 302
rect 2204 246 3554 302
rect 3610 246 3620 302
rect 2138 198 3620 246
rect 2138 142 2148 198
rect 2204 142 3554 198
rect 3610 142 3620 198
rect 2138 132 2214 142
rect 3544 132 3620 142
rect 3704 302 3780 312
rect 4345 302 4421 312
rect 5245 302 9904 350
rect 3704 246 3714 302
rect 3770 246 4355 302
rect 4411 246 5255 302
rect 5311 246 5359 302
rect 5415 246 6259 302
rect 6315 246 6899 302
rect 6955 246 7539 302
rect 7595 246 8942 302
rect 8998 246 9838 302
rect 9894 246 9904 302
rect 3704 198 5425 246
rect 6249 236 6325 246
rect 6889 236 6965 246
rect 7529 236 7605 246
rect 8932 236 9008 246
rect 9828 236 9904 246
rect 18819 369 24687 379
rect 18819 313 20972 369
rect 21028 313 21076 369
rect 21132 313 21180 369
rect 21236 313 22270 369
rect 22326 313 22374 369
rect 22430 313 22478 369
rect 22534 313 24687 369
rect 18819 265 24687 313
rect 3704 142 3714 198
rect 3770 142 4355 198
rect 4411 142 5255 198
rect 5311 142 5359 198
rect 5415 142 5425 198
rect 3704 132 3780 142
rect 4345 132 4421 142
rect 5245 132 5425 142
rect 18819 209 18829 265
rect 18885 209 19469 265
rect 19525 209 20972 265
rect 21028 209 21076 265
rect 21132 209 21180 265
rect 21236 209 22270 265
rect 22326 209 22374 265
rect 22430 209 22478 265
rect 22534 209 23981 265
rect 24037 209 24621 265
rect 24677 209 24687 265
rect 18819 161 24687 209
rect 10885 118 11065 128
rect 11866 118 11942 128
rect 12762 118 12838 128
rect 13658 118 13734 128
rect 10885 62 10895 118
rect 10951 62 10999 118
rect 11055 62 11876 118
rect 11932 62 12772 118
rect 12828 62 13668 118
rect 13724 62 13734 118
rect 18819 105 18829 161
rect 18885 105 19469 161
rect 19525 105 20972 161
rect 21028 105 21076 161
rect 21132 105 21180 161
rect 21236 105 22270 161
rect 22326 105 22374 161
rect 22430 105 22478 161
rect 22534 105 23981 161
rect 24037 105 24621 161
rect 24677 105 24687 161
rect 18819 95 24687 105
rect 27940 369 30367 379
rect 27940 313 30093 369
rect 30149 313 30197 369
rect 30253 313 30301 369
rect 30357 313 30367 369
rect 27940 265 30367 313
rect 27940 209 27950 265
rect 28006 209 28590 265
rect 28646 209 30093 265
rect 30149 209 30197 265
rect 30253 209 30301 265
rect 30357 209 30367 265
rect 31640 333 31650 389
rect 31706 333 31754 389
rect 31810 333 31858 389
rect 31914 333 33247 389
rect 33303 333 33887 389
rect 33943 333 34527 389
rect 34583 333 35167 389
rect 35223 333 37381 389
rect 37437 333 38021 389
rect 38077 333 38661 389
rect 38717 333 39301 389
rect 39357 333 40636 389
rect 40692 333 40740 389
rect 40796 333 40844 389
rect 40900 333 41356 389
rect 41412 333 41460 389
rect 41516 333 41564 389
rect 41620 333 42943 389
rect 42999 333 43583 389
rect 43639 333 44223 389
rect 44279 333 44863 389
rect 44919 333 47077 389
rect 47133 333 47717 389
rect 47773 333 48357 389
rect 48413 333 48997 389
rect 49053 333 50312 389
rect 50368 333 50416 389
rect 50472 333 50520 389
rect 50576 333 51044 389
rect 51100 333 51148 389
rect 51204 333 51252 389
rect 51308 333 52639 389
rect 52695 333 53279 389
rect 53335 333 53919 389
rect 53975 333 54559 389
rect 54615 333 56773 389
rect 56829 333 57413 389
rect 57469 333 58053 389
rect 58109 333 58693 389
rect 58749 333 60028 389
rect 60084 333 60132 389
rect 60188 333 60236 389
rect 60292 333 60792 389
rect 60848 333 60896 389
rect 60952 333 61000 389
rect 61056 333 62335 389
rect 62391 333 62975 389
rect 63031 333 63615 389
rect 63671 333 64255 389
rect 64311 333 64321 389
rect 31640 285 64321 333
rect 31640 229 31650 285
rect 31706 229 31754 285
rect 31810 229 31858 285
rect 31914 229 33247 285
rect 33303 229 33887 285
rect 33943 229 34527 285
rect 34583 229 35167 285
rect 35223 229 37381 285
rect 37437 229 38021 285
rect 38077 229 38661 285
rect 38717 229 39301 285
rect 39357 229 40636 285
rect 40692 229 40740 285
rect 40796 229 40844 285
rect 40900 229 41356 285
rect 41412 229 41460 285
rect 41516 229 41564 285
rect 41620 229 42943 285
rect 42999 229 43583 285
rect 43639 229 44223 285
rect 44279 229 44863 285
rect 44919 229 47077 285
rect 47133 229 47717 285
rect 47773 229 48357 285
rect 48413 229 48997 285
rect 49053 229 50312 285
rect 50368 229 50416 285
rect 50472 229 50520 285
rect 50576 229 51044 285
rect 51100 229 51148 285
rect 51204 229 51252 285
rect 51308 229 52639 285
rect 52695 229 53279 285
rect 53335 229 53919 285
rect 53975 229 54559 285
rect 54615 229 56773 285
rect 56829 229 57413 285
rect 57469 229 58053 285
rect 58109 229 58693 285
rect 58749 229 60028 285
rect 60084 229 60132 285
rect 60188 229 60236 285
rect 60292 229 60792 285
rect 60848 229 60896 285
rect 60952 229 61000 285
rect 61056 229 62335 285
rect 62391 229 62975 285
rect 63031 229 63615 285
rect 63671 229 64255 285
rect 64311 229 64321 285
rect 31640 219 64321 229
rect 27940 161 30367 209
rect 27940 105 27950 161
rect 28006 105 28590 161
rect 28646 105 30093 161
rect 30149 105 30197 161
rect 30253 105 30301 161
rect 30357 105 30367 161
rect 27940 95 30367 105
rect 31260 99 64640 109
rect 10885 14 13734 62
rect 10885 -42 10895 14
rect 10951 -42 10999 14
rect 11055 -42 11876 14
rect 11932 -42 12772 14
rect 12828 -42 13668 14
rect 13724 -42 13734 14
rect 31260 43 31270 99
rect 31326 43 31374 99
rect 31430 43 31478 99
rect 31534 43 40997 99
rect 41053 43 41101 99
rect 41157 43 41205 99
rect 41261 43 50652 99
rect 50708 43 50756 99
rect 50812 43 50860 99
rect 50916 43 60433 99
rect 60489 43 60537 99
rect 60593 43 60641 99
rect 60697 43 64640 99
rect 31260 -5 64640 43
rect 31260 -15 31270 -5
rect 10885 -52 11065 -42
rect 11866 -52 11942 -42
rect 12762 -52 12838 -42
rect 13658 -52 13734 -42
rect 18499 -25 31270 -15
rect 18499 -81 21621 -25
rect 21677 -81 21725 -25
rect 21781 -81 21829 -25
rect 21885 -81 30742 -25
rect 30798 -81 30846 -25
rect 30902 -81 30950 -25
rect 31006 -61 31270 -25
rect 31326 -61 31374 -5
rect 31430 -61 31478 -5
rect 31534 -61 32926 -5
rect 32982 -61 33566 -5
rect 33622 -61 34846 -5
rect 34902 -61 35486 -5
rect 35542 -61 37062 -5
rect 37118 -61 37702 -5
rect 37758 -61 38982 -5
rect 39038 -61 39622 -5
rect 39678 -61 40997 -5
rect 41053 -61 41101 -5
rect 41157 -61 41205 -5
rect 41261 -61 42622 -5
rect 42678 -61 43262 -5
rect 43318 -61 44542 -5
rect 44598 -61 45182 -5
rect 45238 -61 46758 -5
rect 46814 -61 47398 -5
rect 47454 -61 48678 -5
rect 48734 -61 49318 -5
rect 49374 -61 50652 -5
rect 50708 -61 50756 -5
rect 50812 -61 50860 -5
rect 50916 -61 52318 -5
rect 52374 -61 52958 -5
rect 53014 -61 54238 -5
rect 54294 -61 54878 -5
rect 54934 -61 56454 -5
rect 56510 -61 57094 -5
rect 57150 -61 58374 -5
rect 58430 -61 59014 -5
rect 59070 -61 60433 -5
rect 60489 -61 60537 -5
rect 60593 -61 60641 -5
rect 60697 -61 62014 -5
rect 62070 -61 62654 -5
rect 62710 -61 63934 -5
rect 63990 -61 64574 -5
rect 64630 -61 64640 -5
rect 31006 -81 64640 -61
rect 18499 -109 64640 -81
rect 18499 -129 31270 -109
rect 3384 -194 3460 -184
rect 4024 -194 4100 -184
rect 4664 -194 4740 -184
rect 5517 -194 5697 -184
rect 6249 -194 6325 -184
rect 6889 -194 6965 -184
rect 7529 -194 7605 -184
rect 8484 -194 8560 -184
rect 9380 -194 9456 -184
rect 10276 -194 10352 -184
rect 3384 -250 3394 -194
rect 3450 -250 4034 -194
rect 4090 -250 4674 -194
rect 4730 -250 5527 -194
rect 5583 -250 5631 -194
rect 5687 -250 6259 -194
rect 6315 -250 6899 -194
rect 6955 -250 7539 -194
rect 7595 -250 8494 -194
rect 8550 -250 9390 -194
rect 9446 -250 10286 -194
rect 10342 -250 10352 -194
rect 3384 -298 10352 -250
rect 18499 -185 18509 -129
rect 18565 -185 19149 -129
rect 19205 -185 19789 -129
rect 19845 -185 21621 -129
rect 21677 -185 21725 -129
rect 21781 -185 21829 -129
rect 21885 -185 23661 -129
rect 23717 -185 24301 -129
rect 24357 -185 24941 -129
rect 24997 -185 27630 -129
rect 27686 -185 28270 -129
rect 28326 -185 28910 -129
rect 28966 -185 30742 -129
rect 30798 -185 30846 -129
rect 30902 -185 30950 -129
rect 31006 -165 31270 -129
rect 31326 -165 31374 -109
rect 31430 -165 31478 -109
rect 31534 -165 32926 -109
rect 32982 -165 33566 -109
rect 33622 -165 34846 -109
rect 34902 -165 35486 -109
rect 35542 -165 37062 -109
rect 37118 -165 37702 -109
rect 37758 -165 38982 -109
rect 39038 -165 39622 -109
rect 39678 -165 40997 -109
rect 41053 -165 41101 -109
rect 41157 -165 41205 -109
rect 41261 -165 42622 -109
rect 42678 -165 43262 -109
rect 43318 -165 44542 -109
rect 44598 -165 45182 -109
rect 45238 -165 46758 -109
rect 46814 -165 47398 -109
rect 47454 -165 48678 -109
rect 48734 -165 49318 -109
rect 49374 -165 50652 -109
rect 50708 -165 50756 -109
rect 50812 -165 50860 -109
rect 50916 -165 52318 -109
rect 52374 -165 52958 -109
rect 53014 -165 54238 -109
rect 54294 -165 54878 -109
rect 54934 -165 56454 -109
rect 56510 -165 57094 -109
rect 57150 -165 58374 -109
rect 58430 -165 59014 -109
rect 59070 -165 60433 -109
rect 60489 -165 60537 -109
rect 60593 -165 60641 -109
rect 60697 -165 62014 -109
rect 62070 -165 62654 -109
rect 62710 -165 63934 -109
rect 63990 -165 64574 -109
rect 64630 -165 64640 -109
rect 31006 -175 64640 -165
rect 31006 -185 31544 -175
rect 18499 -233 31544 -185
rect 3384 -354 3394 -298
rect 3450 -354 4034 -298
rect 4090 -354 4674 -298
rect 4730 -354 5527 -298
rect 5583 -354 5631 -298
rect 5687 -354 6259 -298
rect 6315 -354 6899 -298
rect 6955 -354 7539 -298
rect 7595 -354 8494 -298
rect 8550 -354 9390 -298
rect 9446 -354 10286 -298
rect 10342 -354 10352 -298
rect 3384 -364 3460 -354
rect 4024 -364 4100 -354
rect 4664 -364 4740 -354
rect 5517 -364 5697 -354
rect 6249 -364 6325 -354
rect 6889 -364 6965 -354
rect 7529 -364 7605 -354
rect 8484 -364 8560 -354
rect 9380 -364 9456 -354
rect 10276 -364 10352 -354
rect 13370 -282 13446 -272
rect 14980 -282 15056 -272
rect 15620 -282 15696 -272
rect 16879 -282 17059 -272
rect 13370 -338 13380 -282
rect 13436 -338 14990 -282
rect 15046 -338 15630 -282
rect 15686 -338 16889 -282
rect 16945 -338 16993 -282
rect 17049 -338 17059 -282
rect 18499 -289 18509 -233
rect 18565 -289 19149 -233
rect 19205 -289 19789 -233
rect 19845 -289 21621 -233
rect 21677 -289 21725 -233
rect 21781 -289 21829 -233
rect 21885 -289 23661 -233
rect 23717 -289 24301 -233
rect 24357 -289 24941 -233
rect 24997 -289 27630 -233
rect 27686 -289 28270 -233
rect 28326 -289 28910 -233
rect 28966 -289 30742 -233
rect 30798 -289 30846 -233
rect 30902 -289 30950 -233
rect 31006 -289 31544 -233
rect 18499 -299 31544 -289
rect 13370 -386 17059 -338
rect 13370 -442 13380 -386
rect 13436 -442 14990 -386
rect 15046 -442 15630 -386
rect 15686 -442 16889 -386
rect 16945 -442 16993 -386
rect 17049 -442 17059 -386
rect 9988 -452 10064 -442
rect 11153 -452 11333 -442
rect 13370 -452 13446 -442
rect 14980 -452 15056 -442
rect 15620 -452 15696 -442
rect 16879 -452 17059 -442
rect 2675 -475 2855 -465
rect 3464 -475 3540 -465
rect 2675 -531 2685 -475
rect 2741 -531 2789 -475
rect 2845 -531 3474 -475
rect 3530 -531 3540 -475
rect 2675 -579 3540 -531
rect 2675 -635 2685 -579
rect 2741 -635 2789 -579
rect 2845 -635 3474 -579
rect 3530 -635 3540 -579
rect 2675 -645 2855 -635
rect 3464 -645 3540 -635
rect 5245 -467 5425 -457
rect 6569 -467 6645 -457
rect 7209 -467 7285 -457
rect 5245 -523 5255 -467
rect 5311 -523 5359 -467
rect 5415 -523 6579 -467
rect 6635 -523 7219 -467
rect 7275 -523 7285 -467
rect 5245 -571 7285 -523
rect 5245 -627 5255 -571
rect 5311 -627 5359 -571
rect 5415 -627 6579 -571
rect 6635 -627 7219 -571
rect 7275 -627 7285 -571
rect 9988 -508 9998 -452
rect 10054 -508 11163 -452
rect 11219 -508 11267 -452
rect 11323 -508 11333 -452
rect 9988 -556 11333 -508
rect 17155 -460 18655 -450
rect 17155 -516 17165 -460
rect 17221 -516 18589 -460
rect 18645 -516 18655 -460
rect 17155 -526 18655 -516
rect 24851 -460 27776 -450
rect 24851 -516 24861 -460
rect 24917 -516 26285 -460
rect 26342 -516 27710 -460
rect 27766 -516 27776 -460
rect 24851 -526 27776 -516
rect 9988 -612 9998 -556
rect 10054 -612 11163 -556
rect 11219 -612 11267 -556
rect 11323 -612 11333 -556
rect 18819 -567 24687 -557
rect 9988 -622 10064 -612
rect 11153 -622 11333 -612
rect 11532 -592 11712 -582
rect 11902 -592 11978 -582
rect 5245 -637 5425 -627
rect 6569 -637 6645 -627
rect 7209 -637 7285 -627
rect 11532 -648 11542 -592
rect 11598 -648 11646 -592
rect 11702 -648 11912 -592
rect 11968 -648 11978 -592
rect 7503 -691 7579 -681
rect 7789 -691 7969 -681
rect 7503 -747 7513 -691
rect 7569 -747 7799 -691
rect 7855 -747 7903 -691
rect 7959 -747 7969 -691
rect 7503 -795 7969 -747
rect 3704 -828 3780 -818
rect 4345 -828 4421 -818
rect 5517 -828 5697 -818
rect 3704 -884 3714 -828
rect 3770 -884 4355 -828
rect 4411 -884 5527 -828
rect 5583 -884 5631 -828
rect 5687 -884 5697 -828
rect 7503 -851 7513 -795
rect 7569 -851 7799 -795
rect 7855 -851 7903 -795
rect 7959 -851 7969 -795
rect 7503 -861 7579 -851
rect 7789 -861 7969 -851
rect 10236 -702 10312 -692
rect 10432 -702 10612 -692
rect 10236 -758 10246 -702
rect 10302 -758 10442 -702
rect 10498 -758 10546 -702
rect 10602 -758 10612 -702
rect 10236 -806 10612 -758
rect 11532 -696 11978 -648
rect 11532 -752 11542 -696
rect 11598 -752 11646 -696
rect 11702 -752 11912 -696
rect 11968 -752 11978 -696
rect 11532 -762 11712 -752
rect 11902 -762 11978 -752
rect 14200 -587 14380 -577
rect 14688 -587 14764 -577
rect 14200 -643 14210 -587
rect 14266 -643 14314 -587
rect 14370 -643 14698 -587
rect 14754 -643 14764 -587
rect 14200 -691 14764 -643
rect 14200 -747 14210 -691
rect 14266 -747 14314 -691
rect 14370 -747 14698 -691
rect 14754 -747 14764 -691
rect 14200 -757 14380 -747
rect 14688 -757 14764 -747
rect 18819 -623 21621 -567
rect 21677 -623 21725 -567
rect 21781 -623 21829 -567
rect 21885 -623 24687 -567
rect 18819 -671 24687 -623
rect 18819 -727 18829 -671
rect 18885 -727 19469 -671
rect 19525 -727 21621 -671
rect 21677 -727 21725 -671
rect 21781 -727 21829 -671
rect 21885 -727 23981 -671
rect 24037 -727 24621 -671
rect 24677 -727 24687 -671
rect 10236 -862 10246 -806
rect 10302 -862 10442 -806
rect 10498 -862 10546 -806
rect 10602 -862 10612 -806
rect 18819 -775 24687 -727
rect 18819 -831 18829 -775
rect 18885 -831 19469 -775
rect 19525 -831 21621 -775
rect 21677 -831 21725 -775
rect 21781 -831 21829 -775
rect 21885 -831 23981 -775
rect 24037 -831 24621 -775
rect 24677 -831 24687 -775
rect 18819 -841 24687 -831
rect 27940 -567 64321 -557
rect 27940 -623 30742 -567
rect 30798 -623 30846 -567
rect 30902 -623 30950 -567
rect 31006 -623 31270 -567
rect 31326 -623 31374 -567
rect 31430 -623 31478 -567
rect 31534 -623 40997 -567
rect 41053 -623 41101 -567
rect 41157 -623 41205 -567
rect 41261 -623 50652 -567
rect 50708 -623 50756 -567
rect 50812 -623 50860 -567
rect 50916 -623 60433 -567
rect 60489 -623 60537 -567
rect 60593 -623 60641 -567
rect 60697 -623 64321 -567
rect 27940 -671 64321 -623
rect 27940 -727 27950 -671
rect 28006 -727 28590 -671
rect 28646 -727 30742 -671
rect 30798 -727 30846 -671
rect 30902 -727 30950 -671
rect 31006 -727 31270 -671
rect 31326 -727 31374 -671
rect 31430 -727 31478 -671
rect 31534 -727 33247 -671
rect 33303 -727 33887 -671
rect 33943 -727 34527 -671
rect 34583 -727 35167 -671
rect 35223 -727 37381 -671
rect 37437 -727 38021 -671
rect 38077 -727 38661 -671
rect 38717 -727 39301 -671
rect 39357 -727 40997 -671
rect 41053 -727 41101 -671
rect 41157 -727 41205 -671
rect 41261 -727 42943 -671
rect 42999 -727 43583 -671
rect 43639 -727 44223 -671
rect 44279 -727 44863 -671
rect 44919 -727 47077 -671
rect 47133 -727 47717 -671
rect 47773 -727 48357 -671
rect 48413 -727 48997 -671
rect 49053 -727 50652 -671
rect 50708 -727 50756 -671
rect 50812 -727 50860 -671
rect 50916 -727 52639 -671
rect 52695 -727 53279 -671
rect 53335 -727 53919 -671
rect 53975 -727 54559 -671
rect 54615 -727 56773 -671
rect 56829 -727 57413 -671
rect 57469 -727 58053 -671
rect 58109 -727 58693 -671
rect 58749 -727 60433 -671
rect 60489 -727 60537 -671
rect 60593 -727 60641 -671
rect 60697 -727 62335 -671
rect 62391 -727 62975 -671
rect 63031 -727 63615 -671
rect 63671 -727 64255 -671
rect 64311 -727 64321 -671
rect 27940 -775 64321 -727
rect 27940 -831 27950 -775
rect 28006 -831 28590 -775
rect 28646 -831 30742 -775
rect 30798 -831 30846 -775
rect 30902 -831 30950 -775
rect 31006 -831 31270 -775
rect 31326 -831 31374 -775
rect 31430 -831 31478 -775
rect 31534 -831 33247 -775
rect 33303 -831 33887 -775
rect 33943 -831 34527 -775
rect 34583 -831 35167 -775
rect 35223 -831 37381 -775
rect 37437 -831 38021 -775
rect 38077 -831 38661 -775
rect 38717 -831 39301 -775
rect 39357 -831 40997 -775
rect 41053 -831 41101 -775
rect 41157 -831 41205 -775
rect 41261 -831 42943 -775
rect 42999 -831 43583 -775
rect 43639 -831 44223 -775
rect 44279 -831 44863 -775
rect 44919 -831 47077 -775
rect 47133 -831 47717 -775
rect 47773 -831 48357 -775
rect 48413 -831 48997 -775
rect 49053 -831 50652 -775
rect 50708 -831 50756 -775
rect 50812 -831 50860 -775
rect 50916 -831 52639 -775
rect 52695 -831 53279 -775
rect 53335 -831 53919 -775
rect 53975 -831 54559 -775
rect 54615 -831 56773 -775
rect 56829 -831 57413 -775
rect 57469 -831 58053 -775
rect 58109 -831 58693 -775
rect 58749 -831 60433 -775
rect 60489 -831 60537 -775
rect 60593 -831 60641 -775
rect 60697 -831 62335 -775
rect 62391 -831 62975 -775
rect 63031 -831 63615 -775
rect 63671 -831 64255 -775
rect 64311 -831 64321 -775
rect 27940 -841 64321 -831
rect 10236 -872 10312 -862
rect 10432 -872 10612 -862
rect 3704 -932 5697 -884
rect 6569 -932 6645 -922
rect 7209 -932 7285 -922
rect 8932 -932 9008 -922
rect 9828 -932 9904 -922
rect 3704 -988 3714 -932
rect 3770 -988 4355 -932
rect 4411 -988 5527 -932
rect 5583 -988 5631 -932
rect 5687 -988 6579 -932
rect 6635 -988 7219 -932
rect 7275 -988 8942 -932
rect 8998 -988 9838 -932
rect 9894 -988 9904 -932
rect 3704 -998 3780 -988
rect 4345 -998 4421 -988
rect 2138 -1028 2214 -1018
rect 3544 -1028 3620 -1018
rect 2138 -1084 2148 -1028
rect 2204 -1084 3554 -1028
rect 3610 -1084 3620 -1028
rect 2138 -1132 3620 -1084
rect 5517 -1036 9904 -988
rect 5517 -1092 5527 -1036
rect 5583 -1092 5631 -1036
rect 5687 -1092 6579 -1036
rect 6635 -1092 7219 -1036
rect 7275 -1092 8942 -1036
rect 8998 -1092 9838 -1036
rect 9894 -1092 9904 -1036
rect 5517 -1102 5697 -1092
rect 6569 -1102 6645 -1092
rect 7209 -1102 7285 -1092
rect 8932 -1102 9008 -1092
rect 9828 -1102 9904 -1092
rect 9988 -932 10064 -922
rect 10885 -932 11065 -922
rect 12314 -932 12390 -922
rect 13210 -932 13286 -922
rect 9988 -988 9998 -932
rect 10054 -988 10895 -932
rect 10951 -988 10999 -932
rect 11055 -988 12324 -932
rect 12380 -988 13220 -932
rect 13276 -988 13286 -932
rect 9988 -1036 13286 -988
rect 9988 -1092 9998 -1036
rect 10054 -1092 10895 -1036
rect 10951 -1092 10999 -1036
rect 11055 -1092 12324 -1036
rect 12380 -1092 13220 -1036
rect 13276 -1092 13286 -1036
rect 9988 -1102 10064 -1092
rect 10885 -1102 11065 -1092
rect 12314 -1102 12390 -1092
rect 13210 -1102 13286 -1092
rect 13370 -932 13446 -922
rect 14980 -932 15056 -922
rect 15620 -932 15696 -922
rect 16617 -932 16797 -922
rect 13370 -988 13380 -932
rect 13436 -988 14990 -932
rect 15046 -988 15630 -932
rect 15686 -988 16627 -932
rect 16683 -988 16731 -932
rect 16787 -988 16797 -932
rect 13370 -1036 16797 -988
rect 13370 -1092 13380 -1036
rect 13436 -1092 14990 -1036
rect 15046 -1092 15630 -1036
rect 15686 -1092 16627 -1036
rect 16683 -1092 16731 -1036
rect 16787 -1092 16797 -1036
rect 13370 -1102 13446 -1092
rect 14980 -1102 15056 -1092
rect 15620 -1102 15696 -1092
rect 16617 -1102 16797 -1092
rect 18499 -961 64640 -951
rect 18499 -1017 20972 -961
rect 21028 -1017 21076 -961
rect 21132 -1017 21180 -961
rect 21236 -1017 22270 -961
rect 22326 -1017 22374 -961
rect 22430 -1017 22478 -961
rect 22534 -1017 30093 -961
rect 30149 -1017 30197 -961
rect 30253 -1017 30301 -961
rect 30357 -1017 31650 -961
rect 31706 -1017 31754 -961
rect 31810 -1017 31858 -961
rect 31914 -1017 40636 -961
rect 40692 -1017 40740 -961
rect 40796 -1017 40844 -961
rect 40900 -1017 41356 -961
rect 41412 -1017 41460 -961
rect 41516 -1017 41564 -961
rect 41620 -1017 50312 -961
rect 50368 -1017 50416 -961
rect 50472 -1017 50520 -961
rect 50576 -1017 51044 -961
rect 51100 -1017 51148 -961
rect 51204 -1017 51252 -961
rect 51308 -1017 60028 -961
rect 60084 -1017 60132 -961
rect 60188 -1017 60236 -961
rect 60292 -1017 60792 -961
rect 60848 -1017 60896 -961
rect 60952 -1017 61000 -961
rect 61056 -1017 64640 -961
rect 18499 -1065 64640 -1017
rect 2138 -1188 2148 -1132
rect 2204 -1188 3554 -1132
rect 3610 -1188 3620 -1132
rect 2138 -1198 2214 -1188
rect 3544 -1198 3620 -1188
rect 18499 -1121 18509 -1065
rect 18565 -1121 19149 -1065
rect 19205 -1121 19789 -1065
rect 19845 -1121 20972 -1065
rect 21028 -1121 21076 -1065
rect 21132 -1121 21180 -1065
rect 21236 -1121 22270 -1065
rect 22326 -1121 22374 -1065
rect 22430 -1121 22478 -1065
rect 22534 -1121 23661 -1065
rect 23717 -1121 24301 -1065
rect 24357 -1121 24941 -1065
rect 24997 -1121 27630 -1065
rect 27686 -1121 28270 -1065
rect 28326 -1121 28910 -1065
rect 28966 -1121 30093 -1065
rect 30149 -1121 30197 -1065
rect 30253 -1121 30301 -1065
rect 30357 -1121 31650 -1065
rect 31706 -1121 31754 -1065
rect 31810 -1121 31858 -1065
rect 31914 -1121 32926 -1065
rect 32982 -1121 33566 -1065
rect 33622 -1121 34846 -1065
rect 34902 -1121 35486 -1065
rect 35542 -1121 37062 -1065
rect 37118 -1121 37702 -1065
rect 37758 -1121 38982 -1065
rect 39038 -1121 39622 -1065
rect 39678 -1121 40636 -1065
rect 40692 -1121 40740 -1065
rect 40796 -1121 40844 -1065
rect 40900 -1121 41356 -1065
rect 41412 -1121 41460 -1065
rect 41516 -1121 41564 -1065
rect 41620 -1121 42622 -1065
rect 42678 -1121 43262 -1065
rect 43318 -1121 44542 -1065
rect 44598 -1121 45182 -1065
rect 45238 -1121 46758 -1065
rect 46814 -1121 47398 -1065
rect 47454 -1121 48678 -1065
rect 48734 -1121 49318 -1065
rect 49374 -1121 50312 -1065
rect 50368 -1121 50416 -1065
rect 50472 -1121 50520 -1065
rect 50576 -1121 51044 -1065
rect 51100 -1121 51148 -1065
rect 51204 -1121 51252 -1065
rect 51308 -1121 52318 -1065
rect 52374 -1121 52958 -1065
rect 53014 -1121 54238 -1065
rect 54294 -1121 54878 -1065
rect 54934 -1121 56454 -1065
rect 56510 -1121 57094 -1065
rect 57150 -1121 58374 -1065
rect 58430 -1121 59014 -1065
rect 59070 -1121 60028 -1065
rect 60084 -1121 60132 -1065
rect 60188 -1121 60236 -1065
rect 60292 -1121 60792 -1065
rect 60848 -1121 60896 -1065
rect 60952 -1121 61000 -1065
rect 61056 -1121 62014 -1065
rect 62070 -1121 62654 -1065
rect 62710 -1121 63934 -1065
rect 63990 -1121 64574 -1065
rect 64630 -1121 64640 -1065
rect 18499 -1169 64640 -1121
rect 18499 -1225 18509 -1169
rect 18565 -1225 19149 -1169
rect 19205 -1225 19789 -1169
rect 19845 -1225 20972 -1169
rect 21028 -1225 21076 -1169
rect 21132 -1225 21180 -1169
rect 21236 -1225 22270 -1169
rect 22326 -1225 22374 -1169
rect 22430 -1225 22478 -1169
rect 22534 -1225 23661 -1169
rect 23717 -1225 24301 -1169
rect 24357 -1225 24941 -1169
rect 24997 -1225 27630 -1169
rect 27686 -1225 28270 -1169
rect 28326 -1225 28910 -1169
rect 28966 -1225 30093 -1169
rect 30149 -1225 30197 -1169
rect 30253 -1225 30301 -1169
rect 30357 -1225 31650 -1169
rect 31706 -1225 31754 -1169
rect 31810 -1225 31858 -1169
rect 31914 -1225 32926 -1169
rect 32982 -1225 33566 -1169
rect 33622 -1225 34846 -1169
rect 34902 -1225 35486 -1169
rect 35542 -1225 37062 -1169
rect 37118 -1225 37702 -1169
rect 37758 -1225 38982 -1169
rect 39038 -1225 39622 -1169
rect 39678 -1225 40636 -1169
rect 40692 -1225 40740 -1169
rect 40796 -1225 40844 -1169
rect 40900 -1225 41356 -1169
rect 41412 -1225 41460 -1169
rect 41516 -1225 41564 -1169
rect 41620 -1225 42622 -1169
rect 42678 -1225 43262 -1169
rect 43318 -1225 44542 -1169
rect 44598 -1225 45182 -1169
rect 45238 -1225 46758 -1169
rect 46814 -1225 47398 -1169
rect 47454 -1225 48678 -1169
rect 48734 -1225 49318 -1169
rect 49374 -1225 50312 -1169
rect 50368 -1225 50416 -1169
rect 50472 -1225 50520 -1169
rect 50576 -1225 51044 -1169
rect 51100 -1225 51148 -1169
rect 51204 -1225 51252 -1169
rect 51308 -1225 52318 -1169
rect 52374 -1225 52958 -1169
rect 53014 -1225 54238 -1169
rect 54294 -1225 54878 -1169
rect 54934 -1225 56454 -1169
rect 56510 -1225 57094 -1169
rect 57150 -1225 58374 -1169
rect 58430 -1225 59014 -1169
rect 59070 -1225 60028 -1169
rect 60084 -1225 60132 -1169
rect 60188 -1225 60236 -1169
rect 60292 -1225 60792 -1169
rect 60848 -1225 60896 -1169
rect 60952 -1225 61000 -1169
rect 61056 -1225 62014 -1169
rect 62070 -1225 62654 -1169
rect 62710 -1225 63934 -1169
rect 63990 -1225 64574 -1169
rect 64630 -1225 64640 -1169
rect 18499 -1235 64640 -1225
rect 3384 -1324 3460 -1314
rect 4024 -1324 4100 -1314
rect 4664 -1324 4740 -1314
rect 5245 -1324 5425 -1314
rect 6249 -1324 6325 -1314
rect 6889 -1324 6965 -1314
rect 7529 -1324 7605 -1314
rect 8484 -1324 8560 -1314
rect 9380 -1324 9456 -1314
rect 10276 -1324 10352 -1314
rect 14660 -1322 14736 -1312
rect 15300 -1322 15376 -1312
rect 15940 -1322 16016 -1312
rect 16879 -1322 17059 -1312
rect 3384 -1380 3394 -1324
rect 3450 -1380 4034 -1324
rect 4090 -1380 4674 -1324
rect 4730 -1380 5255 -1324
rect 5311 -1380 5359 -1324
rect 5415 -1380 6259 -1324
rect 6315 -1380 6899 -1324
rect 6955 -1380 7539 -1324
rect 7595 -1380 8494 -1324
rect 8550 -1380 9390 -1324
rect 9446 -1380 10286 -1324
rect 10342 -1380 10352 -1324
rect 3384 -1428 10352 -1380
rect 3384 -1484 3394 -1428
rect 3450 -1484 4034 -1428
rect 4090 -1484 4674 -1428
rect 4730 -1484 5255 -1428
rect 5311 -1484 5359 -1428
rect 5415 -1484 6259 -1428
rect 6315 -1484 6899 -1428
rect 6955 -1484 7539 -1428
rect 7595 -1484 8494 -1428
rect 8550 -1484 9390 -1428
rect 9446 -1484 10286 -1428
rect 10342 -1484 10352 -1428
rect 3384 -1494 3460 -1484
rect 4024 -1494 4100 -1484
rect 4664 -1494 4740 -1484
rect 5245 -1494 5425 -1484
rect 6249 -1494 6325 -1484
rect 6889 -1494 6965 -1484
rect 7529 -1494 7605 -1484
rect 8484 -1494 8560 -1484
rect 9380 -1494 9456 -1484
rect 10276 -1494 10352 -1484
rect 11153 -1332 11333 -1322
rect 11866 -1332 11942 -1322
rect 12762 -1332 12838 -1322
rect 13658 -1332 13734 -1322
rect 11153 -1388 11163 -1332
rect 11219 -1388 11267 -1332
rect 11323 -1388 11876 -1332
rect 11932 -1388 12772 -1332
rect 12828 -1388 13668 -1332
rect 13724 -1388 13734 -1332
rect 11153 -1436 13734 -1388
rect 11153 -1492 11163 -1436
rect 11219 -1492 11267 -1436
rect 11323 -1492 11876 -1436
rect 11932 -1492 12772 -1436
rect 12828 -1492 13668 -1436
rect 13724 -1492 13734 -1436
rect 14660 -1378 14670 -1322
rect 14726 -1378 15310 -1322
rect 15366 -1378 15950 -1322
rect 16006 -1378 16889 -1322
rect 16945 -1378 16993 -1322
rect 17049 -1378 17059 -1322
rect 14660 -1426 17059 -1378
rect 14660 -1482 14670 -1426
rect 14726 -1482 15310 -1426
rect 15366 -1482 15950 -1426
rect 16006 -1482 16889 -1426
rect 16945 -1482 16993 -1426
rect 17049 -1482 17059 -1426
rect 17355 -1396 18815 -1386
rect 17355 -1452 17365 -1396
rect 17421 -1452 18749 -1396
rect 18805 -1452 18815 -1396
rect 17355 -1462 18815 -1452
rect 19379 -1396 24127 -1386
rect 19379 -1452 19389 -1396
rect 19445 -1452 24061 -1396
rect 24117 -1452 24127 -1396
rect 19379 -1462 24127 -1452
rect 24691 -1396 27936 -1386
rect 24691 -1452 24701 -1396
rect 24757 -1452 26085 -1396
rect 26141 -1452 26486 -1396
rect 26542 -1452 27870 -1396
rect 27926 -1452 27936 -1396
rect 24691 -1462 27936 -1452
rect 14660 -1492 14736 -1482
rect 15300 -1492 15376 -1482
rect 15940 -1492 16016 -1482
rect 16879 -1492 17059 -1482
rect 11153 -1502 11333 -1492
rect 11866 -1502 11942 -1492
rect 12762 -1502 12838 -1492
rect 13658 -1502 13734 -1492
rect -260 -1572 -80 -1562
rect 741 -1572 921 -1562
rect -260 -1628 -250 -1572
rect -194 -1628 -146 -1572
rect -90 -1628 751 -1572
rect 807 -1628 855 -1572
rect 911 -1628 921 -1572
rect -260 -1676 921 -1628
rect -260 -1732 -250 -1676
rect -194 -1732 -146 -1676
rect -90 -1732 751 -1676
rect 807 -1732 855 -1676
rect 911 -1732 921 -1676
rect -260 -1742 -80 -1732
rect 741 -1742 921 -1732
rect 2395 -1663 2575 -1653
rect 3624 -1663 3700 -1653
rect 2395 -1719 2405 -1663
rect 2461 -1719 2509 -1663
rect 2565 -1719 3634 -1663
rect 3690 -1719 3700 -1663
rect 2395 -1767 3700 -1719
rect 2395 -1823 2405 -1767
rect 2461 -1823 2509 -1767
rect 2565 -1823 3634 -1767
rect 3690 -1823 3700 -1767
rect 2395 -1833 2575 -1823
rect 3624 -1833 3700 -1823
rect 16633 -2719 30294 -2709
rect 6896 -2746 7076 -2736
rect 7789 -2746 7969 -2736
rect 6896 -2802 6906 -2746
rect 6962 -2802 7010 -2746
rect 7066 -2802 7799 -2746
rect 7855 -2802 7903 -2746
rect 7959 -2802 7969 -2746
rect 6896 -2850 7969 -2802
rect 6896 -2906 6906 -2850
rect 6962 -2906 7010 -2850
rect 7066 -2906 7799 -2850
rect 7855 -2906 7903 -2850
rect 7959 -2906 7969 -2850
rect 6896 -2916 7076 -2906
rect 7789 -2916 7969 -2906
rect 16633 -2775 16643 -2719
rect 16699 -2775 16747 -2719
rect 16803 -2775 16851 -2719
rect 16907 -2775 29812 -2719
rect 29868 -2775 29916 -2719
rect 29972 -2775 30020 -2719
rect 30076 -2775 30124 -2719
rect 30180 -2775 30228 -2719
rect 30284 -2775 30294 -2719
rect 16633 -2823 30294 -2775
rect 16633 -2879 16643 -2823
rect 16699 -2879 16747 -2823
rect 16803 -2879 16851 -2823
rect 16907 -2879 29812 -2823
rect 29868 -2879 29916 -2823
rect 29972 -2879 30020 -2823
rect 30076 -2879 30124 -2823
rect 30180 -2879 30228 -2823
rect 30284 -2879 30294 -2823
rect 16633 -2927 30294 -2879
rect 16633 -2983 16643 -2927
rect 16699 -2983 16747 -2927
rect 16803 -2983 16851 -2927
rect 16907 -2983 29812 -2927
rect 29868 -2983 29916 -2927
rect 29972 -2983 30020 -2927
rect 30076 -2983 30124 -2927
rect 30180 -2983 30228 -2927
rect 30284 -2983 30294 -2927
rect 16633 -2993 30294 -2983
rect 17070 -3061 29734 -3051
rect 8703 -3113 8779 -3103
rect 9792 -3113 9972 -3103
rect 8703 -3169 8713 -3113
rect 8769 -3169 9802 -3113
rect 9858 -3169 9906 -3113
rect 9962 -3169 9972 -3113
rect 8703 -3217 9972 -3169
rect 8703 -3273 8713 -3217
rect 8769 -3273 9802 -3217
rect 9858 -3273 9906 -3217
rect 9962 -3273 9972 -3217
rect 8703 -3283 8779 -3273
rect 9792 -3283 9972 -3273
rect 17070 -3117 17080 -3061
rect 17136 -3117 17184 -3061
rect 17240 -3117 17288 -3061
rect 17344 -3117 29252 -3061
rect 29308 -3117 29356 -3061
rect 29412 -3117 29460 -3061
rect 29516 -3117 29564 -3061
rect 29620 -3117 29668 -3061
rect 29724 -3117 29734 -3061
rect 17070 -3165 29734 -3117
rect 17070 -3221 17080 -3165
rect 17136 -3221 17184 -3165
rect 17240 -3221 17288 -3165
rect 17344 -3221 29252 -3165
rect 29308 -3221 29356 -3165
rect 29412 -3221 29460 -3165
rect 29516 -3221 29564 -3165
rect 29620 -3221 29668 -3165
rect 29724 -3221 29734 -3165
rect 17070 -3269 29734 -3221
rect 17070 -3325 17080 -3269
rect 17136 -3325 17184 -3269
rect 17240 -3325 17288 -3269
rect 17344 -3325 29252 -3269
rect 29308 -3325 29356 -3269
rect 29412 -3325 29460 -3269
rect 29516 -3325 29564 -3269
rect 29620 -3325 29668 -3269
rect 29724 -3325 29734 -3269
rect 17070 -3335 29734 -3325
rect 7343 -3446 7419 -3436
rect 7663 -3446 7739 -3436
rect 7983 -3446 8059 -3436
rect 8303 -3446 8379 -3436
rect 7343 -3502 7353 -3446
rect 7409 -3502 7673 -3446
rect 7729 -3502 7993 -3446
rect 8049 -3502 8313 -3446
rect 8369 -3502 8379 -3446
rect 7343 -3550 8379 -3502
rect 7343 -3606 7353 -3550
rect 7409 -3606 7673 -3550
rect 7729 -3606 7993 -3550
rect 8049 -3606 8313 -3550
rect 8369 -3606 8379 -3550
rect 7343 -3616 7419 -3606
rect 7663 -3616 7739 -3606
rect 7983 -3616 8059 -3606
rect 8303 -3616 8379 -3606
rect 8463 -3446 8539 -3437
rect 14200 -3446 14380 -3436
rect 8463 -3502 8473 -3446
rect 8529 -3502 14210 -3446
rect 14266 -3502 14314 -3446
rect 14370 -3502 14380 -3446
rect 8463 -3550 14380 -3502
rect 8463 -3606 8473 -3550
rect 8529 -3606 14210 -3550
rect 14266 -3606 14314 -3550
rect 14370 -3606 14380 -3550
rect 8463 -3617 8539 -3606
rect 14200 -3616 14380 -3606
rect 10058 -3711 10238 -3701
rect 8782 -3753 8858 -3743
rect 10058 -3753 10068 -3711
rect 8782 -3809 8792 -3753
rect 8848 -3767 10068 -3753
rect 10124 -3767 10172 -3711
rect 10228 -3767 10238 -3711
rect 8848 -3809 10238 -3767
rect 8782 -3819 8858 -3809
rect 10058 -3815 10238 -3809
rect 10058 -3871 10068 -3815
rect 10124 -3871 10172 -3815
rect 10228 -3871 10238 -3815
rect 10058 -3881 10238 -3871
rect 16848 -3711 17028 -3701
rect 23634 -3711 23814 -3701
rect 16848 -3767 16858 -3711
rect 16914 -3767 16962 -3711
rect 17018 -3767 23644 -3711
rect 23700 -3767 23748 -3711
rect 23804 -3767 23814 -3711
rect 16848 -3815 23814 -3767
rect 16848 -3871 16858 -3815
rect 16914 -3871 16962 -3815
rect 17018 -3871 23644 -3815
rect 23700 -3871 23748 -3815
rect 23804 -3871 23814 -3815
rect 16848 -3881 17028 -3871
rect 23634 -3881 23814 -3871
rect 2561 -3982 2741 -3972
rect 7503 -3982 7579 -3973
rect 2561 -4038 2571 -3982
rect 2627 -4038 2675 -3982
rect 2731 -4038 7513 -3982
rect 7569 -4038 7579 -3982
rect 2561 -4086 7579 -4038
rect 2561 -4142 2571 -4086
rect 2627 -4142 2675 -4086
rect 2731 -4142 7513 -4086
rect 7569 -4142 7579 -4086
rect 2561 -4152 2741 -4142
rect 7503 -4153 7579 -4142
rect 7663 -3982 7739 -3972
rect 7983 -3982 8059 -3972
rect 8303 -3982 8379 -3972
rect 8623 -3982 8699 -3972
rect 7663 -4038 7673 -3982
rect 7729 -4038 7993 -3982
rect 8049 -4038 8313 -3982
rect 8369 -4038 8633 -3982
rect 8689 -4038 8699 -3982
rect 7663 -4086 8699 -4038
rect 7663 -4142 7673 -4086
rect 7729 -4142 7993 -4086
rect 8049 -4142 8313 -4086
rect 8369 -4142 8633 -4086
rect 8689 -4142 8699 -4086
rect 7663 -4152 7739 -4142
rect 7983 -4152 8059 -4142
rect 8303 -4152 8379 -4142
rect 8623 -4152 8699 -4142
rect 9792 -4237 9972 -4227
rect 8585 -4289 8661 -4279
rect 9792 -4289 9802 -4237
rect 8585 -4345 8595 -4289
rect 8651 -4293 9802 -4289
rect 9858 -4293 9906 -4237
rect 9962 -4293 9972 -4237
rect 8651 -4341 9972 -4293
rect 8651 -4345 9802 -4341
rect 8585 -4355 8661 -4345
rect 9792 -4397 9802 -4345
rect 9858 -4397 9906 -4341
rect 9962 -4397 9972 -4341
rect 9792 -4407 9972 -4397
rect 7343 -4518 7419 -4508
rect 7663 -4518 7739 -4508
rect 7983 -4518 8059 -4508
rect 8303 -4518 8379 -4508
rect 8623 -4518 8699 -4508
rect 7343 -4574 7353 -4518
rect 7409 -4574 7673 -4518
rect 7729 -4574 7993 -4518
rect 8049 -4574 8313 -4518
rect 8369 -4574 8633 -4518
rect 8689 -4574 8699 -4518
rect 7343 -4622 8699 -4574
rect 7343 -4678 7353 -4622
rect 7409 -4678 7673 -4622
rect 7729 -4678 7993 -4622
rect 8049 -4678 8313 -4622
rect 8369 -4678 8633 -4622
rect 8689 -4678 8699 -4622
rect 7343 -4688 7419 -4678
rect 7663 -4688 7739 -4678
rect 7983 -4688 8059 -4678
rect 8303 -4688 8379 -4678
rect 8623 -4688 8699 -4678
rect 13726 -4691 21250 -4681
rect 2229 -4736 2305 -4726
rect 5134 -4736 5314 -4726
rect 2229 -4792 2239 -4736
rect 2295 -4792 5144 -4736
rect 5200 -4792 5248 -4736
rect 5304 -4792 5314 -4736
rect 13726 -4747 13736 -4691
rect 13792 -4747 13840 -4691
rect 13896 -4747 13944 -4691
rect 14000 -4747 21184 -4691
rect 21240 -4747 21250 -4691
rect 2229 -4840 5314 -4792
rect 10058 -4771 10238 -4761
rect 2229 -4896 2239 -4840
rect 2295 -4896 5144 -4840
rect 5200 -4896 5248 -4840
rect 5304 -4896 5314 -4840
rect 8703 -4823 8779 -4813
rect 10058 -4823 10068 -4771
rect 8703 -4879 8713 -4823
rect 8769 -4827 10068 -4823
rect 10124 -4827 10172 -4771
rect 10228 -4827 10238 -4771
rect 8769 -4875 10238 -4827
rect 8769 -4879 10068 -4875
rect 8703 -4889 8779 -4879
rect 2229 -4906 2305 -4896
rect 5134 -4906 5314 -4896
rect 10058 -4931 10068 -4879
rect 10124 -4931 10172 -4875
rect 10228 -4931 10238 -4875
rect 10058 -4941 10238 -4931
rect 13726 -4795 21250 -4747
rect 13726 -4851 13736 -4795
rect 13792 -4851 13840 -4795
rect 13896 -4851 13944 -4795
rect 14000 -4851 21184 -4795
rect 21240 -4851 21250 -4795
rect 13726 -4899 21250 -4851
rect 13726 -4955 13736 -4899
rect 13792 -4955 13840 -4899
rect 13896 -4955 13944 -4899
rect 14000 -4955 21184 -4899
rect 21240 -4955 21250 -4899
rect 13726 -4965 21250 -4955
rect 3525 -5026 3601 -5016
rect 5607 -5026 5787 -5016
rect 3525 -5082 3535 -5026
rect 3591 -5082 5617 -5026
rect 5673 -5082 5721 -5026
rect 5777 -5082 5787 -5026
rect 29802 -5018 32080 -5008
rect 3525 -5130 5787 -5082
rect 3525 -5186 3535 -5130
rect 3591 -5186 5617 -5130
rect 5673 -5186 5721 -5130
rect 5777 -5186 5787 -5130
rect 3525 -5196 3601 -5186
rect 5607 -5196 5787 -5186
rect 6058 -5054 6238 -5044
rect 6368 -5054 6548 -5044
rect 7343 -5053 7419 -5044
rect 7663 -5053 7739 -5044
rect 7983 -5053 8059 -5044
rect 8303 -5053 8379 -5044
rect 8623 -5053 8699 -5044
rect 7343 -5054 8699 -5053
rect 6058 -5110 6068 -5054
rect 6124 -5110 6172 -5054
rect 6228 -5110 6378 -5054
rect 6434 -5110 6482 -5054
rect 6538 -5110 7353 -5054
rect 7409 -5110 7673 -5054
rect 7729 -5110 7993 -5054
rect 8049 -5110 8313 -5054
rect 8369 -5110 8633 -5054
rect 8689 -5110 8699 -5054
rect 6058 -5158 8699 -5110
rect 6058 -5214 6068 -5158
rect 6124 -5214 6172 -5158
rect 6228 -5214 6378 -5158
rect 6434 -5214 6482 -5158
rect 6538 -5214 7353 -5158
rect 7409 -5214 7673 -5158
rect 7729 -5214 7993 -5158
rect 8049 -5214 8313 -5158
rect 8369 -5214 8633 -5158
rect 8689 -5214 8699 -5158
rect 6058 -5224 6238 -5214
rect 6368 -5224 6548 -5214
rect 7343 -5224 7419 -5214
rect 7663 -5224 7739 -5214
rect 7983 -5224 8059 -5214
rect 8303 -5224 8379 -5214
rect 8623 -5224 8699 -5214
rect 29802 -5074 29812 -5018
rect 29868 -5074 29916 -5018
rect 29972 -5074 30020 -5018
rect 30076 -5074 30124 -5018
rect 30180 -5074 30228 -5018
rect 30284 -5074 31598 -5018
rect 31654 -5074 31702 -5018
rect 31758 -5074 31806 -5018
rect 31862 -5074 31910 -5018
rect 31966 -5074 32014 -5018
rect 32070 -5074 32080 -5018
rect 29802 -5122 32080 -5074
rect 29802 -5178 29812 -5122
rect 29868 -5178 29916 -5122
rect 29972 -5178 30020 -5122
rect 30076 -5178 30124 -5122
rect 30180 -5178 30228 -5122
rect 30284 -5178 31598 -5122
rect 31654 -5178 31702 -5122
rect 31758 -5178 31806 -5122
rect 31862 -5178 31910 -5122
rect 31966 -5178 32014 -5122
rect 32070 -5178 32080 -5122
rect 29802 -5226 32080 -5178
rect 8782 -5255 8858 -5245
rect 9520 -5255 9700 -5245
rect 9792 -5255 9972 -5247
rect 8782 -5311 8792 -5255
rect 8848 -5311 9530 -5255
rect 9586 -5311 9634 -5255
rect 9690 -5257 9972 -5255
rect 9690 -5311 9802 -5257
rect 8782 -5313 9802 -5311
rect 9858 -5313 9906 -5257
rect 9962 -5313 9972 -5257
rect 3093 -5350 3169 -5340
rect 4898 -5350 5078 -5340
rect 3093 -5406 3103 -5350
rect 3159 -5406 4908 -5350
rect 4964 -5406 5012 -5350
rect 5068 -5406 5078 -5350
rect 3093 -5454 5078 -5406
rect 8782 -5359 9972 -5313
rect 8782 -5415 8792 -5359
rect 8848 -5415 9530 -5359
rect 9586 -5415 9634 -5359
rect 9690 -5361 9972 -5359
rect 9690 -5415 9802 -5361
rect 8782 -5425 8858 -5415
rect 9520 -5425 9700 -5415
rect 9792 -5417 9802 -5415
rect 9858 -5417 9906 -5361
rect 9962 -5417 9972 -5361
rect 9792 -5427 9972 -5417
rect 29802 -5282 29812 -5226
rect 29868 -5282 29916 -5226
rect 29972 -5282 30020 -5226
rect 30076 -5282 30124 -5226
rect 30180 -5282 30228 -5226
rect 30284 -5282 31598 -5226
rect 31654 -5282 31702 -5226
rect 31758 -5282 31806 -5226
rect 31862 -5282 31910 -5226
rect 31966 -5282 32014 -5226
rect 32070 -5282 32080 -5226
rect 29802 -5330 32080 -5282
rect 29802 -5386 29812 -5330
rect 29868 -5386 29916 -5330
rect 29972 -5386 30020 -5330
rect 30076 -5386 30124 -5330
rect 30180 -5386 30228 -5330
rect 30284 -5386 31598 -5330
rect 31654 -5386 31702 -5330
rect 31758 -5386 31806 -5330
rect 31862 -5386 31910 -5330
rect 31966 -5386 32014 -5330
rect 32070 -5386 32080 -5330
rect 3093 -5510 3103 -5454
rect 3159 -5510 4908 -5454
rect 4964 -5510 5012 -5454
rect 5068 -5510 5078 -5454
rect 29802 -5434 32080 -5386
rect 29802 -5490 29812 -5434
rect 29868 -5490 29916 -5434
rect 29972 -5490 30020 -5434
rect 30076 -5490 30124 -5434
rect 30180 -5490 30228 -5434
rect 30284 -5490 31598 -5434
rect 31654 -5490 31702 -5434
rect 31758 -5490 31806 -5434
rect 31862 -5490 31910 -5434
rect 31966 -5490 32014 -5434
rect 32070 -5490 32080 -5434
rect 29802 -5500 32080 -5490
rect 3093 -5520 3169 -5510
rect 4898 -5520 5078 -5510
rect 5365 -5544 5545 -5534
rect 5365 -5600 5375 -5544
rect 5431 -5600 5479 -5544
rect 5535 -5590 5545 -5544
rect 8463 -5590 8539 -5580
rect 5535 -5600 8473 -5590
rect 5365 -5646 8473 -5600
rect 8529 -5646 8539 -5590
rect 5365 -5648 8539 -5646
rect 5365 -5704 5375 -5648
rect 5431 -5704 5479 -5648
rect 5535 -5694 8539 -5648
rect 5535 -5704 8473 -5694
rect 2933 -5752 3113 -5742
rect 5365 -5750 8473 -5704
rect 8529 -5750 8539 -5694
rect 5365 -5752 5545 -5750
rect 2933 -5808 2943 -5752
rect 2999 -5808 3047 -5752
rect 3103 -5808 5375 -5752
rect 5431 -5808 5479 -5752
rect 5535 -5808 5545 -5752
rect 8463 -5761 8539 -5750
rect 14566 -5593 34352 -5583
rect 14566 -5649 14576 -5593
rect 14632 -5649 15184 -5593
rect 15240 -5649 15792 -5593
rect 15848 -5649 34154 -5593
rect 34210 -5649 34258 -5593
rect 34314 -5649 34352 -5593
rect 14566 -5697 34352 -5649
rect 14566 -5753 14576 -5697
rect 14632 -5753 15184 -5697
rect 15240 -5753 15792 -5697
rect 15848 -5753 34154 -5697
rect 34210 -5753 34258 -5697
rect 34314 -5753 34352 -5697
rect 2933 -5856 5545 -5808
rect 2933 -5912 2943 -5856
rect 2999 -5912 3047 -5856
rect 3103 -5912 5375 -5856
rect 5431 -5912 5479 -5856
rect 5535 -5912 5545 -5856
rect 2933 -5922 3113 -5912
rect 5365 -5922 5545 -5912
rect 8782 -5770 8858 -5760
rect 10058 -5770 10238 -5760
rect 14566 -5763 34352 -5753
rect 8782 -5826 8792 -5770
rect 8848 -5826 10068 -5770
rect 10124 -5826 10172 -5770
rect 10228 -5826 10238 -5770
rect 8782 -5874 10238 -5826
rect 8782 -5930 8792 -5874
rect 8848 -5930 10068 -5874
rect 10124 -5930 10172 -5874
rect 10228 -5930 10238 -5874
rect 8782 -5940 8858 -5930
rect 10058 -5940 10238 -5930
rect 741 -5996 921 -5986
rect 2239 -5996 2315 -5986
rect 9253 -5996 9433 -5986
rect 741 -6052 751 -5996
rect 807 -6052 855 -5996
rect 911 -6052 2249 -5996
rect 2305 -6052 9263 -5996
rect 9319 -6052 9367 -5996
rect 9423 -6052 9433 -5996
rect 741 -6100 9433 -6052
rect 741 -6156 751 -6100
rect 807 -6156 855 -6100
rect 911 -6156 2249 -6100
rect 2305 -6156 9263 -6100
rect 9319 -6156 9367 -6100
rect 9423 -6156 9433 -6100
rect 741 -6166 921 -6156
rect 2239 -6166 2315 -6156
rect 9253 -6166 9433 -6156
rect 15070 -5993 20368 -5983
rect 15070 -6049 15080 -5993
rect 15136 -6049 15184 -5993
rect 15240 -6049 15288 -5993
rect 15344 -6049 20094 -5993
rect 20150 -6049 20198 -5993
rect 20254 -6049 20302 -5993
rect 20358 -6049 20368 -5993
rect 15070 -6097 20368 -6049
rect 15070 -6153 15080 -6097
rect 15136 -6153 15184 -6097
rect 15240 -6153 15288 -6097
rect 15344 -6153 20094 -6097
rect 20150 -6153 20198 -6097
rect 20254 -6153 20302 -6097
rect 20358 -6153 20368 -6097
rect 15070 -6201 20368 -6153
rect 15070 -6257 15080 -6201
rect 15136 -6257 15184 -6201
rect 15240 -6257 15288 -6201
rect 15344 -6257 20094 -6201
rect 20150 -6257 20198 -6201
rect 20254 -6257 20302 -6201
rect 20358 -6257 20368 -6201
rect 5607 -6268 5787 -6258
rect 6632 -6268 6812 -6258
rect 15070 -6267 20368 -6257
rect 5607 -6324 5617 -6268
rect 5673 -6324 5721 -6268
rect 5777 -6324 6642 -6268
rect 6698 -6324 6746 -6268
rect 6802 -6324 6812 -6268
rect 5607 -6372 6812 -6324
rect 5607 -6428 5617 -6372
rect 5673 -6428 5721 -6372
rect 5777 -6428 6642 -6372
rect 6698 -6428 6746 -6372
rect 6802 -6428 6812 -6372
rect 5607 -6438 5787 -6428
rect 6632 -6438 6812 -6428
rect 8383 -6446 8459 -6436
rect 9520 -6446 9700 -6436
rect 8383 -6502 8393 -6446
rect 8449 -6502 9530 -6446
rect 9586 -6502 9634 -6446
rect 9690 -6502 9700 -6446
rect 8383 -6550 9700 -6502
rect 3437 -6612 3513 -6602
rect 4658 -6612 4838 -6602
rect 3437 -6668 3447 -6612
rect 3503 -6668 4668 -6612
rect 4724 -6668 4772 -6612
rect 4828 -6668 4838 -6612
rect 8383 -6606 8393 -6550
rect 8449 -6606 9530 -6550
rect 9586 -6606 9634 -6550
rect 9690 -6606 9700 -6550
rect 8383 -6616 8459 -6606
rect 9520 -6616 9700 -6606
rect 3437 -6716 4838 -6668
rect 3437 -6772 3447 -6716
rect 3503 -6772 4668 -6716
rect 4724 -6772 4772 -6716
rect 4828 -6772 4838 -6716
rect 3437 -6782 3513 -6772
rect 4658 -6782 4838 -6772
rect 4898 -6755 5078 -6745
rect 6096 -6755 6172 -6745
rect 4898 -6811 4908 -6755
rect 4964 -6811 5012 -6755
rect 5068 -6811 6106 -6755
rect 6162 -6811 6172 -6755
rect 4898 -6859 6172 -6811
rect 4898 -6915 4908 -6859
rect 4964 -6915 5012 -6859
rect 5068 -6915 6106 -6859
rect 6162 -6915 6172 -6859
rect 4898 -6925 5078 -6915
rect 6096 -6925 6172 -6915
rect 12614 -6861 14687 -6851
rect 12614 -6917 12624 -6861
rect 12680 -6917 14413 -6861
rect 14469 -6917 14517 -6861
rect 14573 -6917 14621 -6861
rect 14677 -6917 14687 -6861
rect 12614 -6965 14687 -6917
rect 12614 -7021 12624 -6965
rect 12680 -7021 14413 -6965
rect 14469 -7021 14517 -6965
rect 14573 -7021 14621 -6965
rect 14677 -7021 14687 -6965
rect 12614 -7069 14687 -7021
rect 12614 -7125 12624 -7069
rect 12680 -7125 14413 -7069
rect 14469 -7125 14517 -7069
rect 14573 -7125 14621 -7069
rect 14677 -7125 14687 -7069
rect 4658 -7141 4838 -7131
rect 6026 -7141 6206 -7131
rect 12614 -7135 14687 -7125
rect 15070 -6861 15354 -6851
rect 15070 -6917 15080 -6861
rect 15136 -6917 15184 -6861
rect 15240 -6917 15288 -6861
rect 15344 -6917 15354 -6861
rect 15070 -6965 15354 -6917
rect 15070 -7021 15080 -6965
rect 15136 -7021 15184 -6965
rect 15240 -7021 15288 -6965
rect 15344 -7021 15354 -6965
rect 15070 -7069 15354 -7021
rect 15070 -7125 15080 -7069
rect 15136 -7125 15184 -7069
rect 15240 -7125 15288 -7069
rect 15344 -7125 15354 -7069
rect 15070 -7135 15354 -7125
rect 15685 -6899 20610 -6889
rect 15685 -6955 15695 -6899
rect 15751 -6955 15799 -6899
rect 15855 -6955 15903 -6899
rect 15959 -6955 18624 -6899
rect 18680 -6955 18944 -6899
rect 19000 -6955 19264 -6899
rect 19320 -6955 19584 -6899
rect 19640 -6955 19904 -6899
rect 19960 -6955 20224 -6899
rect 20280 -6955 20544 -6899
rect 20600 -6955 20610 -6899
rect 15685 -7003 20610 -6955
rect 15685 -7059 15695 -7003
rect 15751 -7059 15799 -7003
rect 15855 -7059 15903 -7003
rect 15959 -7059 18624 -7003
rect 18680 -7059 18944 -7003
rect 19000 -7059 19264 -7003
rect 19320 -7059 19584 -7003
rect 19640 -7059 19904 -7003
rect 19960 -7059 20224 -7003
rect 20280 -7059 20544 -7003
rect 20600 -7059 20610 -7003
rect 15685 -7107 20610 -7059
rect 4658 -7197 4668 -7141
rect 4724 -7197 4772 -7141
rect 4828 -7197 6036 -7141
rect 6092 -7197 6140 -7141
rect 6196 -7197 6206 -7141
rect 4658 -7245 6206 -7197
rect 4658 -7301 4668 -7245
rect 4724 -7301 4772 -7245
rect 4828 -7301 6036 -7245
rect 6092 -7301 6140 -7245
rect 6196 -7301 6206 -7245
rect 4658 -7311 4838 -7301
rect 6026 -7311 6206 -7301
rect 6632 -7151 6812 -7141
rect 8910 -7151 9090 -7141
rect 10432 -7151 10612 -7141
rect 10819 -7151 10999 -7141
rect 6632 -7207 6642 -7151
rect 6698 -7207 6746 -7151
rect 6802 -7207 8920 -7151
rect 8976 -7207 9024 -7151
rect 9080 -7207 10442 -7151
rect 10498 -7207 10546 -7151
rect 10602 -7207 10829 -7151
rect 10885 -7207 10933 -7151
rect 10989 -7207 10999 -7151
rect 15685 -7163 15695 -7107
rect 15751 -7163 15799 -7107
rect 15855 -7163 15903 -7107
rect 15959 -7163 18624 -7107
rect 18680 -7163 18944 -7107
rect 19000 -7163 19264 -7107
rect 19320 -7163 19584 -7107
rect 19640 -7163 19904 -7107
rect 19960 -7163 20224 -7107
rect 20280 -7163 20544 -7107
rect 20600 -7163 20610 -7107
rect 15685 -7173 20610 -7163
rect 29802 -7030 42321 -7020
rect 29802 -7086 29812 -7030
rect 29868 -7086 29916 -7030
rect 29972 -7086 30020 -7030
rect 30076 -7086 30124 -7030
rect 30180 -7086 30228 -7030
rect 30284 -7086 42022 -7030
rect 42078 -7086 42126 -7030
rect 42182 -7086 42230 -7030
rect 42286 -7086 42321 -7030
rect 29802 -7134 42321 -7086
rect 6632 -7255 10999 -7207
rect 6632 -7311 6642 -7255
rect 6698 -7311 6746 -7255
rect 6802 -7311 8920 -7255
rect 8976 -7311 9024 -7255
rect 9080 -7311 10442 -7255
rect 10498 -7311 10546 -7255
rect 10602 -7311 10829 -7255
rect 10885 -7311 10933 -7255
rect 10989 -7311 10999 -7255
rect 6632 -7321 6812 -7311
rect 8910 -7321 9090 -7311
rect 10432 -7321 10612 -7311
rect 10819 -7321 10999 -7311
rect 29802 -7190 29812 -7134
rect 29868 -7190 29916 -7134
rect 29972 -7190 30020 -7134
rect 30076 -7190 30124 -7134
rect 30180 -7190 30228 -7134
rect 30284 -7190 42022 -7134
rect 42078 -7190 42126 -7134
rect 42182 -7190 42230 -7134
rect 42286 -7190 42321 -7134
rect 29802 -7238 42321 -7190
rect 29802 -7294 29812 -7238
rect 29868 -7294 29916 -7238
rect 29972 -7294 30020 -7238
rect 30076 -7294 30124 -7238
rect 30180 -7294 30228 -7238
rect 30284 -7294 42022 -7238
rect 42078 -7294 42126 -7238
rect 42182 -7294 42230 -7238
rect 42286 -7294 42321 -7238
rect 29802 -7342 42321 -7294
rect 3485 -7382 3561 -7372
rect 5936 -7382 6012 -7374
rect 3485 -7438 3495 -7382
rect 3551 -7384 6012 -7382
rect 3551 -7438 5946 -7384
rect 3485 -7440 5946 -7438
rect 6002 -7440 6012 -7384
rect 3485 -7486 6012 -7440
rect 3485 -7542 3495 -7486
rect 3551 -7488 6012 -7486
rect 3551 -7542 5946 -7488
rect 3485 -7552 3561 -7542
rect 5936 -7544 5946 -7542
rect 6002 -7544 6012 -7488
rect 5936 -7554 6012 -7544
rect 6368 -7390 6548 -7380
rect 6368 -7446 6378 -7390
rect 6434 -7446 6482 -7390
rect 6538 -7446 6548 -7390
rect 6368 -7494 6548 -7446
rect 6368 -7550 6378 -7494
rect 6434 -7550 6482 -7494
rect 6538 -7550 6548 -7494
rect 29802 -7398 29812 -7342
rect 29868 -7398 29916 -7342
rect 29972 -7398 30020 -7342
rect 30076 -7398 30124 -7342
rect 30180 -7398 30228 -7342
rect 30284 -7398 42022 -7342
rect 42078 -7398 42126 -7342
rect 42182 -7398 42230 -7342
rect 42286 -7398 42321 -7342
rect 29802 -7446 42321 -7398
rect 29802 -7502 29812 -7446
rect 29868 -7502 29916 -7446
rect 29972 -7502 30020 -7446
rect 30076 -7502 30124 -7446
rect 30180 -7502 30228 -7446
rect 30284 -7502 42022 -7446
rect 42078 -7502 42126 -7446
rect 42182 -7502 42230 -7446
rect 42286 -7502 42321 -7446
rect 29802 -7512 42321 -7502
rect 6368 -7560 6548 -7550
rect 44536 -7954 45028 -7944
rect 44536 -8010 44546 -7954
rect 44602 -8010 44650 -7954
rect 44706 -8010 44754 -7954
rect 44810 -8010 44858 -7954
rect 44914 -8010 44962 -7954
rect 45018 -8010 45028 -7954
rect 5884 -8028 6064 -8018
rect 11532 -8028 11712 -8018
rect 5884 -8084 5894 -8028
rect 5950 -8084 5998 -8028
rect 6054 -8084 11542 -8028
rect 11598 -8084 11646 -8028
rect 11702 -8084 11712 -8028
rect 5884 -8132 11712 -8084
rect 5884 -8188 5894 -8132
rect 5950 -8188 5998 -8132
rect 6054 -8188 11542 -8132
rect 11598 -8188 11646 -8132
rect 11702 -8188 11712 -8132
rect 5884 -8198 6064 -8188
rect 11532 -8198 11712 -8188
rect 34706 -8054 35198 -8044
rect 34706 -8110 34716 -8054
rect 34772 -8110 34820 -8054
rect 34876 -8110 34924 -8054
rect 34980 -8110 35028 -8054
rect 35084 -8110 35132 -8054
rect 35188 -8110 35198 -8054
rect 34706 -8158 35198 -8110
rect 34706 -8214 34716 -8158
rect 34772 -8214 34820 -8158
rect 34876 -8214 34924 -8158
rect 34980 -8214 35028 -8158
rect 35084 -8214 35132 -8158
rect 35188 -8214 35198 -8158
rect 34706 -8262 35198 -8214
rect 5134 -8280 5314 -8270
rect 9827 -8280 10007 -8270
rect 5134 -8336 5144 -8280
rect 5200 -8336 5248 -8280
rect 5304 -8336 9837 -8280
rect 9893 -8336 9941 -8280
rect 9997 -8336 10007 -8280
rect 5134 -8384 10007 -8336
rect 34706 -8318 34716 -8262
rect 34772 -8318 34820 -8262
rect 34876 -8318 34924 -8262
rect 34980 -8318 35028 -8262
rect 35084 -8318 35132 -8262
rect 35188 -8318 35198 -8262
rect 34706 -8360 35198 -8318
rect 39146 -8054 39638 -8044
rect 39146 -8110 39156 -8054
rect 39212 -8110 39260 -8054
rect 39316 -8110 39364 -8054
rect 39420 -8110 39468 -8054
rect 39524 -8110 39572 -8054
rect 39628 -8110 39638 -8054
rect 39146 -8158 39638 -8110
rect 39146 -8214 39156 -8158
rect 39212 -8214 39260 -8158
rect 39316 -8214 39364 -8158
rect 39420 -8214 39468 -8158
rect 39524 -8214 39572 -8158
rect 39628 -8214 39638 -8158
rect 39146 -8262 39638 -8214
rect 39146 -8318 39156 -8262
rect 39212 -8318 39260 -8262
rect 39316 -8318 39364 -8262
rect 39420 -8318 39468 -8262
rect 39524 -8318 39572 -8262
rect 39628 -8318 39638 -8262
rect 39146 -8360 39638 -8318
rect 23632 -8366 39638 -8360
rect 23632 -8370 34716 -8366
rect 5134 -8440 5144 -8384
rect 5200 -8440 5248 -8384
rect 5304 -8440 9837 -8384
rect 9893 -8440 9941 -8384
rect 9997 -8440 10007 -8384
rect 5134 -8450 5314 -8440
rect 9827 -8450 10007 -8440
rect 14403 -8383 21429 -8373
rect 14403 -8439 14413 -8383
rect 14469 -8439 14517 -8383
rect 14573 -8439 14621 -8383
rect 14677 -8439 21155 -8383
rect 21211 -8439 21259 -8383
rect 21315 -8439 21363 -8383
rect 21419 -8439 21429 -8383
rect 14403 -8487 21429 -8439
rect 14403 -8543 14413 -8487
rect 14469 -8543 14517 -8487
rect 14573 -8543 14621 -8487
rect 14677 -8543 21155 -8487
rect 21211 -8543 21259 -8487
rect 21315 -8543 21363 -8487
rect 21419 -8543 21429 -8487
rect 4658 -8600 12894 -8590
rect 4658 -8656 4668 -8600
rect 4724 -8656 4772 -8600
rect 4828 -8656 12724 -8600
rect 12780 -8656 12828 -8600
rect 12884 -8656 12894 -8600
rect 4658 -8704 12894 -8656
rect 14403 -8591 21429 -8543
rect 14403 -8647 14413 -8591
rect 14469 -8647 14517 -8591
rect 14573 -8647 14621 -8591
rect 14677 -8647 21155 -8591
rect 21211 -8647 21259 -8591
rect 21315 -8647 21363 -8591
rect 21419 -8647 21429 -8591
rect 23632 -8426 23642 -8370
rect 23698 -8426 23746 -8370
rect 23802 -8426 30742 -8370
rect 30798 -8426 30846 -8370
rect 30902 -8426 30950 -8370
rect 31006 -8422 34716 -8370
rect 34772 -8422 34820 -8366
rect 34876 -8422 34924 -8366
rect 34980 -8422 35028 -8366
rect 35084 -8422 35132 -8366
rect 35188 -8422 39156 -8366
rect 39212 -8422 39260 -8366
rect 39316 -8422 39364 -8366
rect 39420 -8422 39468 -8366
rect 39524 -8422 39572 -8366
rect 39628 -8422 39638 -8366
rect 31006 -8426 39638 -8422
rect 23632 -8470 39638 -8426
rect 44536 -8058 45028 -8010
rect 44536 -8114 44546 -8058
rect 44602 -8114 44650 -8058
rect 44706 -8114 44754 -8058
rect 44810 -8114 44858 -8058
rect 44914 -8114 44962 -8058
rect 45018 -8114 45028 -8058
rect 44536 -8162 45028 -8114
rect 44536 -8218 44546 -8162
rect 44602 -8218 44650 -8162
rect 44706 -8218 44754 -8162
rect 44810 -8218 44858 -8162
rect 44914 -8218 44962 -8162
rect 45018 -8218 45028 -8162
rect 44536 -8266 45028 -8218
rect 44536 -8322 44546 -8266
rect 44602 -8322 44650 -8266
rect 44706 -8322 44754 -8266
rect 44810 -8322 44858 -8266
rect 44914 -8322 44962 -8266
rect 45018 -8322 45028 -8266
rect 44536 -8370 45028 -8322
rect 44536 -8426 44546 -8370
rect 44602 -8426 44650 -8370
rect 44706 -8426 44754 -8370
rect 44810 -8426 44858 -8370
rect 44914 -8426 44962 -8370
rect 45018 -8426 45028 -8370
rect 44536 -8436 45028 -8426
rect 48976 -7954 49468 -7944
rect 48976 -8010 48986 -7954
rect 49042 -8010 49090 -7954
rect 49146 -8010 49194 -7954
rect 49250 -8010 49298 -7954
rect 49354 -8010 49402 -7954
rect 49458 -8010 49468 -7954
rect 48976 -8058 49468 -8010
rect 48976 -8114 48986 -8058
rect 49042 -8114 49090 -8058
rect 49146 -8114 49194 -8058
rect 49250 -8114 49298 -8058
rect 49354 -8114 49402 -8058
rect 49458 -8114 49468 -8058
rect 48976 -8162 49468 -8114
rect 48976 -8218 48986 -8162
rect 49042 -8218 49090 -8162
rect 49146 -8218 49194 -8162
rect 49250 -8218 49298 -8162
rect 49354 -8218 49402 -8162
rect 49458 -8218 49468 -8162
rect 48976 -8266 49468 -8218
rect 48976 -8322 48986 -8266
rect 49042 -8322 49090 -8266
rect 49146 -8322 49194 -8266
rect 49250 -8322 49298 -8266
rect 49354 -8322 49402 -8266
rect 49458 -8322 49468 -8266
rect 48976 -8370 49468 -8322
rect 48976 -8426 48986 -8370
rect 49042 -8426 49090 -8370
rect 49146 -8426 49194 -8370
rect 49250 -8426 49298 -8370
rect 49354 -8426 49402 -8370
rect 49458 -8426 49468 -8370
rect 48976 -8436 49468 -8426
rect 23632 -8474 34716 -8470
rect 23632 -8530 23642 -8474
rect 23698 -8530 23746 -8474
rect 23802 -8530 30742 -8474
rect 30798 -8530 30846 -8474
rect 30902 -8530 30950 -8474
rect 31006 -8526 34716 -8474
rect 34772 -8526 34820 -8470
rect 34876 -8526 34924 -8470
rect 34980 -8526 35028 -8470
rect 35084 -8526 35132 -8470
rect 35188 -8526 39156 -8470
rect 39212 -8526 39260 -8470
rect 39316 -8526 39364 -8470
rect 39420 -8526 39468 -8470
rect 39524 -8526 39572 -8470
rect 39628 -8526 39638 -8470
rect 31006 -8530 39638 -8526
rect 23632 -8536 39638 -8530
rect 23632 -8578 39620 -8536
rect 23632 -8634 23642 -8578
rect 23698 -8634 23746 -8578
rect 23802 -8634 30742 -8578
rect 30798 -8634 30846 -8578
rect 30902 -8634 30950 -8578
rect 31006 -8634 39620 -8578
rect 23632 -8644 39620 -8634
rect 14403 -8657 21429 -8647
rect 4658 -8760 4668 -8704
rect 4724 -8760 4772 -8704
rect 4828 -8760 12724 -8704
rect 12780 -8760 12828 -8704
rect 12884 -8760 12894 -8704
rect 4658 -8770 12894 -8760
rect 44609 -8761 44893 -8436
rect 49090 -8761 49374 -8436
rect 18953 -8771 49499 -8761
rect 18953 -8827 18963 -8771
rect 19019 -8827 19067 -8771
rect 19123 -8827 19190 -8771
rect 19246 -8827 24092 -8771
rect 24148 -8827 24196 -8771
rect 24252 -8827 31650 -8771
rect 31706 -8827 31754 -8771
rect 31810 -8827 31858 -8771
rect 31914 -8827 49499 -8771
rect 18953 -8875 49499 -8827
rect 18953 -8931 18963 -8875
rect 19019 -8931 19067 -8875
rect 19123 -8931 19190 -8875
rect 19246 -8931 24092 -8875
rect 24148 -8931 24196 -8875
rect 24252 -8931 31650 -8875
rect 31706 -8931 31754 -8875
rect 31810 -8931 31858 -8875
rect 31914 -8931 49499 -8875
rect 18953 -8979 49499 -8931
rect 18953 -9035 18963 -8979
rect 19019 -9035 19067 -8979
rect 19123 -9035 19190 -8979
rect 19246 -9035 24092 -8979
rect 24148 -9035 24196 -8979
rect 24252 -9035 31650 -8979
rect 31706 -9035 31754 -8979
rect 31810 -9035 31858 -8979
rect 31914 -9035 49499 -8979
rect 18953 -9045 49499 -9035
rect 6825 -9391 54425 -9382
rect 6825 -9447 16967 -9391
rect 17023 -9447 17077 -9391
rect 17133 -9447 33967 -9391
rect 34023 -9447 34077 -9391
rect 34133 -9447 54233 -9391
rect 54289 -9447 54343 -9391
rect 54399 -9447 54425 -9391
rect 6825 -9501 54425 -9447
rect 6825 -9557 16967 -9501
rect 17023 -9557 17077 -9501
rect 17133 -9557 33967 -9501
rect 34023 -9557 34077 -9501
rect 34133 -9557 54233 -9501
rect 54289 -9557 54343 -9501
rect 54399 -9557 54425 -9501
rect 6825 -9562 54425 -9557
rect 6825 -9633 54644 -9624
rect 6825 -9689 14946 -9633
rect 15002 -9689 15056 -9633
rect 15112 -9689 31946 -9633
rect 32002 -9689 32056 -9633
rect 32112 -9689 54452 -9633
rect 54508 -9689 54562 -9633
rect 54618 -9689 54644 -9633
rect 6825 -9743 54644 -9689
rect 6825 -9799 14946 -9743
rect 15002 -9799 15056 -9743
rect 15112 -9799 31946 -9743
rect 32002 -9799 32056 -9743
rect 32112 -9799 54452 -9743
rect 54508 -9799 54562 -9743
rect 54618 -9799 54644 -9743
rect 6825 -9804 54644 -9799
rect 6825 -9875 54946 -9866
rect 6825 -9931 12983 -9875
rect 13039 -9931 13093 -9875
rect 13149 -9931 29983 -9875
rect 30039 -9931 30093 -9875
rect 30149 -9931 54754 -9875
rect 54810 -9931 54864 -9875
rect 54920 -9931 54946 -9875
rect 6825 -9985 54946 -9931
rect 6825 -10041 12983 -9985
rect 13039 -10041 13093 -9985
rect 13149 -10041 29983 -9985
rect 30039 -10041 30093 -9985
rect 30149 -10041 54754 -9985
rect 54810 -10041 54864 -9985
rect 54920 -10041 54946 -9985
rect 6825 -10046 54946 -10041
rect 6825 -10120 55182 -10111
rect 6825 -10176 10976 -10120
rect 11032 -10176 11086 -10120
rect 11142 -10176 27976 -10120
rect 28032 -10176 28086 -10120
rect 28142 -10176 54990 -10120
rect 55046 -10176 55100 -10120
rect 55156 -10176 55182 -10120
rect 6825 -10230 55182 -10176
rect 6825 -10286 10976 -10230
rect 11032 -10286 11086 -10230
rect 11142 -10286 27976 -10230
rect 28032 -10286 28086 -10230
rect 28142 -10286 54990 -10230
rect 55046 -10286 55100 -10230
rect 55156 -10286 55182 -10230
rect 6825 -10291 55182 -10286
rect 6825 -10356 55443 -10347
rect 6825 -10412 8941 -10356
rect 8997 -10412 9051 -10356
rect 9107 -10412 25941 -10356
rect 25997 -10412 26051 -10356
rect 26107 -10412 55251 -10356
rect 55307 -10412 55361 -10356
rect 55417 -10412 55443 -10356
rect 6825 -10466 55443 -10412
rect 6825 -10522 8941 -10466
rect 8997 -10522 9051 -10466
rect 9107 -10522 25941 -10466
rect 25997 -10522 26051 -10466
rect 26107 -10522 55251 -10466
rect 55307 -10522 55361 -10466
rect 55417 -10522 55443 -10466
rect 6825 -10527 55443 -10522
rect 55539 -10589 55760 -10588
rect 6825 -10597 55760 -10589
rect 6825 -10598 55568 -10597
rect 6825 -10654 6854 -10598
rect 6910 -10654 6964 -10598
rect 7020 -10654 23854 -10598
rect 23910 -10654 23964 -10598
rect 24020 -10653 55568 -10598
rect 55624 -10653 55678 -10597
rect 55734 -10653 55760 -10597
rect 24020 -10654 55760 -10653
rect 6825 -10707 55760 -10654
rect 6825 -10708 55568 -10707
rect 6825 -10764 6854 -10708
rect 6910 -10764 6964 -10708
rect 7020 -10764 23854 -10708
rect 23910 -10764 23964 -10708
rect 24020 -10763 55568 -10708
rect 55624 -10763 55678 -10707
rect 55734 -10763 55760 -10707
rect 24020 -10764 55760 -10763
rect 6825 -10768 55760 -10764
rect 6825 -10769 55748 -10768
rect -1790 -10933 35772 -10864
rect -1790 -10937 31453 -10933
rect -1790 -10947 29450 -10937
rect -1790 -10977 27397 -10947
rect -1790 -11017 25395 -10977
rect -1790 -11018 -1524 -11017
rect -1790 -11074 -1761 -11018
rect -1705 -11074 -1651 -11018
rect -1595 -11073 -1524 -11018
rect -1468 -11073 -1414 -11017
rect -1358 -11033 25395 -11017
rect 25451 -11033 25505 -10977
rect 25561 -11003 27397 -10977
rect 27453 -11003 27507 -10947
rect 27563 -10993 29450 -10947
rect 29506 -10993 29560 -10937
rect 29616 -10989 31453 -10937
rect 31509 -10989 31563 -10933
rect 31619 -10989 33506 -10933
rect 33562 -10989 33616 -10933
rect 33672 -10989 35557 -10933
rect 35613 -10989 35667 -10933
rect 35723 -10989 35772 -10933
rect 29616 -10993 35772 -10989
rect 27563 -11003 35772 -10993
rect 25561 -11033 35772 -11003
rect -1358 -11043 35772 -11033
rect -1358 -11047 31453 -11043
rect -1358 -11057 29450 -11047
rect -1358 -11073 27397 -11057
rect -1595 -11074 27397 -11073
rect -1790 -11087 27397 -11074
rect -1790 -11127 25395 -11087
rect -1790 -11128 -1524 -11127
rect -1790 -11184 -1761 -11128
rect -1705 -11184 -1651 -11128
rect -1595 -11183 -1524 -11128
rect -1468 -11183 -1414 -11127
rect -1358 -11143 25395 -11127
rect 25451 -11143 25505 -11087
rect 25561 -11113 27397 -11087
rect 27453 -11113 27507 -11057
rect 27563 -11103 29450 -11057
rect 29506 -11103 29560 -11047
rect 29616 -11099 31453 -11047
rect 31509 -11099 31563 -11043
rect 31619 -11099 33506 -11043
rect 33562 -11099 33616 -11043
rect 33672 -11099 35557 -11043
rect 35613 -11099 35667 -11043
rect 35723 -11099 35772 -11043
rect 29616 -11103 35772 -11099
rect 27563 -11113 35772 -11103
rect 25561 -11143 35772 -11113
rect -1358 -11183 35772 -11143
rect -1595 -11184 35772 -11183
rect -1790 -11189 35772 -11184
rect -1108 -11384 18656 -11288
rect -1108 -11387 18448 -11384
rect -1108 -11388 16458 -11387
rect -1108 -11397 14462 -11388
rect -1108 -11401 12428 -11397
rect -1108 -11425 10404 -11401
rect -1108 -11433 8401 -11425
rect -1115 -11442 8401 -11433
rect -1115 -11498 -1086 -11442
rect -1030 -11498 -976 -11442
rect -920 -11498 -858 -11442
rect -802 -11498 -748 -11442
rect -692 -11481 8401 -11442
rect 8457 -11481 8511 -11425
rect 8567 -11457 10404 -11425
rect 10460 -11457 10514 -11401
rect 10570 -11453 12428 -11401
rect 12484 -11453 12538 -11397
rect 12594 -11444 14462 -11397
rect 14518 -11444 14572 -11388
rect 14628 -11443 16458 -11388
rect 16514 -11443 16568 -11387
rect 16624 -11440 18448 -11387
rect 18504 -11440 18558 -11384
rect 18614 -11440 18656 -11384
rect 16624 -11443 18656 -11440
rect 14628 -11444 18656 -11443
rect 12594 -11453 18656 -11444
rect 10570 -11457 18656 -11453
rect 8567 -11481 18656 -11457
rect -692 -11494 18656 -11481
rect -692 -11497 18448 -11494
rect -692 -11498 16458 -11497
rect -1115 -11507 14462 -11498
rect -1115 -11511 12428 -11507
rect -1115 -11535 10404 -11511
rect -1115 -11552 8401 -11535
rect -1115 -11608 -1086 -11552
rect -1030 -11608 -976 -11552
rect -920 -11608 -858 -11552
rect -802 -11608 -748 -11552
rect -692 -11591 8401 -11552
rect 8457 -11591 8511 -11535
rect 8567 -11567 10404 -11535
rect 10460 -11567 10514 -11511
rect 10570 -11563 12428 -11511
rect 12484 -11563 12538 -11507
rect 12594 -11554 14462 -11507
rect 14518 -11554 14572 -11498
rect 14628 -11553 16458 -11498
rect 16514 -11553 16568 -11497
rect 16624 -11550 18448 -11497
rect 18504 -11550 18558 -11494
rect 18614 -11550 18656 -11494
rect 16624 -11553 18656 -11550
rect 14628 -11554 18656 -11553
rect 12594 -11563 18656 -11554
rect 10570 -11567 18656 -11563
rect 8567 -11591 18656 -11567
rect -692 -11608 18656 -11591
rect -1115 -11613 18656 -11608
rect 7127 -12960 17653 -12943
rect 7127 -13016 7132 -12960
rect 7188 -13016 7242 -12960
rect 7298 -13016 17445 -12960
rect 17501 -13016 17555 -12960
rect 17611 -13016 17653 -12960
rect 7127 -13037 17653 -13016
rect 24127 -12960 34653 -12943
rect 24127 -13016 24132 -12960
rect 24188 -13016 24242 -12960
rect 24298 -13016 34445 -12960
rect 34501 -13016 34555 -12960
rect 34611 -13016 34653 -12960
rect 24127 -13037 34653 -13016
rect 7083 -13110 17653 -13093
rect 7083 -13166 7088 -13110
rect 7144 -13166 7198 -13110
rect 7254 -13166 9156 -13110
rect 9212 -13166 9266 -13110
rect 9322 -13166 17653 -13110
rect 7083 -13187 17653 -13166
rect 24083 -13110 34653 -13093
rect 24083 -13166 24088 -13110
rect 24144 -13166 24198 -13110
rect 24254 -13166 26156 -13110
rect 26212 -13166 26266 -13110
rect 26322 -13166 34653 -13110
rect 24083 -13187 34653 -13166
rect 7270 -13260 17808 -13243
rect 7270 -13316 11176 -13260
rect 11232 -13316 11286 -13260
rect 11342 -13316 17628 -13260
rect 17684 -13316 17738 -13260
rect 17794 -13316 17808 -13260
rect 7270 -13337 17808 -13316
rect 24270 -13260 34808 -13243
rect 24270 -13316 28176 -13260
rect 28232 -13316 28286 -13260
rect 28342 -13316 34628 -13260
rect 34684 -13316 34738 -13260
rect 34794 -13316 34808 -13260
rect 24270 -13337 34808 -13316
rect 6699 -13410 17808 -13393
rect 6699 -13466 6704 -13410
rect 6760 -13466 6814 -13410
rect 6870 -13466 13166 -13410
rect 13222 -13466 13276 -13410
rect 13332 -13466 17808 -13410
rect 6699 -13487 17808 -13466
rect 23699 -13410 34808 -13393
rect 23699 -13466 23704 -13410
rect 23760 -13466 23814 -13410
rect 23870 -13466 30166 -13410
rect 30222 -13466 30276 -13410
rect 30332 -13466 34808 -13410
rect 23699 -13487 34808 -13466
rect 7270 -13560 18018 -13543
rect 7270 -13616 15193 -13560
rect 15249 -13616 15303 -13560
rect 15359 -13616 17785 -13560
rect 17841 -13616 17895 -13560
rect 17951 -13616 18018 -13560
rect 7270 -13637 18018 -13616
rect 24270 -13560 35018 -13543
rect 24270 -13616 32193 -13560
rect 32249 -13616 32303 -13560
rect 32359 -13616 34785 -13560
rect 34841 -13616 34895 -13560
rect 34951 -13616 35018 -13560
rect 24270 -13637 35018 -13616
rect 6459 -13710 18018 -13693
rect 6459 -13766 6464 -13710
rect 6520 -13766 6574 -13710
rect 6630 -13766 17122 -13710
rect 17178 -13766 17232 -13710
rect 17288 -13766 18018 -13710
rect 6459 -13787 18018 -13766
rect 23459 -13710 35018 -13693
rect 23459 -13766 23464 -13710
rect 23520 -13766 23574 -13710
rect 23630 -13766 34122 -13710
rect 34178 -13766 34232 -13710
rect 34288 -13766 35018 -13710
rect 23459 -13787 35018 -13766
<< via3 >>
rect 31598 -5074 31654 -5018
rect 31702 -5074 31758 -5018
rect 31806 -5074 31862 -5018
rect 31910 -5074 31966 -5018
rect 32014 -5074 32070 -5018
rect 31598 -5178 31654 -5122
rect 31702 -5178 31758 -5122
rect 31806 -5178 31862 -5122
rect 31910 -5178 31966 -5122
rect 32014 -5178 32070 -5122
rect 31598 -5282 31654 -5226
rect 31702 -5282 31758 -5226
rect 31806 -5282 31862 -5226
rect 31910 -5282 31966 -5226
rect 32014 -5282 32070 -5226
rect 31598 -5386 31654 -5330
rect 31702 -5386 31758 -5330
rect 31806 -5386 31862 -5330
rect 31910 -5386 31966 -5330
rect 32014 -5386 32070 -5330
rect 31598 -5490 31654 -5434
rect 31702 -5490 31758 -5434
rect 31806 -5490 31862 -5434
rect 31910 -5490 31966 -5434
rect 32014 -5490 32070 -5434
rect 42022 -7086 42078 -7030
rect 42126 -7086 42182 -7030
rect 42230 -7086 42286 -7030
rect 42022 -7190 42078 -7134
rect 42126 -7190 42182 -7134
rect 42230 -7190 42286 -7134
rect 42022 -7294 42078 -7238
rect 42126 -7294 42182 -7238
rect 42230 -7294 42286 -7238
rect 42022 -7398 42078 -7342
rect 42126 -7398 42182 -7342
rect 42230 -7398 42286 -7342
rect 42022 -7502 42078 -7446
rect 42126 -7502 42182 -7446
rect 42230 -7502 42286 -7446
rect 44546 -8010 44602 -7954
rect 44650 -8010 44706 -7954
rect 44754 -8010 44810 -7954
rect 44858 -8010 44914 -7954
rect 44962 -8010 45018 -7954
rect 34716 -8110 34772 -8054
rect 34820 -8110 34876 -8054
rect 34924 -8110 34980 -8054
rect 35028 -8110 35084 -8054
rect 35132 -8110 35188 -8054
rect 34716 -8214 34772 -8158
rect 34820 -8214 34876 -8158
rect 34924 -8214 34980 -8158
rect 35028 -8214 35084 -8158
rect 35132 -8214 35188 -8158
rect 34716 -8318 34772 -8262
rect 34820 -8318 34876 -8262
rect 34924 -8318 34980 -8262
rect 35028 -8318 35084 -8262
rect 35132 -8318 35188 -8262
rect 39156 -8110 39212 -8054
rect 39260 -8110 39316 -8054
rect 39364 -8110 39420 -8054
rect 39468 -8110 39524 -8054
rect 39572 -8110 39628 -8054
rect 39156 -8214 39212 -8158
rect 39260 -8214 39316 -8158
rect 39364 -8214 39420 -8158
rect 39468 -8214 39524 -8158
rect 39572 -8214 39628 -8158
rect 39156 -8318 39212 -8262
rect 39260 -8318 39316 -8262
rect 39364 -8318 39420 -8262
rect 39468 -8318 39524 -8262
rect 39572 -8318 39628 -8262
rect 34716 -8422 34772 -8366
rect 34820 -8422 34876 -8366
rect 34924 -8422 34980 -8366
rect 35028 -8422 35084 -8366
rect 35132 -8422 35188 -8366
rect 39156 -8422 39212 -8366
rect 39260 -8422 39316 -8366
rect 39364 -8422 39420 -8366
rect 39468 -8422 39524 -8366
rect 39572 -8422 39628 -8366
rect 44546 -8114 44602 -8058
rect 44650 -8114 44706 -8058
rect 44754 -8114 44810 -8058
rect 44858 -8114 44914 -8058
rect 44962 -8114 45018 -8058
rect 44546 -8218 44602 -8162
rect 44650 -8218 44706 -8162
rect 44754 -8218 44810 -8162
rect 44858 -8218 44914 -8162
rect 44962 -8218 45018 -8162
rect 44546 -8322 44602 -8266
rect 44650 -8322 44706 -8266
rect 44754 -8322 44810 -8266
rect 44858 -8322 44914 -8266
rect 44962 -8322 45018 -8266
rect 44546 -8426 44602 -8370
rect 44650 -8426 44706 -8370
rect 44754 -8426 44810 -8370
rect 44858 -8426 44914 -8370
rect 44962 -8426 45018 -8370
rect 48986 -8010 49042 -7954
rect 49090 -8010 49146 -7954
rect 49194 -8010 49250 -7954
rect 49298 -8010 49354 -7954
rect 49402 -8010 49458 -7954
rect 48986 -8114 49042 -8058
rect 49090 -8114 49146 -8058
rect 49194 -8114 49250 -8058
rect 49298 -8114 49354 -8058
rect 49402 -8114 49458 -8058
rect 48986 -8218 49042 -8162
rect 49090 -8218 49146 -8162
rect 49194 -8218 49250 -8162
rect 49298 -8218 49354 -8162
rect 49402 -8218 49458 -8162
rect 48986 -8322 49042 -8266
rect 49090 -8322 49146 -8266
rect 49194 -8322 49250 -8266
rect 49298 -8322 49354 -8266
rect 49402 -8322 49458 -8266
rect 48986 -8426 49042 -8370
rect 49090 -8426 49146 -8370
rect 49194 -8426 49250 -8370
rect 49298 -8426 49354 -8370
rect 49402 -8426 49458 -8370
rect 34716 -8526 34772 -8470
rect 34820 -8526 34876 -8470
rect 34924 -8526 34980 -8470
rect 35028 -8526 35084 -8470
rect 35132 -8526 35188 -8470
rect 39156 -8526 39212 -8470
rect 39260 -8526 39316 -8470
rect 39364 -8526 39420 -8470
rect 39468 -8526 39524 -8470
rect 39572 -8526 39628 -8470
<< metal4 >>
rect 31588 -5018 32080 -5008
rect 31588 -5074 31598 -5018
rect 31654 -5074 31702 -5018
rect 31758 -5074 31806 -5018
rect 31862 -5074 31910 -5018
rect 31966 -5074 32014 -5018
rect 32070 -5074 32080 -5018
rect 31588 -5122 32080 -5074
rect 31588 -5178 31598 -5122
rect 31654 -5178 31702 -5122
rect 31758 -5178 31806 -5122
rect 31862 -5178 31910 -5122
rect 31966 -5178 32014 -5122
rect 32070 -5178 32080 -5122
rect 31588 -5226 32080 -5178
rect 31588 -5282 31598 -5226
rect 31654 -5282 31702 -5226
rect 31758 -5282 31806 -5226
rect 31862 -5282 31910 -5226
rect 31966 -5282 32014 -5226
rect 32070 -5282 32080 -5226
rect 31588 -5330 32080 -5282
rect 31588 -5386 31598 -5330
rect 31654 -5386 31702 -5330
rect 31758 -5386 31806 -5330
rect 31862 -5386 31910 -5330
rect 31966 -5386 32014 -5330
rect 32070 -5386 32080 -5330
rect 31588 -5434 32080 -5386
rect 31588 -5490 31598 -5434
rect 31654 -5490 31702 -5434
rect 31758 -5490 31806 -5434
rect 31862 -5490 31910 -5434
rect 31966 -5490 32014 -5434
rect 32070 -5490 32080 -5434
rect 31588 -5500 32080 -5490
rect 41977 -5018 42321 -5008
rect 41977 -5074 42022 -5018
rect 42078 -5074 42126 -5018
rect 42182 -5074 42230 -5018
rect 42286 -5074 42321 -5018
rect 41977 -5122 42321 -5074
rect 41977 -5178 42022 -5122
rect 42078 -5178 42126 -5122
rect 42182 -5178 42230 -5122
rect 42286 -5178 42321 -5122
rect 41977 -5226 42321 -5178
rect 41977 -5282 42022 -5226
rect 42078 -5282 42126 -5226
rect 42182 -5282 42230 -5226
rect 42286 -5282 42321 -5226
rect 41977 -5330 42321 -5282
rect 41977 -5386 42022 -5330
rect 42078 -5386 42126 -5330
rect 42182 -5386 42230 -5330
rect 42286 -5386 42321 -5330
rect 41977 -5434 42321 -5386
rect 41977 -5490 42022 -5434
rect 42078 -5490 42126 -5434
rect 42182 -5490 42230 -5434
rect 42286 -5490 42321 -5434
rect 41977 -7030 42321 -5490
rect 41977 -7086 42022 -7030
rect 42078 -7086 42126 -7030
rect 42182 -7086 42230 -7030
rect 42286 -7086 42321 -7030
rect 41977 -7134 42321 -7086
rect 41977 -7190 42022 -7134
rect 42078 -7190 42126 -7134
rect 42182 -7190 42230 -7134
rect 42286 -7190 42321 -7134
rect 41977 -7238 42321 -7190
rect 41977 -7294 42022 -7238
rect 42078 -7294 42126 -7238
rect 42182 -7294 42230 -7238
rect 42286 -7294 42321 -7238
rect 41977 -7342 42321 -7294
rect 41977 -7398 42022 -7342
rect 42078 -7398 42126 -7342
rect 42182 -7398 42230 -7342
rect 42286 -7398 42321 -7342
rect 41977 -7446 42321 -7398
rect 41977 -7502 42022 -7446
rect 42078 -7502 42126 -7446
rect 42182 -7502 42230 -7446
rect 42286 -7502 42321 -7446
rect 41977 -7512 42321 -7502
rect 34706 -8054 35198 -7642
rect 34706 -8110 34716 -8054
rect 34772 -8110 34820 -8054
rect 34876 -8110 34924 -8054
rect 34980 -8110 35028 -8054
rect 35084 -8110 35132 -8054
rect 35188 -8110 35198 -8054
rect 34706 -8158 35198 -8110
rect 34706 -8214 34716 -8158
rect 34772 -8214 34820 -8158
rect 34876 -8214 34924 -8158
rect 34980 -8214 35028 -8158
rect 35084 -8214 35132 -8158
rect 35188 -8214 35198 -8158
rect 34706 -8262 35198 -8214
rect 34706 -8318 34716 -8262
rect 34772 -8318 34820 -8262
rect 34876 -8318 34924 -8262
rect 34980 -8318 35028 -8262
rect 35084 -8318 35132 -8262
rect 35188 -8318 35198 -8262
rect 34706 -8366 35198 -8318
rect 34706 -8422 34716 -8366
rect 34772 -8422 34820 -8366
rect 34876 -8422 34924 -8366
rect 34980 -8422 35028 -8366
rect 35084 -8422 35132 -8366
rect 35188 -8422 35198 -8366
rect 34706 -8470 35198 -8422
rect 34706 -8526 34716 -8470
rect 34772 -8526 34820 -8470
rect 34876 -8526 34924 -8470
rect 34980 -8526 35028 -8470
rect 35084 -8526 35132 -8470
rect 35188 -8526 35198 -8470
rect 34706 -8536 35198 -8526
rect 39146 -8054 39638 -7679
rect 39146 -8110 39156 -8054
rect 39212 -8110 39260 -8054
rect 39316 -8110 39364 -8054
rect 39420 -8110 39468 -8054
rect 39524 -8110 39572 -8054
rect 39628 -8110 39638 -8054
rect 39146 -8158 39638 -8110
rect 39146 -8214 39156 -8158
rect 39212 -8214 39260 -8158
rect 39316 -8214 39364 -8158
rect 39420 -8214 39468 -8158
rect 39524 -8214 39572 -8158
rect 39628 -8214 39638 -8158
rect 39146 -8262 39638 -8214
rect 39146 -8318 39156 -8262
rect 39212 -8318 39260 -8262
rect 39316 -8318 39364 -8262
rect 39420 -8318 39468 -8262
rect 39524 -8318 39572 -8262
rect 39628 -8318 39638 -8262
rect 39146 -8366 39638 -8318
rect 39146 -8422 39156 -8366
rect 39212 -8422 39260 -8366
rect 39316 -8422 39364 -8366
rect 39420 -8422 39468 -8366
rect 39524 -8422 39572 -8366
rect 39628 -8422 39638 -8366
rect 39146 -8470 39638 -8422
rect 44536 -7954 45028 -7704
rect 44536 -8010 44546 -7954
rect 44602 -8010 44650 -7954
rect 44706 -8010 44754 -7954
rect 44810 -8010 44858 -7954
rect 44914 -8010 44962 -7954
rect 45018 -8010 45028 -7954
rect 44536 -8058 45028 -8010
rect 44536 -8114 44546 -8058
rect 44602 -8114 44650 -8058
rect 44706 -8114 44754 -8058
rect 44810 -8114 44858 -8058
rect 44914 -8114 44962 -8058
rect 45018 -8114 45028 -8058
rect 44536 -8162 45028 -8114
rect 44536 -8218 44546 -8162
rect 44602 -8218 44650 -8162
rect 44706 -8218 44754 -8162
rect 44810 -8218 44858 -8162
rect 44914 -8218 44962 -8162
rect 45018 -8218 45028 -8162
rect 44536 -8266 45028 -8218
rect 44536 -8322 44546 -8266
rect 44602 -8322 44650 -8266
rect 44706 -8322 44754 -8266
rect 44810 -8322 44858 -8266
rect 44914 -8322 44962 -8266
rect 45018 -8322 45028 -8266
rect 44536 -8370 45028 -8322
rect 44536 -8426 44546 -8370
rect 44602 -8426 44650 -8370
rect 44706 -8426 44754 -8370
rect 44810 -8426 44858 -8370
rect 44914 -8426 44962 -8370
rect 45018 -8426 45028 -8370
rect 44536 -8436 45028 -8426
rect 48976 -7954 49468 -7704
rect 48976 -8010 48986 -7954
rect 49042 -8010 49090 -7954
rect 49146 -8010 49194 -7954
rect 49250 -8010 49298 -7954
rect 49354 -8010 49402 -7954
rect 49458 -8010 49468 -7954
rect 48976 -8058 49468 -8010
rect 48976 -8114 48986 -8058
rect 49042 -8114 49090 -8058
rect 49146 -8114 49194 -8058
rect 49250 -8114 49298 -8058
rect 49354 -8114 49402 -8058
rect 49458 -8114 49468 -8058
rect 48976 -8162 49468 -8114
rect 48976 -8218 48986 -8162
rect 49042 -8218 49090 -8162
rect 49146 -8218 49194 -8162
rect 49250 -8218 49298 -8162
rect 49354 -8218 49402 -8162
rect 49458 -8218 49468 -8162
rect 48976 -8266 49468 -8218
rect 48976 -8322 48986 -8266
rect 49042 -8322 49090 -8266
rect 49146 -8322 49194 -8266
rect 49250 -8322 49298 -8266
rect 49354 -8322 49402 -8266
rect 49458 -8322 49468 -8266
rect 48976 -8370 49468 -8322
rect 48976 -8426 48986 -8370
rect 49042 -8426 49090 -8370
rect 49146 -8426 49194 -8370
rect 49250 -8426 49298 -8370
rect 49354 -8426 49402 -8370
rect 49458 -8426 49468 -8370
rect 48976 -8436 49468 -8426
rect 39146 -8526 39156 -8470
rect 39212 -8526 39260 -8470
rect 39316 -8526 39364 -8470
rect 39420 -8526 39468 -8470
rect 39524 -8526 39572 -8470
rect 39628 -8526 39638 -8470
rect 39146 -8536 39638 -8526
<< via4 >>
rect 31598 -5074 31654 -5018
rect 31702 -5074 31758 -5018
rect 31806 -5074 31862 -5018
rect 31910 -5074 31966 -5018
rect 32014 -5074 32070 -5018
rect 31598 -5178 31654 -5122
rect 31702 -5178 31758 -5122
rect 31806 -5178 31862 -5122
rect 31910 -5178 31966 -5122
rect 32014 -5178 32070 -5122
rect 31598 -5282 31654 -5226
rect 31702 -5282 31758 -5226
rect 31806 -5282 31862 -5226
rect 31910 -5282 31966 -5226
rect 32014 -5282 32070 -5226
rect 31598 -5386 31654 -5330
rect 31702 -5386 31758 -5330
rect 31806 -5386 31862 -5330
rect 31910 -5386 31966 -5330
rect 32014 -5386 32070 -5330
rect 31598 -5490 31654 -5434
rect 31702 -5490 31758 -5434
rect 31806 -5490 31862 -5434
rect 31910 -5490 31966 -5434
rect 32014 -5490 32070 -5434
rect 42022 -5074 42078 -5018
rect 42126 -5074 42182 -5018
rect 42230 -5074 42286 -5018
rect 42022 -5178 42078 -5122
rect 42126 -5178 42182 -5122
rect 42230 -5178 42286 -5122
rect 42022 -5282 42078 -5226
rect 42126 -5282 42182 -5226
rect 42230 -5282 42286 -5226
rect 42022 -5386 42078 -5330
rect 42126 -5386 42182 -5330
rect 42230 -5386 42286 -5330
rect 42022 -5490 42078 -5434
rect 42126 -5490 42182 -5434
rect 42230 -5490 42286 -5434
rect 42022 -7086 42078 -7030
rect 42126 -7086 42182 -7030
rect 42230 -7086 42286 -7030
rect 42022 -7190 42078 -7134
rect 42126 -7190 42182 -7134
rect 42230 -7190 42286 -7134
rect 42022 -7294 42078 -7238
rect 42126 -7294 42182 -7238
rect 42230 -7294 42286 -7238
rect 42022 -7398 42078 -7342
rect 42126 -7398 42182 -7342
rect 42230 -7398 42286 -7342
rect 42022 -7502 42078 -7446
rect 42126 -7502 42182 -7446
rect 42230 -7502 42286 -7446
<< metal5 >>
rect 31588 -5018 32812 -5008
rect 31588 -5074 31598 -5018
rect 31654 -5074 31702 -5018
rect 31758 -5074 31806 -5018
rect 31862 -5074 31910 -5018
rect 31966 -5074 32014 -5018
rect 32070 -5074 32812 -5018
rect 31588 -5122 32812 -5074
rect 31588 -5178 31598 -5122
rect 31654 -5178 31702 -5122
rect 31758 -5178 31806 -5122
rect 31862 -5178 31910 -5122
rect 31966 -5178 32014 -5122
rect 32070 -5178 32812 -5122
rect 31588 -5226 32812 -5178
rect 31588 -5282 31598 -5226
rect 31654 -5282 31702 -5226
rect 31758 -5282 31806 -5226
rect 31862 -5282 31910 -5226
rect 31966 -5282 32014 -5226
rect 32070 -5282 32812 -5226
rect 31588 -5330 32812 -5282
rect 31588 -5386 31598 -5330
rect 31654 -5386 31702 -5330
rect 31758 -5386 31806 -5330
rect 31862 -5386 31910 -5330
rect 31966 -5386 32014 -5330
rect 32070 -5386 32812 -5330
rect 31588 -5434 32812 -5386
rect 31588 -5490 31598 -5434
rect 31654 -5490 31702 -5434
rect 31758 -5490 31806 -5434
rect 31862 -5490 31910 -5434
rect 31966 -5490 32014 -5434
rect 32070 -5490 32812 -5434
rect 31588 -5500 32812 -5490
rect 41977 -5018 42642 -5008
rect 41977 -5074 42022 -5018
rect 42078 -5074 42126 -5018
rect 42182 -5074 42230 -5018
rect 42286 -5074 42642 -5018
rect 41977 -5122 42642 -5074
rect 41977 -5178 42022 -5122
rect 42078 -5178 42126 -5122
rect 42182 -5178 42230 -5122
rect 42286 -5178 42642 -5122
rect 41977 -5226 42642 -5178
rect 41977 -5282 42022 -5226
rect 42078 -5282 42126 -5226
rect 42182 -5282 42230 -5226
rect 42286 -5282 42642 -5226
rect 41977 -5330 42642 -5282
rect 41977 -5386 42022 -5330
rect 42078 -5386 42126 -5330
rect 42182 -5386 42230 -5330
rect 42286 -5386 42642 -5330
rect 41977 -5434 42642 -5386
rect 41977 -5490 42022 -5434
rect 42078 -5490 42126 -5434
rect 42182 -5490 42230 -5434
rect 42286 -5490 42642 -5434
rect 41977 -5500 42642 -5490
rect 41977 -7030 42321 -7020
rect 41977 -7086 42022 -7030
rect 42078 -7086 42126 -7030
rect 42182 -7086 42230 -7030
rect 42286 -7086 42321 -7030
rect 41977 -7134 42321 -7086
rect 41977 -7190 42022 -7134
rect 42078 -7190 42126 -7134
rect 42182 -7190 42230 -7134
rect 42286 -7190 42321 -7134
rect 41977 -7238 42321 -7190
rect 41977 -7294 42022 -7238
rect 42078 -7294 42126 -7238
rect 42182 -7294 42230 -7238
rect 42286 -7294 42321 -7238
rect 41977 -7342 42321 -7294
rect 41977 -7398 42022 -7342
rect 42078 -7398 42126 -7342
rect 42182 -7398 42230 -7342
rect 42286 -7398 42321 -7342
rect 41977 -7446 42321 -7398
rect 41977 -7502 42022 -7446
rect 42078 -7502 42126 -7446
rect 42182 -7502 42230 -7446
rect 42286 -7502 42321 -7446
rect 41977 -7512 42321 -7502
use cap_mim_2p0fF_3FUNHB  cap_mim_2p0fF_3FUNHB_0
timestamp 1699631467
transform 0 1 37232 -1 0 -5364
box -2340 -4560 2340 4560
use cap_mim_2p0fF_3FUNHB  cap_mim_2p0fF_3FUNHB_1
timestamp 1699631467
transform 0 1 47062 -1 0 -5364
box -2340 -4560 2340 4560
use nmos_3p3_2F3WC4  nmos_3p3_2F3WC4_0
timestamp 1694939250
transform 1 0 15364 0 1 -5844
box -820 -536 820 536
use nmos_3p3_2F3WC4  nmos_3p3_2F3WC4_1
timestamp 1694939250
transform 1 0 13716 0 1 -5844
box -820 -536 820 536
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_0
timestamp 1693995983
transform 1 0 5766 0 1 -6828
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_1
timestamp 1693995983
transform 1 0 10278 0 1 -6828
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_2
timestamp 1693995983
transform 1 0 5766 0 1 -7465
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_3
timestamp 1693995983
transform 1 0 7301 0 1 -5663
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_4
timestamp 1693995983
transform 1 0 7013 0 1 -5663
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_5
timestamp 1693995983
transform 1 0 8741 0 1 -5663
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_6
timestamp 1693995983
transform 1 0 9029 0 1 -5663
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_7
timestamp 1693995983
transform 1 0 7013 0 1 -6199
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_8
timestamp 1693995983
transform 1 0 7301 0 1 -6199
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_9
timestamp 1693995983
transform 1 0 9029 0 1 -6199
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_10
timestamp 1693995983
transform 1 0 8741 0 1 -6199
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_11
timestamp 1693995983
transform 1 0 7301 0 1 -4591
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_12
timestamp 1693995983
transform 1 0 7013 0 1 -4591
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_13
timestamp 1693995983
transform 1 0 8741 0 1 -5127
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_14
timestamp 1693995983
transform 1 0 9029 0 1 -5127
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_15
timestamp 1693995983
transform 1 0 7301 0 1 -5127
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_16
timestamp 1693995983
transform 1 0 7013 0 1 -5127
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_17
timestamp 1693995983
transform 1 0 8741 0 1 -4591
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_18
timestamp 1693995983
transform 1 0 9029 0 1 -4591
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_19
timestamp 1693995983
transform 1 0 7301 0 1 -3519
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_20
timestamp 1693995983
transform 1 0 7013 0 1 -3519
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_21
timestamp 1693995983
transform 1 0 8741 0 1 -3519
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_22
timestamp 1693995983
transform 1 0 9029 0 1 -3519
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_23
timestamp 1693995983
transform 1 0 7301 0 1 -4055
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_24
timestamp 1693995983
transform 1 0 7013 0 1 -4055
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_25
timestamp 1693995983
transform 1 0 9029 0 1 -4055
box -140 -168 140 168
use nmos_3p3_3A6RT2  nmos_3p3_3A6RT2_26
timestamp 1693995983
transform 1 0 8741 0 1 -4055
box -140 -168 140 168
use nmos_3p3_3AEFT2  nmos_3p3_3AEFT2_0
timestamp 1693898117
transform 1 0 8026 0 1 -7465
box -168 -168 168 168
use nmos_3p3_5J7TC4  nmos_3p3_5J7TC4_0
timestamp 1693899127
transform 1 0 9286 0 1 -6828
box -364 -168 364 168
use nmos_3p3_5J7TC4  nmos_3p3_5J7TC4_1
timestamp 1693899127
transform 1 0 9894 0 1 -6828
box -364 -168 364 168
use nmos_3p3_6F3WC4  nmos_3p3_6F3WC4_0
timestamp 1694939532
transform 1 0 12372 0 1 -5844
box -212 -536 212 536
use nmos_3p3_6F3WC4  nmos_3p3_6F3WC4_1
timestamp 1694939532
transform 1 0 16276 0 1 -5844
box -212 -536 212 536
use nmos_3p3_6F3WC4  nmos_3p3_6F3WC4_2
timestamp 1694939532
transform 1 0 12804 0 1 -5844
box -212 -536 212 536
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_0
timestamp 1693069569
transform 1 0 9866 0 1 1364
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_1
timestamp 1693069569
transform 1 0 8970 0 1 1364
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_2
timestamp 1693069569
transform 1 0 9418 0 1 1364
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_3
timestamp 1693069569
transform 1 0 9866 0 1 -1222
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_4
timestamp 1693069569
transform 1 0 9418 0 1 -1222
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_5
timestamp 1693069569
transform 1 0 8970 0 1 -1222
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_6
timestamp 1693069569
transform 1 0 8970 0 1 -360
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_7
timestamp 1693069569
transform 1 0 9418 0 1 -360
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_8
timestamp 1693069569
transform 1 0 9866 0 1 -360
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_9
timestamp 1693069569
transform 1 0 8970 0 1 502
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_10
timestamp 1693069569
transform 1 0 9418 0 1 502
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_11
timestamp 1693069569
transform 1 0 9866 0 1 502
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_12
timestamp 1693069569
transform 1 0 7247 0 1 -341
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_13
timestamp 1693069569
transform 1 0 6607 0 1 -341
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_14
timestamp 1693069569
transform 1 0 6927 0 1 -341
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_15
timestamp 1693069569
transform 1 0 7247 0 1 -1203
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_16
timestamp 1693069569
transform 1 0 6927 0 1 -1203
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_17
timestamp 1693069569
transform 1 0 6607 0 1 -1203
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_18
timestamp 1693069569
transform 1 0 6607 0 1 521
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_19
timestamp 1693069569
transform 1 0 6927 0 1 521
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_20
timestamp 1693069569
transform 1 0 7247 0 1 521
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_21
timestamp 1693069569
transform 1 0 6607 0 1 2245
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_22
timestamp 1693069569
transform 1 0 6927 0 1 2245
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_23
timestamp 1693069569
transform 1 0 7247 0 1 2245
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_24
timestamp 1693069569
transform 1 0 6607 0 1 1383
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_25
timestamp 1693069569
transform 1 0 6927 0 1 1383
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_26
timestamp 1693069569
transform 1 0 7247 0 1 1383
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_27
timestamp 1693069569
transform 1 0 6607 0 1 3107
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_28
timestamp 1693069569
transform 1 0 6927 0 1 3107
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_29
timestamp 1693069569
transform 1 0 7247 0 1 3107
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_30
timestamp 1693069569
transform 1 0 6607 0 1 3969
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_31
timestamp 1693069569
transform 1 0 6927 0 1 3969
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_32
timestamp 1693069569
transform 1 0 7247 0 1 3969
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_33
timestamp 1693069569
transform 1 0 6607 0 1 4831
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_34
timestamp 1693069569
transform 1 0 6927 0 1 4831
box -220 -356 220 356
use nmos_3p3_7WQWW2  nmos_3p3_7WQWW2_35
timestamp 1693069569
transform 1 0 7247 0 1 4831
box -220 -356 220 356
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_0
timestamp 1694765150
transform 1 0 19497 0 1 924
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_1
timestamp 1694765150
transform 1 0 18857 0 1 924
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_2
timestamp 1694765150
transform 1 0 19177 0 1 924
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_3
timestamp 1694765150
transform 1 0 19497 0 1 -948
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_4
timestamp 1694765150
transform 1 0 19177 0 1 -948
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_5
timestamp 1694765150
transform 1 0 18857 0 1 -948
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_6
timestamp 1694765150
transform 1 0 18857 0 1 -12
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_7
timestamp 1694765150
transform 1 0 19177 0 1 -12
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_8
timestamp 1694765150
transform 1 0 19497 0 1 -12
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_9
timestamp 1694765150
transform 1 0 18857 0 1 1860
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_10
timestamp 1694765150
transform 1 0 19177 0 1 1860
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_11
timestamp 1694765150
transform 1 0 19497 0 1 1860
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_12
timestamp 1694765150
transform 1 0 18857 0 1 3732
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_13
timestamp 1694765150
transform 1 0 19177 0 1 3732
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_14
timestamp 1694765150
transform 1 0 19497 0 1 3732
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_15
timestamp 1694765150
transform 1 0 18857 0 1 2796
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_16
timestamp 1694765150
transform 1 0 19177 0 1 2796
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_17
timestamp 1694765150
transform 1 0 19497 0 1 2796
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_18
timestamp 1694765150
transform -1 0 24009 0 1 1860
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_19
timestamp 1694765150
transform -1 0 24649 0 1 1860
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_20
timestamp 1694765150
transform -1 0 24329 0 1 1860
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_21
timestamp 1694765150
transform -1 0 24009 0 1 924
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_22
timestamp 1694765150
transform -1 0 24649 0 1 924
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_23
timestamp 1694765150
transform -1 0 24329 0 1 924
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_24
timestamp 1694765150
transform -1 0 24009 0 1 -12
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_25
timestamp 1694765150
transform -1 0 24649 0 1 -12
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_26
timestamp 1694765150
transform -1 0 24329 0 1 -12
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_27
timestamp 1694765150
transform -1 0 24009 0 1 -948
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_28
timestamp 1694765150
transform -1 0 24329 0 1 -948
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_29
timestamp 1694765150
transform -1 0 24649 0 1 -948
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_30
timestamp 1694765150
transform -1 0 24329 0 1 3732
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_31
timestamp 1694765150
transform -1 0 24009 0 1 3732
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_32
timestamp 1694765150
transform -1 0 24649 0 1 3732
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_33
timestamp 1694765150
transform -1 0 24329 0 1 2796
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_34
timestamp 1694765150
transform -1 0 24009 0 1 2796
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_35
timestamp 1694765150
transform -1 0 24649 0 1 2796
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_36
timestamp 1694765150
transform 1 0 28618 0 1 1860
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_37
timestamp 1694765150
transform 1 0 27978 0 1 1860
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_38
timestamp 1694765150
transform 1 0 28298 0 1 1860
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_39
timestamp 1694765150
transform 1 0 28618 0 1 924
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_40
timestamp 1694765150
transform 1 0 27978 0 1 924
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_41
timestamp 1694765150
transform 1 0 28298 0 1 924
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_42
timestamp 1694765150
transform 1 0 28618 0 1 -12
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_43
timestamp 1694765150
transform 1 0 27978 0 1 -12
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_44
timestamp 1694765150
transform 1 0 28298 0 1 -12
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_45
timestamp 1694765150
transform 1 0 28618 0 1 -948
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_46
timestamp 1694765150
transform 1 0 28298 0 1 -948
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_47
timestamp 1694765150
transform 1 0 27978 0 1 -948
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_48
timestamp 1694765150
transform 1 0 28298 0 1 3732
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_49
timestamp 1694765150
transform 1 0 28618 0 1 3732
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_50
timestamp 1694765150
transform 1 0 27978 0 1 3732
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_51
timestamp 1694765150
transform 1 0 28298 0 1 2796
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_52
timestamp 1694765150
transform 1 0 28618 0 1 2796
box -220 -368 220 368
use nmos_3p3_276RTJ  nmos_3p3_276RTJ_53
timestamp 1694765150
transform 1 0 27978 0 1 2796
box -220 -368 220 368
use nmos_3p3_876RT2  nmos_3p3_876RT2_0
timestamp 1693995983
transform 1 0 7541 0 1 -5663
box -220 -168 220 168
use nmos_3p3_876RT2  nmos_3p3_876RT2_1
timestamp 1693995983
transform 1 0 8501 0 1 -5663
box -220 -168 220 168
use nmos_3p3_876RT2  nmos_3p3_876RT2_2
timestamp 1693995983
transform 1 0 7541 0 1 -6199
box -220 -168 220 168
use nmos_3p3_876RT2  nmos_3p3_876RT2_3
timestamp 1693995983
transform 1 0 8501 0 1 -6199
box -220 -168 220 168
use nmos_3p3_876RT2  nmos_3p3_876RT2_4
timestamp 1693995983
transform 1 0 7541 0 1 -4591
box -220 -168 220 168
use nmos_3p3_876RT2  nmos_3p3_876RT2_5
timestamp 1693995983
transform 1 0 8501 0 1 -5127
box -220 -168 220 168
use nmos_3p3_876RT2  nmos_3p3_876RT2_6
timestamp 1693995983
transform 1 0 7541 0 1 -5127
box -220 -168 220 168
use nmos_3p3_876RT2  nmos_3p3_876RT2_7
timestamp 1693995983
transform 1 0 8501 0 1 -4591
box -220 -168 220 168
use nmos_3p3_876RT2  nmos_3p3_876RT2_8
timestamp 1693995983
transform 1 0 7541 0 1 -3519
box -220 -168 220 168
use nmos_3p3_876RT2  nmos_3p3_876RT2_9
timestamp 1693995983
transform 1 0 8501 0 1 -3519
box -220 -168 220 168
use nmos_3p3_876RT2  nmos_3p3_876RT2_10
timestamp 1693995983
transform 1 0 7541 0 1 -4055
box -220 -168 220 168
use nmos_3p3_876RT2  nmos_3p3_876RT2_11
timestamp 1693995983
transform 1 0 8501 0 1 -4055
box -220 -168 220 168
use nmos_3p3_BSHHD6  nmos_3p3_BSHHD6_0
timestamp 1693895011
transform 1 0 6838 0 1 -7465
box -708 -168 708 168
use nmos_3p3_EA6RT2  nmos_3p3_EA6RT2_0
timestamp 1693995983
transform 1 0 6294 0 1 -6828
box -380 -168 380 168
use nmos_3p3_EA6RT2  nmos_3p3_EA6RT2_1
timestamp 1693995983
transform 1 0 8021 0 1 -5663
box -380 -168 380 168
use nmos_3p3_EA6RT2  nmos_3p3_EA6RT2_2
timestamp 1693995983
transform 1 0 8021 0 1 -6199
box -380 -168 380 168
use nmos_3p3_EA6RT2  nmos_3p3_EA6RT2_3
timestamp 1693995983
transform 1 0 8021 0 1 -5127
box -380 -168 380 168
use nmos_3p3_EA6RT2  nmos_3p3_EA6RT2_4
timestamp 1693995983
transform 1 0 8021 0 1 -4591
box -380 -168 380 168
use nmos_3p3_EA6RT2  nmos_3p3_EA6RT2_5
timestamp 1693995983
transform 1 0 8021 0 1 -3519
box -380 -168 380 168
use nmos_3p3_EA6RT2  nmos_3p3_EA6RT2_6
timestamp 1693995983
transform 1 0 8021 0 1 -4055
box -380 -168 380 168
use nmos_3p3_FSHHD6  nmos_3p3_FSHHD6_0
timestamp 1693895011
transform 1 0 7702 0 1 -7465
box -276 -168 276 168
use nmos_3p3_JE3WC4  nmos_3p3_JE3WC4_0
timestamp 1694938948
transform 1 0 15364 0 1 -6948
box -820 -268 820 268
use nmos_3p3_JE3WC4  nmos_3p3_JE3WC4_1
timestamp 1694938948
transform 1 0 13716 0 1 -6948
box -820 -268 820 268
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_0
timestamp 1694765150
transform 1 0 18617 0 1 924
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_1
timestamp 1694765150
transform 1 0 20025 0 1 1860
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_2
timestamp 1694765150
transform 1 0 18329 0 1 924
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_3
timestamp 1694765150
transform 1 0 19737 0 1 1860
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_4
timestamp 1694765150
transform 1 0 20025 0 1 -948
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_5
timestamp 1694765150
transform 1 0 19737 0 1 -948
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_6
timestamp 1694765150
transform 1 0 18617 0 1 -948
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_7
timestamp 1694765150
transform 1 0 18329 0 1 -948
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_8
timestamp 1694765150
transform 1 0 18329 0 1 -12
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_9
timestamp 1694765150
transform 1 0 18617 0 1 -12
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_10
timestamp 1694765150
transform 1 0 19737 0 1 -12
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_11
timestamp 1694765150
transform 1 0 20025 0 1 -12
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_12
timestamp 1694765150
transform 1 0 18329 0 1 1860
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_13
timestamp 1694765150
transform 1 0 18617 0 1 1860
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_14
timestamp 1694765150
transform 1 0 19737 0 1 924
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_15
timestamp 1694765150
transform 1 0 20025 0 1 924
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_16
timestamp 1694765150
transform 1 0 18329 0 1 3732
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_17
timestamp 1694765150
transform 1 0 18617 0 1 3732
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_18
timestamp 1694765150
transform 1 0 19737 0 1 3732
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_19
timestamp 1694765150
transform 1 0 20025 0 1 3732
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_20
timestamp 1694765150
transform 1 0 18329 0 1 2796
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_21
timestamp 1694765150
transform 1 0 18617 0 1 2796
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_22
timestamp 1694765150
transform 1 0 19737 0 1 2796
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_23
timestamp 1694765150
transform 1 0 20025 0 1 2796
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_24
timestamp 1694765150
transform -1 0 23481 0 1 1860
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_25
timestamp 1694765150
transform -1 0 23769 0 1 1860
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_26
timestamp 1694765150
transform -1 0 24889 0 1 1860
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_27
timestamp 1694765150
transform -1 0 25177 0 1 1860
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_28
timestamp 1694765150
transform -1 0 23769 0 1 924
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_29
timestamp 1694765150
transform -1 0 23481 0 1 924
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_30
timestamp 1694765150
transform -1 0 24889 0 1 924
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_31
timestamp 1694765150
transform -1 0 25177 0 1 924
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_32
timestamp 1694765150
transform -1 0 23769 0 1 -12
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_33
timestamp 1694765150
transform -1 0 23481 0 1 -12
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_34
timestamp 1694765150
transform -1 0 24889 0 1 -12
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_35
timestamp 1694765150
transform -1 0 25177 0 1 -12
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_36
timestamp 1694765150
transform -1 0 23481 0 1 -948
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_37
timestamp 1694765150
transform -1 0 23769 0 1 -948
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_38
timestamp 1694765150
transform -1 0 24889 0 1 -948
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_39
timestamp 1694765150
transform -1 0 25177 0 1 -948
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_40
timestamp 1694765150
transform -1 0 23481 0 1 3732
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_41
timestamp 1694765150
transform -1 0 23769 0 1 3732
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_42
timestamp 1694765150
transform -1 0 25177 0 1 3732
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_43
timestamp 1694765150
transform -1 0 24889 0 1 3732
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_44
timestamp 1694765150
transform -1 0 23481 0 1 2796
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_45
timestamp 1694765150
transform -1 0 23769 0 1 2796
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_46
timestamp 1694765150
transform -1 0 25177 0 1 2796
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_47
timestamp 1694765150
transform -1 0 24889 0 1 2796
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_48
timestamp 1694765150
transform 1 0 27450 0 1 1860
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_49
timestamp 1694765150
transform 1 0 27450 0 1 924
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_50
timestamp 1694765150
transform 1 0 27450 0 1 -12
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_51
timestamp 1694765150
transform 1 0 27450 0 1 -948
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_52
timestamp 1694765150
transform 1 0 29146 0 1 1860
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_53
timestamp 1694765150
transform 1 0 28858 0 1 1860
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_54
timestamp 1694765150
transform 1 0 27738 0 1 1860
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_55
timestamp 1694765150
transform 1 0 28858 0 1 924
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_56
timestamp 1694765150
transform 1 0 29146 0 1 924
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_57
timestamp 1694765150
transform 1 0 27738 0 1 924
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_58
timestamp 1694765150
transform 1 0 28858 0 1 -12
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_59
timestamp 1694765150
transform 1 0 29146 0 1 -12
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_60
timestamp 1694765150
transform 1 0 27738 0 1 -12
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_61
timestamp 1694765150
transform 1 0 29146 0 1 -948
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_62
timestamp 1694765150
transform 1 0 28858 0 1 -948
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_63
timestamp 1694765150
transform 1 0 27738 0 1 -948
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_64
timestamp 1694765150
transform 1 0 27450 0 1 3732
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_65
timestamp 1694765150
transform 1 0 27450 0 1 2796
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_66
timestamp 1694765150
transform 1 0 29146 0 1 3732
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_67
timestamp 1694765150
transform 1 0 28858 0 1 3732
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_68
timestamp 1694765150
transform 1 0 27738 0 1 3732
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_69
timestamp 1694765150
transform 1 0 29146 0 1 2796
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_70
timestamp 1694765150
transform 1 0 28858 0 1 2796
box -140 -368 140 368
use nmos_3p3_M86RTJ  nmos_3p3_M86RTJ_71
timestamp 1694765150
transform 1 0 27738 0 1 2796
box -140 -368 140 368
use nmos_3p3_NE3WC4  nmos_3p3_NE3WC4_0
timestamp 1694939532
transform 1 0 12372 0 1 -6948
box -212 -268 212 268
use nmos_3p3_NE3WC4  nmos_3p3_NE3WC4_1
timestamp 1694939532
transform 1 0 16276 0 1 -6948
box -212 -268 212 268
use nmos_3p3_NE3WC4  nmos_3p3_NE3WC4_2
timestamp 1694939532
transform 1 0 12804 0 1 -6948
box -212 -268 212 268
use nmos_3p3_QNHHD6  nmos_3p3_QNHHD6_0
timestamp 1693895158
transform 1 0 6082 0 1 -7465
box -168 -168 168 168
use nmos_3p3_S75EG7  nmos_3p3_S75EG7_0
timestamp 1693897923
transform 1 0 7734 0 1 -6828
box -1180 -168 1180 168
use nmos_3p3_U56RT2  nmos_3p3_U56RT2_0
timestamp 1693899225
transform 1 0 9878 0 1 -7465
box -540 -168 540 168
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_0
timestamp 1693069569
transform 1 0 8602 0 1 1364
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_1
timestamp 1693069569
transform 1 0 8314 0 1 1364
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_2
timestamp 1693069569
transform 1 0 10522 0 1 1364
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_3
timestamp 1693069569
transform 1 0 10234 0 1 1364
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_4
timestamp 1693069569
transform 1 0 10522 0 1 -1222
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_5
timestamp 1693069569
transform 1 0 10234 0 1 -1222
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_6
timestamp 1693069569
transform 1 0 8602 0 1 -1222
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_7
timestamp 1693069569
transform 1 0 8314 0 1 -1222
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_8
timestamp 1693069569
transform 1 0 8314 0 1 -360
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_9
timestamp 1693069569
transform 1 0 8602 0 1 -360
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_10
timestamp 1693069569
transform 1 0 10234 0 1 -360
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_11
timestamp 1693069569
transform 1 0 10522 0 1 -360
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_12
timestamp 1693069569
transform 1 0 8314 0 1 502
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_13
timestamp 1693069569
transform 1 0 8602 0 1 502
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_14
timestamp 1693069569
transform 1 0 10234 0 1 502
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_15
timestamp 1693069569
transform 1 0 10522 0 1 502
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_16
timestamp 1693069569
transform 1 0 6367 0 1 -341
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_17
timestamp 1693069569
transform 1 0 6079 0 1 -341
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_18
timestamp 1693069569
transform 1 0 7775 0 1 -341
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_19
timestamp 1693069569
transform 1 0 7487 0 1 -341
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_20
timestamp 1693069569
transform 1 0 7775 0 1 -1203
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_21
timestamp 1693069569
transform 1 0 7487 0 1 -1203
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_22
timestamp 1693069569
transform 1 0 6367 0 1 -1203
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_23
timestamp 1693069569
transform 1 0 6079 0 1 -1203
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_24
timestamp 1693069569
transform 1 0 6079 0 1 521
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_25
timestamp 1693069569
transform 1 0 6367 0 1 521
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_26
timestamp 1693069569
transform 1 0 7487 0 1 521
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_27
timestamp 1693069569
transform 1 0 7775 0 1 521
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_28
timestamp 1693069569
transform 1 0 6079 0 1 2245
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_29
timestamp 1693069569
transform 1 0 6367 0 1 2245
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_30
timestamp 1693069569
transform 1 0 7487 0 1 2245
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_31
timestamp 1693069569
transform 1 0 7775 0 1 2245
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_32
timestamp 1693069569
transform 1 0 6079 0 1 1383
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_33
timestamp 1693069569
transform 1 0 6367 0 1 1383
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_34
timestamp 1693069569
transform 1 0 7487 0 1 1383
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_35
timestamp 1693069569
transform 1 0 7775 0 1 1383
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_36
timestamp 1693069569
transform 1 0 6079 0 1 3107
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_37
timestamp 1693069569
transform 1 0 6367 0 1 3107
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_38
timestamp 1693069569
transform 1 0 7487 0 1 3107
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_39
timestamp 1693069569
transform 1 0 7775 0 1 3107
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_40
timestamp 1693069569
transform 1 0 6079 0 1 3969
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_41
timestamp 1693069569
transform 1 0 6367 0 1 3969
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_42
timestamp 1693069569
transform 1 0 7487 0 1 3969
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_43
timestamp 1693069569
transform 1 0 7775 0 1 3969
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_44
timestamp 1693069569
transform 1 0 6079 0 1 4831
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_45
timestamp 1693069569
transform 1 0 6367 0 1 4831
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_46
timestamp 1693069569
transform 1 0 7487 0 1 4831
box -140 -356 140 356
use nmos_3p3_UUQWW2  nmos_3p3_UUQWW2_47
timestamp 1693069569
transform 1 0 7775 0 1 4831
box -140 -356 140 356
use nmos_3p3_V56RT2  nmos_3p3_V56RT2_0
timestamp 1693898117
transform 1 0 8694 0 1 -7465
box -620 -168 620 168
use pfet_03v3_6DHECV  pfet_03v3_6DHECV_0
timestamp 1695292659
transform 1 0 4019 0 1 -5123
box -202 -530 202 530
use PGA_DECODER_magic  PGA_DECODER_magic_0
timestamp 1692798605
transform -1 0 59238 0 1 -9759
box -647 -950 2713 6754
use pga_res_magice_parallel  pga_res_magice_parallel_0
timestamp 1694752906
transform 1 0 6673 0 1 -16352
box 0 -2440 11127 2440
use pga_res_magice_parallel  pga_res_magice_parallel_1
timestamp 1694752906
transform 1 0 23673 0 1 -16352
box 0 -2440 11127 2440
use pmos_3p3_5C3RD7  pmos_3p3_5C3RD7_0
timestamp 1693568584
transform 1 0 2915 0 1 -5123
box -554 -530 554 530
use pmos_3p3_5L6RD7  pmos_3p3_5L6RD7_1
timestamp 1693886538
transform 1 0 3239 0 1 -6383
box -230 -530 230 530
use pmos_3p3_5L6RD7  pmos_3p3_5L6RD7_2
timestamp 1693886538
transform 1 0 3583 0 1 -6383
box -230 -530 230 530
use pmos_3p3_5LZQD7  pmos_3p3_5LZQD7_0
timestamp 1693568584
transform 1 0 1943 0 1 -5123
box -662 -530 662 530
use pmos_3p3_5LZQD7  pmos_3p3_5LZQD7_1
timestamp 1693568584
transform 1 0 1951 0 1 -6383
box -662 -530 662 530
use pmos_3p3_5UYQD7  pmos_3p3_5UYQD7_0
timestamp 1693568584
transform 1 0 3563 0 1 -5123
box -338 -530 338 530
use pmos_3p3_HDY8L7  pmos_3p3_HDY8L7_0
timestamp 1692617267
transform 1 0 556 0 1 -55
box -230 -1586 230 1586
use pmos_3p3_HDY8L7  pmos_3p3_HDY8L7_1
timestamp 1692617267
transform 1 0 2500 0 1 -55
box -230 -1586 230 1586
use pmos_3p3_HMY8L7  pmos_3p3_HMY8L7_0
timestamp 1692617267
transform 1 0 1528 0 1 -55
box -986 -1586 986 1586
use pmos_3p3_K823KY  pmos_3p3_K823KY_0
timestamp 1693883759
transform 1 0 3835 0 1 -7293
box -274 -180 274 180
use pmos_3p3_M2NNAR  pmos_3p3_M2NNAR_0
timestamp 1694922630
transform 1 0 21212 0 1 -5782
box -282 -1534 282 1534
use pmos_3p3_M2NNAR  pmos_3p3_M2NNAR_1
timestamp 1694922630
transform 1 0 20892 0 1 -5782
box -282 -1534 282 1534
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_0
timestamp 1694686376
transform -1 0 62362 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_1
timestamp 1694686376
transform -1 0 64282 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_2
timestamp 1694686376
transform -1 0 63962 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_3
timestamp 1694686376
transform -1 0 63642 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_4
timestamp 1694686376
transform -1 0 63322 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_5
timestamp 1694686376
transform -1 0 63002 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_6
timestamp 1694686376
transform -1 0 62682 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_7
timestamp 1694686376
transform -1 0 63962 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_8
timestamp 1694686376
transform -1 0 64282 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_9
timestamp 1694686376
transform -1 0 62362 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_10
timestamp 1694686376
transform -1 0 62682 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_11
timestamp 1694686376
transform -1 0 63002 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_12
timestamp 1694686376
transform -1 0 63322 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_13
timestamp 1694686376
transform -1 0 63642 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_14
timestamp 1694686376
transform -1 0 63962 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_15
timestamp 1694686376
transform -1 0 64282 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_16
timestamp 1694686376
transform -1 0 63002 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_17
timestamp 1694686376
transform -1 0 63322 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_18
timestamp 1694686376
transform -1 0 63642 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_19
timestamp 1694686376
transform -1 0 62362 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_20
timestamp 1694686376
transform -1 0 62682 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_21
timestamp 1694686376
transform -1 0 63962 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_22
timestamp 1694686376
transform -1 0 64282 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_23
timestamp 1694686376
transform -1 0 62362 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_24
timestamp 1694686376
transform -1 0 62682 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_25
timestamp 1694686376
transform -1 0 63002 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_26
timestamp 1694686376
transform -1 0 63322 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_27
timestamp 1694686376
transform -1 0 63642 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_28
timestamp 1694686376
transform 1 0 56802 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_29
timestamp 1694686376
transform 1 0 57442 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_30
timestamp 1694686376
transform 1 0 57122 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_31
timestamp 1694686376
transform 1 0 58082 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_32
timestamp 1694686376
transform 1 0 57762 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_33
timestamp 1694686376
transform 1 0 58722 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_34
timestamp 1694686376
transform 1 0 58402 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_35
timestamp 1694686376
transform 1 0 56802 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_36
timestamp 1694686376
transform 1 0 57442 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_37
timestamp 1694686376
transform 1 0 57122 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_38
timestamp 1694686376
transform 1 0 58082 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_39
timestamp 1694686376
transform 1 0 57762 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_40
timestamp 1694686376
transform 1 0 58722 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_41
timestamp 1694686376
transform 1 0 58402 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_42
timestamp 1694686376
transform 1 0 56802 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_43
timestamp 1694686376
transform 1 0 57442 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_44
timestamp 1694686376
transform 1 0 57122 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_45
timestamp 1694686376
transform 1 0 58082 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_46
timestamp 1694686376
transform 1 0 57762 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_47
timestamp 1694686376
transform 1 0 58722 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_48
timestamp 1694686376
transform 1 0 58402 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_49
timestamp 1694686376
transform 1 0 57442 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_50
timestamp 1694686376
transform 1 0 57762 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_51
timestamp 1694686376
transform 1 0 58082 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_52
timestamp 1694686376
transform 1 0 58402 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_53
timestamp 1694686376
transform 1 0 58722 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_54
timestamp 1694686376
transform 1 0 56802 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_55
timestamp 1694686376
transform 1 0 57122 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_56
timestamp 1694686376
transform -1 0 54586 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_57
timestamp 1694686376
transform -1 0 54586 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_58
timestamp 1694686376
transform -1 0 54586 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_59
timestamp 1694686376
transform -1 0 53946 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_60
timestamp 1694686376
transform -1 0 54266 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_61
timestamp 1694686376
transform -1 0 53306 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_62
timestamp 1694686376
transform -1 0 53626 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_63
timestamp 1694686376
transform -1 0 52986 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_64
timestamp 1694686376
transform -1 0 53946 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_65
timestamp 1694686376
transform -1 0 54266 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_66
timestamp 1694686376
transform -1 0 53306 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_67
timestamp 1694686376
transform -1 0 53626 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_68
timestamp 1694686376
transform -1 0 52986 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_69
timestamp 1694686376
transform -1 0 53946 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_70
timestamp 1694686376
transform -1 0 54266 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_71
timestamp 1694686376
transform -1 0 53306 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_72
timestamp 1694686376
transform -1 0 53626 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_73
timestamp 1694686376
transform -1 0 52986 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_74
timestamp 1694686376
transform -1 0 54586 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_75
timestamp 1694686376
transform -1 0 53946 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_76
timestamp 1694686376
transform -1 0 53626 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_77
timestamp 1694686376
transform -1 0 53306 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_78
timestamp 1694686376
transform -1 0 52986 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_79
timestamp 1694686376
transform -1 0 54266 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_80
timestamp 1694686376
transform -1 0 52666 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_81
timestamp 1694686376
transform -1 0 52666 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_82
timestamp 1694686376
transform -1 0 52666 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_83
timestamp 1694686376
transform -1 0 52666 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_84
timestamp 1694686376
transform 1 0 49026 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_85
timestamp 1694686376
transform 1 0 48706 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_86
timestamp 1694686376
transform 1 0 48386 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_87
timestamp 1694686376
transform 1 0 48066 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_88
timestamp 1694686376
transform 1 0 47746 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_89
timestamp 1694686376
transform 1 0 47106 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_90
timestamp 1694686376
transform 1 0 47426 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_91
timestamp 1694686376
transform 1 0 49026 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_92
timestamp 1694686376
transform 1 0 48706 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_93
timestamp 1694686376
transform 1 0 48386 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_94
timestamp 1694686376
transform 1 0 47746 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_95
timestamp 1694686376
transform 1 0 48066 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_96
timestamp 1694686376
transform 1 0 47426 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_97
timestamp 1694686376
transform 1 0 47106 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_98
timestamp 1694686376
transform 1 0 49026 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_99
timestamp 1694686376
transform 1 0 48706 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_100
timestamp 1694686376
transform 1 0 48386 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_101
timestamp 1694686376
transform 1 0 48066 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_102
timestamp 1694686376
transform 1 0 47746 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_103
timestamp 1694686376
transform 1 0 47426 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_104
timestamp 1694686376
transform 1 0 47106 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_105
timestamp 1694686376
transform 1 0 47746 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_106
timestamp 1694686376
transform 1 0 48066 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_107
timestamp 1694686376
transform 1 0 48386 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_108
timestamp 1694686376
transform 1 0 48706 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_109
timestamp 1694686376
transform 1 0 49026 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_110
timestamp 1694686376
transform 1 0 47106 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_111
timestamp 1694686376
transform 1 0 47426 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_112
timestamp 1694686376
transform -1 0 42970 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_113
timestamp 1694686376
transform -1 0 43290 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_114
timestamp 1694686376
transform -1 0 43610 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_115
timestamp 1694686376
transform -1 0 43930 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_116
timestamp 1694686376
transform -1 0 44250 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_117
timestamp 1694686376
transform -1 0 44890 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_118
timestamp 1694686376
transform -1 0 44570 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_119
timestamp 1694686376
transform -1 0 42970 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_120
timestamp 1694686376
transform -1 0 43290 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_121
timestamp 1694686376
transform -1 0 43610 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_122
timestamp 1694686376
transform -1 0 44250 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_123
timestamp 1694686376
transform -1 0 43930 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_124
timestamp 1694686376
transform -1 0 44570 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_125
timestamp 1694686376
transform -1 0 44890 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_126
timestamp 1694686376
transform -1 0 42970 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_127
timestamp 1694686376
transform -1 0 43290 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_128
timestamp 1694686376
transform -1 0 43610 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_129
timestamp 1694686376
transform -1 0 43930 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_130
timestamp 1694686376
transform -1 0 44250 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_131
timestamp 1694686376
transform -1 0 44570 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_132
timestamp 1694686376
transform -1 0 44890 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_133
timestamp 1694686376
transform -1 0 44250 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_134
timestamp 1694686376
transform -1 0 43930 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_135
timestamp 1694686376
transform -1 0 43610 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_136
timestamp 1694686376
transform -1 0 43290 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_137
timestamp 1694686376
transform -1 0 42970 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_138
timestamp 1694686376
transform -1 0 44890 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_139
timestamp 1694686376
transform -1 0 44570 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_140
timestamp 1694686376
transform 1 0 39330 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_141
timestamp 1694686376
transform 1 0 39010 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_142
timestamp 1694686376
transform 1 0 38690 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_143
timestamp 1694686376
transform 1 0 38370 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_144
timestamp 1694686376
transform 1 0 38050 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_145
timestamp 1694686376
transform 1 0 37410 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_146
timestamp 1694686376
transform 1 0 37730 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_147
timestamp 1694686376
transform 1 0 39330 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_148
timestamp 1694686376
transform 1 0 39010 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_149
timestamp 1694686376
transform 1 0 38690 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_150
timestamp 1694686376
transform 1 0 38050 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_151
timestamp 1694686376
transform 1 0 38370 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_152
timestamp 1694686376
transform 1 0 37730 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_153
timestamp 1694686376
transform 1 0 37410 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_154
timestamp 1694686376
transform 1 0 39330 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_155
timestamp 1694686376
transform 1 0 39010 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_156
timestamp 1694686376
transform 1 0 38690 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_157
timestamp 1694686376
transform 1 0 38370 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_158
timestamp 1694686376
transform 1 0 38050 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_159
timestamp 1694686376
transform 1 0 37730 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_160
timestamp 1694686376
transform 1 0 37410 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_161
timestamp 1694686376
transform 1 0 38050 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_162
timestamp 1694686376
transform 1 0 38370 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_163
timestamp 1694686376
transform 1 0 38690 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_164
timestamp 1694686376
transform 1 0 39010 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_165
timestamp 1694686376
transform 1 0 39330 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_166
timestamp 1694686376
transform 1 0 37410 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_167
timestamp 1694686376
transform 1 0 37730 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_168
timestamp 1694686376
transform -1 0 34554 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_169
timestamp 1694686376
transform -1 0 34234 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_170
timestamp 1694686376
transform -1 0 33914 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_171
timestamp 1694686376
transform -1 0 33594 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_172
timestamp 1694686376
transform -1 0 33274 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_173
timestamp 1694686376
transform -1 0 35194 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_174
timestamp 1694686376
transform -1 0 34874 0 1 2232
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_175
timestamp 1694686376
transform -1 0 33274 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_176
timestamp 1694686376
transform -1 0 33594 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_177
timestamp 1694686376
transform -1 0 33914 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_178
timestamp 1694686376
transform -1 0 34234 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_179
timestamp 1694686376
transform -1 0 34554 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_180
timestamp 1694686376
transform -1 0 35194 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_181
timestamp 1694686376
transform -1 0 34874 0 1 1172
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_182
timestamp 1694686376
transform -1 0 33274 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_183
timestamp 1694686376
transform -1 0 33594 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_184
timestamp 1694686376
transform -1 0 33914 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_185
timestamp 1694686376
transform -1 0 34554 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_186
timestamp 1694686376
transform -1 0 34234 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_187
timestamp 1694686376
transform -1 0 34874 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_188
timestamp 1694686376
transform -1 0 35194 0 1 112
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_189
timestamp 1694686376
transform -1 0 33274 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_190
timestamp 1694686376
transform -1 0 33594 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_191
timestamp 1694686376
transform -1 0 33914 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_192
timestamp 1694686376
transform -1 0 34234 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_193
timestamp 1694686376
transform -1 0 34554 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_194
timestamp 1694686376
transform -1 0 34874 0 1 -948
box -282 -430 282 430
use pmos_3p3_M22VAR  pmos_3p3_M22VAR_195
timestamp 1694686376
transform -1 0 35194 0 1 -948
box -282 -430 282 430
use pmos_3p3_M82RNG  pmos_3p3_M82RNG_0
timestamp 1693885183
transform 1 0 907 0 1 -7293
box -202 -180 202 180
use pmos_3p3_M82RNG  pmos_3p3_M82RNG_1
timestamp 1693885183
transform 1 0 4067 0 1 -7293
box -202 -180 202 180
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_0
timestamp 1694686376
transform -1 0 64522 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_1
timestamp 1694686376
transform -1 0 64810 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_2
timestamp 1694686376
transform -1 0 61834 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_3
timestamp 1694686376
transform -1 0 62122 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_4
timestamp 1694686376
transform -1 0 64810 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_5
timestamp 1694686376
transform -1 0 64522 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_6
timestamp 1694686376
transform -1 0 61834 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_7
timestamp 1694686376
transform -1 0 62122 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_8
timestamp 1694686376
transform -1 0 64522 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_9
timestamp 1694686376
transform -1 0 64810 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_10
timestamp 1694686376
transform -1 0 62122 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_11
timestamp 1694686376
transform -1 0 61834 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_12
timestamp 1694686376
transform -1 0 64522 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_13
timestamp 1694686376
transform -1 0 64810 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_14
timestamp 1694686376
transform -1 0 61834 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_15
timestamp 1694686376
transform -1 0 62122 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_16
timestamp 1694686376
transform 1 0 56274 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_17
timestamp 1694686376
transform 1 0 56274 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_18
timestamp 1694686376
transform 1 0 56274 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_19
timestamp 1694686376
transform 1 0 56562 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_20
timestamp 1694686376
transform 1 0 58962 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_21
timestamp 1694686376
transform 1 0 59250 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_22
timestamp 1694686376
transform 1 0 56562 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_23
timestamp 1694686376
transform 1 0 58962 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_24
timestamp 1694686376
transform 1 0 59250 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_25
timestamp 1694686376
transform 1 0 56562 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_26
timestamp 1694686376
transform 1 0 59250 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_27
timestamp 1694686376
transform 1 0 58962 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_28
timestamp 1694686376
transform 1 0 56274 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_29
timestamp 1694686376
transform 1 0 58962 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_30
timestamp 1694686376
transform 1 0 59250 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_31
timestamp 1694686376
transform 1 0 56562 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_32
timestamp 1694686376
transform -1 0 55114 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_33
timestamp 1694686376
transform -1 0 54826 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_34
timestamp 1694686376
transform -1 0 55114 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_35
timestamp 1694686376
transform -1 0 54826 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_36
timestamp 1694686376
transform -1 0 55114 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_37
timestamp 1694686376
transform -1 0 54826 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_38
timestamp 1694686376
transform -1 0 55114 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_39
timestamp 1694686376
transform -1 0 54826 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_40
timestamp 1694686376
transform -1 0 52426 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_41
timestamp 1694686376
transform -1 0 52138 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_42
timestamp 1694686376
transform -1 0 52138 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_43
timestamp 1694686376
transform -1 0 52426 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_44
timestamp 1694686376
transform -1 0 52426 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_45
timestamp 1694686376
transform -1 0 52138 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_46
timestamp 1694686376
transform -1 0 52426 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_47
timestamp 1694686376
transform -1 0 52138 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_48
timestamp 1694686376
transform 1 0 46866 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_49
timestamp 1694686376
transform 1 0 46578 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_50
timestamp 1694686376
transform 1 0 46866 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_51
timestamp 1694686376
transform 1 0 46578 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_52
timestamp 1694686376
transform 1 0 46578 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_53
timestamp 1694686376
transform 1 0 46866 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_54
timestamp 1694686376
transform 1 0 49554 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_55
timestamp 1694686376
transform 1 0 49266 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_56
timestamp 1694686376
transform 1 0 49266 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_57
timestamp 1694686376
transform 1 0 49554 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_58
timestamp 1694686376
transform 1 0 49266 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_59
timestamp 1694686376
transform 1 0 49554 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_60
timestamp 1694686376
transform 1 0 46578 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_61
timestamp 1694686376
transform 1 0 46866 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_62
timestamp 1694686376
transform 1 0 49266 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_63
timestamp 1694686376
transform 1 0 49554 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_64
timestamp 1694686376
transform -1 0 45418 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_65
timestamp 1694686376
transform -1 0 45418 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_66
timestamp 1694686376
transform -1 0 45418 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_67
timestamp 1694686376
transform -1 0 42730 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_68
timestamp 1694686376
transform -1 0 42730 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_69
timestamp 1694686376
transform -1 0 42730 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_70
timestamp 1694686376
transform -1 0 45130 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_71
timestamp 1694686376
transform -1 0 45130 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_72
timestamp 1694686376
transform -1 0 45130 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_73
timestamp 1694686376
transform -1 0 42442 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_74
timestamp 1694686376
transform -1 0 42442 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_75
timestamp 1694686376
transform -1 0 42442 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_76
timestamp 1694686376
transform -1 0 45418 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_77
timestamp 1694686376
transform -1 0 42730 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_78
timestamp 1694686376
transform -1 0 45130 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_79
timestamp 1694686376
transform -1 0 42442 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_80
timestamp 1694686376
transform 1 0 37170 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_81
timestamp 1694686376
transform 1 0 36882 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_82
timestamp 1694686376
transform 1 0 37170 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_83
timestamp 1694686376
transform 1 0 36882 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_84
timestamp 1694686376
transform 1 0 36882 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_85
timestamp 1694686376
transform 1 0 37170 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_86
timestamp 1694686376
transform 1 0 39570 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_87
timestamp 1694686376
transform 1 0 39570 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_88
timestamp 1694686376
transform 1 0 39570 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_89
timestamp 1694686376
transform 1 0 36882 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_90
timestamp 1694686376
transform 1 0 37170 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_91
timestamp 1694686376
transform 1 0 39570 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_92
timestamp 1694686376
transform -1 0 32746 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_93
timestamp 1694686376
transform -1 0 32746 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_94
timestamp 1694686376
transform -1 0 32746 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_95
timestamp 1694686376
transform -1 0 32746 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_96
timestamp 1694686376
transform -1 0 33034 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_97
timestamp 1694686376
transform -1 0 35722 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_98
timestamp 1694686376
transform -1 0 35434 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_99
timestamp 1694686376
transform -1 0 33034 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_100
timestamp 1694686376
transform -1 0 33034 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_101
timestamp 1694686376
transform -1 0 33034 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_102
timestamp 1694686376
transform -1 0 35434 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_103
timestamp 1694686376
transform -1 0 35722 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_104
timestamp 1694686376
transform -1 0 35434 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_105
timestamp 1694686376
transform -1 0 35722 0 1 112
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_106
timestamp 1694686376
transform -1 0 35722 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_107
timestamp 1694686376
transform -1 0 35434 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_108
timestamp 1694686376
transform 1 0 39858 0 1 2232
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_109
timestamp 1694686376
transform 1 0 39858 0 1 1172
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_110
timestamp 1694686376
transform 1 0 39858 0 1 -948
box -202 -430 202 430
use pmos_3p3_MA2VAR  pmos_3p3_MA2VAR_111
timestamp 1694686376
transform 1 0 39858 0 1 112
box -202 -430 202 430
use pmos_3p3_MAEVAR  pmos_3p3_MAEVAR_0
timestamp 1694925056
transform 1 0 21580 0 1 -5046
box -202 -798 202 798
use pmos_3p3_MANNAR  pmos_3p3_MANNAR_0
timestamp 1694925645
transform 1 0 21868 0 1 -5782
box -202 -1534 202 1534
use pmos_3p3_MANNAR  pmos_3p3_MANNAR_1
timestamp 1694925645
transform 1 0 18412 0 1 -5782
box -202 -1534 202 1534
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_0
timestamp 1692806196
transform -1 0 14778 0 1 871
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_1
timestamp 1692806196
transform -1 0 15898 0 1 -165
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_2
timestamp 1692806196
transform -1 0 14778 0 1 -1201
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_3
timestamp 1692806196
transform -1 0 16186 0 1 -1201
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_4
timestamp 1692806196
transform -1 0 16186 0 1 -165
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_5
timestamp 1692806196
transform -1 0 14778 0 1 -165
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_6
timestamp 1692806196
transform -1 0 16186 0 1 1907
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_7
timestamp 1692806196
transform -1 0 14778 0 1 1907
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_8
timestamp 1692806196
transform -1 0 14490 0 1 871
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_9
timestamp 1692806196
transform -1 0 14490 0 1 1907
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_10
timestamp 1692806196
transform -1 0 14490 0 1 -165
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_11
timestamp 1692806196
transform -1 0 14490 0 1 -1201
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_12
timestamp 1692806196
transform -1 0 15898 0 1 1907
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_13
timestamp 1692806196
transform -1 0 15898 0 1 871
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_14
timestamp 1692806196
transform -1 0 16186 0 1 871
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_15
timestamp 1692806196
transform -1 0 15898 0 1 -1201
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_16
timestamp 1692806196
transform -1 0 11696 0 1 871
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_17
timestamp 1692806196
transform -1 0 13904 0 1 871
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_18
timestamp 1692806196
transform -1 0 13616 0 1 871
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_19
timestamp 1692806196
transform -1 0 11984 0 1 871
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_20
timestamp 1692806196
transform -1 0 13904 0 1 -1201
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_21
timestamp 1692806196
transform -1 0 13616 0 1 -1201
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_22
timestamp 1692806196
transform -1 0 11696 0 1 -1201
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_23
timestamp 1692806196
transform -1 0 11984 0 1 -1201
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_24
timestamp 1692806196
transform -1 0 13616 0 1 -165
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_25
timestamp 1692806196
transform -1 0 13904 0 1 -165
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_26
timestamp 1692806196
transform -1 0 11984 0 1 -165
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_27
timestamp 1692806196
transform -1 0 11696 0 1 -165
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_28
timestamp 1692806196
transform -1 0 13616 0 1 1907
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_29
timestamp 1692806196
transform -1 0 13904 0 1 1907
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_30
timestamp 1692806196
transform -1 0 11984 0 1 1907
box -202 -443 202 443
use pmos_3p3_ME7U2H  pmos_3p3_ME7U2H_31
timestamp 1692806196
transform -1 0 11696 0 1 1907
box -202 -443 202 443
use pmos_3p3_MEKUKR  pmos_3p3_MEKUKR_0
timestamp 1694924682
transform 1 0 21580 0 1 -6200
box -202 -380 202 380
use pmos_3p3_MEKUKR  pmos_3p3_MEKUKR_1
timestamp 1694924682
transform 1 0 21580 0 1 -6936
box -202 -380 202 380
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_0
timestamp 1692678901
transform 1 0 4622 0 1 1104
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_1
timestamp 1692678901
transform 1 0 3502 0 1 1104
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_2
timestamp 1692678901
transform 1 0 4910 0 1 -26
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_3
timestamp 1692678901
transform 1 0 3214 0 1 -1156
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_4
timestamp 1692678901
transform 1 0 3502 0 1 -26
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_5
timestamp 1692678901
transform 1 0 4622 0 1 -26
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_6
timestamp 1692678901
transform 1 0 4622 0 1 4494
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_7
timestamp 1692678901
transform 1 0 3502 0 1 4494
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_8
timestamp 1692678901
transform 1 0 4622 0 1 2234
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_9
timestamp 1692678901
transform 1 0 3502 0 1 2234
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_10
timestamp 1692678901
transform 1 0 3502 0 1 3364
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_11
timestamp 1692678901
transform 1 0 4622 0 1 3364
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_12
timestamp 1692678901
transform 1 0 4622 0 1 -1156
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_13
timestamp 1692678901
transform 1 0 4910 0 1 -1156
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_14
timestamp 1692678901
transform 1 0 4910 0 1 3364
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_15
timestamp 1692678901
transform 1 0 4910 0 1 1104
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_16
timestamp 1692678901
transform 1 0 4910 0 1 2234
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_17
timestamp 1692678901
transform 1 0 4910 0 1 4494
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_18
timestamp 1692678901
transform 1 0 3502 0 1 -1156
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_19
timestamp 1692678901
transform 1 0 3214 0 1 1104
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_20
timestamp 1692678901
transform 1 0 3214 0 1 -26
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_21
timestamp 1692678901
transform 1 0 3214 0 1 2234
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_22
timestamp 1692678901
transform 1 0 3214 0 1 3364
box -202 -505 202 505
use pmos_3p3_MES6FR  pmos_3p3_MES6FR_23
timestamp 1692678901
transform 1 0 3214 0 1 4494
box -202 -505 202 505
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_0
timestamp 1692877802
transform -1 0 15018 0 1 871
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_1
timestamp 1692877802
transform -1 0 15658 0 1 -165
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_2
timestamp 1692877802
transform -1 0 15338 0 1 -165
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_3
timestamp 1692877802
transform -1 0 15018 0 1 -1201
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_4
timestamp 1692877802
transform -1 0 15338 0 1 -1201
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_5
timestamp 1692877802
transform -1 0 15658 0 1 -1201
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_6
timestamp 1692877802
transform -1 0 15338 0 1 871
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_7
timestamp 1692877802
transform -1 0 15658 0 1 871
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_8
timestamp 1692877802
transform -1 0 15018 0 1 -165
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_9
timestamp 1692877802
transform -1 0 15338 0 1 1907
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_10
timestamp 1692877802
transform -1 0 15658 0 1 1907
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_11
timestamp 1692877802
transform -1 0 15018 0 1 1907
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_12
timestamp 1692877802
transform -1 0 12352 0 1 871
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_13
timestamp 1692877802
transform -1 0 13248 0 1 871
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_14
timestamp 1692877802
transform -1 0 12800 0 1 871
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_15
timestamp 1692877802
transform -1 0 13248 0 1 -1201
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_16
timestamp 1692877802
transform -1 0 12352 0 1 -1201
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_17
timestamp 1692877802
transform -1 0 12800 0 1 -1201
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_18
timestamp 1692877802
transform -1 0 13248 0 1 -165
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_19
timestamp 1692877802
transform -1 0 12800 0 1 -165
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_20
timestamp 1692877802
transform -1 0 12352 0 1 -165
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_21
timestamp 1692877802
transform -1 0 13248 0 1 1907
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_22
timestamp 1692877802
transform -1 0 12800 0 1 1907
box -282 -443 282 443
use pmos_3p3_MN7U2H  pmos_3p3_MN7U2H_23
timestamp 1692877802
transform -1 0 12352 0 1 1907
box -282 -443 282 443
use pmos_3p3_MNS6FR  pmos_3p3_MNS6FR_0
timestamp 1692678901
transform 1 0 4382 0 1 1104
box -282 -505 282 505
use pmos_3p3_MNS6FR  pmos_3p3_MNS6FR_1
timestamp 1692678901
transform 1 0 3742 0 1 1104
box -282 -505 282 505
use pmos_3p3_MNS6FR  pmos_3p3_MNS6FR_2
timestamp 1692678901
transform 1 0 4062 0 1 1104
box -282 -505 282 505
use pmos_3p3_MNS6FR  pmos_3p3_MNS6FR_3
timestamp 1692678901
transform 1 0 4382 0 1 -1156
box -282 -505 282 505
use pmos_3p3_MNS6FR  pmos_3p3_MNS6FR_4
timestamp 1692678901
transform 1 0 4062 0 1 -1156
box -282 -505 282 505
use pmos_3p3_MNS6FR  pmos_3p3_MNS6FR_5
timestamp 1692678901
transform 1 0 3742 0 1 -1156
box -282 -505 282 505
use pmos_3p3_MNS6FR  pmos_3p3_MNS6FR_6
timestamp 1692678901
transform 1 0 4062 0 1 -26
box -282 -505 282 505
use pmos_3p3_MNS6FR  pmos_3p3_MNS6FR_7
timestamp 1692678901
transform 1 0 4382 0 1 -26
box -282 -505 282 505
use pmos_3p3_MNS6FR  pmos_3p3_MNS6FR_8
timestamp 1692678901
transform 1 0 3742 0 1 -26
box -282 -505 282 505
use pmos_3p3_MNS6FR  pmos_3p3_MNS6FR_9
timestamp 1692678901
transform 1 0 3742 0 1 4494
box -282 -505 282 505
use pmos_3p3_MNS6FR  pmos_3p3_MNS6FR_10
timestamp 1692678901
transform 1 0 4382 0 1 4494
box -282 -505 282 505
use pmos_3p3_MNS6FR  pmos_3p3_MNS6FR_11
timestamp 1692678901
transform 1 0 4062 0 1 4494
box -282 -505 282 505
use pmos_3p3_MNS6FR  pmos_3p3_MNS6FR_12
timestamp 1692678901
transform 1 0 3742 0 1 2234
box -282 -505 282 505
use pmos_3p3_MNS6FR  pmos_3p3_MNS6FR_13
timestamp 1692678901
transform 1 0 4382 0 1 2234
box -282 -505 282 505
use pmos_3p3_MNS6FR  pmos_3p3_MNS6FR_14
timestamp 1692678901
transform 1 0 4062 0 1 2234
box -282 -505 282 505
use pmos_3p3_MNS6FR  pmos_3p3_MNS6FR_15
timestamp 1692678901
transform 1 0 3742 0 1 3364
box -282 -505 282 505
use pmos_3p3_MNS6FR  pmos_3p3_MNS6FR_16
timestamp 1692678901
transform 1 0 4062 0 1 3364
box -282 -505 282 505
use pmos_3p3_MNS6FR  pmos_3p3_MNS6FR_17
timestamp 1692678901
transform 1 0 4382 0 1 3364
box -282 -505 282 505
use pmos_3p3_MQ2VAR  pmos_3p3_MQ2VAR_0
timestamp 1693568990
transform 1 0 2651 0 1 -6383
box -282 -530 282 530
use pmos_3p3_MQ2VAR  pmos_3p3_MQ2VAR_1
timestamp 1693568990
transform 1 0 2971 0 1 -6383
box -282 -530 282 530
use pmos_3p3_MYZUAR  pmos_3p3_MYZUAR_0
timestamp 1693886538
transform 1 0 3859 0 1 -5123
box -202 -530 202 530
use pmos_3p3_MYZUAR  pmos_3p3_MYZUAR_1
timestamp 1693886538
transform 1 0 1203 0 1 -6383
box -202 -530 202 530
use pmos_3p3_MYZUAR  pmos_3p3_MYZUAR_2
timestamp 1693886538
transform 1 0 1195 0 1 -5123
box -202 -530 202 530
use pmos_3p3_MYZUAR  pmos_3p3_MYZUAR_3
timestamp 1693886538
transform 1 0 3771 0 1 -6383
box -202 -530 202 530
use pmos_3p3_MYZUAR  pmos_3p3_MYZUAR_4
timestamp 1693886538
transform 1 0 907 0 1 -6383
box -202 -530 202 530
use pmos_3p3_MYZUAR  pmos_3p3_MYZUAR_5
timestamp 1693886538
transform 1 0 4067 0 1 -6383
box -202 -530 202 530
use pmos_3p3_MYZUAR  pmos_3p3_MYZUAR_6
timestamp 1693886538
transform 1 0 907 0 1 -5123
box -202 -530 202 530
use pmos_3p3_Q3NTJU  pmos_3p3_Q3NTJU_0
timestamp 1694921777
transform 1 0 19612 0 1 -5782
box -1242 -1534 1242 1534
use pmos_3p3_RKK9DS  pmos_3p3_RKK9DS_0
timestamp 1693883759
transform 1 0 2403 0 1 -7293
box -1402 -180 1402 180
use ppolyf_u_2V2ZHK  ppolyf_u_2V2ZHK_0
timestamp 1695096662
transform 1 0 26494 0 1 -6812
box -424 -786 424 786
use ppolyf_u_2V2ZHK  ppolyf_u_2V2ZHK_1
timestamp 1695096662
transform 1 0 24310 0 1 -6812
box -424 -786 424 786
use ppolyf_u_2V2ZHK  ppolyf_u_2V2ZHK_2
timestamp 1695096662
transform 1 0 25038 0 1 -6812
box -424 -786 424 786
use ppolyf_u_2V2ZHK  ppolyf_u_2V2ZHK_3
timestamp 1695096662
transform 1 0 25766 0 1 -6812
box -424 -786 424 786
use ppolyf_u_2V2ZHK  ppolyf_u_2V2ZHK_4
timestamp 1695096662
transform 1 0 26494 0 1 -4840
box -424 -786 424 786
use ppolyf_u_2V2ZHK  ppolyf_u_2V2ZHK_5
timestamp 1695096662
transform 1 0 25766 0 1 -4840
box -424 -786 424 786
use ppolyf_u_2V2ZHK  ppolyf_u_2V2ZHK_6
timestamp 1695096662
transform 1 0 25038 0 1 -4840
box -424 -786 424 786
use ppolyf_u_2V2ZHK  ppolyf_u_2V2ZHK_7
timestamp 1695096662
transform 1 0 24310 0 1 -4840
box -424 -786 424 786
use ppolyf_u_2VJWHK  ppolyf_u_2VJWHK_0
timestamp 1695096662
transform 1 0 23722 0 1 -6812
box -284 -786 284 786
use ppolyf_u_2VJWHK  ppolyf_u_2VJWHK_1
timestamp 1695096662
transform 1 0 27554 0 1 -6812
box -284 -786 284 786
use ppolyf_u_2VJWHK  ppolyf_u_2VJWHK_2
timestamp 1695096662
transform 1 0 27082 0 1 -4840
box -284 -786 284 786
use ppolyf_u_2VJWHK  ppolyf_u_2VJWHK_3
timestamp 1695096662
transform 1 0 23722 0 1 -4840
box -284 -786 284 786
use ppolyf_u_2VJWHK  ppolyf_u_2VJWHK_4
timestamp 1695096662
transform 1 0 27082 0 1 -6812
box -284 -786 284 786
use ppolyf_u_2VJWHK  ppolyf_u_2VJWHK_5
timestamp 1695096662
transform 1 0 23274 0 1 -6812
box -284 -786 284 786
use ppolyf_u_2VJWHK  ppolyf_u_2VJWHK_6
timestamp 1695096662
transform 1 0 27554 0 1 -4840
box -284 -786 284 786
use ppolyf_u_2VJWHK  ppolyf_u_2VJWHK_7
timestamp 1695096662
transform 1 0 23274 0 1 -4840
box -284 -786 284 786
use ppolyf_u_RKG95T  ppolyf_u_RKG95T_0
timestamp 1695190274
transform 1 0 28900 0 1 -4776
box -284 -906 284 906
use ppolyf_u_RKG95T  ppolyf_u_RKG95T_1
timestamp 1695190274
transform 1 0 30636 0 1 -6788
box -284 -906 284 906
use ppolyf_u_RKG95T  ppolyf_u_RKG95T_2
timestamp 1695190274
transform 1 0 30636 0 1 -4776
box -284 -906 284 906
use ppolyf_u_RKG95T  ppolyf_u_RKG95T_3
timestamp 1695190274
transform 1 0 28900 0 1 -6788
box -284 -906 284 906
use ppolyf_u_RRG95T  ppolyf_u_RRG95T_0
timestamp 1695189568
transform 1 0 29768 0 1 -6788
box -704 -906 704 906
use ppolyf_u_RRG95T  ppolyf_u_RRG95T_1
timestamp 1695189568
transform 1 0 29768 0 1 -4776
box -704 -906 704 906
use TGATE_PGA_MAGIC  TGATE_PGA_MAGIC_0
timestamp 1699615441
transform 1 0 7854 0 1 -12334
box -534 -578 564 618
use TGATE_PGA_MAGIC  TGATE_PGA_MAGIC_1
timestamp 1699615441
transform 1 0 9854 0 1 -12334
box -534 -578 564 618
use TGATE_PGA_MAGIC  TGATE_PGA_MAGIC_2
timestamp 1699615441
transform 1 0 17854 0 1 -12334
box -534 -578 564 618
use TGATE_PGA_MAGIC  TGATE_PGA_MAGIC_3
timestamp 1699615441
transform 1 0 11854 0 1 -12334
box -534 -578 564 618
use TGATE_PGA_MAGIC  TGATE_PGA_MAGIC_4
timestamp 1699615441
transform 1 0 13854 0 1 -12334
box -534 -578 564 618
use TGATE_PGA_MAGIC  TGATE_PGA_MAGIC_5
timestamp 1699615441
transform 1 0 15854 0 1 -12334
box -534 -578 564 618
use TGATE_PGA_MAGIC  TGATE_PGA_MAGIC_6
timestamp 1699615441
transform 1 0 32854 0 1 -12334
box -534 -578 564 618
use TGATE_PGA_MAGIC  TGATE_PGA_MAGIC_7
timestamp 1699615441
transform 1 0 30854 0 1 -12334
box -534 -578 564 618
use TGATE_PGA_MAGIC  TGATE_PGA_MAGIC_8
timestamp 1699615441
transform 1 0 28854 0 1 -12334
box -534 -578 564 618
use TGATE_PGA_MAGIC  TGATE_PGA_MAGIC_9
timestamp 1699615441
transform 1 0 26854 0 1 -12334
box -534 -578 564 618
use TGATE_PGA_MAGIC  TGATE_PGA_MAGIC_10
timestamp 1699615441
transform 1 0 24854 0 1 -12334
box -534 -578 564 618
use TGATE_PGA_MAGIC  TGATE_PGA_MAGIC_11
timestamp 1699615441
transform 1 0 34854 0 1 -12334
box -534 -578 564 618
<< labels >>
flabel metal1 1932 4742 1932 4742 0 FreeSans 320 0 0 0 BD
port 8 nsew
flabel metal1 5335 5197 5335 5197 0 FreeSans 320 0 0 0 IND
port 10 nsew
flabel metal1 5607 5227 5607 5227 0 FreeSans 320 0 0 0 IPD
port 11 nsew
flabel psubdiffcont 8055 -1856 8055 -1856 0 FreeSans 320 0 0 0 VSS
port 12 nsew
flabel metal1 16969 2368 16969 2368 0 FreeSans 320 0 0 0 VND
port 20 nsew
flabel metal1 16707 2300 16707 2300 0 FreeSans 320 0 0 0 VPD
port 21 nsew
flabel metal1 11850 -8106 11850 -8106 0 FreeSans 320 0 0 0 VB2
port 17 nsew
flabel metal1 2007 -3925 2007 -3925 0 FreeSans 320 0 0 0 IBIAS1
port 24 nsew
flabel metal1 8109 -2826 8109 -2826 0 FreeSans 320 0 0 0 VB4
port 15 nsew
flabel metal1 11141 -7231 11141 -7231 0 FreeSans 320 0 0 0 VB3
port 18 nsew
flabel metal1 10378 -3791 10378 -3791 0 FreeSans 320 0 0 0 VOUT
port 27 nsew
flabel metal1 2651 -3832 2651 -3832 0 FreeSans 320 0 0 0 VBM
port 28 nsew
flabel metal1 6148 -4904 6148 -4904 0 FreeSans 320 0 0 0 VCD
port 29 nsew
flabel metal1 4998 -3774 4998 -3774 0 FreeSans 320 0 0 0 VBIASN
port 25 nsew
flabel metal1 14518 -3524 14518 -3524 0 FreeSans 320 0 0 0 VB1
port 19 nsew
flabel metal1 15604 -9015 15604 -9015 0 FreeSans 320 0 0 0 IBIAS3
port 34 nsew
flabel metal1 21709 -8515 21709 -8515 0 FreeSans 320 0 0 0 IBIAS4
port 33 nsew
flabel nsubdiffcont 1383 1716 1383 1716 0 FreeSans 320 0 0 0 VDD
port 3 nsew
flabel metal3 9672 -8370 9672 -8370 0 FreeSans 1600 0 0 0 IBS
port 37 nsew
flabel metal1 31192 6408 31201 6408 0 FreeSans 1600 0 0 0 OUT_P
port 38 nsew
flabel metal1 66932 3752 66932 3752 0 FreeSans 1600 0 0 0 IBIAS2
port 40 nsew
flabel metal1 -375 -1659 -375 -1659 0 FreeSans 1600 0 0 0 IBIAS
port 41 nsew
flabel metal1 10091 -3206 10091 -3206 0 FreeSans 1600 0 0 0 VCM
port 42 nsew
flabel metal3 17355 -7044 17355 -7044 0 FreeSans 800 0 0 0 IVS
port 43 nsew
flabel metal3 17372 -4830 17372 -4830 0 FreeSans 800 0 0 0 IB4
port 44 nsew
flabel metal1 2786 -7175 2786 -7175 0 FreeSans 800 0 0 0 IB2
port 45 nsew
flabel metal1 8614 -7644 8614 -7644 0 FreeSans 800 0 0 0 IB3
port 46 nsew
flabel metal2 4981 -5653 4981 -5653 0 FreeSans 800 0 0 0 IB5
port 47 nsew
flabel metal1 2226 3953 2226 3953 0 FreeSans 1600 0 0 0 IN_P
port 48 nsew
flabel metal1 2533 5090 2533 5090 0 FreeSans 1600 0 0 0 IN_N
port 49 nsew
flabel metal2 10962 2395 10962 2395 0 FreeSans 1600 0 0 0 OUT2
port 51 nsew
flabel metal1 11163 1796 11323 2518 0 FreeSans 1600 0 0 0 OUT1
port 50 nsew
flabel metal1 32154 5828 32154 5828 0 FreeSans 1600 0 0 0 OUT_N
port 39 nsew
flabel metal1 5455 -18193 5455 -18193 0 FreeSans 4800 0 0 0 VIN_P
port 52 nsew
flabel metal1 22448 -18438 22448 -18438 0 FreeSans 4800 0 0 0 VIN_N
port 53 nsew
flabel metal2 59840 -11085 59840 -11085 0 FreeSans 1600 0 0 0 S_PGA_1
port 55 nsew
flabel metal2 59593 -11442 59593 -11442 0 FreeSans 1600 0 0 0 S_PGA_2
port 56 nsew
flabel metal2 59331 -11758 59331 -11758 0 FreeSans 1600 0 0 0 S_PGA_3
port 58 nsew
<< end >>
