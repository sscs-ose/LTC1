magic
tech gf180mcuC
magscale 1 10
timestamp 1693073856
<< nwell >>
rect -1344 -1287 1344 1287
<< nsubdiff >>
rect -1320 1191 1320 1263
rect -1320 -1191 -1248 1191
rect 1248 -1191 1320 1191
rect -1320 -1263 1320 -1191
<< polysilicon >>
rect -1160 1090 -1000 1103
rect -1160 1044 -1147 1090
rect -1013 1044 -1000 1090
rect -1160 1001 -1000 1044
rect -1160 -1044 -1000 -1001
rect -1160 -1090 -1147 -1044
rect -1013 -1090 -1000 -1044
rect -1160 -1103 -1000 -1090
rect -920 1090 -760 1103
rect -920 1044 -907 1090
rect -773 1044 -760 1090
rect -920 1001 -760 1044
rect -920 -1044 -760 -1001
rect -920 -1090 -907 -1044
rect -773 -1090 -760 -1044
rect -920 -1103 -760 -1090
rect -680 1090 -520 1103
rect -680 1044 -667 1090
rect -533 1044 -520 1090
rect -680 1001 -520 1044
rect -680 -1044 -520 -1001
rect -680 -1090 -667 -1044
rect -533 -1090 -520 -1044
rect -680 -1103 -520 -1090
rect -440 1090 -280 1103
rect -440 1044 -427 1090
rect -293 1044 -280 1090
rect -440 1001 -280 1044
rect -440 -1044 -280 -1001
rect -440 -1090 -427 -1044
rect -293 -1090 -280 -1044
rect -440 -1103 -280 -1090
rect -200 1090 -40 1103
rect -200 1044 -187 1090
rect -53 1044 -40 1090
rect -200 1001 -40 1044
rect -200 -1044 -40 -1001
rect -200 -1090 -187 -1044
rect -53 -1090 -40 -1044
rect -200 -1103 -40 -1090
rect 40 1090 200 1103
rect 40 1044 53 1090
rect 187 1044 200 1090
rect 40 1001 200 1044
rect 40 -1044 200 -1001
rect 40 -1090 53 -1044
rect 187 -1090 200 -1044
rect 40 -1103 200 -1090
rect 280 1090 440 1103
rect 280 1044 293 1090
rect 427 1044 440 1090
rect 280 1001 440 1044
rect 280 -1044 440 -1001
rect 280 -1090 293 -1044
rect 427 -1090 440 -1044
rect 280 -1103 440 -1090
rect 520 1090 680 1103
rect 520 1044 533 1090
rect 667 1044 680 1090
rect 520 1001 680 1044
rect 520 -1044 680 -1001
rect 520 -1090 533 -1044
rect 667 -1090 680 -1044
rect 520 -1103 680 -1090
rect 760 1090 920 1103
rect 760 1044 773 1090
rect 907 1044 920 1090
rect 760 1001 920 1044
rect 760 -1044 920 -1001
rect 760 -1090 773 -1044
rect 907 -1090 920 -1044
rect 760 -1103 920 -1090
rect 1000 1090 1160 1103
rect 1000 1044 1013 1090
rect 1147 1044 1160 1090
rect 1000 1001 1160 1044
rect 1000 -1044 1160 -1001
rect 1000 -1090 1013 -1044
rect 1147 -1090 1160 -1044
rect 1000 -1103 1160 -1090
<< polycontact >>
rect -1147 1044 -1013 1090
rect -1147 -1090 -1013 -1044
rect -907 1044 -773 1090
rect -907 -1090 -773 -1044
rect -667 1044 -533 1090
rect -667 -1090 -533 -1044
rect -427 1044 -293 1090
rect -427 -1090 -293 -1044
rect -187 1044 -53 1090
rect -187 -1090 -53 -1044
rect 53 1044 187 1090
rect 53 -1090 187 -1044
rect 293 1044 427 1090
rect 293 -1090 427 -1044
rect 533 1044 667 1090
rect 533 -1090 667 -1044
rect 773 1044 907 1090
rect 773 -1090 907 -1044
rect 1013 1044 1147 1090
rect 1013 -1090 1147 -1044
<< ppolyres >>
rect -1160 -1001 -1000 1001
rect -920 -1001 -760 1001
rect -680 -1001 -520 1001
rect -440 -1001 -280 1001
rect -200 -1001 -40 1001
rect 40 -1001 200 1001
rect 280 -1001 440 1001
rect 520 -1001 680 1001
rect 760 -1001 920 1001
rect 1000 -1001 1160 1001
<< metal1 >>
rect -1158 1044 -1147 1090
rect -1013 1044 -1002 1090
rect -918 1044 -907 1090
rect -773 1044 -762 1090
rect -678 1044 -667 1090
rect -533 1044 -522 1090
rect -438 1044 -427 1090
rect -293 1044 -282 1090
rect -198 1044 -187 1090
rect -53 1044 -42 1090
rect 42 1044 53 1090
rect 187 1044 198 1090
rect 282 1044 293 1090
rect 427 1044 438 1090
rect 522 1044 533 1090
rect 667 1044 678 1090
rect 762 1044 773 1090
rect 907 1044 918 1090
rect 1002 1044 1013 1090
rect 1147 1044 1158 1090
rect -1158 -1090 -1147 -1044
rect -1013 -1090 -1002 -1044
rect -918 -1090 -907 -1044
rect -773 -1090 -762 -1044
rect -678 -1090 -667 -1044
rect -533 -1090 -522 -1044
rect -438 -1090 -427 -1044
rect -293 -1090 -282 -1044
rect -198 -1090 -187 -1044
rect -53 -1090 -42 -1044
rect 42 -1090 53 -1044
rect 187 -1090 198 -1044
rect 282 -1090 293 -1044
rect 427 -1090 438 -1044
rect 522 -1090 533 -1044
rect 667 -1090 678 -1044
rect 762 -1090 773 -1044
rect 907 -1090 918 -1044
rect 1002 -1090 1013 -1044
rect 1147 -1090 1158 -1044
<< properties >>
string FIXED_BBOX -1284 -1227 1284 1227
string gencell ppolyf_u
string library gf180mcu
string parameters w 0.8 l 10.01 m 1 nx 10 wmin 0.80 lmin 1.00 rho 315 val 4.319k dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0
<< end >>
