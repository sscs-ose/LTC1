magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2032 -2000 17032 72000
use 5LM_METAL_RAIL_PAD_60  5LM_METAL_RAIL_PAD_60_0
timestamp 1713338890
transform 1 0 0 0 1 0
box -32 0 15032 69968
use GF_NI_BI_T_BASE  GF_NI_BI_T_BASE_0
timestamp 1713338890
transform 1 0 -32 0 1 12430
box 0 0 15064 57570
<< labels >>
flabel metal2 s 14202 69950 14202 69950 3 FreeSans 1250 90 0 0 Y
port 1 nsew
flabel metal2 s 14069 69984 14069 69984 3 FreeSans 1250 90 0 0 OE
port 2 nsew
flabel metal2 s 13920 69958 13920 69958 3 FreeSans 1250 90 0 0 A
port 3 nsew
flabel metal2 s 13763 69972 13763 69972 3 FreeSans 1250 90 0 0 SL
port 4 nsew
flabel metal2 s 2321 69975 2321 69975 3 FreeSans 1250 90 0 0 IE
port 5 nsew
flabel metal2 s 2093 69964 2093 69964 3 FreeSans 1250 90 0 0 PD
port 6 nsew
flabel metal2 s 1603 69942 1603 69942 3 FreeSans 1250 90 0 0 PDRV1
port 7 nsew
flabel metal2 s 1463 69946 1463 69946 3 FreeSans 1250 90 0 0 PDRV0
port 8 nsew
flabel metal2 s 1217 69951 1217 69951 3 FreeSans 1250 90 0 0 PU
port 9 nsew
flabel metal2 s 704 69950 704 69950 3 FreeSans 1250 90 0 0 CS
port 10 nsew
rlabel metal5 s 785 37870 785 37870 4 DVDD
port 11 nsew
rlabel metal5 s 785 44279 785 44279 4 DVDD
port 11 nsew
rlabel metal5 s 785 67369 785 67369 4 DVDD
port 11 nsew
rlabel metal5 s 785 59534 785 59534 4 DVDD
port 11 nsew
rlabel metal5 s 785 56334 785 56334 4 DVDD
port 11 nsew
rlabel metal5 s 785 54569 785 54569 4 DVDD
port 11 nsew
rlabel metal5 s 785 53134 785 53134 4 DVDD
port 11 nsew
rlabel metal5 s 785 41888 785 41888 4 DVDD
port 11 nsew
rlabel metal5 s 785 24195 785 24195 4 DVDD
port 11 nsew
rlabel metal5 s 785 28305 785 28305 4 DVDD
port 11 nsew
rlabel metal5 s 785 31520 785 31520 4 DVDD
port 11 nsew
rlabel metal5 s 785 34634 785 34634 4 DVDD
port 11 nsew
rlabel metal4 s 785 37870 785 37870 4 DVDD
port 11 nsew
rlabel metal4 s 785 44279 785 44279 4 DVDD
port 11 nsew
rlabel metal4 s 785 67369 785 67369 4 DVDD
port 11 nsew
rlabel metal4 s 785 59534 785 59534 4 DVDD
port 11 nsew
rlabel metal4 s 785 56334 785 56334 4 DVDD
port 11 nsew
rlabel metal4 s 785 54569 785 54569 4 DVDD
port 11 nsew
rlabel metal4 s 785 53134 785 53134 4 DVDD
port 11 nsew
rlabel metal4 s 785 41888 785 41888 4 DVDD
port 11 nsew
rlabel metal4 s 785 24195 785 24195 4 DVDD
port 11 nsew
rlabel metal4 s 785 28305 785 28305 4 DVDD
port 11 nsew
rlabel metal4 s 785 31520 785 31520 4 DVDD
port 11 nsew
rlabel metal4 s 785 34634 785 34634 4 DVDD
port 11 nsew
rlabel metal3 s 785 37870 785 37870 4 DVDD
port 11 nsew
rlabel metal3 s 785 44279 785 44279 4 DVDD
port 11 nsew
rlabel metal3 s 785 67369 785 67369 4 DVDD
port 11 nsew
rlabel metal3 s 785 59534 785 59534 4 DVDD
port 11 nsew
rlabel metal3 s 785 56334 785 56334 4 DVDD
port 11 nsew
rlabel metal3 s 785 54569 785 54569 4 DVDD
port 11 nsew
rlabel metal3 s 785 53134 785 53134 4 DVDD
port 11 nsew
rlabel metal3 s 785 41888 785 41888 4 DVDD
port 11 nsew
rlabel metal3 s 785 24195 785 24195 4 DVDD
port 11 nsew
rlabel metal3 s 785 28305 785 28305 4 DVDD
port 11 nsew
rlabel metal3 s 785 31520 785 31520 4 DVDD
port 11 nsew
rlabel metal3 s 785 34634 785 34634 4 DVDD
port 11 nsew
rlabel metal5 s 716 18832 716 18832 4 DVSS
port 12 nsew
rlabel metal5 s 763 15661 763 15661 4 DVSS
port 12 nsew
rlabel metal5 s 785 47506 785 47506 4 DVSS
port 12 nsew
rlabel metal5 s 785 40253 785 40253 4 DVSS
port 12 nsew
rlabel metal5 s 785 21818 785 21818 4 DVSS
port 12 nsew
rlabel metal5 s 785 26011 785 26011 4 DVSS
port 12 nsew
rlabel metal5 s 785 57769 785 57769 4 DVSS
port 12 nsew
rlabel metal5 s 785 60969 785 60969 4 DVSS
port 12 nsew
rlabel metal5 s 785 65934 785 65934 4 DVSS
port 12 nsew
rlabel metal5 s 785 68960 785 68960 4 DVSS
port 12 nsew
rlabel metal4 s 716 18832 716 18832 4 DVSS
port 12 nsew
rlabel metal4 s 763 15661 763 15661 4 DVSS
port 12 nsew
rlabel metal4 s 785 47506 785 47506 4 DVSS
port 12 nsew
rlabel metal4 s 785 40253 785 40253 4 DVSS
port 12 nsew
rlabel metal4 s 785 21818 785 21818 4 DVSS
port 12 nsew
rlabel metal4 s 785 26011 785 26011 4 DVSS
port 12 nsew
rlabel metal4 s 785 57769 785 57769 4 DVSS
port 12 nsew
rlabel metal4 s 785 60969 785 60969 4 DVSS
port 12 nsew
rlabel metal4 s 785 65934 785 65934 4 DVSS
port 12 nsew
rlabel metal4 s 785 68960 785 68960 4 DVSS
port 12 nsew
rlabel metal3 s 716 18832 716 18832 4 DVSS
port 12 nsew
rlabel metal3 s 763 15661 763 15661 4 DVSS
port 12 nsew
rlabel metal3 s 785 47506 785 47506 4 DVSS
port 12 nsew
rlabel metal3 s 785 40253 785 40253 4 DVSS
port 12 nsew
rlabel metal3 s 785 21818 785 21818 4 DVSS
port 12 nsew
rlabel metal3 s 785 26011 785 26011 4 DVSS
port 12 nsew
rlabel metal3 s 785 57769 785 57769 4 DVSS
port 12 nsew
rlabel metal3 s 785 60969 785 60969 4 DVSS
port 12 nsew
rlabel metal3 s 785 65934 785 65934 4 DVSS
port 12 nsew
rlabel metal3 s 785 68960 785 68960 4 DVSS
port 12 nsew
rlabel metal5 s 785 51369 785 51369 4 VDD
port 13 nsew
rlabel metal5 s 785 62734 785 62734 4 VDD
port 13 nsew
rlabel metal4 s 785 51369 785 51369 4 VDD
port 13 nsew
rlabel metal4 s 785 62734 785 62734 4 VDD
port 13 nsew
rlabel metal3 s 785 51369 785 51369 4 VDD
port 13 nsew
rlabel metal3 s 785 62734 785 62734 4 VDD
port 13 nsew
rlabel metal5 s 785 64169 785 64169 4 VSS
port 14 nsew
rlabel metal5 s 785 49934 785 49934 4 VSS
port 14 nsew
rlabel metal4 s 785 64169 785 64169 4 VSS
port 14 nsew
rlabel metal4 s 785 49934 785 49934 4 VSS
port 14 nsew
rlabel metal3 s 785 64169 785 64169 4 VSS
port 14 nsew
rlabel metal3 s 785 49934 785 49934 4 VSS
port 14 nsew
rlabel metal5 s 7532 6352 7532 6352 4 PAD
port 15 nsew
<< properties >>
string FIXED_BBOX 0 0 15000 70000
<< end >>
