magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -6311 -2128 6311 2128
<< nwell >>
rect -4311 -128 4311 128
<< nsubdiff >>
rect -4228 23 4228 45
rect -4228 -23 -4206 23
rect 4206 -23 4228 23
rect -4228 -45 4228 -23
<< nsubdiffcont >>
rect -4206 -23 4206 23
<< metal1 >>
rect -4217 23 4217 34
rect -4217 -23 -4206 23
rect 4206 -23 4217 23
rect -4217 -34 4217 -23
<< end >>
