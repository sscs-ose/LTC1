magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1133 -1741 1133 1741
<< metal1 >>
rect -133 735 133 741
rect -133 709 -127 735
rect -101 709 -51 735
rect -25 709 25 735
rect 51 709 101 735
rect 127 709 133 735
rect -133 659 133 709
rect -133 633 -127 659
rect -101 633 -51 659
rect -25 633 25 659
rect 51 633 101 659
rect 127 633 133 659
rect -133 583 133 633
rect -133 557 -127 583
rect -101 557 -51 583
rect -25 557 25 583
rect 51 557 101 583
rect 127 557 133 583
rect -133 507 133 557
rect -133 481 -127 507
rect -101 481 -51 507
rect -25 481 25 507
rect 51 481 101 507
rect 127 481 133 507
rect -133 431 133 481
rect -133 405 -127 431
rect -101 405 -51 431
rect -25 405 25 431
rect 51 405 101 431
rect 127 405 133 431
rect -133 355 133 405
rect -133 329 -127 355
rect -101 329 -51 355
rect -25 329 25 355
rect 51 329 101 355
rect 127 329 133 355
rect -133 279 133 329
rect -133 253 -127 279
rect -101 253 -51 279
rect -25 253 25 279
rect 51 253 101 279
rect 127 253 133 279
rect -133 203 133 253
rect -133 177 -127 203
rect -101 177 -51 203
rect -25 177 25 203
rect 51 177 101 203
rect 127 177 133 203
rect -133 127 133 177
rect -133 101 -127 127
rect -101 101 -51 127
rect -25 101 25 127
rect 51 101 101 127
rect 127 101 133 127
rect -133 51 133 101
rect -133 25 -127 51
rect -101 25 -51 51
rect -25 25 25 51
rect 51 25 101 51
rect 127 25 133 51
rect -133 -25 133 25
rect -133 -51 -127 -25
rect -101 -51 -51 -25
rect -25 -51 25 -25
rect 51 -51 101 -25
rect 127 -51 133 -25
rect -133 -101 133 -51
rect -133 -127 -127 -101
rect -101 -127 -51 -101
rect -25 -127 25 -101
rect 51 -127 101 -101
rect 127 -127 133 -101
rect -133 -177 133 -127
rect -133 -203 -127 -177
rect -101 -203 -51 -177
rect -25 -203 25 -177
rect 51 -203 101 -177
rect 127 -203 133 -177
rect -133 -253 133 -203
rect -133 -279 -127 -253
rect -101 -279 -51 -253
rect -25 -279 25 -253
rect 51 -279 101 -253
rect 127 -279 133 -253
rect -133 -329 133 -279
rect -133 -355 -127 -329
rect -101 -355 -51 -329
rect -25 -355 25 -329
rect 51 -355 101 -329
rect 127 -355 133 -329
rect -133 -405 133 -355
rect -133 -431 -127 -405
rect -101 -431 -51 -405
rect -25 -431 25 -405
rect 51 -431 101 -405
rect 127 -431 133 -405
rect -133 -481 133 -431
rect -133 -507 -127 -481
rect -101 -507 -51 -481
rect -25 -507 25 -481
rect 51 -507 101 -481
rect 127 -507 133 -481
rect -133 -557 133 -507
rect -133 -583 -127 -557
rect -101 -583 -51 -557
rect -25 -583 25 -557
rect 51 -583 101 -557
rect 127 -583 133 -557
rect -133 -633 133 -583
rect -133 -659 -127 -633
rect -101 -659 -51 -633
rect -25 -659 25 -633
rect 51 -659 101 -633
rect 127 -659 133 -633
rect -133 -709 133 -659
rect -133 -735 -127 -709
rect -101 -735 -51 -709
rect -25 -735 25 -709
rect 51 -735 101 -709
rect 127 -735 133 -709
rect -133 -741 133 -735
<< via1 >>
rect -127 709 -101 735
rect -51 709 -25 735
rect 25 709 51 735
rect 101 709 127 735
rect -127 633 -101 659
rect -51 633 -25 659
rect 25 633 51 659
rect 101 633 127 659
rect -127 557 -101 583
rect -51 557 -25 583
rect 25 557 51 583
rect 101 557 127 583
rect -127 481 -101 507
rect -51 481 -25 507
rect 25 481 51 507
rect 101 481 127 507
rect -127 405 -101 431
rect -51 405 -25 431
rect 25 405 51 431
rect 101 405 127 431
rect -127 329 -101 355
rect -51 329 -25 355
rect 25 329 51 355
rect 101 329 127 355
rect -127 253 -101 279
rect -51 253 -25 279
rect 25 253 51 279
rect 101 253 127 279
rect -127 177 -101 203
rect -51 177 -25 203
rect 25 177 51 203
rect 101 177 127 203
rect -127 101 -101 127
rect -51 101 -25 127
rect 25 101 51 127
rect 101 101 127 127
rect -127 25 -101 51
rect -51 25 -25 51
rect 25 25 51 51
rect 101 25 127 51
rect -127 -51 -101 -25
rect -51 -51 -25 -25
rect 25 -51 51 -25
rect 101 -51 127 -25
rect -127 -127 -101 -101
rect -51 -127 -25 -101
rect 25 -127 51 -101
rect 101 -127 127 -101
rect -127 -203 -101 -177
rect -51 -203 -25 -177
rect 25 -203 51 -177
rect 101 -203 127 -177
rect -127 -279 -101 -253
rect -51 -279 -25 -253
rect 25 -279 51 -253
rect 101 -279 127 -253
rect -127 -355 -101 -329
rect -51 -355 -25 -329
rect 25 -355 51 -329
rect 101 -355 127 -329
rect -127 -431 -101 -405
rect -51 -431 -25 -405
rect 25 -431 51 -405
rect 101 -431 127 -405
rect -127 -507 -101 -481
rect -51 -507 -25 -481
rect 25 -507 51 -481
rect 101 -507 127 -481
rect -127 -583 -101 -557
rect -51 -583 -25 -557
rect 25 -583 51 -557
rect 101 -583 127 -557
rect -127 -659 -101 -633
rect -51 -659 -25 -633
rect 25 -659 51 -633
rect 101 -659 127 -633
rect -127 -735 -101 -709
rect -51 -735 -25 -709
rect 25 -735 51 -709
rect 101 -735 127 -709
<< metal2 >>
rect -133 735 133 741
rect -133 709 -127 735
rect -101 709 -51 735
rect -25 709 25 735
rect 51 709 101 735
rect 127 709 133 735
rect -133 659 133 709
rect -133 633 -127 659
rect -101 633 -51 659
rect -25 633 25 659
rect 51 633 101 659
rect 127 633 133 659
rect -133 583 133 633
rect -133 557 -127 583
rect -101 557 -51 583
rect -25 557 25 583
rect 51 557 101 583
rect 127 557 133 583
rect -133 507 133 557
rect -133 481 -127 507
rect -101 481 -51 507
rect -25 481 25 507
rect 51 481 101 507
rect 127 481 133 507
rect -133 431 133 481
rect -133 405 -127 431
rect -101 405 -51 431
rect -25 405 25 431
rect 51 405 101 431
rect 127 405 133 431
rect -133 355 133 405
rect -133 329 -127 355
rect -101 329 -51 355
rect -25 329 25 355
rect 51 329 101 355
rect 127 329 133 355
rect -133 279 133 329
rect -133 253 -127 279
rect -101 253 -51 279
rect -25 253 25 279
rect 51 253 101 279
rect 127 253 133 279
rect -133 203 133 253
rect -133 177 -127 203
rect -101 177 -51 203
rect -25 177 25 203
rect 51 177 101 203
rect 127 177 133 203
rect -133 127 133 177
rect -133 101 -127 127
rect -101 101 -51 127
rect -25 101 25 127
rect 51 101 101 127
rect 127 101 133 127
rect -133 51 133 101
rect -133 25 -127 51
rect -101 25 -51 51
rect -25 25 25 51
rect 51 25 101 51
rect 127 25 133 51
rect -133 -25 133 25
rect -133 -51 -127 -25
rect -101 -51 -51 -25
rect -25 -51 25 -25
rect 51 -51 101 -25
rect 127 -51 133 -25
rect -133 -101 133 -51
rect -133 -127 -127 -101
rect -101 -127 -51 -101
rect -25 -127 25 -101
rect 51 -127 101 -101
rect 127 -127 133 -101
rect -133 -177 133 -127
rect -133 -203 -127 -177
rect -101 -203 -51 -177
rect -25 -203 25 -177
rect 51 -203 101 -177
rect 127 -203 133 -177
rect -133 -253 133 -203
rect -133 -279 -127 -253
rect -101 -279 -51 -253
rect -25 -279 25 -253
rect 51 -279 101 -253
rect 127 -279 133 -253
rect -133 -329 133 -279
rect -133 -355 -127 -329
rect -101 -355 -51 -329
rect -25 -355 25 -329
rect 51 -355 101 -329
rect 127 -355 133 -329
rect -133 -405 133 -355
rect -133 -431 -127 -405
rect -101 -431 -51 -405
rect -25 -431 25 -405
rect 51 -431 101 -405
rect 127 -431 133 -405
rect -133 -481 133 -431
rect -133 -507 -127 -481
rect -101 -507 -51 -481
rect -25 -507 25 -481
rect 51 -507 101 -481
rect 127 -507 133 -481
rect -133 -557 133 -507
rect -133 -583 -127 -557
rect -101 -583 -51 -557
rect -25 -583 25 -557
rect 51 -583 101 -557
rect 127 -583 133 -557
rect -133 -633 133 -583
rect -133 -659 -127 -633
rect -101 -659 -51 -633
rect -25 -659 25 -633
rect 51 -659 101 -633
rect 127 -659 133 -633
rect -133 -709 133 -659
rect -133 -735 -127 -709
rect -101 -735 -51 -709
rect -25 -735 25 -709
rect 51 -735 101 -709
rect 127 -735 133 -709
rect -133 -741 133 -735
<< end >>
