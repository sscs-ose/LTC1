magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -3626 -1382 3626 1382
<< metal1 >>
rect -2626 376 2626 382
rect -2626 350 -2620 376
rect -2594 350 -2554 376
rect -2528 350 -2488 376
rect -2462 350 -2422 376
rect -2396 350 -2356 376
rect -2330 350 -2290 376
rect -2264 350 -2224 376
rect -2198 350 -2158 376
rect -2132 350 -2092 376
rect -2066 350 -2026 376
rect -2000 350 -1960 376
rect -1934 350 -1894 376
rect -1868 350 -1828 376
rect -1802 350 -1762 376
rect -1736 350 -1696 376
rect -1670 350 -1630 376
rect -1604 350 -1564 376
rect -1538 350 -1498 376
rect -1472 350 -1432 376
rect -1406 350 -1366 376
rect -1340 350 -1300 376
rect -1274 350 -1234 376
rect -1208 350 -1168 376
rect -1142 350 -1102 376
rect -1076 350 -1036 376
rect -1010 350 -970 376
rect -944 350 -904 376
rect -878 350 -838 376
rect -812 350 -772 376
rect -746 350 -706 376
rect -680 350 -640 376
rect -614 350 -574 376
rect -548 350 -508 376
rect -482 350 -442 376
rect -416 350 -376 376
rect -350 350 -310 376
rect -284 350 -244 376
rect -218 350 -178 376
rect -152 350 -112 376
rect -86 350 -46 376
rect -20 350 20 376
rect 46 350 86 376
rect 112 350 152 376
rect 178 350 218 376
rect 244 350 284 376
rect 310 350 350 376
rect 376 350 416 376
rect 442 350 482 376
rect 508 350 548 376
rect 574 350 614 376
rect 640 350 680 376
rect 706 350 746 376
rect 772 350 812 376
rect 838 350 878 376
rect 904 350 944 376
rect 970 350 1010 376
rect 1036 350 1076 376
rect 1102 350 1142 376
rect 1168 350 1208 376
rect 1234 350 1274 376
rect 1300 350 1340 376
rect 1366 350 1406 376
rect 1432 350 1472 376
rect 1498 350 1538 376
rect 1564 350 1604 376
rect 1630 350 1670 376
rect 1696 350 1736 376
rect 1762 350 1802 376
rect 1828 350 1868 376
rect 1894 350 1934 376
rect 1960 350 2000 376
rect 2026 350 2066 376
rect 2092 350 2132 376
rect 2158 350 2198 376
rect 2224 350 2264 376
rect 2290 350 2330 376
rect 2356 350 2396 376
rect 2422 350 2462 376
rect 2488 350 2528 376
rect 2554 350 2594 376
rect 2620 350 2626 376
rect -2626 310 2626 350
rect -2626 284 -2620 310
rect -2594 284 -2554 310
rect -2528 284 -2488 310
rect -2462 284 -2422 310
rect -2396 284 -2356 310
rect -2330 284 -2290 310
rect -2264 284 -2224 310
rect -2198 284 -2158 310
rect -2132 284 -2092 310
rect -2066 284 -2026 310
rect -2000 284 -1960 310
rect -1934 284 -1894 310
rect -1868 284 -1828 310
rect -1802 284 -1762 310
rect -1736 284 -1696 310
rect -1670 284 -1630 310
rect -1604 284 -1564 310
rect -1538 284 -1498 310
rect -1472 284 -1432 310
rect -1406 284 -1366 310
rect -1340 284 -1300 310
rect -1274 284 -1234 310
rect -1208 284 -1168 310
rect -1142 284 -1102 310
rect -1076 284 -1036 310
rect -1010 284 -970 310
rect -944 284 -904 310
rect -878 284 -838 310
rect -812 284 -772 310
rect -746 284 -706 310
rect -680 284 -640 310
rect -614 284 -574 310
rect -548 284 -508 310
rect -482 284 -442 310
rect -416 284 -376 310
rect -350 284 -310 310
rect -284 284 -244 310
rect -218 284 -178 310
rect -152 284 -112 310
rect -86 284 -46 310
rect -20 284 20 310
rect 46 284 86 310
rect 112 284 152 310
rect 178 284 218 310
rect 244 284 284 310
rect 310 284 350 310
rect 376 284 416 310
rect 442 284 482 310
rect 508 284 548 310
rect 574 284 614 310
rect 640 284 680 310
rect 706 284 746 310
rect 772 284 812 310
rect 838 284 878 310
rect 904 284 944 310
rect 970 284 1010 310
rect 1036 284 1076 310
rect 1102 284 1142 310
rect 1168 284 1208 310
rect 1234 284 1274 310
rect 1300 284 1340 310
rect 1366 284 1406 310
rect 1432 284 1472 310
rect 1498 284 1538 310
rect 1564 284 1604 310
rect 1630 284 1670 310
rect 1696 284 1736 310
rect 1762 284 1802 310
rect 1828 284 1868 310
rect 1894 284 1934 310
rect 1960 284 2000 310
rect 2026 284 2066 310
rect 2092 284 2132 310
rect 2158 284 2198 310
rect 2224 284 2264 310
rect 2290 284 2330 310
rect 2356 284 2396 310
rect 2422 284 2462 310
rect 2488 284 2528 310
rect 2554 284 2594 310
rect 2620 284 2626 310
rect -2626 244 2626 284
rect -2626 218 -2620 244
rect -2594 218 -2554 244
rect -2528 218 -2488 244
rect -2462 218 -2422 244
rect -2396 218 -2356 244
rect -2330 218 -2290 244
rect -2264 218 -2224 244
rect -2198 218 -2158 244
rect -2132 218 -2092 244
rect -2066 218 -2026 244
rect -2000 218 -1960 244
rect -1934 218 -1894 244
rect -1868 218 -1828 244
rect -1802 218 -1762 244
rect -1736 218 -1696 244
rect -1670 218 -1630 244
rect -1604 218 -1564 244
rect -1538 218 -1498 244
rect -1472 218 -1432 244
rect -1406 218 -1366 244
rect -1340 218 -1300 244
rect -1274 218 -1234 244
rect -1208 218 -1168 244
rect -1142 218 -1102 244
rect -1076 218 -1036 244
rect -1010 218 -970 244
rect -944 218 -904 244
rect -878 218 -838 244
rect -812 218 -772 244
rect -746 218 -706 244
rect -680 218 -640 244
rect -614 218 -574 244
rect -548 218 -508 244
rect -482 218 -442 244
rect -416 218 -376 244
rect -350 218 -310 244
rect -284 218 -244 244
rect -218 218 -178 244
rect -152 218 -112 244
rect -86 218 -46 244
rect -20 218 20 244
rect 46 218 86 244
rect 112 218 152 244
rect 178 218 218 244
rect 244 218 284 244
rect 310 218 350 244
rect 376 218 416 244
rect 442 218 482 244
rect 508 218 548 244
rect 574 218 614 244
rect 640 218 680 244
rect 706 218 746 244
rect 772 218 812 244
rect 838 218 878 244
rect 904 218 944 244
rect 970 218 1010 244
rect 1036 218 1076 244
rect 1102 218 1142 244
rect 1168 218 1208 244
rect 1234 218 1274 244
rect 1300 218 1340 244
rect 1366 218 1406 244
rect 1432 218 1472 244
rect 1498 218 1538 244
rect 1564 218 1604 244
rect 1630 218 1670 244
rect 1696 218 1736 244
rect 1762 218 1802 244
rect 1828 218 1868 244
rect 1894 218 1934 244
rect 1960 218 2000 244
rect 2026 218 2066 244
rect 2092 218 2132 244
rect 2158 218 2198 244
rect 2224 218 2264 244
rect 2290 218 2330 244
rect 2356 218 2396 244
rect 2422 218 2462 244
rect 2488 218 2528 244
rect 2554 218 2594 244
rect 2620 218 2626 244
rect -2626 178 2626 218
rect -2626 152 -2620 178
rect -2594 152 -2554 178
rect -2528 152 -2488 178
rect -2462 152 -2422 178
rect -2396 152 -2356 178
rect -2330 152 -2290 178
rect -2264 152 -2224 178
rect -2198 152 -2158 178
rect -2132 152 -2092 178
rect -2066 152 -2026 178
rect -2000 152 -1960 178
rect -1934 152 -1894 178
rect -1868 152 -1828 178
rect -1802 152 -1762 178
rect -1736 152 -1696 178
rect -1670 152 -1630 178
rect -1604 152 -1564 178
rect -1538 152 -1498 178
rect -1472 152 -1432 178
rect -1406 152 -1366 178
rect -1340 152 -1300 178
rect -1274 152 -1234 178
rect -1208 152 -1168 178
rect -1142 152 -1102 178
rect -1076 152 -1036 178
rect -1010 152 -970 178
rect -944 152 -904 178
rect -878 152 -838 178
rect -812 152 -772 178
rect -746 152 -706 178
rect -680 152 -640 178
rect -614 152 -574 178
rect -548 152 -508 178
rect -482 152 -442 178
rect -416 152 -376 178
rect -350 152 -310 178
rect -284 152 -244 178
rect -218 152 -178 178
rect -152 152 -112 178
rect -86 152 -46 178
rect -20 152 20 178
rect 46 152 86 178
rect 112 152 152 178
rect 178 152 218 178
rect 244 152 284 178
rect 310 152 350 178
rect 376 152 416 178
rect 442 152 482 178
rect 508 152 548 178
rect 574 152 614 178
rect 640 152 680 178
rect 706 152 746 178
rect 772 152 812 178
rect 838 152 878 178
rect 904 152 944 178
rect 970 152 1010 178
rect 1036 152 1076 178
rect 1102 152 1142 178
rect 1168 152 1208 178
rect 1234 152 1274 178
rect 1300 152 1340 178
rect 1366 152 1406 178
rect 1432 152 1472 178
rect 1498 152 1538 178
rect 1564 152 1604 178
rect 1630 152 1670 178
rect 1696 152 1736 178
rect 1762 152 1802 178
rect 1828 152 1868 178
rect 1894 152 1934 178
rect 1960 152 2000 178
rect 2026 152 2066 178
rect 2092 152 2132 178
rect 2158 152 2198 178
rect 2224 152 2264 178
rect 2290 152 2330 178
rect 2356 152 2396 178
rect 2422 152 2462 178
rect 2488 152 2528 178
rect 2554 152 2594 178
rect 2620 152 2626 178
rect -2626 112 2626 152
rect -2626 86 -2620 112
rect -2594 86 -2554 112
rect -2528 86 -2488 112
rect -2462 86 -2422 112
rect -2396 86 -2356 112
rect -2330 86 -2290 112
rect -2264 86 -2224 112
rect -2198 86 -2158 112
rect -2132 86 -2092 112
rect -2066 86 -2026 112
rect -2000 86 -1960 112
rect -1934 86 -1894 112
rect -1868 86 -1828 112
rect -1802 86 -1762 112
rect -1736 86 -1696 112
rect -1670 86 -1630 112
rect -1604 86 -1564 112
rect -1538 86 -1498 112
rect -1472 86 -1432 112
rect -1406 86 -1366 112
rect -1340 86 -1300 112
rect -1274 86 -1234 112
rect -1208 86 -1168 112
rect -1142 86 -1102 112
rect -1076 86 -1036 112
rect -1010 86 -970 112
rect -944 86 -904 112
rect -878 86 -838 112
rect -812 86 -772 112
rect -746 86 -706 112
rect -680 86 -640 112
rect -614 86 -574 112
rect -548 86 -508 112
rect -482 86 -442 112
rect -416 86 -376 112
rect -350 86 -310 112
rect -284 86 -244 112
rect -218 86 -178 112
rect -152 86 -112 112
rect -86 86 -46 112
rect -20 86 20 112
rect 46 86 86 112
rect 112 86 152 112
rect 178 86 218 112
rect 244 86 284 112
rect 310 86 350 112
rect 376 86 416 112
rect 442 86 482 112
rect 508 86 548 112
rect 574 86 614 112
rect 640 86 680 112
rect 706 86 746 112
rect 772 86 812 112
rect 838 86 878 112
rect 904 86 944 112
rect 970 86 1010 112
rect 1036 86 1076 112
rect 1102 86 1142 112
rect 1168 86 1208 112
rect 1234 86 1274 112
rect 1300 86 1340 112
rect 1366 86 1406 112
rect 1432 86 1472 112
rect 1498 86 1538 112
rect 1564 86 1604 112
rect 1630 86 1670 112
rect 1696 86 1736 112
rect 1762 86 1802 112
rect 1828 86 1868 112
rect 1894 86 1934 112
rect 1960 86 2000 112
rect 2026 86 2066 112
rect 2092 86 2132 112
rect 2158 86 2198 112
rect 2224 86 2264 112
rect 2290 86 2330 112
rect 2356 86 2396 112
rect 2422 86 2462 112
rect 2488 86 2528 112
rect 2554 86 2594 112
rect 2620 86 2626 112
rect -2626 46 2626 86
rect -2626 20 -2620 46
rect -2594 20 -2554 46
rect -2528 20 -2488 46
rect -2462 20 -2422 46
rect -2396 20 -2356 46
rect -2330 20 -2290 46
rect -2264 20 -2224 46
rect -2198 20 -2158 46
rect -2132 20 -2092 46
rect -2066 20 -2026 46
rect -2000 20 -1960 46
rect -1934 20 -1894 46
rect -1868 20 -1828 46
rect -1802 20 -1762 46
rect -1736 20 -1696 46
rect -1670 20 -1630 46
rect -1604 20 -1564 46
rect -1538 20 -1498 46
rect -1472 20 -1432 46
rect -1406 20 -1366 46
rect -1340 20 -1300 46
rect -1274 20 -1234 46
rect -1208 20 -1168 46
rect -1142 20 -1102 46
rect -1076 20 -1036 46
rect -1010 20 -970 46
rect -944 20 -904 46
rect -878 20 -838 46
rect -812 20 -772 46
rect -746 20 -706 46
rect -680 20 -640 46
rect -614 20 -574 46
rect -548 20 -508 46
rect -482 20 -442 46
rect -416 20 -376 46
rect -350 20 -310 46
rect -284 20 -244 46
rect -218 20 -178 46
rect -152 20 -112 46
rect -86 20 -46 46
rect -20 20 20 46
rect 46 20 86 46
rect 112 20 152 46
rect 178 20 218 46
rect 244 20 284 46
rect 310 20 350 46
rect 376 20 416 46
rect 442 20 482 46
rect 508 20 548 46
rect 574 20 614 46
rect 640 20 680 46
rect 706 20 746 46
rect 772 20 812 46
rect 838 20 878 46
rect 904 20 944 46
rect 970 20 1010 46
rect 1036 20 1076 46
rect 1102 20 1142 46
rect 1168 20 1208 46
rect 1234 20 1274 46
rect 1300 20 1340 46
rect 1366 20 1406 46
rect 1432 20 1472 46
rect 1498 20 1538 46
rect 1564 20 1604 46
rect 1630 20 1670 46
rect 1696 20 1736 46
rect 1762 20 1802 46
rect 1828 20 1868 46
rect 1894 20 1934 46
rect 1960 20 2000 46
rect 2026 20 2066 46
rect 2092 20 2132 46
rect 2158 20 2198 46
rect 2224 20 2264 46
rect 2290 20 2330 46
rect 2356 20 2396 46
rect 2422 20 2462 46
rect 2488 20 2528 46
rect 2554 20 2594 46
rect 2620 20 2626 46
rect -2626 -20 2626 20
rect -2626 -46 -2620 -20
rect -2594 -46 -2554 -20
rect -2528 -46 -2488 -20
rect -2462 -46 -2422 -20
rect -2396 -46 -2356 -20
rect -2330 -46 -2290 -20
rect -2264 -46 -2224 -20
rect -2198 -46 -2158 -20
rect -2132 -46 -2092 -20
rect -2066 -46 -2026 -20
rect -2000 -46 -1960 -20
rect -1934 -46 -1894 -20
rect -1868 -46 -1828 -20
rect -1802 -46 -1762 -20
rect -1736 -46 -1696 -20
rect -1670 -46 -1630 -20
rect -1604 -46 -1564 -20
rect -1538 -46 -1498 -20
rect -1472 -46 -1432 -20
rect -1406 -46 -1366 -20
rect -1340 -46 -1300 -20
rect -1274 -46 -1234 -20
rect -1208 -46 -1168 -20
rect -1142 -46 -1102 -20
rect -1076 -46 -1036 -20
rect -1010 -46 -970 -20
rect -944 -46 -904 -20
rect -878 -46 -838 -20
rect -812 -46 -772 -20
rect -746 -46 -706 -20
rect -680 -46 -640 -20
rect -614 -46 -574 -20
rect -548 -46 -508 -20
rect -482 -46 -442 -20
rect -416 -46 -376 -20
rect -350 -46 -310 -20
rect -284 -46 -244 -20
rect -218 -46 -178 -20
rect -152 -46 -112 -20
rect -86 -46 -46 -20
rect -20 -46 20 -20
rect 46 -46 86 -20
rect 112 -46 152 -20
rect 178 -46 218 -20
rect 244 -46 284 -20
rect 310 -46 350 -20
rect 376 -46 416 -20
rect 442 -46 482 -20
rect 508 -46 548 -20
rect 574 -46 614 -20
rect 640 -46 680 -20
rect 706 -46 746 -20
rect 772 -46 812 -20
rect 838 -46 878 -20
rect 904 -46 944 -20
rect 970 -46 1010 -20
rect 1036 -46 1076 -20
rect 1102 -46 1142 -20
rect 1168 -46 1208 -20
rect 1234 -46 1274 -20
rect 1300 -46 1340 -20
rect 1366 -46 1406 -20
rect 1432 -46 1472 -20
rect 1498 -46 1538 -20
rect 1564 -46 1604 -20
rect 1630 -46 1670 -20
rect 1696 -46 1736 -20
rect 1762 -46 1802 -20
rect 1828 -46 1868 -20
rect 1894 -46 1934 -20
rect 1960 -46 2000 -20
rect 2026 -46 2066 -20
rect 2092 -46 2132 -20
rect 2158 -46 2198 -20
rect 2224 -46 2264 -20
rect 2290 -46 2330 -20
rect 2356 -46 2396 -20
rect 2422 -46 2462 -20
rect 2488 -46 2528 -20
rect 2554 -46 2594 -20
rect 2620 -46 2626 -20
rect -2626 -86 2626 -46
rect -2626 -112 -2620 -86
rect -2594 -112 -2554 -86
rect -2528 -112 -2488 -86
rect -2462 -112 -2422 -86
rect -2396 -112 -2356 -86
rect -2330 -112 -2290 -86
rect -2264 -112 -2224 -86
rect -2198 -112 -2158 -86
rect -2132 -112 -2092 -86
rect -2066 -112 -2026 -86
rect -2000 -112 -1960 -86
rect -1934 -112 -1894 -86
rect -1868 -112 -1828 -86
rect -1802 -112 -1762 -86
rect -1736 -112 -1696 -86
rect -1670 -112 -1630 -86
rect -1604 -112 -1564 -86
rect -1538 -112 -1498 -86
rect -1472 -112 -1432 -86
rect -1406 -112 -1366 -86
rect -1340 -112 -1300 -86
rect -1274 -112 -1234 -86
rect -1208 -112 -1168 -86
rect -1142 -112 -1102 -86
rect -1076 -112 -1036 -86
rect -1010 -112 -970 -86
rect -944 -112 -904 -86
rect -878 -112 -838 -86
rect -812 -112 -772 -86
rect -746 -112 -706 -86
rect -680 -112 -640 -86
rect -614 -112 -574 -86
rect -548 -112 -508 -86
rect -482 -112 -442 -86
rect -416 -112 -376 -86
rect -350 -112 -310 -86
rect -284 -112 -244 -86
rect -218 -112 -178 -86
rect -152 -112 -112 -86
rect -86 -112 -46 -86
rect -20 -112 20 -86
rect 46 -112 86 -86
rect 112 -112 152 -86
rect 178 -112 218 -86
rect 244 -112 284 -86
rect 310 -112 350 -86
rect 376 -112 416 -86
rect 442 -112 482 -86
rect 508 -112 548 -86
rect 574 -112 614 -86
rect 640 -112 680 -86
rect 706 -112 746 -86
rect 772 -112 812 -86
rect 838 -112 878 -86
rect 904 -112 944 -86
rect 970 -112 1010 -86
rect 1036 -112 1076 -86
rect 1102 -112 1142 -86
rect 1168 -112 1208 -86
rect 1234 -112 1274 -86
rect 1300 -112 1340 -86
rect 1366 -112 1406 -86
rect 1432 -112 1472 -86
rect 1498 -112 1538 -86
rect 1564 -112 1604 -86
rect 1630 -112 1670 -86
rect 1696 -112 1736 -86
rect 1762 -112 1802 -86
rect 1828 -112 1868 -86
rect 1894 -112 1934 -86
rect 1960 -112 2000 -86
rect 2026 -112 2066 -86
rect 2092 -112 2132 -86
rect 2158 -112 2198 -86
rect 2224 -112 2264 -86
rect 2290 -112 2330 -86
rect 2356 -112 2396 -86
rect 2422 -112 2462 -86
rect 2488 -112 2528 -86
rect 2554 -112 2594 -86
rect 2620 -112 2626 -86
rect -2626 -152 2626 -112
rect -2626 -178 -2620 -152
rect -2594 -178 -2554 -152
rect -2528 -178 -2488 -152
rect -2462 -178 -2422 -152
rect -2396 -178 -2356 -152
rect -2330 -178 -2290 -152
rect -2264 -178 -2224 -152
rect -2198 -178 -2158 -152
rect -2132 -178 -2092 -152
rect -2066 -178 -2026 -152
rect -2000 -178 -1960 -152
rect -1934 -178 -1894 -152
rect -1868 -178 -1828 -152
rect -1802 -178 -1762 -152
rect -1736 -178 -1696 -152
rect -1670 -178 -1630 -152
rect -1604 -178 -1564 -152
rect -1538 -178 -1498 -152
rect -1472 -178 -1432 -152
rect -1406 -178 -1366 -152
rect -1340 -178 -1300 -152
rect -1274 -178 -1234 -152
rect -1208 -178 -1168 -152
rect -1142 -178 -1102 -152
rect -1076 -178 -1036 -152
rect -1010 -178 -970 -152
rect -944 -178 -904 -152
rect -878 -178 -838 -152
rect -812 -178 -772 -152
rect -746 -178 -706 -152
rect -680 -178 -640 -152
rect -614 -178 -574 -152
rect -548 -178 -508 -152
rect -482 -178 -442 -152
rect -416 -178 -376 -152
rect -350 -178 -310 -152
rect -284 -178 -244 -152
rect -218 -178 -178 -152
rect -152 -178 -112 -152
rect -86 -178 -46 -152
rect -20 -178 20 -152
rect 46 -178 86 -152
rect 112 -178 152 -152
rect 178 -178 218 -152
rect 244 -178 284 -152
rect 310 -178 350 -152
rect 376 -178 416 -152
rect 442 -178 482 -152
rect 508 -178 548 -152
rect 574 -178 614 -152
rect 640 -178 680 -152
rect 706 -178 746 -152
rect 772 -178 812 -152
rect 838 -178 878 -152
rect 904 -178 944 -152
rect 970 -178 1010 -152
rect 1036 -178 1076 -152
rect 1102 -178 1142 -152
rect 1168 -178 1208 -152
rect 1234 -178 1274 -152
rect 1300 -178 1340 -152
rect 1366 -178 1406 -152
rect 1432 -178 1472 -152
rect 1498 -178 1538 -152
rect 1564 -178 1604 -152
rect 1630 -178 1670 -152
rect 1696 -178 1736 -152
rect 1762 -178 1802 -152
rect 1828 -178 1868 -152
rect 1894 -178 1934 -152
rect 1960 -178 2000 -152
rect 2026 -178 2066 -152
rect 2092 -178 2132 -152
rect 2158 -178 2198 -152
rect 2224 -178 2264 -152
rect 2290 -178 2330 -152
rect 2356 -178 2396 -152
rect 2422 -178 2462 -152
rect 2488 -178 2528 -152
rect 2554 -178 2594 -152
rect 2620 -178 2626 -152
rect -2626 -218 2626 -178
rect -2626 -244 -2620 -218
rect -2594 -244 -2554 -218
rect -2528 -244 -2488 -218
rect -2462 -244 -2422 -218
rect -2396 -244 -2356 -218
rect -2330 -244 -2290 -218
rect -2264 -244 -2224 -218
rect -2198 -244 -2158 -218
rect -2132 -244 -2092 -218
rect -2066 -244 -2026 -218
rect -2000 -244 -1960 -218
rect -1934 -244 -1894 -218
rect -1868 -244 -1828 -218
rect -1802 -244 -1762 -218
rect -1736 -244 -1696 -218
rect -1670 -244 -1630 -218
rect -1604 -244 -1564 -218
rect -1538 -244 -1498 -218
rect -1472 -244 -1432 -218
rect -1406 -244 -1366 -218
rect -1340 -244 -1300 -218
rect -1274 -244 -1234 -218
rect -1208 -244 -1168 -218
rect -1142 -244 -1102 -218
rect -1076 -244 -1036 -218
rect -1010 -244 -970 -218
rect -944 -244 -904 -218
rect -878 -244 -838 -218
rect -812 -244 -772 -218
rect -746 -244 -706 -218
rect -680 -244 -640 -218
rect -614 -244 -574 -218
rect -548 -244 -508 -218
rect -482 -244 -442 -218
rect -416 -244 -376 -218
rect -350 -244 -310 -218
rect -284 -244 -244 -218
rect -218 -244 -178 -218
rect -152 -244 -112 -218
rect -86 -244 -46 -218
rect -20 -244 20 -218
rect 46 -244 86 -218
rect 112 -244 152 -218
rect 178 -244 218 -218
rect 244 -244 284 -218
rect 310 -244 350 -218
rect 376 -244 416 -218
rect 442 -244 482 -218
rect 508 -244 548 -218
rect 574 -244 614 -218
rect 640 -244 680 -218
rect 706 -244 746 -218
rect 772 -244 812 -218
rect 838 -244 878 -218
rect 904 -244 944 -218
rect 970 -244 1010 -218
rect 1036 -244 1076 -218
rect 1102 -244 1142 -218
rect 1168 -244 1208 -218
rect 1234 -244 1274 -218
rect 1300 -244 1340 -218
rect 1366 -244 1406 -218
rect 1432 -244 1472 -218
rect 1498 -244 1538 -218
rect 1564 -244 1604 -218
rect 1630 -244 1670 -218
rect 1696 -244 1736 -218
rect 1762 -244 1802 -218
rect 1828 -244 1868 -218
rect 1894 -244 1934 -218
rect 1960 -244 2000 -218
rect 2026 -244 2066 -218
rect 2092 -244 2132 -218
rect 2158 -244 2198 -218
rect 2224 -244 2264 -218
rect 2290 -244 2330 -218
rect 2356 -244 2396 -218
rect 2422 -244 2462 -218
rect 2488 -244 2528 -218
rect 2554 -244 2594 -218
rect 2620 -244 2626 -218
rect -2626 -284 2626 -244
rect -2626 -310 -2620 -284
rect -2594 -310 -2554 -284
rect -2528 -310 -2488 -284
rect -2462 -310 -2422 -284
rect -2396 -310 -2356 -284
rect -2330 -310 -2290 -284
rect -2264 -310 -2224 -284
rect -2198 -310 -2158 -284
rect -2132 -310 -2092 -284
rect -2066 -310 -2026 -284
rect -2000 -310 -1960 -284
rect -1934 -310 -1894 -284
rect -1868 -310 -1828 -284
rect -1802 -310 -1762 -284
rect -1736 -310 -1696 -284
rect -1670 -310 -1630 -284
rect -1604 -310 -1564 -284
rect -1538 -310 -1498 -284
rect -1472 -310 -1432 -284
rect -1406 -310 -1366 -284
rect -1340 -310 -1300 -284
rect -1274 -310 -1234 -284
rect -1208 -310 -1168 -284
rect -1142 -310 -1102 -284
rect -1076 -310 -1036 -284
rect -1010 -310 -970 -284
rect -944 -310 -904 -284
rect -878 -310 -838 -284
rect -812 -310 -772 -284
rect -746 -310 -706 -284
rect -680 -310 -640 -284
rect -614 -310 -574 -284
rect -548 -310 -508 -284
rect -482 -310 -442 -284
rect -416 -310 -376 -284
rect -350 -310 -310 -284
rect -284 -310 -244 -284
rect -218 -310 -178 -284
rect -152 -310 -112 -284
rect -86 -310 -46 -284
rect -20 -310 20 -284
rect 46 -310 86 -284
rect 112 -310 152 -284
rect 178 -310 218 -284
rect 244 -310 284 -284
rect 310 -310 350 -284
rect 376 -310 416 -284
rect 442 -310 482 -284
rect 508 -310 548 -284
rect 574 -310 614 -284
rect 640 -310 680 -284
rect 706 -310 746 -284
rect 772 -310 812 -284
rect 838 -310 878 -284
rect 904 -310 944 -284
rect 970 -310 1010 -284
rect 1036 -310 1076 -284
rect 1102 -310 1142 -284
rect 1168 -310 1208 -284
rect 1234 -310 1274 -284
rect 1300 -310 1340 -284
rect 1366 -310 1406 -284
rect 1432 -310 1472 -284
rect 1498 -310 1538 -284
rect 1564 -310 1604 -284
rect 1630 -310 1670 -284
rect 1696 -310 1736 -284
rect 1762 -310 1802 -284
rect 1828 -310 1868 -284
rect 1894 -310 1934 -284
rect 1960 -310 2000 -284
rect 2026 -310 2066 -284
rect 2092 -310 2132 -284
rect 2158 -310 2198 -284
rect 2224 -310 2264 -284
rect 2290 -310 2330 -284
rect 2356 -310 2396 -284
rect 2422 -310 2462 -284
rect 2488 -310 2528 -284
rect 2554 -310 2594 -284
rect 2620 -310 2626 -284
rect -2626 -350 2626 -310
rect -2626 -376 -2620 -350
rect -2594 -376 -2554 -350
rect -2528 -376 -2488 -350
rect -2462 -376 -2422 -350
rect -2396 -376 -2356 -350
rect -2330 -376 -2290 -350
rect -2264 -376 -2224 -350
rect -2198 -376 -2158 -350
rect -2132 -376 -2092 -350
rect -2066 -376 -2026 -350
rect -2000 -376 -1960 -350
rect -1934 -376 -1894 -350
rect -1868 -376 -1828 -350
rect -1802 -376 -1762 -350
rect -1736 -376 -1696 -350
rect -1670 -376 -1630 -350
rect -1604 -376 -1564 -350
rect -1538 -376 -1498 -350
rect -1472 -376 -1432 -350
rect -1406 -376 -1366 -350
rect -1340 -376 -1300 -350
rect -1274 -376 -1234 -350
rect -1208 -376 -1168 -350
rect -1142 -376 -1102 -350
rect -1076 -376 -1036 -350
rect -1010 -376 -970 -350
rect -944 -376 -904 -350
rect -878 -376 -838 -350
rect -812 -376 -772 -350
rect -746 -376 -706 -350
rect -680 -376 -640 -350
rect -614 -376 -574 -350
rect -548 -376 -508 -350
rect -482 -376 -442 -350
rect -416 -376 -376 -350
rect -350 -376 -310 -350
rect -284 -376 -244 -350
rect -218 -376 -178 -350
rect -152 -376 -112 -350
rect -86 -376 -46 -350
rect -20 -376 20 -350
rect 46 -376 86 -350
rect 112 -376 152 -350
rect 178 -376 218 -350
rect 244 -376 284 -350
rect 310 -376 350 -350
rect 376 -376 416 -350
rect 442 -376 482 -350
rect 508 -376 548 -350
rect 574 -376 614 -350
rect 640 -376 680 -350
rect 706 -376 746 -350
rect 772 -376 812 -350
rect 838 -376 878 -350
rect 904 -376 944 -350
rect 970 -376 1010 -350
rect 1036 -376 1076 -350
rect 1102 -376 1142 -350
rect 1168 -376 1208 -350
rect 1234 -376 1274 -350
rect 1300 -376 1340 -350
rect 1366 -376 1406 -350
rect 1432 -376 1472 -350
rect 1498 -376 1538 -350
rect 1564 -376 1604 -350
rect 1630 -376 1670 -350
rect 1696 -376 1736 -350
rect 1762 -376 1802 -350
rect 1828 -376 1868 -350
rect 1894 -376 1934 -350
rect 1960 -376 2000 -350
rect 2026 -376 2066 -350
rect 2092 -376 2132 -350
rect 2158 -376 2198 -350
rect 2224 -376 2264 -350
rect 2290 -376 2330 -350
rect 2356 -376 2396 -350
rect 2422 -376 2462 -350
rect 2488 -376 2528 -350
rect 2554 -376 2594 -350
rect 2620 -376 2626 -350
rect -2626 -382 2626 -376
<< via1 >>
rect -2620 350 -2594 376
rect -2554 350 -2528 376
rect -2488 350 -2462 376
rect -2422 350 -2396 376
rect -2356 350 -2330 376
rect -2290 350 -2264 376
rect -2224 350 -2198 376
rect -2158 350 -2132 376
rect -2092 350 -2066 376
rect -2026 350 -2000 376
rect -1960 350 -1934 376
rect -1894 350 -1868 376
rect -1828 350 -1802 376
rect -1762 350 -1736 376
rect -1696 350 -1670 376
rect -1630 350 -1604 376
rect -1564 350 -1538 376
rect -1498 350 -1472 376
rect -1432 350 -1406 376
rect -1366 350 -1340 376
rect -1300 350 -1274 376
rect -1234 350 -1208 376
rect -1168 350 -1142 376
rect -1102 350 -1076 376
rect -1036 350 -1010 376
rect -970 350 -944 376
rect -904 350 -878 376
rect -838 350 -812 376
rect -772 350 -746 376
rect -706 350 -680 376
rect -640 350 -614 376
rect -574 350 -548 376
rect -508 350 -482 376
rect -442 350 -416 376
rect -376 350 -350 376
rect -310 350 -284 376
rect -244 350 -218 376
rect -178 350 -152 376
rect -112 350 -86 376
rect -46 350 -20 376
rect 20 350 46 376
rect 86 350 112 376
rect 152 350 178 376
rect 218 350 244 376
rect 284 350 310 376
rect 350 350 376 376
rect 416 350 442 376
rect 482 350 508 376
rect 548 350 574 376
rect 614 350 640 376
rect 680 350 706 376
rect 746 350 772 376
rect 812 350 838 376
rect 878 350 904 376
rect 944 350 970 376
rect 1010 350 1036 376
rect 1076 350 1102 376
rect 1142 350 1168 376
rect 1208 350 1234 376
rect 1274 350 1300 376
rect 1340 350 1366 376
rect 1406 350 1432 376
rect 1472 350 1498 376
rect 1538 350 1564 376
rect 1604 350 1630 376
rect 1670 350 1696 376
rect 1736 350 1762 376
rect 1802 350 1828 376
rect 1868 350 1894 376
rect 1934 350 1960 376
rect 2000 350 2026 376
rect 2066 350 2092 376
rect 2132 350 2158 376
rect 2198 350 2224 376
rect 2264 350 2290 376
rect 2330 350 2356 376
rect 2396 350 2422 376
rect 2462 350 2488 376
rect 2528 350 2554 376
rect 2594 350 2620 376
rect -2620 284 -2594 310
rect -2554 284 -2528 310
rect -2488 284 -2462 310
rect -2422 284 -2396 310
rect -2356 284 -2330 310
rect -2290 284 -2264 310
rect -2224 284 -2198 310
rect -2158 284 -2132 310
rect -2092 284 -2066 310
rect -2026 284 -2000 310
rect -1960 284 -1934 310
rect -1894 284 -1868 310
rect -1828 284 -1802 310
rect -1762 284 -1736 310
rect -1696 284 -1670 310
rect -1630 284 -1604 310
rect -1564 284 -1538 310
rect -1498 284 -1472 310
rect -1432 284 -1406 310
rect -1366 284 -1340 310
rect -1300 284 -1274 310
rect -1234 284 -1208 310
rect -1168 284 -1142 310
rect -1102 284 -1076 310
rect -1036 284 -1010 310
rect -970 284 -944 310
rect -904 284 -878 310
rect -838 284 -812 310
rect -772 284 -746 310
rect -706 284 -680 310
rect -640 284 -614 310
rect -574 284 -548 310
rect -508 284 -482 310
rect -442 284 -416 310
rect -376 284 -350 310
rect -310 284 -284 310
rect -244 284 -218 310
rect -178 284 -152 310
rect -112 284 -86 310
rect -46 284 -20 310
rect 20 284 46 310
rect 86 284 112 310
rect 152 284 178 310
rect 218 284 244 310
rect 284 284 310 310
rect 350 284 376 310
rect 416 284 442 310
rect 482 284 508 310
rect 548 284 574 310
rect 614 284 640 310
rect 680 284 706 310
rect 746 284 772 310
rect 812 284 838 310
rect 878 284 904 310
rect 944 284 970 310
rect 1010 284 1036 310
rect 1076 284 1102 310
rect 1142 284 1168 310
rect 1208 284 1234 310
rect 1274 284 1300 310
rect 1340 284 1366 310
rect 1406 284 1432 310
rect 1472 284 1498 310
rect 1538 284 1564 310
rect 1604 284 1630 310
rect 1670 284 1696 310
rect 1736 284 1762 310
rect 1802 284 1828 310
rect 1868 284 1894 310
rect 1934 284 1960 310
rect 2000 284 2026 310
rect 2066 284 2092 310
rect 2132 284 2158 310
rect 2198 284 2224 310
rect 2264 284 2290 310
rect 2330 284 2356 310
rect 2396 284 2422 310
rect 2462 284 2488 310
rect 2528 284 2554 310
rect 2594 284 2620 310
rect -2620 218 -2594 244
rect -2554 218 -2528 244
rect -2488 218 -2462 244
rect -2422 218 -2396 244
rect -2356 218 -2330 244
rect -2290 218 -2264 244
rect -2224 218 -2198 244
rect -2158 218 -2132 244
rect -2092 218 -2066 244
rect -2026 218 -2000 244
rect -1960 218 -1934 244
rect -1894 218 -1868 244
rect -1828 218 -1802 244
rect -1762 218 -1736 244
rect -1696 218 -1670 244
rect -1630 218 -1604 244
rect -1564 218 -1538 244
rect -1498 218 -1472 244
rect -1432 218 -1406 244
rect -1366 218 -1340 244
rect -1300 218 -1274 244
rect -1234 218 -1208 244
rect -1168 218 -1142 244
rect -1102 218 -1076 244
rect -1036 218 -1010 244
rect -970 218 -944 244
rect -904 218 -878 244
rect -838 218 -812 244
rect -772 218 -746 244
rect -706 218 -680 244
rect -640 218 -614 244
rect -574 218 -548 244
rect -508 218 -482 244
rect -442 218 -416 244
rect -376 218 -350 244
rect -310 218 -284 244
rect -244 218 -218 244
rect -178 218 -152 244
rect -112 218 -86 244
rect -46 218 -20 244
rect 20 218 46 244
rect 86 218 112 244
rect 152 218 178 244
rect 218 218 244 244
rect 284 218 310 244
rect 350 218 376 244
rect 416 218 442 244
rect 482 218 508 244
rect 548 218 574 244
rect 614 218 640 244
rect 680 218 706 244
rect 746 218 772 244
rect 812 218 838 244
rect 878 218 904 244
rect 944 218 970 244
rect 1010 218 1036 244
rect 1076 218 1102 244
rect 1142 218 1168 244
rect 1208 218 1234 244
rect 1274 218 1300 244
rect 1340 218 1366 244
rect 1406 218 1432 244
rect 1472 218 1498 244
rect 1538 218 1564 244
rect 1604 218 1630 244
rect 1670 218 1696 244
rect 1736 218 1762 244
rect 1802 218 1828 244
rect 1868 218 1894 244
rect 1934 218 1960 244
rect 2000 218 2026 244
rect 2066 218 2092 244
rect 2132 218 2158 244
rect 2198 218 2224 244
rect 2264 218 2290 244
rect 2330 218 2356 244
rect 2396 218 2422 244
rect 2462 218 2488 244
rect 2528 218 2554 244
rect 2594 218 2620 244
rect -2620 152 -2594 178
rect -2554 152 -2528 178
rect -2488 152 -2462 178
rect -2422 152 -2396 178
rect -2356 152 -2330 178
rect -2290 152 -2264 178
rect -2224 152 -2198 178
rect -2158 152 -2132 178
rect -2092 152 -2066 178
rect -2026 152 -2000 178
rect -1960 152 -1934 178
rect -1894 152 -1868 178
rect -1828 152 -1802 178
rect -1762 152 -1736 178
rect -1696 152 -1670 178
rect -1630 152 -1604 178
rect -1564 152 -1538 178
rect -1498 152 -1472 178
rect -1432 152 -1406 178
rect -1366 152 -1340 178
rect -1300 152 -1274 178
rect -1234 152 -1208 178
rect -1168 152 -1142 178
rect -1102 152 -1076 178
rect -1036 152 -1010 178
rect -970 152 -944 178
rect -904 152 -878 178
rect -838 152 -812 178
rect -772 152 -746 178
rect -706 152 -680 178
rect -640 152 -614 178
rect -574 152 -548 178
rect -508 152 -482 178
rect -442 152 -416 178
rect -376 152 -350 178
rect -310 152 -284 178
rect -244 152 -218 178
rect -178 152 -152 178
rect -112 152 -86 178
rect -46 152 -20 178
rect 20 152 46 178
rect 86 152 112 178
rect 152 152 178 178
rect 218 152 244 178
rect 284 152 310 178
rect 350 152 376 178
rect 416 152 442 178
rect 482 152 508 178
rect 548 152 574 178
rect 614 152 640 178
rect 680 152 706 178
rect 746 152 772 178
rect 812 152 838 178
rect 878 152 904 178
rect 944 152 970 178
rect 1010 152 1036 178
rect 1076 152 1102 178
rect 1142 152 1168 178
rect 1208 152 1234 178
rect 1274 152 1300 178
rect 1340 152 1366 178
rect 1406 152 1432 178
rect 1472 152 1498 178
rect 1538 152 1564 178
rect 1604 152 1630 178
rect 1670 152 1696 178
rect 1736 152 1762 178
rect 1802 152 1828 178
rect 1868 152 1894 178
rect 1934 152 1960 178
rect 2000 152 2026 178
rect 2066 152 2092 178
rect 2132 152 2158 178
rect 2198 152 2224 178
rect 2264 152 2290 178
rect 2330 152 2356 178
rect 2396 152 2422 178
rect 2462 152 2488 178
rect 2528 152 2554 178
rect 2594 152 2620 178
rect -2620 86 -2594 112
rect -2554 86 -2528 112
rect -2488 86 -2462 112
rect -2422 86 -2396 112
rect -2356 86 -2330 112
rect -2290 86 -2264 112
rect -2224 86 -2198 112
rect -2158 86 -2132 112
rect -2092 86 -2066 112
rect -2026 86 -2000 112
rect -1960 86 -1934 112
rect -1894 86 -1868 112
rect -1828 86 -1802 112
rect -1762 86 -1736 112
rect -1696 86 -1670 112
rect -1630 86 -1604 112
rect -1564 86 -1538 112
rect -1498 86 -1472 112
rect -1432 86 -1406 112
rect -1366 86 -1340 112
rect -1300 86 -1274 112
rect -1234 86 -1208 112
rect -1168 86 -1142 112
rect -1102 86 -1076 112
rect -1036 86 -1010 112
rect -970 86 -944 112
rect -904 86 -878 112
rect -838 86 -812 112
rect -772 86 -746 112
rect -706 86 -680 112
rect -640 86 -614 112
rect -574 86 -548 112
rect -508 86 -482 112
rect -442 86 -416 112
rect -376 86 -350 112
rect -310 86 -284 112
rect -244 86 -218 112
rect -178 86 -152 112
rect -112 86 -86 112
rect -46 86 -20 112
rect 20 86 46 112
rect 86 86 112 112
rect 152 86 178 112
rect 218 86 244 112
rect 284 86 310 112
rect 350 86 376 112
rect 416 86 442 112
rect 482 86 508 112
rect 548 86 574 112
rect 614 86 640 112
rect 680 86 706 112
rect 746 86 772 112
rect 812 86 838 112
rect 878 86 904 112
rect 944 86 970 112
rect 1010 86 1036 112
rect 1076 86 1102 112
rect 1142 86 1168 112
rect 1208 86 1234 112
rect 1274 86 1300 112
rect 1340 86 1366 112
rect 1406 86 1432 112
rect 1472 86 1498 112
rect 1538 86 1564 112
rect 1604 86 1630 112
rect 1670 86 1696 112
rect 1736 86 1762 112
rect 1802 86 1828 112
rect 1868 86 1894 112
rect 1934 86 1960 112
rect 2000 86 2026 112
rect 2066 86 2092 112
rect 2132 86 2158 112
rect 2198 86 2224 112
rect 2264 86 2290 112
rect 2330 86 2356 112
rect 2396 86 2422 112
rect 2462 86 2488 112
rect 2528 86 2554 112
rect 2594 86 2620 112
rect -2620 20 -2594 46
rect -2554 20 -2528 46
rect -2488 20 -2462 46
rect -2422 20 -2396 46
rect -2356 20 -2330 46
rect -2290 20 -2264 46
rect -2224 20 -2198 46
rect -2158 20 -2132 46
rect -2092 20 -2066 46
rect -2026 20 -2000 46
rect -1960 20 -1934 46
rect -1894 20 -1868 46
rect -1828 20 -1802 46
rect -1762 20 -1736 46
rect -1696 20 -1670 46
rect -1630 20 -1604 46
rect -1564 20 -1538 46
rect -1498 20 -1472 46
rect -1432 20 -1406 46
rect -1366 20 -1340 46
rect -1300 20 -1274 46
rect -1234 20 -1208 46
rect -1168 20 -1142 46
rect -1102 20 -1076 46
rect -1036 20 -1010 46
rect -970 20 -944 46
rect -904 20 -878 46
rect -838 20 -812 46
rect -772 20 -746 46
rect -706 20 -680 46
rect -640 20 -614 46
rect -574 20 -548 46
rect -508 20 -482 46
rect -442 20 -416 46
rect -376 20 -350 46
rect -310 20 -284 46
rect -244 20 -218 46
rect -178 20 -152 46
rect -112 20 -86 46
rect -46 20 -20 46
rect 20 20 46 46
rect 86 20 112 46
rect 152 20 178 46
rect 218 20 244 46
rect 284 20 310 46
rect 350 20 376 46
rect 416 20 442 46
rect 482 20 508 46
rect 548 20 574 46
rect 614 20 640 46
rect 680 20 706 46
rect 746 20 772 46
rect 812 20 838 46
rect 878 20 904 46
rect 944 20 970 46
rect 1010 20 1036 46
rect 1076 20 1102 46
rect 1142 20 1168 46
rect 1208 20 1234 46
rect 1274 20 1300 46
rect 1340 20 1366 46
rect 1406 20 1432 46
rect 1472 20 1498 46
rect 1538 20 1564 46
rect 1604 20 1630 46
rect 1670 20 1696 46
rect 1736 20 1762 46
rect 1802 20 1828 46
rect 1868 20 1894 46
rect 1934 20 1960 46
rect 2000 20 2026 46
rect 2066 20 2092 46
rect 2132 20 2158 46
rect 2198 20 2224 46
rect 2264 20 2290 46
rect 2330 20 2356 46
rect 2396 20 2422 46
rect 2462 20 2488 46
rect 2528 20 2554 46
rect 2594 20 2620 46
rect -2620 -46 -2594 -20
rect -2554 -46 -2528 -20
rect -2488 -46 -2462 -20
rect -2422 -46 -2396 -20
rect -2356 -46 -2330 -20
rect -2290 -46 -2264 -20
rect -2224 -46 -2198 -20
rect -2158 -46 -2132 -20
rect -2092 -46 -2066 -20
rect -2026 -46 -2000 -20
rect -1960 -46 -1934 -20
rect -1894 -46 -1868 -20
rect -1828 -46 -1802 -20
rect -1762 -46 -1736 -20
rect -1696 -46 -1670 -20
rect -1630 -46 -1604 -20
rect -1564 -46 -1538 -20
rect -1498 -46 -1472 -20
rect -1432 -46 -1406 -20
rect -1366 -46 -1340 -20
rect -1300 -46 -1274 -20
rect -1234 -46 -1208 -20
rect -1168 -46 -1142 -20
rect -1102 -46 -1076 -20
rect -1036 -46 -1010 -20
rect -970 -46 -944 -20
rect -904 -46 -878 -20
rect -838 -46 -812 -20
rect -772 -46 -746 -20
rect -706 -46 -680 -20
rect -640 -46 -614 -20
rect -574 -46 -548 -20
rect -508 -46 -482 -20
rect -442 -46 -416 -20
rect -376 -46 -350 -20
rect -310 -46 -284 -20
rect -244 -46 -218 -20
rect -178 -46 -152 -20
rect -112 -46 -86 -20
rect -46 -46 -20 -20
rect 20 -46 46 -20
rect 86 -46 112 -20
rect 152 -46 178 -20
rect 218 -46 244 -20
rect 284 -46 310 -20
rect 350 -46 376 -20
rect 416 -46 442 -20
rect 482 -46 508 -20
rect 548 -46 574 -20
rect 614 -46 640 -20
rect 680 -46 706 -20
rect 746 -46 772 -20
rect 812 -46 838 -20
rect 878 -46 904 -20
rect 944 -46 970 -20
rect 1010 -46 1036 -20
rect 1076 -46 1102 -20
rect 1142 -46 1168 -20
rect 1208 -46 1234 -20
rect 1274 -46 1300 -20
rect 1340 -46 1366 -20
rect 1406 -46 1432 -20
rect 1472 -46 1498 -20
rect 1538 -46 1564 -20
rect 1604 -46 1630 -20
rect 1670 -46 1696 -20
rect 1736 -46 1762 -20
rect 1802 -46 1828 -20
rect 1868 -46 1894 -20
rect 1934 -46 1960 -20
rect 2000 -46 2026 -20
rect 2066 -46 2092 -20
rect 2132 -46 2158 -20
rect 2198 -46 2224 -20
rect 2264 -46 2290 -20
rect 2330 -46 2356 -20
rect 2396 -46 2422 -20
rect 2462 -46 2488 -20
rect 2528 -46 2554 -20
rect 2594 -46 2620 -20
rect -2620 -112 -2594 -86
rect -2554 -112 -2528 -86
rect -2488 -112 -2462 -86
rect -2422 -112 -2396 -86
rect -2356 -112 -2330 -86
rect -2290 -112 -2264 -86
rect -2224 -112 -2198 -86
rect -2158 -112 -2132 -86
rect -2092 -112 -2066 -86
rect -2026 -112 -2000 -86
rect -1960 -112 -1934 -86
rect -1894 -112 -1868 -86
rect -1828 -112 -1802 -86
rect -1762 -112 -1736 -86
rect -1696 -112 -1670 -86
rect -1630 -112 -1604 -86
rect -1564 -112 -1538 -86
rect -1498 -112 -1472 -86
rect -1432 -112 -1406 -86
rect -1366 -112 -1340 -86
rect -1300 -112 -1274 -86
rect -1234 -112 -1208 -86
rect -1168 -112 -1142 -86
rect -1102 -112 -1076 -86
rect -1036 -112 -1010 -86
rect -970 -112 -944 -86
rect -904 -112 -878 -86
rect -838 -112 -812 -86
rect -772 -112 -746 -86
rect -706 -112 -680 -86
rect -640 -112 -614 -86
rect -574 -112 -548 -86
rect -508 -112 -482 -86
rect -442 -112 -416 -86
rect -376 -112 -350 -86
rect -310 -112 -284 -86
rect -244 -112 -218 -86
rect -178 -112 -152 -86
rect -112 -112 -86 -86
rect -46 -112 -20 -86
rect 20 -112 46 -86
rect 86 -112 112 -86
rect 152 -112 178 -86
rect 218 -112 244 -86
rect 284 -112 310 -86
rect 350 -112 376 -86
rect 416 -112 442 -86
rect 482 -112 508 -86
rect 548 -112 574 -86
rect 614 -112 640 -86
rect 680 -112 706 -86
rect 746 -112 772 -86
rect 812 -112 838 -86
rect 878 -112 904 -86
rect 944 -112 970 -86
rect 1010 -112 1036 -86
rect 1076 -112 1102 -86
rect 1142 -112 1168 -86
rect 1208 -112 1234 -86
rect 1274 -112 1300 -86
rect 1340 -112 1366 -86
rect 1406 -112 1432 -86
rect 1472 -112 1498 -86
rect 1538 -112 1564 -86
rect 1604 -112 1630 -86
rect 1670 -112 1696 -86
rect 1736 -112 1762 -86
rect 1802 -112 1828 -86
rect 1868 -112 1894 -86
rect 1934 -112 1960 -86
rect 2000 -112 2026 -86
rect 2066 -112 2092 -86
rect 2132 -112 2158 -86
rect 2198 -112 2224 -86
rect 2264 -112 2290 -86
rect 2330 -112 2356 -86
rect 2396 -112 2422 -86
rect 2462 -112 2488 -86
rect 2528 -112 2554 -86
rect 2594 -112 2620 -86
rect -2620 -178 -2594 -152
rect -2554 -178 -2528 -152
rect -2488 -178 -2462 -152
rect -2422 -178 -2396 -152
rect -2356 -178 -2330 -152
rect -2290 -178 -2264 -152
rect -2224 -178 -2198 -152
rect -2158 -178 -2132 -152
rect -2092 -178 -2066 -152
rect -2026 -178 -2000 -152
rect -1960 -178 -1934 -152
rect -1894 -178 -1868 -152
rect -1828 -178 -1802 -152
rect -1762 -178 -1736 -152
rect -1696 -178 -1670 -152
rect -1630 -178 -1604 -152
rect -1564 -178 -1538 -152
rect -1498 -178 -1472 -152
rect -1432 -178 -1406 -152
rect -1366 -178 -1340 -152
rect -1300 -178 -1274 -152
rect -1234 -178 -1208 -152
rect -1168 -178 -1142 -152
rect -1102 -178 -1076 -152
rect -1036 -178 -1010 -152
rect -970 -178 -944 -152
rect -904 -178 -878 -152
rect -838 -178 -812 -152
rect -772 -178 -746 -152
rect -706 -178 -680 -152
rect -640 -178 -614 -152
rect -574 -178 -548 -152
rect -508 -178 -482 -152
rect -442 -178 -416 -152
rect -376 -178 -350 -152
rect -310 -178 -284 -152
rect -244 -178 -218 -152
rect -178 -178 -152 -152
rect -112 -178 -86 -152
rect -46 -178 -20 -152
rect 20 -178 46 -152
rect 86 -178 112 -152
rect 152 -178 178 -152
rect 218 -178 244 -152
rect 284 -178 310 -152
rect 350 -178 376 -152
rect 416 -178 442 -152
rect 482 -178 508 -152
rect 548 -178 574 -152
rect 614 -178 640 -152
rect 680 -178 706 -152
rect 746 -178 772 -152
rect 812 -178 838 -152
rect 878 -178 904 -152
rect 944 -178 970 -152
rect 1010 -178 1036 -152
rect 1076 -178 1102 -152
rect 1142 -178 1168 -152
rect 1208 -178 1234 -152
rect 1274 -178 1300 -152
rect 1340 -178 1366 -152
rect 1406 -178 1432 -152
rect 1472 -178 1498 -152
rect 1538 -178 1564 -152
rect 1604 -178 1630 -152
rect 1670 -178 1696 -152
rect 1736 -178 1762 -152
rect 1802 -178 1828 -152
rect 1868 -178 1894 -152
rect 1934 -178 1960 -152
rect 2000 -178 2026 -152
rect 2066 -178 2092 -152
rect 2132 -178 2158 -152
rect 2198 -178 2224 -152
rect 2264 -178 2290 -152
rect 2330 -178 2356 -152
rect 2396 -178 2422 -152
rect 2462 -178 2488 -152
rect 2528 -178 2554 -152
rect 2594 -178 2620 -152
rect -2620 -244 -2594 -218
rect -2554 -244 -2528 -218
rect -2488 -244 -2462 -218
rect -2422 -244 -2396 -218
rect -2356 -244 -2330 -218
rect -2290 -244 -2264 -218
rect -2224 -244 -2198 -218
rect -2158 -244 -2132 -218
rect -2092 -244 -2066 -218
rect -2026 -244 -2000 -218
rect -1960 -244 -1934 -218
rect -1894 -244 -1868 -218
rect -1828 -244 -1802 -218
rect -1762 -244 -1736 -218
rect -1696 -244 -1670 -218
rect -1630 -244 -1604 -218
rect -1564 -244 -1538 -218
rect -1498 -244 -1472 -218
rect -1432 -244 -1406 -218
rect -1366 -244 -1340 -218
rect -1300 -244 -1274 -218
rect -1234 -244 -1208 -218
rect -1168 -244 -1142 -218
rect -1102 -244 -1076 -218
rect -1036 -244 -1010 -218
rect -970 -244 -944 -218
rect -904 -244 -878 -218
rect -838 -244 -812 -218
rect -772 -244 -746 -218
rect -706 -244 -680 -218
rect -640 -244 -614 -218
rect -574 -244 -548 -218
rect -508 -244 -482 -218
rect -442 -244 -416 -218
rect -376 -244 -350 -218
rect -310 -244 -284 -218
rect -244 -244 -218 -218
rect -178 -244 -152 -218
rect -112 -244 -86 -218
rect -46 -244 -20 -218
rect 20 -244 46 -218
rect 86 -244 112 -218
rect 152 -244 178 -218
rect 218 -244 244 -218
rect 284 -244 310 -218
rect 350 -244 376 -218
rect 416 -244 442 -218
rect 482 -244 508 -218
rect 548 -244 574 -218
rect 614 -244 640 -218
rect 680 -244 706 -218
rect 746 -244 772 -218
rect 812 -244 838 -218
rect 878 -244 904 -218
rect 944 -244 970 -218
rect 1010 -244 1036 -218
rect 1076 -244 1102 -218
rect 1142 -244 1168 -218
rect 1208 -244 1234 -218
rect 1274 -244 1300 -218
rect 1340 -244 1366 -218
rect 1406 -244 1432 -218
rect 1472 -244 1498 -218
rect 1538 -244 1564 -218
rect 1604 -244 1630 -218
rect 1670 -244 1696 -218
rect 1736 -244 1762 -218
rect 1802 -244 1828 -218
rect 1868 -244 1894 -218
rect 1934 -244 1960 -218
rect 2000 -244 2026 -218
rect 2066 -244 2092 -218
rect 2132 -244 2158 -218
rect 2198 -244 2224 -218
rect 2264 -244 2290 -218
rect 2330 -244 2356 -218
rect 2396 -244 2422 -218
rect 2462 -244 2488 -218
rect 2528 -244 2554 -218
rect 2594 -244 2620 -218
rect -2620 -310 -2594 -284
rect -2554 -310 -2528 -284
rect -2488 -310 -2462 -284
rect -2422 -310 -2396 -284
rect -2356 -310 -2330 -284
rect -2290 -310 -2264 -284
rect -2224 -310 -2198 -284
rect -2158 -310 -2132 -284
rect -2092 -310 -2066 -284
rect -2026 -310 -2000 -284
rect -1960 -310 -1934 -284
rect -1894 -310 -1868 -284
rect -1828 -310 -1802 -284
rect -1762 -310 -1736 -284
rect -1696 -310 -1670 -284
rect -1630 -310 -1604 -284
rect -1564 -310 -1538 -284
rect -1498 -310 -1472 -284
rect -1432 -310 -1406 -284
rect -1366 -310 -1340 -284
rect -1300 -310 -1274 -284
rect -1234 -310 -1208 -284
rect -1168 -310 -1142 -284
rect -1102 -310 -1076 -284
rect -1036 -310 -1010 -284
rect -970 -310 -944 -284
rect -904 -310 -878 -284
rect -838 -310 -812 -284
rect -772 -310 -746 -284
rect -706 -310 -680 -284
rect -640 -310 -614 -284
rect -574 -310 -548 -284
rect -508 -310 -482 -284
rect -442 -310 -416 -284
rect -376 -310 -350 -284
rect -310 -310 -284 -284
rect -244 -310 -218 -284
rect -178 -310 -152 -284
rect -112 -310 -86 -284
rect -46 -310 -20 -284
rect 20 -310 46 -284
rect 86 -310 112 -284
rect 152 -310 178 -284
rect 218 -310 244 -284
rect 284 -310 310 -284
rect 350 -310 376 -284
rect 416 -310 442 -284
rect 482 -310 508 -284
rect 548 -310 574 -284
rect 614 -310 640 -284
rect 680 -310 706 -284
rect 746 -310 772 -284
rect 812 -310 838 -284
rect 878 -310 904 -284
rect 944 -310 970 -284
rect 1010 -310 1036 -284
rect 1076 -310 1102 -284
rect 1142 -310 1168 -284
rect 1208 -310 1234 -284
rect 1274 -310 1300 -284
rect 1340 -310 1366 -284
rect 1406 -310 1432 -284
rect 1472 -310 1498 -284
rect 1538 -310 1564 -284
rect 1604 -310 1630 -284
rect 1670 -310 1696 -284
rect 1736 -310 1762 -284
rect 1802 -310 1828 -284
rect 1868 -310 1894 -284
rect 1934 -310 1960 -284
rect 2000 -310 2026 -284
rect 2066 -310 2092 -284
rect 2132 -310 2158 -284
rect 2198 -310 2224 -284
rect 2264 -310 2290 -284
rect 2330 -310 2356 -284
rect 2396 -310 2422 -284
rect 2462 -310 2488 -284
rect 2528 -310 2554 -284
rect 2594 -310 2620 -284
rect -2620 -376 -2594 -350
rect -2554 -376 -2528 -350
rect -2488 -376 -2462 -350
rect -2422 -376 -2396 -350
rect -2356 -376 -2330 -350
rect -2290 -376 -2264 -350
rect -2224 -376 -2198 -350
rect -2158 -376 -2132 -350
rect -2092 -376 -2066 -350
rect -2026 -376 -2000 -350
rect -1960 -376 -1934 -350
rect -1894 -376 -1868 -350
rect -1828 -376 -1802 -350
rect -1762 -376 -1736 -350
rect -1696 -376 -1670 -350
rect -1630 -376 -1604 -350
rect -1564 -376 -1538 -350
rect -1498 -376 -1472 -350
rect -1432 -376 -1406 -350
rect -1366 -376 -1340 -350
rect -1300 -376 -1274 -350
rect -1234 -376 -1208 -350
rect -1168 -376 -1142 -350
rect -1102 -376 -1076 -350
rect -1036 -376 -1010 -350
rect -970 -376 -944 -350
rect -904 -376 -878 -350
rect -838 -376 -812 -350
rect -772 -376 -746 -350
rect -706 -376 -680 -350
rect -640 -376 -614 -350
rect -574 -376 -548 -350
rect -508 -376 -482 -350
rect -442 -376 -416 -350
rect -376 -376 -350 -350
rect -310 -376 -284 -350
rect -244 -376 -218 -350
rect -178 -376 -152 -350
rect -112 -376 -86 -350
rect -46 -376 -20 -350
rect 20 -376 46 -350
rect 86 -376 112 -350
rect 152 -376 178 -350
rect 218 -376 244 -350
rect 284 -376 310 -350
rect 350 -376 376 -350
rect 416 -376 442 -350
rect 482 -376 508 -350
rect 548 -376 574 -350
rect 614 -376 640 -350
rect 680 -376 706 -350
rect 746 -376 772 -350
rect 812 -376 838 -350
rect 878 -376 904 -350
rect 944 -376 970 -350
rect 1010 -376 1036 -350
rect 1076 -376 1102 -350
rect 1142 -376 1168 -350
rect 1208 -376 1234 -350
rect 1274 -376 1300 -350
rect 1340 -376 1366 -350
rect 1406 -376 1432 -350
rect 1472 -376 1498 -350
rect 1538 -376 1564 -350
rect 1604 -376 1630 -350
rect 1670 -376 1696 -350
rect 1736 -376 1762 -350
rect 1802 -376 1828 -350
rect 1868 -376 1894 -350
rect 1934 -376 1960 -350
rect 2000 -376 2026 -350
rect 2066 -376 2092 -350
rect 2132 -376 2158 -350
rect 2198 -376 2224 -350
rect 2264 -376 2290 -350
rect 2330 -376 2356 -350
rect 2396 -376 2422 -350
rect 2462 -376 2488 -350
rect 2528 -376 2554 -350
rect 2594 -376 2620 -350
<< metal2 >>
rect -2626 376 2626 382
rect -2626 350 -2620 376
rect -2594 350 -2554 376
rect -2528 350 -2488 376
rect -2462 350 -2422 376
rect -2396 350 -2356 376
rect -2330 350 -2290 376
rect -2264 350 -2224 376
rect -2198 350 -2158 376
rect -2132 350 -2092 376
rect -2066 350 -2026 376
rect -2000 350 -1960 376
rect -1934 350 -1894 376
rect -1868 350 -1828 376
rect -1802 350 -1762 376
rect -1736 350 -1696 376
rect -1670 350 -1630 376
rect -1604 350 -1564 376
rect -1538 350 -1498 376
rect -1472 350 -1432 376
rect -1406 350 -1366 376
rect -1340 350 -1300 376
rect -1274 350 -1234 376
rect -1208 350 -1168 376
rect -1142 350 -1102 376
rect -1076 350 -1036 376
rect -1010 350 -970 376
rect -944 350 -904 376
rect -878 350 -838 376
rect -812 350 -772 376
rect -746 350 -706 376
rect -680 350 -640 376
rect -614 350 -574 376
rect -548 350 -508 376
rect -482 350 -442 376
rect -416 350 -376 376
rect -350 350 -310 376
rect -284 350 -244 376
rect -218 350 -178 376
rect -152 350 -112 376
rect -86 350 -46 376
rect -20 350 20 376
rect 46 350 86 376
rect 112 350 152 376
rect 178 350 218 376
rect 244 350 284 376
rect 310 350 350 376
rect 376 350 416 376
rect 442 350 482 376
rect 508 350 548 376
rect 574 350 614 376
rect 640 350 680 376
rect 706 350 746 376
rect 772 350 812 376
rect 838 350 878 376
rect 904 350 944 376
rect 970 350 1010 376
rect 1036 350 1076 376
rect 1102 350 1142 376
rect 1168 350 1208 376
rect 1234 350 1274 376
rect 1300 350 1340 376
rect 1366 350 1406 376
rect 1432 350 1472 376
rect 1498 350 1538 376
rect 1564 350 1604 376
rect 1630 350 1670 376
rect 1696 350 1736 376
rect 1762 350 1802 376
rect 1828 350 1868 376
rect 1894 350 1934 376
rect 1960 350 2000 376
rect 2026 350 2066 376
rect 2092 350 2132 376
rect 2158 350 2198 376
rect 2224 350 2264 376
rect 2290 350 2330 376
rect 2356 350 2396 376
rect 2422 350 2462 376
rect 2488 350 2528 376
rect 2554 350 2594 376
rect 2620 350 2626 376
rect -2626 310 2626 350
rect -2626 284 -2620 310
rect -2594 284 -2554 310
rect -2528 284 -2488 310
rect -2462 284 -2422 310
rect -2396 284 -2356 310
rect -2330 284 -2290 310
rect -2264 284 -2224 310
rect -2198 284 -2158 310
rect -2132 284 -2092 310
rect -2066 284 -2026 310
rect -2000 284 -1960 310
rect -1934 284 -1894 310
rect -1868 284 -1828 310
rect -1802 284 -1762 310
rect -1736 284 -1696 310
rect -1670 284 -1630 310
rect -1604 284 -1564 310
rect -1538 284 -1498 310
rect -1472 284 -1432 310
rect -1406 284 -1366 310
rect -1340 284 -1300 310
rect -1274 284 -1234 310
rect -1208 284 -1168 310
rect -1142 284 -1102 310
rect -1076 284 -1036 310
rect -1010 284 -970 310
rect -944 284 -904 310
rect -878 284 -838 310
rect -812 284 -772 310
rect -746 284 -706 310
rect -680 284 -640 310
rect -614 284 -574 310
rect -548 284 -508 310
rect -482 284 -442 310
rect -416 284 -376 310
rect -350 284 -310 310
rect -284 284 -244 310
rect -218 284 -178 310
rect -152 284 -112 310
rect -86 284 -46 310
rect -20 284 20 310
rect 46 284 86 310
rect 112 284 152 310
rect 178 284 218 310
rect 244 284 284 310
rect 310 284 350 310
rect 376 284 416 310
rect 442 284 482 310
rect 508 284 548 310
rect 574 284 614 310
rect 640 284 680 310
rect 706 284 746 310
rect 772 284 812 310
rect 838 284 878 310
rect 904 284 944 310
rect 970 284 1010 310
rect 1036 284 1076 310
rect 1102 284 1142 310
rect 1168 284 1208 310
rect 1234 284 1274 310
rect 1300 284 1340 310
rect 1366 284 1406 310
rect 1432 284 1472 310
rect 1498 284 1538 310
rect 1564 284 1604 310
rect 1630 284 1670 310
rect 1696 284 1736 310
rect 1762 284 1802 310
rect 1828 284 1868 310
rect 1894 284 1934 310
rect 1960 284 2000 310
rect 2026 284 2066 310
rect 2092 284 2132 310
rect 2158 284 2198 310
rect 2224 284 2264 310
rect 2290 284 2330 310
rect 2356 284 2396 310
rect 2422 284 2462 310
rect 2488 284 2528 310
rect 2554 284 2594 310
rect 2620 284 2626 310
rect -2626 244 2626 284
rect -2626 218 -2620 244
rect -2594 218 -2554 244
rect -2528 218 -2488 244
rect -2462 218 -2422 244
rect -2396 218 -2356 244
rect -2330 218 -2290 244
rect -2264 218 -2224 244
rect -2198 218 -2158 244
rect -2132 218 -2092 244
rect -2066 218 -2026 244
rect -2000 218 -1960 244
rect -1934 218 -1894 244
rect -1868 218 -1828 244
rect -1802 218 -1762 244
rect -1736 218 -1696 244
rect -1670 218 -1630 244
rect -1604 218 -1564 244
rect -1538 218 -1498 244
rect -1472 218 -1432 244
rect -1406 218 -1366 244
rect -1340 218 -1300 244
rect -1274 218 -1234 244
rect -1208 218 -1168 244
rect -1142 218 -1102 244
rect -1076 218 -1036 244
rect -1010 218 -970 244
rect -944 218 -904 244
rect -878 218 -838 244
rect -812 218 -772 244
rect -746 218 -706 244
rect -680 218 -640 244
rect -614 218 -574 244
rect -548 218 -508 244
rect -482 218 -442 244
rect -416 218 -376 244
rect -350 218 -310 244
rect -284 218 -244 244
rect -218 218 -178 244
rect -152 218 -112 244
rect -86 218 -46 244
rect -20 218 20 244
rect 46 218 86 244
rect 112 218 152 244
rect 178 218 218 244
rect 244 218 284 244
rect 310 218 350 244
rect 376 218 416 244
rect 442 218 482 244
rect 508 218 548 244
rect 574 218 614 244
rect 640 218 680 244
rect 706 218 746 244
rect 772 218 812 244
rect 838 218 878 244
rect 904 218 944 244
rect 970 218 1010 244
rect 1036 218 1076 244
rect 1102 218 1142 244
rect 1168 218 1208 244
rect 1234 218 1274 244
rect 1300 218 1340 244
rect 1366 218 1406 244
rect 1432 218 1472 244
rect 1498 218 1538 244
rect 1564 218 1604 244
rect 1630 218 1670 244
rect 1696 218 1736 244
rect 1762 218 1802 244
rect 1828 218 1868 244
rect 1894 218 1934 244
rect 1960 218 2000 244
rect 2026 218 2066 244
rect 2092 218 2132 244
rect 2158 218 2198 244
rect 2224 218 2264 244
rect 2290 218 2330 244
rect 2356 218 2396 244
rect 2422 218 2462 244
rect 2488 218 2528 244
rect 2554 218 2594 244
rect 2620 218 2626 244
rect -2626 178 2626 218
rect -2626 152 -2620 178
rect -2594 152 -2554 178
rect -2528 152 -2488 178
rect -2462 152 -2422 178
rect -2396 152 -2356 178
rect -2330 152 -2290 178
rect -2264 152 -2224 178
rect -2198 152 -2158 178
rect -2132 152 -2092 178
rect -2066 152 -2026 178
rect -2000 152 -1960 178
rect -1934 152 -1894 178
rect -1868 152 -1828 178
rect -1802 152 -1762 178
rect -1736 152 -1696 178
rect -1670 152 -1630 178
rect -1604 152 -1564 178
rect -1538 152 -1498 178
rect -1472 152 -1432 178
rect -1406 152 -1366 178
rect -1340 152 -1300 178
rect -1274 152 -1234 178
rect -1208 152 -1168 178
rect -1142 152 -1102 178
rect -1076 152 -1036 178
rect -1010 152 -970 178
rect -944 152 -904 178
rect -878 152 -838 178
rect -812 152 -772 178
rect -746 152 -706 178
rect -680 152 -640 178
rect -614 152 -574 178
rect -548 152 -508 178
rect -482 152 -442 178
rect -416 152 -376 178
rect -350 152 -310 178
rect -284 152 -244 178
rect -218 152 -178 178
rect -152 152 -112 178
rect -86 152 -46 178
rect -20 152 20 178
rect 46 152 86 178
rect 112 152 152 178
rect 178 152 218 178
rect 244 152 284 178
rect 310 152 350 178
rect 376 152 416 178
rect 442 152 482 178
rect 508 152 548 178
rect 574 152 614 178
rect 640 152 680 178
rect 706 152 746 178
rect 772 152 812 178
rect 838 152 878 178
rect 904 152 944 178
rect 970 152 1010 178
rect 1036 152 1076 178
rect 1102 152 1142 178
rect 1168 152 1208 178
rect 1234 152 1274 178
rect 1300 152 1340 178
rect 1366 152 1406 178
rect 1432 152 1472 178
rect 1498 152 1538 178
rect 1564 152 1604 178
rect 1630 152 1670 178
rect 1696 152 1736 178
rect 1762 152 1802 178
rect 1828 152 1868 178
rect 1894 152 1934 178
rect 1960 152 2000 178
rect 2026 152 2066 178
rect 2092 152 2132 178
rect 2158 152 2198 178
rect 2224 152 2264 178
rect 2290 152 2330 178
rect 2356 152 2396 178
rect 2422 152 2462 178
rect 2488 152 2528 178
rect 2554 152 2594 178
rect 2620 152 2626 178
rect -2626 112 2626 152
rect -2626 86 -2620 112
rect -2594 86 -2554 112
rect -2528 86 -2488 112
rect -2462 86 -2422 112
rect -2396 86 -2356 112
rect -2330 86 -2290 112
rect -2264 86 -2224 112
rect -2198 86 -2158 112
rect -2132 86 -2092 112
rect -2066 86 -2026 112
rect -2000 86 -1960 112
rect -1934 86 -1894 112
rect -1868 86 -1828 112
rect -1802 86 -1762 112
rect -1736 86 -1696 112
rect -1670 86 -1630 112
rect -1604 86 -1564 112
rect -1538 86 -1498 112
rect -1472 86 -1432 112
rect -1406 86 -1366 112
rect -1340 86 -1300 112
rect -1274 86 -1234 112
rect -1208 86 -1168 112
rect -1142 86 -1102 112
rect -1076 86 -1036 112
rect -1010 86 -970 112
rect -944 86 -904 112
rect -878 86 -838 112
rect -812 86 -772 112
rect -746 86 -706 112
rect -680 86 -640 112
rect -614 86 -574 112
rect -548 86 -508 112
rect -482 86 -442 112
rect -416 86 -376 112
rect -350 86 -310 112
rect -284 86 -244 112
rect -218 86 -178 112
rect -152 86 -112 112
rect -86 86 -46 112
rect -20 86 20 112
rect 46 86 86 112
rect 112 86 152 112
rect 178 86 218 112
rect 244 86 284 112
rect 310 86 350 112
rect 376 86 416 112
rect 442 86 482 112
rect 508 86 548 112
rect 574 86 614 112
rect 640 86 680 112
rect 706 86 746 112
rect 772 86 812 112
rect 838 86 878 112
rect 904 86 944 112
rect 970 86 1010 112
rect 1036 86 1076 112
rect 1102 86 1142 112
rect 1168 86 1208 112
rect 1234 86 1274 112
rect 1300 86 1340 112
rect 1366 86 1406 112
rect 1432 86 1472 112
rect 1498 86 1538 112
rect 1564 86 1604 112
rect 1630 86 1670 112
rect 1696 86 1736 112
rect 1762 86 1802 112
rect 1828 86 1868 112
rect 1894 86 1934 112
rect 1960 86 2000 112
rect 2026 86 2066 112
rect 2092 86 2132 112
rect 2158 86 2198 112
rect 2224 86 2264 112
rect 2290 86 2330 112
rect 2356 86 2396 112
rect 2422 86 2462 112
rect 2488 86 2528 112
rect 2554 86 2594 112
rect 2620 86 2626 112
rect -2626 46 2626 86
rect -2626 20 -2620 46
rect -2594 20 -2554 46
rect -2528 20 -2488 46
rect -2462 20 -2422 46
rect -2396 20 -2356 46
rect -2330 20 -2290 46
rect -2264 20 -2224 46
rect -2198 20 -2158 46
rect -2132 20 -2092 46
rect -2066 20 -2026 46
rect -2000 20 -1960 46
rect -1934 20 -1894 46
rect -1868 20 -1828 46
rect -1802 20 -1762 46
rect -1736 20 -1696 46
rect -1670 20 -1630 46
rect -1604 20 -1564 46
rect -1538 20 -1498 46
rect -1472 20 -1432 46
rect -1406 20 -1366 46
rect -1340 20 -1300 46
rect -1274 20 -1234 46
rect -1208 20 -1168 46
rect -1142 20 -1102 46
rect -1076 20 -1036 46
rect -1010 20 -970 46
rect -944 20 -904 46
rect -878 20 -838 46
rect -812 20 -772 46
rect -746 20 -706 46
rect -680 20 -640 46
rect -614 20 -574 46
rect -548 20 -508 46
rect -482 20 -442 46
rect -416 20 -376 46
rect -350 20 -310 46
rect -284 20 -244 46
rect -218 20 -178 46
rect -152 20 -112 46
rect -86 20 -46 46
rect -20 20 20 46
rect 46 20 86 46
rect 112 20 152 46
rect 178 20 218 46
rect 244 20 284 46
rect 310 20 350 46
rect 376 20 416 46
rect 442 20 482 46
rect 508 20 548 46
rect 574 20 614 46
rect 640 20 680 46
rect 706 20 746 46
rect 772 20 812 46
rect 838 20 878 46
rect 904 20 944 46
rect 970 20 1010 46
rect 1036 20 1076 46
rect 1102 20 1142 46
rect 1168 20 1208 46
rect 1234 20 1274 46
rect 1300 20 1340 46
rect 1366 20 1406 46
rect 1432 20 1472 46
rect 1498 20 1538 46
rect 1564 20 1604 46
rect 1630 20 1670 46
rect 1696 20 1736 46
rect 1762 20 1802 46
rect 1828 20 1868 46
rect 1894 20 1934 46
rect 1960 20 2000 46
rect 2026 20 2066 46
rect 2092 20 2132 46
rect 2158 20 2198 46
rect 2224 20 2264 46
rect 2290 20 2330 46
rect 2356 20 2396 46
rect 2422 20 2462 46
rect 2488 20 2528 46
rect 2554 20 2594 46
rect 2620 20 2626 46
rect -2626 -20 2626 20
rect -2626 -46 -2620 -20
rect -2594 -46 -2554 -20
rect -2528 -46 -2488 -20
rect -2462 -46 -2422 -20
rect -2396 -46 -2356 -20
rect -2330 -46 -2290 -20
rect -2264 -46 -2224 -20
rect -2198 -46 -2158 -20
rect -2132 -46 -2092 -20
rect -2066 -46 -2026 -20
rect -2000 -46 -1960 -20
rect -1934 -46 -1894 -20
rect -1868 -46 -1828 -20
rect -1802 -46 -1762 -20
rect -1736 -46 -1696 -20
rect -1670 -46 -1630 -20
rect -1604 -46 -1564 -20
rect -1538 -46 -1498 -20
rect -1472 -46 -1432 -20
rect -1406 -46 -1366 -20
rect -1340 -46 -1300 -20
rect -1274 -46 -1234 -20
rect -1208 -46 -1168 -20
rect -1142 -46 -1102 -20
rect -1076 -46 -1036 -20
rect -1010 -46 -970 -20
rect -944 -46 -904 -20
rect -878 -46 -838 -20
rect -812 -46 -772 -20
rect -746 -46 -706 -20
rect -680 -46 -640 -20
rect -614 -46 -574 -20
rect -548 -46 -508 -20
rect -482 -46 -442 -20
rect -416 -46 -376 -20
rect -350 -46 -310 -20
rect -284 -46 -244 -20
rect -218 -46 -178 -20
rect -152 -46 -112 -20
rect -86 -46 -46 -20
rect -20 -46 20 -20
rect 46 -46 86 -20
rect 112 -46 152 -20
rect 178 -46 218 -20
rect 244 -46 284 -20
rect 310 -46 350 -20
rect 376 -46 416 -20
rect 442 -46 482 -20
rect 508 -46 548 -20
rect 574 -46 614 -20
rect 640 -46 680 -20
rect 706 -46 746 -20
rect 772 -46 812 -20
rect 838 -46 878 -20
rect 904 -46 944 -20
rect 970 -46 1010 -20
rect 1036 -46 1076 -20
rect 1102 -46 1142 -20
rect 1168 -46 1208 -20
rect 1234 -46 1274 -20
rect 1300 -46 1340 -20
rect 1366 -46 1406 -20
rect 1432 -46 1472 -20
rect 1498 -46 1538 -20
rect 1564 -46 1604 -20
rect 1630 -46 1670 -20
rect 1696 -46 1736 -20
rect 1762 -46 1802 -20
rect 1828 -46 1868 -20
rect 1894 -46 1934 -20
rect 1960 -46 2000 -20
rect 2026 -46 2066 -20
rect 2092 -46 2132 -20
rect 2158 -46 2198 -20
rect 2224 -46 2264 -20
rect 2290 -46 2330 -20
rect 2356 -46 2396 -20
rect 2422 -46 2462 -20
rect 2488 -46 2528 -20
rect 2554 -46 2594 -20
rect 2620 -46 2626 -20
rect -2626 -86 2626 -46
rect -2626 -112 -2620 -86
rect -2594 -112 -2554 -86
rect -2528 -112 -2488 -86
rect -2462 -112 -2422 -86
rect -2396 -112 -2356 -86
rect -2330 -112 -2290 -86
rect -2264 -112 -2224 -86
rect -2198 -112 -2158 -86
rect -2132 -112 -2092 -86
rect -2066 -112 -2026 -86
rect -2000 -112 -1960 -86
rect -1934 -112 -1894 -86
rect -1868 -112 -1828 -86
rect -1802 -112 -1762 -86
rect -1736 -112 -1696 -86
rect -1670 -112 -1630 -86
rect -1604 -112 -1564 -86
rect -1538 -112 -1498 -86
rect -1472 -112 -1432 -86
rect -1406 -112 -1366 -86
rect -1340 -112 -1300 -86
rect -1274 -112 -1234 -86
rect -1208 -112 -1168 -86
rect -1142 -112 -1102 -86
rect -1076 -112 -1036 -86
rect -1010 -112 -970 -86
rect -944 -112 -904 -86
rect -878 -112 -838 -86
rect -812 -112 -772 -86
rect -746 -112 -706 -86
rect -680 -112 -640 -86
rect -614 -112 -574 -86
rect -548 -112 -508 -86
rect -482 -112 -442 -86
rect -416 -112 -376 -86
rect -350 -112 -310 -86
rect -284 -112 -244 -86
rect -218 -112 -178 -86
rect -152 -112 -112 -86
rect -86 -112 -46 -86
rect -20 -112 20 -86
rect 46 -112 86 -86
rect 112 -112 152 -86
rect 178 -112 218 -86
rect 244 -112 284 -86
rect 310 -112 350 -86
rect 376 -112 416 -86
rect 442 -112 482 -86
rect 508 -112 548 -86
rect 574 -112 614 -86
rect 640 -112 680 -86
rect 706 -112 746 -86
rect 772 -112 812 -86
rect 838 -112 878 -86
rect 904 -112 944 -86
rect 970 -112 1010 -86
rect 1036 -112 1076 -86
rect 1102 -112 1142 -86
rect 1168 -112 1208 -86
rect 1234 -112 1274 -86
rect 1300 -112 1340 -86
rect 1366 -112 1406 -86
rect 1432 -112 1472 -86
rect 1498 -112 1538 -86
rect 1564 -112 1604 -86
rect 1630 -112 1670 -86
rect 1696 -112 1736 -86
rect 1762 -112 1802 -86
rect 1828 -112 1868 -86
rect 1894 -112 1934 -86
rect 1960 -112 2000 -86
rect 2026 -112 2066 -86
rect 2092 -112 2132 -86
rect 2158 -112 2198 -86
rect 2224 -112 2264 -86
rect 2290 -112 2330 -86
rect 2356 -112 2396 -86
rect 2422 -112 2462 -86
rect 2488 -112 2528 -86
rect 2554 -112 2594 -86
rect 2620 -112 2626 -86
rect -2626 -152 2626 -112
rect -2626 -178 -2620 -152
rect -2594 -178 -2554 -152
rect -2528 -178 -2488 -152
rect -2462 -178 -2422 -152
rect -2396 -178 -2356 -152
rect -2330 -178 -2290 -152
rect -2264 -178 -2224 -152
rect -2198 -178 -2158 -152
rect -2132 -178 -2092 -152
rect -2066 -178 -2026 -152
rect -2000 -178 -1960 -152
rect -1934 -178 -1894 -152
rect -1868 -178 -1828 -152
rect -1802 -178 -1762 -152
rect -1736 -178 -1696 -152
rect -1670 -178 -1630 -152
rect -1604 -178 -1564 -152
rect -1538 -178 -1498 -152
rect -1472 -178 -1432 -152
rect -1406 -178 -1366 -152
rect -1340 -178 -1300 -152
rect -1274 -178 -1234 -152
rect -1208 -178 -1168 -152
rect -1142 -178 -1102 -152
rect -1076 -178 -1036 -152
rect -1010 -178 -970 -152
rect -944 -178 -904 -152
rect -878 -178 -838 -152
rect -812 -178 -772 -152
rect -746 -178 -706 -152
rect -680 -178 -640 -152
rect -614 -178 -574 -152
rect -548 -178 -508 -152
rect -482 -178 -442 -152
rect -416 -178 -376 -152
rect -350 -178 -310 -152
rect -284 -178 -244 -152
rect -218 -178 -178 -152
rect -152 -178 -112 -152
rect -86 -178 -46 -152
rect -20 -178 20 -152
rect 46 -178 86 -152
rect 112 -178 152 -152
rect 178 -178 218 -152
rect 244 -178 284 -152
rect 310 -178 350 -152
rect 376 -178 416 -152
rect 442 -178 482 -152
rect 508 -178 548 -152
rect 574 -178 614 -152
rect 640 -178 680 -152
rect 706 -178 746 -152
rect 772 -178 812 -152
rect 838 -178 878 -152
rect 904 -178 944 -152
rect 970 -178 1010 -152
rect 1036 -178 1076 -152
rect 1102 -178 1142 -152
rect 1168 -178 1208 -152
rect 1234 -178 1274 -152
rect 1300 -178 1340 -152
rect 1366 -178 1406 -152
rect 1432 -178 1472 -152
rect 1498 -178 1538 -152
rect 1564 -178 1604 -152
rect 1630 -178 1670 -152
rect 1696 -178 1736 -152
rect 1762 -178 1802 -152
rect 1828 -178 1868 -152
rect 1894 -178 1934 -152
rect 1960 -178 2000 -152
rect 2026 -178 2066 -152
rect 2092 -178 2132 -152
rect 2158 -178 2198 -152
rect 2224 -178 2264 -152
rect 2290 -178 2330 -152
rect 2356 -178 2396 -152
rect 2422 -178 2462 -152
rect 2488 -178 2528 -152
rect 2554 -178 2594 -152
rect 2620 -178 2626 -152
rect -2626 -218 2626 -178
rect -2626 -244 -2620 -218
rect -2594 -244 -2554 -218
rect -2528 -244 -2488 -218
rect -2462 -244 -2422 -218
rect -2396 -244 -2356 -218
rect -2330 -244 -2290 -218
rect -2264 -244 -2224 -218
rect -2198 -244 -2158 -218
rect -2132 -244 -2092 -218
rect -2066 -244 -2026 -218
rect -2000 -244 -1960 -218
rect -1934 -244 -1894 -218
rect -1868 -244 -1828 -218
rect -1802 -244 -1762 -218
rect -1736 -244 -1696 -218
rect -1670 -244 -1630 -218
rect -1604 -244 -1564 -218
rect -1538 -244 -1498 -218
rect -1472 -244 -1432 -218
rect -1406 -244 -1366 -218
rect -1340 -244 -1300 -218
rect -1274 -244 -1234 -218
rect -1208 -244 -1168 -218
rect -1142 -244 -1102 -218
rect -1076 -244 -1036 -218
rect -1010 -244 -970 -218
rect -944 -244 -904 -218
rect -878 -244 -838 -218
rect -812 -244 -772 -218
rect -746 -244 -706 -218
rect -680 -244 -640 -218
rect -614 -244 -574 -218
rect -548 -244 -508 -218
rect -482 -244 -442 -218
rect -416 -244 -376 -218
rect -350 -244 -310 -218
rect -284 -244 -244 -218
rect -218 -244 -178 -218
rect -152 -244 -112 -218
rect -86 -244 -46 -218
rect -20 -244 20 -218
rect 46 -244 86 -218
rect 112 -244 152 -218
rect 178 -244 218 -218
rect 244 -244 284 -218
rect 310 -244 350 -218
rect 376 -244 416 -218
rect 442 -244 482 -218
rect 508 -244 548 -218
rect 574 -244 614 -218
rect 640 -244 680 -218
rect 706 -244 746 -218
rect 772 -244 812 -218
rect 838 -244 878 -218
rect 904 -244 944 -218
rect 970 -244 1010 -218
rect 1036 -244 1076 -218
rect 1102 -244 1142 -218
rect 1168 -244 1208 -218
rect 1234 -244 1274 -218
rect 1300 -244 1340 -218
rect 1366 -244 1406 -218
rect 1432 -244 1472 -218
rect 1498 -244 1538 -218
rect 1564 -244 1604 -218
rect 1630 -244 1670 -218
rect 1696 -244 1736 -218
rect 1762 -244 1802 -218
rect 1828 -244 1868 -218
rect 1894 -244 1934 -218
rect 1960 -244 2000 -218
rect 2026 -244 2066 -218
rect 2092 -244 2132 -218
rect 2158 -244 2198 -218
rect 2224 -244 2264 -218
rect 2290 -244 2330 -218
rect 2356 -244 2396 -218
rect 2422 -244 2462 -218
rect 2488 -244 2528 -218
rect 2554 -244 2594 -218
rect 2620 -244 2626 -218
rect -2626 -284 2626 -244
rect -2626 -310 -2620 -284
rect -2594 -310 -2554 -284
rect -2528 -310 -2488 -284
rect -2462 -310 -2422 -284
rect -2396 -310 -2356 -284
rect -2330 -310 -2290 -284
rect -2264 -310 -2224 -284
rect -2198 -310 -2158 -284
rect -2132 -310 -2092 -284
rect -2066 -310 -2026 -284
rect -2000 -310 -1960 -284
rect -1934 -310 -1894 -284
rect -1868 -310 -1828 -284
rect -1802 -310 -1762 -284
rect -1736 -310 -1696 -284
rect -1670 -310 -1630 -284
rect -1604 -310 -1564 -284
rect -1538 -310 -1498 -284
rect -1472 -310 -1432 -284
rect -1406 -310 -1366 -284
rect -1340 -310 -1300 -284
rect -1274 -310 -1234 -284
rect -1208 -310 -1168 -284
rect -1142 -310 -1102 -284
rect -1076 -310 -1036 -284
rect -1010 -310 -970 -284
rect -944 -310 -904 -284
rect -878 -310 -838 -284
rect -812 -310 -772 -284
rect -746 -310 -706 -284
rect -680 -310 -640 -284
rect -614 -310 -574 -284
rect -548 -310 -508 -284
rect -482 -310 -442 -284
rect -416 -310 -376 -284
rect -350 -310 -310 -284
rect -284 -310 -244 -284
rect -218 -310 -178 -284
rect -152 -310 -112 -284
rect -86 -310 -46 -284
rect -20 -310 20 -284
rect 46 -310 86 -284
rect 112 -310 152 -284
rect 178 -310 218 -284
rect 244 -310 284 -284
rect 310 -310 350 -284
rect 376 -310 416 -284
rect 442 -310 482 -284
rect 508 -310 548 -284
rect 574 -310 614 -284
rect 640 -310 680 -284
rect 706 -310 746 -284
rect 772 -310 812 -284
rect 838 -310 878 -284
rect 904 -310 944 -284
rect 970 -310 1010 -284
rect 1036 -310 1076 -284
rect 1102 -310 1142 -284
rect 1168 -310 1208 -284
rect 1234 -310 1274 -284
rect 1300 -310 1340 -284
rect 1366 -310 1406 -284
rect 1432 -310 1472 -284
rect 1498 -310 1538 -284
rect 1564 -310 1604 -284
rect 1630 -310 1670 -284
rect 1696 -310 1736 -284
rect 1762 -310 1802 -284
rect 1828 -310 1868 -284
rect 1894 -310 1934 -284
rect 1960 -310 2000 -284
rect 2026 -310 2066 -284
rect 2092 -310 2132 -284
rect 2158 -310 2198 -284
rect 2224 -310 2264 -284
rect 2290 -310 2330 -284
rect 2356 -310 2396 -284
rect 2422 -310 2462 -284
rect 2488 -310 2528 -284
rect 2554 -310 2594 -284
rect 2620 -310 2626 -284
rect -2626 -350 2626 -310
rect -2626 -376 -2620 -350
rect -2594 -376 -2554 -350
rect -2528 -376 -2488 -350
rect -2462 -376 -2422 -350
rect -2396 -376 -2356 -350
rect -2330 -376 -2290 -350
rect -2264 -376 -2224 -350
rect -2198 -376 -2158 -350
rect -2132 -376 -2092 -350
rect -2066 -376 -2026 -350
rect -2000 -376 -1960 -350
rect -1934 -376 -1894 -350
rect -1868 -376 -1828 -350
rect -1802 -376 -1762 -350
rect -1736 -376 -1696 -350
rect -1670 -376 -1630 -350
rect -1604 -376 -1564 -350
rect -1538 -376 -1498 -350
rect -1472 -376 -1432 -350
rect -1406 -376 -1366 -350
rect -1340 -376 -1300 -350
rect -1274 -376 -1234 -350
rect -1208 -376 -1168 -350
rect -1142 -376 -1102 -350
rect -1076 -376 -1036 -350
rect -1010 -376 -970 -350
rect -944 -376 -904 -350
rect -878 -376 -838 -350
rect -812 -376 -772 -350
rect -746 -376 -706 -350
rect -680 -376 -640 -350
rect -614 -376 -574 -350
rect -548 -376 -508 -350
rect -482 -376 -442 -350
rect -416 -376 -376 -350
rect -350 -376 -310 -350
rect -284 -376 -244 -350
rect -218 -376 -178 -350
rect -152 -376 -112 -350
rect -86 -376 -46 -350
rect -20 -376 20 -350
rect 46 -376 86 -350
rect 112 -376 152 -350
rect 178 -376 218 -350
rect 244 -376 284 -350
rect 310 -376 350 -350
rect 376 -376 416 -350
rect 442 -376 482 -350
rect 508 -376 548 -350
rect 574 -376 614 -350
rect 640 -376 680 -350
rect 706 -376 746 -350
rect 772 -376 812 -350
rect 838 -376 878 -350
rect 904 -376 944 -350
rect 970 -376 1010 -350
rect 1036 -376 1076 -350
rect 1102 -376 1142 -350
rect 1168 -376 1208 -350
rect 1234 -376 1274 -350
rect 1300 -376 1340 -350
rect 1366 -376 1406 -350
rect 1432 -376 1472 -350
rect 1498 -376 1538 -350
rect 1564 -376 1604 -350
rect 1630 -376 1670 -350
rect 1696 -376 1736 -350
rect 1762 -376 1802 -350
rect 1828 -376 1868 -350
rect 1894 -376 1934 -350
rect 1960 -376 2000 -350
rect 2026 -376 2066 -350
rect 2092 -376 2132 -350
rect 2158 -376 2198 -350
rect 2224 -376 2264 -350
rect 2290 -376 2330 -350
rect 2356 -376 2396 -350
rect 2422 -376 2462 -350
rect 2488 -376 2528 -350
rect 2554 -376 2594 -350
rect 2620 -376 2626 -350
rect -2626 -382 2626 -376
<< end >>
