magic
tech gf180mcuC
magscale 1 10
timestamp 1683999746
<< error_p >>
rect -34 69 -23 115
rect -118 -23 -107 23
rect 50 -23 61 23
rect -34 -115 -23 -69
<< pwell >>
rect -282 -244 282 244
<< nmos >>
rect -28 -22 28 22
<< ndiff >>
rect -120 23 -48 36
rect -120 -23 -107 23
rect -61 22 -48 23
rect 48 23 120 36
rect 48 22 61 23
rect -61 -22 -28 22
rect 28 -22 61 22
rect -61 -23 -48 -22
rect -120 -36 -48 -23
rect 48 -23 61 -22
rect 107 -23 120 23
rect 48 -36 120 -23
<< ndiffc >>
rect -107 -23 -61 23
rect 61 -23 107 23
<< psubdiff >>
rect -258 148 258 220
rect -258 104 -186 148
rect -258 -104 -245 104
rect -199 -104 -186 104
rect 186 104 258 148
rect -258 -148 -186 -104
rect 186 -104 199 104
rect 245 -104 258 104
rect 186 -148 258 -104
rect -258 -220 258 -148
<< psubdiffcont >>
rect -245 -104 -199 104
rect 199 -104 245 104
<< polysilicon >>
rect -36 115 36 128
rect -36 69 -23 115
rect 23 69 36 115
rect -36 56 36 69
rect -28 22 28 56
rect -28 -56 28 -22
rect -36 -69 36 -56
rect -36 -115 -23 -69
rect 23 -115 36 -69
rect -36 -128 36 -115
<< polycontact >>
rect -23 69 23 115
rect -23 -115 23 -69
<< metal1 >>
rect -245 161 245 207
rect -245 104 -199 161
rect -34 69 -23 115
rect 23 69 34 115
rect 199 104 245 161
rect -118 -23 -107 23
rect -61 -23 -50 23
rect 50 -23 61 23
rect 107 -23 118 23
rect -245 -161 -199 -104
rect -34 -115 -23 -69
rect 23 -115 34 -69
rect 199 -161 245 -104
rect -245 -207 245 -161
<< properties >>
string FIXED_BBOX -222 -184 222 184
string gencell nmos_3p3
string library gf180mcu
string parameters w 0.220 l 0.280 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 1 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
