magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -19343 -2975 19343 2975
<< psubdiff >>
rect -17343 953 17343 975
rect -17343 907 -17321 953
rect -17275 907 -17197 953
rect -17151 907 -17073 953
rect -17027 907 -16949 953
rect -16903 907 -16825 953
rect -16779 907 -16701 953
rect -16655 907 -16577 953
rect -16531 907 -16453 953
rect -16407 907 -16329 953
rect -16283 907 -16205 953
rect -16159 907 -16081 953
rect -16035 907 -15957 953
rect -15911 907 -15833 953
rect -15787 907 -15709 953
rect -15663 907 -15585 953
rect -15539 907 -15461 953
rect -15415 907 -15337 953
rect -15291 907 -15213 953
rect -15167 907 -15089 953
rect -15043 907 -14965 953
rect -14919 907 -14841 953
rect -14795 907 -14717 953
rect -14671 907 -14593 953
rect -14547 907 -14469 953
rect -14423 907 -14345 953
rect -14299 907 -14221 953
rect -14175 907 -14097 953
rect -14051 907 -13973 953
rect -13927 907 -13849 953
rect -13803 907 -13725 953
rect -13679 907 -13601 953
rect -13555 907 -13477 953
rect -13431 907 -13353 953
rect -13307 907 -13229 953
rect -13183 907 -13105 953
rect -13059 907 -12981 953
rect -12935 907 -12857 953
rect -12811 907 -12733 953
rect -12687 907 -12609 953
rect -12563 907 -12485 953
rect -12439 907 -12361 953
rect -12315 907 -12237 953
rect -12191 907 -12113 953
rect -12067 907 -11989 953
rect -11943 907 -11865 953
rect -11819 907 -11741 953
rect -11695 907 -11617 953
rect -11571 907 -11493 953
rect -11447 907 -11369 953
rect -11323 907 -11245 953
rect -11199 907 -11121 953
rect -11075 907 -10997 953
rect -10951 907 -10873 953
rect -10827 907 -10749 953
rect -10703 907 -10625 953
rect -10579 907 -10501 953
rect -10455 907 -10377 953
rect -10331 907 -10253 953
rect -10207 907 -10129 953
rect -10083 907 -10005 953
rect -9959 907 -9881 953
rect -9835 907 -9757 953
rect -9711 907 -9633 953
rect -9587 907 -9509 953
rect -9463 907 -9385 953
rect -9339 907 -9261 953
rect -9215 907 -9137 953
rect -9091 907 -9013 953
rect -8967 907 -8889 953
rect -8843 907 -8765 953
rect -8719 907 -8641 953
rect -8595 907 -8517 953
rect -8471 907 -8393 953
rect -8347 907 -8269 953
rect -8223 907 -8145 953
rect -8099 907 -8021 953
rect -7975 907 -7897 953
rect -7851 907 -7773 953
rect -7727 907 -7649 953
rect -7603 907 -7525 953
rect -7479 907 -7401 953
rect -7355 907 -7277 953
rect -7231 907 -7153 953
rect -7107 907 -7029 953
rect -6983 907 -6905 953
rect -6859 907 -6781 953
rect -6735 907 -6657 953
rect -6611 907 -6533 953
rect -6487 907 -6409 953
rect -6363 907 -6285 953
rect -6239 907 -6161 953
rect -6115 907 -6037 953
rect -5991 907 -5913 953
rect -5867 907 -5789 953
rect -5743 907 -5665 953
rect -5619 907 -5541 953
rect -5495 907 -5417 953
rect -5371 907 -5293 953
rect -5247 907 -5169 953
rect -5123 907 -5045 953
rect -4999 907 -4921 953
rect -4875 907 -4797 953
rect -4751 907 -4673 953
rect -4627 907 -4549 953
rect -4503 907 -4425 953
rect -4379 907 -4301 953
rect -4255 907 -4177 953
rect -4131 907 -4053 953
rect -4007 907 -3929 953
rect -3883 907 -3805 953
rect -3759 907 -3681 953
rect -3635 907 -3557 953
rect -3511 907 -3433 953
rect -3387 907 -3309 953
rect -3263 907 -3185 953
rect -3139 907 -3061 953
rect -3015 907 -2937 953
rect -2891 907 -2813 953
rect -2767 907 -2689 953
rect -2643 907 -2565 953
rect -2519 907 -2441 953
rect -2395 907 -2317 953
rect -2271 907 -2193 953
rect -2147 907 -2069 953
rect -2023 907 -1945 953
rect -1899 907 -1821 953
rect -1775 907 -1697 953
rect -1651 907 -1573 953
rect -1527 907 -1449 953
rect -1403 907 -1325 953
rect -1279 907 -1201 953
rect -1155 907 -1077 953
rect -1031 907 -953 953
rect -907 907 -829 953
rect -783 907 -705 953
rect -659 907 -581 953
rect -535 907 -457 953
rect -411 907 -333 953
rect -287 907 -209 953
rect -163 907 -85 953
rect -39 907 39 953
rect 85 907 163 953
rect 209 907 287 953
rect 333 907 411 953
rect 457 907 535 953
rect 581 907 659 953
rect 705 907 783 953
rect 829 907 907 953
rect 953 907 1031 953
rect 1077 907 1155 953
rect 1201 907 1279 953
rect 1325 907 1403 953
rect 1449 907 1527 953
rect 1573 907 1651 953
rect 1697 907 1775 953
rect 1821 907 1899 953
rect 1945 907 2023 953
rect 2069 907 2147 953
rect 2193 907 2271 953
rect 2317 907 2395 953
rect 2441 907 2519 953
rect 2565 907 2643 953
rect 2689 907 2767 953
rect 2813 907 2891 953
rect 2937 907 3015 953
rect 3061 907 3139 953
rect 3185 907 3263 953
rect 3309 907 3387 953
rect 3433 907 3511 953
rect 3557 907 3635 953
rect 3681 907 3759 953
rect 3805 907 3883 953
rect 3929 907 4007 953
rect 4053 907 4131 953
rect 4177 907 4255 953
rect 4301 907 4379 953
rect 4425 907 4503 953
rect 4549 907 4627 953
rect 4673 907 4751 953
rect 4797 907 4875 953
rect 4921 907 4999 953
rect 5045 907 5123 953
rect 5169 907 5247 953
rect 5293 907 5371 953
rect 5417 907 5495 953
rect 5541 907 5619 953
rect 5665 907 5743 953
rect 5789 907 5867 953
rect 5913 907 5991 953
rect 6037 907 6115 953
rect 6161 907 6239 953
rect 6285 907 6363 953
rect 6409 907 6487 953
rect 6533 907 6611 953
rect 6657 907 6735 953
rect 6781 907 6859 953
rect 6905 907 6983 953
rect 7029 907 7107 953
rect 7153 907 7231 953
rect 7277 907 7355 953
rect 7401 907 7479 953
rect 7525 907 7603 953
rect 7649 907 7727 953
rect 7773 907 7851 953
rect 7897 907 7975 953
rect 8021 907 8099 953
rect 8145 907 8223 953
rect 8269 907 8347 953
rect 8393 907 8471 953
rect 8517 907 8595 953
rect 8641 907 8719 953
rect 8765 907 8843 953
rect 8889 907 8967 953
rect 9013 907 9091 953
rect 9137 907 9215 953
rect 9261 907 9339 953
rect 9385 907 9463 953
rect 9509 907 9587 953
rect 9633 907 9711 953
rect 9757 907 9835 953
rect 9881 907 9959 953
rect 10005 907 10083 953
rect 10129 907 10207 953
rect 10253 907 10331 953
rect 10377 907 10455 953
rect 10501 907 10579 953
rect 10625 907 10703 953
rect 10749 907 10827 953
rect 10873 907 10951 953
rect 10997 907 11075 953
rect 11121 907 11199 953
rect 11245 907 11323 953
rect 11369 907 11447 953
rect 11493 907 11571 953
rect 11617 907 11695 953
rect 11741 907 11819 953
rect 11865 907 11943 953
rect 11989 907 12067 953
rect 12113 907 12191 953
rect 12237 907 12315 953
rect 12361 907 12439 953
rect 12485 907 12563 953
rect 12609 907 12687 953
rect 12733 907 12811 953
rect 12857 907 12935 953
rect 12981 907 13059 953
rect 13105 907 13183 953
rect 13229 907 13307 953
rect 13353 907 13431 953
rect 13477 907 13555 953
rect 13601 907 13679 953
rect 13725 907 13803 953
rect 13849 907 13927 953
rect 13973 907 14051 953
rect 14097 907 14175 953
rect 14221 907 14299 953
rect 14345 907 14423 953
rect 14469 907 14547 953
rect 14593 907 14671 953
rect 14717 907 14795 953
rect 14841 907 14919 953
rect 14965 907 15043 953
rect 15089 907 15167 953
rect 15213 907 15291 953
rect 15337 907 15415 953
rect 15461 907 15539 953
rect 15585 907 15663 953
rect 15709 907 15787 953
rect 15833 907 15911 953
rect 15957 907 16035 953
rect 16081 907 16159 953
rect 16205 907 16283 953
rect 16329 907 16407 953
rect 16453 907 16531 953
rect 16577 907 16655 953
rect 16701 907 16779 953
rect 16825 907 16903 953
rect 16949 907 17027 953
rect 17073 907 17151 953
rect 17197 907 17275 953
rect 17321 907 17343 953
rect -17343 829 17343 907
rect -17343 783 -17321 829
rect -17275 783 -17197 829
rect -17151 783 -17073 829
rect -17027 783 -16949 829
rect -16903 783 -16825 829
rect -16779 783 -16701 829
rect -16655 783 -16577 829
rect -16531 783 -16453 829
rect -16407 783 -16329 829
rect -16283 783 -16205 829
rect -16159 783 -16081 829
rect -16035 783 -15957 829
rect -15911 783 -15833 829
rect -15787 783 -15709 829
rect -15663 783 -15585 829
rect -15539 783 -15461 829
rect -15415 783 -15337 829
rect -15291 783 -15213 829
rect -15167 783 -15089 829
rect -15043 783 -14965 829
rect -14919 783 -14841 829
rect -14795 783 -14717 829
rect -14671 783 -14593 829
rect -14547 783 -14469 829
rect -14423 783 -14345 829
rect -14299 783 -14221 829
rect -14175 783 -14097 829
rect -14051 783 -13973 829
rect -13927 783 -13849 829
rect -13803 783 -13725 829
rect -13679 783 -13601 829
rect -13555 783 -13477 829
rect -13431 783 -13353 829
rect -13307 783 -13229 829
rect -13183 783 -13105 829
rect -13059 783 -12981 829
rect -12935 783 -12857 829
rect -12811 783 -12733 829
rect -12687 783 -12609 829
rect -12563 783 -12485 829
rect -12439 783 -12361 829
rect -12315 783 -12237 829
rect -12191 783 -12113 829
rect -12067 783 -11989 829
rect -11943 783 -11865 829
rect -11819 783 -11741 829
rect -11695 783 -11617 829
rect -11571 783 -11493 829
rect -11447 783 -11369 829
rect -11323 783 -11245 829
rect -11199 783 -11121 829
rect -11075 783 -10997 829
rect -10951 783 -10873 829
rect -10827 783 -10749 829
rect -10703 783 -10625 829
rect -10579 783 -10501 829
rect -10455 783 -10377 829
rect -10331 783 -10253 829
rect -10207 783 -10129 829
rect -10083 783 -10005 829
rect -9959 783 -9881 829
rect -9835 783 -9757 829
rect -9711 783 -9633 829
rect -9587 783 -9509 829
rect -9463 783 -9385 829
rect -9339 783 -9261 829
rect -9215 783 -9137 829
rect -9091 783 -9013 829
rect -8967 783 -8889 829
rect -8843 783 -8765 829
rect -8719 783 -8641 829
rect -8595 783 -8517 829
rect -8471 783 -8393 829
rect -8347 783 -8269 829
rect -8223 783 -8145 829
rect -8099 783 -8021 829
rect -7975 783 -7897 829
rect -7851 783 -7773 829
rect -7727 783 -7649 829
rect -7603 783 -7525 829
rect -7479 783 -7401 829
rect -7355 783 -7277 829
rect -7231 783 -7153 829
rect -7107 783 -7029 829
rect -6983 783 -6905 829
rect -6859 783 -6781 829
rect -6735 783 -6657 829
rect -6611 783 -6533 829
rect -6487 783 -6409 829
rect -6363 783 -6285 829
rect -6239 783 -6161 829
rect -6115 783 -6037 829
rect -5991 783 -5913 829
rect -5867 783 -5789 829
rect -5743 783 -5665 829
rect -5619 783 -5541 829
rect -5495 783 -5417 829
rect -5371 783 -5293 829
rect -5247 783 -5169 829
rect -5123 783 -5045 829
rect -4999 783 -4921 829
rect -4875 783 -4797 829
rect -4751 783 -4673 829
rect -4627 783 -4549 829
rect -4503 783 -4425 829
rect -4379 783 -4301 829
rect -4255 783 -4177 829
rect -4131 783 -4053 829
rect -4007 783 -3929 829
rect -3883 783 -3805 829
rect -3759 783 -3681 829
rect -3635 783 -3557 829
rect -3511 783 -3433 829
rect -3387 783 -3309 829
rect -3263 783 -3185 829
rect -3139 783 -3061 829
rect -3015 783 -2937 829
rect -2891 783 -2813 829
rect -2767 783 -2689 829
rect -2643 783 -2565 829
rect -2519 783 -2441 829
rect -2395 783 -2317 829
rect -2271 783 -2193 829
rect -2147 783 -2069 829
rect -2023 783 -1945 829
rect -1899 783 -1821 829
rect -1775 783 -1697 829
rect -1651 783 -1573 829
rect -1527 783 -1449 829
rect -1403 783 -1325 829
rect -1279 783 -1201 829
rect -1155 783 -1077 829
rect -1031 783 -953 829
rect -907 783 -829 829
rect -783 783 -705 829
rect -659 783 -581 829
rect -535 783 -457 829
rect -411 783 -333 829
rect -287 783 -209 829
rect -163 783 -85 829
rect -39 783 39 829
rect 85 783 163 829
rect 209 783 287 829
rect 333 783 411 829
rect 457 783 535 829
rect 581 783 659 829
rect 705 783 783 829
rect 829 783 907 829
rect 953 783 1031 829
rect 1077 783 1155 829
rect 1201 783 1279 829
rect 1325 783 1403 829
rect 1449 783 1527 829
rect 1573 783 1651 829
rect 1697 783 1775 829
rect 1821 783 1899 829
rect 1945 783 2023 829
rect 2069 783 2147 829
rect 2193 783 2271 829
rect 2317 783 2395 829
rect 2441 783 2519 829
rect 2565 783 2643 829
rect 2689 783 2767 829
rect 2813 783 2891 829
rect 2937 783 3015 829
rect 3061 783 3139 829
rect 3185 783 3263 829
rect 3309 783 3387 829
rect 3433 783 3511 829
rect 3557 783 3635 829
rect 3681 783 3759 829
rect 3805 783 3883 829
rect 3929 783 4007 829
rect 4053 783 4131 829
rect 4177 783 4255 829
rect 4301 783 4379 829
rect 4425 783 4503 829
rect 4549 783 4627 829
rect 4673 783 4751 829
rect 4797 783 4875 829
rect 4921 783 4999 829
rect 5045 783 5123 829
rect 5169 783 5247 829
rect 5293 783 5371 829
rect 5417 783 5495 829
rect 5541 783 5619 829
rect 5665 783 5743 829
rect 5789 783 5867 829
rect 5913 783 5991 829
rect 6037 783 6115 829
rect 6161 783 6239 829
rect 6285 783 6363 829
rect 6409 783 6487 829
rect 6533 783 6611 829
rect 6657 783 6735 829
rect 6781 783 6859 829
rect 6905 783 6983 829
rect 7029 783 7107 829
rect 7153 783 7231 829
rect 7277 783 7355 829
rect 7401 783 7479 829
rect 7525 783 7603 829
rect 7649 783 7727 829
rect 7773 783 7851 829
rect 7897 783 7975 829
rect 8021 783 8099 829
rect 8145 783 8223 829
rect 8269 783 8347 829
rect 8393 783 8471 829
rect 8517 783 8595 829
rect 8641 783 8719 829
rect 8765 783 8843 829
rect 8889 783 8967 829
rect 9013 783 9091 829
rect 9137 783 9215 829
rect 9261 783 9339 829
rect 9385 783 9463 829
rect 9509 783 9587 829
rect 9633 783 9711 829
rect 9757 783 9835 829
rect 9881 783 9959 829
rect 10005 783 10083 829
rect 10129 783 10207 829
rect 10253 783 10331 829
rect 10377 783 10455 829
rect 10501 783 10579 829
rect 10625 783 10703 829
rect 10749 783 10827 829
rect 10873 783 10951 829
rect 10997 783 11075 829
rect 11121 783 11199 829
rect 11245 783 11323 829
rect 11369 783 11447 829
rect 11493 783 11571 829
rect 11617 783 11695 829
rect 11741 783 11819 829
rect 11865 783 11943 829
rect 11989 783 12067 829
rect 12113 783 12191 829
rect 12237 783 12315 829
rect 12361 783 12439 829
rect 12485 783 12563 829
rect 12609 783 12687 829
rect 12733 783 12811 829
rect 12857 783 12935 829
rect 12981 783 13059 829
rect 13105 783 13183 829
rect 13229 783 13307 829
rect 13353 783 13431 829
rect 13477 783 13555 829
rect 13601 783 13679 829
rect 13725 783 13803 829
rect 13849 783 13927 829
rect 13973 783 14051 829
rect 14097 783 14175 829
rect 14221 783 14299 829
rect 14345 783 14423 829
rect 14469 783 14547 829
rect 14593 783 14671 829
rect 14717 783 14795 829
rect 14841 783 14919 829
rect 14965 783 15043 829
rect 15089 783 15167 829
rect 15213 783 15291 829
rect 15337 783 15415 829
rect 15461 783 15539 829
rect 15585 783 15663 829
rect 15709 783 15787 829
rect 15833 783 15911 829
rect 15957 783 16035 829
rect 16081 783 16159 829
rect 16205 783 16283 829
rect 16329 783 16407 829
rect 16453 783 16531 829
rect 16577 783 16655 829
rect 16701 783 16779 829
rect 16825 783 16903 829
rect 16949 783 17027 829
rect 17073 783 17151 829
rect 17197 783 17275 829
rect 17321 783 17343 829
rect -17343 705 17343 783
rect -17343 659 -17321 705
rect -17275 659 -17197 705
rect -17151 659 -17073 705
rect -17027 659 -16949 705
rect -16903 659 -16825 705
rect -16779 659 -16701 705
rect -16655 659 -16577 705
rect -16531 659 -16453 705
rect -16407 659 -16329 705
rect -16283 659 -16205 705
rect -16159 659 -16081 705
rect -16035 659 -15957 705
rect -15911 659 -15833 705
rect -15787 659 -15709 705
rect -15663 659 -15585 705
rect -15539 659 -15461 705
rect -15415 659 -15337 705
rect -15291 659 -15213 705
rect -15167 659 -15089 705
rect -15043 659 -14965 705
rect -14919 659 -14841 705
rect -14795 659 -14717 705
rect -14671 659 -14593 705
rect -14547 659 -14469 705
rect -14423 659 -14345 705
rect -14299 659 -14221 705
rect -14175 659 -14097 705
rect -14051 659 -13973 705
rect -13927 659 -13849 705
rect -13803 659 -13725 705
rect -13679 659 -13601 705
rect -13555 659 -13477 705
rect -13431 659 -13353 705
rect -13307 659 -13229 705
rect -13183 659 -13105 705
rect -13059 659 -12981 705
rect -12935 659 -12857 705
rect -12811 659 -12733 705
rect -12687 659 -12609 705
rect -12563 659 -12485 705
rect -12439 659 -12361 705
rect -12315 659 -12237 705
rect -12191 659 -12113 705
rect -12067 659 -11989 705
rect -11943 659 -11865 705
rect -11819 659 -11741 705
rect -11695 659 -11617 705
rect -11571 659 -11493 705
rect -11447 659 -11369 705
rect -11323 659 -11245 705
rect -11199 659 -11121 705
rect -11075 659 -10997 705
rect -10951 659 -10873 705
rect -10827 659 -10749 705
rect -10703 659 -10625 705
rect -10579 659 -10501 705
rect -10455 659 -10377 705
rect -10331 659 -10253 705
rect -10207 659 -10129 705
rect -10083 659 -10005 705
rect -9959 659 -9881 705
rect -9835 659 -9757 705
rect -9711 659 -9633 705
rect -9587 659 -9509 705
rect -9463 659 -9385 705
rect -9339 659 -9261 705
rect -9215 659 -9137 705
rect -9091 659 -9013 705
rect -8967 659 -8889 705
rect -8843 659 -8765 705
rect -8719 659 -8641 705
rect -8595 659 -8517 705
rect -8471 659 -8393 705
rect -8347 659 -8269 705
rect -8223 659 -8145 705
rect -8099 659 -8021 705
rect -7975 659 -7897 705
rect -7851 659 -7773 705
rect -7727 659 -7649 705
rect -7603 659 -7525 705
rect -7479 659 -7401 705
rect -7355 659 -7277 705
rect -7231 659 -7153 705
rect -7107 659 -7029 705
rect -6983 659 -6905 705
rect -6859 659 -6781 705
rect -6735 659 -6657 705
rect -6611 659 -6533 705
rect -6487 659 -6409 705
rect -6363 659 -6285 705
rect -6239 659 -6161 705
rect -6115 659 -6037 705
rect -5991 659 -5913 705
rect -5867 659 -5789 705
rect -5743 659 -5665 705
rect -5619 659 -5541 705
rect -5495 659 -5417 705
rect -5371 659 -5293 705
rect -5247 659 -5169 705
rect -5123 659 -5045 705
rect -4999 659 -4921 705
rect -4875 659 -4797 705
rect -4751 659 -4673 705
rect -4627 659 -4549 705
rect -4503 659 -4425 705
rect -4379 659 -4301 705
rect -4255 659 -4177 705
rect -4131 659 -4053 705
rect -4007 659 -3929 705
rect -3883 659 -3805 705
rect -3759 659 -3681 705
rect -3635 659 -3557 705
rect -3511 659 -3433 705
rect -3387 659 -3309 705
rect -3263 659 -3185 705
rect -3139 659 -3061 705
rect -3015 659 -2937 705
rect -2891 659 -2813 705
rect -2767 659 -2689 705
rect -2643 659 -2565 705
rect -2519 659 -2441 705
rect -2395 659 -2317 705
rect -2271 659 -2193 705
rect -2147 659 -2069 705
rect -2023 659 -1945 705
rect -1899 659 -1821 705
rect -1775 659 -1697 705
rect -1651 659 -1573 705
rect -1527 659 -1449 705
rect -1403 659 -1325 705
rect -1279 659 -1201 705
rect -1155 659 -1077 705
rect -1031 659 -953 705
rect -907 659 -829 705
rect -783 659 -705 705
rect -659 659 -581 705
rect -535 659 -457 705
rect -411 659 -333 705
rect -287 659 -209 705
rect -163 659 -85 705
rect -39 659 39 705
rect 85 659 163 705
rect 209 659 287 705
rect 333 659 411 705
rect 457 659 535 705
rect 581 659 659 705
rect 705 659 783 705
rect 829 659 907 705
rect 953 659 1031 705
rect 1077 659 1155 705
rect 1201 659 1279 705
rect 1325 659 1403 705
rect 1449 659 1527 705
rect 1573 659 1651 705
rect 1697 659 1775 705
rect 1821 659 1899 705
rect 1945 659 2023 705
rect 2069 659 2147 705
rect 2193 659 2271 705
rect 2317 659 2395 705
rect 2441 659 2519 705
rect 2565 659 2643 705
rect 2689 659 2767 705
rect 2813 659 2891 705
rect 2937 659 3015 705
rect 3061 659 3139 705
rect 3185 659 3263 705
rect 3309 659 3387 705
rect 3433 659 3511 705
rect 3557 659 3635 705
rect 3681 659 3759 705
rect 3805 659 3883 705
rect 3929 659 4007 705
rect 4053 659 4131 705
rect 4177 659 4255 705
rect 4301 659 4379 705
rect 4425 659 4503 705
rect 4549 659 4627 705
rect 4673 659 4751 705
rect 4797 659 4875 705
rect 4921 659 4999 705
rect 5045 659 5123 705
rect 5169 659 5247 705
rect 5293 659 5371 705
rect 5417 659 5495 705
rect 5541 659 5619 705
rect 5665 659 5743 705
rect 5789 659 5867 705
rect 5913 659 5991 705
rect 6037 659 6115 705
rect 6161 659 6239 705
rect 6285 659 6363 705
rect 6409 659 6487 705
rect 6533 659 6611 705
rect 6657 659 6735 705
rect 6781 659 6859 705
rect 6905 659 6983 705
rect 7029 659 7107 705
rect 7153 659 7231 705
rect 7277 659 7355 705
rect 7401 659 7479 705
rect 7525 659 7603 705
rect 7649 659 7727 705
rect 7773 659 7851 705
rect 7897 659 7975 705
rect 8021 659 8099 705
rect 8145 659 8223 705
rect 8269 659 8347 705
rect 8393 659 8471 705
rect 8517 659 8595 705
rect 8641 659 8719 705
rect 8765 659 8843 705
rect 8889 659 8967 705
rect 9013 659 9091 705
rect 9137 659 9215 705
rect 9261 659 9339 705
rect 9385 659 9463 705
rect 9509 659 9587 705
rect 9633 659 9711 705
rect 9757 659 9835 705
rect 9881 659 9959 705
rect 10005 659 10083 705
rect 10129 659 10207 705
rect 10253 659 10331 705
rect 10377 659 10455 705
rect 10501 659 10579 705
rect 10625 659 10703 705
rect 10749 659 10827 705
rect 10873 659 10951 705
rect 10997 659 11075 705
rect 11121 659 11199 705
rect 11245 659 11323 705
rect 11369 659 11447 705
rect 11493 659 11571 705
rect 11617 659 11695 705
rect 11741 659 11819 705
rect 11865 659 11943 705
rect 11989 659 12067 705
rect 12113 659 12191 705
rect 12237 659 12315 705
rect 12361 659 12439 705
rect 12485 659 12563 705
rect 12609 659 12687 705
rect 12733 659 12811 705
rect 12857 659 12935 705
rect 12981 659 13059 705
rect 13105 659 13183 705
rect 13229 659 13307 705
rect 13353 659 13431 705
rect 13477 659 13555 705
rect 13601 659 13679 705
rect 13725 659 13803 705
rect 13849 659 13927 705
rect 13973 659 14051 705
rect 14097 659 14175 705
rect 14221 659 14299 705
rect 14345 659 14423 705
rect 14469 659 14547 705
rect 14593 659 14671 705
rect 14717 659 14795 705
rect 14841 659 14919 705
rect 14965 659 15043 705
rect 15089 659 15167 705
rect 15213 659 15291 705
rect 15337 659 15415 705
rect 15461 659 15539 705
rect 15585 659 15663 705
rect 15709 659 15787 705
rect 15833 659 15911 705
rect 15957 659 16035 705
rect 16081 659 16159 705
rect 16205 659 16283 705
rect 16329 659 16407 705
rect 16453 659 16531 705
rect 16577 659 16655 705
rect 16701 659 16779 705
rect 16825 659 16903 705
rect 16949 659 17027 705
rect 17073 659 17151 705
rect 17197 659 17275 705
rect 17321 659 17343 705
rect -17343 581 17343 659
rect -17343 535 -17321 581
rect -17275 535 -17197 581
rect -17151 535 -17073 581
rect -17027 535 -16949 581
rect -16903 535 -16825 581
rect -16779 535 -16701 581
rect -16655 535 -16577 581
rect -16531 535 -16453 581
rect -16407 535 -16329 581
rect -16283 535 -16205 581
rect -16159 535 -16081 581
rect -16035 535 -15957 581
rect -15911 535 -15833 581
rect -15787 535 -15709 581
rect -15663 535 -15585 581
rect -15539 535 -15461 581
rect -15415 535 -15337 581
rect -15291 535 -15213 581
rect -15167 535 -15089 581
rect -15043 535 -14965 581
rect -14919 535 -14841 581
rect -14795 535 -14717 581
rect -14671 535 -14593 581
rect -14547 535 -14469 581
rect -14423 535 -14345 581
rect -14299 535 -14221 581
rect -14175 535 -14097 581
rect -14051 535 -13973 581
rect -13927 535 -13849 581
rect -13803 535 -13725 581
rect -13679 535 -13601 581
rect -13555 535 -13477 581
rect -13431 535 -13353 581
rect -13307 535 -13229 581
rect -13183 535 -13105 581
rect -13059 535 -12981 581
rect -12935 535 -12857 581
rect -12811 535 -12733 581
rect -12687 535 -12609 581
rect -12563 535 -12485 581
rect -12439 535 -12361 581
rect -12315 535 -12237 581
rect -12191 535 -12113 581
rect -12067 535 -11989 581
rect -11943 535 -11865 581
rect -11819 535 -11741 581
rect -11695 535 -11617 581
rect -11571 535 -11493 581
rect -11447 535 -11369 581
rect -11323 535 -11245 581
rect -11199 535 -11121 581
rect -11075 535 -10997 581
rect -10951 535 -10873 581
rect -10827 535 -10749 581
rect -10703 535 -10625 581
rect -10579 535 -10501 581
rect -10455 535 -10377 581
rect -10331 535 -10253 581
rect -10207 535 -10129 581
rect -10083 535 -10005 581
rect -9959 535 -9881 581
rect -9835 535 -9757 581
rect -9711 535 -9633 581
rect -9587 535 -9509 581
rect -9463 535 -9385 581
rect -9339 535 -9261 581
rect -9215 535 -9137 581
rect -9091 535 -9013 581
rect -8967 535 -8889 581
rect -8843 535 -8765 581
rect -8719 535 -8641 581
rect -8595 535 -8517 581
rect -8471 535 -8393 581
rect -8347 535 -8269 581
rect -8223 535 -8145 581
rect -8099 535 -8021 581
rect -7975 535 -7897 581
rect -7851 535 -7773 581
rect -7727 535 -7649 581
rect -7603 535 -7525 581
rect -7479 535 -7401 581
rect -7355 535 -7277 581
rect -7231 535 -7153 581
rect -7107 535 -7029 581
rect -6983 535 -6905 581
rect -6859 535 -6781 581
rect -6735 535 -6657 581
rect -6611 535 -6533 581
rect -6487 535 -6409 581
rect -6363 535 -6285 581
rect -6239 535 -6161 581
rect -6115 535 -6037 581
rect -5991 535 -5913 581
rect -5867 535 -5789 581
rect -5743 535 -5665 581
rect -5619 535 -5541 581
rect -5495 535 -5417 581
rect -5371 535 -5293 581
rect -5247 535 -5169 581
rect -5123 535 -5045 581
rect -4999 535 -4921 581
rect -4875 535 -4797 581
rect -4751 535 -4673 581
rect -4627 535 -4549 581
rect -4503 535 -4425 581
rect -4379 535 -4301 581
rect -4255 535 -4177 581
rect -4131 535 -4053 581
rect -4007 535 -3929 581
rect -3883 535 -3805 581
rect -3759 535 -3681 581
rect -3635 535 -3557 581
rect -3511 535 -3433 581
rect -3387 535 -3309 581
rect -3263 535 -3185 581
rect -3139 535 -3061 581
rect -3015 535 -2937 581
rect -2891 535 -2813 581
rect -2767 535 -2689 581
rect -2643 535 -2565 581
rect -2519 535 -2441 581
rect -2395 535 -2317 581
rect -2271 535 -2193 581
rect -2147 535 -2069 581
rect -2023 535 -1945 581
rect -1899 535 -1821 581
rect -1775 535 -1697 581
rect -1651 535 -1573 581
rect -1527 535 -1449 581
rect -1403 535 -1325 581
rect -1279 535 -1201 581
rect -1155 535 -1077 581
rect -1031 535 -953 581
rect -907 535 -829 581
rect -783 535 -705 581
rect -659 535 -581 581
rect -535 535 -457 581
rect -411 535 -333 581
rect -287 535 -209 581
rect -163 535 -85 581
rect -39 535 39 581
rect 85 535 163 581
rect 209 535 287 581
rect 333 535 411 581
rect 457 535 535 581
rect 581 535 659 581
rect 705 535 783 581
rect 829 535 907 581
rect 953 535 1031 581
rect 1077 535 1155 581
rect 1201 535 1279 581
rect 1325 535 1403 581
rect 1449 535 1527 581
rect 1573 535 1651 581
rect 1697 535 1775 581
rect 1821 535 1899 581
rect 1945 535 2023 581
rect 2069 535 2147 581
rect 2193 535 2271 581
rect 2317 535 2395 581
rect 2441 535 2519 581
rect 2565 535 2643 581
rect 2689 535 2767 581
rect 2813 535 2891 581
rect 2937 535 3015 581
rect 3061 535 3139 581
rect 3185 535 3263 581
rect 3309 535 3387 581
rect 3433 535 3511 581
rect 3557 535 3635 581
rect 3681 535 3759 581
rect 3805 535 3883 581
rect 3929 535 4007 581
rect 4053 535 4131 581
rect 4177 535 4255 581
rect 4301 535 4379 581
rect 4425 535 4503 581
rect 4549 535 4627 581
rect 4673 535 4751 581
rect 4797 535 4875 581
rect 4921 535 4999 581
rect 5045 535 5123 581
rect 5169 535 5247 581
rect 5293 535 5371 581
rect 5417 535 5495 581
rect 5541 535 5619 581
rect 5665 535 5743 581
rect 5789 535 5867 581
rect 5913 535 5991 581
rect 6037 535 6115 581
rect 6161 535 6239 581
rect 6285 535 6363 581
rect 6409 535 6487 581
rect 6533 535 6611 581
rect 6657 535 6735 581
rect 6781 535 6859 581
rect 6905 535 6983 581
rect 7029 535 7107 581
rect 7153 535 7231 581
rect 7277 535 7355 581
rect 7401 535 7479 581
rect 7525 535 7603 581
rect 7649 535 7727 581
rect 7773 535 7851 581
rect 7897 535 7975 581
rect 8021 535 8099 581
rect 8145 535 8223 581
rect 8269 535 8347 581
rect 8393 535 8471 581
rect 8517 535 8595 581
rect 8641 535 8719 581
rect 8765 535 8843 581
rect 8889 535 8967 581
rect 9013 535 9091 581
rect 9137 535 9215 581
rect 9261 535 9339 581
rect 9385 535 9463 581
rect 9509 535 9587 581
rect 9633 535 9711 581
rect 9757 535 9835 581
rect 9881 535 9959 581
rect 10005 535 10083 581
rect 10129 535 10207 581
rect 10253 535 10331 581
rect 10377 535 10455 581
rect 10501 535 10579 581
rect 10625 535 10703 581
rect 10749 535 10827 581
rect 10873 535 10951 581
rect 10997 535 11075 581
rect 11121 535 11199 581
rect 11245 535 11323 581
rect 11369 535 11447 581
rect 11493 535 11571 581
rect 11617 535 11695 581
rect 11741 535 11819 581
rect 11865 535 11943 581
rect 11989 535 12067 581
rect 12113 535 12191 581
rect 12237 535 12315 581
rect 12361 535 12439 581
rect 12485 535 12563 581
rect 12609 535 12687 581
rect 12733 535 12811 581
rect 12857 535 12935 581
rect 12981 535 13059 581
rect 13105 535 13183 581
rect 13229 535 13307 581
rect 13353 535 13431 581
rect 13477 535 13555 581
rect 13601 535 13679 581
rect 13725 535 13803 581
rect 13849 535 13927 581
rect 13973 535 14051 581
rect 14097 535 14175 581
rect 14221 535 14299 581
rect 14345 535 14423 581
rect 14469 535 14547 581
rect 14593 535 14671 581
rect 14717 535 14795 581
rect 14841 535 14919 581
rect 14965 535 15043 581
rect 15089 535 15167 581
rect 15213 535 15291 581
rect 15337 535 15415 581
rect 15461 535 15539 581
rect 15585 535 15663 581
rect 15709 535 15787 581
rect 15833 535 15911 581
rect 15957 535 16035 581
rect 16081 535 16159 581
rect 16205 535 16283 581
rect 16329 535 16407 581
rect 16453 535 16531 581
rect 16577 535 16655 581
rect 16701 535 16779 581
rect 16825 535 16903 581
rect 16949 535 17027 581
rect 17073 535 17151 581
rect 17197 535 17275 581
rect 17321 535 17343 581
rect -17343 457 17343 535
rect -17343 411 -17321 457
rect -17275 411 -17197 457
rect -17151 411 -17073 457
rect -17027 411 -16949 457
rect -16903 411 -16825 457
rect -16779 411 -16701 457
rect -16655 411 -16577 457
rect -16531 411 -16453 457
rect -16407 411 -16329 457
rect -16283 411 -16205 457
rect -16159 411 -16081 457
rect -16035 411 -15957 457
rect -15911 411 -15833 457
rect -15787 411 -15709 457
rect -15663 411 -15585 457
rect -15539 411 -15461 457
rect -15415 411 -15337 457
rect -15291 411 -15213 457
rect -15167 411 -15089 457
rect -15043 411 -14965 457
rect -14919 411 -14841 457
rect -14795 411 -14717 457
rect -14671 411 -14593 457
rect -14547 411 -14469 457
rect -14423 411 -14345 457
rect -14299 411 -14221 457
rect -14175 411 -14097 457
rect -14051 411 -13973 457
rect -13927 411 -13849 457
rect -13803 411 -13725 457
rect -13679 411 -13601 457
rect -13555 411 -13477 457
rect -13431 411 -13353 457
rect -13307 411 -13229 457
rect -13183 411 -13105 457
rect -13059 411 -12981 457
rect -12935 411 -12857 457
rect -12811 411 -12733 457
rect -12687 411 -12609 457
rect -12563 411 -12485 457
rect -12439 411 -12361 457
rect -12315 411 -12237 457
rect -12191 411 -12113 457
rect -12067 411 -11989 457
rect -11943 411 -11865 457
rect -11819 411 -11741 457
rect -11695 411 -11617 457
rect -11571 411 -11493 457
rect -11447 411 -11369 457
rect -11323 411 -11245 457
rect -11199 411 -11121 457
rect -11075 411 -10997 457
rect -10951 411 -10873 457
rect -10827 411 -10749 457
rect -10703 411 -10625 457
rect -10579 411 -10501 457
rect -10455 411 -10377 457
rect -10331 411 -10253 457
rect -10207 411 -10129 457
rect -10083 411 -10005 457
rect -9959 411 -9881 457
rect -9835 411 -9757 457
rect -9711 411 -9633 457
rect -9587 411 -9509 457
rect -9463 411 -9385 457
rect -9339 411 -9261 457
rect -9215 411 -9137 457
rect -9091 411 -9013 457
rect -8967 411 -8889 457
rect -8843 411 -8765 457
rect -8719 411 -8641 457
rect -8595 411 -8517 457
rect -8471 411 -8393 457
rect -8347 411 -8269 457
rect -8223 411 -8145 457
rect -8099 411 -8021 457
rect -7975 411 -7897 457
rect -7851 411 -7773 457
rect -7727 411 -7649 457
rect -7603 411 -7525 457
rect -7479 411 -7401 457
rect -7355 411 -7277 457
rect -7231 411 -7153 457
rect -7107 411 -7029 457
rect -6983 411 -6905 457
rect -6859 411 -6781 457
rect -6735 411 -6657 457
rect -6611 411 -6533 457
rect -6487 411 -6409 457
rect -6363 411 -6285 457
rect -6239 411 -6161 457
rect -6115 411 -6037 457
rect -5991 411 -5913 457
rect -5867 411 -5789 457
rect -5743 411 -5665 457
rect -5619 411 -5541 457
rect -5495 411 -5417 457
rect -5371 411 -5293 457
rect -5247 411 -5169 457
rect -5123 411 -5045 457
rect -4999 411 -4921 457
rect -4875 411 -4797 457
rect -4751 411 -4673 457
rect -4627 411 -4549 457
rect -4503 411 -4425 457
rect -4379 411 -4301 457
rect -4255 411 -4177 457
rect -4131 411 -4053 457
rect -4007 411 -3929 457
rect -3883 411 -3805 457
rect -3759 411 -3681 457
rect -3635 411 -3557 457
rect -3511 411 -3433 457
rect -3387 411 -3309 457
rect -3263 411 -3185 457
rect -3139 411 -3061 457
rect -3015 411 -2937 457
rect -2891 411 -2813 457
rect -2767 411 -2689 457
rect -2643 411 -2565 457
rect -2519 411 -2441 457
rect -2395 411 -2317 457
rect -2271 411 -2193 457
rect -2147 411 -2069 457
rect -2023 411 -1945 457
rect -1899 411 -1821 457
rect -1775 411 -1697 457
rect -1651 411 -1573 457
rect -1527 411 -1449 457
rect -1403 411 -1325 457
rect -1279 411 -1201 457
rect -1155 411 -1077 457
rect -1031 411 -953 457
rect -907 411 -829 457
rect -783 411 -705 457
rect -659 411 -581 457
rect -535 411 -457 457
rect -411 411 -333 457
rect -287 411 -209 457
rect -163 411 -85 457
rect -39 411 39 457
rect 85 411 163 457
rect 209 411 287 457
rect 333 411 411 457
rect 457 411 535 457
rect 581 411 659 457
rect 705 411 783 457
rect 829 411 907 457
rect 953 411 1031 457
rect 1077 411 1155 457
rect 1201 411 1279 457
rect 1325 411 1403 457
rect 1449 411 1527 457
rect 1573 411 1651 457
rect 1697 411 1775 457
rect 1821 411 1899 457
rect 1945 411 2023 457
rect 2069 411 2147 457
rect 2193 411 2271 457
rect 2317 411 2395 457
rect 2441 411 2519 457
rect 2565 411 2643 457
rect 2689 411 2767 457
rect 2813 411 2891 457
rect 2937 411 3015 457
rect 3061 411 3139 457
rect 3185 411 3263 457
rect 3309 411 3387 457
rect 3433 411 3511 457
rect 3557 411 3635 457
rect 3681 411 3759 457
rect 3805 411 3883 457
rect 3929 411 4007 457
rect 4053 411 4131 457
rect 4177 411 4255 457
rect 4301 411 4379 457
rect 4425 411 4503 457
rect 4549 411 4627 457
rect 4673 411 4751 457
rect 4797 411 4875 457
rect 4921 411 4999 457
rect 5045 411 5123 457
rect 5169 411 5247 457
rect 5293 411 5371 457
rect 5417 411 5495 457
rect 5541 411 5619 457
rect 5665 411 5743 457
rect 5789 411 5867 457
rect 5913 411 5991 457
rect 6037 411 6115 457
rect 6161 411 6239 457
rect 6285 411 6363 457
rect 6409 411 6487 457
rect 6533 411 6611 457
rect 6657 411 6735 457
rect 6781 411 6859 457
rect 6905 411 6983 457
rect 7029 411 7107 457
rect 7153 411 7231 457
rect 7277 411 7355 457
rect 7401 411 7479 457
rect 7525 411 7603 457
rect 7649 411 7727 457
rect 7773 411 7851 457
rect 7897 411 7975 457
rect 8021 411 8099 457
rect 8145 411 8223 457
rect 8269 411 8347 457
rect 8393 411 8471 457
rect 8517 411 8595 457
rect 8641 411 8719 457
rect 8765 411 8843 457
rect 8889 411 8967 457
rect 9013 411 9091 457
rect 9137 411 9215 457
rect 9261 411 9339 457
rect 9385 411 9463 457
rect 9509 411 9587 457
rect 9633 411 9711 457
rect 9757 411 9835 457
rect 9881 411 9959 457
rect 10005 411 10083 457
rect 10129 411 10207 457
rect 10253 411 10331 457
rect 10377 411 10455 457
rect 10501 411 10579 457
rect 10625 411 10703 457
rect 10749 411 10827 457
rect 10873 411 10951 457
rect 10997 411 11075 457
rect 11121 411 11199 457
rect 11245 411 11323 457
rect 11369 411 11447 457
rect 11493 411 11571 457
rect 11617 411 11695 457
rect 11741 411 11819 457
rect 11865 411 11943 457
rect 11989 411 12067 457
rect 12113 411 12191 457
rect 12237 411 12315 457
rect 12361 411 12439 457
rect 12485 411 12563 457
rect 12609 411 12687 457
rect 12733 411 12811 457
rect 12857 411 12935 457
rect 12981 411 13059 457
rect 13105 411 13183 457
rect 13229 411 13307 457
rect 13353 411 13431 457
rect 13477 411 13555 457
rect 13601 411 13679 457
rect 13725 411 13803 457
rect 13849 411 13927 457
rect 13973 411 14051 457
rect 14097 411 14175 457
rect 14221 411 14299 457
rect 14345 411 14423 457
rect 14469 411 14547 457
rect 14593 411 14671 457
rect 14717 411 14795 457
rect 14841 411 14919 457
rect 14965 411 15043 457
rect 15089 411 15167 457
rect 15213 411 15291 457
rect 15337 411 15415 457
rect 15461 411 15539 457
rect 15585 411 15663 457
rect 15709 411 15787 457
rect 15833 411 15911 457
rect 15957 411 16035 457
rect 16081 411 16159 457
rect 16205 411 16283 457
rect 16329 411 16407 457
rect 16453 411 16531 457
rect 16577 411 16655 457
rect 16701 411 16779 457
rect 16825 411 16903 457
rect 16949 411 17027 457
rect 17073 411 17151 457
rect 17197 411 17275 457
rect 17321 411 17343 457
rect -17343 333 17343 411
rect -17343 287 -17321 333
rect -17275 287 -17197 333
rect -17151 287 -17073 333
rect -17027 287 -16949 333
rect -16903 287 -16825 333
rect -16779 287 -16701 333
rect -16655 287 -16577 333
rect -16531 287 -16453 333
rect -16407 287 -16329 333
rect -16283 287 -16205 333
rect -16159 287 -16081 333
rect -16035 287 -15957 333
rect -15911 287 -15833 333
rect -15787 287 -15709 333
rect -15663 287 -15585 333
rect -15539 287 -15461 333
rect -15415 287 -15337 333
rect -15291 287 -15213 333
rect -15167 287 -15089 333
rect -15043 287 -14965 333
rect -14919 287 -14841 333
rect -14795 287 -14717 333
rect -14671 287 -14593 333
rect -14547 287 -14469 333
rect -14423 287 -14345 333
rect -14299 287 -14221 333
rect -14175 287 -14097 333
rect -14051 287 -13973 333
rect -13927 287 -13849 333
rect -13803 287 -13725 333
rect -13679 287 -13601 333
rect -13555 287 -13477 333
rect -13431 287 -13353 333
rect -13307 287 -13229 333
rect -13183 287 -13105 333
rect -13059 287 -12981 333
rect -12935 287 -12857 333
rect -12811 287 -12733 333
rect -12687 287 -12609 333
rect -12563 287 -12485 333
rect -12439 287 -12361 333
rect -12315 287 -12237 333
rect -12191 287 -12113 333
rect -12067 287 -11989 333
rect -11943 287 -11865 333
rect -11819 287 -11741 333
rect -11695 287 -11617 333
rect -11571 287 -11493 333
rect -11447 287 -11369 333
rect -11323 287 -11245 333
rect -11199 287 -11121 333
rect -11075 287 -10997 333
rect -10951 287 -10873 333
rect -10827 287 -10749 333
rect -10703 287 -10625 333
rect -10579 287 -10501 333
rect -10455 287 -10377 333
rect -10331 287 -10253 333
rect -10207 287 -10129 333
rect -10083 287 -10005 333
rect -9959 287 -9881 333
rect -9835 287 -9757 333
rect -9711 287 -9633 333
rect -9587 287 -9509 333
rect -9463 287 -9385 333
rect -9339 287 -9261 333
rect -9215 287 -9137 333
rect -9091 287 -9013 333
rect -8967 287 -8889 333
rect -8843 287 -8765 333
rect -8719 287 -8641 333
rect -8595 287 -8517 333
rect -8471 287 -8393 333
rect -8347 287 -8269 333
rect -8223 287 -8145 333
rect -8099 287 -8021 333
rect -7975 287 -7897 333
rect -7851 287 -7773 333
rect -7727 287 -7649 333
rect -7603 287 -7525 333
rect -7479 287 -7401 333
rect -7355 287 -7277 333
rect -7231 287 -7153 333
rect -7107 287 -7029 333
rect -6983 287 -6905 333
rect -6859 287 -6781 333
rect -6735 287 -6657 333
rect -6611 287 -6533 333
rect -6487 287 -6409 333
rect -6363 287 -6285 333
rect -6239 287 -6161 333
rect -6115 287 -6037 333
rect -5991 287 -5913 333
rect -5867 287 -5789 333
rect -5743 287 -5665 333
rect -5619 287 -5541 333
rect -5495 287 -5417 333
rect -5371 287 -5293 333
rect -5247 287 -5169 333
rect -5123 287 -5045 333
rect -4999 287 -4921 333
rect -4875 287 -4797 333
rect -4751 287 -4673 333
rect -4627 287 -4549 333
rect -4503 287 -4425 333
rect -4379 287 -4301 333
rect -4255 287 -4177 333
rect -4131 287 -4053 333
rect -4007 287 -3929 333
rect -3883 287 -3805 333
rect -3759 287 -3681 333
rect -3635 287 -3557 333
rect -3511 287 -3433 333
rect -3387 287 -3309 333
rect -3263 287 -3185 333
rect -3139 287 -3061 333
rect -3015 287 -2937 333
rect -2891 287 -2813 333
rect -2767 287 -2689 333
rect -2643 287 -2565 333
rect -2519 287 -2441 333
rect -2395 287 -2317 333
rect -2271 287 -2193 333
rect -2147 287 -2069 333
rect -2023 287 -1945 333
rect -1899 287 -1821 333
rect -1775 287 -1697 333
rect -1651 287 -1573 333
rect -1527 287 -1449 333
rect -1403 287 -1325 333
rect -1279 287 -1201 333
rect -1155 287 -1077 333
rect -1031 287 -953 333
rect -907 287 -829 333
rect -783 287 -705 333
rect -659 287 -581 333
rect -535 287 -457 333
rect -411 287 -333 333
rect -287 287 -209 333
rect -163 287 -85 333
rect -39 287 39 333
rect 85 287 163 333
rect 209 287 287 333
rect 333 287 411 333
rect 457 287 535 333
rect 581 287 659 333
rect 705 287 783 333
rect 829 287 907 333
rect 953 287 1031 333
rect 1077 287 1155 333
rect 1201 287 1279 333
rect 1325 287 1403 333
rect 1449 287 1527 333
rect 1573 287 1651 333
rect 1697 287 1775 333
rect 1821 287 1899 333
rect 1945 287 2023 333
rect 2069 287 2147 333
rect 2193 287 2271 333
rect 2317 287 2395 333
rect 2441 287 2519 333
rect 2565 287 2643 333
rect 2689 287 2767 333
rect 2813 287 2891 333
rect 2937 287 3015 333
rect 3061 287 3139 333
rect 3185 287 3263 333
rect 3309 287 3387 333
rect 3433 287 3511 333
rect 3557 287 3635 333
rect 3681 287 3759 333
rect 3805 287 3883 333
rect 3929 287 4007 333
rect 4053 287 4131 333
rect 4177 287 4255 333
rect 4301 287 4379 333
rect 4425 287 4503 333
rect 4549 287 4627 333
rect 4673 287 4751 333
rect 4797 287 4875 333
rect 4921 287 4999 333
rect 5045 287 5123 333
rect 5169 287 5247 333
rect 5293 287 5371 333
rect 5417 287 5495 333
rect 5541 287 5619 333
rect 5665 287 5743 333
rect 5789 287 5867 333
rect 5913 287 5991 333
rect 6037 287 6115 333
rect 6161 287 6239 333
rect 6285 287 6363 333
rect 6409 287 6487 333
rect 6533 287 6611 333
rect 6657 287 6735 333
rect 6781 287 6859 333
rect 6905 287 6983 333
rect 7029 287 7107 333
rect 7153 287 7231 333
rect 7277 287 7355 333
rect 7401 287 7479 333
rect 7525 287 7603 333
rect 7649 287 7727 333
rect 7773 287 7851 333
rect 7897 287 7975 333
rect 8021 287 8099 333
rect 8145 287 8223 333
rect 8269 287 8347 333
rect 8393 287 8471 333
rect 8517 287 8595 333
rect 8641 287 8719 333
rect 8765 287 8843 333
rect 8889 287 8967 333
rect 9013 287 9091 333
rect 9137 287 9215 333
rect 9261 287 9339 333
rect 9385 287 9463 333
rect 9509 287 9587 333
rect 9633 287 9711 333
rect 9757 287 9835 333
rect 9881 287 9959 333
rect 10005 287 10083 333
rect 10129 287 10207 333
rect 10253 287 10331 333
rect 10377 287 10455 333
rect 10501 287 10579 333
rect 10625 287 10703 333
rect 10749 287 10827 333
rect 10873 287 10951 333
rect 10997 287 11075 333
rect 11121 287 11199 333
rect 11245 287 11323 333
rect 11369 287 11447 333
rect 11493 287 11571 333
rect 11617 287 11695 333
rect 11741 287 11819 333
rect 11865 287 11943 333
rect 11989 287 12067 333
rect 12113 287 12191 333
rect 12237 287 12315 333
rect 12361 287 12439 333
rect 12485 287 12563 333
rect 12609 287 12687 333
rect 12733 287 12811 333
rect 12857 287 12935 333
rect 12981 287 13059 333
rect 13105 287 13183 333
rect 13229 287 13307 333
rect 13353 287 13431 333
rect 13477 287 13555 333
rect 13601 287 13679 333
rect 13725 287 13803 333
rect 13849 287 13927 333
rect 13973 287 14051 333
rect 14097 287 14175 333
rect 14221 287 14299 333
rect 14345 287 14423 333
rect 14469 287 14547 333
rect 14593 287 14671 333
rect 14717 287 14795 333
rect 14841 287 14919 333
rect 14965 287 15043 333
rect 15089 287 15167 333
rect 15213 287 15291 333
rect 15337 287 15415 333
rect 15461 287 15539 333
rect 15585 287 15663 333
rect 15709 287 15787 333
rect 15833 287 15911 333
rect 15957 287 16035 333
rect 16081 287 16159 333
rect 16205 287 16283 333
rect 16329 287 16407 333
rect 16453 287 16531 333
rect 16577 287 16655 333
rect 16701 287 16779 333
rect 16825 287 16903 333
rect 16949 287 17027 333
rect 17073 287 17151 333
rect 17197 287 17275 333
rect 17321 287 17343 333
rect -17343 209 17343 287
rect -17343 163 -17321 209
rect -17275 163 -17197 209
rect -17151 163 -17073 209
rect -17027 163 -16949 209
rect -16903 163 -16825 209
rect -16779 163 -16701 209
rect -16655 163 -16577 209
rect -16531 163 -16453 209
rect -16407 163 -16329 209
rect -16283 163 -16205 209
rect -16159 163 -16081 209
rect -16035 163 -15957 209
rect -15911 163 -15833 209
rect -15787 163 -15709 209
rect -15663 163 -15585 209
rect -15539 163 -15461 209
rect -15415 163 -15337 209
rect -15291 163 -15213 209
rect -15167 163 -15089 209
rect -15043 163 -14965 209
rect -14919 163 -14841 209
rect -14795 163 -14717 209
rect -14671 163 -14593 209
rect -14547 163 -14469 209
rect -14423 163 -14345 209
rect -14299 163 -14221 209
rect -14175 163 -14097 209
rect -14051 163 -13973 209
rect -13927 163 -13849 209
rect -13803 163 -13725 209
rect -13679 163 -13601 209
rect -13555 163 -13477 209
rect -13431 163 -13353 209
rect -13307 163 -13229 209
rect -13183 163 -13105 209
rect -13059 163 -12981 209
rect -12935 163 -12857 209
rect -12811 163 -12733 209
rect -12687 163 -12609 209
rect -12563 163 -12485 209
rect -12439 163 -12361 209
rect -12315 163 -12237 209
rect -12191 163 -12113 209
rect -12067 163 -11989 209
rect -11943 163 -11865 209
rect -11819 163 -11741 209
rect -11695 163 -11617 209
rect -11571 163 -11493 209
rect -11447 163 -11369 209
rect -11323 163 -11245 209
rect -11199 163 -11121 209
rect -11075 163 -10997 209
rect -10951 163 -10873 209
rect -10827 163 -10749 209
rect -10703 163 -10625 209
rect -10579 163 -10501 209
rect -10455 163 -10377 209
rect -10331 163 -10253 209
rect -10207 163 -10129 209
rect -10083 163 -10005 209
rect -9959 163 -9881 209
rect -9835 163 -9757 209
rect -9711 163 -9633 209
rect -9587 163 -9509 209
rect -9463 163 -9385 209
rect -9339 163 -9261 209
rect -9215 163 -9137 209
rect -9091 163 -9013 209
rect -8967 163 -8889 209
rect -8843 163 -8765 209
rect -8719 163 -8641 209
rect -8595 163 -8517 209
rect -8471 163 -8393 209
rect -8347 163 -8269 209
rect -8223 163 -8145 209
rect -8099 163 -8021 209
rect -7975 163 -7897 209
rect -7851 163 -7773 209
rect -7727 163 -7649 209
rect -7603 163 -7525 209
rect -7479 163 -7401 209
rect -7355 163 -7277 209
rect -7231 163 -7153 209
rect -7107 163 -7029 209
rect -6983 163 -6905 209
rect -6859 163 -6781 209
rect -6735 163 -6657 209
rect -6611 163 -6533 209
rect -6487 163 -6409 209
rect -6363 163 -6285 209
rect -6239 163 -6161 209
rect -6115 163 -6037 209
rect -5991 163 -5913 209
rect -5867 163 -5789 209
rect -5743 163 -5665 209
rect -5619 163 -5541 209
rect -5495 163 -5417 209
rect -5371 163 -5293 209
rect -5247 163 -5169 209
rect -5123 163 -5045 209
rect -4999 163 -4921 209
rect -4875 163 -4797 209
rect -4751 163 -4673 209
rect -4627 163 -4549 209
rect -4503 163 -4425 209
rect -4379 163 -4301 209
rect -4255 163 -4177 209
rect -4131 163 -4053 209
rect -4007 163 -3929 209
rect -3883 163 -3805 209
rect -3759 163 -3681 209
rect -3635 163 -3557 209
rect -3511 163 -3433 209
rect -3387 163 -3309 209
rect -3263 163 -3185 209
rect -3139 163 -3061 209
rect -3015 163 -2937 209
rect -2891 163 -2813 209
rect -2767 163 -2689 209
rect -2643 163 -2565 209
rect -2519 163 -2441 209
rect -2395 163 -2317 209
rect -2271 163 -2193 209
rect -2147 163 -2069 209
rect -2023 163 -1945 209
rect -1899 163 -1821 209
rect -1775 163 -1697 209
rect -1651 163 -1573 209
rect -1527 163 -1449 209
rect -1403 163 -1325 209
rect -1279 163 -1201 209
rect -1155 163 -1077 209
rect -1031 163 -953 209
rect -907 163 -829 209
rect -783 163 -705 209
rect -659 163 -581 209
rect -535 163 -457 209
rect -411 163 -333 209
rect -287 163 -209 209
rect -163 163 -85 209
rect -39 163 39 209
rect 85 163 163 209
rect 209 163 287 209
rect 333 163 411 209
rect 457 163 535 209
rect 581 163 659 209
rect 705 163 783 209
rect 829 163 907 209
rect 953 163 1031 209
rect 1077 163 1155 209
rect 1201 163 1279 209
rect 1325 163 1403 209
rect 1449 163 1527 209
rect 1573 163 1651 209
rect 1697 163 1775 209
rect 1821 163 1899 209
rect 1945 163 2023 209
rect 2069 163 2147 209
rect 2193 163 2271 209
rect 2317 163 2395 209
rect 2441 163 2519 209
rect 2565 163 2643 209
rect 2689 163 2767 209
rect 2813 163 2891 209
rect 2937 163 3015 209
rect 3061 163 3139 209
rect 3185 163 3263 209
rect 3309 163 3387 209
rect 3433 163 3511 209
rect 3557 163 3635 209
rect 3681 163 3759 209
rect 3805 163 3883 209
rect 3929 163 4007 209
rect 4053 163 4131 209
rect 4177 163 4255 209
rect 4301 163 4379 209
rect 4425 163 4503 209
rect 4549 163 4627 209
rect 4673 163 4751 209
rect 4797 163 4875 209
rect 4921 163 4999 209
rect 5045 163 5123 209
rect 5169 163 5247 209
rect 5293 163 5371 209
rect 5417 163 5495 209
rect 5541 163 5619 209
rect 5665 163 5743 209
rect 5789 163 5867 209
rect 5913 163 5991 209
rect 6037 163 6115 209
rect 6161 163 6239 209
rect 6285 163 6363 209
rect 6409 163 6487 209
rect 6533 163 6611 209
rect 6657 163 6735 209
rect 6781 163 6859 209
rect 6905 163 6983 209
rect 7029 163 7107 209
rect 7153 163 7231 209
rect 7277 163 7355 209
rect 7401 163 7479 209
rect 7525 163 7603 209
rect 7649 163 7727 209
rect 7773 163 7851 209
rect 7897 163 7975 209
rect 8021 163 8099 209
rect 8145 163 8223 209
rect 8269 163 8347 209
rect 8393 163 8471 209
rect 8517 163 8595 209
rect 8641 163 8719 209
rect 8765 163 8843 209
rect 8889 163 8967 209
rect 9013 163 9091 209
rect 9137 163 9215 209
rect 9261 163 9339 209
rect 9385 163 9463 209
rect 9509 163 9587 209
rect 9633 163 9711 209
rect 9757 163 9835 209
rect 9881 163 9959 209
rect 10005 163 10083 209
rect 10129 163 10207 209
rect 10253 163 10331 209
rect 10377 163 10455 209
rect 10501 163 10579 209
rect 10625 163 10703 209
rect 10749 163 10827 209
rect 10873 163 10951 209
rect 10997 163 11075 209
rect 11121 163 11199 209
rect 11245 163 11323 209
rect 11369 163 11447 209
rect 11493 163 11571 209
rect 11617 163 11695 209
rect 11741 163 11819 209
rect 11865 163 11943 209
rect 11989 163 12067 209
rect 12113 163 12191 209
rect 12237 163 12315 209
rect 12361 163 12439 209
rect 12485 163 12563 209
rect 12609 163 12687 209
rect 12733 163 12811 209
rect 12857 163 12935 209
rect 12981 163 13059 209
rect 13105 163 13183 209
rect 13229 163 13307 209
rect 13353 163 13431 209
rect 13477 163 13555 209
rect 13601 163 13679 209
rect 13725 163 13803 209
rect 13849 163 13927 209
rect 13973 163 14051 209
rect 14097 163 14175 209
rect 14221 163 14299 209
rect 14345 163 14423 209
rect 14469 163 14547 209
rect 14593 163 14671 209
rect 14717 163 14795 209
rect 14841 163 14919 209
rect 14965 163 15043 209
rect 15089 163 15167 209
rect 15213 163 15291 209
rect 15337 163 15415 209
rect 15461 163 15539 209
rect 15585 163 15663 209
rect 15709 163 15787 209
rect 15833 163 15911 209
rect 15957 163 16035 209
rect 16081 163 16159 209
rect 16205 163 16283 209
rect 16329 163 16407 209
rect 16453 163 16531 209
rect 16577 163 16655 209
rect 16701 163 16779 209
rect 16825 163 16903 209
rect 16949 163 17027 209
rect 17073 163 17151 209
rect 17197 163 17275 209
rect 17321 163 17343 209
rect -17343 85 17343 163
rect -17343 39 -17321 85
rect -17275 39 -17197 85
rect -17151 39 -17073 85
rect -17027 39 -16949 85
rect -16903 39 -16825 85
rect -16779 39 -16701 85
rect -16655 39 -16577 85
rect -16531 39 -16453 85
rect -16407 39 -16329 85
rect -16283 39 -16205 85
rect -16159 39 -16081 85
rect -16035 39 -15957 85
rect -15911 39 -15833 85
rect -15787 39 -15709 85
rect -15663 39 -15585 85
rect -15539 39 -15461 85
rect -15415 39 -15337 85
rect -15291 39 -15213 85
rect -15167 39 -15089 85
rect -15043 39 -14965 85
rect -14919 39 -14841 85
rect -14795 39 -14717 85
rect -14671 39 -14593 85
rect -14547 39 -14469 85
rect -14423 39 -14345 85
rect -14299 39 -14221 85
rect -14175 39 -14097 85
rect -14051 39 -13973 85
rect -13927 39 -13849 85
rect -13803 39 -13725 85
rect -13679 39 -13601 85
rect -13555 39 -13477 85
rect -13431 39 -13353 85
rect -13307 39 -13229 85
rect -13183 39 -13105 85
rect -13059 39 -12981 85
rect -12935 39 -12857 85
rect -12811 39 -12733 85
rect -12687 39 -12609 85
rect -12563 39 -12485 85
rect -12439 39 -12361 85
rect -12315 39 -12237 85
rect -12191 39 -12113 85
rect -12067 39 -11989 85
rect -11943 39 -11865 85
rect -11819 39 -11741 85
rect -11695 39 -11617 85
rect -11571 39 -11493 85
rect -11447 39 -11369 85
rect -11323 39 -11245 85
rect -11199 39 -11121 85
rect -11075 39 -10997 85
rect -10951 39 -10873 85
rect -10827 39 -10749 85
rect -10703 39 -10625 85
rect -10579 39 -10501 85
rect -10455 39 -10377 85
rect -10331 39 -10253 85
rect -10207 39 -10129 85
rect -10083 39 -10005 85
rect -9959 39 -9881 85
rect -9835 39 -9757 85
rect -9711 39 -9633 85
rect -9587 39 -9509 85
rect -9463 39 -9385 85
rect -9339 39 -9261 85
rect -9215 39 -9137 85
rect -9091 39 -9013 85
rect -8967 39 -8889 85
rect -8843 39 -8765 85
rect -8719 39 -8641 85
rect -8595 39 -8517 85
rect -8471 39 -8393 85
rect -8347 39 -8269 85
rect -8223 39 -8145 85
rect -8099 39 -8021 85
rect -7975 39 -7897 85
rect -7851 39 -7773 85
rect -7727 39 -7649 85
rect -7603 39 -7525 85
rect -7479 39 -7401 85
rect -7355 39 -7277 85
rect -7231 39 -7153 85
rect -7107 39 -7029 85
rect -6983 39 -6905 85
rect -6859 39 -6781 85
rect -6735 39 -6657 85
rect -6611 39 -6533 85
rect -6487 39 -6409 85
rect -6363 39 -6285 85
rect -6239 39 -6161 85
rect -6115 39 -6037 85
rect -5991 39 -5913 85
rect -5867 39 -5789 85
rect -5743 39 -5665 85
rect -5619 39 -5541 85
rect -5495 39 -5417 85
rect -5371 39 -5293 85
rect -5247 39 -5169 85
rect -5123 39 -5045 85
rect -4999 39 -4921 85
rect -4875 39 -4797 85
rect -4751 39 -4673 85
rect -4627 39 -4549 85
rect -4503 39 -4425 85
rect -4379 39 -4301 85
rect -4255 39 -4177 85
rect -4131 39 -4053 85
rect -4007 39 -3929 85
rect -3883 39 -3805 85
rect -3759 39 -3681 85
rect -3635 39 -3557 85
rect -3511 39 -3433 85
rect -3387 39 -3309 85
rect -3263 39 -3185 85
rect -3139 39 -3061 85
rect -3015 39 -2937 85
rect -2891 39 -2813 85
rect -2767 39 -2689 85
rect -2643 39 -2565 85
rect -2519 39 -2441 85
rect -2395 39 -2317 85
rect -2271 39 -2193 85
rect -2147 39 -2069 85
rect -2023 39 -1945 85
rect -1899 39 -1821 85
rect -1775 39 -1697 85
rect -1651 39 -1573 85
rect -1527 39 -1449 85
rect -1403 39 -1325 85
rect -1279 39 -1201 85
rect -1155 39 -1077 85
rect -1031 39 -953 85
rect -907 39 -829 85
rect -783 39 -705 85
rect -659 39 -581 85
rect -535 39 -457 85
rect -411 39 -333 85
rect -287 39 -209 85
rect -163 39 -85 85
rect -39 39 39 85
rect 85 39 163 85
rect 209 39 287 85
rect 333 39 411 85
rect 457 39 535 85
rect 581 39 659 85
rect 705 39 783 85
rect 829 39 907 85
rect 953 39 1031 85
rect 1077 39 1155 85
rect 1201 39 1279 85
rect 1325 39 1403 85
rect 1449 39 1527 85
rect 1573 39 1651 85
rect 1697 39 1775 85
rect 1821 39 1899 85
rect 1945 39 2023 85
rect 2069 39 2147 85
rect 2193 39 2271 85
rect 2317 39 2395 85
rect 2441 39 2519 85
rect 2565 39 2643 85
rect 2689 39 2767 85
rect 2813 39 2891 85
rect 2937 39 3015 85
rect 3061 39 3139 85
rect 3185 39 3263 85
rect 3309 39 3387 85
rect 3433 39 3511 85
rect 3557 39 3635 85
rect 3681 39 3759 85
rect 3805 39 3883 85
rect 3929 39 4007 85
rect 4053 39 4131 85
rect 4177 39 4255 85
rect 4301 39 4379 85
rect 4425 39 4503 85
rect 4549 39 4627 85
rect 4673 39 4751 85
rect 4797 39 4875 85
rect 4921 39 4999 85
rect 5045 39 5123 85
rect 5169 39 5247 85
rect 5293 39 5371 85
rect 5417 39 5495 85
rect 5541 39 5619 85
rect 5665 39 5743 85
rect 5789 39 5867 85
rect 5913 39 5991 85
rect 6037 39 6115 85
rect 6161 39 6239 85
rect 6285 39 6363 85
rect 6409 39 6487 85
rect 6533 39 6611 85
rect 6657 39 6735 85
rect 6781 39 6859 85
rect 6905 39 6983 85
rect 7029 39 7107 85
rect 7153 39 7231 85
rect 7277 39 7355 85
rect 7401 39 7479 85
rect 7525 39 7603 85
rect 7649 39 7727 85
rect 7773 39 7851 85
rect 7897 39 7975 85
rect 8021 39 8099 85
rect 8145 39 8223 85
rect 8269 39 8347 85
rect 8393 39 8471 85
rect 8517 39 8595 85
rect 8641 39 8719 85
rect 8765 39 8843 85
rect 8889 39 8967 85
rect 9013 39 9091 85
rect 9137 39 9215 85
rect 9261 39 9339 85
rect 9385 39 9463 85
rect 9509 39 9587 85
rect 9633 39 9711 85
rect 9757 39 9835 85
rect 9881 39 9959 85
rect 10005 39 10083 85
rect 10129 39 10207 85
rect 10253 39 10331 85
rect 10377 39 10455 85
rect 10501 39 10579 85
rect 10625 39 10703 85
rect 10749 39 10827 85
rect 10873 39 10951 85
rect 10997 39 11075 85
rect 11121 39 11199 85
rect 11245 39 11323 85
rect 11369 39 11447 85
rect 11493 39 11571 85
rect 11617 39 11695 85
rect 11741 39 11819 85
rect 11865 39 11943 85
rect 11989 39 12067 85
rect 12113 39 12191 85
rect 12237 39 12315 85
rect 12361 39 12439 85
rect 12485 39 12563 85
rect 12609 39 12687 85
rect 12733 39 12811 85
rect 12857 39 12935 85
rect 12981 39 13059 85
rect 13105 39 13183 85
rect 13229 39 13307 85
rect 13353 39 13431 85
rect 13477 39 13555 85
rect 13601 39 13679 85
rect 13725 39 13803 85
rect 13849 39 13927 85
rect 13973 39 14051 85
rect 14097 39 14175 85
rect 14221 39 14299 85
rect 14345 39 14423 85
rect 14469 39 14547 85
rect 14593 39 14671 85
rect 14717 39 14795 85
rect 14841 39 14919 85
rect 14965 39 15043 85
rect 15089 39 15167 85
rect 15213 39 15291 85
rect 15337 39 15415 85
rect 15461 39 15539 85
rect 15585 39 15663 85
rect 15709 39 15787 85
rect 15833 39 15911 85
rect 15957 39 16035 85
rect 16081 39 16159 85
rect 16205 39 16283 85
rect 16329 39 16407 85
rect 16453 39 16531 85
rect 16577 39 16655 85
rect 16701 39 16779 85
rect 16825 39 16903 85
rect 16949 39 17027 85
rect 17073 39 17151 85
rect 17197 39 17275 85
rect 17321 39 17343 85
rect -17343 -39 17343 39
rect -17343 -85 -17321 -39
rect -17275 -85 -17197 -39
rect -17151 -85 -17073 -39
rect -17027 -85 -16949 -39
rect -16903 -85 -16825 -39
rect -16779 -85 -16701 -39
rect -16655 -85 -16577 -39
rect -16531 -85 -16453 -39
rect -16407 -85 -16329 -39
rect -16283 -85 -16205 -39
rect -16159 -85 -16081 -39
rect -16035 -85 -15957 -39
rect -15911 -85 -15833 -39
rect -15787 -85 -15709 -39
rect -15663 -85 -15585 -39
rect -15539 -85 -15461 -39
rect -15415 -85 -15337 -39
rect -15291 -85 -15213 -39
rect -15167 -85 -15089 -39
rect -15043 -85 -14965 -39
rect -14919 -85 -14841 -39
rect -14795 -85 -14717 -39
rect -14671 -85 -14593 -39
rect -14547 -85 -14469 -39
rect -14423 -85 -14345 -39
rect -14299 -85 -14221 -39
rect -14175 -85 -14097 -39
rect -14051 -85 -13973 -39
rect -13927 -85 -13849 -39
rect -13803 -85 -13725 -39
rect -13679 -85 -13601 -39
rect -13555 -85 -13477 -39
rect -13431 -85 -13353 -39
rect -13307 -85 -13229 -39
rect -13183 -85 -13105 -39
rect -13059 -85 -12981 -39
rect -12935 -85 -12857 -39
rect -12811 -85 -12733 -39
rect -12687 -85 -12609 -39
rect -12563 -85 -12485 -39
rect -12439 -85 -12361 -39
rect -12315 -85 -12237 -39
rect -12191 -85 -12113 -39
rect -12067 -85 -11989 -39
rect -11943 -85 -11865 -39
rect -11819 -85 -11741 -39
rect -11695 -85 -11617 -39
rect -11571 -85 -11493 -39
rect -11447 -85 -11369 -39
rect -11323 -85 -11245 -39
rect -11199 -85 -11121 -39
rect -11075 -85 -10997 -39
rect -10951 -85 -10873 -39
rect -10827 -85 -10749 -39
rect -10703 -85 -10625 -39
rect -10579 -85 -10501 -39
rect -10455 -85 -10377 -39
rect -10331 -85 -10253 -39
rect -10207 -85 -10129 -39
rect -10083 -85 -10005 -39
rect -9959 -85 -9881 -39
rect -9835 -85 -9757 -39
rect -9711 -85 -9633 -39
rect -9587 -85 -9509 -39
rect -9463 -85 -9385 -39
rect -9339 -85 -9261 -39
rect -9215 -85 -9137 -39
rect -9091 -85 -9013 -39
rect -8967 -85 -8889 -39
rect -8843 -85 -8765 -39
rect -8719 -85 -8641 -39
rect -8595 -85 -8517 -39
rect -8471 -85 -8393 -39
rect -8347 -85 -8269 -39
rect -8223 -85 -8145 -39
rect -8099 -85 -8021 -39
rect -7975 -85 -7897 -39
rect -7851 -85 -7773 -39
rect -7727 -85 -7649 -39
rect -7603 -85 -7525 -39
rect -7479 -85 -7401 -39
rect -7355 -85 -7277 -39
rect -7231 -85 -7153 -39
rect -7107 -85 -7029 -39
rect -6983 -85 -6905 -39
rect -6859 -85 -6781 -39
rect -6735 -85 -6657 -39
rect -6611 -85 -6533 -39
rect -6487 -85 -6409 -39
rect -6363 -85 -6285 -39
rect -6239 -85 -6161 -39
rect -6115 -85 -6037 -39
rect -5991 -85 -5913 -39
rect -5867 -85 -5789 -39
rect -5743 -85 -5665 -39
rect -5619 -85 -5541 -39
rect -5495 -85 -5417 -39
rect -5371 -85 -5293 -39
rect -5247 -85 -5169 -39
rect -5123 -85 -5045 -39
rect -4999 -85 -4921 -39
rect -4875 -85 -4797 -39
rect -4751 -85 -4673 -39
rect -4627 -85 -4549 -39
rect -4503 -85 -4425 -39
rect -4379 -85 -4301 -39
rect -4255 -85 -4177 -39
rect -4131 -85 -4053 -39
rect -4007 -85 -3929 -39
rect -3883 -85 -3805 -39
rect -3759 -85 -3681 -39
rect -3635 -85 -3557 -39
rect -3511 -85 -3433 -39
rect -3387 -85 -3309 -39
rect -3263 -85 -3185 -39
rect -3139 -85 -3061 -39
rect -3015 -85 -2937 -39
rect -2891 -85 -2813 -39
rect -2767 -85 -2689 -39
rect -2643 -85 -2565 -39
rect -2519 -85 -2441 -39
rect -2395 -85 -2317 -39
rect -2271 -85 -2193 -39
rect -2147 -85 -2069 -39
rect -2023 -85 -1945 -39
rect -1899 -85 -1821 -39
rect -1775 -85 -1697 -39
rect -1651 -85 -1573 -39
rect -1527 -85 -1449 -39
rect -1403 -85 -1325 -39
rect -1279 -85 -1201 -39
rect -1155 -85 -1077 -39
rect -1031 -85 -953 -39
rect -907 -85 -829 -39
rect -783 -85 -705 -39
rect -659 -85 -581 -39
rect -535 -85 -457 -39
rect -411 -85 -333 -39
rect -287 -85 -209 -39
rect -163 -85 -85 -39
rect -39 -85 39 -39
rect 85 -85 163 -39
rect 209 -85 287 -39
rect 333 -85 411 -39
rect 457 -85 535 -39
rect 581 -85 659 -39
rect 705 -85 783 -39
rect 829 -85 907 -39
rect 953 -85 1031 -39
rect 1077 -85 1155 -39
rect 1201 -85 1279 -39
rect 1325 -85 1403 -39
rect 1449 -85 1527 -39
rect 1573 -85 1651 -39
rect 1697 -85 1775 -39
rect 1821 -85 1899 -39
rect 1945 -85 2023 -39
rect 2069 -85 2147 -39
rect 2193 -85 2271 -39
rect 2317 -85 2395 -39
rect 2441 -85 2519 -39
rect 2565 -85 2643 -39
rect 2689 -85 2767 -39
rect 2813 -85 2891 -39
rect 2937 -85 3015 -39
rect 3061 -85 3139 -39
rect 3185 -85 3263 -39
rect 3309 -85 3387 -39
rect 3433 -85 3511 -39
rect 3557 -85 3635 -39
rect 3681 -85 3759 -39
rect 3805 -85 3883 -39
rect 3929 -85 4007 -39
rect 4053 -85 4131 -39
rect 4177 -85 4255 -39
rect 4301 -85 4379 -39
rect 4425 -85 4503 -39
rect 4549 -85 4627 -39
rect 4673 -85 4751 -39
rect 4797 -85 4875 -39
rect 4921 -85 4999 -39
rect 5045 -85 5123 -39
rect 5169 -85 5247 -39
rect 5293 -85 5371 -39
rect 5417 -85 5495 -39
rect 5541 -85 5619 -39
rect 5665 -85 5743 -39
rect 5789 -85 5867 -39
rect 5913 -85 5991 -39
rect 6037 -85 6115 -39
rect 6161 -85 6239 -39
rect 6285 -85 6363 -39
rect 6409 -85 6487 -39
rect 6533 -85 6611 -39
rect 6657 -85 6735 -39
rect 6781 -85 6859 -39
rect 6905 -85 6983 -39
rect 7029 -85 7107 -39
rect 7153 -85 7231 -39
rect 7277 -85 7355 -39
rect 7401 -85 7479 -39
rect 7525 -85 7603 -39
rect 7649 -85 7727 -39
rect 7773 -85 7851 -39
rect 7897 -85 7975 -39
rect 8021 -85 8099 -39
rect 8145 -85 8223 -39
rect 8269 -85 8347 -39
rect 8393 -85 8471 -39
rect 8517 -85 8595 -39
rect 8641 -85 8719 -39
rect 8765 -85 8843 -39
rect 8889 -85 8967 -39
rect 9013 -85 9091 -39
rect 9137 -85 9215 -39
rect 9261 -85 9339 -39
rect 9385 -85 9463 -39
rect 9509 -85 9587 -39
rect 9633 -85 9711 -39
rect 9757 -85 9835 -39
rect 9881 -85 9959 -39
rect 10005 -85 10083 -39
rect 10129 -85 10207 -39
rect 10253 -85 10331 -39
rect 10377 -85 10455 -39
rect 10501 -85 10579 -39
rect 10625 -85 10703 -39
rect 10749 -85 10827 -39
rect 10873 -85 10951 -39
rect 10997 -85 11075 -39
rect 11121 -85 11199 -39
rect 11245 -85 11323 -39
rect 11369 -85 11447 -39
rect 11493 -85 11571 -39
rect 11617 -85 11695 -39
rect 11741 -85 11819 -39
rect 11865 -85 11943 -39
rect 11989 -85 12067 -39
rect 12113 -85 12191 -39
rect 12237 -85 12315 -39
rect 12361 -85 12439 -39
rect 12485 -85 12563 -39
rect 12609 -85 12687 -39
rect 12733 -85 12811 -39
rect 12857 -85 12935 -39
rect 12981 -85 13059 -39
rect 13105 -85 13183 -39
rect 13229 -85 13307 -39
rect 13353 -85 13431 -39
rect 13477 -85 13555 -39
rect 13601 -85 13679 -39
rect 13725 -85 13803 -39
rect 13849 -85 13927 -39
rect 13973 -85 14051 -39
rect 14097 -85 14175 -39
rect 14221 -85 14299 -39
rect 14345 -85 14423 -39
rect 14469 -85 14547 -39
rect 14593 -85 14671 -39
rect 14717 -85 14795 -39
rect 14841 -85 14919 -39
rect 14965 -85 15043 -39
rect 15089 -85 15167 -39
rect 15213 -85 15291 -39
rect 15337 -85 15415 -39
rect 15461 -85 15539 -39
rect 15585 -85 15663 -39
rect 15709 -85 15787 -39
rect 15833 -85 15911 -39
rect 15957 -85 16035 -39
rect 16081 -85 16159 -39
rect 16205 -85 16283 -39
rect 16329 -85 16407 -39
rect 16453 -85 16531 -39
rect 16577 -85 16655 -39
rect 16701 -85 16779 -39
rect 16825 -85 16903 -39
rect 16949 -85 17027 -39
rect 17073 -85 17151 -39
rect 17197 -85 17275 -39
rect 17321 -85 17343 -39
rect -17343 -163 17343 -85
rect -17343 -209 -17321 -163
rect -17275 -209 -17197 -163
rect -17151 -209 -17073 -163
rect -17027 -209 -16949 -163
rect -16903 -209 -16825 -163
rect -16779 -209 -16701 -163
rect -16655 -209 -16577 -163
rect -16531 -209 -16453 -163
rect -16407 -209 -16329 -163
rect -16283 -209 -16205 -163
rect -16159 -209 -16081 -163
rect -16035 -209 -15957 -163
rect -15911 -209 -15833 -163
rect -15787 -209 -15709 -163
rect -15663 -209 -15585 -163
rect -15539 -209 -15461 -163
rect -15415 -209 -15337 -163
rect -15291 -209 -15213 -163
rect -15167 -209 -15089 -163
rect -15043 -209 -14965 -163
rect -14919 -209 -14841 -163
rect -14795 -209 -14717 -163
rect -14671 -209 -14593 -163
rect -14547 -209 -14469 -163
rect -14423 -209 -14345 -163
rect -14299 -209 -14221 -163
rect -14175 -209 -14097 -163
rect -14051 -209 -13973 -163
rect -13927 -209 -13849 -163
rect -13803 -209 -13725 -163
rect -13679 -209 -13601 -163
rect -13555 -209 -13477 -163
rect -13431 -209 -13353 -163
rect -13307 -209 -13229 -163
rect -13183 -209 -13105 -163
rect -13059 -209 -12981 -163
rect -12935 -209 -12857 -163
rect -12811 -209 -12733 -163
rect -12687 -209 -12609 -163
rect -12563 -209 -12485 -163
rect -12439 -209 -12361 -163
rect -12315 -209 -12237 -163
rect -12191 -209 -12113 -163
rect -12067 -209 -11989 -163
rect -11943 -209 -11865 -163
rect -11819 -209 -11741 -163
rect -11695 -209 -11617 -163
rect -11571 -209 -11493 -163
rect -11447 -209 -11369 -163
rect -11323 -209 -11245 -163
rect -11199 -209 -11121 -163
rect -11075 -209 -10997 -163
rect -10951 -209 -10873 -163
rect -10827 -209 -10749 -163
rect -10703 -209 -10625 -163
rect -10579 -209 -10501 -163
rect -10455 -209 -10377 -163
rect -10331 -209 -10253 -163
rect -10207 -209 -10129 -163
rect -10083 -209 -10005 -163
rect -9959 -209 -9881 -163
rect -9835 -209 -9757 -163
rect -9711 -209 -9633 -163
rect -9587 -209 -9509 -163
rect -9463 -209 -9385 -163
rect -9339 -209 -9261 -163
rect -9215 -209 -9137 -163
rect -9091 -209 -9013 -163
rect -8967 -209 -8889 -163
rect -8843 -209 -8765 -163
rect -8719 -209 -8641 -163
rect -8595 -209 -8517 -163
rect -8471 -209 -8393 -163
rect -8347 -209 -8269 -163
rect -8223 -209 -8145 -163
rect -8099 -209 -8021 -163
rect -7975 -209 -7897 -163
rect -7851 -209 -7773 -163
rect -7727 -209 -7649 -163
rect -7603 -209 -7525 -163
rect -7479 -209 -7401 -163
rect -7355 -209 -7277 -163
rect -7231 -209 -7153 -163
rect -7107 -209 -7029 -163
rect -6983 -209 -6905 -163
rect -6859 -209 -6781 -163
rect -6735 -209 -6657 -163
rect -6611 -209 -6533 -163
rect -6487 -209 -6409 -163
rect -6363 -209 -6285 -163
rect -6239 -209 -6161 -163
rect -6115 -209 -6037 -163
rect -5991 -209 -5913 -163
rect -5867 -209 -5789 -163
rect -5743 -209 -5665 -163
rect -5619 -209 -5541 -163
rect -5495 -209 -5417 -163
rect -5371 -209 -5293 -163
rect -5247 -209 -5169 -163
rect -5123 -209 -5045 -163
rect -4999 -209 -4921 -163
rect -4875 -209 -4797 -163
rect -4751 -209 -4673 -163
rect -4627 -209 -4549 -163
rect -4503 -209 -4425 -163
rect -4379 -209 -4301 -163
rect -4255 -209 -4177 -163
rect -4131 -209 -4053 -163
rect -4007 -209 -3929 -163
rect -3883 -209 -3805 -163
rect -3759 -209 -3681 -163
rect -3635 -209 -3557 -163
rect -3511 -209 -3433 -163
rect -3387 -209 -3309 -163
rect -3263 -209 -3185 -163
rect -3139 -209 -3061 -163
rect -3015 -209 -2937 -163
rect -2891 -209 -2813 -163
rect -2767 -209 -2689 -163
rect -2643 -209 -2565 -163
rect -2519 -209 -2441 -163
rect -2395 -209 -2317 -163
rect -2271 -209 -2193 -163
rect -2147 -209 -2069 -163
rect -2023 -209 -1945 -163
rect -1899 -209 -1821 -163
rect -1775 -209 -1697 -163
rect -1651 -209 -1573 -163
rect -1527 -209 -1449 -163
rect -1403 -209 -1325 -163
rect -1279 -209 -1201 -163
rect -1155 -209 -1077 -163
rect -1031 -209 -953 -163
rect -907 -209 -829 -163
rect -783 -209 -705 -163
rect -659 -209 -581 -163
rect -535 -209 -457 -163
rect -411 -209 -333 -163
rect -287 -209 -209 -163
rect -163 -209 -85 -163
rect -39 -209 39 -163
rect 85 -209 163 -163
rect 209 -209 287 -163
rect 333 -209 411 -163
rect 457 -209 535 -163
rect 581 -209 659 -163
rect 705 -209 783 -163
rect 829 -209 907 -163
rect 953 -209 1031 -163
rect 1077 -209 1155 -163
rect 1201 -209 1279 -163
rect 1325 -209 1403 -163
rect 1449 -209 1527 -163
rect 1573 -209 1651 -163
rect 1697 -209 1775 -163
rect 1821 -209 1899 -163
rect 1945 -209 2023 -163
rect 2069 -209 2147 -163
rect 2193 -209 2271 -163
rect 2317 -209 2395 -163
rect 2441 -209 2519 -163
rect 2565 -209 2643 -163
rect 2689 -209 2767 -163
rect 2813 -209 2891 -163
rect 2937 -209 3015 -163
rect 3061 -209 3139 -163
rect 3185 -209 3263 -163
rect 3309 -209 3387 -163
rect 3433 -209 3511 -163
rect 3557 -209 3635 -163
rect 3681 -209 3759 -163
rect 3805 -209 3883 -163
rect 3929 -209 4007 -163
rect 4053 -209 4131 -163
rect 4177 -209 4255 -163
rect 4301 -209 4379 -163
rect 4425 -209 4503 -163
rect 4549 -209 4627 -163
rect 4673 -209 4751 -163
rect 4797 -209 4875 -163
rect 4921 -209 4999 -163
rect 5045 -209 5123 -163
rect 5169 -209 5247 -163
rect 5293 -209 5371 -163
rect 5417 -209 5495 -163
rect 5541 -209 5619 -163
rect 5665 -209 5743 -163
rect 5789 -209 5867 -163
rect 5913 -209 5991 -163
rect 6037 -209 6115 -163
rect 6161 -209 6239 -163
rect 6285 -209 6363 -163
rect 6409 -209 6487 -163
rect 6533 -209 6611 -163
rect 6657 -209 6735 -163
rect 6781 -209 6859 -163
rect 6905 -209 6983 -163
rect 7029 -209 7107 -163
rect 7153 -209 7231 -163
rect 7277 -209 7355 -163
rect 7401 -209 7479 -163
rect 7525 -209 7603 -163
rect 7649 -209 7727 -163
rect 7773 -209 7851 -163
rect 7897 -209 7975 -163
rect 8021 -209 8099 -163
rect 8145 -209 8223 -163
rect 8269 -209 8347 -163
rect 8393 -209 8471 -163
rect 8517 -209 8595 -163
rect 8641 -209 8719 -163
rect 8765 -209 8843 -163
rect 8889 -209 8967 -163
rect 9013 -209 9091 -163
rect 9137 -209 9215 -163
rect 9261 -209 9339 -163
rect 9385 -209 9463 -163
rect 9509 -209 9587 -163
rect 9633 -209 9711 -163
rect 9757 -209 9835 -163
rect 9881 -209 9959 -163
rect 10005 -209 10083 -163
rect 10129 -209 10207 -163
rect 10253 -209 10331 -163
rect 10377 -209 10455 -163
rect 10501 -209 10579 -163
rect 10625 -209 10703 -163
rect 10749 -209 10827 -163
rect 10873 -209 10951 -163
rect 10997 -209 11075 -163
rect 11121 -209 11199 -163
rect 11245 -209 11323 -163
rect 11369 -209 11447 -163
rect 11493 -209 11571 -163
rect 11617 -209 11695 -163
rect 11741 -209 11819 -163
rect 11865 -209 11943 -163
rect 11989 -209 12067 -163
rect 12113 -209 12191 -163
rect 12237 -209 12315 -163
rect 12361 -209 12439 -163
rect 12485 -209 12563 -163
rect 12609 -209 12687 -163
rect 12733 -209 12811 -163
rect 12857 -209 12935 -163
rect 12981 -209 13059 -163
rect 13105 -209 13183 -163
rect 13229 -209 13307 -163
rect 13353 -209 13431 -163
rect 13477 -209 13555 -163
rect 13601 -209 13679 -163
rect 13725 -209 13803 -163
rect 13849 -209 13927 -163
rect 13973 -209 14051 -163
rect 14097 -209 14175 -163
rect 14221 -209 14299 -163
rect 14345 -209 14423 -163
rect 14469 -209 14547 -163
rect 14593 -209 14671 -163
rect 14717 -209 14795 -163
rect 14841 -209 14919 -163
rect 14965 -209 15043 -163
rect 15089 -209 15167 -163
rect 15213 -209 15291 -163
rect 15337 -209 15415 -163
rect 15461 -209 15539 -163
rect 15585 -209 15663 -163
rect 15709 -209 15787 -163
rect 15833 -209 15911 -163
rect 15957 -209 16035 -163
rect 16081 -209 16159 -163
rect 16205 -209 16283 -163
rect 16329 -209 16407 -163
rect 16453 -209 16531 -163
rect 16577 -209 16655 -163
rect 16701 -209 16779 -163
rect 16825 -209 16903 -163
rect 16949 -209 17027 -163
rect 17073 -209 17151 -163
rect 17197 -209 17275 -163
rect 17321 -209 17343 -163
rect -17343 -287 17343 -209
rect -17343 -333 -17321 -287
rect -17275 -333 -17197 -287
rect -17151 -333 -17073 -287
rect -17027 -333 -16949 -287
rect -16903 -333 -16825 -287
rect -16779 -333 -16701 -287
rect -16655 -333 -16577 -287
rect -16531 -333 -16453 -287
rect -16407 -333 -16329 -287
rect -16283 -333 -16205 -287
rect -16159 -333 -16081 -287
rect -16035 -333 -15957 -287
rect -15911 -333 -15833 -287
rect -15787 -333 -15709 -287
rect -15663 -333 -15585 -287
rect -15539 -333 -15461 -287
rect -15415 -333 -15337 -287
rect -15291 -333 -15213 -287
rect -15167 -333 -15089 -287
rect -15043 -333 -14965 -287
rect -14919 -333 -14841 -287
rect -14795 -333 -14717 -287
rect -14671 -333 -14593 -287
rect -14547 -333 -14469 -287
rect -14423 -333 -14345 -287
rect -14299 -333 -14221 -287
rect -14175 -333 -14097 -287
rect -14051 -333 -13973 -287
rect -13927 -333 -13849 -287
rect -13803 -333 -13725 -287
rect -13679 -333 -13601 -287
rect -13555 -333 -13477 -287
rect -13431 -333 -13353 -287
rect -13307 -333 -13229 -287
rect -13183 -333 -13105 -287
rect -13059 -333 -12981 -287
rect -12935 -333 -12857 -287
rect -12811 -333 -12733 -287
rect -12687 -333 -12609 -287
rect -12563 -333 -12485 -287
rect -12439 -333 -12361 -287
rect -12315 -333 -12237 -287
rect -12191 -333 -12113 -287
rect -12067 -333 -11989 -287
rect -11943 -333 -11865 -287
rect -11819 -333 -11741 -287
rect -11695 -333 -11617 -287
rect -11571 -333 -11493 -287
rect -11447 -333 -11369 -287
rect -11323 -333 -11245 -287
rect -11199 -333 -11121 -287
rect -11075 -333 -10997 -287
rect -10951 -333 -10873 -287
rect -10827 -333 -10749 -287
rect -10703 -333 -10625 -287
rect -10579 -333 -10501 -287
rect -10455 -333 -10377 -287
rect -10331 -333 -10253 -287
rect -10207 -333 -10129 -287
rect -10083 -333 -10005 -287
rect -9959 -333 -9881 -287
rect -9835 -333 -9757 -287
rect -9711 -333 -9633 -287
rect -9587 -333 -9509 -287
rect -9463 -333 -9385 -287
rect -9339 -333 -9261 -287
rect -9215 -333 -9137 -287
rect -9091 -333 -9013 -287
rect -8967 -333 -8889 -287
rect -8843 -333 -8765 -287
rect -8719 -333 -8641 -287
rect -8595 -333 -8517 -287
rect -8471 -333 -8393 -287
rect -8347 -333 -8269 -287
rect -8223 -333 -8145 -287
rect -8099 -333 -8021 -287
rect -7975 -333 -7897 -287
rect -7851 -333 -7773 -287
rect -7727 -333 -7649 -287
rect -7603 -333 -7525 -287
rect -7479 -333 -7401 -287
rect -7355 -333 -7277 -287
rect -7231 -333 -7153 -287
rect -7107 -333 -7029 -287
rect -6983 -333 -6905 -287
rect -6859 -333 -6781 -287
rect -6735 -333 -6657 -287
rect -6611 -333 -6533 -287
rect -6487 -333 -6409 -287
rect -6363 -333 -6285 -287
rect -6239 -333 -6161 -287
rect -6115 -333 -6037 -287
rect -5991 -333 -5913 -287
rect -5867 -333 -5789 -287
rect -5743 -333 -5665 -287
rect -5619 -333 -5541 -287
rect -5495 -333 -5417 -287
rect -5371 -333 -5293 -287
rect -5247 -333 -5169 -287
rect -5123 -333 -5045 -287
rect -4999 -333 -4921 -287
rect -4875 -333 -4797 -287
rect -4751 -333 -4673 -287
rect -4627 -333 -4549 -287
rect -4503 -333 -4425 -287
rect -4379 -333 -4301 -287
rect -4255 -333 -4177 -287
rect -4131 -333 -4053 -287
rect -4007 -333 -3929 -287
rect -3883 -333 -3805 -287
rect -3759 -333 -3681 -287
rect -3635 -333 -3557 -287
rect -3511 -333 -3433 -287
rect -3387 -333 -3309 -287
rect -3263 -333 -3185 -287
rect -3139 -333 -3061 -287
rect -3015 -333 -2937 -287
rect -2891 -333 -2813 -287
rect -2767 -333 -2689 -287
rect -2643 -333 -2565 -287
rect -2519 -333 -2441 -287
rect -2395 -333 -2317 -287
rect -2271 -333 -2193 -287
rect -2147 -333 -2069 -287
rect -2023 -333 -1945 -287
rect -1899 -333 -1821 -287
rect -1775 -333 -1697 -287
rect -1651 -333 -1573 -287
rect -1527 -333 -1449 -287
rect -1403 -333 -1325 -287
rect -1279 -333 -1201 -287
rect -1155 -333 -1077 -287
rect -1031 -333 -953 -287
rect -907 -333 -829 -287
rect -783 -333 -705 -287
rect -659 -333 -581 -287
rect -535 -333 -457 -287
rect -411 -333 -333 -287
rect -287 -333 -209 -287
rect -163 -333 -85 -287
rect -39 -333 39 -287
rect 85 -333 163 -287
rect 209 -333 287 -287
rect 333 -333 411 -287
rect 457 -333 535 -287
rect 581 -333 659 -287
rect 705 -333 783 -287
rect 829 -333 907 -287
rect 953 -333 1031 -287
rect 1077 -333 1155 -287
rect 1201 -333 1279 -287
rect 1325 -333 1403 -287
rect 1449 -333 1527 -287
rect 1573 -333 1651 -287
rect 1697 -333 1775 -287
rect 1821 -333 1899 -287
rect 1945 -333 2023 -287
rect 2069 -333 2147 -287
rect 2193 -333 2271 -287
rect 2317 -333 2395 -287
rect 2441 -333 2519 -287
rect 2565 -333 2643 -287
rect 2689 -333 2767 -287
rect 2813 -333 2891 -287
rect 2937 -333 3015 -287
rect 3061 -333 3139 -287
rect 3185 -333 3263 -287
rect 3309 -333 3387 -287
rect 3433 -333 3511 -287
rect 3557 -333 3635 -287
rect 3681 -333 3759 -287
rect 3805 -333 3883 -287
rect 3929 -333 4007 -287
rect 4053 -333 4131 -287
rect 4177 -333 4255 -287
rect 4301 -333 4379 -287
rect 4425 -333 4503 -287
rect 4549 -333 4627 -287
rect 4673 -333 4751 -287
rect 4797 -333 4875 -287
rect 4921 -333 4999 -287
rect 5045 -333 5123 -287
rect 5169 -333 5247 -287
rect 5293 -333 5371 -287
rect 5417 -333 5495 -287
rect 5541 -333 5619 -287
rect 5665 -333 5743 -287
rect 5789 -333 5867 -287
rect 5913 -333 5991 -287
rect 6037 -333 6115 -287
rect 6161 -333 6239 -287
rect 6285 -333 6363 -287
rect 6409 -333 6487 -287
rect 6533 -333 6611 -287
rect 6657 -333 6735 -287
rect 6781 -333 6859 -287
rect 6905 -333 6983 -287
rect 7029 -333 7107 -287
rect 7153 -333 7231 -287
rect 7277 -333 7355 -287
rect 7401 -333 7479 -287
rect 7525 -333 7603 -287
rect 7649 -333 7727 -287
rect 7773 -333 7851 -287
rect 7897 -333 7975 -287
rect 8021 -333 8099 -287
rect 8145 -333 8223 -287
rect 8269 -333 8347 -287
rect 8393 -333 8471 -287
rect 8517 -333 8595 -287
rect 8641 -333 8719 -287
rect 8765 -333 8843 -287
rect 8889 -333 8967 -287
rect 9013 -333 9091 -287
rect 9137 -333 9215 -287
rect 9261 -333 9339 -287
rect 9385 -333 9463 -287
rect 9509 -333 9587 -287
rect 9633 -333 9711 -287
rect 9757 -333 9835 -287
rect 9881 -333 9959 -287
rect 10005 -333 10083 -287
rect 10129 -333 10207 -287
rect 10253 -333 10331 -287
rect 10377 -333 10455 -287
rect 10501 -333 10579 -287
rect 10625 -333 10703 -287
rect 10749 -333 10827 -287
rect 10873 -333 10951 -287
rect 10997 -333 11075 -287
rect 11121 -333 11199 -287
rect 11245 -333 11323 -287
rect 11369 -333 11447 -287
rect 11493 -333 11571 -287
rect 11617 -333 11695 -287
rect 11741 -333 11819 -287
rect 11865 -333 11943 -287
rect 11989 -333 12067 -287
rect 12113 -333 12191 -287
rect 12237 -333 12315 -287
rect 12361 -333 12439 -287
rect 12485 -333 12563 -287
rect 12609 -333 12687 -287
rect 12733 -333 12811 -287
rect 12857 -333 12935 -287
rect 12981 -333 13059 -287
rect 13105 -333 13183 -287
rect 13229 -333 13307 -287
rect 13353 -333 13431 -287
rect 13477 -333 13555 -287
rect 13601 -333 13679 -287
rect 13725 -333 13803 -287
rect 13849 -333 13927 -287
rect 13973 -333 14051 -287
rect 14097 -333 14175 -287
rect 14221 -333 14299 -287
rect 14345 -333 14423 -287
rect 14469 -333 14547 -287
rect 14593 -333 14671 -287
rect 14717 -333 14795 -287
rect 14841 -333 14919 -287
rect 14965 -333 15043 -287
rect 15089 -333 15167 -287
rect 15213 -333 15291 -287
rect 15337 -333 15415 -287
rect 15461 -333 15539 -287
rect 15585 -333 15663 -287
rect 15709 -333 15787 -287
rect 15833 -333 15911 -287
rect 15957 -333 16035 -287
rect 16081 -333 16159 -287
rect 16205 -333 16283 -287
rect 16329 -333 16407 -287
rect 16453 -333 16531 -287
rect 16577 -333 16655 -287
rect 16701 -333 16779 -287
rect 16825 -333 16903 -287
rect 16949 -333 17027 -287
rect 17073 -333 17151 -287
rect 17197 -333 17275 -287
rect 17321 -333 17343 -287
rect -17343 -411 17343 -333
rect -17343 -457 -17321 -411
rect -17275 -457 -17197 -411
rect -17151 -457 -17073 -411
rect -17027 -457 -16949 -411
rect -16903 -457 -16825 -411
rect -16779 -457 -16701 -411
rect -16655 -457 -16577 -411
rect -16531 -457 -16453 -411
rect -16407 -457 -16329 -411
rect -16283 -457 -16205 -411
rect -16159 -457 -16081 -411
rect -16035 -457 -15957 -411
rect -15911 -457 -15833 -411
rect -15787 -457 -15709 -411
rect -15663 -457 -15585 -411
rect -15539 -457 -15461 -411
rect -15415 -457 -15337 -411
rect -15291 -457 -15213 -411
rect -15167 -457 -15089 -411
rect -15043 -457 -14965 -411
rect -14919 -457 -14841 -411
rect -14795 -457 -14717 -411
rect -14671 -457 -14593 -411
rect -14547 -457 -14469 -411
rect -14423 -457 -14345 -411
rect -14299 -457 -14221 -411
rect -14175 -457 -14097 -411
rect -14051 -457 -13973 -411
rect -13927 -457 -13849 -411
rect -13803 -457 -13725 -411
rect -13679 -457 -13601 -411
rect -13555 -457 -13477 -411
rect -13431 -457 -13353 -411
rect -13307 -457 -13229 -411
rect -13183 -457 -13105 -411
rect -13059 -457 -12981 -411
rect -12935 -457 -12857 -411
rect -12811 -457 -12733 -411
rect -12687 -457 -12609 -411
rect -12563 -457 -12485 -411
rect -12439 -457 -12361 -411
rect -12315 -457 -12237 -411
rect -12191 -457 -12113 -411
rect -12067 -457 -11989 -411
rect -11943 -457 -11865 -411
rect -11819 -457 -11741 -411
rect -11695 -457 -11617 -411
rect -11571 -457 -11493 -411
rect -11447 -457 -11369 -411
rect -11323 -457 -11245 -411
rect -11199 -457 -11121 -411
rect -11075 -457 -10997 -411
rect -10951 -457 -10873 -411
rect -10827 -457 -10749 -411
rect -10703 -457 -10625 -411
rect -10579 -457 -10501 -411
rect -10455 -457 -10377 -411
rect -10331 -457 -10253 -411
rect -10207 -457 -10129 -411
rect -10083 -457 -10005 -411
rect -9959 -457 -9881 -411
rect -9835 -457 -9757 -411
rect -9711 -457 -9633 -411
rect -9587 -457 -9509 -411
rect -9463 -457 -9385 -411
rect -9339 -457 -9261 -411
rect -9215 -457 -9137 -411
rect -9091 -457 -9013 -411
rect -8967 -457 -8889 -411
rect -8843 -457 -8765 -411
rect -8719 -457 -8641 -411
rect -8595 -457 -8517 -411
rect -8471 -457 -8393 -411
rect -8347 -457 -8269 -411
rect -8223 -457 -8145 -411
rect -8099 -457 -8021 -411
rect -7975 -457 -7897 -411
rect -7851 -457 -7773 -411
rect -7727 -457 -7649 -411
rect -7603 -457 -7525 -411
rect -7479 -457 -7401 -411
rect -7355 -457 -7277 -411
rect -7231 -457 -7153 -411
rect -7107 -457 -7029 -411
rect -6983 -457 -6905 -411
rect -6859 -457 -6781 -411
rect -6735 -457 -6657 -411
rect -6611 -457 -6533 -411
rect -6487 -457 -6409 -411
rect -6363 -457 -6285 -411
rect -6239 -457 -6161 -411
rect -6115 -457 -6037 -411
rect -5991 -457 -5913 -411
rect -5867 -457 -5789 -411
rect -5743 -457 -5665 -411
rect -5619 -457 -5541 -411
rect -5495 -457 -5417 -411
rect -5371 -457 -5293 -411
rect -5247 -457 -5169 -411
rect -5123 -457 -5045 -411
rect -4999 -457 -4921 -411
rect -4875 -457 -4797 -411
rect -4751 -457 -4673 -411
rect -4627 -457 -4549 -411
rect -4503 -457 -4425 -411
rect -4379 -457 -4301 -411
rect -4255 -457 -4177 -411
rect -4131 -457 -4053 -411
rect -4007 -457 -3929 -411
rect -3883 -457 -3805 -411
rect -3759 -457 -3681 -411
rect -3635 -457 -3557 -411
rect -3511 -457 -3433 -411
rect -3387 -457 -3309 -411
rect -3263 -457 -3185 -411
rect -3139 -457 -3061 -411
rect -3015 -457 -2937 -411
rect -2891 -457 -2813 -411
rect -2767 -457 -2689 -411
rect -2643 -457 -2565 -411
rect -2519 -457 -2441 -411
rect -2395 -457 -2317 -411
rect -2271 -457 -2193 -411
rect -2147 -457 -2069 -411
rect -2023 -457 -1945 -411
rect -1899 -457 -1821 -411
rect -1775 -457 -1697 -411
rect -1651 -457 -1573 -411
rect -1527 -457 -1449 -411
rect -1403 -457 -1325 -411
rect -1279 -457 -1201 -411
rect -1155 -457 -1077 -411
rect -1031 -457 -953 -411
rect -907 -457 -829 -411
rect -783 -457 -705 -411
rect -659 -457 -581 -411
rect -535 -457 -457 -411
rect -411 -457 -333 -411
rect -287 -457 -209 -411
rect -163 -457 -85 -411
rect -39 -457 39 -411
rect 85 -457 163 -411
rect 209 -457 287 -411
rect 333 -457 411 -411
rect 457 -457 535 -411
rect 581 -457 659 -411
rect 705 -457 783 -411
rect 829 -457 907 -411
rect 953 -457 1031 -411
rect 1077 -457 1155 -411
rect 1201 -457 1279 -411
rect 1325 -457 1403 -411
rect 1449 -457 1527 -411
rect 1573 -457 1651 -411
rect 1697 -457 1775 -411
rect 1821 -457 1899 -411
rect 1945 -457 2023 -411
rect 2069 -457 2147 -411
rect 2193 -457 2271 -411
rect 2317 -457 2395 -411
rect 2441 -457 2519 -411
rect 2565 -457 2643 -411
rect 2689 -457 2767 -411
rect 2813 -457 2891 -411
rect 2937 -457 3015 -411
rect 3061 -457 3139 -411
rect 3185 -457 3263 -411
rect 3309 -457 3387 -411
rect 3433 -457 3511 -411
rect 3557 -457 3635 -411
rect 3681 -457 3759 -411
rect 3805 -457 3883 -411
rect 3929 -457 4007 -411
rect 4053 -457 4131 -411
rect 4177 -457 4255 -411
rect 4301 -457 4379 -411
rect 4425 -457 4503 -411
rect 4549 -457 4627 -411
rect 4673 -457 4751 -411
rect 4797 -457 4875 -411
rect 4921 -457 4999 -411
rect 5045 -457 5123 -411
rect 5169 -457 5247 -411
rect 5293 -457 5371 -411
rect 5417 -457 5495 -411
rect 5541 -457 5619 -411
rect 5665 -457 5743 -411
rect 5789 -457 5867 -411
rect 5913 -457 5991 -411
rect 6037 -457 6115 -411
rect 6161 -457 6239 -411
rect 6285 -457 6363 -411
rect 6409 -457 6487 -411
rect 6533 -457 6611 -411
rect 6657 -457 6735 -411
rect 6781 -457 6859 -411
rect 6905 -457 6983 -411
rect 7029 -457 7107 -411
rect 7153 -457 7231 -411
rect 7277 -457 7355 -411
rect 7401 -457 7479 -411
rect 7525 -457 7603 -411
rect 7649 -457 7727 -411
rect 7773 -457 7851 -411
rect 7897 -457 7975 -411
rect 8021 -457 8099 -411
rect 8145 -457 8223 -411
rect 8269 -457 8347 -411
rect 8393 -457 8471 -411
rect 8517 -457 8595 -411
rect 8641 -457 8719 -411
rect 8765 -457 8843 -411
rect 8889 -457 8967 -411
rect 9013 -457 9091 -411
rect 9137 -457 9215 -411
rect 9261 -457 9339 -411
rect 9385 -457 9463 -411
rect 9509 -457 9587 -411
rect 9633 -457 9711 -411
rect 9757 -457 9835 -411
rect 9881 -457 9959 -411
rect 10005 -457 10083 -411
rect 10129 -457 10207 -411
rect 10253 -457 10331 -411
rect 10377 -457 10455 -411
rect 10501 -457 10579 -411
rect 10625 -457 10703 -411
rect 10749 -457 10827 -411
rect 10873 -457 10951 -411
rect 10997 -457 11075 -411
rect 11121 -457 11199 -411
rect 11245 -457 11323 -411
rect 11369 -457 11447 -411
rect 11493 -457 11571 -411
rect 11617 -457 11695 -411
rect 11741 -457 11819 -411
rect 11865 -457 11943 -411
rect 11989 -457 12067 -411
rect 12113 -457 12191 -411
rect 12237 -457 12315 -411
rect 12361 -457 12439 -411
rect 12485 -457 12563 -411
rect 12609 -457 12687 -411
rect 12733 -457 12811 -411
rect 12857 -457 12935 -411
rect 12981 -457 13059 -411
rect 13105 -457 13183 -411
rect 13229 -457 13307 -411
rect 13353 -457 13431 -411
rect 13477 -457 13555 -411
rect 13601 -457 13679 -411
rect 13725 -457 13803 -411
rect 13849 -457 13927 -411
rect 13973 -457 14051 -411
rect 14097 -457 14175 -411
rect 14221 -457 14299 -411
rect 14345 -457 14423 -411
rect 14469 -457 14547 -411
rect 14593 -457 14671 -411
rect 14717 -457 14795 -411
rect 14841 -457 14919 -411
rect 14965 -457 15043 -411
rect 15089 -457 15167 -411
rect 15213 -457 15291 -411
rect 15337 -457 15415 -411
rect 15461 -457 15539 -411
rect 15585 -457 15663 -411
rect 15709 -457 15787 -411
rect 15833 -457 15911 -411
rect 15957 -457 16035 -411
rect 16081 -457 16159 -411
rect 16205 -457 16283 -411
rect 16329 -457 16407 -411
rect 16453 -457 16531 -411
rect 16577 -457 16655 -411
rect 16701 -457 16779 -411
rect 16825 -457 16903 -411
rect 16949 -457 17027 -411
rect 17073 -457 17151 -411
rect 17197 -457 17275 -411
rect 17321 -457 17343 -411
rect -17343 -535 17343 -457
rect -17343 -581 -17321 -535
rect -17275 -581 -17197 -535
rect -17151 -581 -17073 -535
rect -17027 -581 -16949 -535
rect -16903 -581 -16825 -535
rect -16779 -581 -16701 -535
rect -16655 -581 -16577 -535
rect -16531 -581 -16453 -535
rect -16407 -581 -16329 -535
rect -16283 -581 -16205 -535
rect -16159 -581 -16081 -535
rect -16035 -581 -15957 -535
rect -15911 -581 -15833 -535
rect -15787 -581 -15709 -535
rect -15663 -581 -15585 -535
rect -15539 -581 -15461 -535
rect -15415 -581 -15337 -535
rect -15291 -581 -15213 -535
rect -15167 -581 -15089 -535
rect -15043 -581 -14965 -535
rect -14919 -581 -14841 -535
rect -14795 -581 -14717 -535
rect -14671 -581 -14593 -535
rect -14547 -581 -14469 -535
rect -14423 -581 -14345 -535
rect -14299 -581 -14221 -535
rect -14175 -581 -14097 -535
rect -14051 -581 -13973 -535
rect -13927 -581 -13849 -535
rect -13803 -581 -13725 -535
rect -13679 -581 -13601 -535
rect -13555 -581 -13477 -535
rect -13431 -581 -13353 -535
rect -13307 -581 -13229 -535
rect -13183 -581 -13105 -535
rect -13059 -581 -12981 -535
rect -12935 -581 -12857 -535
rect -12811 -581 -12733 -535
rect -12687 -581 -12609 -535
rect -12563 -581 -12485 -535
rect -12439 -581 -12361 -535
rect -12315 -581 -12237 -535
rect -12191 -581 -12113 -535
rect -12067 -581 -11989 -535
rect -11943 -581 -11865 -535
rect -11819 -581 -11741 -535
rect -11695 -581 -11617 -535
rect -11571 -581 -11493 -535
rect -11447 -581 -11369 -535
rect -11323 -581 -11245 -535
rect -11199 -581 -11121 -535
rect -11075 -581 -10997 -535
rect -10951 -581 -10873 -535
rect -10827 -581 -10749 -535
rect -10703 -581 -10625 -535
rect -10579 -581 -10501 -535
rect -10455 -581 -10377 -535
rect -10331 -581 -10253 -535
rect -10207 -581 -10129 -535
rect -10083 -581 -10005 -535
rect -9959 -581 -9881 -535
rect -9835 -581 -9757 -535
rect -9711 -581 -9633 -535
rect -9587 -581 -9509 -535
rect -9463 -581 -9385 -535
rect -9339 -581 -9261 -535
rect -9215 -581 -9137 -535
rect -9091 -581 -9013 -535
rect -8967 -581 -8889 -535
rect -8843 -581 -8765 -535
rect -8719 -581 -8641 -535
rect -8595 -581 -8517 -535
rect -8471 -581 -8393 -535
rect -8347 -581 -8269 -535
rect -8223 -581 -8145 -535
rect -8099 -581 -8021 -535
rect -7975 -581 -7897 -535
rect -7851 -581 -7773 -535
rect -7727 -581 -7649 -535
rect -7603 -581 -7525 -535
rect -7479 -581 -7401 -535
rect -7355 -581 -7277 -535
rect -7231 -581 -7153 -535
rect -7107 -581 -7029 -535
rect -6983 -581 -6905 -535
rect -6859 -581 -6781 -535
rect -6735 -581 -6657 -535
rect -6611 -581 -6533 -535
rect -6487 -581 -6409 -535
rect -6363 -581 -6285 -535
rect -6239 -581 -6161 -535
rect -6115 -581 -6037 -535
rect -5991 -581 -5913 -535
rect -5867 -581 -5789 -535
rect -5743 -581 -5665 -535
rect -5619 -581 -5541 -535
rect -5495 -581 -5417 -535
rect -5371 -581 -5293 -535
rect -5247 -581 -5169 -535
rect -5123 -581 -5045 -535
rect -4999 -581 -4921 -535
rect -4875 -581 -4797 -535
rect -4751 -581 -4673 -535
rect -4627 -581 -4549 -535
rect -4503 -581 -4425 -535
rect -4379 -581 -4301 -535
rect -4255 -581 -4177 -535
rect -4131 -581 -4053 -535
rect -4007 -581 -3929 -535
rect -3883 -581 -3805 -535
rect -3759 -581 -3681 -535
rect -3635 -581 -3557 -535
rect -3511 -581 -3433 -535
rect -3387 -581 -3309 -535
rect -3263 -581 -3185 -535
rect -3139 -581 -3061 -535
rect -3015 -581 -2937 -535
rect -2891 -581 -2813 -535
rect -2767 -581 -2689 -535
rect -2643 -581 -2565 -535
rect -2519 -581 -2441 -535
rect -2395 -581 -2317 -535
rect -2271 -581 -2193 -535
rect -2147 -581 -2069 -535
rect -2023 -581 -1945 -535
rect -1899 -581 -1821 -535
rect -1775 -581 -1697 -535
rect -1651 -581 -1573 -535
rect -1527 -581 -1449 -535
rect -1403 -581 -1325 -535
rect -1279 -581 -1201 -535
rect -1155 -581 -1077 -535
rect -1031 -581 -953 -535
rect -907 -581 -829 -535
rect -783 -581 -705 -535
rect -659 -581 -581 -535
rect -535 -581 -457 -535
rect -411 -581 -333 -535
rect -287 -581 -209 -535
rect -163 -581 -85 -535
rect -39 -581 39 -535
rect 85 -581 163 -535
rect 209 -581 287 -535
rect 333 -581 411 -535
rect 457 -581 535 -535
rect 581 -581 659 -535
rect 705 -581 783 -535
rect 829 -581 907 -535
rect 953 -581 1031 -535
rect 1077 -581 1155 -535
rect 1201 -581 1279 -535
rect 1325 -581 1403 -535
rect 1449 -581 1527 -535
rect 1573 -581 1651 -535
rect 1697 -581 1775 -535
rect 1821 -581 1899 -535
rect 1945 -581 2023 -535
rect 2069 -581 2147 -535
rect 2193 -581 2271 -535
rect 2317 -581 2395 -535
rect 2441 -581 2519 -535
rect 2565 -581 2643 -535
rect 2689 -581 2767 -535
rect 2813 -581 2891 -535
rect 2937 -581 3015 -535
rect 3061 -581 3139 -535
rect 3185 -581 3263 -535
rect 3309 -581 3387 -535
rect 3433 -581 3511 -535
rect 3557 -581 3635 -535
rect 3681 -581 3759 -535
rect 3805 -581 3883 -535
rect 3929 -581 4007 -535
rect 4053 -581 4131 -535
rect 4177 -581 4255 -535
rect 4301 -581 4379 -535
rect 4425 -581 4503 -535
rect 4549 -581 4627 -535
rect 4673 -581 4751 -535
rect 4797 -581 4875 -535
rect 4921 -581 4999 -535
rect 5045 -581 5123 -535
rect 5169 -581 5247 -535
rect 5293 -581 5371 -535
rect 5417 -581 5495 -535
rect 5541 -581 5619 -535
rect 5665 -581 5743 -535
rect 5789 -581 5867 -535
rect 5913 -581 5991 -535
rect 6037 -581 6115 -535
rect 6161 -581 6239 -535
rect 6285 -581 6363 -535
rect 6409 -581 6487 -535
rect 6533 -581 6611 -535
rect 6657 -581 6735 -535
rect 6781 -581 6859 -535
rect 6905 -581 6983 -535
rect 7029 -581 7107 -535
rect 7153 -581 7231 -535
rect 7277 -581 7355 -535
rect 7401 -581 7479 -535
rect 7525 -581 7603 -535
rect 7649 -581 7727 -535
rect 7773 -581 7851 -535
rect 7897 -581 7975 -535
rect 8021 -581 8099 -535
rect 8145 -581 8223 -535
rect 8269 -581 8347 -535
rect 8393 -581 8471 -535
rect 8517 -581 8595 -535
rect 8641 -581 8719 -535
rect 8765 -581 8843 -535
rect 8889 -581 8967 -535
rect 9013 -581 9091 -535
rect 9137 -581 9215 -535
rect 9261 -581 9339 -535
rect 9385 -581 9463 -535
rect 9509 -581 9587 -535
rect 9633 -581 9711 -535
rect 9757 -581 9835 -535
rect 9881 -581 9959 -535
rect 10005 -581 10083 -535
rect 10129 -581 10207 -535
rect 10253 -581 10331 -535
rect 10377 -581 10455 -535
rect 10501 -581 10579 -535
rect 10625 -581 10703 -535
rect 10749 -581 10827 -535
rect 10873 -581 10951 -535
rect 10997 -581 11075 -535
rect 11121 -581 11199 -535
rect 11245 -581 11323 -535
rect 11369 -581 11447 -535
rect 11493 -581 11571 -535
rect 11617 -581 11695 -535
rect 11741 -581 11819 -535
rect 11865 -581 11943 -535
rect 11989 -581 12067 -535
rect 12113 -581 12191 -535
rect 12237 -581 12315 -535
rect 12361 -581 12439 -535
rect 12485 -581 12563 -535
rect 12609 -581 12687 -535
rect 12733 -581 12811 -535
rect 12857 -581 12935 -535
rect 12981 -581 13059 -535
rect 13105 -581 13183 -535
rect 13229 -581 13307 -535
rect 13353 -581 13431 -535
rect 13477 -581 13555 -535
rect 13601 -581 13679 -535
rect 13725 -581 13803 -535
rect 13849 -581 13927 -535
rect 13973 -581 14051 -535
rect 14097 -581 14175 -535
rect 14221 -581 14299 -535
rect 14345 -581 14423 -535
rect 14469 -581 14547 -535
rect 14593 -581 14671 -535
rect 14717 -581 14795 -535
rect 14841 -581 14919 -535
rect 14965 -581 15043 -535
rect 15089 -581 15167 -535
rect 15213 -581 15291 -535
rect 15337 -581 15415 -535
rect 15461 -581 15539 -535
rect 15585 -581 15663 -535
rect 15709 -581 15787 -535
rect 15833 -581 15911 -535
rect 15957 -581 16035 -535
rect 16081 -581 16159 -535
rect 16205 -581 16283 -535
rect 16329 -581 16407 -535
rect 16453 -581 16531 -535
rect 16577 -581 16655 -535
rect 16701 -581 16779 -535
rect 16825 -581 16903 -535
rect 16949 -581 17027 -535
rect 17073 -581 17151 -535
rect 17197 -581 17275 -535
rect 17321 -581 17343 -535
rect -17343 -659 17343 -581
rect -17343 -705 -17321 -659
rect -17275 -705 -17197 -659
rect -17151 -705 -17073 -659
rect -17027 -705 -16949 -659
rect -16903 -705 -16825 -659
rect -16779 -705 -16701 -659
rect -16655 -705 -16577 -659
rect -16531 -705 -16453 -659
rect -16407 -705 -16329 -659
rect -16283 -705 -16205 -659
rect -16159 -705 -16081 -659
rect -16035 -705 -15957 -659
rect -15911 -705 -15833 -659
rect -15787 -705 -15709 -659
rect -15663 -705 -15585 -659
rect -15539 -705 -15461 -659
rect -15415 -705 -15337 -659
rect -15291 -705 -15213 -659
rect -15167 -705 -15089 -659
rect -15043 -705 -14965 -659
rect -14919 -705 -14841 -659
rect -14795 -705 -14717 -659
rect -14671 -705 -14593 -659
rect -14547 -705 -14469 -659
rect -14423 -705 -14345 -659
rect -14299 -705 -14221 -659
rect -14175 -705 -14097 -659
rect -14051 -705 -13973 -659
rect -13927 -705 -13849 -659
rect -13803 -705 -13725 -659
rect -13679 -705 -13601 -659
rect -13555 -705 -13477 -659
rect -13431 -705 -13353 -659
rect -13307 -705 -13229 -659
rect -13183 -705 -13105 -659
rect -13059 -705 -12981 -659
rect -12935 -705 -12857 -659
rect -12811 -705 -12733 -659
rect -12687 -705 -12609 -659
rect -12563 -705 -12485 -659
rect -12439 -705 -12361 -659
rect -12315 -705 -12237 -659
rect -12191 -705 -12113 -659
rect -12067 -705 -11989 -659
rect -11943 -705 -11865 -659
rect -11819 -705 -11741 -659
rect -11695 -705 -11617 -659
rect -11571 -705 -11493 -659
rect -11447 -705 -11369 -659
rect -11323 -705 -11245 -659
rect -11199 -705 -11121 -659
rect -11075 -705 -10997 -659
rect -10951 -705 -10873 -659
rect -10827 -705 -10749 -659
rect -10703 -705 -10625 -659
rect -10579 -705 -10501 -659
rect -10455 -705 -10377 -659
rect -10331 -705 -10253 -659
rect -10207 -705 -10129 -659
rect -10083 -705 -10005 -659
rect -9959 -705 -9881 -659
rect -9835 -705 -9757 -659
rect -9711 -705 -9633 -659
rect -9587 -705 -9509 -659
rect -9463 -705 -9385 -659
rect -9339 -705 -9261 -659
rect -9215 -705 -9137 -659
rect -9091 -705 -9013 -659
rect -8967 -705 -8889 -659
rect -8843 -705 -8765 -659
rect -8719 -705 -8641 -659
rect -8595 -705 -8517 -659
rect -8471 -705 -8393 -659
rect -8347 -705 -8269 -659
rect -8223 -705 -8145 -659
rect -8099 -705 -8021 -659
rect -7975 -705 -7897 -659
rect -7851 -705 -7773 -659
rect -7727 -705 -7649 -659
rect -7603 -705 -7525 -659
rect -7479 -705 -7401 -659
rect -7355 -705 -7277 -659
rect -7231 -705 -7153 -659
rect -7107 -705 -7029 -659
rect -6983 -705 -6905 -659
rect -6859 -705 -6781 -659
rect -6735 -705 -6657 -659
rect -6611 -705 -6533 -659
rect -6487 -705 -6409 -659
rect -6363 -705 -6285 -659
rect -6239 -705 -6161 -659
rect -6115 -705 -6037 -659
rect -5991 -705 -5913 -659
rect -5867 -705 -5789 -659
rect -5743 -705 -5665 -659
rect -5619 -705 -5541 -659
rect -5495 -705 -5417 -659
rect -5371 -705 -5293 -659
rect -5247 -705 -5169 -659
rect -5123 -705 -5045 -659
rect -4999 -705 -4921 -659
rect -4875 -705 -4797 -659
rect -4751 -705 -4673 -659
rect -4627 -705 -4549 -659
rect -4503 -705 -4425 -659
rect -4379 -705 -4301 -659
rect -4255 -705 -4177 -659
rect -4131 -705 -4053 -659
rect -4007 -705 -3929 -659
rect -3883 -705 -3805 -659
rect -3759 -705 -3681 -659
rect -3635 -705 -3557 -659
rect -3511 -705 -3433 -659
rect -3387 -705 -3309 -659
rect -3263 -705 -3185 -659
rect -3139 -705 -3061 -659
rect -3015 -705 -2937 -659
rect -2891 -705 -2813 -659
rect -2767 -705 -2689 -659
rect -2643 -705 -2565 -659
rect -2519 -705 -2441 -659
rect -2395 -705 -2317 -659
rect -2271 -705 -2193 -659
rect -2147 -705 -2069 -659
rect -2023 -705 -1945 -659
rect -1899 -705 -1821 -659
rect -1775 -705 -1697 -659
rect -1651 -705 -1573 -659
rect -1527 -705 -1449 -659
rect -1403 -705 -1325 -659
rect -1279 -705 -1201 -659
rect -1155 -705 -1077 -659
rect -1031 -705 -953 -659
rect -907 -705 -829 -659
rect -783 -705 -705 -659
rect -659 -705 -581 -659
rect -535 -705 -457 -659
rect -411 -705 -333 -659
rect -287 -705 -209 -659
rect -163 -705 -85 -659
rect -39 -705 39 -659
rect 85 -705 163 -659
rect 209 -705 287 -659
rect 333 -705 411 -659
rect 457 -705 535 -659
rect 581 -705 659 -659
rect 705 -705 783 -659
rect 829 -705 907 -659
rect 953 -705 1031 -659
rect 1077 -705 1155 -659
rect 1201 -705 1279 -659
rect 1325 -705 1403 -659
rect 1449 -705 1527 -659
rect 1573 -705 1651 -659
rect 1697 -705 1775 -659
rect 1821 -705 1899 -659
rect 1945 -705 2023 -659
rect 2069 -705 2147 -659
rect 2193 -705 2271 -659
rect 2317 -705 2395 -659
rect 2441 -705 2519 -659
rect 2565 -705 2643 -659
rect 2689 -705 2767 -659
rect 2813 -705 2891 -659
rect 2937 -705 3015 -659
rect 3061 -705 3139 -659
rect 3185 -705 3263 -659
rect 3309 -705 3387 -659
rect 3433 -705 3511 -659
rect 3557 -705 3635 -659
rect 3681 -705 3759 -659
rect 3805 -705 3883 -659
rect 3929 -705 4007 -659
rect 4053 -705 4131 -659
rect 4177 -705 4255 -659
rect 4301 -705 4379 -659
rect 4425 -705 4503 -659
rect 4549 -705 4627 -659
rect 4673 -705 4751 -659
rect 4797 -705 4875 -659
rect 4921 -705 4999 -659
rect 5045 -705 5123 -659
rect 5169 -705 5247 -659
rect 5293 -705 5371 -659
rect 5417 -705 5495 -659
rect 5541 -705 5619 -659
rect 5665 -705 5743 -659
rect 5789 -705 5867 -659
rect 5913 -705 5991 -659
rect 6037 -705 6115 -659
rect 6161 -705 6239 -659
rect 6285 -705 6363 -659
rect 6409 -705 6487 -659
rect 6533 -705 6611 -659
rect 6657 -705 6735 -659
rect 6781 -705 6859 -659
rect 6905 -705 6983 -659
rect 7029 -705 7107 -659
rect 7153 -705 7231 -659
rect 7277 -705 7355 -659
rect 7401 -705 7479 -659
rect 7525 -705 7603 -659
rect 7649 -705 7727 -659
rect 7773 -705 7851 -659
rect 7897 -705 7975 -659
rect 8021 -705 8099 -659
rect 8145 -705 8223 -659
rect 8269 -705 8347 -659
rect 8393 -705 8471 -659
rect 8517 -705 8595 -659
rect 8641 -705 8719 -659
rect 8765 -705 8843 -659
rect 8889 -705 8967 -659
rect 9013 -705 9091 -659
rect 9137 -705 9215 -659
rect 9261 -705 9339 -659
rect 9385 -705 9463 -659
rect 9509 -705 9587 -659
rect 9633 -705 9711 -659
rect 9757 -705 9835 -659
rect 9881 -705 9959 -659
rect 10005 -705 10083 -659
rect 10129 -705 10207 -659
rect 10253 -705 10331 -659
rect 10377 -705 10455 -659
rect 10501 -705 10579 -659
rect 10625 -705 10703 -659
rect 10749 -705 10827 -659
rect 10873 -705 10951 -659
rect 10997 -705 11075 -659
rect 11121 -705 11199 -659
rect 11245 -705 11323 -659
rect 11369 -705 11447 -659
rect 11493 -705 11571 -659
rect 11617 -705 11695 -659
rect 11741 -705 11819 -659
rect 11865 -705 11943 -659
rect 11989 -705 12067 -659
rect 12113 -705 12191 -659
rect 12237 -705 12315 -659
rect 12361 -705 12439 -659
rect 12485 -705 12563 -659
rect 12609 -705 12687 -659
rect 12733 -705 12811 -659
rect 12857 -705 12935 -659
rect 12981 -705 13059 -659
rect 13105 -705 13183 -659
rect 13229 -705 13307 -659
rect 13353 -705 13431 -659
rect 13477 -705 13555 -659
rect 13601 -705 13679 -659
rect 13725 -705 13803 -659
rect 13849 -705 13927 -659
rect 13973 -705 14051 -659
rect 14097 -705 14175 -659
rect 14221 -705 14299 -659
rect 14345 -705 14423 -659
rect 14469 -705 14547 -659
rect 14593 -705 14671 -659
rect 14717 -705 14795 -659
rect 14841 -705 14919 -659
rect 14965 -705 15043 -659
rect 15089 -705 15167 -659
rect 15213 -705 15291 -659
rect 15337 -705 15415 -659
rect 15461 -705 15539 -659
rect 15585 -705 15663 -659
rect 15709 -705 15787 -659
rect 15833 -705 15911 -659
rect 15957 -705 16035 -659
rect 16081 -705 16159 -659
rect 16205 -705 16283 -659
rect 16329 -705 16407 -659
rect 16453 -705 16531 -659
rect 16577 -705 16655 -659
rect 16701 -705 16779 -659
rect 16825 -705 16903 -659
rect 16949 -705 17027 -659
rect 17073 -705 17151 -659
rect 17197 -705 17275 -659
rect 17321 -705 17343 -659
rect -17343 -783 17343 -705
rect -17343 -829 -17321 -783
rect -17275 -829 -17197 -783
rect -17151 -829 -17073 -783
rect -17027 -829 -16949 -783
rect -16903 -829 -16825 -783
rect -16779 -829 -16701 -783
rect -16655 -829 -16577 -783
rect -16531 -829 -16453 -783
rect -16407 -829 -16329 -783
rect -16283 -829 -16205 -783
rect -16159 -829 -16081 -783
rect -16035 -829 -15957 -783
rect -15911 -829 -15833 -783
rect -15787 -829 -15709 -783
rect -15663 -829 -15585 -783
rect -15539 -829 -15461 -783
rect -15415 -829 -15337 -783
rect -15291 -829 -15213 -783
rect -15167 -829 -15089 -783
rect -15043 -829 -14965 -783
rect -14919 -829 -14841 -783
rect -14795 -829 -14717 -783
rect -14671 -829 -14593 -783
rect -14547 -829 -14469 -783
rect -14423 -829 -14345 -783
rect -14299 -829 -14221 -783
rect -14175 -829 -14097 -783
rect -14051 -829 -13973 -783
rect -13927 -829 -13849 -783
rect -13803 -829 -13725 -783
rect -13679 -829 -13601 -783
rect -13555 -829 -13477 -783
rect -13431 -829 -13353 -783
rect -13307 -829 -13229 -783
rect -13183 -829 -13105 -783
rect -13059 -829 -12981 -783
rect -12935 -829 -12857 -783
rect -12811 -829 -12733 -783
rect -12687 -829 -12609 -783
rect -12563 -829 -12485 -783
rect -12439 -829 -12361 -783
rect -12315 -829 -12237 -783
rect -12191 -829 -12113 -783
rect -12067 -829 -11989 -783
rect -11943 -829 -11865 -783
rect -11819 -829 -11741 -783
rect -11695 -829 -11617 -783
rect -11571 -829 -11493 -783
rect -11447 -829 -11369 -783
rect -11323 -829 -11245 -783
rect -11199 -829 -11121 -783
rect -11075 -829 -10997 -783
rect -10951 -829 -10873 -783
rect -10827 -829 -10749 -783
rect -10703 -829 -10625 -783
rect -10579 -829 -10501 -783
rect -10455 -829 -10377 -783
rect -10331 -829 -10253 -783
rect -10207 -829 -10129 -783
rect -10083 -829 -10005 -783
rect -9959 -829 -9881 -783
rect -9835 -829 -9757 -783
rect -9711 -829 -9633 -783
rect -9587 -829 -9509 -783
rect -9463 -829 -9385 -783
rect -9339 -829 -9261 -783
rect -9215 -829 -9137 -783
rect -9091 -829 -9013 -783
rect -8967 -829 -8889 -783
rect -8843 -829 -8765 -783
rect -8719 -829 -8641 -783
rect -8595 -829 -8517 -783
rect -8471 -829 -8393 -783
rect -8347 -829 -8269 -783
rect -8223 -829 -8145 -783
rect -8099 -829 -8021 -783
rect -7975 -829 -7897 -783
rect -7851 -829 -7773 -783
rect -7727 -829 -7649 -783
rect -7603 -829 -7525 -783
rect -7479 -829 -7401 -783
rect -7355 -829 -7277 -783
rect -7231 -829 -7153 -783
rect -7107 -829 -7029 -783
rect -6983 -829 -6905 -783
rect -6859 -829 -6781 -783
rect -6735 -829 -6657 -783
rect -6611 -829 -6533 -783
rect -6487 -829 -6409 -783
rect -6363 -829 -6285 -783
rect -6239 -829 -6161 -783
rect -6115 -829 -6037 -783
rect -5991 -829 -5913 -783
rect -5867 -829 -5789 -783
rect -5743 -829 -5665 -783
rect -5619 -829 -5541 -783
rect -5495 -829 -5417 -783
rect -5371 -829 -5293 -783
rect -5247 -829 -5169 -783
rect -5123 -829 -5045 -783
rect -4999 -829 -4921 -783
rect -4875 -829 -4797 -783
rect -4751 -829 -4673 -783
rect -4627 -829 -4549 -783
rect -4503 -829 -4425 -783
rect -4379 -829 -4301 -783
rect -4255 -829 -4177 -783
rect -4131 -829 -4053 -783
rect -4007 -829 -3929 -783
rect -3883 -829 -3805 -783
rect -3759 -829 -3681 -783
rect -3635 -829 -3557 -783
rect -3511 -829 -3433 -783
rect -3387 -829 -3309 -783
rect -3263 -829 -3185 -783
rect -3139 -829 -3061 -783
rect -3015 -829 -2937 -783
rect -2891 -829 -2813 -783
rect -2767 -829 -2689 -783
rect -2643 -829 -2565 -783
rect -2519 -829 -2441 -783
rect -2395 -829 -2317 -783
rect -2271 -829 -2193 -783
rect -2147 -829 -2069 -783
rect -2023 -829 -1945 -783
rect -1899 -829 -1821 -783
rect -1775 -829 -1697 -783
rect -1651 -829 -1573 -783
rect -1527 -829 -1449 -783
rect -1403 -829 -1325 -783
rect -1279 -829 -1201 -783
rect -1155 -829 -1077 -783
rect -1031 -829 -953 -783
rect -907 -829 -829 -783
rect -783 -829 -705 -783
rect -659 -829 -581 -783
rect -535 -829 -457 -783
rect -411 -829 -333 -783
rect -287 -829 -209 -783
rect -163 -829 -85 -783
rect -39 -829 39 -783
rect 85 -829 163 -783
rect 209 -829 287 -783
rect 333 -829 411 -783
rect 457 -829 535 -783
rect 581 -829 659 -783
rect 705 -829 783 -783
rect 829 -829 907 -783
rect 953 -829 1031 -783
rect 1077 -829 1155 -783
rect 1201 -829 1279 -783
rect 1325 -829 1403 -783
rect 1449 -829 1527 -783
rect 1573 -829 1651 -783
rect 1697 -829 1775 -783
rect 1821 -829 1899 -783
rect 1945 -829 2023 -783
rect 2069 -829 2147 -783
rect 2193 -829 2271 -783
rect 2317 -829 2395 -783
rect 2441 -829 2519 -783
rect 2565 -829 2643 -783
rect 2689 -829 2767 -783
rect 2813 -829 2891 -783
rect 2937 -829 3015 -783
rect 3061 -829 3139 -783
rect 3185 -829 3263 -783
rect 3309 -829 3387 -783
rect 3433 -829 3511 -783
rect 3557 -829 3635 -783
rect 3681 -829 3759 -783
rect 3805 -829 3883 -783
rect 3929 -829 4007 -783
rect 4053 -829 4131 -783
rect 4177 -829 4255 -783
rect 4301 -829 4379 -783
rect 4425 -829 4503 -783
rect 4549 -829 4627 -783
rect 4673 -829 4751 -783
rect 4797 -829 4875 -783
rect 4921 -829 4999 -783
rect 5045 -829 5123 -783
rect 5169 -829 5247 -783
rect 5293 -829 5371 -783
rect 5417 -829 5495 -783
rect 5541 -829 5619 -783
rect 5665 -829 5743 -783
rect 5789 -829 5867 -783
rect 5913 -829 5991 -783
rect 6037 -829 6115 -783
rect 6161 -829 6239 -783
rect 6285 -829 6363 -783
rect 6409 -829 6487 -783
rect 6533 -829 6611 -783
rect 6657 -829 6735 -783
rect 6781 -829 6859 -783
rect 6905 -829 6983 -783
rect 7029 -829 7107 -783
rect 7153 -829 7231 -783
rect 7277 -829 7355 -783
rect 7401 -829 7479 -783
rect 7525 -829 7603 -783
rect 7649 -829 7727 -783
rect 7773 -829 7851 -783
rect 7897 -829 7975 -783
rect 8021 -829 8099 -783
rect 8145 -829 8223 -783
rect 8269 -829 8347 -783
rect 8393 -829 8471 -783
rect 8517 -829 8595 -783
rect 8641 -829 8719 -783
rect 8765 -829 8843 -783
rect 8889 -829 8967 -783
rect 9013 -829 9091 -783
rect 9137 -829 9215 -783
rect 9261 -829 9339 -783
rect 9385 -829 9463 -783
rect 9509 -829 9587 -783
rect 9633 -829 9711 -783
rect 9757 -829 9835 -783
rect 9881 -829 9959 -783
rect 10005 -829 10083 -783
rect 10129 -829 10207 -783
rect 10253 -829 10331 -783
rect 10377 -829 10455 -783
rect 10501 -829 10579 -783
rect 10625 -829 10703 -783
rect 10749 -829 10827 -783
rect 10873 -829 10951 -783
rect 10997 -829 11075 -783
rect 11121 -829 11199 -783
rect 11245 -829 11323 -783
rect 11369 -829 11447 -783
rect 11493 -829 11571 -783
rect 11617 -829 11695 -783
rect 11741 -829 11819 -783
rect 11865 -829 11943 -783
rect 11989 -829 12067 -783
rect 12113 -829 12191 -783
rect 12237 -829 12315 -783
rect 12361 -829 12439 -783
rect 12485 -829 12563 -783
rect 12609 -829 12687 -783
rect 12733 -829 12811 -783
rect 12857 -829 12935 -783
rect 12981 -829 13059 -783
rect 13105 -829 13183 -783
rect 13229 -829 13307 -783
rect 13353 -829 13431 -783
rect 13477 -829 13555 -783
rect 13601 -829 13679 -783
rect 13725 -829 13803 -783
rect 13849 -829 13927 -783
rect 13973 -829 14051 -783
rect 14097 -829 14175 -783
rect 14221 -829 14299 -783
rect 14345 -829 14423 -783
rect 14469 -829 14547 -783
rect 14593 -829 14671 -783
rect 14717 -829 14795 -783
rect 14841 -829 14919 -783
rect 14965 -829 15043 -783
rect 15089 -829 15167 -783
rect 15213 -829 15291 -783
rect 15337 -829 15415 -783
rect 15461 -829 15539 -783
rect 15585 -829 15663 -783
rect 15709 -829 15787 -783
rect 15833 -829 15911 -783
rect 15957 -829 16035 -783
rect 16081 -829 16159 -783
rect 16205 -829 16283 -783
rect 16329 -829 16407 -783
rect 16453 -829 16531 -783
rect 16577 -829 16655 -783
rect 16701 -829 16779 -783
rect 16825 -829 16903 -783
rect 16949 -829 17027 -783
rect 17073 -829 17151 -783
rect 17197 -829 17275 -783
rect 17321 -829 17343 -783
rect -17343 -907 17343 -829
rect -17343 -953 -17321 -907
rect -17275 -953 -17197 -907
rect -17151 -953 -17073 -907
rect -17027 -953 -16949 -907
rect -16903 -953 -16825 -907
rect -16779 -953 -16701 -907
rect -16655 -953 -16577 -907
rect -16531 -953 -16453 -907
rect -16407 -953 -16329 -907
rect -16283 -953 -16205 -907
rect -16159 -953 -16081 -907
rect -16035 -953 -15957 -907
rect -15911 -953 -15833 -907
rect -15787 -953 -15709 -907
rect -15663 -953 -15585 -907
rect -15539 -953 -15461 -907
rect -15415 -953 -15337 -907
rect -15291 -953 -15213 -907
rect -15167 -953 -15089 -907
rect -15043 -953 -14965 -907
rect -14919 -953 -14841 -907
rect -14795 -953 -14717 -907
rect -14671 -953 -14593 -907
rect -14547 -953 -14469 -907
rect -14423 -953 -14345 -907
rect -14299 -953 -14221 -907
rect -14175 -953 -14097 -907
rect -14051 -953 -13973 -907
rect -13927 -953 -13849 -907
rect -13803 -953 -13725 -907
rect -13679 -953 -13601 -907
rect -13555 -953 -13477 -907
rect -13431 -953 -13353 -907
rect -13307 -953 -13229 -907
rect -13183 -953 -13105 -907
rect -13059 -953 -12981 -907
rect -12935 -953 -12857 -907
rect -12811 -953 -12733 -907
rect -12687 -953 -12609 -907
rect -12563 -953 -12485 -907
rect -12439 -953 -12361 -907
rect -12315 -953 -12237 -907
rect -12191 -953 -12113 -907
rect -12067 -953 -11989 -907
rect -11943 -953 -11865 -907
rect -11819 -953 -11741 -907
rect -11695 -953 -11617 -907
rect -11571 -953 -11493 -907
rect -11447 -953 -11369 -907
rect -11323 -953 -11245 -907
rect -11199 -953 -11121 -907
rect -11075 -953 -10997 -907
rect -10951 -953 -10873 -907
rect -10827 -953 -10749 -907
rect -10703 -953 -10625 -907
rect -10579 -953 -10501 -907
rect -10455 -953 -10377 -907
rect -10331 -953 -10253 -907
rect -10207 -953 -10129 -907
rect -10083 -953 -10005 -907
rect -9959 -953 -9881 -907
rect -9835 -953 -9757 -907
rect -9711 -953 -9633 -907
rect -9587 -953 -9509 -907
rect -9463 -953 -9385 -907
rect -9339 -953 -9261 -907
rect -9215 -953 -9137 -907
rect -9091 -953 -9013 -907
rect -8967 -953 -8889 -907
rect -8843 -953 -8765 -907
rect -8719 -953 -8641 -907
rect -8595 -953 -8517 -907
rect -8471 -953 -8393 -907
rect -8347 -953 -8269 -907
rect -8223 -953 -8145 -907
rect -8099 -953 -8021 -907
rect -7975 -953 -7897 -907
rect -7851 -953 -7773 -907
rect -7727 -953 -7649 -907
rect -7603 -953 -7525 -907
rect -7479 -953 -7401 -907
rect -7355 -953 -7277 -907
rect -7231 -953 -7153 -907
rect -7107 -953 -7029 -907
rect -6983 -953 -6905 -907
rect -6859 -953 -6781 -907
rect -6735 -953 -6657 -907
rect -6611 -953 -6533 -907
rect -6487 -953 -6409 -907
rect -6363 -953 -6285 -907
rect -6239 -953 -6161 -907
rect -6115 -953 -6037 -907
rect -5991 -953 -5913 -907
rect -5867 -953 -5789 -907
rect -5743 -953 -5665 -907
rect -5619 -953 -5541 -907
rect -5495 -953 -5417 -907
rect -5371 -953 -5293 -907
rect -5247 -953 -5169 -907
rect -5123 -953 -5045 -907
rect -4999 -953 -4921 -907
rect -4875 -953 -4797 -907
rect -4751 -953 -4673 -907
rect -4627 -953 -4549 -907
rect -4503 -953 -4425 -907
rect -4379 -953 -4301 -907
rect -4255 -953 -4177 -907
rect -4131 -953 -4053 -907
rect -4007 -953 -3929 -907
rect -3883 -953 -3805 -907
rect -3759 -953 -3681 -907
rect -3635 -953 -3557 -907
rect -3511 -953 -3433 -907
rect -3387 -953 -3309 -907
rect -3263 -953 -3185 -907
rect -3139 -953 -3061 -907
rect -3015 -953 -2937 -907
rect -2891 -953 -2813 -907
rect -2767 -953 -2689 -907
rect -2643 -953 -2565 -907
rect -2519 -953 -2441 -907
rect -2395 -953 -2317 -907
rect -2271 -953 -2193 -907
rect -2147 -953 -2069 -907
rect -2023 -953 -1945 -907
rect -1899 -953 -1821 -907
rect -1775 -953 -1697 -907
rect -1651 -953 -1573 -907
rect -1527 -953 -1449 -907
rect -1403 -953 -1325 -907
rect -1279 -953 -1201 -907
rect -1155 -953 -1077 -907
rect -1031 -953 -953 -907
rect -907 -953 -829 -907
rect -783 -953 -705 -907
rect -659 -953 -581 -907
rect -535 -953 -457 -907
rect -411 -953 -333 -907
rect -287 -953 -209 -907
rect -163 -953 -85 -907
rect -39 -953 39 -907
rect 85 -953 163 -907
rect 209 -953 287 -907
rect 333 -953 411 -907
rect 457 -953 535 -907
rect 581 -953 659 -907
rect 705 -953 783 -907
rect 829 -953 907 -907
rect 953 -953 1031 -907
rect 1077 -953 1155 -907
rect 1201 -953 1279 -907
rect 1325 -953 1403 -907
rect 1449 -953 1527 -907
rect 1573 -953 1651 -907
rect 1697 -953 1775 -907
rect 1821 -953 1899 -907
rect 1945 -953 2023 -907
rect 2069 -953 2147 -907
rect 2193 -953 2271 -907
rect 2317 -953 2395 -907
rect 2441 -953 2519 -907
rect 2565 -953 2643 -907
rect 2689 -953 2767 -907
rect 2813 -953 2891 -907
rect 2937 -953 3015 -907
rect 3061 -953 3139 -907
rect 3185 -953 3263 -907
rect 3309 -953 3387 -907
rect 3433 -953 3511 -907
rect 3557 -953 3635 -907
rect 3681 -953 3759 -907
rect 3805 -953 3883 -907
rect 3929 -953 4007 -907
rect 4053 -953 4131 -907
rect 4177 -953 4255 -907
rect 4301 -953 4379 -907
rect 4425 -953 4503 -907
rect 4549 -953 4627 -907
rect 4673 -953 4751 -907
rect 4797 -953 4875 -907
rect 4921 -953 4999 -907
rect 5045 -953 5123 -907
rect 5169 -953 5247 -907
rect 5293 -953 5371 -907
rect 5417 -953 5495 -907
rect 5541 -953 5619 -907
rect 5665 -953 5743 -907
rect 5789 -953 5867 -907
rect 5913 -953 5991 -907
rect 6037 -953 6115 -907
rect 6161 -953 6239 -907
rect 6285 -953 6363 -907
rect 6409 -953 6487 -907
rect 6533 -953 6611 -907
rect 6657 -953 6735 -907
rect 6781 -953 6859 -907
rect 6905 -953 6983 -907
rect 7029 -953 7107 -907
rect 7153 -953 7231 -907
rect 7277 -953 7355 -907
rect 7401 -953 7479 -907
rect 7525 -953 7603 -907
rect 7649 -953 7727 -907
rect 7773 -953 7851 -907
rect 7897 -953 7975 -907
rect 8021 -953 8099 -907
rect 8145 -953 8223 -907
rect 8269 -953 8347 -907
rect 8393 -953 8471 -907
rect 8517 -953 8595 -907
rect 8641 -953 8719 -907
rect 8765 -953 8843 -907
rect 8889 -953 8967 -907
rect 9013 -953 9091 -907
rect 9137 -953 9215 -907
rect 9261 -953 9339 -907
rect 9385 -953 9463 -907
rect 9509 -953 9587 -907
rect 9633 -953 9711 -907
rect 9757 -953 9835 -907
rect 9881 -953 9959 -907
rect 10005 -953 10083 -907
rect 10129 -953 10207 -907
rect 10253 -953 10331 -907
rect 10377 -953 10455 -907
rect 10501 -953 10579 -907
rect 10625 -953 10703 -907
rect 10749 -953 10827 -907
rect 10873 -953 10951 -907
rect 10997 -953 11075 -907
rect 11121 -953 11199 -907
rect 11245 -953 11323 -907
rect 11369 -953 11447 -907
rect 11493 -953 11571 -907
rect 11617 -953 11695 -907
rect 11741 -953 11819 -907
rect 11865 -953 11943 -907
rect 11989 -953 12067 -907
rect 12113 -953 12191 -907
rect 12237 -953 12315 -907
rect 12361 -953 12439 -907
rect 12485 -953 12563 -907
rect 12609 -953 12687 -907
rect 12733 -953 12811 -907
rect 12857 -953 12935 -907
rect 12981 -953 13059 -907
rect 13105 -953 13183 -907
rect 13229 -953 13307 -907
rect 13353 -953 13431 -907
rect 13477 -953 13555 -907
rect 13601 -953 13679 -907
rect 13725 -953 13803 -907
rect 13849 -953 13927 -907
rect 13973 -953 14051 -907
rect 14097 -953 14175 -907
rect 14221 -953 14299 -907
rect 14345 -953 14423 -907
rect 14469 -953 14547 -907
rect 14593 -953 14671 -907
rect 14717 -953 14795 -907
rect 14841 -953 14919 -907
rect 14965 -953 15043 -907
rect 15089 -953 15167 -907
rect 15213 -953 15291 -907
rect 15337 -953 15415 -907
rect 15461 -953 15539 -907
rect 15585 -953 15663 -907
rect 15709 -953 15787 -907
rect 15833 -953 15911 -907
rect 15957 -953 16035 -907
rect 16081 -953 16159 -907
rect 16205 -953 16283 -907
rect 16329 -953 16407 -907
rect 16453 -953 16531 -907
rect 16577 -953 16655 -907
rect 16701 -953 16779 -907
rect 16825 -953 16903 -907
rect 16949 -953 17027 -907
rect 17073 -953 17151 -907
rect 17197 -953 17275 -907
rect 17321 -953 17343 -907
rect -17343 -975 17343 -953
<< psubdiffcont >>
rect -17321 907 -17275 953
rect -17197 907 -17151 953
rect -17073 907 -17027 953
rect -16949 907 -16903 953
rect -16825 907 -16779 953
rect -16701 907 -16655 953
rect -16577 907 -16531 953
rect -16453 907 -16407 953
rect -16329 907 -16283 953
rect -16205 907 -16159 953
rect -16081 907 -16035 953
rect -15957 907 -15911 953
rect -15833 907 -15787 953
rect -15709 907 -15663 953
rect -15585 907 -15539 953
rect -15461 907 -15415 953
rect -15337 907 -15291 953
rect -15213 907 -15167 953
rect -15089 907 -15043 953
rect -14965 907 -14919 953
rect -14841 907 -14795 953
rect -14717 907 -14671 953
rect -14593 907 -14547 953
rect -14469 907 -14423 953
rect -14345 907 -14299 953
rect -14221 907 -14175 953
rect -14097 907 -14051 953
rect -13973 907 -13927 953
rect -13849 907 -13803 953
rect -13725 907 -13679 953
rect -13601 907 -13555 953
rect -13477 907 -13431 953
rect -13353 907 -13307 953
rect -13229 907 -13183 953
rect -13105 907 -13059 953
rect -12981 907 -12935 953
rect -12857 907 -12811 953
rect -12733 907 -12687 953
rect -12609 907 -12563 953
rect -12485 907 -12439 953
rect -12361 907 -12315 953
rect -12237 907 -12191 953
rect -12113 907 -12067 953
rect -11989 907 -11943 953
rect -11865 907 -11819 953
rect -11741 907 -11695 953
rect -11617 907 -11571 953
rect -11493 907 -11447 953
rect -11369 907 -11323 953
rect -11245 907 -11199 953
rect -11121 907 -11075 953
rect -10997 907 -10951 953
rect -10873 907 -10827 953
rect -10749 907 -10703 953
rect -10625 907 -10579 953
rect -10501 907 -10455 953
rect -10377 907 -10331 953
rect -10253 907 -10207 953
rect -10129 907 -10083 953
rect -10005 907 -9959 953
rect -9881 907 -9835 953
rect -9757 907 -9711 953
rect -9633 907 -9587 953
rect -9509 907 -9463 953
rect -9385 907 -9339 953
rect -9261 907 -9215 953
rect -9137 907 -9091 953
rect -9013 907 -8967 953
rect -8889 907 -8843 953
rect -8765 907 -8719 953
rect -8641 907 -8595 953
rect -8517 907 -8471 953
rect -8393 907 -8347 953
rect -8269 907 -8223 953
rect -8145 907 -8099 953
rect -8021 907 -7975 953
rect -7897 907 -7851 953
rect -7773 907 -7727 953
rect -7649 907 -7603 953
rect -7525 907 -7479 953
rect -7401 907 -7355 953
rect -7277 907 -7231 953
rect -7153 907 -7107 953
rect -7029 907 -6983 953
rect -6905 907 -6859 953
rect -6781 907 -6735 953
rect -6657 907 -6611 953
rect -6533 907 -6487 953
rect -6409 907 -6363 953
rect -6285 907 -6239 953
rect -6161 907 -6115 953
rect -6037 907 -5991 953
rect -5913 907 -5867 953
rect -5789 907 -5743 953
rect -5665 907 -5619 953
rect -5541 907 -5495 953
rect -5417 907 -5371 953
rect -5293 907 -5247 953
rect -5169 907 -5123 953
rect -5045 907 -4999 953
rect -4921 907 -4875 953
rect -4797 907 -4751 953
rect -4673 907 -4627 953
rect -4549 907 -4503 953
rect -4425 907 -4379 953
rect -4301 907 -4255 953
rect -4177 907 -4131 953
rect -4053 907 -4007 953
rect -3929 907 -3883 953
rect -3805 907 -3759 953
rect -3681 907 -3635 953
rect -3557 907 -3511 953
rect -3433 907 -3387 953
rect -3309 907 -3263 953
rect -3185 907 -3139 953
rect -3061 907 -3015 953
rect -2937 907 -2891 953
rect -2813 907 -2767 953
rect -2689 907 -2643 953
rect -2565 907 -2519 953
rect -2441 907 -2395 953
rect -2317 907 -2271 953
rect -2193 907 -2147 953
rect -2069 907 -2023 953
rect -1945 907 -1899 953
rect -1821 907 -1775 953
rect -1697 907 -1651 953
rect -1573 907 -1527 953
rect -1449 907 -1403 953
rect -1325 907 -1279 953
rect -1201 907 -1155 953
rect -1077 907 -1031 953
rect -953 907 -907 953
rect -829 907 -783 953
rect -705 907 -659 953
rect -581 907 -535 953
rect -457 907 -411 953
rect -333 907 -287 953
rect -209 907 -163 953
rect -85 907 -39 953
rect 39 907 85 953
rect 163 907 209 953
rect 287 907 333 953
rect 411 907 457 953
rect 535 907 581 953
rect 659 907 705 953
rect 783 907 829 953
rect 907 907 953 953
rect 1031 907 1077 953
rect 1155 907 1201 953
rect 1279 907 1325 953
rect 1403 907 1449 953
rect 1527 907 1573 953
rect 1651 907 1697 953
rect 1775 907 1821 953
rect 1899 907 1945 953
rect 2023 907 2069 953
rect 2147 907 2193 953
rect 2271 907 2317 953
rect 2395 907 2441 953
rect 2519 907 2565 953
rect 2643 907 2689 953
rect 2767 907 2813 953
rect 2891 907 2937 953
rect 3015 907 3061 953
rect 3139 907 3185 953
rect 3263 907 3309 953
rect 3387 907 3433 953
rect 3511 907 3557 953
rect 3635 907 3681 953
rect 3759 907 3805 953
rect 3883 907 3929 953
rect 4007 907 4053 953
rect 4131 907 4177 953
rect 4255 907 4301 953
rect 4379 907 4425 953
rect 4503 907 4549 953
rect 4627 907 4673 953
rect 4751 907 4797 953
rect 4875 907 4921 953
rect 4999 907 5045 953
rect 5123 907 5169 953
rect 5247 907 5293 953
rect 5371 907 5417 953
rect 5495 907 5541 953
rect 5619 907 5665 953
rect 5743 907 5789 953
rect 5867 907 5913 953
rect 5991 907 6037 953
rect 6115 907 6161 953
rect 6239 907 6285 953
rect 6363 907 6409 953
rect 6487 907 6533 953
rect 6611 907 6657 953
rect 6735 907 6781 953
rect 6859 907 6905 953
rect 6983 907 7029 953
rect 7107 907 7153 953
rect 7231 907 7277 953
rect 7355 907 7401 953
rect 7479 907 7525 953
rect 7603 907 7649 953
rect 7727 907 7773 953
rect 7851 907 7897 953
rect 7975 907 8021 953
rect 8099 907 8145 953
rect 8223 907 8269 953
rect 8347 907 8393 953
rect 8471 907 8517 953
rect 8595 907 8641 953
rect 8719 907 8765 953
rect 8843 907 8889 953
rect 8967 907 9013 953
rect 9091 907 9137 953
rect 9215 907 9261 953
rect 9339 907 9385 953
rect 9463 907 9509 953
rect 9587 907 9633 953
rect 9711 907 9757 953
rect 9835 907 9881 953
rect 9959 907 10005 953
rect 10083 907 10129 953
rect 10207 907 10253 953
rect 10331 907 10377 953
rect 10455 907 10501 953
rect 10579 907 10625 953
rect 10703 907 10749 953
rect 10827 907 10873 953
rect 10951 907 10997 953
rect 11075 907 11121 953
rect 11199 907 11245 953
rect 11323 907 11369 953
rect 11447 907 11493 953
rect 11571 907 11617 953
rect 11695 907 11741 953
rect 11819 907 11865 953
rect 11943 907 11989 953
rect 12067 907 12113 953
rect 12191 907 12237 953
rect 12315 907 12361 953
rect 12439 907 12485 953
rect 12563 907 12609 953
rect 12687 907 12733 953
rect 12811 907 12857 953
rect 12935 907 12981 953
rect 13059 907 13105 953
rect 13183 907 13229 953
rect 13307 907 13353 953
rect 13431 907 13477 953
rect 13555 907 13601 953
rect 13679 907 13725 953
rect 13803 907 13849 953
rect 13927 907 13973 953
rect 14051 907 14097 953
rect 14175 907 14221 953
rect 14299 907 14345 953
rect 14423 907 14469 953
rect 14547 907 14593 953
rect 14671 907 14717 953
rect 14795 907 14841 953
rect 14919 907 14965 953
rect 15043 907 15089 953
rect 15167 907 15213 953
rect 15291 907 15337 953
rect 15415 907 15461 953
rect 15539 907 15585 953
rect 15663 907 15709 953
rect 15787 907 15833 953
rect 15911 907 15957 953
rect 16035 907 16081 953
rect 16159 907 16205 953
rect 16283 907 16329 953
rect 16407 907 16453 953
rect 16531 907 16577 953
rect 16655 907 16701 953
rect 16779 907 16825 953
rect 16903 907 16949 953
rect 17027 907 17073 953
rect 17151 907 17197 953
rect 17275 907 17321 953
rect -17321 783 -17275 829
rect -17197 783 -17151 829
rect -17073 783 -17027 829
rect -16949 783 -16903 829
rect -16825 783 -16779 829
rect -16701 783 -16655 829
rect -16577 783 -16531 829
rect -16453 783 -16407 829
rect -16329 783 -16283 829
rect -16205 783 -16159 829
rect -16081 783 -16035 829
rect -15957 783 -15911 829
rect -15833 783 -15787 829
rect -15709 783 -15663 829
rect -15585 783 -15539 829
rect -15461 783 -15415 829
rect -15337 783 -15291 829
rect -15213 783 -15167 829
rect -15089 783 -15043 829
rect -14965 783 -14919 829
rect -14841 783 -14795 829
rect -14717 783 -14671 829
rect -14593 783 -14547 829
rect -14469 783 -14423 829
rect -14345 783 -14299 829
rect -14221 783 -14175 829
rect -14097 783 -14051 829
rect -13973 783 -13927 829
rect -13849 783 -13803 829
rect -13725 783 -13679 829
rect -13601 783 -13555 829
rect -13477 783 -13431 829
rect -13353 783 -13307 829
rect -13229 783 -13183 829
rect -13105 783 -13059 829
rect -12981 783 -12935 829
rect -12857 783 -12811 829
rect -12733 783 -12687 829
rect -12609 783 -12563 829
rect -12485 783 -12439 829
rect -12361 783 -12315 829
rect -12237 783 -12191 829
rect -12113 783 -12067 829
rect -11989 783 -11943 829
rect -11865 783 -11819 829
rect -11741 783 -11695 829
rect -11617 783 -11571 829
rect -11493 783 -11447 829
rect -11369 783 -11323 829
rect -11245 783 -11199 829
rect -11121 783 -11075 829
rect -10997 783 -10951 829
rect -10873 783 -10827 829
rect -10749 783 -10703 829
rect -10625 783 -10579 829
rect -10501 783 -10455 829
rect -10377 783 -10331 829
rect -10253 783 -10207 829
rect -10129 783 -10083 829
rect -10005 783 -9959 829
rect -9881 783 -9835 829
rect -9757 783 -9711 829
rect -9633 783 -9587 829
rect -9509 783 -9463 829
rect -9385 783 -9339 829
rect -9261 783 -9215 829
rect -9137 783 -9091 829
rect -9013 783 -8967 829
rect -8889 783 -8843 829
rect -8765 783 -8719 829
rect -8641 783 -8595 829
rect -8517 783 -8471 829
rect -8393 783 -8347 829
rect -8269 783 -8223 829
rect -8145 783 -8099 829
rect -8021 783 -7975 829
rect -7897 783 -7851 829
rect -7773 783 -7727 829
rect -7649 783 -7603 829
rect -7525 783 -7479 829
rect -7401 783 -7355 829
rect -7277 783 -7231 829
rect -7153 783 -7107 829
rect -7029 783 -6983 829
rect -6905 783 -6859 829
rect -6781 783 -6735 829
rect -6657 783 -6611 829
rect -6533 783 -6487 829
rect -6409 783 -6363 829
rect -6285 783 -6239 829
rect -6161 783 -6115 829
rect -6037 783 -5991 829
rect -5913 783 -5867 829
rect -5789 783 -5743 829
rect -5665 783 -5619 829
rect -5541 783 -5495 829
rect -5417 783 -5371 829
rect -5293 783 -5247 829
rect -5169 783 -5123 829
rect -5045 783 -4999 829
rect -4921 783 -4875 829
rect -4797 783 -4751 829
rect -4673 783 -4627 829
rect -4549 783 -4503 829
rect -4425 783 -4379 829
rect -4301 783 -4255 829
rect -4177 783 -4131 829
rect -4053 783 -4007 829
rect -3929 783 -3883 829
rect -3805 783 -3759 829
rect -3681 783 -3635 829
rect -3557 783 -3511 829
rect -3433 783 -3387 829
rect -3309 783 -3263 829
rect -3185 783 -3139 829
rect -3061 783 -3015 829
rect -2937 783 -2891 829
rect -2813 783 -2767 829
rect -2689 783 -2643 829
rect -2565 783 -2519 829
rect -2441 783 -2395 829
rect -2317 783 -2271 829
rect -2193 783 -2147 829
rect -2069 783 -2023 829
rect -1945 783 -1899 829
rect -1821 783 -1775 829
rect -1697 783 -1651 829
rect -1573 783 -1527 829
rect -1449 783 -1403 829
rect -1325 783 -1279 829
rect -1201 783 -1155 829
rect -1077 783 -1031 829
rect -953 783 -907 829
rect -829 783 -783 829
rect -705 783 -659 829
rect -581 783 -535 829
rect -457 783 -411 829
rect -333 783 -287 829
rect -209 783 -163 829
rect -85 783 -39 829
rect 39 783 85 829
rect 163 783 209 829
rect 287 783 333 829
rect 411 783 457 829
rect 535 783 581 829
rect 659 783 705 829
rect 783 783 829 829
rect 907 783 953 829
rect 1031 783 1077 829
rect 1155 783 1201 829
rect 1279 783 1325 829
rect 1403 783 1449 829
rect 1527 783 1573 829
rect 1651 783 1697 829
rect 1775 783 1821 829
rect 1899 783 1945 829
rect 2023 783 2069 829
rect 2147 783 2193 829
rect 2271 783 2317 829
rect 2395 783 2441 829
rect 2519 783 2565 829
rect 2643 783 2689 829
rect 2767 783 2813 829
rect 2891 783 2937 829
rect 3015 783 3061 829
rect 3139 783 3185 829
rect 3263 783 3309 829
rect 3387 783 3433 829
rect 3511 783 3557 829
rect 3635 783 3681 829
rect 3759 783 3805 829
rect 3883 783 3929 829
rect 4007 783 4053 829
rect 4131 783 4177 829
rect 4255 783 4301 829
rect 4379 783 4425 829
rect 4503 783 4549 829
rect 4627 783 4673 829
rect 4751 783 4797 829
rect 4875 783 4921 829
rect 4999 783 5045 829
rect 5123 783 5169 829
rect 5247 783 5293 829
rect 5371 783 5417 829
rect 5495 783 5541 829
rect 5619 783 5665 829
rect 5743 783 5789 829
rect 5867 783 5913 829
rect 5991 783 6037 829
rect 6115 783 6161 829
rect 6239 783 6285 829
rect 6363 783 6409 829
rect 6487 783 6533 829
rect 6611 783 6657 829
rect 6735 783 6781 829
rect 6859 783 6905 829
rect 6983 783 7029 829
rect 7107 783 7153 829
rect 7231 783 7277 829
rect 7355 783 7401 829
rect 7479 783 7525 829
rect 7603 783 7649 829
rect 7727 783 7773 829
rect 7851 783 7897 829
rect 7975 783 8021 829
rect 8099 783 8145 829
rect 8223 783 8269 829
rect 8347 783 8393 829
rect 8471 783 8517 829
rect 8595 783 8641 829
rect 8719 783 8765 829
rect 8843 783 8889 829
rect 8967 783 9013 829
rect 9091 783 9137 829
rect 9215 783 9261 829
rect 9339 783 9385 829
rect 9463 783 9509 829
rect 9587 783 9633 829
rect 9711 783 9757 829
rect 9835 783 9881 829
rect 9959 783 10005 829
rect 10083 783 10129 829
rect 10207 783 10253 829
rect 10331 783 10377 829
rect 10455 783 10501 829
rect 10579 783 10625 829
rect 10703 783 10749 829
rect 10827 783 10873 829
rect 10951 783 10997 829
rect 11075 783 11121 829
rect 11199 783 11245 829
rect 11323 783 11369 829
rect 11447 783 11493 829
rect 11571 783 11617 829
rect 11695 783 11741 829
rect 11819 783 11865 829
rect 11943 783 11989 829
rect 12067 783 12113 829
rect 12191 783 12237 829
rect 12315 783 12361 829
rect 12439 783 12485 829
rect 12563 783 12609 829
rect 12687 783 12733 829
rect 12811 783 12857 829
rect 12935 783 12981 829
rect 13059 783 13105 829
rect 13183 783 13229 829
rect 13307 783 13353 829
rect 13431 783 13477 829
rect 13555 783 13601 829
rect 13679 783 13725 829
rect 13803 783 13849 829
rect 13927 783 13973 829
rect 14051 783 14097 829
rect 14175 783 14221 829
rect 14299 783 14345 829
rect 14423 783 14469 829
rect 14547 783 14593 829
rect 14671 783 14717 829
rect 14795 783 14841 829
rect 14919 783 14965 829
rect 15043 783 15089 829
rect 15167 783 15213 829
rect 15291 783 15337 829
rect 15415 783 15461 829
rect 15539 783 15585 829
rect 15663 783 15709 829
rect 15787 783 15833 829
rect 15911 783 15957 829
rect 16035 783 16081 829
rect 16159 783 16205 829
rect 16283 783 16329 829
rect 16407 783 16453 829
rect 16531 783 16577 829
rect 16655 783 16701 829
rect 16779 783 16825 829
rect 16903 783 16949 829
rect 17027 783 17073 829
rect 17151 783 17197 829
rect 17275 783 17321 829
rect -17321 659 -17275 705
rect -17197 659 -17151 705
rect -17073 659 -17027 705
rect -16949 659 -16903 705
rect -16825 659 -16779 705
rect -16701 659 -16655 705
rect -16577 659 -16531 705
rect -16453 659 -16407 705
rect -16329 659 -16283 705
rect -16205 659 -16159 705
rect -16081 659 -16035 705
rect -15957 659 -15911 705
rect -15833 659 -15787 705
rect -15709 659 -15663 705
rect -15585 659 -15539 705
rect -15461 659 -15415 705
rect -15337 659 -15291 705
rect -15213 659 -15167 705
rect -15089 659 -15043 705
rect -14965 659 -14919 705
rect -14841 659 -14795 705
rect -14717 659 -14671 705
rect -14593 659 -14547 705
rect -14469 659 -14423 705
rect -14345 659 -14299 705
rect -14221 659 -14175 705
rect -14097 659 -14051 705
rect -13973 659 -13927 705
rect -13849 659 -13803 705
rect -13725 659 -13679 705
rect -13601 659 -13555 705
rect -13477 659 -13431 705
rect -13353 659 -13307 705
rect -13229 659 -13183 705
rect -13105 659 -13059 705
rect -12981 659 -12935 705
rect -12857 659 -12811 705
rect -12733 659 -12687 705
rect -12609 659 -12563 705
rect -12485 659 -12439 705
rect -12361 659 -12315 705
rect -12237 659 -12191 705
rect -12113 659 -12067 705
rect -11989 659 -11943 705
rect -11865 659 -11819 705
rect -11741 659 -11695 705
rect -11617 659 -11571 705
rect -11493 659 -11447 705
rect -11369 659 -11323 705
rect -11245 659 -11199 705
rect -11121 659 -11075 705
rect -10997 659 -10951 705
rect -10873 659 -10827 705
rect -10749 659 -10703 705
rect -10625 659 -10579 705
rect -10501 659 -10455 705
rect -10377 659 -10331 705
rect -10253 659 -10207 705
rect -10129 659 -10083 705
rect -10005 659 -9959 705
rect -9881 659 -9835 705
rect -9757 659 -9711 705
rect -9633 659 -9587 705
rect -9509 659 -9463 705
rect -9385 659 -9339 705
rect -9261 659 -9215 705
rect -9137 659 -9091 705
rect -9013 659 -8967 705
rect -8889 659 -8843 705
rect -8765 659 -8719 705
rect -8641 659 -8595 705
rect -8517 659 -8471 705
rect -8393 659 -8347 705
rect -8269 659 -8223 705
rect -8145 659 -8099 705
rect -8021 659 -7975 705
rect -7897 659 -7851 705
rect -7773 659 -7727 705
rect -7649 659 -7603 705
rect -7525 659 -7479 705
rect -7401 659 -7355 705
rect -7277 659 -7231 705
rect -7153 659 -7107 705
rect -7029 659 -6983 705
rect -6905 659 -6859 705
rect -6781 659 -6735 705
rect -6657 659 -6611 705
rect -6533 659 -6487 705
rect -6409 659 -6363 705
rect -6285 659 -6239 705
rect -6161 659 -6115 705
rect -6037 659 -5991 705
rect -5913 659 -5867 705
rect -5789 659 -5743 705
rect -5665 659 -5619 705
rect -5541 659 -5495 705
rect -5417 659 -5371 705
rect -5293 659 -5247 705
rect -5169 659 -5123 705
rect -5045 659 -4999 705
rect -4921 659 -4875 705
rect -4797 659 -4751 705
rect -4673 659 -4627 705
rect -4549 659 -4503 705
rect -4425 659 -4379 705
rect -4301 659 -4255 705
rect -4177 659 -4131 705
rect -4053 659 -4007 705
rect -3929 659 -3883 705
rect -3805 659 -3759 705
rect -3681 659 -3635 705
rect -3557 659 -3511 705
rect -3433 659 -3387 705
rect -3309 659 -3263 705
rect -3185 659 -3139 705
rect -3061 659 -3015 705
rect -2937 659 -2891 705
rect -2813 659 -2767 705
rect -2689 659 -2643 705
rect -2565 659 -2519 705
rect -2441 659 -2395 705
rect -2317 659 -2271 705
rect -2193 659 -2147 705
rect -2069 659 -2023 705
rect -1945 659 -1899 705
rect -1821 659 -1775 705
rect -1697 659 -1651 705
rect -1573 659 -1527 705
rect -1449 659 -1403 705
rect -1325 659 -1279 705
rect -1201 659 -1155 705
rect -1077 659 -1031 705
rect -953 659 -907 705
rect -829 659 -783 705
rect -705 659 -659 705
rect -581 659 -535 705
rect -457 659 -411 705
rect -333 659 -287 705
rect -209 659 -163 705
rect -85 659 -39 705
rect 39 659 85 705
rect 163 659 209 705
rect 287 659 333 705
rect 411 659 457 705
rect 535 659 581 705
rect 659 659 705 705
rect 783 659 829 705
rect 907 659 953 705
rect 1031 659 1077 705
rect 1155 659 1201 705
rect 1279 659 1325 705
rect 1403 659 1449 705
rect 1527 659 1573 705
rect 1651 659 1697 705
rect 1775 659 1821 705
rect 1899 659 1945 705
rect 2023 659 2069 705
rect 2147 659 2193 705
rect 2271 659 2317 705
rect 2395 659 2441 705
rect 2519 659 2565 705
rect 2643 659 2689 705
rect 2767 659 2813 705
rect 2891 659 2937 705
rect 3015 659 3061 705
rect 3139 659 3185 705
rect 3263 659 3309 705
rect 3387 659 3433 705
rect 3511 659 3557 705
rect 3635 659 3681 705
rect 3759 659 3805 705
rect 3883 659 3929 705
rect 4007 659 4053 705
rect 4131 659 4177 705
rect 4255 659 4301 705
rect 4379 659 4425 705
rect 4503 659 4549 705
rect 4627 659 4673 705
rect 4751 659 4797 705
rect 4875 659 4921 705
rect 4999 659 5045 705
rect 5123 659 5169 705
rect 5247 659 5293 705
rect 5371 659 5417 705
rect 5495 659 5541 705
rect 5619 659 5665 705
rect 5743 659 5789 705
rect 5867 659 5913 705
rect 5991 659 6037 705
rect 6115 659 6161 705
rect 6239 659 6285 705
rect 6363 659 6409 705
rect 6487 659 6533 705
rect 6611 659 6657 705
rect 6735 659 6781 705
rect 6859 659 6905 705
rect 6983 659 7029 705
rect 7107 659 7153 705
rect 7231 659 7277 705
rect 7355 659 7401 705
rect 7479 659 7525 705
rect 7603 659 7649 705
rect 7727 659 7773 705
rect 7851 659 7897 705
rect 7975 659 8021 705
rect 8099 659 8145 705
rect 8223 659 8269 705
rect 8347 659 8393 705
rect 8471 659 8517 705
rect 8595 659 8641 705
rect 8719 659 8765 705
rect 8843 659 8889 705
rect 8967 659 9013 705
rect 9091 659 9137 705
rect 9215 659 9261 705
rect 9339 659 9385 705
rect 9463 659 9509 705
rect 9587 659 9633 705
rect 9711 659 9757 705
rect 9835 659 9881 705
rect 9959 659 10005 705
rect 10083 659 10129 705
rect 10207 659 10253 705
rect 10331 659 10377 705
rect 10455 659 10501 705
rect 10579 659 10625 705
rect 10703 659 10749 705
rect 10827 659 10873 705
rect 10951 659 10997 705
rect 11075 659 11121 705
rect 11199 659 11245 705
rect 11323 659 11369 705
rect 11447 659 11493 705
rect 11571 659 11617 705
rect 11695 659 11741 705
rect 11819 659 11865 705
rect 11943 659 11989 705
rect 12067 659 12113 705
rect 12191 659 12237 705
rect 12315 659 12361 705
rect 12439 659 12485 705
rect 12563 659 12609 705
rect 12687 659 12733 705
rect 12811 659 12857 705
rect 12935 659 12981 705
rect 13059 659 13105 705
rect 13183 659 13229 705
rect 13307 659 13353 705
rect 13431 659 13477 705
rect 13555 659 13601 705
rect 13679 659 13725 705
rect 13803 659 13849 705
rect 13927 659 13973 705
rect 14051 659 14097 705
rect 14175 659 14221 705
rect 14299 659 14345 705
rect 14423 659 14469 705
rect 14547 659 14593 705
rect 14671 659 14717 705
rect 14795 659 14841 705
rect 14919 659 14965 705
rect 15043 659 15089 705
rect 15167 659 15213 705
rect 15291 659 15337 705
rect 15415 659 15461 705
rect 15539 659 15585 705
rect 15663 659 15709 705
rect 15787 659 15833 705
rect 15911 659 15957 705
rect 16035 659 16081 705
rect 16159 659 16205 705
rect 16283 659 16329 705
rect 16407 659 16453 705
rect 16531 659 16577 705
rect 16655 659 16701 705
rect 16779 659 16825 705
rect 16903 659 16949 705
rect 17027 659 17073 705
rect 17151 659 17197 705
rect 17275 659 17321 705
rect -17321 535 -17275 581
rect -17197 535 -17151 581
rect -17073 535 -17027 581
rect -16949 535 -16903 581
rect -16825 535 -16779 581
rect -16701 535 -16655 581
rect -16577 535 -16531 581
rect -16453 535 -16407 581
rect -16329 535 -16283 581
rect -16205 535 -16159 581
rect -16081 535 -16035 581
rect -15957 535 -15911 581
rect -15833 535 -15787 581
rect -15709 535 -15663 581
rect -15585 535 -15539 581
rect -15461 535 -15415 581
rect -15337 535 -15291 581
rect -15213 535 -15167 581
rect -15089 535 -15043 581
rect -14965 535 -14919 581
rect -14841 535 -14795 581
rect -14717 535 -14671 581
rect -14593 535 -14547 581
rect -14469 535 -14423 581
rect -14345 535 -14299 581
rect -14221 535 -14175 581
rect -14097 535 -14051 581
rect -13973 535 -13927 581
rect -13849 535 -13803 581
rect -13725 535 -13679 581
rect -13601 535 -13555 581
rect -13477 535 -13431 581
rect -13353 535 -13307 581
rect -13229 535 -13183 581
rect -13105 535 -13059 581
rect -12981 535 -12935 581
rect -12857 535 -12811 581
rect -12733 535 -12687 581
rect -12609 535 -12563 581
rect -12485 535 -12439 581
rect -12361 535 -12315 581
rect -12237 535 -12191 581
rect -12113 535 -12067 581
rect -11989 535 -11943 581
rect -11865 535 -11819 581
rect -11741 535 -11695 581
rect -11617 535 -11571 581
rect -11493 535 -11447 581
rect -11369 535 -11323 581
rect -11245 535 -11199 581
rect -11121 535 -11075 581
rect -10997 535 -10951 581
rect -10873 535 -10827 581
rect -10749 535 -10703 581
rect -10625 535 -10579 581
rect -10501 535 -10455 581
rect -10377 535 -10331 581
rect -10253 535 -10207 581
rect -10129 535 -10083 581
rect -10005 535 -9959 581
rect -9881 535 -9835 581
rect -9757 535 -9711 581
rect -9633 535 -9587 581
rect -9509 535 -9463 581
rect -9385 535 -9339 581
rect -9261 535 -9215 581
rect -9137 535 -9091 581
rect -9013 535 -8967 581
rect -8889 535 -8843 581
rect -8765 535 -8719 581
rect -8641 535 -8595 581
rect -8517 535 -8471 581
rect -8393 535 -8347 581
rect -8269 535 -8223 581
rect -8145 535 -8099 581
rect -8021 535 -7975 581
rect -7897 535 -7851 581
rect -7773 535 -7727 581
rect -7649 535 -7603 581
rect -7525 535 -7479 581
rect -7401 535 -7355 581
rect -7277 535 -7231 581
rect -7153 535 -7107 581
rect -7029 535 -6983 581
rect -6905 535 -6859 581
rect -6781 535 -6735 581
rect -6657 535 -6611 581
rect -6533 535 -6487 581
rect -6409 535 -6363 581
rect -6285 535 -6239 581
rect -6161 535 -6115 581
rect -6037 535 -5991 581
rect -5913 535 -5867 581
rect -5789 535 -5743 581
rect -5665 535 -5619 581
rect -5541 535 -5495 581
rect -5417 535 -5371 581
rect -5293 535 -5247 581
rect -5169 535 -5123 581
rect -5045 535 -4999 581
rect -4921 535 -4875 581
rect -4797 535 -4751 581
rect -4673 535 -4627 581
rect -4549 535 -4503 581
rect -4425 535 -4379 581
rect -4301 535 -4255 581
rect -4177 535 -4131 581
rect -4053 535 -4007 581
rect -3929 535 -3883 581
rect -3805 535 -3759 581
rect -3681 535 -3635 581
rect -3557 535 -3511 581
rect -3433 535 -3387 581
rect -3309 535 -3263 581
rect -3185 535 -3139 581
rect -3061 535 -3015 581
rect -2937 535 -2891 581
rect -2813 535 -2767 581
rect -2689 535 -2643 581
rect -2565 535 -2519 581
rect -2441 535 -2395 581
rect -2317 535 -2271 581
rect -2193 535 -2147 581
rect -2069 535 -2023 581
rect -1945 535 -1899 581
rect -1821 535 -1775 581
rect -1697 535 -1651 581
rect -1573 535 -1527 581
rect -1449 535 -1403 581
rect -1325 535 -1279 581
rect -1201 535 -1155 581
rect -1077 535 -1031 581
rect -953 535 -907 581
rect -829 535 -783 581
rect -705 535 -659 581
rect -581 535 -535 581
rect -457 535 -411 581
rect -333 535 -287 581
rect -209 535 -163 581
rect -85 535 -39 581
rect 39 535 85 581
rect 163 535 209 581
rect 287 535 333 581
rect 411 535 457 581
rect 535 535 581 581
rect 659 535 705 581
rect 783 535 829 581
rect 907 535 953 581
rect 1031 535 1077 581
rect 1155 535 1201 581
rect 1279 535 1325 581
rect 1403 535 1449 581
rect 1527 535 1573 581
rect 1651 535 1697 581
rect 1775 535 1821 581
rect 1899 535 1945 581
rect 2023 535 2069 581
rect 2147 535 2193 581
rect 2271 535 2317 581
rect 2395 535 2441 581
rect 2519 535 2565 581
rect 2643 535 2689 581
rect 2767 535 2813 581
rect 2891 535 2937 581
rect 3015 535 3061 581
rect 3139 535 3185 581
rect 3263 535 3309 581
rect 3387 535 3433 581
rect 3511 535 3557 581
rect 3635 535 3681 581
rect 3759 535 3805 581
rect 3883 535 3929 581
rect 4007 535 4053 581
rect 4131 535 4177 581
rect 4255 535 4301 581
rect 4379 535 4425 581
rect 4503 535 4549 581
rect 4627 535 4673 581
rect 4751 535 4797 581
rect 4875 535 4921 581
rect 4999 535 5045 581
rect 5123 535 5169 581
rect 5247 535 5293 581
rect 5371 535 5417 581
rect 5495 535 5541 581
rect 5619 535 5665 581
rect 5743 535 5789 581
rect 5867 535 5913 581
rect 5991 535 6037 581
rect 6115 535 6161 581
rect 6239 535 6285 581
rect 6363 535 6409 581
rect 6487 535 6533 581
rect 6611 535 6657 581
rect 6735 535 6781 581
rect 6859 535 6905 581
rect 6983 535 7029 581
rect 7107 535 7153 581
rect 7231 535 7277 581
rect 7355 535 7401 581
rect 7479 535 7525 581
rect 7603 535 7649 581
rect 7727 535 7773 581
rect 7851 535 7897 581
rect 7975 535 8021 581
rect 8099 535 8145 581
rect 8223 535 8269 581
rect 8347 535 8393 581
rect 8471 535 8517 581
rect 8595 535 8641 581
rect 8719 535 8765 581
rect 8843 535 8889 581
rect 8967 535 9013 581
rect 9091 535 9137 581
rect 9215 535 9261 581
rect 9339 535 9385 581
rect 9463 535 9509 581
rect 9587 535 9633 581
rect 9711 535 9757 581
rect 9835 535 9881 581
rect 9959 535 10005 581
rect 10083 535 10129 581
rect 10207 535 10253 581
rect 10331 535 10377 581
rect 10455 535 10501 581
rect 10579 535 10625 581
rect 10703 535 10749 581
rect 10827 535 10873 581
rect 10951 535 10997 581
rect 11075 535 11121 581
rect 11199 535 11245 581
rect 11323 535 11369 581
rect 11447 535 11493 581
rect 11571 535 11617 581
rect 11695 535 11741 581
rect 11819 535 11865 581
rect 11943 535 11989 581
rect 12067 535 12113 581
rect 12191 535 12237 581
rect 12315 535 12361 581
rect 12439 535 12485 581
rect 12563 535 12609 581
rect 12687 535 12733 581
rect 12811 535 12857 581
rect 12935 535 12981 581
rect 13059 535 13105 581
rect 13183 535 13229 581
rect 13307 535 13353 581
rect 13431 535 13477 581
rect 13555 535 13601 581
rect 13679 535 13725 581
rect 13803 535 13849 581
rect 13927 535 13973 581
rect 14051 535 14097 581
rect 14175 535 14221 581
rect 14299 535 14345 581
rect 14423 535 14469 581
rect 14547 535 14593 581
rect 14671 535 14717 581
rect 14795 535 14841 581
rect 14919 535 14965 581
rect 15043 535 15089 581
rect 15167 535 15213 581
rect 15291 535 15337 581
rect 15415 535 15461 581
rect 15539 535 15585 581
rect 15663 535 15709 581
rect 15787 535 15833 581
rect 15911 535 15957 581
rect 16035 535 16081 581
rect 16159 535 16205 581
rect 16283 535 16329 581
rect 16407 535 16453 581
rect 16531 535 16577 581
rect 16655 535 16701 581
rect 16779 535 16825 581
rect 16903 535 16949 581
rect 17027 535 17073 581
rect 17151 535 17197 581
rect 17275 535 17321 581
rect -17321 411 -17275 457
rect -17197 411 -17151 457
rect -17073 411 -17027 457
rect -16949 411 -16903 457
rect -16825 411 -16779 457
rect -16701 411 -16655 457
rect -16577 411 -16531 457
rect -16453 411 -16407 457
rect -16329 411 -16283 457
rect -16205 411 -16159 457
rect -16081 411 -16035 457
rect -15957 411 -15911 457
rect -15833 411 -15787 457
rect -15709 411 -15663 457
rect -15585 411 -15539 457
rect -15461 411 -15415 457
rect -15337 411 -15291 457
rect -15213 411 -15167 457
rect -15089 411 -15043 457
rect -14965 411 -14919 457
rect -14841 411 -14795 457
rect -14717 411 -14671 457
rect -14593 411 -14547 457
rect -14469 411 -14423 457
rect -14345 411 -14299 457
rect -14221 411 -14175 457
rect -14097 411 -14051 457
rect -13973 411 -13927 457
rect -13849 411 -13803 457
rect -13725 411 -13679 457
rect -13601 411 -13555 457
rect -13477 411 -13431 457
rect -13353 411 -13307 457
rect -13229 411 -13183 457
rect -13105 411 -13059 457
rect -12981 411 -12935 457
rect -12857 411 -12811 457
rect -12733 411 -12687 457
rect -12609 411 -12563 457
rect -12485 411 -12439 457
rect -12361 411 -12315 457
rect -12237 411 -12191 457
rect -12113 411 -12067 457
rect -11989 411 -11943 457
rect -11865 411 -11819 457
rect -11741 411 -11695 457
rect -11617 411 -11571 457
rect -11493 411 -11447 457
rect -11369 411 -11323 457
rect -11245 411 -11199 457
rect -11121 411 -11075 457
rect -10997 411 -10951 457
rect -10873 411 -10827 457
rect -10749 411 -10703 457
rect -10625 411 -10579 457
rect -10501 411 -10455 457
rect -10377 411 -10331 457
rect -10253 411 -10207 457
rect -10129 411 -10083 457
rect -10005 411 -9959 457
rect -9881 411 -9835 457
rect -9757 411 -9711 457
rect -9633 411 -9587 457
rect -9509 411 -9463 457
rect -9385 411 -9339 457
rect -9261 411 -9215 457
rect -9137 411 -9091 457
rect -9013 411 -8967 457
rect -8889 411 -8843 457
rect -8765 411 -8719 457
rect -8641 411 -8595 457
rect -8517 411 -8471 457
rect -8393 411 -8347 457
rect -8269 411 -8223 457
rect -8145 411 -8099 457
rect -8021 411 -7975 457
rect -7897 411 -7851 457
rect -7773 411 -7727 457
rect -7649 411 -7603 457
rect -7525 411 -7479 457
rect -7401 411 -7355 457
rect -7277 411 -7231 457
rect -7153 411 -7107 457
rect -7029 411 -6983 457
rect -6905 411 -6859 457
rect -6781 411 -6735 457
rect -6657 411 -6611 457
rect -6533 411 -6487 457
rect -6409 411 -6363 457
rect -6285 411 -6239 457
rect -6161 411 -6115 457
rect -6037 411 -5991 457
rect -5913 411 -5867 457
rect -5789 411 -5743 457
rect -5665 411 -5619 457
rect -5541 411 -5495 457
rect -5417 411 -5371 457
rect -5293 411 -5247 457
rect -5169 411 -5123 457
rect -5045 411 -4999 457
rect -4921 411 -4875 457
rect -4797 411 -4751 457
rect -4673 411 -4627 457
rect -4549 411 -4503 457
rect -4425 411 -4379 457
rect -4301 411 -4255 457
rect -4177 411 -4131 457
rect -4053 411 -4007 457
rect -3929 411 -3883 457
rect -3805 411 -3759 457
rect -3681 411 -3635 457
rect -3557 411 -3511 457
rect -3433 411 -3387 457
rect -3309 411 -3263 457
rect -3185 411 -3139 457
rect -3061 411 -3015 457
rect -2937 411 -2891 457
rect -2813 411 -2767 457
rect -2689 411 -2643 457
rect -2565 411 -2519 457
rect -2441 411 -2395 457
rect -2317 411 -2271 457
rect -2193 411 -2147 457
rect -2069 411 -2023 457
rect -1945 411 -1899 457
rect -1821 411 -1775 457
rect -1697 411 -1651 457
rect -1573 411 -1527 457
rect -1449 411 -1403 457
rect -1325 411 -1279 457
rect -1201 411 -1155 457
rect -1077 411 -1031 457
rect -953 411 -907 457
rect -829 411 -783 457
rect -705 411 -659 457
rect -581 411 -535 457
rect -457 411 -411 457
rect -333 411 -287 457
rect -209 411 -163 457
rect -85 411 -39 457
rect 39 411 85 457
rect 163 411 209 457
rect 287 411 333 457
rect 411 411 457 457
rect 535 411 581 457
rect 659 411 705 457
rect 783 411 829 457
rect 907 411 953 457
rect 1031 411 1077 457
rect 1155 411 1201 457
rect 1279 411 1325 457
rect 1403 411 1449 457
rect 1527 411 1573 457
rect 1651 411 1697 457
rect 1775 411 1821 457
rect 1899 411 1945 457
rect 2023 411 2069 457
rect 2147 411 2193 457
rect 2271 411 2317 457
rect 2395 411 2441 457
rect 2519 411 2565 457
rect 2643 411 2689 457
rect 2767 411 2813 457
rect 2891 411 2937 457
rect 3015 411 3061 457
rect 3139 411 3185 457
rect 3263 411 3309 457
rect 3387 411 3433 457
rect 3511 411 3557 457
rect 3635 411 3681 457
rect 3759 411 3805 457
rect 3883 411 3929 457
rect 4007 411 4053 457
rect 4131 411 4177 457
rect 4255 411 4301 457
rect 4379 411 4425 457
rect 4503 411 4549 457
rect 4627 411 4673 457
rect 4751 411 4797 457
rect 4875 411 4921 457
rect 4999 411 5045 457
rect 5123 411 5169 457
rect 5247 411 5293 457
rect 5371 411 5417 457
rect 5495 411 5541 457
rect 5619 411 5665 457
rect 5743 411 5789 457
rect 5867 411 5913 457
rect 5991 411 6037 457
rect 6115 411 6161 457
rect 6239 411 6285 457
rect 6363 411 6409 457
rect 6487 411 6533 457
rect 6611 411 6657 457
rect 6735 411 6781 457
rect 6859 411 6905 457
rect 6983 411 7029 457
rect 7107 411 7153 457
rect 7231 411 7277 457
rect 7355 411 7401 457
rect 7479 411 7525 457
rect 7603 411 7649 457
rect 7727 411 7773 457
rect 7851 411 7897 457
rect 7975 411 8021 457
rect 8099 411 8145 457
rect 8223 411 8269 457
rect 8347 411 8393 457
rect 8471 411 8517 457
rect 8595 411 8641 457
rect 8719 411 8765 457
rect 8843 411 8889 457
rect 8967 411 9013 457
rect 9091 411 9137 457
rect 9215 411 9261 457
rect 9339 411 9385 457
rect 9463 411 9509 457
rect 9587 411 9633 457
rect 9711 411 9757 457
rect 9835 411 9881 457
rect 9959 411 10005 457
rect 10083 411 10129 457
rect 10207 411 10253 457
rect 10331 411 10377 457
rect 10455 411 10501 457
rect 10579 411 10625 457
rect 10703 411 10749 457
rect 10827 411 10873 457
rect 10951 411 10997 457
rect 11075 411 11121 457
rect 11199 411 11245 457
rect 11323 411 11369 457
rect 11447 411 11493 457
rect 11571 411 11617 457
rect 11695 411 11741 457
rect 11819 411 11865 457
rect 11943 411 11989 457
rect 12067 411 12113 457
rect 12191 411 12237 457
rect 12315 411 12361 457
rect 12439 411 12485 457
rect 12563 411 12609 457
rect 12687 411 12733 457
rect 12811 411 12857 457
rect 12935 411 12981 457
rect 13059 411 13105 457
rect 13183 411 13229 457
rect 13307 411 13353 457
rect 13431 411 13477 457
rect 13555 411 13601 457
rect 13679 411 13725 457
rect 13803 411 13849 457
rect 13927 411 13973 457
rect 14051 411 14097 457
rect 14175 411 14221 457
rect 14299 411 14345 457
rect 14423 411 14469 457
rect 14547 411 14593 457
rect 14671 411 14717 457
rect 14795 411 14841 457
rect 14919 411 14965 457
rect 15043 411 15089 457
rect 15167 411 15213 457
rect 15291 411 15337 457
rect 15415 411 15461 457
rect 15539 411 15585 457
rect 15663 411 15709 457
rect 15787 411 15833 457
rect 15911 411 15957 457
rect 16035 411 16081 457
rect 16159 411 16205 457
rect 16283 411 16329 457
rect 16407 411 16453 457
rect 16531 411 16577 457
rect 16655 411 16701 457
rect 16779 411 16825 457
rect 16903 411 16949 457
rect 17027 411 17073 457
rect 17151 411 17197 457
rect 17275 411 17321 457
rect -17321 287 -17275 333
rect -17197 287 -17151 333
rect -17073 287 -17027 333
rect -16949 287 -16903 333
rect -16825 287 -16779 333
rect -16701 287 -16655 333
rect -16577 287 -16531 333
rect -16453 287 -16407 333
rect -16329 287 -16283 333
rect -16205 287 -16159 333
rect -16081 287 -16035 333
rect -15957 287 -15911 333
rect -15833 287 -15787 333
rect -15709 287 -15663 333
rect -15585 287 -15539 333
rect -15461 287 -15415 333
rect -15337 287 -15291 333
rect -15213 287 -15167 333
rect -15089 287 -15043 333
rect -14965 287 -14919 333
rect -14841 287 -14795 333
rect -14717 287 -14671 333
rect -14593 287 -14547 333
rect -14469 287 -14423 333
rect -14345 287 -14299 333
rect -14221 287 -14175 333
rect -14097 287 -14051 333
rect -13973 287 -13927 333
rect -13849 287 -13803 333
rect -13725 287 -13679 333
rect -13601 287 -13555 333
rect -13477 287 -13431 333
rect -13353 287 -13307 333
rect -13229 287 -13183 333
rect -13105 287 -13059 333
rect -12981 287 -12935 333
rect -12857 287 -12811 333
rect -12733 287 -12687 333
rect -12609 287 -12563 333
rect -12485 287 -12439 333
rect -12361 287 -12315 333
rect -12237 287 -12191 333
rect -12113 287 -12067 333
rect -11989 287 -11943 333
rect -11865 287 -11819 333
rect -11741 287 -11695 333
rect -11617 287 -11571 333
rect -11493 287 -11447 333
rect -11369 287 -11323 333
rect -11245 287 -11199 333
rect -11121 287 -11075 333
rect -10997 287 -10951 333
rect -10873 287 -10827 333
rect -10749 287 -10703 333
rect -10625 287 -10579 333
rect -10501 287 -10455 333
rect -10377 287 -10331 333
rect -10253 287 -10207 333
rect -10129 287 -10083 333
rect -10005 287 -9959 333
rect -9881 287 -9835 333
rect -9757 287 -9711 333
rect -9633 287 -9587 333
rect -9509 287 -9463 333
rect -9385 287 -9339 333
rect -9261 287 -9215 333
rect -9137 287 -9091 333
rect -9013 287 -8967 333
rect -8889 287 -8843 333
rect -8765 287 -8719 333
rect -8641 287 -8595 333
rect -8517 287 -8471 333
rect -8393 287 -8347 333
rect -8269 287 -8223 333
rect -8145 287 -8099 333
rect -8021 287 -7975 333
rect -7897 287 -7851 333
rect -7773 287 -7727 333
rect -7649 287 -7603 333
rect -7525 287 -7479 333
rect -7401 287 -7355 333
rect -7277 287 -7231 333
rect -7153 287 -7107 333
rect -7029 287 -6983 333
rect -6905 287 -6859 333
rect -6781 287 -6735 333
rect -6657 287 -6611 333
rect -6533 287 -6487 333
rect -6409 287 -6363 333
rect -6285 287 -6239 333
rect -6161 287 -6115 333
rect -6037 287 -5991 333
rect -5913 287 -5867 333
rect -5789 287 -5743 333
rect -5665 287 -5619 333
rect -5541 287 -5495 333
rect -5417 287 -5371 333
rect -5293 287 -5247 333
rect -5169 287 -5123 333
rect -5045 287 -4999 333
rect -4921 287 -4875 333
rect -4797 287 -4751 333
rect -4673 287 -4627 333
rect -4549 287 -4503 333
rect -4425 287 -4379 333
rect -4301 287 -4255 333
rect -4177 287 -4131 333
rect -4053 287 -4007 333
rect -3929 287 -3883 333
rect -3805 287 -3759 333
rect -3681 287 -3635 333
rect -3557 287 -3511 333
rect -3433 287 -3387 333
rect -3309 287 -3263 333
rect -3185 287 -3139 333
rect -3061 287 -3015 333
rect -2937 287 -2891 333
rect -2813 287 -2767 333
rect -2689 287 -2643 333
rect -2565 287 -2519 333
rect -2441 287 -2395 333
rect -2317 287 -2271 333
rect -2193 287 -2147 333
rect -2069 287 -2023 333
rect -1945 287 -1899 333
rect -1821 287 -1775 333
rect -1697 287 -1651 333
rect -1573 287 -1527 333
rect -1449 287 -1403 333
rect -1325 287 -1279 333
rect -1201 287 -1155 333
rect -1077 287 -1031 333
rect -953 287 -907 333
rect -829 287 -783 333
rect -705 287 -659 333
rect -581 287 -535 333
rect -457 287 -411 333
rect -333 287 -287 333
rect -209 287 -163 333
rect -85 287 -39 333
rect 39 287 85 333
rect 163 287 209 333
rect 287 287 333 333
rect 411 287 457 333
rect 535 287 581 333
rect 659 287 705 333
rect 783 287 829 333
rect 907 287 953 333
rect 1031 287 1077 333
rect 1155 287 1201 333
rect 1279 287 1325 333
rect 1403 287 1449 333
rect 1527 287 1573 333
rect 1651 287 1697 333
rect 1775 287 1821 333
rect 1899 287 1945 333
rect 2023 287 2069 333
rect 2147 287 2193 333
rect 2271 287 2317 333
rect 2395 287 2441 333
rect 2519 287 2565 333
rect 2643 287 2689 333
rect 2767 287 2813 333
rect 2891 287 2937 333
rect 3015 287 3061 333
rect 3139 287 3185 333
rect 3263 287 3309 333
rect 3387 287 3433 333
rect 3511 287 3557 333
rect 3635 287 3681 333
rect 3759 287 3805 333
rect 3883 287 3929 333
rect 4007 287 4053 333
rect 4131 287 4177 333
rect 4255 287 4301 333
rect 4379 287 4425 333
rect 4503 287 4549 333
rect 4627 287 4673 333
rect 4751 287 4797 333
rect 4875 287 4921 333
rect 4999 287 5045 333
rect 5123 287 5169 333
rect 5247 287 5293 333
rect 5371 287 5417 333
rect 5495 287 5541 333
rect 5619 287 5665 333
rect 5743 287 5789 333
rect 5867 287 5913 333
rect 5991 287 6037 333
rect 6115 287 6161 333
rect 6239 287 6285 333
rect 6363 287 6409 333
rect 6487 287 6533 333
rect 6611 287 6657 333
rect 6735 287 6781 333
rect 6859 287 6905 333
rect 6983 287 7029 333
rect 7107 287 7153 333
rect 7231 287 7277 333
rect 7355 287 7401 333
rect 7479 287 7525 333
rect 7603 287 7649 333
rect 7727 287 7773 333
rect 7851 287 7897 333
rect 7975 287 8021 333
rect 8099 287 8145 333
rect 8223 287 8269 333
rect 8347 287 8393 333
rect 8471 287 8517 333
rect 8595 287 8641 333
rect 8719 287 8765 333
rect 8843 287 8889 333
rect 8967 287 9013 333
rect 9091 287 9137 333
rect 9215 287 9261 333
rect 9339 287 9385 333
rect 9463 287 9509 333
rect 9587 287 9633 333
rect 9711 287 9757 333
rect 9835 287 9881 333
rect 9959 287 10005 333
rect 10083 287 10129 333
rect 10207 287 10253 333
rect 10331 287 10377 333
rect 10455 287 10501 333
rect 10579 287 10625 333
rect 10703 287 10749 333
rect 10827 287 10873 333
rect 10951 287 10997 333
rect 11075 287 11121 333
rect 11199 287 11245 333
rect 11323 287 11369 333
rect 11447 287 11493 333
rect 11571 287 11617 333
rect 11695 287 11741 333
rect 11819 287 11865 333
rect 11943 287 11989 333
rect 12067 287 12113 333
rect 12191 287 12237 333
rect 12315 287 12361 333
rect 12439 287 12485 333
rect 12563 287 12609 333
rect 12687 287 12733 333
rect 12811 287 12857 333
rect 12935 287 12981 333
rect 13059 287 13105 333
rect 13183 287 13229 333
rect 13307 287 13353 333
rect 13431 287 13477 333
rect 13555 287 13601 333
rect 13679 287 13725 333
rect 13803 287 13849 333
rect 13927 287 13973 333
rect 14051 287 14097 333
rect 14175 287 14221 333
rect 14299 287 14345 333
rect 14423 287 14469 333
rect 14547 287 14593 333
rect 14671 287 14717 333
rect 14795 287 14841 333
rect 14919 287 14965 333
rect 15043 287 15089 333
rect 15167 287 15213 333
rect 15291 287 15337 333
rect 15415 287 15461 333
rect 15539 287 15585 333
rect 15663 287 15709 333
rect 15787 287 15833 333
rect 15911 287 15957 333
rect 16035 287 16081 333
rect 16159 287 16205 333
rect 16283 287 16329 333
rect 16407 287 16453 333
rect 16531 287 16577 333
rect 16655 287 16701 333
rect 16779 287 16825 333
rect 16903 287 16949 333
rect 17027 287 17073 333
rect 17151 287 17197 333
rect 17275 287 17321 333
rect -17321 163 -17275 209
rect -17197 163 -17151 209
rect -17073 163 -17027 209
rect -16949 163 -16903 209
rect -16825 163 -16779 209
rect -16701 163 -16655 209
rect -16577 163 -16531 209
rect -16453 163 -16407 209
rect -16329 163 -16283 209
rect -16205 163 -16159 209
rect -16081 163 -16035 209
rect -15957 163 -15911 209
rect -15833 163 -15787 209
rect -15709 163 -15663 209
rect -15585 163 -15539 209
rect -15461 163 -15415 209
rect -15337 163 -15291 209
rect -15213 163 -15167 209
rect -15089 163 -15043 209
rect -14965 163 -14919 209
rect -14841 163 -14795 209
rect -14717 163 -14671 209
rect -14593 163 -14547 209
rect -14469 163 -14423 209
rect -14345 163 -14299 209
rect -14221 163 -14175 209
rect -14097 163 -14051 209
rect -13973 163 -13927 209
rect -13849 163 -13803 209
rect -13725 163 -13679 209
rect -13601 163 -13555 209
rect -13477 163 -13431 209
rect -13353 163 -13307 209
rect -13229 163 -13183 209
rect -13105 163 -13059 209
rect -12981 163 -12935 209
rect -12857 163 -12811 209
rect -12733 163 -12687 209
rect -12609 163 -12563 209
rect -12485 163 -12439 209
rect -12361 163 -12315 209
rect -12237 163 -12191 209
rect -12113 163 -12067 209
rect -11989 163 -11943 209
rect -11865 163 -11819 209
rect -11741 163 -11695 209
rect -11617 163 -11571 209
rect -11493 163 -11447 209
rect -11369 163 -11323 209
rect -11245 163 -11199 209
rect -11121 163 -11075 209
rect -10997 163 -10951 209
rect -10873 163 -10827 209
rect -10749 163 -10703 209
rect -10625 163 -10579 209
rect -10501 163 -10455 209
rect -10377 163 -10331 209
rect -10253 163 -10207 209
rect -10129 163 -10083 209
rect -10005 163 -9959 209
rect -9881 163 -9835 209
rect -9757 163 -9711 209
rect -9633 163 -9587 209
rect -9509 163 -9463 209
rect -9385 163 -9339 209
rect -9261 163 -9215 209
rect -9137 163 -9091 209
rect -9013 163 -8967 209
rect -8889 163 -8843 209
rect -8765 163 -8719 209
rect -8641 163 -8595 209
rect -8517 163 -8471 209
rect -8393 163 -8347 209
rect -8269 163 -8223 209
rect -8145 163 -8099 209
rect -8021 163 -7975 209
rect -7897 163 -7851 209
rect -7773 163 -7727 209
rect -7649 163 -7603 209
rect -7525 163 -7479 209
rect -7401 163 -7355 209
rect -7277 163 -7231 209
rect -7153 163 -7107 209
rect -7029 163 -6983 209
rect -6905 163 -6859 209
rect -6781 163 -6735 209
rect -6657 163 -6611 209
rect -6533 163 -6487 209
rect -6409 163 -6363 209
rect -6285 163 -6239 209
rect -6161 163 -6115 209
rect -6037 163 -5991 209
rect -5913 163 -5867 209
rect -5789 163 -5743 209
rect -5665 163 -5619 209
rect -5541 163 -5495 209
rect -5417 163 -5371 209
rect -5293 163 -5247 209
rect -5169 163 -5123 209
rect -5045 163 -4999 209
rect -4921 163 -4875 209
rect -4797 163 -4751 209
rect -4673 163 -4627 209
rect -4549 163 -4503 209
rect -4425 163 -4379 209
rect -4301 163 -4255 209
rect -4177 163 -4131 209
rect -4053 163 -4007 209
rect -3929 163 -3883 209
rect -3805 163 -3759 209
rect -3681 163 -3635 209
rect -3557 163 -3511 209
rect -3433 163 -3387 209
rect -3309 163 -3263 209
rect -3185 163 -3139 209
rect -3061 163 -3015 209
rect -2937 163 -2891 209
rect -2813 163 -2767 209
rect -2689 163 -2643 209
rect -2565 163 -2519 209
rect -2441 163 -2395 209
rect -2317 163 -2271 209
rect -2193 163 -2147 209
rect -2069 163 -2023 209
rect -1945 163 -1899 209
rect -1821 163 -1775 209
rect -1697 163 -1651 209
rect -1573 163 -1527 209
rect -1449 163 -1403 209
rect -1325 163 -1279 209
rect -1201 163 -1155 209
rect -1077 163 -1031 209
rect -953 163 -907 209
rect -829 163 -783 209
rect -705 163 -659 209
rect -581 163 -535 209
rect -457 163 -411 209
rect -333 163 -287 209
rect -209 163 -163 209
rect -85 163 -39 209
rect 39 163 85 209
rect 163 163 209 209
rect 287 163 333 209
rect 411 163 457 209
rect 535 163 581 209
rect 659 163 705 209
rect 783 163 829 209
rect 907 163 953 209
rect 1031 163 1077 209
rect 1155 163 1201 209
rect 1279 163 1325 209
rect 1403 163 1449 209
rect 1527 163 1573 209
rect 1651 163 1697 209
rect 1775 163 1821 209
rect 1899 163 1945 209
rect 2023 163 2069 209
rect 2147 163 2193 209
rect 2271 163 2317 209
rect 2395 163 2441 209
rect 2519 163 2565 209
rect 2643 163 2689 209
rect 2767 163 2813 209
rect 2891 163 2937 209
rect 3015 163 3061 209
rect 3139 163 3185 209
rect 3263 163 3309 209
rect 3387 163 3433 209
rect 3511 163 3557 209
rect 3635 163 3681 209
rect 3759 163 3805 209
rect 3883 163 3929 209
rect 4007 163 4053 209
rect 4131 163 4177 209
rect 4255 163 4301 209
rect 4379 163 4425 209
rect 4503 163 4549 209
rect 4627 163 4673 209
rect 4751 163 4797 209
rect 4875 163 4921 209
rect 4999 163 5045 209
rect 5123 163 5169 209
rect 5247 163 5293 209
rect 5371 163 5417 209
rect 5495 163 5541 209
rect 5619 163 5665 209
rect 5743 163 5789 209
rect 5867 163 5913 209
rect 5991 163 6037 209
rect 6115 163 6161 209
rect 6239 163 6285 209
rect 6363 163 6409 209
rect 6487 163 6533 209
rect 6611 163 6657 209
rect 6735 163 6781 209
rect 6859 163 6905 209
rect 6983 163 7029 209
rect 7107 163 7153 209
rect 7231 163 7277 209
rect 7355 163 7401 209
rect 7479 163 7525 209
rect 7603 163 7649 209
rect 7727 163 7773 209
rect 7851 163 7897 209
rect 7975 163 8021 209
rect 8099 163 8145 209
rect 8223 163 8269 209
rect 8347 163 8393 209
rect 8471 163 8517 209
rect 8595 163 8641 209
rect 8719 163 8765 209
rect 8843 163 8889 209
rect 8967 163 9013 209
rect 9091 163 9137 209
rect 9215 163 9261 209
rect 9339 163 9385 209
rect 9463 163 9509 209
rect 9587 163 9633 209
rect 9711 163 9757 209
rect 9835 163 9881 209
rect 9959 163 10005 209
rect 10083 163 10129 209
rect 10207 163 10253 209
rect 10331 163 10377 209
rect 10455 163 10501 209
rect 10579 163 10625 209
rect 10703 163 10749 209
rect 10827 163 10873 209
rect 10951 163 10997 209
rect 11075 163 11121 209
rect 11199 163 11245 209
rect 11323 163 11369 209
rect 11447 163 11493 209
rect 11571 163 11617 209
rect 11695 163 11741 209
rect 11819 163 11865 209
rect 11943 163 11989 209
rect 12067 163 12113 209
rect 12191 163 12237 209
rect 12315 163 12361 209
rect 12439 163 12485 209
rect 12563 163 12609 209
rect 12687 163 12733 209
rect 12811 163 12857 209
rect 12935 163 12981 209
rect 13059 163 13105 209
rect 13183 163 13229 209
rect 13307 163 13353 209
rect 13431 163 13477 209
rect 13555 163 13601 209
rect 13679 163 13725 209
rect 13803 163 13849 209
rect 13927 163 13973 209
rect 14051 163 14097 209
rect 14175 163 14221 209
rect 14299 163 14345 209
rect 14423 163 14469 209
rect 14547 163 14593 209
rect 14671 163 14717 209
rect 14795 163 14841 209
rect 14919 163 14965 209
rect 15043 163 15089 209
rect 15167 163 15213 209
rect 15291 163 15337 209
rect 15415 163 15461 209
rect 15539 163 15585 209
rect 15663 163 15709 209
rect 15787 163 15833 209
rect 15911 163 15957 209
rect 16035 163 16081 209
rect 16159 163 16205 209
rect 16283 163 16329 209
rect 16407 163 16453 209
rect 16531 163 16577 209
rect 16655 163 16701 209
rect 16779 163 16825 209
rect 16903 163 16949 209
rect 17027 163 17073 209
rect 17151 163 17197 209
rect 17275 163 17321 209
rect -17321 39 -17275 85
rect -17197 39 -17151 85
rect -17073 39 -17027 85
rect -16949 39 -16903 85
rect -16825 39 -16779 85
rect -16701 39 -16655 85
rect -16577 39 -16531 85
rect -16453 39 -16407 85
rect -16329 39 -16283 85
rect -16205 39 -16159 85
rect -16081 39 -16035 85
rect -15957 39 -15911 85
rect -15833 39 -15787 85
rect -15709 39 -15663 85
rect -15585 39 -15539 85
rect -15461 39 -15415 85
rect -15337 39 -15291 85
rect -15213 39 -15167 85
rect -15089 39 -15043 85
rect -14965 39 -14919 85
rect -14841 39 -14795 85
rect -14717 39 -14671 85
rect -14593 39 -14547 85
rect -14469 39 -14423 85
rect -14345 39 -14299 85
rect -14221 39 -14175 85
rect -14097 39 -14051 85
rect -13973 39 -13927 85
rect -13849 39 -13803 85
rect -13725 39 -13679 85
rect -13601 39 -13555 85
rect -13477 39 -13431 85
rect -13353 39 -13307 85
rect -13229 39 -13183 85
rect -13105 39 -13059 85
rect -12981 39 -12935 85
rect -12857 39 -12811 85
rect -12733 39 -12687 85
rect -12609 39 -12563 85
rect -12485 39 -12439 85
rect -12361 39 -12315 85
rect -12237 39 -12191 85
rect -12113 39 -12067 85
rect -11989 39 -11943 85
rect -11865 39 -11819 85
rect -11741 39 -11695 85
rect -11617 39 -11571 85
rect -11493 39 -11447 85
rect -11369 39 -11323 85
rect -11245 39 -11199 85
rect -11121 39 -11075 85
rect -10997 39 -10951 85
rect -10873 39 -10827 85
rect -10749 39 -10703 85
rect -10625 39 -10579 85
rect -10501 39 -10455 85
rect -10377 39 -10331 85
rect -10253 39 -10207 85
rect -10129 39 -10083 85
rect -10005 39 -9959 85
rect -9881 39 -9835 85
rect -9757 39 -9711 85
rect -9633 39 -9587 85
rect -9509 39 -9463 85
rect -9385 39 -9339 85
rect -9261 39 -9215 85
rect -9137 39 -9091 85
rect -9013 39 -8967 85
rect -8889 39 -8843 85
rect -8765 39 -8719 85
rect -8641 39 -8595 85
rect -8517 39 -8471 85
rect -8393 39 -8347 85
rect -8269 39 -8223 85
rect -8145 39 -8099 85
rect -8021 39 -7975 85
rect -7897 39 -7851 85
rect -7773 39 -7727 85
rect -7649 39 -7603 85
rect -7525 39 -7479 85
rect -7401 39 -7355 85
rect -7277 39 -7231 85
rect -7153 39 -7107 85
rect -7029 39 -6983 85
rect -6905 39 -6859 85
rect -6781 39 -6735 85
rect -6657 39 -6611 85
rect -6533 39 -6487 85
rect -6409 39 -6363 85
rect -6285 39 -6239 85
rect -6161 39 -6115 85
rect -6037 39 -5991 85
rect -5913 39 -5867 85
rect -5789 39 -5743 85
rect -5665 39 -5619 85
rect -5541 39 -5495 85
rect -5417 39 -5371 85
rect -5293 39 -5247 85
rect -5169 39 -5123 85
rect -5045 39 -4999 85
rect -4921 39 -4875 85
rect -4797 39 -4751 85
rect -4673 39 -4627 85
rect -4549 39 -4503 85
rect -4425 39 -4379 85
rect -4301 39 -4255 85
rect -4177 39 -4131 85
rect -4053 39 -4007 85
rect -3929 39 -3883 85
rect -3805 39 -3759 85
rect -3681 39 -3635 85
rect -3557 39 -3511 85
rect -3433 39 -3387 85
rect -3309 39 -3263 85
rect -3185 39 -3139 85
rect -3061 39 -3015 85
rect -2937 39 -2891 85
rect -2813 39 -2767 85
rect -2689 39 -2643 85
rect -2565 39 -2519 85
rect -2441 39 -2395 85
rect -2317 39 -2271 85
rect -2193 39 -2147 85
rect -2069 39 -2023 85
rect -1945 39 -1899 85
rect -1821 39 -1775 85
rect -1697 39 -1651 85
rect -1573 39 -1527 85
rect -1449 39 -1403 85
rect -1325 39 -1279 85
rect -1201 39 -1155 85
rect -1077 39 -1031 85
rect -953 39 -907 85
rect -829 39 -783 85
rect -705 39 -659 85
rect -581 39 -535 85
rect -457 39 -411 85
rect -333 39 -287 85
rect -209 39 -163 85
rect -85 39 -39 85
rect 39 39 85 85
rect 163 39 209 85
rect 287 39 333 85
rect 411 39 457 85
rect 535 39 581 85
rect 659 39 705 85
rect 783 39 829 85
rect 907 39 953 85
rect 1031 39 1077 85
rect 1155 39 1201 85
rect 1279 39 1325 85
rect 1403 39 1449 85
rect 1527 39 1573 85
rect 1651 39 1697 85
rect 1775 39 1821 85
rect 1899 39 1945 85
rect 2023 39 2069 85
rect 2147 39 2193 85
rect 2271 39 2317 85
rect 2395 39 2441 85
rect 2519 39 2565 85
rect 2643 39 2689 85
rect 2767 39 2813 85
rect 2891 39 2937 85
rect 3015 39 3061 85
rect 3139 39 3185 85
rect 3263 39 3309 85
rect 3387 39 3433 85
rect 3511 39 3557 85
rect 3635 39 3681 85
rect 3759 39 3805 85
rect 3883 39 3929 85
rect 4007 39 4053 85
rect 4131 39 4177 85
rect 4255 39 4301 85
rect 4379 39 4425 85
rect 4503 39 4549 85
rect 4627 39 4673 85
rect 4751 39 4797 85
rect 4875 39 4921 85
rect 4999 39 5045 85
rect 5123 39 5169 85
rect 5247 39 5293 85
rect 5371 39 5417 85
rect 5495 39 5541 85
rect 5619 39 5665 85
rect 5743 39 5789 85
rect 5867 39 5913 85
rect 5991 39 6037 85
rect 6115 39 6161 85
rect 6239 39 6285 85
rect 6363 39 6409 85
rect 6487 39 6533 85
rect 6611 39 6657 85
rect 6735 39 6781 85
rect 6859 39 6905 85
rect 6983 39 7029 85
rect 7107 39 7153 85
rect 7231 39 7277 85
rect 7355 39 7401 85
rect 7479 39 7525 85
rect 7603 39 7649 85
rect 7727 39 7773 85
rect 7851 39 7897 85
rect 7975 39 8021 85
rect 8099 39 8145 85
rect 8223 39 8269 85
rect 8347 39 8393 85
rect 8471 39 8517 85
rect 8595 39 8641 85
rect 8719 39 8765 85
rect 8843 39 8889 85
rect 8967 39 9013 85
rect 9091 39 9137 85
rect 9215 39 9261 85
rect 9339 39 9385 85
rect 9463 39 9509 85
rect 9587 39 9633 85
rect 9711 39 9757 85
rect 9835 39 9881 85
rect 9959 39 10005 85
rect 10083 39 10129 85
rect 10207 39 10253 85
rect 10331 39 10377 85
rect 10455 39 10501 85
rect 10579 39 10625 85
rect 10703 39 10749 85
rect 10827 39 10873 85
rect 10951 39 10997 85
rect 11075 39 11121 85
rect 11199 39 11245 85
rect 11323 39 11369 85
rect 11447 39 11493 85
rect 11571 39 11617 85
rect 11695 39 11741 85
rect 11819 39 11865 85
rect 11943 39 11989 85
rect 12067 39 12113 85
rect 12191 39 12237 85
rect 12315 39 12361 85
rect 12439 39 12485 85
rect 12563 39 12609 85
rect 12687 39 12733 85
rect 12811 39 12857 85
rect 12935 39 12981 85
rect 13059 39 13105 85
rect 13183 39 13229 85
rect 13307 39 13353 85
rect 13431 39 13477 85
rect 13555 39 13601 85
rect 13679 39 13725 85
rect 13803 39 13849 85
rect 13927 39 13973 85
rect 14051 39 14097 85
rect 14175 39 14221 85
rect 14299 39 14345 85
rect 14423 39 14469 85
rect 14547 39 14593 85
rect 14671 39 14717 85
rect 14795 39 14841 85
rect 14919 39 14965 85
rect 15043 39 15089 85
rect 15167 39 15213 85
rect 15291 39 15337 85
rect 15415 39 15461 85
rect 15539 39 15585 85
rect 15663 39 15709 85
rect 15787 39 15833 85
rect 15911 39 15957 85
rect 16035 39 16081 85
rect 16159 39 16205 85
rect 16283 39 16329 85
rect 16407 39 16453 85
rect 16531 39 16577 85
rect 16655 39 16701 85
rect 16779 39 16825 85
rect 16903 39 16949 85
rect 17027 39 17073 85
rect 17151 39 17197 85
rect 17275 39 17321 85
rect -17321 -85 -17275 -39
rect -17197 -85 -17151 -39
rect -17073 -85 -17027 -39
rect -16949 -85 -16903 -39
rect -16825 -85 -16779 -39
rect -16701 -85 -16655 -39
rect -16577 -85 -16531 -39
rect -16453 -85 -16407 -39
rect -16329 -85 -16283 -39
rect -16205 -85 -16159 -39
rect -16081 -85 -16035 -39
rect -15957 -85 -15911 -39
rect -15833 -85 -15787 -39
rect -15709 -85 -15663 -39
rect -15585 -85 -15539 -39
rect -15461 -85 -15415 -39
rect -15337 -85 -15291 -39
rect -15213 -85 -15167 -39
rect -15089 -85 -15043 -39
rect -14965 -85 -14919 -39
rect -14841 -85 -14795 -39
rect -14717 -85 -14671 -39
rect -14593 -85 -14547 -39
rect -14469 -85 -14423 -39
rect -14345 -85 -14299 -39
rect -14221 -85 -14175 -39
rect -14097 -85 -14051 -39
rect -13973 -85 -13927 -39
rect -13849 -85 -13803 -39
rect -13725 -85 -13679 -39
rect -13601 -85 -13555 -39
rect -13477 -85 -13431 -39
rect -13353 -85 -13307 -39
rect -13229 -85 -13183 -39
rect -13105 -85 -13059 -39
rect -12981 -85 -12935 -39
rect -12857 -85 -12811 -39
rect -12733 -85 -12687 -39
rect -12609 -85 -12563 -39
rect -12485 -85 -12439 -39
rect -12361 -85 -12315 -39
rect -12237 -85 -12191 -39
rect -12113 -85 -12067 -39
rect -11989 -85 -11943 -39
rect -11865 -85 -11819 -39
rect -11741 -85 -11695 -39
rect -11617 -85 -11571 -39
rect -11493 -85 -11447 -39
rect -11369 -85 -11323 -39
rect -11245 -85 -11199 -39
rect -11121 -85 -11075 -39
rect -10997 -85 -10951 -39
rect -10873 -85 -10827 -39
rect -10749 -85 -10703 -39
rect -10625 -85 -10579 -39
rect -10501 -85 -10455 -39
rect -10377 -85 -10331 -39
rect -10253 -85 -10207 -39
rect -10129 -85 -10083 -39
rect -10005 -85 -9959 -39
rect -9881 -85 -9835 -39
rect -9757 -85 -9711 -39
rect -9633 -85 -9587 -39
rect -9509 -85 -9463 -39
rect -9385 -85 -9339 -39
rect -9261 -85 -9215 -39
rect -9137 -85 -9091 -39
rect -9013 -85 -8967 -39
rect -8889 -85 -8843 -39
rect -8765 -85 -8719 -39
rect -8641 -85 -8595 -39
rect -8517 -85 -8471 -39
rect -8393 -85 -8347 -39
rect -8269 -85 -8223 -39
rect -8145 -85 -8099 -39
rect -8021 -85 -7975 -39
rect -7897 -85 -7851 -39
rect -7773 -85 -7727 -39
rect -7649 -85 -7603 -39
rect -7525 -85 -7479 -39
rect -7401 -85 -7355 -39
rect -7277 -85 -7231 -39
rect -7153 -85 -7107 -39
rect -7029 -85 -6983 -39
rect -6905 -85 -6859 -39
rect -6781 -85 -6735 -39
rect -6657 -85 -6611 -39
rect -6533 -85 -6487 -39
rect -6409 -85 -6363 -39
rect -6285 -85 -6239 -39
rect -6161 -85 -6115 -39
rect -6037 -85 -5991 -39
rect -5913 -85 -5867 -39
rect -5789 -85 -5743 -39
rect -5665 -85 -5619 -39
rect -5541 -85 -5495 -39
rect -5417 -85 -5371 -39
rect -5293 -85 -5247 -39
rect -5169 -85 -5123 -39
rect -5045 -85 -4999 -39
rect -4921 -85 -4875 -39
rect -4797 -85 -4751 -39
rect -4673 -85 -4627 -39
rect -4549 -85 -4503 -39
rect -4425 -85 -4379 -39
rect -4301 -85 -4255 -39
rect -4177 -85 -4131 -39
rect -4053 -85 -4007 -39
rect -3929 -85 -3883 -39
rect -3805 -85 -3759 -39
rect -3681 -85 -3635 -39
rect -3557 -85 -3511 -39
rect -3433 -85 -3387 -39
rect -3309 -85 -3263 -39
rect -3185 -85 -3139 -39
rect -3061 -85 -3015 -39
rect -2937 -85 -2891 -39
rect -2813 -85 -2767 -39
rect -2689 -85 -2643 -39
rect -2565 -85 -2519 -39
rect -2441 -85 -2395 -39
rect -2317 -85 -2271 -39
rect -2193 -85 -2147 -39
rect -2069 -85 -2023 -39
rect -1945 -85 -1899 -39
rect -1821 -85 -1775 -39
rect -1697 -85 -1651 -39
rect -1573 -85 -1527 -39
rect -1449 -85 -1403 -39
rect -1325 -85 -1279 -39
rect -1201 -85 -1155 -39
rect -1077 -85 -1031 -39
rect -953 -85 -907 -39
rect -829 -85 -783 -39
rect -705 -85 -659 -39
rect -581 -85 -535 -39
rect -457 -85 -411 -39
rect -333 -85 -287 -39
rect -209 -85 -163 -39
rect -85 -85 -39 -39
rect 39 -85 85 -39
rect 163 -85 209 -39
rect 287 -85 333 -39
rect 411 -85 457 -39
rect 535 -85 581 -39
rect 659 -85 705 -39
rect 783 -85 829 -39
rect 907 -85 953 -39
rect 1031 -85 1077 -39
rect 1155 -85 1201 -39
rect 1279 -85 1325 -39
rect 1403 -85 1449 -39
rect 1527 -85 1573 -39
rect 1651 -85 1697 -39
rect 1775 -85 1821 -39
rect 1899 -85 1945 -39
rect 2023 -85 2069 -39
rect 2147 -85 2193 -39
rect 2271 -85 2317 -39
rect 2395 -85 2441 -39
rect 2519 -85 2565 -39
rect 2643 -85 2689 -39
rect 2767 -85 2813 -39
rect 2891 -85 2937 -39
rect 3015 -85 3061 -39
rect 3139 -85 3185 -39
rect 3263 -85 3309 -39
rect 3387 -85 3433 -39
rect 3511 -85 3557 -39
rect 3635 -85 3681 -39
rect 3759 -85 3805 -39
rect 3883 -85 3929 -39
rect 4007 -85 4053 -39
rect 4131 -85 4177 -39
rect 4255 -85 4301 -39
rect 4379 -85 4425 -39
rect 4503 -85 4549 -39
rect 4627 -85 4673 -39
rect 4751 -85 4797 -39
rect 4875 -85 4921 -39
rect 4999 -85 5045 -39
rect 5123 -85 5169 -39
rect 5247 -85 5293 -39
rect 5371 -85 5417 -39
rect 5495 -85 5541 -39
rect 5619 -85 5665 -39
rect 5743 -85 5789 -39
rect 5867 -85 5913 -39
rect 5991 -85 6037 -39
rect 6115 -85 6161 -39
rect 6239 -85 6285 -39
rect 6363 -85 6409 -39
rect 6487 -85 6533 -39
rect 6611 -85 6657 -39
rect 6735 -85 6781 -39
rect 6859 -85 6905 -39
rect 6983 -85 7029 -39
rect 7107 -85 7153 -39
rect 7231 -85 7277 -39
rect 7355 -85 7401 -39
rect 7479 -85 7525 -39
rect 7603 -85 7649 -39
rect 7727 -85 7773 -39
rect 7851 -85 7897 -39
rect 7975 -85 8021 -39
rect 8099 -85 8145 -39
rect 8223 -85 8269 -39
rect 8347 -85 8393 -39
rect 8471 -85 8517 -39
rect 8595 -85 8641 -39
rect 8719 -85 8765 -39
rect 8843 -85 8889 -39
rect 8967 -85 9013 -39
rect 9091 -85 9137 -39
rect 9215 -85 9261 -39
rect 9339 -85 9385 -39
rect 9463 -85 9509 -39
rect 9587 -85 9633 -39
rect 9711 -85 9757 -39
rect 9835 -85 9881 -39
rect 9959 -85 10005 -39
rect 10083 -85 10129 -39
rect 10207 -85 10253 -39
rect 10331 -85 10377 -39
rect 10455 -85 10501 -39
rect 10579 -85 10625 -39
rect 10703 -85 10749 -39
rect 10827 -85 10873 -39
rect 10951 -85 10997 -39
rect 11075 -85 11121 -39
rect 11199 -85 11245 -39
rect 11323 -85 11369 -39
rect 11447 -85 11493 -39
rect 11571 -85 11617 -39
rect 11695 -85 11741 -39
rect 11819 -85 11865 -39
rect 11943 -85 11989 -39
rect 12067 -85 12113 -39
rect 12191 -85 12237 -39
rect 12315 -85 12361 -39
rect 12439 -85 12485 -39
rect 12563 -85 12609 -39
rect 12687 -85 12733 -39
rect 12811 -85 12857 -39
rect 12935 -85 12981 -39
rect 13059 -85 13105 -39
rect 13183 -85 13229 -39
rect 13307 -85 13353 -39
rect 13431 -85 13477 -39
rect 13555 -85 13601 -39
rect 13679 -85 13725 -39
rect 13803 -85 13849 -39
rect 13927 -85 13973 -39
rect 14051 -85 14097 -39
rect 14175 -85 14221 -39
rect 14299 -85 14345 -39
rect 14423 -85 14469 -39
rect 14547 -85 14593 -39
rect 14671 -85 14717 -39
rect 14795 -85 14841 -39
rect 14919 -85 14965 -39
rect 15043 -85 15089 -39
rect 15167 -85 15213 -39
rect 15291 -85 15337 -39
rect 15415 -85 15461 -39
rect 15539 -85 15585 -39
rect 15663 -85 15709 -39
rect 15787 -85 15833 -39
rect 15911 -85 15957 -39
rect 16035 -85 16081 -39
rect 16159 -85 16205 -39
rect 16283 -85 16329 -39
rect 16407 -85 16453 -39
rect 16531 -85 16577 -39
rect 16655 -85 16701 -39
rect 16779 -85 16825 -39
rect 16903 -85 16949 -39
rect 17027 -85 17073 -39
rect 17151 -85 17197 -39
rect 17275 -85 17321 -39
rect -17321 -209 -17275 -163
rect -17197 -209 -17151 -163
rect -17073 -209 -17027 -163
rect -16949 -209 -16903 -163
rect -16825 -209 -16779 -163
rect -16701 -209 -16655 -163
rect -16577 -209 -16531 -163
rect -16453 -209 -16407 -163
rect -16329 -209 -16283 -163
rect -16205 -209 -16159 -163
rect -16081 -209 -16035 -163
rect -15957 -209 -15911 -163
rect -15833 -209 -15787 -163
rect -15709 -209 -15663 -163
rect -15585 -209 -15539 -163
rect -15461 -209 -15415 -163
rect -15337 -209 -15291 -163
rect -15213 -209 -15167 -163
rect -15089 -209 -15043 -163
rect -14965 -209 -14919 -163
rect -14841 -209 -14795 -163
rect -14717 -209 -14671 -163
rect -14593 -209 -14547 -163
rect -14469 -209 -14423 -163
rect -14345 -209 -14299 -163
rect -14221 -209 -14175 -163
rect -14097 -209 -14051 -163
rect -13973 -209 -13927 -163
rect -13849 -209 -13803 -163
rect -13725 -209 -13679 -163
rect -13601 -209 -13555 -163
rect -13477 -209 -13431 -163
rect -13353 -209 -13307 -163
rect -13229 -209 -13183 -163
rect -13105 -209 -13059 -163
rect -12981 -209 -12935 -163
rect -12857 -209 -12811 -163
rect -12733 -209 -12687 -163
rect -12609 -209 -12563 -163
rect -12485 -209 -12439 -163
rect -12361 -209 -12315 -163
rect -12237 -209 -12191 -163
rect -12113 -209 -12067 -163
rect -11989 -209 -11943 -163
rect -11865 -209 -11819 -163
rect -11741 -209 -11695 -163
rect -11617 -209 -11571 -163
rect -11493 -209 -11447 -163
rect -11369 -209 -11323 -163
rect -11245 -209 -11199 -163
rect -11121 -209 -11075 -163
rect -10997 -209 -10951 -163
rect -10873 -209 -10827 -163
rect -10749 -209 -10703 -163
rect -10625 -209 -10579 -163
rect -10501 -209 -10455 -163
rect -10377 -209 -10331 -163
rect -10253 -209 -10207 -163
rect -10129 -209 -10083 -163
rect -10005 -209 -9959 -163
rect -9881 -209 -9835 -163
rect -9757 -209 -9711 -163
rect -9633 -209 -9587 -163
rect -9509 -209 -9463 -163
rect -9385 -209 -9339 -163
rect -9261 -209 -9215 -163
rect -9137 -209 -9091 -163
rect -9013 -209 -8967 -163
rect -8889 -209 -8843 -163
rect -8765 -209 -8719 -163
rect -8641 -209 -8595 -163
rect -8517 -209 -8471 -163
rect -8393 -209 -8347 -163
rect -8269 -209 -8223 -163
rect -8145 -209 -8099 -163
rect -8021 -209 -7975 -163
rect -7897 -209 -7851 -163
rect -7773 -209 -7727 -163
rect -7649 -209 -7603 -163
rect -7525 -209 -7479 -163
rect -7401 -209 -7355 -163
rect -7277 -209 -7231 -163
rect -7153 -209 -7107 -163
rect -7029 -209 -6983 -163
rect -6905 -209 -6859 -163
rect -6781 -209 -6735 -163
rect -6657 -209 -6611 -163
rect -6533 -209 -6487 -163
rect -6409 -209 -6363 -163
rect -6285 -209 -6239 -163
rect -6161 -209 -6115 -163
rect -6037 -209 -5991 -163
rect -5913 -209 -5867 -163
rect -5789 -209 -5743 -163
rect -5665 -209 -5619 -163
rect -5541 -209 -5495 -163
rect -5417 -209 -5371 -163
rect -5293 -209 -5247 -163
rect -5169 -209 -5123 -163
rect -5045 -209 -4999 -163
rect -4921 -209 -4875 -163
rect -4797 -209 -4751 -163
rect -4673 -209 -4627 -163
rect -4549 -209 -4503 -163
rect -4425 -209 -4379 -163
rect -4301 -209 -4255 -163
rect -4177 -209 -4131 -163
rect -4053 -209 -4007 -163
rect -3929 -209 -3883 -163
rect -3805 -209 -3759 -163
rect -3681 -209 -3635 -163
rect -3557 -209 -3511 -163
rect -3433 -209 -3387 -163
rect -3309 -209 -3263 -163
rect -3185 -209 -3139 -163
rect -3061 -209 -3015 -163
rect -2937 -209 -2891 -163
rect -2813 -209 -2767 -163
rect -2689 -209 -2643 -163
rect -2565 -209 -2519 -163
rect -2441 -209 -2395 -163
rect -2317 -209 -2271 -163
rect -2193 -209 -2147 -163
rect -2069 -209 -2023 -163
rect -1945 -209 -1899 -163
rect -1821 -209 -1775 -163
rect -1697 -209 -1651 -163
rect -1573 -209 -1527 -163
rect -1449 -209 -1403 -163
rect -1325 -209 -1279 -163
rect -1201 -209 -1155 -163
rect -1077 -209 -1031 -163
rect -953 -209 -907 -163
rect -829 -209 -783 -163
rect -705 -209 -659 -163
rect -581 -209 -535 -163
rect -457 -209 -411 -163
rect -333 -209 -287 -163
rect -209 -209 -163 -163
rect -85 -209 -39 -163
rect 39 -209 85 -163
rect 163 -209 209 -163
rect 287 -209 333 -163
rect 411 -209 457 -163
rect 535 -209 581 -163
rect 659 -209 705 -163
rect 783 -209 829 -163
rect 907 -209 953 -163
rect 1031 -209 1077 -163
rect 1155 -209 1201 -163
rect 1279 -209 1325 -163
rect 1403 -209 1449 -163
rect 1527 -209 1573 -163
rect 1651 -209 1697 -163
rect 1775 -209 1821 -163
rect 1899 -209 1945 -163
rect 2023 -209 2069 -163
rect 2147 -209 2193 -163
rect 2271 -209 2317 -163
rect 2395 -209 2441 -163
rect 2519 -209 2565 -163
rect 2643 -209 2689 -163
rect 2767 -209 2813 -163
rect 2891 -209 2937 -163
rect 3015 -209 3061 -163
rect 3139 -209 3185 -163
rect 3263 -209 3309 -163
rect 3387 -209 3433 -163
rect 3511 -209 3557 -163
rect 3635 -209 3681 -163
rect 3759 -209 3805 -163
rect 3883 -209 3929 -163
rect 4007 -209 4053 -163
rect 4131 -209 4177 -163
rect 4255 -209 4301 -163
rect 4379 -209 4425 -163
rect 4503 -209 4549 -163
rect 4627 -209 4673 -163
rect 4751 -209 4797 -163
rect 4875 -209 4921 -163
rect 4999 -209 5045 -163
rect 5123 -209 5169 -163
rect 5247 -209 5293 -163
rect 5371 -209 5417 -163
rect 5495 -209 5541 -163
rect 5619 -209 5665 -163
rect 5743 -209 5789 -163
rect 5867 -209 5913 -163
rect 5991 -209 6037 -163
rect 6115 -209 6161 -163
rect 6239 -209 6285 -163
rect 6363 -209 6409 -163
rect 6487 -209 6533 -163
rect 6611 -209 6657 -163
rect 6735 -209 6781 -163
rect 6859 -209 6905 -163
rect 6983 -209 7029 -163
rect 7107 -209 7153 -163
rect 7231 -209 7277 -163
rect 7355 -209 7401 -163
rect 7479 -209 7525 -163
rect 7603 -209 7649 -163
rect 7727 -209 7773 -163
rect 7851 -209 7897 -163
rect 7975 -209 8021 -163
rect 8099 -209 8145 -163
rect 8223 -209 8269 -163
rect 8347 -209 8393 -163
rect 8471 -209 8517 -163
rect 8595 -209 8641 -163
rect 8719 -209 8765 -163
rect 8843 -209 8889 -163
rect 8967 -209 9013 -163
rect 9091 -209 9137 -163
rect 9215 -209 9261 -163
rect 9339 -209 9385 -163
rect 9463 -209 9509 -163
rect 9587 -209 9633 -163
rect 9711 -209 9757 -163
rect 9835 -209 9881 -163
rect 9959 -209 10005 -163
rect 10083 -209 10129 -163
rect 10207 -209 10253 -163
rect 10331 -209 10377 -163
rect 10455 -209 10501 -163
rect 10579 -209 10625 -163
rect 10703 -209 10749 -163
rect 10827 -209 10873 -163
rect 10951 -209 10997 -163
rect 11075 -209 11121 -163
rect 11199 -209 11245 -163
rect 11323 -209 11369 -163
rect 11447 -209 11493 -163
rect 11571 -209 11617 -163
rect 11695 -209 11741 -163
rect 11819 -209 11865 -163
rect 11943 -209 11989 -163
rect 12067 -209 12113 -163
rect 12191 -209 12237 -163
rect 12315 -209 12361 -163
rect 12439 -209 12485 -163
rect 12563 -209 12609 -163
rect 12687 -209 12733 -163
rect 12811 -209 12857 -163
rect 12935 -209 12981 -163
rect 13059 -209 13105 -163
rect 13183 -209 13229 -163
rect 13307 -209 13353 -163
rect 13431 -209 13477 -163
rect 13555 -209 13601 -163
rect 13679 -209 13725 -163
rect 13803 -209 13849 -163
rect 13927 -209 13973 -163
rect 14051 -209 14097 -163
rect 14175 -209 14221 -163
rect 14299 -209 14345 -163
rect 14423 -209 14469 -163
rect 14547 -209 14593 -163
rect 14671 -209 14717 -163
rect 14795 -209 14841 -163
rect 14919 -209 14965 -163
rect 15043 -209 15089 -163
rect 15167 -209 15213 -163
rect 15291 -209 15337 -163
rect 15415 -209 15461 -163
rect 15539 -209 15585 -163
rect 15663 -209 15709 -163
rect 15787 -209 15833 -163
rect 15911 -209 15957 -163
rect 16035 -209 16081 -163
rect 16159 -209 16205 -163
rect 16283 -209 16329 -163
rect 16407 -209 16453 -163
rect 16531 -209 16577 -163
rect 16655 -209 16701 -163
rect 16779 -209 16825 -163
rect 16903 -209 16949 -163
rect 17027 -209 17073 -163
rect 17151 -209 17197 -163
rect 17275 -209 17321 -163
rect -17321 -333 -17275 -287
rect -17197 -333 -17151 -287
rect -17073 -333 -17027 -287
rect -16949 -333 -16903 -287
rect -16825 -333 -16779 -287
rect -16701 -333 -16655 -287
rect -16577 -333 -16531 -287
rect -16453 -333 -16407 -287
rect -16329 -333 -16283 -287
rect -16205 -333 -16159 -287
rect -16081 -333 -16035 -287
rect -15957 -333 -15911 -287
rect -15833 -333 -15787 -287
rect -15709 -333 -15663 -287
rect -15585 -333 -15539 -287
rect -15461 -333 -15415 -287
rect -15337 -333 -15291 -287
rect -15213 -333 -15167 -287
rect -15089 -333 -15043 -287
rect -14965 -333 -14919 -287
rect -14841 -333 -14795 -287
rect -14717 -333 -14671 -287
rect -14593 -333 -14547 -287
rect -14469 -333 -14423 -287
rect -14345 -333 -14299 -287
rect -14221 -333 -14175 -287
rect -14097 -333 -14051 -287
rect -13973 -333 -13927 -287
rect -13849 -333 -13803 -287
rect -13725 -333 -13679 -287
rect -13601 -333 -13555 -287
rect -13477 -333 -13431 -287
rect -13353 -333 -13307 -287
rect -13229 -333 -13183 -287
rect -13105 -333 -13059 -287
rect -12981 -333 -12935 -287
rect -12857 -333 -12811 -287
rect -12733 -333 -12687 -287
rect -12609 -333 -12563 -287
rect -12485 -333 -12439 -287
rect -12361 -333 -12315 -287
rect -12237 -333 -12191 -287
rect -12113 -333 -12067 -287
rect -11989 -333 -11943 -287
rect -11865 -333 -11819 -287
rect -11741 -333 -11695 -287
rect -11617 -333 -11571 -287
rect -11493 -333 -11447 -287
rect -11369 -333 -11323 -287
rect -11245 -333 -11199 -287
rect -11121 -333 -11075 -287
rect -10997 -333 -10951 -287
rect -10873 -333 -10827 -287
rect -10749 -333 -10703 -287
rect -10625 -333 -10579 -287
rect -10501 -333 -10455 -287
rect -10377 -333 -10331 -287
rect -10253 -333 -10207 -287
rect -10129 -333 -10083 -287
rect -10005 -333 -9959 -287
rect -9881 -333 -9835 -287
rect -9757 -333 -9711 -287
rect -9633 -333 -9587 -287
rect -9509 -333 -9463 -287
rect -9385 -333 -9339 -287
rect -9261 -333 -9215 -287
rect -9137 -333 -9091 -287
rect -9013 -333 -8967 -287
rect -8889 -333 -8843 -287
rect -8765 -333 -8719 -287
rect -8641 -333 -8595 -287
rect -8517 -333 -8471 -287
rect -8393 -333 -8347 -287
rect -8269 -333 -8223 -287
rect -8145 -333 -8099 -287
rect -8021 -333 -7975 -287
rect -7897 -333 -7851 -287
rect -7773 -333 -7727 -287
rect -7649 -333 -7603 -287
rect -7525 -333 -7479 -287
rect -7401 -333 -7355 -287
rect -7277 -333 -7231 -287
rect -7153 -333 -7107 -287
rect -7029 -333 -6983 -287
rect -6905 -333 -6859 -287
rect -6781 -333 -6735 -287
rect -6657 -333 -6611 -287
rect -6533 -333 -6487 -287
rect -6409 -333 -6363 -287
rect -6285 -333 -6239 -287
rect -6161 -333 -6115 -287
rect -6037 -333 -5991 -287
rect -5913 -333 -5867 -287
rect -5789 -333 -5743 -287
rect -5665 -333 -5619 -287
rect -5541 -333 -5495 -287
rect -5417 -333 -5371 -287
rect -5293 -333 -5247 -287
rect -5169 -333 -5123 -287
rect -5045 -333 -4999 -287
rect -4921 -333 -4875 -287
rect -4797 -333 -4751 -287
rect -4673 -333 -4627 -287
rect -4549 -333 -4503 -287
rect -4425 -333 -4379 -287
rect -4301 -333 -4255 -287
rect -4177 -333 -4131 -287
rect -4053 -333 -4007 -287
rect -3929 -333 -3883 -287
rect -3805 -333 -3759 -287
rect -3681 -333 -3635 -287
rect -3557 -333 -3511 -287
rect -3433 -333 -3387 -287
rect -3309 -333 -3263 -287
rect -3185 -333 -3139 -287
rect -3061 -333 -3015 -287
rect -2937 -333 -2891 -287
rect -2813 -333 -2767 -287
rect -2689 -333 -2643 -287
rect -2565 -333 -2519 -287
rect -2441 -333 -2395 -287
rect -2317 -333 -2271 -287
rect -2193 -333 -2147 -287
rect -2069 -333 -2023 -287
rect -1945 -333 -1899 -287
rect -1821 -333 -1775 -287
rect -1697 -333 -1651 -287
rect -1573 -333 -1527 -287
rect -1449 -333 -1403 -287
rect -1325 -333 -1279 -287
rect -1201 -333 -1155 -287
rect -1077 -333 -1031 -287
rect -953 -333 -907 -287
rect -829 -333 -783 -287
rect -705 -333 -659 -287
rect -581 -333 -535 -287
rect -457 -333 -411 -287
rect -333 -333 -287 -287
rect -209 -333 -163 -287
rect -85 -333 -39 -287
rect 39 -333 85 -287
rect 163 -333 209 -287
rect 287 -333 333 -287
rect 411 -333 457 -287
rect 535 -333 581 -287
rect 659 -333 705 -287
rect 783 -333 829 -287
rect 907 -333 953 -287
rect 1031 -333 1077 -287
rect 1155 -333 1201 -287
rect 1279 -333 1325 -287
rect 1403 -333 1449 -287
rect 1527 -333 1573 -287
rect 1651 -333 1697 -287
rect 1775 -333 1821 -287
rect 1899 -333 1945 -287
rect 2023 -333 2069 -287
rect 2147 -333 2193 -287
rect 2271 -333 2317 -287
rect 2395 -333 2441 -287
rect 2519 -333 2565 -287
rect 2643 -333 2689 -287
rect 2767 -333 2813 -287
rect 2891 -333 2937 -287
rect 3015 -333 3061 -287
rect 3139 -333 3185 -287
rect 3263 -333 3309 -287
rect 3387 -333 3433 -287
rect 3511 -333 3557 -287
rect 3635 -333 3681 -287
rect 3759 -333 3805 -287
rect 3883 -333 3929 -287
rect 4007 -333 4053 -287
rect 4131 -333 4177 -287
rect 4255 -333 4301 -287
rect 4379 -333 4425 -287
rect 4503 -333 4549 -287
rect 4627 -333 4673 -287
rect 4751 -333 4797 -287
rect 4875 -333 4921 -287
rect 4999 -333 5045 -287
rect 5123 -333 5169 -287
rect 5247 -333 5293 -287
rect 5371 -333 5417 -287
rect 5495 -333 5541 -287
rect 5619 -333 5665 -287
rect 5743 -333 5789 -287
rect 5867 -333 5913 -287
rect 5991 -333 6037 -287
rect 6115 -333 6161 -287
rect 6239 -333 6285 -287
rect 6363 -333 6409 -287
rect 6487 -333 6533 -287
rect 6611 -333 6657 -287
rect 6735 -333 6781 -287
rect 6859 -333 6905 -287
rect 6983 -333 7029 -287
rect 7107 -333 7153 -287
rect 7231 -333 7277 -287
rect 7355 -333 7401 -287
rect 7479 -333 7525 -287
rect 7603 -333 7649 -287
rect 7727 -333 7773 -287
rect 7851 -333 7897 -287
rect 7975 -333 8021 -287
rect 8099 -333 8145 -287
rect 8223 -333 8269 -287
rect 8347 -333 8393 -287
rect 8471 -333 8517 -287
rect 8595 -333 8641 -287
rect 8719 -333 8765 -287
rect 8843 -333 8889 -287
rect 8967 -333 9013 -287
rect 9091 -333 9137 -287
rect 9215 -333 9261 -287
rect 9339 -333 9385 -287
rect 9463 -333 9509 -287
rect 9587 -333 9633 -287
rect 9711 -333 9757 -287
rect 9835 -333 9881 -287
rect 9959 -333 10005 -287
rect 10083 -333 10129 -287
rect 10207 -333 10253 -287
rect 10331 -333 10377 -287
rect 10455 -333 10501 -287
rect 10579 -333 10625 -287
rect 10703 -333 10749 -287
rect 10827 -333 10873 -287
rect 10951 -333 10997 -287
rect 11075 -333 11121 -287
rect 11199 -333 11245 -287
rect 11323 -333 11369 -287
rect 11447 -333 11493 -287
rect 11571 -333 11617 -287
rect 11695 -333 11741 -287
rect 11819 -333 11865 -287
rect 11943 -333 11989 -287
rect 12067 -333 12113 -287
rect 12191 -333 12237 -287
rect 12315 -333 12361 -287
rect 12439 -333 12485 -287
rect 12563 -333 12609 -287
rect 12687 -333 12733 -287
rect 12811 -333 12857 -287
rect 12935 -333 12981 -287
rect 13059 -333 13105 -287
rect 13183 -333 13229 -287
rect 13307 -333 13353 -287
rect 13431 -333 13477 -287
rect 13555 -333 13601 -287
rect 13679 -333 13725 -287
rect 13803 -333 13849 -287
rect 13927 -333 13973 -287
rect 14051 -333 14097 -287
rect 14175 -333 14221 -287
rect 14299 -333 14345 -287
rect 14423 -333 14469 -287
rect 14547 -333 14593 -287
rect 14671 -333 14717 -287
rect 14795 -333 14841 -287
rect 14919 -333 14965 -287
rect 15043 -333 15089 -287
rect 15167 -333 15213 -287
rect 15291 -333 15337 -287
rect 15415 -333 15461 -287
rect 15539 -333 15585 -287
rect 15663 -333 15709 -287
rect 15787 -333 15833 -287
rect 15911 -333 15957 -287
rect 16035 -333 16081 -287
rect 16159 -333 16205 -287
rect 16283 -333 16329 -287
rect 16407 -333 16453 -287
rect 16531 -333 16577 -287
rect 16655 -333 16701 -287
rect 16779 -333 16825 -287
rect 16903 -333 16949 -287
rect 17027 -333 17073 -287
rect 17151 -333 17197 -287
rect 17275 -333 17321 -287
rect -17321 -457 -17275 -411
rect -17197 -457 -17151 -411
rect -17073 -457 -17027 -411
rect -16949 -457 -16903 -411
rect -16825 -457 -16779 -411
rect -16701 -457 -16655 -411
rect -16577 -457 -16531 -411
rect -16453 -457 -16407 -411
rect -16329 -457 -16283 -411
rect -16205 -457 -16159 -411
rect -16081 -457 -16035 -411
rect -15957 -457 -15911 -411
rect -15833 -457 -15787 -411
rect -15709 -457 -15663 -411
rect -15585 -457 -15539 -411
rect -15461 -457 -15415 -411
rect -15337 -457 -15291 -411
rect -15213 -457 -15167 -411
rect -15089 -457 -15043 -411
rect -14965 -457 -14919 -411
rect -14841 -457 -14795 -411
rect -14717 -457 -14671 -411
rect -14593 -457 -14547 -411
rect -14469 -457 -14423 -411
rect -14345 -457 -14299 -411
rect -14221 -457 -14175 -411
rect -14097 -457 -14051 -411
rect -13973 -457 -13927 -411
rect -13849 -457 -13803 -411
rect -13725 -457 -13679 -411
rect -13601 -457 -13555 -411
rect -13477 -457 -13431 -411
rect -13353 -457 -13307 -411
rect -13229 -457 -13183 -411
rect -13105 -457 -13059 -411
rect -12981 -457 -12935 -411
rect -12857 -457 -12811 -411
rect -12733 -457 -12687 -411
rect -12609 -457 -12563 -411
rect -12485 -457 -12439 -411
rect -12361 -457 -12315 -411
rect -12237 -457 -12191 -411
rect -12113 -457 -12067 -411
rect -11989 -457 -11943 -411
rect -11865 -457 -11819 -411
rect -11741 -457 -11695 -411
rect -11617 -457 -11571 -411
rect -11493 -457 -11447 -411
rect -11369 -457 -11323 -411
rect -11245 -457 -11199 -411
rect -11121 -457 -11075 -411
rect -10997 -457 -10951 -411
rect -10873 -457 -10827 -411
rect -10749 -457 -10703 -411
rect -10625 -457 -10579 -411
rect -10501 -457 -10455 -411
rect -10377 -457 -10331 -411
rect -10253 -457 -10207 -411
rect -10129 -457 -10083 -411
rect -10005 -457 -9959 -411
rect -9881 -457 -9835 -411
rect -9757 -457 -9711 -411
rect -9633 -457 -9587 -411
rect -9509 -457 -9463 -411
rect -9385 -457 -9339 -411
rect -9261 -457 -9215 -411
rect -9137 -457 -9091 -411
rect -9013 -457 -8967 -411
rect -8889 -457 -8843 -411
rect -8765 -457 -8719 -411
rect -8641 -457 -8595 -411
rect -8517 -457 -8471 -411
rect -8393 -457 -8347 -411
rect -8269 -457 -8223 -411
rect -8145 -457 -8099 -411
rect -8021 -457 -7975 -411
rect -7897 -457 -7851 -411
rect -7773 -457 -7727 -411
rect -7649 -457 -7603 -411
rect -7525 -457 -7479 -411
rect -7401 -457 -7355 -411
rect -7277 -457 -7231 -411
rect -7153 -457 -7107 -411
rect -7029 -457 -6983 -411
rect -6905 -457 -6859 -411
rect -6781 -457 -6735 -411
rect -6657 -457 -6611 -411
rect -6533 -457 -6487 -411
rect -6409 -457 -6363 -411
rect -6285 -457 -6239 -411
rect -6161 -457 -6115 -411
rect -6037 -457 -5991 -411
rect -5913 -457 -5867 -411
rect -5789 -457 -5743 -411
rect -5665 -457 -5619 -411
rect -5541 -457 -5495 -411
rect -5417 -457 -5371 -411
rect -5293 -457 -5247 -411
rect -5169 -457 -5123 -411
rect -5045 -457 -4999 -411
rect -4921 -457 -4875 -411
rect -4797 -457 -4751 -411
rect -4673 -457 -4627 -411
rect -4549 -457 -4503 -411
rect -4425 -457 -4379 -411
rect -4301 -457 -4255 -411
rect -4177 -457 -4131 -411
rect -4053 -457 -4007 -411
rect -3929 -457 -3883 -411
rect -3805 -457 -3759 -411
rect -3681 -457 -3635 -411
rect -3557 -457 -3511 -411
rect -3433 -457 -3387 -411
rect -3309 -457 -3263 -411
rect -3185 -457 -3139 -411
rect -3061 -457 -3015 -411
rect -2937 -457 -2891 -411
rect -2813 -457 -2767 -411
rect -2689 -457 -2643 -411
rect -2565 -457 -2519 -411
rect -2441 -457 -2395 -411
rect -2317 -457 -2271 -411
rect -2193 -457 -2147 -411
rect -2069 -457 -2023 -411
rect -1945 -457 -1899 -411
rect -1821 -457 -1775 -411
rect -1697 -457 -1651 -411
rect -1573 -457 -1527 -411
rect -1449 -457 -1403 -411
rect -1325 -457 -1279 -411
rect -1201 -457 -1155 -411
rect -1077 -457 -1031 -411
rect -953 -457 -907 -411
rect -829 -457 -783 -411
rect -705 -457 -659 -411
rect -581 -457 -535 -411
rect -457 -457 -411 -411
rect -333 -457 -287 -411
rect -209 -457 -163 -411
rect -85 -457 -39 -411
rect 39 -457 85 -411
rect 163 -457 209 -411
rect 287 -457 333 -411
rect 411 -457 457 -411
rect 535 -457 581 -411
rect 659 -457 705 -411
rect 783 -457 829 -411
rect 907 -457 953 -411
rect 1031 -457 1077 -411
rect 1155 -457 1201 -411
rect 1279 -457 1325 -411
rect 1403 -457 1449 -411
rect 1527 -457 1573 -411
rect 1651 -457 1697 -411
rect 1775 -457 1821 -411
rect 1899 -457 1945 -411
rect 2023 -457 2069 -411
rect 2147 -457 2193 -411
rect 2271 -457 2317 -411
rect 2395 -457 2441 -411
rect 2519 -457 2565 -411
rect 2643 -457 2689 -411
rect 2767 -457 2813 -411
rect 2891 -457 2937 -411
rect 3015 -457 3061 -411
rect 3139 -457 3185 -411
rect 3263 -457 3309 -411
rect 3387 -457 3433 -411
rect 3511 -457 3557 -411
rect 3635 -457 3681 -411
rect 3759 -457 3805 -411
rect 3883 -457 3929 -411
rect 4007 -457 4053 -411
rect 4131 -457 4177 -411
rect 4255 -457 4301 -411
rect 4379 -457 4425 -411
rect 4503 -457 4549 -411
rect 4627 -457 4673 -411
rect 4751 -457 4797 -411
rect 4875 -457 4921 -411
rect 4999 -457 5045 -411
rect 5123 -457 5169 -411
rect 5247 -457 5293 -411
rect 5371 -457 5417 -411
rect 5495 -457 5541 -411
rect 5619 -457 5665 -411
rect 5743 -457 5789 -411
rect 5867 -457 5913 -411
rect 5991 -457 6037 -411
rect 6115 -457 6161 -411
rect 6239 -457 6285 -411
rect 6363 -457 6409 -411
rect 6487 -457 6533 -411
rect 6611 -457 6657 -411
rect 6735 -457 6781 -411
rect 6859 -457 6905 -411
rect 6983 -457 7029 -411
rect 7107 -457 7153 -411
rect 7231 -457 7277 -411
rect 7355 -457 7401 -411
rect 7479 -457 7525 -411
rect 7603 -457 7649 -411
rect 7727 -457 7773 -411
rect 7851 -457 7897 -411
rect 7975 -457 8021 -411
rect 8099 -457 8145 -411
rect 8223 -457 8269 -411
rect 8347 -457 8393 -411
rect 8471 -457 8517 -411
rect 8595 -457 8641 -411
rect 8719 -457 8765 -411
rect 8843 -457 8889 -411
rect 8967 -457 9013 -411
rect 9091 -457 9137 -411
rect 9215 -457 9261 -411
rect 9339 -457 9385 -411
rect 9463 -457 9509 -411
rect 9587 -457 9633 -411
rect 9711 -457 9757 -411
rect 9835 -457 9881 -411
rect 9959 -457 10005 -411
rect 10083 -457 10129 -411
rect 10207 -457 10253 -411
rect 10331 -457 10377 -411
rect 10455 -457 10501 -411
rect 10579 -457 10625 -411
rect 10703 -457 10749 -411
rect 10827 -457 10873 -411
rect 10951 -457 10997 -411
rect 11075 -457 11121 -411
rect 11199 -457 11245 -411
rect 11323 -457 11369 -411
rect 11447 -457 11493 -411
rect 11571 -457 11617 -411
rect 11695 -457 11741 -411
rect 11819 -457 11865 -411
rect 11943 -457 11989 -411
rect 12067 -457 12113 -411
rect 12191 -457 12237 -411
rect 12315 -457 12361 -411
rect 12439 -457 12485 -411
rect 12563 -457 12609 -411
rect 12687 -457 12733 -411
rect 12811 -457 12857 -411
rect 12935 -457 12981 -411
rect 13059 -457 13105 -411
rect 13183 -457 13229 -411
rect 13307 -457 13353 -411
rect 13431 -457 13477 -411
rect 13555 -457 13601 -411
rect 13679 -457 13725 -411
rect 13803 -457 13849 -411
rect 13927 -457 13973 -411
rect 14051 -457 14097 -411
rect 14175 -457 14221 -411
rect 14299 -457 14345 -411
rect 14423 -457 14469 -411
rect 14547 -457 14593 -411
rect 14671 -457 14717 -411
rect 14795 -457 14841 -411
rect 14919 -457 14965 -411
rect 15043 -457 15089 -411
rect 15167 -457 15213 -411
rect 15291 -457 15337 -411
rect 15415 -457 15461 -411
rect 15539 -457 15585 -411
rect 15663 -457 15709 -411
rect 15787 -457 15833 -411
rect 15911 -457 15957 -411
rect 16035 -457 16081 -411
rect 16159 -457 16205 -411
rect 16283 -457 16329 -411
rect 16407 -457 16453 -411
rect 16531 -457 16577 -411
rect 16655 -457 16701 -411
rect 16779 -457 16825 -411
rect 16903 -457 16949 -411
rect 17027 -457 17073 -411
rect 17151 -457 17197 -411
rect 17275 -457 17321 -411
rect -17321 -581 -17275 -535
rect -17197 -581 -17151 -535
rect -17073 -581 -17027 -535
rect -16949 -581 -16903 -535
rect -16825 -581 -16779 -535
rect -16701 -581 -16655 -535
rect -16577 -581 -16531 -535
rect -16453 -581 -16407 -535
rect -16329 -581 -16283 -535
rect -16205 -581 -16159 -535
rect -16081 -581 -16035 -535
rect -15957 -581 -15911 -535
rect -15833 -581 -15787 -535
rect -15709 -581 -15663 -535
rect -15585 -581 -15539 -535
rect -15461 -581 -15415 -535
rect -15337 -581 -15291 -535
rect -15213 -581 -15167 -535
rect -15089 -581 -15043 -535
rect -14965 -581 -14919 -535
rect -14841 -581 -14795 -535
rect -14717 -581 -14671 -535
rect -14593 -581 -14547 -535
rect -14469 -581 -14423 -535
rect -14345 -581 -14299 -535
rect -14221 -581 -14175 -535
rect -14097 -581 -14051 -535
rect -13973 -581 -13927 -535
rect -13849 -581 -13803 -535
rect -13725 -581 -13679 -535
rect -13601 -581 -13555 -535
rect -13477 -581 -13431 -535
rect -13353 -581 -13307 -535
rect -13229 -581 -13183 -535
rect -13105 -581 -13059 -535
rect -12981 -581 -12935 -535
rect -12857 -581 -12811 -535
rect -12733 -581 -12687 -535
rect -12609 -581 -12563 -535
rect -12485 -581 -12439 -535
rect -12361 -581 -12315 -535
rect -12237 -581 -12191 -535
rect -12113 -581 -12067 -535
rect -11989 -581 -11943 -535
rect -11865 -581 -11819 -535
rect -11741 -581 -11695 -535
rect -11617 -581 -11571 -535
rect -11493 -581 -11447 -535
rect -11369 -581 -11323 -535
rect -11245 -581 -11199 -535
rect -11121 -581 -11075 -535
rect -10997 -581 -10951 -535
rect -10873 -581 -10827 -535
rect -10749 -581 -10703 -535
rect -10625 -581 -10579 -535
rect -10501 -581 -10455 -535
rect -10377 -581 -10331 -535
rect -10253 -581 -10207 -535
rect -10129 -581 -10083 -535
rect -10005 -581 -9959 -535
rect -9881 -581 -9835 -535
rect -9757 -581 -9711 -535
rect -9633 -581 -9587 -535
rect -9509 -581 -9463 -535
rect -9385 -581 -9339 -535
rect -9261 -581 -9215 -535
rect -9137 -581 -9091 -535
rect -9013 -581 -8967 -535
rect -8889 -581 -8843 -535
rect -8765 -581 -8719 -535
rect -8641 -581 -8595 -535
rect -8517 -581 -8471 -535
rect -8393 -581 -8347 -535
rect -8269 -581 -8223 -535
rect -8145 -581 -8099 -535
rect -8021 -581 -7975 -535
rect -7897 -581 -7851 -535
rect -7773 -581 -7727 -535
rect -7649 -581 -7603 -535
rect -7525 -581 -7479 -535
rect -7401 -581 -7355 -535
rect -7277 -581 -7231 -535
rect -7153 -581 -7107 -535
rect -7029 -581 -6983 -535
rect -6905 -581 -6859 -535
rect -6781 -581 -6735 -535
rect -6657 -581 -6611 -535
rect -6533 -581 -6487 -535
rect -6409 -581 -6363 -535
rect -6285 -581 -6239 -535
rect -6161 -581 -6115 -535
rect -6037 -581 -5991 -535
rect -5913 -581 -5867 -535
rect -5789 -581 -5743 -535
rect -5665 -581 -5619 -535
rect -5541 -581 -5495 -535
rect -5417 -581 -5371 -535
rect -5293 -581 -5247 -535
rect -5169 -581 -5123 -535
rect -5045 -581 -4999 -535
rect -4921 -581 -4875 -535
rect -4797 -581 -4751 -535
rect -4673 -581 -4627 -535
rect -4549 -581 -4503 -535
rect -4425 -581 -4379 -535
rect -4301 -581 -4255 -535
rect -4177 -581 -4131 -535
rect -4053 -581 -4007 -535
rect -3929 -581 -3883 -535
rect -3805 -581 -3759 -535
rect -3681 -581 -3635 -535
rect -3557 -581 -3511 -535
rect -3433 -581 -3387 -535
rect -3309 -581 -3263 -535
rect -3185 -581 -3139 -535
rect -3061 -581 -3015 -535
rect -2937 -581 -2891 -535
rect -2813 -581 -2767 -535
rect -2689 -581 -2643 -535
rect -2565 -581 -2519 -535
rect -2441 -581 -2395 -535
rect -2317 -581 -2271 -535
rect -2193 -581 -2147 -535
rect -2069 -581 -2023 -535
rect -1945 -581 -1899 -535
rect -1821 -581 -1775 -535
rect -1697 -581 -1651 -535
rect -1573 -581 -1527 -535
rect -1449 -581 -1403 -535
rect -1325 -581 -1279 -535
rect -1201 -581 -1155 -535
rect -1077 -581 -1031 -535
rect -953 -581 -907 -535
rect -829 -581 -783 -535
rect -705 -581 -659 -535
rect -581 -581 -535 -535
rect -457 -581 -411 -535
rect -333 -581 -287 -535
rect -209 -581 -163 -535
rect -85 -581 -39 -535
rect 39 -581 85 -535
rect 163 -581 209 -535
rect 287 -581 333 -535
rect 411 -581 457 -535
rect 535 -581 581 -535
rect 659 -581 705 -535
rect 783 -581 829 -535
rect 907 -581 953 -535
rect 1031 -581 1077 -535
rect 1155 -581 1201 -535
rect 1279 -581 1325 -535
rect 1403 -581 1449 -535
rect 1527 -581 1573 -535
rect 1651 -581 1697 -535
rect 1775 -581 1821 -535
rect 1899 -581 1945 -535
rect 2023 -581 2069 -535
rect 2147 -581 2193 -535
rect 2271 -581 2317 -535
rect 2395 -581 2441 -535
rect 2519 -581 2565 -535
rect 2643 -581 2689 -535
rect 2767 -581 2813 -535
rect 2891 -581 2937 -535
rect 3015 -581 3061 -535
rect 3139 -581 3185 -535
rect 3263 -581 3309 -535
rect 3387 -581 3433 -535
rect 3511 -581 3557 -535
rect 3635 -581 3681 -535
rect 3759 -581 3805 -535
rect 3883 -581 3929 -535
rect 4007 -581 4053 -535
rect 4131 -581 4177 -535
rect 4255 -581 4301 -535
rect 4379 -581 4425 -535
rect 4503 -581 4549 -535
rect 4627 -581 4673 -535
rect 4751 -581 4797 -535
rect 4875 -581 4921 -535
rect 4999 -581 5045 -535
rect 5123 -581 5169 -535
rect 5247 -581 5293 -535
rect 5371 -581 5417 -535
rect 5495 -581 5541 -535
rect 5619 -581 5665 -535
rect 5743 -581 5789 -535
rect 5867 -581 5913 -535
rect 5991 -581 6037 -535
rect 6115 -581 6161 -535
rect 6239 -581 6285 -535
rect 6363 -581 6409 -535
rect 6487 -581 6533 -535
rect 6611 -581 6657 -535
rect 6735 -581 6781 -535
rect 6859 -581 6905 -535
rect 6983 -581 7029 -535
rect 7107 -581 7153 -535
rect 7231 -581 7277 -535
rect 7355 -581 7401 -535
rect 7479 -581 7525 -535
rect 7603 -581 7649 -535
rect 7727 -581 7773 -535
rect 7851 -581 7897 -535
rect 7975 -581 8021 -535
rect 8099 -581 8145 -535
rect 8223 -581 8269 -535
rect 8347 -581 8393 -535
rect 8471 -581 8517 -535
rect 8595 -581 8641 -535
rect 8719 -581 8765 -535
rect 8843 -581 8889 -535
rect 8967 -581 9013 -535
rect 9091 -581 9137 -535
rect 9215 -581 9261 -535
rect 9339 -581 9385 -535
rect 9463 -581 9509 -535
rect 9587 -581 9633 -535
rect 9711 -581 9757 -535
rect 9835 -581 9881 -535
rect 9959 -581 10005 -535
rect 10083 -581 10129 -535
rect 10207 -581 10253 -535
rect 10331 -581 10377 -535
rect 10455 -581 10501 -535
rect 10579 -581 10625 -535
rect 10703 -581 10749 -535
rect 10827 -581 10873 -535
rect 10951 -581 10997 -535
rect 11075 -581 11121 -535
rect 11199 -581 11245 -535
rect 11323 -581 11369 -535
rect 11447 -581 11493 -535
rect 11571 -581 11617 -535
rect 11695 -581 11741 -535
rect 11819 -581 11865 -535
rect 11943 -581 11989 -535
rect 12067 -581 12113 -535
rect 12191 -581 12237 -535
rect 12315 -581 12361 -535
rect 12439 -581 12485 -535
rect 12563 -581 12609 -535
rect 12687 -581 12733 -535
rect 12811 -581 12857 -535
rect 12935 -581 12981 -535
rect 13059 -581 13105 -535
rect 13183 -581 13229 -535
rect 13307 -581 13353 -535
rect 13431 -581 13477 -535
rect 13555 -581 13601 -535
rect 13679 -581 13725 -535
rect 13803 -581 13849 -535
rect 13927 -581 13973 -535
rect 14051 -581 14097 -535
rect 14175 -581 14221 -535
rect 14299 -581 14345 -535
rect 14423 -581 14469 -535
rect 14547 -581 14593 -535
rect 14671 -581 14717 -535
rect 14795 -581 14841 -535
rect 14919 -581 14965 -535
rect 15043 -581 15089 -535
rect 15167 -581 15213 -535
rect 15291 -581 15337 -535
rect 15415 -581 15461 -535
rect 15539 -581 15585 -535
rect 15663 -581 15709 -535
rect 15787 -581 15833 -535
rect 15911 -581 15957 -535
rect 16035 -581 16081 -535
rect 16159 -581 16205 -535
rect 16283 -581 16329 -535
rect 16407 -581 16453 -535
rect 16531 -581 16577 -535
rect 16655 -581 16701 -535
rect 16779 -581 16825 -535
rect 16903 -581 16949 -535
rect 17027 -581 17073 -535
rect 17151 -581 17197 -535
rect 17275 -581 17321 -535
rect -17321 -705 -17275 -659
rect -17197 -705 -17151 -659
rect -17073 -705 -17027 -659
rect -16949 -705 -16903 -659
rect -16825 -705 -16779 -659
rect -16701 -705 -16655 -659
rect -16577 -705 -16531 -659
rect -16453 -705 -16407 -659
rect -16329 -705 -16283 -659
rect -16205 -705 -16159 -659
rect -16081 -705 -16035 -659
rect -15957 -705 -15911 -659
rect -15833 -705 -15787 -659
rect -15709 -705 -15663 -659
rect -15585 -705 -15539 -659
rect -15461 -705 -15415 -659
rect -15337 -705 -15291 -659
rect -15213 -705 -15167 -659
rect -15089 -705 -15043 -659
rect -14965 -705 -14919 -659
rect -14841 -705 -14795 -659
rect -14717 -705 -14671 -659
rect -14593 -705 -14547 -659
rect -14469 -705 -14423 -659
rect -14345 -705 -14299 -659
rect -14221 -705 -14175 -659
rect -14097 -705 -14051 -659
rect -13973 -705 -13927 -659
rect -13849 -705 -13803 -659
rect -13725 -705 -13679 -659
rect -13601 -705 -13555 -659
rect -13477 -705 -13431 -659
rect -13353 -705 -13307 -659
rect -13229 -705 -13183 -659
rect -13105 -705 -13059 -659
rect -12981 -705 -12935 -659
rect -12857 -705 -12811 -659
rect -12733 -705 -12687 -659
rect -12609 -705 -12563 -659
rect -12485 -705 -12439 -659
rect -12361 -705 -12315 -659
rect -12237 -705 -12191 -659
rect -12113 -705 -12067 -659
rect -11989 -705 -11943 -659
rect -11865 -705 -11819 -659
rect -11741 -705 -11695 -659
rect -11617 -705 -11571 -659
rect -11493 -705 -11447 -659
rect -11369 -705 -11323 -659
rect -11245 -705 -11199 -659
rect -11121 -705 -11075 -659
rect -10997 -705 -10951 -659
rect -10873 -705 -10827 -659
rect -10749 -705 -10703 -659
rect -10625 -705 -10579 -659
rect -10501 -705 -10455 -659
rect -10377 -705 -10331 -659
rect -10253 -705 -10207 -659
rect -10129 -705 -10083 -659
rect -10005 -705 -9959 -659
rect -9881 -705 -9835 -659
rect -9757 -705 -9711 -659
rect -9633 -705 -9587 -659
rect -9509 -705 -9463 -659
rect -9385 -705 -9339 -659
rect -9261 -705 -9215 -659
rect -9137 -705 -9091 -659
rect -9013 -705 -8967 -659
rect -8889 -705 -8843 -659
rect -8765 -705 -8719 -659
rect -8641 -705 -8595 -659
rect -8517 -705 -8471 -659
rect -8393 -705 -8347 -659
rect -8269 -705 -8223 -659
rect -8145 -705 -8099 -659
rect -8021 -705 -7975 -659
rect -7897 -705 -7851 -659
rect -7773 -705 -7727 -659
rect -7649 -705 -7603 -659
rect -7525 -705 -7479 -659
rect -7401 -705 -7355 -659
rect -7277 -705 -7231 -659
rect -7153 -705 -7107 -659
rect -7029 -705 -6983 -659
rect -6905 -705 -6859 -659
rect -6781 -705 -6735 -659
rect -6657 -705 -6611 -659
rect -6533 -705 -6487 -659
rect -6409 -705 -6363 -659
rect -6285 -705 -6239 -659
rect -6161 -705 -6115 -659
rect -6037 -705 -5991 -659
rect -5913 -705 -5867 -659
rect -5789 -705 -5743 -659
rect -5665 -705 -5619 -659
rect -5541 -705 -5495 -659
rect -5417 -705 -5371 -659
rect -5293 -705 -5247 -659
rect -5169 -705 -5123 -659
rect -5045 -705 -4999 -659
rect -4921 -705 -4875 -659
rect -4797 -705 -4751 -659
rect -4673 -705 -4627 -659
rect -4549 -705 -4503 -659
rect -4425 -705 -4379 -659
rect -4301 -705 -4255 -659
rect -4177 -705 -4131 -659
rect -4053 -705 -4007 -659
rect -3929 -705 -3883 -659
rect -3805 -705 -3759 -659
rect -3681 -705 -3635 -659
rect -3557 -705 -3511 -659
rect -3433 -705 -3387 -659
rect -3309 -705 -3263 -659
rect -3185 -705 -3139 -659
rect -3061 -705 -3015 -659
rect -2937 -705 -2891 -659
rect -2813 -705 -2767 -659
rect -2689 -705 -2643 -659
rect -2565 -705 -2519 -659
rect -2441 -705 -2395 -659
rect -2317 -705 -2271 -659
rect -2193 -705 -2147 -659
rect -2069 -705 -2023 -659
rect -1945 -705 -1899 -659
rect -1821 -705 -1775 -659
rect -1697 -705 -1651 -659
rect -1573 -705 -1527 -659
rect -1449 -705 -1403 -659
rect -1325 -705 -1279 -659
rect -1201 -705 -1155 -659
rect -1077 -705 -1031 -659
rect -953 -705 -907 -659
rect -829 -705 -783 -659
rect -705 -705 -659 -659
rect -581 -705 -535 -659
rect -457 -705 -411 -659
rect -333 -705 -287 -659
rect -209 -705 -163 -659
rect -85 -705 -39 -659
rect 39 -705 85 -659
rect 163 -705 209 -659
rect 287 -705 333 -659
rect 411 -705 457 -659
rect 535 -705 581 -659
rect 659 -705 705 -659
rect 783 -705 829 -659
rect 907 -705 953 -659
rect 1031 -705 1077 -659
rect 1155 -705 1201 -659
rect 1279 -705 1325 -659
rect 1403 -705 1449 -659
rect 1527 -705 1573 -659
rect 1651 -705 1697 -659
rect 1775 -705 1821 -659
rect 1899 -705 1945 -659
rect 2023 -705 2069 -659
rect 2147 -705 2193 -659
rect 2271 -705 2317 -659
rect 2395 -705 2441 -659
rect 2519 -705 2565 -659
rect 2643 -705 2689 -659
rect 2767 -705 2813 -659
rect 2891 -705 2937 -659
rect 3015 -705 3061 -659
rect 3139 -705 3185 -659
rect 3263 -705 3309 -659
rect 3387 -705 3433 -659
rect 3511 -705 3557 -659
rect 3635 -705 3681 -659
rect 3759 -705 3805 -659
rect 3883 -705 3929 -659
rect 4007 -705 4053 -659
rect 4131 -705 4177 -659
rect 4255 -705 4301 -659
rect 4379 -705 4425 -659
rect 4503 -705 4549 -659
rect 4627 -705 4673 -659
rect 4751 -705 4797 -659
rect 4875 -705 4921 -659
rect 4999 -705 5045 -659
rect 5123 -705 5169 -659
rect 5247 -705 5293 -659
rect 5371 -705 5417 -659
rect 5495 -705 5541 -659
rect 5619 -705 5665 -659
rect 5743 -705 5789 -659
rect 5867 -705 5913 -659
rect 5991 -705 6037 -659
rect 6115 -705 6161 -659
rect 6239 -705 6285 -659
rect 6363 -705 6409 -659
rect 6487 -705 6533 -659
rect 6611 -705 6657 -659
rect 6735 -705 6781 -659
rect 6859 -705 6905 -659
rect 6983 -705 7029 -659
rect 7107 -705 7153 -659
rect 7231 -705 7277 -659
rect 7355 -705 7401 -659
rect 7479 -705 7525 -659
rect 7603 -705 7649 -659
rect 7727 -705 7773 -659
rect 7851 -705 7897 -659
rect 7975 -705 8021 -659
rect 8099 -705 8145 -659
rect 8223 -705 8269 -659
rect 8347 -705 8393 -659
rect 8471 -705 8517 -659
rect 8595 -705 8641 -659
rect 8719 -705 8765 -659
rect 8843 -705 8889 -659
rect 8967 -705 9013 -659
rect 9091 -705 9137 -659
rect 9215 -705 9261 -659
rect 9339 -705 9385 -659
rect 9463 -705 9509 -659
rect 9587 -705 9633 -659
rect 9711 -705 9757 -659
rect 9835 -705 9881 -659
rect 9959 -705 10005 -659
rect 10083 -705 10129 -659
rect 10207 -705 10253 -659
rect 10331 -705 10377 -659
rect 10455 -705 10501 -659
rect 10579 -705 10625 -659
rect 10703 -705 10749 -659
rect 10827 -705 10873 -659
rect 10951 -705 10997 -659
rect 11075 -705 11121 -659
rect 11199 -705 11245 -659
rect 11323 -705 11369 -659
rect 11447 -705 11493 -659
rect 11571 -705 11617 -659
rect 11695 -705 11741 -659
rect 11819 -705 11865 -659
rect 11943 -705 11989 -659
rect 12067 -705 12113 -659
rect 12191 -705 12237 -659
rect 12315 -705 12361 -659
rect 12439 -705 12485 -659
rect 12563 -705 12609 -659
rect 12687 -705 12733 -659
rect 12811 -705 12857 -659
rect 12935 -705 12981 -659
rect 13059 -705 13105 -659
rect 13183 -705 13229 -659
rect 13307 -705 13353 -659
rect 13431 -705 13477 -659
rect 13555 -705 13601 -659
rect 13679 -705 13725 -659
rect 13803 -705 13849 -659
rect 13927 -705 13973 -659
rect 14051 -705 14097 -659
rect 14175 -705 14221 -659
rect 14299 -705 14345 -659
rect 14423 -705 14469 -659
rect 14547 -705 14593 -659
rect 14671 -705 14717 -659
rect 14795 -705 14841 -659
rect 14919 -705 14965 -659
rect 15043 -705 15089 -659
rect 15167 -705 15213 -659
rect 15291 -705 15337 -659
rect 15415 -705 15461 -659
rect 15539 -705 15585 -659
rect 15663 -705 15709 -659
rect 15787 -705 15833 -659
rect 15911 -705 15957 -659
rect 16035 -705 16081 -659
rect 16159 -705 16205 -659
rect 16283 -705 16329 -659
rect 16407 -705 16453 -659
rect 16531 -705 16577 -659
rect 16655 -705 16701 -659
rect 16779 -705 16825 -659
rect 16903 -705 16949 -659
rect 17027 -705 17073 -659
rect 17151 -705 17197 -659
rect 17275 -705 17321 -659
rect -17321 -829 -17275 -783
rect -17197 -829 -17151 -783
rect -17073 -829 -17027 -783
rect -16949 -829 -16903 -783
rect -16825 -829 -16779 -783
rect -16701 -829 -16655 -783
rect -16577 -829 -16531 -783
rect -16453 -829 -16407 -783
rect -16329 -829 -16283 -783
rect -16205 -829 -16159 -783
rect -16081 -829 -16035 -783
rect -15957 -829 -15911 -783
rect -15833 -829 -15787 -783
rect -15709 -829 -15663 -783
rect -15585 -829 -15539 -783
rect -15461 -829 -15415 -783
rect -15337 -829 -15291 -783
rect -15213 -829 -15167 -783
rect -15089 -829 -15043 -783
rect -14965 -829 -14919 -783
rect -14841 -829 -14795 -783
rect -14717 -829 -14671 -783
rect -14593 -829 -14547 -783
rect -14469 -829 -14423 -783
rect -14345 -829 -14299 -783
rect -14221 -829 -14175 -783
rect -14097 -829 -14051 -783
rect -13973 -829 -13927 -783
rect -13849 -829 -13803 -783
rect -13725 -829 -13679 -783
rect -13601 -829 -13555 -783
rect -13477 -829 -13431 -783
rect -13353 -829 -13307 -783
rect -13229 -829 -13183 -783
rect -13105 -829 -13059 -783
rect -12981 -829 -12935 -783
rect -12857 -829 -12811 -783
rect -12733 -829 -12687 -783
rect -12609 -829 -12563 -783
rect -12485 -829 -12439 -783
rect -12361 -829 -12315 -783
rect -12237 -829 -12191 -783
rect -12113 -829 -12067 -783
rect -11989 -829 -11943 -783
rect -11865 -829 -11819 -783
rect -11741 -829 -11695 -783
rect -11617 -829 -11571 -783
rect -11493 -829 -11447 -783
rect -11369 -829 -11323 -783
rect -11245 -829 -11199 -783
rect -11121 -829 -11075 -783
rect -10997 -829 -10951 -783
rect -10873 -829 -10827 -783
rect -10749 -829 -10703 -783
rect -10625 -829 -10579 -783
rect -10501 -829 -10455 -783
rect -10377 -829 -10331 -783
rect -10253 -829 -10207 -783
rect -10129 -829 -10083 -783
rect -10005 -829 -9959 -783
rect -9881 -829 -9835 -783
rect -9757 -829 -9711 -783
rect -9633 -829 -9587 -783
rect -9509 -829 -9463 -783
rect -9385 -829 -9339 -783
rect -9261 -829 -9215 -783
rect -9137 -829 -9091 -783
rect -9013 -829 -8967 -783
rect -8889 -829 -8843 -783
rect -8765 -829 -8719 -783
rect -8641 -829 -8595 -783
rect -8517 -829 -8471 -783
rect -8393 -829 -8347 -783
rect -8269 -829 -8223 -783
rect -8145 -829 -8099 -783
rect -8021 -829 -7975 -783
rect -7897 -829 -7851 -783
rect -7773 -829 -7727 -783
rect -7649 -829 -7603 -783
rect -7525 -829 -7479 -783
rect -7401 -829 -7355 -783
rect -7277 -829 -7231 -783
rect -7153 -829 -7107 -783
rect -7029 -829 -6983 -783
rect -6905 -829 -6859 -783
rect -6781 -829 -6735 -783
rect -6657 -829 -6611 -783
rect -6533 -829 -6487 -783
rect -6409 -829 -6363 -783
rect -6285 -829 -6239 -783
rect -6161 -829 -6115 -783
rect -6037 -829 -5991 -783
rect -5913 -829 -5867 -783
rect -5789 -829 -5743 -783
rect -5665 -829 -5619 -783
rect -5541 -829 -5495 -783
rect -5417 -829 -5371 -783
rect -5293 -829 -5247 -783
rect -5169 -829 -5123 -783
rect -5045 -829 -4999 -783
rect -4921 -829 -4875 -783
rect -4797 -829 -4751 -783
rect -4673 -829 -4627 -783
rect -4549 -829 -4503 -783
rect -4425 -829 -4379 -783
rect -4301 -829 -4255 -783
rect -4177 -829 -4131 -783
rect -4053 -829 -4007 -783
rect -3929 -829 -3883 -783
rect -3805 -829 -3759 -783
rect -3681 -829 -3635 -783
rect -3557 -829 -3511 -783
rect -3433 -829 -3387 -783
rect -3309 -829 -3263 -783
rect -3185 -829 -3139 -783
rect -3061 -829 -3015 -783
rect -2937 -829 -2891 -783
rect -2813 -829 -2767 -783
rect -2689 -829 -2643 -783
rect -2565 -829 -2519 -783
rect -2441 -829 -2395 -783
rect -2317 -829 -2271 -783
rect -2193 -829 -2147 -783
rect -2069 -829 -2023 -783
rect -1945 -829 -1899 -783
rect -1821 -829 -1775 -783
rect -1697 -829 -1651 -783
rect -1573 -829 -1527 -783
rect -1449 -829 -1403 -783
rect -1325 -829 -1279 -783
rect -1201 -829 -1155 -783
rect -1077 -829 -1031 -783
rect -953 -829 -907 -783
rect -829 -829 -783 -783
rect -705 -829 -659 -783
rect -581 -829 -535 -783
rect -457 -829 -411 -783
rect -333 -829 -287 -783
rect -209 -829 -163 -783
rect -85 -829 -39 -783
rect 39 -829 85 -783
rect 163 -829 209 -783
rect 287 -829 333 -783
rect 411 -829 457 -783
rect 535 -829 581 -783
rect 659 -829 705 -783
rect 783 -829 829 -783
rect 907 -829 953 -783
rect 1031 -829 1077 -783
rect 1155 -829 1201 -783
rect 1279 -829 1325 -783
rect 1403 -829 1449 -783
rect 1527 -829 1573 -783
rect 1651 -829 1697 -783
rect 1775 -829 1821 -783
rect 1899 -829 1945 -783
rect 2023 -829 2069 -783
rect 2147 -829 2193 -783
rect 2271 -829 2317 -783
rect 2395 -829 2441 -783
rect 2519 -829 2565 -783
rect 2643 -829 2689 -783
rect 2767 -829 2813 -783
rect 2891 -829 2937 -783
rect 3015 -829 3061 -783
rect 3139 -829 3185 -783
rect 3263 -829 3309 -783
rect 3387 -829 3433 -783
rect 3511 -829 3557 -783
rect 3635 -829 3681 -783
rect 3759 -829 3805 -783
rect 3883 -829 3929 -783
rect 4007 -829 4053 -783
rect 4131 -829 4177 -783
rect 4255 -829 4301 -783
rect 4379 -829 4425 -783
rect 4503 -829 4549 -783
rect 4627 -829 4673 -783
rect 4751 -829 4797 -783
rect 4875 -829 4921 -783
rect 4999 -829 5045 -783
rect 5123 -829 5169 -783
rect 5247 -829 5293 -783
rect 5371 -829 5417 -783
rect 5495 -829 5541 -783
rect 5619 -829 5665 -783
rect 5743 -829 5789 -783
rect 5867 -829 5913 -783
rect 5991 -829 6037 -783
rect 6115 -829 6161 -783
rect 6239 -829 6285 -783
rect 6363 -829 6409 -783
rect 6487 -829 6533 -783
rect 6611 -829 6657 -783
rect 6735 -829 6781 -783
rect 6859 -829 6905 -783
rect 6983 -829 7029 -783
rect 7107 -829 7153 -783
rect 7231 -829 7277 -783
rect 7355 -829 7401 -783
rect 7479 -829 7525 -783
rect 7603 -829 7649 -783
rect 7727 -829 7773 -783
rect 7851 -829 7897 -783
rect 7975 -829 8021 -783
rect 8099 -829 8145 -783
rect 8223 -829 8269 -783
rect 8347 -829 8393 -783
rect 8471 -829 8517 -783
rect 8595 -829 8641 -783
rect 8719 -829 8765 -783
rect 8843 -829 8889 -783
rect 8967 -829 9013 -783
rect 9091 -829 9137 -783
rect 9215 -829 9261 -783
rect 9339 -829 9385 -783
rect 9463 -829 9509 -783
rect 9587 -829 9633 -783
rect 9711 -829 9757 -783
rect 9835 -829 9881 -783
rect 9959 -829 10005 -783
rect 10083 -829 10129 -783
rect 10207 -829 10253 -783
rect 10331 -829 10377 -783
rect 10455 -829 10501 -783
rect 10579 -829 10625 -783
rect 10703 -829 10749 -783
rect 10827 -829 10873 -783
rect 10951 -829 10997 -783
rect 11075 -829 11121 -783
rect 11199 -829 11245 -783
rect 11323 -829 11369 -783
rect 11447 -829 11493 -783
rect 11571 -829 11617 -783
rect 11695 -829 11741 -783
rect 11819 -829 11865 -783
rect 11943 -829 11989 -783
rect 12067 -829 12113 -783
rect 12191 -829 12237 -783
rect 12315 -829 12361 -783
rect 12439 -829 12485 -783
rect 12563 -829 12609 -783
rect 12687 -829 12733 -783
rect 12811 -829 12857 -783
rect 12935 -829 12981 -783
rect 13059 -829 13105 -783
rect 13183 -829 13229 -783
rect 13307 -829 13353 -783
rect 13431 -829 13477 -783
rect 13555 -829 13601 -783
rect 13679 -829 13725 -783
rect 13803 -829 13849 -783
rect 13927 -829 13973 -783
rect 14051 -829 14097 -783
rect 14175 -829 14221 -783
rect 14299 -829 14345 -783
rect 14423 -829 14469 -783
rect 14547 -829 14593 -783
rect 14671 -829 14717 -783
rect 14795 -829 14841 -783
rect 14919 -829 14965 -783
rect 15043 -829 15089 -783
rect 15167 -829 15213 -783
rect 15291 -829 15337 -783
rect 15415 -829 15461 -783
rect 15539 -829 15585 -783
rect 15663 -829 15709 -783
rect 15787 -829 15833 -783
rect 15911 -829 15957 -783
rect 16035 -829 16081 -783
rect 16159 -829 16205 -783
rect 16283 -829 16329 -783
rect 16407 -829 16453 -783
rect 16531 -829 16577 -783
rect 16655 -829 16701 -783
rect 16779 -829 16825 -783
rect 16903 -829 16949 -783
rect 17027 -829 17073 -783
rect 17151 -829 17197 -783
rect 17275 -829 17321 -783
rect -17321 -953 -17275 -907
rect -17197 -953 -17151 -907
rect -17073 -953 -17027 -907
rect -16949 -953 -16903 -907
rect -16825 -953 -16779 -907
rect -16701 -953 -16655 -907
rect -16577 -953 -16531 -907
rect -16453 -953 -16407 -907
rect -16329 -953 -16283 -907
rect -16205 -953 -16159 -907
rect -16081 -953 -16035 -907
rect -15957 -953 -15911 -907
rect -15833 -953 -15787 -907
rect -15709 -953 -15663 -907
rect -15585 -953 -15539 -907
rect -15461 -953 -15415 -907
rect -15337 -953 -15291 -907
rect -15213 -953 -15167 -907
rect -15089 -953 -15043 -907
rect -14965 -953 -14919 -907
rect -14841 -953 -14795 -907
rect -14717 -953 -14671 -907
rect -14593 -953 -14547 -907
rect -14469 -953 -14423 -907
rect -14345 -953 -14299 -907
rect -14221 -953 -14175 -907
rect -14097 -953 -14051 -907
rect -13973 -953 -13927 -907
rect -13849 -953 -13803 -907
rect -13725 -953 -13679 -907
rect -13601 -953 -13555 -907
rect -13477 -953 -13431 -907
rect -13353 -953 -13307 -907
rect -13229 -953 -13183 -907
rect -13105 -953 -13059 -907
rect -12981 -953 -12935 -907
rect -12857 -953 -12811 -907
rect -12733 -953 -12687 -907
rect -12609 -953 -12563 -907
rect -12485 -953 -12439 -907
rect -12361 -953 -12315 -907
rect -12237 -953 -12191 -907
rect -12113 -953 -12067 -907
rect -11989 -953 -11943 -907
rect -11865 -953 -11819 -907
rect -11741 -953 -11695 -907
rect -11617 -953 -11571 -907
rect -11493 -953 -11447 -907
rect -11369 -953 -11323 -907
rect -11245 -953 -11199 -907
rect -11121 -953 -11075 -907
rect -10997 -953 -10951 -907
rect -10873 -953 -10827 -907
rect -10749 -953 -10703 -907
rect -10625 -953 -10579 -907
rect -10501 -953 -10455 -907
rect -10377 -953 -10331 -907
rect -10253 -953 -10207 -907
rect -10129 -953 -10083 -907
rect -10005 -953 -9959 -907
rect -9881 -953 -9835 -907
rect -9757 -953 -9711 -907
rect -9633 -953 -9587 -907
rect -9509 -953 -9463 -907
rect -9385 -953 -9339 -907
rect -9261 -953 -9215 -907
rect -9137 -953 -9091 -907
rect -9013 -953 -8967 -907
rect -8889 -953 -8843 -907
rect -8765 -953 -8719 -907
rect -8641 -953 -8595 -907
rect -8517 -953 -8471 -907
rect -8393 -953 -8347 -907
rect -8269 -953 -8223 -907
rect -8145 -953 -8099 -907
rect -8021 -953 -7975 -907
rect -7897 -953 -7851 -907
rect -7773 -953 -7727 -907
rect -7649 -953 -7603 -907
rect -7525 -953 -7479 -907
rect -7401 -953 -7355 -907
rect -7277 -953 -7231 -907
rect -7153 -953 -7107 -907
rect -7029 -953 -6983 -907
rect -6905 -953 -6859 -907
rect -6781 -953 -6735 -907
rect -6657 -953 -6611 -907
rect -6533 -953 -6487 -907
rect -6409 -953 -6363 -907
rect -6285 -953 -6239 -907
rect -6161 -953 -6115 -907
rect -6037 -953 -5991 -907
rect -5913 -953 -5867 -907
rect -5789 -953 -5743 -907
rect -5665 -953 -5619 -907
rect -5541 -953 -5495 -907
rect -5417 -953 -5371 -907
rect -5293 -953 -5247 -907
rect -5169 -953 -5123 -907
rect -5045 -953 -4999 -907
rect -4921 -953 -4875 -907
rect -4797 -953 -4751 -907
rect -4673 -953 -4627 -907
rect -4549 -953 -4503 -907
rect -4425 -953 -4379 -907
rect -4301 -953 -4255 -907
rect -4177 -953 -4131 -907
rect -4053 -953 -4007 -907
rect -3929 -953 -3883 -907
rect -3805 -953 -3759 -907
rect -3681 -953 -3635 -907
rect -3557 -953 -3511 -907
rect -3433 -953 -3387 -907
rect -3309 -953 -3263 -907
rect -3185 -953 -3139 -907
rect -3061 -953 -3015 -907
rect -2937 -953 -2891 -907
rect -2813 -953 -2767 -907
rect -2689 -953 -2643 -907
rect -2565 -953 -2519 -907
rect -2441 -953 -2395 -907
rect -2317 -953 -2271 -907
rect -2193 -953 -2147 -907
rect -2069 -953 -2023 -907
rect -1945 -953 -1899 -907
rect -1821 -953 -1775 -907
rect -1697 -953 -1651 -907
rect -1573 -953 -1527 -907
rect -1449 -953 -1403 -907
rect -1325 -953 -1279 -907
rect -1201 -953 -1155 -907
rect -1077 -953 -1031 -907
rect -953 -953 -907 -907
rect -829 -953 -783 -907
rect -705 -953 -659 -907
rect -581 -953 -535 -907
rect -457 -953 -411 -907
rect -333 -953 -287 -907
rect -209 -953 -163 -907
rect -85 -953 -39 -907
rect 39 -953 85 -907
rect 163 -953 209 -907
rect 287 -953 333 -907
rect 411 -953 457 -907
rect 535 -953 581 -907
rect 659 -953 705 -907
rect 783 -953 829 -907
rect 907 -953 953 -907
rect 1031 -953 1077 -907
rect 1155 -953 1201 -907
rect 1279 -953 1325 -907
rect 1403 -953 1449 -907
rect 1527 -953 1573 -907
rect 1651 -953 1697 -907
rect 1775 -953 1821 -907
rect 1899 -953 1945 -907
rect 2023 -953 2069 -907
rect 2147 -953 2193 -907
rect 2271 -953 2317 -907
rect 2395 -953 2441 -907
rect 2519 -953 2565 -907
rect 2643 -953 2689 -907
rect 2767 -953 2813 -907
rect 2891 -953 2937 -907
rect 3015 -953 3061 -907
rect 3139 -953 3185 -907
rect 3263 -953 3309 -907
rect 3387 -953 3433 -907
rect 3511 -953 3557 -907
rect 3635 -953 3681 -907
rect 3759 -953 3805 -907
rect 3883 -953 3929 -907
rect 4007 -953 4053 -907
rect 4131 -953 4177 -907
rect 4255 -953 4301 -907
rect 4379 -953 4425 -907
rect 4503 -953 4549 -907
rect 4627 -953 4673 -907
rect 4751 -953 4797 -907
rect 4875 -953 4921 -907
rect 4999 -953 5045 -907
rect 5123 -953 5169 -907
rect 5247 -953 5293 -907
rect 5371 -953 5417 -907
rect 5495 -953 5541 -907
rect 5619 -953 5665 -907
rect 5743 -953 5789 -907
rect 5867 -953 5913 -907
rect 5991 -953 6037 -907
rect 6115 -953 6161 -907
rect 6239 -953 6285 -907
rect 6363 -953 6409 -907
rect 6487 -953 6533 -907
rect 6611 -953 6657 -907
rect 6735 -953 6781 -907
rect 6859 -953 6905 -907
rect 6983 -953 7029 -907
rect 7107 -953 7153 -907
rect 7231 -953 7277 -907
rect 7355 -953 7401 -907
rect 7479 -953 7525 -907
rect 7603 -953 7649 -907
rect 7727 -953 7773 -907
rect 7851 -953 7897 -907
rect 7975 -953 8021 -907
rect 8099 -953 8145 -907
rect 8223 -953 8269 -907
rect 8347 -953 8393 -907
rect 8471 -953 8517 -907
rect 8595 -953 8641 -907
rect 8719 -953 8765 -907
rect 8843 -953 8889 -907
rect 8967 -953 9013 -907
rect 9091 -953 9137 -907
rect 9215 -953 9261 -907
rect 9339 -953 9385 -907
rect 9463 -953 9509 -907
rect 9587 -953 9633 -907
rect 9711 -953 9757 -907
rect 9835 -953 9881 -907
rect 9959 -953 10005 -907
rect 10083 -953 10129 -907
rect 10207 -953 10253 -907
rect 10331 -953 10377 -907
rect 10455 -953 10501 -907
rect 10579 -953 10625 -907
rect 10703 -953 10749 -907
rect 10827 -953 10873 -907
rect 10951 -953 10997 -907
rect 11075 -953 11121 -907
rect 11199 -953 11245 -907
rect 11323 -953 11369 -907
rect 11447 -953 11493 -907
rect 11571 -953 11617 -907
rect 11695 -953 11741 -907
rect 11819 -953 11865 -907
rect 11943 -953 11989 -907
rect 12067 -953 12113 -907
rect 12191 -953 12237 -907
rect 12315 -953 12361 -907
rect 12439 -953 12485 -907
rect 12563 -953 12609 -907
rect 12687 -953 12733 -907
rect 12811 -953 12857 -907
rect 12935 -953 12981 -907
rect 13059 -953 13105 -907
rect 13183 -953 13229 -907
rect 13307 -953 13353 -907
rect 13431 -953 13477 -907
rect 13555 -953 13601 -907
rect 13679 -953 13725 -907
rect 13803 -953 13849 -907
rect 13927 -953 13973 -907
rect 14051 -953 14097 -907
rect 14175 -953 14221 -907
rect 14299 -953 14345 -907
rect 14423 -953 14469 -907
rect 14547 -953 14593 -907
rect 14671 -953 14717 -907
rect 14795 -953 14841 -907
rect 14919 -953 14965 -907
rect 15043 -953 15089 -907
rect 15167 -953 15213 -907
rect 15291 -953 15337 -907
rect 15415 -953 15461 -907
rect 15539 -953 15585 -907
rect 15663 -953 15709 -907
rect 15787 -953 15833 -907
rect 15911 -953 15957 -907
rect 16035 -953 16081 -907
rect 16159 -953 16205 -907
rect 16283 -953 16329 -907
rect 16407 -953 16453 -907
rect 16531 -953 16577 -907
rect 16655 -953 16701 -907
rect 16779 -953 16825 -907
rect 16903 -953 16949 -907
rect 17027 -953 17073 -907
rect 17151 -953 17197 -907
rect 17275 -953 17321 -907
<< metal1 >>
rect -17332 953 17332 964
rect -17332 907 -17321 953
rect -17275 907 -17197 953
rect -17151 907 -17073 953
rect -17027 907 -16949 953
rect -16903 907 -16825 953
rect -16779 907 -16701 953
rect -16655 907 -16577 953
rect -16531 907 -16453 953
rect -16407 907 -16329 953
rect -16283 907 -16205 953
rect -16159 907 -16081 953
rect -16035 907 -15957 953
rect -15911 907 -15833 953
rect -15787 907 -15709 953
rect -15663 907 -15585 953
rect -15539 907 -15461 953
rect -15415 907 -15337 953
rect -15291 907 -15213 953
rect -15167 907 -15089 953
rect -15043 907 -14965 953
rect -14919 907 -14841 953
rect -14795 907 -14717 953
rect -14671 907 -14593 953
rect -14547 907 -14469 953
rect -14423 907 -14345 953
rect -14299 907 -14221 953
rect -14175 907 -14097 953
rect -14051 907 -13973 953
rect -13927 907 -13849 953
rect -13803 907 -13725 953
rect -13679 907 -13601 953
rect -13555 907 -13477 953
rect -13431 907 -13353 953
rect -13307 907 -13229 953
rect -13183 907 -13105 953
rect -13059 907 -12981 953
rect -12935 907 -12857 953
rect -12811 907 -12733 953
rect -12687 907 -12609 953
rect -12563 907 -12485 953
rect -12439 907 -12361 953
rect -12315 907 -12237 953
rect -12191 907 -12113 953
rect -12067 907 -11989 953
rect -11943 907 -11865 953
rect -11819 907 -11741 953
rect -11695 907 -11617 953
rect -11571 907 -11493 953
rect -11447 907 -11369 953
rect -11323 907 -11245 953
rect -11199 907 -11121 953
rect -11075 907 -10997 953
rect -10951 907 -10873 953
rect -10827 907 -10749 953
rect -10703 907 -10625 953
rect -10579 907 -10501 953
rect -10455 907 -10377 953
rect -10331 907 -10253 953
rect -10207 907 -10129 953
rect -10083 907 -10005 953
rect -9959 907 -9881 953
rect -9835 907 -9757 953
rect -9711 907 -9633 953
rect -9587 907 -9509 953
rect -9463 907 -9385 953
rect -9339 907 -9261 953
rect -9215 907 -9137 953
rect -9091 907 -9013 953
rect -8967 907 -8889 953
rect -8843 907 -8765 953
rect -8719 907 -8641 953
rect -8595 907 -8517 953
rect -8471 907 -8393 953
rect -8347 907 -8269 953
rect -8223 907 -8145 953
rect -8099 907 -8021 953
rect -7975 907 -7897 953
rect -7851 907 -7773 953
rect -7727 907 -7649 953
rect -7603 907 -7525 953
rect -7479 907 -7401 953
rect -7355 907 -7277 953
rect -7231 907 -7153 953
rect -7107 907 -7029 953
rect -6983 907 -6905 953
rect -6859 907 -6781 953
rect -6735 907 -6657 953
rect -6611 907 -6533 953
rect -6487 907 -6409 953
rect -6363 907 -6285 953
rect -6239 907 -6161 953
rect -6115 907 -6037 953
rect -5991 907 -5913 953
rect -5867 907 -5789 953
rect -5743 907 -5665 953
rect -5619 907 -5541 953
rect -5495 907 -5417 953
rect -5371 907 -5293 953
rect -5247 907 -5169 953
rect -5123 907 -5045 953
rect -4999 907 -4921 953
rect -4875 907 -4797 953
rect -4751 907 -4673 953
rect -4627 907 -4549 953
rect -4503 907 -4425 953
rect -4379 907 -4301 953
rect -4255 907 -4177 953
rect -4131 907 -4053 953
rect -4007 907 -3929 953
rect -3883 907 -3805 953
rect -3759 907 -3681 953
rect -3635 907 -3557 953
rect -3511 907 -3433 953
rect -3387 907 -3309 953
rect -3263 907 -3185 953
rect -3139 907 -3061 953
rect -3015 907 -2937 953
rect -2891 907 -2813 953
rect -2767 907 -2689 953
rect -2643 907 -2565 953
rect -2519 907 -2441 953
rect -2395 907 -2317 953
rect -2271 907 -2193 953
rect -2147 907 -2069 953
rect -2023 907 -1945 953
rect -1899 907 -1821 953
rect -1775 907 -1697 953
rect -1651 907 -1573 953
rect -1527 907 -1449 953
rect -1403 907 -1325 953
rect -1279 907 -1201 953
rect -1155 907 -1077 953
rect -1031 907 -953 953
rect -907 907 -829 953
rect -783 907 -705 953
rect -659 907 -581 953
rect -535 907 -457 953
rect -411 907 -333 953
rect -287 907 -209 953
rect -163 907 -85 953
rect -39 907 39 953
rect 85 907 163 953
rect 209 907 287 953
rect 333 907 411 953
rect 457 907 535 953
rect 581 907 659 953
rect 705 907 783 953
rect 829 907 907 953
rect 953 907 1031 953
rect 1077 907 1155 953
rect 1201 907 1279 953
rect 1325 907 1403 953
rect 1449 907 1527 953
rect 1573 907 1651 953
rect 1697 907 1775 953
rect 1821 907 1899 953
rect 1945 907 2023 953
rect 2069 907 2147 953
rect 2193 907 2271 953
rect 2317 907 2395 953
rect 2441 907 2519 953
rect 2565 907 2643 953
rect 2689 907 2767 953
rect 2813 907 2891 953
rect 2937 907 3015 953
rect 3061 907 3139 953
rect 3185 907 3263 953
rect 3309 907 3387 953
rect 3433 907 3511 953
rect 3557 907 3635 953
rect 3681 907 3759 953
rect 3805 907 3883 953
rect 3929 907 4007 953
rect 4053 907 4131 953
rect 4177 907 4255 953
rect 4301 907 4379 953
rect 4425 907 4503 953
rect 4549 907 4627 953
rect 4673 907 4751 953
rect 4797 907 4875 953
rect 4921 907 4999 953
rect 5045 907 5123 953
rect 5169 907 5247 953
rect 5293 907 5371 953
rect 5417 907 5495 953
rect 5541 907 5619 953
rect 5665 907 5743 953
rect 5789 907 5867 953
rect 5913 907 5991 953
rect 6037 907 6115 953
rect 6161 907 6239 953
rect 6285 907 6363 953
rect 6409 907 6487 953
rect 6533 907 6611 953
rect 6657 907 6735 953
rect 6781 907 6859 953
rect 6905 907 6983 953
rect 7029 907 7107 953
rect 7153 907 7231 953
rect 7277 907 7355 953
rect 7401 907 7479 953
rect 7525 907 7603 953
rect 7649 907 7727 953
rect 7773 907 7851 953
rect 7897 907 7975 953
rect 8021 907 8099 953
rect 8145 907 8223 953
rect 8269 907 8347 953
rect 8393 907 8471 953
rect 8517 907 8595 953
rect 8641 907 8719 953
rect 8765 907 8843 953
rect 8889 907 8967 953
rect 9013 907 9091 953
rect 9137 907 9215 953
rect 9261 907 9339 953
rect 9385 907 9463 953
rect 9509 907 9587 953
rect 9633 907 9711 953
rect 9757 907 9835 953
rect 9881 907 9959 953
rect 10005 907 10083 953
rect 10129 907 10207 953
rect 10253 907 10331 953
rect 10377 907 10455 953
rect 10501 907 10579 953
rect 10625 907 10703 953
rect 10749 907 10827 953
rect 10873 907 10951 953
rect 10997 907 11075 953
rect 11121 907 11199 953
rect 11245 907 11323 953
rect 11369 907 11447 953
rect 11493 907 11571 953
rect 11617 907 11695 953
rect 11741 907 11819 953
rect 11865 907 11943 953
rect 11989 907 12067 953
rect 12113 907 12191 953
rect 12237 907 12315 953
rect 12361 907 12439 953
rect 12485 907 12563 953
rect 12609 907 12687 953
rect 12733 907 12811 953
rect 12857 907 12935 953
rect 12981 907 13059 953
rect 13105 907 13183 953
rect 13229 907 13307 953
rect 13353 907 13431 953
rect 13477 907 13555 953
rect 13601 907 13679 953
rect 13725 907 13803 953
rect 13849 907 13927 953
rect 13973 907 14051 953
rect 14097 907 14175 953
rect 14221 907 14299 953
rect 14345 907 14423 953
rect 14469 907 14547 953
rect 14593 907 14671 953
rect 14717 907 14795 953
rect 14841 907 14919 953
rect 14965 907 15043 953
rect 15089 907 15167 953
rect 15213 907 15291 953
rect 15337 907 15415 953
rect 15461 907 15539 953
rect 15585 907 15663 953
rect 15709 907 15787 953
rect 15833 907 15911 953
rect 15957 907 16035 953
rect 16081 907 16159 953
rect 16205 907 16283 953
rect 16329 907 16407 953
rect 16453 907 16531 953
rect 16577 907 16655 953
rect 16701 907 16779 953
rect 16825 907 16903 953
rect 16949 907 17027 953
rect 17073 907 17151 953
rect 17197 907 17275 953
rect 17321 907 17332 953
rect -17332 829 17332 907
rect -17332 783 -17321 829
rect -17275 783 -17197 829
rect -17151 783 -17073 829
rect -17027 783 -16949 829
rect -16903 783 -16825 829
rect -16779 783 -16701 829
rect -16655 783 -16577 829
rect -16531 783 -16453 829
rect -16407 783 -16329 829
rect -16283 783 -16205 829
rect -16159 783 -16081 829
rect -16035 783 -15957 829
rect -15911 783 -15833 829
rect -15787 783 -15709 829
rect -15663 783 -15585 829
rect -15539 783 -15461 829
rect -15415 783 -15337 829
rect -15291 783 -15213 829
rect -15167 783 -15089 829
rect -15043 783 -14965 829
rect -14919 783 -14841 829
rect -14795 783 -14717 829
rect -14671 783 -14593 829
rect -14547 783 -14469 829
rect -14423 783 -14345 829
rect -14299 783 -14221 829
rect -14175 783 -14097 829
rect -14051 783 -13973 829
rect -13927 783 -13849 829
rect -13803 783 -13725 829
rect -13679 783 -13601 829
rect -13555 783 -13477 829
rect -13431 783 -13353 829
rect -13307 783 -13229 829
rect -13183 783 -13105 829
rect -13059 783 -12981 829
rect -12935 783 -12857 829
rect -12811 783 -12733 829
rect -12687 783 -12609 829
rect -12563 783 -12485 829
rect -12439 783 -12361 829
rect -12315 783 -12237 829
rect -12191 783 -12113 829
rect -12067 783 -11989 829
rect -11943 783 -11865 829
rect -11819 783 -11741 829
rect -11695 783 -11617 829
rect -11571 783 -11493 829
rect -11447 783 -11369 829
rect -11323 783 -11245 829
rect -11199 783 -11121 829
rect -11075 783 -10997 829
rect -10951 783 -10873 829
rect -10827 783 -10749 829
rect -10703 783 -10625 829
rect -10579 783 -10501 829
rect -10455 783 -10377 829
rect -10331 783 -10253 829
rect -10207 783 -10129 829
rect -10083 783 -10005 829
rect -9959 783 -9881 829
rect -9835 783 -9757 829
rect -9711 783 -9633 829
rect -9587 783 -9509 829
rect -9463 783 -9385 829
rect -9339 783 -9261 829
rect -9215 783 -9137 829
rect -9091 783 -9013 829
rect -8967 783 -8889 829
rect -8843 783 -8765 829
rect -8719 783 -8641 829
rect -8595 783 -8517 829
rect -8471 783 -8393 829
rect -8347 783 -8269 829
rect -8223 783 -8145 829
rect -8099 783 -8021 829
rect -7975 783 -7897 829
rect -7851 783 -7773 829
rect -7727 783 -7649 829
rect -7603 783 -7525 829
rect -7479 783 -7401 829
rect -7355 783 -7277 829
rect -7231 783 -7153 829
rect -7107 783 -7029 829
rect -6983 783 -6905 829
rect -6859 783 -6781 829
rect -6735 783 -6657 829
rect -6611 783 -6533 829
rect -6487 783 -6409 829
rect -6363 783 -6285 829
rect -6239 783 -6161 829
rect -6115 783 -6037 829
rect -5991 783 -5913 829
rect -5867 783 -5789 829
rect -5743 783 -5665 829
rect -5619 783 -5541 829
rect -5495 783 -5417 829
rect -5371 783 -5293 829
rect -5247 783 -5169 829
rect -5123 783 -5045 829
rect -4999 783 -4921 829
rect -4875 783 -4797 829
rect -4751 783 -4673 829
rect -4627 783 -4549 829
rect -4503 783 -4425 829
rect -4379 783 -4301 829
rect -4255 783 -4177 829
rect -4131 783 -4053 829
rect -4007 783 -3929 829
rect -3883 783 -3805 829
rect -3759 783 -3681 829
rect -3635 783 -3557 829
rect -3511 783 -3433 829
rect -3387 783 -3309 829
rect -3263 783 -3185 829
rect -3139 783 -3061 829
rect -3015 783 -2937 829
rect -2891 783 -2813 829
rect -2767 783 -2689 829
rect -2643 783 -2565 829
rect -2519 783 -2441 829
rect -2395 783 -2317 829
rect -2271 783 -2193 829
rect -2147 783 -2069 829
rect -2023 783 -1945 829
rect -1899 783 -1821 829
rect -1775 783 -1697 829
rect -1651 783 -1573 829
rect -1527 783 -1449 829
rect -1403 783 -1325 829
rect -1279 783 -1201 829
rect -1155 783 -1077 829
rect -1031 783 -953 829
rect -907 783 -829 829
rect -783 783 -705 829
rect -659 783 -581 829
rect -535 783 -457 829
rect -411 783 -333 829
rect -287 783 -209 829
rect -163 783 -85 829
rect -39 783 39 829
rect 85 783 163 829
rect 209 783 287 829
rect 333 783 411 829
rect 457 783 535 829
rect 581 783 659 829
rect 705 783 783 829
rect 829 783 907 829
rect 953 783 1031 829
rect 1077 783 1155 829
rect 1201 783 1279 829
rect 1325 783 1403 829
rect 1449 783 1527 829
rect 1573 783 1651 829
rect 1697 783 1775 829
rect 1821 783 1899 829
rect 1945 783 2023 829
rect 2069 783 2147 829
rect 2193 783 2271 829
rect 2317 783 2395 829
rect 2441 783 2519 829
rect 2565 783 2643 829
rect 2689 783 2767 829
rect 2813 783 2891 829
rect 2937 783 3015 829
rect 3061 783 3139 829
rect 3185 783 3263 829
rect 3309 783 3387 829
rect 3433 783 3511 829
rect 3557 783 3635 829
rect 3681 783 3759 829
rect 3805 783 3883 829
rect 3929 783 4007 829
rect 4053 783 4131 829
rect 4177 783 4255 829
rect 4301 783 4379 829
rect 4425 783 4503 829
rect 4549 783 4627 829
rect 4673 783 4751 829
rect 4797 783 4875 829
rect 4921 783 4999 829
rect 5045 783 5123 829
rect 5169 783 5247 829
rect 5293 783 5371 829
rect 5417 783 5495 829
rect 5541 783 5619 829
rect 5665 783 5743 829
rect 5789 783 5867 829
rect 5913 783 5991 829
rect 6037 783 6115 829
rect 6161 783 6239 829
rect 6285 783 6363 829
rect 6409 783 6487 829
rect 6533 783 6611 829
rect 6657 783 6735 829
rect 6781 783 6859 829
rect 6905 783 6983 829
rect 7029 783 7107 829
rect 7153 783 7231 829
rect 7277 783 7355 829
rect 7401 783 7479 829
rect 7525 783 7603 829
rect 7649 783 7727 829
rect 7773 783 7851 829
rect 7897 783 7975 829
rect 8021 783 8099 829
rect 8145 783 8223 829
rect 8269 783 8347 829
rect 8393 783 8471 829
rect 8517 783 8595 829
rect 8641 783 8719 829
rect 8765 783 8843 829
rect 8889 783 8967 829
rect 9013 783 9091 829
rect 9137 783 9215 829
rect 9261 783 9339 829
rect 9385 783 9463 829
rect 9509 783 9587 829
rect 9633 783 9711 829
rect 9757 783 9835 829
rect 9881 783 9959 829
rect 10005 783 10083 829
rect 10129 783 10207 829
rect 10253 783 10331 829
rect 10377 783 10455 829
rect 10501 783 10579 829
rect 10625 783 10703 829
rect 10749 783 10827 829
rect 10873 783 10951 829
rect 10997 783 11075 829
rect 11121 783 11199 829
rect 11245 783 11323 829
rect 11369 783 11447 829
rect 11493 783 11571 829
rect 11617 783 11695 829
rect 11741 783 11819 829
rect 11865 783 11943 829
rect 11989 783 12067 829
rect 12113 783 12191 829
rect 12237 783 12315 829
rect 12361 783 12439 829
rect 12485 783 12563 829
rect 12609 783 12687 829
rect 12733 783 12811 829
rect 12857 783 12935 829
rect 12981 783 13059 829
rect 13105 783 13183 829
rect 13229 783 13307 829
rect 13353 783 13431 829
rect 13477 783 13555 829
rect 13601 783 13679 829
rect 13725 783 13803 829
rect 13849 783 13927 829
rect 13973 783 14051 829
rect 14097 783 14175 829
rect 14221 783 14299 829
rect 14345 783 14423 829
rect 14469 783 14547 829
rect 14593 783 14671 829
rect 14717 783 14795 829
rect 14841 783 14919 829
rect 14965 783 15043 829
rect 15089 783 15167 829
rect 15213 783 15291 829
rect 15337 783 15415 829
rect 15461 783 15539 829
rect 15585 783 15663 829
rect 15709 783 15787 829
rect 15833 783 15911 829
rect 15957 783 16035 829
rect 16081 783 16159 829
rect 16205 783 16283 829
rect 16329 783 16407 829
rect 16453 783 16531 829
rect 16577 783 16655 829
rect 16701 783 16779 829
rect 16825 783 16903 829
rect 16949 783 17027 829
rect 17073 783 17151 829
rect 17197 783 17275 829
rect 17321 783 17332 829
rect -17332 705 17332 783
rect -17332 659 -17321 705
rect -17275 659 -17197 705
rect -17151 659 -17073 705
rect -17027 659 -16949 705
rect -16903 659 -16825 705
rect -16779 659 -16701 705
rect -16655 659 -16577 705
rect -16531 659 -16453 705
rect -16407 659 -16329 705
rect -16283 659 -16205 705
rect -16159 659 -16081 705
rect -16035 659 -15957 705
rect -15911 659 -15833 705
rect -15787 659 -15709 705
rect -15663 659 -15585 705
rect -15539 659 -15461 705
rect -15415 659 -15337 705
rect -15291 659 -15213 705
rect -15167 659 -15089 705
rect -15043 659 -14965 705
rect -14919 659 -14841 705
rect -14795 659 -14717 705
rect -14671 659 -14593 705
rect -14547 659 -14469 705
rect -14423 659 -14345 705
rect -14299 659 -14221 705
rect -14175 659 -14097 705
rect -14051 659 -13973 705
rect -13927 659 -13849 705
rect -13803 659 -13725 705
rect -13679 659 -13601 705
rect -13555 659 -13477 705
rect -13431 659 -13353 705
rect -13307 659 -13229 705
rect -13183 659 -13105 705
rect -13059 659 -12981 705
rect -12935 659 -12857 705
rect -12811 659 -12733 705
rect -12687 659 -12609 705
rect -12563 659 -12485 705
rect -12439 659 -12361 705
rect -12315 659 -12237 705
rect -12191 659 -12113 705
rect -12067 659 -11989 705
rect -11943 659 -11865 705
rect -11819 659 -11741 705
rect -11695 659 -11617 705
rect -11571 659 -11493 705
rect -11447 659 -11369 705
rect -11323 659 -11245 705
rect -11199 659 -11121 705
rect -11075 659 -10997 705
rect -10951 659 -10873 705
rect -10827 659 -10749 705
rect -10703 659 -10625 705
rect -10579 659 -10501 705
rect -10455 659 -10377 705
rect -10331 659 -10253 705
rect -10207 659 -10129 705
rect -10083 659 -10005 705
rect -9959 659 -9881 705
rect -9835 659 -9757 705
rect -9711 659 -9633 705
rect -9587 659 -9509 705
rect -9463 659 -9385 705
rect -9339 659 -9261 705
rect -9215 659 -9137 705
rect -9091 659 -9013 705
rect -8967 659 -8889 705
rect -8843 659 -8765 705
rect -8719 659 -8641 705
rect -8595 659 -8517 705
rect -8471 659 -8393 705
rect -8347 659 -8269 705
rect -8223 659 -8145 705
rect -8099 659 -8021 705
rect -7975 659 -7897 705
rect -7851 659 -7773 705
rect -7727 659 -7649 705
rect -7603 659 -7525 705
rect -7479 659 -7401 705
rect -7355 659 -7277 705
rect -7231 659 -7153 705
rect -7107 659 -7029 705
rect -6983 659 -6905 705
rect -6859 659 -6781 705
rect -6735 659 -6657 705
rect -6611 659 -6533 705
rect -6487 659 -6409 705
rect -6363 659 -6285 705
rect -6239 659 -6161 705
rect -6115 659 -6037 705
rect -5991 659 -5913 705
rect -5867 659 -5789 705
rect -5743 659 -5665 705
rect -5619 659 -5541 705
rect -5495 659 -5417 705
rect -5371 659 -5293 705
rect -5247 659 -5169 705
rect -5123 659 -5045 705
rect -4999 659 -4921 705
rect -4875 659 -4797 705
rect -4751 659 -4673 705
rect -4627 659 -4549 705
rect -4503 659 -4425 705
rect -4379 659 -4301 705
rect -4255 659 -4177 705
rect -4131 659 -4053 705
rect -4007 659 -3929 705
rect -3883 659 -3805 705
rect -3759 659 -3681 705
rect -3635 659 -3557 705
rect -3511 659 -3433 705
rect -3387 659 -3309 705
rect -3263 659 -3185 705
rect -3139 659 -3061 705
rect -3015 659 -2937 705
rect -2891 659 -2813 705
rect -2767 659 -2689 705
rect -2643 659 -2565 705
rect -2519 659 -2441 705
rect -2395 659 -2317 705
rect -2271 659 -2193 705
rect -2147 659 -2069 705
rect -2023 659 -1945 705
rect -1899 659 -1821 705
rect -1775 659 -1697 705
rect -1651 659 -1573 705
rect -1527 659 -1449 705
rect -1403 659 -1325 705
rect -1279 659 -1201 705
rect -1155 659 -1077 705
rect -1031 659 -953 705
rect -907 659 -829 705
rect -783 659 -705 705
rect -659 659 -581 705
rect -535 659 -457 705
rect -411 659 -333 705
rect -287 659 -209 705
rect -163 659 -85 705
rect -39 659 39 705
rect 85 659 163 705
rect 209 659 287 705
rect 333 659 411 705
rect 457 659 535 705
rect 581 659 659 705
rect 705 659 783 705
rect 829 659 907 705
rect 953 659 1031 705
rect 1077 659 1155 705
rect 1201 659 1279 705
rect 1325 659 1403 705
rect 1449 659 1527 705
rect 1573 659 1651 705
rect 1697 659 1775 705
rect 1821 659 1899 705
rect 1945 659 2023 705
rect 2069 659 2147 705
rect 2193 659 2271 705
rect 2317 659 2395 705
rect 2441 659 2519 705
rect 2565 659 2643 705
rect 2689 659 2767 705
rect 2813 659 2891 705
rect 2937 659 3015 705
rect 3061 659 3139 705
rect 3185 659 3263 705
rect 3309 659 3387 705
rect 3433 659 3511 705
rect 3557 659 3635 705
rect 3681 659 3759 705
rect 3805 659 3883 705
rect 3929 659 4007 705
rect 4053 659 4131 705
rect 4177 659 4255 705
rect 4301 659 4379 705
rect 4425 659 4503 705
rect 4549 659 4627 705
rect 4673 659 4751 705
rect 4797 659 4875 705
rect 4921 659 4999 705
rect 5045 659 5123 705
rect 5169 659 5247 705
rect 5293 659 5371 705
rect 5417 659 5495 705
rect 5541 659 5619 705
rect 5665 659 5743 705
rect 5789 659 5867 705
rect 5913 659 5991 705
rect 6037 659 6115 705
rect 6161 659 6239 705
rect 6285 659 6363 705
rect 6409 659 6487 705
rect 6533 659 6611 705
rect 6657 659 6735 705
rect 6781 659 6859 705
rect 6905 659 6983 705
rect 7029 659 7107 705
rect 7153 659 7231 705
rect 7277 659 7355 705
rect 7401 659 7479 705
rect 7525 659 7603 705
rect 7649 659 7727 705
rect 7773 659 7851 705
rect 7897 659 7975 705
rect 8021 659 8099 705
rect 8145 659 8223 705
rect 8269 659 8347 705
rect 8393 659 8471 705
rect 8517 659 8595 705
rect 8641 659 8719 705
rect 8765 659 8843 705
rect 8889 659 8967 705
rect 9013 659 9091 705
rect 9137 659 9215 705
rect 9261 659 9339 705
rect 9385 659 9463 705
rect 9509 659 9587 705
rect 9633 659 9711 705
rect 9757 659 9835 705
rect 9881 659 9959 705
rect 10005 659 10083 705
rect 10129 659 10207 705
rect 10253 659 10331 705
rect 10377 659 10455 705
rect 10501 659 10579 705
rect 10625 659 10703 705
rect 10749 659 10827 705
rect 10873 659 10951 705
rect 10997 659 11075 705
rect 11121 659 11199 705
rect 11245 659 11323 705
rect 11369 659 11447 705
rect 11493 659 11571 705
rect 11617 659 11695 705
rect 11741 659 11819 705
rect 11865 659 11943 705
rect 11989 659 12067 705
rect 12113 659 12191 705
rect 12237 659 12315 705
rect 12361 659 12439 705
rect 12485 659 12563 705
rect 12609 659 12687 705
rect 12733 659 12811 705
rect 12857 659 12935 705
rect 12981 659 13059 705
rect 13105 659 13183 705
rect 13229 659 13307 705
rect 13353 659 13431 705
rect 13477 659 13555 705
rect 13601 659 13679 705
rect 13725 659 13803 705
rect 13849 659 13927 705
rect 13973 659 14051 705
rect 14097 659 14175 705
rect 14221 659 14299 705
rect 14345 659 14423 705
rect 14469 659 14547 705
rect 14593 659 14671 705
rect 14717 659 14795 705
rect 14841 659 14919 705
rect 14965 659 15043 705
rect 15089 659 15167 705
rect 15213 659 15291 705
rect 15337 659 15415 705
rect 15461 659 15539 705
rect 15585 659 15663 705
rect 15709 659 15787 705
rect 15833 659 15911 705
rect 15957 659 16035 705
rect 16081 659 16159 705
rect 16205 659 16283 705
rect 16329 659 16407 705
rect 16453 659 16531 705
rect 16577 659 16655 705
rect 16701 659 16779 705
rect 16825 659 16903 705
rect 16949 659 17027 705
rect 17073 659 17151 705
rect 17197 659 17275 705
rect 17321 659 17332 705
rect -17332 581 17332 659
rect -17332 535 -17321 581
rect -17275 535 -17197 581
rect -17151 535 -17073 581
rect -17027 535 -16949 581
rect -16903 535 -16825 581
rect -16779 535 -16701 581
rect -16655 535 -16577 581
rect -16531 535 -16453 581
rect -16407 535 -16329 581
rect -16283 535 -16205 581
rect -16159 535 -16081 581
rect -16035 535 -15957 581
rect -15911 535 -15833 581
rect -15787 535 -15709 581
rect -15663 535 -15585 581
rect -15539 535 -15461 581
rect -15415 535 -15337 581
rect -15291 535 -15213 581
rect -15167 535 -15089 581
rect -15043 535 -14965 581
rect -14919 535 -14841 581
rect -14795 535 -14717 581
rect -14671 535 -14593 581
rect -14547 535 -14469 581
rect -14423 535 -14345 581
rect -14299 535 -14221 581
rect -14175 535 -14097 581
rect -14051 535 -13973 581
rect -13927 535 -13849 581
rect -13803 535 -13725 581
rect -13679 535 -13601 581
rect -13555 535 -13477 581
rect -13431 535 -13353 581
rect -13307 535 -13229 581
rect -13183 535 -13105 581
rect -13059 535 -12981 581
rect -12935 535 -12857 581
rect -12811 535 -12733 581
rect -12687 535 -12609 581
rect -12563 535 -12485 581
rect -12439 535 -12361 581
rect -12315 535 -12237 581
rect -12191 535 -12113 581
rect -12067 535 -11989 581
rect -11943 535 -11865 581
rect -11819 535 -11741 581
rect -11695 535 -11617 581
rect -11571 535 -11493 581
rect -11447 535 -11369 581
rect -11323 535 -11245 581
rect -11199 535 -11121 581
rect -11075 535 -10997 581
rect -10951 535 -10873 581
rect -10827 535 -10749 581
rect -10703 535 -10625 581
rect -10579 535 -10501 581
rect -10455 535 -10377 581
rect -10331 535 -10253 581
rect -10207 535 -10129 581
rect -10083 535 -10005 581
rect -9959 535 -9881 581
rect -9835 535 -9757 581
rect -9711 535 -9633 581
rect -9587 535 -9509 581
rect -9463 535 -9385 581
rect -9339 535 -9261 581
rect -9215 535 -9137 581
rect -9091 535 -9013 581
rect -8967 535 -8889 581
rect -8843 535 -8765 581
rect -8719 535 -8641 581
rect -8595 535 -8517 581
rect -8471 535 -8393 581
rect -8347 535 -8269 581
rect -8223 535 -8145 581
rect -8099 535 -8021 581
rect -7975 535 -7897 581
rect -7851 535 -7773 581
rect -7727 535 -7649 581
rect -7603 535 -7525 581
rect -7479 535 -7401 581
rect -7355 535 -7277 581
rect -7231 535 -7153 581
rect -7107 535 -7029 581
rect -6983 535 -6905 581
rect -6859 535 -6781 581
rect -6735 535 -6657 581
rect -6611 535 -6533 581
rect -6487 535 -6409 581
rect -6363 535 -6285 581
rect -6239 535 -6161 581
rect -6115 535 -6037 581
rect -5991 535 -5913 581
rect -5867 535 -5789 581
rect -5743 535 -5665 581
rect -5619 535 -5541 581
rect -5495 535 -5417 581
rect -5371 535 -5293 581
rect -5247 535 -5169 581
rect -5123 535 -5045 581
rect -4999 535 -4921 581
rect -4875 535 -4797 581
rect -4751 535 -4673 581
rect -4627 535 -4549 581
rect -4503 535 -4425 581
rect -4379 535 -4301 581
rect -4255 535 -4177 581
rect -4131 535 -4053 581
rect -4007 535 -3929 581
rect -3883 535 -3805 581
rect -3759 535 -3681 581
rect -3635 535 -3557 581
rect -3511 535 -3433 581
rect -3387 535 -3309 581
rect -3263 535 -3185 581
rect -3139 535 -3061 581
rect -3015 535 -2937 581
rect -2891 535 -2813 581
rect -2767 535 -2689 581
rect -2643 535 -2565 581
rect -2519 535 -2441 581
rect -2395 535 -2317 581
rect -2271 535 -2193 581
rect -2147 535 -2069 581
rect -2023 535 -1945 581
rect -1899 535 -1821 581
rect -1775 535 -1697 581
rect -1651 535 -1573 581
rect -1527 535 -1449 581
rect -1403 535 -1325 581
rect -1279 535 -1201 581
rect -1155 535 -1077 581
rect -1031 535 -953 581
rect -907 535 -829 581
rect -783 535 -705 581
rect -659 535 -581 581
rect -535 535 -457 581
rect -411 535 -333 581
rect -287 535 -209 581
rect -163 535 -85 581
rect -39 535 39 581
rect 85 535 163 581
rect 209 535 287 581
rect 333 535 411 581
rect 457 535 535 581
rect 581 535 659 581
rect 705 535 783 581
rect 829 535 907 581
rect 953 535 1031 581
rect 1077 535 1155 581
rect 1201 535 1279 581
rect 1325 535 1403 581
rect 1449 535 1527 581
rect 1573 535 1651 581
rect 1697 535 1775 581
rect 1821 535 1899 581
rect 1945 535 2023 581
rect 2069 535 2147 581
rect 2193 535 2271 581
rect 2317 535 2395 581
rect 2441 535 2519 581
rect 2565 535 2643 581
rect 2689 535 2767 581
rect 2813 535 2891 581
rect 2937 535 3015 581
rect 3061 535 3139 581
rect 3185 535 3263 581
rect 3309 535 3387 581
rect 3433 535 3511 581
rect 3557 535 3635 581
rect 3681 535 3759 581
rect 3805 535 3883 581
rect 3929 535 4007 581
rect 4053 535 4131 581
rect 4177 535 4255 581
rect 4301 535 4379 581
rect 4425 535 4503 581
rect 4549 535 4627 581
rect 4673 535 4751 581
rect 4797 535 4875 581
rect 4921 535 4999 581
rect 5045 535 5123 581
rect 5169 535 5247 581
rect 5293 535 5371 581
rect 5417 535 5495 581
rect 5541 535 5619 581
rect 5665 535 5743 581
rect 5789 535 5867 581
rect 5913 535 5991 581
rect 6037 535 6115 581
rect 6161 535 6239 581
rect 6285 535 6363 581
rect 6409 535 6487 581
rect 6533 535 6611 581
rect 6657 535 6735 581
rect 6781 535 6859 581
rect 6905 535 6983 581
rect 7029 535 7107 581
rect 7153 535 7231 581
rect 7277 535 7355 581
rect 7401 535 7479 581
rect 7525 535 7603 581
rect 7649 535 7727 581
rect 7773 535 7851 581
rect 7897 535 7975 581
rect 8021 535 8099 581
rect 8145 535 8223 581
rect 8269 535 8347 581
rect 8393 535 8471 581
rect 8517 535 8595 581
rect 8641 535 8719 581
rect 8765 535 8843 581
rect 8889 535 8967 581
rect 9013 535 9091 581
rect 9137 535 9215 581
rect 9261 535 9339 581
rect 9385 535 9463 581
rect 9509 535 9587 581
rect 9633 535 9711 581
rect 9757 535 9835 581
rect 9881 535 9959 581
rect 10005 535 10083 581
rect 10129 535 10207 581
rect 10253 535 10331 581
rect 10377 535 10455 581
rect 10501 535 10579 581
rect 10625 535 10703 581
rect 10749 535 10827 581
rect 10873 535 10951 581
rect 10997 535 11075 581
rect 11121 535 11199 581
rect 11245 535 11323 581
rect 11369 535 11447 581
rect 11493 535 11571 581
rect 11617 535 11695 581
rect 11741 535 11819 581
rect 11865 535 11943 581
rect 11989 535 12067 581
rect 12113 535 12191 581
rect 12237 535 12315 581
rect 12361 535 12439 581
rect 12485 535 12563 581
rect 12609 535 12687 581
rect 12733 535 12811 581
rect 12857 535 12935 581
rect 12981 535 13059 581
rect 13105 535 13183 581
rect 13229 535 13307 581
rect 13353 535 13431 581
rect 13477 535 13555 581
rect 13601 535 13679 581
rect 13725 535 13803 581
rect 13849 535 13927 581
rect 13973 535 14051 581
rect 14097 535 14175 581
rect 14221 535 14299 581
rect 14345 535 14423 581
rect 14469 535 14547 581
rect 14593 535 14671 581
rect 14717 535 14795 581
rect 14841 535 14919 581
rect 14965 535 15043 581
rect 15089 535 15167 581
rect 15213 535 15291 581
rect 15337 535 15415 581
rect 15461 535 15539 581
rect 15585 535 15663 581
rect 15709 535 15787 581
rect 15833 535 15911 581
rect 15957 535 16035 581
rect 16081 535 16159 581
rect 16205 535 16283 581
rect 16329 535 16407 581
rect 16453 535 16531 581
rect 16577 535 16655 581
rect 16701 535 16779 581
rect 16825 535 16903 581
rect 16949 535 17027 581
rect 17073 535 17151 581
rect 17197 535 17275 581
rect 17321 535 17332 581
rect -17332 457 17332 535
rect -17332 411 -17321 457
rect -17275 411 -17197 457
rect -17151 411 -17073 457
rect -17027 411 -16949 457
rect -16903 411 -16825 457
rect -16779 411 -16701 457
rect -16655 411 -16577 457
rect -16531 411 -16453 457
rect -16407 411 -16329 457
rect -16283 411 -16205 457
rect -16159 411 -16081 457
rect -16035 411 -15957 457
rect -15911 411 -15833 457
rect -15787 411 -15709 457
rect -15663 411 -15585 457
rect -15539 411 -15461 457
rect -15415 411 -15337 457
rect -15291 411 -15213 457
rect -15167 411 -15089 457
rect -15043 411 -14965 457
rect -14919 411 -14841 457
rect -14795 411 -14717 457
rect -14671 411 -14593 457
rect -14547 411 -14469 457
rect -14423 411 -14345 457
rect -14299 411 -14221 457
rect -14175 411 -14097 457
rect -14051 411 -13973 457
rect -13927 411 -13849 457
rect -13803 411 -13725 457
rect -13679 411 -13601 457
rect -13555 411 -13477 457
rect -13431 411 -13353 457
rect -13307 411 -13229 457
rect -13183 411 -13105 457
rect -13059 411 -12981 457
rect -12935 411 -12857 457
rect -12811 411 -12733 457
rect -12687 411 -12609 457
rect -12563 411 -12485 457
rect -12439 411 -12361 457
rect -12315 411 -12237 457
rect -12191 411 -12113 457
rect -12067 411 -11989 457
rect -11943 411 -11865 457
rect -11819 411 -11741 457
rect -11695 411 -11617 457
rect -11571 411 -11493 457
rect -11447 411 -11369 457
rect -11323 411 -11245 457
rect -11199 411 -11121 457
rect -11075 411 -10997 457
rect -10951 411 -10873 457
rect -10827 411 -10749 457
rect -10703 411 -10625 457
rect -10579 411 -10501 457
rect -10455 411 -10377 457
rect -10331 411 -10253 457
rect -10207 411 -10129 457
rect -10083 411 -10005 457
rect -9959 411 -9881 457
rect -9835 411 -9757 457
rect -9711 411 -9633 457
rect -9587 411 -9509 457
rect -9463 411 -9385 457
rect -9339 411 -9261 457
rect -9215 411 -9137 457
rect -9091 411 -9013 457
rect -8967 411 -8889 457
rect -8843 411 -8765 457
rect -8719 411 -8641 457
rect -8595 411 -8517 457
rect -8471 411 -8393 457
rect -8347 411 -8269 457
rect -8223 411 -8145 457
rect -8099 411 -8021 457
rect -7975 411 -7897 457
rect -7851 411 -7773 457
rect -7727 411 -7649 457
rect -7603 411 -7525 457
rect -7479 411 -7401 457
rect -7355 411 -7277 457
rect -7231 411 -7153 457
rect -7107 411 -7029 457
rect -6983 411 -6905 457
rect -6859 411 -6781 457
rect -6735 411 -6657 457
rect -6611 411 -6533 457
rect -6487 411 -6409 457
rect -6363 411 -6285 457
rect -6239 411 -6161 457
rect -6115 411 -6037 457
rect -5991 411 -5913 457
rect -5867 411 -5789 457
rect -5743 411 -5665 457
rect -5619 411 -5541 457
rect -5495 411 -5417 457
rect -5371 411 -5293 457
rect -5247 411 -5169 457
rect -5123 411 -5045 457
rect -4999 411 -4921 457
rect -4875 411 -4797 457
rect -4751 411 -4673 457
rect -4627 411 -4549 457
rect -4503 411 -4425 457
rect -4379 411 -4301 457
rect -4255 411 -4177 457
rect -4131 411 -4053 457
rect -4007 411 -3929 457
rect -3883 411 -3805 457
rect -3759 411 -3681 457
rect -3635 411 -3557 457
rect -3511 411 -3433 457
rect -3387 411 -3309 457
rect -3263 411 -3185 457
rect -3139 411 -3061 457
rect -3015 411 -2937 457
rect -2891 411 -2813 457
rect -2767 411 -2689 457
rect -2643 411 -2565 457
rect -2519 411 -2441 457
rect -2395 411 -2317 457
rect -2271 411 -2193 457
rect -2147 411 -2069 457
rect -2023 411 -1945 457
rect -1899 411 -1821 457
rect -1775 411 -1697 457
rect -1651 411 -1573 457
rect -1527 411 -1449 457
rect -1403 411 -1325 457
rect -1279 411 -1201 457
rect -1155 411 -1077 457
rect -1031 411 -953 457
rect -907 411 -829 457
rect -783 411 -705 457
rect -659 411 -581 457
rect -535 411 -457 457
rect -411 411 -333 457
rect -287 411 -209 457
rect -163 411 -85 457
rect -39 411 39 457
rect 85 411 163 457
rect 209 411 287 457
rect 333 411 411 457
rect 457 411 535 457
rect 581 411 659 457
rect 705 411 783 457
rect 829 411 907 457
rect 953 411 1031 457
rect 1077 411 1155 457
rect 1201 411 1279 457
rect 1325 411 1403 457
rect 1449 411 1527 457
rect 1573 411 1651 457
rect 1697 411 1775 457
rect 1821 411 1899 457
rect 1945 411 2023 457
rect 2069 411 2147 457
rect 2193 411 2271 457
rect 2317 411 2395 457
rect 2441 411 2519 457
rect 2565 411 2643 457
rect 2689 411 2767 457
rect 2813 411 2891 457
rect 2937 411 3015 457
rect 3061 411 3139 457
rect 3185 411 3263 457
rect 3309 411 3387 457
rect 3433 411 3511 457
rect 3557 411 3635 457
rect 3681 411 3759 457
rect 3805 411 3883 457
rect 3929 411 4007 457
rect 4053 411 4131 457
rect 4177 411 4255 457
rect 4301 411 4379 457
rect 4425 411 4503 457
rect 4549 411 4627 457
rect 4673 411 4751 457
rect 4797 411 4875 457
rect 4921 411 4999 457
rect 5045 411 5123 457
rect 5169 411 5247 457
rect 5293 411 5371 457
rect 5417 411 5495 457
rect 5541 411 5619 457
rect 5665 411 5743 457
rect 5789 411 5867 457
rect 5913 411 5991 457
rect 6037 411 6115 457
rect 6161 411 6239 457
rect 6285 411 6363 457
rect 6409 411 6487 457
rect 6533 411 6611 457
rect 6657 411 6735 457
rect 6781 411 6859 457
rect 6905 411 6983 457
rect 7029 411 7107 457
rect 7153 411 7231 457
rect 7277 411 7355 457
rect 7401 411 7479 457
rect 7525 411 7603 457
rect 7649 411 7727 457
rect 7773 411 7851 457
rect 7897 411 7975 457
rect 8021 411 8099 457
rect 8145 411 8223 457
rect 8269 411 8347 457
rect 8393 411 8471 457
rect 8517 411 8595 457
rect 8641 411 8719 457
rect 8765 411 8843 457
rect 8889 411 8967 457
rect 9013 411 9091 457
rect 9137 411 9215 457
rect 9261 411 9339 457
rect 9385 411 9463 457
rect 9509 411 9587 457
rect 9633 411 9711 457
rect 9757 411 9835 457
rect 9881 411 9959 457
rect 10005 411 10083 457
rect 10129 411 10207 457
rect 10253 411 10331 457
rect 10377 411 10455 457
rect 10501 411 10579 457
rect 10625 411 10703 457
rect 10749 411 10827 457
rect 10873 411 10951 457
rect 10997 411 11075 457
rect 11121 411 11199 457
rect 11245 411 11323 457
rect 11369 411 11447 457
rect 11493 411 11571 457
rect 11617 411 11695 457
rect 11741 411 11819 457
rect 11865 411 11943 457
rect 11989 411 12067 457
rect 12113 411 12191 457
rect 12237 411 12315 457
rect 12361 411 12439 457
rect 12485 411 12563 457
rect 12609 411 12687 457
rect 12733 411 12811 457
rect 12857 411 12935 457
rect 12981 411 13059 457
rect 13105 411 13183 457
rect 13229 411 13307 457
rect 13353 411 13431 457
rect 13477 411 13555 457
rect 13601 411 13679 457
rect 13725 411 13803 457
rect 13849 411 13927 457
rect 13973 411 14051 457
rect 14097 411 14175 457
rect 14221 411 14299 457
rect 14345 411 14423 457
rect 14469 411 14547 457
rect 14593 411 14671 457
rect 14717 411 14795 457
rect 14841 411 14919 457
rect 14965 411 15043 457
rect 15089 411 15167 457
rect 15213 411 15291 457
rect 15337 411 15415 457
rect 15461 411 15539 457
rect 15585 411 15663 457
rect 15709 411 15787 457
rect 15833 411 15911 457
rect 15957 411 16035 457
rect 16081 411 16159 457
rect 16205 411 16283 457
rect 16329 411 16407 457
rect 16453 411 16531 457
rect 16577 411 16655 457
rect 16701 411 16779 457
rect 16825 411 16903 457
rect 16949 411 17027 457
rect 17073 411 17151 457
rect 17197 411 17275 457
rect 17321 411 17332 457
rect -17332 333 17332 411
rect -17332 287 -17321 333
rect -17275 287 -17197 333
rect -17151 287 -17073 333
rect -17027 287 -16949 333
rect -16903 287 -16825 333
rect -16779 287 -16701 333
rect -16655 287 -16577 333
rect -16531 287 -16453 333
rect -16407 287 -16329 333
rect -16283 287 -16205 333
rect -16159 287 -16081 333
rect -16035 287 -15957 333
rect -15911 287 -15833 333
rect -15787 287 -15709 333
rect -15663 287 -15585 333
rect -15539 287 -15461 333
rect -15415 287 -15337 333
rect -15291 287 -15213 333
rect -15167 287 -15089 333
rect -15043 287 -14965 333
rect -14919 287 -14841 333
rect -14795 287 -14717 333
rect -14671 287 -14593 333
rect -14547 287 -14469 333
rect -14423 287 -14345 333
rect -14299 287 -14221 333
rect -14175 287 -14097 333
rect -14051 287 -13973 333
rect -13927 287 -13849 333
rect -13803 287 -13725 333
rect -13679 287 -13601 333
rect -13555 287 -13477 333
rect -13431 287 -13353 333
rect -13307 287 -13229 333
rect -13183 287 -13105 333
rect -13059 287 -12981 333
rect -12935 287 -12857 333
rect -12811 287 -12733 333
rect -12687 287 -12609 333
rect -12563 287 -12485 333
rect -12439 287 -12361 333
rect -12315 287 -12237 333
rect -12191 287 -12113 333
rect -12067 287 -11989 333
rect -11943 287 -11865 333
rect -11819 287 -11741 333
rect -11695 287 -11617 333
rect -11571 287 -11493 333
rect -11447 287 -11369 333
rect -11323 287 -11245 333
rect -11199 287 -11121 333
rect -11075 287 -10997 333
rect -10951 287 -10873 333
rect -10827 287 -10749 333
rect -10703 287 -10625 333
rect -10579 287 -10501 333
rect -10455 287 -10377 333
rect -10331 287 -10253 333
rect -10207 287 -10129 333
rect -10083 287 -10005 333
rect -9959 287 -9881 333
rect -9835 287 -9757 333
rect -9711 287 -9633 333
rect -9587 287 -9509 333
rect -9463 287 -9385 333
rect -9339 287 -9261 333
rect -9215 287 -9137 333
rect -9091 287 -9013 333
rect -8967 287 -8889 333
rect -8843 287 -8765 333
rect -8719 287 -8641 333
rect -8595 287 -8517 333
rect -8471 287 -8393 333
rect -8347 287 -8269 333
rect -8223 287 -8145 333
rect -8099 287 -8021 333
rect -7975 287 -7897 333
rect -7851 287 -7773 333
rect -7727 287 -7649 333
rect -7603 287 -7525 333
rect -7479 287 -7401 333
rect -7355 287 -7277 333
rect -7231 287 -7153 333
rect -7107 287 -7029 333
rect -6983 287 -6905 333
rect -6859 287 -6781 333
rect -6735 287 -6657 333
rect -6611 287 -6533 333
rect -6487 287 -6409 333
rect -6363 287 -6285 333
rect -6239 287 -6161 333
rect -6115 287 -6037 333
rect -5991 287 -5913 333
rect -5867 287 -5789 333
rect -5743 287 -5665 333
rect -5619 287 -5541 333
rect -5495 287 -5417 333
rect -5371 287 -5293 333
rect -5247 287 -5169 333
rect -5123 287 -5045 333
rect -4999 287 -4921 333
rect -4875 287 -4797 333
rect -4751 287 -4673 333
rect -4627 287 -4549 333
rect -4503 287 -4425 333
rect -4379 287 -4301 333
rect -4255 287 -4177 333
rect -4131 287 -4053 333
rect -4007 287 -3929 333
rect -3883 287 -3805 333
rect -3759 287 -3681 333
rect -3635 287 -3557 333
rect -3511 287 -3433 333
rect -3387 287 -3309 333
rect -3263 287 -3185 333
rect -3139 287 -3061 333
rect -3015 287 -2937 333
rect -2891 287 -2813 333
rect -2767 287 -2689 333
rect -2643 287 -2565 333
rect -2519 287 -2441 333
rect -2395 287 -2317 333
rect -2271 287 -2193 333
rect -2147 287 -2069 333
rect -2023 287 -1945 333
rect -1899 287 -1821 333
rect -1775 287 -1697 333
rect -1651 287 -1573 333
rect -1527 287 -1449 333
rect -1403 287 -1325 333
rect -1279 287 -1201 333
rect -1155 287 -1077 333
rect -1031 287 -953 333
rect -907 287 -829 333
rect -783 287 -705 333
rect -659 287 -581 333
rect -535 287 -457 333
rect -411 287 -333 333
rect -287 287 -209 333
rect -163 287 -85 333
rect -39 287 39 333
rect 85 287 163 333
rect 209 287 287 333
rect 333 287 411 333
rect 457 287 535 333
rect 581 287 659 333
rect 705 287 783 333
rect 829 287 907 333
rect 953 287 1031 333
rect 1077 287 1155 333
rect 1201 287 1279 333
rect 1325 287 1403 333
rect 1449 287 1527 333
rect 1573 287 1651 333
rect 1697 287 1775 333
rect 1821 287 1899 333
rect 1945 287 2023 333
rect 2069 287 2147 333
rect 2193 287 2271 333
rect 2317 287 2395 333
rect 2441 287 2519 333
rect 2565 287 2643 333
rect 2689 287 2767 333
rect 2813 287 2891 333
rect 2937 287 3015 333
rect 3061 287 3139 333
rect 3185 287 3263 333
rect 3309 287 3387 333
rect 3433 287 3511 333
rect 3557 287 3635 333
rect 3681 287 3759 333
rect 3805 287 3883 333
rect 3929 287 4007 333
rect 4053 287 4131 333
rect 4177 287 4255 333
rect 4301 287 4379 333
rect 4425 287 4503 333
rect 4549 287 4627 333
rect 4673 287 4751 333
rect 4797 287 4875 333
rect 4921 287 4999 333
rect 5045 287 5123 333
rect 5169 287 5247 333
rect 5293 287 5371 333
rect 5417 287 5495 333
rect 5541 287 5619 333
rect 5665 287 5743 333
rect 5789 287 5867 333
rect 5913 287 5991 333
rect 6037 287 6115 333
rect 6161 287 6239 333
rect 6285 287 6363 333
rect 6409 287 6487 333
rect 6533 287 6611 333
rect 6657 287 6735 333
rect 6781 287 6859 333
rect 6905 287 6983 333
rect 7029 287 7107 333
rect 7153 287 7231 333
rect 7277 287 7355 333
rect 7401 287 7479 333
rect 7525 287 7603 333
rect 7649 287 7727 333
rect 7773 287 7851 333
rect 7897 287 7975 333
rect 8021 287 8099 333
rect 8145 287 8223 333
rect 8269 287 8347 333
rect 8393 287 8471 333
rect 8517 287 8595 333
rect 8641 287 8719 333
rect 8765 287 8843 333
rect 8889 287 8967 333
rect 9013 287 9091 333
rect 9137 287 9215 333
rect 9261 287 9339 333
rect 9385 287 9463 333
rect 9509 287 9587 333
rect 9633 287 9711 333
rect 9757 287 9835 333
rect 9881 287 9959 333
rect 10005 287 10083 333
rect 10129 287 10207 333
rect 10253 287 10331 333
rect 10377 287 10455 333
rect 10501 287 10579 333
rect 10625 287 10703 333
rect 10749 287 10827 333
rect 10873 287 10951 333
rect 10997 287 11075 333
rect 11121 287 11199 333
rect 11245 287 11323 333
rect 11369 287 11447 333
rect 11493 287 11571 333
rect 11617 287 11695 333
rect 11741 287 11819 333
rect 11865 287 11943 333
rect 11989 287 12067 333
rect 12113 287 12191 333
rect 12237 287 12315 333
rect 12361 287 12439 333
rect 12485 287 12563 333
rect 12609 287 12687 333
rect 12733 287 12811 333
rect 12857 287 12935 333
rect 12981 287 13059 333
rect 13105 287 13183 333
rect 13229 287 13307 333
rect 13353 287 13431 333
rect 13477 287 13555 333
rect 13601 287 13679 333
rect 13725 287 13803 333
rect 13849 287 13927 333
rect 13973 287 14051 333
rect 14097 287 14175 333
rect 14221 287 14299 333
rect 14345 287 14423 333
rect 14469 287 14547 333
rect 14593 287 14671 333
rect 14717 287 14795 333
rect 14841 287 14919 333
rect 14965 287 15043 333
rect 15089 287 15167 333
rect 15213 287 15291 333
rect 15337 287 15415 333
rect 15461 287 15539 333
rect 15585 287 15663 333
rect 15709 287 15787 333
rect 15833 287 15911 333
rect 15957 287 16035 333
rect 16081 287 16159 333
rect 16205 287 16283 333
rect 16329 287 16407 333
rect 16453 287 16531 333
rect 16577 287 16655 333
rect 16701 287 16779 333
rect 16825 287 16903 333
rect 16949 287 17027 333
rect 17073 287 17151 333
rect 17197 287 17275 333
rect 17321 287 17332 333
rect -17332 209 17332 287
rect -17332 163 -17321 209
rect -17275 163 -17197 209
rect -17151 163 -17073 209
rect -17027 163 -16949 209
rect -16903 163 -16825 209
rect -16779 163 -16701 209
rect -16655 163 -16577 209
rect -16531 163 -16453 209
rect -16407 163 -16329 209
rect -16283 163 -16205 209
rect -16159 163 -16081 209
rect -16035 163 -15957 209
rect -15911 163 -15833 209
rect -15787 163 -15709 209
rect -15663 163 -15585 209
rect -15539 163 -15461 209
rect -15415 163 -15337 209
rect -15291 163 -15213 209
rect -15167 163 -15089 209
rect -15043 163 -14965 209
rect -14919 163 -14841 209
rect -14795 163 -14717 209
rect -14671 163 -14593 209
rect -14547 163 -14469 209
rect -14423 163 -14345 209
rect -14299 163 -14221 209
rect -14175 163 -14097 209
rect -14051 163 -13973 209
rect -13927 163 -13849 209
rect -13803 163 -13725 209
rect -13679 163 -13601 209
rect -13555 163 -13477 209
rect -13431 163 -13353 209
rect -13307 163 -13229 209
rect -13183 163 -13105 209
rect -13059 163 -12981 209
rect -12935 163 -12857 209
rect -12811 163 -12733 209
rect -12687 163 -12609 209
rect -12563 163 -12485 209
rect -12439 163 -12361 209
rect -12315 163 -12237 209
rect -12191 163 -12113 209
rect -12067 163 -11989 209
rect -11943 163 -11865 209
rect -11819 163 -11741 209
rect -11695 163 -11617 209
rect -11571 163 -11493 209
rect -11447 163 -11369 209
rect -11323 163 -11245 209
rect -11199 163 -11121 209
rect -11075 163 -10997 209
rect -10951 163 -10873 209
rect -10827 163 -10749 209
rect -10703 163 -10625 209
rect -10579 163 -10501 209
rect -10455 163 -10377 209
rect -10331 163 -10253 209
rect -10207 163 -10129 209
rect -10083 163 -10005 209
rect -9959 163 -9881 209
rect -9835 163 -9757 209
rect -9711 163 -9633 209
rect -9587 163 -9509 209
rect -9463 163 -9385 209
rect -9339 163 -9261 209
rect -9215 163 -9137 209
rect -9091 163 -9013 209
rect -8967 163 -8889 209
rect -8843 163 -8765 209
rect -8719 163 -8641 209
rect -8595 163 -8517 209
rect -8471 163 -8393 209
rect -8347 163 -8269 209
rect -8223 163 -8145 209
rect -8099 163 -8021 209
rect -7975 163 -7897 209
rect -7851 163 -7773 209
rect -7727 163 -7649 209
rect -7603 163 -7525 209
rect -7479 163 -7401 209
rect -7355 163 -7277 209
rect -7231 163 -7153 209
rect -7107 163 -7029 209
rect -6983 163 -6905 209
rect -6859 163 -6781 209
rect -6735 163 -6657 209
rect -6611 163 -6533 209
rect -6487 163 -6409 209
rect -6363 163 -6285 209
rect -6239 163 -6161 209
rect -6115 163 -6037 209
rect -5991 163 -5913 209
rect -5867 163 -5789 209
rect -5743 163 -5665 209
rect -5619 163 -5541 209
rect -5495 163 -5417 209
rect -5371 163 -5293 209
rect -5247 163 -5169 209
rect -5123 163 -5045 209
rect -4999 163 -4921 209
rect -4875 163 -4797 209
rect -4751 163 -4673 209
rect -4627 163 -4549 209
rect -4503 163 -4425 209
rect -4379 163 -4301 209
rect -4255 163 -4177 209
rect -4131 163 -4053 209
rect -4007 163 -3929 209
rect -3883 163 -3805 209
rect -3759 163 -3681 209
rect -3635 163 -3557 209
rect -3511 163 -3433 209
rect -3387 163 -3309 209
rect -3263 163 -3185 209
rect -3139 163 -3061 209
rect -3015 163 -2937 209
rect -2891 163 -2813 209
rect -2767 163 -2689 209
rect -2643 163 -2565 209
rect -2519 163 -2441 209
rect -2395 163 -2317 209
rect -2271 163 -2193 209
rect -2147 163 -2069 209
rect -2023 163 -1945 209
rect -1899 163 -1821 209
rect -1775 163 -1697 209
rect -1651 163 -1573 209
rect -1527 163 -1449 209
rect -1403 163 -1325 209
rect -1279 163 -1201 209
rect -1155 163 -1077 209
rect -1031 163 -953 209
rect -907 163 -829 209
rect -783 163 -705 209
rect -659 163 -581 209
rect -535 163 -457 209
rect -411 163 -333 209
rect -287 163 -209 209
rect -163 163 -85 209
rect -39 163 39 209
rect 85 163 163 209
rect 209 163 287 209
rect 333 163 411 209
rect 457 163 535 209
rect 581 163 659 209
rect 705 163 783 209
rect 829 163 907 209
rect 953 163 1031 209
rect 1077 163 1155 209
rect 1201 163 1279 209
rect 1325 163 1403 209
rect 1449 163 1527 209
rect 1573 163 1651 209
rect 1697 163 1775 209
rect 1821 163 1899 209
rect 1945 163 2023 209
rect 2069 163 2147 209
rect 2193 163 2271 209
rect 2317 163 2395 209
rect 2441 163 2519 209
rect 2565 163 2643 209
rect 2689 163 2767 209
rect 2813 163 2891 209
rect 2937 163 3015 209
rect 3061 163 3139 209
rect 3185 163 3263 209
rect 3309 163 3387 209
rect 3433 163 3511 209
rect 3557 163 3635 209
rect 3681 163 3759 209
rect 3805 163 3883 209
rect 3929 163 4007 209
rect 4053 163 4131 209
rect 4177 163 4255 209
rect 4301 163 4379 209
rect 4425 163 4503 209
rect 4549 163 4627 209
rect 4673 163 4751 209
rect 4797 163 4875 209
rect 4921 163 4999 209
rect 5045 163 5123 209
rect 5169 163 5247 209
rect 5293 163 5371 209
rect 5417 163 5495 209
rect 5541 163 5619 209
rect 5665 163 5743 209
rect 5789 163 5867 209
rect 5913 163 5991 209
rect 6037 163 6115 209
rect 6161 163 6239 209
rect 6285 163 6363 209
rect 6409 163 6487 209
rect 6533 163 6611 209
rect 6657 163 6735 209
rect 6781 163 6859 209
rect 6905 163 6983 209
rect 7029 163 7107 209
rect 7153 163 7231 209
rect 7277 163 7355 209
rect 7401 163 7479 209
rect 7525 163 7603 209
rect 7649 163 7727 209
rect 7773 163 7851 209
rect 7897 163 7975 209
rect 8021 163 8099 209
rect 8145 163 8223 209
rect 8269 163 8347 209
rect 8393 163 8471 209
rect 8517 163 8595 209
rect 8641 163 8719 209
rect 8765 163 8843 209
rect 8889 163 8967 209
rect 9013 163 9091 209
rect 9137 163 9215 209
rect 9261 163 9339 209
rect 9385 163 9463 209
rect 9509 163 9587 209
rect 9633 163 9711 209
rect 9757 163 9835 209
rect 9881 163 9959 209
rect 10005 163 10083 209
rect 10129 163 10207 209
rect 10253 163 10331 209
rect 10377 163 10455 209
rect 10501 163 10579 209
rect 10625 163 10703 209
rect 10749 163 10827 209
rect 10873 163 10951 209
rect 10997 163 11075 209
rect 11121 163 11199 209
rect 11245 163 11323 209
rect 11369 163 11447 209
rect 11493 163 11571 209
rect 11617 163 11695 209
rect 11741 163 11819 209
rect 11865 163 11943 209
rect 11989 163 12067 209
rect 12113 163 12191 209
rect 12237 163 12315 209
rect 12361 163 12439 209
rect 12485 163 12563 209
rect 12609 163 12687 209
rect 12733 163 12811 209
rect 12857 163 12935 209
rect 12981 163 13059 209
rect 13105 163 13183 209
rect 13229 163 13307 209
rect 13353 163 13431 209
rect 13477 163 13555 209
rect 13601 163 13679 209
rect 13725 163 13803 209
rect 13849 163 13927 209
rect 13973 163 14051 209
rect 14097 163 14175 209
rect 14221 163 14299 209
rect 14345 163 14423 209
rect 14469 163 14547 209
rect 14593 163 14671 209
rect 14717 163 14795 209
rect 14841 163 14919 209
rect 14965 163 15043 209
rect 15089 163 15167 209
rect 15213 163 15291 209
rect 15337 163 15415 209
rect 15461 163 15539 209
rect 15585 163 15663 209
rect 15709 163 15787 209
rect 15833 163 15911 209
rect 15957 163 16035 209
rect 16081 163 16159 209
rect 16205 163 16283 209
rect 16329 163 16407 209
rect 16453 163 16531 209
rect 16577 163 16655 209
rect 16701 163 16779 209
rect 16825 163 16903 209
rect 16949 163 17027 209
rect 17073 163 17151 209
rect 17197 163 17275 209
rect 17321 163 17332 209
rect -17332 85 17332 163
rect -17332 39 -17321 85
rect -17275 39 -17197 85
rect -17151 39 -17073 85
rect -17027 39 -16949 85
rect -16903 39 -16825 85
rect -16779 39 -16701 85
rect -16655 39 -16577 85
rect -16531 39 -16453 85
rect -16407 39 -16329 85
rect -16283 39 -16205 85
rect -16159 39 -16081 85
rect -16035 39 -15957 85
rect -15911 39 -15833 85
rect -15787 39 -15709 85
rect -15663 39 -15585 85
rect -15539 39 -15461 85
rect -15415 39 -15337 85
rect -15291 39 -15213 85
rect -15167 39 -15089 85
rect -15043 39 -14965 85
rect -14919 39 -14841 85
rect -14795 39 -14717 85
rect -14671 39 -14593 85
rect -14547 39 -14469 85
rect -14423 39 -14345 85
rect -14299 39 -14221 85
rect -14175 39 -14097 85
rect -14051 39 -13973 85
rect -13927 39 -13849 85
rect -13803 39 -13725 85
rect -13679 39 -13601 85
rect -13555 39 -13477 85
rect -13431 39 -13353 85
rect -13307 39 -13229 85
rect -13183 39 -13105 85
rect -13059 39 -12981 85
rect -12935 39 -12857 85
rect -12811 39 -12733 85
rect -12687 39 -12609 85
rect -12563 39 -12485 85
rect -12439 39 -12361 85
rect -12315 39 -12237 85
rect -12191 39 -12113 85
rect -12067 39 -11989 85
rect -11943 39 -11865 85
rect -11819 39 -11741 85
rect -11695 39 -11617 85
rect -11571 39 -11493 85
rect -11447 39 -11369 85
rect -11323 39 -11245 85
rect -11199 39 -11121 85
rect -11075 39 -10997 85
rect -10951 39 -10873 85
rect -10827 39 -10749 85
rect -10703 39 -10625 85
rect -10579 39 -10501 85
rect -10455 39 -10377 85
rect -10331 39 -10253 85
rect -10207 39 -10129 85
rect -10083 39 -10005 85
rect -9959 39 -9881 85
rect -9835 39 -9757 85
rect -9711 39 -9633 85
rect -9587 39 -9509 85
rect -9463 39 -9385 85
rect -9339 39 -9261 85
rect -9215 39 -9137 85
rect -9091 39 -9013 85
rect -8967 39 -8889 85
rect -8843 39 -8765 85
rect -8719 39 -8641 85
rect -8595 39 -8517 85
rect -8471 39 -8393 85
rect -8347 39 -8269 85
rect -8223 39 -8145 85
rect -8099 39 -8021 85
rect -7975 39 -7897 85
rect -7851 39 -7773 85
rect -7727 39 -7649 85
rect -7603 39 -7525 85
rect -7479 39 -7401 85
rect -7355 39 -7277 85
rect -7231 39 -7153 85
rect -7107 39 -7029 85
rect -6983 39 -6905 85
rect -6859 39 -6781 85
rect -6735 39 -6657 85
rect -6611 39 -6533 85
rect -6487 39 -6409 85
rect -6363 39 -6285 85
rect -6239 39 -6161 85
rect -6115 39 -6037 85
rect -5991 39 -5913 85
rect -5867 39 -5789 85
rect -5743 39 -5665 85
rect -5619 39 -5541 85
rect -5495 39 -5417 85
rect -5371 39 -5293 85
rect -5247 39 -5169 85
rect -5123 39 -5045 85
rect -4999 39 -4921 85
rect -4875 39 -4797 85
rect -4751 39 -4673 85
rect -4627 39 -4549 85
rect -4503 39 -4425 85
rect -4379 39 -4301 85
rect -4255 39 -4177 85
rect -4131 39 -4053 85
rect -4007 39 -3929 85
rect -3883 39 -3805 85
rect -3759 39 -3681 85
rect -3635 39 -3557 85
rect -3511 39 -3433 85
rect -3387 39 -3309 85
rect -3263 39 -3185 85
rect -3139 39 -3061 85
rect -3015 39 -2937 85
rect -2891 39 -2813 85
rect -2767 39 -2689 85
rect -2643 39 -2565 85
rect -2519 39 -2441 85
rect -2395 39 -2317 85
rect -2271 39 -2193 85
rect -2147 39 -2069 85
rect -2023 39 -1945 85
rect -1899 39 -1821 85
rect -1775 39 -1697 85
rect -1651 39 -1573 85
rect -1527 39 -1449 85
rect -1403 39 -1325 85
rect -1279 39 -1201 85
rect -1155 39 -1077 85
rect -1031 39 -953 85
rect -907 39 -829 85
rect -783 39 -705 85
rect -659 39 -581 85
rect -535 39 -457 85
rect -411 39 -333 85
rect -287 39 -209 85
rect -163 39 -85 85
rect -39 39 39 85
rect 85 39 163 85
rect 209 39 287 85
rect 333 39 411 85
rect 457 39 535 85
rect 581 39 659 85
rect 705 39 783 85
rect 829 39 907 85
rect 953 39 1031 85
rect 1077 39 1155 85
rect 1201 39 1279 85
rect 1325 39 1403 85
rect 1449 39 1527 85
rect 1573 39 1651 85
rect 1697 39 1775 85
rect 1821 39 1899 85
rect 1945 39 2023 85
rect 2069 39 2147 85
rect 2193 39 2271 85
rect 2317 39 2395 85
rect 2441 39 2519 85
rect 2565 39 2643 85
rect 2689 39 2767 85
rect 2813 39 2891 85
rect 2937 39 3015 85
rect 3061 39 3139 85
rect 3185 39 3263 85
rect 3309 39 3387 85
rect 3433 39 3511 85
rect 3557 39 3635 85
rect 3681 39 3759 85
rect 3805 39 3883 85
rect 3929 39 4007 85
rect 4053 39 4131 85
rect 4177 39 4255 85
rect 4301 39 4379 85
rect 4425 39 4503 85
rect 4549 39 4627 85
rect 4673 39 4751 85
rect 4797 39 4875 85
rect 4921 39 4999 85
rect 5045 39 5123 85
rect 5169 39 5247 85
rect 5293 39 5371 85
rect 5417 39 5495 85
rect 5541 39 5619 85
rect 5665 39 5743 85
rect 5789 39 5867 85
rect 5913 39 5991 85
rect 6037 39 6115 85
rect 6161 39 6239 85
rect 6285 39 6363 85
rect 6409 39 6487 85
rect 6533 39 6611 85
rect 6657 39 6735 85
rect 6781 39 6859 85
rect 6905 39 6983 85
rect 7029 39 7107 85
rect 7153 39 7231 85
rect 7277 39 7355 85
rect 7401 39 7479 85
rect 7525 39 7603 85
rect 7649 39 7727 85
rect 7773 39 7851 85
rect 7897 39 7975 85
rect 8021 39 8099 85
rect 8145 39 8223 85
rect 8269 39 8347 85
rect 8393 39 8471 85
rect 8517 39 8595 85
rect 8641 39 8719 85
rect 8765 39 8843 85
rect 8889 39 8967 85
rect 9013 39 9091 85
rect 9137 39 9215 85
rect 9261 39 9339 85
rect 9385 39 9463 85
rect 9509 39 9587 85
rect 9633 39 9711 85
rect 9757 39 9835 85
rect 9881 39 9959 85
rect 10005 39 10083 85
rect 10129 39 10207 85
rect 10253 39 10331 85
rect 10377 39 10455 85
rect 10501 39 10579 85
rect 10625 39 10703 85
rect 10749 39 10827 85
rect 10873 39 10951 85
rect 10997 39 11075 85
rect 11121 39 11199 85
rect 11245 39 11323 85
rect 11369 39 11447 85
rect 11493 39 11571 85
rect 11617 39 11695 85
rect 11741 39 11819 85
rect 11865 39 11943 85
rect 11989 39 12067 85
rect 12113 39 12191 85
rect 12237 39 12315 85
rect 12361 39 12439 85
rect 12485 39 12563 85
rect 12609 39 12687 85
rect 12733 39 12811 85
rect 12857 39 12935 85
rect 12981 39 13059 85
rect 13105 39 13183 85
rect 13229 39 13307 85
rect 13353 39 13431 85
rect 13477 39 13555 85
rect 13601 39 13679 85
rect 13725 39 13803 85
rect 13849 39 13927 85
rect 13973 39 14051 85
rect 14097 39 14175 85
rect 14221 39 14299 85
rect 14345 39 14423 85
rect 14469 39 14547 85
rect 14593 39 14671 85
rect 14717 39 14795 85
rect 14841 39 14919 85
rect 14965 39 15043 85
rect 15089 39 15167 85
rect 15213 39 15291 85
rect 15337 39 15415 85
rect 15461 39 15539 85
rect 15585 39 15663 85
rect 15709 39 15787 85
rect 15833 39 15911 85
rect 15957 39 16035 85
rect 16081 39 16159 85
rect 16205 39 16283 85
rect 16329 39 16407 85
rect 16453 39 16531 85
rect 16577 39 16655 85
rect 16701 39 16779 85
rect 16825 39 16903 85
rect 16949 39 17027 85
rect 17073 39 17151 85
rect 17197 39 17275 85
rect 17321 39 17332 85
rect -17332 -39 17332 39
rect -17332 -85 -17321 -39
rect -17275 -85 -17197 -39
rect -17151 -85 -17073 -39
rect -17027 -85 -16949 -39
rect -16903 -85 -16825 -39
rect -16779 -85 -16701 -39
rect -16655 -85 -16577 -39
rect -16531 -85 -16453 -39
rect -16407 -85 -16329 -39
rect -16283 -85 -16205 -39
rect -16159 -85 -16081 -39
rect -16035 -85 -15957 -39
rect -15911 -85 -15833 -39
rect -15787 -85 -15709 -39
rect -15663 -85 -15585 -39
rect -15539 -85 -15461 -39
rect -15415 -85 -15337 -39
rect -15291 -85 -15213 -39
rect -15167 -85 -15089 -39
rect -15043 -85 -14965 -39
rect -14919 -85 -14841 -39
rect -14795 -85 -14717 -39
rect -14671 -85 -14593 -39
rect -14547 -85 -14469 -39
rect -14423 -85 -14345 -39
rect -14299 -85 -14221 -39
rect -14175 -85 -14097 -39
rect -14051 -85 -13973 -39
rect -13927 -85 -13849 -39
rect -13803 -85 -13725 -39
rect -13679 -85 -13601 -39
rect -13555 -85 -13477 -39
rect -13431 -85 -13353 -39
rect -13307 -85 -13229 -39
rect -13183 -85 -13105 -39
rect -13059 -85 -12981 -39
rect -12935 -85 -12857 -39
rect -12811 -85 -12733 -39
rect -12687 -85 -12609 -39
rect -12563 -85 -12485 -39
rect -12439 -85 -12361 -39
rect -12315 -85 -12237 -39
rect -12191 -85 -12113 -39
rect -12067 -85 -11989 -39
rect -11943 -85 -11865 -39
rect -11819 -85 -11741 -39
rect -11695 -85 -11617 -39
rect -11571 -85 -11493 -39
rect -11447 -85 -11369 -39
rect -11323 -85 -11245 -39
rect -11199 -85 -11121 -39
rect -11075 -85 -10997 -39
rect -10951 -85 -10873 -39
rect -10827 -85 -10749 -39
rect -10703 -85 -10625 -39
rect -10579 -85 -10501 -39
rect -10455 -85 -10377 -39
rect -10331 -85 -10253 -39
rect -10207 -85 -10129 -39
rect -10083 -85 -10005 -39
rect -9959 -85 -9881 -39
rect -9835 -85 -9757 -39
rect -9711 -85 -9633 -39
rect -9587 -85 -9509 -39
rect -9463 -85 -9385 -39
rect -9339 -85 -9261 -39
rect -9215 -85 -9137 -39
rect -9091 -85 -9013 -39
rect -8967 -85 -8889 -39
rect -8843 -85 -8765 -39
rect -8719 -85 -8641 -39
rect -8595 -85 -8517 -39
rect -8471 -85 -8393 -39
rect -8347 -85 -8269 -39
rect -8223 -85 -8145 -39
rect -8099 -85 -8021 -39
rect -7975 -85 -7897 -39
rect -7851 -85 -7773 -39
rect -7727 -85 -7649 -39
rect -7603 -85 -7525 -39
rect -7479 -85 -7401 -39
rect -7355 -85 -7277 -39
rect -7231 -85 -7153 -39
rect -7107 -85 -7029 -39
rect -6983 -85 -6905 -39
rect -6859 -85 -6781 -39
rect -6735 -85 -6657 -39
rect -6611 -85 -6533 -39
rect -6487 -85 -6409 -39
rect -6363 -85 -6285 -39
rect -6239 -85 -6161 -39
rect -6115 -85 -6037 -39
rect -5991 -85 -5913 -39
rect -5867 -85 -5789 -39
rect -5743 -85 -5665 -39
rect -5619 -85 -5541 -39
rect -5495 -85 -5417 -39
rect -5371 -85 -5293 -39
rect -5247 -85 -5169 -39
rect -5123 -85 -5045 -39
rect -4999 -85 -4921 -39
rect -4875 -85 -4797 -39
rect -4751 -85 -4673 -39
rect -4627 -85 -4549 -39
rect -4503 -85 -4425 -39
rect -4379 -85 -4301 -39
rect -4255 -85 -4177 -39
rect -4131 -85 -4053 -39
rect -4007 -85 -3929 -39
rect -3883 -85 -3805 -39
rect -3759 -85 -3681 -39
rect -3635 -85 -3557 -39
rect -3511 -85 -3433 -39
rect -3387 -85 -3309 -39
rect -3263 -85 -3185 -39
rect -3139 -85 -3061 -39
rect -3015 -85 -2937 -39
rect -2891 -85 -2813 -39
rect -2767 -85 -2689 -39
rect -2643 -85 -2565 -39
rect -2519 -85 -2441 -39
rect -2395 -85 -2317 -39
rect -2271 -85 -2193 -39
rect -2147 -85 -2069 -39
rect -2023 -85 -1945 -39
rect -1899 -85 -1821 -39
rect -1775 -85 -1697 -39
rect -1651 -85 -1573 -39
rect -1527 -85 -1449 -39
rect -1403 -85 -1325 -39
rect -1279 -85 -1201 -39
rect -1155 -85 -1077 -39
rect -1031 -85 -953 -39
rect -907 -85 -829 -39
rect -783 -85 -705 -39
rect -659 -85 -581 -39
rect -535 -85 -457 -39
rect -411 -85 -333 -39
rect -287 -85 -209 -39
rect -163 -85 -85 -39
rect -39 -85 39 -39
rect 85 -85 163 -39
rect 209 -85 287 -39
rect 333 -85 411 -39
rect 457 -85 535 -39
rect 581 -85 659 -39
rect 705 -85 783 -39
rect 829 -85 907 -39
rect 953 -85 1031 -39
rect 1077 -85 1155 -39
rect 1201 -85 1279 -39
rect 1325 -85 1403 -39
rect 1449 -85 1527 -39
rect 1573 -85 1651 -39
rect 1697 -85 1775 -39
rect 1821 -85 1899 -39
rect 1945 -85 2023 -39
rect 2069 -85 2147 -39
rect 2193 -85 2271 -39
rect 2317 -85 2395 -39
rect 2441 -85 2519 -39
rect 2565 -85 2643 -39
rect 2689 -85 2767 -39
rect 2813 -85 2891 -39
rect 2937 -85 3015 -39
rect 3061 -85 3139 -39
rect 3185 -85 3263 -39
rect 3309 -85 3387 -39
rect 3433 -85 3511 -39
rect 3557 -85 3635 -39
rect 3681 -85 3759 -39
rect 3805 -85 3883 -39
rect 3929 -85 4007 -39
rect 4053 -85 4131 -39
rect 4177 -85 4255 -39
rect 4301 -85 4379 -39
rect 4425 -85 4503 -39
rect 4549 -85 4627 -39
rect 4673 -85 4751 -39
rect 4797 -85 4875 -39
rect 4921 -85 4999 -39
rect 5045 -85 5123 -39
rect 5169 -85 5247 -39
rect 5293 -85 5371 -39
rect 5417 -85 5495 -39
rect 5541 -85 5619 -39
rect 5665 -85 5743 -39
rect 5789 -85 5867 -39
rect 5913 -85 5991 -39
rect 6037 -85 6115 -39
rect 6161 -85 6239 -39
rect 6285 -85 6363 -39
rect 6409 -85 6487 -39
rect 6533 -85 6611 -39
rect 6657 -85 6735 -39
rect 6781 -85 6859 -39
rect 6905 -85 6983 -39
rect 7029 -85 7107 -39
rect 7153 -85 7231 -39
rect 7277 -85 7355 -39
rect 7401 -85 7479 -39
rect 7525 -85 7603 -39
rect 7649 -85 7727 -39
rect 7773 -85 7851 -39
rect 7897 -85 7975 -39
rect 8021 -85 8099 -39
rect 8145 -85 8223 -39
rect 8269 -85 8347 -39
rect 8393 -85 8471 -39
rect 8517 -85 8595 -39
rect 8641 -85 8719 -39
rect 8765 -85 8843 -39
rect 8889 -85 8967 -39
rect 9013 -85 9091 -39
rect 9137 -85 9215 -39
rect 9261 -85 9339 -39
rect 9385 -85 9463 -39
rect 9509 -85 9587 -39
rect 9633 -85 9711 -39
rect 9757 -85 9835 -39
rect 9881 -85 9959 -39
rect 10005 -85 10083 -39
rect 10129 -85 10207 -39
rect 10253 -85 10331 -39
rect 10377 -85 10455 -39
rect 10501 -85 10579 -39
rect 10625 -85 10703 -39
rect 10749 -85 10827 -39
rect 10873 -85 10951 -39
rect 10997 -85 11075 -39
rect 11121 -85 11199 -39
rect 11245 -85 11323 -39
rect 11369 -85 11447 -39
rect 11493 -85 11571 -39
rect 11617 -85 11695 -39
rect 11741 -85 11819 -39
rect 11865 -85 11943 -39
rect 11989 -85 12067 -39
rect 12113 -85 12191 -39
rect 12237 -85 12315 -39
rect 12361 -85 12439 -39
rect 12485 -85 12563 -39
rect 12609 -85 12687 -39
rect 12733 -85 12811 -39
rect 12857 -85 12935 -39
rect 12981 -85 13059 -39
rect 13105 -85 13183 -39
rect 13229 -85 13307 -39
rect 13353 -85 13431 -39
rect 13477 -85 13555 -39
rect 13601 -85 13679 -39
rect 13725 -85 13803 -39
rect 13849 -85 13927 -39
rect 13973 -85 14051 -39
rect 14097 -85 14175 -39
rect 14221 -85 14299 -39
rect 14345 -85 14423 -39
rect 14469 -85 14547 -39
rect 14593 -85 14671 -39
rect 14717 -85 14795 -39
rect 14841 -85 14919 -39
rect 14965 -85 15043 -39
rect 15089 -85 15167 -39
rect 15213 -85 15291 -39
rect 15337 -85 15415 -39
rect 15461 -85 15539 -39
rect 15585 -85 15663 -39
rect 15709 -85 15787 -39
rect 15833 -85 15911 -39
rect 15957 -85 16035 -39
rect 16081 -85 16159 -39
rect 16205 -85 16283 -39
rect 16329 -85 16407 -39
rect 16453 -85 16531 -39
rect 16577 -85 16655 -39
rect 16701 -85 16779 -39
rect 16825 -85 16903 -39
rect 16949 -85 17027 -39
rect 17073 -85 17151 -39
rect 17197 -85 17275 -39
rect 17321 -85 17332 -39
rect -17332 -163 17332 -85
rect -17332 -209 -17321 -163
rect -17275 -209 -17197 -163
rect -17151 -209 -17073 -163
rect -17027 -209 -16949 -163
rect -16903 -209 -16825 -163
rect -16779 -209 -16701 -163
rect -16655 -209 -16577 -163
rect -16531 -209 -16453 -163
rect -16407 -209 -16329 -163
rect -16283 -209 -16205 -163
rect -16159 -209 -16081 -163
rect -16035 -209 -15957 -163
rect -15911 -209 -15833 -163
rect -15787 -209 -15709 -163
rect -15663 -209 -15585 -163
rect -15539 -209 -15461 -163
rect -15415 -209 -15337 -163
rect -15291 -209 -15213 -163
rect -15167 -209 -15089 -163
rect -15043 -209 -14965 -163
rect -14919 -209 -14841 -163
rect -14795 -209 -14717 -163
rect -14671 -209 -14593 -163
rect -14547 -209 -14469 -163
rect -14423 -209 -14345 -163
rect -14299 -209 -14221 -163
rect -14175 -209 -14097 -163
rect -14051 -209 -13973 -163
rect -13927 -209 -13849 -163
rect -13803 -209 -13725 -163
rect -13679 -209 -13601 -163
rect -13555 -209 -13477 -163
rect -13431 -209 -13353 -163
rect -13307 -209 -13229 -163
rect -13183 -209 -13105 -163
rect -13059 -209 -12981 -163
rect -12935 -209 -12857 -163
rect -12811 -209 -12733 -163
rect -12687 -209 -12609 -163
rect -12563 -209 -12485 -163
rect -12439 -209 -12361 -163
rect -12315 -209 -12237 -163
rect -12191 -209 -12113 -163
rect -12067 -209 -11989 -163
rect -11943 -209 -11865 -163
rect -11819 -209 -11741 -163
rect -11695 -209 -11617 -163
rect -11571 -209 -11493 -163
rect -11447 -209 -11369 -163
rect -11323 -209 -11245 -163
rect -11199 -209 -11121 -163
rect -11075 -209 -10997 -163
rect -10951 -209 -10873 -163
rect -10827 -209 -10749 -163
rect -10703 -209 -10625 -163
rect -10579 -209 -10501 -163
rect -10455 -209 -10377 -163
rect -10331 -209 -10253 -163
rect -10207 -209 -10129 -163
rect -10083 -209 -10005 -163
rect -9959 -209 -9881 -163
rect -9835 -209 -9757 -163
rect -9711 -209 -9633 -163
rect -9587 -209 -9509 -163
rect -9463 -209 -9385 -163
rect -9339 -209 -9261 -163
rect -9215 -209 -9137 -163
rect -9091 -209 -9013 -163
rect -8967 -209 -8889 -163
rect -8843 -209 -8765 -163
rect -8719 -209 -8641 -163
rect -8595 -209 -8517 -163
rect -8471 -209 -8393 -163
rect -8347 -209 -8269 -163
rect -8223 -209 -8145 -163
rect -8099 -209 -8021 -163
rect -7975 -209 -7897 -163
rect -7851 -209 -7773 -163
rect -7727 -209 -7649 -163
rect -7603 -209 -7525 -163
rect -7479 -209 -7401 -163
rect -7355 -209 -7277 -163
rect -7231 -209 -7153 -163
rect -7107 -209 -7029 -163
rect -6983 -209 -6905 -163
rect -6859 -209 -6781 -163
rect -6735 -209 -6657 -163
rect -6611 -209 -6533 -163
rect -6487 -209 -6409 -163
rect -6363 -209 -6285 -163
rect -6239 -209 -6161 -163
rect -6115 -209 -6037 -163
rect -5991 -209 -5913 -163
rect -5867 -209 -5789 -163
rect -5743 -209 -5665 -163
rect -5619 -209 -5541 -163
rect -5495 -209 -5417 -163
rect -5371 -209 -5293 -163
rect -5247 -209 -5169 -163
rect -5123 -209 -5045 -163
rect -4999 -209 -4921 -163
rect -4875 -209 -4797 -163
rect -4751 -209 -4673 -163
rect -4627 -209 -4549 -163
rect -4503 -209 -4425 -163
rect -4379 -209 -4301 -163
rect -4255 -209 -4177 -163
rect -4131 -209 -4053 -163
rect -4007 -209 -3929 -163
rect -3883 -209 -3805 -163
rect -3759 -209 -3681 -163
rect -3635 -209 -3557 -163
rect -3511 -209 -3433 -163
rect -3387 -209 -3309 -163
rect -3263 -209 -3185 -163
rect -3139 -209 -3061 -163
rect -3015 -209 -2937 -163
rect -2891 -209 -2813 -163
rect -2767 -209 -2689 -163
rect -2643 -209 -2565 -163
rect -2519 -209 -2441 -163
rect -2395 -209 -2317 -163
rect -2271 -209 -2193 -163
rect -2147 -209 -2069 -163
rect -2023 -209 -1945 -163
rect -1899 -209 -1821 -163
rect -1775 -209 -1697 -163
rect -1651 -209 -1573 -163
rect -1527 -209 -1449 -163
rect -1403 -209 -1325 -163
rect -1279 -209 -1201 -163
rect -1155 -209 -1077 -163
rect -1031 -209 -953 -163
rect -907 -209 -829 -163
rect -783 -209 -705 -163
rect -659 -209 -581 -163
rect -535 -209 -457 -163
rect -411 -209 -333 -163
rect -287 -209 -209 -163
rect -163 -209 -85 -163
rect -39 -209 39 -163
rect 85 -209 163 -163
rect 209 -209 287 -163
rect 333 -209 411 -163
rect 457 -209 535 -163
rect 581 -209 659 -163
rect 705 -209 783 -163
rect 829 -209 907 -163
rect 953 -209 1031 -163
rect 1077 -209 1155 -163
rect 1201 -209 1279 -163
rect 1325 -209 1403 -163
rect 1449 -209 1527 -163
rect 1573 -209 1651 -163
rect 1697 -209 1775 -163
rect 1821 -209 1899 -163
rect 1945 -209 2023 -163
rect 2069 -209 2147 -163
rect 2193 -209 2271 -163
rect 2317 -209 2395 -163
rect 2441 -209 2519 -163
rect 2565 -209 2643 -163
rect 2689 -209 2767 -163
rect 2813 -209 2891 -163
rect 2937 -209 3015 -163
rect 3061 -209 3139 -163
rect 3185 -209 3263 -163
rect 3309 -209 3387 -163
rect 3433 -209 3511 -163
rect 3557 -209 3635 -163
rect 3681 -209 3759 -163
rect 3805 -209 3883 -163
rect 3929 -209 4007 -163
rect 4053 -209 4131 -163
rect 4177 -209 4255 -163
rect 4301 -209 4379 -163
rect 4425 -209 4503 -163
rect 4549 -209 4627 -163
rect 4673 -209 4751 -163
rect 4797 -209 4875 -163
rect 4921 -209 4999 -163
rect 5045 -209 5123 -163
rect 5169 -209 5247 -163
rect 5293 -209 5371 -163
rect 5417 -209 5495 -163
rect 5541 -209 5619 -163
rect 5665 -209 5743 -163
rect 5789 -209 5867 -163
rect 5913 -209 5991 -163
rect 6037 -209 6115 -163
rect 6161 -209 6239 -163
rect 6285 -209 6363 -163
rect 6409 -209 6487 -163
rect 6533 -209 6611 -163
rect 6657 -209 6735 -163
rect 6781 -209 6859 -163
rect 6905 -209 6983 -163
rect 7029 -209 7107 -163
rect 7153 -209 7231 -163
rect 7277 -209 7355 -163
rect 7401 -209 7479 -163
rect 7525 -209 7603 -163
rect 7649 -209 7727 -163
rect 7773 -209 7851 -163
rect 7897 -209 7975 -163
rect 8021 -209 8099 -163
rect 8145 -209 8223 -163
rect 8269 -209 8347 -163
rect 8393 -209 8471 -163
rect 8517 -209 8595 -163
rect 8641 -209 8719 -163
rect 8765 -209 8843 -163
rect 8889 -209 8967 -163
rect 9013 -209 9091 -163
rect 9137 -209 9215 -163
rect 9261 -209 9339 -163
rect 9385 -209 9463 -163
rect 9509 -209 9587 -163
rect 9633 -209 9711 -163
rect 9757 -209 9835 -163
rect 9881 -209 9959 -163
rect 10005 -209 10083 -163
rect 10129 -209 10207 -163
rect 10253 -209 10331 -163
rect 10377 -209 10455 -163
rect 10501 -209 10579 -163
rect 10625 -209 10703 -163
rect 10749 -209 10827 -163
rect 10873 -209 10951 -163
rect 10997 -209 11075 -163
rect 11121 -209 11199 -163
rect 11245 -209 11323 -163
rect 11369 -209 11447 -163
rect 11493 -209 11571 -163
rect 11617 -209 11695 -163
rect 11741 -209 11819 -163
rect 11865 -209 11943 -163
rect 11989 -209 12067 -163
rect 12113 -209 12191 -163
rect 12237 -209 12315 -163
rect 12361 -209 12439 -163
rect 12485 -209 12563 -163
rect 12609 -209 12687 -163
rect 12733 -209 12811 -163
rect 12857 -209 12935 -163
rect 12981 -209 13059 -163
rect 13105 -209 13183 -163
rect 13229 -209 13307 -163
rect 13353 -209 13431 -163
rect 13477 -209 13555 -163
rect 13601 -209 13679 -163
rect 13725 -209 13803 -163
rect 13849 -209 13927 -163
rect 13973 -209 14051 -163
rect 14097 -209 14175 -163
rect 14221 -209 14299 -163
rect 14345 -209 14423 -163
rect 14469 -209 14547 -163
rect 14593 -209 14671 -163
rect 14717 -209 14795 -163
rect 14841 -209 14919 -163
rect 14965 -209 15043 -163
rect 15089 -209 15167 -163
rect 15213 -209 15291 -163
rect 15337 -209 15415 -163
rect 15461 -209 15539 -163
rect 15585 -209 15663 -163
rect 15709 -209 15787 -163
rect 15833 -209 15911 -163
rect 15957 -209 16035 -163
rect 16081 -209 16159 -163
rect 16205 -209 16283 -163
rect 16329 -209 16407 -163
rect 16453 -209 16531 -163
rect 16577 -209 16655 -163
rect 16701 -209 16779 -163
rect 16825 -209 16903 -163
rect 16949 -209 17027 -163
rect 17073 -209 17151 -163
rect 17197 -209 17275 -163
rect 17321 -209 17332 -163
rect -17332 -287 17332 -209
rect -17332 -333 -17321 -287
rect -17275 -333 -17197 -287
rect -17151 -333 -17073 -287
rect -17027 -333 -16949 -287
rect -16903 -333 -16825 -287
rect -16779 -333 -16701 -287
rect -16655 -333 -16577 -287
rect -16531 -333 -16453 -287
rect -16407 -333 -16329 -287
rect -16283 -333 -16205 -287
rect -16159 -333 -16081 -287
rect -16035 -333 -15957 -287
rect -15911 -333 -15833 -287
rect -15787 -333 -15709 -287
rect -15663 -333 -15585 -287
rect -15539 -333 -15461 -287
rect -15415 -333 -15337 -287
rect -15291 -333 -15213 -287
rect -15167 -333 -15089 -287
rect -15043 -333 -14965 -287
rect -14919 -333 -14841 -287
rect -14795 -333 -14717 -287
rect -14671 -333 -14593 -287
rect -14547 -333 -14469 -287
rect -14423 -333 -14345 -287
rect -14299 -333 -14221 -287
rect -14175 -333 -14097 -287
rect -14051 -333 -13973 -287
rect -13927 -333 -13849 -287
rect -13803 -333 -13725 -287
rect -13679 -333 -13601 -287
rect -13555 -333 -13477 -287
rect -13431 -333 -13353 -287
rect -13307 -333 -13229 -287
rect -13183 -333 -13105 -287
rect -13059 -333 -12981 -287
rect -12935 -333 -12857 -287
rect -12811 -333 -12733 -287
rect -12687 -333 -12609 -287
rect -12563 -333 -12485 -287
rect -12439 -333 -12361 -287
rect -12315 -333 -12237 -287
rect -12191 -333 -12113 -287
rect -12067 -333 -11989 -287
rect -11943 -333 -11865 -287
rect -11819 -333 -11741 -287
rect -11695 -333 -11617 -287
rect -11571 -333 -11493 -287
rect -11447 -333 -11369 -287
rect -11323 -333 -11245 -287
rect -11199 -333 -11121 -287
rect -11075 -333 -10997 -287
rect -10951 -333 -10873 -287
rect -10827 -333 -10749 -287
rect -10703 -333 -10625 -287
rect -10579 -333 -10501 -287
rect -10455 -333 -10377 -287
rect -10331 -333 -10253 -287
rect -10207 -333 -10129 -287
rect -10083 -333 -10005 -287
rect -9959 -333 -9881 -287
rect -9835 -333 -9757 -287
rect -9711 -333 -9633 -287
rect -9587 -333 -9509 -287
rect -9463 -333 -9385 -287
rect -9339 -333 -9261 -287
rect -9215 -333 -9137 -287
rect -9091 -333 -9013 -287
rect -8967 -333 -8889 -287
rect -8843 -333 -8765 -287
rect -8719 -333 -8641 -287
rect -8595 -333 -8517 -287
rect -8471 -333 -8393 -287
rect -8347 -333 -8269 -287
rect -8223 -333 -8145 -287
rect -8099 -333 -8021 -287
rect -7975 -333 -7897 -287
rect -7851 -333 -7773 -287
rect -7727 -333 -7649 -287
rect -7603 -333 -7525 -287
rect -7479 -333 -7401 -287
rect -7355 -333 -7277 -287
rect -7231 -333 -7153 -287
rect -7107 -333 -7029 -287
rect -6983 -333 -6905 -287
rect -6859 -333 -6781 -287
rect -6735 -333 -6657 -287
rect -6611 -333 -6533 -287
rect -6487 -333 -6409 -287
rect -6363 -333 -6285 -287
rect -6239 -333 -6161 -287
rect -6115 -333 -6037 -287
rect -5991 -333 -5913 -287
rect -5867 -333 -5789 -287
rect -5743 -333 -5665 -287
rect -5619 -333 -5541 -287
rect -5495 -333 -5417 -287
rect -5371 -333 -5293 -287
rect -5247 -333 -5169 -287
rect -5123 -333 -5045 -287
rect -4999 -333 -4921 -287
rect -4875 -333 -4797 -287
rect -4751 -333 -4673 -287
rect -4627 -333 -4549 -287
rect -4503 -333 -4425 -287
rect -4379 -333 -4301 -287
rect -4255 -333 -4177 -287
rect -4131 -333 -4053 -287
rect -4007 -333 -3929 -287
rect -3883 -333 -3805 -287
rect -3759 -333 -3681 -287
rect -3635 -333 -3557 -287
rect -3511 -333 -3433 -287
rect -3387 -333 -3309 -287
rect -3263 -333 -3185 -287
rect -3139 -333 -3061 -287
rect -3015 -333 -2937 -287
rect -2891 -333 -2813 -287
rect -2767 -333 -2689 -287
rect -2643 -333 -2565 -287
rect -2519 -333 -2441 -287
rect -2395 -333 -2317 -287
rect -2271 -333 -2193 -287
rect -2147 -333 -2069 -287
rect -2023 -333 -1945 -287
rect -1899 -333 -1821 -287
rect -1775 -333 -1697 -287
rect -1651 -333 -1573 -287
rect -1527 -333 -1449 -287
rect -1403 -333 -1325 -287
rect -1279 -333 -1201 -287
rect -1155 -333 -1077 -287
rect -1031 -333 -953 -287
rect -907 -333 -829 -287
rect -783 -333 -705 -287
rect -659 -333 -581 -287
rect -535 -333 -457 -287
rect -411 -333 -333 -287
rect -287 -333 -209 -287
rect -163 -333 -85 -287
rect -39 -333 39 -287
rect 85 -333 163 -287
rect 209 -333 287 -287
rect 333 -333 411 -287
rect 457 -333 535 -287
rect 581 -333 659 -287
rect 705 -333 783 -287
rect 829 -333 907 -287
rect 953 -333 1031 -287
rect 1077 -333 1155 -287
rect 1201 -333 1279 -287
rect 1325 -333 1403 -287
rect 1449 -333 1527 -287
rect 1573 -333 1651 -287
rect 1697 -333 1775 -287
rect 1821 -333 1899 -287
rect 1945 -333 2023 -287
rect 2069 -333 2147 -287
rect 2193 -333 2271 -287
rect 2317 -333 2395 -287
rect 2441 -333 2519 -287
rect 2565 -333 2643 -287
rect 2689 -333 2767 -287
rect 2813 -333 2891 -287
rect 2937 -333 3015 -287
rect 3061 -333 3139 -287
rect 3185 -333 3263 -287
rect 3309 -333 3387 -287
rect 3433 -333 3511 -287
rect 3557 -333 3635 -287
rect 3681 -333 3759 -287
rect 3805 -333 3883 -287
rect 3929 -333 4007 -287
rect 4053 -333 4131 -287
rect 4177 -333 4255 -287
rect 4301 -333 4379 -287
rect 4425 -333 4503 -287
rect 4549 -333 4627 -287
rect 4673 -333 4751 -287
rect 4797 -333 4875 -287
rect 4921 -333 4999 -287
rect 5045 -333 5123 -287
rect 5169 -333 5247 -287
rect 5293 -333 5371 -287
rect 5417 -333 5495 -287
rect 5541 -333 5619 -287
rect 5665 -333 5743 -287
rect 5789 -333 5867 -287
rect 5913 -333 5991 -287
rect 6037 -333 6115 -287
rect 6161 -333 6239 -287
rect 6285 -333 6363 -287
rect 6409 -333 6487 -287
rect 6533 -333 6611 -287
rect 6657 -333 6735 -287
rect 6781 -333 6859 -287
rect 6905 -333 6983 -287
rect 7029 -333 7107 -287
rect 7153 -333 7231 -287
rect 7277 -333 7355 -287
rect 7401 -333 7479 -287
rect 7525 -333 7603 -287
rect 7649 -333 7727 -287
rect 7773 -333 7851 -287
rect 7897 -333 7975 -287
rect 8021 -333 8099 -287
rect 8145 -333 8223 -287
rect 8269 -333 8347 -287
rect 8393 -333 8471 -287
rect 8517 -333 8595 -287
rect 8641 -333 8719 -287
rect 8765 -333 8843 -287
rect 8889 -333 8967 -287
rect 9013 -333 9091 -287
rect 9137 -333 9215 -287
rect 9261 -333 9339 -287
rect 9385 -333 9463 -287
rect 9509 -333 9587 -287
rect 9633 -333 9711 -287
rect 9757 -333 9835 -287
rect 9881 -333 9959 -287
rect 10005 -333 10083 -287
rect 10129 -333 10207 -287
rect 10253 -333 10331 -287
rect 10377 -333 10455 -287
rect 10501 -333 10579 -287
rect 10625 -333 10703 -287
rect 10749 -333 10827 -287
rect 10873 -333 10951 -287
rect 10997 -333 11075 -287
rect 11121 -333 11199 -287
rect 11245 -333 11323 -287
rect 11369 -333 11447 -287
rect 11493 -333 11571 -287
rect 11617 -333 11695 -287
rect 11741 -333 11819 -287
rect 11865 -333 11943 -287
rect 11989 -333 12067 -287
rect 12113 -333 12191 -287
rect 12237 -333 12315 -287
rect 12361 -333 12439 -287
rect 12485 -333 12563 -287
rect 12609 -333 12687 -287
rect 12733 -333 12811 -287
rect 12857 -333 12935 -287
rect 12981 -333 13059 -287
rect 13105 -333 13183 -287
rect 13229 -333 13307 -287
rect 13353 -333 13431 -287
rect 13477 -333 13555 -287
rect 13601 -333 13679 -287
rect 13725 -333 13803 -287
rect 13849 -333 13927 -287
rect 13973 -333 14051 -287
rect 14097 -333 14175 -287
rect 14221 -333 14299 -287
rect 14345 -333 14423 -287
rect 14469 -333 14547 -287
rect 14593 -333 14671 -287
rect 14717 -333 14795 -287
rect 14841 -333 14919 -287
rect 14965 -333 15043 -287
rect 15089 -333 15167 -287
rect 15213 -333 15291 -287
rect 15337 -333 15415 -287
rect 15461 -333 15539 -287
rect 15585 -333 15663 -287
rect 15709 -333 15787 -287
rect 15833 -333 15911 -287
rect 15957 -333 16035 -287
rect 16081 -333 16159 -287
rect 16205 -333 16283 -287
rect 16329 -333 16407 -287
rect 16453 -333 16531 -287
rect 16577 -333 16655 -287
rect 16701 -333 16779 -287
rect 16825 -333 16903 -287
rect 16949 -333 17027 -287
rect 17073 -333 17151 -287
rect 17197 -333 17275 -287
rect 17321 -333 17332 -287
rect -17332 -411 17332 -333
rect -17332 -457 -17321 -411
rect -17275 -457 -17197 -411
rect -17151 -457 -17073 -411
rect -17027 -457 -16949 -411
rect -16903 -457 -16825 -411
rect -16779 -457 -16701 -411
rect -16655 -457 -16577 -411
rect -16531 -457 -16453 -411
rect -16407 -457 -16329 -411
rect -16283 -457 -16205 -411
rect -16159 -457 -16081 -411
rect -16035 -457 -15957 -411
rect -15911 -457 -15833 -411
rect -15787 -457 -15709 -411
rect -15663 -457 -15585 -411
rect -15539 -457 -15461 -411
rect -15415 -457 -15337 -411
rect -15291 -457 -15213 -411
rect -15167 -457 -15089 -411
rect -15043 -457 -14965 -411
rect -14919 -457 -14841 -411
rect -14795 -457 -14717 -411
rect -14671 -457 -14593 -411
rect -14547 -457 -14469 -411
rect -14423 -457 -14345 -411
rect -14299 -457 -14221 -411
rect -14175 -457 -14097 -411
rect -14051 -457 -13973 -411
rect -13927 -457 -13849 -411
rect -13803 -457 -13725 -411
rect -13679 -457 -13601 -411
rect -13555 -457 -13477 -411
rect -13431 -457 -13353 -411
rect -13307 -457 -13229 -411
rect -13183 -457 -13105 -411
rect -13059 -457 -12981 -411
rect -12935 -457 -12857 -411
rect -12811 -457 -12733 -411
rect -12687 -457 -12609 -411
rect -12563 -457 -12485 -411
rect -12439 -457 -12361 -411
rect -12315 -457 -12237 -411
rect -12191 -457 -12113 -411
rect -12067 -457 -11989 -411
rect -11943 -457 -11865 -411
rect -11819 -457 -11741 -411
rect -11695 -457 -11617 -411
rect -11571 -457 -11493 -411
rect -11447 -457 -11369 -411
rect -11323 -457 -11245 -411
rect -11199 -457 -11121 -411
rect -11075 -457 -10997 -411
rect -10951 -457 -10873 -411
rect -10827 -457 -10749 -411
rect -10703 -457 -10625 -411
rect -10579 -457 -10501 -411
rect -10455 -457 -10377 -411
rect -10331 -457 -10253 -411
rect -10207 -457 -10129 -411
rect -10083 -457 -10005 -411
rect -9959 -457 -9881 -411
rect -9835 -457 -9757 -411
rect -9711 -457 -9633 -411
rect -9587 -457 -9509 -411
rect -9463 -457 -9385 -411
rect -9339 -457 -9261 -411
rect -9215 -457 -9137 -411
rect -9091 -457 -9013 -411
rect -8967 -457 -8889 -411
rect -8843 -457 -8765 -411
rect -8719 -457 -8641 -411
rect -8595 -457 -8517 -411
rect -8471 -457 -8393 -411
rect -8347 -457 -8269 -411
rect -8223 -457 -8145 -411
rect -8099 -457 -8021 -411
rect -7975 -457 -7897 -411
rect -7851 -457 -7773 -411
rect -7727 -457 -7649 -411
rect -7603 -457 -7525 -411
rect -7479 -457 -7401 -411
rect -7355 -457 -7277 -411
rect -7231 -457 -7153 -411
rect -7107 -457 -7029 -411
rect -6983 -457 -6905 -411
rect -6859 -457 -6781 -411
rect -6735 -457 -6657 -411
rect -6611 -457 -6533 -411
rect -6487 -457 -6409 -411
rect -6363 -457 -6285 -411
rect -6239 -457 -6161 -411
rect -6115 -457 -6037 -411
rect -5991 -457 -5913 -411
rect -5867 -457 -5789 -411
rect -5743 -457 -5665 -411
rect -5619 -457 -5541 -411
rect -5495 -457 -5417 -411
rect -5371 -457 -5293 -411
rect -5247 -457 -5169 -411
rect -5123 -457 -5045 -411
rect -4999 -457 -4921 -411
rect -4875 -457 -4797 -411
rect -4751 -457 -4673 -411
rect -4627 -457 -4549 -411
rect -4503 -457 -4425 -411
rect -4379 -457 -4301 -411
rect -4255 -457 -4177 -411
rect -4131 -457 -4053 -411
rect -4007 -457 -3929 -411
rect -3883 -457 -3805 -411
rect -3759 -457 -3681 -411
rect -3635 -457 -3557 -411
rect -3511 -457 -3433 -411
rect -3387 -457 -3309 -411
rect -3263 -457 -3185 -411
rect -3139 -457 -3061 -411
rect -3015 -457 -2937 -411
rect -2891 -457 -2813 -411
rect -2767 -457 -2689 -411
rect -2643 -457 -2565 -411
rect -2519 -457 -2441 -411
rect -2395 -457 -2317 -411
rect -2271 -457 -2193 -411
rect -2147 -457 -2069 -411
rect -2023 -457 -1945 -411
rect -1899 -457 -1821 -411
rect -1775 -457 -1697 -411
rect -1651 -457 -1573 -411
rect -1527 -457 -1449 -411
rect -1403 -457 -1325 -411
rect -1279 -457 -1201 -411
rect -1155 -457 -1077 -411
rect -1031 -457 -953 -411
rect -907 -457 -829 -411
rect -783 -457 -705 -411
rect -659 -457 -581 -411
rect -535 -457 -457 -411
rect -411 -457 -333 -411
rect -287 -457 -209 -411
rect -163 -457 -85 -411
rect -39 -457 39 -411
rect 85 -457 163 -411
rect 209 -457 287 -411
rect 333 -457 411 -411
rect 457 -457 535 -411
rect 581 -457 659 -411
rect 705 -457 783 -411
rect 829 -457 907 -411
rect 953 -457 1031 -411
rect 1077 -457 1155 -411
rect 1201 -457 1279 -411
rect 1325 -457 1403 -411
rect 1449 -457 1527 -411
rect 1573 -457 1651 -411
rect 1697 -457 1775 -411
rect 1821 -457 1899 -411
rect 1945 -457 2023 -411
rect 2069 -457 2147 -411
rect 2193 -457 2271 -411
rect 2317 -457 2395 -411
rect 2441 -457 2519 -411
rect 2565 -457 2643 -411
rect 2689 -457 2767 -411
rect 2813 -457 2891 -411
rect 2937 -457 3015 -411
rect 3061 -457 3139 -411
rect 3185 -457 3263 -411
rect 3309 -457 3387 -411
rect 3433 -457 3511 -411
rect 3557 -457 3635 -411
rect 3681 -457 3759 -411
rect 3805 -457 3883 -411
rect 3929 -457 4007 -411
rect 4053 -457 4131 -411
rect 4177 -457 4255 -411
rect 4301 -457 4379 -411
rect 4425 -457 4503 -411
rect 4549 -457 4627 -411
rect 4673 -457 4751 -411
rect 4797 -457 4875 -411
rect 4921 -457 4999 -411
rect 5045 -457 5123 -411
rect 5169 -457 5247 -411
rect 5293 -457 5371 -411
rect 5417 -457 5495 -411
rect 5541 -457 5619 -411
rect 5665 -457 5743 -411
rect 5789 -457 5867 -411
rect 5913 -457 5991 -411
rect 6037 -457 6115 -411
rect 6161 -457 6239 -411
rect 6285 -457 6363 -411
rect 6409 -457 6487 -411
rect 6533 -457 6611 -411
rect 6657 -457 6735 -411
rect 6781 -457 6859 -411
rect 6905 -457 6983 -411
rect 7029 -457 7107 -411
rect 7153 -457 7231 -411
rect 7277 -457 7355 -411
rect 7401 -457 7479 -411
rect 7525 -457 7603 -411
rect 7649 -457 7727 -411
rect 7773 -457 7851 -411
rect 7897 -457 7975 -411
rect 8021 -457 8099 -411
rect 8145 -457 8223 -411
rect 8269 -457 8347 -411
rect 8393 -457 8471 -411
rect 8517 -457 8595 -411
rect 8641 -457 8719 -411
rect 8765 -457 8843 -411
rect 8889 -457 8967 -411
rect 9013 -457 9091 -411
rect 9137 -457 9215 -411
rect 9261 -457 9339 -411
rect 9385 -457 9463 -411
rect 9509 -457 9587 -411
rect 9633 -457 9711 -411
rect 9757 -457 9835 -411
rect 9881 -457 9959 -411
rect 10005 -457 10083 -411
rect 10129 -457 10207 -411
rect 10253 -457 10331 -411
rect 10377 -457 10455 -411
rect 10501 -457 10579 -411
rect 10625 -457 10703 -411
rect 10749 -457 10827 -411
rect 10873 -457 10951 -411
rect 10997 -457 11075 -411
rect 11121 -457 11199 -411
rect 11245 -457 11323 -411
rect 11369 -457 11447 -411
rect 11493 -457 11571 -411
rect 11617 -457 11695 -411
rect 11741 -457 11819 -411
rect 11865 -457 11943 -411
rect 11989 -457 12067 -411
rect 12113 -457 12191 -411
rect 12237 -457 12315 -411
rect 12361 -457 12439 -411
rect 12485 -457 12563 -411
rect 12609 -457 12687 -411
rect 12733 -457 12811 -411
rect 12857 -457 12935 -411
rect 12981 -457 13059 -411
rect 13105 -457 13183 -411
rect 13229 -457 13307 -411
rect 13353 -457 13431 -411
rect 13477 -457 13555 -411
rect 13601 -457 13679 -411
rect 13725 -457 13803 -411
rect 13849 -457 13927 -411
rect 13973 -457 14051 -411
rect 14097 -457 14175 -411
rect 14221 -457 14299 -411
rect 14345 -457 14423 -411
rect 14469 -457 14547 -411
rect 14593 -457 14671 -411
rect 14717 -457 14795 -411
rect 14841 -457 14919 -411
rect 14965 -457 15043 -411
rect 15089 -457 15167 -411
rect 15213 -457 15291 -411
rect 15337 -457 15415 -411
rect 15461 -457 15539 -411
rect 15585 -457 15663 -411
rect 15709 -457 15787 -411
rect 15833 -457 15911 -411
rect 15957 -457 16035 -411
rect 16081 -457 16159 -411
rect 16205 -457 16283 -411
rect 16329 -457 16407 -411
rect 16453 -457 16531 -411
rect 16577 -457 16655 -411
rect 16701 -457 16779 -411
rect 16825 -457 16903 -411
rect 16949 -457 17027 -411
rect 17073 -457 17151 -411
rect 17197 -457 17275 -411
rect 17321 -457 17332 -411
rect -17332 -535 17332 -457
rect -17332 -581 -17321 -535
rect -17275 -581 -17197 -535
rect -17151 -581 -17073 -535
rect -17027 -581 -16949 -535
rect -16903 -581 -16825 -535
rect -16779 -581 -16701 -535
rect -16655 -581 -16577 -535
rect -16531 -581 -16453 -535
rect -16407 -581 -16329 -535
rect -16283 -581 -16205 -535
rect -16159 -581 -16081 -535
rect -16035 -581 -15957 -535
rect -15911 -581 -15833 -535
rect -15787 -581 -15709 -535
rect -15663 -581 -15585 -535
rect -15539 -581 -15461 -535
rect -15415 -581 -15337 -535
rect -15291 -581 -15213 -535
rect -15167 -581 -15089 -535
rect -15043 -581 -14965 -535
rect -14919 -581 -14841 -535
rect -14795 -581 -14717 -535
rect -14671 -581 -14593 -535
rect -14547 -581 -14469 -535
rect -14423 -581 -14345 -535
rect -14299 -581 -14221 -535
rect -14175 -581 -14097 -535
rect -14051 -581 -13973 -535
rect -13927 -581 -13849 -535
rect -13803 -581 -13725 -535
rect -13679 -581 -13601 -535
rect -13555 -581 -13477 -535
rect -13431 -581 -13353 -535
rect -13307 -581 -13229 -535
rect -13183 -581 -13105 -535
rect -13059 -581 -12981 -535
rect -12935 -581 -12857 -535
rect -12811 -581 -12733 -535
rect -12687 -581 -12609 -535
rect -12563 -581 -12485 -535
rect -12439 -581 -12361 -535
rect -12315 -581 -12237 -535
rect -12191 -581 -12113 -535
rect -12067 -581 -11989 -535
rect -11943 -581 -11865 -535
rect -11819 -581 -11741 -535
rect -11695 -581 -11617 -535
rect -11571 -581 -11493 -535
rect -11447 -581 -11369 -535
rect -11323 -581 -11245 -535
rect -11199 -581 -11121 -535
rect -11075 -581 -10997 -535
rect -10951 -581 -10873 -535
rect -10827 -581 -10749 -535
rect -10703 -581 -10625 -535
rect -10579 -581 -10501 -535
rect -10455 -581 -10377 -535
rect -10331 -581 -10253 -535
rect -10207 -581 -10129 -535
rect -10083 -581 -10005 -535
rect -9959 -581 -9881 -535
rect -9835 -581 -9757 -535
rect -9711 -581 -9633 -535
rect -9587 -581 -9509 -535
rect -9463 -581 -9385 -535
rect -9339 -581 -9261 -535
rect -9215 -581 -9137 -535
rect -9091 -581 -9013 -535
rect -8967 -581 -8889 -535
rect -8843 -581 -8765 -535
rect -8719 -581 -8641 -535
rect -8595 -581 -8517 -535
rect -8471 -581 -8393 -535
rect -8347 -581 -8269 -535
rect -8223 -581 -8145 -535
rect -8099 -581 -8021 -535
rect -7975 -581 -7897 -535
rect -7851 -581 -7773 -535
rect -7727 -581 -7649 -535
rect -7603 -581 -7525 -535
rect -7479 -581 -7401 -535
rect -7355 -581 -7277 -535
rect -7231 -581 -7153 -535
rect -7107 -581 -7029 -535
rect -6983 -581 -6905 -535
rect -6859 -581 -6781 -535
rect -6735 -581 -6657 -535
rect -6611 -581 -6533 -535
rect -6487 -581 -6409 -535
rect -6363 -581 -6285 -535
rect -6239 -581 -6161 -535
rect -6115 -581 -6037 -535
rect -5991 -581 -5913 -535
rect -5867 -581 -5789 -535
rect -5743 -581 -5665 -535
rect -5619 -581 -5541 -535
rect -5495 -581 -5417 -535
rect -5371 -581 -5293 -535
rect -5247 -581 -5169 -535
rect -5123 -581 -5045 -535
rect -4999 -581 -4921 -535
rect -4875 -581 -4797 -535
rect -4751 -581 -4673 -535
rect -4627 -581 -4549 -535
rect -4503 -581 -4425 -535
rect -4379 -581 -4301 -535
rect -4255 -581 -4177 -535
rect -4131 -581 -4053 -535
rect -4007 -581 -3929 -535
rect -3883 -581 -3805 -535
rect -3759 -581 -3681 -535
rect -3635 -581 -3557 -535
rect -3511 -581 -3433 -535
rect -3387 -581 -3309 -535
rect -3263 -581 -3185 -535
rect -3139 -581 -3061 -535
rect -3015 -581 -2937 -535
rect -2891 -581 -2813 -535
rect -2767 -581 -2689 -535
rect -2643 -581 -2565 -535
rect -2519 -581 -2441 -535
rect -2395 -581 -2317 -535
rect -2271 -581 -2193 -535
rect -2147 -581 -2069 -535
rect -2023 -581 -1945 -535
rect -1899 -581 -1821 -535
rect -1775 -581 -1697 -535
rect -1651 -581 -1573 -535
rect -1527 -581 -1449 -535
rect -1403 -581 -1325 -535
rect -1279 -581 -1201 -535
rect -1155 -581 -1077 -535
rect -1031 -581 -953 -535
rect -907 -581 -829 -535
rect -783 -581 -705 -535
rect -659 -581 -581 -535
rect -535 -581 -457 -535
rect -411 -581 -333 -535
rect -287 -581 -209 -535
rect -163 -581 -85 -535
rect -39 -581 39 -535
rect 85 -581 163 -535
rect 209 -581 287 -535
rect 333 -581 411 -535
rect 457 -581 535 -535
rect 581 -581 659 -535
rect 705 -581 783 -535
rect 829 -581 907 -535
rect 953 -581 1031 -535
rect 1077 -581 1155 -535
rect 1201 -581 1279 -535
rect 1325 -581 1403 -535
rect 1449 -581 1527 -535
rect 1573 -581 1651 -535
rect 1697 -581 1775 -535
rect 1821 -581 1899 -535
rect 1945 -581 2023 -535
rect 2069 -581 2147 -535
rect 2193 -581 2271 -535
rect 2317 -581 2395 -535
rect 2441 -581 2519 -535
rect 2565 -581 2643 -535
rect 2689 -581 2767 -535
rect 2813 -581 2891 -535
rect 2937 -581 3015 -535
rect 3061 -581 3139 -535
rect 3185 -581 3263 -535
rect 3309 -581 3387 -535
rect 3433 -581 3511 -535
rect 3557 -581 3635 -535
rect 3681 -581 3759 -535
rect 3805 -581 3883 -535
rect 3929 -581 4007 -535
rect 4053 -581 4131 -535
rect 4177 -581 4255 -535
rect 4301 -581 4379 -535
rect 4425 -581 4503 -535
rect 4549 -581 4627 -535
rect 4673 -581 4751 -535
rect 4797 -581 4875 -535
rect 4921 -581 4999 -535
rect 5045 -581 5123 -535
rect 5169 -581 5247 -535
rect 5293 -581 5371 -535
rect 5417 -581 5495 -535
rect 5541 -581 5619 -535
rect 5665 -581 5743 -535
rect 5789 -581 5867 -535
rect 5913 -581 5991 -535
rect 6037 -581 6115 -535
rect 6161 -581 6239 -535
rect 6285 -581 6363 -535
rect 6409 -581 6487 -535
rect 6533 -581 6611 -535
rect 6657 -581 6735 -535
rect 6781 -581 6859 -535
rect 6905 -581 6983 -535
rect 7029 -581 7107 -535
rect 7153 -581 7231 -535
rect 7277 -581 7355 -535
rect 7401 -581 7479 -535
rect 7525 -581 7603 -535
rect 7649 -581 7727 -535
rect 7773 -581 7851 -535
rect 7897 -581 7975 -535
rect 8021 -581 8099 -535
rect 8145 -581 8223 -535
rect 8269 -581 8347 -535
rect 8393 -581 8471 -535
rect 8517 -581 8595 -535
rect 8641 -581 8719 -535
rect 8765 -581 8843 -535
rect 8889 -581 8967 -535
rect 9013 -581 9091 -535
rect 9137 -581 9215 -535
rect 9261 -581 9339 -535
rect 9385 -581 9463 -535
rect 9509 -581 9587 -535
rect 9633 -581 9711 -535
rect 9757 -581 9835 -535
rect 9881 -581 9959 -535
rect 10005 -581 10083 -535
rect 10129 -581 10207 -535
rect 10253 -581 10331 -535
rect 10377 -581 10455 -535
rect 10501 -581 10579 -535
rect 10625 -581 10703 -535
rect 10749 -581 10827 -535
rect 10873 -581 10951 -535
rect 10997 -581 11075 -535
rect 11121 -581 11199 -535
rect 11245 -581 11323 -535
rect 11369 -581 11447 -535
rect 11493 -581 11571 -535
rect 11617 -581 11695 -535
rect 11741 -581 11819 -535
rect 11865 -581 11943 -535
rect 11989 -581 12067 -535
rect 12113 -581 12191 -535
rect 12237 -581 12315 -535
rect 12361 -581 12439 -535
rect 12485 -581 12563 -535
rect 12609 -581 12687 -535
rect 12733 -581 12811 -535
rect 12857 -581 12935 -535
rect 12981 -581 13059 -535
rect 13105 -581 13183 -535
rect 13229 -581 13307 -535
rect 13353 -581 13431 -535
rect 13477 -581 13555 -535
rect 13601 -581 13679 -535
rect 13725 -581 13803 -535
rect 13849 -581 13927 -535
rect 13973 -581 14051 -535
rect 14097 -581 14175 -535
rect 14221 -581 14299 -535
rect 14345 -581 14423 -535
rect 14469 -581 14547 -535
rect 14593 -581 14671 -535
rect 14717 -581 14795 -535
rect 14841 -581 14919 -535
rect 14965 -581 15043 -535
rect 15089 -581 15167 -535
rect 15213 -581 15291 -535
rect 15337 -581 15415 -535
rect 15461 -581 15539 -535
rect 15585 -581 15663 -535
rect 15709 -581 15787 -535
rect 15833 -581 15911 -535
rect 15957 -581 16035 -535
rect 16081 -581 16159 -535
rect 16205 -581 16283 -535
rect 16329 -581 16407 -535
rect 16453 -581 16531 -535
rect 16577 -581 16655 -535
rect 16701 -581 16779 -535
rect 16825 -581 16903 -535
rect 16949 -581 17027 -535
rect 17073 -581 17151 -535
rect 17197 -581 17275 -535
rect 17321 -581 17332 -535
rect -17332 -659 17332 -581
rect -17332 -705 -17321 -659
rect -17275 -705 -17197 -659
rect -17151 -705 -17073 -659
rect -17027 -705 -16949 -659
rect -16903 -705 -16825 -659
rect -16779 -705 -16701 -659
rect -16655 -705 -16577 -659
rect -16531 -705 -16453 -659
rect -16407 -705 -16329 -659
rect -16283 -705 -16205 -659
rect -16159 -705 -16081 -659
rect -16035 -705 -15957 -659
rect -15911 -705 -15833 -659
rect -15787 -705 -15709 -659
rect -15663 -705 -15585 -659
rect -15539 -705 -15461 -659
rect -15415 -705 -15337 -659
rect -15291 -705 -15213 -659
rect -15167 -705 -15089 -659
rect -15043 -705 -14965 -659
rect -14919 -705 -14841 -659
rect -14795 -705 -14717 -659
rect -14671 -705 -14593 -659
rect -14547 -705 -14469 -659
rect -14423 -705 -14345 -659
rect -14299 -705 -14221 -659
rect -14175 -705 -14097 -659
rect -14051 -705 -13973 -659
rect -13927 -705 -13849 -659
rect -13803 -705 -13725 -659
rect -13679 -705 -13601 -659
rect -13555 -705 -13477 -659
rect -13431 -705 -13353 -659
rect -13307 -705 -13229 -659
rect -13183 -705 -13105 -659
rect -13059 -705 -12981 -659
rect -12935 -705 -12857 -659
rect -12811 -705 -12733 -659
rect -12687 -705 -12609 -659
rect -12563 -705 -12485 -659
rect -12439 -705 -12361 -659
rect -12315 -705 -12237 -659
rect -12191 -705 -12113 -659
rect -12067 -705 -11989 -659
rect -11943 -705 -11865 -659
rect -11819 -705 -11741 -659
rect -11695 -705 -11617 -659
rect -11571 -705 -11493 -659
rect -11447 -705 -11369 -659
rect -11323 -705 -11245 -659
rect -11199 -705 -11121 -659
rect -11075 -705 -10997 -659
rect -10951 -705 -10873 -659
rect -10827 -705 -10749 -659
rect -10703 -705 -10625 -659
rect -10579 -705 -10501 -659
rect -10455 -705 -10377 -659
rect -10331 -705 -10253 -659
rect -10207 -705 -10129 -659
rect -10083 -705 -10005 -659
rect -9959 -705 -9881 -659
rect -9835 -705 -9757 -659
rect -9711 -705 -9633 -659
rect -9587 -705 -9509 -659
rect -9463 -705 -9385 -659
rect -9339 -705 -9261 -659
rect -9215 -705 -9137 -659
rect -9091 -705 -9013 -659
rect -8967 -705 -8889 -659
rect -8843 -705 -8765 -659
rect -8719 -705 -8641 -659
rect -8595 -705 -8517 -659
rect -8471 -705 -8393 -659
rect -8347 -705 -8269 -659
rect -8223 -705 -8145 -659
rect -8099 -705 -8021 -659
rect -7975 -705 -7897 -659
rect -7851 -705 -7773 -659
rect -7727 -705 -7649 -659
rect -7603 -705 -7525 -659
rect -7479 -705 -7401 -659
rect -7355 -705 -7277 -659
rect -7231 -705 -7153 -659
rect -7107 -705 -7029 -659
rect -6983 -705 -6905 -659
rect -6859 -705 -6781 -659
rect -6735 -705 -6657 -659
rect -6611 -705 -6533 -659
rect -6487 -705 -6409 -659
rect -6363 -705 -6285 -659
rect -6239 -705 -6161 -659
rect -6115 -705 -6037 -659
rect -5991 -705 -5913 -659
rect -5867 -705 -5789 -659
rect -5743 -705 -5665 -659
rect -5619 -705 -5541 -659
rect -5495 -705 -5417 -659
rect -5371 -705 -5293 -659
rect -5247 -705 -5169 -659
rect -5123 -705 -5045 -659
rect -4999 -705 -4921 -659
rect -4875 -705 -4797 -659
rect -4751 -705 -4673 -659
rect -4627 -705 -4549 -659
rect -4503 -705 -4425 -659
rect -4379 -705 -4301 -659
rect -4255 -705 -4177 -659
rect -4131 -705 -4053 -659
rect -4007 -705 -3929 -659
rect -3883 -705 -3805 -659
rect -3759 -705 -3681 -659
rect -3635 -705 -3557 -659
rect -3511 -705 -3433 -659
rect -3387 -705 -3309 -659
rect -3263 -705 -3185 -659
rect -3139 -705 -3061 -659
rect -3015 -705 -2937 -659
rect -2891 -705 -2813 -659
rect -2767 -705 -2689 -659
rect -2643 -705 -2565 -659
rect -2519 -705 -2441 -659
rect -2395 -705 -2317 -659
rect -2271 -705 -2193 -659
rect -2147 -705 -2069 -659
rect -2023 -705 -1945 -659
rect -1899 -705 -1821 -659
rect -1775 -705 -1697 -659
rect -1651 -705 -1573 -659
rect -1527 -705 -1449 -659
rect -1403 -705 -1325 -659
rect -1279 -705 -1201 -659
rect -1155 -705 -1077 -659
rect -1031 -705 -953 -659
rect -907 -705 -829 -659
rect -783 -705 -705 -659
rect -659 -705 -581 -659
rect -535 -705 -457 -659
rect -411 -705 -333 -659
rect -287 -705 -209 -659
rect -163 -705 -85 -659
rect -39 -705 39 -659
rect 85 -705 163 -659
rect 209 -705 287 -659
rect 333 -705 411 -659
rect 457 -705 535 -659
rect 581 -705 659 -659
rect 705 -705 783 -659
rect 829 -705 907 -659
rect 953 -705 1031 -659
rect 1077 -705 1155 -659
rect 1201 -705 1279 -659
rect 1325 -705 1403 -659
rect 1449 -705 1527 -659
rect 1573 -705 1651 -659
rect 1697 -705 1775 -659
rect 1821 -705 1899 -659
rect 1945 -705 2023 -659
rect 2069 -705 2147 -659
rect 2193 -705 2271 -659
rect 2317 -705 2395 -659
rect 2441 -705 2519 -659
rect 2565 -705 2643 -659
rect 2689 -705 2767 -659
rect 2813 -705 2891 -659
rect 2937 -705 3015 -659
rect 3061 -705 3139 -659
rect 3185 -705 3263 -659
rect 3309 -705 3387 -659
rect 3433 -705 3511 -659
rect 3557 -705 3635 -659
rect 3681 -705 3759 -659
rect 3805 -705 3883 -659
rect 3929 -705 4007 -659
rect 4053 -705 4131 -659
rect 4177 -705 4255 -659
rect 4301 -705 4379 -659
rect 4425 -705 4503 -659
rect 4549 -705 4627 -659
rect 4673 -705 4751 -659
rect 4797 -705 4875 -659
rect 4921 -705 4999 -659
rect 5045 -705 5123 -659
rect 5169 -705 5247 -659
rect 5293 -705 5371 -659
rect 5417 -705 5495 -659
rect 5541 -705 5619 -659
rect 5665 -705 5743 -659
rect 5789 -705 5867 -659
rect 5913 -705 5991 -659
rect 6037 -705 6115 -659
rect 6161 -705 6239 -659
rect 6285 -705 6363 -659
rect 6409 -705 6487 -659
rect 6533 -705 6611 -659
rect 6657 -705 6735 -659
rect 6781 -705 6859 -659
rect 6905 -705 6983 -659
rect 7029 -705 7107 -659
rect 7153 -705 7231 -659
rect 7277 -705 7355 -659
rect 7401 -705 7479 -659
rect 7525 -705 7603 -659
rect 7649 -705 7727 -659
rect 7773 -705 7851 -659
rect 7897 -705 7975 -659
rect 8021 -705 8099 -659
rect 8145 -705 8223 -659
rect 8269 -705 8347 -659
rect 8393 -705 8471 -659
rect 8517 -705 8595 -659
rect 8641 -705 8719 -659
rect 8765 -705 8843 -659
rect 8889 -705 8967 -659
rect 9013 -705 9091 -659
rect 9137 -705 9215 -659
rect 9261 -705 9339 -659
rect 9385 -705 9463 -659
rect 9509 -705 9587 -659
rect 9633 -705 9711 -659
rect 9757 -705 9835 -659
rect 9881 -705 9959 -659
rect 10005 -705 10083 -659
rect 10129 -705 10207 -659
rect 10253 -705 10331 -659
rect 10377 -705 10455 -659
rect 10501 -705 10579 -659
rect 10625 -705 10703 -659
rect 10749 -705 10827 -659
rect 10873 -705 10951 -659
rect 10997 -705 11075 -659
rect 11121 -705 11199 -659
rect 11245 -705 11323 -659
rect 11369 -705 11447 -659
rect 11493 -705 11571 -659
rect 11617 -705 11695 -659
rect 11741 -705 11819 -659
rect 11865 -705 11943 -659
rect 11989 -705 12067 -659
rect 12113 -705 12191 -659
rect 12237 -705 12315 -659
rect 12361 -705 12439 -659
rect 12485 -705 12563 -659
rect 12609 -705 12687 -659
rect 12733 -705 12811 -659
rect 12857 -705 12935 -659
rect 12981 -705 13059 -659
rect 13105 -705 13183 -659
rect 13229 -705 13307 -659
rect 13353 -705 13431 -659
rect 13477 -705 13555 -659
rect 13601 -705 13679 -659
rect 13725 -705 13803 -659
rect 13849 -705 13927 -659
rect 13973 -705 14051 -659
rect 14097 -705 14175 -659
rect 14221 -705 14299 -659
rect 14345 -705 14423 -659
rect 14469 -705 14547 -659
rect 14593 -705 14671 -659
rect 14717 -705 14795 -659
rect 14841 -705 14919 -659
rect 14965 -705 15043 -659
rect 15089 -705 15167 -659
rect 15213 -705 15291 -659
rect 15337 -705 15415 -659
rect 15461 -705 15539 -659
rect 15585 -705 15663 -659
rect 15709 -705 15787 -659
rect 15833 -705 15911 -659
rect 15957 -705 16035 -659
rect 16081 -705 16159 -659
rect 16205 -705 16283 -659
rect 16329 -705 16407 -659
rect 16453 -705 16531 -659
rect 16577 -705 16655 -659
rect 16701 -705 16779 -659
rect 16825 -705 16903 -659
rect 16949 -705 17027 -659
rect 17073 -705 17151 -659
rect 17197 -705 17275 -659
rect 17321 -705 17332 -659
rect -17332 -783 17332 -705
rect -17332 -829 -17321 -783
rect -17275 -829 -17197 -783
rect -17151 -829 -17073 -783
rect -17027 -829 -16949 -783
rect -16903 -829 -16825 -783
rect -16779 -829 -16701 -783
rect -16655 -829 -16577 -783
rect -16531 -829 -16453 -783
rect -16407 -829 -16329 -783
rect -16283 -829 -16205 -783
rect -16159 -829 -16081 -783
rect -16035 -829 -15957 -783
rect -15911 -829 -15833 -783
rect -15787 -829 -15709 -783
rect -15663 -829 -15585 -783
rect -15539 -829 -15461 -783
rect -15415 -829 -15337 -783
rect -15291 -829 -15213 -783
rect -15167 -829 -15089 -783
rect -15043 -829 -14965 -783
rect -14919 -829 -14841 -783
rect -14795 -829 -14717 -783
rect -14671 -829 -14593 -783
rect -14547 -829 -14469 -783
rect -14423 -829 -14345 -783
rect -14299 -829 -14221 -783
rect -14175 -829 -14097 -783
rect -14051 -829 -13973 -783
rect -13927 -829 -13849 -783
rect -13803 -829 -13725 -783
rect -13679 -829 -13601 -783
rect -13555 -829 -13477 -783
rect -13431 -829 -13353 -783
rect -13307 -829 -13229 -783
rect -13183 -829 -13105 -783
rect -13059 -829 -12981 -783
rect -12935 -829 -12857 -783
rect -12811 -829 -12733 -783
rect -12687 -829 -12609 -783
rect -12563 -829 -12485 -783
rect -12439 -829 -12361 -783
rect -12315 -829 -12237 -783
rect -12191 -829 -12113 -783
rect -12067 -829 -11989 -783
rect -11943 -829 -11865 -783
rect -11819 -829 -11741 -783
rect -11695 -829 -11617 -783
rect -11571 -829 -11493 -783
rect -11447 -829 -11369 -783
rect -11323 -829 -11245 -783
rect -11199 -829 -11121 -783
rect -11075 -829 -10997 -783
rect -10951 -829 -10873 -783
rect -10827 -829 -10749 -783
rect -10703 -829 -10625 -783
rect -10579 -829 -10501 -783
rect -10455 -829 -10377 -783
rect -10331 -829 -10253 -783
rect -10207 -829 -10129 -783
rect -10083 -829 -10005 -783
rect -9959 -829 -9881 -783
rect -9835 -829 -9757 -783
rect -9711 -829 -9633 -783
rect -9587 -829 -9509 -783
rect -9463 -829 -9385 -783
rect -9339 -829 -9261 -783
rect -9215 -829 -9137 -783
rect -9091 -829 -9013 -783
rect -8967 -829 -8889 -783
rect -8843 -829 -8765 -783
rect -8719 -829 -8641 -783
rect -8595 -829 -8517 -783
rect -8471 -829 -8393 -783
rect -8347 -829 -8269 -783
rect -8223 -829 -8145 -783
rect -8099 -829 -8021 -783
rect -7975 -829 -7897 -783
rect -7851 -829 -7773 -783
rect -7727 -829 -7649 -783
rect -7603 -829 -7525 -783
rect -7479 -829 -7401 -783
rect -7355 -829 -7277 -783
rect -7231 -829 -7153 -783
rect -7107 -829 -7029 -783
rect -6983 -829 -6905 -783
rect -6859 -829 -6781 -783
rect -6735 -829 -6657 -783
rect -6611 -829 -6533 -783
rect -6487 -829 -6409 -783
rect -6363 -829 -6285 -783
rect -6239 -829 -6161 -783
rect -6115 -829 -6037 -783
rect -5991 -829 -5913 -783
rect -5867 -829 -5789 -783
rect -5743 -829 -5665 -783
rect -5619 -829 -5541 -783
rect -5495 -829 -5417 -783
rect -5371 -829 -5293 -783
rect -5247 -829 -5169 -783
rect -5123 -829 -5045 -783
rect -4999 -829 -4921 -783
rect -4875 -829 -4797 -783
rect -4751 -829 -4673 -783
rect -4627 -829 -4549 -783
rect -4503 -829 -4425 -783
rect -4379 -829 -4301 -783
rect -4255 -829 -4177 -783
rect -4131 -829 -4053 -783
rect -4007 -829 -3929 -783
rect -3883 -829 -3805 -783
rect -3759 -829 -3681 -783
rect -3635 -829 -3557 -783
rect -3511 -829 -3433 -783
rect -3387 -829 -3309 -783
rect -3263 -829 -3185 -783
rect -3139 -829 -3061 -783
rect -3015 -829 -2937 -783
rect -2891 -829 -2813 -783
rect -2767 -829 -2689 -783
rect -2643 -829 -2565 -783
rect -2519 -829 -2441 -783
rect -2395 -829 -2317 -783
rect -2271 -829 -2193 -783
rect -2147 -829 -2069 -783
rect -2023 -829 -1945 -783
rect -1899 -829 -1821 -783
rect -1775 -829 -1697 -783
rect -1651 -829 -1573 -783
rect -1527 -829 -1449 -783
rect -1403 -829 -1325 -783
rect -1279 -829 -1201 -783
rect -1155 -829 -1077 -783
rect -1031 -829 -953 -783
rect -907 -829 -829 -783
rect -783 -829 -705 -783
rect -659 -829 -581 -783
rect -535 -829 -457 -783
rect -411 -829 -333 -783
rect -287 -829 -209 -783
rect -163 -829 -85 -783
rect -39 -829 39 -783
rect 85 -829 163 -783
rect 209 -829 287 -783
rect 333 -829 411 -783
rect 457 -829 535 -783
rect 581 -829 659 -783
rect 705 -829 783 -783
rect 829 -829 907 -783
rect 953 -829 1031 -783
rect 1077 -829 1155 -783
rect 1201 -829 1279 -783
rect 1325 -829 1403 -783
rect 1449 -829 1527 -783
rect 1573 -829 1651 -783
rect 1697 -829 1775 -783
rect 1821 -829 1899 -783
rect 1945 -829 2023 -783
rect 2069 -829 2147 -783
rect 2193 -829 2271 -783
rect 2317 -829 2395 -783
rect 2441 -829 2519 -783
rect 2565 -829 2643 -783
rect 2689 -829 2767 -783
rect 2813 -829 2891 -783
rect 2937 -829 3015 -783
rect 3061 -829 3139 -783
rect 3185 -829 3263 -783
rect 3309 -829 3387 -783
rect 3433 -829 3511 -783
rect 3557 -829 3635 -783
rect 3681 -829 3759 -783
rect 3805 -829 3883 -783
rect 3929 -829 4007 -783
rect 4053 -829 4131 -783
rect 4177 -829 4255 -783
rect 4301 -829 4379 -783
rect 4425 -829 4503 -783
rect 4549 -829 4627 -783
rect 4673 -829 4751 -783
rect 4797 -829 4875 -783
rect 4921 -829 4999 -783
rect 5045 -829 5123 -783
rect 5169 -829 5247 -783
rect 5293 -829 5371 -783
rect 5417 -829 5495 -783
rect 5541 -829 5619 -783
rect 5665 -829 5743 -783
rect 5789 -829 5867 -783
rect 5913 -829 5991 -783
rect 6037 -829 6115 -783
rect 6161 -829 6239 -783
rect 6285 -829 6363 -783
rect 6409 -829 6487 -783
rect 6533 -829 6611 -783
rect 6657 -829 6735 -783
rect 6781 -829 6859 -783
rect 6905 -829 6983 -783
rect 7029 -829 7107 -783
rect 7153 -829 7231 -783
rect 7277 -829 7355 -783
rect 7401 -829 7479 -783
rect 7525 -829 7603 -783
rect 7649 -829 7727 -783
rect 7773 -829 7851 -783
rect 7897 -829 7975 -783
rect 8021 -829 8099 -783
rect 8145 -829 8223 -783
rect 8269 -829 8347 -783
rect 8393 -829 8471 -783
rect 8517 -829 8595 -783
rect 8641 -829 8719 -783
rect 8765 -829 8843 -783
rect 8889 -829 8967 -783
rect 9013 -829 9091 -783
rect 9137 -829 9215 -783
rect 9261 -829 9339 -783
rect 9385 -829 9463 -783
rect 9509 -829 9587 -783
rect 9633 -829 9711 -783
rect 9757 -829 9835 -783
rect 9881 -829 9959 -783
rect 10005 -829 10083 -783
rect 10129 -829 10207 -783
rect 10253 -829 10331 -783
rect 10377 -829 10455 -783
rect 10501 -829 10579 -783
rect 10625 -829 10703 -783
rect 10749 -829 10827 -783
rect 10873 -829 10951 -783
rect 10997 -829 11075 -783
rect 11121 -829 11199 -783
rect 11245 -829 11323 -783
rect 11369 -829 11447 -783
rect 11493 -829 11571 -783
rect 11617 -829 11695 -783
rect 11741 -829 11819 -783
rect 11865 -829 11943 -783
rect 11989 -829 12067 -783
rect 12113 -829 12191 -783
rect 12237 -829 12315 -783
rect 12361 -829 12439 -783
rect 12485 -829 12563 -783
rect 12609 -829 12687 -783
rect 12733 -829 12811 -783
rect 12857 -829 12935 -783
rect 12981 -829 13059 -783
rect 13105 -829 13183 -783
rect 13229 -829 13307 -783
rect 13353 -829 13431 -783
rect 13477 -829 13555 -783
rect 13601 -829 13679 -783
rect 13725 -829 13803 -783
rect 13849 -829 13927 -783
rect 13973 -829 14051 -783
rect 14097 -829 14175 -783
rect 14221 -829 14299 -783
rect 14345 -829 14423 -783
rect 14469 -829 14547 -783
rect 14593 -829 14671 -783
rect 14717 -829 14795 -783
rect 14841 -829 14919 -783
rect 14965 -829 15043 -783
rect 15089 -829 15167 -783
rect 15213 -829 15291 -783
rect 15337 -829 15415 -783
rect 15461 -829 15539 -783
rect 15585 -829 15663 -783
rect 15709 -829 15787 -783
rect 15833 -829 15911 -783
rect 15957 -829 16035 -783
rect 16081 -829 16159 -783
rect 16205 -829 16283 -783
rect 16329 -829 16407 -783
rect 16453 -829 16531 -783
rect 16577 -829 16655 -783
rect 16701 -829 16779 -783
rect 16825 -829 16903 -783
rect 16949 -829 17027 -783
rect 17073 -829 17151 -783
rect 17197 -829 17275 -783
rect 17321 -829 17332 -783
rect -17332 -907 17332 -829
rect -17332 -953 -17321 -907
rect -17275 -953 -17197 -907
rect -17151 -953 -17073 -907
rect -17027 -953 -16949 -907
rect -16903 -953 -16825 -907
rect -16779 -953 -16701 -907
rect -16655 -953 -16577 -907
rect -16531 -953 -16453 -907
rect -16407 -953 -16329 -907
rect -16283 -953 -16205 -907
rect -16159 -953 -16081 -907
rect -16035 -953 -15957 -907
rect -15911 -953 -15833 -907
rect -15787 -953 -15709 -907
rect -15663 -953 -15585 -907
rect -15539 -953 -15461 -907
rect -15415 -953 -15337 -907
rect -15291 -953 -15213 -907
rect -15167 -953 -15089 -907
rect -15043 -953 -14965 -907
rect -14919 -953 -14841 -907
rect -14795 -953 -14717 -907
rect -14671 -953 -14593 -907
rect -14547 -953 -14469 -907
rect -14423 -953 -14345 -907
rect -14299 -953 -14221 -907
rect -14175 -953 -14097 -907
rect -14051 -953 -13973 -907
rect -13927 -953 -13849 -907
rect -13803 -953 -13725 -907
rect -13679 -953 -13601 -907
rect -13555 -953 -13477 -907
rect -13431 -953 -13353 -907
rect -13307 -953 -13229 -907
rect -13183 -953 -13105 -907
rect -13059 -953 -12981 -907
rect -12935 -953 -12857 -907
rect -12811 -953 -12733 -907
rect -12687 -953 -12609 -907
rect -12563 -953 -12485 -907
rect -12439 -953 -12361 -907
rect -12315 -953 -12237 -907
rect -12191 -953 -12113 -907
rect -12067 -953 -11989 -907
rect -11943 -953 -11865 -907
rect -11819 -953 -11741 -907
rect -11695 -953 -11617 -907
rect -11571 -953 -11493 -907
rect -11447 -953 -11369 -907
rect -11323 -953 -11245 -907
rect -11199 -953 -11121 -907
rect -11075 -953 -10997 -907
rect -10951 -953 -10873 -907
rect -10827 -953 -10749 -907
rect -10703 -953 -10625 -907
rect -10579 -953 -10501 -907
rect -10455 -953 -10377 -907
rect -10331 -953 -10253 -907
rect -10207 -953 -10129 -907
rect -10083 -953 -10005 -907
rect -9959 -953 -9881 -907
rect -9835 -953 -9757 -907
rect -9711 -953 -9633 -907
rect -9587 -953 -9509 -907
rect -9463 -953 -9385 -907
rect -9339 -953 -9261 -907
rect -9215 -953 -9137 -907
rect -9091 -953 -9013 -907
rect -8967 -953 -8889 -907
rect -8843 -953 -8765 -907
rect -8719 -953 -8641 -907
rect -8595 -953 -8517 -907
rect -8471 -953 -8393 -907
rect -8347 -953 -8269 -907
rect -8223 -953 -8145 -907
rect -8099 -953 -8021 -907
rect -7975 -953 -7897 -907
rect -7851 -953 -7773 -907
rect -7727 -953 -7649 -907
rect -7603 -953 -7525 -907
rect -7479 -953 -7401 -907
rect -7355 -953 -7277 -907
rect -7231 -953 -7153 -907
rect -7107 -953 -7029 -907
rect -6983 -953 -6905 -907
rect -6859 -953 -6781 -907
rect -6735 -953 -6657 -907
rect -6611 -953 -6533 -907
rect -6487 -953 -6409 -907
rect -6363 -953 -6285 -907
rect -6239 -953 -6161 -907
rect -6115 -953 -6037 -907
rect -5991 -953 -5913 -907
rect -5867 -953 -5789 -907
rect -5743 -953 -5665 -907
rect -5619 -953 -5541 -907
rect -5495 -953 -5417 -907
rect -5371 -953 -5293 -907
rect -5247 -953 -5169 -907
rect -5123 -953 -5045 -907
rect -4999 -953 -4921 -907
rect -4875 -953 -4797 -907
rect -4751 -953 -4673 -907
rect -4627 -953 -4549 -907
rect -4503 -953 -4425 -907
rect -4379 -953 -4301 -907
rect -4255 -953 -4177 -907
rect -4131 -953 -4053 -907
rect -4007 -953 -3929 -907
rect -3883 -953 -3805 -907
rect -3759 -953 -3681 -907
rect -3635 -953 -3557 -907
rect -3511 -953 -3433 -907
rect -3387 -953 -3309 -907
rect -3263 -953 -3185 -907
rect -3139 -953 -3061 -907
rect -3015 -953 -2937 -907
rect -2891 -953 -2813 -907
rect -2767 -953 -2689 -907
rect -2643 -953 -2565 -907
rect -2519 -953 -2441 -907
rect -2395 -953 -2317 -907
rect -2271 -953 -2193 -907
rect -2147 -953 -2069 -907
rect -2023 -953 -1945 -907
rect -1899 -953 -1821 -907
rect -1775 -953 -1697 -907
rect -1651 -953 -1573 -907
rect -1527 -953 -1449 -907
rect -1403 -953 -1325 -907
rect -1279 -953 -1201 -907
rect -1155 -953 -1077 -907
rect -1031 -953 -953 -907
rect -907 -953 -829 -907
rect -783 -953 -705 -907
rect -659 -953 -581 -907
rect -535 -953 -457 -907
rect -411 -953 -333 -907
rect -287 -953 -209 -907
rect -163 -953 -85 -907
rect -39 -953 39 -907
rect 85 -953 163 -907
rect 209 -953 287 -907
rect 333 -953 411 -907
rect 457 -953 535 -907
rect 581 -953 659 -907
rect 705 -953 783 -907
rect 829 -953 907 -907
rect 953 -953 1031 -907
rect 1077 -953 1155 -907
rect 1201 -953 1279 -907
rect 1325 -953 1403 -907
rect 1449 -953 1527 -907
rect 1573 -953 1651 -907
rect 1697 -953 1775 -907
rect 1821 -953 1899 -907
rect 1945 -953 2023 -907
rect 2069 -953 2147 -907
rect 2193 -953 2271 -907
rect 2317 -953 2395 -907
rect 2441 -953 2519 -907
rect 2565 -953 2643 -907
rect 2689 -953 2767 -907
rect 2813 -953 2891 -907
rect 2937 -953 3015 -907
rect 3061 -953 3139 -907
rect 3185 -953 3263 -907
rect 3309 -953 3387 -907
rect 3433 -953 3511 -907
rect 3557 -953 3635 -907
rect 3681 -953 3759 -907
rect 3805 -953 3883 -907
rect 3929 -953 4007 -907
rect 4053 -953 4131 -907
rect 4177 -953 4255 -907
rect 4301 -953 4379 -907
rect 4425 -953 4503 -907
rect 4549 -953 4627 -907
rect 4673 -953 4751 -907
rect 4797 -953 4875 -907
rect 4921 -953 4999 -907
rect 5045 -953 5123 -907
rect 5169 -953 5247 -907
rect 5293 -953 5371 -907
rect 5417 -953 5495 -907
rect 5541 -953 5619 -907
rect 5665 -953 5743 -907
rect 5789 -953 5867 -907
rect 5913 -953 5991 -907
rect 6037 -953 6115 -907
rect 6161 -953 6239 -907
rect 6285 -953 6363 -907
rect 6409 -953 6487 -907
rect 6533 -953 6611 -907
rect 6657 -953 6735 -907
rect 6781 -953 6859 -907
rect 6905 -953 6983 -907
rect 7029 -953 7107 -907
rect 7153 -953 7231 -907
rect 7277 -953 7355 -907
rect 7401 -953 7479 -907
rect 7525 -953 7603 -907
rect 7649 -953 7727 -907
rect 7773 -953 7851 -907
rect 7897 -953 7975 -907
rect 8021 -953 8099 -907
rect 8145 -953 8223 -907
rect 8269 -953 8347 -907
rect 8393 -953 8471 -907
rect 8517 -953 8595 -907
rect 8641 -953 8719 -907
rect 8765 -953 8843 -907
rect 8889 -953 8967 -907
rect 9013 -953 9091 -907
rect 9137 -953 9215 -907
rect 9261 -953 9339 -907
rect 9385 -953 9463 -907
rect 9509 -953 9587 -907
rect 9633 -953 9711 -907
rect 9757 -953 9835 -907
rect 9881 -953 9959 -907
rect 10005 -953 10083 -907
rect 10129 -953 10207 -907
rect 10253 -953 10331 -907
rect 10377 -953 10455 -907
rect 10501 -953 10579 -907
rect 10625 -953 10703 -907
rect 10749 -953 10827 -907
rect 10873 -953 10951 -907
rect 10997 -953 11075 -907
rect 11121 -953 11199 -907
rect 11245 -953 11323 -907
rect 11369 -953 11447 -907
rect 11493 -953 11571 -907
rect 11617 -953 11695 -907
rect 11741 -953 11819 -907
rect 11865 -953 11943 -907
rect 11989 -953 12067 -907
rect 12113 -953 12191 -907
rect 12237 -953 12315 -907
rect 12361 -953 12439 -907
rect 12485 -953 12563 -907
rect 12609 -953 12687 -907
rect 12733 -953 12811 -907
rect 12857 -953 12935 -907
rect 12981 -953 13059 -907
rect 13105 -953 13183 -907
rect 13229 -953 13307 -907
rect 13353 -953 13431 -907
rect 13477 -953 13555 -907
rect 13601 -953 13679 -907
rect 13725 -953 13803 -907
rect 13849 -953 13927 -907
rect 13973 -953 14051 -907
rect 14097 -953 14175 -907
rect 14221 -953 14299 -907
rect 14345 -953 14423 -907
rect 14469 -953 14547 -907
rect 14593 -953 14671 -907
rect 14717 -953 14795 -907
rect 14841 -953 14919 -907
rect 14965 -953 15043 -907
rect 15089 -953 15167 -907
rect 15213 -953 15291 -907
rect 15337 -953 15415 -907
rect 15461 -953 15539 -907
rect 15585 -953 15663 -907
rect 15709 -953 15787 -907
rect 15833 -953 15911 -907
rect 15957 -953 16035 -907
rect 16081 -953 16159 -907
rect 16205 -953 16283 -907
rect 16329 -953 16407 -907
rect 16453 -953 16531 -907
rect 16577 -953 16655 -907
rect 16701 -953 16779 -907
rect 16825 -953 16903 -907
rect 16949 -953 17027 -907
rect 17073 -953 17151 -907
rect 17197 -953 17275 -907
rect 17321 -953 17332 -907
rect -17332 -964 17332 -953
<< end >>
