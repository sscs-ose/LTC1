** sch_path: /home/shahid/GF180Projects/Top_test/top/xschem/untitled-11.sch
**.subckt untitled-11
V1 VDD VSS 3.3
.save i(v1)
V2 VSS GND 0
.save i(v2)
V3 CLK VSS pulse(3.3 0 0 100p 100p 2.50n 5n)
.save i(v3)
C5 Vdiv VSS 10f m=1
V5 RST VSS PWL( 0 0 10n 0 10.001n 3)
.save i(v5)
V6 P1 VSS pulse(3.3 0 0 100p 100p 80n 160n)
.save i(v6)
V7 P0 VSS pulse(3.3 0 0 100p 100p 40n 80n)
.save i(v7)
x1 VSS VDD RST Vdiv P1 P0 CLK pex_Output_Divider_Mag
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.inlcude pex_Output_Divider_Mag.spice
.control
save all
tran 1n 200n
plot v(CLK) v(Vdiv)+3.5 v(RST)+7 v(P0)+10.5 v(P1)+14
**write Output_Divider_TB.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
