magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2208 -2120 3568 2820
<< nwell >>
rect -208 -120 1568 820
<< mvpmos >>
rect 0 0 140 700
rect 244 0 384 700
rect 488 0 628 700
rect 732 0 872 700
rect 976 0 1116 700
rect 1220 0 1360 700
<< mvpdiff >>
rect -88 687 0 700
rect -88 641 -75 687
rect -29 641 0 687
rect -88 583 0 641
rect -88 537 -75 583
rect -29 537 0 583
rect -88 479 0 537
rect -88 433 -75 479
rect -29 433 0 479
rect -88 374 0 433
rect -88 328 -75 374
rect -29 328 0 374
rect -88 269 0 328
rect -88 223 -75 269
rect -29 223 0 269
rect -88 164 0 223
rect -88 118 -75 164
rect -29 118 0 164
rect -88 59 0 118
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 140 687 244 700
rect 140 641 169 687
rect 215 641 244 687
rect 140 583 244 641
rect 140 537 169 583
rect 215 537 244 583
rect 140 479 244 537
rect 140 433 169 479
rect 215 433 244 479
rect 140 374 244 433
rect 140 328 169 374
rect 215 328 244 374
rect 140 269 244 328
rect 140 223 169 269
rect 215 223 244 269
rect 140 164 244 223
rect 140 118 169 164
rect 215 118 244 164
rect 140 59 244 118
rect 140 13 169 59
rect 215 13 244 59
rect 140 0 244 13
rect 384 687 488 700
rect 384 641 413 687
rect 459 641 488 687
rect 384 583 488 641
rect 384 537 413 583
rect 459 537 488 583
rect 384 479 488 537
rect 384 433 413 479
rect 459 433 488 479
rect 384 374 488 433
rect 384 328 413 374
rect 459 328 488 374
rect 384 269 488 328
rect 384 223 413 269
rect 459 223 488 269
rect 384 164 488 223
rect 384 118 413 164
rect 459 118 488 164
rect 384 59 488 118
rect 384 13 413 59
rect 459 13 488 59
rect 384 0 488 13
rect 628 687 732 700
rect 628 641 657 687
rect 703 641 732 687
rect 628 583 732 641
rect 628 537 657 583
rect 703 537 732 583
rect 628 479 732 537
rect 628 433 657 479
rect 703 433 732 479
rect 628 374 732 433
rect 628 328 657 374
rect 703 328 732 374
rect 628 269 732 328
rect 628 223 657 269
rect 703 223 732 269
rect 628 164 732 223
rect 628 118 657 164
rect 703 118 732 164
rect 628 59 732 118
rect 628 13 657 59
rect 703 13 732 59
rect 628 0 732 13
rect 872 687 976 700
rect 872 641 901 687
rect 947 641 976 687
rect 872 583 976 641
rect 872 537 901 583
rect 947 537 976 583
rect 872 479 976 537
rect 872 433 901 479
rect 947 433 976 479
rect 872 374 976 433
rect 872 328 901 374
rect 947 328 976 374
rect 872 269 976 328
rect 872 223 901 269
rect 947 223 976 269
rect 872 164 976 223
rect 872 118 901 164
rect 947 118 976 164
rect 872 59 976 118
rect 872 13 901 59
rect 947 13 976 59
rect 872 0 976 13
rect 1116 687 1220 700
rect 1116 641 1145 687
rect 1191 641 1220 687
rect 1116 583 1220 641
rect 1116 537 1145 583
rect 1191 537 1220 583
rect 1116 479 1220 537
rect 1116 433 1145 479
rect 1191 433 1220 479
rect 1116 374 1220 433
rect 1116 328 1145 374
rect 1191 328 1220 374
rect 1116 269 1220 328
rect 1116 223 1145 269
rect 1191 223 1220 269
rect 1116 164 1220 223
rect 1116 118 1145 164
rect 1191 118 1220 164
rect 1116 59 1220 118
rect 1116 13 1145 59
rect 1191 13 1220 59
rect 1116 0 1220 13
rect 1360 687 1448 700
rect 1360 641 1389 687
rect 1435 641 1448 687
rect 1360 583 1448 641
rect 1360 537 1389 583
rect 1435 537 1448 583
rect 1360 479 1448 537
rect 1360 433 1389 479
rect 1435 433 1448 479
rect 1360 374 1448 433
rect 1360 328 1389 374
rect 1435 328 1448 374
rect 1360 269 1448 328
rect 1360 223 1389 269
rect 1435 223 1448 269
rect 1360 164 1448 223
rect 1360 118 1389 164
rect 1435 118 1448 164
rect 1360 59 1448 118
rect 1360 13 1389 59
rect 1435 13 1448 59
rect 1360 0 1448 13
<< mvpdiffc >>
rect -75 641 -29 687
rect -75 537 -29 583
rect -75 433 -29 479
rect -75 328 -29 374
rect -75 223 -29 269
rect -75 118 -29 164
rect -75 13 -29 59
rect 169 641 215 687
rect 169 537 215 583
rect 169 433 215 479
rect 169 328 215 374
rect 169 223 215 269
rect 169 118 215 164
rect 169 13 215 59
rect 413 641 459 687
rect 413 537 459 583
rect 413 433 459 479
rect 413 328 459 374
rect 413 223 459 269
rect 413 118 459 164
rect 413 13 459 59
rect 657 641 703 687
rect 657 537 703 583
rect 657 433 703 479
rect 657 328 703 374
rect 657 223 703 269
rect 657 118 703 164
rect 657 13 703 59
rect 901 641 947 687
rect 901 537 947 583
rect 901 433 947 479
rect 901 328 947 374
rect 901 223 947 269
rect 901 118 947 164
rect 901 13 947 59
rect 1145 641 1191 687
rect 1145 537 1191 583
rect 1145 433 1191 479
rect 1145 328 1191 374
rect 1145 223 1191 269
rect 1145 118 1191 164
rect 1145 13 1191 59
rect 1389 641 1435 687
rect 1389 537 1435 583
rect 1389 433 1435 479
rect 1389 328 1435 374
rect 1389 223 1435 269
rect 1389 118 1435 164
rect 1389 13 1435 59
<< polysilicon >>
rect 0 700 140 744
rect 244 700 384 744
rect 488 700 628 744
rect 732 700 872 744
rect 976 700 1116 744
rect 1220 700 1360 744
rect 0 -44 140 0
rect 244 -44 384 0
rect 488 -44 628 0
rect 732 -44 872 0
rect 976 -44 1116 0
rect 1220 -44 1360 0
<< metal1 >>
rect -75 687 -29 700
rect -75 583 -29 641
rect -75 479 -29 537
rect -75 374 -29 433
rect -75 269 -29 328
rect -75 164 -29 223
rect -75 59 -29 118
rect -75 0 -29 13
rect 169 687 215 700
rect 169 583 215 641
rect 169 479 215 537
rect 169 374 215 433
rect 169 269 215 328
rect 169 164 215 223
rect 169 59 215 118
rect 169 0 215 13
rect 413 687 459 700
rect 413 583 459 641
rect 413 479 459 537
rect 413 374 459 433
rect 413 269 459 328
rect 413 164 459 223
rect 413 59 459 118
rect 413 0 459 13
rect 657 687 703 700
rect 657 583 703 641
rect 657 479 703 537
rect 657 374 703 433
rect 657 269 703 328
rect 657 164 703 223
rect 657 59 703 118
rect 657 0 703 13
rect 901 687 947 700
rect 901 583 947 641
rect 901 479 947 537
rect 901 374 947 433
rect 901 269 947 328
rect 901 164 947 223
rect 901 59 947 118
rect 901 0 947 13
rect 1145 687 1191 700
rect 1145 583 1191 641
rect 1145 479 1191 537
rect 1145 374 1191 433
rect 1145 269 1191 328
rect 1145 164 1191 223
rect 1145 59 1191 118
rect 1145 0 1191 13
rect 1389 687 1435 700
rect 1389 583 1435 641
rect 1389 479 1435 537
rect 1389 374 1435 433
rect 1389 269 1435 328
rect 1389 164 1435 223
rect 1389 59 1435 118
rect 1389 0 1435 13
<< labels >>
rlabel mvpdiffc 1168 350 1168 350 4 D
rlabel mvpdiffc 924 350 924 350 4 S
rlabel mvpdiffc 680 350 680 350 4 D
rlabel mvpdiffc 436 350 436 350 4 S
rlabel mvpdiffc 192 350 192 350 4 D
rlabel mvpdiffc 1412 350 1412 350 4 S
rlabel mvpdiffc -52 350 -52 350 4 S
<< end >>
