magic
tech gf180mcuC
magscale 1 10
timestamp 1711086265
<< nwell >>
rect -2726 -3062 2726 3062
<< nsubdiff >>
rect -2702 3025 2702 3038
rect -2702 2979 -2586 3025
rect 2586 2979 2702 3025
rect -2702 2966 2702 2979
rect -2702 2922 -2630 2966
rect -2702 -2922 -2689 2922
rect -2643 -2922 -2630 2922
rect 2630 2922 2702 2966
rect -2702 -2966 -2630 -2922
rect 2630 -2922 2643 2922
rect 2689 -2922 2702 2922
rect 2630 -2966 2702 -2922
rect -2702 -2979 2702 -2966
rect -2702 -3025 -2586 -2979
rect 2586 -3025 2702 -2979
rect -2702 -3038 2702 -3025
<< nsubdiffcont >>
rect -2586 2979 2586 3025
rect -2689 -2922 -2643 2922
rect 2643 -2922 2689 2922
rect -2586 -3025 2586 -2979
<< polysilicon >>
rect -2510 2833 -2290 2846
rect -2510 2787 -2497 2833
rect -2303 2787 -2290 2833
rect -2510 2744 -2290 2787
rect -2510 2181 -2290 2224
rect -2510 2135 -2497 2181
rect -2303 2135 -2290 2181
rect -2510 2122 -2290 2135
rect -2210 2833 -1990 2846
rect -2210 2787 -2197 2833
rect -2003 2787 -1990 2833
rect -2210 2744 -1990 2787
rect -2210 2181 -1990 2224
rect -2210 2135 -2197 2181
rect -2003 2135 -1990 2181
rect -2210 2122 -1990 2135
rect -1910 2833 -1690 2846
rect -1910 2787 -1897 2833
rect -1703 2787 -1690 2833
rect -1910 2744 -1690 2787
rect -1910 2181 -1690 2224
rect -1910 2135 -1897 2181
rect -1703 2135 -1690 2181
rect -1910 2122 -1690 2135
rect -1610 2833 -1390 2846
rect -1610 2787 -1597 2833
rect -1403 2787 -1390 2833
rect -1610 2744 -1390 2787
rect -1610 2181 -1390 2224
rect -1610 2135 -1597 2181
rect -1403 2135 -1390 2181
rect -1610 2122 -1390 2135
rect -1310 2833 -1090 2846
rect -1310 2787 -1297 2833
rect -1103 2787 -1090 2833
rect -1310 2744 -1090 2787
rect -1310 2181 -1090 2224
rect -1310 2135 -1297 2181
rect -1103 2135 -1090 2181
rect -1310 2122 -1090 2135
rect -1010 2833 -790 2846
rect -1010 2787 -997 2833
rect -803 2787 -790 2833
rect -1010 2744 -790 2787
rect -1010 2181 -790 2224
rect -1010 2135 -997 2181
rect -803 2135 -790 2181
rect -1010 2122 -790 2135
rect -710 2833 -490 2846
rect -710 2787 -697 2833
rect -503 2787 -490 2833
rect -710 2744 -490 2787
rect -710 2181 -490 2224
rect -710 2135 -697 2181
rect -503 2135 -490 2181
rect -710 2122 -490 2135
rect -410 2833 -190 2846
rect -410 2787 -397 2833
rect -203 2787 -190 2833
rect -410 2744 -190 2787
rect -410 2181 -190 2224
rect -410 2135 -397 2181
rect -203 2135 -190 2181
rect -410 2122 -190 2135
rect -110 2833 110 2846
rect -110 2787 -97 2833
rect 97 2787 110 2833
rect -110 2744 110 2787
rect -110 2181 110 2224
rect -110 2135 -97 2181
rect 97 2135 110 2181
rect -110 2122 110 2135
rect 190 2833 410 2846
rect 190 2787 203 2833
rect 397 2787 410 2833
rect 190 2744 410 2787
rect 190 2181 410 2224
rect 190 2135 203 2181
rect 397 2135 410 2181
rect 190 2122 410 2135
rect 490 2833 710 2846
rect 490 2787 503 2833
rect 697 2787 710 2833
rect 490 2744 710 2787
rect 490 2181 710 2224
rect 490 2135 503 2181
rect 697 2135 710 2181
rect 490 2122 710 2135
rect 790 2833 1010 2846
rect 790 2787 803 2833
rect 997 2787 1010 2833
rect 790 2744 1010 2787
rect 790 2181 1010 2224
rect 790 2135 803 2181
rect 997 2135 1010 2181
rect 790 2122 1010 2135
rect 1090 2833 1310 2846
rect 1090 2787 1103 2833
rect 1297 2787 1310 2833
rect 1090 2744 1310 2787
rect 1090 2181 1310 2224
rect 1090 2135 1103 2181
rect 1297 2135 1310 2181
rect 1090 2122 1310 2135
rect 1390 2833 1610 2846
rect 1390 2787 1403 2833
rect 1597 2787 1610 2833
rect 1390 2744 1610 2787
rect 1390 2181 1610 2224
rect 1390 2135 1403 2181
rect 1597 2135 1610 2181
rect 1390 2122 1610 2135
rect 1690 2833 1910 2846
rect 1690 2787 1703 2833
rect 1897 2787 1910 2833
rect 1690 2744 1910 2787
rect 1690 2181 1910 2224
rect 1690 2135 1703 2181
rect 1897 2135 1910 2181
rect 1690 2122 1910 2135
rect 1990 2833 2210 2846
rect 1990 2787 2003 2833
rect 2197 2787 2210 2833
rect 1990 2744 2210 2787
rect 1990 2181 2210 2224
rect 1990 2135 2003 2181
rect 2197 2135 2210 2181
rect 1990 2122 2210 2135
rect 2290 2833 2510 2846
rect 2290 2787 2303 2833
rect 2497 2787 2510 2833
rect 2290 2744 2510 2787
rect 2290 2181 2510 2224
rect 2290 2135 2303 2181
rect 2497 2135 2510 2181
rect 2290 2122 2510 2135
rect -2510 2005 -2290 2018
rect -2510 1959 -2497 2005
rect -2303 1959 -2290 2005
rect -2510 1916 -2290 1959
rect -2510 1353 -2290 1396
rect -2510 1307 -2497 1353
rect -2303 1307 -2290 1353
rect -2510 1294 -2290 1307
rect -2210 2005 -1990 2018
rect -2210 1959 -2197 2005
rect -2003 1959 -1990 2005
rect -2210 1916 -1990 1959
rect -2210 1353 -1990 1396
rect -2210 1307 -2197 1353
rect -2003 1307 -1990 1353
rect -2210 1294 -1990 1307
rect -1910 2005 -1690 2018
rect -1910 1959 -1897 2005
rect -1703 1959 -1690 2005
rect -1910 1916 -1690 1959
rect -1910 1353 -1690 1396
rect -1910 1307 -1897 1353
rect -1703 1307 -1690 1353
rect -1910 1294 -1690 1307
rect -1610 2005 -1390 2018
rect -1610 1959 -1597 2005
rect -1403 1959 -1390 2005
rect -1610 1916 -1390 1959
rect -1610 1353 -1390 1396
rect -1610 1307 -1597 1353
rect -1403 1307 -1390 1353
rect -1610 1294 -1390 1307
rect -1310 2005 -1090 2018
rect -1310 1959 -1297 2005
rect -1103 1959 -1090 2005
rect -1310 1916 -1090 1959
rect -1310 1353 -1090 1396
rect -1310 1307 -1297 1353
rect -1103 1307 -1090 1353
rect -1310 1294 -1090 1307
rect -1010 2005 -790 2018
rect -1010 1959 -997 2005
rect -803 1959 -790 2005
rect -1010 1916 -790 1959
rect -1010 1353 -790 1396
rect -1010 1307 -997 1353
rect -803 1307 -790 1353
rect -1010 1294 -790 1307
rect -710 2005 -490 2018
rect -710 1959 -697 2005
rect -503 1959 -490 2005
rect -710 1916 -490 1959
rect -710 1353 -490 1396
rect -710 1307 -697 1353
rect -503 1307 -490 1353
rect -710 1294 -490 1307
rect -410 2005 -190 2018
rect -410 1959 -397 2005
rect -203 1959 -190 2005
rect -410 1916 -190 1959
rect -410 1353 -190 1396
rect -410 1307 -397 1353
rect -203 1307 -190 1353
rect -410 1294 -190 1307
rect -110 2005 110 2018
rect -110 1959 -97 2005
rect 97 1959 110 2005
rect -110 1916 110 1959
rect -110 1353 110 1396
rect -110 1307 -97 1353
rect 97 1307 110 1353
rect -110 1294 110 1307
rect 190 2005 410 2018
rect 190 1959 203 2005
rect 397 1959 410 2005
rect 190 1916 410 1959
rect 190 1353 410 1396
rect 190 1307 203 1353
rect 397 1307 410 1353
rect 190 1294 410 1307
rect 490 2005 710 2018
rect 490 1959 503 2005
rect 697 1959 710 2005
rect 490 1916 710 1959
rect 490 1353 710 1396
rect 490 1307 503 1353
rect 697 1307 710 1353
rect 490 1294 710 1307
rect 790 2005 1010 2018
rect 790 1959 803 2005
rect 997 1959 1010 2005
rect 790 1916 1010 1959
rect 790 1353 1010 1396
rect 790 1307 803 1353
rect 997 1307 1010 1353
rect 790 1294 1010 1307
rect 1090 2005 1310 2018
rect 1090 1959 1103 2005
rect 1297 1959 1310 2005
rect 1090 1916 1310 1959
rect 1090 1353 1310 1396
rect 1090 1307 1103 1353
rect 1297 1307 1310 1353
rect 1090 1294 1310 1307
rect 1390 2005 1610 2018
rect 1390 1959 1403 2005
rect 1597 1959 1610 2005
rect 1390 1916 1610 1959
rect 1390 1353 1610 1396
rect 1390 1307 1403 1353
rect 1597 1307 1610 1353
rect 1390 1294 1610 1307
rect 1690 2005 1910 2018
rect 1690 1959 1703 2005
rect 1897 1959 1910 2005
rect 1690 1916 1910 1959
rect 1690 1353 1910 1396
rect 1690 1307 1703 1353
rect 1897 1307 1910 1353
rect 1690 1294 1910 1307
rect 1990 2005 2210 2018
rect 1990 1959 2003 2005
rect 2197 1959 2210 2005
rect 1990 1916 2210 1959
rect 1990 1353 2210 1396
rect 1990 1307 2003 1353
rect 2197 1307 2210 1353
rect 1990 1294 2210 1307
rect 2290 2005 2510 2018
rect 2290 1959 2303 2005
rect 2497 1959 2510 2005
rect 2290 1916 2510 1959
rect 2290 1353 2510 1396
rect 2290 1307 2303 1353
rect 2497 1307 2510 1353
rect 2290 1294 2510 1307
rect -2510 1177 -2290 1190
rect -2510 1131 -2497 1177
rect -2303 1131 -2290 1177
rect -2510 1088 -2290 1131
rect -2510 525 -2290 568
rect -2510 479 -2497 525
rect -2303 479 -2290 525
rect -2510 466 -2290 479
rect -2210 1177 -1990 1190
rect -2210 1131 -2197 1177
rect -2003 1131 -1990 1177
rect -2210 1088 -1990 1131
rect -2210 525 -1990 568
rect -2210 479 -2197 525
rect -2003 479 -1990 525
rect -2210 466 -1990 479
rect -1910 1177 -1690 1190
rect -1910 1131 -1897 1177
rect -1703 1131 -1690 1177
rect -1910 1088 -1690 1131
rect -1910 525 -1690 568
rect -1910 479 -1897 525
rect -1703 479 -1690 525
rect -1910 466 -1690 479
rect -1610 1177 -1390 1190
rect -1610 1131 -1597 1177
rect -1403 1131 -1390 1177
rect -1610 1088 -1390 1131
rect -1610 525 -1390 568
rect -1610 479 -1597 525
rect -1403 479 -1390 525
rect -1610 466 -1390 479
rect -1310 1177 -1090 1190
rect -1310 1131 -1297 1177
rect -1103 1131 -1090 1177
rect -1310 1088 -1090 1131
rect -1310 525 -1090 568
rect -1310 479 -1297 525
rect -1103 479 -1090 525
rect -1310 466 -1090 479
rect -1010 1177 -790 1190
rect -1010 1131 -997 1177
rect -803 1131 -790 1177
rect -1010 1088 -790 1131
rect -1010 525 -790 568
rect -1010 479 -997 525
rect -803 479 -790 525
rect -1010 466 -790 479
rect -710 1177 -490 1190
rect -710 1131 -697 1177
rect -503 1131 -490 1177
rect -710 1088 -490 1131
rect -710 525 -490 568
rect -710 479 -697 525
rect -503 479 -490 525
rect -710 466 -490 479
rect -410 1177 -190 1190
rect -410 1131 -397 1177
rect -203 1131 -190 1177
rect -410 1088 -190 1131
rect -410 525 -190 568
rect -410 479 -397 525
rect -203 479 -190 525
rect -410 466 -190 479
rect -110 1177 110 1190
rect -110 1131 -97 1177
rect 97 1131 110 1177
rect -110 1088 110 1131
rect -110 525 110 568
rect -110 479 -97 525
rect 97 479 110 525
rect -110 466 110 479
rect 190 1177 410 1190
rect 190 1131 203 1177
rect 397 1131 410 1177
rect 190 1088 410 1131
rect 190 525 410 568
rect 190 479 203 525
rect 397 479 410 525
rect 190 466 410 479
rect 490 1177 710 1190
rect 490 1131 503 1177
rect 697 1131 710 1177
rect 490 1088 710 1131
rect 490 525 710 568
rect 490 479 503 525
rect 697 479 710 525
rect 490 466 710 479
rect 790 1177 1010 1190
rect 790 1131 803 1177
rect 997 1131 1010 1177
rect 790 1088 1010 1131
rect 790 525 1010 568
rect 790 479 803 525
rect 997 479 1010 525
rect 790 466 1010 479
rect 1090 1177 1310 1190
rect 1090 1131 1103 1177
rect 1297 1131 1310 1177
rect 1090 1088 1310 1131
rect 1090 525 1310 568
rect 1090 479 1103 525
rect 1297 479 1310 525
rect 1090 466 1310 479
rect 1390 1177 1610 1190
rect 1390 1131 1403 1177
rect 1597 1131 1610 1177
rect 1390 1088 1610 1131
rect 1390 525 1610 568
rect 1390 479 1403 525
rect 1597 479 1610 525
rect 1390 466 1610 479
rect 1690 1177 1910 1190
rect 1690 1131 1703 1177
rect 1897 1131 1910 1177
rect 1690 1088 1910 1131
rect 1690 525 1910 568
rect 1690 479 1703 525
rect 1897 479 1910 525
rect 1690 466 1910 479
rect 1990 1177 2210 1190
rect 1990 1131 2003 1177
rect 2197 1131 2210 1177
rect 1990 1088 2210 1131
rect 1990 525 2210 568
rect 1990 479 2003 525
rect 2197 479 2210 525
rect 1990 466 2210 479
rect 2290 1177 2510 1190
rect 2290 1131 2303 1177
rect 2497 1131 2510 1177
rect 2290 1088 2510 1131
rect 2290 525 2510 568
rect 2290 479 2303 525
rect 2497 479 2510 525
rect 2290 466 2510 479
rect -2510 349 -2290 362
rect -2510 303 -2497 349
rect -2303 303 -2290 349
rect -2510 260 -2290 303
rect -2510 -303 -2290 -260
rect -2510 -349 -2497 -303
rect -2303 -349 -2290 -303
rect -2510 -362 -2290 -349
rect -2210 349 -1990 362
rect -2210 303 -2197 349
rect -2003 303 -1990 349
rect -2210 260 -1990 303
rect -2210 -303 -1990 -260
rect -2210 -349 -2197 -303
rect -2003 -349 -1990 -303
rect -2210 -362 -1990 -349
rect -1910 349 -1690 362
rect -1910 303 -1897 349
rect -1703 303 -1690 349
rect -1910 260 -1690 303
rect -1910 -303 -1690 -260
rect -1910 -349 -1897 -303
rect -1703 -349 -1690 -303
rect -1910 -362 -1690 -349
rect -1610 349 -1390 362
rect -1610 303 -1597 349
rect -1403 303 -1390 349
rect -1610 260 -1390 303
rect -1610 -303 -1390 -260
rect -1610 -349 -1597 -303
rect -1403 -349 -1390 -303
rect -1610 -362 -1390 -349
rect -1310 349 -1090 362
rect -1310 303 -1297 349
rect -1103 303 -1090 349
rect -1310 260 -1090 303
rect -1310 -303 -1090 -260
rect -1310 -349 -1297 -303
rect -1103 -349 -1090 -303
rect -1310 -362 -1090 -349
rect -1010 349 -790 362
rect -1010 303 -997 349
rect -803 303 -790 349
rect -1010 260 -790 303
rect -1010 -303 -790 -260
rect -1010 -349 -997 -303
rect -803 -349 -790 -303
rect -1010 -362 -790 -349
rect -710 349 -490 362
rect -710 303 -697 349
rect -503 303 -490 349
rect -710 260 -490 303
rect -710 -303 -490 -260
rect -710 -349 -697 -303
rect -503 -349 -490 -303
rect -710 -362 -490 -349
rect -410 349 -190 362
rect -410 303 -397 349
rect -203 303 -190 349
rect -410 260 -190 303
rect -410 -303 -190 -260
rect -410 -349 -397 -303
rect -203 -349 -190 -303
rect -410 -362 -190 -349
rect -110 349 110 362
rect -110 303 -97 349
rect 97 303 110 349
rect -110 260 110 303
rect -110 -303 110 -260
rect -110 -349 -97 -303
rect 97 -349 110 -303
rect -110 -362 110 -349
rect 190 349 410 362
rect 190 303 203 349
rect 397 303 410 349
rect 190 260 410 303
rect 190 -303 410 -260
rect 190 -349 203 -303
rect 397 -349 410 -303
rect 190 -362 410 -349
rect 490 349 710 362
rect 490 303 503 349
rect 697 303 710 349
rect 490 260 710 303
rect 490 -303 710 -260
rect 490 -349 503 -303
rect 697 -349 710 -303
rect 490 -362 710 -349
rect 790 349 1010 362
rect 790 303 803 349
rect 997 303 1010 349
rect 790 260 1010 303
rect 790 -303 1010 -260
rect 790 -349 803 -303
rect 997 -349 1010 -303
rect 790 -362 1010 -349
rect 1090 349 1310 362
rect 1090 303 1103 349
rect 1297 303 1310 349
rect 1090 260 1310 303
rect 1090 -303 1310 -260
rect 1090 -349 1103 -303
rect 1297 -349 1310 -303
rect 1090 -362 1310 -349
rect 1390 349 1610 362
rect 1390 303 1403 349
rect 1597 303 1610 349
rect 1390 260 1610 303
rect 1390 -303 1610 -260
rect 1390 -349 1403 -303
rect 1597 -349 1610 -303
rect 1390 -362 1610 -349
rect 1690 349 1910 362
rect 1690 303 1703 349
rect 1897 303 1910 349
rect 1690 260 1910 303
rect 1690 -303 1910 -260
rect 1690 -349 1703 -303
rect 1897 -349 1910 -303
rect 1690 -362 1910 -349
rect 1990 349 2210 362
rect 1990 303 2003 349
rect 2197 303 2210 349
rect 1990 260 2210 303
rect 1990 -303 2210 -260
rect 1990 -349 2003 -303
rect 2197 -349 2210 -303
rect 1990 -362 2210 -349
rect 2290 349 2510 362
rect 2290 303 2303 349
rect 2497 303 2510 349
rect 2290 260 2510 303
rect 2290 -303 2510 -260
rect 2290 -349 2303 -303
rect 2497 -349 2510 -303
rect 2290 -362 2510 -349
rect -2510 -479 -2290 -466
rect -2510 -525 -2497 -479
rect -2303 -525 -2290 -479
rect -2510 -568 -2290 -525
rect -2510 -1131 -2290 -1088
rect -2510 -1177 -2497 -1131
rect -2303 -1177 -2290 -1131
rect -2510 -1190 -2290 -1177
rect -2210 -479 -1990 -466
rect -2210 -525 -2197 -479
rect -2003 -525 -1990 -479
rect -2210 -568 -1990 -525
rect -2210 -1131 -1990 -1088
rect -2210 -1177 -2197 -1131
rect -2003 -1177 -1990 -1131
rect -2210 -1190 -1990 -1177
rect -1910 -479 -1690 -466
rect -1910 -525 -1897 -479
rect -1703 -525 -1690 -479
rect -1910 -568 -1690 -525
rect -1910 -1131 -1690 -1088
rect -1910 -1177 -1897 -1131
rect -1703 -1177 -1690 -1131
rect -1910 -1190 -1690 -1177
rect -1610 -479 -1390 -466
rect -1610 -525 -1597 -479
rect -1403 -525 -1390 -479
rect -1610 -568 -1390 -525
rect -1610 -1131 -1390 -1088
rect -1610 -1177 -1597 -1131
rect -1403 -1177 -1390 -1131
rect -1610 -1190 -1390 -1177
rect -1310 -479 -1090 -466
rect -1310 -525 -1297 -479
rect -1103 -525 -1090 -479
rect -1310 -568 -1090 -525
rect -1310 -1131 -1090 -1088
rect -1310 -1177 -1297 -1131
rect -1103 -1177 -1090 -1131
rect -1310 -1190 -1090 -1177
rect -1010 -479 -790 -466
rect -1010 -525 -997 -479
rect -803 -525 -790 -479
rect -1010 -568 -790 -525
rect -1010 -1131 -790 -1088
rect -1010 -1177 -997 -1131
rect -803 -1177 -790 -1131
rect -1010 -1190 -790 -1177
rect -710 -479 -490 -466
rect -710 -525 -697 -479
rect -503 -525 -490 -479
rect -710 -568 -490 -525
rect -710 -1131 -490 -1088
rect -710 -1177 -697 -1131
rect -503 -1177 -490 -1131
rect -710 -1190 -490 -1177
rect -410 -479 -190 -466
rect -410 -525 -397 -479
rect -203 -525 -190 -479
rect -410 -568 -190 -525
rect -410 -1131 -190 -1088
rect -410 -1177 -397 -1131
rect -203 -1177 -190 -1131
rect -410 -1190 -190 -1177
rect -110 -479 110 -466
rect -110 -525 -97 -479
rect 97 -525 110 -479
rect -110 -568 110 -525
rect -110 -1131 110 -1088
rect -110 -1177 -97 -1131
rect 97 -1177 110 -1131
rect -110 -1190 110 -1177
rect 190 -479 410 -466
rect 190 -525 203 -479
rect 397 -525 410 -479
rect 190 -568 410 -525
rect 190 -1131 410 -1088
rect 190 -1177 203 -1131
rect 397 -1177 410 -1131
rect 190 -1190 410 -1177
rect 490 -479 710 -466
rect 490 -525 503 -479
rect 697 -525 710 -479
rect 490 -568 710 -525
rect 490 -1131 710 -1088
rect 490 -1177 503 -1131
rect 697 -1177 710 -1131
rect 490 -1190 710 -1177
rect 790 -479 1010 -466
rect 790 -525 803 -479
rect 997 -525 1010 -479
rect 790 -568 1010 -525
rect 790 -1131 1010 -1088
rect 790 -1177 803 -1131
rect 997 -1177 1010 -1131
rect 790 -1190 1010 -1177
rect 1090 -479 1310 -466
rect 1090 -525 1103 -479
rect 1297 -525 1310 -479
rect 1090 -568 1310 -525
rect 1090 -1131 1310 -1088
rect 1090 -1177 1103 -1131
rect 1297 -1177 1310 -1131
rect 1090 -1190 1310 -1177
rect 1390 -479 1610 -466
rect 1390 -525 1403 -479
rect 1597 -525 1610 -479
rect 1390 -568 1610 -525
rect 1390 -1131 1610 -1088
rect 1390 -1177 1403 -1131
rect 1597 -1177 1610 -1131
rect 1390 -1190 1610 -1177
rect 1690 -479 1910 -466
rect 1690 -525 1703 -479
rect 1897 -525 1910 -479
rect 1690 -568 1910 -525
rect 1690 -1131 1910 -1088
rect 1690 -1177 1703 -1131
rect 1897 -1177 1910 -1131
rect 1690 -1190 1910 -1177
rect 1990 -479 2210 -466
rect 1990 -525 2003 -479
rect 2197 -525 2210 -479
rect 1990 -568 2210 -525
rect 1990 -1131 2210 -1088
rect 1990 -1177 2003 -1131
rect 2197 -1177 2210 -1131
rect 1990 -1190 2210 -1177
rect 2290 -479 2510 -466
rect 2290 -525 2303 -479
rect 2497 -525 2510 -479
rect 2290 -568 2510 -525
rect 2290 -1131 2510 -1088
rect 2290 -1177 2303 -1131
rect 2497 -1177 2510 -1131
rect 2290 -1190 2510 -1177
rect -2510 -1307 -2290 -1294
rect -2510 -1353 -2497 -1307
rect -2303 -1353 -2290 -1307
rect -2510 -1396 -2290 -1353
rect -2510 -1959 -2290 -1916
rect -2510 -2005 -2497 -1959
rect -2303 -2005 -2290 -1959
rect -2510 -2018 -2290 -2005
rect -2210 -1307 -1990 -1294
rect -2210 -1353 -2197 -1307
rect -2003 -1353 -1990 -1307
rect -2210 -1396 -1990 -1353
rect -2210 -1959 -1990 -1916
rect -2210 -2005 -2197 -1959
rect -2003 -2005 -1990 -1959
rect -2210 -2018 -1990 -2005
rect -1910 -1307 -1690 -1294
rect -1910 -1353 -1897 -1307
rect -1703 -1353 -1690 -1307
rect -1910 -1396 -1690 -1353
rect -1910 -1959 -1690 -1916
rect -1910 -2005 -1897 -1959
rect -1703 -2005 -1690 -1959
rect -1910 -2018 -1690 -2005
rect -1610 -1307 -1390 -1294
rect -1610 -1353 -1597 -1307
rect -1403 -1353 -1390 -1307
rect -1610 -1396 -1390 -1353
rect -1610 -1959 -1390 -1916
rect -1610 -2005 -1597 -1959
rect -1403 -2005 -1390 -1959
rect -1610 -2018 -1390 -2005
rect -1310 -1307 -1090 -1294
rect -1310 -1353 -1297 -1307
rect -1103 -1353 -1090 -1307
rect -1310 -1396 -1090 -1353
rect -1310 -1959 -1090 -1916
rect -1310 -2005 -1297 -1959
rect -1103 -2005 -1090 -1959
rect -1310 -2018 -1090 -2005
rect -1010 -1307 -790 -1294
rect -1010 -1353 -997 -1307
rect -803 -1353 -790 -1307
rect -1010 -1396 -790 -1353
rect -1010 -1959 -790 -1916
rect -1010 -2005 -997 -1959
rect -803 -2005 -790 -1959
rect -1010 -2018 -790 -2005
rect -710 -1307 -490 -1294
rect -710 -1353 -697 -1307
rect -503 -1353 -490 -1307
rect -710 -1396 -490 -1353
rect -710 -1959 -490 -1916
rect -710 -2005 -697 -1959
rect -503 -2005 -490 -1959
rect -710 -2018 -490 -2005
rect -410 -1307 -190 -1294
rect -410 -1353 -397 -1307
rect -203 -1353 -190 -1307
rect -410 -1396 -190 -1353
rect -410 -1959 -190 -1916
rect -410 -2005 -397 -1959
rect -203 -2005 -190 -1959
rect -410 -2018 -190 -2005
rect -110 -1307 110 -1294
rect -110 -1353 -97 -1307
rect 97 -1353 110 -1307
rect -110 -1396 110 -1353
rect -110 -1959 110 -1916
rect -110 -2005 -97 -1959
rect 97 -2005 110 -1959
rect -110 -2018 110 -2005
rect 190 -1307 410 -1294
rect 190 -1353 203 -1307
rect 397 -1353 410 -1307
rect 190 -1396 410 -1353
rect 190 -1959 410 -1916
rect 190 -2005 203 -1959
rect 397 -2005 410 -1959
rect 190 -2018 410 -2005
rect 490 -1307 710 -1294
rect 490 -1353 503 -1307
rect 697 -1353 710 -1307
rect 490 -1396 710 -1353
rect 490 -1959 710 -1916
rect 490 -2005 503 -1959
rect 697 -2005 710 -1959
rect 490 -2018 710 -2005
rect 790 -1307 1010 -1294
rect 790 -1353 803 -1307
rect 997 -1353 1010 -1307
rect 790 -1396 1010 -1353
rect 790 -1959 1010 -1916
rect 790 -2005 803 -1959
rect 997 -2005 1010 -1959
rect 790 -2018 1010 -2005
rect 1090 -1307 1310 -1294
rect 1090 -1353 1103 -1307
rect 1297 -1353 1310 -1307
rect 1090 -1396 1310 -1353
rect 1090 -1959 1310 -1916
rect 1090 -2005 1103 -1959
rect 1297 -2005 1310 -1959
rect 1090 -2018 1310 -2005
rect 1390 -1307 1610 -1294
rect 1390 -1353 1403 -1307
rect 1597 -1353 1610 -1307
rect 1390 -1396 1610 -1353
rect 1390 -1959 1610 -1916
rect 1390 -2005 1403 -1959
rect 1597 -2005 1610 -1959
rect 1390 -2018 1610 -2005
rect 1690 -1307 1910 -1294
rect 1690 -1353 1703 -1307
rect 1897 -1353 1910 -1307
rect 1690 -1396 1910 -1353
rect 1690 -1959 1910 -1916
rect 1690 -2005 1703 -1959
rect 1897 -2005 1910 -1959
rect 1690 -2018 1910 -2005
rect 1990 -1307 2210 -1294
rect 1990 -1353 2003 -1307
rect 2197 -1353 2210 -1307
rect 1990 -1396 2210 -1353
rect 1990 -1959 2210 -1916
rect 1990 -2005 2003 -1959
rect 2197 -2005 2210 -1959
rect 1990 -2018 2210 -2005
rect 2290 -1307 2510 -1294
rect 2290 -1353 2303 -1307
rect 2497 -1353 2510 -1307
rect 2290 -1396 2510 -1353
rect 2290 -1959 2510 -1916
rect 2290 -2005 2303 -1959
rect 2497 -2005 2510 -1959
rect 2290 -2018 2510 -2005
rect -2510 -2135 -2290 -2122
rect -2510 -2181 -2497 -2135
rect -2303 -2181 -2290 -2135
rect -2510 -2224 -2290 -2181
rect -2510 -2787 -2290 -2744
rect -2510 -2833 -2497 -2787
rect -2303 -2833 -2290 -2787
rect -2510 -2846 -2290 -2833
rect -2210 -2135 -1990 -2122
rect -2210 -2181 -2197 -2135
rect -2003 -2181 -1990 -2135
rect -2210 -2224 -1990 -2181
rect -2210 -2787 -1990 -2744
rect -2210 -2833 -2197 -2787
rect -2003 -2833 -1990 -2787
rect -2210 -2846 -1990 -2833
rect -1910 -2135 -1690 -2122
rect -1910 -2181 -1897 -2135
rect -1703 -2181 -1690 -2135
rect -1910 -2224 -1690 -2181
rect -1910 -2787 -1690 -2744
rect -1910 -2833 -1897 -2787
rect -1703 -2833 -1690 -2787
rect -1910 -2846 -1690 -2833
rect -1610 -2135 -1390 -2122
rect -1610 -2181 -1597 -2135
rect -1403 -2181 -1390 -2135
rect -1610 -2224 -1390 -2181
rect -1610 -2787 -1390 -2744
rect -1610 -2833 -1597 -2787
rect -1403 -2833 -1390 -2787
rect -1610 -2846 -1390 -2833
rect -1310 -2135 -1090 -2122
rect -1310 -2181 -1297 -2135
rect -1103 -2181 -1090 -2135
rect -1310 -2224 -1090 -2181
rect -1310 -2787 -1090 -2744
rect -1310 -2833 -1297 -2787
rect -1103 -2833 -1090 -2787
rect -1310 -2846 -1090 -2833
rect -1010 -2135 -790 -2122
rect -1010 -2181 -997 -2135
rect -803 -2181 -790 -2135
rect -1010 -2224 -790 -2181
rect -1010 -2787 -790 -2744
rect -1010 -2833 -997 -2787
rect -803 -2833 -790 -2787
rect -1010 -2846 -790 -2833
rect -710 -2135 -490 -2122
rect -710 -2181 -697 -2135
rect -503 -2181 -490 -2135
rect -710 -2224 -490 -2181
rect -710 -2787 -490 -2744
rect -710 -2833 -697 -2787
rect -503 -2833 -490 -2787
rect -710 -2846 -490 -2833
rect -410 -2135 -190 -2122
rect -410 -2181 -397 -2135
rect -203 -2181 -190 -2135
rect -410 -2224 -190 -2181
rect -410 -2787 -190 -2744
rect -410 -2833 -397 -2787
rect -203 -2833 -190 -2787
rect -410 -2846 -190 -2833
rect -110 -2135 110 -2122
rect -110 -2181 -97 -2135
rect 97 -2181 110 -2135
rect -110 -2224 110 -2181
rect -110 -2787 110 -2744
rect -110 -2833 -97 -2787
rect 97 -2833 110 -2787
rect -110 -2846 110 -2833
rect 190 -2135 410 -2122
rect 190 -2181 203 -2135
rect 397 -2181 410 -2135
rect 190 -2224 410 -2181
rect 190 -2787 410 -2744
rect 190 -2833 203 -2787
rect 397 -2833 410 -2787
rect 190 -2846 410 -2833
rect 490 -2135 710 -2122
rect 490 -2181 503 -2135
rect 697 -2181 710 -2135
rect 490 -2224 710 -2181
rect 490 -2787 710 -2744
rect 490 -2833 503 -2787
rect 697 -2833 710 -2787
rect 490 -2846 710 -2833
rect 790 -2135 1010 -2122
rect 790 -2181 803 -2135
rect 997 -2181 1010 -2135
rect 790 -2224 1010 -2181
rect 790 -2787 1010 -2744
rect 790 -2833 803 -2787
rect 997 -2833 1010 -2787
rect 790 -2846 1010 -2833
rect 1090 -2135 1310 -2122
rect 1090 -2181 1103 -2135
rect 1297 -2181 1310 -2135
rect 1090 -2224 1310 -2181
rect 1090 -2787 1310 -2744
rect 1090 -2833 1103 -2787
rect 1297 -2833 1310 -2787
rect 1090 -2846 1310 -2833
rect 1390 -2135 1610 -2122
rect 1390 -2181 1403 -2135
rect 1597 -2181 1610 -2135
rect 1390 -2224 1610 -2181
rect 1390 -2787 1610 -2744
rect 1390 -2833 1403 -2787
rect 1597 -2833 1610 -2787
rect 1390 -2846 1610 -2833
rect 1690 -2135 1910 -2122
rect 1690 -2181 1703 -2135
rect 1897 -2181 1910 -2135
rect 1690 -2224 1910 -2181
rect 1690 -2787 1910 -2744
rect 1690 -2833 1703 -2787
rect 1897 -2833 1910 -2787
rect 1690 -2846 1910 -2833
rect 1990 -2135 2210 -2122
rect 1990 -2181 2003 -2135
rect 2197 -2181 2210 -2135
rect 1990 -2224 2210 -2181
rect 1990 -2787 2210 -2744
rect 1990 -2833 2003 -2787
rect 2197 -2833 2210 -2787
rect 1990 -2846 2210 -2833
rect 2290 -2135 2510 -2122
rect 2290 -2181 2303 -2135
rect 2497 -2181 2510 -2135
rect 2290 -2224 2510 -2181
rect 2290 -2787 2510 -2744
rect 2290 -2833 2303 -2787
rect 2497 -2833 2510 -2787
rect 2290 -2846 2510 -2833
<< polycontact >>
rect -2497 2787 -2303 2833
rect -2497 2135 -2303 2181
rect -2197 2787 -2003 2833
rect -2197 2135 -2003 2181
rect -1897 2787 -1703 2833
rect -1897 2135 -1703 2181
rect -1597 2787 -1403 2833
rect -1597 2135 -1403 2181
rect -1297 2787 -1103 2833
rect -1297 2135 -1103 2181
rect -997 2787 -803 2833
rect -997 2135 -803 2181
rect -697 2787 -503 2833
rect -697 2135 -503 2181
rect -397 2787 -203 2833
rect -397 2135 -203 2181
rect -97 2787 97 2833
rect -97 2135 97 2181
rect 203 2787 397 2833
rect 203 2135 397 2181
rect 503 2787 697 2833
rect 503 2135 697 2181
rect 803 2787 997 2833
rect 803 2135 997 2181
rect 1103 2787 1297 2833
rect 1103 2135 1297 2181
rect 1403 2787 1597 2833
rect 1403 2135 1597 2181
rect 1703 2787 1897 2833
rect 1703 2135 1897 2181
rect 2003 2787 2197 2833
rect 2003 2135 2197 2181
rect 2303 2787 2497 2833
rect 2303 2135 2497 2181
rect -2497 1959 -2303 2005
rect -2497 1307 -2303 1353
rect -2197 1959 -2003 2005
rect -2197 1307 -2003 1353
rect -1897 1959 -1703 2005
rect -1897 1307 -1703 1353
rect -1597 1959 -1403 2005
rect -1597 1307 -1403 1353
rect -1297 1959 -1103 2005
rect -1297 1307 -1103 1353
rect -997 1959 -803 2005
rect -997 1307 -803 1353
rect -697 1959 -503 2005
rect -697 1307 -503 1353
rect -397 1959 -203 2005
rect -397 1307 -203 1353
rect -97 1959 97 2005
rect -97 1307 97 1353
rect 203 1959 397 2005
rect 203 1307 397 1353
rect 503 1959 697 2005
rect 503 1307 697 1353
rect 803 1959 997 2005
rect 803 1307 997 1353
rect 1103 1959 1297 2005
rect 1103 1307 1297 1353
rect 1403 1959 1597 2005
rect 1403 1307 1597 1353
rect 1703 1959 1897 2005
rect 1703 1307 1897 1353
rect 2003 1959 2197 2005
rect 2003 1307 2197 1353
rect 2303 1959 2497 2005
rect 2303 1307 2497 1353
rect -2497 1131 -2303 1177
rect -2497 479 -2303 525
rect -2197 1131 -2003 1177
rect -2197 479 -2003 525
rect -1897 1131 -1703 1177
rect -1897 479 -1703 525
rect -1597 1131 -1403 1177
rect -1597 479 -1403 525
rect -1297 1131 -1103 1177
rect -1297 479 -1103 525
rect -997 1131 -803 1177
rect -997 479 -803 525
rect -697 1131 -503 1177
rect -697 479 -503 525
rect -397 1131 -203 1177
rect -397 479 -203 525
rect -97 1131 97 1177
rect -97 479 97 525
rect 203 1131 397 1177
rect 203 479 397 525
rect 503 1131 697 1177
rect 503 479 697 525
rect 803 1131 997 1177
rect 803 479 997 525
rect 1103 1131 1297 1177
rect 1103 479 1297 525
rect 1403 1131 1597 1177
rect 1403 479 1597 525
rect 1703 1131 1897 1177
rect 1703 479 1897 525
rect 2003 1131 2197 1177
rect 2003 479 2197 525
rect 2303 1131 2497 1177
rect 2303 479 2497 525
rect -2497 303 -2303 349
rect -2497 -349 -2303 -303
rect -2197 303 -2003 349
rect -2197 -349 -2003 -303
rect -1897 303 -1703 349
rect -1897 -349 -1703 -303
rect -1597 303 -1403 349
rect -1597 -349 -1403 -303
rect -1297 303 -1103 349
rect -1297 -349 -1103 -303
rect -997 303 -803 349
rect -997 -349 -803 -303
rect -697 303 -503 349
rect -697 -349 -503 -303
rect -397 303 -203 349
rect -397 -349 -203 -303
rect -97 303 97 349
rect -97 -349 97 -303
rect 203 303 397 349
rect 203 -349 397 -303
rect 503 303 697 349
rect 503 -349 697 -303
rect 803 303 997 349
rect 803 -349 997 -303
rect 1103 303 1297 349
rect 1103 -349 1297 -303
rect 1403 303 1597 349
rect 1403 -349 1597 -303
rect 1703 303 1897 349
rect 1703 -349 1897 -303
rect 2003 303 2197 349
rect 2003 -349 2197 -303
rect 2303 303 2497 349
rect 2303 -349 2497 -303
rect -2497 -525 -2303 -479
rect -2497 -1177 -2303 -1131
rect -2197 -525 -2003 -479
rect -2197 -1177 -2003 -1131
rect -1897 -525 -1703 -479
rect -1897 -1177 -1703 -1131
rect -1597 -525 -1403 -479
rect -1597 -1177 -1403 -1131
rect -1297 -525 -1103 -479
rect -1297 -1177 -1103 -1131
rect -997 -525 -803 -479
rect -997 -1177 -803 -1131
rect -697 -525 -503 -479
rect -697 -1177 -503 -1131
rect -397 -525 -203 -479
rect -397 -1177 -203 -1131
rect -97 -525 97 -479
rect -97 -1177 97 -1131
rect 203 -525 397 -479
rect 203 -1177 397 -1131
rect 503 -525 697 -479
rect 503 -1177 697 -1131
rect 803 -525 997 -479
rect 803 -1177 997 -1131
rect 1103 -525 1297 -479
rect 1103 -1177 1297 -1131
rect 1403 -525 1597 -479
rect 1403 -1177 1597 -1131
rect 1703 -525 1897 -479
rect 1703 -1177 1897 -1131
rect 2003 -525 2197 -479
rect 2003 -1177 2197 -1131
rect 2303 -525 2497 -479
rect 2303 -1177 2497 -1131
rect -2497 -1353 -2303 -1307
rect -2497 -2005 -2303 -1959
rect -2197 -1353 -2003 -1307
rect -2197 -2005 -2003 -1959
rect -1897 -1353 -1703 -1307
rect -1897 -2005 -1703 -1959
rect -1597 -1353 -1403 -1307
rect -1597 -2005 -1403 -1959
rect -1297 -1353 -1103 -1307
rect -1297 -2005 -1103 -1959
rect -997 -1353 -803 -1307
rect -997 -2005 -803 -1959
rect -697 -1353 -503 -1307
rect -697 -2005 -503 -1959
rect -397 -1353 -203 -1307
rect -397 -2005 -203 -1959
rect -97 -1353 97 -1307
rect -97 -2005 97 -1959
rect 203 -1353 397 -1307
rect 203 -2005 397 -1959
rect 503 -1353 697 -1307
rect 503 -2005 697 -1959
rect 803 -1353 997 -1307
rect 803 -2005 997 -1959
rect 1103 -1353 1297 -1307
rect 1103 -2005 1297 -1959
rect 1403 -1353 1597 -1307
rect 1403 -2005 1597 -1959
rect 1703 -1353 1897 -1307
rect 1703 -2005 1897 -1959
rect 2003 -1353 2197 -1307
rect 2003 -2005 2197 -1959
rect 2303 -1353 2497 -1307
rect 2303 -2005 2497 -1959
rect -2497 -2181 -2303 -2135
rect -2497 -2833 -2303 -2787
rect -2197 -2181 -2003 -2135
rect -2197 -2833 -2003 -2787
rect -1897 -2181 -1703 -2135
rect -1897 -2833 -1703 -2787
rect -1597 -2181 -1403 -2135
rect -1597 -2833 -1403 -2787
rect -1297 -2181 -1103 -2135
rect -1297 -2833 -1103 -2787
rect -997 -2181 -803 -2135
rect -997 -2833 -803 -2787
rect -697 -2181 -503 -2135
rect -697 -2833 -503 -2787
rect -397 -2181 -203 -2135
rect -397 -2833 -203 -2787
rect -97 -2181 97 -2135
rect -97 -2833 97 -2787
rect 203 -2181 397 -2135
rect 203 -2833 397 -2787
rect 503 -2181 697 -2135
rect 503 -2833 697 -2787
rect 803 -2181 997 -2135
rect 803 -2833 997 -2787
rect 1103 -2181 1297 -2135
rect 1103 -2833 1297 -2787
rect 1403 -2181 1597 -2135
rect 1403 -2833 1597 -2787
rect 1703 -2181 1897 -2135
rect 1703 -2833 1897 -2787
rect 2003 -2181 2197 -2135
rect 2003 -2833 2197 -2787
rect 2303 -2181 2497 -2135
rect 2303 -2833 2497 -2787
<< ppolyres >>
rect -2510 2224 -2290 2744
rect -2210 2224 -1990 2744
rect -1910 2224 -1690 2744
rect -1610 2224 -1390 2744
rect -1310 2224 -1090 2744
rect -1010 2224 -790 2744
rect -710 2224 -490 2744
rect -410 2224 -190 2744
rect -110 2224 110 2744
rect 190 2224 410 2744
rect 490 2224 710 2744
rect 790 2224 1010 2744
rect 1090 2224 1310 2744
rect 1390 2224 1610 2744
rect 1690 2224 1910 2744
rect 1990 2224 2210 2744
rect 2290 2224 2510 2744
rect -2510 1396 -2290 1916
rect -2210 1396 -1990 1916
rect -1910 1396 -1690 1916
rect -1610 1396 -1390 1916
rect -1310 1396 -1090 1916
rect -1010 1396 -790 1916
rect -710 1396 -490 1916
rect -410 1396 -190 1916
rect -110 1396 110 1916
rect 190 1396 410 1916
rect 490 1396 710 1916
rect 790 1396 1010 1916
rect 1090 1396 1310 1916
rect 1390 1396 1610 1916
rect 1690 1396 1910 1916
rect 1990 1396 2210 1916
rect 2290 1396 2510 1916
rect -2510 568 -2290 1088
rect -2210 568 -1990 1088
rect -1910 568 -1690 1088
rect -1610 568 -1390 1088
rect -1310 568 -1090 1088
rect -1010 568 -790 1088
rect -710 568 -490 1088
rect -410 568 -190 1088
rect -110 568 110 1088
rect 190 568 410 1088
rect 490 568 710 1088
rect 790 568 1010 1088
rect 1090 568 1310 1088
rect 1390 568 1610 1088
rect 1690 568 1910 1088
rect 1990 568 2210 1088
rect 2290 568 2510 1088
rect -2510 -260 -2290 260
rect -2210 -260 -1990 260
rect -1910 -260 -1690 260
rect -1610 -260 -1390 260
rect -1310 -260 -1090 260
rect -1010 -260 -790 260
rect -710 -260 -490 260
rect -410 -260 -190 260
rect -110 -260 110 260
rect 190 -260 410 260
rect 490 -260 710 260
rect 790 -260 1010 260
rect 1090 -260 1310 260
rect 1390 -260 1610 260
rect 1690 -260 1910 260
rect 1990 -260 2210 260
rect 2290 -260 2510 260
rect -2510 -1088 -2290 -568
rect -2210 -1088 -1990 -568
rect -1910 -1088 -1690 -568
rect -1610 -1088 -1390 -568
rect -1310 -1088 -1090 -568
rect -1010 -1088 -790 -568
rect -710 -1088 -490 -568
rect -410 -1088 -190 -568
rect -110 -1088 110 -568
rect 190 -1088 410 -568
rect 490 -1088 710 -568
rect 790 -1088 1010 -568
rect 1090 -1088 1310 -568
rect 1390 -1088 1610 -568
rect 1690 -1088 1910 -568
rect 1990 -1088 2210 -568
rect 2290 -1088 2510 -568
rect -2510 -1916 -2290 -1396
rect -2210 -1916 -1990 -1396
rect -1910 -1916 -1690 -1396
rect -1610 -1916 -1390 -1396
rect -1310 -1916 -1090 -1396
rect -1010 -1916 -790 -1396
rect -710 -1916 -490 -1396
rect -410 -1916 -190 -1396
rect -110 -1916 110 -1396
rect 190 -1916 410 -1396
rect 490 -1916 710 -1396
rect 790 -1916 1010 -1396
rect 1090 -1916 1310 -1396
rect 1390 -1916 1610 -1396
rect 1690 -1916 1910 -1396
rect 1990 -1916 2210 -1396
rect 2290 -1916 2510 -1396
rect -2510 -2744 -2290 -2224
rect -2210 -2744 -1990 -2224
rect -1910 -2744 -1690 -2224
rect -1610 -2744 -1390 -2224
rect -1310 -2744 -1090 -2224
rect -1010 -2744 -790 -2224
rect -710 -2744 -490 -2224
rect -410 -2744 -190 -2224
rect -110 -2744 110 -2224
rect 190 -2744 410 -2224
rect 490 -2744 710 -2224
rect 790 -2744 1010 -2224
rect 1090 -2744 1310 -2224
rect 1390 -2744 1610 -2224
rect 1690 -2744 1910 -2224
rect 1990 -2744 2210 -2224
rect 2290 -2744 2510 -2224
<< metal1 >>
rect -2689 2979 -2586 3025
rect 2586 2979 2689 3025
rect -2689 2922 -2643 2979
rect 2643 2922 2689 2979
rect -2508 2787 -2497 2833
rect -2303 2787 -2292 2833
rect -2208 2787 -2197 2833
rect -2003 2787 -1992 2833
rect -1908 2787 -1897 2833
rect -1703 2787 -1692 2833
rect -1608 2787 -1597 2833
rect -1403 2787 -1392 2833
rect -1308 2787 -1297 2833
rect -1103 2787 -1092 2833
rect -1008 2787 -997 2833
rect -803 2787 -792 2833
rect -708 2787 -697 2833
rect -503 2787 -492 2833
rect -408 2787 -397 2833
rect -203 2787 -192 2833
rect -108 2787 -97 2833
rect 97 2787 108 2833
rect 192 2787 203 2833
rect 397 2787 408 2833
rect 492 2787 503 2833
rect 697 2787 708 2833
rect 792 2787 803 2833
rect 997 2787 1008 2833
rect 1092 2787 1103 2833
rect 1297 2787 1308 2833
rect 1392 2787 1403 2833
rect 1597 2787 1608 2833
rect 1692 2787 1703 2833
rect 1897 2787 1908 2833
rect 1992 2787 2003 2833
rect 2197 2787 2208 2833
rect 2292 2787 2303 2833
rect 2497 2787 2508 2833
rect -2508 2135 -2497 2181
rect -2303 2135 -2292 2181
rect -2208 2135 -2197 2181
rect -2003 2135 -1992 2181
rect -1908 2135 -1897 2181
rect -1703 2135 -1692 2181
rect -1608 2135 -1597 2181
rect -1403 2135 -1392 2181
rect -1308 2135 -1297 2181
rect -1103 2135 -1092 2181
rect -1008 2135 -997 2181
rect -803 2135 -792 2181
rect -708 2135 -697 2181
rect -503 2135 -492 2181
rect -408 2135 -397 2181
rect -203 2135 -192 2181
rect -108 2135 -97 2181
rect 97 2135 108 2181
rect 192 2135 203 2181
rect 397 2135 408 2181
rect 492 2135 503 2181
rect 697 2135 708 2181
rect 792 2135 803 2181
rect 997 2135 1008 2181
rect 1092 2135 1103 2181
rect 1297 2135 1308 2181
rect 1392 2135 1403 2181
rect 1597 2135 1608 2181
rect 1692 2135 1703 2181
rect 1897 2135 1908 2181
rect 1992 2135 2003 2181
rect 2197 2135 2208 2181
rect 2292 2135 2303 2181
rect 2497 2135 2508 2181
rect -2508 1959 -2497 2005
rect -2303 1959 -2292 2005
rect -2208 1959 -2197 2005
rect -2003 1959 -1992 2005
rect -1908 1959 -1897 2005
rect -1703 1959 -1692 2005
rect -1608 1959 -1597 2005
rect -1403 1959 -1392 2005
rect -1308 1959 -1297 2005
rect -1103 1959 -1092 2005
rect -1008 1959 -997 2005
rect -803 1959 -792 2005
rect -708 1959 -697 2005
rect -503 1959 -492 2005
rect -408 1959 -397 2005
rect -203 1959 -192 2005
rect -108 1959 -97 2005
rect 97 1959 108 2005
rect 192 1959 203 2005
rect 397 1959 408 2005
rect 492 1959 503 2005
rect 697 1959 708 2005
rect 792 1959 803 2005
rect 997 1959 1008 2005
rect 1092 1959 1103 2005
rect 1297 1959 1308 2005
rect 1392 1959 1403 2005
rect 1597 1959 1608 2005
rect 1692 1959 1703 2005
rect 1897 1959 1908 2005
rect 1992 1959 2003 2005
rect 2197 1959 2208 2005
rect 2292 1959 2303 2005
rect 2497 1959 2508 2005
rect -2508 1307 -2497 1353
rect -2303 1307 -2292 1353
rect -2208 1307 -2197 1353
rect -2003 1307 -1992 1353
rect -1908 1307 -1897 1353
rect -1703 1307 -1692 1353
rect -1608 1307 -1597 1353
rect -1403 1307 -1392 1353
rect -1308 1307 -1297 1353
rect -1103 1307 -1092 1353
rect -1008 1307 -997 1353
rect -803 1307 -792 1353
rect -708 1307 -697 1353
rect -503 1307 -492 1353
rect -408 1307 -397 1353
rect -203 1307 -192 1353
rect -108 1307 -97 1353
rect 97 1307 108 1353
rect 192 1307 203 1353
rect 397 1307 408 1353
rect 492 1307 503 1353
rect 697 1307 708 1353
rect 792 1307 803 1353
rect 997 1307 1008 1353
rect 1092 1307 1103 1353
rect 1297 1307 1308 1353
rect 1392 1307 1403 1353
rect 1597 1307 1608 1353
rect 1692 1307 1703 1353
rect 1897 1307 1908 1353
rect 1992 1307 2003 1353
rect 2197 1307 2208 1353
rect 2292 1307 2303 1353
rect 2497 1307 2508 1353
rect -2508 1131 -2497 1177
rect -2303 1131 -2292 1177
rect -2208 1131 -2197 1177
rect -2003 1131 -1992 1177
rect -1908 1131 -1897 1177
rect -1703 1131 -1692 1177
rect -1608 1131 -1597 1177
rect -1403 1131 -1392 1177
rect -1308 1131 -1297 1177
rect -1103 1131 -1092 1177
rect -1008 1131 -997 1177
rect -803 1131 -792 1177
rect -708 1131 -697 1177
rect -503 1131 -492 1177
rect -408 1131 -397 1177
rect -203 1131 -192 1177
rect -108 1131 -97 1177
rect 97 1131 108 1177
rect 192 1131 203 1177
rect 397 1131 408 1177
rect 492 1131 503 1177
rect 697 1131 708 1177
rect 792 1131 803 1177
rect 997 1131 1008 1177
rect 1092 1131 1103 1177
rect 1297 1131 1308 1177
rect 1392 1131 1403 1177
rect 1597 1131 1608 1177
rect 1692 1131 1703 1177
rect 1897 1131 1908 1177
rect 1992 1131 2003 1177
rect 2197 1131 2208 1177
rect 2292 1131 2303 1177
rect 2497 1131 2508 1177
rect -2508 479 -2497 525
rect -2303 479 -2292 525
rect -2208 479 -2197 525
rect -2003 479 -1992 525
rect -1908 479 -1897 525
rect -1703 479 -1692 525
rect -1608 479 -1597 525
rect -1403 479 -1392 525
rect -1308 479 -1297 525
rect -1103 479 -1092 525
rect -1008 479 -997 525
rect -803 479 -792 525
rect -708 479 -697 525
rect -503 479 -492 525
rect -408 479 -397 525
rect -203 479 -192 525
rect -108 479 -97 525
rect 97 479 108 525
rect 192 479 203 525
rect 397 479 408 525
rect 492 479 503 525
rect 697 479 708 525
rect 792 479 803 525
rect 997 479 1008 525
rect 1092 479 1103 525
rect 1297 479 1308 525
rect 1392 479 1403 525
rect 1597 479 1608 525
rect 1692 479 1703 525
rect 1897 479 1908 525
rect 1992 479 2003 525
rect 2197 479 2208 525
rect 2292 479 2303 525
rect 2497 479 2508 525
rect -2508 303 -2497 349
rect -2303 303 -2292 349
rect -2208 303 -2197 349
rect -2003 303 -1992 349
rect -1908 303 -1897 349
rect -1703 303 -1692 349
rect -1608 303 -1597 349
rect -1403 303 -1392 349
rect -1308 303 -1297 349
rect -1103 303 -1092 349
rect -1008 303 -997 349
rect -803 303 -792 349
rect -708 303 -697 349
rect -503 303 -492 349
rect -408 303 -397 349
rect -203 303 -192 349
rect -108 303 -97 349
rect 97 303 108 349
rect 192 303 203 349
rect 397 303 408 349
rect 492 303 503 349
rect 697 303 708 349
rect 792 303 803 349
rect 997 303 1008 349
rect 1092 303 1103 349
rect 1297 303 1308 349
rect 1392 303 1403 349
rect 1597 303 1608 349
rect 1692 303 1703 349
rect 1897 303 1908 349
rect 1992 303 2003 349
rect 2197 303 2208 349
rect 2292 303 2303 349
rect 2497 303 2508 349
rect -2508 -349 -2497 -303
rect -2303 -349 -2292 -303
rect -2208 -349 -2197 -303
rect -2003 -349 -1992 -303
rect -1908 -349 -1897 -303
rect -1703 -349 -1692 -303
rect -1608 -349 -1597 -303
rect -1403 -349 -1392 -303
rect -1308 -349 -1297 -303
rect -1103 -349 -1092 -303
rect -1008 -349 -997 -303
rect -803 -349 -792 -303
rect -708 -349 -697 -303
rect -503 -349 -492 -303
rect -408 -349 -397 -303
rect -203 -349 -192 -303
rect -108 -349 -97 -303
rect 97 -349 108 -303
rect 192 -349 203 -303
rect 397 -349 408 -303
rect 492 -349 503 -303
rect 697 -349 708 -303
rect 792 -349 803 -303
rect 997 -349 1008 -303
rect 1092 -349 1103 -303
rect 1297 -349 1308 -303
rect 1392 -349 1403 -303
rect 1597 -349 1608 -303
rect 1692 -349 1703 -303
rect 1897 -349 1908 -303
rect 1992 -349 2003 -303
rect 2197 -349 2208 -303
rect 2292 -349 2303 -303
rect 2497 -349 2508 -303
rect -2508 -525 -2497 -479
rect -2303 -525 -2292 -479
rect -2208 -525 -2197 -479
rect -2003 -525 -1992 -479
rect -1908 -525 -1897 -479
rect -1703 -525 -1692 -479
rect -1608 -525 -1597 -479
rect -1403 -525 -1392 -479
rect -1308 -525 -1297 -479
rect -1103 -525 -1092 -479
rect -1008 -525 -997 -479
rect -803 -525 -792 -479
rect -708 -525 -697 -479
rect -503 -525 -492 -479
rect -408 -525 -397 -479
rect -203 -525 -192 -479
rect -108 -525 -97 -479
rect 97 -525 108 -479
rect 192 -525 203 -479
rect 397 -525 408 -479
rect 492 -525 503 -479
rect 697 -525 708 -479
rect 792 -525 803 -479
rect 997 -525 1008 -479
rect 1092 -525 1103 -479
rect 1297 -525 1308 -479
rect 1392 -525 1403 -479
rect 1597 -525 1608 -479
rect 1692 -525 1703 -479
rect 1897 -525 1908 -479
rect 1992 -525 2003 -479
rect 2197 -525 2208 -479
rect 2292 -525 2303 -479
rect 2497 -525 2508 -479
rect -2508 -1177 -2497 -1131
rect -2303 -1177 -2292 -1131
rect -2208 -1177 -2197 -1131
rect -2003 -1177 -1992 -1131
rect -1908 -1177 -1897 -1131
rect -1703 -1177 -1692 -1131
rect -1608 -1177 -1597 -1131
rect -1403 -1177 -1392 -1131
rect -1308 -1177 -1297 -1131
rect -1103 -1177 -1092 -1131
rect -1008 -1177 -997 -1131
rect -803 -1177 -792 -1131
rect -708 -1177 -697 -1131
rect -503 -1177 -492 -1131
rect -408 -1177 -397 -1131
rect -203 -1177 -192 -1131
rect -108 -1177 -97 -1131
rect 97 -1177 108 -1131
rect 192 -1177 203 -1131
rect 397 -1177 408 -1131
rect 492 -1177 503 -1131
rect 697 -1177 708 -1131
rect 792 -1177 803 -1131
rect 997 -1177 1008 -1131
rect 1092 -1177 1103 -1131
rect 1297 -1177 1308 -1131
rect 1392 -1177 1403 -1131
rect 1597 -1177 1608 -1131
rect 1692 -1177 1703 -1131
rect 1897 -1177 1908 -1131
rect 1992 -1177 2003 -1131
rect 2197 -1177 2208 -1131
rect 2292 -1177 2303 -1131
rect 2497 -1177 2508 -1131
rect -2508 -1353 -2497 -1307
rect -2303 -1353 -2292 -1307
rect -2208 -1353 -2197 -1307
rect -2003 -1353 -1992 -1307
rect -1908 -1353 -1897 -1307
rect -1703 -1353 -1692 -1307
rect -1608 -1353 -1597 -1307
rect -1403 -1353 -1392 -1307
rect -1308 -1353 -1297 -1307
rect -1103 -1353 -1092 -1307
rect -1008 -1353 -997 -1307
rect -803 -1353 -792 -1307
rect -708 -1353 -697 -1307
rect -503 -1353 -492 -1307
rect -408 -1353 -397 -1307
rect -203 -1353 -192 -1307
rect -108 -1353 -97 -1307
rect 97 -1353 108 -1307
rect 192 -1353 203 -1307
rect 397 -1353 408 -1307
rect 492 -1353 503 -1307
rect 697 -1353 708 -1307
rect 792 -1353 803 -1307
rect 997 -1353 1008 -1307
rect 1092 -1353 1103 -1307
rect 1297 -1353 1308 -1307
rect 1392 -1353 1403 -1307
rect 1597 -1353 1608 -1307
rect 1692 -1353 1703 -1307
rect 1897 -1353 1908 -1307
rect 1992 -1353 2003 -1307
rect 2197 -1353 2208 -1307
rect 2292 -1353 2303 -1307
rect 2497 -1353 2508 -1307
rect -2508 -2005 -2497 -1959
rect -2303 -2005 -2292 -1959
rect -2208 -2005 -2197 -1959
rect -2003 -2005 -1992 -1959
rect -1908 -2005 -1897 -1959
rect -1703 -2005 -1692 -1959
rect -1608 -2005 -1597 -1959
rect -1403 -2005 -1392 -1959
rect -1308 -2005 -1297 -1959
rect -1103 -2005 -1092 -1959
rect -1008 -2005 -997 -1959
rect -803 -2005 -792 -1959
rect -708 -2005 -697 -1959
rect -503 -2005 -492 -1959
rect -408 -2005 -397 -1959
rect -203 -2005 -192 -1959
rect -108 -2005 -97 -1959
rect 97 -2005 108 -1959
rect 192 -2005 203 -1959
rect 397 -2005 408 -1959
rect 492 -2005 503 -1959
rect 697 -2005 708 -1959
rect 792 -2005 803 -1959
rect 997 -2005 1008 -1959
rect 1092 -2005 1103 -1959
rect 1297 -2005 1308 -1959
rect 1392 -2005 1403 -1959
rect 1597 -2005 1608 -1959
rect 1692 -2005 1703 -1959
rect 1897 -2005 1908 -1959
rect 1992 -2005 2003 -1959
rect 2197 -2005 2208 -1959
rect 2292 -2005 2303 -1959
rect 2497 -2005 2508 -1959
rect -2508 -2181 -2497 -2135
rect -2303 -2181 -2292 -2135
rect -2208 -2181 -2197 -2135
rect -2003 -2181 -1992 -2135
rect -1908 -2181 -1897 -2135
rect -1703 -2181 -1692 -2135
rect -1608 -2181 -1597 -2135
rect -1403 -2181 -1392 -2135
rect -1308 -2181 -1297 -2135
rect -1103 -2181 -1092 -2135
rect -1008 -2181 -997 -2135
rect -803 -2181 -792 -2135
rect -708 -2181 -697 -2135
rect -503 -2181 -492 -2135
rect -408 -2181 -397 -2135
rect -203 -2181 -192 -2135
rect -108 -2181 -97 -2135
rect 97 -2181 108 -2135
rect 192 -2181 203 -2135
rect 397 -2181 408 -2135
rect 492 -2181 503 -2135
rect 697 -2181 708 -2135
rect 792 -2181 803 -2135
rect 997 -2181 1008 -2135
rect 1092 -2181 1103 -2135
rect 1297 -2181 1308 -2135
rect 1392 -2181 1403 -2135
rect 1597 -2181 1608 -2135
rect 1692 -2181 1703 -2135
rect 1897 -2181 1908 -2135
rect 1992 -2181 2003 -2135
rect 2197 -2181 2208 -2135
rect 2292 -2181 2303 -2135
rect 2497 -2181 2508 -2135
rect -2508 -2833 -2497 -2787
rect -2303 -2833 -2292 -2787
rect -2208 -2833 -2197 -2787
rect -2003 -2833 -1992 -2787
rect -1908 -2833 -1897 -2787
rect -1703 -2833 -1692 -2787
rect -1608 -2833 -1597 -2787
rect -1403 -2833 -1392 -2787
rect -1308 -2833 -1297 -2787
rect -1103 -2833 -1092 -2787
rect -1008 -2833 -997 -2787
rect -803 -2833 -792 -2787
rect -708 -2833 -697 -2787
rect -503 -2833 -492 -2787
rect -408 -2833 -397 -2787
rect -203 -2833 -192 -2787
rect -108 -2833 -97 -2787
rect 97 -2833 108 -2787
rect 192 -2833 203 -2787
rect 397 -2833 408 -2787
rect 492 -2833 503 -2787
rect 697 -2833 708 -2787
rect 792 -2833 803 -2787
rect 997 -2833 1008 -2787
rect 1092 -2833 1103 -2787
rect 1297 -2833 1308 -2787
rect 1392 -2833 1403 -2787
rect 1597 -2833 1608 -2787
rect 1692 -2833 1703 -2787
rect 1897 -2833 1908 -2787
rect 1992 -2833 2003 -2787
rect 2197 -2833 2208 -2787
rect 2292 -2833 2303 -2787
rect 2497 -2833 2508 -2787
rect -2689 -2979 -2643 -2922
rect 2643 -2979 2689 -2922
rect -2689 -3025 -2586 -2979
rect 2586 -3025 2689 -2979
<< properties >>
string FIXED_BBOX -2666 -3002 2666 3002
string gencell ppolyf_u
string library gf180mcu
string parameters w 1.10 l 2.6 m 7 nx 17 wmin 0.80 lmin 1.00 rho 315 val 795.145 dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1
<< end >>
