* NGSPICE file created from INVERTER_magic_flat.ext - technology: gf180mcuC

.subckt INVERTER_magic_flat IN OUT VDD VSS
X0 OUT IN.t0 VSS.t1 VSS.t0 nfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X1 VSS.t4 VSS.t2 VSS.t4 VSS.t3 nfet_03v3 ad=0 pd=0 as=0.155p ps=1.64u w=0.25u l=0.28u
X2 OUT IN.t1 VDD.t4 VDD.t3 pfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X3 VDD IN.t2 OUT.t1 VDD.t0 pfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
R0 IN.t2 IN.n0 31.2628
R1 IN.n0 IN.t0 27.5059
R2 IN IN.t2 18.8858
R3 IN.n0 IN.t1 10.2987
R4 VSS.n1 VSS.t0 755.814
R5 VSS.n5 VSS.t3 279.721
R6 VSS.t0 VSS.n0 178.946
R7 VSS.n4 VSS.t2 16.6451
R8 VSS.n2 VSS.n0 10.7975
R9 VSS.n5 VSS.n2 10.7975
R10 VSS.n3 VSS.t1 6.73354
R11 VSS VSS.n2 5.2005
R12 VSS VSS.n2 5.2005
R13 VSS.n3 VSS.t4 2.836
R14 VSS.n2 VSS.n1 2.6005
R15 VSS VSS.n0 2.2994
R16 VSS.n6 VSS.n5 2.21164
R17 VSS.n4 VSS.n3 1.70051
R18 VSS.n6 VSS.n4 0.0905
R19 VSS VSS.n6 0.08825
R20 OUT.n1 OUT.t1 9.68225
R21 OUT.n3 OUT.n2 9.04464
R22 OUT.n1 OUT.n0 9.02485
R23 OUT OUT.n3 0.182457
R24 OUT.n3 OUT.n1 0.0102826
R25 VDD.n4 VDD.t3 192.309
R26 VDD.n6 VDD.t0 73.5996
R27 VDD.t3 VDD.n3 47.9603
R28 VDD.n5 VDD.n3 9.73809
R29 VDD.n6 VDD.n5 9.73765
R30 VDD.n1 VDD.n0 6.3005
R31 VDD.n1 VDD.t4 6.3005
R32 VDD VDD.n5 6.3005
R33 VDD VDD.n5 6.3005
R34 VDD.n5 VDD.n4 3.1505
R35 VDD.n2 VDD.n1 2.99094
R36 VDD VDD.n6 2.62331
R37 VDD.n3 VDD.n2 2.61557
R38 VDD VDD.n2 0.00725
C0 OUT VDD 0.221f
C1 OUT IN 0.115f
C2 VDD IN 0.58f
.ends

