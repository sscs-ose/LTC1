magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2371 -2042 2371 2042
<< polysilicon >>
rect -371 23 371 42
rect -371 -23 -352 23
rect 352 -23 371 23
rect -371 -42 371 -23
<< polycontact >>
rect -352 -23 352 23
<< metal1 >>
rect -363 23 363 34
rect -363 -23 -352 23
rect 352 -23 363 23
rect -363 -34 363 -23
<< end >>
