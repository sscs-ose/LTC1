* NGSPICE file created from Inv_16x_Layout_flat.ext - technology: gf180mcuC

.subckt INV_16x_PEX VDD OUT IN VSS
X0 OUT IN.t0 VDD.t1 VDD.t0 pfet_03v3 ad=0.194p pd=1.76u as=0.194p ps=1.76u w=0.44u l=2.24u
X1 OUT IN.t1 VSS.t1 VSS.t0 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=2.24u
R0 IN.n0 IN.t0 20.6254
R1 IN IN.n0 14.0348
R2 IN.n0 IN.t1 12.9662
R3 VDD.t0 VDD.n0 112.05
R4 VDD.n1 VDD.t0 91.8808
R5 VDD.n2 VDD.n0 8.25406
R6 VDD.n8 VDD.n2 8.2255
R7 VDD.n3 VDD.t1 7.06752
R8 VDD VDD.n2 6.3005
R9 VDD VDD.n2 6.3005
R10 VDD.n2 VDD.n1 3.1505
R11 VDD.n9 VDD.n8 3.1505
R12 VDD.n8 VDD.n7 3.1505
R13 VDD.n6 VDD.n5 3.1505
R14 VDD VDD.n0 2.46788
R15 VDD.n5 VDD.n4 0.121293
R16 VDD VDD.n9 0.0760357
R17 VDD.n9 VDD.n6 0.0760357
R18 VDD.n6 VDD.n3 0.0366607
R19 OUT OUT.n1 9.42306
R20 OUT OUT.n0 7.41143
R21 VSS.n1 VSS.t0 604.271
R22 VSS.n5 VSS.t1 9.32958
R23 VSS.n8 VSS.n3 9.13939
R24 VSS VSS.n3 5.2005
R25 VSS VSS.n3 5.2005
R26 VSS.n5 VSS.n4 2.60371
R27 VSS.n9 VSS.n8 2.6005
R28 VSS.n7 VSS.n6 2.6005
R29 VSS.n3 VSS.n2 1.92228
R30 VSS VSS.n2 1.62146
R31 VSS.n1 VSS.n0 0.472445
R32 VSS.n2 VSS.n1 0.173689
R33 VSS VSS.n9 0.0760357
R34 VSS.n9 VSS.n7 0.0760357
R35 VSS.n7 VSS.n5 0.0728214
C0 OUT IN 0.05f
C1 VDD IN 0.416f
C2 OUT VDD 0.0609f
.ends

