magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1154 -1073 1154 1073
<< metal1 >>
rect -154 67 154 73
rect -154 41 -148 67
rect -122 41 -94 67
rect -68 41 -40 67
rect -14 41 14 67
rect 40 41 68 67
rect 94 41 122 67
rect 148 41 154 67
rect -154 13 154 41
rect -154 -13 -148 13
rect -122 -13 -94 13
rect -68 -13 -40 13
rect -14 -13 14 13
rect 40 -13 68 13
rect 94 -13 122 13
rect 148 -13 154 13
rect -154 -41 154 -13
rect -154 -67 -148 -41
rect -122 -67 -94 -41
rect -68 -67 -40 -41
rect -14 -67 14 -41
rect 40 -67 68 -41
rect 94 -67 122 -41
rect 148 -67 154 -41
rect -154 -73 154 -67
<< via1 >>
rect -148 41 -122 67
rect -94 41 -68 67
rect -40 41 -14 67
rect 14 41 40 67
rect 68 41 94 67
rect 122 41 148 67
rect -148 -13 -122 13
rect -94 -13 -68 13
rect -40 -13 -14 13
rect 14 -13 40 13
rect 68 -13 94 13
rect 122 -13 148 13
rect -148 -67 -122 -41
rect -94 -67 -68 -41
rect -40 -67 -14 -41
rect 14 -67 40 -41
rect 68 -67 94 -41
rect 122 -67 148 -41
<< metal2 >>
rect -154 67 154 73
rect -154 41 -148 67
rect -122 41 -94 67
rect -68 41 -40 67
rect -14 41 14 67
rect 40 41 68 67
rect 94 41 122 67
rect 148 41 154 67
rect -154 13 154 41
rect -154 -13 -148 13
rect -122 -13 -94 13
rect -68 -13 -40 13
rect -14 -13 14 13
rect 40 -13 68 13
rect 94 -13 122 13
rect 148 -13 154 13
rect -154 -41 154 -13
rect -154 -67 -148 -41
rect -122 -67 -94 -41
rect -68 -67 -40 -41
rect -14 -67 14 -41
rect 40 -67 68 -41
rect 94 -67 122 -41
rect 148 -67 154 -41
rect -154 -73 154 -67
<< end >>
