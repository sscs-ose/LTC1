magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1343 1019 1343
<< metal2 >>
rect -19 326 19 343
rect -19 -326 -14 326
rect 14 -326 19 326
rect -19 -343 19 -326
<< via2 >>
rect -14 -326 14 326
<< metal3 >>
rect -19 326 19 343
rect -19 -326 -14 326
rect 14 -326 19 326
rect -19 -343 19 -326
<< end >>
