magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1045 -1253 1045 1253
<< metal2 >>
rect -45 248 45 253
rect -45 -248 -40 248
rect 40 -248 45 248
rect -45 -253 45 -248
<< via2 >>
rect -40 -248 40 248
<< metal3 >>
rect -45 248 45 253
rect -45 -248 -40 248
rect 40 -248 45 248
rect -45 -253 45 -248
<< end >>
