magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2044 -1600 4074 10000
<< metal1 >>
rect -44 400 200 8000
rect 430 401 2074 8000
<< metal2 >>
rect -44 400 200 8000
rect 430 401 2074 8000
use M2_M1_CDNS_69033583165673  M2_M1_CDNS_69033583165673_0
timestamp 1713338890
transform 1 0 1252 0 1 4199
box -782 -3758 782 3758
use M2_M1_CDNS_69033583165674  M2_M1_CDNS_69033583165674_0
timestamp 1713338890
transform 1 0 78 0 1 4207
box -90 -3758 90 3758
use M3_M2_CDNS_69033583165670  M3_M2_CDNS_69033583165670_0
timestamp 1713338890
transform 1 0 80 0 1 6840
box -90 -818 90 818
use M3_M2_CDNS_69033583165671  M3_M2_CDNS_69033583165671_0
timestamp 1713338890
transform 1 0 80 0 1 3979
box -90 -1078 90 1078
use M3_M2_CDNS_69033583165672  M3_M2_CDNS_69033583165672_0
timestamp 1713338890
transform 1 0 80 0 1 1340
box -90 -662 90 662
<< end >>
