magic
tech gf180mcuC
magscale 1 10
timestamp 1694585882
<< nwell >>
rect 2610 372 2715 813
rect 1570 -1476 1734 -988
rect 2863 -1528 2896 -1087
rect 1249 -2045 1327 -1946
rect 1250 -2414 1327 -2045
rect 2859 -2486 2896 -2045
rect 1570 -3427 1590 -2906
rect 1570 -4169 1618 -3868
rect 1535 -4240 1618 -4169
rect 1570 -4336 1618 -4240
<< metal1 >>
rect -821 847 -747 856
rect 51 847 3508 891
rect -821 791 -812 847
rect -756 791 3508 847
rect -821 781 -747 791
rect 51 773 3508 791
rect 2610 700 3508 773
rect -655 576 -581 585
rect -10 576 89 579
rect -655 520 -646 576
rect -590 520 89 576
rect -655 511 -581 520
rect -10 492 89 520
rect -489 426 -417 435
rect -489 372 -480 426
rect -426 422 -417 426
rect -426 376 36 422
rect 1314 418 1360 422
rect -426 372 -417 376
rect -489 363 -417 372
rect 1234 371 1360 418
rect 3558 371 3568 418
rect -12 299 68 308
rect -12 243 0 299
rect 56 243 68 299
rect -12 234 68 243
rect 1250 113 1398 118
rect -198 100 -126 109
rect -198 46 -189 100
rect -135 97 -126 100
rect 54 97 3486 113
rect -135 48 3486 97
rect -135 46 -126 48
rect -198 37 -126 46
rect 54 0 3486 48
rect -822 -84 -748 -75
rect 41 -84 3311 -48
rect -822 -140 -812 -84
rect -756 -126 3311 -84
rect -756 -140 50 -126
rect -822 -149 -748 -140
rect 1250 -239 2179 -126
rect 3333 -344 3410 -329
rect -658 -375 -587 -363
rect -4 -370 79 -360
rect -21 -375 79 -370
rect -658 -431 -646 -375
rect -590 -376 79 -375
rect -590 -430 7 -376
rect 61 -430 79 -376
rect 3333 -400 3340 -344
rect 3396 -400 3410 -344
rect 3333 -414 3410 -400
rect -590 -431 79 -430
rect -658 -443 -587 -431
rect -21 -446 79 -431
rect -4 -447 79 -446
rect -500 -513 -428 -504
rect -500 -567 -491 -513
rect -437 -517 -428 -513
rect 2380 -509 2466 -501
rect -437 -563 46 -517
rect 2208 -521 2255 -520
rect -437 -567 -428 -563
rect -500 -576 -428 -567
rect 2182 -568 2264 -521
rect 2380 -565 2399 -509
rect 2455 -565 2466 -509
rect 2208 -657 2255 -568
rect 2380 -577 2466 -565
rect 3314 -568 3407 -521
rect 2358 -653 2452 -635
rect 2358 -657 2382 -653
rect 2208 -704 2382 -657
rect 2358 -707 2382 -704
rect 2436 -707 2452 -653
rect 2358 -726 2452 -707
rect -201 -854 -127 -846
rect 44 -849 3296 -826
rect -19 -854 3296 -849
rect -201 -910 -190 -854
rect -134 -910 3296 -854
rect -201 -918 -127 -910
rect -19 -913 3296 -910
rect 44 -939 3296 -913
rect -825 -1013 -747 -1005
rect 41 -1013 3682 -988
rect -825 -1069 -812 -1013
rect -756 -1069 3682 -1013
rect -825 -1081 -747 -1069
rect 41 -1087 3682 -1069
rect -658 -1193 -583 -1187
rect -57 -1193 19 -1185
rect -658 -1194 19 -1193
rect -658 -1249 -646 -1194
rect -591 -1249 -48 -1194
rect -658 -1250 -48 -1249
rect -658 -1260 -583 -1250
rect -57 -1251 -48 -1250
rect 9 -1251 19 -1194
rect -57 -1260 19 -1251
rect -502 -1370 -424 -1361
rect -502 -1424 -491 -1370
rect -437 -1374 -424 -1370
rect -437 -1420 84 -1374
rect -437 -1424 -424 -1420
rect -502 -1433 -424 -1424
rect -354 -1505 -274 -1496
rect -354 -1559 -344 -1505
rect -290 -1509 -274 -1505
rect -290 -1555 84 -1509
rect 1557 -1529 1676 -1482
rect 2772 -1492 2818 -1447
rect 3685 -1529 3759 -1482
rect -290 -1559 -274 -1555
rect -354 -1569 -274 -1559
rect -200 -1809 -127 -1800
rect -200 -1863 -191 -1809
rect -137 -1812 -127 -1809
rect 51 -1812 3669 -1782
rect -137 -1861 3669 -1812
rect -137 -1863 -127 -1861
rect -200 -1873 -127 -1863
rect 51 -1900 3669 -1861
rect -823 -1980 -749 -1969
rect 51 -1980 3678 -1946
rect -823 -2036 -812 -1980
rect -756 -2036 3678 -1980
rect -823 -2046 -749 -2036
rect 51 -2045 3678 -2036
rect 1253 -2250 1328 -2240
rect 1253 -2251 1329 -2250
rect -499 -2269 -421 -2258
rect -499 -2325 -487 -2269
rect -431 -2325 33 -2269
rect 1253 -2305 1266 -2251
rect 1320 -2255 1329 -2251
rect 1320 -2305 1373 -2255
rect 1253 -2315 1373 -2305
rect -499 -2334 -421 -2325
rect 1327 -2378 1373 -2315
rect -356 -2411 -275 -2401
rect -356 -2465 -343 -2411
rect -289 -2415 -275 -2411
rect -289 -2461 46 -2415
rect -289 -2465 -275 -2461
rect -356 -2474 -275 -2465
rect 1233 -2464 1280 -2419
rect 2758 -2440 2780 -2405
rect 1233 -2511 1370 -2464
rect 3681 -2487 3761 -2440
rect -662 -2551 -583 -2541
rect -15 -2547 67 -2532
rect -15 -2551 2 -2547
rect -662 -2607 -646 -2551
rect -590 -2603 2 -2551
rect 58 -2603 67 -2547
rect -590 -2607 67 -2603
rect -662 -2617 -583 -2607
rect -15 -2623 67 -2607
rect -202 -2750 -121 -2738
rect 44 -2750 3656 -2745
rect -202 -2806 -190 -2750
rect -134 -2806 3656 -2750
rect -202 -2817 -121 -2806
rect 44 -2834 3656 -2806
rect 38 -2858 3656 -2834
rect -842 -2925 -744 -2912
rect 1570 -2925 2389 -2906
rect -842 -2981 -812 -2925
rect -756 -2981 2389 -2925
rect -842 -2999 -744 -2981
rect 1570 -3005 2389 -2981
rect -664 -3288 -582 -3278
rect -664 -3342 -649 -3288
rect -595 -3292 -582 -3288
rect -595 -3338 84 -3292
rect -595 -3342 -582 -3338
rect -664 -3351 -582 -3342
rect 1471 -3404 1524 -3365
rect -503 -3423 -422 -3413
rect -503 -3477 -490 -3423
rect -436 -3427 -422 -3423
rect -436 -3473 84 -3427
rect 2392 -3447 2485 -3400
rect -436 -3477 -422 -3473
rect -503 -3488 -422 -3477
rect -202 -3742 -127 -3733
rect -202 -3798 -190 -3742
rect -134 -3748 46 -3742
rect -134 -3798 2382 -3748
rect -202 -3814 -127 -3798
rect 38 -3812 2382 -3798
rect -825 -3896 -750 -3884
rect 41 -3896 4110 -3868
rect -825 -3952 -812 -3896
rect -756 -3952 4110 -3896
rect -825 -3967 -750 -3952
rect 41 -3967 4110 -3952
rect 2999 -4011 4110 -3967
rect 1534 -4174 1607 -4163
rect 1534 -4228 1543 -4174
rect 1597 -4228 1607 -4174
rect -664 -4250 -583 -4241
rect -664 -4304 -651 -4250
rect -597 -4254 -583 -4250
rect 1534 -4254 1607 -4228
rect -597 -4300 84 -4254
rect 1534 -4255 1616 -4254
rect 1543 -4300 1616 -4255
rect -597 -4304 -583 -4300
rect -664 -4315 -583 -4304
rect -508 -4385 -428 -4375
rect -508 -4439 -493 -4385
rect -439 -4389 -428 -4385
rect -439 -4435 84 -4389
rect 1534 -4435 1616 -4389
rect 3129 -4409 3244 -4362
rect 4114 -4409 4210 -4362
rect -439 -4439 -428 -4435
rect -508 -4450 -428 -4439
rect -355 -4502 -274 -4490
rect 19 -4502 92 -4500
rect -355 -4558 -340 -4502
rect -284 -4512 92 -4502
rect -284 -4558 30 -4512
rect -355 -4572 -274 -4558
rect 19 -4568 30 -4558
rect 86 -4568 92 -4512
rect 19 -4580 92 -4568
rect -204 -4670 -124 -4658
rect 54 -4670 4100 -4667
rect -204 -4726 -190 -4670
rect -134 -4726 4100 -4670
rect -204 -4742 -124 -4726
rect 54 -4780 4100 -4726
<< via1 >>
rect -812 791 -756 847
rect -646 520 -590 576
rect 1373 507 1436 566
rect -480 372 -426 426
rect 0 243 56 299
rect -189 46 -135 100
rect -812 -140 -756 -84
rect -646 -431 -590 -375
rect 7 -430 61 -376
rect 3340 -400 3396 -344
rect -491 -567 -437 -513
rect 2399 -565 2455 -509
rect 2382 -707 2436 -653
rect -190 -910 -134 -854
rect -812 -1069 -756 -1013
rect -646 -1249 -591 -1194
rect -48 -1251 9 -1194
rect -491 -1424 -437 -1370
rect 1626 -1393 1689 -1334
rect -344 -1559 -290 -1505
rect -191 -1863 -137 -1809
rect -812 -2036 -756 -1980
rect -487 -2325 -431 -2269
rect 1266 -2305 1320 -2251
rect -343 -2465 -289 -2411
rect -646 -2607 -590 -2551
rect 2 -2603 58 -2547
rect -190 -2806 -134 -2750
rect -812 -2981 -756 -2925
rect -649 -3342 -595 -3288
rect -490 -3477 -436 -3423
rect -190 -3798 -134 -3742
rect -812 -3952 -756 -3896
rect 1543 -4228 1597 -4174
rect -651 -4304 -597 -4250
rect -493 -4439 -439 -4385
rect -340 -4558 -284 -4502
rect 30 -4568 86 -4512
rect -190 -4726 -134 -4670
<< metal2 >>
rect -821 847 -747 856
rect -821 791 -812 847
rect -756 791 -747 847
rect -821 781 -747 791
rect -812 -75 -756 781
rect -655 576 -581 585
rect -655 520 -646 576
rect -590 520 -581 576
rect -655 511 -581 520
rect 200 566 1449 579
rect 200 523 1373 566
rect -822 -84 -748 -75
rect -822 -140 -812 -84
rect -756 -140 -748 -84
rect -822 -149 -748 -140
rect -812 -1005 -756 -149
rect -646 -363 -590 511
rect -489 426 -417 435
rect -489 372 -480 426
rect -426 372 -417 426
rect -489 363 -417 372
rect -658 -375 -587 -363
rect -658 -431 -646 -375
rect -590 -431 -587 -375
rect -658 -443 -587 -431
rect -825 -1013 -747 -1005
rect -825 -1069 -812 -1013
rect -756 -1069 -747 -1013
rect -825 -1081 -747 -1069
rect -812 -1969 -756 -1081
rect -646 -1187 -590 -443
rect -487 -504 -431 363
rect -12 299 68 308
rect 200 299 256 523
rect 1329 521 1373 523
rect 1360 507 1373 521
rect 1436 507 1449 566
rect 1360 492 1449 507
rect -340 243 0 299
rect 56 243 256 299
rect -500 -513 -428 -504
rect -500 -567 -491 -513
rect -437 -567 -428 -513
rect -500 -576 -428 -567
rect -658 -1194 -583 -1187
rect -658 -1249 -646 -1194
rect -591 -1249 -583 -1194
rect -658 -1260 -583 -1249
rect -823 -1980 -749 -1969
rect -823 -2036 -812 -1980
rect -756 -2036 -749 -1980
rect -823 -2046 -749 -2036
rect -812 -2912 -756 -2046
rect -646 -2541 -590 -1260
rect -487 -1361 -431 -576
rect -502 -1370 -424 -1361
rect -502 -1424 -491 -1370
rect -437 -1424 -424 -1370
rect -502 -1433 -424 -1424
rect -487 -2258 -431 -1433
rect -340 -1496 -284 243
rect -12 234 68 243
rect -198 100 -126 109
rect -198 46 -189 100
rect -135 46 -126 100
rect -198 37 -126 46
rect -190 -846 -134 37
rect 6 -312 2455 -256
rect 6 -370 62 -312
rect -21 -376 73 -370
rect -21 -430 7 -376
rect 61 -430 73 -376
rect -21 -446 73 -430
rect 2399 -501 2455 -312
rect 3333 -344 3410 -329
rect 2648 -400 3340 -344
rect 3396 -400 3410 -344
rect 2380 -509 2466 -501
rect 2380 -565 2399 -509
rect 2455 -565 2466 -509
rect 2380 -577 2466 -565
rect 2358 -652 2452 -635
rect 2648 -652 2704 -400
rect 3333 -414 3410 -400
rect 2358 -653 2704 -652
rect 2358 -707 2382 -653
rect 2436 -707 2704 -653
rect 2358 -708 2704 -707
rect 2358 -726 2452 -708
rect -201 -854 -127 -846
rect -201 -910 -190 -854
rect -134 -910 -127 -854
rect -201 -918 -127 -910
rect -354 -1505 -274 -1496
rect -354 -1559 -344 -1505
rect -290 -1559 -274 -1505
rect -354 -1569 -274 -1559
rect -499 -2269 -421 -2258
rect -499 -2325 -487 -2269
rect -431 -2325 -421 -2269
rect -499 -2334 -421 -2325
rect -662 -2551 -583 -2541
rect -662 -2607 -646 -2551
rect -590 -2607 -583 -2551
rect -662 -2617 -583 -2607
rect -842 -2925 -744 -2912
rect -842 -2981 -812 -2925
rect -756 -2981 -744 -2925
rect -842 -2999 -744 -2981
rect -812 -3884 -756 -2999
rect -646 -3278 -590 -2617
rect -664 -3288 -582 -3278
rect -664 -3342 -649 -3288
rect -595 -3342 -582 -3288
rect -664 -3351 -582 -3342
rect -825 -3896 -750 -3884
rect -825 -3952 -812 -3896
rect -756 -3952 -750 -3896
rect -825 -3967 -750 -3952
rect -646 -4241 -590 -3351
rect -487 -3413 -431 -2334
rect -340 -2401 -284 -1569
rect -190 -1800 -134 -918
rect -57 -1194 19 -1185
rect -57 -1251 -48 -1194
rect 9 -1251 130 -1194
rect -57 -1260 130 -1251
rect 73 -1332 130 -1260
rect 1613 -1332 1702 -1321
rect 73 -1334 1702 -1332
rect 73 -1389 1626 -1334
rect 1613 -1393 1626 -1389
rect 1689 -1393 1702 -1334
rect 1613 -1408 1702 -1393
rect -200 -1809 -127 -1800
rect -200 -1863 -191 -1809
rect -137 -1863 -127 -1809
rect -200 -1873 -127 -1863
rect -356 -2411 -275 -2401
rect -356 -2465 -343 -2411
rect -289 -2465 -275 -2411
rect -356 -2474 -275 -2465
rect -503 -3423 -422 -3413
rect -503 -3477 -490 -3423
rect -436 -3477 -422 -3423
rect -503 -3488 -422 -3477
rect -664 -4250 -583 -4241
rect -664 -4304 -651 -4250
rect -597 -4304 -583 -4250
rect -664 -4315 -583 -4304
rect -487 -4371 -431 -3488
rect -509 -4385 -426 -4371
rect -509 -4439 -493 -4385
rect -439 -4439 -426 -4385
rect -509 -4453 -426 -4439
rect -340 -4490 -284 -2474
rect -190 -2738 -134 -1873
rect 1253 -2250 1328 -2240
rect 258 -2251 1328 -2250
rect 258 -2305 1266 -2251
rect 1320 -2305 1328 -2251
rect 258 -2306 1328 -2305
rect -15 -2547 67 -2532
rect 258 -2547 314 -2306
rect 1253 -2315 1328 -2306
rect -15 -2603 2 -2547
rect 58 -2603 314 -2547
rect -15 -2623 67 -2603
rect -202 -2750 -121 -2738
rect -202 -2806 -190 -2750
rect -134 -2806 -121 -2750
rect -202 -2817 -121 -2806
rect -190 -3733 -134 -2817
rect -202 -3742 -127 -3733
rect -202 -3798 -190 -3742
rect -134 -3798 -127 -3742
rect -202 -3814 -127 -3798
rect -355 -4502 -274 -4490
rect -355 -4558 -340 -4502
rect -284 -4558 -274 -4502
rect -355 -4572 -274 -4558
rect -190 -4658 -134 -3814
rect 1533 -4174 1607 -4163
rect 1533 -4200 1543 -4174
rect 261 -4228 1543 -4200
rect 1597 -4228 1607 -4174
rect 261 -4255 1607 -4228
rect 261 -4256 1570 -4255
rect 19 -4512 92 -4500
rect 261 -4512 317 -4256
rect 19 -4568 30 -4512
rect 86 -4568 317 -4512
rect 19 -4580 92 -4568
rect -204 -4670 -124 -4658
rect -204 -4726 -190 -4670
rect -134 -4726 -124 -4670
rect -204 -4742 -124 -4726
use AND  AND_0
timestamp 1694585703
transform 1 0 1378 0 1 137
box -18 -137 1263 754
use AND  AND_1
timestamp 1694585703
transform 1 0 18 0 1 137
box -18 -137 1263 754
use AND  AND_2
timestamp 1694585703
transform 1 0 18 0 1 -802
box -18 -137 1263 754
use AND  AND_3
timestamp 1694585703
transform 1 0 1631 0 1 -1763
box -18 -137 1263 754
use AND  AND_4
timestamp 1694585703
transform 1 0 18 0 1 -2700
box -18 -137 1263 754
use INV_BUFF  INV_BUFF_0
timestamp 1694585882
transform 1 0 2700 0 1 0
box -90 0 858 813
use INV_BUFF  INV_BUFF_1
timestamp 1694585882
transform 1 0 1371 0 1 -939
box -90 0 858 813
use INV_BUFF  INV_BUFF_2
timestamp 1694585882
transform 1 0 2874 0 1 -1900
box -90 0 858 813
use INV_BUFF  INV_BUFF_3
timestamp 1694585882
transform 1 0 2503 0 1 -939
box -90 0 858 813
use INV_BUFF  INV_BUFF_4
timestamp 1694585882
transform 1 0 2870 0 1 -2858
box -90 0 858 813
use INV_BUFF  INV_BUFF_5
timestamp 1694585882
transform 1 0 1581 0 1 -3818
box -90 0 858 813
use INV_BUFF  INV_BUFF_6
timestamp 1694585882
transform 1 0 3303 0 1 -4780
box -90 0 858 813
use OR  OR_0
timestamp 1694585780
transform 1 0 38 0 1 -1750
box 0 -150 1566 762
use OR  OR_1
timestamp 1694585780
transform 1 0 1327 0 1 -2708
box 0 -150 1566 762
use OR  OR_2
timestamp 1694585780
transform 1 0 38 0 1 -3668
box 0 -150 1566 762
use OR  OR_3
timestamp 1694585780
transform 1 0 1610 0 1 -4630
box 0 -150 1566 762
use OR  OR_4
timestamp 1694585780
transform 1 0 38 0 1 -4630
box 0 -150 1566 762
<< labels >>
flabel metal1 34 536 34 536 0 FreeSans 640 0 0 0 B1
port 0 nsew
flabel metal1 4 398 4 398 0 FreeSans 640 0 0 0 B2
port 1 nsew
flabel via1 18 270 18 270 0 FreeSans 640 0 0 0 B3
port 2 nsew
flabel metal1 1320 841 1320 841 0 FreeSans 640 0 0 0 VDD
port 3 nsew
flabel metal1 1314 46 1314 46 0 FreeSans 640 0 0 0 VSS
port 4 nsew
flabel metal1 3562 396 3562 396 0 FreeSans 640 0 0 0 D1
port 5 nsew
flabel via1 3367 -373 3367 -373 0 FreeSans 640 0 0 0 D2
port 6 nsew
flabel metal1 3372 -543 3372 -543 0 FreeSans 640 0 0 0 D4
port 7 nsew
flabel metal1 3741 -1506 3741 -1506 0 FreeSans 640 0 0 0 D3
port 8 nsew
flabel metal1 3737 -2461 3737 -2461 0 FreeSans 640 0 0 0 D5
port 9 nsew
flabel metal1 2471 -3426 2471 -3426 0 FreeSans 640 0 0 0 D6
port 11 nsew
flabel metal1 4200 -4382 4200 -4382 0 FreeSans 640 0 0 0 D7
port 12 nsew
<< end >>
