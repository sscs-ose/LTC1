magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1143 -1267 1143 1267
<< metal2 >>
rect -143 262 143 267
rect -143 234 -138 262
rect -110 234 -76 262
rect -48 234 -14 262
rect 14 234 48 262
rect 76 234 110 262
rect 138 234 143 262
rect -143 200 143 234
rect -143 172 -138 200
rect -110 172 -76 200
rect -48 172 -14 200
rect 14 172 48 200
rect 76 172 110 200
rect 138 172 143 200
rect -143 138 143 172
rect -143 110 -138 138
rect -110 110 -76 138
rect -48 110 -14 138
rect 14 110 48 138
rect 76 110 110 138
rect 138 110 143 138
rect -143 76 143 110
rect -143 48 -138 76
rect -110 48 -76 76
rect -48 48 -14 76
rect 14 48 48 76
rect 76 48 110 76
rect 138 48 143 76
rect -143 14 143 48
rect -143 -14 -138 14
rect -110 -14 -76 14
rect -48 -14 -14 14
rect 14 -14 48 14
rect 76 -14 110 14
rect 138 -14 143 14
rect -143 -48 143 -14
rect -143 -76 -138 -48
rect -110 -76 -76 -48
rect -48 -76 -14 -48
rect 14 -76 48 -48
rect 76 -76 110 -48
rect 138 -76 143 -48
rect -143 -110 143 -76
rect -143 -138 -138 -110
rect -110 -138 -76 -110
rect -48 -138 -14 -110
rect 14 -138 48 -110
rect 76 -138 110 -110
rect 138 -138 143 -110
rect -143 -172 143 -138
rect -143 -200 -138 -172
rect -110 -200 -76 -172
rect -48 -200 -14 -172
rect 14 -200 48 -172
rect 76 -200 110 -172
rect 138 -200 143 -172
rect -143 -234 143 -200
rect -143 -262 -138 -234
rect -110 -262 -76 -234
rect -48 -262 -14 -234
rect 14 -262 48 -234
rect 76 -262 110 -234
rect 138 -262 143 -234
rect -143 -267 143 -262
<< via2 >>
rect -138 234 -110 262
rect -76 234 -48 262
rect -14 234 14 262
rect 48 234 76 262
rect 110 234 138 262
rect -138 172 -110 200
rect -76 172 -48 200
rect -14 172 14 200
rect 48 172 76 200
rect 110 172 138 200
rect -138 110 -110 138
rect -76 110 -48 138
rect -14 110 14 138
rect 48 110 76 138
rect 110 110 138 138
rect -138 48 -110 76
rect -76 48 -48 76
rect -14 48 14 76
rect 48 48 76 76
rect 110 48 138 76
rect -138 -14 -110 14
rect -76 -14 -48 14
rect -14 -14 14 14
rect 48 -14 76 14
rect 110 -14 138 14
rect -138 -76 -110 -48
rect -76 -76 -48 -48
rect -14 -76 14 -48
rect 48 -76 76 -48
rect 110 -76 138 -48
rect -138 -138 -110 -110
rect -76 -138 -48 -110
rect -14 -138 14 -110
rect 48 -138 76 -110
rect 110 -138 138 -110
rect -138 -200 -110 -172
rect -76 -200 -48 -172
rect -14 -200 14 -172
rect 48 -200 76 -172
rect 110 -200 138 -172
rect -138 -262 -110 -234
rect -76 -262 -48 -234
rect -14 -262 14 -234
rect 48 -262 76 -234
rect 110 -262 138 -234
<< metal3 >>
rect -143 262 143 267
rect -143 234 -138 262
rect -110 234 -76 262
rect -48 234 -14 262
rect 14 234 48 262
rect 76 234 110 262
rect 138 234 143 262
rect -143 200 143 234
rect -143 172 -138 200
rect -110 172 -76 200
rect -48 172 -14 200
rect 14 172 48 200
rect 76 172 110 200
rect 138 172 143 200
rect -143 138 143 172
rect -143 110 -138 138
rect -110 110 -76 138
rect -48 110 -14 138
rect 14 110 48 138
rect 76 110 110 138
rect 138 110 143 138
rect -143 76 143 110
rect -143 48 -138 76
rect -110 48 -76 76
rect -48 48 -14 76
rect 14 48 48 76
rect 76 48 110 76
rect 138 48 143 76
rect -143 14 143 48
rect -143 -14 -138 14
rect -110 -14 -76 14
rect -48 -14 -14 14
rect 14 -14 48 14
rect 76 -14 110 14
rect 138 -14 143 14
rect -143 -48 143 -14
rect -143 -76 -138 -48
rect -110 -76 -76 -48
rect -48 -76 -14 -48
rect 14 -76 48 -48
rect 76 -76 110 -48
rect 138 -76 143 -48
rect -143 -110 143 -76
rect -143 -138 -138 -110
rect -110 -138 -76 -110
rect -48 -138 -14 -110
rect 14 -138 48 -110
rect 76 -138 110 -110
rect 138 -138 143 -110
rect -143 -172 143 -138
rect -143 -200 -138 -172
rect -110 -200 -76 -172
rect -48 -200 -14 -172
rect 14 -200 48 -172
rect 76 -200 110 -172
rect 138 -200 143 -172
rect -143 -234 143 -200
rect -143 -262 -138 -234
rect -110 -262 -76 -234
rect -48 -262 -14 -234
rect 14 -262 48 -234
rect 76 -262 110 -234
rect 138 -262 143 -234
rect -143 -267 143 -262
<< end >>
