magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1745 -4880 1745 4880
<< metal3 >>
rect -745 3875 745 3880
rect -745 3847 -740 3875
rect -712 3847 -674 3875
rect -646 3847 -608 3875
rect -580 3847 -542 3875
rect -514 3847 -476 3875
rect -448 3847 -410 3875
rect -382 3847 -344 3875
rect -316 3847 -278 3875
rect -250 3847 -212 3875
rect -184 3847 -146 3875
rect -118 3847 -80 3875
rect -52 3847 -14 3875
rect 14 3847 52 3875
rect 80 3847 118 3875
rect 146 3847 184 3875
rect 212 3847 250 3875
rect 278 3847 316 3875
rect 344 3847 382 3875
rect 410 3847 448 3875
rect 476 3847 514 3875
rect 542 3847 580 3875
rect 608 3847 646 3875
rect 674 3847 712 3875
rect 740 3847 745 3875
rect -745 3809 745 3847
rect -745 3781 -740 3809
rect -712 3781 -674 3809
rect -646 3781 -608 3809
rect -580 3781 -542 3809
rect -514 3781 -476 3809
rect -448 3781 -410 3809
rect -382 3781 -344 3809
rect -316 3781 -278 3809
rect -250 3781 -212 3809
rect -184 3781 -146 3809
rect -118 3781 -80 3809
rect -52 3781 -14 3809
rect 14 3781 52 3809
rect 80 3781 118 3809
rect 146 3781 184 3809
rect 212 3781 250 3809
rect 278 3781 316 3809
rect 344 3781 382 3809
rect 410 3781 448 3809
rect 476 3781 514 3809
rect 542 3781 580 3809
rect 608 3781 646 3809
rect 674 3781 712 3809
rect 740 3781 745 3809
rect -745 3743 745 3781
rect -745 3715 -740 3743
rect -712 3715 -674 3743
rect -646 3715 -608 3743
rect -580 3715 -542 3743
rect -514 3715 -476 3743
rect -448 3715 -410 3743
rect -382 3715 -344 3743
rect -316 3715 -278 3743
rect -250 3715 -212 3743
rect -184 3715 -146 3743
rect -118 3715 -80 3743
rect -52 3715 -14 3743
rect 14 3715 52 3743
rect 80 3715 118 3743
rect 146 3715 184 3743
rect 212 3715 250 3743
rect 278 3715 316 3743
rect 344 3715 382 3743
rect 410 3715 448 3743
rect 476 3715 514 3743
rect 542 3715 580 3743
rect 608 3715 646 3743
rect 674 3715 712 3743
rect 740 3715 745 3743
rect -745 3677 745 3715
rect -745 3649 -740 3677
rect -712 3649 -674 3677
rect -646 3649 -608 3677
rect -580 3649 -542 3677
rect -514 3649 -476 3677
rect -448 3649 -410 3677
rect -382 3649 -344 3677
rect -316 3649 -278 3677
rect -250 3649 -212 3677
rect -184 3649 -146 3677
rect -118 3649 -80 3677
rect -52 3649 -14 3677
rect 14 3649 52 3677
rect 80 3649 118 3677
rect 146 3649 184 3677
rect 212 3649 250 3677
rect 278 3649 316 3677
rect 344 3649 382 3677
rect 410 3649 448 3677
rect 476 3649 514 3677
rect 542 3649 580 3677
rect 608 3649 646 3677
rect 674 3649 712 3677
rect 740 3649 745 3677
rect -745 3611 745 3649
rect -745 3583 -740 3611
rect -712 3583 -674 3611
rect -646 3583 -608 3611
rect -580 3583 -542 3611
rect -514 3583 -476 3611
rect -448 3583 -410 3611
rect -382 3583 -344 3611
rect -316 3583 -278 3611
rect -250 3583 -212 3611
rect -184 3583 -146 3611
rect -118 3583 -80 3611
rect -52 3583 -14 3611
rect 14 3583 52 3611
rect 80 3583 118 3611
rect 146 3583 184 3611
rect 212 3583 250 3611
rect 278 3583 316 3611
rect 344 3583 382 3611
rect 410 3583 448 3611
rect 476 3583 514 3611
rect 542 3583 580 3611
rect 608 3583 646 3611
rect 674 3583 712 3611
rect 740 3583 745 3611
rect -745 3545 745 3583
rect -745 3517 -740 3545
rect -712 3517 -674 3545
rect -646 3517 -608 3545
rect -580 3517 -542 3545
rect -514 3517 -476 3545
rect -448 3517 -410 3545
rect -382 3517 -344 3545
rect -316 3517 -278 3545
rect -250 3517 -212 3545
rect -184 3517 -146 3545
rect -118 3517 -80 3545
rect -52 3517 -14 3545
rect 14 3517 52 3545
rect 80 3517 118 3545
rect 146 3517 184 3545
rect 212 3517 250 3545
rect 278 3517 316 3545
rect 344 3517 382 3545
rect 410 3517 448 3545
rect 476 3517 514 3545
rect 542 3517 580 3545
rect 608 3517 646 3545
rect 674 3517 712 3545
rect 740 3517 745 3545
rect -745 3479 745 3517
rect -745 3451 -740 3479
rect -712 3451 -674 3479
rect -646 3451 -608 3479
rect -580 3451 -542 3479
rect -514 3451 -476 3479
rect -448 3451 -410 3479
rect -382 3451 -344 3479
rect -316 3451 -278 3479
rect -250 3451 -212 3479
rect -184 3451 -146 3479
rect -118 3451 -80 3479
rect -52 3451 -14 3479
rect 14 3451 52 3479
rect 80 3451 118 3479
rect 146 3451 184 3479
rect 212 3451 250 3479
rect 278 3451 316 3479
rect 344 3451 382 3479
rect 410 3451 448 3479
rect 476 3451 514 3479
rect 542 3451 580 3479
rect 608 3451 646 3479
rect 674 3451 712 3479
rect 740 3451 745 3479
rect -745 3413 745 3451
rect -745 3385 -740 3413
rect -712 3385 -674 3413
rect -646 3385 -608 3413
rect -580 3385 -542 3413
rect -514 3385 -476 3413
rect -448 3385 -410 3413
rect -382 3385 -344 3413
rect -316 3385 -278 3413
rect -250 3385 -212 3413
rect -184 3385 -146 3413
rect -118 3385 -80 3413
rect -52 3385 -14 3413
rect 14 3385 52 3413
rect 80 3385 118 3413
rect 146 3385 184 3413
rect 212 3385 250 3413
rect 278 3385 316 3413
rect 344 3385 382 3413
rect 410 3385 448 3413
rect 476 3385 514 3413
rect 542 3385 580 3413
rect 608 3385 646 3413
rect 674 3385 712 3413
rect 740 3385 745 3413
rect -745 3347 745 3385
rect -745 3319 -740 3347
rect -712 3319 -674 3347
rect -646 3319 -608 3347
rect -580 3319 -542 3347
rect -514 3319 -476 3347
rect -448 3319 -410 3347
rect -382 3319 -344 3347
rect -316 3319 -278 3347
rect -250 3319 -212 3347
rect -184 3319 -146 3347
rect -118 3319 -80 3347
rect -52 3319 -14 3347
rect 14 3319 52 3347
rect 80 3319 118 3347
rect 146 3319 184 3347
rect 212 3319 250 3347
rect 278 3319 316 3347
rect 344 3319 382 3347
rect 410 3319 448 3347
rect 476 3319 514 3347
rect 542 3319 580 3347
rect 608 3319 646 3347
rect 674 3319 712 3347
rect 740 3319 745 3347
rect -745 3281 745 3319
rect -745 3253 -740 3281
rect -712 3253 -674 3281
rect -646 3253 -608 3281
rect -580 3253 -542 3281
rect -514 3253 -476 3281
rect -448 3253 -410 3281
rect -382 3253 -344 3281
rect -316 3253 -278 3281
rect -250 3253 -212 3281
rect -184 3253 -146 3281
rect -118 3253 -80 3281
rect -52 3253 -14 3281
rect 14 3253 52 3281
rect 80 3253 118 3281
rect 146 3253 184 3281
rect 212 3253 250 3281
rect 278 3253 316 3281
rect 344 3253 382 3281
rect 410 3253 448 3281
rect 476 3253 514 3281
rect 542 3253 580 3281
rect 608 3253 646 3281
rect 674 3253 712 3281
rect 740 3253 745 3281
rect -745 3215 745 3253
rect -745 3187 -740 3215
rect -712 3187 -674 3215
rect -646 3187 -608 3215
rect -580 3187 -542 3215
rect -514 3187 -476 3215
rect -448 3187 -410 3215
rect -382 3187 -344 3215
rect -316 3187 -278 3215
rect -250 3187 -212 3215
rect -184 3187 -146 3215
rect -118 3187 -80 3215
rect -52 3187 -14 3215
rect 14 3187 52 3215
rect 80 3187 118 3215
rect 146 3187 184 3215
rect 212 3187 250 3215
rect 278 3187 316 3215
rect 344 3187 382 3215
rect 410 3187 448 3215
rect 476 3187 514 3215
rect 542 3187 580 3215
rect 608 3187 646 3215
rect 674 3187 712 3215
rect 740 3187 745 3215
rect -745 3149 745 3187
rect -745 3121 -740 3149
rect -712 3121 -674 3149
rect -646 3121 -608 3149
rect -580 3121 -542 3149
rect -514 3121 -476 3149
rect -448 3121 -410 3149
rect -382 3121 -344 3149
rect -316 3121 -278 3149
rect -250 3121 -212 3149
rect -184 3121 -146 3149
rect -118 3121 -80 3149
rect -52 3121 -14 3149
rect 14 3121 52 3149
rect 80 3121 118 3149
rect 146 3121 184 3149
rect 212 3121 250 3149
rect 278 3121 316 3149
rect 344 3121 382 3149
rect 410 3121 448 3149
rect 476 3121 514 3149
rect 542 3121 580 3149
rect 608 3121 646 3149
rect 674 3121 712 3149
rect 740 3121 745 3149
rect -745 3083 745 3121
rect -745 3055 -740 3083
rect -712 3055 -674 3083
rect -646 3055 -608 3083
rect -580 3055 -542 3083
rect -514 3055 -476 3083
rect -448 3055 -410 3083
rect -382 3055 -344 3083
rect -316 3055 -278 3083
rect -250 3055 -212 3083
rect -184 3055 -146 3083
rect -118 3055 -80 3083
rect -52 3055 -14 3083
rect 14 3055 52 3083
rect 80 3055 118 3083
rect 146 3055 184 3083
rect 212 3055 250 3083
rect 278 3055 316 3083
rect 344 3055 382 3083
rect 410 3055 448 3083
rect 476 3055 514 3083
rect 542 3055 580 3083
rect 608 3055 646 3083
rect 674 3055 712 3083
rect 740 3055 745 3083
rect -745 3017 745 3055
rect -745 2989 -740 3017
rect -712 2989 -674 3017
rect -646 2989 -608 3017
rect -580 2989 -542 3017
rect -514 2989 -476 3017
rect -448 2989 -410 3017
rect -382 2989 -344 3017
rect -316 2989 -278 3017
rect -250 2989 -212 3017
rect -184 2989 -146 3017
rect -118 2989 -80 3017
rect -52 2989 -14 3017
rect 14 2989 52 3017
rect 80 2989 118 3017
rect 146 2989 184 3017
rect 212 2989 250 3017
rect 278 2989 316 3017
rect 344 2989 382 3017
rect 410 2989 448 3017
rect 476 2989 514 3017
rect 542 2989 580 3017
rect 608 2989 646 3017
rect 674 2989 712 3017
rect 740 2989 745 3017
rect -745 2951 745 2989
rect -745 2923 -740 2951
rect -712 2923 -674 2951
rect -646 2923 -608 2951
rect -580 2923 -542 2951
rect -514 2923 -476 2951
rect -448 2923 -410 2951
rect -382 2923 -344 2951
rect -316 2923 -278 2951
rect -250 2923 -212 2951
rect -184 2923 -146 2951
rect -118 2923 -80 2951
rect -52 2923 -14 2951
rect 14 2923 52 2951
rect 80 2923 118 2951
rect 146 2923 184 2951
rect 212 2923 250 2951
rect 278 2923 316 2951
rect 344 2923 382 2951
rect 410 2923 448 2951
rect 476 2923 514 2951
rect 542 2923 580 2951
rect 608 2923 646 2951
rect 674 2923 712 2951
rect 740 2923 745 2951
rect -745 2885 745 2923
rect -745 2857 -740 2885
rect -712 2857 -674 2885
rect -646 2857 -608 2885
rect -580 2857 -542 2885
rect -514 2857 -476 2885
rect -448 2857 -410 2885
rect -382 2857 -344 2885
rect -316 2857 -278 2885
rect -250 2857 -212 2885
rect -184 2857 -146 2885
rect -118 2857 -80 2885
rect -52 2857 -14 2885
rect 14 2857 52 2885
rect 80 2857 118 2885
rect 146 2857 184 2885
rect 212 2857 250 2885
rect 278 2857 316 2885
rect 344 2857 382 2885
rect 410 2857 448 2885
rect 476 2857 514 2885
rect 542 2857 580 2885
rect 608 2857 646 2885
rect 674 2857 712 2885
rect 740 2857 745 2885
rect -745 2819 745 2857
rect -745 2791 -740 2819
rect -712 2791 -674 2819
rect -646 2791 -608 2819
rect -580 2791 -542 2819
rect -514 2791 -476 2819
rect -448 2791 -410 2819
rect -382 2791 -344 2819
rect -316 2791 -278 2819
rect -250 2791 -212 2819
rect -184 2791 -146 2819
rect -118 2791 -80 2819
rect -52 2791 -14 2819
rect 14 2791 52 2819
rect 80 2791 118 2819
rect 146 2791 184 2819
rect 212 2791 250 2819
rect 278 2791 316 2819
rect 344 2791 382 2819
rect 410 2791 448 2819
rect 476 2791 514 2819
rect 542 2791 580 2819
rect 608 2791 646 2819
rect 674 2791 712 2819
rect 740 2791 745 2819
rect -745 2753 745 2791
rect -745 2725 -740 2753
rect -712 2725 -674 2753
rect -646 2725 -608 2753
rect -580 2725 -542 2753
rect -514 2725 -476 2753
rect -448 2725 -410 2753
rect -382 2725 -344 2753
rect -316 2725 -278 2753
rect -250 2725 -212 2753
rect -184 2725 -146 2753
rect -118 2725 -80 2753
rect -52 2725 -14 2753
rect 14 2725 52 2753
rect 80 2725 118 2753
rect 146 2725 184 2753
rect 212 2725 250 2753
rect 278 2725 316 2753
rect 344 2725 382 2753
rect 410 2725 448 2753
rect 476 2725 514 2753
rect 542 2725 580 2753
rect 608 2725 646 2753
rect 674 2725 712 2753
rect 740 2725 745 2753
rect -745 2687 745 2725
rect -745 2659 -740 2687
rect -712 2659 -674 2687
rect -646 2659 -608 2687
rect -580 2659 -542 2687
rect -514 2659 -476 2687
rect -448 2659 -410 2687
rect -382 2659 -344 2687
rect -316 2659 -278 2687
rect -250 2659 -212 2687
rect -184 2659 -146 2687
rect -118 2659 -80 2687
rect -52 2659 -14 2687
rect 14 2659 52 2687
rect 80 2659 118 2687
rect 146 2659 184 2687
rect 212 2659 250 2687
rect 278 2659 316 2687
rect 344 2659 382 2687
rect 410 2659 448 2687
rect 476 2659 514 2687
rect 542 2659 580 2687
rect 608 2659 646 2687
rect 674 2659 712 2687
rect 740 2659 745 2687
rect -745 2621 745 2659
rect -745 2593 -740 2621
rect -712 2593 -674 2621
rect -646 2593 -608 2621
rect -580 2593 -542 2621
rect -514 2593 -476 2621
rect -448 2593 -410 2621
rect -382 2593 -344 2621
rect -316 2593 -278 2621
rect -250 2593 -212 2621
rect -184 2593 -146 2621
rect -118 2593 -80 2621
rect -52 2593 -14 2621
rect 14 2593 52 2621
rect 80 2593 118 2621
rect 146 2593 184 2621
rect 212 2593 250 2621
rect 278 2593 316 2621
rect 344 2593 382 2621
rect 410 2593 448 2621
rect 476 2593 514 2621
rect 542 2593 580 2621
rect 608 2593 646 2621
rect 674 2593 712 2621
rect 740 2593 745 2621
rect -745 2555 745 2593
rect -745 2527 -740 2555
rect -712 2527 -674 2555
rect -646 2527 -608 2555
rect -580 2527 -542 2555
rect -514 2527 -476 2555
rect -448 2527 -410 2555
rect -382 2527 -344 2555
rect -316 2527 -278 2555
rect -250 2527 -212 2555
rect -184 2527 -146 2555
rect -118 2527 -80 2555
rect -52 2527 -14 2555
rect 14 2527 52 2555
rect 80 2527 118 2555
rect 146 2527 184 2555
rect 212 2527 250 2555
rect 278 2527 316 2555
rect 344 2527 382 2555
rect 410 2527 448 2555
rect 476 2527 514 2555
rect 542 2527 580 2555
rect 608 2527 646 2555
rect 674 2527 712 2555
rect 740 2527 745 2555
rect -745 2489 745 2527
rect -745 2461 -740 2489
rect -712 2461 -674 2489
rect -646 2461 -608 2489
rect -580 2461 -542 2489
rect -514 2461 -476 2489
rect -448 2461 -410 2489
rect -382 2461 -344 2489
rect -316 2461 -278 2489
rect -250 2461 -212 2489
rect -184 2461 -146 2489
rect -118 2461 -80 2489
rect -52 2461 -14 2489
rect 14 2461 52 2489
rect 80 2461 118 2489
rect 146 2461 184 2489
rect 212 2461 250 2489
rect 278 2461 316 2489
rect 344 2461 382 2489
rect 410 2461 448 2489
rect 476 2461 514 2489
rect 542 2461 580 2489
rect 608 2461 646 2489
rect 674 2461 712 2489
rect 740 2461 745 2489
rect -745 2423 745 2461
rect -745 2395 -740 2423
rect -712 2395 -674 2423
rect -646 2395 -608 2423
rect -580 2395 -542 2423
rect -514 2395 -476 2423
rect -448 2395 -410 2423
rect -382 2395 -344 2423
rect -316 2395 -278 2423
rect -250 2395 -212 2423
rect -184 2395 -146 2423
rect -118 2395 -80 2423
rect -52 2395 -14 2423
rect 14 2395 52 2423
rect 80 2395 118 2423
rect 146 2395 184 2423
rect 212 2395 250 2423
rect 278 2395 316 2423
rect 344 2395 382 2423
rect 410 2395 448 2423
rect 476 2395 514 2423
rect 542 2395 580 2423
rect 608 2395 646 2423
rect 674 2395 712 2423
rect 740 2395 745 2423
rect -745 2357 745 2395
rect -745 2329 -740 2357
rect -712 2329 -674 2357
rect -646 2329 -608 2357
rect -580 2329 -542 2357
rect -514 2329 -476 2357
rect -448 2329 -410 2357
rect -382 2329 -344 2357
rect -316 2329 -278 2357
rect -250 2329 -212 2357
rect -184 2329 -146 2357
rect -118 2329 -80 2357
rect -52 2329 -14 2357
rect 14 2329 52 2357
rect 80 2329 118 2357
rect 146 2329 184 2357
rect 212 2329 250 2357
rect 278 2329 316 2357
rect 344 2329 382 2357
rect 410 2329 448 2357
rect 476 2329 514 2357
rect 542 2329 580 2357
rect 608 2329 646 2357
rect 674 2329 712 2357
rect 740 2329 745 2357
rect -745 2291 745 2329
rect -745 2263 -740 2291
rect -712 2263 -674 2291
rect -646 2263 -608 2291
rect -580 2263 -542 2291
rect -514 2263 -476 2291
rect -448 2263 -410 2291
rect -382 2263 -344 2291
rect -316 2263 -278 2291
rect -250 2263 -212 2291
rect -184 2263 -146 2291
rect -118 2263 -80 2291
rect -52 2263 -14 2291
rect 14 2263 52 2291
rect 80 2263 118 2291
rect 146 2263 184 2291
rect 212 2263 250 2291
rect 278 2263 316 2291
rect 344 2263 382 2291
rect 410 2263 448 2291
rect 476 2263 514 2291
rect 542 2263 580 2291
rect 608 2263 646 2291
rect 674 2263 712 2291
rect 740 2263 745 2291
rect -745 2225 745 2263
rect -745 2197 -740 2225
rect -712 2197 -674 2225
rect -646 2197 -608 2225
rect -580 2197 -542 2225
rect -514 2197 -476 2225
rect -448 2197 -410 2225
rect -382 2197 -344 2225
rect -316 2197 -278 2225
rect -250 2197 -212 2225
rect -184 2197 -146 2225
rect -118 2197 -80 2225
rect -52 2197 -14 2225
rect 14 2197 52 2225
rect 80 2197 118 2225
rect 146 2197 184 2225
rect 212 2197 250 2225
rect 278 2197 316 2225
rect 344 2197 382 2225
rect 410 2197 448 2225
rect 476 2197 514 2225
rect 542 2197 580 2225
rect 608 2197 646 2225
rect 674 2197 712 2225
rect 740 2197 745 2225
rect -745 2159 745 2197
rect -745 2131 -740 2159
rect -712 2131 -674 2159
rect -646 2131 -608 2159
rect -580 2131 -542 2159
rect -514 2131 -476 2159
rect -448 2131 -410 2159
rect -382 2131 -344 2159
rect -316 2131 -278 2159
rect -250 2131 -212 2159
rect -184 2131 -146 2159
rect -118 2131 -80 2159
rect -52 2131 -14 2159
rect 14 2131 52 2159
rect 80 2131 118 2159
rect 146 2131 184 2159
rect 212 2131 250 2159
rect 278 2131 316 2159
rect 344 2131 382 2159
rect 410 2131 448 2159
rect 476 2131 514 2159
rect 542 2131 580 2159
rect 608 2131 646 2159
rect 674 2131 712 2159
rect 740 2131 745 2159
rect -745 2093 745 2131
rect -745 2065 -740 2093
rect -712 2065 -674 2093
rect -646 2065 -608 2093
rect -580 2065 -542 2093
rect -514 2065 -476 2093
rect -448 2065 -410 2093
rect -382 2065 -344 2093
rect -316 2065 -278 2093
rect -250 2065 -212 2093
rect -184 2065 -146 2093
rect -118 2065 -80 2093
rect -52 2065 -14 2093
rect 14 2065 52 2093
rect 80 2065 118 2093
rect 146 2065 184 2093
rect 212 2065 250 2093
rect 278 2065 316 2093
rect 344 2065 382 2093
rect 410 2065 448 2093
rect 476 2065 514 2093
rect 542 2065 580 2093
rect 608 2065 646 2093
rect 674 2065 712 2093
rect 740 2065 745 2093
rect -745 2027 745 2065
rect -745 1999 -740 2027
rect -712 1999 -674 2027
rect -646 1999 -608 2027
rect -580 1999 -542 2027
rect -514 1999 -476 2027
rect -448 1999 -410 2027
rect -382 1999 -344 2027
rect -316 1999 -278 2027
rect -250 1999 -212 2027
rect -184 1999 -146 2027
rect -118 1999 -80 2027
rect -52 1999 -14 2027
rect 14 1999 52 2027
rect 80 1999 118 2027
rect 146 1999 184 2027
rect 212 1999 250 2027
rect 278 1999 316 2027
rect 344 1999 382 2027
rect 410 1999 448 2027
rect 476 1999 514 2027
rect 542 1999 580 2027
rect 608 1999 646 2027
rect 674 1999 712 2027
rect 740 1999 745 2027
rect -745 1961 745 1999
rect -745 1933 -740 1961
rect -712 1933 -674 1961
rect -646 1933 -608 1961
rect -580 1933 -542 1961
rect -514 1933 -476 1961
rect -448 1933 -410 1961
rect -382 1933 -344 1961
rect -316 1933 -278 1961
rect -250 1933 -212 1961
rect -184 1933 -146 1961
rect -118 1933 -80 1961
rect -52 1933 -14 1961
rect 14 1933 52 1961
rect 80 1933 118 1961
rect 146 1933 184 1961
rect 212 1933 250 1961
rect 278 1933 316 1961
rect 344 1933 382 1961
rect 410 1933 448 1961
rect 476 1933 514 1961
rect 542 1933 580 1961
rect 608 1933 646 1961
rect 674 1933 712 1961
rect 740 1933 745 1961
rect -745 1895 745 1933
rect -745 1867 -740 1895
rect -712 1867 -674 1895
rect -646 1867 -608 1895
rect -580 1867 -542 1895
rect -514 1867 -476 1895
rect -448 1867 -410 1895
rect -382 1867 -344 1895
rect -316 1867 -278 1895
rect -250 1867 -212 1895
rect -184 1867 -146 1895
rect -118 1867 -80 1895
rect -52 1867 -14 1895
rect 14 1867 52 1895
rect 80 1867 118 1895
rect 146 1867 184 1895
rect 212 1867 250 1895
rect 278 1867 316 1895
rect 344 1867 382 1895
rect 410 1867 448 1895
rect 476 1867 514 1895
rect 542 1867 580 1895
rect 608 1867 646 1895
rect 674 1867 712 1895
rect 740 1867 745 1895
rect -745 1829 745 1867
rect -745 1801 -740 1829
rect -712 1801 -674 1829
rect -646 1801 -608 1829
rect -580 1801 -542 1829
rect -514 1801 -476 1829
rect -448 1801 -410 1829
rect -382 1801 -344 1829
rect -316 1801 -278 1829
rect -250 1801 -212 1829
rect -184 1801 -146 1829
rect -118 1801 -80 1829
rect -52 1801 -14 1829
rect 14 1801 52 1829
rect 80 1801 118 1829
rect 146 1801 184 1829
rect 212 1801 250 1829
rect 278 1801 316 1829
rect 344 1801 382 1829
rect 410 1801 448 1829
rect 476 1801 514 1829
rect 542 1801 580 1829
rect 608 1801 646 1829
rect 674 1801 712 1829
rect 740 1801 745 1829
rect -745 1763 745 1801
rect -745 1735 -740 1763
rect -712 1735 -674 1763
rect -646 1735 -608 1763
rect -580 1735 -542 1763
rect -514 1735 -476 1763
rect -448 1735 -410 1763
rect -382 1735 -344 1763
rect -316 1735 -278 1763
rect -250 1735 -212 1763
rect -184 1735 -146 1763
rect -118 1735 -80 1763
rect -52 1735 -14 1763
rect 14 1735 52 1763
rect 80 1735 118 1763
rect 146 1735 184 1763
rect 212 1735 250 1763
rect 278 1735 316 1763
rect 344 1735 382 1763
rect 410 1735 448 1763
rect 476 1735 514 1763
rect 542 1735 580 1763
rect 608 1735 646 1763
rect 674 1735 712 1763
rect 740 1735 745 1763
rect -745 1697 745 1735
rect -745 1669 -740 1697
rect -712 1669 -674 1697
rect -646 1669 -608 1697
rect -580 1669 -542 1697
rect -514 1669 -476 1697
rect -448 1669 -410 1697
rect -382 1669 -344 1697
rect -316 1669 -278 1697
rect -250 1669 -212 1697
rect -184 1669 -146 1697
rect -118 1669 -80 1697
rect -52 1669 -14 1697
rect 14 1669 52 1697
rect 80 1669 118 1697
rect 146 1669 184 1697
rect 212 1669 250 1697
rect 278 1669 316 1697
rect 344 1669 382 1697
rect 410 1669 448 1697
rect 476 1669 514 1697
rect 542 1669 580 1697
rect 608 1669 646 1697
rect 674 1669 712 1697
rect 740 1669 745 1697
rect -745 1631 745 1669
rect -745 1603 -740 1631
rect -712 1603 -674 1631
rect -646 1603 -608 1631
rect -580 1603 -542 1631
rect -514 1603 -476 1631
rect -448 1603 -410 1631
rect -382 1603 -344 1631
rect -316 1603 -278 1631
rect -250 1603 -212 1631
rect -184 1603 -146 1631
rect -118 1603 -80 1631
rect -52 1603 -14 1631
rect 14 1603 52 1631
rect 80 1603 118 1631
rect 146 1603 184 1631
rect 212 1603 250 1631
rect 278 1603 316 1631
rect 344 1603 382 1631
rect 410 1603 448 1631
rect 476 1603 514 1631
rect 542 1603 580 1631
rect 608 1603 646 1631
rect 674 1603 712 1631
rect 740 1603 745 1631
rect -745 1565 745 1603
rect -745 1537 -740 1565
rect -712 1537 -674 1565
rect -646 1537 -608 1565
rect -580 1537 -542 1565
rect -514 1537 -476 1565
rect -448 1537 -410 1565
rect -382 1537 -344 1565
rect -316 1537 -278 1565
rect -250 1537 -212 1565
rect -184 1537 -146 1565
rect -118 1537 -80 1565
rect -52 1537 -14 1565
rect 14 1537 52 1565
rect 80 1537 118 1565
rect 146 1537 184 1565
rect 212 1537 250 1565
rect 278 1537 316 1565
rect 344 1537 382 1565
rect 410 1537 448 1565
rect 476 1537 514 1565
rect 542 1537 580 1565
rect 608 1537 646 1565
rect 674 1537 712 1565
rect 740 1537 745 1565
rect -745 1499 745 1537
rect -745 1471 -740 1499
rect -712 1471 -674 1499
rect -646 1471 -608 1499
rect -580 1471 -542 1499
rect -514 1471 -476 1499
rect -448 1471 -410 1499
rect -382 1471 -344 1499
rect -316 1471 -278 1499
rect -250 1471 -212 1499
rect -184 1471 -146 1499
rect -118 1471 -80 1499
rect -52 1471 -14 1499
rect 14 1471 52 1499
rect 80 1471 118 1499
rect 146 1471 184 1499
rect 212 1471 250 1499
rect 278 1471 316 1499
rect 344 1471 382 1499
rect 410 1471 448 1499
rect 476 1471 514 1499
rect 542 1471 580 1499
rect 608 1471 646 1499
rect 674 1471 712 1499
rect 740 1471 745 1499
rect -745 1433 745 1471
rect -745 1405 -740 1433
rect -712 1405 -674 1433
rect -646 1405 -608 1433
rect -580 1405 -542 1433
rect -514 1405 -476 1433
rect -448 1405 -410 1433
rect -382 1405 -344 1433
rect -316 1405 -278 1433
rect -250 1405 -212 1433
rect -184 1405 -146 1433
rect -118 1405 -80 1433
rect -52 1405 -14 1433
rect 14 1405 52 1433
rect 80 1405 118 1433
rect 146 1405 184 1433
rect 212 1405 250 1433
rect 278 1405 316 1433
rect 344 1405 382 1433
rect 410 1405 448 1433
rect 476 1405 514 1433
rect 542 1405 580 1433
rect 608 1405 646 1433
rect 674 1405 712 1433
rect 740 1405 745 1433
rect -745 1367 745 1405
rect -745 1339 -740 1367
rect -712 1339 -674 1367
rect -646 1339 -608 1367
rect -580 1339 -542 1367
rect -514 1339 -476 1367
rect -448 1339 -410 1367
rect -382 1339 -344 1367
rect -316 1339 -278 1367
rect -250 1339 -212 1367
rect -184 1339 -146 1367
rect -118 1339 -80 1367
rect -52 1339 -14 1367
rect 14 1339 52 1367
rect 80 1339 118 1367
rect 146 1339 184 1367
rect 212 1339 250 1367
rect 278 1339 316 1367
rect 344 1339 382 1367
rect 410 1339 448 1367
rect 476 1339 514 1367
rect 542 1339 580 1367
rect 608 1339 646 1367
rect 674 1339 712 1367
rect 740 1339 745 1367
rect -745 1301 745 1339
rect -745 1273 -740 1301
rect -712 1273 -674 1301
rect -646 1273 -608 1301
rect -580 1273 -542 1301
rect -514 1273 -476 1301
rect -448 1273 -410 1301
rect -382 1273 -344 1301
rect -316 1273 -278 1301
rect -250 1273 -212 1301
rect -184 1273 -146 1301
rect -118 1273 -80 1301
rect -52 1273 -14 1301
rect 14 1273 52 1301
rect 80 1273 118 1301
rect 146 1273 184 1301
rect 212 1273 250 1301
rect 278 1273 316 1301
rect 344 1273 382 1301
rect 410 1273 448 1301
rect 476 1273 514 1301
rect 542 1273 580 1301
rect 608 1273 646 1301
rect 674 1273 712 1301
rect 740 1273 745 1301
rect -745 1235 745 1273
rect -745 1207 -740 1235
rect -712 1207 -674 1235
rect -646 1207 -608 1235
rect -580 1207 -542 1235
rect -514 1207 -476 1235
rect -448 1207 -410 1235
rect -382 1207 -344 1235
rect -316 1207 -278 1235
rect -250 1207 -212 1235
rect -184 1207 -146 1235
rect -118 1207 -80 1235
rect -52 1207 -14 1235
rect 14 1207 52 1235
rect 80 1207 118 1235
rect 146 1207 184 1235
rect 212 1207 250 1235
rect 278 1207 316 1235
rect 344 1207 382 1235
rect 410 1207 448 1235
rect 476 1207 514 1235
rect 542 1207 580 1235
rect 608 1207 646 1235
rect 674 1207 712 1235
rect 740 1207 745 1235
rect -745 1169 745 1207
rect -745 1141 -740 1169
rect -712 1141 -674 1169
rect -646 1141 -608 1169
rect -580 1141 -542 1169
rect -514 1141 -476 1169
rect -448 1141 -410 1169
rect -382 1141 -344 1169
rect -316 1141 -278 1169
rect -250 1141 -212 1169
rect -184 1141 -146 1169
rect -118 1141 -80 1169
rect -52 1141 -14 1169
rect 14 1141 52 1169
rect 80 1141 118 1169
rect 146 1141 184 1169
rect 212 1141 250 1169
rect 278 1141 316 1169
rect 344 1141 382 1169
rect 410 1141 448 1169
rect 476 1141 514 1169
rect 542 1141 580 1169
rect 608 1141 646 1169
rect 674 1141 712 1169
rect 740 1141 745 1169
rect -745 1103 745 1141
rect -745 1075 -740 1103
rect -712 1075 -674 1103
rect -646 1075 -608 1103
rect -580 1075 -542 1103
rect -514 1075 -476 1103
rect -448 1075 -410 1103
rect -382 1075 -344 1103
rect -316 1075 -278 1103
rect -250 1075 -212 1103
rect -184 1075 -146 1103
rect -118 1075 -80 1103
rect -52 1075 -14 1103
rect 14 1075 52 1103
rect 80 1075 118 1103
rect 146 1075 184 1103
rect 212 1075 250 1103
rect 278 1075 316 1103
rect 344 1075 382 1103
rect 410 1075 448 1103
rect 476 1075 514 1103
rect 542 1075 580 1103
rect 608 1075 646 1103
rect 674 1075 712 1103
rect 740 1075 745 1103
rect -745 1037 745 1075
rect -745 1009 -740 1037
rect -712 1009 -674 1037
rect -646 1009 -608 1037
rect -580 1009 -542 1037
rect -514 1009 -476 1037
rect -448 1009 -410 1037
rect -382 1009 -344 1037
rect -316 1009 -278 1037
rect -250 1009 -212 1037
rect -184 1009 -146 1037
rect -118 1009 -80 1037
rect -52 1009 -14 1037
rect 14 1009 52 1037
rect 80 1009 118 1037
rect 146 1009 184 1037
rect 212 1009 250 1037
rect 278 1009 316 1037
rect 344 1009 382 1037
rect 410 1009 448 1037
rect 476 1009 514 1037
rect 542 1009 580 1037
rect 608 1009 646 1037
rect 674 1009 712 1037
rect 740 1009 745 1037
rect -745 971 745 1009
rect -745 943 -740 971
rect -712 943 -674 971
rect -646 943 -608 971
rect -580 943 -542 971
rect -514 943 -476 971
rect -448 943 -410 971
rect -382 943 -344 971
rect -316 943 -278 971
rect -250 943 -212 971
rect -184 943 -146 971
rect -118 943 -80 971
rect -52 943 -14 971
rect 14 943 52 971
rect 80 943 118 971
rect 146 943 184 971
rect 212 943 250 971
rect 278 943 316 971
rect 344 943 382 971
rect 410 943 448 971
rect 476 943 514 971
rect 542 943 580 971
rect 608 943 646 971
rect 674 943 712 971
rect 740 943 745 971
rect -745 905 745 943
rect -745 877 -740 905
rect -712 877 -674 905
rect -646 877 -608 905
rect -580 877 -542 905
rect -514 877 -476 905
rect -448 877 -410 905
rect -382 877 -344 905
rect -316 877 -278 905
rect -250 877 -212 905
rect -184 877 -146 905
rect -118 877 -80 905
rect -52 877 -14 905
rect 14 877 52 905
rect 80 877 118 905
rect 146 877 184 905
rect 212 877 250 905
rect 278 877 316 905
rect 344 877 382 905
rect 410 877 448 905
rect 476 877 514 905
rect 542 877 580 905
rect 608 877 646 905
rect 674 877 712 905
rect 740 877 745 905
rect -745 839 745 877
rect -745 811 -740 839
rect -712 811 -674 839
rect -646 811 -608 839
rect -580 811 -542 839
rect -514 811 -476 839
rect -448 811 -410 839
rect -382 811 -344 839
rect -316 811 -278 839
rect -250 811 -212 839
rect -184 811 -146 839
rect -118 811 -80 839
rect -52 811 -14 839
rect 14 811 52 839
rect 80 811 118 839
rect 146 811 184 839
rect 212 811 250 839
rect 278 811 316 839
rect 344 811 382 839
rect 410 811 448 839
rect 476 811 514 839
rect 542 811 580 839
rect 608 811 646 839
rect 674 811 712 839
rect 740 811 745 839
rect -745 773 745 811
rect -745 745 -740 773
rect -712 745 -674 773
rect -646 745 -608 773
rect -580 745 -542 773
rect -514 745 -476 773
rect -448 745 -410 773
rect -382 745 -344 773
rect -316 745 -278 773
rect -250 745 -212 773
rect -184 745 -146 773
rect -118 745 -80 773
rect -52 745 -14 773
rect 14 745 52 773
rect 80 745 118 773
rect 146 745 184 773
rect 212 745 250 773
rect 278 745 316 773
rect 344 745 382 773
rect 410 745 448 773
rect 476 745 514 773
rect 542 745 580 773
rect 608 745 646 773
rect 674 745 712 773
rect 740 745 745 773
rect -745 707 745 745
rect -745 679 -740 707
rect -712 679 -674 707
rect -646 679 -608 707
rect -580 679 -542 707
rect -514 679 -476 707
rect -448 679 -410 707
rect -382 679 -344 707
rect -316 679 -278 707
rect -250 679 -212 707
rect -184 679 -146 707
rect -118 679 -80 707
rect -52 679 -14 707
rect 14 679 52 707
rect 80 679 118 707
rect 146 679 184 707
rect 212 679 250 707
rect 278 679 316 707
rect 344 679 382 707
rect 410 679 448 707
rect 476 679 514 707
rect 542 679 580 707
rect 608 679 646 707
rect 674 679 712 707
rect 740 679 745 707
rect -745 641 745 679
rect -745 613 -740 641
rect -712 613 -674 641
rect -646 613 -608 641
rect -580 613 -542 641
rect -514 613 -476 641
rect -448 613 -410 641
rect -382 613 -344 641
rect -316 613 -278 641
rect -250 613 -212 641
rect -184 613 -146 641
rect -118 613 -80 641
rect -52 613 -14 641
rect 14 613 52 641
rect 80 613 118 641
rect 146 613 184 641
rect 212 613 250 641
rect 278 613 316 641
rect 344 613 382 641
rect 410 613 448 641
rect 476 613 514 641
rect 542 613 580 641
rect 608 613 646 641
rect 674 613 712 641
rect 740 613 745 641
rect -745 575 745 613
rect -745 547 -740 575
rect -712 547 -674 575
rect -646 547 -608 575
rect -580 547 -542 575
rect -514 547 -476 575
rect -448 547 -410 575
rect -382 547 -344 575
rect -316 547 -278 575
rect -250 547 -212 575
rect -184 547 -146 575
rect -118 547 -80 575
rect -52 547 -14 575
rect 14 547 52 575
rect 80 547 118 575
rect 146 547 184 575
rect 212 547 250 575
rect 278 547 316 575
rect 344 547 382 575
rect 410 547 448 575
rect 476 547 514 575
rect 542 547 580 575
rect 608 547 646 575
rect 674 547 712 575
rect 740 547 745 575
rect -745 509 745 547
rect -745 481 -740 509
rect -712 481 -674 509
rect -646 481 -608 509
rect -580 481 -542 509
rect -514 481 -476 509
rect -448 481 -410 509
rect -382 481 -344 509
rect -316 481 -278 509
rect -250 481 -212 509
rect -184 481 -146 509
rect -118 481 -80 509
rect -52 481 -14 509
rect 14 481 52 509
rect 80 481 118 509
rect 146 481 184 509
rect 212 481 250 509
rect 278 481 316 509
rect 344 481 382 509
rect 410 481 448 509
rect 476 481 514 509
rect 542 481 580 509
rect 608 481 646 509
rect 674 481 712 509
rect 740 481 745 509
rect -745 443 745 481
rect -745 415 -740 443
rect -712 415 -674 443
rect -646 415 -608 443
rect -580 415 -542 443
rect -514 415 -476 443
rect -448 415 -410 443
rect -382 415 -344 443
rect -316 415 -278 443
rect -250 415 -212 443
rect -184 415 -146 443
rect -118 415 -80 443
rect -52 415 -14 443
rect 14 415 52 443
rect 80 415 118 443
rect 146 415 184 443
rect 212 415 250 443
rect 278 415 316 443
rect 344 415 382 443
rect 410 415 448 443
rect 476 415 514 443
rect 542 415 580 443
rect 608 415 646 443
rect 674 415 712 443
rect 740 415 745 443
rect -745 377 745 415
rect -745 349 -740 377
rect -712 349 -674 377
rect -646 349 -608 377
rect -580 349 -542 377
rect -514 349 -476 377
rect -448 349 -410 377
rect -382 349 -344 377
rect -316 349 -278 377
rect -250 349 -212 377
rect -184 349 -146 377
rect -118 349 -80 377
rect -52 349 -14 377
rect 14 349 52 377
rect 80 349 118 377
rect 146 349 184 377
rect 212 349 250 377
rect 278 349 316 377
rect 344 349 382 377
rect 410 349 448 377
rect 476 349 514 377
rect 542 349 580 377
rect 608 349 646 377
rect 674 349 712 377
rect 740 349 745 377
rect -745 311 745 349
rect -745 283 -740 311
rect -712 283 -674 311
rect -646 283 -608 311
rect -580 283 -542 311
rect -514 283 -476 311
rect -448 283 -410 311
rect -382 283 -344 311
rect -316 283 -278 311
rect -250 283 -212 311
rect -184 283 -146 311
rect -118 283 -80 311
rect -52 283 -14 311
rect 14 283 52 311
rect 80 283 118 311
rect 146 283 184 311
rect 212 283 250 311
rect 278 283 316 311
rect 344 283 382 311
rect 410 283 448 311
rect 476 283 514 311
rect 542 283 580 311
rect 608 283 646 311
rect 674 283 712 311
rect 740 283 745 311
rect -745 245 745 283
rect -745 217 -740 245
rect -712 217 -674 245
rect -646 217 -608 245
rect -580 217 -542 245
rect -514 217 -476 245
rect -448 217 -410 245
rect -382 217 -344 245
rect -316 217 -278 245
rect -250 217 -212 245
rect -184 217 -146 245
rect -118 217 -80 245
rect -52 217 -14 245
rect 14 217 52 245
rect 80 217 118 245
rect 146 217 184 245
rect 212 217 250 245
rect 278 217 316 245
rect 344 217 382 245
rect 410 217 448 245
rect 476 217 514 245
rect 542 217 580 245
rect 608 217 646 245
rect 674 217 712 245
rect 740 217 745 245
rect -745 179 745 217
rect -745 151 -740 179
rect -712 151 -674 179
rect -646 151 -608 179
rect -580 151 -542 179
rect -514 151 -476 179
rect -448 151 -410 179
rect -382 151 -344 179
rect -316 151 -278 179
rect -250 151 -212 179
rect -184 151 -146 179
rect -118 151 -80 179
rect -52 151 -14 179
rect 14 151 52 179
rect 80 151 118 179
rect 146 151 184 179
rect 212 151 250 179
rect 278 151 316 179
rect 344 151 382 179
rect 410 151 448 179
rect 476 151 514 179
rect 542 151 580 179
rect 608 151 646 179
rect 674 151 712 179
rect 740 151 745 179
rect -745 113 745 151
rect -745 85 -740 113
rect -712 85 -674 113
rect -646 85 -608 113
rect -580 85 -542 113
rect -514 85 -476 113
rect -448 85 -410 113
rect -382 85 -344 113
rect -316 85 -278 113
rect -250 85 -212 113
rect -184 85 -146 113
rect -118 85 -80 113
rect -52 85 -14 113
rect 14 85 52 113
rect 80 85 118 113
rect 146 85 184 113
rect 212 85 250 113
rect 278 85 316 113
rect 344 85 382 113
rect 410 85 448 113
rect 476 85 514 113
rect 542 85 580 113
rect 608 85 646 113
rect 674 85 712 113
rect 740 85 745 113
rect -745 47 745 85
rect -745 19 -740 47
rect -712 19 -674 47
rect -646 19 -608 47
rect -580 19 -542 47
rect -514 19 -476 47
rect -448 19 -410 47
rect -382 19 -344 47
rect -316 19 -278 47
rect -250 19 -212 47
rect -184 19 -146 47
rect -118 19 -80 47
rect -52 19 -14 47
rect 14 19 52 47
rect 80 19 118 47
rect 146 19 184 47
rect 212 19 250 47
rect 278 19 316 47
rect 344 19 382 47
rect 410 19 448 47
rect 476 19 514 47
rect 542 19 580 47
rect 608 19 646 47
rect 674 19 712 47
rect 740 19 745 47
rect -745 -19 745 19
rect -745 -47 -740 -19
rect -712 -47 -674 -19
rect -646 -47 -608 -19
rect -580 -47 -542 -19
rect -514 -47 -476 -19
rect -448 -47 -410 -19
rect -382 -47 -344 -19
rect -316 -47 -278 -19
rect -250 -47 -212 -19
rect -184 -47 -146 -19
rect -118 -47 -80 -19
rect -52 -47 -14 -19
rect 14 -47 52 -19
rect 80 -47 118 -19
rect 146 -47 184 -19
rect 212 -47 250 -19
rect 278 -47 316 -19
rect 344 -47 382 -19
rect 410 -47 448 -19
rect 476 -47 514 -19
rect 542 -47 580 -19
rect 608 -47 646 -19
rect 674 -47 712 -19
rect 740 -47 745 -19
rect -745 -85 745 -47
rect -745 -113 -740 -85
rect -712 -113 -674 -85
rect -646 -113 -608 -85
rect -580 -113 -542 -85
rect -514 -113 -476 -85
rect -448 -113 -410 -85
rect -382 -113 -344 -85
rect -316 -113 -278 -85
rect -250 -113 -212 -85
rect -184 -113 -146 -85
rect -118 -113 -80 -85
rect -52 -113 -14 -85
rect 14 -113 52 -85
rect 80 -113 118 -85
rect 146 -113 184 -85
rect 212 -113 250 -85
rect 278 -113 316 -85
rect 344 -113 382 -85
rect 410 -113 448 -85
rect 476 -113 514 -85
rect 542 -113 580 -85
rect 608 -113 646 -85
rect 674 -113 712 -85
rect 740 -113 745 -85
rect -745 -151 745 -113
rect -745 -179 -740 -151
rect -712 -179 -674 -151
rect -646 -179 -608 -151
rect -580 -179 -542 -151
rect -514 -179 -476 -151
rect -448 -179 -410 -151
rect -382 -179 -344 -151
rect -316 -179 -278 -151
rect -250 -179 -212 -151
rect -184 -179 -146 -151
rect -118 -179 -80 -151
rect -52 -179 -14 -151
rect 14 -179 52 -151
rect 80 -179 118 -151
rect 146 -179 184 -151
rect 212 -179 250 -151
rect 278 -179 316 -151
rect 344 -179 382 -151
rect 410 -179 448 -151
rect 476 -179 514 -151
rect 542 -179 580 -151
rect 608 -179 646 -151
rect 674 -179 712 -151
rect 740 -179 745 -151
rect -745 -217 745 -179
rect -745 -245 -740 -217
rect -712 -245 -674 -217
rect -646 -245 -608 -217
rect -580 -245 -542 -217
rect -514 -245 -476 -217
rect -448 -245 -410 -217
rect -382 -245 -344 -217
rect -316 -245 -278 -217
rect -250 -245 -212 -217
rect -184 -245 -146 -217
rect -118 -245 -80 -217
rect -52 -245 -14 -217
rect 14 -245 52 -217
rect 80 -245 118 -217
rect 146 -245 184 -217
rect 212 -245 250 -217
rect 278 -245 316 -217
rect 344 -245 382 -217
rect 410 -245 448 -217
rect 476 -245 514 -217
rect 542 -245 580 -217
rect 608 -245 646 -217
rect 674 -245 712 -217
rect 740 -245 745 -217
rect -745 -283 745 -245
rect -745 -311 -740 -283
rect -712 -311 -674 -283
rect -646 -311 -608 -283
rect -580 -311 -542 -283
rect -514 -311 -476 -283
rect -448 -311 -410 -283
rect -382 -311 -344 -283
rect -316 -311 -278 -283
rect -250 -311 -212 -283
rect -184 -311 -146 -283
rect -118 -311 -80 -283
rect -52 -311 -14 -283
rect 14 -311 52 -283
rect 80 -311 118 -283
rect 146 -311 184 -283
rect 212 -311 250 -283
rect 278 -311 316 -283
rect 344 -311 382 -283
rect 410 -311 448 -283
rect 476 -311 514 -283
rect 542 -311 580 -283
rect 608 -311 646 -283
rect 674 -311 712 -283
rect 740 -311 745 -283
rect -745 -349 745 -311
rect -745 -377 -740 -349
rect -712 -377 -674 -349
rect -646 -377 -608 -349
rect -580 -377 -542 -349
rect -514 -377 -476 -349
rect -448 -377 -410 -349
rect -382 -377 -344 -349
rect -316 -377 -278 -349
rect -250 -377 -212 -349
rect -184 -377 -146 -349
rect -118 -377 -80 -349
rect -52 -377 -14 -349
rect 14 -377 52 -349
rect 80 -377 118 -349
rect 146 -377 184 -349
rect 212 -377 250 -349
rect 278 -377 316 -349
rect 344 -377 382 -349
rect 410 -377 448 -349
rect 476 -377 514 -349
rect 542 -377 580 -349
rect 608 -377 646 -349
rect 674 -377 712 -349
rect 740 -377 745 -349
rect -745 -415 745 -377
rect -745 -443 -740 -415
rect -712 -443 -674 -415
rect -646 -443 -608 -415
rect -580 -443 -542 -415
rect -514 -443 -476 -415
rect -448 -443 -410 -415
rect -382 -443 -344 -415
rect -316 -443 -278 -415
rect -250 -443 -212 -415
rect -184 -443 -146 -415
rect -118 -443 -80 -415
rect -52 -443 -14 -415
rect 14 -443 52 -415
rect 80 -443 118 -415
rect 146 -443 184 -415
rect 212 -443 250 -415
rect 278 -443 316 -415
rect 344 -443 382 -415
rect 410 -443 448 -415
rect 476 -443 514 -415
rect 542 -443 580 -415
rect 608 -443 646 -415
rect 674 -443 712 -415
rect 740 -443 745 -415
rect -745 -481 745 -443
rect -745 -509 -740 -481
rect -712 -509 -674 -481
rect -646 -509 -608 -481
rect -580 -509 -542 -481
rect -514 -509 -476 -481
rect -448 -509 -410 -481
rect -382 -509 -344 -481
rect -316 -509 -278 -481
rect -250 -509 -212 -481
rect -184 -509 -146 -481
rect -118 -509 -80 -481
rect -52 -509 -14 -481
rect 14 -509 52 -481
rect 80 -509 118 -481
rect 146 -509 184 -481
rect 212 -509 250 -481
rect 278 -509 316 -481
rect 344 -509 382 -481
rect 410 -509 448 -481
rect 476 -509 514 -481
rect 542 -509 580 -481
rect 608 -509 646 -481
rect 674 -509 712 -481
rect 740 -509 745 -481
rect -745 -547 745 -509
rect -745 -575 -740 -547
rect -712 -575 -674 -547
rect -646 -575 -608 -547
rect -580 -575 -542 -547
rect -514 -575 -476 -547
rect -448 -575 -410 -547
rect -382 -575 -344 -547
rect -316 -575 -278 -547
rect -250 -575 -212 -547
rect -184 -575 -146 -547
rect -118 -575 -80 -547
rect -52 -575 -14 -547
rect 14 -575 52 -547
rect 80 -575 118 -547
rect 146 -575 184 -547
rect 212 -575 250 -547
rect 278 -575 316 -547
rect 344 -575 382 -547
rect 410 -575 448 -547
rect 476 -575 514 -547
rect 542 -575 580 -547
rect 608 -575 646 -547
rect 674 -575 712 -547
rect 740 -575 745 -547
rect -745 -613 745 -575
rect -745 -641 -740 -613
rect -712 -641 -674 -613
rect -646 -641 -608 -613
rect -580 -641 -542 -613
rect -514 -641 -476 -613
rect -448 -641 -410 -613
rect -382 -641 -344 -613
rect -316 -641 -278 -613
rect -250 -641 -212 -613
rect -184 -641 -146 -613
rect -118 -641 -80 -613
rect -52 -641 -14 -613
rect 14 -641 52 -613
rect 80 -641 118 -613
rect 146 -641 184 -613
rect 212 -641 250 -613
rect 278 -641 316 -613
rect 344 -641 382 -613
rect 410 -641 448 -613
rect 476 -641 514 -613
rect 542 -641 580 -613
rect 608 -641 646 -613
rect 674 -641 712 -613
rect 740 -641 745 -613
rect -745 -679 745 -641
rect -745 -707 -740 -679
rect -712 -707 -674 -679
rect -646 -707 -608 -679
rect -580 -707 -542 -679
rect -514 -707 -476 -679
rect -448 -707 -410 -679
rect -382 -707 -344 -679
rect -316 -707 -278 -679
rect -250 -707 -212 -679
rect -184 -707 -146 -679
rect -118 -707 -80 -679
rect -52 -707 -14 -679
rect 14 -707 52 -679
rect 80 -707 118 -679
rect 146 -707 184 -679
rect 212 -707 250 -679
rect 278 -707 316 -679
rect 344 -707 382 -679
rect 410 -707 448 -679
rect 476 -707 514 -679
rect 542 -707 580 -679
rect 608 -707 646 -679
rect 674 -707 712 -679
rect 740 -707 745 -679
rect -745 -745 745 -707
rect -745 -773 -740 -745
rect -712 -773 -674 -745
rect -646 -773 -608 -745
rect -580 -773 -542 -745
rect -514 -773 -476 -745
rect -448 -773 -410 -745
rect -382 -773 -344 -745
rect -316 -773 -278 -745
rect -250 -773 -212 -745
rect -184 -773 -146 -745
rect -118 -773 -80 -745
rect -52 -773 -14 -745
rect 14 -773 52 -745
rect 80 -773 118 -745
rect 146 -773 184 -745
rect 212 -773 250 -745
rect 278 -773 316 -745
rect 344 -773 382 -745
rect 410 -773 448 -745
rect 476 -773 514 -745
rect 542 -773 580 -745
rect 608 -773 646 -745
rect 674 -773 712 -745
rect 740 -773 745 -745
rect -745 -811 745 -773
rect -745 -839 -740 -811
rect -712 -839 -674 -811
rect -646 -839 -608 -811
rect -580 -839 -542 -811
rect -514 -839 -476 -811
rect -448 -839 -410 -811
rect -382 -839 -344 -811
rect -316 -839 -278 -811
rect -250 -839 -212 -811
rect -184 -839 -146 -811
rect -118 -839 -80 -811
rect -52 -839 -14 -811
rect 14 -839 52 -811
rect 80 -839 118 -811
rect 146 -839 184 -811
rect 212 -839 250 -811
rect 278 -839 316 -811
rect 344 -839 382 -811
rect 410 -839 448 -811
rect 476 -839 514 -811
rect 542 -839 580 -811
rect 608 -839 646 -811
rect 674 -839 712 -811
rect 740 -839 745 -811
rect -745 -877 745 -839
rect -745 -905 -740 -877
rect -712 -905 -674 -877
rect -646 -905 -608 -877
rect -580 -905 -542 -877
rect -514 -905 -476 -877
rect -448 -905 -410 -877
rect -382 -905 -344 -877
rect -316 -905 -278 -877
rect -250 -905 -212 -877
rect -184 -905 -146 -877
rect -118 -905 -80 -877
rect -52 -905 -14 -877
rect 14 -905 52 -877
rect 80 -905 118 -877
rect 146 -905 184 -877
rect 212 -905 250 -877
rect 278 -905 316 -877
rect 344 -905 382 -877
rect 410 -905 448 -877
rect 476 -905 514 -877
rect 542 -905 580 -877
rect 608 -905 646 -877
rect 674 -905 712 -877
rect 740 -905 745 -877
rect -745 -943 745 -905
rect -745 -971 -740 -943
rect -712 -971 -674 -943
rect -646 -971 -608 -943
rect -580 -971 -542 -943
rect -514 -971 -476 -943
rect -448 -971 -410 -943
rect -382 -971 -344 -943
rect -316 -971 -278 -943
rect -250 -971 -212 -943
rect -184 -971 -146 -943
rect -118 -971 -80 -943
rect -52 -971 -14 -943
rect 14 -971 52 -943
rect 80 -971 118 -943
rect 146 -971 184 -943
rect 212 -971 250 -943
rect 278 -971 316 -943
rect 344 -971 382 -943
rect 410 -971 448 -943
rect 476 -971 514 -943
rect 542 -971 580 -943
rect 608 -971 646 -943
rect 674 -971 712 -943
rect 740 -971 745 -943
rect -745 -1009 745 -971
rect -745 -1037 -740 -1009
rect -712 -1037 -674 -1009
rect -646 -1037 -608 -1009
rect -580 -1037 -542 -1009
rect -514 -1037 -476 -1009
rect -448 -1037 -410 -1009
rect -382 -1037 -344 -1009
rect -316 -1037 -278 -1009
rect -250 -1037 -212 -1009
rect -184 -1037 -146 -1009
rect -118 -1037 -80 -1009
rect -52 -1037 -14 -1009
rect 14 -1037 52 -1009
rect 80 -1037 118 -1009
rect 146 -1037 184 -1009
rect 212 -1037 250 -1009
rect 278 -1037 316 -1009
rect 344 -1037 382 -1009
rect 410 -1037 448 -1009
rect 476 -1037 514 -1009
rect 542 -1037 580 -1009
rect 608 -1037 646 -1009
rect 674 -1037 712 -1009
rect 740 -1037 745 -1009
rect -745 -1075 745 -1037
rect -745 -1103 -740 -1075
rect -712 -1103 -674 -1075
rect -646 -1103 -608 -1075
rect -580 -1103 -542 -1075
rect -514 -1103 -476 -1075
rect -448 -1103 -410 -1075
rect -382 -1103 -344 -1075
rect -316 -1103 -278 -1075
rect -250 -1103 -212 -1075
rect -184 -1103 -146 -1075
rect -118 -1103 -80 -1075
rect -52 -1103 -14 -1075
rect 14 -1103 52 -1075
rect 80 -1103 118 -1075
rect 146 -1103 184 -1075
rect 212 -1103 250 -1075
rect 278 -1103 316 -1075
rect 344 -1103 382 -1075
rect 410 -1103 448 -1075
rect 476 -1103 514 -1075
rect 542 -1103 580 -1075
rect 608 -1103 646 -1075
rect 674 -1103 712 -1075
rect 740 -1103 745 -1075
rect -745 -1141 745 -1103
rect -745 -1169 -740 -1141
rect -712 -1169 -674 -1141
rect -646 -1169 -608 -1141
rect -580 -1169 -542 -1141
rect -514 -1169 -476 -1141
rect -448 -1169 -410 -1141
rect -382 -1169 -344 -1141
rect -316 -1169 -278 -1141
rect -250 -1169 -212 -1141
rect -184 -1169 -146 -1141
rect -118 -1169 -80 -1141
rect -52 -1169 -14 -1141
rect 14 -1169 52 -1141
rect 80 -1169 118 -1141
rect 146 -1169 184 -1141
rect 212 -1169 250 -1141
rect 278 -1169 316 -1141
rect 344 -1169 382 -1141
rect 410 -1169 448 -1141
rect 476 -1169 514 -1141
rect 542 -1169 580 -1141
rect 608 -1169 646 -1141
rect 674 -1169 712 -1141
rect 740 -1169 745 -1141
rect -745 -1207 745 -1169
rect -745 -1235 -740 -1207
rect -712 -1235 -674 -1207
rect -646 -1235 -608 -1207
rect -580 -1235 -542 -1207
rect -514 -1235 -476 -1207
rect -448 -1235 -410 -1207
rect -382 -1235 -344 -1207
rect -316 -1235 -278 -1207
rect -250 -1235 -212 -1207
rect -184 -1235 -146 -1207
rect -118 -1235 -80 -1207
rect -52 -1235 -14 -1207
rect 14 -1235 52 -1207
rect 80 -1235 118 -1207
rect 146 -1235 184 -1207
rect 212 -1235 250 -1207
rect 278 -1235 316 -1207
rect 344 -1235 382 -1207
rect 410 -1235 448 -1207
rect 476 -1235 514 -1207
rect 542 -1235 580 -1207
rect 608 -1235 646 -1207
rect 674 -1235 712 -1207
rect 740 -1235 745 -1207
rect -745 -1273 745 -1235
rect -745 -1301 -740 -1273
rect -712 -1301 -674 -1273
rect -646 -1301 -608 -1273
rect -580 -1301 -542 -1273
rect -514 -1301 -476 -1273
rect -448 -1301 -410 -1273
rect -382 -1301 -344 -1273
rect -316 -1301 -278 -1273
rect -250 -1301 -212 -1273
rect -184 -1301 -146 -1273
rect -118 -1301 -80 -1273
rect -52 -1301 -14 -1273
rect 14 -1301 52 -1273
rect 80 -1301 118 -1273
rect 146 -1301 184 -1273
rect 212 -1301 250 -1273
rect 278 -1301 316 -1273
rect 344 -1301 382 -1273
rect 410 -1301 448 -1273
rect 476 -1301 514 -1273
rect 542 -1301 580 -1273
rect 608 -1301 646 -1273
rect 674 -1301 712 -1273
rect 740 -1301 745 -1273
rect -745 -1339 745 -1301
rect -745 -1367 -740 -1339
rect -712 -1367 -674 -1339
rect -646 -1367 -608 -1339
rect -580 -1367 -542 -1339
rect -514 -1367 -476 -1339
rect -448 -1367 -410 -1339
rect -382 -1367 -344 -1339
rect -316 -1367 -278 -1339
rect -250 -1367 -212 -1339
rect -184 -1367 -146 -1339
rect -118 -1367 -80 -1339
rect -52 -1367 -14 -1339
rect 14 -1367 52 -1339
rect 80 -1367 118 -1339
rect 146 -1367 184 -1339
rect 212 -1367 250 -1339
rect 278 -1367 316 -1339
rect 344 -1367 382 -1339
rect 410 -1367 448 -1339
rect 476 -1367 514 -1339
rect 542 -1367 580 -1339
rect 608 -1367 646 -1339
rect 674 -1367 712 -1339
rect 740 -1367 745 -1339
rect -745 -1405 745 -1367
rect -745 -1433 -740 -1405
rect -712 -1433 -674 -1405
rect -646 -1433 -608 -1405
rect -580 -1433 -542 -1405
rect -514 -1433 -476 -1405
rect -448 -1433 -410 -1405
rect -382 -1433 -344 -1405
rect -316 -1433 -278 -1405
rect -250 -1433 -212 -1405
rect -184 -1433 -146 -1405
rect -118 -1433 -80 -1405
rect -52 -1433 -14 -1405
rect 14 -1433 52 -1405
rect 80 -1433 118 -1405
rect 146 -1433 184 -1405
rect 212 -1433 250 -1405
rect 278 -1433 316 -1405
rect 344 -1433 382 -1405
rect 410 -1433 448 -1405
rect 476 -1433 514 -1405
rect 542 -1433 580 -1405
rect 608 -1433 646 -1405
rect 674 -1433 712 -1405
rect 740 -1433 745 -1405
rect -745 -1471 745 -1433
rect -745 -1499 -740 -1471
rect -712 -1499 -674 -1471
rect -646 -1499 -608 -1471
rect -580 -1499 -542 -1471
rect -514 -1499 -476 -1471
rect -448 -1499 -410 -1471
rect -382 -1499 -344 -1471
rect -316 -1499 -278 -1471
rect -250 -1499 -212 -1471
rect -184 -1499 -146 -1471
rect -118 -1499 -80 -1471
rect -52 -1499 -14 -1471
rect 14 -1499 52 -1471
rect 80 -1499 118 -1471
rect 146 -1499 184 -1471
rect 212 -1499 250 -1471
rect 278 -1499 316 -1471
rect 344 -1499 382 -1471
rect 410 -1499 448 -1471
rect 476 -1499 514 -1471
rect 542 -1499 580 -1471
rect 608 -1499 646 -1471
rect 674 -1499 712 -1471
rect 740 -1499 745 -1471
rect -745 -1537 745 -1499
rect -745 -1565 -740 -1537
rect -712 -1565 -674 -1537
rect -646 -1565 -608 -1537
rect -580 -1565 -542 -1537
rect -514 -1565 -476 -1537
rect -448 -1565 -410 -1537
rect -382 -1565 -344 -1537
rect -316 -1565 -278 -1537
rect -250 -1565 -212 -1537
rect -184 -1565 -146 -1537
rect -118 -1565 -80 -1537
rect -52 -1565 -14 -1537
rect 14 -1565 52 -1537
rect 80 -1565 118 -1537
rect 146 -1565 184 -1537
rect 212 -1565 250 -1537
rect 278 -1565 316 -1537
rect 344 -1565 382 -1537
rect 410 -1565 448 -1537
rect 476 -1565 514 -1537
rect 542 -1565 580 -1537
rect 608 -1565 646 -1537
rect 674 -1565 712 -1537
rect 740 -1565 745 -1537
rect -745 -1603 745 -1565
rect -745 -1631 -740 -1603
rect -712 -1631 -674 -1603
rect -646 -1631 -608 -1603
rect -580 -1631 -542 -1603
rect -514 -1631 -476 -1603
rect -448 -1631 -410 -1603
rect -382 -1631 -344 -1603
rect -316 -1631 -278 -1603
rect -250 -1631 -212 -1603
rect -184 -1631 -146 -1603
rect -118 -1631 -80 -1603
rect -52 -1631 -14 -1603
rect 14 -1631 52 -1603
rect 80 -1631 118 -1603
rect 146 -1631 184 -1603
rect 212 -1631 250 -1603
rect 278 -1631 316 -1603
rect 344 -1631 382 -1603
rect 410 -1631 448 -1603
rect 476 -1631 514 -1603
rect 542 -1631 580 -1603
rect 608 -1631 646 -1603
rect 674 -1631 712 -1603
rect 740 -1631 745 -1603
rect -745 -1669 745 -1631
rect -745 -1697 -740 -1669
rect -712 -1697 -674 -1669
rect -646 -1697 -608 -1669
rect -580 -1697 -542 -1669
rect -514 -1697 -476 -1669
rect -448 -1697 -410 -1669
rect -382 -1697 -344 -1669
rect -316 -1697 -278 -1669
rect -250 -1697 -212 -1669
rect -184 -1697 -146 -1669
rect -118 -1697 -80 -1669
rect -52 -1697 -14 -1669
rect 14 -1697 52 -1669
rect 80 -1697 118 -1669
rect 146 -1697 184 -1669
rect 212 -1697 250 -1669
rect 278 -1697 316 -1669
rect 344 -1697 382 -1669
rect 410 -1697 448 -1669
rect 476 -1697 514 -1669
rect 542 -1697 580 -1669
rect 608 -1697 646 -1669
rect 674 -1697 712 -1669
rect 740 -1697 745 -1669
rect -745 -1735 745 -1697
rect -745 -1763 -740 -1735
rect -712 -1763 -674 -1735
rect -646 -1763 -608 -1735
rect -580 -1763 -542 -1735
rect -514 -1763 -476 -1735
rect -448 -1763 -410 -1735
rect -382 -1763 -344 -1735
rect -316 -1763 -278 -1735
rect -250 -1763 -212 -1735
rect -184 -1763 -146 -1735
rect -118 -1763 -80 -1735
rect -52 -1763 -14 -1735
rect 14 -1763 52 -1735
rect 80 -1763 118 -1735
rect 146 -1763 184 -1735
rect 212 -1763 250 -1735
rect 278 -1763 316 -1735
rect 344 -1763 382 -1735
rect 410 -1763 448 -1735
rect 476 -1763 514 -1735
rect 542 -1763 580 -1735
rect 608 -1763 646 -1735
rect 674 -1763 712 -1735
rect 740 -1763 745 -1735
rect -745 -1801 745 -1763
rect -745 -1829 -740 -1801
rect -712 -1829 -674 -1801
rect -646 -1829 -608 -1801
rect -580 -1829 -542 -1801
rect -514 -1829 -476 -1801
rect -448 -1829 -410 -1801
rect -382 -1829 -344 -1801
rect -316 -1829 -278 -1801
rect -250 -1829 -212 -1801
rect -184 -1829 -146 -1801
rect -118 -1829 -80 -1801
rect -52 -1829 -14 -1801
rect 14 -1829 52 -1801
rect 80 -1829 118 -1801
rect 146 -1829 184 -1801
rect 212 -1829 250 -1801
rect 278 -1829 316 -1801
rect 344 -1829 382 -1801
rect 410 -1829 448 -1801
rect 476 -1829 514 -1801
rect 542 -1829 580 -1801
rect 608 -1829 646 -1801
rect 674 -1829 712 -1801
rect 740 -1829 745 -1801
rect -745 -1867 745 -1829
rect -745 -1895 -740 -1867
rect -712 -1895 -674 -1867
rect -646 -1895 -608 -1867
rect -580 -1895 -542 -1867
rect -514 -1895 -476 -1867
rect -448 -1895 -410 -1867
rect -382 -1895 -344 -1867
rect -316 -1895 -278 -1867
rect -250 -1895 -212 -1867
rect -184 -1895 -146 -1867
rect -118 -1895 -80 -1867
rect -52 -1895 -14 -1867
rect 14 -1895 52 -1867
rect 80 -1895 118 -1867
rect 146 -1895 184 -1867
rect 212 -1895 250 -1867
rect 278 -1895 316 -1867
rect 344 -1895 382 -1867
rect 410 -1895 448 -1867
rect 476 -1895 514 -1867
rect 542 -1895 580 -1867
rect 608 -1895 646 -1867
rect 674 -1895 712 -1867
rect 740 -1895 745 -1867
rect -745 -1933 745 -1895
rect -745 -1961 -740 -1933
rect -712 -1961 -674 -1933
rect -646 -1961 -608 -1933
rect -580 -1961 -542 -1933
rect -514 -1961 -476 -1933
rect -448 -1961 -410 -1933
rect -382 -1961 -344 -1933
rect -316 -1961 -278 -1933
rect -250 -1961 -212 -1933
rect -184 -1961 -146 -1933
rect -118 -1961 -80 -1933
rect -52 -1961 -14 -1933
rect 14 -1961 52 -1933
rect 80 -1961 118 -1933
rect 146 -1961 184 -1933
rect 212 -1961 250 -1933
rect 278 -1961 316 -1933
rect 344 -1961 382 -1933
rect 410 -1961 448 -1933
rect 476 -1961 514 -1933
rect 542 -1961 580 -1933
rect 608 -1961 646 -1933
rect 674 -1961 712 -1933
rect 740 -1961 745 -1933
rect -745 -1999 745 -1961
rect -745 -2027 -740 -1999
rect -712 -2027 -674 -1999
rect -646 -2027 -608 -1999
rect -580 -2027 -542 -1999
rect -514 -2027 -476 -1999
rect -448 -2027 -410 -1999
rect -382 -2027 -344 -1999
rect -316 -2027 -278 -1999
rect -250 -2027 -212 -1999
rect -184 -2027 -146 -1999
rect -118 -2027 -80 -1999
rect -52 -2027 -14 -1999
rect 14 -2027 52 -1999
rect 80 -2027 118 -1999
rect 146 -2027 184 -1999
rect 212 -2027 250 -1999
rect 278 -2027 316 -1999
rect 344 -2027 382 -1999
rect 410 -2027 448 -1999
rect 476 -2027 514 -1999
rect 542 -2027 580 -1999
rect 608 -2027 646 -1999
rect 674 -2027 712 -1999
rect 740 -2027 745 -1999
rect -745 -2065 745 -2027
rect -745 -2093 -740 -2065
rect -712 -2093 -674 -2065
rect -646 -2093 -608 -2065
rect -580 -2093 -542 -2065
rect -514 -2093 -476 -2065
rect -448 -2093 -410 -2065
rect -382 -2093 -344 -2065
rect -316 -2093 -278 -2065
rect -250 -2093 -212 -2065
rect -184 -2093 -146 -2065
rect -118 -2093 -80 -2065
rect -52 -2093 -14 -2065
rect 14 -2093 52 -2065
rect 80 -2093 118 -2065
rect 146 -2093 184 -2065
rect 212 -2093 250 -2065
rect 278 -2093 316 -2065
rect 344 -2093 382 -2065
rect 410 -2093 448 -2065
rect 476 -2093 514 -2065
rect 542 -2093 580 -2065
rect 608 -2093 646 -2065
rect 674 -2093 712 -2065
rect 740 -2093 745 -2065
rect -745 -2131 745 -2093
rect -745 -2159 -740 -2131
rect -712 -2159 -674 -2131
rect -646 -2159 -608 -2131
rect -580 -2159 -542 -2131
rect -514 -2159 -476 -2131
rect -448 -2159 -410 -2131
rect -382 -2159 -344 -2131
rect -316 -2159 -278 -2131
rect -250 -2159 -212 -2131
rect -184 -2159 -146 -2131
rect -118 -2159 -80 -2131
rect -52 -2159 -14 -2131
rect 14 -2159 52 -2131
rect 80 -2159 118 -2131
rect 146 -2159 184 -2131
rect 212 -2159 250 -2131
rect 278 -2159 316 -2131
rect 344 -2159 382 -2131
rect 410 -2159 448 -2131
rect 476 -2159 514 -2131
rect 542 -2159 580 -2131
rect 608 -2159 646 -2131
rect 674 -2159 712 -2131
rect 740 -2159 745 -2131
rect -745 -2197 745 -2159
rect -745 -2225 -740 -2197
rect -712 -2225 -674 -2197
rect -646 -2225 -608 -2197
rect -580 -2225 -542 -2197
rect -514 -2225 -476 -2197
rect -448 -2225 -410 -2197
rect -382 -2225 -344 -2197
rect -316 -2225 -278 -2197
rect -250 -2225 -212 -2197
rect -184 -2225 -146 -2197
rect -118 -2225 -80 -2197
rect -52 -2225 -14 -2197
rect 14 -2225 52 -2197
rect 80 -2225 118 -2197
rect 146 -2225 184 -2197
rect 212 -2225 250 -2197
rect 278 -2225 316 -2197
rect 344 -2225 382 -2197
rect 410 -2225 448 -2197
rect 476 -2225 514 -2197
rect 542 -2225 580 -2197
rect 608 -2225 646 -2197
rect 674 -2225 712 -2197
rect 740 -2225 745 -2197
rect -745 -2263 745 -2225
rect -745 -2291 -740 -2263
rect -712 -2291 -674 -2263
rect -646 -2291 -608 -2263
rect -580 -2291 -542 -2263
rect -514 -2291 -476 -2263
rect -448 -2291 -410 -2263
rect -382 -2291 -344 -2263
rect -316 -2291 -278 -2263
rect -250 -2291 -212 -2263
rect -184 -2291 -146 -2263
rect -118 -2291 -80 -2263
rect -52 -2291 -14 -2263
rect 14 -2291 52 -2263
rect 80 -2291 118 -2263
rect 146 -2291 184 -2263
rect 212 -2291 250 -2263
rect 278 -2291 316 -2263
rect 344 -2291 382 -2263
rect 410 -2291 448 -2263
rect 476 -2291 514 -2263
rect 542 -2291 580 -2263
rect 608 -2291 646 -2263
rect 674 -2291 712 -2263
rect 740 -2291 745 -2263
rect -745 -2329 745 -2291
rect -745 -2357 -740 -2329
rect -712 -2357 -674 -2329
rect -646 -2357 -608 -2329
rect -580 -2357 -542 -2329
rect -514 -2357 -476 -2329
rect -448 -2357 -410 -2329
rect -382 -2357 -344 -2329
rect -316 -2357 -278 -2329
rect -250 -2357 -212 -2329
rect -184 -2357 -146 -2329
rect -118 -2357 -80 -2329
rect -52 -2357 -14 -2329
rect 14 -2357 52 -2329
rect 80 -2357 118 -2329
rect 146 -2357 184 -2329
rect 212 -2357 250 -2329
rect 278 -2357 316 -2329
rect 344 -2357 382 -2329
rect 410 -2357 448 -2329
rect 476 -2357 514 -2329
rect 542 -2357 580 -2329
rect 608 -2357 646 -2329
rect 674 -2357 712 -2329
rect 740 -2357 745 -2329
rect -745 -2395 745 -2357
rect -745 -2423 -740 -2395
rect -712 -2423 -674 -2395
rect -646 -2423 -608 -2395
rect -580 -2423 -542 -2395
rect -514 -2423 -476 -2395
rect -448 -2423 -410 -2395
rect -382 -2423 -344 -2395
rect -316 -2423 -278 -2395
rect -250 -2423 -212 -2395
rect -184 -2423 -146 -2395
rect -118 -2423 -80 -2395
rect -52 -2423 -14 -2395
rect 14 -2423 52 -2395
rect 80 -2423 118 -2395
rect 146 -2423 184 -2395
rect 212 -2423 250 -2395
rect 278 -2423 316 -2395
rect 344 -2423 382 -2395
rect 410 -2423 448 -2395
rect 476 -2423 514 -2395
rect 542 -2423 580 -2395
rect 608 -2423 646 -2395
rect 674 -2423 712 -2395
rect 740 -2423 745 -2395
rect -745 -2461 745 -2423
rect -745 -2489 -740 -2461
rect -712 -2489 -674 -2461
rect -646 -2489 -608 -2461
rect -580 -2489 -542 -2461
rect -514 -2489 -476 -2461
rect -448 -2489 -410 -2461
rect -382 -2489 -344 -2461
rect -316 -2489 -278 -2461
rect -250 -2489 -212 -2461
rect -184 -2489 -146 -2461
rect -118 -2489 -80 -2461
rect -52 -2489 -14 -2461
rect 14 -2489 52 -2461
rect 80 -2489 118 -2461
rect 146 -2489 184 -2461
rect 212 -2489 250 -2461
rect 278 -2489 316 -2461
rect 344 -2489 382 -2461
rect 410 -2489 448 -2461
rect 476 -2489 514 -2461
rect 542 -2489 580 -2461
rect 608 -2489 646 -2461
rect 674 -2489 712 -2461
rect 740 -2489 745 -2461
rect -745 -2527 745 -2489
rect -745 -2555 -740 -2527
rect -712 -2555 -674 -2527
rect -646 -2555 -608 -2527
rect -580 -2555 -542 -2527
rect -514 -2555 -476 -2527
rect -448 -2555 -410 -2527
rect -382 -2555 -344 -2527
rect -316 -2555 -278 -2527
rect -250 -2555 -212 -2527
rect -184 -2555 -146 -2527
rect -118 -2555 -80 -2527
rect -52 -2555 -14 -2527
rect 14 -2555 52 -2527
rect 80 -2555 118 -2527
rect 146 -2555 184 -2527
rect 212 -2555 250 -2527
rect 278 -2555 316 -2527
rect 344 -2555 382 -2527
rect 410 -2555 448 -2527
rect 476 -2555 514 -2527
rect 542 -2555 580 -2527
rect 608 -2555 646 -2527
rect 674 -2555 712 -2527
rect 740 -2555 745 -2527
rect -745 -2593 745 -2555
rect -745 -2621 -740 -2593
rect -712 -2621 -674 -2593
rect -646 -2621 -608 -2593
rect -580 -2621 -542 -2593
rect -514 -2621 -476 -2593
rect -448 -2621 -410 -2593
rect -382 -2621 -344 -2593
rect -316 -2621 -278 -2593
rect -250 -2621 -212 -2593
rect -184 -2621 -146 -2593
rect -118 -2621 -80 -2593
rect -52 -2621 -14 -2593
rect 14 -2621 52 -2593
rect 80 -2621 118 -2593
rect 146 -2621 184 -2593
rect 212 -2621 250 -2593
rect 278 -2621 316 -2593
rect 344 -2621 382 -2593
rect 410 -2621 448 -2593
rect 476 -2621 514 -2593
rect 542 -2621 580 -2593
rect 608 -2621 646 -2593
rect 674 -2621 712 -2593
rect 740 -2621 745 -2593
rect -745 -2659 745 -2621
rect -745 -2687 -740 -2659
rect -712 -2687 -674 -2659
rect -646 -2687 -608 -2659
rect -580 -2687 -542 -2659
rect -514 -2687 -476 -2659
rect -448 -2687 -410 -2659
rect -382 -2687 -344 -2659
rect -316 -2687 -278 -2659
rect -250 -2687 -212 -2659
rect -184 -2687 -146 -2659
rect -118 -2687 -80 -2659
rect -52 -2687 -14 -2659
rect 14 -2687 52 -2659
rect 80 -2687 118 -2659
rect 146 -2687 184 -2659
rect 212 -2687 250 -2659
rect 278 -2687 316 -2659
rect 344 -2687 382 -2659
rect 410 -2687 448 -2659
rect 476 -2687 514 -2659
rect 542 -2687 580 -2659
rect 608 -2687 646 -2659
rect 674 -2687 712 -2659
rect 740 -2687 745 -2659
rect -745 -2725 745 -2687
rect -745 -2753 -740 -2725
rect -712 -2753 -674 -2725
rect -646 -2753 -608 -2725
rect -580 -2753 -542 -2725
rect -514 -2753 -476 -2725
rect -448 -2753 -410 -2725
rect -382 -2753 -344 -2725
rect -316 -2753 -278 -2725
rect -250 -2753 -212 -2725
rect -184 -2753 -146 -2725
rect -118 -2753 -80 -2725
rect -52 -2753 -14 -2725
rect 14 -2753 52 -2725
rect 80 -2753 118 -2725
rect 146 -2753 184 -2725
rect 212 -2753 250 -2725
rect 278 -2753 316 -2725
rect 344 -2753 382 -2725
rect 410 -2753 448 -2725
rect 476 -2753 514 -2725
rect 542 -2753 580 -2725
rect 608 -2753 646 -2725
rect 674 -2753 712 -2725
rect 740 -2753 745 -2725
rect -745 -2791 745 -2753
rect -745 -2819 -740 -2791
rect -712 -2819 -674 -2791
rect -646 -2819 -608 -2791
rect -580 -2819 -542 -2791
rect -514 -2819 -476 -2791
rect -448 -2819 -410 -2791
rect -382 -2819 -344 -2791
rect -316 -2819 -278 -2791
rect -250 -2819 -212 -2791
rect -184 -2819 -146 -2791
rect -118 -2819 -80 -2791
rect -52 -2819 -14 -2791
rect 14 -2819 52 -2791
rect 80 -2819 118 -2791
rect 146 -2819 184 -2791
rect 212 -2819 250 -2791
rect 278 -2819 316 -2791
rect 344 -2819 382 -2791
rect 410 -2819 448 -2791
rect 476 -2819 514 -2791
rect 542 -2819 580 -2791
rect 608 -2819 646 -2791
rect 674 -2819 712 -2791
rect 740 -2819 745 -2791
rect -745 -2857 745 -2819
rect -745 -2885 -740 -2857
rect -712 -2885 -674 -2857
rect -646 -2885 -608 -2857
rect -580 -2885 -542 -2857
rect -514 -2885 -476 -2857
rect -448 -2885 -410 -2857
rect -382 -2885 -344 -2857
rect -316 -2885 -278 -2857
rect -250 -2885 -212 -2857
rect -184 -2885 -146 -2857
rect -118 -2885 -80 -2857
rect -52 -2885 -14 -2857
rect 14 -2885 52 -2857
rect 80 -2885 118 -2857
rect 146 -2885 184 -2857
rect 212 -2885 250 -2857
rect 278 -2885 316 -2857
rect 344 -2885 382 -2857
rect 410 -2885 448 -2857
rect 476 -2885 514 -2857
rect 542 -2885 580 -2857
rect 608 -2885 646 -2857
rect 674 -2885 712 -2857
rect 740 -2885 745 -2857
rect -745 -2923 745 -2885
rect -745 -2951 -740 -2923
rect -712 -2951 -674 -2923
rect -646 -2951 -608 -2923
rect -580 -2951 -542 -2923
rect -514 -2951 -476 -2923
rect -448 -2951 -410 -2923
rect -382 -2951 -344 -2923
rect -316 -2951 -278 -2923
rect -250 -2951 -212 -2923
rect -184 -2951 -146 -2923
rect -118 -2951 -80 -2923
rect -52 -2951 -14 -2923
rect 14 -2951 52 -2923
rect 80 -2951 118 -2923
rect 146 -2951 184 -2923
rect 212 -2951 250 -2923
rect 278 -2951 316 -2923
rect 344 -2951 382 -2923
rect 410 -2951 448 -2923
rect 476 -2951 514 -2923
rect 542 -2951 580 -2923
rect 608 -2951 646 -2923
rect 674 -2951 712 -2923
rect 740 -2951 745 -2923
rect -745 -2989 745 -2951
rect -745 -3017 -740 -2989
rect -712 -3017 -674 -2989
rect -646 -3017 -608 -2989
rect -580 -3017 -542 -2989
rect -514 -3017 -476 -2989
rect -448 -3017 -410 -2989
rect -382 -3017 -344 -2989
rect -316 -3017 -278 -2989
rect -250 -3017 -212 -2989
rect -184 -3017 -146 -2989
rect -118 -3017 -80 -2989
rect -52 -3017 -14 -2989
rect 14 -3017 52 -2989
rect 80 -3017 118 -2989
rect 146 -3017 184 -2989
rect 212 -3017 250 -2989
rect 278 -3017 316 -2989
rect 344 -3017 382 -2989
rect 410 -3017 448 -2989
rect 476 -3017 514 -2989
rect 542 -3017 580 -2989
rect 608 -3017 646 -2989
rect 674 -3017 712 -2989
rect 740 -3017 745 -2989
rect -745 -3055 745 -3017
rect -745 -3083 -740 -3055
rect -712 -3083 -674 -3055
rect -646 -3083 -608 -3055
rect -580 -3083 -542 -3055
rect -514 -3083 -476 -3055
rect -448 -3083 -410 -3055
rect -382 -3083 -344 -3055
rect -316 -3083 -278 -3055
rect -250 -3083 -212 -3055
rect -184 -3083 -146 -3055
rect -118 -3083 -80 -3055
rect -52 -3083 -14 -3055
rect 14 -3083 52 -3055
rect 80 -3083 118 -3055
rect 146 -3083 184 -3055
rect 212 -3083 250 -3055
rect 278 -3083 316 -3055
rect 344 -3083 382 -3055
rect 410 -3083 448 -3055
rect 476 -3083 514 -3055
rect 542 -3083 580 -3055
rect 608 -3083 646 -3055
rect 674 -3083 712 -3055
rect 740 -3083 745 -3055
rect -745 -3121 745 -3083
rect -745 -3149 -740 -3121
rect -712 -3149 -674 -3121
rect -646 -3149 -608 -3121
rect -580 -3149 -542 -3121
rect -514 -3149 -476 -3121
rect -448 -3149 -410 -3121
rect -382 -3149 -344 -3121
rect -316 -3149 -278 -3121
rect -250 -3149 -212 -3121
rect -184 -3149 -146 -3121
rect -118 -3149 -80 -3121
rect -52 -3149 -14 -3121
rect 14 -3149 52 -3121
rect 80 -3149 118 -3121
rect 146 -3149 184 -3121
rect 212 -3149 250 -3121
rect 278 -3149 316 -3121
rect 344 -3149 382 -3121
rect 410 -3149 448 -3121
rect 476 -3149 514 -3121
rect 542 -3149 580 -3121
rect 608 -3149 646 -3121
rect 674 -3149 712 -3121
rect 740 -3149 745 -3121
rect -745 -3187 745 -3149
rect -745 -3215 -740 -3187
rect -712 -3215 -674 -3187
rect -646 -3215 -608 -3187
rect -580 -3215 -542 -3187
rect -514 -3215 -476 -3187
rect -448 -3215 -410 -3187
rect -382 -3215 -344 -3187
rect -316 -3215 -278 -3187
rect -250 -3215 -212 -3187
rect -184 -3215 -146 -3187
rect -118 -3215 -80 -3187
rect -52 -3215 -14 -3187
rect 14 -3215 52 -3187
rect 80 -3215 118 -3187
rect 146 -3215 184 -3187
rect 212 -3215 250 -3187
rect 278 -3215 316 -3187
rect 344 -3215 382 -3187
rect 410 -3215 448 -3187
rect 476 -3215 514 -3187
rect 542 -3215 580 -3187
rect 608 -3215 646 -3187
rect 674 -3215 712 -3187
rect 740 -3215 745 -3187
rect -745 -3253 745 -3215
rect -745 -3281 -740 -3253
rect -712 -3281 -674 -3253
rect -646 -3281 -608 -3253
rect -580 -3281 -542 -3253
rect -514 -3281 -476 -3253
rect -448 -3281 -410 -3253
rect -382 -3281 -344 -3253
rect -316 -3281 -278 -3253
rect -250 -3281 -212 -3253
rect -184 -3281 -146 -3253
rect -118 -3281 -80 -3253
rect -52 -3281 -14 -3253
rect 14 -3281 52 -3253
rect 80 -3281 118 -3253
rect 146 -3281 184 -3253
rect 212 -3281 250 -3253
rect 278 -3281 316 -3253
rect 344 -3281 382 -3253
rect 410 -3281 448 -3253
rect 476 -3281 514 -3253
rect 542 -3281 580 -3253
rect 608 -3281 646 -3253
rect 674 -3281 712 -3253
rect 740 -3281 745 -3253
rect -745 -3319 745 -3281
rect -745 -3347 -740 -3319
rect -712 -3347 -674 -3319
rect -646 -3347 -608 -3319
rect -580 -3347 -542 -3319
rect -514 -3347 -476 -3319
rect -448 -3347 -410 -3319
rect -382 -3347 -344 -3319
rect -316 -3347 -278 -3319
rect -250 -3347 -212 -3319
rect -184 -3347 -146 -3319
rect -118 -3347 -80 -3319
rect -52 -3347 -14 -3319
rect 14 -3347 52 -3319
rect 80 -3347 118 -3319
rect 146 -3347 184 -3319
rect 212 -3347 250 -3319
rect 278 -3347 316 -3319
rect 344 -3347 382 -3319
rect 410 -3347 448 -3319
rect 476 -3347 514 -3319
rect 542 -3347 580 -3319
rect 608 -3347 646 -3319
rect 674 -3347 712 -3319
rect 740 -3347 745 -3319
rect -745 -3385 745 -3347
rect -745 -3413 -740 -3385
rect -712 -3413 -674 -3385
rect -646 -3413 -608 -3385
rect -580 -3413 -542 -3385
rect -514 -3413 -476 -3385
rect -448 -3413 -410 -3385
rect -382 -3413 -344 -3385
rect -316 -3413 -278 -3385
rect -250 -3413 -212 -3385
rect -184 -3413 -146 -3385
rect -118 -3413 -80 -3385
rect -52 -3413 -14 -3385
rect 14 -3413 52 -3385
rect 80 -3413 118 -3385
rect 146 -3413 184 -3385
rect 212 -3413 250 -3385
rect 278 -3413 316 -3385
rect 344 -3413 382 -3385
rect 410 -3413 448 -3385
rect 476 -3413 514 -3385
rect 542 -3413 580 -3385
rect 608 -3413 646 -3385
rect 674 -3413 712 -3385
rect 740 -3413 745 -3385
rect -745 -3451 745 -3413
rect -745 -3479 -740 -3451
rect -712 -3479 -674 -3451
rect -646 -3479 -608 -3451
rect -580 -3479 -542 -3451
rect -514 -3479 -476 -3451
rect -448 -3479 -410 -3451
rect -382 -3479 -344 -3451
rect -316 -3479 -278 -3451
rect -250 -3479 -212 -3451
rect -184 -3479 -146 -3451
rect -118 -3479 -80 -3451
rect -52 -3479 -14 -3451
rect 14 -3479 52 -3451
rect 80 -3479 118 -3451
rect 146 -3479 184 -3451
rect 212 -3479 250 -3451
rect 278 -3479 316 -3451
rect 344 -3479 382 -3451
rect 410 -3479 448 -3451
rect 476 -3479 514 -3451
rect 542 -3479 580 -3451
rect 608 -3479 646 -3451
rect 674 -3479 712 -3451
rect 740 -3479 745 -3451
rect -745 -3517 745 -3479
rect -745 -3545 -740 -3517
rect -712 -3545 -674 -3517
rect -646 -3545 -608 -3517
rect -580 -3545 -542 -3517
rect -514 -3545 -476 -3517
rect -448 -3545 -410 -3517
rect -382 -3545 -344 -3517
rect -316 -3545 -278 -3517
rect -250 -3545 -212 -3517
rect -184 -3545 -146 -3517
rect -118 -3545 -80 -3517
rect -52 -3545 -14 -3517
rect 14 -3545 52 -3517
rect 80 -3545 118 -3517
rect 146 -3545 184 -3517
rect 212 -3545 250 -3517
rect 278 -3545 316 -3517
rect 344 -3545 382 -3517
rect 410 -3545 448 -3517
rect 476 -3545 514 -3517
rect 542 -3545 580 -3517
rect 608 -3545 646 -3517
rect 674 -3545 712 -3517
rect 740 -3545 745 -3517
rect -745 -3583 745 -3545
rect -745 -3611 -740 -3583
rect -712 -3611 -674 -3583
rect -646 -3611 -608 -3583
rect -580 -3611 -542 -3583
rect -514 -3611 -476 -3583
rect -448 -3611 -410 -3583
rect -382 -3611 -344 -3583
rect -316 -3611 -278 -3583
rect -250 -3611 -212 -3583
rect -184 -3611 -146 -3583
rect -118 -3611 -80 -3583
rect -52 -3611 -14 -3583
rect 14 -3611 52 -3583
rect 80 -3611 118 -3583
rect 146 -3611 184 -3583
rect 212 -3611 250 -3583
rect 278 -3611 316 -3583
rect 344 -3611 382 -3583
rect 410 -3611 448 -3583
rect 476 -3611 514 -3583
rect 542 -3611 580 -3583
rect 608 -3611 646 -3583
rect 674 -3611 712 -3583
rect 740 -3611 745 -3583
rect -745 -3649 745 -3611
rect -745 -3677 -740 -3649
rect -712 -3677 -674 -3649
rect -646 -3677 -608 -3649
rect -580 -3677 -542 -3649
rect -514 -3677 -476 -3649
rect -448 -3677 -410 -3649
rect -382 -3677 -344 -3649
rect -316 -3677 -278 -3649
rect -250 -3677 -212 -3649
rect -184 -3677 -146 -3649
rect -118 -3677 -80 -3649
rect -52 -3677 -14 -3649
rect 14 -3677 52 -3649
rect 80 -3677 118 -3649
rect 146 -3677 184 -3649
rect 212 -3677 250 -3649
rect 278 -3677 316 -3649
rect 344 -3677 382 -3649
rect 410 -3677 448 -3649
rect 476 -3677 514 -3649
rect 542 -3677 580 -3649
rect 608 -3677 646 -3649
rect 674 -3677 712 -3649
rect 740 -3677 745 -3649
rect -745 -3715 745 -3677
rect -745 -3743 -740 -3715
rect -712 -3743 -674 -3715
rect -646 -3743 -608 -3715
rect -580 -3743 -542 -3715
rect -514 -3743 -476 -3715
rect -448 -3743 -410 -3715
rect -382 -3743 -344 -3715
rect -316 -3743 -278 -3715
rect -250 -3743 -212 -3715
rect -184 -3743 -146 -3715
rect -118 -3743 -80 -3715
rect -52 -3743 -14 -3715
rect 14 -3743 52 -3715
rect 80 -3743 118 -3715
rect 146 -3743 184 -3715
rect 212 -3743 250 -3715
rect 278 -3743 316 -3715
rect 344 -3743 382 -3715
rect 410 -3743 448 -3715
rect 476 -3743 514 -3715
rect 542 -3743 580 -3715
rect 608 -3743 646 -3715
rect 674 -3743 712 -3715
rect 740 -3743 745 -3715
rect -745 -3781 745 -3743
rect -745 -3809 -740 -3781
rect -712 -3809 -674 -3781
rect -646 -3809 -608 -3781
rect -580 -3809 -542 -3781
rect -514 -3809 -476 -3781
rect -448 -3809 -410 -3781
rect -382 -3809 -344 -3781
rect -316 -3809 -278 -3781
rect -250 -3809 -212 -3781
rect -184 -3809 -146 -3781
rect -118 -3809 -80 -3781
rect -52 -3809 -14 -3781
rect 14 -3809 52 -3781
rect 80 -3809 118 -3781
rect 146 -3809 184 -3781
rect 212 -3809 250 -3781
rect 278 -3809 316 -3781
rect 344 -3809 382 -3781
rect 410 -3809 448 -3781
rect 476 -3809 514 -3781
rect 542 -3809 580 -3781
rect 608 -3809 646 -3781
rect 674 -3809 712 -3781
rect 740 -3809 745 -3781
rect -745 -3847 745 -3809
rect -745 -3875 -740 -3847
rect -712 -3875 -674 -3847
rect -646 -3875 -608 -3847
rect -580 -3875 -542 -3847
rect -514 -3875 -476 -3847
rect -448 -3875 -410 -3847
rect -382 -3875 -344 -3847
rect -316 -3875 -278 -3847
rect -250 -3875 -212 -3847
rect -184 -3875 -146 -3847
rect -118 -3875 -80 -3847
rect -52 -3875 -14 -3847
rect 14 -3875 52 -3847
rect 80 -3875 118 -3847
rect 146 -3875 184 -3847
rect 212 -3875 250 -3847
rect 278 -3875 316 -3847
rect 344 -3875 382 -3847
rect 410 -3875 448 -3847
rect 476 -3875 514 -3847
rect 542 -3875 580 -3847
rect 608 -3875 646 -3847
rect 674 -3875 712 -3847
rect 740 -3875 745 -3847
rect -745 -3880 745 -3875
<< via3 >>
rect -740 3847 -712 3875
rect -674 3847 -646 3875
rect -608 3847 -580 3875
rect -542 3847 -514 3875
rect -476 3847 -448 3875
rect -410 3847 -382 3875
rect -344 3847 -316 3875
rect -278 3847 -250 3875
rect -212 3847 -184 3875
rect -146 3847 -118 3875
rect -80 3847 -52 3875
rect -14 3847 14 3875
rect 52 3847 80 3875
rect 118 3847 146 3875
rect 184 3847 212 3875
rect 250 3847 278 3875
rect 316 3847 344 3875
rect 382 3847 410 3875
rect 448 3847 476 3875
rect 514 3847 542 3875
rect 580 3847 608 3875
rect 646 3847 674 3875
rect 712 3847 740 3875
rect -740 3781 -712 3809
rect -674 3781 -646 3809
rect -608 3781 -580 3809
rect -542 3781 -514 3809
rect -476 3781 -448 3809
rect -410 3781 -382 3809
rect -344 3781 -316 3809
rect -278 3781 -250 3809
rect -212 3781 -184 3809
rect -146 3781 -118 3809
rect -80 3781 -52 3809
rect -14 3781 14 3809
rect 52 3781 80 3809
rect 118 3781 146 3809
rect 184 3781 212 3809
rect 250 3781 278 3809
rect 316 3781 344 3809
rect 382 3781 410 3809
rect 448 3781 476 3809
rect 514 3781 542 3809
rect 580 3781 608 3809
rect 646 3781 674 3809
rect 712 3781 740 3809
rect -740 3715 -712 3743
rect -674 3715 -646 3743
rect -608 3715 -580 3743
rect -542 3715 -514 3743
rect -476 3715 -448 3743
rect -410 3715 -382 3743
rect -344 3715 -316 3743
rect -278 3715 -250 3743
rect -212 3715 -184 3743
rect -146 3715 -118 3743
rect -80 3715 -52 3743
rect -14 3715 14 3743
rect 52 3715 80 3743
rect 118 3715 146 3743
rect 184 3715 212 3743
rect 250 3715 278 3743
rect 316 3715 344 3743
rect 382 3715 410 3743
rect 448 3715 476 3743
rect 514 3715 542 3743
rect 580 3715 608 3743
rect 646 3715 674 3743
rect 712 3715 740 3743
rect -740 3649 -712 3677
rect -674 3649 -646 3677
rect -608 3649 -580 3677
rect -542 3649 -514 3677
rect -476 3649 -448 3677
rect -410 3649 -382 3677
rect -344 3649 -316 3677
rect -278 3649 -250 3677
rect -212 3649 -184 3677
rect -146 3649 -118 3677
rect -80 3649 -52 3677
rect -14 3649 14 3677
rect 52 3649 80 3677
rect 118 3649 146 3677
rect 184 3649 212 3677
rect 250 3649 278 3677
rect 316 3649 344 3677
rect 382 3649 410 3677
rect 448 3649 476 3677
rect 514 3649 542 3677
rect 580 3649 608 3677
rect 646 3649 674 3677
rect 712 3649 740 3677
rect -740 3583 -712 3611
rect -674 3583 -646 3611
rect -608 3583 -580 3611
rect -542 3583 -514 3611
rect -476 3583 -448 3611
rect -410 3583 -382 3611
rect -344 3583 -316 3611
rect -278 3583 -250 3611
rect -212 3583 -184 3611
rect -146 3583 -118 3611
rect -80 3583 -52 3611
rect -14 3583 14 3611
rect 52 3583 80 3611
rect 118 3583 146 3611
rect 184 3583 212 3611
rect 250 3583 278 3611
rect 316 3583 344 3611
rect 382 3583 410 3611
rect 448 3583 476 3611
rect 514 3583 542 3611
rect 580 3583 608 3611
rect 646 3583 674 3611
rect 712 3583 740 3611
rect -740 3517 -712 3545
rect -674 3517 -646 3545
rect -608 3517 -580 3545
rect -542 3517 -514 3545
rect -476 3517 -448 3545
rect -410 3517 -382 3545
rect -344 3517 -316 3545
rect -278 3517 -250 3545
rect -212 3517 -184 3545
rect -146 3517 -118 3545
rect -80 3517 -52 3545
rect -14 3517 14 3545
rect 52 3517 80 3545
rect 118 3517 146 3545
rect 184 3517 212 3545
rect 250 3517 278 3545
rect 316 3517 344 3545
rect 382 3517 410 3545
rect 448 3517 476 3545
rect 514 3517 542 3545
rect 580 3517 608 3545
rect 646 3517 674 3545
rect 712 3517 740 3545
rect -740 3451 -712 3479
rect -674 3451 -646 3479
rect -608 3451 -580 3479
rect -542 3451 -514 3479
rect -476 3451 -448 3479
rect -410 3451 -382 3479
rect -344 3451 -316 3479
rect -278 3451 -250 3479
rect -212 3451 -184 3479
rect -146 3451 -118 3479
rect -80 3451 -52 3479
rect -14 3451 14 3479
rect 52 3451 80 3479
rect 118 3451 146 3479
rect 184 3451 212 3479
rect 250 3451 278 3479
rect 316 3451 344 3479
rect 382 3451 410 3479
rect 448 3451 476 3479
rect 514 3451 542 3479
rect 580 3451 608 3479
rect 646 3451 674 3479
rect 712 3451 740 3479
rect -740 3385 -712 3413
rect -674 3385 -646 3413
rect -608 3385 -580 3413
rect -542 3385 -514 3413
rect -476 3385 -448 3413
rect -410 3385 -382 3413
rect -344 3385 -316 3413
rect -278 3385 -250 3413
rect -212 3385 -184 3413
rect -146 3385 -118 3413
rect -80 3385 -52 3413
rect -14 3385 14 3413
rect 52 3385 80 3413
rect 118 3385 146 3413
rect 184 3385 212 3413
rect 250 3385 278 3413
rect 316 3385 344 3413
rect 382 3385 410 3413
rect 448 3385 476 3413
rect 514 3385 542 3413
rect 580 3385 608 3413
rect 646 3385 674 3413
rect 712 3385 740 3413
rect -740 3319 -712 3347
rect -674 3319 -646 3347
rect -608 3319 -580 3347
rect -542 3319 -514 3347
rect -476 3319 -448 3347
rect -410 3319 -382 3347
rect -344 3319 -316 3347
rect -278 3319 -250 3347
rect -212 3319 -184 3347
rect -146 3319 -118 3347
rect -80 3319 -52 3347
rect -14 3319 14 3347
rect 52 3319 80 3347
rect 118 3319 146 3347
rect 184 3319 212 3347
rect 250 3319 278 3347
rect 316 3319 344 3347
rect 382 3319 410 3347
rect 448 3319 476 3347
rect 514 3319 542 3347
rect 580 3319 608 3347
rect 646 3319 674 3347
rect 712 3319 740 3347
rect -740 3253 -712 3281
rect -674 3253 -646 3281
rect -608 3253 -580 3281
rect -542 3253 -514 3281
rect -476 3253 -448 3281
rect -410 3253 -382 3281
rect -344 3253 -316 3281
rect -278 3253 -250 3281
rect -212 3253 -184 3281
rect -146 3253 -118 3281
rect -80 3253 -52 3281
rect -14 3253 14 3281
rect 52 3253 80 3281
rect 118 3253 146 3281
rect 184 3253 212 3281
rect 250 3253 278 3281
rect 316 3253 344 3281
rect 382 3253 410 3281
rect 448 3253 476 3281
rect 514 3253 542 3281
rect 580 3253 608 3281
rect 646 3253 674 3281
rect 712 3253 740 3281
rect -740 3187 -712 3215
rect -674 3187 -646 3215
rect -608 3187 -580 3215
rect -542 3187 -514 3215
rect -476 3187 -448 3215
rect -410 3187 -382 3215
rect -344 3187 -316 3215
rect -278 3187 -250 3215
rect -212 3187 -184 3215
rect -146 3187 -118 3215
rect -80 3187 -52 3215
rect -14 3187 14 3215
rect 52 3187 80 3215
rect 118 3187 146 3215
rect 184 3187 212 3215
rect 250 3187 278 3215
rect 316 3187 344 3215
rect 382 3187 410 3215
rect 448 3187 476 3215
rect 514 3187 542 3215
rect 580 3187 608 3215
rect 646 3187 674 3215
rect 712 3187 740 3215
rect -740 3121 -712 3149
rect -674 3121 -646 3149
rect -608 3121 -580 3149
rect -542 3121 -514 3149
rect -476 3121 -448 3149
rect -410 3121 -382 3149
rect -344 3121 -316 3149
rect -278 3121 -250 3149
rect -212 3121 -184 3149
rect -146 3121 -118 3149
rect -80 3121 -52 3149
rect -14 3121 14 3149
rect 52 3121 80 3149
rect 118 3121 146 3149
rect 184 3121 212 3149
rect 250 3121 278 3149
rect 316 3121 344 3149
rect 382 3121 410 3149
rect 448 3121 476 3149
rect 514 3121 542 3149
rect 580 3121 608 3149
rect 646 3121 674 3149
rect 712 3121 740 3149
rect -740 3055 -712 3083
rect -674 3055 -646 3083
rect -608 3055 -580 3083
rect -542 3055 -514 3083
rect -476 3055 -448 3083
rect -410 3055 -382 3083
rect -344 3055 -316 3083
rect -278 3055 -250 3083
rect -212 3055 -184 3083
rect -146 3055 -118 3083
rect -80 3055 -52 3083
rect -14 3055 14 3083
rect 52 3055 80 3083
rect 118 3055 146 3083
rect 184 3055 212 3083
rect 250 3055 278 3083
rect 316 3055 344 3083
rect 382 3055 410 3083
rect 448 3055 476 3083
rect 514 3055 542 3083
rect 580 3055 608 3083
rect 646 3055 674 3083
rect 712 3055 740 3083
rect -740 2989 -712 3017
rect -674 2989 -646 3017
rect -608 2989 -580 3017
rect -542 2989 -514 3017
rect -476 2989 -448 3017
rect -410 2989 -382 3017
rect -344 2989 -316 3017
rect -278 2989 -250 3017
rect -212 2989 -184 3017
rect -146 2989 -118 3017
rect -80 2989 -52 3017
rect -14 2989 14 3017
rect 52 2989 80 3017
rect 118 2989 146 3017
rect 184 2989 212 3017
rect 250 2989 278 3017
rect 316 2989 344 3017
rect 382 2989 410 3017
rect 448 2989 476 3017
rect 514 2989 542 3017
rect 580 2989 608 3017
rect 646 2989 674 3017
rect 712 2989 740 3017
rect -740 2923 -712 2951
rect -674 2923 -646 2951
rect -608 2923 -580 2951
rect -542 2923 -514 2951
rect -476 2923 -448 2951
rect -410 2923 -382 2951
rect -344 2923 -316 2951
rect -278 2923 -250 2951
rect -212 2923 -184 2951
rect -146 2923 -118 2951
rect -80 2923 -52 2951
rect -14 2923 14 2951
rect 52 2923 80 2951
rect 118 2923 146 2951
rect 184 2923 212 2951
rect 250 2923 278 2951
rect 316 2923 344 2951
rect 382 2923 410 2951
rect 448 2923 476 2951
rect 514 2923 542 2951
rect 580 2923 608 2951
rect 646 2923 674 2951
rect 712 2923 740 2951
rect -740 2857 -712 2885
rect -674 2857 -646 2885
rect -608 2857 -580 2885
rect -542 2857 -514 2885
rect -476 2857 -448 2885
rect -410 2857 -382 2885
rect -344 2857 -316 2885
rect -278 2857 -250 2885
rect -212 2857 -184 2885
rect -146 2857 -118 2885
rect -80 2857 -52 2885
rect -14 2857 14 2885
rect 52 2857 80 2885
rect 118 2857 146 2885
rect 184 2857 212 2885
rect 250 2857 278 2885
rect 316 2857 344 2885
rect 382 2857 410 2885
rect 448 2857 476 2885
rect 514 2857 542 2885
rect 580 2857 608 2885
rect 646 2857 674 2885
rect 712 2857 740 2885
rect -740 2791 -712 2819
rect -674 2791 -646 2819
rect -608 2791 -580 2819
rect -542 2791 -514 2819
rect -476 2791 -448 2819
rect -410 2791 -382 2819
rect -344 2791 -316 2819
rect -278 2791 -250 2819
rect -212 2791 -184 2819
rect -146 2791 -118 2819
rect -80 2791 -52 2819
rect -14 2791 14 2819
rect 52 2791 80 2819
rect 118 2791 146 2819
rect 184 2791 212 2819
rect 250 2791 278 2819
rect 316 2791 344 2819
rect 382 2791 410 2819
rect 448 2791 476 2819
rect 514 2791 542 2819
rect 580 2791 608 2819
rect 646 2791 674 2819
rect 712 2791 740 2819
rect -740 2725 -712 2753
rect -674 2725 -646 2753
rect -608 2725 -580 2753
rect -542 2725 -514 2753
rect -476 2725 -448 2753
rect -410 2725 -382 2753
rect -344 2725 -316 2753
rect -278 2725 -250 2753
rect -212 2725 -184 2753
rect -146 2725 -118 2753
rect -80 2725 -52 2753
rect -14 2725 14 2753
rect 52 2725 80 2753
rect 118 2725 146 2753
rect 184 2725 212 2753
rect 250 2725 278 2753
rect 316 2725 344 2753
rect 382 2725 410 2753
rect 448 2725 476 2753
rect 514 2725 542 2753
rect 580 2725 608 2753
rect 646 2725 674 2753
rect 712 2725 740 2753
rect -740 2659 -712 2687
rect -674 2659 -646 2687
rect -608 2659 -580 2687
rect -542 2659 -514 2687
rect -476 2659 -448 2687
rect -410 2659 -382 2687
rect -344 2659 -316 2687
rect -278 2659 -250 2687
rect -212 2659 -184 2687
rect -146 2659 -118 2687
rect -80 2659 -52 2687
rect -14 2659 14 2687
rect 52 2659 80 2687
rect 118 2659 146 2687
rect 184 2659 212 2687
rect 250 2659 278 2687
rect 316 2659 344 2687
rect 382 2659 410 2687
rect 448 2659 476 2687
rect 514 2659 542 2687
rect 580 2659 608 2687
rect 646 2659 674 2687
rect 712 2659 740 2687
rect -740 2593 -712 2621
rect -674 2593 -646 2621
rect -608 2593 -580 2621
rect -542 2593 -514 2621
rect -476 2593 -448 2621
rect -410 2593 -382 2621
rect -344 2593 -316 2621
rect -278 2593 -250 2621
rect -212 2593 -184 2621
rect -146 2593 -118 2621
rect -80 2593 -52 2621
rect -14 2593 14 2621
rect 52 2593 80 2621
rect 118 2593 146 2621
rect 184 2593 212 2621
rect 250 2593 278 2621
rect 316 2593 344 2621
rect 382 2593 410 2621
rect 448 2593 476 2621
rect 514 2593 542 2621
rect 580 2593 608 2621
rect 646 2593 674 2621
rect 712 2593 740 2621
rect -740 2527 -712 2555
rect -674 2527 -646 2555
rect -608 2527 -580 2555
rect -542 2527 -514 2555
rect -476 2527 -448 2555
rect -410 2527 -382 2555
rect -344 2527 -316 2555
rect -278 2527 -250 2555
rect -212 2527 -184 2555
rect -146 2527 -118 2555
rect -80 2527 -52 2555
rect -14 2527 14 2555
rect 52 2527 80 2555
rect 118 2527 146 2555
rect 184 2527 212 2555
rect 250 2527 278 2555
rect 316 2527 344 2555
rect 382 2527 410 2555
rect 448 2527 476 2555
rect 514 2527 542 2555
rect 580 2527 608 2555
rect 646 2527 674 2555
rect 712 2527 740 2555
rect -740 2461 -712 2489
rect -674 2461 -646 2489
rect -608 2461 -580 2489
rect -542 2461 -514 2489
rect -476 2461 -448 2489
rect -410 2461 -382 2489
rect -344 2461 -316 2489
rect -278 2461 -250 2489
rect -212 2461 -184 2489
rect -146 2461 -118 2489
rect -80 2461 -52 2489
rect -14 2461 14 2489
rect 52 2461 80 2489
rect 118 2461 146 2489
rect 184 2461 212 2489
rect 250 2461 278 2489
rect 316 2461 344 2489
rect 382 2461 410 2489
rect 448 2461 476 2489
rect 514 2461 542 2489
rect 580 2461 608 2489
rect 646 2461 674 2489
rect 712 2461 740 2489
rect -740 2395 -712 2423
rect -674 2395 -646 2423
rect -608 2395 -580 2423
rect -542 2395 -514 2423
rect -476 2395 -448 2423
rect -410 2395 -382 2423
rect -344 2395 -316 2423
rect -278 2395 -250 2423
rect -212 2395 -184 2423
rect -146 2395 -118 2423
rect -80 2395 -52 2423
rect -14 2395 14 2423
rect 52 2395 80 2423
rect 118 2395 146 2423
rect 184 2395 212 2423
rect 250 2395 278 2423
rect 316 2395 344 2423
rect 382 2395 410 2423
rect 448 2395 476 2423
rect 514 2395 542 2423
rect 580 2395 608 2423
rect 646 2395 674 2423
rect 712 2395 740 2423
rect -740 2329 -712 2357
rect -674 2329 -646 2357
rect -608 2329 -580 2357
rect -542 2329 -514 2357
rect -476 2329 -448 2357
rect -410 2329 -382 2357
rect -344 2329 -316 2357
rect -278 2329 -250 2357
rect -212 2329 -184 2357
rect -146 2329 -118 2357
rect -80 2329 -52 2357
rect -14 2329 14 2357
rect 52 2329 80 2357
rect 118 2329 146 2357
rect 184 2329 212 2357
rect 250 2329 278 2357
rect 316 2329 344 2357
rect 382 2329 410 2357
rect 448 2329 476 2357
rect 514 2329 542 2357
rect 580 2329 608 2357
rect 646 2329 674 2357
rect 712 2329 740 2357
rect -740 2263 -712 2291
rect -674 2263 -646 2291
rect -608 2263 -580 2291
rect -542 2263 -514 2291
rect -476 2263 -448 2291
rect -410 2263 -382 2291
rect -344 2263 -316 2291
rect -278 2263 -250 2291
rect -212 2263 -184 2291
rect -146 2263 -118 2291
rect -80 2263 -52 2291
rect -14 2263 14 2291
rect 52 2263 80 2291
rect 118 2263 146 2291
rect 184 2263 212 2291
rect 250 2263 278 2291
rect 316 2263 344 2291
rect 382 2263 410 2291
rect 448 2263 476 2291
rect 514 2263 542 2291
rect 580 2263 608 2291
rect 646 2263 674 2291
rect 712 2263 740 2291
rect -740 2197 -712 2225
rect -674 2197 -646 2225
rect -608 2197 -580 2225
rect -542 2197 -514 2225
rect -476 2197 -448 2225
rect -410 2197 -382 2225
rect -344 2197 -316 2225
rect -278 2197 -250 2225
rect -212 2197 -184 2225
rect -146 2197 -118 2225
rect -80 2197 -52 2225
rect -14 2197 14 2225
rect 52 2197 80 2225
rect 118 2197 146 2225
rect 184 2197 212 2225
rect 250 2197 278 2225
rect 316 2197 344 2225
rect 382 2197 410 2225
rect 448 2197 476 2225
rect 514 2197 542 2225
rect 580 2197 608 2225
rect 646 2197 674 2225
rect 712 2197 740 2225
rect -740 2131 -712 2159
rect -674 2131 -646 2159
rect -608 2131 -580 2159
rect -542 2131 -514 2159
rect -476 2131 -448 2159
rect -410 2131 -382 2159
rect -344 2131 -316 2159
rect -278 2131 -250 2159
rect -212 2131 -184 2159
rect -146 2131 -118 2159
rect -80 2131 -52 2159
rect -14 2131 14 2159
rect 52 2131 80 2159
rect 118 2131 146 2159
rect 184 2131 212 2159
rect 250 2131 278 2159
rect 316 2131 344 2159
rect 382 2131 410 2159
rect 448 2131 476 2159
rect 514 2131 542 2159
rect 580 2131 608 2159
rect 646 2131 674 2159
rect 712 2131 740 2159
rect -740 2065 -712 2093
rect -674 2065 -646 2093
rect -608 2065 -580 2093
rect -542 2065 -514 2093
rect -476 2065 -448 2093
rect -410 2065 -382 2093
rect -344 2065 -316 2093
rect -278 2065 -250 2093
rect -212 2065 -184 2093
rect -146 2065 -118 2093
rect -80 2065 -52 2093
rect -14 2065 14 2093
rect 52 2065 80 2093
rect 118 2065 146 2093
rect 184 2065 212 2093
rect 250 2065 278 2093
rect 316 2065 344 2093
rect 382 2065 410 2093
rect 448 2065 476 2093
rect 514 2065 542 2093
rect 580 2065 608 2093
rect 646 2065 674 2093
rect 712 2065 740 2093
rect -740 1999 -712 2027
rect -674 1999 -646 2027
rect -608 1999 -580 2027
rect -542 1999 -514 2027
rect -476 1999 -448 2027
rect -410 1999 -382 2027
rect -344 1999 -316 2027
rect -278 1999 -250 2027
rect -212 1999 -184 2027
rect -146 1999 -118 2027
rect -80 1999 -52 2027
rect -14 1999 14 2027
rect 52 1999 80 2027
rect 118 1999 146 2027
rect 184 1999 212 2027
rect 250 1999 278 2027
rect 316 1999 344 2027
rect 382 1999 410 2027
rect 448 1999 476 2027
rect 514 1999 542 2027
rect 580 1999 608 2027
rect 646 1999 674 2027
rect 712 1999 740 2027
rect -740 1933 -712 1961
rect -674 1933 -646 1961
rect -608 1933 -580 1961
rect -542 1933 -514 1961
rect -476 1933 -448 1961
rect -410 1933 -382 1961
rect -344 1933 -316 1961
rect -278 1933 -250 1961
rect -212 1933 -184 1961
rect -146 1933 -118 1961
rect -80 1933 -52 1961
rect -14 1933 14 1961
rect 52 1933 80 1961
rect 118 1933 146 1961
rect 184 1933 212 1961
rect 250 1933 278 1961
rect 316 1933 344 1961
rect 382 1933 410 1961
rect 448 1933 476 1961
rect 514 1933 542 1961
rect 580 1933 608 1961
rect 646 1933 674 1961
rect 712 1933 740 1961
rect -740 1867 -712 1895
rect -674 1867 -646 1895
rect -608 1867 -580 1895
rect -542 1867 -514 1895
rect -476 1867 -448 1895
rect -410 1867 -382 1895
rect -344 1867 -316 1895
rect -278 1867 -250 1895
rect -212 1867 -184 1895
rect -146 1867 -118 1895
rect -80 1867 -52 1895
rect -14 1867 14 1895
rect 52 1867 80 1895
rect 118 1867 146 1895
rect 184 1867 212 1895
rect 250 1867 278 1895
rect 316 1867 344 1895
rect 382 1867 410 1895
rect 448 1867 476 1895
rect 514 1867 542 1895
rect 580 1867 608 1895
rect 646 1867 674 1895
rect 712 1867 740 1895
rect -740 1801 -712 1829
rect -674 1801 -646 1829
rect -608 1801 -580 1829
rect -542 1801 -514 1829
rect -476 1801 -448 1829
rect -410 1801 -382 1829
rect -344 1801 -316 1829
rect -278 1801 -250 1829
rect -212 1801 -184 1829
rect -146 1801 -118 1829
rect -80 1801 -52 1829
rect -14 1801 14 1829
rect 52 1801 80 1829
rect 118 1801 146 1829
rect 184 1801 212 1829
rect 250 1801 278 1829
rect 316 1801 344 1829
rect 382 1801 410 1829
rect 448 1801 476 1829
rect 514 1801 542 1829
rect 580 1801 608 1829
rect 646 1801 674 1829
rect 712 1801 740 1829
rect -740 1735 -712 1763
rect -674 1735 -646 1763
rect -608 1735 -580 1763
rect -542 1735 -514 1763
rect -476 1735 -448 1763
rect -410 1735 -382 1763
rect -344 1735 -316 1763
rect -278 1735 -250 1763
rect -212 1735 -184 1763
rect -146 1735 -118 1763
rect -80 1735 -52 1763
rect -14 1735 14 1763
rect 52 1735 80 1763
rect 118 1735 146 1763
rect 184 1735 212 1763
rect 250 1735 278 1763
rect 316 1735 344 1763
rect 382 1735 410 1763
rect 448 1735 476 1763
rect 514 1735 542 1763
rect 580 1735 608 1763
rect 646 1735 674 1763
rect 712 1735 740 1763
rect -740 1669 -712 1697
rect -674 1669 -646 1697
rect -608 1669 -580 1697
rect -542 1669 -514 1697
rect -476 1669 -448 1697
rect -410 1669 -382 1697
rect -344 1669 -316 1697
rect -278 1669 -250 1697
rect -212 1669 -184 1697
rect -146 1669 -118 1697
rect -80 1669 -52 1697
rect -14 1669 14 1697
rect 52 1669 80 1697
rect 118 1669 146 1697
rect 184 1669 212 1697
rect 250 1669 278 1697
rect 316 1669 344 1697
rect 382 1669 410 1697
rect 448 1669 476 1697
rect 514 1669 542 1697
rect 580 1669 608 1697
rect 646 1669 674 1697
rect 712 1669 740 1697
rect -740 1603 -712 1631
rect -674 1603 -646 1631
rect -608 1603 -580 1631
rect -542 1603 -514 1631
rect -476 1603 -448 1631
rect -410 1603 -382 1631
rect -344 1603 -316 1631
rect -278 1603 -250 1631
rect -212 1603 -184 1631
rect -146 1603 -118 1631
rect -80 1603 -52 1631
rect -14 1603 14 1631
rect 52 1603 80 1631
rect 118 1603 146 1631
rect 184 1603 212 1631
rect 250 1603 278 1631
rect 316 1603 344 1631
rect 382 1603 410 1631
rect 448 1603 476 1631
rect 514 1603 542 1631
rect 580 1603 608 1631
rect 646 1603 674 1631
rect 712 1603 740 1631
rect -740 1537 -712 1565
rect -674 1537 -646 1565
rect -608 1537 -580 1565
rect -542 1537 -514 1565
rect -476 1537 -448 1565
rect -410 1537 -382 1565
rect -344 1537 -316 1565
rect -278 1537 -250 1565
rect -212 1537 -184 1565
rect -146 1537 -118 1565
rect -80 1537 -52 1565
rect -14 1537 14 1565
rect 52 1537 80 1565
rect 118 1537 146 1565
rect 184 1537 212 1565
rect 250 1537 278 1565
rect 316 1537 344 1565
rect 382 1537 410 1565
rect 448 1537 476 1565
rect 514 1537 542 1565
rect 580 1537 608 1565
rect 646 1537 674 1565
rect 712 1537 740 1565
rect -740 1471 -712 1499
rect -674 1471 -646 1499
rect -608 1471 -580 1499
rect -542 1471 -514 1499
rect -476 1471 -448 1499
rect -410 1471 -382 1499
rect -344 1471 -316 1499
rect -278 1471 -250 1499
rect -212 1471 -184 1499
rect -146 1471 -118 1499
rect -80 1471 -52 1499
rect -14 1471 14 1499
rect 52 1471 80 1499
rect 118 1471 146 1499
rect 184 1471 212 1499
rect 250 1471 278 1499
rect 316 1471 344 1499
rect 382 1471 410 1499
rect 448 1471 476 1499
rect 514 1471 542 1499
rect 580 1471 608 1499
rect 646 1471 674 1499
rect 712 1471 740 1499
rect -740 1405 -712 1433
rect -674 1405 -646 1433
rect -608 1405 -580 1433
rect -542 1405 -514 1433
rect -476 1405 -448 1433
rect -410 1405 -382 1433
rect -344 1405 -316 1433
rect -278 1405 -250 1433
rect -212 1405 -184 1433
rect -146 1405 -118 1433
rect -80 1405 -52 1433
rect -14 1405 14 1433
rect 52 1405 80 1433
rect 118 1405 146 1433
rect 184 1405 212 1433
rect 250 1405 278 1433
rect 316 1405 344 1433
rect 382 1405 410 1433
rect 448 1405 476 1433
rect 514 1405 542 1433
rect 580 1405 608 1433
rect 646 1405 674 1433
rect 712 1405 740 1433
rect -740 1339 -712 1367
rect -674 1339 -646 1367
rect -608 1339 -580 1367
rect -542 1339 -514 1367
rect -476 1339 -448 1367
rect -410 1339 -382 1367
rect -344 1339 -316 1367
rect -278 1339 -250 1367
rect -212 1339 -184 1367
rect -146 1339 -118 1367
rect -80 1339 -52 1367
rect -14 1339 14 1367
rect 52 1339 80 1367
rect 118 1339 146 1367
rect 184 1339 212 1367
rect 250 1339 278 1367
rect 316 1339 344 1367
rect 382 1339 410 1367
rect 448 1339 476 1367
rect 514 1339 542 1367
rect 580 1339 608 1367
rect 646 1339 674 1367
rect 712 1339 740 1367
rect -740 1273 -712 1301
rect -674 1273 -646 1301
rect -608 1273 -580 1301
rect -542 1273 -514 1301
rect -476 1273 -448 1301
rect -410 1273 -382 1301
rect -344 1273 -316 1301
rect -278 1273 -250 1301
rect -212 1273 -184 1301
rect -146 1273 -118 1301
rect -80 1273 -52 1301
rect -14 1273 14 1301
rect 52 1273 80 1301
rect 118 1273 146 1301
rect 184 1273 212 1301
rect 250 1273 278 1301
rect 316 1273 344 1301
rect 382 1273 410 1301
rect 448 1273 476 1301
rect 514 1273 542 1301
rect 580 1273 608 1301
rect 646 1273 674 1301
rect 712 1273 740 1301
rect -740 1207 -712 1235
rect -674 1207 -646 1235
rect -608 1207 -580 1235
rect -542 1207 -514 1235
rect -476 1207 -448 1235
rect -410 1207 -382 1235
rect -344 1207 -316 1235
rect -278 1207 -250 1235
rect -212 1207 -184 1235
rect -146 1207 -118 1235
rect -80 1207 -52 1235
rect -14 1207 14 1235
rect 52 1207 80 1235
rect 118 1207 146 1235
rect 184 1207 212 1235
rect 250 1207 278 1235
rect 316 1207 344 1235
rect 382 1207 410 1235
rect 448 1207 476 1235
rect 514 1207 542 1235
rect 580 1207 608 1235
rect 646 1207 674 1235
rect 712 1207 740 1235
rect -740 1141 -712 1169
rect -674 1141 -646 1169
rect -608 1141 -580 1169
rect -542 1141 -514 1169
rect -476 1141 -448 1169
rect -410 1141 -382 1169
rect -344 1141 -316 1169
rect -278 1141 -250 1169
rect -212 1141 -184 1169
rect -146 1141 -118 1169
rect -80 1141 -52 1169
rect -14 1141 14 1169
rect 52 1141 80 1169
rect 118 1141 146 1169
rect 184 1141 212 1169
rect 250 1141 278 1169
rect 316 1141 344 1169
rect 382 1141 410 1169
rect 448 1141 476 1169
rect 514 1141 542 1169
rect 580 1141 608 1169
rect 646 1141 674 1169
rect 712 1141 740 1169
rect -740 1075 -712 1103
rect -674 1075 -646 1103
rect -608 1075 -580 1103
rect -542 1075 -514 1103
rect -476 1075 -448 1103
rect -410 1075 -382 1103
rect -344 1075 -316 1103
rect -278 1075 -250 1103
rect -212 1075 -184 1103
rect -146 1075 -118 1103
rect -80 1075 -52 1103
rect -14 1075 14 1103
rect 52 1075 80 1103
rect 118 1075 146 1103
rect 184 1075 212 1103
rect 250 1075 278 1103
rect 316 1075 344 1103
rect 382 1075 410 1103
rect 448 1075 476 1103
rect 514 1075 542 1103
rect 580 1075 608 1103
rect 646 1075 674 1103
rect 712 1075 740 1103
rect -740 1009 -712 1037
rect -674 1009 -646 1037
rect -608 1009 -580 1037
rect -542 1009 -514 1037
rect -476 1009 -448 1037
rect -410 1009 -382 1037
rect -344 1009 -316 1037
rect -278 1009 -250 1037
rect -212 1009 -184 1037
rect -146 1009 -118 1037
rect -80 1009 -52 1037
rect -14 1009 14 1037
rect 52 1009 80 1037
rect 118 1009 146 1037
rect 184 1009 212 1037
rect 250 1009 278 1037
rect 316 1009 344 1037
rect 382 1009 410 1037
rect 448 1009 476 1037
rect 514 1009 542 1037
rect 580 1009 608 1037
rect 646 1009 674 1037
rect 712 1009 740 1037
rect -740 943 -712 971
rect -674 943 -646 971
rect -608 943 -580 971
rect -542 943 -514 971
rect -476 943 -448 971
rect -410 943 -382 971
rect -344 943 -316 971
rect -278 943 -250 971
rect -212 943 -184 971
rect -146 943 -118 971
rect -80 943 -52 971
rect -14 943 14 971
rect 52 943 80 971
rect 118 943 146 971
rect 184 943 212 971
rect 250 943 278 971
rect 316 943 344 971
rect 382 943 410 971
rect 448 943 476 971
rect 514 943 542 971
rect 580 943 608 971
rect 646 943 674 971
rect 712 943 740 971
rect -740 877 -712 905
rect -674 877 -646 905
rect -608 877 -580 905
rect -542 877 -514 905
rect -476 877 -448 905
rect -410 877 -382 905
rect -344 877 -316 905
rect -278 877 -250 905
rect -212 877 -184 905
rect -146 877 -118 905
rect -80 877 -52 905
rect -14 877 14 905
rect 52 877 80 905
rect 118 877 146 905
rect 184 877 212 905
rect 250 877 278 905
rect 316 877 344 905
rect 382 877 410 905
rect 448 877 476 905
rect 514 877 542 905
rect 580 877 608 905
rect 646 877 674 905
rect 712 877 740 905
rect -740 811 -712 839
rect -674 811 -646 839
rect -608 811 -580 839
rect -542 811 -514 839
rect -476 811 -448 839
rect -410 811 -382 839
rect -344 811 -316 839
rect -278 811 -250 839
rect -212 811 -184 839
rect -146 811 -118 839
rect -80 811 -52 839
rect -14 811 14 839
rect 52 811 80 839
rect 118 811 146 839
rect 184 811 212 839
rect 250 811 278 839
rect 316 811 344 839
rect 382 811 410 839
rect 448 811 476 839
rect 514 811 542 839
rect 580 811 608 839
rect 646 811 674 839
rect 712 811 740 839
rect -740 745 -712 773
rect -674 745 -646 773
rect -608 745 -580 773
rect -542 745 -514 773
rect -476 745 -448 773
rect -410 745 -382 773
rect -344 745 -316 773
rect -278 745 -250 773
rect -212 745 -184 773
rect -146 745 -118 773
rect -80 745 -52 773
rect -14 745 14 773
rect 52 745 80 773
rect 118 745 146 773
rect 184 745 212 773
rect 250 745 278 773
rect 316 745 344 773
rect 382 745 410 773
rect 448 745 476 773
rect 514 745 542 773
rect 580 745 608 773
rect 646 745 674 773
rect 712 745 740 773
rect -740 679 -712 707
rect -674 679 -646 707
rect -608 679 -580 707
rect -542 679 -514 707
rect -476 679 -448 707
rect -410 679 -382 707
rect -344 679 -316 707
rect -278 679 -250 707
rect -212 679 -184 707
rect -146 679 -118 707
rect -80 679 -52 707
rect -14 679 14 707
rect 52 679 80 707
rect 118 679 146 707
rect 184 679 212 707
rect 250 679 278 707
rect 316 679 344 707
rect 382 679 410 707
rect 448 679 476 707
rect 514 679 542 707
rect 580 679 608 707
rect 646 679 674 707
rect 712 679 740 707
rect -740 613 -712 641
rect -674 613 -646 641
rect -608 613 -580 641
rect -542 613 -514 641
rect -476 613 -448 641
rect -410 613 -382 641
rect -344 613 -316 641
rect -278 613 -250 641
rect -212 613 -184 641
rect -146 613 -118 641
rect -80 613 -52 641
rect -14 613 14 641
rect 52 613 80 641
rect 118 613 146 641
rect 184 613 212 641
rect 250 613 278 641
rect 316 613 344 641
rect 382 613 410 641
rect 448 613 476 641
rect 514 613 542 641
rect 580 613 608 641
rect 646 613 674 641
rect 712 613 740 641
rect -740 547 -712 575
rect -674 547 -646 575
rect -608 547 -580 575
rect -542 547 -514 575
rect -476 547 -448 575
rect -410 547 -382 575
rect -344 547 -316 575
rect -278 547 -250 575
rect -212 547 -184 575
rect -146 547 -118 575
rect -80 547 -52 575
rect -14 547 14 575
rect 52 547 80 575
rect 118 547 146 575
rect 184 547 212 575
rect 250 547 278 575
rect 316 547 344 575
rect 382 547 410 575
rect 448 547 476 575
rect 514 547 542 575
rect 580 547 608 575
rect 646 547 674 575
rect 712 547 740 575
rect -740 481 -712 509
rect -674 481 -646 509
rect -608 481 -580 509
rect -542 481 -514 509
rect -476 481 -448 509
rect -410 481 -382 509
rect -344 481 -316 509
rect -278 481 -250 509
rect -212 481 -184 509
rect -146 481 -118 509
rect -80 481 -52 509
rect -14 481 14 509
rect 52 481 80 509
rect 118 481 146 509
rect 184 481 212 509
rect 250 481 278 509
rect 316 481 344 509
rect 382 481 410 509
rect 448 481 476 509
rect 514 481 542 509
rect 580 481 608 509
rect 646 481 674 509
rect 712 481 740 509
rect -740 415 -712 443
rect -674 415 -646 443
rect -608 415 -580 443
rect -542 415 -514 443
rect -476 415 -448 443
rect -410 415 -382 443
rect -344 415 -316 443
rect -278 415 -250 443
rect -212 415 -184 443
rect -146 415 -118 443
rect -80 415 -52 443
rect -14 415 14 443
rect 52 415 80 443
rect 118 415 146 443
rect 184 415 212 443
rect 250 415 278 443
rect 316 415 344 443
rect 382 415 410 443
rect 448 415 476 443
rect 514 415 542 443
rect 580 415 608 443
rect 646 415 674 443
rect 712 415 740 443
rect -740 349 -712 377
rect -674 349 -646 377
rect -608 349 -580 377
rect -542 349 -514 377
rect -476 349 -448 377
rect -410 349 -382 377
rect -344 349 -316 377
rect -278 349 -250 377
rect -212 349 -184 377
rect -146 349 -118 377
rect -80 349 -52 377
rect -14 349 14 377
rect 52 349 80 377
rect 118 349 146 377
rect 184 349 212 377
rect 250 349 278 377
rect 316 349 344 377
rect 382 349 410 377
rect 448 349 476 377
rect 514 349 542 377
rect 580 349 608 377
rect 646 349 674 377
rect 712 349 740 377
rect -740 283 -712 311
rect -674 283 -646 311
rect -608 283 -580 311
rect -542 283 -514 311
rect -476 283 -448 311
rect -410 283 -382 311
rect -344 283 -316 311
rect -278 283 -250 311
rect -212 283 -184 311
rect -146 283 -118 311
rect -80 283 -52 311
rect -14 283 14 311
rect 52 283 80 311
rect 118 283 146 311
rect 184 283 212 311
rect 250 283 278 311
rect 316 283 344 311
rect 382 283 410 311
rect 448 283 476 311
rect 514 283 542 311
rect 580 283 608 311
rect 646 283 674 311
rect 712 283 740 311
rect -740 217 -712 245
rect -674 217 -646 245
rect -608 217 -580 245
rect -542 217 -514 245
rect -476 217 -448 245
rect -410 217 -382 245
rect -344 217 -316 245
rect -278 217 -250 245
rect -212 217 -184 245
rect -146 217 -118 245
rect -80 217 -52 245
rect -14 217 14 245
rect 52 217 80 245
rect 118 217 146 245
rect 184 217 212 245
rect 250 217 278 245
rect 316 217 344 245
rect 382 217 410 245
rect 448 217 476 245
rect 514 217 542 245
rect 580 217 608 245
rect 646 217 674 245
rect 712 217 740 245
rect -740 151 -712 179
rect -674 151 -646 179
rect -608 151 -580 179
rect -542 151 -514 179
rect -476 151 -448 179
rect -410 151 -382 179
rect -344 151 -316 179
rect -278 151 -250 179
rect -212 151 -184 179
rect -146 151 -118 179
rect -80 151 -52 179
rect -14 151 14 179
rect 52 151 80 179
rect 118 151 146 179
rect 184 151 212 179
rect 250 151 278 179
rect 316 151 344 179
rect 382 151 410 179
rect 448 151 476 179
rect 514 151 542 179
rect 580 151 608 179
rect 646 151 674 179
rect 712 151 740 179
rect -740 85 -712 113
rect -674 85 -646 113
rect -608 85 -580 113
rect -542 85 -514 113
rect -476 85 -448 113
rect -410 85 -382 113
rect -344 85 -316 113
rect -278 85 -250 113
rect -212 85 -184 113
rect -146 85 -118 113
rect -80 85 -52 113
rect -14 85 14 113
rect 52 85 80 113
rect 118 85 146 113
rect 184 85 212 113
rect 250 85 278 113
rect 316 85 344 113
rect 382 85 410 113
rect 448 85 476 113
rect 514 85 542 113
rect 580 85 608 113
rect 646 85 674 113
rect 712 85 740 113
rect -740 19 -712 47
rect -674 19 -646 47
rect -608 19 -580 47
rect -542 19 -514 47
rect -476 19 -448 47
rect -410 19 -382 47
rect -344 19 -316 47
rect -278 19 -250 47
rect -212 19 -184 47
rect -146 19 -118 47
rect -80 19 -52 47
rect -14 19 14 47
rect 52 19 80 47
rect 118 19 146 47
rect 184 19 212 47
rect 250 19 278 47
rect 316 19 344 47
rect 382 19 410 47
rect 448 19 476 47
rect 514 19 542 47
rect 580 19 608 47
rect 646 19 674 47
rect 712 19 740 47
rect -740 -47 -712 -19
rect -674 -47 -646 -19
rect -608 -47 -580 -19
rect -542 -47 -514 -19
rect -476 -47 -448 -19
rect -410 -47 -382 -19
rect -344 -47 -316 -19
rect -278 -47 -250 -19
rect -212 -47 -184 -19
rect -146 -47 -118 -19
rect -80 -47 -52 -19
rect -14 -47 14 -19
rect 52 -47 80 -19
rect 118 -47 146 -19
rect 184 -47 212 -19
rect 250 -47 278 -19
rect 316 -47 344 -19
rect 382 -47 410 -19
rect 448 -47 476 -19
rect 514 -47 542 -19
rect 580 -47 608 -19
rect 646 -47 674 -19
rect 712 -47 740 -19
rect -740 -113 -712 -85
rect -674 -113 -646 -85
rect -608 -113 -580 -85
rect -542 -113 -514 -85
rect -476 -113 -448 -85
rect -410 -113 -382 -85
rect -344 -113 -316 -85
rect -278 -113 -250 -85
rect -212 -113 -184 -85
rect -146 -113 -118 -85
rect -80 -113 -52 -85
rect -14 -113 14 -85
rect 52 -113 80 -85
rect 118 -113 146 -85
rect 184 -113 212 -85
rect 250 -113 278 -85
rect 316 -113 344 -85
rect 382 -113 410 -85
rect 448 -113 476 -85
rect 514 -113 542 -85
rect 580 -113 608 -85
rect 646 -113 674 -85
rect 712 -113 740 -85
rect -740 -179 -712 -151
rect -674 -179 -646 -151
rect -608 -179 -580 -151
rect -542 -179 -514 -151
rect -476 -179 -448 -151
rect -410 -179 -382 -151
rect -344 -179 -316 -151
rect -278 -179 -250 -151
rect -212 -179 -184 -151
rect -146 -179 -118 -151
rect -80 -179 -52 -151
rect -14 -179 14 -151
rect 52 -179 80 -151
rect 118 -179 146 -151
rect 184 -179 212 -151
rect 250 -179 278 -151
rect 316 -179 344 -151
rect 382 -179 410 -151
rect 448 -179 476 -151
rect 514 -179 542 -151
rect 580 -179 608 -151
rect 646 -179 674 -151
rect 712 -179 740 -151
rect -740 -245 -712 -217
rect -674 -245 -646 -217
rect -608 -245 -580 -217
rect -542 -245 -514 -217
rect -476 -245 -448 -217
rect -410 -245 -382 -217
rect -344 -245 -316 -217
rect -278 -245 -250 -217
rect -212 -245 -184 -217
rect -146 -245 -118 -217
rect -80 -245 -52 -217
rect -14 -245 14 -217
rect 52 -245 80 -217
rect 118 -245 146 -217
rect 184 -245 212 -217
rect 250 -245 278 -217
rect 316 -245 344 -217
rect 382 -245 410 -217
rect 448 -245 476 -217
rect 514 -245 542 -217
rect 580 -245 608 -217
rect 646 -245 674 -217
rect 712 -245 740 -217
rect -740 -311 -712 -283
rect -674 -311 -646 -283
rect -608 -311 -580 -283
rect -542 -311 -514 -283
rect -476 -311 -448 -283
rect -410 -311 -382 -283
rect -344 -311 -316 -283
rect -278 -311 -250 -283
rect -212 -311 -184 -283
rect -146 -311 -118 -283
rect -80 -311 -52 -283
rect -14 -311 14 -283
rect 52 -311 80 -283
rect 118 -311 146 -283
rect 184 -311 212 -283
rect 250 -311 278 -283
rect 316 -311 344 -283
rect 382 -311 410 -283
rect 448 -311 476 -283
rect 514 -311 542 -283
rect 580 -311 608 -283
rect 646 -311 674 -283
rect 712 -311 740 -283
rect -740 -377 -712 -349
rect -674 -377 -646 -349
rect -608 -377 -580 -349
rect -542 -377 -514 -349
rect -476 -377 -448 -349
rect -410 -377 -382 -349
rect -344 -377 -316 -349
rect -278 -377 -250 -349
rect -212 -377 -184 -349
rect -146 -377 -118 -349
rect -80 -377 -52 -349
rect -14 -377 14 -349
rect 52 -377 80 -349
rect 118 -377 146 -349
rect 184 -377 212 -349
rect 250 -377 278 -349
rect 316 -377 344 -349
rect 382 -377 410 -349
rect 448 -377 476 -349
rect 514 -377 542 -349
rect 580 -377 608 -349
rect 646 -377 674 -349
rect 712 -377 740 -349
rect -740 -443 -712 -415
rect -674 -443 -646 -415
rect -608 -443 -580 -415
rect -542 -443 -514 -415
rect -476 -443 -448 -415
rect -410 -443 -382 -415
rect -344 -443 -316 -415
rect -278 -443 -250 -415
rect -212 -443 -184 -415
rect -146 -443 -118 -415
rect -80 -443 -52 -415
rect -14 -443 14 -415
rect 52 -443 80 -415
rect 118 -443 146 -415
rect 184 -443 212 -415
rect 250 -443 278 -415
rect 316 -443 344 -415
rect 382 -443 410 -415
rect 448 -443 476 -415
rect 514 -443 542 -415
rect 580 -443 608 -415
rect 646 -443 674 -415
rect 712 -443 740 -415
rect -740 -509 -712 -481
rect -674 -509 -646 -481
rect -608 -509 -580 -481
rect -542 -509 -514 -481
rect -476 -509 -448 -481
rect -410 -509 -382 -481
rect -344 -509 -316 -481
rect -278 -509 -250 -481
rect -212 -509 -184 -481
rect -146 -509 -118 -481
rect -80 -509 -52 -481
rect -14 -509 14 -481
rect 52 -509 80 -481
rect 118 -509 146 -481
rect 184 -509 212 -481
rect 250 -509 278 -481
rect 316 -509 344 -481
rect 382 -509 410 -481
rect 448 -509 476 -481
rect 514 -509 542 -481
rect 580 -509 608 -481
rect 646 -509 674 -481
rect 712 -509 740 -481
rect -740 -575 -712 -547
rect -674 -575 -646 -547
rect -608 -575 -580 -547
rect -542 -575 -514 -547
rect -476 -575 -448 -547
rect -410 -575 -382 -547
rect -344 -575 -316 -547
rect -278 -575 -250 -547
rect -212 -575 -184 -547
rect -146 -575 -118 -547
rect -80 -575 -52 -547
rect -14 -575 14 -547
rect 52 -575 80 -547
rect 118 -575 146 -547
rect 184 -575 212 -547
rect 250 -575 278 -547
rect 316 -575 344 -547
rect 382 -575 410 -547
rect 448 -575 476 -547
rect 514 -575 542 -547
rect 580 -575 608 -547
rect 646 -575 674 -547
rect 712 -575 740 -547
rect -740 -641 -712 -613
rect -674 -641 -646 -613
rect -608 -641 -580 -613
rect -542 -641 -514 -613
rect -476 -641 -448 -613
rect -410 -641 -382 -613
rect -344 -641 -316 -613
rect -278 -641 -250 -613
rect -212 -641 -184 -613
rect -146 -641 -118 -613
rect -80 -641 -52 -613
rect -14 -641 14 -613
rect 52 -641 80 -613
rect 118 -641 146 -613
rect 184 -641 212 -613
rect 250 -641 278 -613
rect 316 -641 344 -613
rect 382 -641 410 -613
rect 448 -641 476 -613
rect 514 -641 542 -613
rect 580 -641 608 -613
rect 646 -641 674 -613
rect 712 -641 740 -613
rect -740 -707 -712 -679
rect -674 -707 -646 -679
rect -608 -707 -580 -679
rect -542 -707 -514 -679
rect -476 -707 -448 -679
rect -410 -707 -382 -679
rect -344 -707 -316 -679
rect -278 -707 -250 -679
rect -212 -707 -184 -679
rect -146 -707 -118 -679
rect -80 -707 -52 -679
rect -14 -707 14 -679
rect 52 -707 80 -679
rect 118 -707 146 -679
rect 184 -707 212 -679
rect 250 -707 278 -679
rect 316 -707 344 -679
rect 382 -707 410 -679
rect 448 -707 476 -679
rect 514 -707 542 -679
rect 580 -707 608 -679
rect 646 -707 674 -679
rect 712 -707 740 -679
rect -740 -773 -712 -745
rect -674 -773 -646 -745
rect -608 -773 -580 -745
rect -542 -773 -514 -745
rect -476 -773 -448 -745
rect -410 -773 -382 -745
rect -344 -773 -316 -745
rect -278 -773 -250 -745
rect -212 -773 -184 -745
rect -146 -773 -118 -745
rect -80 -773 -52 -745
rect -14 -773 14 -745
rect 52 -773 80 -745
rect 118 -773 146 -745
rect 184 -773 212 -745
rect 250 -773 278 -745
rect 316 -773 344 -745
rect 382 -773 410 -745
rect 448 -773 476 -745
rect 514 -773 542 -745
rect 580 -773 608 -745
rect 646 -773 674 -745
rect 712 -773 740 -745
rect -740 -839 -712 -811
rect -674 -839 -646 -811
rect -608 -839 -580 -811
rect -542 -839 -514 -811
rect -476 -839 -448 -811
rect -410 -839 -382 -811
rect -344 -839 -316 -811
rect -278 -839 -250 -811
rect -212 -839 -184 -811
rect -146 -839 -118 -811
rect -80 -839 -52 -811
rect -14 -839 14 -811
rect 52 -839 80 -811
rect 118 -839 146 -811
rect 184 -839 212 -811
rect 250 -839 278 -811
rect 316 -839 344 -811
rect 382 -839 410 -811
rect 448 -839 476 -811
rect 514 -839 542 -811
rect 580 -839 608 -811
rect 646 -839 674 -811
rect 712 -839 740 -811
rect -740 -905 -712 -877
rect -674 -905 -646 -877
rect -608 -905 -580 -877
rect -542 -905 -514 -877
rect -476 -905 -448 -877
rect -410 -905 -382 -877
rect -344 -905 -316 -877
rect -278 -905 -250 -877
rect -212 -905 -184 -877
rect -146 -905 -118 -877
rect -80 -905 -52 -877
rect -14 -905 14 -877
rect 52 -905 80 -877
rect 118 -905 146 -877
rect 184 -905 212 -877
rect 250 -905 278 -877
rect 316 -905 344 -877
rect 382 -905 410 -877
rect 448 -905 476 -877
rect 514 -905 542 -877
rect 580 -905 608 -877
rect 646 -905 674 -877
rect 712 -905 740 -877
rect -740 -971 -712 -943
rect -674 -971 -646 -943
rect -608 -971 -580 -943
rect -542 -971 -514 -943
rect -476 -971 -448 -943
rect -410 -971 -382 -943
rect -344 -971 -316 -943
rect -278 -971 -250 -943
rect -212 -971 -184 -943
rect -146 -971 -118 -943
rect -80 -971 -52 -943
rect -14 -971 14 -943
rect 52 -971 80 -943
rect 118 -971 146 -943
rect 184 -971 212 -943
rect 250 -971 278 -943
rect 316 -971 344 -943
rect 382 -971 410 -943
rect 448 -971 476 -943
rect 514 -971 542 -943
rect 580 -971 608 -943
rect 646 -971 674 -943
rect 712 -971 740 -943
rect -740 -1037 -712 -1009
rect -674 -1037 -646 -1009
rect -608 -1037 -580 -1009
rect -542 -1037 -514 -1009
rect -476 -1037 -448 -1009
rect -410 -1037 -382 -1009
rect -344 -1037 -316 -1009
rect -278 -1037 -250 -1009
rect -212 -1037 -184 -1009
rect -146 -1037 -118 -1009
rect -80 -1037 -52 -1009
rect -14 -1037 14 -1009
rect 52 -1037 80 -1009
rect 118 -1037 146 -1009
rect 184 -1037 212 -1009
rect 250 -1037 278 -1009
rect 316 -1037 344 -1009
rect 382 -1037 410 -1009
rect 448 -1037 476 -1009
rect 514 -1037 542 -1009
rect 580 -1037 608 -1009
rect 646 -1037 674 -1009
rect 712 -1037 740 -1009
rect -740 -1103 -712 -1075
rect -674 -1103 -646 -1075
rect -608 -1103 -580 -1075
rect -542 -1103 -514 -1075
rect -476 -1103 -448 -1075
rect -410 -1103 -382 -1075
rect -344 -1103 -316 -1075
rect -278 -1103 -250 -1075
rect -212 -1103 -184 -1075
rect -146 -1103 -118 -1075
rect -80 -1103 -52 -1075
rect -14 -1103 14 -1075
rect 52 -1103 80 -1075
rect 118 -1103 146 -1075
rect 184 -1103 212 -1075
rect 250 -1103 278 -1075
rect 316 -1103 344 -1075
rect 382 -1103 410 -1075
rect 448 -1103 476 -1075
rect 514 -1103 542 -1075
rect 580 -1103 608 -1075
rect 646 -1103 674 -1075
rect 712 -1103 740 -1075
rect -740 -1169 -712 -1141
rect -674 -1169 -646 -1141
rect -608 -1169 -580 -1141
rect -542 -1169 -514 -1141
rect -476 -1169 -448 -1141
rect -410 -1169 -382 -1141
rect -344 -1169 -316 -1141
rect -278 -1169 -250 -1141
rect -212 -1169 -184 -1141
rect -146 -1169 -118 -1141
rect -80 -1169 -52 -1141
rect -14 -1169 14 -1141
rect 52 -1169 80 -1141
rect 118 -1169 146 -1141
rect 184 -1169 212 -1141
rect 250 -1169 278 -1141
rect 316 -1169 344 -1141
rect 382 -1169 410 -1141
rect 448 -1169 476 -1141
rect 514 -1169 542 -1141
rect 580 -1169 608 -1141
rect 646 -1169 674 -1141
rect 712 -1169 740 -1141
rect -740 -1235 -712 -1207
rect -674 -1235 -646 -1207
rect -608 -1235 -580 -1207
rect -542 -1235 -514 -1207
rect -476 -1235 -448 -1207
rect -410 -1235 -382 -1207
rect -344 -1235 -316 -1207
rect -278 -1235 -250 -1207
rect -212 -1235 -184 -1207
rect -146 -1235 -118 -1207
rect -80 -1235 -52 -1207
rect -14 -1235 14 -1207
rect 52 -1235 80 -1207
rect 118 -1235 146 -1207
rect 184 -1235 212 -1207
rect 250 -1235 278 -1207
rect 316 -1235 344 -1207
rect 382 -1235 410 -1207
rect 448 -1235 476 -1207
rect 514 -1235 542 -1207
rect 580 -1235 608 -1207
rect 646 -1235 674 -1207
rect 712 -1235 740 -1207
rect -740 -1301 -712 -1273
rect -674 -1301 -646 -1273
rect -608 -1301 -580 -1273
rect -542 -1301 -514 -1273
rect -476 -1301 -448 -1273
rect -410 -1301 -382 -1273
rect -344 -1301 -316 -1273
rect -278 -1301 -250 -1273
rect -212 -1301 -184 -1273
rect -146 -1301 -118 -1273
rect -80 -1301 -52 -1273
rect -14 -1301 14 -1273
rect 52 -1301 80 -1273
rect 118 -1301 146 -1273
rect 184 -1301 212 -1273
rect 250 -1301 278 -1273
rect 316 -1301 344 -1273
rect 382 -1301 410 -1273
rect 448 -1301 476 -1273
rect 514 -1301 542 -1273
rect 580 -1301 608 -1273
rect 646 -1301 674 -1273
rect 712 -1301 740 -1273
rect -740 -1367 -712 -1339
rect -674 -1367 -646 -1339
rect -608 -1367 -580 -1339
rect -542 -1367 -514 -1339
rect -476 -1367 -448 -1339
rect -410 -1367 -382 -1339
rect -344 -1367 -316 -1339
rect -278 -1367 -250 -1339
rect -212 -1367 -184 -1339
rect -146 -1367 -118 -1339
rect -80 -1367 -52 -1339
rect -14 -1367 14 -1339
rect 52 -1367 80 -1339
rect 118 -1367 146 -1339
rect 184 -1367 212 -1339
rect 250 -1367 278 -1339
rect 316 -1367 344 -1339
rect 382 -1367 410 -1339
rect 448 -1367 476 -1339
rect 514 -1367 542 -1339
rect 580 -1367 608 -1339
rect 646 -1367 674 -1339
rect 712 -1367 740 -1339
rect -740 -1433 -712 -1405
rect -674 -1433 -646 -1405
rect -608 -1433 -580 -1405
rect -542 -1433 -514 -1405
rect -476 -1433 -448 -1405
rect -410 -1433 -382 -1405
rect -344 -1433 -316 -1405
rect -278 -1433 -250 -1405
rect -212 -1433 -184 -1405
rect -146 -1433 -118 -1405
rect -80 -1433 -52 -1405
rect -14 -1433 14 -1405
rect 52 -1433 80 -1405
rect 118 -1433 146 -1405
rect 184 -1433 212 -1405
rect 250 -1433 278 -1405
rect 316 -1433 344 -1405
rect 382 -1433 410 -1405
rect 448 -1433 476 -1405
rect 514 -1433 542 -1405
rect 580 -1433 608 -1405
rect 646 -1433 674 -1405
rect 712 -1433 740 -1405
rect -740 -1499 -712 -1471
rect -674 -1499 -646 -1471
rect -608 -1499 -580 -1471
rect -542 -1499 -514 -1471
rect -476 -1499 -448 -1471
rect -410 -1499 -382 -1471
rect -344 -1499 -316 -1471
rect -278 -1499 -250 -1471
rect -212 -1499 -184 -1471
rect -146 -1499 -118 -1471
rect -80 -1499 -52 -1471
rect -14 -1499 14 -1471
rect 52 -1499 80 -1471
rect 118 -1499 146 -1471
rect 184 -1499 212 -1471
rect 250 -1499 278 -1471
rect 316 -1499 344 -1471
rect 382 -1499 410 -1471
rect 448 -1499 476 -1471
rect 514 -1499 542 -1471
rect 580 -1499 608 -1471
rect 646 -1499 674 -1471
rect 712 -1499 740 -1471
rect -740 -1565 -712 -1537
rect -674 -1565 -646 -1537
rect -608 -1565 -580 -1537
rect -542 -1565 -514 -1537
rect -476 -1565 -448 -1537
rect -410 -1565 -382 -1537
rect -344 -1565 -316 -1537
rect -278 -1565 -250 -1537
rect -212 -1565 -184 -1537
rect -146 -1565 -118 -1537
rect -80 -1565 -52 -1537
rect -14 -1565 14 -1537
rect 52 -1565 80 -1537
rect 118 -1565 146 -1537
rect 184 -1565 212 -1537
rect 250 -1565 278 -1537
rect 316 -1565 344 -1537
rect 382 -1565 410 -1537
rect 448 -1565 476 -1537
rect 514 -1565 542 -1537
rect 580 -1565 608 -1537
rect 646 -1565 674 -1537
rect 712 -1565 740 -1537
rect -740 -1631 -712 -1603
rect -674 -1631 -646 -1603
rect -608 -1631 -580 -1603
rect -542 -1631 -514 -1603
rect -476 -1631 -448 -1603
rect -410 -1631 -382 -1603
rect -344 -1631 -316 -1603
rect -278 -1631 -250 -1603
rect -212 -1631 -184 -1603
rect -146 -1631 -118 -1603
rect -80 -1631 -52 -1603
rect -14 -1631 14 -1603
rect 52 -1631 80 -1603
rect 118 -1631 146 -1603
rect 184 -1631 212 -1603
rect 250 -1631 278 -1603
rect 316 -1631 344 -1603
rect 382 -1631 410 -1603
rect 448 -1631 476 -1603
rect 514 -1631 542 -1603
rect 580 -1631 608 -1603
rect 646 -1631 674 -1603
rect 712 -1631 740 -1603
rect -740 -1697 -712 -1669
rect -674 -1697 -646 -1669
rect -608 -1697 -580 -1669
rect -542 -1697 -514 -1669
rect -476 -1697 -448 -1669
rect -410 -1697 -382 -1669
rect -344 -1697 -316 -1669
rect -278 -1697 -250 -1669
rect -212 -1697 -184 -1669
rect -146 -1697 -118 -1669
rect -80 -1697 -52 -1669
rect -14 -1697 14 -1669
rect 52 -1697 80 -1669
rect 118 -1697 146 -1669
rect 184 -1697 212 -1669
rect 250 -1697 278 -1669
rect 316 -1697 344 -1669
rect 382 -1697 410 -1669
rect 448 -1697 476 -1669
rect 514 -1697 542 -1669
rect 580 -1697 608 -1669
rect 646 -1697 674 -1669
rect 712 -1697 740 -1669
rect -740 -1763 -712 -1735
rect -674 -1763 -646 -1735
rect -608 -1763 -580 -1735
rect -542 -1763 -514 -1735
rect -476 -1763 -448 -1735
rect -410 -1763 -382 -1735
rect -344 -1763 -316 -1735
rect -278 -1763 -250 -1735
rect -212 -1763 -184 -1735
rect -146 -1763 -118 -1735
rect -80 -1763 -52 -1735
rect -14 -1763 14 -1735
rect 52 -1763 80 -1735
rect 118 -1763 146 -1735
rect 184 -1763 212 -1735
rect 250 -1763 278 -1735
rect 316 -1763 344 -1735
rect 382 -1763 410 -1735
rect 448 -1763 476 -1735
rect 514 -1763 542 -1735
rect 580 -1763 608 -1735
rect 646 -1763 674 -1735
rect 712 -1763 740 -1735
rect -740 -1829 -712 -1801
rect -674 -1829 -646 -1801
rect -608 -1829 -580 -1801
rect -542 -1829 -514 -1801
rect -476 -1829 -448 -1801
rect -410 -1829 -382 -1801
rect -344 -1829 -316 -1801
rect -278 -1829 -250 -1801
rect -212 -1829 -184 -1801
rect -146 -1829 -118 -1801
rect -80 -1829 -52 -1801
rect -14 -1829 14 -1801
rect 52 -1829 80 -1801
rect 118 -1829 146 -1801
rect 184 -1829 212 -1801
rect 250 -1829 278 -1801
rect 316 -1829 344 -1801
rect 382 -1829 410 -1801
rect 448 -1829 476 -1801
rect 514 -1829 542 -1801
rect 580 -1829 608 -1801
rect 646 -1829 674 -1801
rect 712 -1829 740 -1801
rect -740 -1895 -712 -1867
rect -674 -1895 -646 -1867
rect -608 -1895 -580 -1867
rect -542 -1895 -514 -1867
rect -476 -1895 -448 -1867
rect -410 -1895 -382 -1867
rect -344 -1895 -316 -1867
rect -278 -1895 -250 -1867
rect -212 -1895 -184 -1867
rect -146 -1895 -118 -1867
rect -80 -1895 -52 -1867
rect -14 -1895 14 -1867
rect 52 -1895 80 -1867
rect 118 -1895 146 -1867
rect 184 -1895 212 -1867
rect 250 -1895 278 -1867
rect 316 -1895 344 -1867
rect 382 -1895 410 -1867
rect 448 -1895 476 -1867
rect 514 -1895 542 -1867
rect 580 -1895 608 -1867
rect 646 -1895 674 -1867
rect 712 -1895 740 -1867
rect -740 -1961 -712 -1933
rect -674 -1961 -646 -1933
rect -608 -1961 -580 -1933
rect -542 -1961 -514 -1933
rect -476 -1961 -448 -1933
rect -410 -1961 -382 -1933
rect -344 -1961 -316 -1933
rect -278 -1961 -250 -1933
rect -212 -1961 -184 -1933
rect -146 -1961 -118 -1933
rect -80 -1961 -52 -1933
rect -14 -1961 14 -1933
rect 52 -1961 80 -1933
rect 118 -1961 146 -1933
rect 184 -1961 212 -1933
rect 250 -1961 278 -1933
rect 316 -1961 344 -1933
rect 382 -1961 410 -1933
rect 448 -1961 476 -1933
rect 514 -1961 542 -1933
rect 580 -1961 608 -1933
rect 646 -1961 674 -1933
rect 712 -1961 740 -1933
rect -740 -2027 -712 -1999
rect -674 -2027 -646 -1999
rect -608 -2027 -580 -1999
rect -542 -2027 -514 -1999
rect -476 -2027 -448 -1999
rect -410 -2027 -382 -1999
rect -344 -2027 -316 -1999
rect -278 -2027 -250 -1999
rect -212 -2027 -184 -1999
rect -146 -2027 -118 -1999
rect -80 -2027 -52 -1999
rect -14 -2027 14 -1999
rect 52 -2027 80 -1999
rect 118 -2027 146 -1999
rect 184 -2027 212 -1999
rect 250 -2027 278 -1999
rect 316 -2027 344 -1999
rect 382 -2027 410 -1999
rect 448 -2027 476 -1999
rect 514 -2027 542 -1999
rect 580 -2027 608 -1999
rect 646 -2027 674 -1999
rect 712 -2027 740 -1999
rect -740 -2093 -712 -2065
rect -674 -2093 -646 -2065
rect -608 -2093 -580 -2065
rect -542 -2093 -514 -2065
rect -476 -2093 -448 -2065
rect -410 -2093 -382 -2065
rect -344 -2093 -316 -2065
rect -278 -2093 -250 -2065
rect -212 -2093 -184 -2065
rect -146 -2093 -118 -2065
rect -80 -2093 -52 -2065
rect -14 -2093 14 -2065
rect 52 -2093 80 -2065
rect 118 -2093 146 -2065
rect 184 -2093 212 -2065
rect 250 -2093 278 -2065
rect 316 -2093 344 -2065
rect 382 -2093 410 -2065
rect 448 -2093 476 -2065
rect 514 -2093 542 -2065
rect 580 -2093 608 -2065
rect 646 -2093 674 -2065
rect 712 -2093 740 -2065
rect -740 -2159 -712 -2131
rect -674 -2159 -646 -2131
rect -608 -2159 -580 -2131
rect -542 -2159 -514 -2131
rect -476 -2159 -448 -2131
rect -410 -2159 -382 -2131
rect -344 -2159 -316 -2131
rect -278 -2159 -250 -2131
rect -212 -2159 -184 -2131
rect -146 -2159 -118 -2131
rect -80 -2159 -52 -2131
rect -14 -2159 14 -2131
rect 52 -2159 80 -2131
rect 118 -2159 146 -2131
rect 184 -2159 212 -2131
rect 250 -2159 278 -2131
rect 316 -2159 344 -2131
rect 382 -2159 410 -2131
rect 448 -2159 476 -2131
rect 514 -2159 542 -2131
rect 580 -2159 608 -2131
rect 646 -2159 674 -2131
rect 712 -2159 740 -2131
rect -740 -2225 -712 -2197
rect -674 -2225 -646 -2197
rect -608 -2225 -580 -2197
rect -542 -2225 -514 -2197
rect -476 -2225 -448 -2197
rect -410 -2225 -382 -2197
rect -344 -2225 -316 -2197
rect -278 -2225 -250 -2197
rect -212 -2225 -184 -2197
rect -146 -2225 -118 -2197
rect -80 -2225 -52 -2197
rect -14 -2225 14 -2197
rect 52 -2225 80 -2197
rect 118 -2225 146 -2197
rect 184 -2225 212 -2197
rect 250 -2225 278 -2197
rect 316 -2225 344 -2197
rect 382 -2225 410 -2197
rect 448 -2225 476 -2197
rect 514 -2225 542 -2197
rect 580 -2225 608 -2197
rect 646 -2225 674 -2197
rect 712 -2225 740 -2197
rect -740 -2291 -712 -2263
rect -674 -2291 -646 -2263
rect -608 -2291 -580 -2263
rect -542 -2291 -514 -2263
rect -476 -2291 -448 -2263
rect -410 -2291 -382 -2263
rect -344 -2291 -316 -2263
rect -278 -2291 -250 -2263
rect -212 -2291 -184 -2263
rect -146 -2291 -118 -2263
rect -80 -2291 -52 -2263
rect -14 -2291 14 -2263
rect 52 -2291 80 -2263
rect 118 -2291 146 -2263
rect 184 -2291 212 -2263
rect 250 -2291 278 -2263
rect 316 -2291 344 -2263
rect 382 -2291 410 -2263
rect 448 -2291 476 -2263
rect 514 -2291 542 -2263
rect 580 -2291 608 -2263
rect 646 -2291 674 -2263
rect 712 -2291 740 -2263
rect -740 -2357 -712 -2329
rect -674 -2357 -646 -2329
rect -608 -2357 -580 -2329
rect -542 -2357 -514 -2329
rect -476 -2357 -448 -2329
rect -410 -2357 -382 -2329
rect -344 -2357 -316 -2329
rect -278 -2357 -250 -2329
rect -212 -2357 -184 -2329
rect -146 -2357 -118 -2329
rect -80 -2357 -52 -2329
rect -14 -2357 14 -2329
rect 52 -2357 80 -2329
rect 118 -2357 146 -2329
rect 184 -2357 212 -2329
rect 250 -2357 278 -2329
rect 316 -2357 344 -2329
rect 382 -2357 410 -2329
rect 448 -2357 476 -2329
rect 514 -2357 542 -2329
rect 580 -2357 608 -2329
rect 646 -2357 674 -2329
rect 712 -2357 740 -2329
rect -740 -2423 -712 -2395
rect -674 -2423 -646 -2395
rect -608 -2423 -580 -2395
rect -542 -2423 -514 -2395
rect -476 -2423 -448 -2395
rect -410 -2423 -382 -2395
rect -344 -2423 -316 -2395
rect -278 -2423 -250 -2395
rect -212 -2423 -184 -2395
rect -146 -2423 -118 -2395
rect -80 -2423 -52 -2395
rect -14 -2423 14 -2395
rect 52 -2423 80 -2395
rect 118 -2423 146 -2395
rect 184 -2423 212 -2395
rect 250 -2423 278 -2395
rect 316 -2423 344 -2395
rect 382 -2423 410 -2395
rect 448 -2423 476 -2395
rect 514 -2423 542 -2395
rect 580 -2423 608 -2395
rect 646 -2423 674 -2395
rect 712 -2423 740 -2395
rect -740 -2489 -712 -2461
rect -674 -2489 -646 -2461
rect -608 -2489 -580 -2461
rect -542 -2489 -514 -2461
rect -476 -2489 -448 -2461
rect -410 -2489 -382 -2461
rect -344 -2489 -316 -2461
rect -278 -2489 -250 -2461
rect -212 -2489 -184 -2461
rect -146 -2489 -118 -2461
rect -80 -2489 -52 -2461
rect -14 -2489 14 -2461
rect 52 -2489 80 -2461
rect 118 -2489 146 -2461
rect 184 -2489 212 -2461
rect 250 -2489 278 -2461
rect 316 -2489 344 -2461
rect 382 -2489 410 -2461
rect 448 -2489 476 -2461
rect 514 -2489 542 -2461
rect 580 -2489 608 -2461
rect 646 -2489 674 -2461
rect 712 -2489 740 -2461
rect -740 -2555 -712 -2527
rect -674 -2555 -646 -2527
rect -608 -2555 -580 -2527
rect -542 -2555 -514 -2527
rect -476 -2555 -448 -2527
rect -410 -2555 -382 -2527
rect -344 -2555 -316 -2527
rect -278 -2555 -250 -2527
rect -212 -2555 -184 -2527
rect -146 -2555 -118 -2527
rect -80 -2555 -52 -2527
rect -14 -2555 14 -2527
rect 52 -2555 80 -2527
rect 118 -2555 146 -2527
rect 184 -2555 212 -2527
rect 250 -2555 278 -2527
rect 316 -2555 344 -2527
rect 382 -2555 410 -2527
rect 448 -2555 476 -2527
rect 514 -2555 542 -2527
rect 580 -2555 608 -2527
rect 646 -2555 674 -2527
rect 712 -2555 740 -2527
rect -740 -2621 -712 -2593
rect -674 -2621 -646 -2593
rect -608 -2621 -580 -2593
rect -542 -2621 -514 -2593
rect -476 -2621 -448 -2593
rect -410 -2621 -382 -2593
rect -344 -2621 -316 -2593
rect -278 -2621 -250 -2593
rect -212 -2621 -184 -2593
rect -146 -2621 -118 -2593
rect -80 -2621 -52 -2593
rect -14 -2621 14 -2593
rect 52 -2621 80 -2593
rect 118 -2621 146 -2593
rect 184 -2621 212 -2593
rect 250 -2621 278 -2593
rect 316 -2621 344 -2593
rect 382 -2621 410 -2593
rect 448 -2621 476 -2593
rect 514 -2621 542 -2593
rect 580 -2621 608 -2593
rect 646 -2621 674 -2593
rect 712 -2621 740 -2593
rect -740 -2687 -712 -2659
rect -674 -2687 -646 -2659
rect -608 -2687 -580 -2659
rect -542 -2687 -514 -2659
rect -476 -2687 -448 -2659
rect -410 -2687 -382 -2659
rect -344 -2687 -316 -2659
rect -278 -2687 -250 -2659
rect -212 -2687 -184 -2659
rect -146 -2687 -118 -2659
rect -80 -2687 -52 -2659
rect -14 -2687 14 -2659
rect 52 -2687 80 -2659
rect 118 -2687 146 -2659
rect 184 -2687 212 -2659
rect 250 -2687 278 -2659
rect 316 -2687 344 -2659
rect 382 -2687 410 -2659
rect 448 -2687 476 -2659
rect 514 -2687 542 -2659
rect 580 -2687 608 -2659
rect 646 -2687 674 -2659
rect 712 -2687 740 -2659
rect -740 -2753 -712 -2725
rect -674 -2753 -646 -2725
rect -608 -2753 -580 -2725
rect -542 -2753 -514 -2725
rect -476 -2753 -448 -2725
rect -410 -2753 -382 -2725
rect -344 -2753 -316 -2725
rect -278 -2753 -250 -2725
rect -212 -2753 -184 -2725
rect -146 -2753 -118 -2725
rect -80 -2753 -52 -2725
rect -14 -2753 14 -2725
rect 52 -2753 80 -2725
rect 118 -2753 146 -2725
rect 184 -2753 212 -2725
rect 250 -2753 278 -2725
rect 316 -2753 344 -2725
rect 382 -2753 410 -2725
rect 448 -2753 476 -2725
rect 514 -2753 542 -2725
rect 580 -2753 608 -2725
rect 646 -2753 674 -2725
rect 712 -2753 740 -2725
rect -740 -2819 -712 -2791
rect -674 -2819 -646 -2791
rect -608 -2819 -580 -2791
rect -542 -2819 -514 -2791
rect -476 -2819 -448 -2791
rect -410 -2819 -382 -2791
rect -344 -2819 -316 -2791
rect -278 -2819 -250 -2791
rect -212 -2819 -184 -2791
rect -146 -2819 -118 -2791
rect -80 -2819 -52 -2791
rect -14 -2819 14 -2791
rect 52 -2819 80 -2791
rect 118 -2819 146 -2791
rect 184 -2819 212 -2791
rect 250 -2819 278 -2791
rect 316 -2819 344 -2791
rect 382 -2819 410 -2791
rect 448 -2819 476 -2791
rect 514 -2819 542 -2791
rect 580 -2819 608 -2791
rect 646 -2819 674 -2791
rect 712 -2819 740 -2791
rect -740 -2885 -712 -2857
rect -674 -2885 -646 -2857
rect -608 -2885 -580 -2857
rect -542 -2885 -514 -2857
rect -476 -2885 -448 -2857
rect -410 -2885 -382 -2857
rect -344 -2885 -316 -2857
rect -278 -2885 -250 -2857
rect -212 -2885 -184 -2857
rect -146 -2885 -118 -2857
rect -80 -2885 -52 -2857
rect -14 -2885 14 -2857
rect 52 -2885 80 -2857
rect 118 -2885 146 -2857
rect 184 -2885 212 -2857
rect 250 -2885 278 -2857
rect 316 -2885 344 -2857
rect 382 -2885 410 -2857
rect 448 -2885 476 -2857
rect 514 -2885 542 -2857
rect 580 -2885 608 -2857
rect 646 -2885 674 -2857
rect 712 -2885 740 -2857
rect -740 -2951 -712 -2923
rect -674 -2951 -646 -2923
rect -608 -2951 -580 -2923
rect -542 -2951 -514 -2923
rect -476 -2951 -448 -2923
rect -410 -2951 -382 -2923
rect -344 -2951 -316 -2923
rect -278 -2951 -250 -2923
rect -212 -2951 -184 -2923
rect -146 -2951 -118 -2923
rect -80 -2951 -52 -2923
rect -14 -2951 14 -2923
rect 52 -2951 80 -2923
rect 118 -2951 146 -2923
rect 184 -2951 212 -2923
rect 250 -2951 278 -2923
rect 316 -2951 344 -2923
rect 382 -2951 410 -2923
rect 448 -2951 476 -2923
rect 514 -2951 542 -2923
rect 580 -2951 608 -2923
rect 646 -2951 674 -2923
rect 712 -2951 740 -2923
rect -740 -3017 -712 -2989
rect -674 -3017 -646 -2989
rect -608 -3017 -580 -2989
rect -542 -3017 -514 -2989
rect -476 -3017 -448 -2989
rect -410 -3017 -382 -2989
rect -344 -3017 -316 -2989
rect -278 -3017 -250 -2989
rect -212 -3017 -184 -2989
rect -146 -3017 -118 -2989
rect -80 -3017 -52 -2989
rect -14 -3017 14 -2989
rect 52 -3017 80 -2989
rect 118 -3017 146 -2989
rect 184 -3017 212 -2989
rect 250 -3017 278 -2989
rect 316 -3017 344 -2989
rect 382 -3017 410 -2989
rect 448 -3017 476 -2989
rect 514 -3017 542 -2989
rect 580 -3017 608 -2989
rect 646 -3017 674 -2989
rect 712 -3017 740 -2989
rect -740 -3083 -712 -3055
rect -674 -3083 -646 -3055
rect -608 -3083 -580 -3055
rect -542 -3083 -514 -3055
rect -476 -3083 -448 -3055
rect -410 -3083 -382 -3055
rect -344 -3083 -316 -3055
rect -278 -3083 -250 -3055
rect -212 -3083 -184 -3055
rect -146 -3083 -118 -3055
rect -80 -3083 -52 -3055
rect -14 -3083 14 -3055
rect 52 -3083 80 -3055
rect 118 -3083 146 -3055
rect 184 -3083 212 -3055
rect 250 -3083 278 -3055
rect 316 -3083 344 -3055
rect 382 -3083 410 -3055
rect 448 -3083 476 -3055
rect 514 -3083 542 -3055
rect 580 -3083 608 -3055
rect 646 -3083 674 -3055
rect 712 -3083 740 -3055
rect -740 -3149 -712 -3121
rect -674 -3149 -646 -3121
rect -608 -3149 -580 -3121
rect -542 -3149 -514 -3121
rect -476 -3149 -448 -3121
rect -410 -3149 -382 -3121
rect -344 -3149 -316 -3121
rect -278 -3149 -250 -3121
rect -212 -3149 -184 -3121
rect -146 -3149 -118 -3121
rect -80 -3149 -52 -3121
rect -14 -3149 14 -3121
rect 52 -3149 80 -3121
rect 118 -3149 146 -3121
rect 184 -3149 212 -3121
rect 250 -3149 278 -3121
rect 316 -3149 344 -3121
rect 382 -3149 410 -3121
rect 448 -3149 476 -3121
rect 514 -3149 542 -3121
rect 580 -3149 608 -3121
rect 646 -3149 674 -3121
rect 712 -3149 740 -3121
rect -740 -3215 -712 -3187
rect -674 -3215 -646 -3187
rect -608 -3215 -580 -3187
rect -542 -3215 -514 -3187
rect -476 -3215 -448 -3187
rect -410 -3215 -382 -3187
rect -344 -3215 -316 -3187
rect -278 -3215 -250 -3187
rect -212 -3215 -184 -3187
rect -146 -3215 -118 -3187
rect -80 -3215 -52 -3187
rect -14 -3215 14 -3187
rect 52 -3215 80 -3187
rect 118 -3215 146 -3187
rect 184 -3215 212 -3187
rect 250 -3215 278 -3187
rect 316 -3215 344 -3187
rect 382 -3215 410 -3187
rect 448 -3215 476 -3187
rect 514 -3215 542 -3187
rect 580 -3215 608 -3187
rect 646 -3215 674 -3187
rect 712 -3215 740 -3187
rect -740 -3281 -712 -3253
rect -674 -3281 -646 -3253
rect -608 -3281 -580 -3253
rect -542 -3281 -514 -3253
rect -476 -3281 -448 -3253
rect -410 -3281 -382 -3253
rect -344 -3281 -316 -3253
rect -278 -3281 -250 -3253
rect -212 -3281 -184 -3253
rect -146 -3281 -118 -3253
rect -80 -3281 -52 -3253
rect -14 -3281 14 -3253
rect 52 -3281 80 -3253
rect 118 -3281 146 -3253
rect 184 -3281 212 -3253
rect 250 -3281 278 -3253
rect 316 -3281 344 -3253
rect 382 -3281 410 -3253
rect 448 -3281 476 -3253
rect 514 -3281 542 -3253
rect 580 -3281 608 -3253
rect 646 -3281 674 -3253
rect 712 -3281 740 -3253
rect -740 -3347 -712 -3319
rect -674 -3347 -646 -3319
rect -608 -3347 -580 -3319
rect -542 -3347 -514 -3319
rect -476 -3347 -448 -3319
rect -410 -3347 -382 -3319
rect -344 -3347 -316 -3319
rect -278 -3347 -250 -3319
rect -212 -3347 -184 -3319
rect -146 -3347 -118 -3319
rect -80 -3347 -52 -3319
rect -14 -3347 14 -3319
rect 52 -3347 80 -3319
rect 118 -3347 146 -3319
rect 184 -3347 212 -3319
rect 250 -3347 278 -3319
rect 316 -3347 344 -3319
rect 382 -3347 410 -3319
rect 448 -3347 476 -3319
rect 514 -3347 542 -3319
rect 580 -3347 608 -3319
rect 646 -3347 674 -3319
rect 712 -3347 740 -3319
rect -740 -3413 -712 -3385
rect -674 -3413 -646 -3385
rect -608 -3413 -580 -3385
rect -542 -3413 -514 -3385
rect -476 -3413 -448 -3385
rect -410 -3413 -382 -3385
rect -344 -3413 -316 -3385
rect -278 -3413 -250 -3385
rect -212 -3413 -184 -3385
rect -146 -3413 -118 -3385
rect -80 -3413 -52 -3385
rect -14 -3413 14 -3385
rect 52 -3413 80 -3385
rect 118 -3413 146 -3385
rect 184 -3413 212 -3385
rect 250 -3413 278 -3385
rect 316 -3413 344 -3385
rect 382 -3413 410 -3385
rect 448 -3413 476 -3385
rect 514 -3413 542 -3385
rect 580 -3413 608 -3385
rect 646 -3413 674 -3385
rect 712 -3413 740 -3385
rect -740 -3479 -712 -3451
rect -674 -3479 -646 -3451
rect -608 -3479 -580 -3451
rect -542 -3479 -514 -3451
rect -476 -3479 -448 -3451
rect -410 -3479 -382 -3451
rect -344 -3479 -316 -3451
rect -278 -3479 -250 -3451
rect -212 -3479 -184 -3451
rect -146 -3479 -118 -3451
rect -80 -3479 -52 -3451
rect -14 -3479 14 -3451
rect 52 -3479 80 -3451
rect 118 -3479 146 -3451
rect 184 -3479 212 -3451
rect 250 -3479 278 -3451
rect 316 -3479 344 -3451
rect 382 -3479 410 -3451
rect 448 -3479 476 -3451
rect 514 -3479 542 -3451
rect 580 -3479 608 -3451
rect 646 -3479 674 -3451
rect 712 -3479 740 -3451
rect -740 -3545 -712 -3517
rect -674 -3545 -646 -3517
rect -608 -3545 -580 -3517
rect -542 -3545 -514 -3517
rect -476 -3545 -448 -3517
rect -410 -3545 -382 -3517
rect -344 -3545 -316 -3517
rect -278 -3545 -250 -3517
rect -212 -3545 -184 -3517
rect -146 -3545 -118 -3517
rect -80 -3545 -52 -3517
rect -14 -3545 14 -3517
rect 52 -3545 80 -3517
rect 118 -3545 146 -3517
rect 184 -3545 212 -3517
rect 250 -3545 278 -3517
rect 316 -3545 344 -3517
rect 382 -3545 410 -3517
rect 448 -3545 476 -3517
rect 514 -3545 542 -3517
rect 580 -3545 608 -3517
rect 646 -3545 674 -3517
rect 712 -3545 740 -3517
rect -740 -3611 -712 -3583
rect -674 -3611 -646 -3583
rect -608 -3611 -580 -3583
rect -542 -3611 -514 -3583
rect -476 -3611 -448 -3583
rect -410 -3611 -382 -3583
rect -344 -3611 -316 -3583
rect -278 -3611 -250 -3583
rect -212 -3611 -184 -3583
rect -146 -3611 -118 -3583
rect -80 -3611 -52 -3583
rect -14 -3611 14 -3583
rect 52 -3611 80 -3583
rect 118 -3611 146 -3583
rect 184 -3611 212 -3583
rect 250 -3611 278 -3583
rect 316 -3611 344 -3583
rect 382 -3611 410 -3583
rect 448 -3611 476 -3583
rect 514 -3611 542 -3583
rect 580 -3611 608 -3583
rect 646 -3611 674 -3583
rect 712 -3611 740 -3583
rect -740 -3677 -712 -3649
rect -674 -3677 -646 -3649
rect -608 -3677 -580 -3649
rect -542 -3677 -514 -3649
rect -476 -3677 -448 -3649
rect -410 -3677 -382 -3649
rect -344 -3677 -316 -3649
rect -278 -3677 -250 -3649
rect -212 -3677 -184 -3649
rect -146 -3677 -118 -3649
rect -80 -3677 -52 -3649
rect -14 -3677 14 -3649
rect 52 -3677 80 -3649
rect 118 -3677 146 -3649
rect 184 -3677 212 -3649
rect 250 -3677 278 -3649
rect 316 -3677 344 -3649
rect 382 -3677 410 -3649
rect 448 -3677 476 -3649
rect 514 -3677 542 -3649
rect 580 -3677 608 -3649
rect 646 -3677 674 -3649
rect 712 -3677 740 -3649
rect -740 -3743 -712 -3715
rect -674 -3743 -646 -3715
rect -608 -3743 -580 -3715
rect -542 -3743 -514 -3715
rect -476 -3743 -448 -3715
rect -410 -3743 -382 -3715
rect -344 -3743 -316 -3715
rect -278 -3743 -250 -3715
rect -212 -3743 -184 -3715
rect -146 -3743 -118 -3715
rect -80 -3743 -52 -3715
rect -14 -3743 14 -3715
rect 52 -3743 80 -3715
rect 118 -3743 146 -3715
rect 184 -3743 212 -3715
rect 250 -3743 278 -3715
rect 316 -3743 344 -3715
rect 382 -3743 410 -3715
rect 448 -3743 476 -3715
rect 514 -3743 542 -3715
rect 580 -3743 608 -3715
rect 646 -3743 674 -3715
rect 712 -3743 740 -3715
rect -740 -3809 -712 -3781
rect -674 -3809 -646 -3781
rect -608 -3809 -580 -3781
rect -542 -3809 -514 -3781
rect -476 -3809 -448 -3781
rect -410 -3809 -382 -3781
rect -344 -3809 -316 -3781
rect -278 -3809 -250 -3781
rect -212 -3809 -184 -3781
rect -146 -3809 -118 -3781
rect -80 -3809 -52 -3781
rect -14 -3809 14 -3781
rect 52 -3809 80 -3781
rect 118 -3809 146 -3781
rect 184 -3809 212 -3781
rect 250 -3809 278 -3781
rect 316 -3809 344 -3781
rect 382 -3809 410 -3781
rect 448 -3809 476 -3781
rect 514 -3809 542 -3781
rect 580 -3809 608 -3781
rect 646 -3809 674 -3781
rect 712 -3809 740 -3781
rect -740 -3875 -712 -3847
rect -674 -3875 -646 -3847
rect -608 -3875 -580 -3847
rect -542 -3875 -514 -3847
rect -476 -3875 -448 -3847
rect -410 -3875 -382 -3847
rect -344 -3875 -316 -3847
rect -278 -3875 -250 -3847
rect -212 -3875 -184 -3847
rect -146 -3875 -118 -3847
rect -80 -3875 -52 -3847
rect -14 -3875 14 -3847
rect 52 -3875 80 -3847
rect 118 -3875 146 -3847
rect 184 -3875 212 -3847
rect 250 -3875 278 -3847
rect 316 -3875 344 -3847
rect 382 -3875 410 -3847
rect 448 -3875 476 -3847
rect 514 -3875 542 -3847
rect 580 -3875 608 -3847
rect 646 -3875 674 -3847
rect 712 -3875 740 -3847
<< metal4 >>
rect -745 3875 745 3880
rect -745 3847 -740 3875
rect -712 3847 -674 3875
rect -646 3847 -608 3875
rect -580 3847 -542 3875
rect -514 3847 -476 3875
rect -448 3847 -410 3875
rect -382 3847 -344 3875
rect -316 3847 -278 3875
rect -250 3847 -212 3875
rect -184 3847 -146 3875
rect -118 3847 -80 3875
rect -52 3847 -14 3875
rect 14 3847 52 3875
rect 80 3847 118 3875
rect 146 3847 184 3875
rect 212 3847 250 3875
rect 278 3847 316 3875
rect 344 3847 382 3875
rect 410 3847 448 3875
rect 476 3847 514 3875
rect 542 3847 580 3875
rect 608 3847 646 3875
rect 674 3847 712 3875
rect 740 3847 745 3875
rect -745 3809 745 3847
rect -745 3781 -740 3809
rect -712 3781 -674 3809
rect -646 3781 -608 3809
rect -580 3781 -542 3809
rect -514 3781 -476 3809
rect -448 3781 -410 3809
rect -382 3781 -344 3809
rect -316 3781 -278 3809
rect -250 3781 -212 3809
rect -184 3781 -146 3809
rect -118 3781 -80 3809
rect -52 3781 -14 3809
rect 14 3781 52 3809
rect 80 3781 118 3809
rect 146 3781 184 3809
rect 212 3781 250 3809
rect 278 3781 316 3809
rect 344 3781 382 3809
rect 410 3781 448 3809
rect 476 3781 514 3809
rect 542 3781 580 3809
rect 608 3781 646 3809
rect 674 3781 712 3809
rect 740 3781 745 3809
rect -745 3743 745 3781
rect -745 3715 -740 3743
rect -712 3715 -674 3743
rect -646 3715 -608 3743
rect -580 3715 -542 3743
rect -514 3715 -476 3743
rect -448 3715 -410 3743
rect -382 3715 -344 3743
rect -316 3715 -278 3743
rect -250 3715 -212 3743
rect -184 3715 -146 3743
rect -118 3715 -80 3743
rect -52 3715 -14 3743
rect 14 3715 52 3743
rect 80 3715 118 3743
rect 146 3715 184 3743
rect 212 3715 250 3743
rect 278 3715 316 3743
rect 344 3715 382 3743
rect 410 3715 448 3743
rect 476 3715 514 3743
rect 542 3715 580 3743
rect 608 3715 646 3743
rect 674 3715 712 3743
rect 740 3715 745 3743
rect -745 3677 745 3715
rect -745 3649 -740 3677
rect -712 3649 -674 3677
rect -646 3649 -608 3677
rect -580 3649 -542 3677
rect -514 3649 -476 3677
rect -448 3649 -410 3677
rect -382 3649 -344 3677
rect -316 3649 -278 3677
rect -250 3649 -212 3677
rect -184 3649 -146 3677
rect -118 3649 -80 3677
rect -52 3649 -14 3677
rect 14 3649 52 3677
rect 80 3649 118 3677
rect 146 3649 184 3677
rect 212 3649 250 3677
rect 278 3649 316 3677
rect 344 3649 382 3677
rect 410 3649 448 3677
rect 476 3649 514 3677
rect 542 3649 580 3677
rect 608 3649 646 3677
rect 674 3649 712 3677
rect 740 3649 745 3677
rect -745 3611 745 3649
rect -745 3583 -740 3611
rect -712 3583 -674 3611
rect -646 3583 -608 3611
rect -580 3583 -542 3611
rect -514 3583 -476 3611
rect -448 3583 -410 3611
rect -382 3583 -344 3611
rect -316 3583 -278 3611
rect -250 3583 -212 3611
rect -184 3583 -146 3611
rect -118 3583 -80 3611
rect -52 3583 -14 3611
rect 14 3583 52 3611
rect 80 3583 118 3611
rect 146 3583 184 3611
rect 212 3583 250 3611
rect 278 3583 316 3611
rect 344 3583 382 3611
rect 410 3583 448 3611
rect 476 3583 514 3611
rect 542 3583 580 3611
rect 608 3583 646 3611
rect 674 3583 712 3611
rect 740 3583 745 3611
rect -745 3545 745 3583
rect -745 3517 -740 3545
rect -712 3517 -674 3545
rect -646 3517 -608 3545
rect -580 3517 -542 3545
rect -514 3517 -476 3545
rect -448 3517 -410 3545
rect -382 3517 -344 3545
rect -316 3517 -278 3545
rect -250 3517 -212 3545
rect -184 3517 -146 3545
rect -118 3517 -80 3545
rect -52 3517 -14 3545
rect 14 3517 52 3545
rect 80 3517 118 3545
rect 146 3517 184 3545
rect 212 3517 250 3545
rect 278 3517 316 3545
rect 344 3517 382 3545
rect 410 3517 448 3545
rect 476 3517 514 3545
rect 542 3517 580 3545
rect 608 3517 646 3545
rect 674 3517 712 3545
rect 740 3517 745 3545
rect -745 3479 745 3517
rect -745 3451 -740 3479
rect -712 3451 -674 3479
rect -646 3451 -608 3479
rect -580 3451 -542 3479
rect -514 3451 -476 3479
rect -448 3451 -410 3479
rect -382 3451 -344 3479
rect -316 3451 -278 3479
rect -250 3451 -212 3479
rect -184 3451 -146 3479
rect -118 3451 -80 3479
rect -52 3451 -14 3479
rect 14 3451 52 3479
rect 80 3451 118 3479
rect 146 3451 184 3479
rect 212 3451 250 3479
rect 278 3451 316 3479
rect 344 3451 382 3479
rect 410 3451 448 3479
rect 476 3451 514 3479
rect 542 3451 580 3479
rect 608 3451 646 3479
rect 674 3451 712 3479
rect 740 3451 745 3479
rect -745 3413 745 3451
rect -745 3385 -740 3413
rect -712 3385 -674 3413
rect -646 3385 -608 3413
rect -580 3385 -542 3413
rect -514 3385 -476 3413
rect -448 3385 -410 3413
rect -382 3385 -344 3413
rect -316 3385 -278 3413
rect -250 3385 -212 3413
rect -184 3385 -146 3413
rect -118 3385 -80 3413
rect -52 3385 -14 3413
rect 14 3385 52 3413
rect 80 3385 118 3413
rect 146 3385 184 3413
rect 212 3385 250 3413
rect 278 3385 316 3413
rect 344 3385 382 3413
rect 410 3385 448 3413
rect 476 3385 514 3413
rect 542 3385 580 3413
rect 608 3385 646 3413
rect 674 3385 712 3413
rect 740 3385 745 3413
rect -745 3347 745 3385
rect -745 3319 -740 3347
rect -712 3319 -674 3347
rect -646 3319 -608 3347
rect -580 3319 -542 3347
rect -514 3319 -476 3347
rect -448 3319 -410 3347
rect -382 3319 -344 3347
rect -316 3319 -278 3347
rect -250 3319 -212 3347
rect -184 3319 -146 3347
rect -118 3319 -80 3347
rect -52 3319 -14 3347
rect 14 3319 52 3347
rect 80 3319 118 3347
rect 146 3319 184 3347
rect 212 3319 250 3347
rect 278 3319 316 3347
rect 344 3319 382 3347
rect 410 3319 448 3347
rect 476 3319 514 3347
rect 542 3319 580 3347
rect 608 3319 646 3347
rect 674 3319 712 3347
rect 740 3319 745 3347
rect -745 3281 745 3319
rect -745 3253 -740 3281
rect -712 3253 -674 3281
rect -646 3253 -608 3281
rect -580 3253 -542 3281
rect -514 3253 -476 3281
rect -448 3253 -410 3281
rect -382 3253 -344 3281
rect -316 3253 -278 3281
rect -250 3253 -212 3281
rect -184 3253 -146 3281
rect -118 3253 -80 3281
rect -52 3253 -14 3281
rect 14 3253 52 3281
rect 80 3253 118 3281
rect 146 3253 184 3281
rect 212 3253 250 3281
rect 278 3253 316 3281
rect 344 3253 382 3281
rect 410 3253 448 3281
rect 476 3253 514 3281
rect 542 3253 580 3281
rect 608 3253 646 3281
rect 674 3253 712 3281
rect 740 3253 745 3281
rect -745 3215 745 3253
rect -745 3187 -740 3215
rect -712 3187 -674 3215
rect -646 3187 -608 3215
rect -580 3187 -542 3215
rect -514 3187 -476 3215
rect -448 3187 -410 3215
rect -382 3187 -344 3215
rect -316 3187 -278 3215
rect -250 3187 -212 3215
rect -184 3187 -146 3215
rect -118 3187 -80 3215
rect -52 3187 -14 3215
rect 14 3187 52 3215
rect 80 3187 118 3215
rect 146 3187 184 3215
rect 212 3187 250 3215
rect 278 3187 316 3215
rect 344 3187 382 3215
rect 410 3187 448 3215
rect 476 3187 514 3215
rect 542 3187 580 3215
rect 608 3187 646 3215
rect 674 3187 712 3215
rect 740 3187 745 3215
rect -745 3149 745 3187
rect -745 3121 -740 3149
rect -712 3121 -674 3149
rect -646 3121 -608 3149
rect -580 3121 -542 3149
rect -514 3121 -476 3149
rect -448 3121 -410 3149
rect -382 3121 -344 3149
rect -316 3121 -278 3149
rect -250 3121 -212 3149
rect -184 3121 -146 3149
rect -118 3121 -80 3149
rect -52 3121 -14 3149
rect 14 3121 52 3149
rect 80 3121 118 3149
rect 146 3121 184 3149
rect 212 3121 250 3149
rect 278 3121 316 3149
rect 344 3121 382 3149
rect 410 3121 448 3149
rect 476 3121 514 3149
rect 542 3121 580 3149
rect 608 3121 646 3149
rect 674 3121 712 3149
rect 740 3121 745 3149
rect -745 3083 745 3121
rect -745 3055 -740 3083
rect -712 3055 -674 3083
rect -646 3055 -608 3083
rect -580 3055 -542 3083
rect -514 3055 -476 3083
rect -448 3055 -410 3083
rect -382 3055 -344 3083
rect -316 3055 -278 3083
rect -250 3055 -212 3083
rect -184 3055 -146 3083
rect -118 3055 -80 3083
rect -52 3055 -14 3083
rect 14 3055 52 3083
rect 80 3055 118 3083
rect 146 3055 184 3083
rect 212 3055 250 3083
rect 278 3055 316 3083
rect 344 3055 382 3083
rect 410 3055 448 3083
rect 476 3055 514 3083
rect 542 3055 580 3083
rect 608 3055 646 3083
rect 674 3055 712 3083
rect 740 3055 745 3083
rect -745 3017 745 3055
rect -745 2989 -740 3017
rect -712 2989 -674 3017
rect -646 2989 -608 3017
rect -580 2989 -542 3017
rect -514 2989 -476 3017
rect -448 2989 -410 3017
rect -382 2989 -344 3017
rect -316 2989 -278 3017
rect -250 2989 -212 3017
rect -184 2989 -146 3017
rect -118 2989 -80 3017
rect -52 2989 -14 3017
rect 14 2989 52 3017
rect 80 2989 118 3017
rect 146 2989 184 3017
rect 212 2989 250 3017
rect 278 2989 316 3017
rect 344 2989 382 3017
rect 410 2989 448 3017
rect 476 2989 514 3017
rect 542 2989 580 3017
rect 608 2989 646 3017
rect 674 2989 712 3017
rect 740 2989 745 3017
rect -745 2951 745 2989
rect -745 2923 -740 2951
rect -712 2923 -674 2951
rect -646 2923 -608 2951
rect -580 2923 -542 2951
rect -514 2923 -476 2951
rect -448 2923 -410 2951
rect -382 2923 -344 2951
rect -316 2923 -278 2951
rect -250 2923 -212 2951
rect -184 2923 -146 2951
rect -118 2923 -80 2951
rect -52 2923 -14 2951
rect 14 2923 52 2951
rect 80 2923 118 2951
rect 146 2923 184 2951
rect 212 2923 250 2951
rect 278 2923 316 2951
rect 344 2923 382 2951
rect 410 2923 448 2951
rect 476 2923 514 2951
rect 542 2923 580 2951
rect 608 2923 646 2951
rect 674 2923 712 2951
rect 740 2923 745 2951
rect -745 2885 745 2923
rect -745 2857 -740 2885
rect -712 2857 -674 2885
rect -646 2857 -608 2885
rect -580 2857 -542 2885
rect -514 2857 -476 2885
rect -448 2857 -410 2885
rect -382 2857 -344 2885
rect -316 2857 -278 2885
rect -250 2857 -212 2885
rect -184 2857 -146 2885
rect -118 2857 -80 2885
rect -52 2857 -14 2885
rect 14 2857 52 2885
rect 80 2857 118 2885
rect 146 2857 184 2885
rect 212 2857 250 2885
rect 278 2857 316 2885
rect 344 2857 382 2885
rect 410 2857 448 2885
rect 476 2857 514 2885
rect 542 2857 580 2885
rect 608 2857 646 2885
rect 674 2857 712 2885
rect 740 2857 745 2885
rect -745 2819 745 2857
rect -745 2791 -740 2819
rect -712 2791 -674 2819
rect -646 2791 -608 2819
rect -580 2791 -542 2819
rect -514 2791 -476 2819
rect -448 2791 -410 2819
rect -382 2791 -344 2819
rect -316 2791 -278 2819
rect -250 2791 -212 2819
rect -184 2791 -146 2819
rect -118 2791 -80 2819
rect -52 2791 -14 2819
rect 14 2791 52 2819
rect 80 2791 118 2819
rect 146 2791 184 2819
rect 212 2791 250 2819
rect 278 2791 316 2819
rect 344 2791 382 2819
rect 410 2791 448 2819
rect 476 2791 514 2819
rect 542 2791 580 2819
rect 608 2791 646 2819
rect 674 2791 712 2819
rect 740 2791 745 2819
rect -745 2753 745 2791
rect -745 2725 -740 2753
rect -712 2725 -674 2753
rect -646 2725 -608 2753
rect -580 2725 -542 2753
rect -514 2725 -476 2753
rect -448 2725 -410 2753
rect -382 2725 -344 2753
rect -316 2725 -278 2753
rect -250 2725 -212 2753
rect -184 2725 -146 2753
rect -118 2725 -80 2753
rect -52 2725 -14 2753
rect 14 2725 52 2753
rect 80 2725 118 2753
rect 146 2725 184 2753
rect 212 2725 250 2753
rect 278 2725 316 2753
rect 344 2725 382 2753
rect 410 2725 448 2753
rect 476 2725 514 2753
rect 542 2725 580 2753
rect 608 2725 646 2753
rect 674 2725 712 2753
rect 740 2725 745 2753
rect -745 2687 745 2725
rect -745 2659 -740 2687
rect -712 2659 -674 2687
rect -646 2659 -608 2687
rect -580 2659 -542 2687
rect -514 2659 -476 2687
rect -448 2659 -410 2687
rect -382 2659 -344 2687
rect -316 2659 -278 2687
rect -250 2659 -212 2687
rect -184 2659 -146 2687
rect -118 2659 -80 2687
rect -52 2659 -14 2687
rect 14 2659 52 2687
rect 80 2659 118 2687
rect 146 2659 184 2687
rect 212 2659 250 2687
rect 278 2659 316 2687
rect 344 2659 382 2687
rect 410 2659 448 2687
rect 476 2659 514 2687
rect 542 2659 580 2687
rect 608 2659 646 2687
rect 674 2659 712 2687
rect 740 2659 745 2687
rect -745 2621 745 2659
rect -745 2593 -740 2621
rect -712 2593 -674 2621
rect -646 2593 -608 2621
rect -580 2593 -542 2621
rect -514 2593 -476 2621
rect -448 2593 -410 2621
rect -382 2593 -344 2621
rect -316 2593 -278 2621
rect -250 2593 -212 2621
rect -184 2593 -146 2621
rect -118 2593 -80 2621
rect -52 2593 -14 2621
rect 14 2593 52 2621
rect 80 2593 118 2621
rect 146 2593 184 2621
rect 212 2593 250 2621
rect 278 2593 316 2621
rect 344 2593 382 2621
rect 410 2593 448 2621
rect 476 2593 514 2621
rect 542 2593 580 2621
rect 608 2593 646 2621
rect 674 2593 712 2621
rect 740 2593 745 2621
rect -745 2555 745 2593
rect -745 2527 -740 2555
rect -712 2527 -674 2555
rect -646 2527 -608 2555
rect -580 2527 -542 2555
rect -514 2527 -476 2555
rect -448 2527 -410 2555
rect -382 2527 -344 2555
rect -316 2527 -278 2555
rect -250 2527 -212 2555
rect -184 2527 -146 2555
rect -118 2527 -80 2555
rect -52 2527 -14 2555
rect 14 2527 52 2555
rect 80 2527 118 2555
rect 146 2527 184 2555
rect 212 2527 250 2555
rect 278 2527 316 2555
rect 344 2527 382 2555
rect 410 2527 448 2555
rect 476 2527 514 2555
rect 542 2527 580 2555
rect 608 2527 646 2555
rect 674 2527 712 2555
rect 740 2527 745 2555
rect -745 2489 745 2527
rect -745 2461 -740 2489
rect -712 2461 -674 2489
rect -646 2461 -608 2489
rect -580 2461 -542 2489
rect -514 2461 -476 2489
rect -448 2461 -410 2489
rect -382 2461 -344 2489
rect -316 2461 -278 2489
rect -250 2461 -212 2489
rect -184 2461 -146 2489
rect -118 2461 -80 2489
rect -52 2461 -14 2489
rect 14 2461 52 2489
rect 80 2461 118 2489
rect 146 2461 184 2489
rect 212 2461 250 2489
rect 278 2461 316 2489
rect 344 2461 382 2489
rect 410 2461 448 2489
rect 476 2461 514 2489
rect 542 2461 580 2489
rect 608 2461 646 2489
rect 674 2461 712 2489
rect 740 2461 745 2489
rect -745 2423 745 2461
rect -745 2395 -740 2423
rect -712 2395 -674 2423
rect -646 2395 -608 2423
rect -580 2395 -542 2423
rect -514 2395 -476 2423
rect -448 2395 -410 2423
rect -382 2395 -344 2423
rect -316 2395 -278 2423
rect -250 2395 -212 2423
rect -184 2395 -146 2423
rect -118 2395 -80 2423
rect -52 2395 -14 2423
rect 14 2395 52 2423
rect 80 2395 118 2423
rect 146 2395 184 2423
rect 212 2395 250 2423
rect 278 2395 316 2423
rect 344 2395 382 2423
rect 410 2395 448 2423
rect 476 2395 514 2423
rect 542 2395 580 2423
rect 608 2395 646 2423
rect 674 2395 712 2423
rect 740 2395 745 2423
rect -745 2357 745 2395
rect -745 2329 -740 2357
rect -712 2329 -674 2357
rect -646 2329 -608 2357
rect -580 2329 -542 2357
rect -514 2329 -476 2357
rect -448 2329 -410 2357
rect -382 2329 -344 2357
rect -316 2329 -278 2357
rect -250 2329 -212 2357
rect -184 2329 -146 2357
rect -118 2329 -80 2357
rect -52 2329 -14 2357
rect 14 2329 52 2357
rect 80 2329 118 2357
rect 146 2329 184 2357
rect 212 2329 250 2357
rect 278 2329 316 2357
rect 344 2329 382 2357
rect 410 2329 448 2357
rect 476 2329 514 2357
rect 542 2329 580 2357
rect 608 2329 646 2357
rect 674 2329 712 2357
rect 740 2329 745 2357
rect -745 2291 745 2329
rect -745 2263 -740 2291
rect -712 2263 -674 2291
rect -646 2263 -608 2291
rect -580 2263 -542 2291
rect -514 2263 -476 2291
rect -448 2263 -410 2291
rect -382 2263 -344 2291
rect -316 2263 -278 2291
rect -250 2263 -212 2291
rect -184 2263 -146 2291
rect -118 2263 -80 2291
rect -52 2263 -14 2291
rect 14 2263 52 2291
rect 80 2263 118 2291
rect 146 2263 184 2291
rect 212 2263 250 2291
rect 278 2263 316 2291
rect 344 2263 382 2291
rect 410 2263 448 2291
rect 476 2263 514 2291
rect 542 2263 580 2291
rect 608 2263 646 2291
rect 674 2263 712 2291
rect 740 2263 745 2291
rect -745 2225 745 2263
rect -745 2197 -740 2225
rect -712 2197 -674 2225
rect -646 2197 -608 2225
rect -580 2197 -542 2225
rect -514 2197 -476 2225
rect -448 2197 -410 2225
rect -382 2197 -344 2225
rect -316 2197 -278 2225
rect -250 2197 -212 2225
rect -184 2197 -146 2225
rect -118 2197 -80 2225
rect -52 2197 -14 2225
rect 14 2197 52 2225
rect 80 2197 118 2225
rect 146 2197 184 2225
rect 212 2197 250 2225
rect 278 2197 316 2225
rect 344 2197 382 2225
rect 410 2197 448 2225
rect 476 2197 514 2225
rect 542 2197 580 2225
rect 608 2197 646 2225
rect 674 2197 712 2225
rect 740 2197 745 2225
rect -745 2159 745 2197
rect -745 2131 -740 2159
rect -712 2131 -674 2159
rect -646 2131 -608 2159
rect -580 2131 -542 2159
rect -514 2131 -476 2159
rect -448 2131 -410 2159
rect -382 2131 -344 2159
rect -316 2131 -278 2159
rect -250 2131 -212 2159
rect -184 2131 -146 2159
rect -118 2131 -80 2159
rect -52 2131 -14 2159
rect 14 2131 52 2159
rect 80 2131 118 2159
rect 146 2131 184 2159
rect 212 2131 250 2159
rect 278 2131 316 2159
rect 344 2131 382 2159
rect 410 2131 448 2159
rect 476 2131 514 2159
rect 542 2131 580 2159
rect 608 2131 646 2159
rect 674 2131 712 2159
rect 740 2131 745 2159
rect -745 2093 745 2131
rect -745 2065 -740 2093
rect -712 2065 -674 2093
rect -646 2065 -608 2093
rect -580 2065 -542 2093
rect -514 2065 -476 2093
rect -448 2065 -410 2093
rect -382 2065 -344 2093
rect -316 2065 -278 2093
rect -250 2065 -212 2093
rect -184 2065 -146 2093
rect -118 2065 -80 2093
rect -52 2065 -14 2093
rect 14 2065 52 2093
rect 80 2065 118 2093
rect 146 2065 184 2093
rect 212 2065 250 2093
rect 278 2065 316 2093
rect 344 2065 382 2093
rect 410 2065 448 2093
rect 476 2065 514 2093
rect 542 2065 580 2093
rect 608 2065 646 2093
rect 674 2065 712 2093
rect 740 2065 745 2093
rect -745 2027 745 2065
rect -745 1999 -740 2027
rect -712 1999 -674 2027
rect -646 1999 -608 2027
rect -580 1999 -542 2027
rect -514 1999 -476 2027
rect -448 1999 -410 2027
rect -382 1999 -344 2027
rect -316 1999 -278 2027
rect -250 1999 -212 2027
rect -184 1999 -146 2027
rect -118 1999 -80 2027
rect -52 1999 -14 2027
rect 14 1999 52 2027
rect 80 1999 118 2027
rect 146 1999 184 2027
rect 212 1999 250 2027
rect 278 1999 316 2027
rect 344 1999 382 2027
rect 410 1999 448 2027
rect 476 1999 514 2027
rect 542 1999 580 2027
rect 608 1999 646 2027
rect 674 1999 712 2027
rect 740 1999 745 2027
rect -745 1961 745 1999
rect -745 1933 -740 1961
rect -712 1933 -674 1961
rect -646 1933 -608 1961
rect -580 1933 -542 1961
rect -514 1933 -476 1961
rect -448 1933 -410 1961
rect -382 1933 -344 1961
rect -316 1933 -278 1961
rect -250 1933 -212 1961
rect -184 1933 -146 1961
rect -118 1933 -80 1961
rect -52 1933 -14 1961
rect 14 1933 52 1961
rect 80 1933 118 1961
rect 146 1933 184 1961
rect 212 1933 250 1961
rect 278 1933 316 1961
rect 344 1933 382 1961
rect 410 1933 448 1961
rect 476 1933 514 1961
rect 542 1933 580 1961
rect 608 1933 646 1961
rect 674 1933 712 1961
rect 740 1933 745 1961
rect -745 1895 745 1933
rect -745 1867 -740 1895
rect -712 1867 -674 1895
rect -646 1867 -608 1895
rect -580 1867 -542 1895
rect -514 1867 -476 1895
rect -448 1867 -410 1895
rect -382 1867 -344 1895
rect -316 1867 -278 1895
rect -250 1867 -212 1895
rect -184 1867 -146 1895
rect -118 1867 -80 1895
rect -52 1867 -14 1895
rect 14 1867 52 1895
rect 80 1867 118 1895
rect 146 1867 184 1895
rect 212 1867 250 1895
rect 278 1867 316 1895
rect 344 1867 382 1895
rect 410 1867 448 1895
rect 476 1867 514 1895
rect 542 1867 580 1895
rect 608 1867 646 1895
rect 674 1867 712 1895
rect 740 1867 745 1895
rect -745 1829 745 1867
rect -745 1801 -740 1829
rect -712 1801 -674 1829
rect -646 1801 -608 1829
rect -580 1801 -542 1829
rect -514 1801 -476 1829
rect -448 1801 -410 1829
rect -382 1801 -344 1829
rect -316 1801 -278 1829
rect -250 1801 -212 1829
rect -184 1801 -146 1829
rect -118 1801 -80 1829
rect -52 1801 -14 1829
rect 14 1801 52 1829
rect 80 1801 118 1829
rect 146 1801 184 1829
rect 212 1801 250 1829
rect 278 1801 316 1829
rect 344 1801 382 1829
rect 410 1801 448 1829
rect 476 1801 514 1829
rect 542 1801 580 1829
rect 608 1801 646 1829
rect 674 1801 712 1829
rect 740 1801 745 1829
rect -745 1763 745 1801
rect -745 1735 -740 1763
rect -712 1735 -674 1763
rect -646 1735 -608 1763
rect -580 1735 -542 1763
rect -514 1735 -476 1763
rect -448 1735 -410 1763
rect -382 1735 -344 1763
rect -316 1735 -278 1763
rect -250 1735 -212 1763
rect -184 1735 -146 1763
rect -118 1735 -80 1763
rect -52 1735 -14 1763
rect 14 1735 52 1763
rect 80 1735 118 1763
rect 146 1735 184 1763
rect 212 1735 250 1763
rect 278 1735 316 1763
rect 344 1735 382 1763
rect 410 1735 448 1763
rect 476 1735 514 1763
rect 542 1735 580 1763
rect 608 1735 646 1763
rect 674 1735 712 1763
rect 740 1735 745 1763
rect -745 1697 745 1735
rect -745 1669 -740 1697
rect -712 1669 -674 1697
rect -646 1669 -608 1697
rect -580 1669 -542 1697
rect -514 1669 -476 1697
rect -448 1669 -410 1697
rect -382 1669 -344 1697
rect -316 1669 -278 1697
rect -250 1669 -212 1697
rect -184 1669 -146 1697
rect -118 1669 -80 1697
rect -52 1669 -14 1697
rect 14 1669 52 1697
rect 80 1669 118 1697
rect 146 1669 184 1697
rect 212 1669 250 1697
rect 278 1669 316 1697
rect 344 1669 382 1697
rect 410 1669 448 1697
rect 476 1669 514 1697
rect 542 1669 580 1697
rect 608 1669 646 1697
rect 674 1669 712 1697
rect 740 1669 745 1697
rect -745 1631 745 1669
rect -745 1603 -740 1631
rect -712 1603 -674 1631
rect -646 1603 -608 1631
rect -580 1603 -542 1631
rect -514 1603 -476 1631
rect -448 1603 -410 1631
rect -382 1603 -344 1631
rect -316 1603 -278 1631
rect -250 1603 -212 1631
rect -184 1603 -146 1631
rect -118 1603 -80 1631
rect -52 1603 -14 1631
rect 14 1603 52 1631
rect 80 1603 118 1631
rect 146 1603 184 1631
rect 212 1603 250 1631
rect 278 1603 316 1631
rect 344 1603 382 1631
rect 410 1603 448 1631
rect 476 1603 514 1631
rect 542 1603 580 1631
rect 608 1603 646 1631
rect 674 1603 712 1631
rect 740 1603 745 1631
rect -745 1565 745 1603
rect -745 1537 -740 1565
rect -712 1537 -674 1565
rect -646 1537 -608 1565
rect -580 1537 -542 1565
rect -514 1537 -476 1565
rect -448 1537 -410 1565
rect -382 1537 -344 1565
rect -316 1537 -278 1565
rect -250 1537 -212 1565
rect -184 1537 -146 1565
rect -118 1537 -80 1565
rect -52 1537 -14 1565
rect 14 1537 52 1565
rect 80 1537 118 1565
rect 146 1537 184 1565
rect 212 1537 250 1565
rect 278 1537 316 1565
rect 344 1537 382 1565
rect 410 1537 448 1565
rect 476 1537 514 1565
rect 542 1537 580 1565
rect 608 1537 646 1565
rect 674 1537 712 1565
rect 740 1537 745 1565
rect -745 1499 745 1537
rect -745 1471 -740 1499
rect -712 1471 -674 1499
rect -646 1471 -608 1499
rect -580 1471 -542 1499
rect -514 1471 -476 1499
rect -448 1471 -410 1499
rect -382 1471 -344 1499
rect -316 1471 -278 1499
rect -250 1471 -212 1499
rect -184 1471 -146 1499
rect -118 1471 -80 1499
rect -52 1471 -14 1499
rect 14 1471 52 1499
rect 80 1471 118 1499
rect 146 1471 184 1499
rect 212 1471 250 1499
rect 278 1471 316 1499
rect 344 1471 382 1499
rect 410 1471 448 1499
rect 476 1471 514 1499
rect 542 1471 580 1499
rect 608 1471 646 1499
rect 674 1471 712 1499
rect 740 1471 745 1499
rect -745 1433 745 1471
rect -745 1405 -740 1433
rect -712 1405 -674 1433
rect -646 1405 -608 1433
rect -580 1405 -542 1433
rect -514 1405 -476 1433
rect -448 1405 -410 1433
rect -382 1405 -344 1433
rect -316 1405 -278 1433
rect -250 1405 -212 1433
rect -184 1405 -146 1433
rect -118 1405 -80 1433
rect -52 1405 -14 1433
rect 14 1405 52 1433
rect 80 1405 118 1433
rect 146 1405 184 1433
rect 212 1405 250 1433
rect 278 1405 316 1433
rect 344 1405 382 1433
rect 410 1405 448 1433
rect 476 1405 514 1433
rect 542 1405 580 1433
rect 608 1405 646 1433
rect 674 1405 712 1433
rect 740 1405 745 1433
rect -745 1367 745 1405
rect -745 1339 -740 1367
rect -712 1339 -674 1367
rect -646 1339 -608 1367
rect -580 1339 -542 1367
rect -514 1339 -476 1367
rect -448 1339 -410 1367
rect -382 1339 -344 1367
rect -316 1339 -278 1367
rect -250 1339 -212 1367
rect -184 1339 -146 1367
rect -118 1339 -80 1367
rect -52 1339 -14 1367
rect 14 1339 52 1367
rect 80 1339 118 1367
rect 146 1339 184 1367
rect 212 1339 250 1367
rect 278 1339 316 1367
rect 344 1339 382 1367
rect 410 1339 448 1367
rect 476 1339 514 1367
rect 542 1339 580 1367
rect 608 1339 646 1367
rect 674 1339 712 1367
rect 740 1339 745 1367
rect -745 1301 745 1339
rect -745 1273 -740 1301
rect -712 1273 -674 1301
rect -646 1273 -608 1301
rect -580 1273 -542 1301
rect -514 1273 -476 1301
rect -448 1273 -410 1301
rect -382 1273 -344 1301
rect -316 1273 -278 1301
rect -250 1273 -212 1301
rect -184 1273 -146 1301
rect -118 1273 -80 1301
rect -52 1273 -14 1301
rect 14 1273 52 1301
rect 80 1273 118 1301
rect 146 1273 184 1301
rect 212 1273 250 1301
rect 278 1273 316 1301
rect 344 1273 382 1301
rect 410 1273 448 1301
rect 476 1273 514 1301
rect 542 1273 580 1301
rect 608 1273 646 1301
rect 674 1273 712 1301
rect 740 1273 745 1301
rect -745 1235 745 1273
rect -745 1207 -740 1235
rect -712 1207 -674 1235
rect -646 1207 -608 1235
rect -580 1207 -542 1235
rect -514 1207 -476 1235
rect -448 1207 -410 1235
rect -382 1207 -344 1235
rect -316 1207 -278 1235
rect -250 1207 -212 1235
rect -184 1207 -146 1235
rect -118 1207 -80 1235
rect -52 1207 -14 1235
rect 14 1207 52 1235
rect 80 1207 118 1235
rect 146 1207 184 1235
rect 212 1207 250 1235
rect 278 1207 316 1235
rect 344 1207 382 1235
rect 410 1207 448 1235
rect 476 1207 514 1235
rect 542 1207 580 1235
rect 608 1207 646 1235
rect 674 1207 712 1235
rect 740 1207 745 1235
rect -745 1169 745 1207
rect -745 1141 -740 1169
rect -712 1141 -674 1169
rect -646 1141 -608 1169
rect -580 1141 -542 1169
rect -514 1141 -476 1169
rect -448 1141 -410 1169
rect -382 1141 -344 1169
rect -316 1141 -278 1169
rect -250 1141 -212 1169
rect -184 1141 -146 1169
rect -118 1141 -80 1169
rect -52 1141 -14 1169
rect 14 1141 52 1169
rect 80 1141 118 1169
rect 146 1141 184 1169
rect 212 1141 250 1169
rect 278 1141 316 1169
rect 344 1141 382 1169
rect 410 1141 448 1169
rect 476 1141 514 1169
rect 542 1141 580 1169
rect 608 1141 646 1169
rect 674 1141 712 1169
rect 740 1141 745 1169
rect -745 1103 745 1141
rect -745 1075 -740 1103
rect -712 1075 -674 1103
rect -646 1075 -608 1103
rect -580 1075 -542 1103
rect -514 1075 -476 1103
rect -448 1075 -410 1103
rect -382 1075 -344 1103
rect -316 1075 -278 1103
rect -250 1075 -212 1103
rect -184 1075 -146 1103
rect -118 1075 -80 1103
rect -52 1075 -14 1103
rect 14 1075 52 1103
rect 80 1075 118 1103
rect 146 1075 184 1103
rect 212 1075 250 1103
rect 278 1075 316 1103
rect 344 1075 382 1103
rect 410 1075 448 1103
rect 476 1075 514 1103
rect 542 1075 580 1103
rect 608 1075 646 1103
rect 674 1075 712 1103
rect 740 1075 745 1103
rect -745 1037 745 1075
rect -745 1009 -740 1037
rect -712 1009 -674 1037
rect -646 1009 -608 1037
rect -580 1009 -542 1037
rect -514 1009 -476 1037
rect -448 1009 -410 1037
rect -382 1009 -344 1037
rect -316 1009 -278 1037
rect -250 1009 -212 1037
rect -184 1009 -146 1037
rect -118 1009 -80 1037
rect -52 1009 -14 1037
rect 14 1009 52 1037
rect 80 1009 118 1037
rect 146 1009 184 1037
rect 212 1009 250 1037
rect 278 1009 316 1037
rect 344 1009 382 1037
rect 410 1009 448 1037
rect 476 1009 514 1037
rect 542 1009 580 1037
rect 608 1009 646 1037
rect 674 1009 712 1037
rect 740 1009 745 1037
rect -745 971 745 1009
rect -745 943 -740 971
rect -712 943 -674 971
rect -646 943 -608 971
rect -580 943 -542 971
rect -514 943 -476 971
rect -448 943 -410 971
rect -382 943 -344 971
rect -316 943 -278 971
rect -250 943 -212 971
rect -184 943 -146 971
rect -118 943 -80 971
rect -52 943 -14 971
rect 14 943 52 971
rect 80 943 118 971
rect 146 943 184 971
rect 212 943 250 971
rect 278 943 316 971
rect 344 943 382 971
rect 410 943 448 971
rect 476 943 514 971
rect 542 943 580 971
rect 608 943 646 971
rect 674 943 712 971
rect 740 943 745 971
rect -745 905 745 943
rect -745 877 -740 905
rect -712 877 -674 905
rect -646 877 -608 905
rect -580 877 -542 905
rect -514 877 -476 905
rect -448 877 -410 905
rect -382 877 -344 905
rect -316 877 -278 905
rect -250 877 -212 905
rect -184 877 -146 905
rect -118 877 -80 905
rect -52 877 -14 905
rect 14 877 52 905
rect 80 877 118 905
rect 146 877 184 905
rect 212 877 250 905
rect 278 877 316 905
rect 344 877 382 905
rect 410 877 448 905
rect 476 877 514 905
rect 542 877 580 905
rect 608 877 646 905
rect 674 877 712 905
rect 740 877 745 905
rect -745 839 745 877
rect -745 811 -740 839
rect -712 811 -674 839
rect -646 811 -608 839
rect -580 811 -542 839
rect -514 811 -476 839
rect -448 811 -410 839
rect -382 811 -344 839
rect -316 811 -278 839
rect -250 811 -212 839
rect -184 811 -146 839
rect -118 811 -80 839
rect -52 811 -14 839
rect 14 811 52 839
rect 80 811 118 839
rect 146 811 184 839
rect 212 811 250 839
rect 278 811 316 839
rect 344 811 382 839
rect 410 811 448 839
rect 476 811 514 839
rect 542 811 580 839
rect 608 811 646 839
rect 674 811 712 839
rect 740 811 745 839
rect -745 773 745 811
rect -745 745 -740 773
rect -712 745 -674 773
rect -646 745 -608 773
rect -580 745 -542 773
rect -514 745 -476 773
rect -448 745 -410 773
rect -382 745 -344 773
rect -316 745 -278 773
rect -250 745 -212 773
rect -184 745 -146 773
rect -118 745 -80 773
rect -52 745 -14 773
rect 14 745 52 773
rect 80 745 118 773
rect 146 745 184 773
rect 212 745 250 773
rect 278 745 316 773
rect 344 745 382 773
rect 410 745 448 773
rect 476 745 514 773
rect 542 745 580 773
rect 608 745 646 773
rect 674 745 712 773
rect 740 745 745 773
rect -745 707 745 745
rect -745 679 -740 707
rect -712 679 -674 707
rect -646 679 -608 707
rect -580 679 -542 707
rect -514 679 -476 707
rect -448 679 -410 707
rect -382 679 -344 707
rect -316 679 -278 707
rect -250 679 -212 707
rect -184 679 -146 707
rect -118 679 -80 707
rect -52 679 -14 707
rect 14 679 52 707
rect 80 679 118 707
rect 146 679 184 707
rect 212 679 250 707
rect 278 679 316 707
rect 344 679 382 707
rect 410 679 448 707
rect 476 679 514 707
rect 542 679 580 707
rect 608 679 646 707
rect 674 679 712 707
rect 740 679 745 707
rect -745 641 745 679
rect -745 613 -740 641
rect -712 613 -674 641
rect -646 613 -608 641
rect -580 613 -542 641
rect -514 613 -476 641
rect -448 613 -410 641
rect -382 613 -344 641
rect -316 613 -278 641
rect -250 613 -212 641
rect -184 613 -146 641
rect -118 613 -80 641
rect -52 613 -14 641
rect 14 613 52 641
rect 80 613 118 641
rect 146 613 184 641
rect 212 613 250 641
rect 278 613 316 641
rect 344 613 382 641
rect 410 613 448 641
rect 476 613 514 641
rect 542 613 580 641
rect 608 613 646 641
rect 674 613 712 641
rect 740 613 745 641
rect -745 575 745 613
rect -745 547 -740 575
rect -712 547 -674 575
rect -646 547 -608 575
rect -580 547 -542 575
rect -514 547 -476 575
rect -448 547 -410 575
rect -382 547 -344 575
rect -316 547 -278 575
rect -250 547 -212 575
rect -184 547 -146 575
rect -118 547 -80 575
rect -52 547 -14 575
rect 14 547 52 575
rect 80 547 118 575
rect 146 547 184 575
rect 212 547 250 575
rect 278 547 316 575
rect 344 547 382 575
rect 410 547 448 575
rect 476 547 514 575
rect 542 547 580 575
rect 608 547 646 575
rect 674 547 712 575
rect 740 547 745 575
rect -745 509 745 547
rect -745 481 -740 509
rect -712 481 -674 509
rect -646 481 -608 509
rect -580 481 -542 509
rect -514 481 -476 509
rect -448 481 -410 509
rect -382 481 -344 509
rect -316 481 -278 509
rect -250 481 -212 509
rect -184 481 -146 509
rect -118 481 -80 509
rect -52 481 -14 509
rect 14 481 52 509
rect 80 481 118 509
rect 146 481 184 509
rect 212 481 250 509
rect 278 481 316 509
rect 344 481 382 509
rect 410 481 448 509
rect 476 481 514 509
rect 542 481 580 509
rect 608 481 646 509
rect 674 481 712 509
rect 740 481 745 509
rect -745 443 745 481
rect -745 415 -740 443
rect -712 415 -674 443
rect -646 415 -608 443
rect -580 415 -542 443
rect -514 415 -476 443
rect -448 415 -410 443
rect -382 415 -344 443
rect -316 415 -278 443
rect -250 415 -212 443
rect -184 415 -146 443
rect -118 415 -80 443
rect -52 415 -14 443
rect 14 415 52 443
rect 80 415 118 443
rect 146 415 184 443
rect 212 415 250 443
rect 278 415 316 443
rect 344 415 382 443
rect 410 415 448 443
rect 476 415 514 443
rect 542 415 580 443
rect 608 415 646 443
rect 674 415 712 443
rect 740 415 745 443
rect -745 377 745 415
rect -745 349 -740 377
rect -712 349 -674 377
rect -646 349 -608 377
rect -580 349 -542 377
rect -514 349 -476 377
rect -448 349 -410 377
rect -382 349 -344 377
rect -316 349 -278 377
rect -250 349 -212 377
rect -184 349 -146 377
rect -118 349 -80 377
rect -52 349 -14 377
rect 14 349 52 377
rect 80 349 118 377
rect 146 349 184 377
rect 212 349 250 377
rect 278 349 316 377
rect 344 349 382 377
rect 410 349 448 377
rect 476 349 514 377
rect 542 349 580 377
rect 608 349 646 377
rect 674 349 712 377
rect 740 349 745 377
rect -745 311 745 349
rect -745 283 -740 311
rect -712 283 -674 311
rect -646 283 -608 311
rect -580 283 -542 311
rect -514 283 -476 311
rect -448 283 -410 311
rect -382 283 -344 311
rect -316 283 -278 311
rect -250 283 -212 311
rect -184 283 -146 311
rect -118 283 -80 311
rect -52 283 -14 311
rect 14 283 52 311
rect 80 283 118 311
rect 146 283 184 311
rect 212 283 250 311
rect 278 283 316 311
rect 344 283 382 311
rect 410 283 448 311
rect 476 283 514 311
rect 542 283 580 311
rect 608 283 646 311
rect 674 283 712 311
rect 740 283 745 311
rect -745 245 745 283
rect -745 217 -740 245
rect -712 217 -674 245
rect -646 217 -608 245
rect -580 217 -542 245
rect -514 217 -476 245
rect -448 217 -410 245
rect -382 217 -344 245
rect -316 217 -278 245
rect -250 217 -212 245
rect -184 217 -146 245
rect -118 217 -80 245
rect -52 217 -14 245
rect 14 217 52 245
rect 80 217 118 245
rect 146 217 184 245
rect 212 217 250 245
rect 278 217 316 245
rect 344 217 382 245
rect 410 217 448 245
rect 476 217 514 245
rect 542 217 580 245
rect 608 217 646 245
rect 674 217 712 245
rect 740 217 745 245
rect -745 179 745 217
rect -745 151 -740 179
rect -712 151 -674 179
rect -646 151 -608 179
rect -580 151 -542 179
rect -514 151 -476 179
rect -448 151 -410 179
rect -382 151 -344 179
rect -316 151 -278 179
rect -250 151 -212 179
rect -184 151 -146 179
rect -118 151 -80 179
rect -52 151 -14 179
rect 14 151 52 179
rect 80 151 118 179
rect 146 151 184 179
rect 212 151 250 179
rect 278 151 316 179
rect 344 151 382 179
rect 410 151 448 179
rect 476 151 514 179
rect 542 151 580 179
rect 608 151 646 179
rect 674 151 712 179
rect 740 151 745 179
rect -745 113 745 151
rect -745 85 -740 113
rect -712 85 -674 113
rect -646 85 -608 113
rect -580 85 -542 113
rect -514 85 -476 113
rect -448 85 -410 113
rect -382 85 -344 113
rect -316 85 -278 113
rect -250 85 -212 113
rect -184 85 -146 113
rect -118 85 -80 113
rect -52 85 -14 113
rect 14 85 52 113
rect 80 85 118 113
rect 146 85 184 113
rect 212 85 250 113
rect 278 85 316 113
rect 344 85 382 113
rect 410 85 448 113
rect 476 85 514 113
rect 542 85 580 113
rect 608 85 646 113
rect 674 85 712 113
rect 740 85 745 113
rect -745 47 745 85
rect -745 19 -740 47
rect -712 19 -674 47
rect -646 19 -608 47
rect -580 19 -542 47
rect -514 19 -476 47
rect -448 19 -410 47
rect -382 19 -344 47
rect -316 19 -278 47
rect -250 19 -212 47
rect -184 19 -146 47
rect -118 19 -80 47
rect -52 19 -14 47
rect 14 19 52 47
rect 80 19 118 47
rect 146 19 184 47
rect 212 19 250 47
rect 278 19 316 47
rect 344 19 382 47
rect 410 19 448 47
rect 476 19 514 47
rect 542 19 580 47
rect 608 19 646 47
rect 674 19 712 47
rect 740 19 745 47
rect -745 -19 745 19
rect -745 -47 -740 -19
rect -712 -47 -674 -19
rect -646 -47 -608 -19
rect -580 -47 -542 -19
rect -514 -47 -476 -19
rect -448 -47 -410 -19
rect -382 -47 -344 -19
rect -316 -47 -278 -19
rect -250 -47 -212 -19
rect -184 -47 -146 -19
rect -118 -47 -80 -19
rect -52 -47 -14 -19
rect 14 -47 52 -19
rect 80 -47 118 -19
rect 146 -47 184 -19
rect 212 -47 250 -19
rect 278 -47 316 -19
rect 344 -47 382 -19
rect 410 -47 448 -19
rect 476 -47 514 -19
rect 542 -47 580 -19
rect 608 -47 646 -19
rect 674 -47 712 -19
rect 740 -47 745 -19
rect -745 -85 745 -47
rect -745 -113 -740 -85
rect -712 -113 -674 -85
rect -646 -113 -608 -85
rect -580 -113 -542 -85
rect -514 -113 -476 -85
rect -448 -113 -410 -85
rect -382 -113 -344 -85
rect -316 -113 -278 -85
rect -250 -113 -212 -85
rect -184 -113 -146 -85
rect -118 -113 -80 -85
rect -52 -113 -14 -85
rect 14 -113 52 -85
rect 80 -113 118 -85
rect 146 -113 184 -85
rect 212 -113 250 -85
rect 278 -113 316 -85
rect 344 -113 382 -85
rect 410 -113 448 -85
rect 476 -113 514 -85
rect 542 -113 580 -85
rect 608 -113 646 -85
rect 674 -113 712 -85
rect 740 -113 745 -85
rect -745 -151 745 -113
rect -745 -179 -740 -151
rect -712 -179 -674 -151
rect -646 -179 -608 -151
rect -580 -179 -542 -151
rect -514 -179 -476 -151
rect -448 -179 -410 -151
rect -382 -179 -344 -151
rect -316 -179 -278 -151
rect -250 -179 -212 -151
rect -184 -179 -146 -151
rect -118 -179 -80 -151
rect -52 -179 -14 -151
rect 14 -179 52 -151
rect 80 -179 118 -151
rect 146 -179 184 -151
rect 212 -179 250 -151
rect 278 -179 316 -151
rect 344 -179 382 -151
rect 410 -179 448 -151
rect 476 -179 514 -151
rect 542 -179 580 -151
rect 608 -179 646 -151
rect 674 -179 712 -151
rect 740 -179 745 -151
rect -745 -217 745 -179
rect -745 -245 -740 -217
rect -712 -245 -674 -217
rect -646 -245 -608 -217
rect -580 -245 -542 -217
rect -514 -245 -476 -217
rect -448 -245 -410 -217
rect -382 -245 -344 -217
rect -316 -245 -278 -217
rect -250 -245 -212 -217
rect -184 -245 -146 -217
rect -118 -245 -80 -217
rect -52 -245 -14 -217
rect 14 -245 52 -217
rect 80 -245 118 -217
rect 146 -245 184 -217
rect 212 -245 250 -217
rect 278 -245 316 -217
rect 344 -245 382 -217
rect 410 -245 448 -217
rect 476 -245 514 -217
rect 542 -245 580 -217
rect 608 -245 646 -217
rect 674 -245 712 -217
rect 740 -245 745 -217
rect -745 -283 745 -245
rect -745 -311 -740 -283
rect -712 -311 -674 -283
rect -646 -311 -608 -283
rect -580 -311 -542 -283
rect -514 -311 -476 -283
rect -448 -311 -410 -283
rect -382 -311 -344 -283
rect -316 -311 -278 -283
rect -250 -311 -212 -283
rect -184 -311 -146 -283
rect -118 -311 -80 -283
rect -52 -311 -14 -283
rect 14 -311 52 -283
rect 80 -311 118 -283
rect 146 -311 184 -283
rect 212 -311 250 -283
rect 278 -311 316 -283
rect 344 -311 382 -283
rect 410 -311 448 -283
rect 476 -311 514 -283
rect 542 -311 580 -283
rect 608 -311 646 -283
rect 674 -311 712 -283
rect 740 -311 745 -283
rect -745 -349 745 -311
rect -745 -377 -740 -349
rect -712 -377 -674 -349
rect -646 -377 -608 -349
rect -580 -377 -542 -349
rect -514 -377 -476 -349
rect -448 -377 -410 -349
rect -382 -377 -344 -349
rect -316 -377 -278 -349
rect -250 -377 -212 -349
rect -184 -377 -146 -349
rect -118 -377 -80 -349
rect -52 -377 -14 -349
rect 14 -377 52 -349
rect 80 -377 118 -349
rect 146 -377 184 -349
rect 212 -377 250 -349
rect 278 -377 316 -349
rect 344 -377 382 -349
rect 410 -377 448 -349
rect 476 -377 514 -349
rect 542 -377 580 -349
rect 608 -377 646 -349
rect 674 -377 712 -349
rect 740 -377 745 -349
rect -745 -415 745 -377
rect -745 -443 -740 -415
rect -712 -443 -674 -415
rect -646 -443 -608 -415
rect -580 -443 -542 -415
rect -514 -443 -476 -415
rect -448 -443 -410 -415
rect -382 -443 -344 -415
rect -316 -443 -278 -415
rect -250 -443 -212 -415
rect -184 -443 -146 -415
rect -118 -443 -80 -415
rect -52 -443 -14 -415
rect 14 -443 52 -415
rect 80 -443 118 -415
rect 146 -443 184 -415
rect 212 -443 250 -415
rect 278 -443 316 -415
rect 344 -443 382 -415
rect 410 -443 448 -415
rect 476 -443 514 -415
rect 542 -443 580 -415
rect 608 -443 646 -415
rect 674 -443 712 -415
rect 740 -443 745 -415
rect -745 -481 745 -443
rect -745 -509 -740 -481
rect -712 -509 -674 -481
rect -646 -509 -608 -481
rect -580 -509 -542 -481
rect -514 -509 -476 -481
rect -448 -509 -410 -481
rect -382 -509 -344 -481
rect -316 -509 -278 -481
rect -250 -509 -212 -481
rect -184 -509 -146 -481
rect -118 -509 -80 -481
rect -52 -509 -14 -481
rect 14 -509 52 -481
rect 80 -509 118 -481
rect 146 -509 184 -481
rect 212 -509 250 -481
rect 278 -509 316 -481
rect 344 -509 382 -481
rect 410 -509 448 -481
rect 476 -509 514 -481
rect 542 -509 580 -481
rect 608 -509 646 -481
rect 674 -509 712 -481
rect 740 -509 745 -481
rect -745 -547 745 -509
rect -745 -575 -740 -547
rect -712 -575 -674 -547
rect -646 -575 -608 -547
rect -580 -575 -542 -547
rect -514 -575 -476 -547
rect -448 -575 -410 -547
rect -382 -575 -344 -547
rect -316 -575 -278 -547
rect -250 -575 -212 -547
rect -184 -575 -146 -547
rect -118 -575 -80 -547
rect -52 -575 -14 -547
rect 14 -575 52 -547
rect 80 -575 118 -547
rect 146 -575 184 -547
rect 212 -575 250 -547
rect 278 -575 316 -547
rect 344 -575 382 -547
rect 410 -575 448 -547
rect 476 -575 514 -547
rect 542 -575 580 -547
rect 608 -575 646 -547
rect 674 -575 712 -547
rect 740 -575 745 -547
rect -745 -613 745 -575
rect -745 -641 -740 -613
rect -712 -641 -674 -613
rect -646 -641 -608 -613
rect -580 -641 -542 -613
rect -514 -641 -476 -613
rect -448 -641 -410 -613
rect -382 -641 -344 -613
rect -316 -641 -278 -613
rect -250 -641 -212 -613
rect -184 -641 -146 -613
rect -118 -641 -80 -613
rect -52 -641 -14 -613
rect 14 -641 52 -613
rect 80 -641 118 -613
rect 146 -641 184 -613
rect 212 -641 250 -613
rect 278 -641 316 -613
rect 344 -641 382 -613
rect 410 -641 448 -613
rect 476 -641 514 -613
rect 542 -641 580 -613
rect 608 -641 646 -613
rect 674 -641 712 -613
rect 740 -641 745 -613
rect -745 -679 745 -641
rect -745 -707 -740 -679
rect -712 -707 -674 -679
rect -646 -707 -608 -679
rect -580 -707 -542 -679
rect -514 -707 -476 -679
rect -448 -707 -410 -679
rect -382 -707 -344 -679
rect -316 -707 -278 -679
rect -250 -707 -212 -679
rect -184 -707 -146 -679
rect -118 -707 -80 -679
rect -52 -707 -14 -679
rect 14 -707 52 -679
rect 80 -707 118 -679
rect 146 -707 184 -679
rect 212 -707 250 -679
rect 278 -707 316 -679
rect 344 -707 382 -679
rect 410 -707 448 -679
rect 476 -707 514 -679
rect 542 -707 580 -679
rect 608 -707 646 -679
rect 674 -707 712 -679
rect 740 -707 745 -679
rect -745 -745 745 -707
rect -745 -773 -740 -745
rect -712 -773 -674 -745
rect -646 -773 -608 -745
rect -580 -773 -542 -745
rect -514 -773 -476 -745
rect -448 -773 -410 -745
rect -382 -773 -344 -745
rect -316 -773 -278 -745
rect -250 -773 -212 -745
rect -184 -773 -146 -745
rect -118 -773 -80 -745
rect -52 -773 -14 -745
rect 14 -773 52 -745
rect 80 -773 118 -745
rect 146 -773 184 -745
rect 212 -773 250 -745
rect 278 -773 316 -745
rect 344 -773 382 -745
rect 410 -773 448 -745
rect 476 -773 514 -745
rect 542 -773 580 -745
rect 608 -773 646 -745
rect 674 -773 712 -745
rect 740 -773 745 -745
rect -745 -811 745 -773
rect -745 -839 -740 -811
rect -712 -839 -674 -811
rect -646 -839 -608 -811
rect -580 -839 -542 -811
rect -514 -839 -476 -811
rect -448 -839 -410 -811
rect -382 -839 -344 -811
rect -316 -839 -278 -811
rect -250 -839 -212 -811
rect -184 -839 -146 -811
rect -118 -839 -80 -811
rect -52 -839 -14 -811
rect 14 -839 52 -811
rect 80 -839 118 -811
rect 146 -839 184 -811
rect 212 -839 250 -811
rect 278 -839 316 -811
rect 344 -839 382 -811
rect 410 -839 448 -811
rect 476 -839 514 -811
rect 542 -839 580 -811
rect 608 -839 646 -811
rect 674 -839 712 -811
rect 740 -839 745 -811
rect -745 -877 745 -839
rect -745 -905 -740 -877
rect -712 -905 -674 -877
rect -646 -905 -608 -877
rect -580 -905 -542 -877
rect -514 -905 -476 -877
rect -448 -905 -410 -877
rect -382 -905 -344 -877
rect -316 -905 -278 -877
rect -250 -905 -212 -877
rect -184 -905 -146 -877
rect -118 -905 -80 -877
rect -52 -905 -14 -877
rect 14 -905 52 -877
rect 80 -905 118 -877
rect 146 -905 184 -877
rect 212 -905 250 -877
rect 278 -905 316 -877
rect 344 -905 382 -877
rect 410 -905 448 -877
rect 476 -905 514 -877
rect 542 -905 580 -877
rect 608 -905 646 -877
rect 674 -905 712 -877
rect 740 -905 745 -877
rect -745 -943 745 -905
rect -745 -971 -740 -943
rect -712 -971 -674 -943
rect -646 -971 -608 -943
rect -580 -971 -542 -943
rect -514 -971 -476 -943
rect -448 -971 -410 -943
rect -382 -971 -344 -943
rect -316 -971 -278 -943
rect -250 -971 -212 -943
rect -184 -971 -146 -943
rect -118 -971 -80 -943
rect -52 -971 -14 -943
rect 14 -971 52 -943
rect 80 -971 118 -943
rect 146 -971 184 -943
rect 212 -971 250 -943
rect 278 -971 316 -943
rect 344 -971 382 -943
rect 410 -971 448 -943
rect 476 -971 514 -943
rect 542 -971 580 -943
rect 608 -971 646 -943
rect 674 -971 712 -943
rect 740 -971 745 -943
rect -745 -1009 745 -971
rect -745 -1037 -740 -1009
rect -712 -1037 -674 -1009
rect -646 -1037 -608 -1009
rect -580 -1037 -542 -1009
rect -514 -1037 -476 -1009
rect -448 -1037 -410 -1009
rect -382 -1037 -344 -1009
rect -316 -1037 -278 -1009
rect -250 -1037 -212 -1009
rect -184 -1037 -146 -1009
rect -118 -1037 -80 -1009
rect -52 -1037 -14 -1009
rect 14 -1037 52 -1009
rect 80 -1037 118 -1009
rect 146 -1037 184 -1009
rect 212 -1037 250 -1009
rect 278 -1037 316 -1009
rect 344 -1037 382 -1009
rect 410 -1037 448 -1009
rect 476 -1037 514 -1009
rect 542 -1037 580 -1009
rect 608 -1037 646 -1009
rect 674 -1037 712 -1009
rect 740 -1037 745 -1009
rect -745 -1075 745 -1037
rect -745 -1103 -740 -1075
rect -712 -1103 -674 -1075
rect -646 -1103 -608 -1075
rect -580 -1103 -542 -1075
rect -514 -1103 -476 -1075
rect -448 -1103 -410 -1075
rect -382 -1103 -344 -1075
rect -316 -1103 -278 -1075
rect -250 -1103 -212 -1075
rect -184 -1103 -146 -1075
rect -118 -1103 -80 -1075
rect -52 -1103 -14 -1075
rect 14 -1103 52 -1075
rect 80 -1103 118 -1075
rect 146 -1103 184 -1075
rect 212 -1103 250 -1075
rect 278 -1103 316 -1075
rect 344 -1103 382 -1075
rect 410 -1103 448 -1075
rect 476 -1103 514 -1075
rect 542 -1103 580 -1075
rect 608 -1103 646 -1075
rect 674 -1103 712 -1075
rect 740 -1103 745 -1075
rect -745 -1141 745 -1103
rect -745 -1169 -740 -1141
rect -712 -1169 -674 -1141
rect -646 -1169 -608 -1141
rect -580 -1169 -542 -1141
rect -514 -1169 -476 -1141
rect -448 -1169 -410 -1141
rect -382 -1169 -344 -1141
rect -316 -1169 -278 -1141
rect -250 -1169 -212 -1141
rect -184 -1169 -146 -1141
rect -118 -1169 -80 -1141
rect -52 -1169 -14 -1141
rect 14 -1169 52 -1141
rect 80 -1169 118 -1141
rect 146 -1169 184 -1141
rect 212 -1169 250 -1141
rect 278 -1169 316 -1141
rect 344 -1169 382 -1141
rect 410 -1169 448 -1141
rect 476 -1169 514 -1141
rect 542 -1169 580 -1141
rect 608 -1169 646 -1141
rect 674 -1169 712 -1141
rect 740 -1169 745 -1141
rect -745 -1207 745 -1169
rect -745 -1235 -740 -1207
rect -712 -1235 -674 -1207
rect -646 -1235 -608 -1207
rect -580 -1235 -542 -1207
rect -514 -1235 -476 -1207
rect -448 -1235 -410 -1207
rect -382 -1235 -344 -1207
rect -316 -1235 -278 -1207
rect -250 -1235 -212 -1207
rect -184 -1235 -146 -1207
rect -118 -1235 -80 -1207
rect -52 -1235 -14 -1207
rect 14 -1235 52 -1207
rect 80 -1235 118 -1207
rect 146 -1235 184 -1207
rect 212 -1235 250 -1207
rect 278 -1235 316 -1207
rect 344 -1235 382 -1207
rect 410 -1235 448 -1207
rect 476 -1235 514 -1207
rect 542 -1235 580 -1207
rect 608 -1235 646 -1207
rect 674 -1235 712 -1207
rect 740 -1235 745 -1207
rect -745 -1273 745 -1235
rect -745 -1301 -740 -1273
rect -712 -1301 -674 -1273
rect -646 -1301 -608 -1273
rect -580 -1301 -542 -1273
rect -514 -1301 -476 -1273
rect -448 -1301 -410 -1273
rect -382 -1301 -344 -1273
rect -316 -1301 -278 -1273
rect -250 -1301 -212 -1273
rect -184 -1301 -146 -1273
rect -118 -1301 -80 -1273
rect -52 -1301 -14 -1273
rect 14 -1301 52 -1273
rect 80 -1301 118 -1273
rect 146 -1301 184 -1273
rect 212 -1301 250 -1273
rect 278 -1301 316 -1273
rect 344 -1301 382 -1273
rect 410 -1301 448 -1273
rect 476 -1301 514 -1273
rect 542 -1301 580 -1273
rect 608 -1301 646 -1273
rect 674 -1301 712 -1273
rect 740 -1301 745 -1273
rect -745 -1339 745 -1301
rect -745 -1367 -740 -1339
rect -712 -1367 -674 -1339
rect -646 -1367 -608 -1339
rect -580 -1367 -542 -1339
rect -514 -1367 -476 -1339
rect -448 -1367 -410 -1339
rect -382 -1367 -344 -1339
rect -316 -1367 -278 -1339
rect -250 -1367 -212 -1339
rect -184 -1367 -146 -1339
rect -118 -1367 -80 -1339
rect -52 -1367 -14 -1339
rect 14 -1367 52 -1339
rect 80 -1367 118 -1339
rect 146 -1367 184 -1339
rect 212 -1367 250 -1339
rect 278 -1367 316 -1339
rect 344 -1367 382 -1339
rect 410 -1367 448 -1339
rect 476 -1367 514 -1339
rect 542 -1367 580 -1339
rect 608 -1367 646 -1339
rect 674 -1367 712 -1339
rect 740 -1367 745 -1339
rect -745 -1405 745 -1367
rect -745 -1433 -740 -1405
rect -712 -1433 -674 -1405
rect -646 -1433 -608 -1405
rect -580 -1433 -542 -1405
rect -514 -1433 -476 -1405
rect -448 -1433 -410 -1405
rect -382 -1433 -344 -1405
rect -316 -1433 -278 -1405
rect -250 -1433 -212 -1405
rect -184 -1433 -146 -1405
rect -118 -1433 -80 -1405
rect -52 -1433 -14 -1405
rect 14 -1433 52 -1405
rect 80 -1433 118 -1405
rect 146 -1433 184 -1405
rect 212 -1433 250 -1405
rect 278 -1433 316 -1405
rect 344 -1433 382 -1405
rect 410 -1433 448 -1405
rect 476 -1433 514 -1405
rect 542 -1433 580 -1405
rect 608 -1433 646 -1405
rect 674 -1433 712 -1405
rect 740 -1433 745 -1405
rect -745 -1471 745 -1433
rect -745 -1499 -740 -1471
rect -712 -1499 -674 -1471
rect -646 -1499 -608 -1471
rect -580 -1499 -542 -1471
rect -514 -1499 -476 -1471
rect -448 -1499 -410 -1471
rect -382 -1499 -344 -1471
rect -316 -1499 -278 -1471
rect -250 -1499 -212 -1471
rect -184 -1499 -146 -1471
rect -118 -1499 -80 -1471
rect -52 -1499 -14 -1471
rect 14 -1499 52 -1471
rect 80 -1499 118 -1471
rect 146 -1499 184 -1471
rect 212 -1499 250 -1471
rect 278 -1499 316 -1471
rect 344 -1499 382 -1471
rect 410 -1499 448 -1471
rect 476 -1499 514 -1471
rect 542 -1499 580 -1471
rect 608 -1499 646 -1471
rect 674 -1499 712 -1471
rect 740 -1499 745 -1471
rect -745 -1537 745 -1499
rect -745 -1565 -740 -1537
rect -712 -1565 -674 -1537
rect -646 -1565 -608 -1537
rect -580 -1565 -542 -1537
rect -514 -1565 -476 -1537
rect -448 -1565 -410 -1537
rect -382 -1565 -344 -1537
rect -316 -1565 -278 -1537
rect -250 -1565 -212 -1537
rect -184 -1565 -146 -1537
rect -118 -1565 -80 -1537
rect -52 -1565 -14 -1537
rect 14 -1565 52 -1537
rect 80 -1565 118 -1537
rect 146 -1565 184 -1537
rect 212 -1565 250 -1537
rect 278 -1565 316 -1537
rect 344 -1565 382 -1537
rect 410 -1565 448 -1537
rect 476 -1565 514 -1537
rect 542 -1565 580 -1537
rect 608 -1565 646 -1537
rect 674 -1565 712 -1537
rect 740 -1565 745 -1537
rect -745 -1603 745 -1565
rect -745 -1631 -740 -1603
rect -712 -1631 -674 -1603
rect -646 -1631 -608 -1603
rect -580 -1631 -542 -1603
rect -514 -1631 -476 -1603
rect -448 -1631 -410 -1603
rect -382 -1631 -344 -1603
rect -316 -1631 -278 -1603
rect -250 -1631 -212 -1603
rect -184 -1631 -146 -1603
rect -118 -1631 -80 -1603
rect -52 -1631 -14 -1603
rect 14 -1631 52 -1603
rect 80 -1631 118 -1603
rect 146 -1631 184 -1603
rect 212 -1631 250 -1603
rect 278 -1631 316 -1603
rect 344 -1631 382 -1603
rect 410 -1631 448 -1603
rect 476 -1631 514 -1603
rect 542 -1631 580 -1603
rect 608 -1631 646 -1603
rect 674 -1631 712 -1603
rect 740 -1631 745 -1603
rect -745 -1669 745 -1631
rect -745 -1697 -740 -1669
rect -712 -1697 -674 -1669
rect -646 -1697 -608 -1669
rect -580 -1697 -542 -1669
rect -514 -1697 -476 -1669
rect -448 -1697 -410 -1669
rect -382 -1697 -344 -1669
rect -316 -1697 -278 -1669
rect -250 -1697 -212 -1669
rect -184 -1697 -146 -1669
rect -118 -1697 -80 -1669
rect -52 -1697 -14 -1669
rect 14 -1697 52 -1669
rect 80 -1697 118 -1669
rect 146 -1697 184 -1669
rect 212 -1697 250 -1669
rect 278 -1697 316 -1669
rect 344 -1697 382 -1669
rect 410 -1697 448 -1669
rect 476 -1697 514 -1669
rect 542 -1697 580 -1669
rect 608 -1697 646 -1669
rect 674 -1697 712 -1669
rect 740 -1697 745 -1669
rect -745 -1735 745 -1697
rect -745 -1763 -740 -1735
rect -712 -1763 -674 -1735
rect -646 -1763 -608 -1735
rect -580 -1763 -542 -1735
rect -514 -1763 -476 -1735
rect -448 -1763 -410 -1735
rect -382 -1763 -344 -1735
rect -316 -1763 -278 -1735
rect -250 -1763 -212 -1735
rect -184 -1763 -146 -1735
rect -118 -1763 -80 -1735
rect -52 -1763 -14 -1735
rect 14 -1763 52 -1735
rect 80 -1763 118 -1735
rect 146 -1763 184 -1735
rect 212 -1763 250 -1735
rect 278 -1763 316 -1735
rect 344 -1763 382 -1735
rect 410 -1763 448 -1735
rect 476 -1763 514 -1735
rect 542 -1763 580 -1735
rect 608 -1763 646 -1735
rect 674 -1763 712 -1735
rect 740 -1763 745 -1735
rect -745 -1801 745 -1763
rect -745 -1829 -740 -1801
rect -712 -1829 -674 -1801
rect -646 -1829 -608 -1801
rect -580 -1829 -542 -1801
rect -514 -1829 -476 -1801
rect -448 -1829 -410 -1801
rect -382 -1829 -344 -1801
rect -316 -1829 -278 -1801
rect -250 -1829 -212 -1801
rect -184 -1829 -146 -1801
rect -118 -1829 -80 -1801
rect -52 -1829 -14 -1801
rect 14 -1829 52 -1801
rect 80 -1829 118 -1801
rect 146 -1829 184 -1801
rect 212 -1829 250 -1801
rect 278 -1829 316 -1801
rect 344 -1829 382 -1801
rect 410 -1829 448 -1801
rect 476 -1829 514 -1801
rect 542 -1829 580 -1801
rect 608 -1829 646 -1801
rect 674 -1829 712 -1801
rect 740 -1829 745 -1801
rect -745 -1867 745 -1829
rect -745 -1895 -740 -1867
rect -712 -1895 -674 -1867
rect -646 -1895 -608 -1867
rect -580 -1895 -542 -1867
rect -514 -1895 -476 -1867
rect -448 -1895 -410 -1867
rect -382 -1895 -344 -1867
rect -316 -1895 -278 -1867
rect -250 -1895 -212 -1867
rect -184 -1895 -146 -1867
rect -118 -1895 -80 -1867
rect -52 -1895 -14 -1867
rect 14 -1895 52 -1867
rect 80 -1895 118 -1867
rect 146 -1895 184 -1867
rect 212 -1895 250 -1867
rect 278 -1895 316 -1867
rect 344 -1895 382 -1867
rect 410 -1895 448 -1867
rect 476 -1895 514 -1867
rect 542 -1895 580 -1867
rect 608 -1895 646 -1867
rect 674 -1895 712 -1867
rect 740 -1895 745 -1867
rect -745 -1933 745 -1895
rect -745 -1961 -740 -1933
rect -712 -1961 -674 -1933
rect -646 -1961 -608 -1933
rect -580 -1961 -542 -1933
rect -514 -1961 -476 -1933
rect -448 -1961 -410 -1933
rect -382 -1961 -344 -1933
rect -316 -1961 -278 -1933
rect -250 -1961 -212 -1933
rect -184 -1961 -146 -1933
rect -118 -1961 -80 -1933
rect -52 -1961 -14 -1933
rect 14 -1961 52 -1933
rect 80 -1961 118 -1933
rect 146 -1961 184 -1933
rect 212 -1961 250 -1933
rect 278 -1961 316 -1933
rect 344 -1961 382 -1933
rect 410 -1961 448 -1933
rect 476 -1961 514 -1933
rect 542 -1961 580 -1933
rect 608 -1961 646 -1933
rect 674 -1961 712 -1933
rect 740 -1961 745 -1933
rect -745 -1999 745 -1961
rect -745 -2027 -740 -1999
rect -712 -2027 -674 -1999
rect -646 -2027 -608 -1999
rect -580 -2027 -542 -1999
rect -514 -2027 -476 -1999
rect -448 -2027 -410 -1999
rect -382 -2027 -344 -1999
rect -316 -2027 -278 -1999
rect -250 -2027 -212 -1999
rect -184 -2027 -146 -1999
rect -118 -2027 -80 -1999
rect -52 -2027 -14 -1999
rect 14 -2027 52 -1999
rect 80 -2027 118 -1999
rect 146 -2027 184 -1999
rect 212 -2027 250 -1999
rect 278 -2027 316 -1999
rect 344 -2027 382 -1999
rect 410 -2027 448 -1999
rect 476 -2027 514 -1999
rect 542 -2027 580 -1999
rect 608 -2027 646 -1999
rect 674 -2027 712 -1999
rect 740 -2027 745 -1999
rect -745 -2065 745 -2027
rect -745 -2093 -740 -2065
rect -712 -2093 -674 -2065
rect -646 -2093 -608 -2065
rect -580 -2093 -542 -2065
rect -514 -2093 -476 -2065
rect -448 -2093 -410 -2065
rect -382 -2093 -344 -2065
rect -316 -2093 -278 -2065
rect -250 -2093 -212 -2065
rect -184 -2093 -146 -2065
rect -118 -2093 -80 -2065
rect -52 -2093 -14 -2065
rect 14 -2093 52 -2065
rect 80 -2093 118 -2065
rect 146 -2093 184 -2065
rect 212 -2093 250 -2065
rect 278 -2093 316 -2065
rect 344 -2093 382 -2065
rect 410 -2093 448 -2065
rect 476 -2093 514 -2065
rect 542 -2093 580 -2065
rect 608 -2093 646 -2065
rect 674 -2093 712 -2065
rect 740 -2093 745 -2065
rect -745 -2131 745 -2093
rect -745 -2159 -740 -2131
rect -712 -2159 -674 -2131
rect -646 -2159 -608 -2131
rect -580 -2159 -542 -2131
rect -514 -2159 -476 -2131
rect -448 -2159 -410 -2131
rect -382 -2159 -344 -2131
rect -316 -2159 -278 -2131
rect -250 -2159 -212 -2131
rect -184 -2159 -146 -2131
rect -118 -2159 -80 -2131
rect -52 -2159 -14 -2131
rect 14 -2159 52 -2131
rect 80 -2159 118 -2131
rect 146 -2159 184 -2131
rect 212 -2159 250 -2131
rect 278 -2159 316 -2131
rect 344 -2159 382 -2131
rect 410 -2159 448 -2131
rect 476 -2159 514 -2131
rect 542 -2159 580 -2131
rect 608 -2159 646 -2131
rect 674 -2159 712 -2131
rect 740 -2159 745 -2131
rect -745 -2197 745 -2159
rect -745 -2225 -740 -2197
rect -712 -2225 -674 -2197
rect -646 -2225 -608 -2197
rect -580 -2225 -542 -2197
rect -514 -2225 -476 -2197
rect -448 -2225 -410 -2197
rect -382 -2225 -344 -2197
rect -316 -2225 -278 -2197
rect -250 -2225 -212 -2197
rect -184 -2225 -146 -2197
rect -118 -2225 -80 -2197
rect -52 -2225 -14 -2197
rect 14 -2225 52 -2197
rect 80 -2225 118 -2197
rect 146 -2225 184 -2197
rect 212 -2225 250 -2197
rect 278 -2225 316 -2197
rect 344 -2225 382 -2197
rect 410 -2225 448 -2197
rect 476 -2225 514 -2197
rect 542 -2225 580 -2197
rect 608 -2225 646 -2197
rect 674 -2225 712 -2197
rect 740 -2225 745 -2197
rect -745 -2263 745 -2225
rect -745 -2291 -740 -2263
rect -712 -2291 -674 -2263
rect -646 -2291 -608 -2263
rect -580 -2291 -542 -2263
rect -514 -2291 -476 -2263
rect -448 -2291 -410 -2263
rect -382 -2291 -344 -2263
rect -316 -2291 -278 -2263
rect -250 -2291 -212 -2263
rect -184 -2291 -146 -2263
rect -118 -2291 -80 -2263
rect -52 -2291 -14 -2263
rect 14 -2291 52 -2263
rect 80 -2291 118 -2263
rect 146 -2291 184 -2263
rect 212 -2291 250 -2263
rect 278 -2291 316 -2263
rect 344 -2291 382 -2263
rect 410 -2291 448 -2263
rect 476 -2291 514 -2263
rect 542 -2291 580 -2263
rect 608 -2291 646 -2263
rect 674 -2291 712 -2263
rect 740 -2291 745 -2263
rect -745 -2329 745 -2291
rect -745 -2357 -740 -2329
rect -712 -2357 -674 -2329
rect -646 -2357 -608 -2329
rect -580 -2357 -542 -2329
rect -514 -2357 -476 -2329
rect -448 -2357 -410 -2329
rect -382 -2357 -344 -2329
rect -316 -2357 -278 -2329
rect -250 -2357 -212 -2329
rect -184 -2357 -146 -2329
rect -118 -2357 -80 -2329
rect -52 -2357 -14 -2329
rect 14 -2357 52 -2329
rect 80 -2357 118 -2329
rect 146 -2357 184 -2329
rect 212 -2357 250 -2329
rect 278 -2357 316 -2329
rect 344 -2357 382 -2329
rect 410 -2357 448 -2329
rect 476 -2357 514 -2329
rect 542 -2357 580 -2329
rect 608 -2357 646 -2329
rect 674 -2357 712 -2329
rect 740 -2357 745 -2329
rect -745 -2395 745 -2357
rect -745 -2423 -740 -2395
rect -712 -2423 -674 -2395
rect -646 -2423 -608 -2395
rect -580 -2423 -542 -2395
rect -514 -2423 -476 -2395
rect -448 -2423 -410 -2395
rect -382 -2423 -344 -2395
rect -316 -2423 -278 -2395
rect -250 -2423 -212 -2395
rect -184 -2423 -146 -2395
rect -118 -2423 -80 -2395
rect -52 -2423 -14 -2395
rect 14 -2423 52 -2395
rect 80 -2423 118 -2395
rect 146 -2423 184 -2395
rect 212 -2423 250 -2395
rect 278 -2423 316 -2395
rect 344 -2423 382 -2395
rect 410 -2423 448 -2395
rect 476 -2423 514 -2395
rect 542 -2423 580 -2395
rect 608 -2423 646 -2395
rect 674 -2423 712 -2395
rect 740 -2423 745 -2395
rect -745 -2461 745 -2423
rect -745 -2489 -740 -2461
rect -712 -2489 -674 -2461
rect -646 -2489 -608 -2461
rect -580 -2489 -542 -2461
rect -514 -2489 -476 -2461
rect -448 -2489 -410 -2461
rect -382 -2489 -344 -2461
rect -316 -2489 -278 -2461
rect -250 -2489 -212 -2461
rect -184 -2489 -146 -2461
rect -118 -2489 -80 -2461
rect -52 -2489 -14 -2461
rect 14 -2489 52 -2461
rect 80 -2489 118 -2461
rect 146 -2489 184 -2461
rect 212 -2489 250 -2461
rect 278 -2489 316 -2461
rect 344 -2489 382 -2461
rect 410 -2489 448 -2461
rect 476 -2489 514 -2461
rect 542 -2489 580 -2461
rect 608 -2489 646 -2461
rect 674 -2489 712 -2461
rect 740 -2489 745 -2461
rect -745 -2527 745 -2489
rect -745 -2555 -740 -2527
rect -712 -2555 -674 -2527
rect -646 -2555 -608 -2527
rect -580 -2555 -542 -2527
rect -514 -2555 -476 -2527
rect -448 -2555 -410 -2527
rect -382 -2555 -344 -2527
rect -316 -2555 -278 -2527
rect -250 -2555 -212 -2527
rect -184 -2555 -146 -2527
rect -118 -2555 -80 -2527
rect -52 -2555 -14 -2527
rect 14 -2555 52 -2527
rect 80 -2555 118 -2527
rect 146 -2555 184 -2527
rect 212 -2555 250 -2527
rect 278 -2555 316 -2527
rect 344 -2555 382 -2527
rect 410 -2555 448 -2527
rect 476 -2555 514 -2527
rect 542 -2555 580 -2527
rect 608 -2555 646 -2527
rect 674 -2555 712 -2527
rect 740 -2555 745 -2527
rect -745 -2593 745 -2555
rect -745 -2621 -740 -2593
rect -712 -2621 -674 -2593
rect -646 -2621 -608 -2593
rect -580 -2621 -542 -2593
rect -514 -2621 -476 -2593
rect -448 -2621 -410 -2593
rect -382 -2621 -344 -2593
rect -316 -2621 -278 -2593
rect -250 -2621 -212 -2593
rect -184 -2621 -146 -2593
rect -118 -2621 -80 -2593
rect -52 -2621 -14 -2593
rect 14 -2621 52 -2593
rect 80 -2621 118 -2593
rect 146 -2621 184 -2593
rect 212 -2621 250 -2593
rect 278 -2621 316 -2593
rect 344 -2621 382 -2593
rect 410 -2621 448 -2593
rect 476 -2621 514 -2593
rect 542 -2621 580 -2593
rect 608 -2621 646 -2593
rect 674 -2621 712 -2593
rect 740 -2621 745 -2593
rect -745 -2659 745 -2621
rect -745 -2687 -740 -2659
rect -712 -2687 -674 -2659
rect -646 -2687 -608 -2659
rect -580 -2687 -542 -2659
rect -514 -2687 -476 -2659
rect -448 -2687 -410 -2659
rect -382 -2687 -344 -2659
rect -316 -2687 -278 -2659
rect -250 -2687 -212 -2659
rect -184 -2687 -146 -2659
rect -118 -2687 -80 -2659
rect -52 -2687 -14 -2659
rect 14 -2687 52 -2659
rect 80 -2687 118 -2659
rect 146 -2687 184 -2659
rect 212 -2687 250 -2659
rect 278 -2687 316 -2659
rect 344 -2687 382 -2659
rect 410 -2687 448 -2659
rect 476 -2687 514 -2659
rect 542 -2687 580 -2659
rect 608 -2687 646 -2659
rect 674 -2687 712 -2659
rect 740 -2687 745 -2659
rect -745 -2725 745 -2687
rect -745 -2753 -740 -2725
rect -712 -2753 -674 -2725
rect -646 -2753 -608 -2725
rect -580 -2753 -542 -2725
rect -514 -2753 -476 -2725
rect -448 -2753 -410 -2725
rect -382 -2753 -344 -2725
rect -316 -2753 -278 -2725
rect -250 -2753 -212 -2725
rect -184 -2753 -146 -2725
rect -118 -2753 -80 -2725
rect -52 -2753 -14 -2725
rect 14 -2753 52 -2725
rect 80 -2753 118 -2725
rect 146 -2753 184 -2725
rect 212 -2753 250 -2725
rect 278 -2753 316 -2725
rect 344 -2753 382 -2725
rect 410 -2753 448 -2725
rect 476 -2753 514 -2725
rect 542 -2753 580 -2725
rect 608 -2753 646 -2725
rect 674 -2753 712 -2725
rect 740 -2753 745 -2725
rect -745 -2791 745 -2753
rect -745 -2819 -740 -2791
rect -712 -2819 -674 -2791
rect -646 -2819 -608 -2791
rect -580 -2819 -542 -2791
rect -514 -2819 -476 -2791
rect -448 -2819 -410 -2791
rect -382 -2819 -344 -2791
rect -316 -2819 -278 -2791
rect -250 -2819 -212 -2791
rect -184 -2819 -146 -2791
rect -118 -2819 -80 -2791
rect -52 -2819 -14 -2791
rect 14 -2819 52 -2791
rect 80 -2819 118 -2791
rect 146 -2819 184 -2791
rect 212 -2819 250 -2791
rect 278 -2819 316 -2791
rect 344 -2819 382 -2791
rect 410 -2819 448 -2791
rect 476 -2819 514 -2791
rect 542 -2819 580 -2791
rect 608 -2819 646 -2791
rect 674 -2819 712 -2791
rect 740 -2819 745 -2791
rect -745 -2857 745 -2819
rect -745 -2885 -740 -2857
rect -712 -2885 -674 -2857
rect -646 -2885 -608 -2857
rect -580 -2885 -542 -2857
rect -514 -2885 -476 -2857
rect -448 -2885 -410 -2857
rect -382 -2885 -344 -2857
rect -316 -2885 -278 -2857
rect -250 -2885 -212 -2857
rect -184 -2885 -146 -2857
rect -118 -2885 -80 -2857
rect -52 -2885 -14 -2857
rect 14 -2885 52 -2857
rect 80 -2885 118 -2857
rect 146 -2885 184 -2857
rect 212 -2885 250 -2857
rect 278 -2885 316 -2857
rect 344 -2885 382 -2857
rect 410 -2885 448 -2857
rect 476 -2885 514 -2857
rect 542 -2885 580 -2857
rect 608 -2885 646 -2857
rect 674 -2885 712 -2857
rect 740 -2885 745 -2857
rect -745 -2923 745 -2885
rect -745 -2951 -740 -2923
rect -712 -2951 -674 -2923
rect -646 -2951 -608 -2923
rect -580 -2951 -542 -2923
rect -514 -2951 -476 -2923
rect -448 -2951 -410 -2923
rect -382 -2951 -344 -2923
rect -316 -2951 -278 -2923
rect -250 -2951 -212 -2923
rect -184 -2951 -146 -2923
rect -118 -2951 -80 -2923
rect -52 -2951 -14 -2923
rect 14 -2951 52 -2923
rect 80 -2951 118 -2923
rect 146 -2951 184 -2923
rect 212 -2951 250 -2923
rect 278 -2951 316 -2923
rect 344 -2951 382 -2923
rect 410 -2951 448 -2923
rect 476 -2951 514 -2923
rect 542 -2951 580 -2923
rect 608 -2951 646 -2923
rect 674 -2951 712 -2923
rect 740 -2951 745 -2923
rect -745 -2989 745 -2951
rect -745 -3017 -740 -2989
rect -712 -3017 -674 -2989
rect -646 -3017 -608 -2989
rect -580 -3017 -542 -2989
rect -514 -3017 -476 -2989
rect -448 -3017 -410 -2989
rect -382 -3017 -344 -2989
rect -316 -3017 -278 -2989
rect -250 -3017 -212 -2989
rect -184 -3017 -146 -2989
rect -118 -3017 -80 -2989
rect -52 -3017 -14 -2989
rect 14 -3017 52 -2989
rect 80 -3017 118 -2989
rect 146 -3017 184 -2989
rect 212 -3017 250 -2989
rect 278 -3017 316 -2989
rect 344 -3017 382 -2989
rect 410 -3017 448 -2989
rect 476 -3017 514 -2989
rect 542 -3017 580 -2989
rect 608 -3017 646 -2989
rect 674 -3017 712 -2989
rect 740 -3017 745 -2989
rect -745 -3055 745 -3017
rect -745 -3083 -740 -3055
rect -712 -3083 -674 -3055
rect -646 -3083 -608 -3055
rect -580 -3083 -542 -3055
rect -514 -3083 -476 -3055
rect -448 -3083 -410 -3055
rect -382 -3083 -344 -3055
rect -316 -3083 -278 -3055
rect -250 -3083 -212 -3055
rect -184 -3083 -146 -3055
rect -118 -3083 -80 -3055
rect -52 -3083 -14 -3055
rect 14 -3083 52 -3055
rect 80 -3083 118 -3055
rect 146 -3083 184 -3055
rect 212 -3083 250 -3055
rect 278 -3083 316 -3055
rect 344 -3083 382 -3055
rect 410 -3083 448 -3055
rect 476 -3083 514 -3055
rect 542 -3083 580 -3055
rect 608 -3083 646 -3055
rect 674 -3083 712 -3055
rect 740 -3083 745 -3055
rect -745 -3121 745 -3083
rect -745 -3149 -740 -3121
rect -712 -3149 -674 -3121
rect -646 -3149 -608 -3121
rect -580 -3149 -542 -3121
rect -514 -3149 -476 -3121
rect -448 -3149 -410 -3121
rect -382 -3149 -344 -3121
rect -316 -3149 -278 -3121
rect -250 -3149 -212 -3121
rect -184 -3149 -146 -3121
rect -118 -3149 -80 -3121
rect -52 -3149 -14 -3121
rect 14 -3149 52 -3121
rect 80 -3149 118 -3121
rect 146 -3149 184 -3121
rect 212 -3149 250 -3121
rect 278 -3149 316 -3121
rect 344 -3149 382 -3121
rect 410 -3149 448 -3121
rect 476 -3149 514 -3121
rect 542 -3149 580 -3121
rect 608 -3149 646 -3121
rect 674 -3149 712 -3121
rect 740 -3149 745 -3121
rect -745 -3187 745 -3149
rect -745 -3215 -740 -3187
rect -712 -3215 -674 -3187
rect -646 -3215 -608 -3187
rect -580 -3215 -542 -3187
rect -514 -3215 -476 -3187
rect -448 -3215 -410 -3187
rect -382 -3215 -344 -3187
rect -316 -3215 -278 -3187
rect -250 -3215 -212 -3187
rect -184 -3215 -146 -3187
rect -118 -3215 -80 -3187
rect -52 -3215 -14 -3187
rect 14 -3215 52 -3187
rect 80 -3215 118 -3187
rect 146 -3215 184 -3187
rect 212 -3215 250 -3187
rect 278 -3215 316 -3187
rect 344 -3215 382 -3187
rect 410 -3215 448 -3187
rect 476 -3215 514 -3187
rect 542 -3215 580 -3187
rect 608 -3215 646 -3187
rect 674 -3215 712 -3187
rect 740 -3215 745 -3187
rect -745 -3253 745 -3215
rect -745 -3281 -740 -3253
rect -712 -3281 -674 -3253
rect -646 -3281 -608 -3253
rect -580 -3281 -542 -3253
rect -514 -3281 -476 -3253
rect -448 -3281 -410 -3253
rect -382 -3281 -344 -3253
rect -316 -3281 -278 -3253
rect -250 -3281 -212 -3253
rect -184 -3281 -146 -3253
rect -118 -3281 -80 -3253
rect -52 -3281 -14 -3253
rect 14 -3281 52 -3253
rect 80 -3281 118 -3253
rect 146 -3281 184 -3253
rect 212 -3281 250 -3253
rect 278 -3281 316 -3253
rect 344 -3281 382 -3253
rect 410 -3281 448 -3253
rect 476 -3281 514 -3253
rect 542 -3281 580 -3253
rect 608 -3281 646 -3253
rect 674 -3281 712 -3253
rect 740 -3281 745 -3253
rect -745 -3319 745 -3281
rect -745 -3347 -740 -3319
rect -712 -3347 -674 -3319
rect -646 -3347 -608 -3319
rect -580 -3347 -542 -3319
rect -514 -3347 -476 -3319
rect -448 -3347 -410 -3319
rect -382 -3347 -344 -3319
rect -316 -3347 -278 -3319
rect -250 -3347 -212 -3319
rect -184 -3347 -146 -3319
rect -118 -3347 -80 -3319
rect -52 -3347 -14 -3319
rect 14 -3347 52 -3319
rect 80 -3347 118 -3319
rect 146 -3347 184 -3319
rect 212 -3347 250 -3319
rect 278 -3347 316 -3319
rect 344 -3347 382 -3319
rect 410 -3347 448 -3319
rect 476 -3347 514 -3319
rect 542 -3347 580 -3319
rect 608 -3347 646 -3319
rect 674 -3347 712 -3319
rect 740 -3347 745 -3319
rect -745 -3385 745 -3347
rect -745 -3413 -740 -3385
rect -712 -3413 -674 -3385
rect -646 -3413 -608 -3385
rect -580 -3413 -542 -3385
rect -514 -3413 -476 -3385
rect -448 -3413 -410 -3385
rect -382 -3413 -344 -3385
rect -316 -3413 -278 -3385
rect -250 -3413 -212 -3385
rect -184 -3413 -146 -3385
rect -118 -3413 -80 -3385
rect -52 -3413 -14 -3385
rect 14 -3413 52 -3385
rect 80 -3413 118 -3385
rect 146 -3413 184 -3385
rect 212 -3413 250 -3385
rect 278 -3413 316 -3385
rect 344 -3413 382 -3385
rect 410 -3413 448 -3385
rect 476 -3413 514 -3385
rect 542 -3413 580 -3385
rect 608 -3413 646 -3385
rect 674 -3413 712 -3385
rect 740 -3413 745 -3385
rect -745 -3451 745 -3413
rect -745 -3479 -740 -3451
rect -712 -3479 -674 -3451
rect -646 -3479 -608 -3451
rect -580 -3479 -542 -3451
rect -514 -3479 -476 -3451
rect -448 -3479 -410 -3451
rect -382 -3479 -344 -3451
rect -316 -3479 -278 -3451
rect -250 -3479 -212 -3451
rect -184 -3479 -146 -3451
rect -118 -3479 -80 -3451
rect -52 -3479 -14 -3451
rect 14 -3479 52 -3451
rect 80 -3479 118 -3451
rect 146 -3479 184 -3451
rect 212 -3479 250 -3451
rect 278 -3479 316 -3451
rect 344 -3479 382 -3451
rect 410 -3479 448 -3451
rect 476 -3479 514 -3451
rect 542 -3479 580 -3451
rect 608 -3479 646 -3451
rect 674 -3479 712 -3451
rect 740 -3479 745 -3451
rect -745 -3517 745 -3479
rect -745 -3545 -740 -3517
rect -712 -3545 -674 -3517
rect -646 -3545 -608 -3517
rect -580 -3545 -542 -3517
rect -514 -3545 -476 -3517
rect -448 -3545 -410 -3517
rect -382 -3545 -344 -3517
rect -316 -3545 -278 -3517
rect -250 -3545 -212 -3517
rect -184 -3545 -146 -3517
rect -118 -3545 -80 -3517
rect -52 -3545 -14 -3517
rect 14 -3545 52 -3517
rect 80 -3545 118 -3517
rect 146 -3545 184 -3517
rect 212 -3545 250 -3517
rect 278 -3545 316 -3517
rect 344 -3545 382 -3517
rect 410 -3545 448 -3517
rect 476 -3545 514 -3517
rect 542 -3545 580 -3517
rect 608 -3545 646 -3517
rect 674 -3545 712 -3517
rect 740 -3545 745 -3517
rect -745 -3583 745 -3545
rect -745 -3611 -740 -3583
rect -712 -3611 -674 -3583
rect -646 -3611 -608 -3583
rect -580 -3611 -542 -3583
rect -514 -3611 -476 -3583
rect -448 -3611 -410 -3583
rect -382 -3611 -344 -3583
rect -316 -3611 -278 -3583
rect -250 -3611 -212 -3583
rect -184 -3611 -146 -3583
rect -118 -3611 -80 -3583
rect -52 -3611 -14 -3583
rect 14 -3611 52 -3583
rect 80 -3611 118 -3583
rect 146 -3611 184 -3583
rect 212 -3611 250 -3583
rect 278 -3611 316 -3583
rect 344 -3611 382 -3583
rect 410 -3611 448 -3583
rect 476 -3611 514 -3583
rect 542 -3611 580 -3583
rect 608 -3611 646 -3583
rect 674 -3611 712 -3583
rect 740 -3611 745 -3583
rect -745 -3649 745 -3611
rect -745 -3677 -740 -3649
rect -712 -3677 -674 -3649
rect -646 -3677 -608 -3649
rect -580 -3677 -542 -3649
rect -514 -3677 -476 -3649
rect -448 -3677 -410 -3649
rect -382 -3677 -344 -3649
rect -316 -3677 -278 -3649
rect -250 -3677 -212 -3649
rect -184 -3677 -146 -3649
rect -118 -3677 -80 -3649
rect -52 -3677 -14 -3649
rect 14 -3677 52 -3649
rect 80 -3677 118 -3649
rect 146 -3677 184 -3649
rect 212 -3677 250 -3649
rect 278 -3677 316 -3649
rect 344 -3677 382 -3649
rect 410 -3677 448 -3649
rect 476 -3677 514 -3649
rect 542 -3677 580 -3649
rect 608 -3677 646 -3649
rect 674 -3677 712 -3649
rect 740 -3677 745 -3649
rect -745 -3715 745 -3677
rect -745 -3743 -740 -3715
rect -712 -3743 -674 -3715
rect -646 -3743 -608 -3715
rect -580 -3743 -542 -3715
rect -514 -3743 -476 -3715
rect -448 -3743 -410 -3715
rect -382 -3743 -344 -3715
rect -316 -3743 -278 -3715
rect -250 -3743 -212 -3715
rect -184 -3743 -146 -3715
rect -118 -3743 -80 -3715
rect -52 -3743 -14 -3715
rect 14 -3743 52 -3715
rect 80 -3743 118 -3715
rect 146 -3743 184 -3715
rect 212 -3743 250 -3715
rect 278 -3743 316 -3715
rect 344 -3743 382 -3715
rect 410 -3743 448 -3715
rect 476 -3743 514 -3715
rect 542 -3743 580 -3715
rect 608 -3743 646 -3715
rect 674 -3743 712 -3715
rect 740 -3743 745 -3715
rect -745 -3781 745 -3743
rect -745 -3809 -740 -3781
rect -712 -3809 -674 -3781
rect -646 -3809 -608 -3781
rect -580 -3809 -542 -3781
rect -514 -3809 -476 -3781
rect -448 -3809 -410 -3781
rect -382 -3809 -344 -3781
rect -316 -3809 -278 -3781
rect -250 -3809 -212 -3781
rect -184 -3809 -146 -3781
rect -118 -3809 -80 -3781
rect -52 -3809 -14 -3781
rect 14 -3809 52 -3781
rect 80 -3809 118 -3781
rect 146 -3809 184 -3781
rect 212 -3809 250 -3781
rect 278 -3809 316 -3781
rect 344 -3809 382 -3781
rect 410 -3809 448 -3781
rect 476 -3809 514 -3781
rect 542 -3809 580 -3781
rect 608 -3809 646 -3781
rect 674 -3809 712 -3781
rect 740 -3809 745 -3781
rect -745 -3847 745 -3809
rect -745 -3875 -740 -3847
rect -712 -3875 -674 -3847
rect -646 -3875 -608 -3847
rect -580 -3875 -542 -3847
rect -514 -3875 -476 -3847
rect -448 -3875 -410 -3847
rect -382 -3875 -344 -3847
rect -316 -3875 -278 -3847
rect -250 -3875 -212 -3847
rect -184 -3875 -146 -3847
rect -118 -3875 -80 -3847
rect -52 -3875 -14 -3847
rect 14 -3875 52 -3847
rect 80 -3875 118 -3847
rect 146 -3875 184 -3847
rect 212 -3875 250 -3847
rect 278 -3875 316 -3847
rect 344 -3875 382 -3847
rect 410 -3875 448 -3847
rect 476 -3875 514 -3847
rect 542 -3875 580 -3847
rect 608 -3875 646 -3847
rect 674 -3875 712 -3847
rect 740 -3875 745 -3847
rect -745 -3880 745 -3875
<< end >>
