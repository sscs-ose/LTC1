magic
tech gf180mcuC
magscale 1 10
timestamp 1699967350
<< nwell >>
rect -707 3813 3491 4009
rect -707 1481 -507 3813
rect 104 1481 221 1482
rect 3265 1481 3491 3813
rect -707 1281 3491 1481
<< pwell >>
rect -534 -1300 3084 1134
<< psubdiff >>
rect -484 1067 3034 1084
rect -484 1021 -467 1067
rect -421 1021 -369 1067
rect -323 1021 -271 1067
rect -225 1021 -173 1067
rect -127 1021 -75 1067
rect -29 1021 23 1067
rect 69 1021 121 1067
rect 167 1021 219 1067
rect 265 1021 317 1067
rect 363 1021 415 1067
rect 461 1021 513 1067
rect 559 1021 611 1067
rect 657 1021 709 1067
rect 755 1021 807 1067
rect 853 1021 905 1067
rect 951 1021 1003 1067
rect 1049 1021 1101 1067
rect 1147 1021 1199 1067
rect 1245 1021 1297 1067
rect 1343 1021 1395 1067
rect 1441 1021 1493 1067
rect 1539 1021 1591 1067
rect 1637 1021 1689 1067
rect 1735 1021 1787 1067
rect 1833 1021 1885 1067
rect 1931 1021 1983 1067
rect 2029 1021 2081 1067
rect 2127 1021 2179 1067
rect 2225 1021 2277 1067
rect 2323 1021 2375 1067
rect 2421 1021 2473 1067
rect 2519 1021 2579 1067
rect 2625 1021 2677 1067
rect 2723 1021 2775 1067
rect 2821 1021 2873 1067
rect 2919 1021 2971 1067
rect 3017 1021 3034 1067
rect -484 1004 3034 1021
rect -484 969 -404 1004
rect -484 923 -467 969
rect -421 923 -404 969
rect -484 871 -404 923
rect -484 825 -467 871
rect -421 825 -404 871
rect -484 773 -404 825
rect -484 727 -467 773
rect -421 727 -404 773
rect -484 675 -404 727
rect -484 629 -467 675
rect -421 629 -404 675
rect -484 577 -404 629
rect -484 531 -467 577
rect -421 531 -404 577
rect -484 479 -404 531
rect -484 433 -467 479
rect -421 433 -404 479
rect -484 381 -404 433
rect -484 335 -467 381
rect -421 335 -404 381
rect -484 283 -404 335
rect -484 237 -467 283
rect -421 237 -404 283
rect -484 185 -404 237
rect -484 139 -467 185
rect -421 139 -404 185
rect -484 87 -404 139
rect -484 41 -467 87
rect -421 41 -404 87
rect 2954 969 3034 1004
rect 2954 923 2971 969
rect 3017 923 3034 969
rect 2954 871 3034 923
rect 2954 825 2971 871
rect 3017 825 3034 871
rect 2954 773 3034 825
rect 2954 727 2971 773
rect 3017 727 3034 773
rect 2954 675 3034 727
rect 2954 629 2971 675
rect 3017 629 3034 675
rect 2954 577 3034 629
rect 2954 531 2971 577
rect 3017 531 3034 577
rect 2954 479 3034 531
rect 2954 433 2971 479
rect 3017 433 3034 479
rect 2954 381 3034 433
rect 2954 335 2971 381
rect 3017 335 3034 381
rect 2954 283 3034 335
rect 2954 237 2971 283
rect 3017 237 3034 283
rect 2954 185 3034 237
rect 2954 139 2971 185
rect 3017 139 3034 185
rect 2954 87 3034 139
rect -484 -11 -404 41
rect -484 -57 -467 -11
rect -421 -57 -404 -11
rect -484 -109 -404 -57
rect -484 -155 -467 -109
rect -421 -155 -404 -109
rect 2954 41 2971 87
rect 3017 41 3034 87
rect 2954 -11 3034 41
rect 2954 -57 2971 -11
rect 3017 -57 3034 -11
rect -484 -207 -404 -155
rect -484 -253 -467 -207
rect -421 -253 -404 -207
rect -484 -305 -404 -253
rect 2954 -109 3034 -57
rect 2954 -155 2971 -109
rect 3017 -155 3034 -109
rect 2954 -207 3034 -155
rect -484 -351 -467 -305
rect -421 -351 -404 -305
rect -484 -403 -404 -351
rect -484 -449 -467 -403
rect -421 -449 -404 -403
rect 2954 -253 2971 -207
rect 3017 -253 3034 -207
rect 2954 -305 3034 -253
rect 2954 -351 2971 -305
rect 3017 -351 3034 -305
rect 2954 -403 3034 -351
rect -484 -501 -404 -449
rect -484 -547 -467 -501
rect -421 -547 -404 -501
rect -484 -599 -404 -547
rect -484 -645 -467 -599
rect -421 -645 -404 -599
rect -484 -697 -404 -645
rect -484 -743 -467 -697
rect -421 -743 -404 -697
rect -484 -795 -404 -743
rect -484 -841 -467 -795
rect -421 -841 -404 -795
rect -484 -893 -404 -841
rect -484 -939 -467 -893
rect -421 -939 -404 -893
rect -484 -991 -404 -939
rect -484 -1037 -467 -991
rect -421 -1037 -404 -991
rect -484 -1089 -404 -1037
rect -484 -1135 -467 -1089
rect -421 -1135 -404 -1089
rect -484 -1170 -404 -1135
rect 2954 -449 2971 -403
rect 3017 -449 3034 -403
rect 2954 -501 3034 -449
rect 2954 -547 2971 -501
rect 3017 -547 3034 -501
rect 2954 -599 3034 -547
rect 2954 -645 2971 -599
rect 3017 -645 3034 -599
rect 2954 -697 3034 -645
rect 2954 -743 2971 -697
rect 3017 -743 3034 -697
rect 2954 -795 3034 -743
rect 2954 -841 2971 -795
rect 3017 -841 3034 -795
rect 2954 -893 3034 -841
rect 2954 -939 2971 -893
rect 3017 -939 3034 -893
rect 2954 -991 3034 -939
rect 2954 -1037 2971 -991
rect 3017 -1037 3034 -991
rect 2954 -1089 3034 -1037
rect 2954 -1135 2971 -1089
rect 3017 -1135 3034 -1089
rect 2954 -1170 3034 -1135
rect -484 -1187 3034 -1170
rect -484 -1233 -467 -1187
rect -421 -1233 -369 -1187
rect -323 -1233 -271 -1187
rect -225 -1233 -173 -1187
rect -127 -1233 -75 -1187
rect -29 -1233 23 -1187
rect 69 -1233 121 -1187
rect 167 -1233 219 -1187
rect 265 -1233 317 -1187
rect 363 -1233 415 -1187
rect 461 -1233 513 -1187
rect 559 -1233 611 -1187
rect 657 -1233 709 -1187
rect 755 -1233 807 -1187
rect 853 -1233 905 -1187
rect 951 -1233 1003 -1187
rect 1049 -1233 1101 -1187
rect 1147 -1233 1199 -1187
rect 1245 -1233 1297 -1187
rect 1343 -1233 1395 -1187
rect 1441 -1233 1493 -1187
rect 1539 -1233 1591 -1187
rect 1637 -1233 1689 -1187
rect 1735 -1233 1787 -1187
rect 1833 -1233 1885 -1187
rect 1931 -1233 1983 -1187
rect 2029 -1233 2081 -1187
rect 2127 -1233 2179 -1187
rect 2225 -1233 2277 -1187
rect 2323 -1233 2375 -1187
rect 2421 -1233 2473 -1187
rect 2519 -1233 2579 -1187
rect 2625 -1233 2677 -1187
rect 2723 -1233 2775 -1187
rect 2821 -1233 2873 -1187
rect 2919 -1233 2971 -1187
rect 3017 -1233 3034 -1187
rect -484 -1250 3034 -1233
<< nsubdiff >>
rect -657 3942 3441 3959
rect -657 3896 -640 3942
rect -594 3896 -542 3942
rect -496 3896 -444 3942
rect -398 3896 -346 3942
rect -300 3896 -248 3942
rect -202 3896 -150 3942
rect -104 3896 -52 3942
rect -6 3896 46 3942
rect 92 3896 144 3942
rect 190 3896 242 3942
rect 288 3896 340 3942
rect 386 3896 438 3942
rect 484 3896 536 3942
rect 582 3896 634 3942
rect 680 3896 732 3942
rect 778 3896 830 3942
rect 876 3896 928 3942
rect 974 3896 1026 3942
rect 1072 3896 1124 3942
rect 1170 3896 1222 3942
rect 1268 3896 1320 3942
rect 1366 3896 1418 3942
rect 1464 3896 1516 3942
rect 1562 3896 1614 3942
rect 1660 3896 1712 3942
rect 1758 3896 1810 3942
rect 1856 3896 1908 3942
rect 1954 3896 2006 3942
rect 2052 3896 2104 3942
rect 2150 3896 2202 3942
rect 2248 3896 2300 3942
rect 2346 3896 2398 3942
rect 2444 3896 2496 3942
rect 2542 3896 2594 3942
rect 2640 3896 2692 3942
rect 2738 3896 2790 3942
rect 2836 3896 2888 3942
rect 2934 3896 2986 3942
rect 3032 3896 3084 3942
rect 3130 3896 3182 3942
rect 3228 3896 3280 3942
rect 3326 3896 3378 3942
rect 3424 3896 3441 3942
rect -657 3879 3441 3896
rect -657 3844 -577 3879
rect -657 3798 -640 3844
rect -594 3798 -577 3844
rect 3361 3844 3441 3879
rect -657 3746 -577 3798
rect -657 3700 -640 3746
rect -594 3700 -577 3746
rect 3361 3798 3378 3844
rect 3424 3798 3441 3844
rect 3361 3746 3441 3798
rect -657 3648 -577 3700
rect -657 3602 -640 3648
rect -594 3602 -577 3648
rect -657 3550 -577 3602
rect -657 3504 -640 3550
rect -594 3504 -577 3550
rect -657 3452 -577 3504
rect -657 3406 -640 3452
rect -594 3406 -577 3452
rect -657 3354 -577 3406
rect -657 3308 -640 3354
rect -594 3308 -577 3354
rect -657 3256 -577 3308
rect -657 3210 -640 3256
rect -594 3210 -577 3256
rect -657 3158 -577 3210
rect -657 3112 -640 3158
rect -594 3112 -577 3158
rect -657 3060 -577 3112
rect -657 3014 -640 3060
rect -594 3014 -577 3060
rect -657 2962 -577 3014
rect -657 2916 -640 2962
rect -594 2916 -577 2962
rect -657 2864 -577 2916
rect -657 2818 -640 2864
rect -594 2818 -577 2864
rect -657 2766 -577 2818
rect -657 2720 -640 2766
rect -594 2720 -577 2766
rect -657 2668 -577 2720
rect -657 2622 -640 2668
rect -594 2622 -577 2668
rect -657 2570 -577 2622
rect -657 2524 -640 2570
rect -594 2524 -577 2570
rect -657 2472 -577 2524
rect -657 2426 -640 2472
rect -594 2426 -577 2472
rect -657 2374 -577 2426
rect -657 2328 -640 2374
rect -594 2328 -577 2374
rect -657 2276 -577 2328
rect -657 2230 -640 2276
rect -594 2230 -577 2276
rect -657 2178 -577 2230
rect -657 2132 -640 2178
rect -594 2132 -577 2178
rect -657 2080 -577 2132
rect -657 2034 -640 2080
rect -594 2034 -577 2080
rect -657 1982 -577 2034
rect -657 1936 -640 1982
rect -594 1936 -577 1982
rect -657 1884 -577 1936
rect -657 1838 -640 1884
rect -594 1838 -577 1884
rect -657 1786 -577 1838
rect -657 1740 -640 1786
rect -594 1740 -577 1786
rect -657 1688 -577 1740
rect -657 1642 -640 1688
rect -594 1642 -577 1688
rect -657 1590 -577 1642
rect -657 1544 -640 1590
rect -594 1544 -577 1590
rect 3361 3700 3378 3746
rect 3424 3700 3441 3746
rect 3361 3648 3441 3700
rect 3361 3602 3378 3648
rect 3424 3602 3441 3648
rect 3361 3550 3441 3602
rect 3361 3504 3378 3550
rect 3424 3504 3441 3550
rect 3361 3452 3441 3504
rect 3361 3406 3378 3452
rect 3424 3406 3441 3452
rect 3361 3354 3441 3406
rect 3361 3308 3378 3354
rect 3424 3308 3441 3354
rect 3361 3256 3441 3308
rect 3361 3210 3378 3256
rect 3424 3210 3441 3256
rect 3361 3158 3441 3210
rect 3361 3112 3378 3158
rect 3424 3112 3441 3158
rect 3361 3060 3441 3112
rect 3361 3014 3378 3060
rect 3424 3014 3441 3060
rect 3361 2962 3441 3014
rect 3361 2916 3378 2962
rect 3424 2916 3441 2962
rect 3361 2864 3441 2916
rect 3361 2818 3378 2864
rect 3424 2818 3441 2864
rect 3361 2766 3441 2818
rect 3361 2720 3378 2766
rect 3424 2720 3441 2766
rect 3361 2668 3441 2720
rect 3361 2622 3378 2668
rect 3424 2622 3441 2668
rect 3361 2570 3441 2622
rect 3361 2524 3378 2570
rect 3424 2524 3441 2570
rect 3361 2472 3441 2524
rect 3361 2426 3378 2472
rect 3424 2426 3441 2472
rect 3361 2374 3441 2426
rect 3361 2328 3378 2374
rect 3424 2328 3441 2374
rect 3361 2276 3441 2328
rect 3361 2230 3378 2276
rect 3424 2230 3441 2276
rect 3361 2178 3441 2230
rect 3361 2132 3378 2178
rect 3424 2132 3441 2178
rect 3361 2080 3441 2132
rect 3361 2034 3378 2080
rect 3424 2034 3441 2080
rect 3361 1982 3441 2034
rect 3361 1936 3378 1982
rect 3424 1936 3441 1982
rect 3361 1884 3441 1936
rect 3361 1838 3378 1884
rect 3424 1838 3441 1884
rect 3361 1786 3441 1838
rect 3361 1740 3378 1786
rect 3424 1740 3441 1786
rect 3361 1688 3441 1740
rect 3361 1642 3378 1688
rect 3424 1642 3441 1688
rect 3361 1590 3441 1642
rect -657 1492 -577 1544
rect -657 1446 -640 1492
rect -594 1446 -577 1492
rect 3361 1544 3378 1590
rect 3424 1544 3441 1590
rect 3361 1492 3441 1544
rect -657 1411 -577 1446
rect 3361 1446 3378 1492
rect 3424 1446 3441 1492
rect 3361 1411 3441 1446
rect -657 1394 3441 1411
rect -657 1348 -640 1394
rect -594 1348 -542 1394
rect -496 1348 -444 1394
rect -398 1348 -346 1394
rect -300 1348 -248 1394
rect -202 1348 -150 1394
rect -104 1348 -52 1394
rect -6 1348 46 1394
rect 92 1348 144 1394
rect 190 1348 242 1394
rect 288 1348 340 1394
rect 386 1348 438 1394
rect 484 1348 536 1394
rect 582 1348 634 1394
rect 680 1348 732 1394
rect 778 1348 830 1394
rect 876 1348 928 1394
rect 974 1348 1026 1394
rect 1072 1348 1124 1394
rect 1170 1348 1222 1394
rect 1268 1348 1320 1394
rect 1366 1348 1418 1394
rect 1464 1348 1516 1394
rect 1562 1348 1614 1394
rect 1660 1348 1712 1394
rect 1758 1348 1810 1394
rect 1856 1348 1908 1394
rect 1954 1348 2006 1394
rect 2052 1348 2104 1394
rect 2150 1348 2202 1394
rect 2248 1348 2300 1394
rect 2346 1348 2398 1394
rect 2444 1348 2496 1394
rect 2542 1348 2594 1394
rect 2640 1348 2692 1394
rect 2738 1348 2790 1394
rect 2836 1348 2888 1394
rect 2934 1348 2986 1394
rect 3032 1348 3084 1394
rect 3130 1348 3182 1394
rect 3228 1348 3280 1394
rect 3326 1348 3378 1394
rect 3424 1348 3441 1394
rect -657 1331 3441 1348
<< psubdiffcont >>
rect -467 1021 -421 1067
rect -369 1021 -323 1067
rect -271 1021 -225 1067
rect -173 1021 -127 1067
rect -75 1021 -29 1067
rect 23 1021 69 1067
rect 121 1021 167 1067
rect 219 1021 265 1067
rect 317 1021 363 1067
rect 415 1021 461 1067
rect 513 1021 559 1067
rect 611 1021 657 1067
rect 709 1021 755 1067
rect 807 1021 853 1067
rect 905 1021 951 1067
rect 1003 1021 1049 1067
rect 1101 1021 1147 1067
rect 1199 1021 1245 1067
rect 1297 1021 1343 1067
rect 1395 1021 1441 1067
rect 1493 1021 1539 1067
rect 1591 1021 1637 1067
rect 1689 1021 1735 1067
rect 1787 1021 1833 1067
rect 1885 1021 1931 1067
rect 1983 1021 2029 1067
rect 2081 1021 2127 1067
rect 2179 1021 2225 1067
rect 2277 1021 2323 1067
rect 2375 1021 2421 1067
rect 2473 1021 2519 1067
rect 2579 1021 2625 1067
rect 2677 1021 2723 1067
rect 2775 1021 2821 1067
rect 2873 1021 2919 1067
rect 2971 1021 3017 1067
rect -467 923 -421 969
rect -467 825 -421 871
rect -467 727 -421 773
rect -467 629 -421 675
rect -467 531 -421 577
rect -467 433 -421 479
rect -467 335 -421 381
rect -467 237 -421 283
rect -467 139 -421 185
rect -467 41 -421 87
rect 2971 923 3017 969
rect 2971 825 3017 871
rect 2971 727 3017 773
rect 2971 629 3017 675
rect 2971 531 3017 577
rect 2971 433 3017 479
rect 2971 335 3017 381
rect 2971 237 3017 283
rect 2971 139 3017 185
rect -467 -57 -421 -11
rect -467 -155 -421 -109
rect 2971 41 3017 87
rect 2971 -57 3017 -11
rect -467 -253 -421 -207
rect 2971 -155 3017 -109
rect -467 -351 -421 -305
rect -467 -449 -421 -403
rect 2971 -253 3017 -207
rect 2971 -351 3017 -305
rect -467 -547 -421 -501
rect -467 -645 -421 -599
rect -467 -743 -421 -697
rect -467 -841 -421 -795
rect -467 -939 -421 -893
rect -467 -1037 -421 -991
rect -467 -1135 -421 -1089
rect 2971 -449 3017 -403
rect 2971 -547 3017 -501
rect 2971 -645 3017 -599
rect 2971 -743 3017 -697
rect 2971 -841 3017 -795
rect 2971 -939 3017 -893
rect 2971 -1037 3017 -991
rect 2971 -1135 3017 -1089
rect -467 -1233 -421 -1187
rect -369 -1233 -323 -1187
rect -271 -1233 -225 -1187
rect -173 -1233 -127 -1187
rect -75 -1233 -29 -1187
rect 23 -1233 69 -1187
rect 121 -1233 167 -1187
rect 219 -1233 265 -1187
rect 317 -1233 363 -1187
rect 415 -1233 461 -1187
rect 513 -1233 559 -1187
rect 611 -1233 657 -1187
rect 709 -1233 755 -1187
rect 807 -1233 853 -1187
rect 905 -1233 951 -1187
rect 1003 -1233 1049 -1187
rect 1101 -1233 1147 -1187
rect 1199 -1233 1245 -1187
rect 1297 -1233 1343 -1187
rect 1395 -1233 1441 -1187
rect 1493 -1233 1539 -1187
rect 1591 -1233 1637 -1187
rect 1689 -1233 1735 -1187
rect 1787 -1233 1833 -1187
rect 1885 -1233 1931 -1187
rect 1983 -1233 2029 -1187
rect 2081 -1233 2127 -1187
rect 2179 -1233 2225 -1187
rect 2277 -1233 2323 -1187
rect 2375 -1233 2421 -1187
rect 2473 -1233 2519 -1187
rect 2579 -1233 2625 -1187
rect 2677 -1233 2723 -1187
rect 2775 -1233 2821 -1187
rect 2873 -1233 2919 -1187
rect 2971 -1233 3017 -1187
<< nsubdiffcont >>
rect -640 3896 -594 3942
rect -542 3896 -496 3942
rect -444 3896 -398 3942
rect -346 3896 -300 3942
rect -248 3896 -202 3942
rect -150 3896 -104 3942
rect -52 3896 -6 3942
rect 46 3896 92 3942
rect 144 3896 190 3942
rect 242 3896 288 3942
rect 340 3896 386 3942
rect 438 3896 484 3942
rect 536 3896 582 3942
rect 634 3896 680 3942
rect 732 3896 778 3942
rect 830 3896 876 3942
rect 928 3896 974 3942
rect 1026 3896 1072 3942
rect 1124 3896 1170 3942
rect 1222 3896 1268 3942
rect 1320 3896 1366 3942
rect 1418 3896 1464 3942
rect 1516 3896 1562 3942
rect 1614 3896 1660 3942
rect 1712 3896 1758 3942
rect 1810 3896 1856 3942
rect 1908 3896 1954 3942
rect 2006 3896 2052 3942
rect 2104 3896 2150 3942
rect 2202 3896 2248 3942
rect 2300 3896 2346 3942
rect 2398 3896 2444 3942
rect 2496 3896 2542 3942
rect 2594 3896 2640 3942
rect 2692 3896 2738 3942
rect 2790 3896 2836 3942
rect 2888 3896 2934 3942
rect 2986 3896 3032 3942
rect 3084 3896 3130 3942
rect 3182 3896 3228 3942
rect 3280 3896 3326 3942
rect 3378 3896 3424 3942
rect -640 3798 -594 3844
rect -640 3700 -594 3746
rect 3378 3798 3424 3844
rect -640 3602 -594 3648
rect -640 3504 -594 3550
rect -640 3406 -594 3452
rect -640 3308 -594 3354
rect -640 3210 -594 3256
rect -640 3112 -594 3158
rect -640 3014 -594 3060
rect -640 2916 -594 2962
rect -640 2818 -594 2864
rect -640 2720 -594 2766
rect -640 2622 -594 2668
rect -640 2524 -594 2570
rect -640 2426 -594 2472
rect -640 2328 -594 2374
rect -640 2230 -594 2276
rect -640 2132 -594 2178
rect -640 2034 -594 2080
rect -640 1936 -594 1982
rect -640 1838 -594 1884
rect -640 1740 -594 1786
rect -640 1642 -594 1688
rect -640 1544 -594 1590
rect 3378 3700 3424 3746
rect 3378 3602 3424 3648
rect 3378 3504 3424 3550
rect 3378 3406 3424 3452
rect 3378 3308 3424 3354
rect 3378 3210 3424 3256
rect 3378 3112 3424 3158
rect 3378 3014 3424 3060
rect 3378 2916 3424 2962
rect 3378 2818 3424 2864
rect 3378 2720 3424 2766
rect 3378 2622 3424 2668
rect 3378 2524 3424 2570
rect 3378 2426 3424 2472
rect 3378 2328 3424 2374
rect 3378 2230 3424 2276
rect 3378 2132 3424 2178
rect 3378 2034 3424 2080
rect 3378 1936 3424 1982
rect 3378 1838 3424 1884
rect 3378 1740 3424 1786
rect 3378 1642 3424 1688
rect -640 1446 -594 1492
rect 3378 1544 3424 1590
rect 3378 1446 3424 1492
rect -640 1348 -594 1394
rect -542 1348 -496 1394
rect -444 1348 -398 1394
rect -346 1348 -300 1394
rect -248 1348 -202 1394
rect -150 1348 -104 1394
rect -52 1348 -6 1394
rect 46 1348 92 1394
rect 144 1348 190 1394
rect 242 1348 288 1394
rect 340 1348 386 1394
rect 438 1348 484 1394
rect 536 1348 582 1394
rect 634 1348 680 1394
rect 732 1348 778 1394
rect 830 1348 876 1394
rect 928 1348 974 1394
rect 1026 1348 1072 1394
rect 1124 1348 1170 1394
rect 1222 1348 1268 1394
rect 1320 1348 1366 1394
rect 1418 1348 1464 1394
rect 1516 1348 1562 1394
rect 1614 1348 1660 1394
rect 1712 1348 1758 1394
rect 1810 1348 1856 1394
rect 1908 1348 1954 1394
rect 2006 1348 2052 1394
rect 2104 1348 2150 1394
rect 2202 1348 2248 1394
rect 2300 1348 2346 1394
rect 2398 1348 2444 1394
rect 2496 1348 2542 1394
rect 2594 1348 2640 1394
rect 2692 1348 2738 1394
rect 2790 1348 2836 1394
rect 2888 1348 2934 1394
rect 2986 1348 3032 1394
rect 3084 1348 3130 1394
rect 3182 1348 3228 1394
rect 3280 1348 3326 1394
rect 3378 1348 3424 1394
<< polysilicon >>
rect 215 3795 2551 3809
rect 215 3749 263 3795
rect 309 3749 2551 3795
rect 215 3727 2551 3749
rect -333 3039 -133 3727
rect 215 3040 415 3727
rect 519 3703 719 3727
rect 823 3703 1023 3727
rect 1127 3703 1327 3727
rect 1431 3703 1631 3727
rect 1735 3703 1935 3727
rect 2039 3703 2239 3727
rect 2343 3703 2543 3727
rect 519 3654 718 3703
rect 519 3040 719 3654
rect 823 3040 1023 3654
rect 1127 3040 1327 3654
rect 1431 3040 1631 3654
rect 1735 3040 1935 3654
rect 2039 3040 2239 3654
rect 2343 3040 2543 3654
rect -333 2993 -260 3039
rect -214 2993 -133 3039
rect -333 2304 -133 2993
rect 214 3038 2543 3040
rect 214 2992 296 3038
rect 342 2992 2543 3038
rect 214 2990 2543 2992
rect 215 2305 415 2990
rect 519 2305 719 2990
rect 823 2305 1023 2990
rect 1127 2305 1327 2990
rect 1431 2305 1631 2990
rect 1735 2305 1935 2990
rect 2039 2305 2239 2990
rect 2343 2305 2543 2990
rect -333 2258 -266 2304
rect -220 2258 -133 2304
rect -333 1567 -133 2258
rect 214 2302 2543 2305
rect 214 2256 265 2302
rect 311 2256 2543 2302
rect 214 2255 2543 2256
rect 215 1567 415 2255
rect 519 1567 719 2255
rect 823 1567 1023 2255
rect 1127 1567 1327 2255
rect 1431 1567 1631 2255
rect 1735 1567 1935 2255
rect 2039 1567 2239 2255
rect 2343 1567 2543 2255
rect 2891 3039 3091 3727
rect 2891 2993 2963 3039
rect 3009 2993 3091 3039
rect 2891 2302 3091 2993
rect 2891 2256 2957 2302
rect 3003 2256 3091 2302
rect 2891 1567 3091 2256
rect 207 1550 2543 1567
rect 207 1504 276 1550
rect 322 1504 2543 1550
rect 207 1485 2543 1504
rect -222 40 -178 61
rect -166 40 -122 50
rect -222 -153 -122 40
rect 2455 24 2456 36
rect 2746 31 2790 57
rect 112 6 2456 24
rect 112 -7 2476 6
rect 84 -8 1273 -7
rect 84 -20 453 -8
rect 84 -76 101 -20
rect 157 -64 453 -20
rect 509 -9 1273 -8
rect 509 -64 857 -9
rect 157 -65 857 -64
rect 913 -63 1273 -9
rect 1329 -8 2087 -7
rect 1329 -63 1691 -8
rect 913 -64 1691 -63
rect 1747 -63 2087 -8
rect 2143 -63 2406 -7
rect 2462 -63 2476 -7
rect 1747 -64 2476 -63
rect 913 -65 2476 -64
rect 157 -76 2476 -65
rect 84 -77 2476 -76
rect 84 -78 2455 -77
rect 84 -90 171 -78
rect 840 -79 927 -78
rect 2690 -82 2790 31
rect 2594 -126 2894 -82
rect 2594 -129 2818 -126
rect 2594 -132 2718 -129
rect -323 -197 -23 -153
rect -323 -200 -99 -197
rect -323 -203 -199 -200
rect -323 -249 -296 -203
rect -250 -246 -199 -203
rect -153 -243 -99 -200
rect -53 -243 -23 -197
rect 2594 -178 2621 -132
rect 2667 -175 2718 -132
rect 2764 -172 2818 -129
rect 2864 -172 2894 -126
rect 2764 -175 2894 -172
rect 2667 -178 2894 -175
rect 2594 -226 2894 -178
rect -153 -246 -23 -243
rect -250 -249 -23 -246
rect -323 -297 -23 -249
rect 87 -286 174 -281
rect 427 -286 514 -280
rect 832 -286 919 -281
rect 1654 -286 1741 -283
rect 2057 -286 2144 -283
rect 87 -293 2457 -286
rect 87 -294 444 -293
rect -222 -432 -122 -297
rect 87 -350 104 -294
rect 160 -349 444 -294
rect 500 -294 2457 -293
rect 500 -349 849 -294
rect 160 -350 849 -349
rect 905 -295 2457 -294
rect 905 -296 2477 -295
rect 905 -300 1671 -296
rect 905 -350 1254 -300
rect 87 -356 1254 -350
rect 1310 -352 1671 -300
rect 1727 -352 2074 -296
rect 2130 -308 2477 -296
rect 2130 -352 2407 -308
rect 1310 -356 2407 -352
rect 87 -364 2407 -356
rect 2463 -364 2477 -308
rect 112 -378 2477 -364
rect 112 -388 2457 -378
rect 2690 -432 2790 -226
<< polycontact >>
rect 263 3749 309 3795
rect -260 2993 -214 3039
rect 296 2992 342 3038
rect -266 2258 -220 2304
rect 265 2256 311 2302
rect 2963 2993 3009 3039
rect 2957 2256 3003 2302
rect 276 1504 322 1550
rect 101 -76 157 -20
rect 453 -64 509 -8
rect 857 -65 913 -9
rect 1273 -63 1329 -7
rect 1691 -64 1747 -8
rect 2087 -63 2143 -7
rect 2406 -63 2462 -7
rect -296 -249 -250 -203
rect -199 -246 -153 -200
rect -99 -243 -53 -197
rect 2621 -178 2667 -132
rect 2718 -175 2764 -129
rect 2818 -172 2864 -126
rect 104 -350 160 -294
rect 444 -349 500 -293
rect 849 -350 905 -294
rect 1254 -356 1310 -300
rect 1671 -352 1727 -296
rect 2074 -352 2130 -296
rect 2407 -364 2463 -308
<< metal1 >>
rect -657 3942 3441 3959
rect -657 3896 -640 3942
rect -594 3896 -542 3942
rect -496 3896 -444 3942
rect -398 3896 -346 3942
rect -300 3896 -248 3942
rect -202 3896 -150 3942
rect -104 3896 -52 3942
rect -6 3896 46 3942
rect 92 3896 144 3942
rect 190 3896 242 3942
rect 288 3896 340 3942
rect 386 3896 438 3942
rect 484 3896 536 3942
rect 582 3896 634 3942
rect 680 3896 732 3942
rect 778 3896 830 3942
rect 876 3896 928 3942
rect 974 3896 1026 3942
rect 1072 3896 1124 3942
rect 1170 3896 1222 3942
rect 1268 3896 1320 3942
rect 1366 3896 1418 3942
rect 1464 3896 1516 3942
rect 1562 3896 1614 3942
rect 1660 3896 1712 3942
rect 1758 3896 1810 3942
rect 1856 3896 1908 3942
rect 1954 3896 2006 3942
rect 2052 3896 2104 3942
rect 2150 3896 2202 3942
rect 2248 3896 2300 3942
rect 2346 3896 2398 3942
rect 2444 3896 2496 3942
rect 2542 3896 2594 3942
rect 2640 3896 2692 3942
rect 2738 3896 2790 3942
rect 2836 3896 2888 3942
rect 2934 3896 2986 3942
rect 3032 3896 3084 3942
rect 3130 3896 3182 3942
rect 3228 3896 3280 3942
rect 3326 3896 3378 3942
rect 3424 3896 3441 3942
rect -657 3879 3441 3896
rect -657 3844 -577 3879
rect -657 3798 -640 3844
rect -594 3798 -577 3844
rect -657 3746 -577 3798
rect -657 3700 -640 3746
rect -594 3700 -577 3746
rect -657 3648 -577 3700
rect -657 3602 -640 3648
rect -594 3602 -577 3648
rect -657 3550 -577 3602
rect -657 3504 -640 3550
rect -594 3504 -577 3550
rect -657 3452 -577 3504
rect -657 3406 -640 3452
rect -594 3406 -577 3452
rect -657 3354 -577 3406
rect -657 3308 -640 3354
rect -594 3308 -577 3354
rect -657 3256 -577 3308
rect -657 3210 -640 3256
rect -594 3210 -577 3256
rect -657 3158 -577 3210
rect -657 3112 -640 3158
rect -594 3112 -577 3158
rect -657 3060 -577 3112
rect -657 3014 -640 3060
rect -594 3035 -577 3060
rect -427 3054 -343 3879
rect -120 3054 -36 3879
rect 110 3795 345 3811
rect 110 3749 263 3795
rect 309 3749 345 3795
rect 110 3726 345 3749
rect 110 3671 195 3726
rect -427 3039 -36 3054
rect -427 3035 -260 3039
rect -594 3014 -260 3035
rect -657 2993 -260 3014
rect -214 2993 -36 3039
rect -657 2970 -36 2993
rect -657 2962 -343 2970
rect -657 2916 -640 2962
rect -594 2951 -343 2962
rect -594 2916 -577 2951
rect -657 2864 -577 2916
rect -657 2818 -640 2864
rect -594 2818 -577 2864
rect -657 2766 -577 2818
rect -657 2720 -640 2766
rect -594 2720 -577 2766
rect -657 2668 -577 2720
rect -657 2622 -640 2668
rect -594 2622 -577 2668
rect -657 2570 -577 2622
rect -657 2524 -640 2570
rect -594 2524 -577 2570
rect -657 2472 -577 2524
rect -657 2426 -640 2472
rect -594 2426 -577 2472
rect -657 2374 -577 2426
rect -657 2328 -640 2374
rect -594 2328 -577 2374
rect -657 2319 -577 2328
rect -427 2319 -343 2951
rect -657 2314 -343 2319
rect -120 2314 -36 2970
rect -657 2304 -36 2314
rect -657 2276 -266 2304
rect -657 2230 -640 2276
rect -594 2258 -266 2276
rect -220 2258 -36 2304
rect -594 2235 -36 2258
rect -594 2230 -577 2235
rect -657 2178 -577 2230
rect -657 2132 -640 2178
rect -594 2132 -577 2178
rect -657 2080 -577 2132
rect -657 2034 -640 2080
rect -594 2034 -577 2080
rect -657 1982 -577 2034
rect -657 1936 -640 1982
rect -594 1936 -577 1982
rect -657 1884 -577 1936
rect -657 1838 -640 1884
rect -594 1838 -577 1884
rect -657 1786 -577 1838
rect -657 1740 -640 1786
rect -594 1740 -577 1786
rect -657 1688 -577 1740
rect -657 1642 -640 1688
rect -594 1642 -577 1688
rect -657 1590 -577 1642
rect -657 1544 -640 1590
rect -594 1544 -577 1590
rect -657 1492 -577 1544
rect -657 1446 -640 1492
rect -594 1446 -577 1492
rect -657 1411 -577 1446
rect -427 2230 -36 2235
rect -427 1411 -343 2230
rect -120 1411 -36 2230
rect 92 3663 198 3671
rect 92 3607 110 3663
rect 166 3607 198 3663
rect 92 3553 198 3607
rect 92 3497 110 3553
rect 166 3497 198 3553
rect 92 3443 198 3497
rect 92 3387 110 3443
rect 166 3387 198 3443
rect 92 3333 198 3387
rect 92 3277 110 3333
rect 166 3277 198 3333
rect 92 3223 198 3277
rect 92 3167 110 3223
rect 166 3167 198 3223
rect 92 3113 198 3167
rect 92 3057 110 3113
rect 166 3106 198 3113
rect 168 3065 198 3106
rect 92 3050 112 3057
rect 168 3050 366 3065
rect 92 3038 366 3050
rect 92 2996 296 3038
rect 92 2940 112 2996
rect 168 2992 296 2996
rect 342 2992 366 3038
rect 168 2980 366 2992
rect 168 2940 198 2980
rect 92 2886 198 2940
rect 92 2830 112 2886
rect 168 2830 198 2886
rect 92 2776 198 2830
rect 92 2720 112 2776
rect 168 2720 198 2776
rect 92 2666 198 2720
rect 92 2610 112 2666
rect 168 2610 198 2666
rect 92 2556 198 2610
rect 92 2500 112 2556
rect 168 2500 198 2556
rect 92 2436 198 2500
rect 92 2380 108 2436
rect 164 2380 198 2436
rect 92 2326 198 2380
rect 92 2270 108 2326
rect 164 2322 198 2326
rect 164 2302 357 2322
rect 164 2270 265 2302
rect 92 2256 265 2270
rect 311 2256 357 2302
rect 92 2237 357 2256
rect 92 2216 198 2237
rect 92 2160 108 2216
rect 164 2160 198 2216
rect 92 2106 198 2160
rect 92 2050 108 2106
rect 164 2050 198 2106
rect 92 1996 198 2050
rect 92 1940 108 1996
rect 164 1940 198 1996
rect 92 1886 198 1940
rect 92 1830 108 1886
rect 164 1830 198 1886
rect 92 1778 198 1830
rect 92 1722 111 1778
rect 167 1722 198 1778
rect 92 1668 198 1722
rect 92 1612 111 1668
rect 167 1612 198 1668
rect 92 1567 198 1612
rect 92 1558 368 1567
rect 92 1502 111 1558
rect 167 1550 368 1558
rect 167 1504 276 1550
rect 322 1504 368 1550
rect 167 1502 368 1504
rect 92 1482 368 1502
rect 420 1411 504 3691
rect 719 3603 821 3654
rect 719 3549 735 3603
rect 790 3549 821 3603
rect 719 3495 821 3549
rect 719 3439 735 3495
rect 790 3439 821 3495
rect 719 3385 821 3439
rect 719 3329 735 3385
rect 790 3329 821 3385
rect 719 3275 821 3329
rect 719 3219 735 3275
rect 790 3219 821 3275
rect 719 3165 821 3219
rect 719 3109 735 3165
rect 790 3109 821 3165
rect 719 2961 821 3109
rect 719 2905 738 2961
rect 794 2905 821 2961
rect 719 2851 821 2905
rect 719 2795 738 2851
rect 794 2795 821 2851
rect 719 2741 821 2795
rect 719 2685 738 2741
rect 794 2685 821 2741
rect 719 2631 821 2685
rect 719 2575 738 2631
rect 794 2575 821 2631
rect 719 2521 821 2575
rect 719 2465 738 2521
rect 794 2465 821 2521
rect 719 2411 821 2465
rect 719 2355 738 2411
rect 794 2355 821 2411
rect 719 2224 821 2355
rect 719 2168 743 2224
rect 799 2168 821 2224
rect 719 2114 821 2168
rect 719 2058 743 2114
rect 799 2058 821 2114
rect 719 2004 821 2058
rect 719 1948 743 2004
rect 799 1948 821 2004
rect 719 1894 821 1948
rect 719 1838 743 1894
rect 799 1838 821 1894
rect 719 1784 821 1838
rect 719 1728 743 1784
rect 799 1728 821 1784
rect 719 1674 821 1728
rect 719 1618 743 1674
rect 799 1618 821 1674
rect 719 1597 821 1618
rect 722 1595 810 1597
rect 1031 1411 1112 3654
rect 1327 3615 1429 3667
rect 1327 3561 1350 3615
rect 1405 3561 1429 3615
rect 1327 3507 1429 3561
rect 1327 3451 1350 3507
rect 1405 3451 1429 3507
rect 1327 3397 1429 3451
rect 1327 3341 1350 3397
rect 1405 3341 1429 3397
rect 1327 3287 1429 3341
rect 1327 3231 1350 3287
rect 1405 3231 1429 3287
rect 1327 3177 1429 3231
rect 1327 3121 1350 3177
rect 1405 3121 1429 3177
rect 1327 2962 1429 3121
rect 1327 2906 1342 2962
rect 1398 2906 1429 2962
rect 1327 2852 1429 2906
rect 1327 2796 1342 2852
rect 1398 2796 1429 2852
rect 1327 2742 1429 2796
rect 1327 2686 1342 2742
rect 1398 2686 1429 2742
rect 1327 2632 1429 2686
rect 1327 2576 1342 2632
rect 1398 2576 1429 2632
rect 1327 2522 1429 2576
rect 1327 2466 1342 2522
rect 1398 2466 1429 2522
rect 1327 2412 1429 2466
rect 1327 2356 1342 2412
rect 1398 2356 1429 2412
rect 1327 2221 1429 2356
rect 1327 2165 1345 2221
rect 1401 2165 1429 2221
rect 1327 2111 1429 2165
rect 1327 2055 1345 2111
rect 1401 2055 1429 2111
rect 1327 2001 1429 2055
rect 1327 1945 1345 2001
rect 1401 1945 1429 2001
rect 1327 1891 1429 1945
rect 1327 1835 1345 1891
rect 1401 1835 1429 1891
rect 1327 1781 1429 1835
rect 1327 1725 1345 1781
rect 1401 1725 1429 1781
rect 1327 1671 1429 1725
rect 1327 1615 1345 1671
rect 1401 1615 1429 1671
rect 1327 1610 1429 1615
rect 1642 1411 1723 3654
rect 1935 3627 2037 3667
rect 1935 3573 1955 3627
rect 2010 3573 2037 3627
rect 1935 3519 2037 3573
rect 1935 3463 1955 3519
rect 2010 3463 2037 3519
rect 1935 3409 2037 3463
rect 1935 3353 1955 3409
rect 2010 3353 2037 3409
rect 1935 3299 2037 3353
rect 1935 3243 1955 3299
rect 2010 3243 2037 3299
rect 1935 3189 2037 3243
rect 1935 3133 1955 3189
rect 2010 3133 2037 3189
rect 1935 2963 2037 3133
rect 1935 2907 1956 2963
rect 2012 2907 2037 2963
rect 1935 2853 2037 2907
rect 1935 2797 1956 2853
rect 2012 2797 2037 2853
rect 1935 2743 2037 2797
rect 1935 2687 1956 2743
rect 2012 2687 2037 2743
rect 1935 2633 2037 2687
rect 1935 2577 1956 2633
rect 2012 2577 2037 2633
rect 1935 2523 2037 2577
rect 1935 2467 1956 2523
rect 2012 2467 2037 2523
rect 1935 2413 2037 2467
rect 1935 2357 1956 2413
rect 2012 2357 2037 2413
rect 1935 2231 2037 2357
rect 1935 2175 1953 2231
rect 2009 2175 2037 2231
rect 1935 2121 2037 2175
rect 1935 2065 1953 2121
rect 2009 2065 2037 2121
rect 1935 2011 2037 2065
rect 1935 1955 1953 2011
rect 2009 1955 2037 2011
rect 1935 1901 2037 1955
rect 1935 1845 1953 1901
rect 2009 1845 2037 1901
rect 1935 1791 2037 1845
rect 1935 1735 1953 1791
rect 2009 1735 2037 1791
rect 1935 1681 2037 1735
rect 1935 1625 1953 1681
rect 2009 1625 2037 1681
rect 1935 1610 2037 1625
rect 2250 1411 2331 3654
rect 2543 3624 2645 3668
rect 2543 3570 2566 3624
rect 2621 3570 2645 3624
rect 2543 3516 2645 3570
rect 2543 3460 2566 3516
rect 2621 3460 2645 3516
rect 2543 3406 2645 3460
rect 2543 3350 2566 3406
rect 2621 3350 2645 3406
rect 2543 3296 2645 3350
rect 2543 3240 2566 3296
rect 2621 3240 2645 3296
rect 2543 3186 2645 3240
rect 2543 3130 2566 3186
rect 2621 3130 2645 3186
rect 2543 2960 2645 3130
rect 2543 2904 2560 2960
rect 2616 2904 2645 2960
rect 2543 2850 2645 2904
rect 2543 2794 2560 2850
rect 2616 2794 2645 2850
rect 2543 2740 2645 2794
rect 2543 2684 2560 2740
rect 2616 2684 2645 2740
rect 2543 2630 2645 2684
rect 2543 2574 2560 2630
rect 2616 2574 2645 2630
rect 2543 2520 2645 2574
rect 2543 2464 2560 2520
rect 2616 2464 2645 2520
rect 2543 2410 2645 2464
rect 2543 2354 2560 2410
rect 2616 2354 2645 2410
rect 2543 2223 2645 2354
rect 2543 2167 2567 2223
rect 2623 2167 2645 2223
rect 2543 2113 2645 2167
rect 2543 2057 2567 2113
rect 2623 2057 2645 2113
rect 2543 2003 2645 2057
rect 2543 1947 2567 2003
rect 2623 1947 2645 2003
rect 2543 1893 2645 1947
rect 2543 1837 2567 1893
rect 2623 1837 2645 1893
rect 2543 1783 2645 1837
rect 2543 1727 2567 1783
rect 2623 1727 2645 1783
rect 2543 1673 2645 1727
rect 2543 1617 2567 1673
rect 2623 1617 2645 1673
rect 2543 1611 2645 1617
rect 2795 3057 2879 3879
rect 3108 3057 3192 3879
rect 2795 3051 3192 3057
rect 3361 3844 3441 3879
rect 3361 3798 3378 3844
rect 3424 3798 3441 3844
rect 3361 3746 3441 3798
rect 3361 3700 3378 3746
rect 3424 3700 3441 3746
rect 3361 3648 3441 3700
rect 3361 3602 3378 3648
rect 3424 3602 3441 3648
rect 3361 3550 3441 3602
rect 3361 3504 3378 3550
rect 3424 3504 3441 3550
rect 3361 3452 3441 3504
rect 3361 3406 3378 3452
rect 3424 3406 3441 3452
rect 3361 3354 3441 3406
rect 3361 3308 3378 3354
rect 3424 3308 3441 3354
rect 3361 3256 3441 3308
rect 3361 3210 3378 3256
rect 3424 3210 3441 3256
rect 3361 3158 3441 3210
rect 3361 3112 3378 3158
rect 3424 3112 3441 3158
rect 3361 3060 3441 3112
rect 3361 3051 3378 3060
rect 2795 3039 3378 3051
rect 2795 2993 2963 3039
rect 3009 3014 3378 3039
rect 3424 3051 3441 3060
rect 3424 3014 3449 3051
rect 3009 2993 3449 3014
rect 2795 2973 3449 2993
rect 2795 2325 2879 2973
rect 3108 2967 3449 2973
rect 3108 2325 3192 2967
rect 2795 2302 3192 2325
rect 2795 2256 2957 2302
rect 3003 2296 3192 2302
rect 3361 2962 3441 2967
rect 3361 2916 3378 2962
rect 3424 2916 3441 2962
rect 3361 2864 3441 2916
rect 3361 2818 3378 2864
rect 3424 2818 3441 2864
rect 3361 2766 3441 2818
rect 3361 2720 3378 2766
rect 3424 2720 3441 2766
rect 3361 2668 3441 2720
rect 3361 2622 3378 2668
rect 3424 2622 3441 2668
rect 3361 2570 3441 2622
rect 3361 2524 3378 2570
rect 3424 2524 3441 2570
rect 3361 2472 3441 2524
rect 3361 2426 3378 2472
rect 3424 2426 3441 2472
rect 3361 2374 3441 2426
rect 3361 2328 3378 2374
rect 3424 2328 3441 2374
rect 3361 2296 3441 2328
rect 3003 2276 3441 2296
rect 3003 2256 3378 2276
rect 2795 2241 3378 2256
rect 2795 1411 2879 2241
rect 3108 2230 3378 2241
rect 3424 2230 3441 2276
rect 3108 2212 3441 2230
rect 3108 1411 3192 2212
rect 3361 2178 3441 2212
rect 3361 2132 3378 2178
rect 3424 2132 3441 2178
rect 3361 2080 3441 2132
rect 3361 2034 3378 2080
rect 3424 2034 3441 2080
rect 3361 1982 3441 2034
rect 3361 1936 3378 1982
rect 3424 1936 3441 1982
rect 3361 1884 3441 1936
rect 3361 1838 3378 1884
rect 3424 1838 3441 1884
rect 3361 1786 3441 1838
rect 3361 1740 3378 1786
rect 3424 1740 3441 1786
rect 3361 1688 3441 1740
rect 3361 1642 3378 1688
rect 3424 1642 3441 1688
rect 3361 1590 3441 1642
rect 3361 1544 3378 1590
rect 3424 1544 3441 1590
rect 3361 1492 3441 1544
rect 3361 1446 3378 1492
rect 3424 1446 3441 1492
rect 3361 1411 3441 1446
rect -657 1394 3441 1411
rect -657 1348 -640 1394
rect -594 1348 -542 1394
rect -496 1348 -444 1394
rect -398 1348 -346 1394
rect -300 1348 -248 1394
rect -202 1348 -150 1394
rect -104 1348 -52 1394
rect -6 1348 46 1394
rect 92 1348 144 1394
rect 190 1348 242 1394
rect 288 1348 340 1394
rect 386 1348 438 1394
rect 484 1348 536 1394
rect 582 1348 634 1394
rect 680 1348 732 1394
rect 778 1348 830 1394
rect 876 1348 928 1394
rect 974 1348 1026 1394
rect 1072 1348 1124 1394
rect 1170 1348 1222 1394
rect 1268 1348 1320 1394
rect 1366 1348 1418 1394
rect 1464 1348 1516 1394
rect 1562 1348 1614 1394
rect 1660 1348 1712 1394
rect 1758 1348 1810 1394
rect 1856 1348 1908 1394
rect 1954 1348 2006 1394
rect 2052 1348 2104 1394
rect 2150 1348 2202 1394
rect 2248 1348 2300 1394
rect 2346 1348 2398 1394
rect 2444 1348 2496 1394
rect 2542 1348 2594 1394
rect 2640 1348 2692 1394
rect 2738 1348 2790 1394
rect 2836 1348 2888 1394
rect 2934 1348 2986 1394
rect 3032 1348 3084 1394
rect 3130 1348 3182 1394
rect 3228 1348 3280 1394
rect 3326 1348 3378 1394
rect 3424 1348 3441 1394
rect -657 1331 3441 1348
rect -484 1067 3034 1084
rect -484 1021 -467 1067
rect -421 1021 -369 1067
rect -323 1021 -271 1067
rect -225 1021 -173 1067
rect -127 1021 -75 1067
rect -29 1021 23 1067
rect 69 1021 121 1067
rect 167 1021 219 1067
rect 265 1021 317 1067
rect 363 1021 415 1067
rect 461 1021 513 1067
rect 559 1021 611 1067
rect 657 1021 709 1067
rect 755 1021 807 1067
rect 853 1021 905 1067
rect 951 1021 1003 1067
rect 1049 1021 1101 1067
rect 1147 1021 1199 1067
rect 1245 1021 1297 1067
rect 1343 1021 1395 1067
rect 1441 1021 1493 1067
rect 1539 1021 1591 1067
rect 1637 1021 1689 1067
rect 1735 1021 1787 1067
rect 1833 1021 1885 1067
rect 1931 1021 1983 1067
rect 2029 1021 2081 1067
rect 2127 1021 2179 1067
rect 2225 1021 2277 1067
rect 2323 1021 2375 1067
rect 2421 1021 2473 1067
rect 2519 1021 2579 1067
rect 2625 1021 2677 1067
rect 2723 1021 2775 1067
rect 2821 1021 2873 1067
rect 2919 1021 2971 1067
rect 3017 1021 3034 1067
rect -484 1004 3034 1021
rect -484 969 -404 1004
rect -484 923 -467 969
rect -421 923 -404 969
rect -484 871 -404 923
rect -484 825 -467 871
rect -421 825 -404 871
rect -484 773 -404 825
rect -484 727 -467 773
rect -421 727 -404 773
rect -484 675 -404 727
rect -484 629 -467 675
rect -421 629 -404 675
rect -484 577 -404 629
rect -484 531 -467 577
rect -421 531 -404 577
rect -484 479 -404 531
rect -484 433 -467 479
rect -421 433 -404 479
rect -484 381 -404 433
rect -484 335 -467 381
rect -421 335 -404 381
rect -484 283 -404 335
rect -484 237 -467 283
rect -421 237 -404 283
rect -484 185 -404 237
rect -484 139 -467 185
rect -421 139 -404 185
rect -484 87 -404 139
rect -484 41 -467 87
rect -421 41 -404 87
rect -484 -11 -404 41
rect -484 -57 -467 -11
rect -421 -57 -404 -11
rect -484 -109 -404 -57
rect -484 -155 -467 -109
rect -421 -155 -404 -109
rect -484 -207 -404 -155
rect -484 -253 -467 -207
rect -421 -253 -404 -207
rect -484 -305 -404 -253
rect -484 -351 -467 -305
rect -421 -351 -404 -305
rect -484 -403 -404 -351
rect -484 -449 -467 -403
rect -421 -449 -404 -403
rect -484 -501 -404 -449
rect -484 -547 -467 -501
rect -421 -547 -404 -501
rect -484 -599 -404 -547
rect -484 -645 -467 -599
rect -421 -645 -404 -599
rect -484 -697 -404 -645
rect -484 -743 -467 -697
rect -421 -743 -404 -697
rect -484 -795 -404 -743
rect -484 -841 -467 -795
rect -421 -841 -404 -795
rect -484 -893 -404 -841
rect -484 -939 -467 -893
rect -421 -939 -404 -893
rect -484 -991 -404 -939
rect -484 -1037 -467 -991
rect -421 -1037 -404 -991
rect -484 -1089 -404 -1037
rect -484 -1135 -467 -1089
rect -421 -1135 -404 -1089
rect -484 -1170 -404 -1135
rect -323 -153 -230 1004
rect -116 -153 -23 1004
rect 2469 880 2543 881
rect 28 844 2543 880
rect 28 788 63 844
rect 119 788 173 844
rect 229 788 283 844
rect 339 788 393 844
rect 449 788 503 844
rect 559 788 613 844
rect 669 837 2543 844
rect 669 788 724 837
rect 28 781 724 788
rect 780 781 834 837
rect 890 781 944 837
rect 1000 781 1054 837
rect 1110 781 1164 837
rect 1220 781 1274 837
rect 1330 835 2156 837
rect 1330 781 1404 835
rect 28 779 1404 781
rect 1460 779 1514 835
rect 1570 779 1624 835
rect 1680 779 1734 835
rect 1790 779 1844 835
rect 1900 779 1954 835
rect 2010 781 2156 835
rect 2212 781 2266 837
rect 2322 781 2376 837
rect 2432 781 2543 837
rect 2010 779 2543 781
rect 28 774 2543 779
rect 28 736 2541 774
rect 33 73 101 736
rect 84 -20 171 -7
rect 84 -76 101 -20
rect 157 -76 171 -20
rect 84 -90 171 -76
rect -323 -197 -23 -153
rect -323 -200 -99 -197
rect -323 -203 -199 -200
rect -323 -249 -296 -203
rect -250 -246 -199 -203
rect -153 -243 -99 -200
rect -53 -243 -23 -197
rect -153 -246 -23 -243
rect -250 -249 -23 -246
rect -323 -297 -23 -249
rect 221 -129 304 668
rect 425 70 511 736
rect 436 -8 523 5
rect 436 -64 453 -8
rect 509 -64 523 -8
rect 436 -78 523 -64
rect 626 -129 709 677
rect 831 73 917 736
rect 840 -9 927 4
rect 840 -65 857 -9
rect 913 -65 927 -9
rect 840 -79 927 -65
rect 1037 -129 1120 665
rect 1240 68 1326 736
rect 1256 -7 1343 6
rect 1256 -63 1273 -7
rect 1329 -63 1343 -7
rect 1256 -77 1343 -63
rect 1440 -129 1523 673
rect 1647 64 1733 736
rect 1674 -8 1761 5
rect 1674 -64 1691 -8
rect 1747 -64 1761 -8
rect 1674 -78 1761 -64
rect 1855 -129 1938 671
rect 2060 73 2146 736
rect 2070 -7 2157 6
rect 2070 -63 2087 -7
rect 2143 -63 2157 -7
rect 2070 -77 2157 -63
rect 2254 -129 2328 670
rect 2474 70 2541 736
rect 2389 -7 2476 6
rect 2389 -63 2406 -7
rect 2462 -63 2476 -7
rect 2389 -77 2476 -63
rect 2594 -82 2687 1004
rect 2800 -82 2893 1004
rect 2954 969 3034 1004
rect 2954 923 2971 969
rect 3017 923 3034 969
rect 2954 871 3034 923
rect 2954 825 2971 871
rect 3017 825 3034 871
rect 2954 773 3034 825
rect 2954 727 2971 773
rect 3017 727 3034 773
rect 2954 675 3034 727
rect 2954 629 2971 675
rect 3017 629 3034 675
rect 2954 577 3034 629
rect 2954 531 2971 577
rect 3017 531 3034 577
rect 2954 479 3034 531
rect 2954 433 2971 479
rect 3017 433 3034 479
rect 2954 381 3034 433
rect 2954 335 2971 381
rect 3017 335 3034 381
rect 2954 283 3034 335
rect 2954 237 2971 283
rect 3017 237 3034 283
rect 2954 185 3034 237
rect 2954 139 2971 185
rect 3017 139 3034 185
rect 2954 87 3034 139
rect 2954 41 2971 87
rect 3017 41 3034 87
rect 2954 -11 3034 41
rect 2954 -57 2971 -11
rect 3017 -57 3034 -11
rect 2594 -126 2894 -82
rect 2594 -129 2818 -126
rect 221 -216 2333 -129
rect 2594 -132 2718 -129
rect 2594 -178 2621 -132
rect 2667 -175 2718 -132
rect 2764 -172 2818 -129
rect 2864 -172 2894 -126
rect 2764 -175 2894 -172
rect 2667 -178 2894 -175
rect -323 -1170 -230 -297
rect -116 -1170 -23 -297
rect 87 -294 174 -281
rect 87 -350 104 -294
rect 160 -350 174 -294
rect 87 -364 174 -350
rect 24 -1170 102 -433
rect 221 -1033 304 -216
rect 427 -293 514 -280
rect 427 -349 444 -293
rect 500 -349 514 -293
rect 427 -363 514 -349
rect 427 -1170 505 -437
rect 626 -1024 709 -216
rect 832 -294 919 -281
rect 832 -350 849 -294
rect 905 -350 919 -294
rect 832 -364 919 -350
rect 838 -1170 916 -437
rect 1037 -1036 1120 -216
rect 1237 -300 1324 -287
rect 1237 -356 1254 -300
rect 1310 -356 1324 -300
rect 1237 -370 1324 -356
rect 1250 -1170 1328 -441
rect 1440 -1028 1523 -216
rect 1654 -296 1741 -283
rect 1654 -352 1671 -296
rect 1727 -352 1741 -296
rect 1654 -366 1741 -352
rect 1652 -1170 1730 -441
rect 1855 -1030 1938 -216
rect 2057 -296 2144 -283
rect 2057 -352 2074 -296
rect 2130 -352 2144 -296
rect 2057 -366 2144 -352
rect 2060 -1170 2138 -441
rect 2254 -1030 2328 -216
rect 2594 -226 2894 -178
rect 2954 -109 3034 -57
rect 2954 -155 2971 -109
rect 3017 -155 3034 -109
rect 2954 -207 3034 -155
rect 2390 -308 2477 -295
rect 2390 -364 2407 -308
rect 2463 -364 2477 -308
rect 2390 -378 2477 -364
rect 2462 -1170 2540 -437
rect 2594 -1170 2687 -226
rect 2800 -1170 2893 -226
rect 2954 -253 2971 -207
rect 3017 -253 3034 -207
rect 2954 -305 3034 -253
rect 2954 -351 2971 -305
rect 3017 -351 3034 -305
rect 2954 -403 3034 -351
rect 2954 -449 2971 -403
rect 3017 -449 3034 -403
rect 2954 -501 3034 -449
rect 2954 -547 2971 -501
rect 3017 -547 3034 -501
rect 2954 -599 3034 -547
rect 2954 -645 2971 -599
rect 3017 -645 3034 -599
rect 2954 -697 3034 -645
rect 2954 -743 2971 -697
rect 3017 -743 3034 -697
rect 2954 -795 3034 -743
rect 2954 -841 2971 -795
rect 3017 -841 3034 -795
rect 2954 -893 3034 -841
rect 2954 -939 2971 -893
rect 3017 -939 3034 -893
rect 2954 -991 3034 -939
rect 2954 -1037 2971 -991
rect 3017 -1037 3034 -991
rect 2954 -1089 3034 -1037
rect 2954 -1135 2971 -1089
rect 3017 -1135 3034 -1089
rect 2954 -1170 3034 -1135
rect -484 -1187 3034 -1170
rect -484 -1233 -467 -1187
rect -421 -1233 -369 -1187
rect -323 -1233 -271 -1187
rect -225 -1233 -173 -1187
rect -127 -1233 -75 -1187
rect -29 -1233 23 -1187
rect 69 -1233 121 -1187
rect 167 -1233 219 -1187
rect 265 -1233 317 -1187
rect 363 -1233 415 -1187
rect 461 -1233 513 -1187
rect 559 -1233 611 -1187
rect 657 -1233 709 -1187
rect 755 -1233 807 -1187
rect 853 -1233 905 -1187
rect 951 -1233 1003 -1187
rect 1049 -1233 1101 -1187
rect 1147 -1233 1199 -1187
rect 1245 -1233 1297 -1187
rect 1343 -1233 1395 -1187
rect 1441 -1233 1493 -1187
rect 1539 -1233 1591 -1187
rect 1637 -1233 1689 -1187
rect 1735 -1233 1787 -1187
rect 1833 -1233 1885 -1187
rect 1931 -1233 1983 -1187
rect 2029 -1233 2081 -1187
rect 2127 -1233 2179 -1187
rect 2225 -1233 2277 -1187
rect 2323 -1233 2375 -1187
rect 2421 -1233 2473 -1187
rect 2519 -1233 2579 -1187
rect 2625 -1233 2677 -1187
rect 2723 -1233 2775 -1187
rect 2821 -1233 2873 -1187
rect 2919 -1233 2971 -1187
rect 3017 -1233 3034 -1187
rect -484 -1250 3034 -1233
<< via1 >>
rect 110 3607 166 3663
rect 110 3497 166 3553
rect 110 3387 166 3443
rect 110 3277 166 3333
rect 110 3167 166 3223
rect 110 3106 166 3113
rect 110 3057 168 3106
rect 112 3050 168 3057
rect 112 2940 168 2996
rect 112 2830 168 2886
rect 112 2720 168 2776
rect 112 2610 168 2666
rect 112 2500 168 2556
rect 108 2380 164 2436
rect 108 2270 164 2326
rect 108 2160 164 2216
rect 108 2050 164 2106
rect 108 1940 164 1996
rect 108 1830 164 1886
rect 111 1722 167 1778
rect 111 1612 167 1668
rect 111 1502 167 1558
rect 735 3549 790 3603
rect 735 3439 790 3495
rect 735 3329 790 3385
rect 735 3219 790 3275
rect 735 3109 790 3165
rect 738 2905 794 2961
rect 738 2795 794 2851
rect 738 2685 794 2741
rect 738 2575 794 2631
rect 738 2465 794 2521
rect 738 2355 794 2411
rect 743 2168 799 2224
rect 743 2058 799 2114
rect 743 1948 799 2004
rect 743 1838 799 1894
rect 743 1728 799 1784
rect 743 1618 799 1674
rect 1350 3561 1405 3615
rect 1350 3451 1405 3507
rect 1350 3341 1405 3397
rect 1350 3231 1405 3287
rect 1350 3121 1405 3177
rect 1342 2906 1398 2962
rect 1342 2796 1398 2852
rect 1342 2686 1398 2742
rect 1342 2576 1398 2632
rect 1342 2466 1398 2522
rect 1342 2356 1398 2412
rect 1345 2165 1401 2221
rect 1345 2055 1401 2111
rect 1345 1945 1401 2001
rect 1345 1835 1401 1891
rect 1345 1725 1401 1781
rect 1345 1615 1401 1671
rect 1955 3573 2010 3627
rect 1955 3463 2010 3519
rect 1955 3353 2010 3409
rect 1955 3243 2010 3299
rect 1955 3133 2010 3189
rect 1956 2907 2012 2963
rect 1956 2797 2012 2853
rect 1956 2687 2012 2743
rect 1956 2577 2012 2633
rect 1956 2467 2012 2523
rect 1956 2357 2012 2413
rect 1953 2175 2009 2231
rect 1953 2065 2009 2121
rect 1953 1955 2009 2011
rect 1953 1845 2009 1901
rect 1953 1735 2009 1791
rect 1953 1625 2009 1681
rect 2566 3570 2621 3624
rect 2566 3460 2621 3516
rect 2566 3350 2621 3406
rect 2566 3240 2621 3296
rect 2566 3130 2621 3186
rect 2560 2904 2616 2960
rect 2560 2794 2616 2850
rect 2560 2684 2616 2740
rect 2560 2574 2616 2630
rect 2560 2464 2616 2520
rect 2560 2354 2616 2410
rect 2567 2167 2623 2223
rect 2567 2057 2623 2113
rect 2567 1947 2623 2003
rect 2567 1837 2623 1893
rect 2567 1727 2623 1783
rect 2567 1617 2623 1673
rect 63 788 119 844
rect 173 788 229 844
rect 283 788 339 844
rect 393 788 449 844
rect 503 788 559 844
rect 613 788 669 844
rect 724 781 780 837
rect 834 781 890 837
rect 944 781 1000 837
rect 1054 781 1110 837
rect 1164 781 1220 837
rect 1274 781 1330 837
rect 1404 779 1460 835
rect 1514 779 1570 835
rect 1624 779 1680 835
rect 1734 779 1790 835
rect 1844 779 1900 835
rect 1954 779 2010 835
rect 2156 781 2212 837
rect 2266 781 2322 837
rect 2376 781 2432 837
rect 101 -76 157 -20
rect 453 -64 509 -8
rect 857 -65 913 -9
rect 1273 -63 1329 -7
rect 1691 -64 1747 -8
rect 2087 -63 2143 -7
rect 2406 -63 2462 -7
rect 104 -350 160 -294
rect 444 -349 500 -293
rect 849 -350 905 -294
rect 1254 -356 1310 -300
rect 1671 -352 1727 -296
rect 2074 -352 2130 -296
rect 2407 -364 2463 -308
<< metal2 >>
rect 713 3790 2638 3914
rect 713 3725 2645 3790
rect 29 3663 199 3678
rect 29 3607 110 3663
rect 166 3607 199 3663
rect 29 3553 199 3607
rect 29 3497 110 3553
rect 166 3497 199 3553
rect 29 3443 199 3497
rect 29 3387 110 3443
rect 166 3387 199 3443
rect 29 3333 199 3387
rect 29 3277 110 3333
rect 166 3277 199 3333
rect 29 3223 199 3277
rect 29 3167 110 3223
rect 166 3167 199 3223
rect 29 3113 199 3167
rect 29 3057 110 3113
rect 166 3106 199 3113
rect 29 3050 112 3057
rect 168 3050 199 3106
rect 29 2996 199 3050
rect 29 2940 112 2996
rect 168 2940 199 2996
rect 29 2886 199 2940
rect 29 2830 112 2886
rect 168 2830 199 2886
rect 29 2776 199 2830
rect 29 2720 112 2776
rect 168 2720 199 2776
rect 29 2666 199 2720
rect 29 2610 112 2666
rect 168 2610 199 2666
rect 29 2556 199 2610
rect 29 2500 112 2556
rect 168 2500 199 2556
rect 29 2436 199 2500
rect 29 2380 108 2436
rect 164 2380 199 2436
rect 29 2326 199 2380
rect 29 2270 108 2326
rect 164 2270 199 2326
rect 29 2216 199 2270
rect 29 2160 108 2216
rect 164 2160 199 2216
rect 29 2106 199 2160
rect 29 2050 108 2106
rect 164 2050 199 2106
rect 29 1996 199 2050
rect 29 1940 108 1996
rect 164 1940 199 1996
rect 29 1886 199 1940
rect 29 1830 108 1886
rect 164 1830 199 1886
rect 29 1807 199 1830
rect 719 3603 821 3725
rect 719 3549 735 3603
rect 790 3549 821 3603
rect 719 3495 821 3549
rect 719 3439 735 3495
rect 790 3439 821 3495
rect 719 3385 821 3439
rect 719 3329 735 3385
rect 790 3329 821 3385
rect 719 3275 821 3329
rect 719 3219 735 3275
rect 790 3219 821 3275
rect 719 3165 821 3219
rect 719 3109 735 3165
rect 790 3109 821 3165
rect 719 2961 821 3109
rect 719 2905 738 2961
rect 794 2905 821 2961
rect 719 2851 821 2905
rect 719 2795 738 2851
rect 794 2795 821 2851
rect 719 2741 821 2795
rect 719 2685 738 2741
rect 794 2685 821 2741
rect 719 2631 821 2685
rect 719 2575 738 2631
rect 794 2575 821 2631
rect 719 2521 821 2575
rect 719 2465 738 2521
rect 794 2465 821 2521
rect 719 2411 821 2465
rect 719 2355 738 2411
rect 794 2355 821 2411
rect 719 2224 821 2355
rect 719 2168 743 2224
rect 799 2168 821 2224
rect 719 2114 821 2168
rect 719 2058 743 2114
rect 799 2058 821 2114
rect 719 2004 821 2058
rect 719 1948 743 2004
rect 799 1948 821 2004
rect 719 1894 821 1948
rect 719 1838 743 1894
rect 799 1838 821 1894
rect 29 1778 218 1807
rect 29 1722 111 1778
rect 167 1722 218 1778
rect 29 1668 218 1722
rect 29 1612 111 1668
rect 167 1612 218 1668
rect 29 1558 218 1612
rect 719 1784 821 1838
rect 719 1728 743 1784
rect 799 1728 821 1784
rect 719 1674 821 1728
rect 719 1618 743 1674
rect 799 1618 821 1674
rect 719 1597 821 1618
rect 1327 3615 1429 3725
rect 1327 3561 1350 3615
rect 1405 3561 1429 3615
rect 1327 3507 1429 3561
rect 1327 3451 1350 3507
rect 1405 3451 1429 3507
rect 1327 3397 1429 3451
rect 1327 3341 1350 3397
rect 1405 3341 1429 3397
rect 1327 3287 1429 3341
rect 1327 3231 1350 3287
rect 1405 3231 1429 3287
rect 1327 3177 1429 3231
rect 1327 3121 1350 3177
rect 1405 3121 1429 3177
rect 1327 2962 1429 3121
rect 1327 2906 1342 2962
rect 1398 2906 1429 2962
rect 1327 2852 1429 2906
rect 1327 2796 1342 2852
rect 1398 2796 1429 2852
rect 1327 2742 1429 2796
rect 1327 2686 1342 2742
rect 1398 2686 1429 2742
rect 1327 2632 1429 2686
rect 1327 2576 1342 2632
rect 1398 2576 1429 2632
rect 1327 2522 1429 2576
rect 1327 2466 1342 2522
rect 1398 2466 1429 2522
rect 1327 2412 1429 2466
rect 1327 2356 1342 2412
rect 1398 2356 1429 2412
rect 1327 2221 1429 2356
rect 1327 2165 1345 2221
rect 1401 2165 1429 2221
rect 1327 2111 1429 2165
rect 1327 2055 1345 2111
rect 1401 2055 1429 2111
rect 1327 2001 1429 2055
rect 1327 1945 1345 2001
rect 1401 1945 1429 2001
rect 1327 1891 1429 1945
rect 1327 1835 1345 1891
rect 1401 1835 1429 1891
rect 1327 1781 1429 1835
rect 1327 1725 1345 1781
rect 1401 1725 1429 1781
rect 1327 1671 1429 1725
rect 1327 1615 1345 1671
rect 1401 1615 1429 1671
rect 1327 1610 1429 1615
rect 1935 3627 2037 3725
rect 1935 3573 1955 3627
rect 2010 3573 2037 3627
rect 1935 3519 2037 3573
rect 1935 3463 1955 3519
rect 2010 3463 2037 3519
rect 1935 3409 2037 3463
rect 1935 3353 1955 3409
rect 2010 3353 2037 3409
rect 1935 3299 2037 3353
rect 1935 3243 1955 3299
rect 2010 3243 2037 3299
rect 1935 3189 2037 3243
rect 1935 3133 1955 3189
rect 2010 3133 2037 3189
rect 1935 2963 2037 3133
rect 1935 2907 1956 2963
rect 2012 2907 2037 2963
rect 1935 2853 2037 2907
rect 1935 2797 1956 2853
rect 2012 2797 2037 2853
rect 1935 2743 2037 2797
rect 1935 2687 1956 2743
rect 2012 2687 2037 2743
rect 1935 2633 2037 2687
rect 1935 2577 1956 2633
rect 2012 2577 2037 2633
rect 1935 2523 2037 2577
rect 1935 2467 1956 2523
rect 2012 2467 2037 2523
rect 1935 2413 2037 2467
rect 1935 2357 1956 2413
rect 2012 2357 2037 2413
rect 1935 2231 2037 2357
rect 1935 2175 1953 2231
rect 2009 2175 2037 2231
rect 1935 2121 2037 2175
rect 1935 2065 1953 2121
rect 2009 2065 2037 2121
rect 1935 2011 2037 2065
rect 1935 1955 1953 2011
rect 2009 1955 2037 2011
rect 1935 1901 2037 1955
rect 1935 1845 1953 1901
rect 2009 1845 2037 1901
rect 1935 1791 2037 1845
rect 1935 1735 1953 1791
rect 2009 1735 2037 1791
rect 1935 1681 2037 1735
rect 1935 1625 1953 1681
rect 2009 1625 2037 1681
rect 1935 1610 2037 1625
rect 2543 3624 2645 3725
rect 2543 3570 2566 3624
rect 2621 3570 2645 3624
rect 2543 3516 2645 3570
rect 2543 3460 2566 3516
rect 2621 3460 2645 3516
rect 2543 3406 2645 3460
rect 2543 3350 2566 3406
rect 2621 3350 2645 3406
rect 2543 3296 2645 3350
rect 2543 3240 2566 3296
rect 2621 3240 2645 3296
rect 2543 3186 2645 3240
rect 2543 3130 2566 3186
rect 2621 3130 2645 3186
rect 2543 2960 2645 3130
rect 2543 2904 2560 2960
rect 2616 2904 2645 2960
rect 2543 2850 2645 2904
rect 2543 2794 2560 2850
rect 2616 2794 2645 2850
rect 2543 2740 2645 2794
rect 2543 2684 2560 2740
rect 2616 2684 2645 2740
rect 2543 2630 2645 2684
rect 2543 2574 2560 2630
rect 2616 2574 2645 2630
rect 2543 2520 2645 2574
rect 2543 2464 2560 2520
rect 2616 2464 2645 2520
rect 2543 2410 2645 2464
rect 2543 2354 2560 2410
rect 2616 2354 2645 2410
rect 2543 2223 2645 2354
rect 2543 2167 2567 2223
rect 2623 2167 2645 2223
rect 2543 2113 2645 2167
rect 2543 2057 2567 2113
rect 2623 2057 2645 2113
rect 2543 2003 2645 2057
rect 2543 1947 2567 2003
rect 2623 1947 2645 2003
rect 2543 1893 2645 1947
rect 2543 1837 2567 1893
rect 2623 1837 2645 1893
rect 2543 1783 2645 1837
rect 2543 1727 2567 1783
rect 2623 1727 2645 1783
rect 2543 1673 2645 1727
rect 2543 1617 2567 1673
rect 2623 1617 2645 1673
rect 2543 1611 2645 1617
rect 29 1502 111 1558
rect 167 1502 218 1558
rect 29 881 218 1502
rect 26 844 2543 881
rect 26 788 63 844
rect 119 788 173 844
rect 229 788 283 844
rect 339 788 393 844
rect 449 788 503 844
rect 559 788 613 844
rect 669 837 2543 844
rect 669 788 724 837
rect 26 781 724 788
rect 780 781 834 837
rect 890 781 944 837
rect 1000 781 1054 837
rect 1110 781 1164 837
rect 1220 781 1274 837
rect 1330 835 2156 837
rect 1330 781 1404 835
rect 26 779 1404 781
rect 1460 779 1514 835
rect 1570 779 1624 835
rect 1680 779 1734 835
rect 1790 779 1844 835
rect 1900 779 1954 835
rect 2010 781 2156 835
rect 2212 781 2266 837
rect 2322 781 2376 837
rect 2432 781 2543 837
rect 2010 779 2543 781
rect 26 738 2543 779
rect -605 6 2453 20
rect -605 -7 2476 6
rect -605 -8 1273 -7
rect -605 -20 453 -8
rect -605 -76 101 -20
rect 157 -64 453 -20
rect 509 -9 1273 -8
rect 509 -64 857 -9
rect 157 -65 857 -64
rect 913 -63 1273 -9
rect 1329 -8 2087 -7
rect 1329 -63 1691 -8
rect 913 -64 1691 -63
rect 1747 -63 2087 -8
rect 2143 -63 2406 -7
rect 2462 -63 2476 -7
rect 1747 -64 2476 -63
rect 913 -65 2476 -64
rect 157 -76 2476 -65
rect -605 -77 2476 -76
rect -605 -99 2453 -77
rect -605 -293 2454 -259
rect -605 -294 444 -293
rect -605 -350 104 -294
rect 160 -349 444 -294
rect 500 -294 2454 -293
rect 500 -349 849 -294
rect 160 -350 849 -349
rect 905 -295 2454 -294
rect 905 -296 2477 -295
rect 905 -300 1671 -296
rect 905 -350 1254 -300
rect -605 -356 1254 -350
rect 1310 -352 1671 -300
rect 1727 -352 2074 -296
rect 2130 -308 2477 -296
rect 2130 -352 2407 -308
rect 1310 -356 2407 -352
rect -605 -364 2407 -356
rect 2463 -364 2477 -308
rect -605 -378 2477 -364
use nfet_03v3_8Z2ENZ  nfet_03v3_8Z2ENZ_0
timestamp 1699956126
transform 1 0 -172 0 1 368
box -162 -368 162 368
use nfet_03v3_8Z2ENZ  nfet_03v3_8Z2ENZ_1
timestamp 1699956126
transform 1 0 2406 0 1 368
box -162 -368 162 368
use nfet_03v3_8Z2ENZ  nfet_03v3_8Z2ENZ_2
timestamp 1699956126
transform 1 0 -172 0 1 -732
box -162 -368 162 368
use nfet_03v3_8Z2ENZ  nfet_03v3_8Z2ENZ_3
timestamp 1699956126
transform 1 0 2740 0 1 368
box -162 -368 162 368
use nfet_03v3_8Z2ENZ  nfet_03v3_8Z2ENZ_4
timestamp 1699956126
transform 1 0 2406 0 1 -732
box -162 -368 162 368
use nfet_03v3_8Z2ENZ  nfet_03v3_8Z2ENZ_5
timestamp 1699956126
transform 1 0 2740 0 1 -732
box -162 -368 162 368
use nfet_03v3_U5DXAV  nfet_03v3_U5DXAV_0
timestamp 1699956126
transform 1 0 1182 0 1 368
box -1182 -368 1182 368
use nfet_03v3_U5DXAV  nfet_03v3_U5DXAV_1
timestamp 1699956126
transform 1 0 1182 0 1 -732
box -1182 -368 1182 368
use pfet_03v3_GKYJHF  pfet_03v3_GKYJHF_0
timestamp 1699963945
transform 1 0 -233 0 1 2647
box -274 -1166 274 1166
use pfet_03v3_GKYJHF  pfet_03v3_GKYJHF_1
timestamp 1699963945
transform 1 0 315 0 1 2647
box -274 -1166 274 1166
use pfet_03v3_GKYJHF  pfet_03v3_GKYJHF_2
timestamp 1699963945
transform 1 0 2991 0 1 2647
box -274 -1166 274 1166
use pfet_03v3_GKYWHF  pfet_03v3_GKYWHF_0
timestamp 1699963945
transform 1 0 1531 0 1 2647
box -1186 -1166 1186 1166
<< labels >>
flabel metal1 13 3915 13 3915 0 FreeSans 800 0 0 0 VDD
port 0 nsew
flabel metal2 952 3828 952 3828 0 FreeSans 800 0 0 0 IOUT
port 2 nsew
flabel metal2 -555 -52 -555 -52 0 FreeSans 800 0 0 0 G_SINK_UP
port 3 nsew
flabel metal2 -590 -331 -590 -331 0 FreeSans 800 0 0 0 G_SINK_DOWN
port 4 nsew
flabel metal1 -116 -1213 -116 -1213 0 FreeSans 800 0 0 0 VSS
port 6 nsew
<< end >>
