magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -5906 -1319 5906 1319
<< metal4 >>
rect -4903 311 4903 316
rect -4903 283 -4898 311
rect -4870 283 -4832 311
rect -4804 283 -4766 311
rect -4738 283 -4700 311
rect -4672 283 -4634 311
rect -4606 283 -4568 311
rect -4540 283 -4502 311
rect -4474 283 -4436 311
rect -4408 283 -4370 311
rect -4342 283 -4304 311
rect -4276 283 -4238 311
rect -4210 283 -4172 311
rect -4144 283 -4106 311
rect -4078 283 -4040 311
rect -4012 283 -3974 311
rect -3946 283 -3908 311
rect -3880 283 -3842 311
rect -3814 283 -3776 311
rect -3748 283 -3710 311
rect -3682 283 -3644 311
rect -3616 283 -3578 311
rect -3550 283 -3512 311
rect -3484 283 -3446 311
rect -3418 283 -3380 311
rect -3352 283 -3314 311
rect -3286 283 -3248 311
rect -3220 283 -3182 311
rect -3154 283 -3116 311
rect -3088 283 -3050 311
rect -3022 283 -2984 311
rect -2956 283 -2918 311
rect -2890 283 -2852 311
rect -2824 283 -2786 311
rect -2758 283 -2720 311
rect -2692 283 -2654 311
rect -2626 283 -2588 311
rect -2560 283 -2522 311
rect -2494 283 -2456 311
rect -2428 283 -2390 311
rect -2362 283 -2324 311
rect -2296 283 -2258 311
rect -2230 283 -2192 311
rect -2164 283 -2126 311
rect -2098 283 -2060 311
rect -2032 283 -1994 311
rect -1966 283 -1928 311
rect -1900 283 -1862 311
rect -1834 283 -1796 311
rect -1768 283 -1730 311
rect -1702 283 -1664 311
rect -1636 283 -1598 311
rect -1570 283 -1532 311
rect -1504 283 -1466 311
rect -1438 283 -1400 311
rect -1372 283 -1334 311
rect -1306 283 -1268 311
rect -1240 283 -1202 311
rect -1174 283 -1136 311
rect -1108 283 -1070 311
rect -1042 283 -1004 311
rect -976 283 -938 311
rect -910 283 -872 311
rect -844 283 -806 311
rect -778 283 -740 311
rect -712 283 -674 311
rect -646 283 -608 311
rect -580 283 -542 311
rect -514 283 -476 311
rect -448 283 -410 311
rect -382 283 -344 311
rect -316 283 -278 311
rect -250 283 -212 311
rect -184 283 -146 311
rect -118 283 -80 311
rect -52 283 -14 311
rect 14 283 52 311
rect 80 283 118 311
rect 146 283 184 311
rect 212 283 250 311
rect 278 283 316 311
rect 344 283 382 311
rect 410 283 448 311
rect 476 283 514 311
rect 542 283 580 311
rect 608 283 646 311
rect 674 283 712 311
rect 740 283 778 311
rect 806 283 844 311
rect 872 283 910 311
rect 938 283 976 311
rect 1004 283 1042 311
rect 1070 283 1108 311
rect 1136 283 1174 311
rect 1202 283 1240 311
rect 1268 283 1306 311
rect 1334 283 1372 311
rect 1400 283 1438 311
rect 1466 283 1504 311
rect 1532 283 1570 311
rect 1598 283 1636 311
rect 1664 283 1702 311
rect 1730 283 1768 311
rect 1796 283 1834 311
rect 1862 283 1900 311
rect 1928 283 1966 311
rect 1994 283 2032 311
rect 2060 283 2098 311
rect 2126 283 2164 311
rect 2192 283 2230 311
rect 2258 283 2296 311
rect 2324 283 2362 311
rect 2390 283 2428 311
rect 2456 283 2494 311
rect 2522 283 2560 311
rect 2588 283 2626 311
rect 2654 283 2692 311
rect 2720 283 2758 311
rect 2786 283 2824 311
rect 2852 283 2890 311
rect 2918 283 2956 311
rect 2984 283 3022 311
rect 3050 283 3088 311
rect 3116 283 3154 311
rect 3182 283 3220 311
rect 3248 283 3286 311
rect 3314 283 3352 311
rect 3380 283 3418 311
rect 3446 283 3484 311
rect 3512 283 3550 311
rect 3578 283 3616 311
rect 3644 283 3682 311
rect 3710 283 3748 311
rect 3776 283 3814 311
rect 3842 283 3880 311
rect 3908 283 3946 311
rect 3974 283 4012 311
rect 4040 283 4078 311
rect 4106 283 4144 311
rect 4172 283 4210 311
rect 4238 283 4276 311
rect 4304 283 4342 311
rect 4370 283 4408 311
rect 4436 283 4474 311
rect 4502 283 4540 311
rect 4568 283 4606 311
rect 4634 283 4672 311
rect 4700 283 4738 311
rect 4766 283 4804 311
rect 4832 283 4870 311
rect 4898 283 4903 311
rect -4903 245 4903 283
rect -4903 217 -4898 245
rect -4870 217 -4832 245
rect -4804 217 -4766 245
rect -4738 217 -4700 245
rect -4672 217 -4634 245
rect -4606 217 -4568 245
rect -4540 217 -4502 245
rect -4474 217 -4436 245
rect -4408 217 -4370 245
rect -4342 217 -4304 245
rect -4276 217 -4238 245
rect -4210 217 -4172 245
rect -4144 217 -4106 245
rect -4078 217 -4040 245
rect -4012 217 -3974 245
rect -3946 217 -3908 245
rect -3880 217 -3842 245
rect -3814 217 -3776 245
rect -3748 217 -3710 245
rect -3682 217 -3644 245
rect -3616 217 -3578 245
rect -3550 217 -3512 245
rect -3484 217 -3446 245
rect -3418 217 -3380 245
rect -3352 217 -3314 245
rect -3286 217 -3248 245
rect -3220 217 -3182 245
rect -3154 217 -3116 245
rect -3088 217 -3050 245
rect -3022 217 -2984 245
rect -2956 217 -2918 245
rect -2890 217 -2852 245
rect -2824 217 -2786 245
rect -2758 217 -2720 245
rect -2692 217 -2654 245
rect -2626 217 -2588 245
rect -2560 217 -2522 245
rect -2494 217 -2456 245
rect -2428 217 -2390 245
rect -2362 217 -2324 245
rect -2296 217 -2258 245
rect -2230 217 -2192 245
rect -2164 217 -2126 245
rect -2098 217 -2060 245
rect -2032 217 -1994 245
rect -1966 217 -1928 245
rect -1900 217 -1862 245
rect -1834 217 -1796 245
rect -1768 217 -1730 245
rect -1702 217 -1664 245
rect -1636 217 -1598 245
rect -1570 217 -1532 245
rect -1504 217 -1466 245
rect -1438 217 -1400 245
rect -1372 217 -1334 245
rect -1306 217 -1268 245
rect -1240 217 -1202 245
rect -1174 217 -1136 245
rect -1108 217 -1070 245
rect -1042 217 -1004 245
rect -976 217 -938 245
rect -910 217 -872 245
rect -844 217 -806 245
rect -778 217 -740 245
rect -712 217 -674 245
rect -646 217 -608 245
rect -580 217 -542 245
rect -514 217 -476 245
rect -448 217 -410 245
rect -382 217 -344 245
rect -316 217 -278 245
rect -250 217 -212 245
rect -184 217 -146 245
rect -118 217 -80 245
rect -52 217 -14 245
rect 14 217 52 245
rect 80 217 118 245
rect 146 217 184 245
rect 212 217 250 245
rect 278 217 316 245
rect 344 217 382 245
rect 410 217 448 245
rect 476 217 514 245
rect 542 217 580 245
rect 608 217 646 245
rect 674 217 712 245
rect 740 217 778 245
rect 806 217 844 245
rect 872 217 910 245
rect 938 217 976 245
rect 1004 217 1042 245
rect 1070 217 1108 245
rect 1136 217 1174 245
rect 1202 217 1240 245
rect 1268 217 1306 245
rect 1334 217 1372 245
rect 1400 217 1438 245
rect 1466 217 1504 245
rect 1532 217 1570 245
rect 1598 217 1636 245
rect 1664 217 1702 245
rect 1730 217 1768 245
rect 1796 217 1834 245
rect 1862 217 1900 245
rect 1928 217 1966 245
rect 1994 217 2032 245
rect 2060 217 2098 245
rect 2126 217 2164 245
rect 2192 217 2230 245
rect 2258 217 2296 245
rect 2324 217 2362 245
rect 2390 217 2428 245
rect 2456 217 2494 245
rect 2522 217 2560 245
rect 2588 217 2626 245
rect 2654 217 2692 245
rect 2720 217 2758 245
rect 2786 217 2824 245
rect 2852 217 2890 245
rect 2918 217 2956 245
rect 2984 217 3022 245
rect 3050 217 3088 245
rect 3116 217 3154 245
rect 3182 217 3220 245
rect 3248 217 3286 245
rect 3314 217 3352 245
rect 3380 217 3418 245
rect 3446 217 3484 245
rect 3512 217 3550 245
rect 3578 217 3616 245
rect 3644 217 3682 245
rect 3710 217 3748 245
rect 3776 217 3814 245
rect 3842 217 3880 245
rect 3908 217 3946 245
rect 3974 217 4012 245
rect 4040 217 4078 245
rect 4106 217 4144 245
rect 4172 217 4210 245
rect 4238 217 4276 245
rect 4304 217 4342 245
rect 4370 217 4408 245
rect 4436 217 4474 245
rect 4502 217 4540 245
rect 4568 217 4606 245
rect 4634 217 4672 245
rect 4700 217 4738 245
rect 4766 217 4804 245
rect 4832 217 4870 245
rect 4898 217 4903 245
rect -4903 179 4903 217
rect -4903 151 -4898 179
rect -4870 151 -4832 179
rect -4804 151 -4766 179
rect -4738 151 -4700 179
rect -4672 151 -4634 179
rect -4606 151 -4568 179
rect -4540 151 -4502 179
rect -4474 151 -4436 179
rect -4408 151 -4370 179
rect -4342 151 -4304 179
rect -4276 151 -4238 179
rect -4210 151 -4172 179
rect -4144 151 -4106 179
rect -4078 151 -4040 179
rect -4012 151 -3974 179
rect -3946 151 -3908 179
rect -3880 151 -3842 179
rect -3814 151 -3776 179
rect -3748 151 -3710 179
rect -3682 151 -3644 179
rect -3616 151 -3578 179
rect -3550 151 -3512 179
rect -3484 151 -3446 179
rect -3418 151 -3380 179
rect -3352 151 -3314 179
rect -3286 151 -3248 179
rect -3220 151 -3182 179
rect -3154 151 -3116 179
rect -3088 151 -3050 179
rect -3022 151 -2984 179
rect -2956 151 -2918 179
rect -2890 151 -2852 179
rect -2824 151 -2786 179
rect -2758 151 -2720 179
rect -2692 151 -2654 179
rect -2626 151 -2588 179
rect -2560 151 -2522 179
rect -2494 151 -2456 179
rect -2428 151 -2390 179
rect -2362 151 -2324 179
rect -2296 151 -2258 179
rect -2230 151 -2192 179
rect -2164 151 -2126 179
rect -2098 151 -2060 179
rect -2032 151 -1994 179
rect -1966 151 -1928 179
rect -1900 151 -1862 179
rect -1834 151 -1796 179
rect -1768 151 -1730 179
rect -1702 151 -1664 179
rect -1636 151 -1598 179
rect -1570 151 -1532 179
rect -1504 151 -1466 179
rect -1438 151 -1400 179
rect -1372 151 -1334 179
rect -1306 151 -1268 179
rect -1240 151 -1202 179
rect -1174 151 -1136 179
rect -1108 151 -1070 179
rect -1042 151 -1004 179
rect -976 151 -938 179
rect -910 151 -872 179
rect -844 151 -806 179
rect -778 151 -740 179
rect -712 151 -674 179
rect -646 151 -608 179
rect -580 151 -542 179
rect -514 151 -476 179
rect -448 151 -410 179
rect -382 151 -344 179
rect -316 151 -278 179
rect -250 151 -212 179
rect -184 151 -146 179
rect -118 151 -80 179
rect -52 151 -14 179
rect 14 151 52 179
rect 80 151 118 179
rect 146 151 184 179
rect 212 151 250 179
rect 278 151 316 179
rect 344 151 382 179
rect 410 151 448 179
rect 476 151 514 179
rect 542 151 580 179
rect 608 151 646 179
rect 674 151 712 179
rect 740 151 778 179
rect 806 151 844 179
rect 872 151 910 179
rect 938 151 976 179
rect 1004 151 1042 179
rect 1070 151 1108 179
rect 1136 151 1174 179
rect 1202 151 1240 179
rect 1268 151 1306 179
rect 1334 151 1372 179
rect 1400 151 1438 179
rect 1466 151 1504 179
rect 1532 151 1570 179
rect 1598 151 1636 179
rect 1664 151 1702 179
rect 1730 151 1768 179
rect 1796 151 1834 179
rect 1862 151 1900 179
rect 1928 151 1966 179
rect 1994 151 2032 179
rect 2060 151 2098 179
rect 2126 151 2164 179
rect 2192 151 2230 179
rect 2258 151 2296 179
rect 2324 151 2362 179
rect 2390 151 2428 179
rect 2456 151 2494 179
rect 2522 151 2560 179
rect 2588 151 2626 179
rect 2654 151 2692 179
rect 2720 151 2758 179
rect 2786 151 2824 179
rect 2852 151 2890 179
rect 2918 151 2956 179
rect 2984 151 3022 179
rect 3050 151 3088 179
rect 3116 151 3154 179
rect 3182 151 3220 179
rect 3248 151 3286 179
rect 3314 151 3352 179
rect 3380 151 3418 179
rect 3446 151 3484 179
rect 3512 151 3550 179
rect 3578 151 3616 179
rect 3644 151 3682 179
rect 3710 151 3748 179
rect 3776 151 3814 179
rect 3842 151 3880 179
rect 3908 151 3946 179
rect 3974 151 4012 179
rect 4040 151 4078 179
rect 4106 151 4144 179
rect 4172 151 4210 179
rect 4238 151 4276 179
rect 4304 151 4342 179
rect 4370 151 4408 179
rect 4436 151 4474 179
rect 4502 151 4540 179
rect 4568 151 4606 179
rect 4634 151 4672 179
rect 4700 151 4738 179
rect 4766 151 4804 179
rect 4832 151 4870 179
rect 4898 151 4903 179
rect -4903 113 4903 151
rect -4903 85 -4898 113
rect -4870 85 -4832 113
rect -4804 85 -4766 113
rect -4738 85 -4700 113
rect -4672 85 -4634 113
rect -4606 85 -4568 113
rect -4540 85 -4502 113
rect -4474 85 -4436 113
rect -4408 85 -4370 113
rect -4342 85 -4304 113
rect -4276 85 -4238 113
rect -4210 85 -4172 113
rect -4144 85 -4106 113
rect -4078 85 -4040 113
rect -4012 85 -3974 113
rect -3946 85 -3908 113
rect -3880 85 -3842 113
rect -3814 85 -3776 113
rect -3748 85 -3710 113
rect -3682 85 -3644 113
rect -3616 85 -3578 113
rect -3550 85 -3512 113
rect -3484 85 -3446 113
rect -3418 85 -3380 113
rect -3352 85 -3314 113
rect -3286 85 -3248 113
rect -3220 85 -3182 113
rect -3154 85 -3116 113
rect -3088 85 -3050 113
rect -3022 85 -2984 113
rect -2956 85 -2918 113
rect -2890 85 -2852 113
rect -2824 85 -2786 113
rect -2758 85 -2720 113
rect -2692 85 -2654 113
rect -2626 85 -2588 113
rect -2560 85 -2522 113
rect -2494 85 -2456 113
rect -2428 85 -2390 113
rect -2362 85 -2324 113
rect -2296 85 -2258 113
rect -2230 85 -2192 113
rect -2164 85 -2126 113
rect -2098 85 -2060 113
rect -2032 85 -1994 113
rect -1966 85 -1928 113
rect -1900 85 -1862 113
rect -1834 85 -1796 113
rect -1768 85 -1730 113
rect -1702 85 -1664 113
rect -1636 85 -1598 113
rect -1570 85 -1532 113
rect -1504 85 -1466 113
rect -1438 85 -1400 113
rect -1372 85 -1334 113
rect -1306 85 -1268 113
rect -1240 85 -1202 113
rect -1174 85 -1136 113
rect -1108 85 -1070 113
rect -1042 85 -1004 113
rect -976 85 -938 113
rect -910 85 -872 113
rect -844 85 -806 113
rect -778 85 -740 113
rect -712 85 -674 113
rect -646 85 -608 113
rect -580 85 -542 113
rect -514 85 -476 113
rect -448 85 -410 113
rect -382 85 -344 113
rect -316 85 -278 113
rect -250 85 -212 113
rect -184 85 -146 113
rect -118 85 -80 113
rect -52 85 -14 113
rect 14 85 52 113
rect 80 85 118 113
rect 146 85 184 113
rect 212 85 250 113
rect 278 85 316 113
rect 344 85 382 113
rect 410 85 448 113
rect 476 85 514 113
rect 542 85 580 113
rect 608 85 646 113
rect 674 85 712 113
rect 740 85 778 113
rect 806 85 844 113
rect 872 85 910 113
rect 938 85 976 113
rect 1004 85 1042 113
rect 1070 85 1108 113
rect 1136 85 1174 113
rect 1202 85 1240 113
rect 1268 85 1306 113
rect 1334 85 1372 113
rect 1400 85 1438 113
rect 1466 85 1504 113
rect 1532 85 1570 113
rect 1598 85 1636 113
rect 1664 85 1702 113
rect 1730 85 1768 113
rect 1796 85 1834 113
rect 1862 85 1900 113
rect 1928 85 1966 113
rect 1994 85 2032 113
rect 2060 85 2098 113
rect 2126 85 2164 113
rect 2192 85 2230 113
rect 2258 85 2296 113
rect 2324 85 2362 113
rect 2390 85 2428 113
rect 2456 85 2494 113
rect 2522 85 2560 113
rect 2588 85 2626 113
rect 2654 85 2692 113
rect 2720 85 2758 113
rect 2786 85 2824 113
rect 2852 85 2890 113
rect 2918 85 2956 113
rect 2984 85 3022 113
rect 3050 85 3088 113
rect 3116 85 3154 113
rect 3182 85 3220 113
rect 3248 85 3286 113
rect 3314 85 3352 113
rect 3380 85 3418 113
rect 3446 85 3484 113
rect 3512 85 3550 113
rect 3578 85 3616 113
rect 3644 85 3682 113
rect 3710 85 3748 113
rect 3776 85 3814 113
rect 3842 85 3880 113
rect 3908 85 3946 113
rect 3974 85 4012 113
rect 4040 85 4078 113
rect 4106 85 4144 113
rect 4172 85 4210 113
rect 4238 85 4276 113
rect 4304 85 4342 113
rect 4370 85 4408 113
rect 4436 85 4474 113
rect 4502 85 4540 113
rect 4568 85 4606 113
rect 4634 85 4672 113
rect 4700 85 4738 113
rect 4766 85 4804 113
rect 4832 85 4870 113
rect 4898 85 4903 113
rect -4903 47 4903 85
rect -4903 19 -4898 47
rect -4870 19 -4832 47
rect -4804 19 -4766 47
rect -4738 19 -4700 47
rect -4672 19 -4634 47
rect -4606 19 -4568 47
rect -4540 19 -4502 47
rect -4474 19 -4436 47
rect -4408 19 -4370 47
rect -4342 19 -4304 47
rect -4276 19 -4238 47
rect -4210 19 -4172 47
rect -4144 19 -4106 47
rect -4078 19 -4040 47
rect -4012 19 -3974 47
rect -3946 19 -3908 47
rect -3880 19 -3842 47
rect -3814 19 -3776 47
rect -3748 19 -3710 47
rect -3682 19 -3644 47
rect -3616 19 -3578 47
rect -3550 19 -3512 47
rect -3484 19 -3446 47
rect -3418 19 -3380 47
rect -3352 19 -3314 47
rect -3286 19 -3248 47
rect -3220 19 -3182 47
rect -3154 19 -3116 47
rect -3088 19 -3050 47
rect -3022 19 -2984 47
rect -2956 19 -2918 47
rect -2890 19 -2852 47
rect -2824 19 -2786 47
rect -2758 19 -2720 47
rect -2692 19 -2654 47
rect -2626 19 -2588 47
rect -2560 19 -2522 47
rect -2494 19 -2456 47
rect -2428 19 -2390 47
rect -2362 19 -2324 47
rect -2296 19 -2258 47
rect -2230 19 -2192 47
rect -2164 19 -2126 47
rect -2098 19 -2060 47
rect -2032 19 -1994 47
rect -1966 19 -1928 47
rect -1900 19 -1862 47
rect -1834 19 -1796 47
rect -1768 19 -1730 47
rect -1702 19 -1664 47
rect -1636 19 -1598 47
rect -1570 19 -1532 47
rect -1504 19 -1466 47
rect -1438 19 -1400 47
rect -1372 19 -1334 47
rect -1306 19 -1268 47
rect -1240 19 -1202 47
rect -1174 19 -1136 47
rect -1108 19 -1070 47
rect -1042 19 -1004 47
rect -976 19 -938 47
rect -910 19 -872 47
rect -844 19 -806 47
rect -778 19 -740 47
rect -712 19 -674 47
rect -646 19 -608 47
rect -580 19 -542 47
rect -514 19 -476 47
rect -448 19 -410 47
rect -382 19 -344 47
rect -316 19 -278 47
rect -250 19 -212 47
rect -184 19 -146 47
rect -118 19 -80 47
rect -52 19 -14 47
rect 14 19 52 47
rect 80 19 118 47
rect 146 19 184 47
rect 212 19 250 47
rect 278 19 316 47
rect 344 19 382 47
rect 410 19 448 47
rect 476 19 514 47
rect 542 19 580 47
rect 608 19 646 47
rect 674 19 712 47
rect 740 19 778 47
rect 806 19 844 47
rect 872 19 910 47
rect 938 19 976 47
rect 1004 19 1042 47
rect 1070 19 1108 47
rect 1136 19 1174 47
rect 1202 19 1240 47
rect 1268 19 1306 47
rect 1334 19 1372 47
rect 1400 19 1438 47
rect 1466 19 1504 47
rect 1532 19 1570 47
rect 1598 19 1636 47
rect 1664 19 1702 47
rect 1730 19 1768 47
rect 1796 19 1834 47
rect 1862 19 1900 47
rect 1928 19 1966 47
rect 1994 19 2032 47
rect 2060 19 2098 47
rect 2126 19 2164 47
rect 2192 19 2230 47
rect 2258 19 2296 47
rect 2324 19 2362 47
rect 2390 19 2428 47
rect 2456 19 2494 47
rect 2522 19 2560 47
rect 2588 19 2626 47
rect 2654 19 2692 47
rect 2720 19 2758 47
rect 2786 19 2824 47
rect 2852 19 2890 47
rect 2918 19 2956 47
rect 2984 19 3022 47
rect 3050 19 3088 47
rect 3116 19 3154 47
rect 3182 19 3220 47
rect 3248 19 3286 47
rect 3314 19 3352 47
rect 3380 19 3418 47
rect 3446 19 3484 47
rect 3512 19 3550 47
rect 3578 19 3616 47
rect 3644 19 3682 47
rect 3710 19 3748 47
rect 3776 19 3814 47
rect 3842 19 3880 47
rect 3908 19 3946 47
rect 3974 19 4012 47
rect 4040 19 4078 47
rect 4106 19 4144 47
rect 4172 19 4210 47
rect 4238 19 4276 47
rect 4304 19 4342 47
rect 4370 19 4408 47
rect 4436 19 4474 47
rect 4502 19 4540 47
rect 4568 19 4606 47
rect 4634 19 4672 47
rect 4700 19 4738 47
rect 4766 19 4804 47
rect 4832 19 4870 47
rect 4898 19 4903 47
rect -4903 -19 4903 19
rect -4903 -47 -4898 -19
rect -4870 -47 -4832 -19
rect -4804 -47 -4766 -19
rect -4738 -47 -4700 -19
rect -4672 -47 -4634 -19
rect -4606 -47 -4568 -19
rect -4540 -47 -4502 -19
rect -4474 -47 -4436 -19
rect -4408 -47 -4370 -19
rect -4342 -47 -4304 -19
rect -4276 -47 -4238 -19
rect -4210 -47 -4172 -19
rect -4144 -47 -4106 -19
rect -4078 -47 -4040 -19
rect -4012 -47 -3974 -19
rect -3946 -47 -3908 -19
rect -3880 -47 -3842 -19
rect -3814 -47 -3776 -19
rect -3748 -47 -3710 -19
rect -3682 -47 -3644 -19
rect -3616 -47 -3578 -19
rect -3550 -47 -3512 -19
rect -3484 -47 -3446 -19
rect -3418 -47 -3380 -19
rect -3352 -47 -3314 -19
rect -3286 -47 -3248 -19
rect -3220 -47 -3182 -19
rect -3154 -47 -3116 -19
rect -3088 -47 -3050 -19
rect -3022 -47 -2984 -19
rect -2956 -47 -2918 -19
rect -2890 -47 -2852 -19
rect -2824 -47 -2786 -19
rect -2758 -47 -2720 -19
rect -2692 -47 -2654 -19
rect -2626 -47 -2588 -19
rect -2560 -47 -2522 -19
rect -2494 -47 -2456 -19
rect -2428 -47 -2390 -19
rect -2362 -47 -2324 -19
rect -2296 -47 -2258 -19
rect -2230 -47 -2192 -19
rect -2164 -47 -2126 -19
rect -2098 -47 -2060 -19
rect -2032 -47 -1994 -19
rect -1966 -47 -1928 -19
rect -1900 -47 -1862 -19
rect -1834 -47 -1796 -19
rect -1768 -47 -1730 -19
rect -1702 -47 -1664 -19
rect -1636 -47 -1598 -19
rect -1570 -47 -1532 -19
rect -1504 -47 -1466 -19
rect -1438 -47 -1400 -19
rect -1372 -47 -1334 -19
rect -1306 -47 -1268 -19
rect -1240 -47 -1202 -19
rect -1174 -47 -1136 -19
rect -1108 -47 -1070 -19
rect -1042 -47 -1004 -19
rect -976 -47 -938 -19
rect -910 -47 -872 -19
rect -844 -47 -806 -19
rect -778 -47 -740 -19
rect -712 -47 -674 -19
rect -646 -47 -608 -19
rect -580 -47 -542 -19
rect -514 -47 -476 -19
rect -448 -47 -410 -19
rect -382 -47 -344 -19
rect -316 -47 -278 -19
rect -250 -47 -212 -19
rect -184 -47 -146 -19
rect -118 -47 -80 -19
rect -52 -47 -14 -19
rect 14 -47 52 -19
rect 80 -47 118 -19
rect 146 -47 184 -19
rect 212 -47 250 -19
rect 278 -47 316 -19
rect 344 -47 382 -19
rect 410 -47 448 -19
rect 476 -47 514 -19
rect 542 -47 580 -19
rect 608 -47 646 -19
rect 674 -47 712 -19
rect 740 -47 778 -19
rect 806 -47 844 -19
rect 872 -47 910 -19
rect 938 -47 976 -19
rect 1004 -47 1042 -19
rect 1070 -47 1108 -19
rect 1136 -47 1174 -19
rect 1202 -47 1240 -19
rect 1268 -47 1306 -19
rect 1334 -47 1372 -19
rect 1400 -47 1438 -19
rect 1466 -47 1504 -19
rect 1532 -47 1570 -19
rect 1598 -47 1636 -19
rect 1664 -47 1702 -19
rect 1730 -47 1768 -19
rect 1796 -47 1834 -19
rect 1862 -47 1900 -19
rect 1928 -47 1966 -19
rect 1994 -47 2032 -19
rect 2060 -47 2098 -19
rect 2126 -47 2164 -19
rect 2192 -47 2230 -19
rect 2258 -47 2296 -19
rect 2324 -47 2362 -19
rect 2390 -47 2428 -19
rect 2456 -47 2494 -19
rect 2522 -47 2560 -19
rect 2588 -47 2626 -19
rect 2654 -47 2692 -19
rect 2720 -47 2758 -19
rect 2786 -47 2824 -19
rect 2852 -47 2890 -19
rect 2918 -47 2956 -19
rect 2984 -47 3022 -19
rect 3050 -47 3088 -19
rect 3116 -47 3154 -19
rect 3182 -47 3220 -19
rect 3248 -47 3286 -19
rect 3314 -47 3352 -19
rect 3380 -47 3418 -19
rect 3446 -47 3484 -19
rect 3512 -47 3550 -19
rect 3578 -47 3616 -19
rect 3644 -47 3682 -19
rect 3710 -47 3748 -19
rect 3776 -47 3814 -19
rect 3842 -47 3880 -19
rect 3908 -47 3946 -19
rect 3974 -47 4012 -19
rect 4040 -47 4078 -19
rect 4106 -47 4144 -19
rect 4172 -47 4210 -19
rect 4238 -47 4276 -19
rect 4304 -47 4342 -19
rect 4370 -47 4408 -19
rect 4436 -47 4474 -19
rect 4502 -47 4540 -19
rect 4568 -47 4606 -19
rect 4634 -47 4672 -19
rect 4700 -47 4738 -19
rect 4766 -47 4804 -19
rect 4832 -47 4870 -19
rect 4898 -47 4903 -19
rect -4903 -85 4903 -47
rect -4903 -113 -4898 -85
rect -4870 -113 -4832 -85
rect -4804 -113 -4766 -85
rect -4738 -113 -4700 -85
rect -4672 -113 -4634 -85
rect -4606 -113 -4568 -85
rect -4540 -113 -4502 -85
rect -4474 -113 -4436 -85
rect -4408 -113 -4370 -85
rect -4342 -113 -4304 -85
rect -4276 -113 -4238 -85
rect -4210 -113 -4172 -85
rect -4144 -113 -4106 -85
rect -4078 -113 -4040 -85
rect -4012 -113 -3974 -85
rect -3946 -113 -3908 -85
rect -3880 -113 -3842 -85
rect -3814 -113 -3776 -85
rect -3748 -113 -3710 -85
rect -3682 -113 -3644 -85
rect -3616 -113 -3578 -85
rect -3550 -113 -3512 -85
rect -3484 -113 -3446 -85
rect -3418 -113 -3380 -85
rect -3352 -113 -3314 -85
rect -3286 -113 -3248 -85
rect -3220 -113 -3182 -85
rect -3154 -113 -3116 -85
rect -3088 -113 -3050 -85
rect -3022 -113 -2984 -85
rect -2956 -113 -2918 -85
rect -2890 -113 -2852 -85
rect -2824 -113 -2786 -85
rect -2758 -113 -2720 -85
rect -2692 -113 -2654 -85
rect -2626 -113 -2588 -85
rect -2560 -113 -2522 -85
rect -2494 -113 -2456 -85
rect -2428 -113 -2390 -85
rect -2362 -113 -2324 -85
rect -2296 -113 -2258 -85
rect -2230 -113 -2192 -85
rect -2164 -113 -2126 -85
rect -2098 -113 -2060 -85
rect -2032 -113 -1994 -85
rect -1966 -113 -1928 -85
rect -1900 -113 -1862 -85
rect -1834 -113 -1796 -85
rect -1768 -113 -1730 -85
rect -1702 -113 -1664 -85
rect -1636 -113 -1598 -85
rect -1570 -113 -1532 -85
rect -1504 -113 -1466 -85
rect -1438 -113 -1400 -85
rect -1372 -113 -1334 -85
rect -1306 -113 -1268 -85
rect -1240 -113 -1202 -85
rect -1174 -113 -1136 -85
rect -1108 -113 -1070 -85
rect -1042 -113 -1004 -85
rect -976 -113 -938 -85
rect -910 -113 -872 -85
rect -844 -113 -806 -85
rect -778 -113 -740 -85
rect -712 -113 -674 -85
rect -646 -113 -608 -85
rect -580 -113 -542 -85
rect -514 -113 -476 -85
rect -448 -113 -410 -85
rect -382 -113 -344 -85
rect -316 -113 -278 -85
rect -250 -113 -212 -85
rect -184 -113 -146 -85
rect -118 -113 -80 -85
rect -52 -113 -14 -85
rect 14 -113 52 -85
rect 80 -113 118 -85
rect 146 -113 184 -85
rect 212 -113 250 -85
rect 278 -113 316 -85
rect 344 -113 382 -85
rect 410 -113 448 -85
rect 476 -113 514 -85
rect 542 -113 580 -85
rect 608 -113 646 -85
rect 674 -113 712 -85
rect 740 -113 778 -85
rect 806 -113 844 -85
rect 872 -113 910 -85
rect 938 -113 976 -85
rect 1004 -113 1042 -85
rect 1070 -113 1108 -85
rect 1136 -113 1174 -85
rect 1202 -113 1240 -85
rect 1268 -113 1306 -85
rect 1334 -113 1372 -85
rect 1400 -113 1438 -85
rect 1466 -113 1504 -85
rect 1532 -113 1570 -85
rect 1598 -113 1636 -85
rect 1664 -113 1702 -85
rect 1730 -113 1768 -85
rect 1796 -113 1834 -85
rect 1862 -113 1900 -85
rect 1928 -113 1966 -85
rect 1994 -113 2032 -85
rect 2060 -113 2098 -85
rect 2126 -113 2164 -85
rect 2192 -113 2230 -85
rect 2258 -113 2296 -85
rect 2324 -113 2362 -85
rect 2390 -113 2428 -85
rect 2456 -113 2494 -85
rect 2522 -113 2560 -85
rect 2588 -113 2626 -85
rect 2654 -113 2692 -85
rect 2720 -113 2758 -85
rect 2786 -113 2824 -85
rect 2852 -113 2890 -85
rect 2918 -113 2956 -85
rect 2984 -113 3022 -85
rect 3050 -113 3088 -85
rect 3116 -113 3154 -85
rect 3182 -113 3220 -85
rect 3248 -113 3286 -85
rect 3314 -113 3352 -85
rect 3380 -113 3418 -85
rect 3446 -113 3484 -85
rect 3512 -113 3550 -85
rect 3578 -113 3616 -85
rect 3644 -113 3682 -85
rect 3710 -113 3748 -85
rect 3776 -113 3814 -85
rect 3842 -113 3880 -85
rect 3908 -113 3946 -85
rect 3974 -113 4012 -85
rect 4040 -113 4078 -85
rect 4106 -113 4144 -85
rect 4172 -113 4210 -85
rect 4238 -113 4276 -85
rect 4304 -113 4342 -85
rect 4370 -113 4408 -85
rect 4436 -113 4474 -85
rect 4502 -113 4540 -85
rect 4568 -113 4606 -85
rect 4634 -113 4672 -85
rect 4700 -113 4738 -85
rect 4766 -113 4804 -85
rect 4832 -113 4870 -85
rect 4898 -113 4903 -85
rect -4903 -151 4903 -113
rect -4903 -179 -4898 -151
rect -4870 -179 -4832 -151
rect -4804 -179 -4766 -151
rect -4738 -179 -4700 -151
rect -4672 -179 -4634 -151
rect -4606 -179 -4568 -151
rect -4540 -179 -4502 -151
rect -4474 -179 -4436 -151
rect -4408 -179 -4370 -151
rect -4342 -179 -4304 -151
rect -4276 -179 -4238 -151
rect -4210 -179 -4172 -151
rect -4144 -179 -4106 -151
rect -4078 -179 -4040 -151
rect -4012 -179 -3974 -151
rect -3946 -179 -3908 -151
rect -3880 -179 -3842 -151
rect -3814 -179 -3776 -151
rect -3748 -179 -3710 -151
rect -3682 -179 -3644 -151
rect -3616 -179 -3578 -151
rect -3550 -179 -3512 -151
rect -3484 -179 -3446 -151
rect -3418 -179 -3380 -151
rect -3352 -179 -3314 -151
rect -3286 -179 -3248 -151
rect -3220 -179 -3182 -151
rect -3154 -179 -3116 -151
rect -3088 -179 -3050 -151
rect -3022 -179 -2984 -151
rect -2956 -179 -2918 -151
rect -2890 -179 -2852 -151
rect -2824 -179 -2786 -151
rect -2758 -179 -2720 -151
rect -2692 -179 -2654 -151
rect -2626 -179 -2588 -151
rect -2560 -179 -2522 -151
rect -2494 -179 -2456 -151
rect -2428 -179 -2390 -151
rect -2362 -179 -2324 -151
rect -2296 -179 -2258 -151
rect -2230 -179 -2192 -151
rect -2164 -179 -2126 -151
rect -2098 -179 -2060 -151
rect -2032 -179 -1994 -151
rect -1966 -179 -1928 -151
rect -1900 -179 -1862 -151
rect -1834 -179 -1796 -151
rect -1768 -179 -1730 -151
rect -1702 -179 -1664 -151
rect -1636 -179 -1598 -151
rect -1570 -179 -1532 -151
rect -1504 -179 -1466 -151
rect -1438 -179 -1400 -151
rect -1372 -179 -1334 -151
rect -1306 -179 -1268 -151
rect -1240 -179 -1202 -151
rect -1174 -179 -1136 -151
rect -1108 -179 -1070 -151
rect -1042 -179 -1004 -151
rect -976 -179 -938 -151
rect -910 -179 -872 -151
rect -844 -179 -806 -151
rect -778 -179 -740 -151
rect -712 -179 -674 -151
rect -646 -179 -608 -151
rect -580 -179 -542 -151
rect -514 -179 -476 -151
rect -448 -179 -410 -151
rect -382 -179 -344 -151
rect -316 -179 -278 -151
rect -250 -179 -212 -151
rect -184 -179 -146 -151
rect -118 -179 -80 -151
rect -52 -179 -14 -151
rect 14 -179 52 -151
rect 80 -179 118 -151
rect 146 -179 184 -151
rect 212 -179 250 -151
rect 278 -179 316 -151
rect 344 -179 382 -151
rect 410 -179 448 -151
rect 476 -179 514 -151
rect 542 -179 580 -151
rect 608 -179 646 -151
rect 674 -179 712 -151
rect 740 -179 778 -151
rect 806 -179 844 -151
rect 872 -179 910 -151
rect 938 -179 976 -151
rect 1004 -179 1042 -151
rect 1070 -179 1108 -151
rect 1136 -179 1174 -151
rect 1202 -179 1240 -151
rect 1268 -179 1306 -151
rect 1334 -179 1372 -151
rect 1400 -179 1438 -151
rect 1466 -179 1504 -151
rect 1532 -179 1570 -151
rect 1598 -179 1636 -151
rect 1664 -179 1702 -151
rect 1730 -179 1768 -151
rect 1796 -179 1834 -151
rect 1862 -179 1900 -151
rect 1928 -179 1966 -151
rect 1994 -179 2032 -151
rect 2060 -179 2098 -151
rect 2126 -179 2164 -151
rect 2192 -179 2230 -151
rect 2258 -179 2296 -151
rect 2324 -179 2362 -151
rect 2390 -179 2428 -151
rect 2456 -179 2494 -151
rect 2522 -179 2560 -151
rect 2588 -179 2626 -151
rect 2654 -179 2692 -151
rect 2720 -179 2758 -151
rect 2786 -179 2824 -151
rect 2852 -179 2890 -151
rect 2918 -179 2956 -151
rect 2984 -179 3022 -151
rect 3050 -179 3088 -151
rect 3116 -179 3154 -151
rect 3182 -179 3220 -151
rect 3248 -179 3286 -151
rect 3314 -179 3352 -151
rect 3380 -179 3418 -151
rect 3446 -179 3484 -151
rect 3512 -179 3550 -151
rect 3578 -179 3616 -151
rect 3644 -179 3682 -151
rect 3710 -179 3748 -151
rect 3776 -179 3814 -151
rect 3842 -179 3880 -151
rect 3908 -179 3946 -151
rect 3974 -179 4012 -151
rect 4040 -179 4078 -151
rect 4106 -179 4144 -151
rect 4172 -179 4210 -151
rect 4238 -179 4276 -151
rect 4304 -179 4342 -151
rect 4370 -179 4408 -151
rect 4436 -179 4474 -151
rect 4502 -179 4540 -151
rect 4568 -179 4606 -151
rect 4634 -179 4672 -151
rect 4700 -179 4738 -151
rect 4766 -179 4804 -151
rect 4832 -179 4870 -151
rect 4898 -179 4903 -151
rect -4903 -217 4903 -179
rect -4903 -245 -4898 -217
rect -4870 -245 -4832 -217
rect -4804 -245 -4766 -217
rect -4738 -245 -4700 -217
rect -4672 -245 -4634 -217
rect -4606 -245 -4568 -217
rect -4540 -245 -4502 -217
rect -4474 -245 -4436 -217
rect -4408 -245 -4370 -217
rect -4342 -245 -4304 -217
rect -4276 -245 -4238 -217
rect -4210 -245 -4172 -217
rect -4144 -245 -4106 -217
rect -4078 -245 -4040 -217
rect -4012 -245 -3974 -217
rect -3946 -245 -3908 -217
rect -3880 -245 -3842 -217
rect -3814 -245 -3776 -217
rect -3748 -245 -3710 -217
rect -3682 -245 -3644 -217
rect -3616 -245 -3578 -217
rect -3550 -245 -3512 -217
rect -3484 -245 -3446 -217
rect -3418 -245 -3380 -217
rect -3352 -245 -3314 -217
rect -3286 -245 -3248 -217
rect -3220 -245 -3182 -217
rect -3154 -245 -3116 -217
rect -3088 -245 -3050 -217
rect -3022 -245 -2984 -217
rect -2956 -245 -2918 -217
rect -2890 -245 -2852 -217
rect -2824 -245 -2786 -217
rect -2758 -245 -2720 -217
rect -2692 -245 -2654 -217
rect -2626 -245 -2588 -217
rect -2560 -245 -2522 -217
rect -2494 -245 -2456 -217
rect -2428 -245 -2390 -217
rect -2362 -245 -2324 -217
rect -2296 -245 -2258 -217
rect -2230 -245 -2192 -217
rect -2164 -245 -2126 -217
rect -2098 -245 -2060 -217
rect -2032 -245 -1994 -217
rect -1966 -245 -1928 -217
rect -1900 -245 -1862 -217
rect -1834 -245 -1796 -217
rect -1768 -245 -1730 -217
rect -1702 -245 -1664 -217
rect -1636 -245 -1598 -217
rect -1570 -245 -1532 -217
rect -1504 -245 -1466 -217
rect -1438 -245 -1400 -217
rect -1372 -245 -1334 -217
rect -1306 -245 -1268 -217
rect -1240 -245 -1202 -217
rect -1174 -245 -1136 -217
rect -1108 -245 -1070 -217
rect -1042 -245 -1004 -217
rect -976 -245 -938 -217
rect -910 -245 -872 -217
rect -844 -245 -806 -217
rect -778 -245 -740 -217
rect -712 -245 -674 -217
rect -646 -245 -608 -217
rect -580 -245 -542 -217
rect -514 -245 -476 -217
rect -448 -245 -410 -217
rect -382 -245 -344 -217
rect -316 -245 -278 -217
rect -250 -245 -212 -217
rect -184 -245 -146 -217
rect -118 -245 -80 -217
rect -52 -245 -14 -217
rect 14 -245 52 -217
rect 80 -245 118 -217
rect 146 -245 184 -217
rect 212 -245 250 -217
rect 278 -245 316 -217
rect 344 -245 382 -217
rect 410 -245 448 -217
rect 476 -245 514 -217
rect 542 -245 580 -217
rect 608 -245 646 -217
rect 674 -245 712 -217
rect 740 -245 778 -217
rect 806 -245 844 -217
rect 872 -245 910 -217
rect 938 -245 976 -217
rect 1004 -245 1042 -217
rect 1070 -245 1108 -217
rect 1136 -245 1174 -217
rect 1202 -245 1240 -217
rect 1268 -245 1306 -217
rect 1334 -245 1372 -217
rect 1400 -245 1438 -217
rect 1466 -245 1504 -217
rect 1532 -245 1570 -217
rect 1598 -245 1636 -217
rect 1664 -245 1702 -217
rect 1730 -245 1768 -217
rect 1796 -245 1834 -217
rect 1862 -245 1900 -217
rect 1928 -245 1966 -217
rect 1994 -245 2032 -217
rect 2060 -245 2098 -217
rect 2126 -245 2164 -217
rect 2192 -245 2230 -217
rect 2258 -245 2296 -217
rect 2324 -245 2362 -217
rect 2390 -245 2428 -217
rect 2456 -245 2494 -217
rect 2522 -245 2560 -217
rect 2588 -245 2626 -217
rect 2654 -245 2692 -217
rect 2720 -245 2758 -217
rect 2786 -245 2824 -217
rect 2852 -245 2890 -217
rect 2918 -245 2956 -217
rect 2984 -245 3022 -217
rect 3050 -245 3088 -217
rect 3116 -245 3154 -217
rect 3182 -245 3220 -217
rect 3248 -245 3286 -217
rect 3314 -245 3352 -217
rect 3380 -245 3418 -217
rect 3446 -245 3484 -217
rect 3512 -245 3550 -217
rect 3578 -245 3616 -217
rect 3644 -245 3682 -217
rect 3710 -245 3748 -217
rect 3776 -245 3814 -217
rect 3842 -245 3880 -217
rect 3908 -245 3946 -217
rect 3974 -245 4012 -217
rect 4040 -245 4078 -217
rect 4106 -245 4144 -217
rect 4172 -245 4210 -217
rect 4238 -245 4276 -217
rect 4304 -245 4342 -217
rect 4370 -245 4408 -217
rect 4436 -245 4474 -217
rect 4502 -245 4540 -217
rect 4568 -245 4606 -217
rect 4634 -245 4672 -217
rect 4700 -245 4738 -217
rect 4766 -245 4804 -217
rect 4832 -245 4870 -217
rect 4898 -245 4903 -217
rect -4903 -283 4903 -245
rect -4903 -311 -4898 -283
rect -4870 -311 -4832 -283
rect -4804 -311 -4766 -283
rect -4738 -311 -4700 -283
rect -4672 -311 -4634 -283
rect -4606 -311 -4568 -283
rect -4540 -311 -4502 -283
rect -4474 -311 -4436 -283
rect -4408 -311 -4370 -283
rect -4342 -311 -4304 -283
rect -4276 -311 -4238 -283
rect -4210 -311 -4172 -283
rect -4144 -311 -4106 -283
rect -4078 -311 -4040 -283
rect -4012 -311 -3974 -283
rect -3946 -311 -3908 -283
rect -3880 -311 -3842 -283
rect -3814 -311 -3776 -283
rect -3748 -311 -3710 -283
rect -3682 -311 -3644 -283
rect -3616 -311 -3578 -283
rect -3550 -311 -3512 -283
rect -3484 -311 -3446 -283
rect -3418 -311 -3380 -283
rect -3352 -311 -3314 -283
rect -3286 -311 -3248 -283
rect -3220 -311 -3182 -283
rect -3154 -311 -3116 -283
rect -3088 -311 -3050 -283
rect -3022 -311 -2984 -283
rect -2956 -311 -2918 -283
rect -2890 -311 -2852 -283
rect -2824 -311 -2786 -283
rect -2758 -311 -2720 -283
rect -2692 -311 -2654 -283
rect -2626 -311 -2588 -283
rect -2560 -311 -2522 -283
rect -2494 -311 -2456 -283
rect -2428 -311 -2390 -283
rect -2362 -311 -2324 -283
rect -2296 -311 -2258 -283
rect -2230 -311 -2192 -283
rect -2164 -311 -2126 -283
rect -2098 -311 -2060 -283
rect -2032 -311 -1994 -283
rect -1966 -311 -1928 -283
rect -1900 -311 -1862 -283
rect -1834 -311 -1796 -283
rect -1768 -311 -1730 -283
rect -1702 -311 -1664 -283
rect -1636 -311 -1598 -283
rect -1570 -311 -1532 -283
rect -1504 -311 -1466 -283
rect -1438 -311 -1400 -283
rect -1372 -311 -1334 -283
rect -1306 -311 -1268 -283
rect -1240 -311 -1202 -283
rect -1174 -311 -1136 -283
rect -1108 -311 -1070 -283
rect -1042 -311 -1004 -283
rect -976 -311 -938 -283
rect -910 -311 -872 -283
rect -844 -311 -806 -283
rect -778 -311 -740 -283
rect -712 -311 -674 -283
rect -646 -311 -608 -283
rect -580 -311 -542 -283
rect -514 -311 -476 -283
rect -448 -311 -410 -283
rect -382 -311 -344 -283
rect -316 -311 -278 -283
rect -250 -311 -212 -283
rect -184 -311 -146 -283
rect -118 -311 -80 -283
rect -52 -311 -14 -283
rect 14 -311 52 -283
rect 80 -311 118 -283
rect 146 -311 184 -283
rect 212 -311 250 -283
rect 278 -311 316 -283
rect 344 -311 382 -283
rect 410 -311 448 -283
rect 476 -311 514 -283
rect 542 -311 580 -283
rect 608 -311 646 -283
rect 674 -311 712 -283
rect 740 -311 778 -283
rect 806 -311 844 -283
rect 872 -311 910 -283
rect 938 -311 976 -283
rect 1004 -311 1042 -283
rect 1070 -311 1108 -283
rect 1136 -311 1174 -283
rect 1202 -311 1240 -283
rect 1268 -311 1306 -283
rect 1334 -311 1372 -283
rect 1400 -311 1438 -283
rect 1466 -311 1504 -283
rect 1532 -311 1570 -283
rect 1598 -311 1636 -283
rect 1664 -311 1702 -283
rect 1730 -311 1768 -283
rect 1796 -311 1834 -283
rect 1862 -311 1900 -283
rect 1928 -311 1966 -283
rect 1994 -311 2032 -283
rect 2060 -311 2098 -283
rect 2126 -311 2164 -283
rect 2192 -311 2230 -283
rect 2258 -311 2296 -283
rect 2324 -311 2362 -283
rect 2390 -311 2428 -283
rect 2456 -311 2494 -283
rect 2522 -311 2560 -283
rect 2588 -311 2626 -283
rect 2654 -311 2692 -283
rect 2720 -311 2758 -283
rect 2786 -311 2824 -283
rect 2852 -311 2890 -283
rect 2918 -311 2956 -283
rect 2984 -311 3022 -283
rect 3050 -311 3088 -283
rect 3116 -311 3154 -283
rect 3182 -311 3220 -283
rect 3248 -311 3286 -283
rect 3314 -311 3352 -283
rect 3380 -311 3418 -283
rect 3446 -311 3484 -283
rect 3512 -311 3550 -283
rect 3578 -311 3616 -283
rect 3644 -311 3682 -283
rect 3710 -311 3748 -283
rect 3776 -311 3814 -283
rect 3842 -311 3880 -283
rect 3908 -311 3946 -283
rect 3974 -311 4012 -283
rect 4040 -311 4078 -283
rect 4106 -311 4144 -283
rect 4172 -311 4210 -283
rect 4238 -311 4276 -283
rect 4304 -311 4342 -283
rect 4370 -311 4408 -283
rect 4436 -311 4474 -283
rect 4502 -311 4540 -283
rect 4568 -311 4606 -283
rect 4634 -311 4672 -283
rect 4700 -311 4738 -283
rect 4766 -311 4804 -283
rect 4832 -311 4870 -283
rect 4898 -311 4903 -283
rect -4903 -316 4903 -311
<< via4 >>
rect -4898 283 -4870 311
rect -4832 283 -4804 311
rect -4766 283 -4738 311
rect -4700 283 -4672 311
rect -4634 283 -4606 311
rect -4568 283 -4540 311
rect -4502 283 -4474 311
rect -4436 283 -4408 311
rect -4370 283 -4342 311
rect -4304 283 -4276 311
rect -4238 283 -4210 311
rect -4172 283 -4144 311
rect -4106 283 -4078 311
rect -4040 283 -4012 311
rect -3974 283 -3946 311
rect -3908 283 -3880 311
rect -3842 283 -3814 311
rect -3776 283 -3748 311
rect -3710 283 -3682 311
rect -3644 283 -3616 311
rect -3578 283 -3550 311
rect -3512 283 -3484 311
rect -3446 283 -3418 311
rect -3380 283 -3352 311
rect -3314 283 -3286 311
rect -3248 283 -3220 311
rect -3182 283 -3154 311
rect -3116 283 -3088 311
rect -3050 283 -3022 311
rect -2984 283 -2956 311
rect -2918 283 -2890 311
rect -2852 283 -2824 311
rect -2786 283 -2758 311
rect -2720 283 -2692 311
rect -2654 283 -2626 311
rect -2588 283 -2560 311
rect -2522 283 -2494 311
rect -2456 283 -2428 311
rect -2390 283 -2362 311
rect -2324 283 -2296 311
rect -2258 283 -2230 311
rect -2192 283 -2164 311
rect -2126 283 -2098 311
rect -2060 283 -2032 311
rect -1994 283 -1966 311
rect -1928 283 -1900 311
rect -1862 283 -1834 311
rect -1796 283 -1768 311
rect -1730 283 -1702 311
rect -1664 283 -1636 311
rect -1598 283 -1570 311
rect -1532 283 -1504 311
rect -1466 283 -1438 311
rect -1400 283 -1372 311
rect -1334 283 -1306 311
rect -1268 283 -1240 311
rect -1202 283 -1174 311
rect -1136 283 -1108 311
rect -1070 283 -1042 311
rect -1004 283 -976 311
rect -938 283 -910 311
rect -872 283 -844 311
rect -806 283 -778 311
rect -740 283 -712 311
rect -674 283 -646 311
rect -608 283 -580 311
rect -542 283 -514 311
rect -476 283 -448 311
rect -410 283 -382 311
rect -344 283 -316 311
rect -278 283 -250 311
rect -212 283 -184 311
rect -146 283 -118 311
rect -80 283 -52 311
rect -14 283 14 311
rect 52 283 80 311
rect 118 283 146 311
rect 184 283 212 311
rect 250 283 278 311
rect 316 283 344 311
rect 382 283 410 311
rect 448 283 476 311
rect 514 283 542 311
rect 580 283 608 311
rect 646 283 674 311
rect 712 283 740 311
rect 778 283 806 311
rect 844 283 872 311
rect 910 283 938 311
rect 976 283 1004 311
rect 1042 283 1070 311
rect 1108 283 1136 311
rect 1174 283 1202 311
rect 1240 283 1268 311
rect 1306 283 1334 311
rect 1372 283 1400 311
rect 1438 283 1466 311
rect 1504 283 1532 311
rect 1570 283 1598 311
rect 1636 283 1664 311
rect 1702 283 1730 311
rect 1768 283 1796 311
rect 1834 283 1862 311
rect 1900 283 1928 311
rect 1966 283 1994 311
rect 2032 283 2060 311
rect 2098 283 2126 311
rect 2164 283 2192 311
rect 2230 283 2258 311
rect 2296 283 2324 311
rect 2362 283 2390 311
rect 2428 283 2456 311
rect 2494 283 2522 311
rect 2560 283 2588 311
rect 2626 283 2654 311
rect 2692 283 2720 311
rect 2758 283 2786 311
rect 2824 283 2852 311
rect 2890 283 2918 311
rect 2956 283 2984 311
rect 3022 283 3050 311
rect 3088 283 3116 311
rect 3154 283 3182 311
rect 3220 283 3248 311
rect 3286 283 3314 311
rect 3352 283 3380 311
rect 3418 283 3446 311
rect 3484 283 3512 311
rect 3550 283 3578 311
rect 3616 283 3644 311
rect 3682 283 3710 311
rect 3748 283 3776 311
rect 3814 283 3842 311
rect 3880 283 3908 311
rect 3946 283 3974 311
rect 4012 283 4040 311
rect 4078 283 4106 311
rect 4144 283 4172 311
rect 4210 283 4238 311
rect 4276 283 4304 311
rect 4342 283 4370 311
rect 4408 283 4436 311
rect 4474 283 4502 311
rect 4540 283 4568 311
rect 4606 283 4634 311
rect 4672 283 4700 311
rect 4738 283 4766 311
rect 4804 283 4832 311
rect 4870 283 4898 311
rect -4898 217 -4870 245
rect -4832 217 -4804 245
rect -4766 217 -4738 245
rect -4700 217 -4672 245
rect -4634 217 -4606 245
rect -4568 217 -4540 245
rect -4502 217 -4474 245
rect -4436 217 -4408 245
rect -4370 217 -4342 245
rect -4304 217 -4276 245
rect -4238 217 -4210 245
rect -4172 217 -4144 245
rect -4106 217 -4078 245
rect -4040 217 -4012 245
rect -3974 217 -3946 245
rect -3908 217 -3880 245
rect -3842 217 -3814 245
rect -3776 217 -3748 245
rect -3710 217 -3682 245
rect -3644 217 -3616 245
rect -3578 217 -3550 245
rect -3512 217 -3484 245
rect -3446 217 -3418 245
rect -3380 217 -3352 245
rect -3314 217 -3286 245
rect -3248 217 -3220 245
rect -3182 217 -3154 245
rect -3116 217 -3088 245
rect -3050 217 -3022 245
rect -2984 217 -2956 245
rect -2918 217 -2890 245
rect -2852 217 -2824 245
rect -2786 217 -2758 245
rect -2720 217 -2692 245
rect -2654 217 -2626 245
rect -2588 217 -2560 245
rect -2522 217 -2494 245
rect -2456 217 -2428 245
rect -2390 217 -2362 245
rect -2324 217 -2296 245
rect -2258 217 -2230 245
rect -2192 217 -2164 245
rect -2126 217 -2098 245
rect -2060 217 -2032 245
rect -1994 217 -1966 245
rect -1928 217 -1900 245
rect -1862 217 -1834 245
rect -1796 217 -1768 245
rect -1730 217 -1702 245
rect -1664 217 -1636 245
rect -1598 217 -1570 245
rect -1532 217 -1504 245
rect -1466 217 -1438 245
rect -1400 217 -1372 245
rect -1334 217 -1306 245
rect -1268 217 -1240 245
rect -1202 217 -1174 245
rect -1136 217 -1108 245
rect -1070 217 -1042 245
rect -1004 217 -976 245
rect -938 217 -910 245
rect -872 217 -844 245
rect -806 217 -778 245
rect -740 217 -712 245
rect -674 217 -646 245
rect -608 217 -580 245
rect -542 217 -514 245
rect -476 217 -448 245
rect -410 217 -382 245
rect -344 217 -316 245
rect -278 217 -250 245
rect -212 217 -184 245
rect -146 217 -118 245
rect -80 217 -52 245
rect -14 217 14 245
rect 52 217 80 245
rect 118 217 146 245
rect 184 217 212 245
rect 250 217 278 245
rect 316 217 344 245
rect 382 217 410 245
rect 448 217 476 245
rect 514 217 542 245
rect 580 217 608 245
rect 646 217 674 245
rect 712 217 740 245
rect 778 217 806 245
rect 844 217 872 245
rect 910 217 938 245
rect 976 217 1004 245
rect 1042 217 1070 245
rect 1108 217 1136 245
rect 1174 217 1202 245
rect 1240 217 1268 245
rect 1306 217 1334 245
rect 1372 217 1400 245
rect 1438 217 1466 245
rect 1504 217 1532 245
rect 1570 217 1598 245
rect 1636 217 1664 245
rect 1702 217 1730 245
rect 1768 217 1796 245
rect 1834 217 1862 245
rect 1900 217 1928 245
rect 1966 217 1994 245
rect 2032 217 2060 245
rect 2098 217 2126 245
rect 2164 217 2192 245
rect 2230 217 2258 245
rect 2296 217 2324 245
rect 2362 217 2390 245
rect 2428 217 2456 245
rect 2494 217 2522 245
rect 2560 217 2588 245
rect 2626 217 2654 245
rect 2692 217 2720 245
rect 2758 217 2786 245
rect 2824 217 2852 245
rect 2890 217 2918 245
rect 2956 217 2984 245
rect 3022 217 3050 245
rect 3088 217 3116 245
rect 3154 217 3182 245
rect 3220 217 3248 245
rect 3286 217 3314 245
rect 3352 217 3380 245
rect 3418 217 3446 245
rect 3484 217 3512 245
rect 3550 217 3578 245
rect 3616 217 3644 245
rect 3682 217 3710 245
rect 3748 217 3776 245
rect 3814 217 3842 245
rect 3880 217 3908 245
rect 3946 217 3974 245
rect 4012 217 4040 245
rect 4078 217 4106 245
rect 4144 217 4172 245
rect 4210 217 4238 245
rect 4276 217 4304 245
rect 4342 217 4370 245
rect 4408 217 4436 245
rect 4474 217 4502 245
rect 4540 217 4568 245
rect 4606 217 4634 245
rect 4672 217 4700 245
rect 4738 217 4766 245
rect 4804 217 4832 245
rect 4870 217 4898 245
rect -4898 151 -4870 179
rect -4832 151 -4804 179
rect -4766 151 -4738 179
rect -4700 151 -4672 179
rect -4634 151 -4606 179
rect -4568 151 -4540 179
rect -4502 151 -4474 179
rect -4436 151 -4408 179
rect -4370 151 -4342 179
rect -4304 151 -4276 179
rect -4238 151 -4210 179
rect -4172 151 -4144 179
rect -4106 151 -4078 179
rect -4040 151 -4012 179
rect -3974 151 -3946 179
rect -3908 151 -3880 179
rect -3842 151 -3814 179
rect -3776 151 -3748 179
rect -3710 151 -3682 179
rect -3644 151 -3616 179
rect -3578 151 -3550 179
rect -3512 151 -3484 179
rect -3446 151 -3418 179
rect -3380 151 -3352 179
rect -3314 151 -3286 179
rect -3248 151 -3220 179
rect -3182 151 -3154 179
rect -3116 151 -3088 179
rect -3050 151 -3022 179
rect -2984 151 -2956 179
rect -2918 151 -2890 179
rect -2852 151 -2824 179
rect -2786 151 -2758 179
rect -2720 151 -2692 179
rect -2654 151 -2626 179
rect -2588 151 -2560 179
rect -2522 151 -2494 179
rect -2456 151 -2428 179
rect -2390 151 -2362 179
rect -2324 151 -2296 179
rect -2258 151 -2230 179
rect -2192 151 -2164 179
rect -2126 151 -2098 179
rect -2060 151 -2032 179
rect -1994 151 -1966 179
rect -1928 151 -1900 179
rect -1862 151 -1834 179
rect -1796 151 -1768 179
rect -1730 151 -1702 179
rect -1664 151 -1636 179
rect -1598 151 -1570 179
rect -1532 151 -1504 179
rect -1466 151 -1438 179
rect -1400 151 -1372 179
rect -1334 151 -1306 179
rect -1268 151 -1240 179
rect -1202 151 -1174 179
rect -1136 151 -1108 179
rect -1070 151 -1042 179
rect -1004 151 -976 179
rect -938 151 -910 179
rect -872 151 -844 179
rect -806 151 -778 179
rect -740 151 -712 179
rect -674 151 -646 179
rect -608 151 -580 179
rect -542 151 -514 179
rect -476 151 -448 179
rect -410 151 -382 179
rect -344 151 -316 179
rect -278 151 -250 179
rect -212 151 -184 179
rect -146 151 -118 179
rect -80 151 -52 179
rect -14 151 14 179
rect 52 151 80 179
rect 118 151 146 179
rect 184 151 212 179
rect 250 151 278 179
rect 316 151 344 179
rect 382 151 410 179
rect 448 151 476 179
rect 514 151 542 179
rect 580 151 608 179
rect 646 151 674 179
rect 712 151 740 179
rect 778 151 806 179
rect 844 151 872 179
rect 910 151 938 179
rect 976 151 1004 179
rect 1042 151 1070 179
rect 1108 151 1136 179
rect 1174 151 1202 179
rect 1240 151 1268 179
rect 1306 151 1334 179
rect 1372 151 1400 179
rect 1438 151 1466 179
rect 1504 151 1532 179
rect 1570 151 1598 179
rect 1636 151 1664 179
rect 1702 151 1730 179
rect 1768 151 1796 179
rect 1834 151 1862 179
rect 1900 151 1928 179
rect 1966 151 1994 179
rect 2032 151 2060 179
rect 2098 151 2126 179
rect 2164 151 2192 179
rect 2230 151 2258 179
rect 2296 151 2324 179
rect 2362 151 2390 179
rect 2428 151 2456 179
rect 2494 151 2522 179
rect 2560 151 2588 179
rect 2626 151 2654 179
rect 2692 151 2720 179
rect 2758 151 2786 179
rect 2824 151 2852 179
rect 2890 151 2918 179
rect 2956 151 2984 179
rect 3022 151 3050 179
rect 3088 151 3116 179
rect 3154 151 3182 179
rect 3220 151 3248 179
rect 3286 151 3314 179
rect 3352 151 3380 179
rect 3418 151 3446 179
rect 3484 151 3512 179
rect 3550 151 3578 179
rect 3616 151 3644 179
rect 3682 151 3710 179
rect 3748 151 3776 179
rect 3814 151 3842 179
rect 3880 151 3908 179
rect 3946 151 3974 179
rect 4012 151 4040 179
rect 4078 151 4106 179
rect 4144 151 4172 179
rect 4210 151 4238 179
rect 4276 151 4304 179
rect 4342 151 4370 179
rect 4408 151 4436 179
rect 4474 151 4502 179
rect 4540 151 4568 179
rect 4606 151 4634 179
rect 4672 151 4700 179
rect 4738 151 4766 179
rect 4804 151 4832 179
rect 4870 151 4898 179
rect -4898 85 -4870 113
rect -4832 85 -4804 113
rect -4766 85 -4738 113
rect -4700 85 -4672 113
rect -4634 85 -4606 113
rect -4568 85 -4540 113
rect -4502 85 -4474 113
rect -4436 85 -4408 113
rect -4370 85 -4342 113
rect -4304 85 -4276 113
rect -4238 85 -4210 113
rect -4172 85 -4144 113
rect -4106 85 -4078 113
rect -4040 85 -4012 113
rect -3974 85 -3946 113
rect -3908 85 -3880 113
rect -3842 85 -3814 113
rect -3776 85 -3748 113
rect -3710 85 -3682 113
rect -3644 85 -3616 113
rect -3578 85 -3550 113
rect -3512 85 -3484 113
rect -3446 85 -3418 113
rect -3380 85 -3352 113
rect -3314 85 -3286 113
rect -3248 85 -3220 113
rect -3182 85 -3154 113
rect -3116 85 -3088 113
rect -3050 85 -3022 113
rect -2984 85 -2956 113
rect -2918 85 -2890 113
rect -2852 85 -2824 113
rect -2786 85 -2758 113
rect -2720 85 -2692 113
rect -2654 85 -2626 113
rect -2588 85 -2560 113
rect -2522 85 -2494 113
rect -2456 85 -2428 113
rect -2390 85 -2362 113
rect -2324 85 -2296 113
rect -2258 85 -2230 113
rect -2192 85 -2164 113
rect -2126 85 -2098 113
rect -2060 85 -2032 113
rect -1994 85 -1966 113
rect -1928 85 -1900 113
rect -1862 85 -1834 113
rect -1796 85 -1768 113
rect -1730 85 -1702 113
rect -1664 85 -1636 113
rect -1598 85 -1570 113
rect -1532 85 -1504 113
rect -1466 85 -1438 113
rect -1400 85 -1372 113
rect -1334 85 -1306 113
rect -1268 85 -1240 113
rect -1202 85 -1174 113
rect -1136 85 -1108 113
rect -1070 85 -1042 113
rect -1004 85 -976 113
rect -938 85 -910 113
rect -872 85 -844 113
rect -806 85 -778 113
rect -740 85 -712 113
rect -674 85 -646 113
rect -608 85 -580 113
rect -542 85 -514 113
rect -476 85 -448 113
rect -410 85 -382 113
rect -344 85 -316 113
rect -278 85 -250 113
rect -212 85 -184 113
rect -146 85 -118 113
rect -80 85 -52 113
rect -14 85 14 113
rect 52 85 80 113
rect 118 85 146 113
rect 184 85 212 113
rect 250 85 278 113
rect 316 85 344 113
rect 382 85 410 113
rect 448 85 476 113
rect 514 85 542 113
rect 580 85 608 113
rect 646 85 674 113
rect 712 85 740 113
rect 778 85 806 113
rect 844 85 872 113
rect 910 85 938 113
rect 976 85 1004 113
rect 1042 85 1070 113
rect 1108 85 1136 113
rect 1174 85 1202 113
rect 1240 85 1268 113
rect 1306 85 1334 113
rect 1372 85 1400 113
rect 1438 85 1466 113
rect 1504 85 1532 113
rect 1570 85 1598 113
rect 1636 85 1664 113
rect 1702 85 1730 113
rect 1768 85 1796 113
rect 1834 85 1862 113
rect 1900 85 1928 113
rect 1966 85 1994 113
rect 2032 85 2060 113
rect 2098 85 2126 113
rect 2164 85 2192 113
rect 2230 85 2258 113
rect 2296 85 2324 113
rect 2362 85 2390 113
rect 2428 85 2456 113
rect 2494 85 2522 113
rect 2560 85 2588 113
rect 2626 85 2654 113
rect 2692 85 2720 113
rect 2758 85 2786 113
rect 2824 85 2852 113
rect 2890 85 2918 113
rect 2956 85 2984 113
rect 3022 85 3050 113
rect 3088 85 3116 113
rect 3154 85 3182 113
rect 3220 85 3248 113
rect 3286 85 3314 113
rect 3352 85 3380 113
rect 3418 85 3446 113
rect 3484 85 3512 113
rect 3550 85 3578 113
rect 3616 85 3644 113
rect 3682 85 3710 113
rect 3748 85 3776 113
rect 3814 85 3842 113
rect 3880 85 3908 113
rect 3946 85 3974 113
rect 4012 85 4040 113
rect 4078 85 4106 113
rect 4144 85 4172 113
rect 4210 85 4238 113
rect 4276 85 4304 113
rect 4342 85 4370 113
rect 4408 85 4436 113
rect 4474 85 4502 113
rect 4540 85 4568 113
rect 4606 85 4634 113
rect 4672 85 4700 113
rect 4738 85 4766 113
rect 4804 85 4832 113
rect 4870 85 4898 113
rect -4898 19 -4870 47
rect -4832 19 -4804 47
rect -4766 19 -4738 47
rect -4700 19 -4672 47
rect -4634 19 -4606 47
rect -4568 19 -4540 47
rect -4502 19 -4474 47
rect -4436 19 -4408 47
rect -4370 19 -4342 47
rect -4304 19 -4276 47
rect -4238 19 -4210 47
rect -4172 19 -4144 47
rect -4106 19 -4078 47
rect -4040 19 -4012 47
rect -3974 19 -3946 47
rect -3908 19 -3880 47
rect -3842 19 -3814 47
rect -3776 19 -3748 47
rect -3710 19 -3682 47
rect -3644 19 -3616 47
rect -3578 19 -3550 47
rect -3512 19 -3484 47
rect -3446 19 -3418 47
rect -3380 19 -3352 47
rect -3314 19 -3286 47
rect -3248 19 -3220 47
rect -3182 19 -3154 47
rect -3116 19 -3088 47
rect -3050 19 -3022 47
rect -2984 19 -2956 47
rect -2918 19 -2890 47
rect -2852 19 -2824 47
rect -2786 19 -2758 47
rect -2720 19 -2692 47
rect -2654 19 -2626 47
rect -2588 19 -2560 47
rect -2522 19 -2494 47
rect -2456 19 -2428 47
rect -2390 19 -2362 47
rect -2324 19 -2296 47
rect -2258 19 -2230 47
rect -2192 19 -2164 47
rect -2126 19 -2098 47
rect -2060 19 -2032 47
rect -1994 19 -1966 47
rect -1928 19 -1900 47
rect -1862 19 -1834 47
rect -1796 19 -1768 47
rect -1730 19 -1702 47
rect -1664 19 -1636 47
rect -1598 19 -1570 47
rect -1532 19 -1504 47
rect -1466 19 -1438 47
rect -1400 19 -1372 47
rect -1334 19 -1306 47
rect -1268 19 -1240 47
rect -1202 19 -1174 47
rect -1136 19 -1108 47
rect -1070 19 -1042 47
rect -1004 19 -976 47
rect -938 19 -910 47
rect -872 19 -844 47
rect -806 19 -778 47
rect -740 19 -712 47
rect -674 19 -646 47
rect -608 19 -580 47
rect -542 19 -514 47
rect -476 19 -448 47
rect -410 19 -382 47
rect -344 19 -316 47
rect -278 19 -250 47
rect -212 19 -184 47
rect -146 19 -118 47
rect -80 19 -52 47
rect -14 19 14 47
rect 52 19 80 47
rect 118 19 146 47
rect 184 19 212 47
rect 250 19 278 47
rect 316 19 344 47
rect 382 19 410 47
rect 448 19 476 47
rect 514 19 542 47
rect 580 19 608 47
rect 646 19 674 47
rect 712 19 740 47
rect 778 19 806 47
rect 844 19 872 47
rect 910 19 938 47
rect 976 19 1004 47
rect 1042 19 1070 47
rect 1108 19 1136 47
rect 1174 19 1202 47
rect 1240 19 1268 47
rect 1306 19 1334 47
rect 1372 19 1400 47
rect 1438 19 1466 47
rect 1504 19 1532 47
rect 1570 19 1598 47
rect 1636 19 1664 47
rect 1702 19 1730 47
rect 1768 19 1796 47
rect 1834 19 1862 47
rect 1900 19 1928 47
rect 1966 19 1994 47
rect 2032 19 2060 47
rect 2098 19 2126 47
rect 2164 19 2192 47
rect 2230 19 2258 47
rect 2296 19 2324 47
rect 2362 19 2390 47
rect 2428 19 2456 47
rect 2494 19 2522 47
rect 2560 19 2588 47
rect 2626 19 2654 47
rect 2692 19 2720 47
rect 2758 19 2786 47
rect 2824 19 2852 47
rect 2890 19 2918 47
rect 2956 19 2984 47
rect 3022 19 3050 47
rect 3088 19 3116 47
rect 3154 19 3182 47
rect 3220 19 3248 47
rect 3286 19 3314 47
rect 3352 19 3380 47
rect 3418 19 3446 47
rect 3484 19 3512 47
rect 3550 19 3578 47
rect 3616 19 3644 47
rect 3682 19 3710 47
rect 3748 19 3776 47
rect 3814 19 3842 47
rect 3880 19 3908 47
rect 3946 19 3974 47
rect 4012 19 4040 47
rect 4078 19 4106 47
rect 4144 19 4172 47
rect 4210 19 4238 47
rect 4276 19 4304 47
rect 4342 19 4370 47
rect 4408 19 4436 47
rect 4474 19 4502 47
rect 4540 19 4568 47
rect 4606 19 4634 47
rect 4672 19 4700 47
rect 4738 19 4766 47
rect 4804 19 4832 47
rect 4870 19 4898 47
rect -4898 -47 -4870 -19
rect -4832 -47 -4804 -19
rect -4766 -47 -4738 -19
rect -4700 -47 -4672 -19
rect -4634 -47 -4606 -19
rect -4568 -47 -4540 -19
rect -4502 -47 -4474 -19
rect -4436 -47 -4408 -19
rect -4370 -47 -4342 -19
rect -4304 -47 -4276 -19
rect -4238 -47 -4210 -19
rect -4172 -47 -4144 -19
rect -4106 -47 -4078 -19
rect -4040 -47 -4012 -19
rect -3974 -47 -3946 -19
rect -3908 -47 -3880 -19
rect -3842 -47 -3814 -19
rect -3776 -47 -3748 -19
rect -3710 -47 -3682 -19
rect -3644 -47 -3616 -19
rect -3578 -47 -3550 -19
rect -3512 -47 -3484 -19
rect -3446 -47 -3418 -19
rect -3380 -47 -3352 -19
rect -3314 -47 -3286 -19
rect -3248 -47 -3220 -19
rect -3182 -47 -3154 -19
rect -3116 -47 -3088 -19
rect -3050 -47 -3022 -19
rect -2984 -47 -2956 -19
rect -2918 -47 -2890 -19
rect -2852 -47 -2824 -19
rect -2786 -47 -2758 -19
rect -2720 -47 -2692 -19
rect -2654 -47 -2626 -19
rect -2588 -47 -2560 -19
rect -2522 -47 -2494 -19
rect -2456 -47 -2428 -19
rect -2390 -47 -2362 -19
rect -2324 -47 -2296 -19
rect -2258 -47 -2230 -19
rect -2192 -47 -2164 -19
rect -2126 -47 -2098 -19
rect -2060 -47 -2032 -19
rect -1994 -47 -1966 -19
rect -1928 -47 -1900 -19
rect -1862 -47 -1834 -19
rect -1796 -47 -1768 -19
rect -1730 -47 -1702 -19
rect -1664 -47 -1636 -19
rect -1598 -47 -1570 -19
rect -1532 -47 -1504 -19
rect -1466 -47 -1438 -19
rect -1400 -47 -1372 -19
rect -1334 -47 -1306 -19
rect -1268 -47 -1240 -19
rect -1202 -47 -1174 -19
rect -1136 -47 -1108 -19
rect -1070 -47 -1042 -19
rect -1004 -47 -976 -19
rect -938 -47 -910 -19
rect -872 -47 -844 -19
rect -806 -47 -778 -19
rect -740 -47 -712 -19
rect -674 -47 -646 -19
rect -608 -47 -580 -19
rect -542 -47 -514 -19
rect -476 -47 -448 -19
rect -410 -47 -382 -19
rect -344 -47 -316 -19
rect -278 -47 -250 -19
rect -212 -47 -184 -19
rect -146 -47 -118 -19
rect -80 -47 -52 -19
rect -14 -47 14 -19
rect 52 -47 80 -19
rect 118 -47 146 -19
rect 184 -47 212 -19
rect 250 -47 278 -19
rect 316 -47 344 -19
rect 382 -47 410 -19
rect 448 -47 476 -19
rect 514 -47 542 -19
rect 580 -47 608 -19
rect 646 -47 674 -19
rect 712 -47 740 -19
rect 778 -47 806 -19
rect 844 -47 872 -19
rect 910 -47 938 -19
rect 976 -47 1004 -19
rect 1042 -47 1070 -19
rect 1108 -47 1136 -19
rect 1174 -47 1202 -19
rect 1240 -47 1268 -19
rect 1306 -47 1334 -19
rect 1372 -47 1400 -19
rect 1438 -47 1466 -19
rect 1504 -47 1532 -19
rect 1570 -47 1598 -19
rect 1636 -47 1664 -19
rect 1702 -47 1730 -19
rect 1768 -47 1796 -19
rect 1834 -47 1862 -19
rect 1900 -47 1928 -19
rect 1966 -47 1994 -19
rect 2032 -47 2060 -19
rect 2098 -47 2126 -19
rect 2164 -47 2192 -19
rect 2230 -47 2258 -19
rect 2296 -47 2324 -19
rect 2362 -47 2390 -19
rect 2428 -47 2456 -19
rect 2494 -47 2522 -19
rect 2560 -47 2588 -19
rect 2626 -47 2654 -19
rect 2692 -47 2720 -19
rect 2758 -47 2786 -19
rect 2824 -47 2852 -19
rect 2890 -47 2918 -19
rect 2956 -47 2984 -19
rect 3022 -47 3050 -19
rect 3088 -47 3116 -19
rect 3154 -47 3182 -19
rect 3220 -47 3248 -19
rect 3286 -47 3314 -19
rect 3352 -47 3380 -19
rect 3418 -47 3446 -19
rect 3484 -47 3512 -19
rect 3550 -47 3578 -19
rect 3616 -47 3644 -19
rect 3682 -47 3710 -19
rect 3748 -47 3776 -19
rect 3814 -47 3842 -19
rect 3880 -47 3908 -19
rect 3946 -47 3974 -19
rect 4012 -47 4040 -19
rect 4078 -47 4106 -19
rect 4144 -47 4172 -19
rect 4210 -47 4238 -19
rect 4276 -47 4304 -19
rect 4342 -47 4370 -19
rect 4408 -47 4436 -19
rect 4474 -47 4502 -19
rect 4540 -47 4568 -19
rect 4606 -47 4634 -19
rect 4672 -47 4700 -19
rect 4738 -47 4766 -19
rect 4804 -47 4832 -19
rect 4870 -47 4898 -19
rect -4898 -113 -4870 -85
rect -4832 -113 -4804 -85
rect -4766 -113 -4738 -85
rect -4700 -113 -4672 -85
rect -4634 -113 -4606 -85
rect -4568 -113 -4540 -85
rect -4502 -113 -4474 -85
rect -4436 -113 -4408 -85
rect -4370 -113 -4342 -85
rect -4304 -113 -4276 -85
rect -4238 -113 -4210 -85
rect -4172 -113 -4144 -85
rect -4106 -113 -4078 -85
rect -4040 -113 -4012 -85
rect -3974 -113 -3946 -85
rect -3908 -113 -3880 -85
rect -3842 -113 -3814 -85
rect -3776 -113 -3748 -85
rect -3710 -113 -3682 -85
rect -3644 -113 -3616 -85
rect -3578 -113 -3550 -85
rect -3512 -113 -3484 -85
rect -3446 -113 -3418 -85
rect -3380 -113 -3352 -85
rect -3314 -113 -3286 -85
rect -3248 -113 -3220 -85
rect -3182 -113 -3154 -85
rect -3116 -113 -3088 -85
rect -3050 -113 -3022 -85
rect -2984 -113 -2956 -85
rect -2918 -113 -2890 -85
rect -2852 -113 -2824 -85
rect -2786 -113 -2758 -85
rect -2720 -113 -2692 -85
rect -2654 -113 -2626 -85
rect -2588 -113 -2560 -85
rect -2522 -113 -2494 -85
rect -2456 -113 -2428 -85
rect -2390 -113 -2362 -85
rect -2324 -113 -2296 -85
rect -2258 -113 -2230 -85
rect -2192 -113 -2164 -85
rect -2126 -113 -2098 -85
rect -2060 -113 -2032 -85
rect -1994 -113 -1966 -85
rect -1928 -113 -1900 -85
rect -1862 -113 -1834 -85
rect -1796 -113 -1768 -85
rect -1730 -113 -1702 -85
rect -1664 -113 -1636 -85
rect -1598 -113 -1570 -85
rect -1532 -113 -1504 -85
rect -1466 -113 -1438 -85
rect -1400 -113 -1372 -85
rect -1334 -113 -1306 -85
rect -1268 -113 -1240 -85
rect -1202 -113 -1174 -85
rect -1136 -113 -1108 -85
rect -1070 -113 -1042 -85
rect -1004 -113 -976 -85
rect -938 -113 -910 -85
rect -872 -113 -844 -85
rect -806 -113 -778 -85
rect -740 -113 -712 -85
rect -674 -113 -646 -85
rect -608 -113 -580 -85
rect -542 -113 -514 -85
rect -476 -113 -448 -85
rect -410 -113 -382 -85
rect -344 -113 -316 -85
rect -278 -113 -250 -85
rect -212 -113 -184 -85
rect -146 -113 -118 -85
rect -80 -113 -52 -85
rect -14 -113 14 -85
rect 52 -113 80 -85
rect 118 -113 146 -85
rect 184 -113 212 -85
rect 250 -113 278 -85
rect 316 -113 344 -85
rect 382 -113 410 -85
rect 448 -113 476 -85
rect 514 -113 542 -85
rect 580 -113 608 -85
rect 646 -113 674 -85
rect 712 -113 740 -85
rect 778 -113 806 -85
rect 844 -113 872 -85
rect 910 -113 938 -85
rect 976 -113 1004 -85
rect 1042 -113 1070 -85
rect 1108 -113 1136 -85
rect 1174 -113 1202 -85
rect 1240 -113 1268 -85
rect 1306 -113 1334 -85
rect 1372 -113 1400 -85
rect 1438 -113 1466 -85
rect 1504 -113 1532 -85
rect 1570 -113 1598 -85
rect 1636 -113 1664 -85
rect 1702 -113 1730 -85
rect 1768 -113 1796 -85
rect 1834 -113 1862 -85
rect 1900 -113 1928 -85
rect 1966 -113 1994 -85
rect 2032 -113 2060 -85
rect 2098 -113 2126 -85
rect 2164 -113 2192 -85
rect 2230 -113 2258 -85
rect 2296 -113 2324 -85
rect 2362 -113 2390 -85
rect 2428 -113 2456 -85
rect 2494 -113 2522 -85
rect 2560 -113 2588 -85
rect 2626 -113 2654 -85
rect 2692 -113 2720 -85
rect 2758 -113 2786 -85
rect 2824 -113 2852 -85
rect 2890 -113 2918 -85
rect 2956 -113 2984 -85
rect 3022 -113 3050 -85
rect 3088 -113 3116 -85
rect 3154 -113 3182 -85
rect 3220 -113 3248 -85
rect 3286 -113 3314 -85
rect 3352 -113 3380 -85
rect 3418 -113 3446 -85
rect 3484 -113 3512 -85
rect 3550 -113 3578 -85
rect 3616 -113 3644 -85
rect 3682 -113 3710 -85
rect 3748 -113 3776 -85
rect 3814 -113 3842 -85
rect 3880 -113 3908 -85
rect 3946 -113 3974 -85
rect 4012 -113 4040 -85
rect 4078 -113 4106 -85
rect 4144 -113 4172 -85
rect 4210 -113 4238 -85
rect 4276 -113 4304 -85
rect 4342 -113 4370 -85
rect 4408 -113 4436 -85
rect 4474 -113 4502 -85
rect 4540 -113 4568 -85
rect 4606 -113 4634 -85
rect 4672 -113 4700 -85
rect 4738 -113 4766 -85
rect 4804 -113 4832 -85
rect 4870 -113 4898 -85
rect -4898 -179 -4870 -151
rect -4832 -179 -4804 -151
rect -4766 -179 -4738 -151
rect -4700 -179 -4672 -151
rect -4634 -179 -4606 -151
rect -4568 -179 -4540 -151
rect -4502 -179 -4474 -151
rect -4436 -179 -4408 -151
rect -4370 -179 -4342 -151
rect -4304 -179 -4276 -151
rect -4238 -179 -4210 -151
rect -4172 -179 -4144 -151
rect -4106 -179 -4078 -151
rect -4040 -179 -4012 -151
rect -3974 -179 -3946 -151
rect -3908 -179 -3880 -151
rect -3842 -179 -3814 -151
rect -3776 -179 -3748 -151
rect -3710 -179 -3682 -151
rect -3644 -179 -3616 -151
rect -3578 -179 -3550 -151
rect -3512 -179 -3484 -151
rect -3446 -179 -3418 -151
rect -3380 -179 -3352 -151
rect -3314 -179 -3286 -151
rect -3248 -179 -3220 -151
rect -3182 -179 -3154 -151
rect -3116 -179 -3088 -151
rect -3050 -179 -3022 -151
rect -2984 -179 -2956 -151
rect -2918 -179 -2890 -151
rect -2852 -179 -2824 -151
rect -2786 -179 -2758 -151
rect -2720 -179 -2692 -151
rect -2654 -179 -2626 -151
rect -2588 -179 -2560 -151
rect -2522 -179 -2494 -151
rect -2456 -179 -2428 -151
rect -2390 -179 -2362 -151
rect -2324 -179 -2296 -151
rect -2258 -179 -2230 -151
rect -2192 -179 -2164 -151
rect -2126 -179 -2098 -151
rect -2060 -179 -2032 -151
rect -1994 -179 -1966 -151
rect -1928 -179 -1900 -151
rect -1862 -179 -1834 -151
rect -1796 -179 -1768 -151
rect -1730 -179 -1702 -151
rect -1664 -179 -1636 -151
rect -1598 -179 -1570 -151
rect -1532 -179 -1504 -151
rect -1466 -179 -1438 -151
rect -1400 -179 -1372 -151
rect -1334 -179 -1306 -151
rect -1268 -179 -1240 -151
rect -1202 -179 -1174 -151
rect -1136 -179 -1108 -151
rect -1070 -179 -1042 -151
rect -1004 -179 -976 -151
rect -938 -179 -910 -151
rect -872 -179 -844 -151
rect -806 -179 -778 -151
rect -740 -179 -712 -151
rect -674 -179 -646 -151
rect -608 -179 -580 -151
rect -542 -179 -514 -151
rect -476 -179 -448 -151
rect -410 -179 -382 -151
rect -344 -179 -316 -151
rect -278 -179 -250 -151
rect -212 -179 -184 -151
rect -146 -179 -118 -151
rect -80 -179 -52 -151
rect -14 -179 14 -151
rect 52 -179 80 -151
rect 118 -179 146 -151
rect 184 -179 212 -151
rect 250 -179 278 -151
rect 316 -179 344 -151
rect 382 -179 410 -151
rect 448 -179 476 -151
rect 514 -179 542 -151
rect 580 -179 608 -151
rect 646 -179 674 -151
rect 712 -179 740 -151
rect 778 -179 806 -151
rect 844 -179 872 -151
rect 910 -179 938 -151
rect 976 -179 1004 -151
rect 1042 -179 1070 -151
rect 1108 -179 1136 -151
rect 1174 -179 1202 -151
rect 1240 -179 1268 -151
rect 1306 -179 1334 -151
rect 1372 -179 1400 -151
rect 1438 -179 1466 -151
rect 1504 -179 1532 -151
rect 1570 -179 1598 -151
rect 1636 -179 1664 -151
rect 1702 -179 1730 -151
rect 1768 -179 1796 -151
rect 1834 -179 1862 -151
rect 1900 -179 1928 -151
rect 1966 -179 1994 -151
rect 2032 -179 2060 -151
rect 2098 -179 2126 -151
rect 2164 -179 2192 -151
rect 2230 -179 2258 -151
rect 2296 -179 2324 -151
rect 2362 -179 2390 -151
rect 2428 -179 2456 -151
rect 2494 -179 2522 -151
rect 2560 -179 2588 -151
rect 2626 -179 2654 -151
rect 2692 -179 2720 -151
rect 2758 -179 2786 -151
rect 2824 -179 2852 -151
rect 2890 -179 2918 -151
rect 2956 -179 2984 -151
rect 3022 -179 3050 -151
rect 3088 -179 3116 -151
rect 3154 -179 3182 -151
rect 3220 -179 3248 -151
rect 3286 -179 3314 -151
rect 3352 -179 3380 -151
rect 3418 -179 3446 -151
rect 3484 -179 3512 -151
rect 3550 -179 3578 -151
rect 3616 -179 3644 -151
rect 3682 -179 3710 -151
rect 3748 -179 3776 -151
rect 3814 -179 3842 -151
rect 3880 -179 3908 -151
rect 3946 -179 3974 -151
rect 4012 -179 4040 -151
rect 4078 -179 4106 -151
rect 4144 -179 4172 -151
rect 4210 -179 4238 -151
rect 4276 -179 4304 -151
rect 4342 -179 4370 -151
rect 4408 -179 4436 -151
rect 4474 -179 4502 -151
rect 4540 -179 4568 -151
rect 4606 -179 4634 -151
rect 4672 -179 4700 -151
rect 4738 -179 4766 -151
rect 4804 -179 4832 -151
rect 4870 -179 4898 -151
rect -4898 -245 -4870 -217
rect -4832 -245 -4804 -217
rect -4766 -245 -4738 -217
rect -4700 -245 -4672 -217
rect -4634 -245 -4606 -217
rect -4568 -245 -4540 -217
rect -4502 -245 -4474 -217
rect -4436 -245 -4408 -217
rect -4370 -245 -4342 -217
rect -4304 -245 -4276 -217
rect -4238 -245 -4210 -217
rect -4172 -245 -4144 -217
rect -4106 -245 -4078 -217
rect -4040 -245 -4012 -217
rect -3974 -245 -3946 -217
rect -3908 -245 -3880 -217
rect -3842 -245 -3814 -217
rect -3776 -245 -3748 -217
rect -3710 -245 -3682 -217
rect -3644 -245 -3616 -217
rect -3578 -245 -3550 -217
rect -3512 -245 -3484 -217
rect -3446 -245 -3418 -217
rect -3380 -245 -3352 -217
rect -3314 -245 -3286 -217
rect -3248 -245 -3220 -217
rect -3182 -245 -3154 -217
rect -3116 -245 -3088 -217
rect -3050 -245 -3022 -217
rect -2984 -245 -2956 -217
rect -2918 -245 -2890 -217
rect -2852 -245 -2824 -217
rect -2786 -245 -2758 -217
rect -2720 -245 -2692 -217
rect -2654 -245 -2626 -217
rect -2588 -245 -2560 -217
rect -2522 -245 -2494 -217
rect -2456 -245 -2428 -217
rect -2390 -245 -2362 -217
rect -2324 -245 -2296 -217
rect -2258 -245 -2230 -217
rect -2192 -245 -2164 -217
rect -2126 -245 -2098 -217
rect -2060 -245 -2032 -217
rect -1994 -245 -1966 -217
rect -1928 -245 -1900 -217
rect -1862 -245 -1834 -217
rect -1796 -245 -1768 -217
rect -1730 -245 -1702 -217
rect -1664 -245 -1636 -217
rect -1598 -245 -1570 -217
rect -1532 -245 -1504 -217
rect -1466 -245 -1438 -217
rect -1400 -245 -1372 -217
rect -1334 -245 -1306 -217
rect -1268 -245 -1240 -217
rect -1202 -245 -1174 -217
rect -1136 -245 -1108 -217
rect -1070 -245 -1042 -217
rect -1004 -245 -976 -217
rect -938 -245 -910 -217
rect -872 -245 -844 -217
rect -806 -245 -778 -217
rect -740 -245 -712 -217
rect -674 -245 -646 -217
rect -608 -245 -580 -217
rect -542 -245 -514 -217
rect -476 -245 -448 -217
rect -410 -245 -382 -217
rect -344 -245 -316 -217
rect -278 -245 -250 -217
rect -212 -245 -184 -217
rect -146 -245 -118 -217
rect -80 -245 -52 -217
rect -14 -245 14 -217
rect 52 -245 80 -217
rect 118 -245 146 -217
rect 184 -245 212 -217
rect 250 -245 278 -217
rect 316 -245 344 -217
rect 382 -245 410 -217
rect 448 -245 476 -217
rect 514 -245 542 -217
rect 580 -245 608 -217
rect 646 -245 674 -217
rect 712 -245 740 -217
rect 778 -245 806 -217
rect 844 -245 872 -217
rect 910 -245 938 -217
rect 976 -245 1004 -217
rect 1042 -245 1070 -217
rect 1108 -245 1136 -217
rect 1174 -245 1202 -217
rect 1240 -245 1268 -217
rect 1306 -245 1334 -217
rect 1372 -245 1400 -217
rect 1438 -245 1466 -217
rect 1504 -245 1532 -217
rect 1570 -245 1598 -217
rect 1636 -245 1664 -217
rect 1702 -245 1730 -217
rect 1768 -245 1796 -217
rect 1834 -245 1862 -217
rect 1900 -245 1928 -217
rect 1966 -245 1994 -217
rect 2032 -245 2060 -217
rect 2098 -245 2126 -217
rect 2164 -245 2192 -217
rect 2230 -245 2258 -217
rect 2296 -245 2324 -217
rect 2362 -245 2390 -217
rect 2428 -245 2456 -217
rect 2494 -245 2522 -217
rect 2560 -245 2588 -217
rect 2626 -245 2654 -217
rect 2692 -245 2720 -217
rect 2758 -245 2786 -217
rect 2824 -245 2852 -217
rect 2890 -245 2918 -217
rect 2956 -245 2984 -217
rect 3022 -245 3050 -217
rect 3088 -245 3116 -217
rect 3154 -245 3182 -217
rect 3220 -245 3248 -217
rect 3286 -245 3314 -217
rect 3352 -245 3380 -217
rect 3418 -245 3446 -217
rect 3484 -245 3512 -217
rect 3550 -245 3578 -217
rect 3616 -245 3644 -217
rect 3682 -245 3710 -217
rect 3748 -245 3776 -217
rect 3814 -245 3842 -217
rect 3880 -245 3908 -217
rect 3946 -245 3974 -217
rect 4012 -245 4040 -217
rect 4078 -245 4106 -217
rect 4144 -245 4172 -217
rect 4210 -245 4238 -217
rect 4276 -245 4304 -217
rect 4342 -245 4370 -217
rect 4408 -245 4436 -217
rect 4474 -245 4502 -217
rect 4540 -245 4568 -217
rect 4606 -245 4634 -217
rect 4672 -245 4700 -217
rect 4738 -245 4766 -217
rect 4804 -245 4832 -217
rect 4870 -245 4898 -217
rect -4898 -311 -4870 -283
rect -4832 -311 -4804 -283
rect -4766 -311 -4738 -283
rect -4700 -311 -4672 -283
rect -4634 -311 -4606 -283
rect -4568 -311 -4540 -283
rect -4502 -311 -4474 -283
rect -4436 -311 -4408 -283
rect -4370 -311 -4342 -283
rect -4304 -311 -4276 -283
rect -4238 -311 -4210 -283
rect -4172 -311 -4144 -283
rect -4106 -311 -4078 -283
rect -4040 -311 -4012 -283
rect -3974 -311 -3946 -283
rect -3908 -311 -3880 -283
rect -3842 -311 -3814 -283
rect -3776 -311 -3748 -283
rect -3710 -311 -3682 -283
rect -3644 -311 -3616 -283
rect -3578 -311 -3550 -283
rect -3512 -311 -3484 -283
rect -3446 -311 -3418 -283
rect -3380 -311 -3352 -283
rect -3314 -311 -3286 -283
rect -3248 -311 -3220 -283
rect -3182 -311 -3154 -283
rect -3116 -311 -3088 -283
rect -3050 -311 -3022 -283
rect -2984 -311 -2956 -283
rect -2918 -311 -2890 -283
rect -2852 -311 -2824 -283
rect -2786 -311 -2758 -283
rect -2720 -311 -2692 -283
rect -2654 -311 -2626 -283
rect -2588 -311 -2560 -283
rect -2522 -311 -2494 -283
rect -2456 -311 -2428 -283
rect -2390 -311 -2362 -283
rect -2324 -311 -2296 -283
rect -2258 -311 -2230 -283
rect -2192 -311 -2164 -283
rect -2126 -311 -2098 -283
rect -2060 -311 -2032 -283
rect -1994 -311 -1966 -283
rect -1928 -311 -1900 -283
rect -1862 -311 -1834 -283
rect -1796 -311 -1768 -283
rect -1730 -311 -1702 -283
rect -1664 -311 -1636 -283
rect -1598 -311 -1570 -283
rect -1532 -311 -1504 -283
rect -1466 -311 -1438 -283
rect -1400 -311 -1372 -283
rect -1334 -311 -1306 -283
rect -1268 -311 -1240 -283
rect -1202 -311 -1174 -283
rect -1136 -311 -1108 -283
rect -1070 -311 -1042 -283
rect -1004 -311 -976 -283
rect -938 -311 -910 -283
rect -872 -311 -844 -283
rect -806 -311 -778 -283
rect -740 -311 -712 -283
rect -674 -311 -646 -283
rect -608 -311 -580 -283
rect -542 -311 -514 -283
rect -476 -311 -448 -283
rect -410 -311 -382 -283
rect -344 -311 -316 -283
rect -278 -311 -250 -283
rect -212 -311 -184 -283
rect -146 -311 -118 -283
rect -80 -311 -52 -283
rect -14 -311 14 -283
rect 52 -311 80 -283
rect 118 -311 146 -283
rect 184 -311 212 -283
rect 250 -311 278 -283
rect 316 -311 344 -283
rect 382 -311 410 -283
rect 448 -311 476 -283
rect 514 -311 542 -283
rect 580 -311 608 -283
rect 646 -311 674 -283
rect 712 -311 740 -283
rect 778 -311 806 -283
rect 844 -311 872 -283
rect 910 -311 938 -283
rect 976 -311 1004 -283
rect 1042 -311 1070 -283
rect 1108 -311 1136 -283
rect 1174 -311 1202 -283
rect 1240 -311 1268 -283
rect 1306 -311 1334 -283
rect 1372 -311 1400 -283
rect 1438 -311 1466 -283
rect 1504 -311 1532 -283
rect 1570 -311 1598 -283
rect 1636 -311 1664 -283
rect 1702 -311 1730 -283
rect 1768 -311 1796 -283
rect 1834 -311 1862 -283
rect 1900 -311 1928 -283
rect 1966 -311 1994 -283
rect 2032 -311 2060 -283
rect 2098 -311 2126 -283
rect 2164 -311 2192 -283
rect 2230 -311 2258 -283
rect 2296 -311 2324 -283
rect 2362 -311 2390 -283
rect 2428 -311 2456 -283
rect 2494 -311 2522 -283
rect 2560 -311 2588 -283
rect 2626 -311 2654 -283
rect 2692 -311 2720 -283
rect 2758 -311 2786 -283
rect 2824 -311 2852 -283
rect 2890 -311 2918 -283
rect 2956 -311 2984 -283
rect 3022 -311 3050 -283
rect 3088 -311 3116 -283
rect 3154 -311 3182 -283
rect 3220 -311 3248 -283
rect 3286 -311 3314 -283
rect 3352 -311 3380 -283
rect 3418 -311 3446 -283
rect 3484 -311 3512 -283
rect 3550 -311 3578 -283
rect 3616 -311 3644 -283
rect 3682 -311 3710 -283
rect 3748 -311 3776 -283
rect 3814 -311 3842 -283
rect 3880 -311 3908 -283
rect 3946 -311 3974 -283
rect 4012 -311 4040 -283
rect 4078 -311 4106 -283
rect 4144 -311 4172 -283
rect 4210 -311 4238 -283
rect 4276 -311 4304 -283
rect 4342 -311 4370 -283
rect 4408 -311 4436 -283
rect 4474 -311 4502 -283
rect 4540 -311 4568 -283
rect 4606 -311 4634 -283
rect 4672 -311 4700 -283
rect 4738 -311 4766 -283
rect 4804 -311 4832 -283
rect 4870 -311 4898 -283
<< metal5 >>
rect -4906 311 4906 319
rect -4906 283 -4898 311
rect -4870 283 -4832 311
rect -4804 283 -4766 311
rect -4738 283 -4700 311
rect -4672 283 -4634 311
rect -4606 283 -4568 311
rect -4540 283 -4502 311
rect -4474 283 -4436 311
rect -4408 283 -4370 311
rect -4342 283 -4304 311
rect -4276 283 -4238 311
rect -4210 283 -4172 311
rect -4144 283 -4106 311
rect -4078 283 -4040 311
rect -4012 283 -3974 311
rect -3946 283 -3908 311
rect -3880 283 -3842 311
rect -3814 283 -3776 311
rect -3748 283 -3710 311
rect -3682 283 -3644 311
rect -3616 283 -3578 311
rect -3550 283 -3512 311
rect -3484 283 -3446 311
rect -3418 283 -3380 311
rect -3352 283 -3314 311
rect -3286 283 -3248 311
rect -3220 283 -3182 311
rect -3154 283 -3116 311
rect -3088 283 -3050 311
rect -3022 283 -2984 311
rect -2956 283 -2918 311
rect -2890 283 -2852 311
rect -2824 283 -2786 311
rect -2758 283 -2720 311
rect -2692 283 -2654 311
rect -2626 283 -2588 311
rect -2560 283 -2522 311
rect -2494 283 -2456 311
rect -2428 283 -2390 311
rect -2362 283 -2324 311
rect -2296 283 -2258 311
rect -2230 283 -2192 311
rect -2164 283 -2126 311
rect -2098 283 -2060 311
rect -2032 283 -1994 311
rect -1966 283 -1928 311
rect -1900 283 -1862 311
rect -1834 283 -1796 311
rect -1768 283 -1730 311
rect -1702 283 -1664 311
rect -1636 283 -1598 311
rect -1570 283 -1532 311
rect -1504 283 -1466 311
rect -1438 283 -1400 311
rect -1372 283 -1334 311
rect -1306 283 -1268 311
rect -1240 283 -1202 311
rect -1174 283 -1136 311
rect -1108 283 -1070 311
rect -1042 283 -1004 311
rect -976 283 -938 311
rect -910 283 -872 311
rect -844 283 -806 311
rect -778 283 -740 311
rect -712 283 -674 311
rect -646 283 -608 311
rect -580 283 -542 311
rect -514 283 -476 311
rect -448 283 -410 311
rect -382 283 -344 311
rect -316 283 -278 311
rect -250 283 -212 311
rect -184 283 -146 311
rect -118 283 -80 311
rect -52 283 -14 311
rect 14 283 52 311
rect 80 283 118 311
rect 146 283 184 311
rect 212 283 250 311
rect 278 283 316 311
rect 344 283 382 311
rect 410 283 448 311
rect 476 283 514 311
rect 542 283 580 311
rect 608 283 646 311
rect 674 283 712 311
rect 740 283 778 311
rect 806 283 844 311
rect 872 283 910 311
rect 938 283 976 311
rect 1004 283 1042 311
rect 1070 283 1108 311
rect 1136 283 1174 311
rect 1202 283 1240 311
rect 1268 283 1306 311
rect 1334 283 1372 311
rect 1400 283 1438 311
rect 1466 283 1504 311
rect 1532 283 1570 311
rect 1598 283 1636 311
rect 1664 283 1702 311
rect 1730 283 1768 311
rect 1796 283 1834 311
rect 1862 283 1900 311
rect 1928 283 1966 311
rect 1994 283 2032 311
rect 2060 283 2098 311
rect 2126 283 2164 311
rect 2192 283 2230 311
rect 2258 283 2296 311
rect 2324 283 2362 311
rect 2390 283 2428 311
rect 2456 283 2494 311
rect 2522 283 2560 311
rect 2588 283 2626 311
rect 2654 283 2692 311
rect 2720 283 2758 311
rect 2786 283 2824 311
rect 2852 283 2890 311
rect 2918 283 2956 311
rect 2984 283 3022 311
rect 3050 283 3088 311
rect 3116 283 3154 311
rect 3182 283 3220 311
rect 3248 283 3286 311
rect 3314 283 3352 311
rect 3380 283 3418 311
rect 3446 283 3484 311
rect 3512 283 3550 311
rect 3578 283 3616 311
rect 3644 283 3682 311
rect 3710 283 3748 311
rect 3776 283 3814 311
rect 3842 283 3880 311
rect 3908 283 3946 311
rect 3974 283 4012 311
rect 4040 283 4078 311
rect 4106 283 4144 311
rect 4172 283 4210 311
rect 4238 283 4276 311
rect 4304 283 4342 311
rect 4370 283 4408 311
rect 4436 283 4474 311
rect 4502 283 4540 311
rect 4568 283 4606 311
rect 4634 283 4672 311
rect 4700 283 4738 311
rect 4766 283 4804 311
rect 4832 283 4870 311
rect 4898 283 4906 311
rect -4906 245 4906 283
rect -4906 217 -4898 245
rect -4870 217 -4832 245
rect -4804 217 -4766 245
rect -4738 217 -4700 245
rect -4672 217 -4634 245
rect -4606 217 -4568 245
rect -4540 217 -4502 245
rect -4474 217 -4436 245
rect -4408 217 -4370 245
rect -4342 217 -4304 245
rect -4276 217 -4238 245
rect -4210 217 -4172 245
rect -4144 217 -4106 245
rect -4078 217 -4040 245
rect -4012 217 -3974 245
rect -3946 217 -3908 245
rect -3880 217 -3842 245
rect -3814 217 -3776 245
rect -3748 217 -3710 245
rect -3682 217 -3644 245
rect -3616 217 -3578 245
rect -3550 217 -3512 245
rect -3484 217 -3446 245
rect -3418 217 -3380 245
rect -3352 217 -3314 245
rect -3286 217 -3248 245
rect -3220 217 -3182 245
rect -3154 217 -3116 245
rect -3088 217 -3050 245
rect -3022 217 -2984 245
rect -2956 217 -2918 245
rect -2890 217 -2852 245
rect -2824 217 -2786 245
rect -2758 217 -2720 245
rect -2692 217 -2654 245
rect -2626 217 -2588 245
rect -2560 217 -2522 245
rect -2494 217 -2456 245
rect -2428 217 -2390 245
rect -2362 217 -2324 245
rect -2296 217 -2258 245
rect -2230 217 -2192 245
rect -2164 217 -2126 245
rect -2098 217 -2060 245
rect -2032 217 -1994 245
rect -1966 217 -1928 245
rect -1900 217 -1862 245
rect -1834 217 -1796 245
rect -1768 217 -1730 245
rect -1702 217 -1664 245
rect -1636 217 -1598 245
rect -1570 217 -1532 245
rect -1504 217 -1466 245
rect -1438 217 -1400 245
rect -1372 217 -1334 245
rect -1306 217 -1268 245
rect -1240 217 -1202 245
rect -1174 217 -1136 245
rect -1108 217 -1070 245
rect -1042 217 -1004 245
rect -976 217 -938 245
rect -910 217 -872 245
rect -844 217 -806 245
rect -778 217 -740 245
rect -712 217 -674 245
rect -646 217 -608 245
rect -580 217 -542 245
rect -514 217 -476 245
rect -448 217 -410 245
rect -382 217 -344 245
rect -316 217 -278 245
rect -250 217 -212 245
rect -184 217 -146 245
rect -118 217 -80 245
rect -52 217 -14 245
rect 14 217 52 245
rect 80 217 118 245
rect 146 217 184 245
rect 212 217 250 245
rect 278 217 316 245
rect 344 217 382 245
rect 410 217 448 245
rect 476 217 514 245
rect 542 217 580 245
rect 608 217 646 245
rect 674 217 712 245
rect 740 217 778 245
rect 806 217 844 245
rect 872 217 910 245
rect 938 217 976 245
rect 1004 217 1042 245
rect 1070 217 1108 245
rect 1136 217 1174 245
rect 1202 217 1240 245
rect 1268 217 1306 245
rect 1334 217 1372 245
rect 1400 217 1438 245
rect 1466 217 1504 245
rect 1532 217 1570 245
rect 1598 217 1636 245
rect 1664 217 1702 245
rect 1730 217 1768 245
rect 1796 217 1834 245
rect 1862 217 1900 245
rect 1928 217 1966 245
rect 1994 217 2032 245
rect 2060 217 2098 245
rect 2126 217 2164 245
rect 2192 217 2230 245
rect 2258 217 2296 245
rect 2324 217 2362 245
rect 2390 217 2428 245
rect 2456 217 2494 245
rect 2522 217 2560 245
rect 2588 217 2626 245
rect 2654 217 2692 245
rect 2720 217 2758 245
rect 2786 217 2824 245
rect 2852 217 2890 245
rect 2918 217 2956 245
rect 2984 217 3022 245
rect 3050 217 3088 245
rect 3116 217 3154 245
rect 3182 217 3220 245
rect 3248 217 3286 245
rect 3314 217 3352 245
rect 3380 217 3418 245
rect 3446 217 3484 245
rect 3512 217 3550 245
rect 3578 217 3616 245
rect 3644 217 3682 245
rect 3710 217 3748 245
rect 3776 217 3814 245
rect 3842 217 3880 245
rect 3908 217 3946 245
rect 3974 217 4012 245
rect 4040 217 4078 245
rect 4106 217 4144 245
rect 4172 217 4210 245
rect 4238 217 4276 245
rect 4304 217 4342 245
rect 4370 217 4408 245
rect 4436 217 4474 245
rect 4502 217 4540 245
rect 4568 217 4606 245
rect 4634 217 4672 245
rect 4700 217 4738 245
rect 4766 217 4804 245
rect 4832 217 4870 245
rect 4898 217 4906 245
rect -4906 179 4906 217
rect -4906 151 -4898 179
rect -4870 151 -4832 179
rect -4804 151 -4766 179
rect -4738 151 -4700 179
rect -4672 151 -4634 179
rect -4606 151 -4568 179
rect -4540 151 -4502 179
rect -4474 151 -4436 179
rect -4408 151 -4370 179
rect -4342 151 -4304 179
rect -4276 151 -4238 179
rect -4210 151 -4172 179
rect -4144 151 -4106 179
rect -4078 151 -4040 179
rect -4012 151 -3974 179
rect -3946 151 -3908 179
rect -3880 151 -3842 179
rect -3814 151 -3776 179
rect -3748 151 -3710 179
rect -3682 151 -3644 179
rect -3616 151 -3578 179
rect -3550 151 -3512 179
rect -3484 151 -3446 179
rect -3418 151 -3380 179
rect -3352 151 -3314 179
rect -3286 151 -3248 179
rect -3220 151 -3182 179
rect -3154 151 -3116 179
rect -3088 151 -3050 179
rect -3022 151 -2984 179
rect -2956 151 -2918 179
rect -2890 151 -2852 179
rect -2824 151 -2786 179
rect -2758 151 -2720 179
rect -2692 151 -2654 179
rect -2626 151 -2588 179
rect -2560 151 -2522 179
rect -2494 151 -2456 179
rect -2428 151 -2390 179
rect -2362 151 -2324 179
rect -2296 151 -2258 179
rect -2230 151 -2192 179
rect -2164 151 -2126 179
rect -2098 151 -2060 179
rect -2032 151 -1994 179
rect -1966 151 -1928 179
rect -1900 151 -1862 179
rect -1834 151 -1796 179
rect -1768 151 -1730 179
rect -1702 151 -1664 179
rect -1636 151 -1598 179
rect -1570 151 -1532 179
rect -1504 151 -1466 179
rect -1438 151 -1400 179
rect -1372 151 -1334 179
rect -1306 151 -1268 179
rect -1240 151 -1202 179
rect -1174 151 -1136 179
rect -1108 151 -1070 179
rect -1042 151 -1004 179
rect -976 151 -938 179
rect -910 151 -872 179
rect -844 151 -806 179
rect -778 151 -740 179
rect -712 151 -674 179
rect -646 151 -608 179
rect -580 151 -542 179
rect -514 151 -476 179
rect -448 151 -410 179
rect -382 151 -344 179
rect -316 151 -278 179
rect -250 151 -212 179
rect -184 151 -146 179
rect -118 151 -80 179
rect -52 151 -14 179
rect 14 151 52 179
rect 80 151 118 179
rect 146 151 184 179
rect 212 151 250 179
rect 278 151 316 179
rect 344 151 382 179
rect 410 151 448 179
rect 476 151 514 179
rect 542 151 580 179
rect 608 151 646 179
rect 674 151 712 179
rect 740 151 778 179
rect 806 151 844 179
rect 872 151 910 179
rect 938 151 976 179
rect 1004 151 1042 179
rect 1070 151 1108 179
rect 1136 151 1174 179
rect 1202 151 1240 179
rect 1268 151 1306 179
rect 1334 151 1372 179
rect 1400 151 1438 179
rect 1466 151 1504 179
rect 1532 151 1570 179
rect 1598 151 1636 179
rect 1664 151 1702 179
rect 1730 151 1768 179
rect 1796 151 1834 179
rect 1862 151 1900 179
rect 1928 151 1966 179
rect 1994 151 2032 179
rect 2060 151 2098 179
rect 2126 151 2164 179
rect 2192 151 2230 179
rect 2258 151 2296 179
rect 2324 151 2362 179
rect 2390 151 2428 179
rect 2456 151 2494 179
rect 2522 151 2560 179
rect 2588 151 2626 179
rect 2654 151 2692 179
rect 2720 151 2758 179
rect 2786 151 2824 179
rect 2852 151 2890 179
rect 2918 151 2956 179
rect 2984 151 3022 179
rect 3050 151 3088 179
rect 3116 151 3154 179
rect 3182 151 3220 179
rect 3248 151 3286 179
rect 3314 151 3352 179
rect 3380 151 3418 179
rect 3446 151 3484 179
rect 3512 151 3550 179
rect 3578 151 3616 179
rect 3644 151 3682 179
rect 3710 151 3748 179
rect 3776 151 3814 179
rect 3842 151 3880 179
rect 3908 151 3946 179
rect 3974 151 4012 179
rect 4040 151 4078 179
rect 4106 151 4144 179
rect 4172 151 4210 179
rect 4238 151 4276 179
rect 4304 151 4342 179
rect 4370 151 4408 179
rect 4436 151 4474 179
rect 4502 151 4540 179
rect 4568 151 4606 179
rect 4634 151 4672 179
rect 4700 151 4738 179
rect 4766 151 4804 179
rect 4832 151 4870 179
rect 4898 151 4906 179
rect -4906 113 4906 151
rect -4906 85 -4898 113
rect -4870 85 -4832 113
rect -4804 85 -4766 113
rect -4738 85 -4700 113
rect -4672 85 -4634 113
rect -4606 85 -4568 113
rect -4540 85 -4502 113
rect -4474 85 -4436 113
rect -4408 85 -4370 113
rect -4342 85 -4304 113
rect -4276 85 -4238 113
rect -4210 85 -4172 113
rect -4144 85 -4106 113
rect -4078 85 -4040 113
rect -4012 85 -3974 113
rect -3946 85 -3908 113
rect -3880 85 -3842 113
rect -3814 85 -3776 113
rect -3748 85 -3710 113
rect -3682 85 -3644 113
rect -3616 85 -3578 113
rect -3550 85 -3512 113
rect -3484 85 -3446 113
rect -3418 85 -3380 113
rect -3352 85 -3314 113
rect -3286 85 -3248 113
rect -3220 85 -3182 113
rect -3154 85 -3116 113
rect -3088 85 -3050 113
rect -3022 85 -2984 113
rect -2956 85 -2918 113
rect -2890 85 -2852 113
rect -2824 85 -2786 113
rect -2758 85 -2720 113
rect -2692 85 -2654 113
rect -2626 85 -2588 113
rect -2560 85 -2522 113
rect -2494 85 -2456 113
rect -2428 85 -2390 113
rect -2362 85 -2324 113
rect -2296 85 -2258 113
rect -2230 85 -2192 113
rect -2164 85 -2126 113
rect -2098 85 -2060 113
rect -2032 85 -1994 113
rect -1966 85 -1928 113
rect -1900 85 -1862 113
rect -1834 85 -1796 113
rect -1768 85 -1730 113
rect -1702 85 -1664 113
rect -1636 85 -1598 113
rect -1570 85 -1532 113
rect -1504 85 -1466 113
rect -1438 85 -1400 113
rect -1372 85 -1334 113
rect -1306 85 -1268 113
rect -1240 85 -1202 113
rect -1174 85 -1136 113
rect -1108 85 -1070 113
rect -1042 85 -1004 113
rect -976 85 -938 113
rect -910 85 -872 113
rect -844 85 -806 113
rect -778 85 -740 113
rect -712 85 -674 113
rect -646 85 -608 113
rect -580 85 -542 113
rect -514 85 -476 113
rect -448 85 -410 113
rect -382 85 -344 113
rect -316 85 -278 113
rect -250 85 -212 113
rect -184 85 -146 113
rect -118 85 -80 113
rect -52 85 -14 113
rect 14 85 52 113
rect 80 85 118 113
rect 146 85 184 113
rect 212 85 250 113
rect 278 85 316 113
rect 344 85 382 113
rect 410 85 448 113
rect 476 85 514 113
rect 542 85 580 113
rect 608 85 646 113
rect 674 85 712 113
rect 740 85 778 113
rect 806 85 844 113
rect 872 85 910 113
rect 938 85 976 113
rect 1004 85 1042 113
rect 1070 85 1108 113
rect 1136 85 1174 113
rect 1202 85 1240 113
rect 1268 85 1306 113
rect 1334 85 1372 113
rect 1400 85 1438 113
rect 1466 85 1504 113
rect 1532 85 1570 113
rect 1598 85 1636 113
rect 1664 85 1702 113
rect 1730 85 1768 113
rect 1796 85 1834 113
rect 1862 85 1900 113
rect 1928 85 1966 113
rect 1994 85 2032 113
rect 2060 85 2098 113
rect 2126 85 2164 113
rect 2192 85 2230 113
rect 2258 85 2296 113
rect 2324 85 2362 113
rect 2390 85 2428 113
rect 2456 85 2494 113
rect 2522 85 2560 113
rect 2588 85 2626 113
rect 2654 85 2692 113
rect 2720 85 2758 113
rect 2786 85 2824 113
rect 2852 85 2890 113
rect 2918 85 2956 113
rect 2984 85 3022 113
rect 3050 85 3088 113
rect 3116 85 3154 113
rect 3182 85 3220 113
rect 3248 85 3286 113
rect 3314 85 3352 113
rect 3380 85 3418 113
rect 3446 85 3484 113
rect 3512 85 3550 113
rect 3578 85 3616 113
rect 3644 85 3682 113
rect 3710 85 3748 113
rect 3776 85 3814 113
rect 3842 85 3880 113
rect 3908 85 3946 113
rect 3974 85 4012 113
rect 4040 85 4078 113
rect 4106 85 4144 113
rect 4172 85 4210 113
rect 4238 85 4276 113
rect 4304 85 4342 113
rect 4370 85 4408 113
rect 4436 85 4474 113
rect 4502 85 4540 113
rect 4568 85 4606 113
rect 4634 85 4672 113
rect 4700 85 4738 113
rect 4766 85 4804 113
rect 4832 85 4870 113
rect 4898 85 4906 113
rect -4906 47 4906 85
rect -4906 19 -4898 47
rect -4870 19 -4832 47
rect -4804 19 -4766 47
rect -4738 19 -4700 47
rect -4672 19 -4634 47
rect -4606 19 -4568 47
rect -4540 19 -4502 47
rect -4474 19 -4436 47
rect -4408 19 -4370 47
rect -4342 19 -4304 47
rect -4276 19 -4238 47
rect -4210 19 -4172 47
rect -4144 19 -4106 47
rect -4078 19 -4040 47
rect -4012 19 -3974 47
rect -3946 19 -3908 47
rect -3880 19 -3842 47
rect -3814 19 -3776 47
rect -3748 19 -3710 47
rect -3682 19 -3644 47
rect -3616 19 -3578 47
rect -3550 19 -3512 47
rect -3484 19 -3446 47
rect -3418 19 -3380 47
rect -3352 19 -3314 47
rect -3286 19 -3248 47
rect -3220 19 -3182 47
rect -3154 19 -3116 47
rect -3088 19 -3050 47
rect -3022 19 -2984 47
rect -2956 19 -2918 47
rect -2890 19 -2852 47
rect -2824 19 -2786 47
rect -2758 19 -2720 47
rect -2692 19 -2654 47
rect -2626 19 -2588 47
rect -2560 19 -2522 47
rect -2494 19 -2456 47
rect -2428 19 -2390 47
rect -2362 19 -2324 47
rect -2296 19 -2258 47
rect -2230 19 -2192 47
rect -2164 19 -2126 47
rect -2098 19 -2060 47
rect -2032 19 -1994 47
rect -1966 19 -1928 47
rect -1900 19 -1862 47
rect -1834 19 -1796 47
rect -1768 19 -1730 47
rect -1702 19 -1664 47
rect -1636 19 -1598 47
rect -1570 19 -1532 47
rect -1504 19 -1466 47
rect -1438 19 -1400 47
rect -1372 19 -1334 47
rect -1306 19 -1268 47
rect -1240 19 -1202 47
rect -1174 19 -1136 47
rect -1108 19 -1070 47
rect -1042 19 -1004 47
rect -976 19 -938 47
rect -910 19 -872 47
rect -844 19 -806 47
rect -778 19 -740 47
rect -712 19 -674 47
rect -646 19 -608 47
rect -580 19 -542 47
rect -514 19 -476 47
rect -448 19 -410 47
rect -382 19 -344 47
rect -316 19 -278 47
rect -250 19 -212 47
rect -184 19 -146 47
rect -118 19 -80 47
rect -52 19 -14 47
rect 14 19 52 47
rect 80 19 118 47
rect 146 19 184 47
rect 212 19 250 47
rect 278 19 316 47
rect 344 19 382 47
rect 410 19 448 47
rect 476 19 514 47
rect 542 19 580 47
rect 608 19 646 47
rect 674 19 712 47
rect 740 19 778 47
rect 806 19 844 47
rect 872 19 910 47
rect 938 19 976 47
rect 1004 19 1042 47
rect 1070 19 1108 47
rect 1136 19 1174 47
rect 1202 19 1240 47
rect 1268 19 1306 47
rect 1334 19 1372 47
rect 1400 19 1438 47
rect 1466 19 1504 47
rect 1532 19 1570 47
rect 1598 19 1636 47
rect 1664 19 1702 47
rect 1730 19 1768 47
rect 1796 19 1834 47
rect 1862 19 1900 47
rect 1928 19 1966 47
rect 1994 19 2032 47
rect 2060 19 2098 47
rect 2126 19 2164 47
rect 2192 19 2230 47
rect 2258 19 2296 47
rect 2324 19 2362 47
rect 2390 19 2428 47
rect 2456 19 2494 47
rect 2522 19 2560 47
rect 2588 19 2626 47
rect 2654 19 2692 47
rect 2720 19 2758 47
rect 2786 19 2824 47
rect 2852 19 2890 47
rect 2918 19 2956 47
rect 2984 19 3022 47
rect 3050 19 3088 47
rect 3116 19 3154 47
rect 3182 19 3220 47
rect 3248 19 3286 47
rect 3314 19 3352 47
rect 3380 19 3418 47
rect 3446 19 3484 47
rect 3512 19 3550 47
rect 3578 19 3616 47
rect 3644 19 3682 47
rect 3710 19 3748 47
rect 3776 19 3814 47
rect 3842 19 3880 47
rect 3908 19 3946 47
rect 3974 19 4012 47
rect 4040 19 4078 47
rect 4106 19 4144 47
rect 4172 19 4210 47
rect 4238 19 4276 47
rect 4304 19 4342 47
rect 4370 19 4408 47
rect 4436 19 4474 47
rect 4502 19 4540 47
rect 4568 19 4606 47
rect 4634 19 4672 47
rect 4700 19 4738 47
rect 4766 19 4804 47
rect 4832 19 4870 47
rect 4898 19 4906 47
rect -4906 -19 4906 19
rect -4906 -47 -4898 -19
rect -4870 -47 -4832 -19
rect -4804 -47 -4766 -19
rect -4738 -47 -4700 -19
rect -4672 -47 -4634 -19
rect -4606 -47 -4568 -19
rect -4540 -47 -4502 -19
rect -4474 -47 -4436 -19
rect -4408 -47 -4370 -19
rect -4342 -47 -4304 -19
rect -4276 -47 -4238 -19
rect -4210 -47 -4172 -19
rect -4144 -47 -4106 -19
rect -4078 -47 -4040 -19
rect -4012 -47 -3974 -19
rect -3946 -47 -3908 -19
rect -3880 -47 -3842 -19
rect -3814 -47 -3776 -19
rect -3748 -47 -3710 -19
rect -3682 -47 -3644 -19
rect -3616 -47 -3578 -19
rect -3550 -47 -3512 -19
rect -3484 -47 -3446 -19
rect -3418 -47 -3380 -19
rect -3352 -47 -3314 -19
rect -3286 -47 -3248 -19
rect -3220 -47 -3182 -19
rect -3154 -47 -3116 -19
rect -3088 -47 -3050 -19
rect -3022 -47 -2984 -19
rect -2956 -47 -2918 -19
rect -2890 -47 -2852 -19
rect -2824 -47 -2786 -19
rect -2758 -47 -2720 -19
rect -2692 -47 -2654 -19
rect -2626 -47 -2588 -19
rect -2560 -47 -2522 -19
rect -2494 -47 -2456 -19
rect -2428 -47 -2390 -19
rect -2362 -47 -2324 -19
rect -2296 -47 -2258 -19
rect -2230 -47 -2192 -19
rect -2164 -47 -2126 -19
rect -2098 -47 -2060 -19
rect -2032 -47 -1994 -19
rect -1966 -47 -1928 -19
rect -1900 -47 -1862 -19
rect -1834 -47 -1796 -19
rect -1768 -47 -1730 -19
rect -1702 -47 -1664 -19
rect -1636 -47 -1598 -19
rect -1570 -47 -1532 -19
rect -1504 -47 -1466 -19
rect -1438 -47 -1400 -19
rect -1372 -47 -1334 -19
rect -1306 -47 -1268 -19
rect -1240 -47 -1202 -19
rect -1174 -47 -1136 -19
rect -1108 -47 -1070 -19
rect -1042 -47 -1004 -19
rect -976 -47 -938 -19
rect -910 -47 -872 -19
rect -844 -47 -806 -19
rect -778 -47 -740 -19
rect -712 -47 -674 -19
rect -646 -47 -608 -19
rect -580 -47 -542 -19
rect -514 -47 -476 -19
rect -448 -47 -410 -19
rect -382 -47 -344 -19
rect -316 -47 -278 -19
rect -250 -47 -212 -19
rect -184 -47 -146 -19
rect -118 -47 -80 -19
rect -52 -47 -14 -19
rect 14 -47 52 -19
rect 80 -47 118 -19
rect 146 -47 184 -19
rect 212 -47 250 -19
rect 278 -47 316 -19
rect 344 -47 382 -19
rect 410 -47 448 -19
rect 476 -47 514 -19
rect 542 -47 580 -19
rect 608 -47 646 -19
rect 674 -47 712 -19
rect 740 -47 778 -19
rect 806 -47 844 -19
rect 872 -47 910 -19
rect 938 -47 976 -19
rect 1004 -47 1042 -19
rect 1070 -47 1108 -19
rect 1136 -47 1174 -19
rect 1202 -47 1240 -19
rect 1268 -47 1306 -19
rect 1334 -47 1372 -19
rect 1400 -47 1438 -19
rect 1466 -47 1504 -19
rect 1532 -47 1570 -19
rect 1598 -47 1636 -19
rect 1664 -47 1702 -19
rect 1730 -47 1768 -19
rect 1796 -47 1834 -19
rect 1862 -47 1900 -19
rect 1928 -47 1966 -19
rect 1994 -47 2032 -19
rect 2060 -47 2098 -19
rect 2126 -47 2164 -19
rect 2192 -47 2230 -19
rect 2258 -47 2296 -19
rect 2324 -47 2362 -19
rect 2390 -47 2428 -19
rect 2456 -47 2494 -19
rect 2522 -47 2560 -19
rect 2588 -47 2626 -19
rect 2654 -47 2692 -19
rect 2720 -47 2758 -19
rect 2786 -47 2824 -19
rect 2852 -47 2890 -19
rect 2918 -47 2956 -19
rect 2984 -47 3022 -19
rect 3050 -47 3088 -19
rect 3116 -47 3154 -19
rect 3182 -47 3220 -19
rect 3248 -47 3286 -19
rect 3314 -47 3352 -19
rect 3380 -47 3418 -19
rect 3446 -47 3484 -19
rect 3512 -47 3550 -19
rect 3578 -47 3616 -19
rect 3644 -47 3682 -19
rect 3710 -47 3748 -19
rect 3776 -47 3814 -19
rect 3842 -47 3880 -19
rect 3908 -47 3946 -19
rect 3974 -47 4012 -19
rect 4040 -47 4078 -19
rect 4106 -47 4144 -19
rect 4172 -47 4210 -19
rect 4238 -47 4276 -19
rect 4304 -47 4342 -19
rect 4370 -47 4408 -19
rect 4436 -47 4474 -19
rect 4502 -47 4540 -19
rect 4568 -47 4606 -19
rect 4634 -47 4672 -19
rect 4700 -47 4738 -19
rect 4766 -47 4804 -19
rect 4832 -47 4870 -19
rect 4898 -47 4906 -19
rect -4906 -85 4906 -47
rect -4906 -113 -4898 -85
rect -4870 -113 -4832 -85
rect -4804 -113 -4766 -85
rect -4738 -113 -4700 -85
rect -4672 -113 -4634 -85
rect -4606 -113 -4568 -85
rect -4540 -113 -4502 -85
rect -4474 -113 -4436 -85
rect -4408 -113 -4370 -85
rect -4342 -113 -4304 -85
rect -4276 -113 -4238 -85
rect -4210 -113 -4172 -85
rect -4144 -113 -4106 -85
rect -4078 -113 -4040 -85
rect -4012 -113 -3974 -85
rect -3946 -113 -3908 -85
rect -3880 -113 -3842 -85
rect -3814 -113 -3776 -85
rect -3748 -113 -3710 -85
rect -3682 -113 -3644 -85
rect -3616 -113 -3578 -85
rect -3550 -113 -3512 -85
rect -3484 -113 -3446 -85
rect -3418 -113 -3380 -85
rect -3352 -113 -3314 -85
rect -3286 -113 -3248 -85
rect -3220 -113 -3182 -85
rect -3154 -113 -3116 -85
rect -3088 -113 -3050 -85
rect -3022 -113 -2984 -85
rect -2956 -113 -2918 -85
rect -2890 -113 -2852 -85
rect -2824 -113 -2786 -85
rect -2758 -113 -2720 -85
rect -2692 -113 -2654 -85
rect -2626 -113 -2588 -85
rect -2560 -113 -2522 -85
rect -2494 -113 -2456 -85
rect -2428 -113 -2390 -85
rect -2362 -113 -2324 -85
rect -2296 -113 -2258 -85
rect -2230 -113 -2192 -85
rect -2164 -113 -2126 -85
rect -2098 -113 -2060 -85
rect -2032 -113 -1994 -85
rect -1966 -113 -1928 -85
rect -1900 -113 -1862 -85
rect -1834 -113 -1796 -85
rect -1768 -113 -1730 -85
rect -1702 -113 -1664 -85
rect -1636 -113 -1598 -85
rect -1570 -113 -1532 -85
rect -1504 -113 -1466 -85
rect -1438 -113 -1400 -85
rect -1372 -113 -1334 -85
rect -1306 -113 -1268 -85
rect -1240 -113 -1202 -85
rect -1174 -113 -1136 -85
rect -1108 -113 -1070 -85
rect -1042 -113 -1004 -85
rect -976 -113 -938 -85
rect -910 -113 -872 -85
rect -844 -113 -806 -85
rect -778 -113 -740 -85
rect -712 -113 -674 -85
rect -646 -113 -608 -85
rect -580 -113 -542 -85
rect -514 -113 -476 -85
rect -448 -113 -410 -85
rect -382 -113 -344 -85
rect -316 -113 -278 -85
rect -250 -113 -212 -85
rect -184 -113 -146 -85
rect -118 -113 -80 -85
rect -52 -113 -14 -85
rect 14 -113 52 -85
rect 80 -113 118 -85
rect 146 -113 184 -85
rect 212 -113 250 -85
rect 278 -113 316 -85
rect 344 -113 382 -85
rect 410 -113 448 -85
rect 476 -113 514 -85
rect 542 -113 580 -85
rect 608 -113 646 -85
rect 674 -113 712 -85
rect 740 -113 778 -85
rect 806 -113 844 -85
rect 872 -113 910 -85
rect 938 -113 976 -85
rect 1004 -113 1042 -85
rect 1070 -113 1108 -85
rect 1136 -113 1174 -85
rect 1202 -113 1240 -85
rect 1268 -113 1306 -85
rect 1334 -113 1372 -85
rect 1400 -113 1438 -85
rect 1466 -113 1504 -85
rect 1532 -113 1570 -85
rect 1598 -113 1636 -85
rect 1664 -113 1702 -85
rect 1730 -113 1768 -85
rect 1796 -113 1834 -85
rect 1862 -113 1900 -85
rect 1928 -113 1966 -85
rect 1994 -113 2032 -85
rect 2060 -113 2098 -85
rect 2126 -113 2164 -85
rect 2192 -113 2230 -85
rect 2258 -113 2296 -85
rect 2324 -113 2362 -85
rect 2390 -113 2428 -85
rect 2456 -113 2494 -85
rect 2522 -113 2560 -85
rect 2588 -113 2626 -85
rect 2654 -113 2692 -85
rect 2720 -113 2758 -85
rect 2786 -113 2824 -85
rect 2852 -113 2890 -85
rect 2918 -113 2956 -85
rect 2984 -113 3022 -85
rect 3050 -113 3088 -85
rect 3116 -113 3154 -85
rect 3182 -113 3220 -85
rect 3248 -113 3286 -85
rect 3314 -113 3352 -85
rect 3380 -113 3418 -85
rect 3446 -113 3484 -85
rect 3512 -113 3550 -85
rect 3578 -113 3616 -85
rect 3644 -113 3682 -85
rect 3710 -113 3748 -85
rect 3776 -113 3814 -85
rect 3842 -113 3880 -85
rect 3908 -113 3946 -85
rect 3974 -113 4012 -85
rect 4040 -113 4078 -85
rect 4106 -113 4144 -85
rect 4172 -113 4210 -85
rect 4238 -113 4276 -85
rect 4304 -113 4342 -85
rect 4370 -113 4408 -85
rect 4436 -113 4474 -85
rect 4502 -113 4540 -85
rect 4568 -113 4606 -85
rect 4634 -113 4672 -85
rect 4700 -113 4738 -85
rect 4766 -113 4804 -85
rect 4832 -113 4870 -85
rect 4898 -113 4906 -85
rect -4906 -151 4906 -113
rect -4906 -179 -4898 -151
rect -4870 -179 -4832 -151
rect -4804 -179 -4766 -151
rect -4738 -179 -4700 -151
rect -4672 -179 -4634 -151
rect -4606 -179 -4568 -151
rect -4540 -179 -4502 -151
rect -4474 -179 -4436 -151
rect -4408 -179 -4370 -151
rect -4342 -179 -4304 -151
rect -4276 -179 -4238 -151
rect -4210 -179 -4172 -151
rect -4144 -179 -4106 -151
rect -4078 -179 -4040 -151
rect -4012 -179 -3974 -151
rect -3946 -179 -3908 -151
rect -3880 -179 -3842 -151
rect -3814 -179 -3776 -151
rect -3748 -179 -3710 -151
rect -3682 -179 -3644 -151
rect -3616 -179 -3578 -151
rect -3550 -179 -3512 -151
rect -3484 -179 -3446 -151
rect -3418 -179 -3380 -151
rect -3352 -179 -3314 -151
rect -3286 -179 -3248 -151
rect -3220 -179 -3182 -151
rect -3154 -179 -3116 -151
rect -3088 -179 -3050 -151
rect -3022 -179 -2984 -151
rect -2956 -179 -2918 -151
rect -2890 -179 -2852 -151
rect -2824 -179 -2786 -151
rect -2758 -179 -2720 -151
rect -2692 -179 -2654 -151
rect -2626 -179 -2588 -151
rect -2560 -179 -2522 -151
rect -2494 -179 -2456 -151
rect -2428 -179 -2390 -151
rect -2362 -179 -2324 -151
rect -2296 -179 -2258 -151
rect -2230 -179 -2192 -151
rect -2164 -179 -2126 -151
rect -2098 -179 -2060 -151
rect -2032 -179 -1994 -151
rect -1966 -179 -1928 -151
rect -1900 -179 -1862 -151
rect -1834 -179 -1796 -151
rect -1768 -179 -1730 -151
rect -1702 -179 -1664 -151
rect -1636 -179 -1598 -151
rect -1570 -179 -1532 -151
rect -1504 -179 -1466 -151
rect -1438 -179 -1400 -151
rect -1372 -179 -1334 -151
rect -1306 -179 -1268 -151
rect -1240 -179 -1202 -151
rect -1174 -179 -1136 -151
rect -1108 -179 -1070 -151
rect -1042 -179 -1004 -151
rect -976 -179 -938 -151
rect -910 -179 -872 -151
rect -844 -179 -806 -151
rect -778 -179 -740 -151
rect -712 -179 -674 -151
rect -646 -179 -608 -151
rect -580 -179 -542 -151
rect -514 -179 -476 -151
rect -448 -179 -410 -151
rect -382 -179 -344 -151
rect -316 -179 -278 -151
rect -250 -179 -212 -151
rect -184 -179 -146 -151
rect -118 -179 -80 -151
rect -52 -179 -14 -151
rect 14 -179 52 -151
rect 80 -179 118 -151
rect 146 -179 184 -151
rect 212 -179 250 -151
rect 278 -179 316 -151
rect 344 -179 382 -151
rect 410 -179 448 -151
rect 476 -179 514 -151
rect 542 -179 580 -151
rect 608 -179 646 -151
rect 674 -179 712 -151
rect 740 -179 778 -151
rect 806 -179 844 -151
rect 872 -179 910 -151
rect 938 -179 976 -151
rect 1004 -179 1042 -151
rect 1070 -179 1108 -151
rect 1136 -179 1174 -151
rect 1202 -179 1240 -151
rect 1268 -179 1306 -151
rect 1334 -179 1372 -151
rect 1400 -179 1438 -151
rect 1466 -179 1504 -151
rect 1532 -179 1570 -151
rect 1598 -179 1636 -151
rect 1664 -179 1702 -151
rect 1730 -179 1768 -151
rect 1796 -179 1834 -151
rect 1862 -179 1900 -151
rect 1928 -179 1966 -151
rect 1994 -179 2032 -151
rect 2060 -179 2098 -151
rect 2126 -179 2164 -151
rect 2192 -179 2230 -151
rect 2258 -179 2296 -151
rect 2324 -179 2362 -151
rect 2390 -179 2428 -151
rect 2456 -179 2494 -151
rect 2522 -179 2560 -151
rect 2588 -179 2626 -151
rect 2654 -179 2692 -151
rect 2720 -179 2758 -151
rect 2786 -179 2824 -151
rect 2852 -179 2890 -151
rect 2918 -179 2956 -151
rect 2984 -179 3022 -151
rect 3050 -179 3088 -151
rect 3116 -179 3154 -151
rect 3182 -179 3220 -151
rect 3248 -179 3286 -151
rect 3314 -179 3352 -151
rect 3380 -179 3418 -151
rect 3446 -179 3484 -151
rect 3512 -179 3550 -151
rect 3578 -179 3616 -151
rect 3644 -179 3682 -151
rect 3710 -179 3748 -151
rect 3776 -179 3814 -151
rect 3842 -179 3880 -151
rect 3908 -179 3946 -151
rect 3974 -179 4012 -151
rect 4040 -179 4078 -151
rect 4106 -179 4144 -151
rect 4172 -179 4210 -151
rect 4238 -179 4276 -151
rect 4304 -179 4342 -151
rect 4370 -179 4408 -151
rect 4436 -179 4474 -151
rect 4502 -179 4540 -151
rect 4568 -179 4606 -151
rect 4634 -179 4672 -151
rect 4700 -179 4738 -151
rect 4766 -179 4804 -151
rect 4832 -179 4870 -151
rect 4898 -179 4906 -151
rect -4906 -217 4906 -179
rect -4906 -245 -4898 -217
rect -4870 -245 -4832 -217
rect -4804 -245 -4766 -217
rect -4738 -245 -4700 -217
rect -4672 -245 -4634 -217
rect -4606 -245 -4568 -217
rect -4540 -245 -4502 -217
rect -4474 -245 -4436 -217
rect -4408 -245 -4370 -217
rect -4342 -245 -4304 -217
rect -4276 -245 -4238 -217
rect -4210 -245 -4172 -217
rect -4144 -245 -4106 -217
rect -4078 -245 -4040 -217
rect -4012 -245 -3974 -217
rect -3946 -245 -3908 -217
rect -3880 -245 -3842 -217
rect -3814 -245 -3776 -217
rect -3748 -245 -3710 -217
rect -3682 -245 -3644 -217
rect -3616 -245 -3578 -217
rect -3550 -245 -3512 -217
rect -3484 -245 -3446 -217
rect -3418 -245 -3380 -217
rect -3352 -245 -3314 -217
rect -3286 -245 -3248 -217
rect -3220 -245 -3182 -217
rect -3154 -245 -3116 -217
rect -3088 -245 -3050 -217
rect -3022 -245 -2984 -217
rect -2956 -245 -2918 -217
rect -2890 -245 -2852 -217
rect -2824 -245 -2786 -217
rect -2758 -245 -2720 -217
rect -2692 -245 -2654 -217
rect -2626 -245 -2588 -217
rect -2560 -245 -2522 -217
rect -2494 -245 -2456 -217
rect -2428 -245 -2390 -217
rect -2362 -245 -2324 -217
rect -2296 -245 -2258 -217
rect -2230 -245 -2192 -217
rect -2164 -245 -2126 -217
rect -2098 -245 -2060 -217
rect -2032 -245 -1994 -217
rect -1966 -245 -1928 -217
rect -1900 -245 -1862 -217
rect -1834 -245 -1796 -217
rect -1768 -245 -1730 -217
rect -1702 -245 -1664 -217
rect -1636 -245 -1598 -217
rect -1570 -245 -1532 -217
rect -1504 -245 -1466 -217
rect -1438 -245 -1400 -217
rect -1372 -245 -1334 -217
rect -1306 -245 -1268 -217
rect -1240 -245 -1202 -217
rect -1174 -245 -1136 -217
rect -1108 -245 -1070 -217
rect -1042 -245 -1004 -217
rect -976 -245 -938 -217
rect -910 -245 -872 -217
rect -844 -245 -806 -217
rect -778 -245 -740 -217
rect -712 -245 -674 -217
rect -646 -245 -608 -217
rect -580 -245 -542 -217
rect -514 -245 -476 -217
rect -448 -245 -410 -217
rect -382 -245 -344 -217
rect -316 -245 -278 -217
rect -250 -245 -212 -217
rect -184 -245 -146 -217
rect -118 -245 -80 -217
rect -52 -245 -14 -217
rect 14 -245 52 -217
rect 80 -245 118 -217
rect 146 -245 184 -217
rect 212 -245 250 -217
rect 278 -245 316 -217
rect 344 -245 382 -217
rect 410 -245 448 -217
rect 476 -245 514 -217
rect 542 -245 580 -217
rect 608 -245 646 -217
rect 674 -245 712 -217
rect 740 -245 778 -217
rect 806 -245 844 -217
rect 872 -245 910 -217
rect 938 -245 976 -217
rect 1004 -245 1042 -217
rect 1070 -245 1108 -217
rect 1136 -245 1174 -217
rect 1202 -245 1240 -217
rect 1268 -245 1306 -217
rect 1334 -245 1372 -217
rect 1400 -245 1438 -217
rect 1466 -245 1504 -217
rect 1532 -245 1570 -217
rect 1598 -245 1636 -217
rect 1664 -245 1702 -217
rect 1730 -245 1768 -217
rect 1796 -245 1834 -217
rect 1862 -245 1900 -217
rect 1928 -245 1966 -217
rect 1994 -245 2032 -217
rect 2060 -245 2098 -217
rect 2126 -245 2164 -217
rect 2192 -245 2230 -217
rect 2258 -245 2296 -217
rect 2324 -245 2362 -217
rect 2390 -245 2428 -217
rect 2456 -245 2494 -217
rect 2522 -245 2560 -217
rect 2588 -245 2626 -217
rect 2654 -245 2692 -217
rect 2720 -245 2758 -217
rect 2786 -245 2824 -217
rect 2852 -245 2890 -217
rect 2918 -245 2956 -217
rect 2984 -245 3022 -217
rect 3050 -245 3088 -217
rect 3116 -245 3154 -217
rect 3182 -245 3220 -217
rect 3248 -245 3286 -217
rect 3314 -245 3352 -217
rect 3380 -245 3418 -217
rect 3446 -245 3484 -217
rect 3512 -245 3550 -217
rect 3578 -245 3616 -217
rect 3644 -245 3682 -217
rect 3710 -245 3748 -217
rect 3776 -245 3814 -217
rect 3842 -245 3880 -217
rect 3908 -245 3946 -217
rect 3974 -245 4012 -217
rect 4040 -245 4078 -217
rect 4106 -245 4144 -217
rect 4172 -245 4210 -217
rect 4238 -245 4276 -217
rect 4304 -245 4342 -217
rect 4370 -245 4408 -217
rect 4436 -245 4474 -217
rect 4502 -245 4540 -217
rect 4568 -245 4606 -217
rect 4634 -245 4672 -217
rect 4700 -245 4738 -217
rect 4766 -245 4804 -217
rect 4832 -245 4870 -217
rect 4898 -245 4906 -217
rect -4906 -283 4906 -245
rect -4906 -311 -4898 -283
rect -4870 -311 -4832 -283
rect -4804 -311 -4766 -283
rect -4738 -311 -4700 -283
rect -4672 -311 -4634 -283
rect -4606 -311 -4568 -283
rect -4540 -311 -4502 -283
rect -4474 -311 -4436 -283
rect -4408 -311 -4370 -283
rect -4342 -311 -4304 -283
rect -4276 -311 -4238 -283
rect -4210 -311 -4172 -283
rect -4144 -311 -4106 -283
rect -4078 -311 -4040 -283
rect -4012 -311 -3974 -283
rect -3946 -311 -3908 -283
rect -3880 -311 -3842 -283
rect -3814 -311 -3776 -283
rect -3748 -311 -3710 -283
rect -3682 -311 -3644 -283
rect -3616 -311 -3578 -283
rect -3550 -311 -3512 -283
rect -3484 -311 -3446 -283
rect -3418 -311 -3380 -283
rect -3352 -311 -3314 -283
rect -3286 -311 -3248 -283
rect -3220 -311 -3182 -283
rect -3154 -311 -3116 -283
rect -3088 -311 -3050 -283
rect -3022 -311 -2984 -283
rect -2956 -311 -2918 -283
rect -2890 -311 -2852 -283
rect -2824 -311 -2786 -283
rect -2758 -311 -2720 -283
rect -2692 -311 -2654 -283
rect -2626 -311 -2588 -283
rect -2560 -311 -2522 -283
rect -2494 -311 -2456 -283
rect -2428 -311 -2390 -283
rect -2362 -311 -2324 -283
rect -2296 -311 -2258 -283
rect -2230 -311 -2192 -283
rect -2164 -311 -2126 -283
rect -2098 -311 -2060 -283
rect -2032 -311 -1994 -283
rect -1966 -311 -1928 -283
rect -1900 -311 -1862 -283
rect -1834 -311 -1796 -283
rect -1768 -311 -1730 -283
rect -1702 -311 -1664 -283
rect -1636 -311 -1598 -283
rect -1570 -311 -1532 -283
rect -1504 -311 -1466 -283
rect -1438 -311 -1400 -283
rect -1372 -311 -1334 -283
rect -1306 -311 -1268 -283
rect -1240 -311 -1202 -283
rect -1174 -311 -1136 -283
rect -1108 -311 -1070 -283
rect -1042 -311 -1004 -283
rect -976 -311 -938 -283
rect -910 -311 -872 -283
rect -844 -311 -806 -283
rect -778 -311 -740 -283
rect -712 -311 -674 -283
rect -646 -311 -608 -283
rect -580 -311 -542 -283
rect -514 -311 -476 -283
rect -448 -311 -410 -283
rect -382 -311 -344 -283
rect -316 -311 -278 -283
rect -250 -311 -212 -283
rect -184 -311 -146 -283
rect -118 -311 -80 -283
rect -52 -311 -14 -283
rect 14 -311 52 -283
rect 80 -311 118 -283
rect 146 -311 184 -283
rect 212 -311 250 -283
rect 278 -311 316 -283
rect 344 -311 382 -283
rect 410 -311 448 -283
rect 476 -311 514 -283
rect 542 -311 580 -283
rect 608 -311 646 -283
rect 674 -311 712 -283
rect 740 -311 778 -283
rect 806 -311 844 -283
rect 872 -311 910 -283
rect 938 -311 976 -283
rect 1004 -311 1042 -283
rect 1070 -311 1108 -283
rect 1136 -311 1174 -283
rect 1202 -311 1240 -283
rect 1268 -311 1306 -283
rect 1334 -311 1372 -283
rect 1400 -311 1438 -283
rect 1466 -311 1504 -283
rect 1532 -311 1570 -283
rect 1598 -311 1636 -283
rect 1664 -311 1702 -283
rect 1730 -311 1768 -283
rect 1796 -311 1834 -283
rect 1862 -311 1900 -283
rect 1928 -311 1966 -283
rect 1994 -311 2032 -283
rect 2060 -311 2098 -283
rect 2126 -311 2164 -283
rect 2192 -311 2230 -283
rect 2258 -311 2296 -283
rect 2324 -311 2362 -283
rect 2390 -311 2428 -283
rect 2456 -311 2494 -283
rect 2522 -311 2560 -283
rect 2588 -311 2626 -283
rect 2654 -311 2692 -283
rect 2720 -311 2758 -283
rect 2786 -311 2824 -283
rect 2852 -311 2890 -283
rect 2918 -311 2956 -283
rect 2984 -311 3022 -283
rect 3050 -311 3088 -283
rect 3116 -311 3154 -283
rect 3182 -311 3220 -283
rect 3248 -311 3286 -283
rect 3314 -311 3352 -283
rect 3380 -311 3418 -283
rect 3446 -311 3484 -283
rect 3512 -311 3550 -283
rect 3578 -311 3616 -283
rect 3644 -311 3682 -283
rect 3710 -311 3748 -283
rect 3776 -311 3814 -283
rect 3842 -311 3880 -283
rect 3908 -311 3946 -283
rect 3974 -311 4012 -283
rect 4040 -311 4078 -283
rect 4106 -311 4144 -283
rect 4172 -311 4210 -283
rect 4238 -311 4276 -283
rect 4304 -311 4342 -283
rect 4370 -311 4408 -283
rect 4436 -311 4474 -283
rect 4502 -311 4540 -283
rect 4568 -311 4606 -283
rect 4634 -311 4672 -283
rect 4700 -311 4738 -283
rect 4766 -311 4804 -283
rect 4832 -311 4870 -283
rect 4898 -311 4906 -283
rect -4906 -319 4906 -311
<< end >>
