* NGSPICE file created from nmos_3p3_GGGST2_flat.ext - technology: gf180mcuC

.subckt nmos_3p3_GGGST2_flat CLK VIN VOUT
X0 VOUT Inverter_Layout_0.OUT.t0 VIN.t58 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1 VOUT Inverter_Layout_0.OUT.t1 VIN.t57 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X2 VIN CLK.t0 VOUT.t70 Inverter_Layout_0.VSS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X3 VOUT CLK.t1 VIN.t8 Inverter_Layout_0.VSS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X4 VOUT CLK.t2 VIN.t16 Inverter_Layout_0.VSS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X5 Inverter_Layout_0.VSS CLK.t3 Inverter_Layout_0.OUT Inverter_Layout_0.VSS nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X6 VIN Inverter_Layout_0.OUT.t2 VOUT.t64 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X7 VOUT Inverter_Layout_0.OUT.t3 VIN.t56 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X8 VOUT Inverter_Layout_0.OUT.t4 VIN.t55 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X9 VOUT Inverter_Layout_0.OUT.t5 VIN.t54 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X10 VIN Inverter_Layout_0.OUT.t6 VOUT.t60 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X11 VOUT CLK.t4 VIN.t1 Inverter_Layout_0.VSS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X12 VIN CLK.t5 VOUT.t15 Inverter_Layout_0.VSS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X13 VIN Inverter_Layout_0.OUT.t7 VOUT.t59 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X14 VIN Inverter_Layout_0.OUT.t8 VOUT.t58 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X15 VIN CLK.t6 VOUT.t6 Inverter_Layout_0.VSS nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X16 VOUT CLK.t7 VIN.t68 Inverter_Layout_0.VSS nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X17 VOUT Inverter_Layout_0.OUT.t9 VIN.t53 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X18 VOUT Inverter_Layout_0.OUT.t10 VIN.t52 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X19 VOUT Inverter_Layout_0.OUT.t11 VIN.t51 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X20 VOUT Inverter_Layout_0.OUT.t12 VIN.t50 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X21 VIN Inverter_Layout_0.OUT.t13 VOUT.t53 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X22 VIN Inverter_Layout_0.OUT.t14 VOUT.t52 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X23 VIN CLK.t8 VOUT.t4 Inverter_Layout_0.VSS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X24 VIN Inverter_Layout_0.OUT.t15 VOUT.t51 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X25 VOUT CLK.t9 VIN.t67 Inverter_Layout_0.VSS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X26 VOUT Inverter_Layout_0.OUT.t16 VIN.t49 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X27 VIN Inverter_Layout_0.OUT.t17 VOUT.t49 Inverter_Layout_0.VDD pfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X28 VIN Inverter_Layout_0.OUT.t18 VOUT.t48 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X29 VIN CLK.t10 VOUT.t14 Inverter_Layout_0.VSS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X30 VOUT Inverter_Layout_0.OUT.t19 VIN.t48 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X31 VOUT Inverter_Layout_0.OUT.t20 VIN.t47 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X32 VOUT CLK.t11 VIN.t5 Inverter_Layout_0.VSS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X33 Inverter_Layout_0.VDD CLK.t12 Inverter_Layout_0.OUT Inverter_Layout_0.VDD pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X34 VIN Inverter_Layout_0.OUT.t21 VOUT.t45 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X35 VIN CLK.t13 VOUT.t2 Inverter_Layout_0.VSS nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X36 VOUT CLK.t14 VIN.t0 Inverter_Layout_0.VSS nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X37 VOUT Inverter_Layout_0.OUT.t22 VIN.t46 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X38 VIN Inverter_Layout_0.OUT.t23 VOUT.t43 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X39 VIN Inverter_Layout_0.OUT.t24 VOUT.t42 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X40 VIN Inverter_Layout_0.OUT.t25 VOUT.t41 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X41 VOUT Inverter_Layout_0.OUT.t26 VIN.t45 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X42 VOUT Inverter_Layout_0.OUT.t27 VIN.t44 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X43 VOUT Inverter_Layout_0.OUT.t28 VIN.t43 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X44 VOUT CLK.t15 VIN.t7 Inverter_Layout_0.VSS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X45 VIN CLK.t16 VOUT.t13 Inverter_Layout_0.VSS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X46 VOUT Inverter_Layout_0.OUT.t29 VIN.t42 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X47 VIN CLK.t17 VOUT.t18 Inverter_Layout_0.VSS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X48 VOUT CLK.t18 VIN.t69 Inverter_Layout_0.VSS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X49 VIN Inverter_Layout_0.OUT.t30 VOUT.t36 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X50 VIN Inverter_Layout_0.OUT.t31 VOUT.t35 Inverter_Layout_0.VDD pfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X51 VOUT Inverter_Layout_0.OUT.t32 VIN.t41 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X52 VIN CLK.t19 VOUT.t9 Inverter_Layout_0.VSS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X53 VIN Inverter_Layout_0.OUT.t33 VOUT.t33 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X54 VOUT CLK.t20 VIN.t10 Inverter_Layout_0.VSS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X55 VIN CLK.t21 VOUT.t3 Inverter_Layout_0.VSS nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X56 VOUT Inverter_Layout_0.OUT.t34 VIN.t40 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X57 VOUT Inverter_Layout_0.OUT.t35 VIN.t39 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X58 VIN Inverter_Layout_0.OUT.t36 VOUT.t30 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X59 VIN Inverter_Layout_0.OUT.t37 VOUT.t29 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X60 VIN Inverter_Layout_0.OUT.t38 VOUT.t28 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X61 VOUT Inverter_Layout_0.OUT.t39 VIN.t38 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X62 VOUT CLK.t22 VIN.t12 Inverter_Layout_0.VSS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X63 VIN Inverter_Layout_0.OUT.t40 VOUT.t26 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X64 VIN CLK.t23 VOUT.t11 Inverter_Layout_0.VSS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X65 VOUT Inverter_Layout_0.OUT.t41 VIN.t37 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X66 VOUT Inverter_Layout_0.OUT.t42 VIN.t36 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X67 VIN Inverter_Layout_0.OUT.t43 VOUT.t23 Inverter_Layout_0.VDD pfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X68 VOUT CLK.t24 VIN.t71 Inverter_Layout_0.VSS nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X69 VIN Inverter_Layout_0.OUT.t44 VOUT.t22 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X70 VOUT Inverter_Layout_0.OUT.t45 VIN.t35 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X71 VIN Inverter_Layout_0.OUT.t46 VOUT.t20 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X72 VIN Inverter_Layout_0.OUT.t47 VOUT.t19 Inverter_Layout_0.VDD pfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X73 VIN CLK.t25 VOUT.t17 Inverter_Layout_0.VSS nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
R0 Inverter_Layout_0.OUT.t2 Inverter_Layout_0.OUT.t18 50.3184
R1 Inverter_Layout_0.OUT.t40 Inverter_Layout_0.OUT.t2 50.3184
R2 Inverter_Layout_0.OUT.t35 Inverter_Layout_0.OUT.t3 50.3184
R3 Inverter_Layout_0.OUT.t29 Inverter_Layout_0.OUT.t35 50.3184
R4 Inverter_Layout_0.OUT.t24 Inverter_Layout_0.OUT.t36 50.3184
R5 Inverter_Layout_0.OUT.t15 Inverter_Layout_0.OUT.t24 50.3184
R6 Inverter_Layout_0.OUT.t22 Inverter_Layout_0.OUT.t34 50.3184
R7 Inverter_Layout_0.OUT.t10 Inverter_Layout_0.OUT.t22 50.3184
R8 Inverter_Layout_0.OUT.t7 Inverter_Layout_0.OUT.t21 50.3184
R9 Inverter_Layout_0.OUT.t44 Inverter_Layout_0.OUT.t7 50.3184
R10 Inverter_Layout_0.OUT.t5 Inverter_Layout_0.OUT.t20 50.3184
R11 Inverter_Layout_0.OUT.t42 Inverter_Layout_0.OUT.t5 50.3184
R12 Inverter_Layout_0.OUT.t38 Inverter_Layout_0.OUT.t6 50.3184
R13 Inverter_Layout_0.OUT.t30 Inverter_Layout_0.OUT.t38 50.3184
R14 Inverter_Layout_0.OUT.t28 Inverter_Layout_0.OUT.t39 50.3184
R15 Inverter_Layout_0.OUT.t16 Inverter_Layout_0.OUT.t28 50.3184
R16 Inverter_Layout_0.OUT.t25 Inverter_Layout_0.OUT.t37 50.3184
R17 Inverter_Layout_0.OUT.t14 Inverter_Layout_0.OUT.t25 50.3184
R18 Inverter_Layout_0.OUT.t11 Inverter_Layout_0.OUT.t26 50.3184
R19 Inverter_Layout_0.OUT.t0 Inverter_Layout_0.OUT.t11 50.3184
R20 Inverter_Layout_0.OUT.t8 Inverter_Layout_0.OUT.t23 50.3184
R21 Inverter_Layout_0.OUT.t46 Inverter_Layout_0.OUT.t8 50.3184
R22 Inverter_Layout_0.OUT.t12 Inverter_Layout_0.OUT.t27 50.3184
R23 Inverter_Layout_0.OUT.t1 Inverter_Layout_0.OUT.t12 50.3184
R24 Inverter_Layout_0.OUT.t47 Inverter_Layout_0.OUT.t13 50.3184
R25 Inverter_Layout_0.OUT.t33 Inverter_Layout_0.OUT.t47 50.3184
R26 Inverter_Layout_0.OUT.t45 Inverter_Layout_0.OUT.t9 50.3184
R27 Inverter_Layout_0.OUT.t32 Inverter_Layout_0.OUT.t45 50.3184
R28 Inverter_Layout_0.OUT.t31 Inverter_Layout_0.OUT.t43 50.3184
R29 Inverter_Layout_0.OUT.t17 Inverter_Layout_0.OUT.t31 50.3184
R30 Inverter_Layout_0.OUT.t4 Inverter_Layout_0.OUT.t41 50.3184
R31 Inverter_Layout_0.OUT.t19 Inverter_Layout_0.OUT.t4 50.3184
R32 Inverter_Layout_0.OUT Inverter_Layout_0.OUT.t19 49.2314
R33 Inverter_Layout_0.OUT.n0 Inverter_Layout_0.OUT.t17 39.7594
R34 Inverter_Layout_0.OUT.t41 Inverter_Layout_0.OUT.n13 39.7594
R35 Inverter_Layout_0.OUT.n1 Inverter_Layout_0.OUT.n0 20.8576
R36 Inverter_Layout_0.OUT.n2 Inverter_Layout_0.OUT.n1 20.8576
R37 Inverter_Layout_0.OUT.n3 Inverter_Layout_0.OUT.n2 20.8576
R38 Inverter_Layout_0.OUT.n4 Inverter_Layout_0.OUT.n3 20.8576
R39 Inverter_Layout_0.OUT.n5 Inverter_Layout_0.OUT.n4 20.8576
R40 Inverter_Layout_0.OUT.n6 Inverter_Layout_0.OUT.n5 20.8576
R41 Inverter_Layout_0.OUT.n7 Inverter_Layout_0.OUT.n6 20.8576
R42 Inverter_Layout_0.OUT.n8 Inverter_Layout_0.OUT.n7 20.8576
R43 Inverter_Layout_0.OUT.n9 Inverter_Layout_0.OUT.n8 20.8576
R44 Inverter_Layout_0.OUT.n10 Inverter_Layout_0.OUT.n9 20.8576
R45 Inverter_Layout_0.OUT.n11 Inverter_Layout_0.OUT.n10 20.8576
R46 Inverter_Layout_0.OUT.n12 Inverter_Layout_0.OUT.n11 20.8576
R47 Inverter_Layout_0.OUT.n13 Inverter_Layout_0.OUT.n12 20.8576
R48 Inverter_Layout_0.OUT.n13 Inverter_Layout_0.OUT.t40 18.9023
R49 Inverter_Layout_0.OUT.n12 Inverter_Layout_0.OUT.t29 18.9023
R50 Inverter_Layout_0.OUT.n11 Inverter_Layout_0.OUT.t15 18.9023
R51 Inverter_Layout_0.OUT.n10 Inverter_Layout_0.OUT.t10 18.9023
R52 Inverter_Layout_0.OUT.n9 Inverter_Layout_0.OUT.t44 18.9023
R53 Inverter_Layout_0.OUT.n8 Inverter_Layout_0.OUT.t42 18.9023
R54 Inverter_Layout_0.OUT.n7 Inverter_Layout_0.OUT.t30 18.9023
R55 Inverter_Layout_0.OUT.n6 Inverter_Layout_0.OUT.t16 18.9023
R56 Inverter_Layout_0.OUT.n5 Inverter_Layout_0.OUT.t14 18.9023
R57 Inverter_Layout_0.OUT.n4 Inverter_Layout_0.OUT.t0 18.9023
R58 Inverter_Layout_0.OUT.n3 Inverter_Layout_0.OUT.t46 18.9023
R59 Inverter_Layout_0.OUT.n2 Inverter_Layout_0.OUT.t1 18.9023
R60 Inverter_Layout_0.OUT.n1 Inverter_Layout_0.OUT.t33 18.9023
R61 Inverter_Layout_0.OUT.n0 Inverter_Layout_0.OUT.t32 18.9023
R62 VIN.n73 VIN.n72 4.81172
R63 VIN.n104 VIN.n2 4.4609
R64 VIN.n105 VIN.n1 4.4609
R65 VIN.n106 VIN.n0 4.4609
R66 VIN.n100 VIN.t71 4.4609
R67 VIN.n101 VIN.t68 4.4609
R68 VIN.n102 VIN.t0 4.4609
R69 VIN.n95 VIN.t37 4.0565
R70 VIN.n96 VIN.t55 4.0565
R71 VIN.n97 VIN.t48 4.0565
R72 VIN.n74 VIN.n70 4.0565
R73 VIN.n73 VIN.n71 4.0565
R74 VIN.n26 VIN.n25 3.90572
R75 VIN.n9 VIN.n8 3.90572
R76 VIN.n32 VIN.n29 3.35572
R77 VIN.n46 VIN.n43 3.35572
R78 VIN.n86 VIN.n83 3.35572
R79 VIN.n63 VIN.n60 3.35572
R80 VIN.n26 VIN.n23 3.1505
R81 VIN.n27 VIN.n21 3.1505
R82 VIN.n9 VIN.n6 3.1505
R83 VIN.n10 VIN.n4 3.1505
R84 VIN.n13 VIN.n12 3.1505
R85 VIN.n16 VIN.n15 3.1505
R86 VIN.n19 VIN.n18 3.1505
R87 VIN.n32 VIN.n31 2.6005
R88 VIN.n35 VIN.n34 2.6005
R89 VIN.n46 VIN.n45 2.6005
R90 VIN.n49 VIN.n48 2.6005
R91 VIN.n50 VIN.n41 2.6005
R92 VIN.n51 VIN.n39 2.6005
R93 VIN.n52 VIN.n37 2.6005
R94 VIN.n86 VIN.n85 2.6005
R95 VIN.n89 VIN.n88 2.6005
R96 VIN.n63 VIN.n62 2.6005
R97 VIN.n66 VIN.n65 2.6005
R98 VIN.n67 VIN.n58 2.6005
R99 VIN.n68 VIN.n56 2.6005
R100 VIN.n69 VIN.n54 2.6005
R101 VIN.n90 VIN.n81 2.6005
R102 VIN.n91 VIN.n79 2.6005
R103 VIN.n92 VIN.n77 2.6005
R104 VIN.n95 VIN.n94 2.47941
R105 VIN.n103 VIN.n102 2.47941
R106 VIN.n93 VIN.n75 2.05876
R107 VIN.n34 VIN.t56 1.4565
R108 VIN.n34 VIN.n33 1.4565
R109 VIN.n31 VIN.t39 1.4565
R110 VIN.n31 VIN.n30 1.4565
R111 VIN.n29 VIN.t42 1.4565
R112 VIN.n29 VIN.n28 1.4565
R113 VIN.n37 VIN.t36 1.4565
R114 VIN.n37 VIN.n36 1.4565
R115 VIN.n39 VIN.t54 1.4565
R116 VIN.n39 VIN.n38 1.4565
R117 VIN.n41 VIN.t47 1.4565
R118 VIN.n41 VIN.n40 1.4565
R119 VIN.n48 VIN.t40 1.4565
R120 VIN.n48 VIN.n47 1.4565
R121 VIN.n45 VIN.t46 1.4565
R122 VIN.n45 VIN.n44 1.4565
R123 VIN.n43 VIN.t52 1.4565
R124 VIN.n43 VIN.n42 1.4565
R125 VIN.n77 VIN.t49 1.4565
R126 VIN.n77 VIN.n76 1.4565
R127 VIN.n79 VIN.t43 1.4565
R128 VIN.n79 VIN.n78 1.4565
R129 VIN.n81 VIN.t38 1.4565
R130 VIN.n81 VIN.n80 1.4565
R131 VIN.n88 VIN.t45 1.4565
R132 VIN.n88 VIN.n87 1.4565
R133 VIN.n85 VIN.t51 1.4565
R134 VIN.n85 VIN.n84 1.4565
R135 VIN.n83 VIN.t58 1.4565
R136 VIN.n83 VIN.n82 1.4565
R137 VIN.n54 VIN.t41 1.4565
R138 VIN.n54 VIN.n53 1.4565
R139 VIN.n56 VIN.t35 1.4565
R140 VIN.n56 VIN.n55 1.4565
R141 VIN.n58 VIN.t53 1.4565
R142 VIN.n58 VIN.n57 1.4565
R143 VIN.n65 VIN.t44 1.4565
R144 VIN.n65 VIN.n64 1.4565
R145 VIN.n62 VIN.t50 1.4565
R146 VIN.n62 VIN.n61 1.4565
R147 VIN.n60 VIN.t57 1.4565
R148 VIN.n60 VIN.n59 1.4565
R149 VIN.n21 VIN.t7 1.3109
R150 VIN.n21 VIN.n20 1.3109
R151 VIN.n23 VIN.t12 1.3109
R152 VIN.n23 VIN.n22 1.3109
R153 VIN.n25 VIN.t1 1.3109
R154 VIN.n25 VIN.n24 1.3109
R155 VIN.n18 VIN.t69 1.3109
R156 VIN.n18 VIN.n17 1.3109
R157 VIN.n15 VIN.t67 1.3109
R158 VIN.n15 VIN.n14 1.3109
R159 VIN.n12 VIN.t8 1.3109
R160 VIN.n12 VIN.n11 1.3109
R161 VIN.n4 VIN.t5 1.3109
R162 VIN.n4 VIN.n3 1.3109
R163 VIN.n6 VIN.t10 1.3109
R164 VIN.n6 VIN.n5 1.3109
R165 VIN.n8 VIN.t16 1.3109
R166 VIN.n8 VIN.n7 1.3109
R167 VIN.n50 VIN.n49 1.28789
R168 VIN.n90 VIN.n89 1.28789
R169 VIN.n67 VIN.n66 1.28789
R170 VIN.n13 VIN.n10 1.28789
R171 VIN.n75 VIN.n74 0.957239
R172 VIN.n98 VIN.n97 0.957239
R173 VIN.n99 VIN.n27 0.957239
R174 VIN.n104 VIN.n103 0.957239
R175 VIN.n99 VIN.n98 0.896587
R176 VIN.n35 VIN.n32 0.755717
R177 VIN.n49 VIN.n46 0.755717
R178 VIN.n52 VIN.n51 0.755717
R179 VIN.n51 VIN.n50 0.755717
R180 VIN.n89 VIN.n86 0.755717
R181 VIN.n66 VIN.n63 0.755717
R182 VIN.n69 VIN.n68 0.755717
R183 VIN.n68 VIN.n67 0.755717
R184 VIN.n74 VIN.n73 0.755717
R185 VIN.n92 VIN.n91 0.755717
R186 VIN.n91 VIN.n90 0.755717
R187 VIN.n96 VIN.n95 0.755717
R188 VIN.n97 VIN.n96 0.755717
R189 VIN.n27 VIN.n26 0.755717
R190 VIN.n101 VIN.n100 0.755717
R191 VIN.n102 VIN.n101 0.755717
R192 VIN.n10 VIN.n9 0.755717
R193 VIN.n16 VIN.n13 0.755717
R194 VIN.n19 VIN.n16 0.755717
R195 VIN.n106 VIN.n105 0.755717
R196 VIN.n105 VIN.n104 0.755717
R197 VIN.n94 VIN.n93 0.626587
R198 VIN VIN.n106 0.513109
R199 VIN.n98 VIN.n35 0.331152
R200 VIN.n94 VIN.n52 0.331152
R201 VIN.n75 VIN.n69 0.331152
R202 VIN.n93 VIN.n92 0.331152
R203 VIN.n100 VIN.n99 0.331152
R204 VIN.n103 VIN.n19 0.331152
R205 VOUT.n40 VOUT.n39 3.90572
R206 VOUT.n60 VOUT.n57 3.90572
R207 VOUT.n68 VOUT.n65 3.90572
R208 VOUT.n4 VOUT.n1 3.35572
R209 VOUT.n22 VOUT.n21 3.35572
R210 VOUT.n14 VOUT.n13 3.35572
R211 VOUT.n46 VOUT.n43 3.35572
R212 VOUT.n90 VOUT.n89 3.35572
R213 VOUT.n82 VOUT.n81 3.35572
R214 VOUT.n40 VOUT.n37 3.1505
R215 VOUT.n41 VOUT.n35 3.1505
R216 VOUT.n60 VOUT.n59 3.1505
R217 VOUT.n63 VOUT.n62 3.1505
R218 VOUT.n68 VOUT.n67 3.1505
R219 VOUT.n71 VOUT.n70 3.1505
R220 VOUT.n73 VOUT.n55 3.1505
R221 VOUT.n74 VOUT.n53 3.1505
R222 VOUT.n75 VOUT.n51 3.1505
R223 VOUT.n4 VOUT.n3 2.6005
R224 VOUT.n7 VOUT.n6 2.6005
R225 VOUT.n22 VOUT.n19 2.6005
R226 VOUT.n23 VOUT.n17 2.6005
R227 VOUT.n14 VOUT.n11 2.6005
R228 VOUT.n15 VOUT.n9 2.6005
R229 VOUT.n27 VOUT.n26 2.6005
R230 VOUT.n30 VOUT.n29 2.6005
R231 VOUT.n33 VOUT.n32 2.6005
R232 VOUT.n46 VOUT.n45 2.6005
R233 VOUT.n49 VOUT.n48 2.6005
R234 VOUT.n90 VOUT.n87 2.6005
R235 VOUT.n91 VOUT.n85 2.6005
R236 VOUT.n82 VOUT.n79 2.6005
R237 VOUT.n83 VOUT.n77 2.6005
R238 VOUT.n101 VOUT.n100 2.6005
R239 VOUT.n98 VOUT.n97 2.6005
R240 VOUT.n95 VOUT.n94 2.6005
R241 VOUT.n102 VOUT.n101 1.76333
R242 VOUT.n6 VOUT.t23 1.4565
R243 VOUT.n6 VOUT.n5 1.4565
R244 VOUT.n3 VOUT.t35 1.4565
R245 VOUT.n3 VOUT.n2 1.4565
R246 VOUT.n1 VOUT.t49 1.4565
R247 VOUT.n1 VOUT.n0 1.4565
R248 VOUT.n32 VOUT.t43 1.4565
R249 VOUT.n32 VOUT.n31 1.4565
R250 VOUT.n29 VOUT.t58 1.4565
R251 VOUT.n29 VOUT.n28 1.4565
R252 VOUT.n26 VOUT.t20 1.4565
R253 VOUT.n26 VOUT.n25 1.4565
R254 VOUT.n17 VOUT.t52 1.4565
R255 VOUT.n17 VOUT.n16 1.4565
R256 VOUT.n19 VOUT.t41 1.4565
R257 VOUT.n19 VOUT.n18 1.4565
R258 VOUT.n21 VOUT.t29 1.4565
R259 VOUT.n21 VOUT.n20 1.4565
R260 VOUT.n9 VOUT.t33 1.4565
R261 VOUT.n9 VOUT.n8 1.4565
R262 VOUT.n11 VOUT.t19 1.4565
R263 VOUT.n11 VOUT.n10 1.4565
R264 VOUT.n13 VOUT.t53 1.4565
R265 VOUT.n13 VOUT.n12 1.4565
R266 VOUT.n48 VOUT.t60 1.4565
R267 VOUT.n48 VOUT.n47 1.4565
R268 VOUT.n45 VOUT.t28 1.4565
R269 VOUT.n45 VOUT.n44 1.4565
R270 VOUT.n43 VOUT.t36 1.4565
R271 VOUT.n43 VOUT.n42 1.4565
R272 VOUT.n94 VOUT.t51 1.4565
R273 VOUT.n94 VOUT.n93 1.4565
R274 VOUT.n97 VOUT.t42 1.4565
R275 VOUT.n97 VOUT.n96 1.4565
R276 VOUT.n100 VOUT.t30 1.4565
R277 VOUT.n100 VOUT.n99 1.4565
R278 VOUT.n85 VOUT.t26 1.4565
R279 VOUT.n85 VOUT.n84 1.4565
R280 VOUT.n87 VOUT.t64 1.4565
R281 VOUT.n87 VOUT.n86 1.4565
R282 VOUT.n89 VOUT.t48 1.4565
R283 VOUT.n89 VOUT.n88 1.4565
R284 VOUT.n77 VOUT.t22 1.4565
R285 VOUT.n77 VOUT.n76 1.4565
R286 VOUT.n79 VOUT.t59 1.4565
R287 VOUT.n79 VOUT.n78 1.4565
R288 VOUT.n81 VOUT.t45 1.4565
R289 VOUT.n81 VOUT.n80 1.4565
R290 VOUT.n35 VOUT.t6 1.3109
R291 VOUT.n35 VOUT.n34 1.3109
R292 VOUT.n37 VOUT.t2 1.3109
R293 VOUT.n37 VOUT.n36 1.3109
R294 VOUT.n39 VOUT.t3 1.3109
R295 VOUT.n39 VOUT.n38 1.3109
R296 VOUT.n51 VOUT.t70 1.3109
R297 VOUT.n51 VOUT.n50 1.3109
R298 VOUT.n53 VOUT.t4 1.3109
R299 VOUT.n53 VOUT.n52 1.3109
R300 VOUT.n55 VOUT.t13 1.3109
R301 VOUT.n55 VOUT.n54 1.3109
R302 VOUT.n62 VOUT.t15 1.3109
R303 VOUT.n62 VOUT.n61 1.3109
R304 VOUT.n59 VOUT.t11 1.3109
R305 VOUT.n59 VOUT.n58 1.3109
R306 VOUT.n57 VOUT.t18 1.3109
R307 VOUT.n57 VOUT.n56 1.3109
R308 VOUT.n70 VOUT.t17 1.3109
R309 VOUT.n70 VOUT.n69 1.3109
R310 VOUT.n67 VOUT.t9 1.3109
R311 VOUT.n67 VOUT.n66 1.3109
R312 VOUT.n65 VOUT.t14 1.3109
R313 VOUT.n65 VOUT.n64 1.3109
R314 VOUT.n104 VOUT.n103 1.25267
R315 VOUT.n103 VOUT.n102 1.25267
R316 VOUT.n24 VOUT.n23 0.957239
R317 VOUT.n24 VOUT.n15 0.957239
R318 VOUT.n72 VOUT.n63 0.957239
R319 VOUT.n72 VOUT.n71 0.957239
R320 VOUT.n92 VOUT.n91 0.957239
R321 VOUT.n92 VOUT.n83 0.957239
R322 VOUT.n7 VOUT.n4 0.755717
R323 VOUT.n23 VOUT.n22 0.755717
R324 VOUT.n15 VOUT.n14 0.755717
R325 VOUT.n30 VOUT.n27 0.755717
R326 VOUT.n33 VOUT.n30 0.755717
R327 VOUT.n41 VOUT.n40 0.755717
R328 VOUT.n63 VOUT.n60 0.755717
R329 VOUT.n71 VOUT.n68 0.755717
R330 VOUT.n49 VOUT.n46 0.755717
R331 VOUT.n75 VOUT.n74 0.755717
R332 VOUT.n74 VOUT.n73 0.755717
R333 VOUT.n91 VOUT.n90 0.755717
R334 VOUT.n83 VOUT.n82 0.755717
R335 VOUT.n98 VOUT.n95 0.755717
R336 VOUT.n101 VOUT.n98 0.755717
R337 VOUT.n104 VOUT.n7 0.511152
R338 VOUT.n103 VOUT.n33 0.511152
R339 VOUT.n103 VOUT.n41 0.511152
R340 VOUT.n102 VOUT.n49 0.511152
R341 VOUT.n102 VOUT.n75 0.511152
R342 VOUT.n27 VOUT.n24 0.331152
R343 VOUT.n73 VOUT.n72 0.331152
R344 VOUT.n95 VOUT.n92 0.331152
R345 VOUT VOUT.n104 0.0885435
R346 CLK.t13 CLK.t6 50.3184
R347 CLK.t21 CLK.t13 50.3184
R348 CLK.t9 CLK.t1 50.3184
R349 CLK.t18 CLK.t9 50.3184
R350 CLK.t23 CLK.t17 50.3184
R351 CLK.t5 CLK.t23 50.3184
R352 CLK.t20 CLK.t11 50.3184
R353 CLK.t2 CLK.t20 50.3184
R354 CLK.t8 CLK.t0 50.3184
R355 CLK.t16 CLK.t8 50.3184
R356 CLK.t22 CLK.t15 50.3184
R357 CLK.t4 CLK.t22 50.3184
R358 CLK.t19 CLK.t10 50.3184
R359 CLK.t25 CLK.t19 50.3184
R360 CLK.t7 CLK.t24 50.3184
R361 CLK.t14 CLK.t7 50.3184
R362 CLK CLK.n6 48.0321
R363 CLK.n0 CLK.t21 39.7594
R364 CLK.n7 CLK.t12 34.6755
R365 CLK.n1 CLK.n0 20.8576
R366 CLK.n2 CLK.n1 20.8576
R367 CLK.n3 CLK.n2 20.8576
R368 CLK.n4 CLK.n3 20.8576
R369 CLK.n5 CLK.n4 20.8576
R370 CLK.n6 CLK.n5 20.8576
R371 CLK.n0 CLK.t18 18.9023
R372 CLK.n1 CLK.t5 18.9023
R373 CLK.n2 CLK.t2 18.9023
R374 CLK.n3 CLK.t16 18.9023
R375 CLK.n4 CLK.t4 18.9023
R376 CLK.n5 CLK.t25 18.9023
R377 CLK.n6 CLK.t14 18.9023
R378 CLK CLK.n7 17.6692
R379 CLK.n7 CLK.t3 13.0362
C0 VOUT CLK 0.318f
C1 Inverter_Layout_0.OUT Inverter_Layout_0.VDD 4.02f
C2 VOUT Inverter_Layout_0.VDD 0.379f
C3 VIN Inverter_Layout_0.OUT 0.755f
C4 VOUT VIN 15.9f
C5 CLK Inverter_Layout_0.VDD 0.198f
C6 VOUT Inverter_Layout_0.OUT 0.623f
C7 VIN CLK 0.543f
C8 CLK Inverter_Layout_0.OUT 0.0739f
C9 VIN Inverter_Layout_0.VDD 0.722f
C10 VOUT Inverter_Layout_0.VSS 1.1f
C11 VIN Inverter_Layout_0.VSS 2.77f
C12 CLK Inverter_Layout_0.VSS 3.37f
C13 Inverter_Layout_0.OUT Inverter_Layout_0.VSS 2.63f
C14 Inverter_Layout_0.VDD Inverter_Layout_0.VSS 12.3f
C15 VOUT.t49 Inverter_Layout_0.VSS 0.0592f
C16 VOUT.n0 Inverter_Layout_0.VSS 0.0592f
C17 VOUT.n1 Inverter_Layout_0.VSS 0.148f
C18 VOUT.t35 Inverter_Layout_0.VSS 0.0592f
C19 VOUT.n2 Inverter_Layout_0.VSS 0.0592f
C20 VOUT.n3 Inverter_Layout_0.VSS 0.118f
C21 VOUT.n4 Inverter_Layout_0.VSS 0.264f
C22 VOUT.t23 Inverter_Layout_0.VSS 0.0592f
C23 VOUT.n5 Inverter_Layout_0.VSS 0.0592f
C24 VOUT.n6 Inverter_Layout_0.VSS 0.118f
C25 VOUT.n7 Inverter_Layout_0.VSS 0.136f
C26 VOUT.t33 Inverter_Layout_0.VSS 0.0592f
C27 VOUT.n8 Inverter_Layout_0.VSS 0.0592f
C28 VOUT.n9 Inverter_Layout_0.VSS 0.118f
C29 VOUT.t19 Inverter_Layout_0.VSS 0.0592f
C30 VOUT.n10 Inverter_Layout_0.VSS 0.0592f
C31 VOUT.n11 Inverter_Layout_0.VSS 0.118f
C32 VOUT.t53 Inverter_Layout_0.VSS 0.0592f
C33 VOUT.n12 Inverter_Layout_0.VSS 0.0592f
C34 VOUT.n13 Inverter_Layout_0.VSS 0.148f
C35 VOUT.n14 Inverter_Layout_0.VSS 0.264f
C36 VOUT.n15 Inverter_Layout_0.VSS 0.19f
C37 VOUT.t52 Inverter_Layout_0.VSS 0.0592f
C38 VOUT.n16 Inverter_Layout_0.VSS 0.0592f
C39 VOUT.n17 Inverter_Layout_0.VSS 0.118f
C40 VOUT.t41 Inverter_Layout_0.VSS 0.0592f
C41 VOUT.n18 Inverter_Layout_0.VSS 0.0592f
C42 VOUT.n19 Inverter_Layout_0.VSS 0.118f
C43 VOUT.t29 Inverter_Layout_0.VSS 0.0592f
C44 VOUT.n20 Inverter_Layout_0.VSS 0.0592f
C45 VOUT.n21 Inverter_Layout_0.VSS 0.148f
C46 VOUT.n22 Inverter_Layout_0.VSS 0.264f
C47 VOUT.n23 Inverter_Layout_0.VSS 0.19f
C48 VOUT.n24 Inverter_Layout_0.VSS 0.247f
C49 VOUT.t20 Inverter_Layout_0.VSS 0.0592f
C50 VOUT.n25 Inverter_Layout_0.VSS 0.0592f
C51 VOUT.n26 Inverter_Layout_0.VSS 0.118f
C52 VOUT.n27 Inverter_Layout_0.VSS 0.116f
C53 VOUT.t58 Inverter_Layout_0.VSS 0.0592f
C54 VOUT.n28 Inverter_Layout_0.VSS 0.0592f
C55 VOUT.n29 Inverter_Layout_0.VSS 0.118f
C56 VOUT.n30 Inverter_Layout_0.VSS 0.162f
C57 VOUT.t43 Inverter_Layout_0.VSS 0.0592f
C58 VOUT.n31 Inverter_Layout_0.VSS 0.0592f
C59 VOUT.n32 Inverter_Layout_0.VSS 0.118f
C60 VOUT.n33 Inverter_Layout_0.VSS 0.136f
C61 VOUT.t6 Inverter_Layout_0.VSS 0.0592f
C62 VOUT.n34 Inverter_Layout_0.VSS 0.0592f
C63 VOUT.n35 Inverter_Layout_0.VSS 0.118f
C64 VOUT.t2 Inverter_Layout_0.VSS 0.0592f
C65 VOUT.n36 Inverter_Layout_0.VSS 0.0592f
C66 VOUT.n37 Inverter_Layout_0.VSS 0.118f
C67 VOUT.t3 Inverter_Layout_0.VSS 0.0592f
C68 VOUT.n38 Inverter_Layout_0.VSS 0.0592f
C69 VOUT.n39 Inverter_Layout_0.VSS 0.144f
C70 VOUT.n40 Inverter_Layout_0.VSS 0.269f
C71 VOUT.n41 Inverter_Layout_0.VSS 0.136f
C72 VOUT.t36 Inverter_Layout_0.VSS 0.0592f
C73 VOUT.n42 Inverter_Layout_0.VSS 0.0592f
C74 VOUT.n43 Inverter_Layout_0.VSS 0.148f
C75 VOUT.t28 Inverter_Layout_0.VSS 0.0592f
C76 VOUT.n44 Inverter_Layout_0.VSS 0.0592f
C77 VOUT.n45 Inverter_Layout_0.VSS 0.118f
C78 VOUT.n46 Inverter_Layout_0.VSS 0.264f
C79 VOUT.t60 Inverter_Layout_0.VSS 0.0592f
C80 VOUT.n47 Inverter_Layout_0.VSS 0.0592f
C81 VOUT.n48 Inverter_Layout_0.VSS 0.118f
C82 VOUT.n49 Inverter_Layout_0.VSS 0.136f
C83 VOUT.t70 Inverter_Layout_0.VSS 0.0592f
C84 VOUT.n50 Inverter_Layout_0.VSS 0.0592f
C85 VOUT.n51 Inverter_Layout_0.VSS 0.118f
C86 VOUT.t4 Inverter_Layout_0.VSS 0.0592f
C87 VOUT.n52 Inverter_Layout_0.VSS 0.0592f
C88 VOUT.n53 Inverter_Layout_0.VSS 0.118f
C89 VOUT.t13 Inverter_Layout_0.VSS 0.0592f
C90 VOUT.n54 Inverter_Layout_0.VSS 0.0592f
C91 VOUT.n55 Inverter_Layout_0.VSS 0.118f
C92 VOUT.t18 Inverter_Layout_0.VSS 0.0592f
C93 VOUT.n56 Inverter_Layout_0.VSS 0.0592f
C94 VOUT.n57 Inverter_Layout_0.VSS 0.144f
C95 VOUT.t11 Inverter_Layout_0.VSS 0.0592f
C96 VOUT.n58 Inverter_Layout_0.VSS 0.0592f
C97 VOUT.n59 Inverter_Layout_0.VSS 0.118f
C98 VOUT.n60 Inverter_Layout_0.VSS 0.269f
C99 VOUT.t15 Inverter_Layout_0.VSS 0.0592f
C100 VOUT.n61 Inverter_Layout_0.VSS 0.0592f
C101 VOUT.n62 Inverter_Layout_0.VSS 0.118f
C102 VOUT.n63 Inverter_Layout_0.VSS 0.19f
C103 VOUT.t14 Inverter_Layout_0.VSS 0.0592f
C104 VOUT.n64 Inverter_Layout_0.VSS 0.0592f
C105 VOUT.n65 Inverter_Layout_0.VSS 0.144f
C106 VOUT.t9 Inverter_Layout_0.VSS 0.0592f
C107 VOUT.n66 Inverter_Layout_0.VSS 0.0592f
C108 VOUT.n67 Inverter_Layout_0.VSS 0.118f
C109 VOUT.n68 Inverter_Layout_0.VSS 0.269f
C110 VOUT.t17 Inverter_Layout_0.VSS 0.0592f
C111 VOUT.n69 Inverter_Layout_0.VSS 0.0592f
C112 VOUT.n70 Inverter_Layout_0.VSS 0.118f
C113 VOUT.n71 Inverter_Layout_0.VSS 0.19f
C114 VOUT.n72 Inverter_Layout_0.VSS 0.247f
C115 VOUT.n73 Inverter_Layout_0.VSS 0.116f
C116 VOUT.n74 Inverter_Layout_0.VSS 0.162f
C117 VOUT.n75 Inverter_Layout_0.VSS 0.136f
C118 VOUT.t22 Inverter_Layout_0.VSS 0.0592f
C119 VOUT.n76 Inverter_Layout_0.VSS 0.0592f
C120 VOUT.n77 Inverter_Layout_0.VSS 0.118f
C121 VOUT.t59 Inverter_Layout_0.VSS 0.0592f
C122 VOUT.n78 Inverter_Layout_0.VSS 0.0592f
C123 VOUT.n79 Inverter_Layout_0.VSS 0.118f
C124 VOUT.t45 Inverter_Layout_0.VSS 0.0592f
C125 VOUT.n80 Inverter_Layout_0.VSS 0.0592f
C126 VOUT.n81 Inverter_Layout_0.VSS 0.148f
C127 VOUT.n82 Inverter_Layout_0.VSS 0.264f
C128 VOUT.n83 Inverter_Layout_0.VSS 0.19f
C129 VOUT.t26 Inverter_Layout_0.VSS 0.0592f
C130 VOUT.n84 Inverter_Layout_0.VSS 0.0592f
C131 VOUT.n85 Inverter_Layout_0.VSS 0.118f
C132 VOUT.t64 Inverter_Layout_0.VSS 0.0592f
C133 VOUT.n86 Inverter_Layout_0.VSS 0.0592f
C134 VOUT.n87 Inverter_Layout_0.VSS 0.118f
C135 VOUT.t48 Inverter_Layout_0.VSS 0.0592f
C136 VOUT.n88 Inverter_Layout_0.VSS 0.0592f
C137 VOUT.n89 Inverter_Layout_0.VSS 0.148f
C138 VOUT.n90 Inverter_Layout_0.VSS 0.264f
C139 VOUT.n91 Inverter_Layout_0.VSS 0.19f
C140 VOUT.n92 Inverter_Layout_0.VSS 0.247f
C141 VOUT.t51 Inverter_Layout_0.VSS 0.0592f
C142 VOUT.n93 Inverter_Layout_0.VSS 0.0592f
C143 VOUT.n94 Inverter_Layout_0.VSS 0.118f
C144 VOUT.n95 Inverter_Layout_0.VSS 0.116f
C145 VOUT.t42 Inverter_Layout_0.VSS 0.0592f
C146 VOUT.n96 Inverter_Layout_0.VSS 0.0592f
C147 VOUT.n97 Inverter_Layout_0.VSS 0.118f
C148 VOUT.n98 Inverter_Layout_0.VSS 0.162f
C149 VOUT.t30 Inverter_Layout_0.VSS 0.0592f
C150 VOUT.n99 Inverter_Layout_0.VSS 0.0592f
C151 VOUT.n100 Inverter_Layout_0.VSS 0.118f
C152 VOUT.n101 Inverter_Layout_0.VSS 0.277f
C153 VOUT.n102 Inverter_Layout_0.VSS 0.435f
C154 VOUT.n103 Inverter_Layout_0.VSS 0.378f
C155 VOUT.n104 Inverter_Layout_0.VSS 0.198f
C156 VIN.n0 Inverter_Layout_0.VSS 0.133f
C157 VIN.n1 Inverter_Layout_0.VSS 0.133f
C158 VIN.n2 Inverter_Layout_0.VSS 0.133f
C159 VIN.t5 Inverter_Layout_0.VSS 0.0496f
C160 VIN.n3 Inverter_Layout_0.VSS 0.0496f
C161 VIN.n4 Inverter_Layout_0.VSS 0.0993f
C162 VIN.t10 Inverter_Layout_0.VSS 0.0496f
C163 VIN.n5 Inverter_Layout_0.VSS 0.0496f
C164 VIN.n6 Inverter_Layout_0.VSS 0.0993f
C165 VIN.t16 Inverter_Layout_0.VSS 0.0496f
C166 VIN.n7 Inverter_Layout_0.VSS 0.0496f
C167 VIN.n8 Inverter_Layout_0.VSS 0.121f
C168 VIN.n9 Inverter_Layout_0.VSS 0.225f
C169 VIN.n10 Inverter_Layout_0.VSS 0.191f
C170 VIN.t8 Inverter_Layout_0.VSS 0.0496f
C171 VIN.n11 Inverter_Layout_0.VSS 0.0496f
C172 VIN.n12 Inverter_Layout_0.VSS 0.0993f
C173 VIN.n13 Inverter_Layout_0.VSS 0.191f
C174 VIN.t67 Inverter_Layout_0.VSS 0.0496f
C175 VIN.n14 Inverter_Layout_0.VSS 0.0496f
C176 VIN.n15 Inverter_Layout_0.VSS 0.0993f
C177 VIN.n16 Inverter_Layout_0.VSS 0.136f
C178 VIN.t69 Inverter_Layout_0.VSS 0.0496f
C179 VIN.n17 Inverter_Layout_0.VSS 0.0496f
C180 VIN.n18 Inverter_Layout_0.VSS 0.0993f
C181 VIN.n19 Inverter_Layout_0.VSS 0.0975f
C182 VIN.t7 Inverter_Layout_0.VSS 0.0496f
C183 VIN.n20 Inverter_Layout_0.VSS 0.0496f
C184 VIN.n21 Inverter_Layout_0.VSS 0.0993f
C185 VIN.t12 Inverter_Layout_0.VSS 0.0496f
C186 VIN.n22 Inverter_Layout_0.VSS 0.0496f
C187 VIN.n23 Inverter_Layout_0.VSS 0.0993f
C188 VIN.t1 Inverter_Layout_0.VSS 0.0496f
C189 VIN.n24 Inverter_Layout_0.VSS 0.0496f
C190 VIN.n25 Inverter_Layout_0.VSS 0.121f
C191 VIN.n26 Inverter_Layout_0.VSS 0.225f
C192 VIN.n27 Inverter_Layout_0.VSS 0.159f
C193 VIN.t42 Inverter_Layout_0.VSS 0.0496f
C194 VIN.n28 Inverter_Layout_0.VSS 0.0496f
C195 VIN.n29 Inverter_Layout_0.VSS 0.124f
C196 VIN.t39 Inverter_Layout_0.VSS 0.0496f
C197 VIN.n30 Inverter_Layout_0.VSS 0.0496f
C198 VIN.n31 Inverter_Layout_0.VSS 0.0993f
C199 VIN.n32 Inverter_Layout_0.VSS 0.222f
C200 VIN.t56 Inverter_Layout_0.VSS 0.0496f
C201 VIN.n33 Inverter_Layout_0.VSS 0.0496f
C202 VIN.n34 Inverter_Layout_0.VSS 0.0993f
C203 VIN.n35 Inverter_Layout_0.VSS 0.0975f
C204 VIN.t36 Inverter_Layout_0.VSS 0.0496f
C205 VIN.n36 Inverter_Layout_0.VSS 0.0496f
C206 VIN.n37 Inverter_Layout_0.VSS 0.0993f
C207 VIN.t54 Inverter_Layout_0.VSS 0.0496f
C208 VIN.n38 Inverter_Layout_0.VSS 0.0496f
C209 VIN.n39 Inverter_Layout_0.VSS 0.0993f
C210 VIN.t47 Inverter_Layout_0.VSS 0.0496f
C211 VIN.n40 Inverter_Layout_0.VSS 0.0496f
C212 VIN.n41 Inverter_Layout_0.VSS 0.0993f
C213 VIN.t52 Inverter_Layout_0.VSS 0.0496f
C214 VIN.n42 Inverter_Layout_0.VSS 0.0496f
C215 VIN.n43 Inverter_Layout_0.VSS 0.124f
C216 VIN.t46 Inverter_Layout_0.VSS 0.0496f
C217 VIN.n44 Inverter_Layout_0.VSS 0.0496f
C218 VIN.n45 Inverter_Layout_0.VSS 0.0993f
C219 VIN.n46 Inverter_Layout_0.VSS 0.222f
C220 VIN.t40 Inverter_Layout_0.VSS 0.0496f
C221 VIN.n47 Inverter_Layout_0.VSS 0.0496f
C222 VIN.n48 Inverter_Layout_0.VSS 0.0993f
C223 VIN.n49 Inverter_Layout_0.VSS 0.191f
C224 VIN.n50 Inverter_Layout_0.VSS 0.191f
C225 VIN.n51 Inverter_Layout_0.VSS 0.136f
C226 VIN.n52 Inverter_Layout_0.VSS 0.0975f
C227 VIN.t41 Inverter_Layout_0.VSS 0.0496f
C228 VIN.n53 Inverter_Layout_0.VSS 0.0496f
C229 VIN.n54 Inverter_Layout_0.VSS 0.0993f
C230 VIN.t35 Inverter_Layout_0.VSS 0.0496f
C231 VIN.n55 Inverter_Layout_0.VSS 0.0496f
C232 VIN.n56 Inverter_Layout_0.VSS 0.0993f
C233 VIN.t53 Inverter_Layout_0.VSS 0.0496f
C234 VIN.n57 Inverter_Layout_0.VSS 0.0496f
C235 VIN.n58 Inverter_Layout_0.VSS 0.0993f
C236 VIN.t57 Inverter_Layout_0.VSS 0.0496f
C237 VIN.n59 Inverter_Layout_0.VSS 0.0496f
C238 VIN.n60 Inverter_Layout_0.VSS 0.124f
C239 VIN.t50 Inverter_Layout_0.VSS 0.0496f
C240 VIN.n61 Inverter_Layout_0.VSS 0.0496f
C241 VIN.n62 Inverter_Layout_0.VSS 0.0993f
C242 VIN.n63 Inverter_Layout_0.VSS 0.222f
C243 VIN.t44 Inverter_Layout_0.VSS 0.0496f
C244 VIN.n64 Inverter_Layout_0.VSS 0.0496f
C245 VIN.n65 Inverter_Layout_0.VSS 0.0993f
C246 VIN.n66 Inverter_Layout_0.VSS 0.192f
C247 VIN.n67 Inverter_Layout_0.VSS 0.192f
C248 VIN.n68 Inverter_Layout_0.VSS 0.136f
C249 VIN.n69 Inverter_Layout_0.VSS 0.0975f
C250 VIN.n70 Inverter_Layout_0.VSS 0.126f
C251 VIN.n71 Inverter_Layout_0.VSS 0.126f
C252 VIN.n72 Inverter_Layout_0.VSS 0.15f
C253 VIN.n73 Inverter_Layout_0.VSS 0.307f
C254 VIN.n74 Inverter_Layout_0.VSS 0.201f
C255 VIN.n75 Inverter_Layout_0.VSS 0.319f
C256 VIN.t49 Inverter_Layout_0.VSS 0.0496f
C257 VIN.n76 Inverter_Layout_0.VSS 0.0496f
C258 VIN.n77 Inverter_Layout_0.VSS 0.0993f
C259 VIN.t43 Inverter_Layout_0.VSS 0.0496f
C260 VIN.n78 Inverter_Layout_0.VSS 0.0496f
C261 VIN.n79 Inverter_Layout_0.VSS 0.0993f
C262 VIN.t38 Inverter_Layout_0.VSS 0.0496f
C263 VIN.n80 Inverter_Layout_0.VSS 0.0496f
C264 VIN.n81 Inverter_Layout_0.VSS 0.0993f
C265 VIN.t58 Inverter_Layout_0.VSS 0.0496f
C266 VIN.n82 Inverter_Layout_0.VSS 0.0496f
C267 VIN.n83 Inverter_Layout_0.VSS 0.124f
C268 VIN.t51 Inverter_Layout_0.VSS 0.0496f
C269 VIN.n84 Inverter_Layout_0.VSS 0.0496f
C270 VIN.n85 Inverter_Layout_0.VSS 0.0993f
C271 VIN.n86 Inverter_Layout_0.VSS 0.222f
C272 VIN.t45 Inverter_Layout_0.VSS 0.0496f
C273 VIN.n87 Inverter_Layout_0.VSS 0.0496f
C274 VIN.n88 Inverter_Layout_0.VSS 0.0993f
C275 VIN.n89 Inverter_Layout_0.VSS 0.191f
C276 VIN.n90 Inverter_Layout_0.VSS 0.191f
C277 VIN.n91 Inverter_Layout_0.VSS 0.136f
C278 VIN.n92 Inverter_Layout_0.VSS 0.0975f
C279 VIN.n93 Inverter_Layout_0.VSS 0.287f
C280 VIN.n94 Inverter_Layout_0.VSS 0.326f
C281 VIN.t37 Inverter_Layout_0.VSS 0.126f
C282 VIN.n95 Inverter_Layout_0.VSS 0.34f
C283 VIN.t55 Inverter_Layout_0.VSS 0.126f
C284 VIN.n96 Inverter_Layout_0.VSS 0.178f
C285 VIN.t48 Inverter_Layout_0.VSS 0.126f
C286 VIN.n97 Inverter_Layout_0.VSS 0.201f
C287 VIN.n98 Inverter_Layout_0.VSS 0.213f
C288 VIN.n99 Inverter_Layout_0.VSS 0.201f
C289 VIN.t71 Inverter_Layout_0.VSS 0.133f
C290 VIN.n100 Inverter_Layout_0.VSS 0.132f
C291 VIN.t68 Inverter_Layout_0.VSS 0.133f
C292 VIN.n101 Inverter_Layout_0.VSS 0.17f
C293 VIN.t0 Inverter_Layout_0.VSS 0.133f
C294 VIN.n102 Inverter_Layout_0.VSS 0.332f
C295 VIN.n103 Inverter_Layout_0.VSS 0.358f
C296 VIN.n104 Inverter_Layout_0.VSS 0.194f
C297 VIN.n105 Inverter_Layout_0.VSS 0.17f
C298 VIN.n106 Inverter_Layout_0.VSS 0.152f
C299 Inverter_Layout_0.OUT.t18 Inverter_Layout_0.VSS 0.0535f
C300 Inverter_Layout_0.OUT.t2 Inverter_Layout_0.VSS 0.0754f
C301 Inverter_Layout_0.OUT.t40 Inverter_Layout_0.VSS 0.0518f
C302 Inverter_Layout_0.OUT.t3 Inverter_Layout_0.VSS 0.0535f
C303 Inverter_Layout_0.OUT.t35 Inverter_Layout_0.VSS 0.0754f
C304 Inverter_Layout_0.OUT.t29 Inverter_Layout_0.VSS 0.0518f
C305 Inverter_Layout_0.OUT.t36 Inverter_Layout_0.VSS 0.0535f
C306 Inverter_Layout_0.OUT.t24 Inverter_Layout_0.VSS 0.0754f
C307 Inverter_Layout_0.OUT.t15 Inverter_Layout_0.VSS 0.0518f
C308 Inverter_Layout_0.OUT.t34 Inverter_Layout_0.VSS 0.0535f
C309 Inverter_Layout_0.OUT.t22 Inverter_Layout_0.VSS 0.0754f
C310 Inverter_Layout_0.OUT.t10 Inverter_Layout_0.VSS 0.0518f
C311 Inverter_Layout_0.OUT.t21 Inverter_Layout_0.VSS 0.0535f
C312 Inverter_Layout_0.OUT.t7 Inverter_Layout_0.VSS 0.0754f
C313 Inverter_Layout_0.OUT.t44 Inverter_Layout_0.VSS 0.0518f
C314 Inverter_Layout_0.OUT.t20 Inverter_Layout_0.VSS 0.0535f
C315 Inverter_Layout_0.OUT.t5 Inverter_Layout_0.VSS 0.0754f
C316 Inverter_Layout_0.OUT.t42 Inverter_Layout_0.VSS 0.0518f
C317 Inverter_Layout_0.OUT.t6 Inverter_Layout_0.VSS 0.0535f
C318 Inverter_Layout_0.OUT.t38 Inverter_Layout_0.VSS 0.0754f
C319 Inverter_Layout_0.OUT.t30 Inverter_Layout_0.VSS 0.0518f
C320 Inverter_Layout_0.OUT.t39 Inverter_Layout_0.VSS 0.0535f
C321 Inverter_Layout_0.OUT.t28 Inverter_Layout_0.VSS 0.0754f
C322 Inverter_Layout_0.OUT.t16 Inverter_Layout_0.VSS 0.0518f
C323 Inverter_Layout_0.OUT.t37 Inverter_Layout_0.VSS 0.0535f
C324 Inverter_Layout_0.OUT.t25 Inverter_Layout_0.VSS 0.0754f
C325 Inverter_Layout_0.OUT.t14 Inverter_Layout_0.VSS 0.0518f
C326 Inverter_Layout_0.OUT.t26 Inverter_Layout_0.VSS 0.0535f
C327 Inverter_Layout_0.OUT.t11 Inverter_Layout_0.VSS 0.0754f
C328 Inverter_Layout_0.OUT.t0 Inverter_Layout_0.VSS 0.0518f
C329 Inverter_Layout_0.OUT.t23 Inverter_Layout_0.VSS 0.0535f
C330 Inverter_Layout_0.OUT.t8 Inverter_Layout_0.VSS 0.0754f
C331 Inverter_Layout_0.OUT.t46 Inverter_Layout_0.VSS 0.0518f
C332 Inverter_Layout_0.OUT.t27 Inverter_Layout_0.VSS 0.0535f
C333 Inverter_Layout_0.OUT.t12 Inverter_Layout_0.VSS 0.0754f
C334 Inverter_Layout_0.OUT.t1 Inverter_Layout_0.VSS 0.0518f
C335 Inverter_Layout_0.OUT.t13 Inverter_Layout_0.VSS 0.0535f
C336 Inverter_Layout_0.OUT.t47 Inverter_Layout_0.VSS 0.0754f
C337 Inverter_Layout_0.OUT.t33 Inverter_Layout_0.VSS 0.0518f
C338 Inverter_Layout_0.OUT.t9 Inverter_Layout_0.VSS 0.0535f
C339 Inverter_Layout_0.OUT.t45 Inverter_Layout_0.VSS 0.0754f
C340 Inverter_Layout_0.OUT.t32 Inverter_Layout_0.VSS 0.0518f
C341 Inverter_Layout_0.OUT.t43 Inverter_Layout_0.VSS 0.0535f
C342 Inverter_Layout_0.OUT.t31 Inverter_Layout_0.VSS 0.0754f
C343 Inverter_Layout_0.OUT.t17 Inverter_Layout_0.VSS 0.0703f
C344 Inverter_Layout_0.OUT.n0 Inverter_Layout_0.VSS 0.0622f
C345 Inverter_Layout_0.OUT.n1 Inverter_Layout_0.VSS 0.0454f
C346 Inverter_Layout_0.OUT.n2 Inverter_Layout_0.VSS 0.0454f
C347 Inverter_Layout_0.OUT.n3 Inverter_Layout_0.VSS 0.0454f
C348 Inverter_Layout_0.OUT.n4 Inverter_Layout_0.VSS 0.0454f
C349 Inverter_Layout_0.OUT.n5 Inverter_Layout_0.VSS 0.0454f
C350 Inverter_Layout_0.OUT.n6 Inverter_Layout_0.VSS 0.0454f
C351 Inverter_Layout_0.OUT.n7 Inverter_Layout_0.VSS 0.0454f
C352 Inverter_Layout_0.OUT.n8 Inverter_Layout_0.VSS 0.0454f
C353 Inverter_Layout_0.OUT.n9 Inverter_Layout_0.VSS 0.0454f
C354 Inverter_Layout_0.OUT.n10 Inverter_Layout_0.VSS 0.0454f
C355 Inverter_Layout_0.OUT.n11 Inverter_Layout_0.VSS 0.0454f
C356 Inverter_Layout_0.OUT.n12 Inverter_Layout_0.VSS 0.0454f
C357 Inverter_Layout_0.OUT.n13 Inverter_Layout_0.VSS 0.0622f
C358 Inverter_Layout_0.OUT.t41 Inverter_Layout_0.VSS 0.0703f
C359 Inverter_Layout_0.OUT.t4 Inverter_Layout_0.VSS 0.0754f
C360 Inverter_Layout_0.OUT.t19 Inverter_Layout_0.VSS 0.0783f
.ends

