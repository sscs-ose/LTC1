magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1133 -1741 1133 1741
<< metal2 >>
rect -133 736 133 741
rect -133 708 -128 736
rect -100 708 -52 736
rect -24 708 24 736
rect 52 708 100 736
rect 128 708 133 736
rect -133 660 133 708
rect -133 632 -128 660
rect -100 632 -52 660
rect -24 632 24 660
rect 52 632 100 660
rect 128 632 133 660
rect -133 584 133 632
rect -133 556 -128 584
rect -100 556 -52 584
rect -24 556 24 584
rect 52 556 100 584
rect 128 556 133 584
rect -133 508 133 556
rect -133 480 -128 508
rect -100 480 -52 508
rect -24 480 24 508
rect 52 480 100 508
rect 128 480 133 508
rect -133 432 133 480
rect -133 404 -128 432
rect -100 404 -52 432
rect -24 404 24 432
rect 52 404 100 432
rect 128 404 133 432
rect -133 356 133 404
rect -133 328 -128 356
rect -100 328 -52 356
rect -24 328 24 356
rect 52 328 100 356
rect 128 328 133 356
rect -133 280 133 328
rect -133 252 -128 280
rect -100 252 -52 280
rect -24 252 24 280
rect 52 252 100 280
rect 128 252 133 280
rect -133 204 133 252
rect -133 176 -128 204
rect -100 176 -52 204
rect -24 176 24 204
rect 52 176 100 204
rect 128 176 133 204
rect -133 128 133 176
rect -133 100 -128 128
rect -100 100 -52 128
rect -24 100 24 128
rect 52 100 100 128
rect 128 100 133 128
rect -133 52 133 100
rect -133 24 -128 52
rect -100 24 -52 52
rect -24 24 24 52
rect 52 24 100 52
rect 128 24 133 52
rect -133 -24 133 24
rect -133 -52 -128 -24
rect -100 -52 -52 -24
rect -24 -52 24 -24
rect 52 -52 100 -24
rect 128 -52 133 -24
rect -133 -100 133 -52
rect -133 -128 -128 -100
rect -100 -128 -52 -100
rect -24 -128 24 -100
rect 52 -128 100 -100
rect 128 -128 133 -100
rect -133 -176 133 -128
rect -133 -204 -128 -176
rect -100 -204 -52 -176
rect -24 -204 24 -176
rect 52 -204 100 -176
rect 128 -204 133 -176
rect -133 -252 133 -204
rect -133 -280 -128 -252
rect -100 -280 -52 -252
rect -24 -280 24 -252
rect 52 -280 100 -252
rect 128 -280 133 -252
rect -133 -328 133 -280
rect -133 -356 -128 -328
rect -100 -356 -52 -328
rect -24 -356 24 -328
rect 52 -356 100 -328
rect 128 -356 133 -328
rect -133 -404 133 -356
rect -133 -432 -128 -404
rect -100 -432 -52 -404
rect -24 -432 24 -404
rect 52 -432 100 -404
rect 128 -432 133 -404
rect -133 -480 133 -432
rect -133 -508 -128 -480
rect -100 -508 -52 -480
rect -24 -508 24 -480
rect 52 -508 100 -480
rect 128 -508 133 -480
rect -133 -556 133 -508
rect -133 -584 -128 -556
rect -100 -584 -52 -556
rect -24 -584 24 -556
rect 52 -584 100 -556
rect 128 -584 133 -556
rect -133 -632 133 -584
rect -133 -660 -128 -632
rect -100 -660 -52 -632
rect -24 -660 24 -632
rect 52 -660 100 -632
rect 128 -660 133 -632
rect -133 -708 133 -660
rect -133 -736 -128 -708
rect -100 -736 -52 -708
rect -24 -736 24 -708
rect 52 -736 100 -708
rect 128 -736 133 -708
rect -133 -741 133 -736
<< via2 >>
rect -128 708 -100 736
rect -52 708 -24 736
rect 24 708 52 736
rect 100 708 128 736
rect -128 632 -100 660
rect -52 632 -24 660
rect 24 632 52 660
rect 100 632 128 660
rect -128 556 -100 584
rect -52 556 -24 584
rect 24 556 52 584
rect 100 556 128 584
rect -128 480 -100 508
rect -52 480 -24 508
rect 24 480 52 508
rect 100 480 128 508
rect -128 404 -100 432
rect -52 404 -24 432
rect 24 404 52 432
rect 100 404 128 432
rect -128 328 -100 356
rect -52 328 -24 356
rect 24 328 52 356
rect 100 328 128 356
rect -128 252 -100 280
rect -52 252 -24 280
rect 24 252 52 280
rect 100 252 128 280
rect -128 176 -100 204
rect -52 176 -24 204
rect 24 176 52 204
rect 100 176 128 204
rect -128 100 -100 128
rect -52 100 -24 128
rect 24 100 52 128
rect 100 100 128 128
rect -128 24 -100 52
rect -52 24 -24 52
rect 24 24 52 52
rect 100 24 128 52
rect -128 -52 -100 -24
rect -52 -52 -24 -24
rect 24 -52 52 -24
rect 100 -52 128 -24
rect -128 -128 -100 -100
rect -52 -128 -24 -100
rect 24 -128 52 -100
rect 100 -128 128 -100
rect -128 -204 -100 -176
rect -52 -204 -24 -176
rect 24 -204 52 -176
rect 100 -204 128 -176
rect -128 -280 -100 -252
rect -52 -280 -24 -252
rect 24 -280 52 -252
rect 100 -280 128 -252
rect -128 -356 -100 -328
rect -52 -356 -24 -328
rect 24 -356 52 -328
rect 100 -356 128 -328
rect -128 -432 -100 -404
rect -52 -432 -24 -404
rect 24 -432 52 -404
rect 100 -432 128 -404
rect -128 -508 -100 -480
rect -52 -508 -24 -480
rect 24 -508 52 -480
rect 100 -508 128 -480
rect -128 -584 -100 -556
rect -52 -584 -24 -556
rect 24 -584 52 -556
rect 100 -584 128 -556
rect -128 -660 -100 -632
rect -52 -660 -24 -632
rect 24 -660 52 -632
rect 100 -660 128 -632
rect -128 -736 -100 -708
rect -52 -736 -24 -708
rect 24 -736 52 -708
rect 100 -736 128 -708
<< metal3 >>
rect -133 736 133 741
rect -133 708 -128 736
rect -100 708 -52 736
rect -24 708 24 736
rect 52 708 100 736
rect 128 708 133 736
rect -133 660 133 708
rect -133 632 -128 660
rect -100 632 -52 660
rect -24 632 24 660
rect 52 632 100 660
rect 128 632 133 660
rect -133 584 133 632
rect -133 556 -128 584
rect -100 556 -52 584
rect -24 556 24 584
rect 52 556 100 584
rect 128 556 133 584
rect -133 508 133 556
rect -133 480 -128 508
rect -100 480 -52 508
rect -24 480 24 508
rect 52 480 100 508
rect 128 480 133 508
rect -133 432 133 480
rect -133 404 -128 432
rect -100 404 -52 432
rect -24 404 24 432
rect 52 404 100 432
rect 128 404 133 432
rect -133 356 133 404
rect -133 328 -128 356
rect -100 328 -52 356
rect -24 328 24 356
rect 52 328 100 356
rect 128 328 133 356
rect -133 280 133 328
rect -133 252 -128 280
rect -100 252 -52 280
rect -24 252 24 280
rect 52 252 100 280
rect 128 252 133 280
rect -133 204 133 252
rect -133 176 -128 204
rect -100 176 -52 204
rect -24 176 24 204
rect 52 176 100 204
rect 128 176 133 204
rect -133 128 133 176
rect -133 100 -128 128
rect -100 100 -52 128
rect -24 100 24 128
rect 52 100 100 128
rect 128 100 133 128
rect -133 52 133 100
rect -133 24 -128 52
rect -100 24 -52 52
rect -24 24 24 52
rect 52 24 100 52
rect 128 24 133 52
rect -133 -24 133 24
rect -133 -52 -128 -24
rect -100 -52 -52 -24
rect -24 -52 24 -24
rect 52 -52 100 -24
rect 128 -52 133 -24
rect -133 -100 133 -52
rect -133 -128 -128 -100
rect -100 -128 -52 -100
rect -24 -128 24 -100
rect 52 -128 100 -100
rect 128 -128 133 -100
rect -133 -176 133 -128
rect -133 -204 -128 -176
rect -100 -204 -52 -176
rect -24 -204 24 -176
rect 52 -204 100 -176
rect 128 -204 133 -176
rect -133 -252 133 -204
rect -133 -280 -128 -252
rect -100 -280 -52 -252
rect -24 -280 24 -252
rect 52 -280 100 -252
rect 128 -280 133 -252
rect -133 -328 133 -280
rect -133 -356 -128 -328
rect -100 -356 -52 -328
rect -24 -356 24 -328
rect 52 -356 100 -328
rect 128 -356 133 -328
rect -133 -404 133 -356
rect -133 -432 -128 -404
rect -100 -432 -52 -404
rect -24 -432 24 -404
rect 52 -432 100 -404
rect 128 -432 133 -404
rect -133 -480 133 -432
rect -133 -508 -128 -480
rect -100 -508 -52 -480
rect -24 -508 24 -480
rect 52 -508 100 -480
rect 128 -508 133 -480
rect -133 -556 133 -508
rect -133 -584 -128 -556
rect -100 -584 -52 -556
rect -24 -584 24 -556
rect 52 -584 100 -556
rect 128 -584 133 -556
rect -133 -632 133 -584
rect -133 -660 -128 -632
rect -100 -660 -52 -632
rect -24 -660 24 -632
rect 52 -660 100 -632
rect 128 -660 133 -632
rect -133 -708 133 -660
rect -133 -736 -128 -708
rect -100 -736 -52 -708
rect -24 -736 24 -708
rect 52 -736 100 -708
rect 128 -736 133 -708
rect -133 -741 133 -736
<< end >>
