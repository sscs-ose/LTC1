magic
tech gf180mcuC
magscale 1 10
timestamp 1690971400
<< nwell >>
rect -602 -734 602 734
<< pmos >>
rect -428 404 -372 604
rect -268 404 -212 604
rect -108 404 -52 604
rect 52 404 108 604
rect 212 404 268 604
rect 372 404 428 604
rect -428 68 -372 268
rect -268 68 -212 268
rect -108 68 -52 268
rect 52 68 108 268
rect 212 68 268 268
rect 372 68 428 268
rect -428 -268 -372 -68
rect -268 -268 -212 -68
rect -108 -268 -52 -68
rect 52 -268 108 -68
rect 212 -268 268 -68
rect 372 -268 428 -68
rect -428 -604 -372 -404
rect -268 -604 -212 -404
rect -108 -604 -52 -404
rect 52 -604 108 -404
rect 212 -604 268 -404
rect 372 -604 428 -404
<< pdiff >>
rect -516 591 -428 604
rect -516 417 -503 591
rect -457 417 -428 591
rect -516 404 -428 417
rect -372 591 -268 604
rect -372 417 -343 591
rect -297 417 -268 591
rect -372 404 -268 417
rect -212 591 -108 604
rect -212 417 -183 591
rect -137 417 -108 591
rect -212 404 -108 417
rect -52 591 52 604
rect -52 417 -23 591
rect 23 417 52 591
rect -52 404 52 417
rect 108 591 212 604
rect 108 417 137 591
rect 183 417 212 591
rect 108 404 212 417
rect 268 591 372 604
rect 268 417 297 591
rect 343 417 372 591
rect 268 404 372 417
rect 428 591 516 604
rect 428 417 457 591
rect 503 417 516 591
rect 428 404 516 417
rect -516 255 -428 268
rect -516 81 -503 255
rect -457 81 -428 255
rect -516 68 -428 81
rect -372 255 -268 268
rect -372 81 -343 255
rect -297 81 -268 255
rect -372 68 -268 81
rect -212 255 -108 268
rect -212 81 -183 255
rect -137 81 -108 255
rect -212 68 -108 81
rect -52 255 52 268
rect -52 81 -23 255
rect 23 81 52 255
rect -52 68 52 81
rect 108 255 212 268
rect 108 81 137 255
rect 183 81 212 255
rect 108 68 212 81
rect 268 255 372 268
rect 268 81 297 255
rect 343 81 372 255
rect 268 68 372 81
rect 428 255 516 268
rect 428 81 457 255
rect 503 81 516 255
rect 428 68 516 81
rect -516 -81 -428 -68
rect -516 -255 -503 -81
rect -457 -255 -428 -81
rect -516 -268 -428 -255
rect -372 -81 -268 -68
rect -372 -255 -343 -81
rect -297 -255 -268 -81
rect -372 -268 -268 -255
rect -212 -81 -108 -68
rect -212 -255 -183 -81
rect -137 -255 -108 -81
rect -212 -268 -108 -255
rect -52 -81 52 -68
rect -52 -255 -23 -81
rect 23 -255 52 -81
rect -52 -268 52 -255
rect 108 -81 212 -68
rect 108 -255 137 -81
rect 183 -255 212 -81
rect 108 -268 212 -255
rect 268 -81 372 -68
rect 268 -255 297 -81
rect 343 -255 372 -81
rect 268 -268 372 -255
rect 428 -81 516 -68
rect 428 -255 457 -81
rect 503 -255 516 -81
rect 428 -268 516 -255
rect -516 -417 -428 -404
rect -516 -591 -503 -417
rect -457 -591 -428 -417
rect -516 -604 -428 -591
rect -372 -417 -268 -404
rect -372 -591 -343 -417
rect -297 -591 -268 -417
rect -372 -604 -268 -591
rect -212 -417 -108 -404
rect -212 -591 -183 -417
rect -137 -591 -108 -417
rect -212 -604 -108 -591
rect -52 -417 52 -404
rect -52 -591 -23 -417
rect 23 -591 52 -417
rect -52 -604 52 -591
rect 108 -417 212 -404
rect 108 -591 137 -417
rect 183 -591 212 -417
rect 108 -604 212 -591
rect 268 -417 372 -404
rect 268 -591 297 -417
rect 343 -591 372 -417
rect 268 -604 372 -591
rect 428 -417 516 -404
rect 428 -591 457 -417
rect 503 -591 516 -417
rect 428 -604 516 -591
<< pdiffc >>
rect -503 417 -457 591
rect -343 417 -297 591
rect -183 417 -137 591
rect -23 417 23 591
rect 137 417 183 591
rect 297 417 343 591
rect 457 417 503 591
rect -503 81 -457 255
rect -343 81 -297 255
rect -183 81 -137 255
rect -23 81 23 255
rect 137 81 183 255
rect 297 81 343 255
rect 457 81 503 255
rect -503 -255 -457 -81
rect -343 -255 -297 -81
rect -183 -255 -137 -81
rect -23 -255 23 -81
rect 137 -255 183 -81
rect 297 -255 343 -81
rect 457 -255 503 -81
rect -503 -591 -457 -417
rect -343 -591 -297 -417
rect -183 -591 -137 -417
rect -23 -591 23 -417
rect 137 -591 183 -417
rect 297 -591 343 -417
rect 457 -591 503 -417
<< polysilicon >>
rect -428 604 -372 648
rect -268 604 -212 648
rect -108 604 -52 648
rect 52 604 108 648
rect 212 604 268 648
rect 372 604 428 648
rect -428 360 -372 404
rect -268 360 -212 404
rect -108 360 -52 404
rect 52 360 108 404
rect 212 360 268 404
rect 372 360 428 404
rect -428 268 -372 312
rect -268 268 -212 312
rect -108 268 -52 312
rect 52 268 108 312
rect 212 268 268 312
rect 372 268 428 312
rect -428 24 -372 68
rect -268 24 -212 68
rect -108 24 -52 68
rect 52 24 108 68
rect 212 24 268 68
rect 372 24 428 68
rect -428 -68 -372 -24
rect -268 -68 -212 -24
rect -108 -68 -52 -24
rect 52 -68 108 -24
rect 212 -68 268 -24
rect 372 -68 428 -24
rect -428 -312 -372 -268
rect -268 -312 -212 -268
rect -108 -312 -52 -268
rect 52 -312 108 -268
rect 212 -312 268 -268
rect 372 -312 428 -268
rect -428 -404 -372 -360
rect -268 -404 -212 -360
rect -108 -404 -52 -360
rect 52 -404 108 -360
rect 212 -404 268 -360
rect 372 -404 428 -360
rect -428 -648 -372 -604
rect -268 -648 -212 -604
rect -108 -648 -52 -604
rect 52 -648 108 -604
rect 212 -648 268 -604
rect 372 -648 428 -604
<< metal1 >>
rect -503 591 -457 602
rect -503 406 -457 417
rect -343 591 -297 602
rect -343 406 -297 417
rect -183 591 -137 602
rect -183 406 -137 417
rect -23 591 23 602
rect -23 406 23 417
rect 137 591 183 602
rect 137 406 183 417
rect 297 591 343 602
rect 297 406 343 417
rect 457 591 503 602
rect 457 406 503 417
rect -503 255 -457 266
rect -503 70 -457 81
rect -343 255 -297 266
rect -343 70 -297 81
rect -183 255 -137 266
rect -183 70 -137 81
rect -23 255 23 266
rect -23 70 23 81
rect 137 255 183 266
rect 137 70 183 81
rect 297 255 343 266
rect 297 70 343 81
rect 457 255 503 266
rect 457 70 503 81
rect -503 -81 -457 -70
rect -503 -266 -457 -255
rect -343 -81 -297 -70
rect -343 -266 -297 -255
rect -183 -81 -137 -70
rect -183 -266 -137 -255
rect -23 -81 23 -70
rect -23 -266 23 -255
rect 137 -81 183 -70
rect 137 -266 183 -255
rect 297 -81 343 -70
rect 297 -266 343 -255
rect 457 -81 503 -70
rect 457 -266 503 -255
rect -503 -417 -457 -406
rect -503 -602 -457 -591
rect -343 -417 -297 -406
rect -343 -602 -297 -591
rect -183 -417 -137 -406
rect -183 -602 -137 -591
rect -23 -417 23 -406
rect -23 -602 23 -591
rect 137 -417 183 -406
rect 137 -602 183 -591
rect 297 -417 343 -406
rect 297 -602 343 -591
rect 457 -417 503 -406
rect 457 -602 503 -591
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 1 l 0.280 m 4 nf 6 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
