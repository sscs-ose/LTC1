** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/MSB_CELL_TB.sch
**.subckt MSB_CELL_TB
V1 VSS GND 0
.save i(v1)
V2 VDD VSS 3.3
.save i(v2)
I0 VDD IM_T 80u
XM1 IM_T IM_T IM VSS nfet_03v3 L=0.5u W=19.2u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 IM IM VSS VSS nfet_03v3 L=0.5u W=19.2u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
V4 Ri-1 VSS pulse(0 3.3 0 10p 10p 3200n 6400n )
.save i(v4)
V3 Ri VSS pulse(0 3.3 100n 10p 10p 6400n 12800n)
.save i(v3)
V5 Ci VSS pulse(0 3.3 200 10p 10p 12800n 25600n)
.save i(v5)
R1 IOUT- VDD 10k m=1
R2 IOUT+ VDD 10k m=1
x1 IOUT+ IOUT- VDD Ri-1 Ri Ci IM_T IM VSS pex_MSB_Unit_Cell
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.include pex_MSB_Unit_Cell.spice
.options savecurrents

.control
save all
tran 10n 20.6u

plot v(IOUT+) v(IOUT-)
*write test_nfet_03v3.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
