magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1286 -1319 1286 1319
<< metal4 >>
rect -283 311 283 316
rect -283 283 -278 311
rect -250 283 -212 311
rect -184 283 -146 311
rect -118 283 -80 311
rect -52 283 -14 311
rect 14 283 52 311
rect 80 283 118 311
rect 146 283 184 311
rect 212 283 250 311
rect 278 283 283 311
rect -283 245 283 283
rect -283 217 -278 245
rect -250 217 -212 245
rect -184 217 -146 245
rect -118 217 -80 245
rect -52 217 -14 245
rect 14 217 52 245
rect 80 217 118 245
rect 146 217 184 245
rect 212 217 250 245
rect 278 217 283 245
rect -283 179 283 217
rect -283 151 -278 179
rect -250 151 -212 179
rect -184 151 -146 179
rect -118 151 -80 179
rect -52 151 -14 179
rect 14 151 52 179
rect 80 151 118 179
rect 146 151 184 179
rect 212 151 250 179
rect 278 151 283 179
rect -283 113 283 151
rect -283 85 -278 113
rect -250 85 -212 113
rect -184 85 -146 113
rect -118 85 -80 113
rect -52 85 -14 113
rect 14 85 52 113
rect 80 85 118 113
rect 146 85 184 113
rect 212 85 250 113
rect 278 85 283 113
rect -283 47 283 85
rect -283 19 -278 47
rect -250 19 -212 47
rect -184 19 -146 47
rect -118 19 -80 47
rect -52 19 -14 47
rect 14 19 52 47
rect 80 19 118 47
rect 146 19 184 47
rect 212 19 250 47
rect 278 19 283 47
rect -283 -19 283 19
rect -283 -47 -278 -19
rect -250 -47 -212 -19
rect -184 -47 -146 -19
rect -118 -47 -80 -19
rect -52 -47 -14 -19
rect 14 -47 52 -19
rect 80 -47 118 -19
rect 146 -47 184 -19
rect 212 -47 250 -19
rect 278 -47 283 -19
rect -283 -85 283 -47
rect -283 -113 -278 -85
rect -250 -113 -212 -85
rect -184 -113 -146 -85
rect -118 -113 -80 -85
rect -52 -113 -14 -85
rect 14 -113 52 -85
rect 80 -113 118 -85
rect 146 -113 184 -85
rect 212 -113 250 -85
rect 278 -113 283 -85
rect -283 -151 283 -113
rect -283 -179 -278 -151
rect -250 -179 -212 -151
rect -184 -179 -146 -151
rect -118 -179 -80 -151
rect -52 -179 -14 -151
rect 14 -179 52 -151
rect 80 -179 118 -151
rect 146 -179 184 -151
rect 212 -179 250 -151
rect 278 -179 283 -151
rect -283 -217 283 -179
rect -283 -245 -278 -217
rect -250 -245 -212 -217
rect -184 -245 -146 -217
rect -118 -245 -80 -217
rect -52 -245 -14 -217
rect 14 -245 52 -217
rect 80 -245 118 -217
rect 146 -245 184 -217
rect 212 -245 250 -217
rect 278 -245 283 -217
rect -283 -283 283 -245
rect -283 -311 -278 -283
rect -250 -311 -212 -283
rect -184 -311 -146 -283
rect -118 -311 -80 -283
rect -52 -311 -14 -283
rect 14 -311 52 -283
rect 80 -311 118 -283
rect 146 -311 184 -283
rect 212 -311 250 -283
rect 278 -311 283 -283
rect -283 -316 283 -311
<< via4 >>
rect -278 283 -250 311
rect -212 283 -184 311
rect -146 283 -118 311
rect -80 283 -52 311
rect -14 283 14 311
rect 52 283 80 311
rect 118 283 146 311
rect 184 283 212 311
rect 250 283 278 311
rect -278 217 -250 245
rect -212 217 -184 245
rect -146 217 -118 245
rect -80 217 -52 245
rect -14 217 14 245
rect 52 217 80 245
rect 118 217 146 245
rect 184 217 212 245
rect 250 217 278 245
rect -278 151 -250 179
rect -212 151 -184 179
rect -146 151 -118 179
rect -80 151 -52 179
rect -14 151 14 179
rect 52 151 80 179
rect 118 151 146 179
rect 184 151 212 179
rect 250 151 278 179
rect -278 85 -250 113
rect -212 85 -184 113
rect -146 85 -118 113
rect -80 85 -52 113
rect -14 85 14 113
rect 52 85 80 113
rect 118 85 146 113
rect 184 85 212 113
rect 250 85 278 113
rect -278 19 -250 47
rect -212 19 -184 47
rect -146 19 -118 47
rect -80 19 -52 47
rect -14 19 14 47
rect 52 19 80 47
rect 118 19 146 47
rect 184 19 212 47
rect 250 19 278 47
rect -278 -47 -250 -19
rect -212 -47 -184 -19
rect -146 -47 -118 -19
rect -80 -47 -52 -19
rect -14 -47 14 -19
rect 52 -47 80 -19
rect 118 -47 146 -19
rect 184 -47 212 -19
rect 250 -47 278 -19
rect -278 -113 -250 -85
rect -212 -113 -184 -85
rect -146 -113 -118 -85
rect -80 -113 -52 -85
rect -14 -113 14 -85
rect 52 -113 80 -85
rect 118 -113 146 -85
rect 184 -113 212 -85
rect 250 -113 278 -85
rect -278 -179 -250 -151
rect -212 -179 -184 -151
rect -146 -179 -118 -151
rect -80 -179 -52 -151
rect -14 -179 14 -151
rect 52 -179 80 -151
rect 118 -179 146 -151
rect 184 -179 212 -151
rect 250 -179 278 -151
rect -278 -245 -250 -217
rect -212 -245 -184 -217
rect -146 -245 -118 -217
rect -80 -245 -52 -217
rect -14 -245 14 -217
rect 52 -245 80 -217
rect 118 -245 146 -217
rect 184 -245 212 -217
rect 250 -245 278 -217
rect -278 -311 -250 -283
rect -212 -311 -184 -283
rect -146 -311 -118 -283
rect -80 -311 -52 -283
rect -14 -311 14 -283
rect 52 -311 80 -283
rect 118 -311 146 -283
rect 184 -311 212 -283
rect 250 -311 278 -283
<< metal5 >>
rect -286 311 286 319
rect -286 283 -278 311
rect -250 283 -212 311
rect -184 283 -146 311
rect -118 283 -80 311
rect -52 283 -14 311
rect 14 283 52 311
rect 80 283 118 311
rect 146 283 184 311
rect 212 283 250 311
rect 278 283 286 311
rect -286 245 286 283
rect -286 217 -278 245
rect -250 217 -212 245
rect -184 217 -146 245
rect -118 217 -80 245
rect -52 217 -14 245
rect 14 217 52 245
rect 80 217 118 245
rect 146 217 184 245
rect 212 217 250 245
rect 278 217 286 245
rect -286 179 286 217
rect -286 151 -278 179
rect -250 151 -212 179
rect -184 151 -146 179
rect -118 151 -80 179
rect -52 151 -14 179
rect 14 151 52 179
rect 80 151 118 179
rect 146 151 184 179
rect 212 151 250 179
rect 278 151 286 179
rect -286 113 286 151
rect -286 85 -278 113
rect -250 85 -212 113
rect -184 85 -146 113
rect -118 85 -80 113
rect -52 85 -14 113
rect 14 85 52 113
rect 80 85 118 113
rect 146 85 184 113
rect 212 85 250 113
rect 278 85 286 113
rect -286 47 286 85
rect -286 19 -278 47
rect -250 19 -212 47
rect -184 19 -146 47
rect -118 19 -80 47
rect -52 19 -14 47
rect 14 19 52 47
rect 80 19 118 47
rect 146 19 184 47
rect 212 19 250 47
rect 278 19 286 47
rect -286 -19 286 19
rect -286 -47 -278 -19
rect -250 -47 -212 -19
rect -184 -47 -146 -19
rect -118 -47 -80 -19
rect -52 -47 -14 -19
rect 14 -47 52 -19
rect 80 -47 118 -19
rect 146 -47 184 -19
rect 212 -47 250 -19
rect 278 -47 286 -19
rect -286 -85 286 -47
rect -286 -113 -278 -85
rect -250 -113 -212 -85
rect -184 -113 -146 -85
rect -118 -113 -80 -85
rect -52 -113 -14 -85
rect 14 -113 52 -85
rect 80 -113 118 -85
rect 146 -113 184 -85
rect 212 -113 250 -85
rect 278 -113 286 -85
rect -286 -151 286 -113
rect -286 -179 -278 -151
rect -250 -179 -212 -151
rect -184 -179 -146 -151
rect -118 -179 -80 -151
rect -52 -179 -14 -151
rect 14 -179 52 -151
rect 80 -179 118 -151
rect 146 -179 184 -151
rect 212 -179 250 -151
rect 278 -179 286 -151
rect -286 -217 286 -179
rect -286 -245 -278 -217
rect -250 -245 -212 -217
rect -184 -245 -146 -217
rect -118 -245 -80 -217
rect -52 -245 -14 -217
rect 14 -245 52 -217
rect 80 -245 118 -217
rect 146 -245 184 -217
rect 212 -245 250 -217
rect 278 -245 286 -217
rect -286 -283 286 -245
rect -286 -311 -278 -283
rect -250 -311 -212 -283
rect -184 -311 -146 -283
rect -118 -311 -80 -283
rect -52 -311 -14 -283
rect 14 -311 52 -283
rect 80 -311 118 -283
rect 146 -311 184 -283
rect 212 -311 250 -283
rect 278 -311 286 -283
rect -286 -319 286 -311
<< end >>
