magic
tech gf180mcuC
magscale 1 10
timestamp 1699963945
<< nwell >>
rect -1186 -1166 1186 1166
<< pmos >>
rect -1012 436 -812 1036
rect -708 436 -508 1036
rect -404 436 -204 1036
rect -100 436 100 1036
rect 204 436 404 1036
rect 508 436 708 1036
rect 812 436 1012 1036
rect -1012 -300 -812 300
rect -708 -300 -508 300
rect -404 -300 -204 300
rect -100 -300 100 300
rect 204 -300 404 300
rect 508 -300 708 300
rect 812 -300 1012 300
rect -1012 -1036 -812 -436
rect -708 -1036 -508 -436
rect -404 -1036 -204 -436
rect -100 -1036 100 -436
rect 204 -1036 404 -436
rect 508 -1036 708 -436
rect 812 -1036 1012 -436
<< pdiff >>
rect -1100 1023 -1012 1036
rect -1100 449 -1087 1023
rect -1041 449 -1012 1023
rect -1100 436 -1012 449
rect -812 1023 -708 1036
rect -812 449 -783 1023
rect -737 449 -708 1023
rect -812 436 -708 449
rect -508 1023 -404 1036
rect -508 449 -479 1023
rect -433 449 -404 1023
rect -508 436 -404 449
rect -204 1023 -100 1036
rect -204 449 -175 1023
rect -129 449 -100 1023
rect -204 436 -100 449
rect 100 1023 204 1036
rect 100 449 129 1023
rect 175 449 204 1023
rect 100 436 204 449
rect 404 1023 508 1036
rect 404 449 433 1023
rect 479 449 508 1023
rect 404 436 508 449
rect 708 1023 812 1036
rect 708 449 737 1023
rect 783 449 812 1023
rect 708 436 812 449
rect 1012 1023 1100 1036
rect 1012 449 1041 1023
rect 1087 449 1100 1023
rect 1012 436 1100 449
rect -1100 287 -1012 300
rect -1100 -287 -1087 287
rect -1041 -287 -1012 287
rect -1100 -300 -1012 -287
rect -812 287 -708 300
rect -812 -287 -783 287
rect -737 -287 -708 287
rect -812 -300 -708 -287
rect -508 287 -404 300
rect -508 -287 -479 287
rect -433 -287 -404 287
rect -508 -300 -404 -287
rect -204 287 -100 300
rect -204 -287 -175 287
rect -129 -287 -100 287
rect -204 -300 -100 -287
rect 100 287 204 300
rect 100 -287 129 287
rect 175 -287 204 287
rect 100 -300 204 -287
rect 404 287 508 300
rect 404 -287 433 287
rect 479 -287 508 287
rect 404 -300 508 -287
rect 708 287 812 300
rect 708 -287 737 287
rect 783 -287 812 287
rect 708 -300 812 -287
rect 1012 287 1100 300
rect 1012 -287 1041 287
rect 1087 -287 1100 287
rect 1012 -300 1100 -287
rect -1100 -449 -1012 -436
rect -1100 -1023 -1087 -449
rect -1041 -1023 -1012 -449
rect -1100 -1036 -1012 -1023
rect -812 -449 -708 -436
rect -812 -1023 -783 -449
rect -737 -1023 -708 -449
rect -812 -1036 -708 -1023
rect -508 -449 -404 -436
rect -508 -1023 -479 -449
rect -433 -1023 -404 -449
rect -508 -1036 -404 -1023
rect -204 -449 -100 -436
rect -204 -1023 -175 -449
rect -129 -1023 -100 -449
rect -204 -1036 -100 -1023
rect 100 -449 204 -436
rect 100 -1023 129 -449
rect 175 -1023 204 -449
rect 100 -1036 204 -1023
rect 404 -449 508 -436
rect 404 -1023 433 -449
rect 479 -1023 508 -449
rect 404 -1036 508 -1023
rect 708 -449 812 -436
rect 708 -1023 737 -449
rect 783 -1023 812 -449
rect 708 -1036 812 -1023
rect 1012 -449 1100 -436
rect 1012 -1023 1041 -449
rect 1087 -1023 1100 -449
rect 1012 -1036 1100 -1023
<< pdiffc >>
rect -1087 449 -1041 1023
rect -783 449 -737 1023
rect -479 449 -433 1023
rect -175 449 -129 1023
rect 129 449 175 1023
rect 433 449 479 1023
rect 737 449 783 1023
rect 1041 449 1087 1023
rect -1087 -287 -1041 287
rect -783 -287 -737 287
rect -479 -287 -433 287
rect -175 -287 -129 287
rect 129 -287 175 287
rect 433 -287 479 287
rect 737 -287 783 287
rect 1041 -287 1087 287
rect -1087 -1023 -1041 -449
rect -783 -1023 -737 -449
rect -479 -1023 -433 -449
rect -175 -1023 -129 -449
rect 129 -1023 175 -449
rect 433 -1023 479 -449
rect 737 -1023 783 -449
rect 1041 -1023 1087 -449
<< polysilicon >>
rect -1012 1036 -812 1080
rect -708 1036 -508 1080
rect -404 1036 -204 1080
rect -100 1036 100 1080
rect 204 1036 404 1080
rect 508 1036 708 1080
rect 812 1036 1012 1080
rect -1012 392 -812 436
rect -708 392 -508 436
rect -404 392 -204 436
rect -100 392 100 436
rect 204 392 404 436
rect 508 392 708 436
rect 812 392 1012 436
rect -1012 300 -812 344
rect -708 300 -508 344
rect -404 300 -204 344
rect -100 300 100 344
rect 204 300 404 344
rect 508 300 708 344
rect 812 300 1012 344
rect -1012 -344 -812 -300
rect -708 -344 -508 -300
rect -404 -344 -204 -300
rect -100 -344 100 -300
rect 204 -344 404 -300
rect 508 -344 708 -300
rect 812 -344 1012 -300
rect -1012 -436 -812 -392
rect -708 -436 -508 -392
rect -404 -436 -204 -392
rect -100 -436 100 -392
rect 204 -436 404 -392
rect 508 -436 708 -392
rect 812 -436 1012 -392
rect -1012 -1080 -812 -1036
rect -708 -1080 -508 -1036
rect -404 -1080 -204 -1036
rect -100 -1080 100 -1036
rect 204 -1080 404 -1036
rect 508 -1080 708 -1036
rect 812 -1080 1012 -1036
<< metal1 >>
rect -1087 1023 -1041 1034
rect -1087 438 -1041 449
rect -783 1023 -737 1034
rect -783 438 -737 449
rect -479 1023 -433 1034
rect -479 438 -433 449
rect -175 1023 -129 1034
rect -175 438 -129 449
rect 129 1023 175 1034
rect 129 438 175 449
rect 433 1023 479 1034
rect 433 438 479 449
rect 737 1023 783 1034
rect 737 438 783 449
rect 1041 1023 1087 1034
rect 1041 438 1087 449
rect -1087 287 -1041 298
rect -1087 -298 -1041 -287
rect -783 287 -737 298
rect -783 -298 -737 -287
rect -479 287 -433 298
rect -479 -298 -433 -287
rect -175 287 -129 298
rect -175 -298 -129 -287
rect 129 287 175 298
rect 129 -298 175 -287
rect 433 287 479 298
rect 433 -298 479 -287
rect 737 287 783 298
rect 737 -298 783 -287
rect 1041 287 1087 298
rect 1041 -298 1087 -287
rect -1087 -449 -1041 -438
rect -1087 -1034 -1041 -1023
rect -783 -449 -737 -438
rect -783 -1034 -737 -1023
rect -479 -449 -433 -438
rect -479 -1034 -433 -1023
rect -175 -449 -129 -438
rect -175 -1034 -129 -1023
rect 129 -449 175 -438
rect 129 -1034 175 -1023
rect 433 -449 479 -438
rect 433 -1034 479 -1023
rect 737 -449 783 -438
rect 737 -1034 783 -1023
rect 1041 -449 1087 -438
rect 1041 -1034 1087 -1023
<< properties >>
string gencell pfet_03v3
string library gf180mcu
string parameters w 3 l 1 m 3 nf 7 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>
