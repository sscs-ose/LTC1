magic
tech gf180mcuC
magscale 1 10
timestamp 1692016503
<< nwell >>
rect -58 405 738 873
<< pwell >>
rect -4 0 676 194
<< nmos >>
rect 112 75 560 119
<< pmos >>
rect 116 535 564 623
<< ndiff >>
rect 20 120 92 133
rect 20 74 33 120
rect 79 119 92 120
rect 580 120 652 133
rect 580 119 593 120
rect 79 75 112 119
rect 560 75 593 119
rect 79 74 92 75
rect 20 61 92 74
rect 580 74 593 75
rect 639 74 652 120
rect 580 61 652 74
<< pdiff >>
rect 28 610 116 623
rect 28 548 41 610
rect 87 548 116 610
rect 28 535 116 548
rect 564 610 652 623
rect 564 548 593 610
rect 639 548 652 610
rect 564 535 652 548
<< ndiffc >>
rect 33 74 79 120
rect 593 74 639 120
<< pdiffc >>
rect 41 548 87 610
rect 593 548 639 610
<< psubdiff >>
rect 16 -28 656 -15
rect 16 -74 29 -28
rect 75 -74 123 -28
rect 169 -74 217 -28
rect 263 -74 311 -28
rect 357 -74 405 -28
rect 451 -74 499 -28
rect 545 -74 593 -28
rect 639 -74 656 -28
rect 16 -87 656 -74
<< nsubdiff >>
rect -21 827 709 840
rect -21 781 -8 827
rect 38 781 86 827
rect 132 781 180 827
rect 226 781 274 827
rect 320 781 368 827
rect 414 781 462 827
rect 508 781 556 827
rect 602 781 650 827
rect 696 781 709 827
rect -21 768 709 781
<< psubdiffcont >>
rect 29 -74 75 -28
rect 123 -74 169 -28
rect 217 -74 263 -28
rect 311 -74 357 -28
rect 405 -74 451 -28
rect 499 -74 545 -28
rect 593 -74 639 -28
<< nsubdiffcont >>
rect -8 781 38 827
rect 86 781 132 827
rect 180 781 226 827
rect 274 781 320 827
rect 368 781 414 827
rect 462 781 508 827
rect 556 781 602 827
rect 650 781 696 827
<< polysilicon >>
rect 116 623 564 667
rect 116 491 564 535
rect 183 373 255 381
rect 303 373 415 491
rect 183 368 415 373
rect 183 322 196 368
rect 242 322 415 368
rect 183 317 415 322
rect 183 309 255 317
rect 303 163 415 317
rect 112 119 560 163
rect 112 31 560 75
<< polycontact >>
rect 196 322 242 368
<< metal1 >>
rect -58 827 738 860
rect -58 781 -8 827
rect 38 781 86 827
rect 132 781 180 827
rect 226 781 274 827
rect 320 781 368 827
rect 414 781 462 827
rect 508 781 556 827
rect 602 781 650 827
rect 696 781 738 827
rect -58 748 738 781
rect 41 610 87 748
rect 41 537 87 548
rect 593 610 639 621
rect 183 368 253 379
rect 117 322 196 368
rect 242 322 253 368
rect 183 315 253 322
rect 185 311 253 315
rect 593 368 639 548
rect 593 322 729 368
rect 593 120 639 322
rect 22 74 33 120
rect 79 74 90 120
rect 582 74 593 120
rect 639 74 650 120
rect 33 5 79 74
rect -4 -28 676 5
rect -4 -74 29 -28
rect 75 -74 123 -28
rect 169 -74 217 -28
rect 263 -74 311 -28
rect 357 -74 405 -28
rect 451 -74 499 -28
rect 545 -74 593 -28
rect 639 -74 676 -28
rect -4 -107 676 -74
<< labels >>
flabel psubdiffcont 334 -51 334 -51 0 FreeSans 320 0 0 0 VSS
port 4 nsew
flabel nsubdiffcont 297 804 297 804 0 FreeSans 320 0 0 0 VDD
port 5 nsew
flabel metal1 143 345 143 345 0 FreeSans 320 0 0 0 IN
port 2 nsew
flabel metal1 651 345 651 345 0 FreeSans 320 0 0 0 OUT
port 3 nsew
<< end >>
