* NGSPICE file created from OR_magic_flat.ext - technology: gf180mcuC

.subckt OR_magic_flat A B OUT VDD VSS
X0 OUT a_86_n570# VDD.t7 VDD.t4 pfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X1 a_86_n570# B.t0 a_234_n257# VDD.t2 pfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X2 a_234_n257# A.t0 VDD.t1 VDD.t0 pfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X3 VDD.t5 VDD.t3 VDD.t5 VDD.t4 pfet_03v3 ad=0.155p pd=1.64u as=0 ps=0 w=0.25u l=0.28u
X4 a_86_n570# B.t1 a_234_n257# VDD.t2 pfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X5 a_234_n257# A.t1 VDD.t10 VDD.t0 pfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X6 a_234_n257# A.t2 VDD.t8 VDD.t0 pfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X7 a_86_n570# B.t2 a_234_n257# VDD.t2 pfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X8 OUT a_86_n570# VSS.t1 VSS.t0 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X9 a_86_n570# B.t3 a_234_n257# VDD.t2 pfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X10 a_86_n570# B.t4 VSS.t3 VSS.t2 nfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X11 OUT a_86_n570# VDD.t6 VDD.t4 pfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X12 VSS A.t3 a_86_n570# VSS.t4 nfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X13 a_234_n257# A.t4 VDD.t9 VDD.t0 pfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
R0 VDD.n13 VDD.t2 64.9948
R1 VDD.n2 VDD.t3 17.4273
R2 VDD.n10 VDD.t0 16.5878
R3 VDD.n3 VDD.t4 14.4507
R4 VDD.n6 VDD.t1 9.12573
R5 VDD.n0 VDD.t6 9.12573
R6 VDD.n8 VDD.t9 8.9005
R7 VDD.n7 VDD.t8 8.9005
R8 VDD.n6 VDD.t10 8.9005
R9 VDD.n0 VDD.t7 8.9005
R10 VDD.n18 VDD.n17 8.86445
R11 VDD.n1 VDD.t5 4.451
R12 VDD.n17 VDD.n5 3.1505
R13 VDD.n17 VDD.n16 3.1505
R14 VDD.n21 VDD.n20 3.1505
R15 VDD.n20 VDD.n19 3.1505
R16 VDD.n15 VDD.n14 3.1505
R17 VDD.n14 VDD.n13 3.1505
R18 VDD.n12 VDD.n11 3.1505
R19 VDD.n4 VDD.n3 2.45371
R20 VDD.n1 VDD.n0 0.60793
R21 VDD.n9 VDD.n8 0.367463
R22 VDD.n7 VDD.n6 0.2316
R23 VDD.n8 VDD.n7 0.22573
R24 VDD.n11 VDD.n10 0.183455
R25 VDD.n20 VDD.n18 0.147012
R26 VDD.n2 VDD.n1 0.125892
R27 VDD.n21 VDD.n15 0.0976053
R28 VDD.n15 VDD.n12 0.0976053
R29 VDD VDD.n5 0.0960263
R30 VDD.n4 VDD.n2 0.0924565
R31 VDD.n5 VDD.n4 0.0897105
R32 VDD.n12 VDD.n9 0.0573421
R33 VDD VDD.n21 0.00207895
R34 OUT.n3 OUT.n2 9.38225
R35 OUT.n4 OUT.n0 8.9005
R36 OUT.n3 OUT.n1 8.9005
R37 OUT OUT.n4 0.293115
R38 OUT.n4 OUT.n3 0.22573
R39 B.n0 B.t4 23.8759
R40 B.t1 B.t2 17.338
R41 B.t2 B.t3 16.9469
R42 B.t0 B.t1 16.9469
R43 B.n0 B.t0 11.8831
R44 B B.n0 4.77137
R45 A.t0 A.t3 39.3684
R46 A A.t4 36.6468
R47 A.t2 A.t1 17.338
R48 A.t1 A.t0 16.9469
R49 A.t4 A.t2 16.9469
R50 VSS.n7 VSS.t2 494
R51 VSS.n5 VSS.t4 106.591
R52 VSS.n0 VSS.t0 89.2573
R53 VSS.n12 VSS.n11 9.84934
R54 VSS.n1 VSS.t1 9.04072
R55 VSS.n4 VSS.n3 5.6705
R56 VSS.n4 VSS.t3 5.6705
R57 VSS.n6 VSS.n4 3.37072
R58 VSS.n11 VSS.n2 2.6005
R59 VSS.n11 VSS.n10 2.6005
R60 VSS.n15 VSS.n14 2.6005
R61 VSS.n14 VSS.n13 2.6005
R62 VSS.n9 VSS.n8 2.6005
R63 VSS.n8 VSS.n7 2.6005
R64 VSS.n6 VSS.n5 2.2294
R65 VSS.n1 VSS.n0 2.22783
R66 VSS.n14 VSS.n12 0.163291
R67 VSS.n15 VSS.n9 0.0976053
R68 VSS VSS.n2 0.0960263
R69 VSS.n2 VSS.n1 0.0233947
R70 VSS.n9 VSS.n6 0.0218158
R71 VSS VSS.n15 0.00207895
C0 OUT VDD 0.21f
C1 A B 0.0969f
C2 A a_234_n257# 0.0203f
C3 A a_86_n570# 0.0201f
C4 OUT B 2.43e-19
C5 OUT a_86_n570# 0.115f
C6 VDD B 0.357f
C7 VDD a_234_n257# 0.219f
C8 VDD a_86_n570# 0.606f
C9 B a_234_n257# 0.0835f
C10 B a_86_n570# 0.399f
C11 a_86_n570# a_234_n257# 0.18f
C12 A VDD 0.472f
.ends

