** sch_path: /home/shahid/GF180Projects/PFD/xschem/analog_mux_test.sch
**.subckt analog_mux_test
x1 S VSS VDD OUT I1 I0 analog_mux
V1 VDD VSS 3.3
.save i(v1)
V2 VSS GND 0
.save i(v2)
V4 S VSS pulse(3.3 0 0 100p 100p 400n 800n)
.save i(v4)
V6 I1 VSS PWL(0 2 400n 3 600n 2.5 700n 3.3)
.save i(v6)
V7 I0 VSS PWL(0 0 50n 1 100n 2 200n 3.3)
.save i(v7)
**** begin user architecture code


.control
save all
tran 50p 800n
plot v(S)  v(I0)+5 v(I1)+10 v(OUT)+15


*write test_nfet_03v3.raw
.endc



.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical

**** end user architecture code
**.ends

* expanding   symbol:  analog_mux.sym # of pins=6
** sym_path: /home/shahid/GF180Projects/PFD/xschem/analog_mux.sym
** sch_path: /home/shahid/GF180Projects/PFD/xschem/analog_mux.sch
.subckt analog_mux S VSS VDD OUT I1 I0
*.ipin I0
*.ipin I1
*.ipin S
*.iopin VSS
*.iopin VDD
*.opin OUT
x1 VDD SB VSS OUT I0 tg
x2 VDD S VSS OUT I1 tg
x3 VSS S SB VSS inv_my
.ends


* expanding   symbol:  tg.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/PFD/xschem/tg.sym
** sch_path: /home/shahid/GF180Projects/PFD/xschem/tg.sch
.subckt tg OUT S VSS VDD IN
*.iopin IN
*.iopin OUT
*.ipin S
*.iopin VSS
*.iopin VDD
x1 VSS S net1 VDD inv_my
XM1 IN net1 OUT VDD pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 IN S OUT VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  inv_my.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/PFD/xschem/inv_my.sym
** sch_path: /home/shahid/GF180Projects/PFD/xschem/inv_my.sch
.subckt inv_my VSS IN OUT VDD
*.iopin VDD
*.iopin VSS
*.ipin IN
*.opin OUT
XM1 OUT IN VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT IN VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends

.GLOBAL GND
.end
