magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2767 -3312 15147 17294
<< nwell >>
rect -2 111 12382 13618
<< psubdiff >>
rect -767 13666 13147 15294
rect -767 13534 -53 13666
rect 12433 13534 13147 13666
rect -121 63 -53 163
rect 12433 63 12501 163
rect -121 -805 12501 63
rect -767 -910 13147 -805
rect -767 -1312 -53 -910
rect 12433 -1312 13147 -910
<< nsubdiff >>
rect 81 13500 12299 13540
rect 81 12958 1318 13500
rect 81 11596 624 12958
rect 858 11596 1318 12958
rect 81 11554 1318 11596
rect 2264 11554 3018 13500
rect 4064 11554 4818 13500
rect 5764 11554 6618 13500
rect 7564 11554 8318 13500
rect 9364 11554 10118 13500
rect 11064 12958 12299 13500
rect 11064 11596 11524 12958
rect 11758 11596 12299 12958
rect 11064 11554 12299 11596
rect 81 11504 12299 11554
rect 81 2431 451 11504
rect 11931 2431 12299 11504
rect 81 246 12299 2431
<< nsubdiffcont >>
rect 624 11596 858 12958
rect 1318 11554 2264 13500
rect 3018 11554 4064 13500
rect 4818 11554 5764 13500
rect 6618 11554 7564 13500
rect 8318 11554 9364 13500
rect 10118 11554 11064 13500
rect 11524 11596 11758 12958
<< polysilicon >>
rect 974 11060 1185 11144
rect 2360 11060 2571 11144
rect 2746 11060 2957 11144
rect 4120 11060 4331 11144
rect 4511 11060 4722 11144
rect 5892 11060 6103 11144
rect 6280 11060 6491 11144
rect 7662 11060 7873 11144
rect 8049 11060 8260 11144
rect 9428 11060 9639 11144
rect 9815 11060 10026 11144
rect 11201 11060 11412 11144
rect 974 2800 1185 2884
rect 2360 2800 2571 2884
rect 2746 2800 2957 2884
rect 4120 2800 4331 2884
rect 4511 2800 4722 2884
rect 5892 2800 6103 2884
rect 6280 2800 6491 2884
rect 7662 2800 7873 2884
rect 8049 2800 8260 2884
rect 9428 2800 9639 2884
rect 9815 2800 10026 2884
rect 11201 2800 11412 2884
<< metal1 >>
rect -756 52 -64 14582
rect 1267 13500 2286 13540
rect 376 13122 889 13490
rect 92 13029 889 13122
rect 376 12958 889 13029
rect 376 11596 624 12958
rect 858 11596 889 12958
rect 376 11543 889 11596
rect 1267 11554 1318 13500
rect 2264 11554 2286 13500
rect 1267 11543 2286 11554
rect 2983 13500 4093 13540
rect 2983 11554 3018 13500
rect 4064 11554 4093 13500
rect 2983 11543 4093 11554
rect 4768 13500 5799 13540
rect 4768 11554 4818 13500
rect 5764 11554 5799 13500
rect 4768 11543 5799 11554
rect 6570 13500 7605 13540
rect 6570 11554 6618 13500
rect 7564 11554 7605 13500
rect 6570 11543 7605 11554
rect 8286 13500 9398 13540
rect 8286 11554 8318 13500
rect 9364 11554 9398 13500
rect 8286 11543 9398 11554
rect 10079 13500 11105 13540
rect 10079 11554 10118 13500
rect 11064 11554 11105 13500
rect 10079 11543 11105 11554
rect 11498 13122 11976 13490
rect 11498 13029 12288 13122
rect 11498 12958 11976 13029
rect 11498 11596 11524 12958
rect 11758 11596 11976 12958
rect 11498 11543 11976 11596
rect 373 2972 765 10972
rect 1055 2876 1101 11071
rect 2441 2876 2487 11071
rect 2823 2876 2869 11071
rect 4209 2876 4255 11071
rect 4591 2876 4637 11071
rect 5977 2876 6023 11071
rect 6359 2876 6405 11071
rect 7745 2876 7791 11071
rect 8127 2876 8173 11071
rect 9513 2876 9559 11071
rect 9895 2876 9941 11071
rect 11281 2876 11327 11071
rect 11615 2972 11989 10972
rect 400 1061 12013 2420
rect 92 1025 12288 1061
rect 92 257 460 1025
rect 11920 257 12288 1025
rect 12444 52 13136 14577
rect -756 -921 13136 52
rect -756 -1301 -64 -921
rect 12444 -1301 13136 -921
<< metal2 >>
rect -756 13411 -439 14820
rect 416 13388 816 15250
rect 1306 14563 2246 14820
rect 3078 14563 4018 14820
rect 4843 14563 5783 14820
rect 6612 14563 7552 14820
rect 8381 14563 9321 14820
rect 10147 14563 11087 14820
rect 11545 13388 11945 15250
rect 428 11472 816 13188
rect 11557 11472 11945 13188
rect 428 10188 1009 10972
rect 11373 10188 11954 10972
rect 428 6988 1009 9988
rect 11373 6988 11954 9988
rect 428 3788 1009 6788
rect 11373 3788 11954 6788
rect 428 2972 1009 3588
rect 11373 2972 11954 3588
rect 428 602 816 2414
rect 11557 602 11945 2414
use comp018green_out_drv_pleg_4T_X  comp018green_out_drv_pleg_4T_X_0
timestamp 1713338890
transform 1 0 731 0 1 2840
box 0 12 2080 8252
use comp018green_out_drv_pleg_4T_X  comp018green_out_drv_pleg_4T_X_1
timestamp 1713338890
transform -1 0 6347 0 1 2840
box 0 12 2080 8252
use comp018green_out_drv_pleg_4T_X  comp018green_out_drv_pleg_4T_X_2
timestamp 1713338890
transform 1 0 6035 0 1 2840
box 0 12 2080 8252
use comp018green_out_drv_pleg_4T_X  comp018green_out_drv_pleg_4T_X_3
timestamp 1713338890
transform -1 0 11651 0 1 2840
box 0 12 2080 8252
use comp018green_out_drv_pleg_4T_Y  comp018green_out_drv_pleg_4T_Y_0
timestamp 1713338890
transform 1 0 2499 0 1 2840
box 0 12 1196 8252
use comp018green_out_drv_pleg_4T_Y  comp018green_out_drv_pleg_4T_Y_1
timestamp 1713338890
transform -1 0 4579 0 1 2840
box 0 12 1196 8252
use comp018green_out_drv_pleg_4T_Y  comp018green_out_drv_pleg_4T_Y_2
timestamp 1713338890
transform 1 0 7803 0 1 2840
box 0 12 1196 8252
use comp018green_out_drv_pleg_4T_Y  comp018green_out_drv_pleg_4T_Y_3
timestamp 1713338890
transform -1 0 9883 0 1 2840
box 0 12 1196 8252
use M1_NWELL_CDNS_40661953145286  M1_NWELL_CDNS_40661953145286_0
timestamp 1713338890
transform 0 -1 6191 1 0 641
box -478 -6178 478 6178
use M1_NWELL_CDNS_40661953145345  M1_NWELL_CDNS_40661953145345_0
timestamp 1713338890
transform 1 0 476 0 1 13306
box -478 -278 478 278
use M1_NWELL_CDNS_40661953145345  M1_NWELL_CDNS_40661953145345_1
timestamp 1713338890
transform 1 0 11904 0 1 13306
box -478 -278 478 278
use M1_NWELL_CDNS_40661953145352  M1_NWELL_CDNS_40661953145352_0
timestamp 1713338890
transform 1 0 6209 0 1 1786
box -5678 -728 5678 728
use M1_NWELL_CDNS_40661953145361  M1_NWELL_CDNS_40661953145361_0
timestamp 1713338890
transform -1 0 276 0 1 7045
box -228 -6078 228 6078
use M1_NWELL_CDNS_40661953145361  M1_NWELL_CDNS_40661953145361_1
timestamp 1713338890
transform 1 0 12104 0 1 7045
box -228 -6078 228 6078
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_0
timestamp 1713338890
transform 1 0 1079 0 1 2842
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_1
timestamp 1713338890
transform 1 0 1079 0 1 11102
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_2
timestamp 1713338890
transform 1 0 2851 0 1 2842
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_3
timestamp 1713338890
transform 1 0 2465 0 1 2842
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_4
timestamp 1713338890
transform 1 0 2851 0 1 11102
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_5
timestamp 1713338890
transform 1 0 2465 0 1 11102
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_6
timestamp 1713338890
transform 1 0 4616 0 1 11102
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_7
timestamp 1713338890
transform 1 0 4225 0 1 11102
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_8
timestamp 1713338890
transform 1 0 4225 0 1 2842
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_9
timestamp 1713338890
transform 1 0 4616 0 1 2842
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_10
timestamp 1713338890
transform 1 0 5997 0 1 11102
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_11
timestamp 1713338890
transform 1 0 5997 0 1 2842
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_12
timestamp 1713338890
transform 1 0 6385 0 1 2842
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_13
timestamp 1713338890
transform 1 0 7767 0 1 2842
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_14
timestamp 1713338890
transform 1 0 8154 0 1 2842
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_15
timestamp 1713338890
transform 1 0 8154 0 1 11102
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_16
timestamp 1713338890
transform 1 0 6385 0 1 11102
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_17
timestamp 1713338890
transform 1 0 7767 0 1 11102
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_18
timestamp 1713338890
transform 1 0 9533 0 1 2842
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_19
timestamp 1713338890
transform 1 0 9920 0 1 2842
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_20
timestamp 1713338890
transform 1 0 9533 0 1 11102
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_21
timestamp 1713338890
transform 1 0 9920 0 1 11102
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_22
timestamp 1713338890
transform 1 0 11306 0 1 2842
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_23
timestamp 1713338890
transform 1 0 11306 0 1 11102
box -89 -42 89 42
use M1_PSUB_CDNS_69033583165675  M1_PSUB_CDNS_69033583165675_0
timestamp 1713338890
transform -1 0 -254 0 1 6808
box -201 -7695 201 7695
use M1_PSUB_CDNS_69033583165675  M1_PSUB_CDNS_69033583165675_1
timestamp 1713338890
transform -1 0 -566 0 1 6808
box -201 -7695 201 7695
use M1_PSUB_CDNS_69033583165675  M1_PSUB_CDNS_69033583165675_2
timestamp 1713338890
transform 1 0 12634 0 1 6808
box -201 -7695 201 7695
use M1_PSUB_CDNS_69033583165675  M1_PSUB_CDNS_69033583165675_3
timestamp 1713338890
transform -1 0 12946 0 1 6808
box -201 -7695 201 7695
use M1_PSUB_CDNS_69033583165676  M1_PSUB_CDNS_69033583165676_0
timestamp 1713338890
transform 0 -1 6191 1 0 -382
box -445 -6095 445 6095
use M1_PSUB_CDNS_69033583165677  M1_PSUB_CDNS_69033583165677_0
timestamp 1713338890
transform 0 -1 6190 1 0 -1111
box -201 -6945 201 6945
use M1_PSUB_CDNS_69033583165683  M1_PSUB_CDNS_69033583165683_0
timestamp 1713338890
transform 1 0 78 0 1 14916
box -845 -345 845 345
use M1_PSUB_CDNS_69033583165683  M1_PSUB_CDNS_69033583165683_1
timestamp 1713338890
transform 1 0 12302 0 1 14911
box -845 -345 845 345
use M1_PSUB_CDNS_69033583165684  M1_PSUB_CDNS_69033583165684_0
timestamp 1713338890
transform 1 0 1772 0 1 14466
box -495 -795 495 795
use M1_PSUB_CDNS_69033583165684  M1_PSUB_CDNS_69033583165684_1
timestamp 1713338890
transform 1 0 3544 0 1 14466
box -495 -795 495 795
use M1_PSUB_CDNS_69033583165684  M1_PSUB_CDNS_69033583165684_2
timestamp 1713338890
transform 1 0 5309 0 1 14466
box -495 -795 495 795
use M1_PSUB_CDNS_69033583165684  M1_PSUB_CDNS_69033583165684_3
timestamp 1713338890
transform 1 0 7078 0 1 14466
box -495 -795 495 795
use M1_PSUB_CDNS_69033583165684  M1_PSUB_CDNS_69033583165684_4
timestamp 1713338890
transform 1 0 10613 0 1 14466
box -495 -795 495 795
use M1_PSUB_CDNS_69033583165684  M1_PSUB_CDNS_69033583165684_5
timestamp 1713338890
transform 1 0 8847 0 1 14466
box -495 -795 495 795
use M2_M1_CDNS_6903358316539  M2_M1_CDNS_6903358316539_0
timestamp 1713338890
transform 1 0 616 0 1 14909
box -162 -286 162 286
use M2_M1_CDNS_6903358316539  M2_M1_CDNS_6903358316539_1
timestamp 1713338890
transform 1 0 11745 0 1 14909
box -162 -286 162 286
use M2_M1_CDNS_69033583165596  M2_M1_CDNS_69033583165596_0
timestamp 1713338890
transform 1 0 622 0 1 12339
box -162 -782 162 782
use M2_M1_CDNS_69033583165596  M2_M1_CDNS_69033583165596_1
timestamp 1713338890
transform 1 0 11751 0 1 12339
box -162 -782 162 782
use M2_M1_CDNS_69033583165679  M2_M1_CDNS_69033583165679_0
timestamp 1713338890
transform 1 0 570 0 1 5304
box -142 -1390 142 1390
use M2_M1_CDNS_69033583165679  M2_M1_CDNS_69033583165679_1
timestamp 1713338890
transform 1 0 570 0 1 8474
box -142 -1390 142 1390
use M2_M1_CDNS_69033583165679  M2_M1_CDNS_69033583165679_2
timestamp 1713338890
transform 1 0 11812 0 1 5304
box -142 -1390 142 1390
use M2_M1_CDNS_69033583165679  M2_M1_CDNS_69033583165679_3
timestamp 1713338890
transform 1 0 11812 0 1 8474
box -142 -1390 142 1390
use M2_M1_CDNS_69033583165680  M2_M1_CDNS_69033583165680_0
timestamp 1713338890
transform 1 0 570 0 1 10575
box -142 -298 142 298
use M2_M1_CDNS_69033583165680  M2_M1_CDNS_69033583165680_1
timestamp 1713338890
transform 1 0 11812 0 1 10575
box -142 -298 142 298
use M2_M1_CDNS_69033583165681  M2_M1_CDNS_69033583165681_0
timestamp 1713338890
transform 1 0 1776 0 1 14801
box -472 -410 472 410
use M2_M1_CDNS_69033583165681  M2_M1_CDNS_69033583165681_1
timestamp 1713338890
transform 1 0 3548 0 1 14801
box -472 -410 472 410
use M2_M1_CDNS_69033583165681  M2_M1_CDNS_69033583165681_2
timestamp 1713338890
transform 1 0 5313 0 1 14801
box -472 -410 472 410
use M2_M1_CDNS_69033583165681  M2_M1_CDNS_69033583165681_3
timestamp 1713338890
transform 1 0 7082 0 1 14801
box -472 -410 472 410
use M2_M1_CDNS_69033583165681  M2_M1_CDNS_69033583165681_4
timestamp 1713338890
transform 1 0 8851 0 1 14801
box -472 -410 472 410
use M2_M1_CDNS_69033583165681  M2_M1_CDNS_69033583165681_5
timestamp 1713338890
transform 1 0 10617 0 1 14801
box -472 -410 472 410
use M2_M1_CDNS_69033583165686  M2_M1_CDNS_69033583165686_0
timestamp 1713338890
transform 1 0 -585 0 1 14088
box -146 -632 146 632
use M2_M1_CDNS_69033583165687  M2_M1_CDNS_69033583165687_0
timestamp 1713338890
transform 1 0 570 0 1 3271
box -142 -246 142 246
use M2_M1_CDNS_69033583165687  M2_M1_CDNS_69033583165687_1
timestamp 1713338890
transform 1 0 11812 0 1 3271
box -142 -246 142 246
use M2_M1_CDNS_69033583165688  M2_M1_CDNS_69033583165688_0
timestamp 1713338890
transform 1 0 -618 0 1 -308
box -90 -610 90 610
use M2_M1_CDNS_69033583165689  M2_M1_CDNS_69033583165689_0
timestamp 1713338890
transform 1 0 622 0 1 1508
box -162 -906 162 906
use M2_M1_CDNS_69033583165689  M2_M1_CDNS_69033583165689_1
timestamp 1713338890
transform 1 0 11751 0 1 1508
box -162 -906 162 906
use M2_M1_CDNS_69033583165691  M2_M1_CDNS_69033583165691_0
timestamp 1713338890
transform -1 0 12969 0 1 -311
box -90 -662 90 662
use M3_M2_CDNS_69033583165560  M3_M2_CDNS_69033583165560_0
timestamp 1713338890
transform 1 0 616 0 1 14088
box -180 -677 180 677
use M3_M2_CDNS_69033583165560  M3_M2_CDNS_69033583165560_1
timestamp 1713338890
transform 1 0 11745 0 1 14088
box -180 -677 180 677
use M3_M2_CDNS_69033583165590  M3_M2_CDNS_69033583165590_0
timestamp 1713338890
transform 1 0 -585 0 1 14088
box -109 -677 109 677
use M3_M2_CDNS_69033583165590  M3_M2_CDNS_69033583165590_1
timestamp 1713338890
transform -1 0 12969 0 1 -311
box -109 -677 109 677
use M3_M2_CDNS_69033583165605  M3_M2_CDNS_69033583165605_0
timestamp 1713338890
transform 1 0 570 0 1 5292
box -109 -1458 109 1458
use M3_M2_CDNS_69033583165605  M3_M2_CDNS_69033583165605_1
timestamp 1713338890
transform 1 0 570 0 1 8474
box -109 -1458 109 1458
use M3_M2_CDNS_69033583165605  M3_M2_CDNS_69033583165605_2
timestamp 1713338890
transform 1 0 11812 0 1 5292
box -109 -1458 109 1458
use M3_M2_CDNS_69033583165605  M3_M2_CDNS_69033583165605_3
timestamp 1713338890
transform 1 0 11812 0 1 8474
box -109 -1458 109 1458
use M3_M2_CDNS_69033583165657  M3_M2_CDNS_69033583165657_0
timestamp 1713338890
transform 1 0 570 0 1 3281
box -109 -251 109 251
use M3_M2_CDNS_69033583165657  M3_M2_CDNS_69033583165657_1
timestamp 1713338890
transform 1 0 11812 0 1 3281
box -109 -251 109 251
use M3_M2_CDNS_69033583165678  M3_M2_CDNS_69033583165678_0
timestamp 1713338890
transform 1 0 1776 0 1 14578
box -464 -180 464 180
use M3_M2_CDNS_69033583165678  M3_M2_CDNS_69033583165678_1
timestamp 1713338890
transform 1 0 3548 0 1 14578
box -464 -180 464 180
use M3_M2_CDNS_69033583165678  M3_M2_CDNS_69033583165678_2
timestamp 1713338890
transform 1 0 5313 0 1 14578
box -464 -180 464 180
use M3_M2_CDNS_69033583165678  M3_M2_CDNS_69033583165678_3
timestamp 1713338890
transform 1 0 7082 0 1 14578
box -464 -180 464 180
use M3_M2_CDNS_69033583165678  M3_M2_CDNS_69033583165678_4
timestamp 1713338890
transform 1 0 8851 0 1 14578
box -464 -180 464 180
use M3_M2_CDNS_69033583165678  M3_M2_CDNS_69033583165678_5
timestamp 1713338890
transform 1 0 10617 0 1 14578
box -464 -180 464 180
use M3_M2_CDNS_69033583165682  M3_M2_CDNS_69033583165682_0
timestamp 1713338890
transform 1 0 622 0 1 1508
box -180 -819 180 819
use M3_M2_CDNS_69033583165682  M3_M2_CDNS_69033583165682_1
timestamp 1713338890
transform 1 0 622 0 1 12339
box -180 -819 180 819
use M3_M2_CDNS_69033583165682  M3_M2_CDNS_69033583165682_2
timestamp 1713338890
transform 1 0 11751 0 1 1508
box -180 -819 180 819
use M3_M2_CDNS_69033583165682  M3_M2_CDNS_69033583165682_3
timestamp 1713338890
transform 1 0 11751 0 1 12339
box -180 -819 180 819
use M3_M2_CDNS_69033583165685  M3_M2_CDNS_69033583165685_0
timestamp 1713338890
transform 1 0 570 0 1 10575
box -109 -322 109 322
use M3_M2_CDNS_69033583165685  M3_M2_CDNS_69033583165685_1
timestamp 1713338890
transform 1 0 11812 0 1 10575
box -109 -322 109 322
use M3_M2_CDNS_69033583165690  M3_M2_CDNS_69033583165690_0
timestamp 1713338890
transform 1 0 -618 0 1 -308
box -109 -606 109 606
use PMOS_4T_metal_stack  PMOS_4T_metal_stack_0
timestamp 1713338890
transform 1 0 809 0 1 2972
box -44 0 1584 8000
use PMOS_4T_metal_stack  PMOS_4T_metal_stack_1
timestamp 1713338890
transform 1 0 2577 0 1 2972
box -44 0 1584 8000
use PMOS_4T_metal_stack  PMOS_4T_metal_stack_2
timestamp 1713338890
transform 1 0 4345 0 1 2972
box -44 0 1584 8000
use PMOS_4T_metal_stack  PMOS_4T_metal_stack_3
timestamp 1713338890
transform 1 0 6113 0 1 2972
box -44 0 1584 8000
use PMOS_4T_metal_stack  PMOS_4T_metal_stack_4
timestamp 1713338890
transform 1 0 7881 0 1 2972
box -44 0 1584 8000
use PMOS_4T_metal_stack  PMOS_4T_metal_stack_5
timestamp 1713338890
transform 1 0 9649 0 1 2972
box -44 0 1584 8000
use PMOS_4T_metal_stack  PMOS_4T_metal_stack_6
timestamp 1713338890
transform -1 0 11573 0 1 2972
box -44 0 1584 8000
<< end >>
