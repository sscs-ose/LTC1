* NGSPICE file created from PFD_layout_flat.ext - technology: gf180mcuC

.subckt pex_PFD_layout VSS VREF VDIV PU PD VDD 
X0 DFF__1.CLK VREF.t0 VDD.t154 VDD.t153 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1 PD a_4617_1139# VDD.t152 VDD.t151 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X2 VDD buffer_mag_0.OUT DFF__0.nand2_3.OUT VDD.t9 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3 VSS buffer_mag_0.gf_inv_mag_1.IN buffer_mag_0.OUT VSS.t48 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X4 VSS nand2_0.IN1 a_4478_3188# VSS.t78 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X5 VSS buffer_mag_0.gf_inv_mag_1.IN buffer_mag_0.OUT VSS.t45 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.35u
X6 DFF__1.inv_0.OUT DFF__1.nand2_3.OUT VSS.t83 VSS.t82 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X7 a_3455_3092# DFF__1.nand2_5.OUT DFF__1.QB VSS.t106 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X8 DFF__1.nand2_3.OUT DFF__1.nand2_2.OUT VDD.t78 VDD.t77 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X9 a_4617_1139# buffer_loading_mag_1.IN VSS.t40 VSS.t39 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X10 DFF__0.nand2_1.IN1 buffer_mag_0.OUT a_1331_1976# VSS.t3 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X11 a_1327_4537# DFF__1.nand2_2.OUT VSS.t62 VSS.t61 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X12 VDD buffer_loading_mag_1.IN DFF__0.QB VDD.t54 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X13 DFF__1.nand2_1.IN1 buffer_mag_0.OUT a_1330_2902# VSS.t2 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X14 DFF__0.nand2_2.IN1 VDD.t15 VDD.t17 VDD.t16 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X15 nand2_0.IN1 DFF__1.QB a_3459_4589# VSS.t99 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X16 a_1328_341# DFF__0.nand2_2.OUT VSS.t54 VSS.t53 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X17 VSS a_4617_1139# PD.t5 VSS.t117 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X18 VSS buffer_loading_mag_1.IN a_4617_1139# VSS.t36 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X19 DFF__0.nand2_1.IN1 DFF__0.CLK VDD.t124 VDD.t123 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X20 VSS buffer_loading_mag_1.IN a_4617_1139# VSS.t33 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X21 buffer_mag_0.gf_inv_mag_1.IN buffer_mag_0.IN VDD.t29 VDD.t28 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X22 DFF__0.QB DFF__0.nand2_5.OUT VDD.t132 VDD.t131 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X23 DFF__1.nand2_2.IN1 DFF__1.nand2_5.OUT a_444_2859# VSS.t105 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X24 buffer_loading_mag_1.IN DFF__0.QB a_3460_289# VSS.t21 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X25 buffer_mag_0.IN nand2_0.IN1 VDD.t97 VDD.t96 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X26 a_3459_4589# DFF__1.nand2_2.IN2 VSS.t66 VSS.t65 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X27 a_6234_2632# nand2_0.IN1 buffer_mag_0.IN VSS.t77 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X28 DFF__1.nand2_1.IN1 DFF__1.CLK VDD.t19 VDD.t18 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X29 VDD DFF__1.QB nand2_0.IN1 VDD.t120 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X30 DFF__0.nand2_5.OUT DFF__0.nand2_3.OUT a_2560_1786# VSS.t86 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X31 VSS buffer_mag_0.IN buffer_mag_0.gf_inv_mag_1.IN VSS.t17 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X32 VDD a_4478_3188# PU.t3 VDD.t117 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X33 nand2_0.IN1 DFF__1.nand2_2.IN2 VDD.t82 VDD.t81 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X34 VSS buffer_mag_0.IN buffer_mag_0.gf_inv_mag_1.IN VSS.t14 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.35u
X35 a_2560_1786# DFF__0.nand2_1.IN1 VSS.t24 VSS.t23 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X36 PU a_4478_3188# VSS.t98 VSS.t97 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X37 VDD nand2_0.IN1 DFF__1.QB VDD.t93 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X38 DFF__1.nand2_2.IN1 VDD.t12 VDD.t14 VDD.t13 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X39 DFF__1.nand2_2.OUT DFF__1.nand2_2.IN2 VDD.t80 VDD.t79 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X40 DFF__1.CLK VREF.t1 VSS.t121 VSS.t120 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X41 a_610_4530# DFF__1.nand2_2.IN2 VSS.t64 VSS.t63 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X42 VDD nand2_0.IN1 a_4478_3188# VDD.t90 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X43 DFF__0.nand2_2.OUT DFF__0.nand2_2.IN2 VDD.t76 VDD.t75 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X44 a_4478_3188# nand2_0.IN1 VSS.t76 VSS.t75 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X45 VDD DFF__1.nand2_3.OUT DFF__1.nand2_5.OUT VDD.t100 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X46 a_4617_1139# buffer_loading_mag_1.IN VDD.t53 VDD.t52 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X47 VDD buffer_mag_0.gf_inv_mag_1.IN buffer_mag_0.OUT VDD.t64 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X48 VSS buffer_loading_mag_1.IN a_3456_1786# VSS.t30 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X49 DFF__1.nand2_5.OUT DFF__1.nand2_1.IN1 VDD.t142 VDD.t141 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X50 a_1331_1976# DFF__0.CLK VSS.t101 VSS.t100 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X51 VDD a_4617_1139# PD.t2 VDD.t148 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X52 VDD buffer_loading_mag_1.IN a_4617_1139# VDD.t49 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X53 buffer_mag_0.OUT buffer_mag_0.gf_inv_mag_1.IN VSS.t44 VSS.t43 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.35u
X54 VDD buffer_loading_mag_1.IN a_4617_1139# VDD.t46 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X55 a_3456_1786# DFF__0.nand2_5.OUT DFF__0.QB VSS.t104 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X56 a_1330_2902# DFF__1.CLK VSS.t9 VSS.t8 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X57 PD a_4617_1139# VSS.t116 VSS.t115 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X58 a_4617_1139# buffer_loading_mag_1.IN VSS.t29 VSS.t28 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X59 a_444_2859# VDD.t155 VSS.t7 VSS.t6 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X60 PU a_4478_3188# VDD.t116 VDD.t115 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X61 VDD buffer_mag_0.IN buffer_mag_0.gf_inv_mag_1.IN VDD.t25 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X62 buffer_mag_0.gf_inv_mag_1.IN buffer_mag_0.IN VSS.t13 VSS.t12 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.35u
X63 DFF__1.QB DFF__1.nand2_5.OUT VDD.t137 VDD.t136 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X64 DFF__0.nand2_3.OUT buffer_mag_0.OUT a_1328_341# VSS.t1 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X65 a_611_348# DFF__0.nand2_2.IN2 VSS.t60 VSS.t59 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X66 DFF__0.nand2_2.IN2 DFF__0.inv_0.OUT VDD.t72 VDD.t71 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X67 DFF__0.nand2_2.IN1 DFF__0.nand2_5.OUT a_445_2019# VSS.t103 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X68 a_4478_3188# nand2_0.IN1 VDD.t89 VDD.t88 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X69 VDD DFF__1.nand2_1.IN1 DFF__1.nand2_2.IN2 VDD.t138 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X70 DFF__0.nand2_3.OUT DFF__0.nand2_2.OUT VDD.t70 VDD.t69 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X71 VSS a_4478_3188# PU.t6 VSS.t94 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X72 VSS nand2_0.IN1 a_4478_3188# VSS.t72 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X73 DFF__1.nand2_2.IN2 DFF__1.inv_0.OUT VDD.t68 VDD.t67 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X74 VDD buffer_mag_0.gf_inv_mag_1.IN buffer_mag_0.OUT VDD.t61 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.35u
X75 PU a_4478_3188# VSS.t93 VSS.t92 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X76 a_4478_3188# nand2_0.IN1 VSS.t71 VSS.t70 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X77 DFF__1.inv_0.OUT DFF__1.nand2_3.OUT VDD.t99 VDD.t98 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X78 buffer_mag_0.OUT buffer_mag_0.gf_inv_mag_1.IN VSS.t42 VSS.t41 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X79 PD a_4617_1139# VDD.t147 VDD.t146 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X80 a_4617_1139# buffer_loading_mag_1.IN VDD.t45 VDD.t44 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X81 buffer_mag_0.OUT buffer_mag_0.gf_inv_mag_1.IN VDD.t60 VDD.t59 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.35u
X82 VSS a_4617_1139# PD.t4 VSS.t112 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X83 VDD DFF__0.nand2_1.IN1 DFF__0.nand2_2.IN2 VDD.t38 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X84 PD a_4617_1139# VSS.t111 VSS.t110 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X85 buffer_loading_mag_1.IN DFF__0.nand2_2.IN2 VDD.t74 VDD.t73 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X86 VDD DFF__0.nand2_2.IN1 DFF__0.nand2_2.OUT VDD.t30 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X87 VSS nand2_0.IN1 a_3455_3092# VSS.t67 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X88 VDD buffer_mag_0.IN buffer_mag_0.gf_inv_mag_1.IN VDD.t22 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.35u
X89 VDD buffer_mag_0.OUT DFF__1.nand2_3.OUT VDD.t6 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X90 a_2564_407# DFF__0.inv_0.OUT VSS.t56 VSS.t55 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X91 DFF__1.nand2_3.OUT buffer_mag_0.OUT a_1327_4537# VSS.t0 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X92 VDD DFF__0.nand2_5.OUT DFF__0.nand2_2.IN1 VDD.t128 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X93 buffer_mag_0.gf_inv_mag_1.IN buffer_mag_0.IN VSS.t11 VSS.t10 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X94 VDD buffer_mag_0.OUT DFF__0.nand2_1.IN1 VDD.t3 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X95 DFF__0.CLK VDIV.t0 VSS.t88 VSS.t87 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X96 DFF__1.nand2_2.IN2 DFF__1.nand2_1.IN1 a_2563_4471# VSS.t109 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X97 buffer_mag_0.gf_inv_mag_1.IN buffer_mag_0.IN VDD.t21 VDD.t20 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.35u
X98 VDD buffer_loading_mag_1.IN buffer_mag_0.IN VDD.t41 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X99 DFF__1.nand2_5.OUT DFF__1.nand2_3.OUT a_2559_3092# VSS.t81 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X100 a_445_2019# VDD.t156 VSS.t5 VSS.t4 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X101 VSS buffer_loading_mag_1.IN a_6234_2632# VSS.t25 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X102 VDD buffer_mag_0.OUT DFF__1.nand2_1.IN1 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X103 VDD a_4478_3188# PU.t1 VDD.t112 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X104 VDD nand2_0.IN1 a_4478_3188# VDD.t85 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X105 a_2563_4471# DFF__1.inv_0.OUT VSS.t52 VSS.t51 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X106 a_2559_3092# DFF__1.nand2_1.IN1 VSS.t108 VSS.t107 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X107 PU a_4478_3188# VDD.t111 VDD.t110 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X108 a_4478_3188# nand2_0.IN1 VDD.t84 VDD.t83 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X109 VDD DFF__0.QB buffer_loading_mag_1.IN VDD.t33 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X110 VDD DFF__0.nand2_3.OUT DFF__0.nand2_5.OUT VDD.t105 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X111 VSS a_4478_3188# PU.t4 VSS.t89 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X112 DFF__0.inv_0.OUT DFF__0.nand2_3.OUT VDD.t104 VDD.t103 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X113 DFF__0.CLK VDIV.t1 VDD.t109 VDD.t108 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X114 DFF__0.nand2_2.IN2 DFF__0.nand2_1.IN1 a_2564_407# VSS.t22 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X115 VDD a_4617_1139# PD.t0 VDD.t143 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X116 DFF__0.nand2_5.OUT DFF__0.nand2_1.IN1 VDD.t37 VDD.t36 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X117 VDD DFF__1.nand2_5.OUT DFF__1.nand2_2.IN1 VDD.t133 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X118 VDD DFF__1.nand2_2.IN1 DFF__1.nand2_2.OUT VDD.t125 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X119 DFF__0.nand2_2.OUT DFF__0.nand2_2.IN1 a_611_348# VSS.t20 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X120 a_3460_289# DFF__0.nand2_2.IN2 VSS.t58 VSS.t57 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X121 buffer_mag_0.OUT buffer_mag_0.gf_inv_mag_1.IN VDD.t58 VDD.t57 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X122 DFF__1.nand2_2.OUT DFF__1.nand2_2.IN1 a_610_4530# VSS.t102 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X123 DFF__0.inv_0.OUT DFF__0.nand2_3.OUT VSS.t85 VSS.t84 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
R0 VREF.n0 VREF.t0 25.4398
R1 VREF.n0 VREF.t1 17.6975
R2 VREF VREF.n0 4.24656
R3 VDD.n134 VDD.n133 91983.3
R4 VDD.t96 VDD.t148 9544.02
R5 VDD VDD.t108 551.043
R6 VDD.n149 VDD.n134 533.333
R7 VDD.n133 VDD.t153 443.07
R8 VDD.t67 VDD.n167 354.539
R9 VDD.t71 VDD.n44 354.539
R10 VDD.n1 VDD.t115 289.017
R11 VDD.n167 VDD 288.426
R12 VDD.n44 VDD 285.887
R13 VDD.n167 VDD.t98 280.245
R14 VDD.n44 VDD.t103 280.245
R15 VDD.n1 VDD.t90 265.897
R16 VDD.n92 VDD.t33 232.809
R17 VDD.n7 VDD.t120 232.809
R18 VDD.n95 VDD.t131 232.803
R19 VDD.n10 VDD.t136 232.803
R20 VDD.t110 VDD.t112 231.214
R21 VDD.t117 VDD.t110 231.214
R22 VDD.t115 VDD.t117 231.214
R23 VDD.t90 VDD.t88 231.214
R24 VDD.t88 VDD.t85 231.214
R25 VDD.t85 VDD.t83 231.214
R26 VDD.n15 VDD.t100 230.548
R27 VDD.n15 VDD.t141 230.548
R28 VDD.n43 VDD.t105 230.548
R29 VDD.n43 VDD.t36 230.548
R30 VDD.n94 VDD.t54 227.667
R31 VDD.n93 VDD.t73 227.667
R32 VDD.n8 VDD.t81 227.667
R33 VDD.n9 VDD.t93 227.667
R34 VDD.n22 VDD.t6 193.183
R35 VDD.n24 VDD.t125 193.183
R36 VDD.n117 VDD.t30 193.183
R37 VDD.n123 VDD.t128 193.183
R38 VDD.n111 VDD.t9 193.183
R39 VDD.n107 VDD.t3 193.183
R40 VDD.n28 VDD.t133 193.183
R41 VDD.n20 VDD.t0 193.183
R42 VDD.n64 VDD.t96 191.288
R43 VDD.t46 VDD.n83 175.573
R44 VDD.t64 VDD.t59 165.977
R45 VDD.t151 VDD.t20 164.123
R46 VDD.n150 VDD.n149 158.333
R47 VDD.t52 VDD.t46 152.673
R48 VDD.t49 VDD.t61 146.947
R49 VDD.n15 VDD.t138 143.345
R50 VDD.n43 VDD.t38 143.345
R51 VDD.t146 VDD.t28 137.405
R52 VDD.t148 VDD.t22 124.046
R53 VDD.n64 VDD.t41 111.743
R54 VDD.n22 VDD.t77 109.849
R55 VDD.n24 VDD.t79 109.849
R56 VDD.n117 VDD.t75 109.849
R57 VDD.n123 VDD.t16 109.849
R58 VDD.n111 VDD.t69 109.849
R59 VDD.n107 VDD.t123 109.849
R60 VDD.n28 VDD.t13 109.849
R61 VDD.n20 VDD.t18 109.849
R62 VDD.n63 VDD.t25 92.5578
R63 VDD.n168 VDD.t67 92.1507
R64 VDD.n45 VDD.t71 92.1507
R65 VDD.n150 VDD.n133 76.7332
R66 VDD.n84 VDD.t57 73.4738
R67 VDD.n84 VDD.t44 60.115
R68 VDD.n96 VDD.n95 59.3792
R69 VDD.n176 VDD.n10 59.3792
R70 VDD.t143 VDD.n63 58.2066
R71 VDD.n92 VDD.n91 56.5869
R72 VDD.n177 VDD.n7 56.5869
R73 VDD.t44 VDD.t64 32.4432
R74 VDD.n35 VDD.t15 30.9379
R75 VDD.n34 VDD.t12 30.9379
R76 VDD.n16 VDD.n15 30.7172
R77 VDD.n46 VDD.n43 30.7172
R78 VDD.t22 VDD.t146 28.6265
R79 VDD.n151 VDD.n150 28.1049
R80 VDD.n83 VDD.t20 26.7181
R81 VDD.n35 VDD.t156 21.6422
R82 VDD.n34 VDD.t155 21.6422
R83 VDD.t57 VDD.t49 19.0845
R84 VDD.n32 VDD.n25 17.9105
R85 VDD.t28 VDD.t143 15.2677
R86 VDD.n82 VDD.n55 12.9385
R87 VDD.n89 VDD.n88 11.1336
R88 VDD.n152 VDD.n151 11.0878
R89 VDD.n119 VDD.n116 10.7307
R90 VDD.n114 VDD.n113 8.95925
R91 VDD.n120 VDD.n119 7.3805
R92 VDD.n142 VDD.n137 7.026
R93 VDD.n168 VDD.n16 6.82644
R94 VDD.n46 VDD.n45 6.82644
R95 VDD.n182 VDD.n4 6.5905
R96 VDD.n0 VDD.t116 6.5805
R97 VDD.n68 VDD.n60 6.45726
R98 VDD.n80 VDD.t21 6.45726
R99 VDD.n78 VDD.n74 6.45726
R100 VDD.n88 VDD.t60 6.45726
R101 VDD.n116 VDD.t76 6.45146
R102 VDD.n124 VDD.n123 6.3005
R103 VDD.n85 VDD.n84 6.3005
R104 VDD.n65 VDD.n64 6.3005
R105 VDD.n108 VDD.n107 6.3005
R106 VDD.n112 VDD.n111 6.3005
R107 VDD.n118 VDD.n117 6.3005
R108 VDD.n136 VDD.n135 6.3005
R109 VDD.n135 VDD.n134 6.3005
R110 VDD.n29 VDD.n28 6.3005
R111 VDD.n157 VDD.n24 6.3005
R112 VDD.n21 VDD.n20 6.3005
R113 VDD.n160 VDD.n22 6.3005
R114 VDD.n185 VDD.n1 6.3005
R115 VDD.n101 VDD.n100 6.00445
R116 VDD.n129 VDD.n128 5.84038
R117 VDD.n127 VDD.n126 5.78069
R118 VDD.t61 VDD.t52 5.72569
R119 VDD.n94 VDD.n93 5.60274
R120 VDD.n9 VDD.n8 5.60274
R121 VDD.n50 VDD.n49 5.59693
R122 VDD.n110 VDD.n109 5.43849
R123 VDD.n105 VDD.t104 5.26145
R124 VDD VDD.t109 5.22218
R125 VDD.n21 VDD.t19 5.21805
R126 VDD.n124 VDD.t17 5.21701
R127 VDD.n164 VDD.n163 5.21429
R128 VDD.n27 VDD.n26 5.20057
R129 VDD.n122 VDD.n121 5.18056
R130 VDD.n136 VDD.t154 5.17584
R131 VDD.n166 VDD.t99 5.17584
R132 VDD.n30 VDD.t14 5.16674
R133 VDD.n65 VDD.n62 5.13813
R134 VDD.n40 VDD.t37 5.13746
R135 VDD.n38 VDD.t124 5.13746
R136 VDD.n113 VDD.t70 5.13746
R137 VDD.n155 VDD.t80 5.13746
R138 VDD.n159 VDD.t78 5.13746
R139 VDD.n17 VDD.t142 5.13746
R140 VDD.n90 VDD.n51 5.13586
R141 VDD.n97 VDD.t74 5.13586
R142 VDD.n175 VDD.t82 5.13586
R143 VDD.n178 VDD.n6 5.13586
R144 VDD.n106 VDD.n39 5.13287
R145 VDD.n115 VDD.n37 5.13287
R146 VDD.n158 VDD.n23 5.13287
R147 VDD.n19 VDD.n18 5.13287
R148 VDD.n172 VDD.n12 5.13287
R149 VDD.n98 VDD.t132 5.13129
R150 VDD.n89 VDD.n52 5.13129
R151 VDD.n179 VDD.n5 5.13129
R152 VDD.n174 VDD.t137 5.13129
R153 VDD.n102 VDD.t72 5.10854
R154 VDD.n14 VDD.t68 5.10854
R155 VDD.n173 VDD.n11 5.10445
R156 VDD.n66 VDD.t97 5.08866
R157 VDD.n99 VDD.n98 5.05272
R158 VDD.n147 VDD.n146 4.97759
R159 VDD.n174 VDD.n173 4.88931
R160 VDD.n148 VDD.n135 4.85833
R161 VDD.n180 VDD.t84 4.7565
R162 VDD.n184 VDD.n2 4.7565
R163 VDD.n87 VDD.t45 4.713
R164 VDD.n79 VDD.n73 4.713
R165 VDD.n72 VDD.t152 4.713
R166 VDD.n67 VDD.n61 4.713
R167 VDD.n120 VDD.n115 4.69819
R168 VDD.n141 VDD.n139 4.6705
R169 VDD.n154 VDD.n33 4.56932
R170 VDD.n148 VDD.n147 4.5005
R171 VDD.n149 VDD.n148 4.5005
R172 VDD.n106 VDD.n105 4.3827
R173 VDD.n114 VDD.n38 4.34898
R174 VDD.n166 VDD.n165 4.21364
R175 VDD VDD.n35 4.005
R176 VDD VDD.n34 4.005
R177 VDD.n180 VDD.n179 3.78851
R178 VDD.n57 VDD.t29 3.6405
R179 VDD.n57 VDD.n56 3.6405
R180 VDD.n54 VDD.t58 3.6405
R181 VDD.n54 VDD.n53 3.6405
R182 VDD.n146 VDD.n131 3.48009
R183 VDD.n122 VDD.n120 3.24518
R184 VDD.n70 VDD.n55 3.1505
R185 VDD.n63 VDD.n55 3.1505
R186 VDD.n82 VDD.n81 3.1505
R187 VDD.n83 VDD.n82 3.1505
R188 VDD.n42 VDD.n41 3.1505
R189 VDD.n45 VDD.n42 3.1505
R190 VDD.n48 VDD.n47 3.1505
R191 VDD.n47 VDD.n46 3.1505
R192 VDD.n132 VDD 3.1505
R193 VDD.n171 VDD.n13 3.1505
R194 VDD.n16 VDD.n13 3.1505
R195 VDD.n170 VDD.n169 3.1505
R196 VDD.n169 VDD.n168 3.1505
R197 VDD.n131 VDD.n130 3.13856
R198 VDD.n77 VDD.n76 2.893
R199 VDD.n69 VDD.n59 2.893
R200 VDD.n71 VDD.n57 2.81726
R201 VDD.n86 VDD.n54 2.81726
R202 VDD.n143 VDD.n142 2.73472
R203 VDD.n165 VDD.n164 2.72534
R204 VDD.n153 VDD.n131 2.2505
R205 VDD.t25 VDD.t151 1.9089
R206 VDD.n76 VDD.t53 1.8205
R207 VDD.n76 VDD.n75 1.8205
R208 VDD.n59 VDD.t147 1.8205
R209 VDD.n59 VDD.n58 1.8205
R210 VDD.n4 VDD.t89 1.8205
R211 VDD.n4 VDD.n3 1.8205
R212 VDD.n139 VDD.t111 1.8205
R213 VDD.n139 VDD.n138 1.8205
R214 VDD.n148 VDD.n132 1.67038
R215 VDD.n165 VDD.n19 1.39383
R216 VDD.n116 VDD.n36 0.7205
R217 VDD.n102 VDD.n101 0.7055
R218 VDD.n31 VDD.n27 0.636929
R219 VDD.n103 VDD.n102 0.6255
R220 VDD.n103 VDD 0.619037
R221 VDD VDD.n17 0.57316
R222 VDD.n146 VDD 0.566214
R223 VDD.n128 VDD 0.56151
R224 VDD.n129 VDD 0.550028
R225 VDD.n104 VDD.n41 0.513109
R226 VDD.n50 VDD.n40 0.43925
R227 VDD VDD.n145 0.372092
R228 VDD.n104 VDD.n40 0.352062
R229 VDD.n126 VDD.n125 0.336214
R230 VDD.n113 VDD.n112 0.257375
R231 VDD.n115 VDD.n114 0.238698
R232 VDD.n104 VDD.n48 0.220133
R233 VDD.n156 VDD.n33 0.171929
R234 VDD.n126 VDD 0.15032
R235 VDD.n159 VDD.n158 0.149994
R236 VDD.n169 VDD.n13 0.138205
R237 VDD.n47 VDD.n42 0.138205
R238 VDD.n182 VDD.n181 0.128315
R239 VDD.n126 VDD.n36 0.122835
R240 VDD.n141 VDD.n140 0.119239
R241 VDD.n95 VDD.n94 0.117546
R242 VDD.n10 VDD.n9 0.117546
R243 VDD.n154 VDD 0.117041
R244 VDD.n93 VDD.n92 0.111412
R245 VDD.n8 VDD.n7 0.111412
R246 VDD.n144 VDD.n143 0.0999848
R247 VDD.n105 VDD.n104 0.0918846
R248 VDD.n156 VDD.n25 0.0905
R249 VDD.n153 VDD.n152 0.0869056
R250 VDD VDD.n27 0.0830688
R251 VDD.n184 VDD.n183 0.0818025
R252 VDD.n30 VDD.n29 0.079766
R253 VDD.n145 VDD.n144 0.0789075
R254 VDD.n172 VDD 0.0786463
R255 VDD.n119 VDD 0.0721766
R256 VDD.n88 VDD.n87 0.0716397
R257 VDD.n158 VDD 0.0699068
R258 VDD.n69 VDD.n68 0.0653529
R259 VDD.n161 VDD.n19 0.0612407
R260 VDD.n66 VDD 0.0610515
R261 VDD.n142 VDD.n141 0.0594643
R262 VDD.n170 VDD.n14 0.0588902
R263 VDD.n125 VDD 0.0585645
R264 VDD.n72 VDD.n71 0.0574118
R265 VDD.n77 VDD 0.0570809
R266 VDD.n78 VDD.n77 0.0534412
R267 VDD.n79 VDD.n78 0.0531103
R268 VDD VDD.n0 0.0515504
R269 VDD.n160 VDD.n159 0.0512407
R270 VDD.n155 VDD.n154 0.0481695
R271 VDD.n87 VDD.n86 0.0455
R272 VDD VDD.n69 0.0451691
R273 VDD.n68 VDD.n67 0.0411985
R274 VDD.n185 VDD.n184 0.0409622
R275 VDD.n91 VDD.n90 0.040956
R276 VDD.n178 VDD.n177 0.040956
R277 VDD.n97 VDD.n96 0.0406629
R278 VDD.n176 VDD.n175 0.0406629
R279 VDD.n118 VDD.n36 0.0393024
R280 VDD.n110 VDD.n106 0.0383228
R281 VDD VDD.n72 0.0382206
R282 VDD VDD.n153 0.0380335
R283 VDD.n31 VDD.n30 0.0379096
R284 VDD.n67 VDD.n66 0.0372279
R285 VDD VDD.n110 0.036125
R286 VDD.n152 VDD 0.0341842
R287 VDD.n147 VDD.n136 0.0341842
R288 VDD.n50 VDD 0.0337609
R289 VDD.n108 VDD.n38 0.0317152
R290 VDD.n156 VDD.n155 0.0291017
R291 VDD.n151 VDD.n132 0.028942
R292 VDD VDD.n166 0.0284422
R293 VDD.n157 VDD.n156 0.0241441
R294 VDD.n128 VDD.n127 0.023
R295 VDD.n104 VDD.n103 0.0205
R296 VDD.n181 VDD.n180 0.0201639
R297 VDD.n130 VDD.n129 0.0200181
R298 VDD.n80 VDD.n79 0.0157206
R299 VDD.n164 VDD.n162 0.0151468
R300 VDD VDD.n80 0.0140662
R301 VDD.n183 VDD.n182 0.0133571
R302 VDD.n147 VDD 0.0120789
R303 VDD.n101 VDD.n99 0.0112339
R304 VDD.n162 VDD 0.00991177
R305 VDD.n105 VDD 0.00928049
R306 VDD.n127 VDD 0.00844118
R307 VDD.n32 VDD.n31 0.00809036
R308 VDD.n161 VDD 0.00716667
R309 VDD.n81 VDD 0.00711765
R310 VDD.n130 VDD 0.00700602
R311 VDD.n33 VDD.n32 0.00537952
R312 VDD.n140 VDD.n0 0.00465966
R313 VDD.n99 VDD.n50 0.00441304
R314 VDD VDD.n41 0.00441304
R315 VDD.n112 VDD 0.00425
R316 VDD.n110 VDD 0.00414557
R317 VDD.n27 VDD.n25 0.00371429
R318 VDD.n71 VDD.n70 0.00347794
R319 VDD.n86 VDD.n85 0.00347794
R320 VDD.n98 VDD.n97 0.00284528
R321 VDD.n175 VDD.n174 0.00284528
R322 VDD.n90 VDD.n89 0.00255212
R323 VDD.n179 VDD.n178 0.00255212
R324 VDD.n162 VDD.n161 0.00241489
R325 VDD.n173 VDD.n172 0.0022561
R326 VDD.n17 VDD.n14 0.0022561
R327 VDD.n101 VDD 0.00215138
R328 VDD VDD.n48 0.00215138
R329 VDD.n29 VDD 0.00215138
R330 VDD VDD.n185 0.00201261
R331 VDD.n70 VDD 0.00182353
R332 VDD.n81 VDD 0.00182353
R333 VDD.n85 VDD 0.00182353
R334 VDD VDD.n21 0.00167647
R335 VDD VDD.n124 0.00166129
R336 VDD VDD.n118 0.00157784
R337 VDD VDD.n171 0.00137805
R338 VDD.n171 VDD 0.00137805
R339 VDD VDD.n170 0.00137805
R340 VDD VDD.n157 0.00126271
R341 VDD VDD.n160 0.00124074
R342 VDD.n96 VDD 0.00108632
R343 VDD VDD.n176 0.00108632
R344 VDD.n125 VDD.n122 0.00106301
R345 VDD VDD.n108 0.000955696
R346 VDD VDD.n65 0.000830882
R347 VDD.n91 VDD 0.00079316
R348 VDD.n177 VDD 0.00079316
R349 PD.n4 PD.n3 3.416
R350 PD.n9 PD.n8 3.416
R351 PD.n3 PD.t4 3.2765
R352 PD.n3 PD.n2 3.2765
R353 PD.n8 PD.t5 3.2765
R354 PD.n8 PD.n7 3.2765
R355 PD.n4 PD.n1 3.013
R356 PD.n9 PD.n6 3.013
R357 PD.n1 PD.t0 1.8205
R358 PD.n1 PD.n0 1.8205
R359 PD.n6 PD.t2 1.8205
R360 PD.n6 PD.n5 1.8205
R361 PD.n9 PD.n4 0.445308
R362 PD PD.n9 0.310308
R363 VSS.n84 VSS.n83 127235
R364 VSS.n49 VSS.n48 118311
R365 VSS.n132 VSS.t59 16491.1
R366 VSS.n84 VSS.n49 14762
R367 VSS.n12 VSS.n11 12018.1
R368 VSS.n107 VSS.n106 9145.5
R369 VSS.n86 VSS.n85 8817.76
R370 VSS.n122 VSS.n121 6498.67
R371 VSS.n4 VSS.n3 6477.06
R372 VSS.t104 VSS.n107 6294.74
R373 VSS.n107 VSS.n26 5696.05
R374 VSS.n123 VSS.n122 5431.91
R375 VSS.t120 VSS.n133 3589.9
R376 VSS.t87 VSS.n132 3546.01
R377 VSS.n8 VSS.n7 3506.18
R378 VSS.n10 VSS.n9 3502.33
R379 VSS.n85 VSS.n84 3339.89
R380 VSS.n89 VSS.n86 3205.07
R381 VSS.n88 VSS.t21 2738.08
R382 VSS.n88 VSS.n87 2052.63
R383 VSS.n112 VSS.t65 1813.76
R384 VSS.n83 VSS.t43 1739.89
R385 VSS.n2 VSS.t84 1608.91
R386 VSS.n106 VSS.t57 1588.85
R387 VSS.n106 VSS.t22 1454.99
R388 VSS.t1 VSS.n4 1453.04
R389 VSS.t6 VSS.n144 1430.4
R390 VSS.t77 VSS.t14 1308.44
R391 VSS.n12 VSS.t53 1196.37
R392 VSS.t20 VSS.n12 1184.14
R393 VSS.n123 VSS.t3 1166.91
R394 VSS.t51 VSS.t82 1120.59
R395 VSS.t107 VSS.n123 1113.16
R396 VSS.n121 VSS.t0 908.602
R397 VSS.n121 VSS.n19 902.135
R398 VSS.n7 VSS.n6 870.861
R399 VSS.n11 VSS.n10 868.078
R400 VSS.t61 VSS.n119 748.808
R401 VSS.n119 VSS.t102 743.01
R402 VSS.n26 VSS.n25 690.782
R403 VSS.n70 VSS.t12 688.312
R404 VSS.t28 VSS.n89 644.163
R405 VSS.n135 VSS.t87 586.688
R406 VSS.n4 VSS.n2 584.657
R407 VSS.n134 VSS.t120 579
R408 VSS.t94 VSS.t92 519.481
R409 VSS.t97 VSS.t17 457.793
R410 VSS.n30 VSS.t110 456.543
R411 VSS.n70 VSS.t78 451.3
R412 VSS.n105 VSS.t21 443.183
R413 VSS.t45 VSS.t75 431.818
R414 VSS.n5 VSS.t1 412.699
R415 VSS.n13 VSS.t20 408.913
R416 VSS.t89 VSS.n69 399.351
R417 VSS.t22 VSS.n0 379.562
R418 VSS.t70 VSS.t48 340.909
R419 VSS.t115 VSS.t117 333.548
R420 VSS.t112 VSS.t115 333.548
R421 VSS.t110 VSS.t112 333.548
R422 VSS.t33 VSS.t39 333.548
R423 VSS.t39 VSS.t36 333.548
R424 VSS.t36 VSS.t28 333.548
R425 VSS.t57 VSS.n105 295.455
R426 VSS.t72 VSS.n82 282.469
R427 VSS.n54 VSS.t77 279.221
R428 VSS.t53 VSS.n5 275.132
R429 VSS.t59 VSS.n13 272.608
R430 VSS.n111 VSS.t99 269.663
R431 VSS.n113 VSS.t109 268.272
R432 VSS.t0 VSS.n120 258.065
R433 VSS.t102 VSS.n118 256.579
R434 VSS.n0 VSS.t55 253.042
R435 VSS.t109 VSS.n112 245.917
R436 VSS.n146 VSS.t105 240.087
R437 VSS.n90 VSS.t33 231.399
R438 VSS.n89 VSS.n88 225.144
R439 VSS.n127 VSS.t2 225.036
R440 VSS.t43 VSS.t70 224.026
R441 VSS.n56 VSS.t25 207.792
R442 VSS.n108 VSS.t104 197.663
R443 VSS.n125 VSS.t81 197.663
R444 VSS.t65 VSS.n111 179.775
R445 VSS.n113 VSS.t51 178.849
R446 VSS.t48 VSS.t72 178.571
R447 VSS.n120 VSS.t61 172.043
R448 VSS.n118 VSS.t63 171.054
R449 VSS.n145 VSS.t4 159.215
R450 VSS.n128 VSS.t100 149.236
R451 VSS.t75 VSS.t41 133.118
R452 VSS.n24 VSS.t67 131.083
R453 VSS.n124 VSS.t23 131.083
R454 VSS.t12 VSS.t97 107.144
R455 VSS.n69 VSS.t10 103.897
R456 VSS.n82 VSS.t41 103.897
R457 VSS.t78 VSS.t45 87.6628
R458 VSS.n26 VSS.t86 64.9263
R459 VSS.t17 VSS.t89 61.6888
R460 VSS.n144 VSS.n135 50.5448
R461 VSS.t14 VSS.t94 29.2213
R462 VSS.n55 VSS.n54 25.9745
R463 VSS.t82 VSS.n19 25.151
R464 VSS.t92 VSS.t10 16.2343
R465 VSS.n143 VSS.n142 10.5926
R466 VSS.n1 VSS.t85 9.36866
R467 VSS.n138 VSS.t121 9.36804
R468 VSS.n155 VSS.t88 9.36804
R469 VSS.n116 VSS.t83 9.36804
R470 VSS VSS.n53 7.23958
R471 VSS.n169 VSS.t56 7.19156
R472 VSS.n17 VSS.t101 7.19156
R473 VSS.n114 VSS.t52 7.19156
R474 VSS.n129 VSS.t9 7.19156
R475 VSS.n126 VSS.t24 7.18989
R476 VSS.n102 VSS.n101 7.18989
R477 VSS.n109 VSS.n22 7.18989
R478 VSS.n18 VSS.t108 7.18989
R479 VSS VSS.t64 7.18966
R480 VSS.n117 VSS.t62 7.12323
R481 VSS.n164 VSS.t60 7.12323
R482 VSS.n131 VSS.t7 7.12156
R483 VSS.n147 VSS.t5 7.11989
R484 VSS.n165 VSS.t54 7.11156
R485 VSS.n20 VSS.t66 7.03656
R486 VSS.n104 VSS.t58 7.02489
R487 VSS.n59 VSS.n52 6.64949
R488 VSS.n35 VSS.n34 6.61132
R489 VSS.n38 VSS.t111 6.61132
R490 VSS.n93 VSS.n29 6.61132
R491 VSS.n96 VSS.t29 6.61132
R492 VSS.n65 VSS.t98 6.59043
R493 VSS.n72 VSS.n51 6.59043
R494 VSS.n78 VSS.t71 6.59043
R495 VSS.n56 VSS.n55 6.49401
R496 VSS.n103 VSS.n102 6.46225
R497 VSS VSS.n110 6.32556
R498 VSS.n168 VSS.n1 5.8505
R499 VSS.n111 VSS 5.2005
R500 VSS VSS.n113 5.2005
R501 VSS.n115 VSS.n19 5.2005
R502 VSS.n120 VSS 5.2005
R503 VSS VSS.n125 5.2005
R504 VSS.n24 VSS 5.2005
R505 VSS.n105 VSS 5.2005
R506 VSS.n92 VSS.n91 5.2005
R507 VSS.n91 VSS.n90 5.2005
R508 VSS.n47 VSS.n45 5.2005
R509 VSS.n47 VSS.n46 5.2005
R510 VSS VSS.n56 5.2005
R511 VSS.n71 VSS.n70 5.2005
R512 VSS.n82 VSS.n81 5.2005
R513 VSS.n69 VSS.n68 5.2005
R514 VSS.n124 VSS 5.2005
R515 VSS VSS.n108 5.2005
R516 VSS.n145 VSS 5.2005
R517 VSS VSS.n146 5.2005
R518 VSS.n161 VSS.n160 5.2005
R519 VSS.n160 VSS.n159 5.2005
R520 VSS.n142 VSS.n140 5.2005
R521 VSS.n142 VSS.n141 5.2005
R522 VSS.n137 VSS.n136 5.2005
R523 VSS.n118 VSS 5.2005
R524 VSS VSS.n128 5.2005
R525 VSS.n127 VSS 5.2005
R526 VSS VSS.n13 5.2005
R527 VSS VSS.n5 5.2005
R528 VSS VSS.n0 5.2005
R529 VSS.n167 VSS.n2 5.2005
R530 VSS.n99 VSS.n98 5.07824
R531 VSS.n58 VSS.n57 5.06621
R532 VSS.n64 VSS.t13 5.04745
R533 VSS.n73 VSS.n50 5.02656
R534 VSS.n21 VSS.t44 4.99985
R535 VSS.n31 VSS.n30 4.5005
R536 VSS.n143 VSS.n15 4.5005
R537 VSS.n144 VSS.n143 4.5005
R538 VSS.n163 VSS.n14 3.90872
R539 VSS.n163 VSS.n162 3.69451
R540 VSS.n79 VSS.n77 3.37758
R541 VSS.n66 VSS.n63 3.37758
R542 VSS.n36 VSS.n33 3.33532
R543 VSS.n97 VSS.n95 3.33532
R544 VSS.n67 VSS.n61 3.31443
R545 VSS.n80 VSS.n75 3.31443
R546 VSS.n33 VSS.t116 3.2765
R547 VSS.n33 VSS.n32 3.2765
R548 VSS.n95 VSS.t40 3.2765
R549 VSS.n95 VSS.n94 3.2765
R550 VSS.n61 VSS.t93 3.2765
R551 VSS.n61 VSS.n60 3.2765
R552 VSS.n75 VSS.t76 3.2765
R553 VSS.n75 VSS.n74 3.2765
R554 VSS.n130 VSS.n16 2.85704
R555 VSS.n149 VSS.n148 2.69391
R556 VSS.n9 VSS.n8 2.61336
R557 VSS.t105 VSS.t103 2.52772
R558 VSS.n146 VSS.n145 2.52772
R559 VSS.t4 VSS.t6 2.52772
R560 VSS.n135 VSS.n134 2.52772
R561 VSS.n162 VSS.n161 2.37524
R562 VSS.t3 VSS.t2 2.3693
R563 VSS.n128 VSS.n127 2.3693
R564 VSS.t100 VSS.t8 2.3693
R565 VSS.t67 VSS.t30 2.08117
R566 VSS.n108 VSS.n24 2.08117
R567 VSS.t104 VSS.t106 2.08117
R568 VSS.t86 VSS.t81 2.08117
R569 VSS.n125 VSS.n124 2.08117
R570 VSS.t23 VSS.t107 2.08117
R571 VSS.n162 VSS.n15 1.80706
R572 VSS.n77 VSS.t42 1.6385
R573 VSS.n77 VSS.n76 1.6385
R574 VSS.n63 VSS.t11 1.6385
R575 VSS.n63 VSS.n62 1.6385
R576 VSS.t30 VSS.n23 1.51003
R577 VSS.n43 VSS.n42 1.50472
R578 VSS.n153 VSS.n151 1.49578
R579 VSS.n91 VSS.n47 1.48535
R580 VSS.n47 VSS.n31 1.37929
R581 VSS VSS.n18 0.841511
R582 VSS VSS.n126 0.840934
R583 VSS VSS.n17 0.545498
R584 VSS VSS.n129 0.545498
R585 VSS.n160 VSS.n158 0.368921
R586 VSS.n149 VSS.n16 0.349591
R587 VSS.n150 VSS.n149 0.325955
R588 VSS VSS.n20 0.278241
R589 VSS VSS.n116 0.256849
R590 VSS VSS.n117 0.22033
R591 VSS.n110 VSS.n109 0.206733
R592 VSS.n158 VSS.n157 0.178049
R593 VSS.n164 VSS.n163 0.165962
R594 VSS.n97 VSS.n96 0.161394
R595 VSS.n36 VSS.n35 0.160891
R596 VSS.n98 VSS.n93 0.158377
R597 VSS.n104 VSS 0.152356
R598 VSS.n66 VSS.n65 0.137706
R599 VSS.n166 VSS 0.137163
R600 VSS.n38 VSS.n37 0.136757
R601 VSS.n165 VSS 0.132962
R602 VSS.n166 VSS.n1 0.127741
R603 VSS VSS.n73 0.125794
R604 VSS.n79 VSS.n78 0.121824
R605 VSS VSS.n17 0.118573
R606 VSS.n129 VSS 0.118573
R607 VSS.n58 VSS 0.118373
R608 VSS VSS.n114 0.114176
R609 VSS VSS.n59 0.110913
R610 VSS.n99 VSS.n28 0.0983462
R611 VSS.n103 VSS.n100 0.0976538
R612 VSS.n142 VSS.n137 0.0926053
R613 VSS VSS.n15 0.0905
R614 VSS.n28 VSS.n27 0.0895769
R615 VSS.n78 VSS.n21 0.0881535
R616 VSS.n102 VSS 0.0874595
R617 VSS.n126 VSS 0.0874595
R618 VSS.n109 VSS 0.0874595
R619 VSS VSS.n18 0.0874595
R620 VSS.n100 VSS.n99 0.0861154
R621 VSS VSS.n131 0.0857318
R622 VSS.n147 VSS 0.0856259
R623 VSS.n156 VSS.n155 0.0644474
R624 VSS.n139 VSS.n138 0.0636579
R625 VSS.n169 VSS.n168 0.0556471
R626 VSS.n117 VSS 0.055266
R627 VSS VSS.n20 0.055266
R628 VSS VSS.n103 0.0533462
R629 VSS.n110 VSS.n21 0.0530664
R630 VSS.n114 VSS 0.05
R631 VSS.n131 VSS.n130 0.0499702
R632 VSS.n148 VSS.n147 0.0496447
R633 VSS.n39 VSS.n38 0.044243
R634 VSS.n71 VSS 0.0362353
R635 VSS.n59 VSS.n58 0.0356813
R636 VSS VSS.n104 0.0335
R637 VSS VSS.n165 0.0335
R638 VSS VSS.n164 0.0335
R639 VSS VSS.n169 0.0320441
R640 VSS.n42 VSS.n41 0.0315345
R641 VSS.n151 VSS.n150 0.0295909
R642 VSS.n151 VSS.n14 0.0286818
R643 VSS.n116 VSS.n115 0.0283244
R644 VSS.n155 VSS.n154 0.0257632
R645 VSS.n37 VSS.n36 0.0251369
R646 VSS.n72 VSS 0.0238824
R647 VSS.n68 VSS.n67 0.0203529
R648 VSS.n64 VSS 0.0203529
R649 VSS.n80 VSS.n79 0.0203529
R650 VSS.n154 VSS.n153 0.0184442
R651 VSS.n168 VSS 0.0181471
R652 VSS.n93 VSS.n92 0.017595
R653 VSS.n65 VSS.n64 0.0168235
R654 VSS.n40 VSS.n39 0.0145782
R655 VSS.n45 VSS.n44 0.0135726
R656 VSS.n167 VSS.n166 0.0113088
R657 VSS.n92 VSS 0.0100531
R658 VSS.n153 VSS.n152 0.00972292
R659 VSS.n44 VSS.n43 0.00834709
R660 VSS.n73 VSS.n72 0.00711765
R661 VSS.n68 VSS 0.00535294
R662 VSS.n81 VSS 0.00535294
R663 VSS.n45 VSS 0.00502514
R664 VSS.n43 VSS.n40 0.0046963
R665 VSS.n67 VSS.n66 0.00447059
R666 VSS VSS.n71 0.00447059
R667 VSS.n81 VSS.n80 0.00447059
R668 VSS.n98 VSS.n97 0.00301397
R669 VSS.n161 VSS 0.00286842
R670 VSS.n140 VSS 0.00128947
R671 VSS.n140 VSS.n139 0.00128947
R672 VSS VSS.n156 0.00128947
R673 VSS.n115 VSS 0.000843511
R674 VSS VSS.n167 0.000720588
R675 PU.n4 PU.n3 3.416
R676 PU.n9 PU.n8 3.416
R677 PU.n3 PU.t4 3.2765
R678 PU.n3 PU.n2 3.2765
R679 PU.n8 PU.t6 3.2765
R680 PU.n8 PU.n7 3.2765
R681 PU.n4 PU.n1 3.013
R682 PU.n9 PU.n6 3.013
R683 PU.n1 PU.t3 1.8205
R684 PU.n1 PU.n0 1.8205
R685 PU.n6 PU.t1 1.8205
R686 PU.n6 PU.n5 1.8205
R687 PU.n9 PU.n4 0.445308
R688 PU PU.n9 0.310308
R689 VDIV.n0 VDIV.t1 25.4398
R690 VDIV.n0 VDIV.t0 17.6975
R691 VDIV VDIV.n0 4.24656
C0 DFF__0.nand2_2.IN1 buffer_mag_0.OUT 0.0963f
C1 a_610_4530# VDD 5.14e-19
C2 DFF__1.nand2_3.OUT DFF__1.nand2_2.IN2 0.0986f
C3 a_445_2019# DFF__1.CLK 1.82e-19
C4 buffer_mag_0.gf_inv_mag_1.IN a_4617_1139# 8.3e-19
C5 DFF__1.nand2_5.OUT DFF__1.inv_0.OUT 1.02e-21
C6 DFF__1.QB buffer_mag_0.OUT 1.19e-19
C7 VREF VDD 0.211f
C8 buffer_mag_0.OUT DFF__1.CLK 0.0528f
C9 a_1327_4537# DFF__1.nand2_2.IN2 0.0144f
C10 a_3460_289# DFF__0.nand2_3.OUT 9.07e-21
C11 DFF__1.nand2_2.OUT DFF__1.nand2_3.OUT 0.106f
C12 DFF__0.nand2_2.IN1 VDD 0.918f
C13 a_3460_289# buffer_loading_mag_1.IN 0.069f
C14 DFF__0.CLK VDIV 0.115f
C15 DFF__0.nand2_1.IN1 DFF__1.nand2_5.OUT 2.09e-19
C16 DFF__1.nand2_3.OUT DFF__1.inv_0.OUT 0.142f
C17 DFF__1.nand2_2.OUT a_1327_4537# 0.00364f
C18 buffer_loading_mag_1.IN PD 0.0238f
C19 buffer_mag_0.OUT buffer_mag_0.gf_inv_mag_1.IN 0.389f
C20 DFF__0.CLK DFF__0.nand2_1.IN1 0.114f
C21 DFF__1.QB VDD 1.14f
C22 DFF__0.nand2_2.OUT DFF__0.nand2_5.OUT 1.33e-19
C23 DFF__1.CLK VDD 1.12f
C24 DFF__1.nand2_2.IN1 DFF__1.nand2_2.IN2 0.0753f
C25 a_1327_4537# DFF__1.inv_0.OUT 1.29e-20
C26 DFF__1.QB nand2_0.IN1 0.618f
C27 DFF__1.nand2_5.OUT DFF__1.nand2_1.IN1 0.176f
C28 DFF__0.CLK a_1331_1976# 0.00347f
C29 buffer_mag_0.OUT a_1330_2902# 0.00519f
C30 a_4478_3188# VDD 1.2f
C31 DFF__0.nand2_5.OUT DFF__1.inv_0.OUT 8.72e-22
C32 a_611_348# DFF__0.nand2_2.IN1 0.00348f
C33 DFF__1.QB a_3459_4589# 0.00619f
C34 nand2_0.IN1 a_4478_3188# 0.365f
C35 DFF__0.nand2_1.IN1 DFF__1.nand2_3.OUT 4.77e-22
C36 a_2563_4471# VDD 3.22e-19
C37 DFF__1.nand2_2.IN1 DFF__1.nand2_2.OUT 0.451f
C38 buffer_mag_0.gf_inv_mag_1.IN VDD 1f
C39 nand2_0.IN1 a_2563_4471# 1.06e-19
C40 DFF__0.nand2_3.OUT DFF__1.nand2_5.OUT 1.36e-19
C41 buffer_mag_0.gf_inv_mag_1.IN nand2_0.IN1 0.292f
C42 buffer_mag_0.OUT DFF__1.nand2_2.IN2 0.0259f
C43 DFF__1.nand2_3.OUT DFF__1.nand2_1.IN1 0.39f
C44 DFF__1.nand2_2.IN1 DFF__1.inv_0.OUT 4.23e-20
C45 a_1330_2902# VDD 4.86e-19
C46 DFF__0.nand2_1.IN1 DFF__0.nand2_5.OUT 0.176f
C47 DFF__0.nand2_1.IN1 DFF__0.inv_0.OUT 0.0551f
C48 a_2559_3092# DFF__1.nand2_1.IN1 0.00376f
C49 DFF__0.nand2_2.OUT DFF__0.nand2_2.IN2 0.159f
C50 DFF__0.nand2_2.OUT buffer_mag_0.OUT 0.0494f
C51 a_1331_1976# DFF__0.nand2_5.OUT 3.83e-19
C52 DFF__1.nand2_2.OUT buffer_mag_0.OUT 0.0494f
C53 DFF__0.nand2_5.OUT DFF__1.nand2_1.IN1 1.69e-19
C54 DFF__0.nand2_3.OUT DFF__1.nand2_3.OUT 5.53e-19
C55 buffer_mag_0.IN a_6234_2632# 0.0691f
C56 DFF__1.nand2_2.IN2 VDD 0.803f
C57 buffer_mag_0.OUT DFF__1.inv_0.OUT 0.00685f
C58 buffer_mag_0.IN a_4617_1139# 0.0088f
C59 DFF__1.nand2_2.IN2 nand2_0.IN1 0.117f
C60 PU VDD 0.588f
C61 DFF__1.nand2_2.IN1 DFF__1.nand2_1.IN1 0.00714f
C62 PU nand2_0.IN1 0.00662f
C63 DFF__0.nand2_2.OUT VDD 0.39f
C64 DFF__0.nand2_3.OUT DFF__0.nand2_5.OUT 0.42f
C65 DFF__1.nand2_2.IN2 a_3459_4589# 0.00411f
C66 DFF__1.nand2_2.OUT VDD 0.396f
C67 DFF__0.nand2_3.OUT DFF__0.inv_0.OUT 0.142f
C68 DFF__0.nand2_1.IN1 DFF__0.nand2_2.IN2 0.459f
C69 DFF__0.nand2_1.IN1 buffer_mag_0.OUT 0.487f
C70 buffer_loading_mag_1.IN DFF__0.nand2_5.OUT 0.0652f
C71 DFF__1.inv_0.OUT VDD 0.347f
C72 a_610_4530# DFF__1.CLK 1.27e-19
C73 a_1331_1976# DFF__0.nand2_2.IN2 2.82e-20
C74 buffer_loading_mag_1.IN DFF__0.inv_0.OUT 5.29e-19
C75 a_1328_341# DFF__0.inv_0.OUT 1.29e-20
C76 DFF__1.inv_0.OUT nand2_0.IN1 5.29e-19
C77 a_1331_1976# buffer_mag_0.OUT 0.00519f
C78 buffer_mag_0.OUT buffer_mag_0.IN 0.00294f
C79 buffer_loading_mag_1.IN a_6234_2632# 0.00403f
C80 buffer_mag_0.OUT DFF__1.nand2_1.IN1 0.487f
C81 VREF DFF__1.CLK 0.115f
C82 DFF__0.nand2_2.OUT a_611_348# 0.069f
C83 buffer_loading_mag_1.IN a_4617_1139# 0.453f
C84 VDIV VDD 0.196f
C85 DFF__0.nand2_1.IN1 VDD 1.3f
C86 buffer_loading_mag_1.IN a_3456_1786# 0.00347f
C87 DFF__0.nand2_2.IN1 DFF__1.CLK 4.28e-19
C88 DFF__0.nand2_3.OUT DFF__0.nand2_2.IN2 0.0984f
C89 DFF__0.nand2_3.OUT buffer_mag_0.OUT 0.889f
C90 buffer_mag_0.IN VDD 0.838f
C91 a_1331_1976# VDD 4.85e-19
C92 DFF__1.nand2_1.IN1 VDD 1.3f
C93 buffer_mag_0.IN nand2_0.IN1 0.44f
C94 DFF__0.CLK DFF__1.nand2_5.OUT 6.58e-19
C95 buffer_loading_mag_1.IN DFF__0.nand2_2.IN2 0.117f
C96 a_1328_341# DFF__0.nand2_2.IN2 0.0144f
C97 DFF__1.nand2_1.IN1 nand2_0.IN1 0.0119f
C98 buffer_mag_0.OUT buffer_loading_mag_1.IN 0.0112f
C99 a_1328_341# buffer_mag_0.OUT 0.00348f
C100 DFF__1.QB a_4478_3188# 0.00174f
C101 DFF__1.nand2_5.OUT a_444_2859# 0.00432f
C102 PD a_4617_1139# 0.332f
C103 DFF__1.nand2_1.IN1 a_3459_4589# 1.63e-20
C104 DFF__0.nand2_1.IN1 a_2560_1786# 0.00376f
C105 DFF__0.CLK a_444_2859# 1.82e-19
C106 a_610_4530# DFF__1.nand2_2.IN2 0.0175f
C107 DFF__0.nand2_3.OUT VDD 0.886f
C108 DFF__1.nand2_5.OUT DFF__1.nand2_3.OUT 0.42f
C109 DFF__1.nand2_5.OUT a_3455_3092# 0.00454f
C110 buffer_loading_mag_1.IN VDD 2.79f
C111 a_1330_2902# DFF__1.CLK 0.00347f
C112 buffer_mag_0.gf_inv_mag_1.IN a_4478_3188# 0.002f
C113 a_1328_341# VDD 3.14e-19
C114 DFF__1.nand2_5.OUT a_2559_3092# 0.0703f
C115 a_3460_289# DFF__0.nand2_2.IN2 0.00411f
C116 buffer_loading_mag_1.IN nand2_0.IN1 0.28f
C117 DFF__1.nand2_2.OUT a_610_4530# 0.069f
C118 a_2564_407# DFF__0.nand2_1.IN1 0.00384f
C119 DFF__0.nand2_5.OUT DFF__1.nand2_5.OUT 1.45f
C120 a_611_348# DFF__0.nand2_3.OUT 1.26e-20
C121 DFF__0.CLK DFF__0.nand2_5.OUT 0.115f
C122 DFF__1.nand2_5.OUT DFF__0.inv_0.OUT 8.72e-22
C123 DFF__0.nand2_3.OUT a_2560_1786# 0.00594f
C124 DFF__1.QB DFF__1.nand2_2.IN2 0.147f
C125 DFF__1.nand2_2.IN2 DFF__1.CLK 0.0318f
C126 a_1327_4537# DFF__1.nand2_3.OUT 0.069f
C127 DFF__0.nand2_1.IN1 DFF__0.QB 0.273f
C128 a_2559_3092# DFF__1.nand2_3.OUT 0.00594f
C129 DFF__1.nand2_2.IN1 DFF__1.nand2_5.OUT 0.492f
C130 DFF__0.nand2_2.OUT DFF__0.nand2_2.IN1 0.451f
C131 DFF__0.CLK DFF__1.nand2_2.IN1 4.55e-19
C132 a_3460_289# VDD 3.15e-19
C133 DFF__0.nand2_5.OUT DFF__1.nand2_3.OUT 1.35e-19
C134 PD VDD 0.645f
C135 PU a_4478_3188# 0.332f
C136 VREF VDIV 3.36e-19
C137 DFF__1.nand2_2.OUT DFF__1.CLK 0.00375f
C138 PD nand2_0.IN1 8.89e-20
C139 DFF__1.nand2_2.IN2 a_2563_4471# 0.0769f
C140 DFF__1.nand2_2.IN1 a_444_2859# 0.069f
C141 a_2564_407# DFF__0.nand2_3.OUT 2.09e-19
C142 DFF__1.QB DFF__1.inv_0.OUT 0.00316f
C143 DFF__0.CLK a_445_2019# 9.59e-19
C144 DFF__1.nand2_2.IN1 DFF__1.nand2_3.OUT 0.0185f
C145 buffer_mag_0.OUT DFF__1.nand2_5.OUT 0.391f
C146 a_1330_2902# DFF__1.nand2_2.IN2 2.82e-20
C147 a_2564_407# buffer_loading_mag_1.IN 1.06e-19
C148 DFF__0.CLK DFF__0.nand2_2.IN2 0.0318f
C149 DFF__0.CLK buffer_mag_0.OUT 0.0528f
C150 DFF__0.nand2_2.IN1 VDIV 2.43e-19
C151 DFF__0.nand2_5.OUT DFF__0.inv_0.OUT 1.02e-21
C152 VREF DFF__1.nand2_1.IN1 1.13e-20
C153 DFF__1.nand2_2.IN1 a_1327_4537# 9.39e-21
C154 DFF__0.nand2_3.OUT DFF__0.QB 0.0138f
C155 DFF__0.nand2_2.IN1 DFF__0.nand2_1.IN1 0.00714f
C156 buffer_mag_0.OUT a_444_2859# 8.75e-20
C157 DFF__1.inv_0.OUT a_2563_4471# 0.00372f
C158 DFF__1.nand2_2.IN1 DFF__0.nand2_5.OUT 4.96e-19
C159 buffer_loading_mag_1.IN DFF__0.QB 0.62f
C160 buffer_mag_0.OUT DFF__1.nand2_3.OUT 0.889f
C161 DFF__0.nand2_5.OUT a_3456_1786# 0.00454f
C162 DFF__1.nand2_5.OUT VDD 0.802f
C163 DFF__0.CLK VDD 1f
C164 DFF__1.nand2_5.OUT nand2_0.IN1 0.0678f
C165 DFF__1.QB DFF__1.nand2_1.IN1 0.273f
C166 DFF__1.nand2_1.IN1 DFF__1.CLK 0.114f
C167 buffer_mag_0.OUT a_1327_4537# 0.00348f
C168 DFF__0.nand2_5.OUT a_445_2019# 0.00432f
C169 buffer_mag_0.OUT a_2559_3092# 0.00168f
C170 buffer_mag_0.IN a_4478_3188# 0.0158f
C171 DFF__0.nand2_5.OUT DFF__0.nand2_2.IN2 0.0065f
C172 a_444_2859# VDD 0.00503f
C173 DFF__1.nand2_2.OUT DFF__1.nand2_2.IN2 0.159f
C174 buffer_mag_0.OUT DFF__0.nand2_5.OUT 0.389f
C175 DFF__0.nand2_2.IN1 DFF__0.nand2_3.OUT 0.0185f
C176 DFF__0.inv_0.OUT DFF__0.nand2_2.IN2 0.155f
C177 buffer_mag_0.OUT DFF__0.inv_0.OUT 0.00685f
C178 buffer_mag_0.IN buffer_mag_0.gf_inv_mag_1.IN 0.393f
C179 DFF__1.nand2_3.OUT VDD 0.887f
C180 a_3455_3092# VDD 3.15e-19
C181 DFF__1.inv_0.OUT DFF__1.nand2_2.IN2 0.155f
C182 a_3460_289# DFF__0.QB 0.00619f
C183 DFF__1.nand2_1.IN1 a_2563_4471# 0.00384f
C184 a_611_348# DFF__0.CLK 1.27e-19
C185 DFF__1.nand2_3.OUT nand2_0.IN1 2.23e-19
C186 a_1328_341# DFF__0.nand2_2.IN1 9.39e-21
C187 a_3455_3092# nand2_0.IN1 0.00351f
C188 a_1327_4537# VDD 3.56e-19
C189 DFF__1.nand2_2.IN1 buffer_mag_0.OUT 0.0963f
C190 a_2559_3092# VDD 3.14e-19
C191 a_1330_2902# DFF__1.nand2_1.IN1 0.069f
C192 DFF__1.nand2_3.OUT a_3459_4589# 9.07e-21
C193 DFF__0.nand2_5.OUT VDD 0.803f
C194 DFF__0.inv_0.OUT VDD 0.346f
C195 a_445_2019# DFF__0.nand2_2.IN2 1.16e-20
C196 a_6234_2632# VDD 3.26e-19
C197 buffer_mag_0.OUT a_445_2019# 8.75e-20
C198 buffer_mag_0.OUT DFF__0.nand2_2.IN2 0.0259f
C199 a_6234_2632# nand2_0.IN1 0.00348f
C200 a_4617_1139# VDD 1.21f
C201 buffer_loading_mag_1.IN buffer_mag_0.gf_inv_mag_1.IN 0.0224f
C202 DFF__1.nand2_2.IN1 VDD 0.942f
C203 DFF__1.nand2_1.IN1 DFF__1.nand2_2.IN2 0.459f
C204 buffer_mag_0.IN PU 5.63e-19
C205 a_4617_1139# nand2_0.IN1 5.62e-19
C206 a_611_348# DFF__0.nand2_5.OUT 1.99e-20
C207 a_3456_1786# VDD 4.2e-19
C208 DFF__1.nand2_5.OUT DFF__0.QB 1.82e-20
C209 DFF__0.nand2_5.OUT a_2560_1786# 0.0703f
C210 a_445_2019# VDD 0.00503f
C211 DFF__1.nand2_5.OUT a_610_4530# 1.99e-20
C212 DFF__0.nand2_2.IN2 VDD 0.71f
C213 buffer_mag_0.OUT VDD 1.9f
C214 DFF__1.inv_0.OUT DFF__1.nand2_1.IN1 0.0551f
C215 buffer_mag_0.OUT nand2_0.IN1 0.375f
C216 DFF__0.nand2_1.IN1 VDIV 4.13e-21
C217 DFF__0.nand2_2.OUT DFF__0.nand2_3.OUT 0.106f
C218 buffer_loading_mag_1.IN PU 5.72e-19
C219 a_2564_407# DFF__0.inv_0.OUT 0.00372f
C220 a_1331_1976# DFF__0.nand2_1.IN1 0.069f
C221 a_611_348# DFF__0.nand2_2.IN2 0.0175f
C222 a_610_4530# DFF__1.nand2_3.OUT 1.26e-20
C223 DFF__0.nand2_2.IN1 DFF__1.nand2_5.OUT 4.94e-19
C224 DFF__0.nand2_2.OUT a_1328_341# 0.00364f
C225 DFF__0.nand2_1.IN1 DFF__1.nand2_1.IN1 8.9e-19
C226 DFF__0.nand2_2.IN1 DFF__0.CLK 0.145f
C227 DFF__0.nand2_5.OUT DFF__0.QB 0.581f
C228 DFF__1.QB DFF__1.nand2_5.OUT 0.581f
C229 buffer_mag_0.OUT a_2560_1786# 0.00168f
C230 nand2_0.IN1 VDD 1.99f
C231 DFF__1.nand2_5.OUT DFF__1.CLK 0.115f
C232 DFF__0.QB DFF__0.inv_0.OUT 0.00316f
C233 DFF__0.CLK DFF__1.CLK 0.00128f
C234 a_3459_4589# VDD 3.15e-19
C235 DFF__0.nand2_1.IN1 DFF__0.nand2_3.OUT 0.39f
C236 a_3459_4589# nand2_0.IN1 0.069f
C237 a_444_2859# DFF__1.CLK 9.59e-19
C238 a_611_348# VDD 3.14e-19
C239 a_2564_407# DFF__0.nand2_2.IN2 0.0769f
C240 DFF__1.nand2_5.OUT buffer_mag_0.gf_inv_mag_1.IN 1.23e-19
C241 DFF__0.QB a_3456_1786# 0.0692f
C242 DFF__1.QB DFF__1.nand2_3.OUT 0.0138f
C243 DFF__0.nand2_1.IN1 buffer_loading_mag_1.IN 0.0119f
C244 DFF__1.QB a_3455_3092# 0.0692f
C245 a_2560_1786# VDD 3.14e-19
C246 DFF__1.nand2_2.IN1 a_610_4530# 0.00348f
C247 DFF__1.nand2_5.OUT a_1330_2902# 3.83e-19
C248 DFF__1.nand2_2.IN1 VREF 3.73e-19
C249 DFF__0.nand2_2.IN1 DFF__0.nand2_5.OUT 0.492f
C250 buffer_mag_0.IN buffer_loading_mag_1.IN 0.137f
C251 DFF__0.QB DFF__0.nand2_2.IN2 0.147f
C252 DFF__0.nand2_2.IN1 DFF__0.inv_0.OUT 4.23e-20
C253 buffer_mag_0.OUT DFF__0.QB 9.68e-20
C254 DFF__1.QB DFF__0.nand2_5.OUT 1.73e-20
C255 DFF__0.nand2_5.OUT DFF__1.CLK 6.57e-19
C256 DFF__1.nand2_3.OUT a_2563_4471# 2.09e-19
C257 a_2564_407# VDD 3.22e-19
C258 DFF__0.nand2_2.IN1 DFF__1.nand2_2.IN1 0.00935f
C259 DFF__1.nand2_5.OUT DFF__1.nand2_2.IN2 0.0065f
C260 a_3460_289# DFF__0.nand2_1.IN1 1.63e-20
C261 DFF__0.nand2_3.OUT buffer_loading_mag_1.IN 2.23e-19
C262 a_1328_341# DFF__0.nand2_3.OUT 0.069f
C263 DFF__1.nand2_2.IN1 DFF__1.CLK 0.146f
C264 DFF__0.nand2_5.OUT buffer_mag_0.gf_inv_mag_1.IN 3.54e-19
C265 DFF__0.QB VDD 1.11f
C266 DFF__0.nand2_2.IN1 a_445_2019# 0.069f
C267 a_444_2859# DFF__1.nand2_2.IN2 1.16e-20
C268 buffer_mag_0.IN PD 6.68e-19
C269 DFF__1.nand2_2.OUT DFF__1.nand2_5.OUT 1.33e-19
C270 DFF__0.nand2_2.OUT DFF__0.CLK 0.00375f
C271 DFF__0.nand2_2.IN1 DFF__0.nand2_2.IN2 0.0753f
.ends

