* NGSPICE file created from Current_Mirror_Top_flat.ext - technology: gf180mcuC

.subckt pex_Current_Mirror_Top VDD ITAIL ITAIL_SRC ITAIL_SINK  VSS
X0 VDD G_source_up.t6 G_source_up.t7 VDD.t50 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 VDD G1_2.t60 SD1_1.t11 VDD.t67 pfet_03v3 ad=0.176p pd=1.68u as=0.104p ps=0.92u w=0.4u l=0.5u
X2 VSS G2_1.t37 G2_1.t38 VSS.t44 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X3 ITAIL ITAIL.t38 G2_1.t7 VSS.t40 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X4 ITAIL_SRC G_source_dn.t24 A1.t14 VDD.t20 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X5 G_source_dn G_source_dn.t22 G_source_up.t21 VDD.t80 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X6 G_sink_up G1_1.t60 SD1_1.t12 VDD.t3 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X7 VDD G1_2.t45 G1_2.t46 VDD.t98 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X8 VSS G_sink_dn.t24 SD0_1.t15 VSS.t32 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X9 VDD G1_2.t43 G1_2.t44 VDD.t95 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X10 SD0_1 G_sink_dn.t25 VSS.t134 VSS.t15 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X11 SD2_1 G2_1.t60 VSS.t129 VSS.t60 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X12 VSS G2_1.t35 G2_1.t36 VSS.t54 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X13 G2_1 ITAIL.t36 ITAIL.t37 VSS.t43 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X14 VDD G1_2.t41 G1_2.t42 VDD.t67 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X15 G2_1 ITAIL.t34 ITAIL.t35 VSS.t46 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X16 G1_2 G1_2.t39 VDD.t109 VDD.t55 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X17 ITAIL ITAIL.t32 G2_1.t12 VSS.t64 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X18 SD2_1 G2_1.t61 VSS.t126 VSS.t18 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X19 SD0_1 G_sink_dn.t26 VSS.t68 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X20 G_sink_dn G_sink_dn.t22 VSS.t49 VSS.t48 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X21 G1_1 G1_1.t38 G1_2.t53 VDD.t3 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X22 G1_2 G1_2.t37 VDD.t14 VDD.t13 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X23 A2 G_sink_up.t26 ITAIL_SINK.t5 VSS.t3 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X24 VDD G1_2.t35 G1_2.t36 VDD.t10 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X25 ITAIL ITAIL.t30 G2_1.t8 VSS.t45 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X26 G1_2 G1_1.t36 G1_1.t37 VDD.t88 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X27 ITAIL_SINK G_sink_up.t27 A2.t6 VSS.t8 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X28 G_sink_dn G_sink_up.t20 G_sink_up.t21 VSS.t58 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X29 VSS G2_1.t62 SD2_1.t37 VSS.t16 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X30 ITAIL_SINK G_sink_up.t28 A2.t5 VSS.t37 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X31 G_sink_up G1_1.t62 SD1_1.t13 VDD.t7 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X32 VSS G2_1.t63 SD2_1.t36 VSS.t40 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X33 ITAIL_SRC G_source_dn.t26 A1.t13 VDD.t45 pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X34 VSS G_sink_dn.t28 SD0_1.t12 VSS.t4 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X35 VSS G2_1.t33 G2_1.t34 VSS.t41 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X36 SD2_1 G2_1.t64 VSS.t119 VSS.t61 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X37 A1 G_source_up.t24 VDD.t49 VDD.t48 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X38 VSS G2_1.t31 G2_1.t32 VSS.t62 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X39 G_source_dn G_source_dn.t20 G_source_up.t20 VDD.t79 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X40 G_sink_up G1_1.t63 SD1_1.t18 VDD.t6 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X41 VSS G2_1.t65 SD2_1.t34 VSS.t44 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X42 G_sink_up G_sink_up.t10 G_sink_dn.t6 VSS.t2 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X43 G2_1 ITAIL.t28 ITAIL.t29 VSS.t61 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X44 G1_1 G1_1.t34 G1_2.t50 VDD.t83 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X45 VSS G_sink_dn.t20 G_sink_dn.t21 VSS.t34 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X46 VSS G_sink_dn.t29 SD0_1.t11 VSS.t47 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X47 SD1_1 G1_2.t63 VDD.t71 VDD.t70 pfet_03v3 ad=0.104p pd=0.92u as=0.176p ps=1.68u w=0.4u l=0.5u
X48 G1_1 ITAIL.t43 SD2_1.t19 VSS.t24 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X49 SD2_1 G2_1.t66 VSS.t114 VSS.t0 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X50 G1_1 G1_1.t32 G1_2.t1 VDD.t7 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X51 VSS G2_1.t67 SD2_1.t32 VSS.t41 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X52 VDD G_source_up.t25 A1.t6 VDD.t45 pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X53 SD2_1 ITAIL G1_1.t59 VSS.t46 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X54 G2_1 ITAIL.t26 ITAIL.t27 VSS.t22 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X55 G2_1 G2_1.t17 VSS.t111 VSS.t65 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X56 A1 G_source_dn.t28 ITAIL_SRC.t5 VDD.t48 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X57 G_source_up G_source_up.t14 VDD.t41 VDD.t40 pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X58 G_source_up G_source_up.t8 VDD.t44 VDD.t43 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X59 SD1_1 G1_2.t64 VDD.t59 VDD.t58 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X60 G_sink_dn G_sink_up.t18 G_sink_up.t19 VSS.t1 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X61 G1_1 G1_1.t30 G1_2.t0 VDD.t6 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X62 VSS G2_1.t29 G2_1.t30 VSS.t23 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X63 SD0_1 G_sink_up.t30 G_source_dn.t4 VSS.t55 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X64 G1_2 G1_2.t33 VDD.t103 VDD.t70 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X65 G2_1 G2_1.t41 VSS.t108 VSS.t0 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X66 G1_1 ITAIL SD2_1.t17 VSS.t45 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X67 G1_2 G1_1.t28 G1_1.t29 VDD.t86 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X68 VSS G2_1.t27 G2_1.t28 VSS.t24 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X69 G_source_up G_source_dn.t18 G_source_dn.t19 VDD.t64 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X70 G2_1 ITAIL.t24 ITAIL.t25 VSS.t17 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X71 G_sink_dn G_sink_up.t16 G_sink_up.t17 VSS.t50 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X72 VSS G_sink_dn.t30 SD0_1.t10 VSS.t29 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X73 G1_2 G1_2.t31 VDD.t102 VDD.t58 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X74 A2 G_sink_dn.t31 VSS.t66 VSS.t3 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X75 G1_1 ITAIL.t44 SD2_1.t16 VSS.t64 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X76 A2 G_sink_dn.t32 VSS.t53 VSS.t52 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X77 ITAIL ITAIL.t22 G2_1.t1 VSS.t16 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X78 G1_1 G1_1.t26 G1_2.t57 VDD.t98 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X79 VSS G_sink_dn.t33 A2.t13 VSS.t19 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X80 G_sink_up G1_1.t68 SD1_1.t19 VDD.t78 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X81 VSS G_sink_dn.t34 A2.t12 VSS.t37 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X82 G1_1 G1_1.t24 G1_2.t56 VDD.t95 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X83 G_sink_up G_sink_up.t22 G_sink_dn.t3 VSS.t12 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X84 G2_1 G2_1.t47 VSS.t105 VSS.t18 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X85 VDD G_source_up.t28 A1.t5 VDD.t8 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X86 G_source_dn G_sink_up.t32 SD0_1.t6 VSS.t32 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X87 A2 G_sink_up.t33 ITAIL_SINK.t4 VSS.t33 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X88 VDD G1_2.t67 SD1_1.t8 VDD.t0 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X89 G1_1 ITAIL.t46 SD2_1.t15 VSS.t62 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X90 SD2_1 G2_1.t71 VSS.t104 VSS.t43 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X91 SD0_1 G_sink_up.t34 G_source_dn.t1 VSS.t15 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X92 SD2_1 ITAIL G1_1.t58 VSS.t18 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X93 G1_1 G1_1.t22 G1_2.t48 VDD.t67 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X94 A1 G_source_dn.t29 ITAIL_SRC.t4 VDD.t34 pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X95 SD1_1 G1_2.t68 VDD.t63 VDD.t62 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X96 VDD G_source_up.t4 G_source_up.t5 VDD.t36 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X97 G2_1 G2_1.t49 VSS.t103 VSS.t60 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X98 VSS G2_1.t25 G2_1.t26 VSS.t40 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X99 VDD G1_2.t29 G1_2.t30 VDD.t3 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X100 SD1_1 G1_1.t71 G_sink_up.t5 VDD.t81 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X101 G1_1 G1_1.t20 G1_2.t47 VDD.t78 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X102 G_sink_dn G_sink_up.t14 G_sink_up.t15 VSS.t48 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X103 SD2_1 G2_1.t73 VSS.t100 VSS.t22 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X104 ITAIL_SRC G_source_dn.t30 A1.t12 VDD.t8 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X105 SD1_1 G1_1.t73 G_sink_up.t4 VDD.t53 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X106 VDD G1_2.t27 G1_2.t28 VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X107 G1_1 ITAIL SD2_1.t13 VSS.t16 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X108 G2_1 ITAIL.t20 ITAIL.t21 VSS.t42 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X109 SD0_1 G_sink_dn.t35 VSS.t67 VSS.t63 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X110 G1_1 ITAIL SD2_1.t12 VSS.t40 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X111 G_source_up G_source_dn.t16 G_source_dn.t17 VDD.t101 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X112 A1 G_source_up.t29 VDD.t35 VDD.t34 pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X113 G2_1 G2_1.t43 VSS.t99 VSS.t43 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X114 G_source_up G_source_dn.t14 G_source_dn.t15 VDD.t104 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X115 G_sink_dn G_sink_dn.t18 VSS.t137 VSS.t58 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X116 SD1_1 G1_1.t74 G_sink_up.t3 VDD.t54 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X117 G1_2 G1_2.t25 VDD.t74 VDD.t62 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X118 ITAIL ITAIL.t18 G2_1.t10 VSS.t54 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X119 G1_2 G1_1.t18 G1_1.t19 VDD.t81 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X120 G2_1 G2_1.t51 VSS.t98 VSS.t46 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X121 G1_1 ITAIL SD2_1.t11 VSS.t44 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X122 G1_2 G1_1.t16 G1_1.t17 VDD.t53 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X123 ITAIL ITAIL.t16 G2_1.t9 VSS.t44 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X124 VSS G2_1.t76 SD2_1.t29 VSS.t24 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X125 G_source_dn G_source_dn.t12 G_source_up.t19 VDD.t77 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X126 G_source_dn G_sink_up.t35 SD0_1.t4 VSS.t47 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X127 VSS G2_1.t23 G2_1.t24 VSS.t45 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X128 G1_1 ITAIL.t49 SD2_1.t10 VSS.t54 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X129 VDD G1_2.t23 G1_2.t24 VDD.t7 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X130 G1_2 G1_1.t14 G1_1.t15 VDD.t54 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X131 A2 G_sink_up.t36 ITAIL_SINK.t3 VSS.t52 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X132 VSS G2_1.t77 SD2_1.t28 VSS.t23 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X133 ITAIL_SINK G_sink_up.t37 A2.t2 VSS.t19 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X134 VSS G_sink_dn.t16 G_sink_dn.t17 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X135 ITAIL_SINK G_sink_up.t38 A2.t1 VSS.t69 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X136 ITAIL ITAIL.t14 G2_1.t15 VSS.t41 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X137 VDD G1_2.t21 G1_2.t22 VDD.t6 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X138 A2 G_sink_dn.t37 VSS.t57 VSS.t33 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X139 ITAIL ITAIL.t12 G2_1.t14 VSS.t62 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X140 SD2_1 G2_1.t78 VSS.t91 VSS.t42 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X141 A2 G_sink_dn.t38 VSS.t26 VSS.t25 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X142 G1_2 G1_1.t12 G1_1.t13 VDD.t70 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X143 VSS G2_1.t21 G2_1.t22 VSS.t64 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X144 SD0_1 G_sink_dn.t39 VSS.t56 VSS.t55 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X145 SD1_1 G1_1.t75 G_sink_up.t2 VDD.t55 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X146 SD2_1 ITAIL.t52 G1_1.t57 VSS.t65 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X147 SD2_1 ITAIL.t53 G1_1.t56 VSS.t17 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X148 G_source_up G_source_dn.t10 G_source_dn.t11 VDD.t57 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X149 SD1_1 G1_1.t76 G_sink_up.t1 VDD.t13 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X150 G2_1 G2_1.t55 VSS.t88 VSS.t22 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X151 VSS G2_1.t80 SD2_1.t26 VSS.t64 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X152 ITAIL_SRC G_source_dn.t32 A1.t11 VDD.t9 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X153 G2_1 ITAIL.t10 ITAIL.t11 VSS.t65 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X154 G1_2 G1_1.t10 G1_1.t11 VDD.t58 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X155 G_sink_dn G_sink_dn.t14 VSS.t51 VSS.t50 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X156 G_sink_up G1_1.t77 SD1_1.t17 VDD.t10 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X157 SD1_1 G1_2.t70 VDD.t89 VDD.t88 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X158 SD2_1 ITAIL.t54 G1_1.t55 VSS.t60 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X159 G_source_up G_source_up.t12 VDD.t33 VDD.t32 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X160 SD0_1 G_sink_up.t39 G_source_dn.t0 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X161 G1_2 G1_1.t8 G1_1.t9 VDD.t55 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X162 VSS G2_1.t81 SD2_1.t25 VSS.t62 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X163 G_source_dn G_source_dn.t8 G_source_up.t16 VDD.t56 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X164 SD2_1 ITAIL G1_1.t54 VSS.t43 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X165 G_source_up G_source_up.t10 VDD.t31 VDD.t30 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X166 G2_1 ITAIL.t8 ITAIL.t9 VSS.t0 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X167 G2_1 G2_1.t45 VSS.t83 VSS.t61 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X168 VSS G_sink_dn.t12 G_sink_dn.t13 VSS.t12 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X169 G1_2 G1_1.t6 G1_1.t7 VDD.t13 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X170 ITAIL ITAIL.t6 G2_1.t6 VSS.t24 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X171 VDD G_source_up.t32 A1.t3 VDD.t9 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X172 VDD G1_2.t71 SD1_1.t5 VDD.t83 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X173 G1_1 G1_1.t4 G1_2.t6 VDD.t10 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X174 G1_2 G1_2.t19 VDD.t112 VDD.t88 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X175 G_source_dn G_sink_up.t40 SD0_1.t2 VSS.t4 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X176 SD2_1 ITAIL G1_1.t53 VSS.t22 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X177 VDD G1_2.t17 G1_2.t18 VDD.t78 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X178 VSS G2_1.t19 G2_1.t20 VSS.t16 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X179 VDD G_source_up.t2 G_source_up.t3 VDD.t25 pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X180 G1_1 G1_1.t2 G1_2.t5 VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X181 ITAIL ITAIL.t4 G2_1.t5 VSS.t23 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X182 VSS G_sink_dn.t10 G_sink_dn.t11 VSS.t2 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X183 VSS G_sink_dn.t41 A2.t9 VSS.t69 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X184 G_sink_up G_sink_up.t12 G_sink_dn.t1 VSS.t34 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X185 SD2_1 ITAIL.t57 G1_1.t52 VSS.t61 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X186 SD0_1 G_sink_up.t42 G_source_dn.t6 VSS.t63 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X187 VDD G1_2.t15 G1_2.t16 VDD.t83 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X188 G1_2 G1_1.t0 G1_1.t1 VDD.t62 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X189 A2 G_sink_up.t43 ITAIL_SINK.t2 VSS.t25 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X190 G1_2 G1_2.t13 VDD.t82 VDD.t81 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X191 G2_1 ITAIL.t2 ITAIL.t3 VSS.t60 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X192 G2_1 G2_1.t39 VSS.t74 VSS.t17 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X193 SD2_1 ITAIL.t58 G1_1.t51 VSS.t0 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X194 A1 G_source_dn.t34 ITAIL_SRC.t1 VDD.t18 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X195 SD1_1 G1_2.t74 VDD.t92 VDD.t86 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X196 G1_2 G1_2.t11 VDD.t76 VDD.t53 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X197 G_sink_dn G_sink_dn.t8 VSS.t59 VSS.t1 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X198 G1_1 ITAIL.t59 SD2_1.t2 VSS.t41 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X199 SD2_1 G2_1.t84 VSS.t80 VSS.t46 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X200 VSS G2_1.t85 SD2_1.t23 VSS.t54 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X201 A1 G_source_up.t33 VDD.t24 VDD.t23 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X202 VSS G_sink_dn.t43 A2.t8 VSS.t8 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X203 G2_1 G2_1.t53 VSS.t73 VSS.t42 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X204 G1_1 ITAIL SD2_1.t1 VSS.t23 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X205 VDD G_source_up.t34 A1.t1 VDD.t20 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X206 G1_2 G1_2.t9 VDD.t75 VDD.t54 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X207 VDD G1_2.t77 SD1_1.t3 VDD.t98 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X208 G2_1 ITAIL.t0 ITAIL.t1 VSS.t18 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X209 VDD G1_2.t78 SD1_1.t2 VDD.t95 pfet_03v3 ad=0.104p pd=0.92u as=0.104p ps=0.92u w=0.4u l=0.5u
X210 A1 G_source_up.t35 VDD.t19 VDD.t18 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X211 VDD G_source_up.t0 G_source_up.t1 VDD.t15 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X212 G1_2 G1_2.t7 VDD.t87 VDD.t86 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X213 SD2_1 ITAIL G1_1.t50 VSS.t42 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X214 G_source_dn G_sink_up.t44 SD0_1.t0 VSS.t29 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X215 G_sink_up G_sink_up.t24 G_sink_dn.t0 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X216 VSS G2_1.t87 SD2_1.t22 VSS.t45 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X217 SD2_1 G2_1.t88 VSS.t75 VSS.t65 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X218 A1 G_source_dn.t35 ITAIL_SRC.t0 VDD.t23 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X219 SD2_1 G2_1.t89 VSS.t72 VSS.t17 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
R0 G_source_up.n38 G_source_up.n37 95.8364
R1 G_source_up.n34 G_source_up.t29 84.6824
R2 G_source_up.n36 G_source_up.n35 68.6827
R3 G_source_up.n37 G_source_up.t33 32.5342
R4 G_source_up.n13 G_source_up.n12 27.2758
R5 G_source_up.n21 G_source_up.n20 27.2758
R6 G_source_up.n29 G_source_up.n28 27.2758
R7 G_source_up.n39 G_source_up.n38 20.988
R8 G_source_up.n35 G_source_up.n34 14.325
R9 G_source_up.n34 G_source_up.t32 13.9435
R10 G_source_up.n35 G_source_up.t35 13.9435
R11 G_source_up.n37 G_source_up.t28 13.0675
R12 G_source_up.n38 G_source_up.t24 13.0675
R13 G_source_up.n36 G_source_up.t25 12.6295
R14 G_source_up.n39 G_source_up.t34 11.5326
R15 G_source_up.n6 G_source_up.t2 10.4831
R16 G_source_up.n41 G_source_up.t14 9.08115
R17 G_source_up.n12 G_source_up.t10 7.5925
R18 G_source_up.n13 G_source_up.t6 7.5925
R19 G_source_up.n20 G_source_up.t8 7.5925
R20 G_source_up.n21 G_source_up.t4 7.5925
R21 G_source_up.n28 G_source_up.t12 7.5925
R22 G_source_up.n29 G_source_up.t0 7.5925
R23 G_source_up.n40 G_source_up.n39 7.36467
R24 G_source_up.n40 G_source_up.n36 5.1305
R25 G_source_up.n42 G_source_up.n40 4.28043
R26 G_source_up.n7 G_source_up.n6 4.0005
R27 G_source_up.n11 G_source_up.n10 4.0005
R28 G_source_up.n15 G_source_up.n14 4.0005
R29 G_source_up.n19 G_source_up.n18 4.0005
R30 G_source_up.n23 G_source_up.n22 4.0005
R31 G_source_up.n27 G_source_up.n26 4.0005
R32 G_source_up.n33 G_source_up.n30 4.0005
R33 G_source_up.n49 G_source_up.t16 3.03383
R34 G_source_up.n49 G_source_up.n48 3.03383
R35 G_source_up.n25 G_source_up.t20 3.03383
R36 G_source_up.n25 G_source_up.n24 3.03383
R37 G_source_up.n1 G_source_up.t5 3.03383
R38 G_source_up.n1 G_source_up.n0 3.03383
R39 G_source_up.n17 G_source_up.t21 3.03383
R40 G_source_up.n17 G_source_up.n16 3.03383
R41 G_source_up.n3 G_source_up.t7 3.03383
R42 G_source_up.n3 G_source_up.n2 3.03383
R43 G_source_up.n9 G_source_up.t19 3.03383
R44 G_source_up.n9 G_source_up.n8 3.03383
R45 G_source_up.n5 G_source_up.t3 3.03383
R46 G_source_up.n5 G_source_up.n4 3.03383
R47 G_source_up.n32 G_source_up.t1 3.03383
R48 G_source_up.n32 G_source_up.n31 3.03383
R49 G_source_up.n26 G_source_up.n25 2.84924
R50 G_source_up.n23 G_source_up.n1 2.84924
R51 G_source_up.n18 G_source_up.n17 2.84924
R52 G_source_up.n15 G_source_up.n3 2.84924
R53 G_source_up.n10 G_source_up.n9 2.84924
R54 G_source_up.n33 G_source_up.n32 2.84924
R55 G_source_up.n7 G_source_up.n5 2.84872
R56 G_source_up.n45 G_source_up.n44 2.66717
R57 G_source_up.n50 G_source_up.n49 2.6005
R58 G_source_up.n12 G_source_up.n11 2.59881
R59 G_source_up.n14 G_source_up.n13 2.59881
R60 G_source_up.n20 G_source_up.n19 2.59881
R61 G_source_up.n22 G_source_up.n21 2.59881
R62 G_source_up.n28 G_source_up.n27 2.59881
R63 G_source_up.n30 G_source_up.n29 2.59881
R64 G_source_up.n42 G_source_up.n41 2.44013
R65 G_source_up.n44 G_source_up.n43 2.28948
R66 G_source_up.n47 G_source_up.n33 0.742375
R67 G_source_up.n10 G_source_up.n7 0.728327
R68 G_source_up.n26 G_source_up.n23 0.724527
R69 G_source_up.n18 G_source_up.n15 0.720586
R70 G_source_up.n50 G_source_up.n47 0.213761
R71 G_source_up G_source_up.n50 0.203898
R72 G_source_up.n46 G_source_up.n45 0.0355526
R73 G_source_up.n47 G_source_up.n46 0.0222895
R74 G_source_up.n45 G_source_up.n42 0.00144737
R75 VDD.n151 VDD.t43 151.695
R76 VDD.n151 VDD.t36 148.749
R77 VDD.n136 VDD.t25 122.648
R78 VDD.n203 VDD.t40 122.444
R79 VDD.n148 VDD.t80 113.403
R80 VDD.n153 VDD.t57 110.457
R81 VDD.n164 VDD.t56 81.002
R82 VDD.n137 VDD.t64 78.0565
R83 VDD.n179 VDD.t45 76.1029
R84 VDD.n146 VDD.t104 75.111
R85 VDD.n155 VDD.t79 72.1654
R86 VDD.n190 VDD.t34 64.0119
R87 VDD.n76 VDD.t78 56.5849
R88 VDD.n60 VDD.t54 54.5272
R89 VDD.n60 VDD.t3 50.412
R90 VDD.n76 VDD.t86 48.3544
R91 VDD.n180 VDD.t23 46.9422
R92 VDD.n189 VDD.t20 45.5197
R93 VDD.n91 VDD.t10 45.268
R94 VDD.n75 VDD.t53 43.2104
R95 VDD.n162 VDD.t101 42.7104
R96 VDD.n59 VDD.t67 41.1528
R97 VDD.n139 VDD.t77 39.7649
R98 VDD.n61 VDD.t58 37.0375
R99 VDD.n144 VDD.t50 36.8194
R100 VDD.n81 VDD.t0 34.9799
R101 VDD.n157 VDD.t32 33.8738
R102 VDD.n93 VDD.t70 32.4079
R103 VDD.n90 VDD.t81 31.8935
R104 VDD.n74 VDD.t95 29.8359
R105 VDD.n183 VDD.t8 28.45
R106 VDD.n186 VDD.t48 27.0275
R107 VDD.n66 VDD.t83 23.663
R108 VDD.n82 VDD.t55 21.6054
R109 VDD.n89 VDD.t98 18.519
R110 VDD.n69 VDD.t88 16.4614
R111 VDD.n67 VDD.t13 10.2886
R112 VDD.n184 VDD.t18 9.95783
R113 VDD.n185 VDD.t9 8.53535
R114 VDD.n83 VDD.t7 8.23095
R115 VDD.n108 VDD.t71 7.62593
R116 VDD.n134 VDD.n7 7.1505
R117 VDD.n57 VDD.n56 6.54575
R118 VDD.n102 VDD.n101 6.50606
R119 VDD.n191 VDD.n190 6.40831
R120 VDD.n110 VDD.n91 6.3005
R121 VDD.n111 VDD.n90 6.3005
R122 VDD.n112 VDD.n89 6.3005
R123 VDD.n114 VDD.n84 6.3005
R124 VDD.n115 VDD.n83 6.3005
R125 VDD.n116 VDD.n82 6.3005
R126 VDD.n117 VDD.n81 6.3005
R127 VDD.n119 VDD.n76 6.3005
R128 VDD.n120 VDD.n75 6.3005
R129 VDD.n121 VDD.n74 6.3005
R130 VDD.n123 VDD.n69 6.3005
R131 VDD.n124 VDD.n68 6.3005
R132 VDD.n125 VDD.n67 6.3005
R133 VDD.n126 VDD.n66 6.3005
R134 VDD.n128 VDD.n61 6.3005
R135 VDD.n129 VDD.n60 6.3005
R136 VDD.n130 VDD.n59 6.3005
R137 VDD.n12 VDD.n10 6.3005
R138 VDD.n96 VDD.n94 6.3005
R139 VDD.n12 VDD.n9 6.3005
R140 VDD.n191 VDD.n189 6.3005
R141 VDD.n193 VDD.n186 6.3005
R142 VDD.n194 VDD.n185 6.3005
R143 VDD.n195 VDD.n184 6.3005
R144 VDD.n196 VDD.n183 6.3005
R145 VDD.n198 VDD.n180 6.3005
R146 VDD.n199 VDD.n179 6.3005
R147 VDD.n165 VDD.n164 6.3005
R148 VDD.n163 VDD.n162 6.3005
R149 VDD.n161 VDD.n160 6.3005
R150 VDD.n158 VDD.n157 6.3005
R151 VDD.n156 VDD.n155 6.3005
R152 VDD.n154 VDD.n153 6.3005
R153 VDD.n152 VDD.n151 6.3005
R154 VDD.n149 VDD.n148 6.3005
R155 VDD.n147 VDD.n146 6.3005
R156 VDD.n145 VDD.n144 6.3005
R157 VDD.n142 VDD.n141 6.3005
R158 VDD.n140 VDD.n139 6.3005
R159 VDD.n138 VDD.n137 6.3005
R160 VDD.n201 VDD.t41 6.21492
R161 VDD.n135 VDD.n6 6.21492
R162 VDD.n169 VDD.t35 6.18924
R163 VDD.n177 VDD.n166 6.18362
R164 VDD.n84 VDD.t62 5.14453
R165 VDD.n94 VDD.n93 5.14453
R166 VDD.n108 VDD.t103 5.00941
R167 VDD.n132 VDD.n58 5.00941
R168 VDD.n63 VDD.t59 4.5505
R169 VDD.n63 VDD.n62 4.5505
R170 VDD.n71 VDD.t89 4.5505
R171 VDD.n71 VDD.n70 4.5505
R172 VDD.n78 VDD.t92 4.5505
R173 VDD.n78 VDD.n77 4.5505
R174 VDD.n86 VDD.t63 4.5505
R175 VDD.n86 VDD.n85 4.5505
R176 VDD.n12 VDD.n11 4.5005
R177 VDD.n160 VDD.t15 4.41876
R178 VDD.n16 VDD.n15 3.60132
R179 VDD.n53 VDD.n23 3.18941
R180 VDD.n48 VDD.n25 3.18941
R181 VDD.n43 VDD.n27 3.18941
R182 VDD.n39 VDD.n29 3.18941
R183 VDD.n34 VDD.n31 3.18941
R184 VDD.n127 VDD.n65 3.18941
R185 VDD.n122 VDD.n73 3.18941
R186 VDD.n118 VDD.n80 3.18941
R187 VDD.n113 VDD.n88 3.18941
R188 VDD.n159 VDD.n1 3.18159
R189 VDD.n150 VDD.n3 3.18159
R190 VDD.n143 VDD.n5 3.18159
R191 VDD.n107 VDD.n106 3.15175
R192 VDD.n18 VDD.n17 3.15175
R193 VDD.n17 VDD.n16 3.151
R194 VDD.n106 VDD.n105 3.151
R195 VDD.n16 VDD.n14 3.151
R196 VDD.n105 VDD.n104 3.151
R197 VDD.n204 VDD.n203 3.1505
R198 VDD.n173 VDD.n168 3.15028
R199 VDD.n197 VDD.n182 3.11115
R200 VDD.n192 VDD.n188 3.11115
R201 VDD.n68 VDD.t6 3.08692
R202 VDD.n127 VDD.n63 3.07593
R203 VDD.n122 VDD.n71 3.07593
R204 VDD.n118 VDD.n78 3.07593
R205 VDD.n113 VDD.n86 3.07593
R206 VDD.n182 VDD.t24 3.03383
R207 VDD.n182 VDD.n181 3.03383
R208 VDD.n188 VDD.t49 3.03383
R209 VDD.n188 VDD.n187 3.03383
R210 VDD.n168 VDD.t19 3.03383
R211 VDD.n168 VDD.n167 3.03383
R212 VDD.n1 VDD.t33 3.03383
R213 VDD.n1 VDD.n0 3.03383
R214 VDD.n3 VDD.t44 3.03383
R215 VDD.n3 VDD.n2 3.03383
R216 VDD.n5 VDD.t31 3.03383
R217 VDD.n5 VDD.n4 3.03383
R218 VDD.n18 VDD.n13 2.76626
R219 VDD.n20 VDD.n19 2.75233
R220 VDD.n102 VDD.n96 2.62983
R221 VDD.n100 VDD.n98 2.62936
R222 VDD.n55 VDD.n21 2.62088
R223 VDD.n135 VDD.n134 2.24061
R224 VDD.n105 VDD.n103 2.05811
R225 VDD.n23 VDD.t75 1.8205
R226 VDD.n23 VDD.n22 1.8205
R227 VDD.n25 VDD.t14 1.8205
R228 VDD.n25 VDD.n24 1.8205
R229 VDD.n27 VDD.t76 1.8205
R230 VDD.n27 VDD.n26 1.8205
R231 VDD.n29 VDD.t109 1.8205
R232 VDD.n29 VDD.n28 1.8205
R233 VDD.n31 VDD.t82 1.8205
R234 VDD.n31 VDD.n30 1.8205
R235 VDD.n65 VDD.t102 1.8205
R236 VDD.n65 VDD.n64 1.8205
R237 VDD.n73 VDD.t112 1.8205
R238 VDD.n73 VDD.n72 1.8205
R239 VDD.n80 VDD.t87 1.8205
R240 VDD.n80 VDD.n79 1.8205
R241 VDD.n88 VDD.t74 1.8205
R242 VDD.n88 VDD.n87 1.8205
R243 VDD.n96 VDD.n92 1.77932
R244 VDD.n96 VDD.n95 1.61584
R245 VDD.n98 VDD.n97 1.48285
R246 VDD.n141 VDD.t30 1.47325
R247 VDD.n9 VDD.n8 1.02931
R248 VDD.n13 VDD.n12 0.78178
R249 VDD.n200 VDD.n178 0.449005
R250 VDD.n200 VDD.n199 0.350061
R251 VDD.n134 VDD.n133 0.19404
R252 VDD.n199 VDD.n198 0.115344
R253 VDD.n201 VDD.n200 0.113938
R254 VDD.n177 VDD.n176 0.113
R255 VDD.n203 VDD.n202 0.111676
R256 VDD.n52 VDD.n51 0.108313
R257 VDD.n51 VDD.n50 0.108313
R258 VDD.n50 VDD.n49 0.108313
R259 VDD.n47 VDD.n46 0.108313
R260 VDD.n46 VDD.n45 0.108313
R261 VDD.n45 VDD.n44 0.108313
R262 VDD.n42 VDD.n41 0.108313
R263 VDD.n41 VDD.n40 0.108313
R264 VDD.n38 VDD.n37 0.108313
R265 VDD.n37 VDD.n36 0.108313
R266 VDD.n36 VDD.n35 0.108313
R267 VDD.n130 VDD.n129 0.108313
R268 VDD.n129 VDD.n128 0.108313
R269 VDD.n126 VDD.n125 0.108313
R270 VDD.n125 VDD.n124 0.108313
R271 VDD.n124 VDD.n123 0.108313
R272 VDD.n121 VDD.n120 0.108313
R273 VDD.n120 VDD.n119 0.108313
R274 VDD.n117 VDD.n116 0.108313
R275 VDD.n116 VDD.n115 0.108313
R276 VDD.n115 VDD.n114 0.108313
R277 VDD.n112 VDD.n111 0.108313
R278 VDD.n111 VDD.n110 0.108313
R279 VDD.n196 VDD.n195 0.108313
R280 VDD.n195 VDD.n194 0.108313
R281 VDD.n194 VDD.n193 0.108313
R282 VDD.n176 VDD.n175 0.108313
R283 VDD.n175 VDD.n174 0.108313
R284 VDD.n172 VDD.n171 0.108313
R285 VDD.n171 VDD.n170 0.108313
R286 VDD.n170 VDD.n169 0.108313
R287 VDD.n138 VDD.n136 0.108313
R288 VDD.n140 VDD.n138 0.108313
R289 VDD.n142 VDD.n140 0.108313
R290 VDD.n147 VDD.n145 0.108313
R291 VDD.n149 VDD.n147 0.108313
R292 VDD.n154 VDD.n152 0.108313
R293 VDD.n156 VDD.n154 0.108313
R294 VDD.n158 VDD.n156 0.108313
R295 VDD.n163 VDD.n161 0.108313
R296 VDD.n165 VDD.n163 0.108313
R297 VDD.n150 VDD.n149 0.107844
R298 VDD VDD.n165 0.107375
R299 VDD.n54 VDD.n53 0.106438
R300 VDD.n43 VDD.n42 0.099875
R301 VDD.n55 VDD.n54 0.0967182
R302 VDD.n119 VDD.n118 0.092375
R303 VDD.n34 VDD.n33 0.0895625
R304 VDD.n110 VDD.n109 0.0890938
R305 VDD.n33 VDD.n32 0.0844062
R306 VDD.n131 VDD.n130 0.083
R307 VDD.n128 VDD.n127 0.0820625
R308 VDD.n198 VDD.n197 0.07925
R309 VDD.n192 VDD.n191 0.0783125
R310 VDD.n122 VDD.n121 0.0755
R311 VDD.n40 VDD.n39 0.068
R312 VDD.n113 VDD.n112 0.0651875
R313 VDD.n145 VDD.n143 0.0600312
R314 VDD.n159 VDD.n158 0.0590938
R315 VDD.n49 VDD.n48 0.0576875
R316 VDD.n174 VDD.n173 0.054875
R317 VDD.n173 VDD.n172 0.0539375
R318 VDD.n48 VDD.n47 0.051125
R319 VDD.n161 VDD.n159 0.0497188
R320 VDD.n143 VDD.n142 0.0487812
R321 VDD.n114 VDD.n113 0.043625
R322 VDD.n39 VDD.n38 0.0408125
R323 VDD.n123 VDD.n122 0.0333125
R324 VDD.n193 VDD.n192 0.0305
R325 VDD.n197 VDD.n196 0.0295625
R326 VDD.n127 VDD.n126 0.02675
R327 VDD.n35 VDD.n34 0.01925
R328 VDD.n118 VDD.n117 0.0164375
R329 VDD.n133 VDD.n132 0.0159688
R330 VDD.n109 VDD.n108 0.0140938
R331 VDD.n136 VDD.n135 0.0112812
R332 VDD.n204 VDD.n201 0.0103438
R333 VDD.n56 VDD.n55 0.00977193
R334 VDD.n44 VDD.n43 0.0089375
R335 VDD.n107 VDD.n102 0.008
R336 VDD.n108 VDD.n107 0.006125
R337 VDD.n57 VDD.n18 0.00565625
R338 VDD.n56 VDD.n20 0.00378125
R339 VDD.n132 VDD.n131 0.0033125
R340 VDD.n178 VDD.n177 0.00284375
R341 VDD.n53 VDD.n52 0.002375
R342 VDD.n133 VDD.n57 0.002375
R343 VDD.n100 VDD.n99 0.00209515
R344 VDD.n101 VDD.n100 0.00177952
R345 VDD VDD.n204 0.0014375
R346 VDD.n152 VDD.n150 0.00096875
R347 G1_2.n130 G1_2.n129 103.823
R348 G1_2.n128 G1_2.n127 103.823
R349 G1_2.n126 G1_2.n125 103.823
R350 G1_2.n124 G1_2.n123 103.823
R351 G1_2.n108 G1_2.n105 90.2366
R352 G1_2.n54 G1_2.n51 90.0338
R353 G1_2.n21 G1_2.n18 89.6266
R354 G1_2.n113 G1_2.n112 89.2199
R355 G1_2.n86 G1_2.n85 86.0167
R356 G1_2.n46 G1_2.n43 85.9783
R357 G1_2.n48 G1_2.n47 25.6154
R358 G1_2.n102 G1_2.n101 25.6154
R359 G1_2.n112 G1_2.n109 25.6154
R360 G1_2.n59 G1_2.n55 25.5424
R361 G1_2.n91 G1_2.n90 25.3234
R362 G1_2.n84 G1_2.n83 25.3234
R363 G1_2.n70 G1_2.n69 25.3234
R364 G1_2.n25 G1_2.n22 25.3234
R365 G1_2.n15 G1_2.n14 25.1774
R366 G1_2.n129 G1_2.n128 21.0894
R367 G1_2.n127 G1_2.n126 21.0894
R368 G1_2.n125 G1_2.n124 21.0894
R369 G1_2.n123 G1_2.n122 21.0894
R370 G1_2.n15 G1_2.t29 14.1625
R371 G1_2.n47 G1_2.t31 14.0895
R372 G1_2.n48 G1_2.t15 14.0895
R373 G1_2.n55 G1_2.t19 14.0895
R374 G1_2.n58 G1_2.t43 14.0895
R375 G1_2.n101 G1_2.t7 14.0895
R376 G1_2.n102 G1_2.t27 14.0895
R377 G1_2.n109 G1_2.t25 14.0895
R378 G1_2.n112 G1_2.t45 14.0895
R379 G1_2.n41 G1_2.t41 14.0535
R380 G1_2.n90 G1_2.t39 14.0165
R381 G1_2.n83 G1_2.t35 14.0165
R382 G1_2.n84 G1_2.t13 14.0165
R383 G1_2.n70 G1_2.t17 14.0165
R384 G1_2.n69 G1_2.t11 14.0165
R385 G1_2.n14 G1_2.t9 14.0165
R386 G1_2.n22 G1_2.t37 14.0165
R387 G1_2.n118 G1_2.t33 14.0165
R388 G1_2.n92 G1_2.t23 13.8688
R389 G1_2.n26 G1_2.t21 13.6515
R390 G1_2.n129 G1_2.t77 13.4325
R391 G1_2.n128 G1_2.t68 13.4325
R392 G1_2.n127 G1_2.t67 13.4325
R393 G1_2.n126 G1_2.t74 13.4325
R394 G1_2.n125 G1_2.t78 13.4325
R395 G1_2.n124 G1_2.t70 13.4325
R396 G1_2.n123 G1_2.t71 13.4325
R397 G1_2.n122 G1_2.t64 13.4325
R398 G1_2.n33 G1_2.t60 9.73306
R399 G1_2.n133 G1_2.t63 8.6145
R400 G1_2.n94 G1_2.n86 8.02477
R401 G1_2.n130 G1_2.n0 8.0005
R402 G1_2.n83 G1_2.n82 7.31048
R403 G1_2.n14 G1_2.n13 7.28939
R404 G1_2.n112 G1_2.n111 6.99488
R405 G1_2.n18 G1_2.n17 6.98985
R406 G1_2.n89 G1_2.n88 6.98577
R407 G1_2.n105 G1_2.n104 6.9857
R408 G1_2.n46 G1_2.n45 6.98386
R409 G1_2.n54 G1_2.n53 6.98202
R410 G1_2.n51 G1_2.n50 6.98202
R411 G1_2.n68 G1_2.n67 6.92657
R412 G1_2.n85 G1_2.n80 6.92657
R413 G1_2.n21 G1_2.n20 6.92657
R414 G1_2.n108 G1_2.n107 6.92646
R415 G1_2.n38 G1_2.n37 5.62918
R416 G1_2.n135 G1_2.n121 5.6219
R417 G1_2.n96 G1_2.n95 4.5005
R418 G1_2.n121 G1_2.n120 4.5005
R419 G1_2.n57 G1_2.n56 4.3805
R420 G1_2.n43 G1_2.n42 4.11505
R421 G1_2.n93 G1_2.n92 3.94099
R422 G1_2.n35 G1_2.n34 3.4914
R423 G1_2.n35 G1_2.n33 3.48541
R424 G1_2.n117 G1_2.n113 3.152
R425 G1_2.n74 G1_2.n73 2.96161
R426 G1_2.n39 G1_2.n31 2.95451
R427 G1_2.n116 G1_2.n115 2.94775
R428 G1_2.n97 G1_2.n78 2.94616
R429 G1_2.n62 G1_2.n61 2.93059
R430 G1_2.n4 G1_2.n3 2.92692
R431 G1_2.n9 G1_2.n8 2.9268
R432 G1_2.n29 G1_2.n28 2.91729
R433 G1_2.n64 G1_2.n59 2.88761
R434 G1_2.n101 G1_2.n100 2.88761
R435 G1_2.n135 G1_2.n134 2.88564
R436 G1_2.n37 G1_2.n36 2.88464
R437 G1_2.n27 G1_2.n26 2.86878
R438 G1_2.n40 G1_2.n39 2.86794
R439 G1_2.n98 G1_2.n97 2.62905
R440 G1_2.n134 G1_2.n133 2.3365
R441 G1_2.n76 G1_2.n75 2.2505
R442 G1_2.n65 G1_2.n64 2.2505
R443 G1_2.n100 G1_2.n99 2.2505
R444 G1_2.n24 G1_2.n23 2.22892
R445 G1_2.n131 G1_2.n130 2.1175
R446 G1_2.n111 G1_2.t46 1.8205
R447 G1_2.n111 G1_2.n110 1.8205
R448 G1_2.n107 G1_2.t1 1.8205
R449 G1_2.n107 G1_2.n106 1.8205
R450 G1_2.n104 G1_2.t28 1.8205
R451 G1_2.n104 G1_2.n103 1.8205
R452 G1_2.n8 G1_2.t22 1.8205
R453 G1_2.n8 G1_2.n7 1.8205
R454 G1_2.n67 G1_2.t56 1.8205
R455 G1_2.n67 G1_2.n66 1.8205
R456 G1_2.n88 G1_2.t5 1.8205
R457 G1_2.n88 G1_2.n87 1.8205
R458 G1_2.n78 G1_2.t24 1.8205
R459 G1_2.n78 G1_2.n77 1.8205
R460 G1_2.n80 G1_2.t57 1.8205
R461 G1_2.n80 G1_2.n79 1.8205
R462 G1_2.n82 G1_2.t36 1.8205
R463 G1_2.n82 G1_2.n81 1.8205
R464 G1_2.n73 G1_2.t18 1.8205
R465 G1_2.n73 G1_2.n72 1.8205
R466 G1_2.n20 G1_2.t50 1.8205
R467 G1_2.n20 G1_2.n19 1.8205
R468 G1_2.n17 G1_2.t30 1.8205
R469 G1_2.n17 G1_2.n16 1.8205
R470 G1_2.n13 G1_2.t48 1.8205
R471 G1_2.n13 G1_2.n12 1.8205
R472 G1_2.n53 G1_2.t0 1.8205
R473 G1_2.n53 G1_2.n52 1.8205
R474 G1_2.n50 G1_2.t16 1.8205
R475 G1_2.n50 G1_2.n49 1.8205
R476 G1_2.n45 G1_2.t53 1.8205
R477 G1_2.n45 G1_2.n44 1.8205
R478 G1_2.n31 G1_2.t42 1.8205
R479 G1_2.n31 G1_2.n30 1.8205
R480 G1_2.n61 G1_2.t44 1.8205
R481 G1_2.n61 G1_2.n60 1.8205
R482 G1_2.n3 G1_2.t47 1.8205
R483 G1_2.n3 G1_2.n2 1.8205
R484 G1_2.n115 G1_2.t6 1.8205
R485 G1_2.n115 G1_2.n114 1.8205
R486 G1_2.n75 G1_2.n71 1.61816
R487 G1_2.n65 G1_2.n29 1.41264
R488 G1_2.n99 G1_2.n98 1.38535
R489 G1_2.n101 G1_2.n1 1.20181
R490 G1_2.n71 G1_2.n70 0.853387
R491 G1_2.n99 G1_2.n65 0.696503
R492 G1_2.n18 G1_2.n15 0.642258
R493 G1_2.n85 G1_2.n84 0.384711
R494 G1_2.n69 G1_2.n68 0.384711
R495 G1_2.n22 G1_2.n21 0.384711
R496 G1_2.n26 G1_2.n25 0.3655
R497 G1_2.n109 G1_2.n108 0.298459
R498 G1_2.n132 G1_2.n131 0.292201
R499 G1_2.n25 G1_2.n24 0.231026
R500 G1_2.n51 G1_2.n48 0.223969
R501 G1_2.n55 G1_2.n54 0.223969
R502 G1_2.n90 G1_2.n89 0.154184
R503 G1_2.n47 G1_2.n46 0.14948
R504 G1_2.n58 G1_2.n57 0.1465
R505 G1_2.n92 G1_2.n91 0.143972
R506 G1_2.n120 G1_2.n119 0.140885
R507 G1_2.n42 G1_2.n40 0.133227
R508 G1_2.n98 G1_2.n76 0.120105
R509 G1_2.n105 G1_2.n102 0.0749898
R510 G1_2.n59 G1_2.n58 0.0735
R511 G1_2.n119 G1_2.n118 0.0735
R512 G1_2.n134 G1_2.n132 0.0734811
R513 G1_2.n63 G1_2.n62 0.055602
R514 G1_2.n5 G1_2.n4 0.0537653
R515 G1_2.n10 G1_2.n9 0.0519286
R516 G1_2.n42 G1_2.n41 0.037206
R517 G1_2.n117 G1_2.n116 0.0356143
R518 G1_2.n39 G1_2.n38 0.021405
R519 G1_2.n28 G1_2.n27 0.0200941
R520 G1_2.n75 G1_2.n74 0.019821
R521 G1_2.n97 G1_2.n96 0.019259
R522 G1_2.n96 G1_2.n94 0.01175
R523 G1_2.n28 G1_2.n11 0.0060102
R524 G1_2.n100 G1_2.n5 0.0060102
R525 G1_2.n94 G1_2.n93 0.00425
R526 G1_2.n64 G1_2.n63 0.00417347
R527 G1_2.n121 G1_2.n117 0.00417347
R528 G1_2.n10 G1_2.n6 0.00293243
R529 G1_2 G1_2.n0 0.0025
R530 G1_2.n11 G1_2.n10 0.00233673
R531 G1_2.n38 G1_2.n32 0.00233673
R532 G1_2.n37 G1_2.n35 0.0015
R533 G1_2 G1_2.n135 0.0015
R534 SD1_1.n28 SD1_1.t17 4.5505
R535 SD1_1.n28 SD1_1.n27 4.5505
R536 SD1_1.n1 SD1_1.t3 4.5505
R537 SD1_1.n1 SD1_1.n0 4.5505
R538 SD1_1.n3 SD1_1.t13 4.5505
R539 SD1_1.n3 SD1_1.n2 4.5505
R540 SD1_1.n5 SD1_1.t8 4.5505
R541 SD1_1.n5 SD1_1.n4 4.5505
R542 SD1_1.n7 SD1_1.t19 4.5505
R543 SD1_1.n7 SD1_1.n6 4.5505
R544 SD1_1.n9 SD1_1.t2 4.5505
R545 SD1_1.n9 SD1_1.n8 4.5505
R546 SD1_1.n11 SD1_1.t18 4.5505
R547 SD1_1.n11 SD1_1.n10 4.5505
R548 SD1_1.n13 SD1_1.t5 4.5505
R549 SD1_1.n13 SD1_1.n12 4.5505
R550 SD1_1.n15 SD1_1.t12 4.5505
R551 SD1_1.n15 SD1_1.n14 4.5505
R552 SD1_1.n17 SD1_1.t11 4.5505
R553 SD1_1.n17 SD1_1.n16 4.5505
R554 SD1_1.n18 SD1_1.n17 3.17149
R555 SD1_1.n19 SD1_1.n13 2.77857
R556 SD1_1.n25 SD1_1.n1 2.54881
R557 SD1_1.n18 SD1_1.n15 2.54881
R558 SD1_1.n24 SD1_1.n3 2.54872
R559 SD1_1.n23 SD1_1.n5 2.54872
R560 SD1_1.n22 SD1_1.n7 2.54872
R561 SD1_1.n20 SD1_1.n11 2.54872
R562 SD1_1.n21 SD1_1.n9 2.54854
R563 SD1_1.n31 SD1_1.n30 2.25795
R564 SD1_1.n29 SD1_1.n26 2.2439
R565 SD1_1.n29 SD1_1.n28 1.65397
R566 SD1_1.n19 SD1_1.n18 0.635915
R567 SD1_1.n24 SD1_1.n23 0.627793
R568 SD1_1.n21 SD1_1.n20 0.626983
R569 SD1_1.n25 SD1_1.n24 0.623305
R570 SD1_1.n22 SD1_1.n21 0.622387
R571 SD1_1.n23 SD1_1.n22 0.621579
R572 SD1_1.n20 SD1_1.n19 0.614074
R573 SD1_1.n26 SD1_1.n25 0.609182
R574 SD1_1.n31 SD1_1.n26 0.0151956
R575 SD1_1.n30 SD1_1.n29 0.010363
R576 SD1_1 SD1_1.n31 0.00163924
R577 G2_1.n133 G2_1.n132 74.2622
R578 G2_1.n26 G2_1.n23 71.202
R579 G2_1.n28 G2_1.t37 37.4414
R580 G2_1.n116 G2_1.t43 37.4414
R581 G2_1.n132 G2_1.n131 21.0894
R582 G2_1.n131 G2_1.n130 21.0894
R583 G2_1.n130 G2_1.n129 21.0894
R584 G2_1.n129 G2_1.n128 21.0894
R585 G2_1.n128 G2_1.n127 21.0894
R586 G2_1.n127 G2_1.n126 21.0894
R587 G2_1.n126 G2_1.n125 21.0894
R588 G2_1.n125 G2_1.n124 21.0894
R589 G2_1.n124 G2_1.n123 21.0894
R590 G2_1.n15 G2_1.n14 21.0894
R591 G2_1.n16 G2_1.n15 21.0894
R592 G2_1.n17 G2_1.n16 21.0894
R593 G2_1.n18 G2_1.n17 21.0894
R594 G2_1.n19 G2_1.n18 21.0894
R595 G2_1.n20 G2_1.n19 21.0894
R596 G2_1.n21 G2_1.n20 21.0894
R597 G2_1.n22 G2_1.n21 21.0894
R598 G2_1.n23 G2_1.n22 21.0894
R599 G2_1.n131 G2_1.t67 16.5715
R600 G2_1.n130 G2_1.t88 16.5715
R601 G2_1.n127 G2_1.t80 16.5715
R602 G2_1.n126 G2_1.t64 16.5715
R603 G2_1.n123 G2_1.t85 16.5715
R604 G2_1.n14 G2_1.t89 16.5715
R605 G2_1.n17 G2_1.t81 16.5715
R606 G2_1.n18 G2_1.t66 16.5715
R607 G2_1.n21 G2_1.t76 16.5715
R608 G2_1.n22 G2_1.t60 16.5715
R609 G2_1.n132 G2_1.t71 16.3525
R610 G2_1.n129 G2_1.t62 16.3525
R611 G2_1.n128 G2_1.t78 16.3525
R612 G2_1.n125 G2_1.t77 16.3525
R613 G2_1.n124 G2_1.t61 16.3525
R614 G2_1.n15 G2_1.t63 16.3525
R615 G2_1.n16 G2_1.t84 16.3525
R616 G2_1.n19 G2_1.t87 16.3525
R617 G2_1.n20 G2_1.t73 16.3525
R618 G2_1.n23 G2_1.t65 16.3525
R619 G2_1.n104 G2_1.t19 14.0165
R620 G2_1.n101 G2_1.t53 14.0165
R621 G2_1.n92 G2_1.t21 14.0165
R622 G2_1.n89 G2_1.t45 14.0165
R623 G2_1.n82 G2_1.t29 14.0165
R624 G2_1.n79 G2_1.t47 14.0165
R625 G2_1.n70 G2_1.t35 14.0165
R626 G2_1.n67 G2_1.t39 14.0165
R627 G2_1.n62 G2_1.t25 14.0165
R628 G2_1.n59 G2_1.t51 14.0165
R629 G2_1.n52 G2_1.t31 14.0165
R630 G2_1.n49 G2_1.t41 14.0165
R631 G2_1.n44 G2_1.t23 14.0165
R632 G2_1.n41 G2_1.t55 14.0165
R633 G2_1.n32 G2_1.t27 14.0165
R634 G2_1.n29 G2_1.t49 14.0165
R635 G2_1.n113 G2_1.t17 14.0165
R636 G2_1.n115 G2_1.t33 13.7245
R637 G2_1.n30 G2_1.n29 4.0005
R638 G2_1.n33 G2_1.n32 4.0005
R639 G2_1.n42 G2_1.n41 4.0005
R640 G2_1.n45 G2_1.n44 4.0005
R641 G2_1.n50 G2_1.n49 4.0005
R642 G2_1.n53 G2_1.n52 4.0005
R643 G2_1.n60 G2_1.n59 4.0005
R644 G2_1.n63 G2_1.n62 4.0005
R645 G2_1.n68 G2_1.n67 4.0005
R646 G2_1.n71 G2_1.n70 4.0005
R647 G2_1.n80 G2_1.n79 4.0005
R648 G2_1.n83 G2_1.n82 4.0005
R649 G2_1.n90 G2_1.n89 4.0005
R650 G2_1.n93 G2_1.n92 4.0005
R651 G2_1.n102 G2_1.n101 4.0005
R652 G2_1.n105 G2_1.n104 4.0005
R653 G2_1.n114 G2_1.n113 4.0005
R654 G2_1.n118 G2_1.n117 4.0005
R655 G2_1.n26 G2_1.n25 3.58493
R656 G2_1.n108 G2_1.n107 3.57898
R657 G2_1.n86 G2_1.n85 3.57507
R658 G2_1.n133 G2_1.n122 3.5665
R659 G2_1.n46 G2_1.n11 3.53988
R660 G2_1.n99 G2_1.n98 3.53861
R661 G2_1.n77 G2_1.n76 3.53721
R662 G2_1.n74 G2_1.n73 3.53202
R663 G2_1.n96 G2_1.n95 3.53202
R664 G2_1.n87 G2_1.n1 3.52224
R665 G2_1.n65 G2_1.n3 3.51637
R666 G2_1.n47 G2_1.n9 3.51246
R667 G2_1.n57 G2_1.n56 3.51057
R668 G2_1.n36 G2_1.n35 3.50854
R669 G2_1.n111 G2_1.n110 3.50645
R670 G2_1.n39 G2_1.n38 3.49699
R671 G2_1.n64 G2_1.n5 3.49116
R672 G2_1.n54 G2_1.n7 3.4806
R673 G2_1.n134 G2_1.n120 3.46399
R674 G2_1.n27 G2_1.n13 3.45496
R675 G2_1.n104 G2_1.n103 2.3365
R676 G2_1.n101 G2_1.n100 2.3365
R677 G2_1.n92 G2_1.n91 2.3365
R678 G2_1.n89 G2_1.n88 2.3365
R679 G2_1.n82 G2_1.n81 2.3365
R680 G2_1.n79 G2_1.n78 2.3365
R681 G2_1.n70 G2_1.n69 2.3365
R682 G2_1.n67 G2_1.n66 2.3365
R683 G2_1.n62 G2_1.n61 2.3365
R684 G2_1.n59 G2_1.n58 2.3365
R685 G2_1.n52 G2_1.n51 2.3365
R686 G2_1.n49 G2_1.n48 2.3365
R687 G2_1.n44 G2_1.n43 2.3365
R688 G2_1.n41 G2_1.n40 2.3365
R689 G2_1.n32 G2_1.n31 2.3365
R690 G2_1.n29 G2_1.n28 2.3365
R691 G2_1.n113 G2_1.n112 2.3365
R692 G2_1.n117 G2_1.n116 2.3365
R693 G2_1.n107 G2_1.t20 1.6385
R694 G2_1.n107 G2_1.n106 1.6385
R695 G2_1.n110 G2_1.t1 1.6385
R696 G2_1.n110 G2_1.n109 1.6385
R697 G2_1.n95 G2_1.t22 1.6385
R698 G2_1.n95 G2_1.n94 1.6385
R699 G2_1.n98 G2_1.t12 1.6385
R700 G2_1.n98 G2_1.n97 1.6385
R701 G2_1.n85 G2_1.t30 1.6385
R702 G2_1.n85 G2_1.n84 1.6385
R703 G2_1.n1 G2_1.t5 1.6385
R704 G2_1.n1 G2_1.n0 1.6385
R705 G2_1.n73 G2_1.t36 1.6385
R706 G2_1.n73 G2_1.n72 1.6385
R707 G2_1.n76 G2_1.t10 1.6385
R708 G2_1.n76 G2_1.n75 1.6385
R709 G2_1.n5 G2_1.t26 1.6385
R710 G2_1.n5 G2_1.n4 1.6385
R711 G2_1.n3 G2_1.t7 1.6385
R712 G2_1.n3 G2_1.n2 1.6385
R713 G2_1.n7 G2_1.t32 1.6385
R714 G2_1.n7 G2_1.n6 1.6385
R715 G2_1.n56 G2_1.t14 1.6385
R716 G2_1.n56 G2_1.n55 1.6385
R717 G2_1.n11 G2_1.t24 1.6385
R718 G2_1.n11 G2_1.n10 1.6385
R719 G2_1.n9 G2_1.t8 1.6385
R720 G2_1.n9 G2_1.n8 1.6385
R721 G2_1.n35 G2_1.t28 1.6385
R722 G2_1.n35 G2_1.n34 1.6385
R723 G2_1.n38 G2_1.t6 1.6385
R724 G2_1.n38 G2_1.n37 1.6385
R725 G2_1.n120 G2_1.t34 1.6385
R726 G2_1.n120 G2_1.n119 1.6385
R727 G2_1.n122 G2_1.t15 1.6385
R728 G2_1.n122 G2_1.n121 1.6385
R729 G2_1.n13 G2_1.t9 1.6385
R730 G2_1.n13 G2_1.n12 1.6385
R731 G2_1.n25 G2_1.t38 1.6385
R732 G2_1.n25 G2_1.n24 1.6385
R733 G2_1 G2_1.n134 0.362318
R734 G2_1.n117 G2_1.n115 0.2925
R735 G2_1.n83 G2_1.n80 0.253351
R736 G2_1.n118 G2_1.n114 0.197599
R737 G2_1.n33 G2_1.n30 0.197599
R738 G2_1.n53 G2_1.n50 0.197599
R739 G2_1.n71 G2_1.n68 0.197599
R740 G2_1.n93 G2_1.n90 0.197599
R741 G2_1.n45 G2_1.n42 0.172031
R742 G2_1.n63 G2_1.n60 0.172031
R743 G2_1.n105 G2_1.n102 0.172031
R744 G2_1.n39 G2_1.n36 0.100499
R745 G2_1.n47 G2_1.n46 0.093148
R746 G2_1.n65 G2_1.n64 0.0926899
R747 G2_1.n57 G2_1.n54 0.0817532
R748 G2_1.n87 G2_1.n86 0.0807174
R749 G2_1.n77 G2_1.n74 0.0742956
R750 G2_1.n99 G2_1.n96 0.0727632
R751 G2_1.n74 G2_1.n71 0.0708476
R752 G2_1.n96 G2_1.n93 0.0705535
R753 G2_1.n111 G2_1.n108 0.0688207
R754 G2_1.n114 G2_1.n111 0.0665096
R755 G2_1.n90 G2_1.n87 0.0655603
R756 G2_1.n68 G2_1.n65 0.0636092
R757 G2_1.n54 G2_1.n53 0.061636
R758 G2_1.n50 G2_1.n47 0.0606109
R759 G2_1.n36 G2_1.n33 0.0579026
R760 G2_1.n108 G2_1.n105 0.049875
R761 G2_1.n86 G2_1.n83 0.0488673
R762 G2_1.n102 G2_1.n99 0.0443624
R763 G2_1.n46 G2_1.n45 0.0432184
R764 G2_1.n80 G2_1.n77 0.0423084
R765 G2_1.n60 G2_1.n57 0.0409019
R766 G2_1.n64 G2_1.n63 0.0397098
R767 G2_1.n42 G2_1.n39 0.0396398
R768 G2_1.n30 G2_1.n27 0.0223182
R769 G2_1.n134 G2_1.n133 0.00742308
R770 G2_1 G2_1.n118 0.00504545
R771 G2_1.n27 G2_1.n26 0.00495545
R772 VSS.n12 VSS.n11 869.582
R773 VSS.n137 VSS.n136 393.498
R774 VSS.n106 VSS.t12 223.469
R775 VSS.n103 VSS.t58 208.894
R776 VSS.n101 VSS.t7 194.321
R777 VSS.n99 VSS.t48 179.746
R778 VSS.n97 VSS.t34 165.173
R779 VSS.n94 VSS.t50 150.599
R780 VSS.n135 VSS.t1 150.599
R781 VSS.n74 VSS.t55 138.453
R782 VSS.n92 VSS.t2 136.024
R783 VSS.n77 VSS.t4 123.879
R784 VSS.n218 VSS.t41 114.472
R785 VSS.n79 VSS.t15 109.305
R786 VSS.n215 VSS.t65 107.007
R787 VSS.n213 VSS.t16 99.5411
R788 VSS.n81 VSS.t47 94.7314
R789 VSS.n211 VSS.t42 92.0755
R790 VSS.n209 VSS.t64 84.61
R791 VSS.n83 VSS.t11 80.1575
R792 VSS.n206 VSS.t61 77.1445
R793 VSS.n228 VSS.t43 77.1445
R794 VSS.n204 VSS.t23 69.6789
R795 VSS.n86 VSS.t29 65.5835
R796 VSS.n202 VSS.t18 62.2134
R797 VSS.n10 VSS.t32 58.2965
R798 VSS.n155 VSS.t25 54.815
R799 VSS.n200 VSS.t54 54.7478
R800 VSS.n88 VSS.t63 51.0095
R801 VSS.n197 VSS.t17 47.2823
R802 VSS.n195 VSS.t40 39.8167
R803 VSS.n193 VSS.t46 32.3512
R804 VSS.n191 VSS.t62 24.8856
R805 VSS.n124 VSS.t37 22.9229
R806 VSS.n188 VSS.t0 17.4201
R807 VSS.n121 VSS.t33 16.9432
R808 VSS.n35 VSS.t44 13.6873
R809 VSS.n114 VSS.t19 12.9566
R810 VSS.n179 VSS.t60 12.4431
R811 VSS.n120 VSS.t8 10.9634
R812 VSS.n186 VSS.t45 9.95456
R813 VSS.n115 VSS.t3 6.97689
R814 VSS.n156 VSS.t26 6.44293
R815 VSS.n22 VSS.n21 6.40927
R816 VSS.n335 VSS.t59 6.40764
R817 VSS.n322 VSS.t67 6.4068
R818 VSS.n324 VSS.n311 6.4068
R819 VSS.n306 VSS.n252 6.35296
R820 VSS.n146 VSS.n145 6.34765
R821 VSS.n62 VSS.n61 5.4245
R822 VSS.n40 VSS.n39 5.41019
R823 VSS.n304 VSS.t104 5.3939
R824 VSS.n251 VSS.t99 5.3802
R825 VSS.n224 VSS.n221 5.2005
R826 VSS.n231 VSS.n229 5.2005
R827 VSS.n36 VSS.n34 5.2005
R828 VSS.n36 VSS.n32 5.2005
R829 VSS.n180 VSS.n179 5.2005
R830 VSS.n183 VSS.n182 5.2005
R831 VSS.n185 VSS.n184 5.2005
R832 VSS.n187 VSS.n186 5.2005
R833 VSS.n189 VSS.n188 5.2005
R834 VSS.n192 VSS.n191 5.2005
R835 VSS.n194 VSS.n193 5.2005
R836 VSS.n196 VSS.n195 5.2005
R837 VSS.n198 VSS.n197 5.2005
R838 VSS.n201 VSS.n200 5.2005
R839 VSS.n203 VSS.n202 5.2005
R840 VSS.n205 VSS.n204 5.2005
R841 VSS.n207 VSS.n206 5.2005
R842 VSS.n210 VSS.n209 5.2005
R843 VSS.n212 VSS.n211 5.2005
R844 VSS.n214 VSS.n213 5.2005
R845 VSS.n216 VSS.n215 5.2005
R846 VSS.n219 VSS.n218 5.2005
R847 VSS.n231 VSS.n228 5.2005
R848 VSS.n112 VSS.n111 5.2005
R849 VSS.n18 VSS.n17 5.2005
R850 VSS.n144 VSS.n143 5.2005
R851 VSS.n163 VSS.n147 5.2005
R852 VSS.n162 VSS.n148 5.2005
R853 VSS.n161 VSS.n149 5.2005
R854 VSS.n159 VSS.n152 5.2005
R855 VSS.n158 VSS.n153 5.2005
R856 VSS.n157 VSS.n154 5.2005
R857 VSS.n156 VSS.n155 5.2005
R858 VSS.n133 VSS.n114 5.2005
R859 VSS.n132 VSS.n115 5.2005
R860 VSS.n130 VSS.n118 5.2005
R861 VSS.n129 VSS.n119 5.2005
R862 VSS.n128 VSS.n120 5.2005
R863 VSS.n127 VSS.n121 5.2005
R864 VSS.n125 VSS.n124 5.2005
R865 VSS.n139 VSS.n137 5.2005
R866 VSS.n75 VSS.n74 5.2005
R867 VSS.n78 VSS.n77 5.2005
R868 VSS.n80 VSS.n79 5.2005
R869 VSS.n82 VSS.n81 5.2005
R870 VSS.n84 VSS.n83 5.2005
R871 VSS.n87 VSS.n86 5.2005
R872 VSS.n89 VSS.n88 5.2005
R873 VSS.n91 VSS.n90 5.2005
R874 VSS.n93 VSS.n92 5.2005
R875 VSS.n95 VSS.n94 5.2005
R876 VSS.n98 VSS.n97 5.2005
R877 VSS.n100 VSS.n99 5.2005
R878 VSS.n102 VSS.n101 5.2005
R879 VSS.n104 VSS.n103 5.2005
R880 VSS.n107 VSS.n106 5.2005
R881 VSS.n139 VSS.n135 5.2005
R882 VSS.n13 VSS.n10 5.2005
R883 VSS.n13 VSS.n12 5.2005
R884 VSS.n119 VSS.t52 4.98363
R885 VSS.n182 VSS.t24 4.97753
R886 VSS.n36 VSS.n35 4.5005
R887 VSS.n231 VSS.n230 4.5005
R888 VSS.n139 VSS.n138 4.5005
R889 VSS.n13 VSS.n8 4.5005
R890 VSS.n69 VSS.n60 4.1554
R891 VSS.n71 VSS.n70 3.92314
R892 VSS.n72 VSS.n71 3.84637
R893 VSS.n338 VSS.n337 3.83363
R894 VSS.n217 VSS.n170 3.75507
R895 VSS.n208 VSS.n172 3.75507
R896 VSS.n199 VSS.n174 3.75507
R897 VSS.n190 VSS.n176 3.75507
R898 VSS.n181 VSS.n178 3.75507
R899 VSS.n275 VSS.n268 3.75507
R900 VSS.n281 VSS.n264 3.75507
R901 VSS.n287 VSS.n260 3.75507
R902 VSS.n293 VSS.n256 3.75507
R903 VSS.n296 VSS.n254 3.75507
R904 VSS.n290 VSS.n258 3.75507
R905 VSS.n284 VSS.n262 3.75507
R906 VSS.n278 VSS.n266 3.75507
R907 VSS.n272 VSS.n270 3.75507
R908 VSS.n55 VSS.n46 3.74137
R909 VSS.n50 VSS.n48 3.74137
R910 VSS.n240 VSS.n236 3.74137
R911 VSS.n245 VSS.n234 3.74137
R912 VSS.n126 VSS.n123 3.68072
R913 VSS.n131 VSS.n117 3.68072
R914 VSS.n317 VSS.n313 3.6768
R915 VSS.n329 VSS.n310 3.6768
R916 VSS.n105 VSS.n1 3.64159
R917 VSS.n96 VSS.n3 3.64159
R918 VSS.n85 VSS.n5 3.64159
R919 VSS.n76 VSS.n7 3.64159
R920 VSS.n160 VSS.n151 3.61615
R921 VSS.n308 VSS.n307 2.89175
R922 VSS.n19 VSS.n18 2.86051
R923 VSS.n151 VSS.t53 2.7305
R924 VSS.n151 VSS.n150 2.7305
R925 VSS.n313 VSS.t134 2.7305
R926 VSS.n313 VSS.n312 2.7305
R927 VSS.n310 VSS.t49 2.7305
R928 VSS.n310 VSS.n309 2.7305
R929 VSS.n123 VSS.t57 2.7305
R930 VSS.n123 VSS.n122 2.7305
R931 VSS.n117 VSS.t66 2.7305
R932 VSS.n117 VSS.n116 2.7305
R933 VSS.n1 VSS.t137 2.7305
R934 VSS.n1 VSS.n0 2.7305
R935 VSS.n3 VSS.t51 2.7305
R936 VSS.n3 VSS.n2 2.7305
R937 VSS.n5 VSS.t68 2.7305
R938 VSS.n5 VSS.n4 2.7305
R939 VSS.n7 VSS.t56 2.7305
R940 VSS.n7 VSS.n6 2.7305
R941 VSS.n42 VSS.n41 2.60175
R942 VSS.n225 VSS.n224 2.60175
R943 VSS.n64 VSS.n63 2.60175
R944 VSS.n300 VSS.n299 2.60175
R945 VSS.n30 VSS.n28 2.60175
R946 VSS.n167 VSS.n166 2.60175
R947 VSS.n113 VSS.n112 2.60175
R948 VSS.n166 VSS.n165 2.601
R949 VSS.n18 VSS.n16 2.601
R950 VSS.n112 VSS.n110 2.601
R951 VSS.n28 VSS.n27 2.601
R952 VSS.n224 VSS.n223 2.601
R953 VSS.n226 VSS.n225 2.601
R954 VSS.n339 VSS.n113 2.601
R955 VSS.n27 VSS.n26 2.48901
R956 VSS.n34 VSS.n33 2.48901
R957 VSS.n184 VSS.t22 2.48901
R958 VSS.n304 VSS.n303 2.41785
R959 VSS.n232 VSS.n231 2.41764
R960 VSS.n146 VSS.n144 2.41728
R961 VSS.n67 VSS.n66 2.40802
R962 VSS.n37 VSS.n36 2.40802
R963 VSS.n140 VSS.n139 2.40798
R964 VSS.n59 VSS.n44 2.40786
R965 VSS.n70 VSS.n38 2.25997
R966 VSS.n307 VSS.n232 2.25167
R967 VSS.n308 VSS.n168 2.2505
R968 VSS.n337 VSS.n336 2.2505
R969 VSS.n71 VSS.n25 2.2505
R970 VSS.n69 VSS.n68 2.2505
R971 VSS.n306 VSS.n305 2.2505
R972 VSS.n144 VSS.n142 2.188
R973 VSS.n30 VSS.n29 2.16377
R974 VSS.n66 VSS.n65 2.13331
R975 VSS.n44 VSS.n43 2.13331
R976 VSS.n13 VSS.n9 2.07862
R977 VSS.n139 VSS.n134 2.02394
R978 VSS.n231 VSS.n227 2.02394
R979 VSS.n303 VSS.n301 2.02394
R980 VSS.n70 VSS.n69 1.87545
R981 VSS.n307 VSS.n306 1.87428
R982 VSS.n170 VSS.t75 1.6385
R983 VSS.n170 VSS.n169 1.6385
R984 VSS.n172 VSS.t119 1.6385
R985 VSS.n172 VSS.n171 1.6385
R986 VSS.n174 VSS.t72 1.6385
R987 VSS.n174 VSS.n173 1.6385
R988 VSS.n176 VSS.t114 1.6385
R989 VSS.n176 VSS.n175 1.6385
R990 VSS.n178 VSS.t129 1.6385
R991 VSS.n178 VSS.n177 1.6385
R992 VSS.n268 VSS.t100 1.6385
R993 VSS.n268 VSS.n267 1.6385
R994 VSS.n264 VSS.t80 1.6385
R995 VSS.n264 VSS.n263 1.6385
R996 VSS.n260 VSS.t126 1.6385
R997 VSS.n260 VSS.n259 1.6385
R998 VSS.n256 VSS.t91 1.6385
R999 VSS.n256 VSS.n255 1.6385
R1000 VSS.n254 VSS.t111 1.6385
R1001 VSS.n254 VSS.n253 1.6385
R1002 VSS.n258 VSS.t83 1.6385
R1003 VSS.n258 VSS.n257 1.6385
R1004 VSS.n262 VSS.t74 1.6385
R1005 VSS.n262 VSS.n261 1.6385
R1006 VSS.n266 VSS.t108 1.6385
R1007 VSS.n266 VSS.n265 1.6385
R1008 VSS.n270 VSS.t103 1.6385
R1009 VSS.n270 VSS.n269 1.6385
R1010 VSS.n46 VSS.t88 1.6385
R1011 VSS.n46 VSS.n45 1.6385
R1012 VSS.n48 VSS.t98 1.6385
R1013 VSS.n48 VSS.n47 1.6385
R1014 VSS.n236 VSS.t105 1.6385
R1015 VSS.n236 VSS.n235 1.6385
R1016 VSS.n234 VSS.t73 1.6385
R1017 VSS.n234 VSS.n233 1.6385
R1018 VSS.n20 VSS.n19 1.56429
R1019 VSS.n32 VSS.n31 1.24476
R1020 VSS.n118 VSS.t69 0.997127
R1021 VSS.n337 VSS.n308 0.650577
R1022 VSS.n16 VSS.n15 0.556908
R1023 VSS.n19 VSS.n13 0.520836
R1024 VSS.n144 VSS.n141 0.514399
R1025 VSS.n110 VSS.n109 0.447533
R1026 VSS.n223 VSS.n222 0.447533
R1027 VSS.n303 VSS.n302 0.430411
R1028 VSS.n140 VSS.n133 0.364923
R1029 VSS.n15 VSS.n14 0.248057
R1030 VSS.n109 VSS.n108 0.24188
R1031 VSS.n163 VSS.n162 0.129952
R1032 VSS.n162 VSS.n161 0.129952
R1033 VSS.n159 VSS.n158 0.129952
R1034 VSS.n158 VSS.n157 0.129952
R1035 VSS.n157 VSS.n156 0.129952
R1036 VSS.n185 VSS.n183 0.129952
R1037 VSS.n187 VSS.n185 0.129952
R1038 VSS.n189 VSS.n187 0.129952
R1039 VSS.n194 VSS.n192 0.129952
R1040 VSS.n196 VSS.n194 0.129952
R1041 VSS.n198 VSS.n196 0.129952
R1042 VSS.n203 VSS.n201 0.129952
R1043 VSS.n205 VSS.n203 0.129952
R1044 VSS.n207 VSS.n205 0.129952
R1045 VSS.n212 VSS.n210 0.129952
R1046 VSS.n214 VSS.n212 0.129952
R1047 VSS.n216 VSS.n214 0.129952
R1048 VSS.n315 VSS.n314 0.129952
R1049 VSS.n316 VSS.n315 0.129952
R1050 VSS.n319 VSS.n318 0.129952
R1051 VSS.n320 VSS.n319 0.129952
R1052 VSS.n321 VSS.n320 0.129952
R1053 VSS.n326 VSS.n325 0.129952
R1054 VSS.n327 VSS.n326 0.129952
R1055 VSS.n328 VSS.n327 0.129952
R1056 VSS.n331 VSS.n330 0.129952
R1057 VSS.n332 VSS.n331 0.129952
R1058 VSS.n274 VSS.n273 0.129952
R1059 VSS.n277 VSS.n276 0.129952
R1060 VSS.n280 VSS.n279 0.129952
R1061 VSS.n283 VSS.n282 0.129952
R1062 VSS.n286 VSS.n285 0.129952
R1063 VSS.n289 VSS.n288 0.129952
R1064 VSS.n292 VSS.n291 0.129952
R1065 VSS.n295 VSS.n294 0.129952
R1066 VSS.n58 VSS.n57 0.129952
R1067 VSS.n57 VSS.n56 0.129952
R1068 VSS.n54 VSS.n53 0.129952
R1069 VSS.n53 VSS.n52 0.129952
R1070 VSS.n52 VSS.n51 0.129952
R1071 VSS.n238 VSS.n237 0.129952
R1072 VSS.n239 VSS.n238 0.129952
R1073 VSS.n242 VSS.n241 0.129952
R1074 VSS.n243 VSS.n242 0.129952
R1075 VSS.n244 VSS.n243 0.129952
R1076 VSS.n247 VSS.n246 0.129952
R1077 VSS.n248 VSS.n247 0.129952
R1078 VSS.n133 VSS.n132 0.129952
R1079 VSS.n130 VSS.n129 0.129952
R1080 VSS.n129 VSS.n128 0.129952
R1081 VSS.n128 VSS.n127 0.129952
R1082 VSS.n80 VSS.n78 0.129952
R1083 VSS.n82 VSS.n80 0.129952
R1084 VSS.n84 VSS.n82 0.129952
R1085 VSS.n89 VSS.n87 0.129952
R1086 VSS.n91 VSS.n89 0.129952
R1087 VSS.n93 VSS.n91 0.129952
R1088 VSS.n95 VSS.n93 0.129952
R1089 VSS.n100 VSS.n98 0.129952
R1090 VSS.n102 VSS.n100 0.129952
R1091 VSS.n104 VSS.n102 0.129952
R1092 VSS.n219 VSS.n217 0.120089
R1093 VSS.n297 VSS.n296 0.120089
R1094 VSS.n107 VSS.n105 0.120089
R1095 VSS.n59 VSS.n58 0.118897
R1096 VSS.n75 VSS.n73 0.117951
R1097 VSS.n330 VSS.n329 0.112692
R1098 VSS.n294 VSS.n293 0.112692
R1099 VSS.n246 VSS.n245 0.112692
R1100 VSS.n161 VSS.n160 0.112075
R1101 VSS.n164 VSS.n163 0.10776
R1102 VSS.n220 VSS.n219 0.10776
R1103 VSS.n333 VSS.n332 0.10776
R1104 VSS.n298 VSS.n297 0.10776
R1105 VSS.n249 VSS.n248 0.10776
R1106 VSS.n210 VSS.n208 0.105295
R1107 VSS.n291 VSS.n290 0.105295
R1108 VSS.n98 VSS.n96 0.105295
R1109 VSS.n76 VSS.n75 0.0985137
R1110 VSS.n325 VSS.n324 0.0978973
R1111 VSS.n288 VSS.n287 0.0978973
R1112 VSS.n241 VSS.n240 0.0978973
R1113 VSS.n317 VSS.n316 0.0911164
R1114 VSS.n201 VSS.n199 0.0905
R1115 VSS.n285 VSS.n284 0.0905
R1116 VSS.n85 VSS.n84 0.0837192
R1117 VSS.n282 VSS.n281 0.0831027
R1118 VSS.n50 VSS.n49 0.0831027
R1119 VSS.n126 VSS.n125 0.0775548
R1120 VSS.n322 VSS.n321 0.0763219
R1121 VSS.n192 VSS.n190 0.0757055
R1122 VSS.n279 VSS.n278 0.0757055
R1123 VSS VSS.n107 0.075089
R1124 VSS.n181 VSS.n180 0.0695411
R1125 VSS.n272 VSS.n271 0.0695411
R1126 VSS.n276 VSS.n275 0.0683082
R1127 VSS.n55 VSS.n54 0.0683082
R1128 VSS.n132 VSS.n131 0.0676918
R1129 VSS.n131 VSS.n130 0.0627603
R1130 VSS.n275 VSS.n274 0.0621438
R1131 VSS.n56 VSS.n55 0.0621438
R1132 VSS.n183 VSS.n181 0.060911
R1133 VSS.n273 VSS.n272 0.060911
R1134 VSS.n190 VSS.n189 0.0547466
R1135 VSS.n278 VSS.n277 0.0547466
R1136 VSS.n323 VSS.n322 0.0541301
R1137 VSS.n127 VSS.n126 0.0528973
R1138 VSS.n281 VSS.n280 0.0473493
R1139 VSS.n51 VSS.n50 0.0473493
R1140 VSS.n87 VSS.n85 0.0467329
R1141 VSS.n199 VSS.n198 0.0399521
R1142 VSS.n284 VSS.n283 0.0399521
R1143 VSS.n318 VSS.n317 0.0393356
R1144 VSS VSS.n340 0.0331712
R1145 VSS.n324 VSS.n323 0.0325548
R1146 VSS.n287 VSS.n286 0.0325548
R1147 VSS.n240 VSS.n239 0.0325548
R1148 VSS.n78 VSS.n76 0.0319384
R1149 VSS.n208 VSS.n207 0.0251575
R1150 VSS.n290 VSS.n289 0.0251575
R1151 VSS.n96 VSS.n95 0.0251575
R1152 VSS.n167 VSS.n164 0.0226918
R1153 VSS.n226 VSS.n220 0.0226918
R1154 VSS.n334 VSS.n333 0.0226918
R1155 VSS.n300 VSS.n298 0.0226918
R1156 VSS.n42 VSS.n40 0.0226918
R1157 VSS.n250 VSS.n249 0.0226918
R1158 VSS.n340 VSS.n339 0.0223939
R1159 VSS.n23 VSS.n22 0.0220753
R1160 VSS.n64 VSS.n62 0.0220753
R1161 VSS.n160 VSS.n159 0.0183767
R1162 VSS.n329 VSS.n328 0.0177603
R1163 VSS.n293 VSS.n292 0.0177603
R1164 VSS.n245 VSS.n244 0.0177603
R1165 VSS.n60 VSS.n59 0.0112717
R1166 VSS.n338 VSS.n140 0.0110653
R1167 VSS.n68 VSS.n67 0.010987
R1168 VSS.n38 VSS.n37 0.010987
R1169 VSS.n25 VSS.n24 0.010987
R1170 VSS.n73 VSS.n72 0.010987
R1171 VSS.n217 VSS.n216 0.010363
R1172 VSS.n296 VSS.n295 0.010363
R1173 VSS.n105 VSS.n104 0.010363
R1174 VSS.n38 VSS.n30 0.00358219
R1175 VSS.n68 VSS.n64 0.00358219
R1176 VSS.n25 VSS.n23 0.00296575
R1177 VSS.n72 VSS.n20 0.00296575
R1178 VSS.n232 VSS.n226 0.00234932
R1179 VSS.n336 VSS.n334 0.00234932
R1180 VSS.n305 VSS.n300 0.00234932
R1181 VSS.n252 VSS.n250 0.00234932
R1182 VSS.n339 VSS.n338 0.00231208
R1183 VSS.n168 VSS.n146 0.00185597
R1184 VSS.n168 VSS.n167 0.00173288
R1185 VSS.n60 VSS.n42 0.00173288
R1186 VSS.n305 VSS.n304 0.00128532
R1187 VSS.n252 VSS.n251 0.00128532
R1188 VSS.n336 VSS.n335 0.00128532
R1189 ITAIL.n52 ITAIL.n51 106.159
R1190 ITAIL.n124 ITAIL.n123 103.823
R1191 ITAIL.n40 ITAIL.n39 103.823
R1192 ITAIL.n23 ITAIL.n22 103.823
R1193 ITAIL.n31 ITAIL.n30 103.823
R1194 ITAIL.n41 ITAIL.n38 103.823
R1195 ITAIL.n87 ITAIL.n86 103.823
R1196 ITAIL.n57 ITAIL.n56 103.823
R1197 ITAIL.n134 ITAIL.n133 103.823
R1198 ITAIL.n139 ITAIL.n138 103.823
R1199 ITAIL.n39 ITAIL.t54 37.2224
R1200 ITAIL.n22 ITAIL.t59 37.2224
R1201 ITAIL.n30 ITAIL.n23 21.0894
R1202 ITAIL.n38 ITAIL.n31 21.0894
R1203 ITAIL.n41 ITAIL.n40 21.0894
R1204 ITAIL.n39 ITAIL.t43 16.1335
R1205 ITAIL.n40 ITAIL.t58 16.1335
R1206 ITAIL.n22 ITAIL.t52 16.1335
R1207 ITAIL.n23 ITAIL.t44 16.1335
R1208 ITAIL.n31 ITAIL.t49 16.1335
R1209 ITAIL.n51 ITAIL.t16 14.0165
R1210 ITAIL.n53 ITAIL.t26 14.0165
R1211 ITAIL.n55 ITAIL.t30 14.0165
R1212 ITAIL.n58 ITAIL.t34 14.0165
R1213 ITAIL.n7 ITAIL.t0 14.0165
R1214 ITAIL.n135 ITAIL.t20 14.0165
R1215 ITAIL.n137 ITAIL.t22 13.9435
R1216 ITAIL.n83 ITAIL.t2 13.7975
R1217 ITAIL.n85 ITAIL.t6 13.7975
R1218 ITAIL.n120 ITAIL.t14 13.7975
R1219 ITAIL.n122 ITAIL.t10 13.7975
R1220 ITAIL.n113 ITAIL.t28 13.7975
R1221 ITAIL.n105 ITAIL.t24 13.7975
R1222 ITAIL.n88 ITAIL.t8 13.7975
R1223 ITAIL.n141 ITAIL.t36 12.7902
R1224 ITAIL.n20 ITAIL.t46 12.7836
R1225 ITAIL.n62 ITAIL.t38 12.7453
R1226 ITAIL.n116 ITAIL.t32 12.5263
R1227 ITAIL.n99 ITAIL.t18 12.4795
R1228 ITAIL.n91 ITAIL.t12 12.4359
R1229 ITAIL.n2 ITAIL.t4 11.6805
R1230 ITAIL.n24 ITAIL.t57 11.5345
R1231 ITAIL.n32 ITAIL.t53 11.4615
R1232 ITAIL.n51 ITAIL.n50 9.23263
R1233 ITAIL.n38 ITAIL.n37 8.0053
R1234 ITAIL.n30 ITAIL.n29 8.0005
R1235 ITAIL.n142 ITAIL.t37 5.20163
R1236 ITAIL.n84 ITAIL.n83 4.15465
R1237 ITAIL.n85 ITAIL.n84 4.15465
R1238 ITAIL.n121 ITAIL.n120 4.15465
R1239 ITAIL.n122 ITAIL.n121 4.15465
R1240 ITAIL.n114 ITAIL.n113 4.15465
R1241 ITAIL.n106 ITAIL.n105 4.15465
R1242 ITAIL.n89 ITAIL.n88 4.15465
R1243 ITAIL.n54 ITAIL.n53 4.15465
R1244 ITAIL.n55 ITAIL.n54 4.15465
R1245 ITAIL.n59 ITAIL.n58 4.15465
R1246 ITAIL.n8 ITAIL.n7 4.15465
R1247 ITAIL.n136 ITAIL.n135 4.15465
R1248 ITAIL.n137 ITAIL.n136 4.15465
R1249 ITAIL.n143 ITAIL.n141 3.51942
R1250 ITAIL.n100 ITAIL.n98 3.50928
R1251 ITAIL.n117 ITAIL.n116 3.50535
R1252 ITAIL.n132 ITAIL.n131 3.50535
R1253 ITAIL.n100 ITAIL.n99 3.49877
R1254 ITAIL.n92 ITAIL.n91 3.47756
R1255 ITAIL.n146 ITAIL.n144 3.46513
R1256 ITAIL.n54 ITAIL.n49 3.43811
R1257 ITAIL.n59 ITAIL.n47 3.43811
R1258 ITAIL.n8 ITAIL.n5 3.43811
R1259 ITAIL.n136 ITAIL.n1 3.43615
R1260 ITAIL.n84 ITAIL.n82 3.43224
R1261 ITAIL.n121 ITAIL.n119 3.43224
R1262 ITAIL.n114 ITAIL.n111 3.43224
R1263 ITAIL.n106 ITAIL.n103 3.43224
R1264 ITAIL.n89 ITAIL.n80 3.43224
R1265 ITAIL.n96 ITAIL.n95 2.90675
R1266 ITAIL.n43 ITAIL.n42 2.88564
R1267 ITAIL.n95 ITAIL.n94 2.88464
R1268 ITAIL.n144 ITAIL.n140 2.88451
R1269 ITAIL.n126 ITAIL.n125 2.88438
R1270 ITAIL.n127 ITAIL.n126 2.87461
R1271 ITAIL.n107 ITAIL.n101 2.8741
R1272 ITAIL.n138 ITAIL.n137 2.4095
R1273 ITAIL.n86 ITAIL.n85 2.3365
R1274 ITAIL.n123 ITAIL.n122 2.3365
R1275 ITAIL.n113 ITAIL.n112 2.3365
R1276 ITAIL.n25 ITAIL.n24 2.3365
R1277 ITAIL.n33 ITAIL.n32 2.3365
R1278 ITAIL.n38 ITAIL.n33 2.3365
R1279 ITAIL.n105 ITAIL.n104 2.3365
R1280 ITAIL.n94 ITAIL.n93 2.3365
R1281 ITAIL.n88 ITAIL.n87 2.3365
R1282 ITAIL.n53 ITAIL.n52 2.3365
R1283 ITAIL.n56 ITAIL.n55 2.3365
R1284 ITAIL.n58 ITAIL.n57 2.3365
R1285 ITAIL.n7 ITAIL.n6 2.3365
R1286 ITAIL.n135 ITAIL.n134 2.3365
R1287 ITAIL.n125 ITAIL.n124 2.2635
R1288 ITAIL.n30 ITAIL.n25 2.2635
R1289 ITAIL.n42 ITAIL.n41 2.2635
R1290 ITAIL.n3 ITAIL.n2 2.2635
R1291 ITAIL.n146 ITAIL.n145 2.2565
R1292 ITAIL.n44 ITAIL.n43 2.2505
R1293 ITAIL.n109 ITAIL.n108 2.2505
R1294 ITAIL.n66 ITAIL.n65 2.2505
R1295 ITAIL.n130 ITAIL.n129 2.2505
R1296 ITAIL.n21 ITAIL.n20 2.22354
R1297 ITAIL.n63 ITAIL.n61 2.1905
R1298 ITAIL.n140 ITAIL.n139 2.1175
R1299 ITAIL.n64 ITAIL.n63 2.11497
R1300 ITAIL.n82 ITAIL.t3 1.6385
R1301 ITAIL.n82 ITAIL.n81 1.6385
R1302 ITAIL.n119 ITAIL.t11 1.6385
R1303 ITAIL.n119 ITAIL.n118 1.6385
R1304 ITAIL.n111 ITAIL.t29 1.6385
R1305 ITAIL.n111 ITAIL.n110 1.6385
R1306 ITAIL.n103 ITAIL.t25 1.6385
R1307 ITAIL.n103 ITAIL.n102 1.6385
R1308 ITAIL.n80 ITAIL.t9 1.6385
R1309 ITAIL.n80 ITAIL.n79 1.6385
R1310 ITAIL.n49 ITAIL.t27 1.6385
R1311 ITAIL.n49 ITAIL.n48 1.6385
R1312 ITAIL.n47 ITAIL.t35 1.6385
R1313 ITAIL.n47 ITAIL.n46 1.6385
R1314 ITAIL.n5 ITAIL.t1 1.6385
R1315 ITAIL.n5 ITAIL.n4 1.6385
R1316 ITAIL.n1 ITAIL.t21 1.6385
R1317 ITAIL.n1 ITAIL.n0 1.6385
R1318 ITAIL.n75 ITAIL.n74 1.54118
R1319 ITAIL.n128 ITAIL.n127 1.22514
R1320 ITAIL.n66 ITAIL.n45 1.20852
R1321 ITAIL.n45 ITAIL.n18 1.12208
R1322 ITAIL.n63 ITAIL.n62 1.06529
R1323 ITAIL.n133 ITAIL.n132 1.06529
R1324 ITAIL.n132 ITAIL.n3 1.06529
R1325 ITAIL.n98 ITAIL.n97 1.02542
R1326 ITAIL.n129 ITAIL.n68 1.01647
R1327 ITAIL.n128 ITAIL.n78 0.807879
R1328 ITAIL.n127 ITAIL.n109 0.652981
R1329 ITAIL.n109 ITAIL.n96 0.604805
R1330 ITAIL.n74 ITAIL.n73 0.558332
R1331 ITAIL.n73 ITAIL.n72 0.543697
R1332 ITAIL.n17 ITAIL.n16 0.526864
R1333 ITAIL.n68 ITAIL.n17 0.255717
R1334 ITAIL.n70 ITAIL.n69 0.249615
R1335 ITAIL.n68 ITAIL.n67 0.246164
R1336 ITAIL.n64 ITAIL.n59 0.147502
R1337 ITAIL.n107 ITAIL.n106 0.141303
R1338 ITAIL.n115 ITAIL.n114 0.124649
R1339 ITAIL.n9 ITAIL.n8 0.123649
R1340 ITAIL.n90 ITAIL.n89 0.122649
R1341 ITAIL.n61 ITAIL.n60 0.0735
R1342 ITAIL.n27 ITAIL.n26 0.0419159
R1343 ITAIL.n37 ITAIL.n34 0.0418237
R1344 ITAIL.n15 ITAIL.n11 0.037926
R1345 ITAIL.n78 ITAIL.n77 0.0329299
R1346 ITAIL.n92 ITAIL.n90 0.0325
R1347 ITAIL.n131 ITAIL.n9 0.0315
R1348 ITAIL.n143 ITAIL.n142 0.0315
R1349 ITAIL.n117 ITAIL.n115 0.0305
R1350 ITAIL.n71 ITAIL.n70 0.0305
R1351 ITAIL.n11 ITAIL.n10 0.0305
R1352 ITAIL.n72 ITAIL.n71 0.0295
R1353 ITAIL.n15 ITAIL.n14 0.024689
R1354 ITAIL.n13 ITAIL.n12 0.0235087
R1355 ITAIL.n67 ITAIL.n66 0.0215938
R1356 ITAIL.n14 ITAIL.n13 0.0178976
R1357 ITAIL.n16 ITAIL.n15 0.0177217
R1358 ITAIL.n108 ITAIL.n107 0.0117741
R1359 ITAIL.n65 ITAIL.n64 0.00955805
R1360 ITAIL.n78 ITAIL.n75 0.00955501
R1361 ITAIL.n45 ITAIL.n44 0.00872297
R1362 ITAIL.n129 ITAIL.n128 0.00692857
R1363 ITAIL ITAIL.n146 0.0065
R1364 ITAIL.n29 ITAIL.n28 0.00579412
R1365 ITAIL.n36 ITAIL.n35 0.00579412
R1366 ITAIL.n77 ITAIL.n76 0.00579412
R1367 ITAIL.n108 ITAIL.n100 0.0035
R1368 ITAIL.n126 ITAIL.n117 0.0025
R1369 ITAIL.n43 ITAIL.n21 0.0025
R1370 ITAIL.n131 ITAIL.n130 0.0025
R1371 ITAIL.n37 ITAIL.n36 0.00163206
R1372 ITAIL.n28 ITAIL.n27 0.00162327
R1373 ITAIL.n44 ITAIL.n19 0.0015
R1374 ITAIL.n95 ITAIL.n92 0.0015
R1375 ITAIL.n144 ITAIL.n143 0.0015
R1376 G_source_dn.n54 G_source_dn.t8 34.3024
R1377 G_source_dn.n39 G_source_dn.t29 31.8591
R1378 G_source_dn.t26 G_source_dn.n44 31.6095
R1379 G_source_dn.n39 G_source_dn.t24 22.4115
R1380 G_source_dn.n40 G_source_dn.t28 22.4115
R1381 G_source_dn.n43 G_source_dn.t30 22.4115
R1382 G_source_dn.n44 G_source_dn.t35 22.4115
R1383 G_source_dn.n40 G_source_dn.n39 18.9805
R1384 G_source_dn.n41 G_source_dn.n40 18.9805
R1385 G_source_dn.n42 G_source_dn.n41 18.9805
R1386 G_source_dn.n43 G_source_dn.n42 18.9805
R1387 G_source_dn.n44 G_source_dn.n43 18.9805
R1388 G_source_dn.n45 G_source_dn.t26 15.4821
R1389 G_source_dn.n41 G_source_dn.t32 12.6295
R1390 G_source_dn.n42 G_source_dn.t34 12.6295
R1391 G_source_dn.n55 G_source_dn.t16 10.8775
R1392 G_source_dn.n52 G_source_dn.t20 10.8775
R1393 G_source_dn.n16 G_source_dn.t14 10.8775
R1394 G_source_dn.n13 G_source_dn.t12 10.8775
R1395 G_source_dn.n10 G_source_dn.t18 10.8775
R1396 G_source_dn.n25 G_source_dn.t10 9.65117
R1397 G_source_dn.n21 G_source_dn.t22 9.65117
R1398 G_source_dn.n34 G_source_dn.n33 6.96833
R1399 G_source_dn.n37 G_source_dn.t6 6.17107
R1400 G_source_dn.n11 G_source_dn.n10 4.15702
R1401 G_source_dn.n14 G_source_dn.n13 4.0005
R1402 G_source_dn.n17 G_source_dn.n16 4.0005
R1403 G_source_dn.n53 G_source_dn.n52 4.0005
R1404 G_source_dn.n56 G_source_dn.n55 4.0005
R1405 G_source_dn.n22 G_source_dn.n21 3.51942
R1406 G_source_dn.n26 G_source_dn.n25 3.51942
R1407 G_source_dn.n36 G_source_dn.n28 3.46159
R1408 G_source_dn.n34 G_source_dn.n32 3.46159
R1409 G_source_dn.n35 G_source_dn.n30 3.44007
R1410 G_source_dn.n38 G_source_dn.n37 3.34436
R1411 G_source_dn.n1 G_source_dn.t17 3.03383
R1412 G_source_dn.n1 G_source_dn.n0 3.03383
R1413 G_source_dn.n9 G_source_dn.t19 3.03383
R1414 G_source_dn.n9 G_source_dn.n8 3.03383
R1415 G_source_dn.n7 G_source_dn.t15 3.03383
R1416 G_source_dn.n7 G_source_dn.n6 3.03383
R1417 G_source_dn.n3 G_source_dn.t11 3.03383
R1418 G_source_dn.n3 G_source_dn.n2 3.03383
R1419 G_source_dn.n19 G_source_dn.n5 2.8741
R1420 G_source_dn.n49 G_source_dn.n48 2.8741
R1421 G_source_dn.n57 G_source_dn.n1 2.80398
R1422 G_source_dn.n11 G_source_dn.n9 2.80398
R1423 G_source_dn.n18 G_source_dn.n7 2.80398
R1424 G_source_dn.n50 G_source_dn.n3 2.80398
R1425 G_source_dn.n30 G_source_dn.t1 2.7305
R1426 G_source_dn.n30 G_source_dn.n29 2.7305
R1427 G_source_dn.n28 G_source_dn.t0 2.7305
R1428 G_source_dn.n28 G_source_dn.n27 2.7305
R1429 G_source_dn.n32 G_source_dn.t4 2.7305
R1430 G_source_dn.n32 G_source_dn.n31 2.7305
R1431 G_source_dn.n55 G_source_dn.n54 2.3365
R1432 G_source_dn.n52 G_source_dn.n51 2.3365
R1433 G_source_dn.n16 G_source_dn.n15 2.3365
R1434 G_source_dn.n13 G_source_dn.n12 2.3365
R1435 G_source_dn.n46 G_source_dn.n45 2.2505
R1436 G_source_dn.n48 G_source_dn.n47 2.1175
R1437 G_source_dn.n5 G_source_dn.n4 2.1175
R1438 G_source_dn.n17 G_source_dn.n14 1.1118
R1439 G_source_dn.n56 G_source_dn.n53 1.1118
R1440 G_source_dn.n24 G_source_dn.n23 1.0508
R1441 G_source_dn.n35 G_source_dn.n34 0.798761
R1442 G_source_dn.n36 G_source_dn.n35 0.798761
R1443 G_source_dn.n37 G_source_dn.n36 0.710717
R1444 G_source_dn.n45 G_source_dn.n38 0.592714
R1445 G_source_dn.n14 G_source_dn.n11 0.157022
R1446 G_source_dn.n18 G_source_dn.n17 0.157022
R1447 G_source_dn.n53 G_source_dn.n50 0.157022
R1448 G_source_dn.n19 G_source_dn.n18 0.143676
R1449 G_source_dn.n50 G_source_dn.n49 0.142676
R1450 G_source_dn.n57 G_source_dn.n56 0.1025
R1451 G_source_dn G_source_dn.n57 0.0434485
R1452 G_source_dn.n23 G_source_dn.n22 0.0315
R1453 G_source_dn.n26 G_source_dn.n24 0.0305
R1454 G_source_dn.n20 G_source_dn.n19 0.0117741
R1455 G_source_dn.n49 G_source_dn.n46 0.0117741
R1456 G_source_dn.n46 G_source_dn.n26 0.0045
R1457 G_source_dn.n22 G_source_dn.n20 0.0035
R1458 A1.n3 A1.n2 3.22739
R1459 A1.n9 A1.n8 3.22703
R1460 A1.n19 A1.n18 3.22692
R1461 A1.n28 A1.t12 3.03383
R1462 A1.n28 A1.n27 3.03383
R1463 A1.n1 A1.t13 3.03383
R1464 A1.n1 A1.n0 3.03383
R1465 A1.n6 A1.t11 3.03383
R1466 A1.n6 A1.n5 3.03383
R1467 A1.n22 A1.t3 3.03383
R1468 A1.n22 A1.n21 3.03383
R1469 A1.n15 A1.t6 3.03383
R1470 A1.n15 A1.n14 3.03383
R1471 A1.n11 A1.n1 2.81935
R1472 A1.n9 A1.t5 2.62488
R1473 A1.n3 A1.t1 2.62459
R1474 A1.n19 A1.t14 2.62411
R1475 A1.n7 A1.n6 2.44998
R1476 A1.n10 A1.n9 2.40501
R1477 A1.n4 A1.n3 2.39877
R1478 A1.n20 A1.n19 2.33972
R1479 A1.n33 A1.n17 2.2443
R1480 A1.n24 A1.n23 1.49465
R1481 A1.n30 A1.n29 1.49465
R1482 A1.n16 A1.n15 1.25784
R1483 A1.n29 A1.n28 1.2574
R1484 A1.n23 A1.n22 1.2574
R1485 A1.n24 A1.n20 0.609831
R1486 A1.n12 A1.n11 0.595697
R1487 A1.n30 A1.n26 0.576036
R1488 A1.n33 A1.n32 0.567771
R1489 A1.n7 A1.n4 0.527868
R1490 A1.n11 A1.n10 0.524711
R1491 A1.n10 A1.n7 0.518395
R1492 A1.n32 A1.n31 0.0273831
R1493 A1.n26 A1.n25 0.0238766
R1494 A1 A1.n33 0.0167392
R1495 A1.n25 A1.n24 0.0160953
R1496 A1.n31 A1.n30 0.0125888
R1497 A1.n16 A1.n13 0.00188827
R1498 A1 A1.n12 0.00166883
R1499 A1.n17 A1.n16 0.00128036
R1500 ITAIL_SRC.n7 ITAIL_SRC.n6 6.40267
R1501 ITAIL_SRC.n10 ITAIL_SRC.t4 6.02318
R1502 ITAIL_SRC.n5 ITAIL_SRC.t0 3.03383
R1503 ITAIL_SRC.n5 ITAIL_SRC.n4 3.03383
R1504 ITAIL_SRC.n1 ITAIL_SRC.t5 3.03383
R1505 ITAIL_SRC.n1 ITAIL_SRC.n0 3.03383
R1506 ITAIL_SRC.n3 ITAIL_SRC.t1 3.03383
R1507 ITAIL_SRC.n3 ITAIL_SRC.n2 3.03383
R1508 ITAIL_SRC.n8 ITAIL_SRC.n3 2.98985
R1509 ITAIL_SRC.n9 ITAIL_SRC.n1 2.9605
R1510 ITAIL_SRC.n7 ITAIL_SRC.n5 2.95975
R1511 ITAIL_SRC.n9 ITAIL_SRC.n8 0.379057
R1512 ITAIL_SRC.n10 ITAIL_SRC.n9 0.379057
R1513 ITAIL_SRC.n8 ITAIL_SRC.n7 0.378129
R1514 ITAIL_SRC ITAIL_SRC.n10 0.256582
R1515 G1_1.n5 G1_1.n2 103.823
R1516 G1_1.n54 G1_1.n53 103.823
R1517 G1_1.n4 G1_1.n3 103.823
R1518 G1_1.n55 G1_1.n52 103.823
R1519 G1_1.n2 G1_1.t77 32.8424
R1520 G1_1.n53 G1_1.t74 32.8424
R1521 G1_1.n117 G1_1.t12 31.6661
R1522 G1_1.n33 G1_1.t22 31.5165
R1523 G1_1.n5 G1_1.n4 21.0894
R1524 G1_1.n55 G1_1.n54 21.0894
R1525 G1_1.n116 G1_1.t18 15.4035
R1526 G1_1.n117 G1_1.t4 15.4035
R1527 G1_1.n69 G1_1.t16 15.1845
R1528 G1_1.n70 G1_1.t20 15.1845
R1529 G1_1.n33 G1_1.t14 15.0385
R1530 G1_1.n34 G1_1.t38 15.0385
R1531 G1_1.n79 G1_1.t8 15.0385
R1532 G1_1.n81 G1_1.t32 15.0385
R1533 G1_1.n45 G1_1.t6 14.8925
R1534 G1_1.n47 G1_1.t30 14.8925
R1535 G1_1.n65 G1_1.t24 12.0455
R1536 G1_1.n64 G1_1.t36 12.0455
R1537 G1_1.n89 G1_1.t26 11.9725
R1538 G1_1.n88 G1_1.t0 11.9725
R1539 G1_1.n39 G1_1.t34 11.8995
R1540 G1_1.n38 G1_1.t10 11.8995
R1541 G1_1.n2 G1_1.t71 11.7535
R1542 G1_1.n53 G1_1.t60 11.7535
R1543 G1_1.n54 G1_1.t76 11.7535
R1544 G1_1.n4 G1_1.t75 11.7535
R1545 G1_1.n3 G1_1.t68 11.7535
R1546 G1_1.n52 G1_1.t73 11.7535
R1547 G1_1.n74 G1_1.t2 11.6805
R1548 G1_1.n73 G1_1.t28 11.6805
R1549 G1_1.n57 G1_1.t63 8.14629
R1550 G1_1.n0 G1_1.t62 8.14629
R1551 G1_1.n5 G1_1.n1 8.0005
R1552 G1_1.n118 G1_1.n116 7.97643
R1553 G1_1.n66 G1_1.n64 7.49604
R1554 G1_1.n35 G1_1.n34 7.2359
R1555 G1_1.n90 G1_1.n88 6.91289
R1556 G1_1.n71 G1_1.n69 6.84014
R1557 G1_1.n75 G1_1.n74 6.80135
R1558 G1_1.n40 G1_1.n39 6.66015
R1559 G1_1.n71 G1_1.n70 6.57708
R1560 G1_1.n40 G1_1.n38 6.40401
R1561 G1_1.n90 G1_1.n89 6.26687
R1562 G1_1.n35 G1_1.n33 5.94386
R1563 G1_1.n75 G1_1.n73 5.92785
R1564 G1_1.n61 G1_1.n60 5.92398
R1565 G1_1.n125 G1_1.n124 5.90903
R1566 G1_1.n118 G1_1.n117 5.81346
R1567 G1_1.n66 G1_1.n65 5.80139
R1568 G1_1.n30 G1_1.n23 5.1485
R1569 G1_1.n114 G1_1.t54 5.1485
R1570 G1_1.n32 G1_1.n31 4.4205
R1571 G1_1.n115 G1_1.t13 4.4205
R1572 G1_1.n46 G1_1.n45 4.19007
R1573 G1_1.n80 G1_1.n79 4.07041
R1574 G1_1.n82 G1_1.n81 4.07041
R1575 G1_1.n121 G1_1.n90 4.0005
R1576 G1_1.n119 G1_1.n118 4.0005
R1577 G1_1.n36 G1_1.n35 4.0005
R1578 G1_1.n41 G1_1.n40 4.0005
R1579 G1_1.n67 G1_1.n66 4.0005
R1580 G1_1.n72 G1_1.n71 4.0005
R1581 G1_1.n76 G1_1.n75 4.0005
R1582 G1_1.n48 G1_1.n47 3.8092
R1583 G1_1.n113 G1_1.n94 3.54572
R1584 G1_1.n111 G1_1.n98 3.54572
R1585 G1_1.n109 G1_1.n102 3.54572
R1586 G1_1.n107 G1_1.n106 3.54572
R1587 G1_1.n29 G1_1.n25 3.54572
R1588 G1_1.n58 G1_1.n56 3.53093
R1589 G1_1.n28 G1_1.n27 3.5105
R1590 G1_1.n108 G1_1.n104 3.5105
R1591 G1_1.n110 G1_1.n100 3.5105
R1592 G1_1.n112 G1_1.n96 3.5105
R1593 G1_1.n58 G1_1.n57 3.50535
R1594 G1_1.n1 G1_1.n0 3.50535
R1595 G1_1.n120 G1_1.n92 3.02311
R1596 G1_1.n68 G1_1.n14 3.01724
R1597 G1_1.n124 G1_1.n10 3.01333
R1598 G1_1.n37 G1_1.n22 3.01333
R1599 G1_1.n44 G1_1.n18 3.00941
R1600 G1_1.n63 G1_1.n16 2.93311
R1601 G1_1.n122 G1_1.n87 2.93115
R1602 G1_1.n42 G1_1.n20 2.9292
R1603 G1_1.n77 G1_1.n12 2.92333
R1604 G1_1.n8 G1_1.n7 2.88455
R1605 G1_1.n60 G1_1.n59 2.88451
R1606 G1_1.n51 G1_1.n50 2.66717
R1607 G1_1.n85 G1_1.n84 2.66717
R1608 G1_1.n83 G1_1.n82 2.51997
R1609 G1_1.n84 G1_1.n80 2.45537
R1610 G1_1.n32 G1_1.n30 2.44296
R1611 G1_1.n50 G1_1.n46 2.41267
R1612 G1_1.n49 G1_1.n48 2.41267
R1613 G1_1.n115 G1_1.n114 2.14942
R1614 G1_1.n6 G1_1.n5 1.9715
R1615 G1_1.n10 G1_1.t9 1.8205
R1616 G1_1.n10 G1_1.n9 1.8205
R1617 G1_1.n87 G1_1.t1 1.8205
R1618 G1_1.n87 G1_1.n86 1.8205
R1619 G1_1.n92 G1_1.t19 1.8205
R1620 G1_1.n92 G1_1.n91 1.8205
R1621 G1_1.n22 G1_1.t15 1.8205
R1622 G1_1.n22 G1_1.n21 1.8205
R1623 G1_1.n20 G1_1.t11 1.8205
R1624 G1_1.n20 G1_1.n19 1.8205
R1625 G1_1.n18 G1_1.t7 1.8205
R1626 G1_1.n18 G1_1.n17 1.8205
R1627 G1_1.n16 G1_1.t37 1.8205
R1628 G1_1.n16 G1_1.n15 1.8205
R1629 G1_1.n14 G1_1.t17 1.8205
R1630 G1_1.n14 G1_1.n13 1.8205
R1631 G1_1.n12 G1_1.t29 1.8205
R1632 G1_1.n12 G1_1.n11 1.8205
R1633 G1_1.n27 G1_1.t53 1.6385
R1634 G1_1.n27 G1_1.n26 1.6385
R1635 G1_1.n104 G1_1.t59 1.6385
R1636 G1_1.n104 G1_1.n103 1.6385
R1637 G1_1.n100 G1_1.t58 1.6385
R1638 G1_1.n100 G1_1.n99 1.6385
R1639 G1_1.n96 G1_1.t50 1.6385
R1640 G1_1.n96 G1_1.n95 1.6385
R1641 G1_1.n94 G1_1.t57 1.6385
R1642 G1_1.n94 G1_1.n93 1.6385
R1643 G1_1.n98 G1_1.t52 1.6385
R1644 G1_1.n98 G1_1.n97 1.6385
R1645 G1_1.n102 G1_1.t56 1.6385
R1646 G1_1.n102 G1_1.n101 1.6385
R1647 G1_1.n106 G1_1.t51 1.6385
R1648 G1_1.n106 G1_1.n105 1.6385
R1649 G1_1.n25 G1_1.t55 1.6385
R1650 G1_1.n25 G1_1.n24 1.6385
R1651 G1_1.n119 G1_1.n115 1.14702
R1652 G1_1.n36 G1_1.n32 1.14051
R1653 G1_1.n56 G1_1.n55 0.995675
R1654 G1_1.n121 G1_1.n120 0.692144
R1655 G1_1.n41 G1_1.n37 0.686551
R1656 G1_1.n68 G1_1.n67 0.660185
R1657 G1_1.n76 G1_1.n72 0.659391
R1658 G1_1.n63 G1_1.n62 0.656587
R1659 G1_1.n123 G1_1.n122 0.651709
R1660 G1_1.n43 G1_1.n42 0.651372
R1661 G1_1.n78 G1_1.n77 0.648302
R1662 G1_1.n30 G1_1.n29 0.565423
R1663 G1_1.n29 G1_1.n28 0.565423
R1664 G1_1.n108 G1_1.n107 0.565423
R1665 G1_1.n109 G1_1.n108 0.565423
R1666 G1_1.n110 G1_1.n109 0.565423
R1667 G1_1.n111 G1_1.n110 0.565423
R1668 G1_1.n112 G1_1.n111 0.565423
R1669 G1_1.n113 G1_1.n112 0.565423
R1670 G1_1.n114 G1_1.n113 0.565423
R1671 G1_1.n7 G1_1.n6 0.3655
R1672 G1_1.n50 G1_1.n49 0.127457
R1673 G1_1.n84 G1_1.n83 0.0651018
R1674 G1_1.n124 G1_1.n123 0.0345777
R1675 G1_1.n85 G1_1.n78 0.0337039
R1676 G1_1.n62 G1_1.n61 0.0330714
R1677 G1_1.n44 G1_1.n43 0.0313571
R1678 G1_1.n120 G1_1.n119 0.0151939
R1679 G1_1.n67 G1_1.n63 0.0106739
R1680 G1_1.n37 G1_1.n36 0.00923786
R1681 G1_1.n77 G1_1.n76 0.00575
R1682 G1_1 G1_1.n125 0.0055
R1683 G1_1.n122 G1_1.n121 0.00437931
R1684 G1_1.n60 G1_1.n58 0.0025
R1685 G1_1.n72 G1_1.n68 0.00228218
R1686 G1_1.n8 G1_1.n1 0.00228158
R1687 G1_1.n51 G1_1.n44 0.00221429
R1688 G1_1.n61 G1_1.n51 0.00221429
R1689 G1_1.n42 G1_1.n41 0.00203846
R1690 G1_1.n125 G1_1.n8 0.0017181
R1691 G1_1.n124 G1_1.n85 0.00137379
R1692 G_sink_up.n29 G_sink_up.n19 143.595
R1693 G_sink_up.n26 G_sink_up.n22 132.008
R1694 G_sink_up.n0 G_sink_up.t32 116.525
R1695 G_sink_up.n56 G_sink_up.n51 106.903
R1696 G_sink_up.n2 G_sink_up.n1 103.823
R1697 G_sink_up.n6 G_sink_up.n5 103.823
R1698 G_sink_up.n21 G_sink_up.n20 103.823
R1699 G_sink_up.n28 G_sink_up.n27 103.823
R1700 G_sink_up.n18 G_sink_up.n17 95.8364
R1701 G_sink_up.n55 G_sink_up.n54 94.1889
R1702 G_sink_up.n52 G_sink_up.t43 84.6824
R1703 G_sink_up.n54 G_sink_up.n53 70.5213
R1704 G_sink_up.n5 G_sink_up.n2 49.2755
R1705 G_sink_up.n20 G_sink_up.t30 33.7914
R1706 G_sink_up.n17 G_sink_up.t28 32.6802
R1707 G_sink_up.n29 G_sink_up.n28 30.4172
R1708 G_sink_up.n1 G_sink_up.n0 21.0894
R1709 G_sink_up.n51 G_sink_up.n6 21.0894
R1710 G_sink_up.n22 G_sink_up.n21 21.0894
R1711 G_sink_up.n27 G_sink_up.n26 21.0894
R1712 G_sink_up.n19 G_sink_up.n18 19.4672
R1713 G_sink_up.n53 G_sink_up.n52 14.325
R1714 G_sink_up.n52 G_sink_up.t27 13.9435
R1715 G_sink_up.n53 G_sink_up.t36 13.9435
R1716 G_sink_up.n54 G_sink_up.t37 13.9435
R1717 G_sink_up.n17 G_sink_up.t33 13.2135
R1718 G_sink_up.n18 G_sink_up.t38 13.2135
R1719 G_sink_up.n19 G_sink_up.t26 13.2135
R1720 G_sink_up.n0 G_sink_up.t34 12.7025
R1721 G_sink_up.n1 G_sink_up.t35 12.7025
R1722 G_sink_up.n2 G_sink_up.t42 12.7025
R1723 G_sink_up.n6 G_sink_up.t14 12.7025
R1724 G_sink_up.n20 G_sink_up.t40 12.7025
R1725 G_sink_up.n21 G_sink_up.t39 12.7025
R1726 G_sink_up.n22 G_sink_up.t44 12.7025
R1727 G_sink_up.n27 G_sink_up.t12 12.7025
R1728 G_sink_up.n28 G_sink_up.t20 12.7025
R1729 G_sink_up.n4 G_sink_up.t10 10.3665
R1730 G_sink_up.n25 G_sink_up.t16 10.3665
R1731 G_sink_up.n4 G_sink_up.n3 10.2268
R1732 G_sink_up.n55 G_sink_up.t18 9.1985
R1733 G_sink_up.n15 G_sink_up.t22 9.14017
R1734 G_sink_up.n7 G_sink_up.t24 7.9575
R1735 G_sink_up.n25 G_sink_up.n24 7.48719
R1736 G_sink_up.n57 G_sink_up.t19 6.05659
R1737 G_sink_up.n34 G_sink_up.t2 4.5505
R1738 G_sink_up.n34 G_sink_up.n33 4.5505
R1739 G_sink_up.n36 G_sink_up.t4 4.5505
R1740 G_sink_up.n36 G_sink_up.n35 4.5505
R1741 G_sink_up.n38 G_sink_up.t1 4.5505
R1742 G_sink_up.n38 G_sink_up.n37 4.5505
R1743 G_sink_up.n40 G_sink_up.t3 4.5505
R1744 G_sink_up.n40 G_sink_up.n39 4.5505
R1745 G_sink_up.n45 G_sink_up.t5 4.5505
R1746 G_sink_up.n45 G_sink_up.n44 4.5505
R1747 G_sink_up.n48 G_sink_up.n47 4.36782
R1748 G_sink_up.n57 G_sink_up.n56 4.13903
R1749 G_sink_up.n47 G_sink_up.n46 4.11987
R1750 G_sink_up.n41 G_sink_up.n40 3.98849
R1751 G_sink_up.n16 G_sink_up.n15 3.51942
R1752 G_sink_up.n50 G_sink_up.n49 3.50535
R1753 G_sink_up.n14 G_sink_up.n13 3.47497
R1754 G_sink_up.n11 G_sink_up.n10 3.45688
R1755 G_sink_up.n32 G_sink_up.n31 2.88447
R1756 G_sink_up.n43 G_sink_up.n34 2.80398
R1757 G_sink_up.n42 G_sink_up.n36 2.80398
R1758 G_sink_up.n41 G_sink_up.n38 2.80398
R1759 G_sink_up.n46 G_sink_up.n45 2.78907
R1760 G_sink_up.n24 G_sink_up.t17 2.7305
R1761 G_sink_up.n24 G_sink_up.n23 2.7305
R1762 G_sink_up.n13 G_sink_up.t21 2.7305
R1763 G_sink_up.n13 G_sink_up.n12 2.7305
R1764 G_sink_up.n10 G_sink_up.t15 2.7305
R1765 G_sink_up.n10 G_sink_up.n9 2.7305
R1766 G_sink_up.n56 G_sink_up.n55 2.39581
R1767 G_sink_up.n5 G_sink_up.n4 2.3365
R1768 G_sink_up.n26 G_sink_up.n25 2.3365
R1769 G_sink_up.n8 G_sink_up.n7 2.2635
R1770 G_sink_up.n47 G_sink_up.n32 2.2505
R1771 G_sink_up.n31 G_sink_up.n30 2.1905
R1772 G_sink_up.n42 G_sink_up.n41 1.18502
R1773 G_sink_up.n43 G_sink_up.n42 1.18502
R1774 G_sink_up.n46 G_sink_up.n43 1.1582
R1775 G_sink_up.n50 G_sink_up.n8 1.13829
R1776 G_sink_up.n51 G_sink_up.n50 1.06529
R1777 G_sink_up.n30 G_sink_up.n29 0.8035
R1778 G_sink_up G_sink_up.n57 0.1805
R1779 G_sink_up.n49 G_sink_up.n11 0.0315
R1780 G_sink_up.n16 G_sink_up.n14 0.0311818
R1781 G_sink_up.n32 G_sink_up.n16 0.00356818
R1782 G_sink_up.n49 G_sink_up.n48 0.0035
R1783 G_sink_dn.n11 G_sink_dn.n10 56.0573
R1784 G_sink_dn.n19 G_sink_dn.n18 49.2755
R1785 G_sink_dn.n12 G_sink_dn.t24 33.7914
R1786 G_sink_dn.n4 G_sink_dn.t38 31.8591
R1787 G_sink_dn.n43 G_sink_dn.n11 23.8634
R1788 G_sink_dn.n13 G_sink_dn.n12 21.0894
R1789 G_sink_dn.n14 G_sink_dn.n13 21.0894
R1790 G_sink_dn.n15 G_sink_dn.n14 21.0894
R1791 G_sink_dn.n16 G_sink_dn.n15 21.0894
R1792 G_sink_dn.n17 G_sink_dn.n16 21.0894
R1793 G_sink_dn.n18 G_sink_dn.n17 21.0894
R1794 G_sink_dn.n26 G_sink_dn.n19 21.0894
R1795 G_sink_dn.n33 G_sink_dn.n26 21.0894
R1796 G_sink_dn.n34 G_sink_dn.n33 21.0894
R1797 G_sink_dn.n35 G_sink_dn.n34 21.0894
R1798 G_sink_dn.n42 G_sink_dn.n35 21.0894
R1799 G_sink_dn.n43 G_sink_dn.n42 21.0894
R1800 G_sink_dn.n10 G_sink_dn.n9 20.5135
R1801 G_sink_dn.n5 G_sink_dn.n4 18.9805
R1802 G_sink_dn.n6 G_sink_dn.n5 18.9805
R1803 G_sink_dn.n7 G_sink_dn.n6 18.9805
R1804 G_sink_dn.n8 G_sink_dn.n7 18.9805
R1805 G_sink_dn.n9 G_sink_dn.n8 18.9805
R1806 G_sink_dn.n12 G_sink_dn.t39 13.0675
R1807 G_sink_dn.n13 G_sink_dn.t28 13.0675
R1808 G_sink_dn.n16 G_sink_dn.t26 13.0675
R1809 G_sink_dn.n17 G_sink_dn.t30 13.0675
R1810 G_sink_dn.n14 G_sink_dn.t25 12.7025
R1811 G_sink_dn.n15 G_sink_dn.t29 12.7025
R1812 G_sink_dn.n18 G_sink_dn.t35 12.7025
R1813 G_sink_dn.n19 G_sink_dn.t10 12.7025
R1814 G_sink_dn.n34 G_sink_dn.t22 12.7025
R1815 G_sink_dn.n35 G_sink_dn.t16 12.7025
R1816 G_sink_dn.n4 G_sink_dn.t34 12.6295
R1817 G_sink_dn.n5 G_sink_dn.t37 12.6295
R1818 G_sink_dn.n6 G_sink_dn.t43 12.6295
R1819 G_sink_dn.n7 G_sink_dn.t32 12.6295
R1820 G_sink_dn.n8 G_sink_dn.t41 12.6295
R1821 G_sink_dn.n9 G_sink_dn.t31 12.6295
R1822 G_sink_dn.n10 G_sink_dn.t33 11.0965
R1823 G_sink_dn.n41 G_sink_dn.t18 10.9505
R1824 G_sink_dn.n44 G_sink_dn.t12 10.9505
R1825 G_sink_dn.n25 G_sink_dn.t14 10.7315
R1826 G_sink_dn.n32 G_sink_dn.t20 10.7315
R1827 G_sink_dn.n11 G_sink_dn.t8 9.9285
R1828 G_sink_dn.n25 G_sink_dn.n24 4.1025
R1829 G_sink_dn.n32 G_sink_dn.n31 4.1025
R1830 G_sink_dn.n41 G_sink_dn.n40 4.09824
R1831 G_sink_dn.n45 G_sink_dn.n44 4.09446
R1832 G_sink_dn.n24 G_sink_dn.n23 3.4655
R1833 G_sink_dn.n31 G_sink_dn.n30 3.4655
R1834 G_sink_dn.n45 G_sink_dn.n3 3.4655
R1835 G_sink_dn.n40 G_sink_dn.n39 3.45572
R1836 G_sink_dn.n40 G_sink_dn.n37 3.35398
R1837 G_sink_dn.n24 G_sink_dn.n21 3.35007
R1838 G_sink_dn.n31 G_sink_dn.n28 3.35007
R1839 G_sink_dn.n45 G_sink_dn.n1 3.34811
R1840 G_sink_dn.n23 G_sink_dn.t11 2.7305
R1841 G_sink_dn.n23 G_sink_dn.n22 2.7305
R1842 G_sink_dn.n21 G_sink_dn.t6 2.7305
R1843 G_sink_dn.n21 G_sink_dn.n20 2.7305
R1844 G_sink_dn.n30 G_sink_dn.t1 2.7305
R1845 G_sink_dn.n30 G_sink_dn.n29 2.7305
R1846 G_sink_dn.n28 G_sink_dn.t21 2.7305
R1847 G_sink_dn.n28 G_sink_dn.n27 2.7305
R1848 G_sink_dn.n39 G_sink_dn.t17 2.7305
R1849 G_sink_dn.n39 G_sink_dn.n38 2.7305
R1850 G_sink_dn.n37 G_sink_dn.t0 2.7305
R1851 G_sink_dn.n37 G_sink_dn.n36 2.7305
R1852 G_sink_dn.n3 G_sink_dn.t3 2.7305
R1853 G_sink_dn.n3 G_sink_dn.n2 2.7305
R1854 G_sink_dn.n1 G_sink_dn.t13 2.7305
R1855 G_sink_dn.n1 G_sink_dn.n0 2.7305
R1856 G_sink_dn.n26 G_sink_dn.n25 2.3365
R1857 G_sink_dn.n33 G_sink_dn.n32 2.3365
R1858 G_sink_dn.n42 G_sink_dn.n41 2.1175
R1859 G_sink_dn.n44 G_sink_dn.n43 2.1175
R1860 G_sink_dn G_sink_dn.n45 0.495747
R1861 SD0_1.n18 SD0_1.n3 3.41579
R1862 SD0_1.n13 SD0_1.n10 3.00682
R1863 SD0_1.n24 SD0_1.n1 3.0043
R1864 SD0_1.n15 SD0_1.n5 3.00256
R1865 SD0_1.n27 SD0_1.t10 2.7305
R1866 SD0_1.n27 SD0_1.n26 2.7305
R1867 SD0_1.n3 SD0_1.t11 2.7305
R1868 SD0_1.n3 SD0_1.n2 2.7305
R1869 SD0_1.n20 SD0_1.t4 2.7305
R1870 SD0_1.n20 SD0_1.n19 2.7305
R1871 SD0_1.n7 SD0_1.t12 2.7305
R1872 SD0_1.n7 SD0_1.n6 2.7305
R1873 SD0_1.n12 SD0_1.t6 2.7305
R1874 SD0_1.n12 SD0_1.n11 2.7305
R1875 SD0_1.n10 SD0_1.t15 2.7305
R1876 SD0_1.n10 SD0_1.n9 2.7305
R1877 SD0_1.n5 SD0_1.t2 2.7305
R1878 SD0_1.n5 SD0_1.n4 2.7305
R1879 SD0_1.n1 SD0_1.t0 2.7305
R1880 SD0_1.n1 SD0_1.n0 2.7305
R1881 SD0_1.n13 SD0_1.n12 2.56463
R1882 SD0_1.n22 SD0_1.n21 2.24419
R1883 SD0_1 SD0_1.n29 1.50504
R1884 SD0_1.n14 SD0_1.n8 1.4943
R1885 SD0_1.n8 SD0_1.n7 1.43801
R1886 SD0_1.n28 SD0_1.n27 1.43776
R1887 SD0_1.n21 SD0_1.n20 1.43749
R1888 SD0_1.n14 SD0_1.n13 0.603471
R1889 SD0_1.n23 SD0_1.n22 0.57715
R1890 SD0_1.n17 SD0_1.n16 0.576682
R1891 SD0_1.n16 SD0_1.n15 0.0255633
R1892 SD0_1.n24 SD0_1.n23 0.0244241
R1893 SD0_1.n18 SD0_1.n17 0.0180472
R1894 SD0_1.n22 SD0_1.n18 0.0146295
R1895 SD0_1.n15 SD0_1.n14 0.0145334
R1896 SD0_1 SD0_1.n24 0.00391772
R1897 SD0_1.n28 SD0_1.n25 0.00358243
R1898 SD0_1.n29 SD0_1.n28 0.00181665
R1899 SD2_1.n68 SD2_1.n1 3.5764
R1900 SD2_1.n26 SD2_1.n25 3.18472
R1901 SD2_1.n30 SD2_1.n17 3.17597
R1902 SD2_1.n39 SD2_1.n15 3.17588
R1903 SD2_1.n41 SD2_1.n13 3.17454
R1904 SD2_1.n44 SD2_1.n9 3.17453
R1905 SD2_1.n56 SD2_1.n5 3.1741
R1906 SD2_1.n27 SD2_1.n21 3.17375
R1907 SD2_1.n72 SD2_1.n69 3.17335
R1908 SD2_1.n50 SD2_1.n7 3.17318
R1909 SD2_1.n65 SD2_1.n3 3.17219
R1910 SD2_1.n74 SD2_1.n73 3.01386
R1911 SD2_1.n42 SD2_1.n11 2.93559
R1912 SD2_1.n26 SD2_1.n23 2.56337
R1913 SD2_1.n28 SD2_1.n19 2.56302
R1914 SD2_1.n75 SD2_1.n74 2.25469
R1915 SD2_1.n64 SD2_1.n63 2.24989
R1916 SD2_1.n38 SD2_1.n37 2.24988
R1917 SD2_1.n34 SD2_1.n33 2.24511
R1918 SD2_1.n48 SD2_1.n47 2.24483
R1919 SD2_1.n60 SD2_1.n59 2.24483
R1920 SD2_1.n54 SD2_1.n53 2.24455
R1921 SD2_1.n62 SD2_1.n61 1.74882
R1922 SD2_1.n58 SD2_1.n57 1.74881
R1923 SD2_1.n46 SD2_1.n45 1.74881
R1924 SD2_1.n36 SD2_1.n35 1.74881
R1925 SD2_1.n19 SD2_1.n18 1.74881
R1926 SD2_1.n32 SD2_1.n31 1.73459
R1927 SD2_1.n52 SD2_1.t1 1.6385
R1928 SD2_1.n52 SD2_1.n51 1.6385
R1929 SD2_1.n11 SD2_1.t12 1.6385
R1930 SD2_1.n11 SD2_1.n10 1.6385
R1931 SD2_1.n23 SD2_1.t11 1.6385
R1932 SD2_1.n23 SD2_1.n22 1.6385
R1933 SD2_1.n25 SD2_1.t34 1.6385
R1934 SD2_1.n25 SD2_1.n24 1.6385
R1935 SD2_1.n21 SD2_1.t19 1.6385
R1936 SD2_1.n21 SD2_1.n20 1.6385
R1937 SD2_1.n17 SD2_1.t22 1.6385
R1938 SD2_1.n17 SD2_1.n16 1.6385
R1939 SD2_1.n15 SD2_1.t15 1.6385
R1940 SD2_1.n15 SD2_1.n14 1.6385
R1941 SD2_1.n13 SD2_1.t36 1.6385
R1942 SD2_1.n13 SD2_1.n12 1.6385
R1943 SD2_1.n9 SD2_1.t10 1.6385
R1944 SD2_1.n9 SD2_1.n8 1.6385
R1945 SD2_1.n7 SD2_1.t28 1.6385
R1946 SD2_1.n7 SD2_1.n6 1.6385
R1947 SD2_1.n5 SD2_1.t16 1.6385
R1948 SD2_1.n5 SD2_1.n4 1.6385
R1949 SD2_1.n3 SD2_1.t37 1.6385
R1950 SD2_1.n3 SD2_1.n2 1.6385
R1951 SD2_1.n1 SD2_1.t2 1.6385
R1952 SD2_1.n1 SD2_1.n0 1.6385
R1953 SD2_1.n71 SD2_1.n70 1.5755
R1954 SD2_1.n32 SD2_1.t17 1.48949
R1955 SD2_1.n58 SD2_1.t26 1.47237
R1956 SD2_1.n46 SD2_1.t23 1.47237
R1957 SD2_1.n36 SD2_1.t25 1.47237
R1958 SD2_1.n19 SD2_1.t29 1.47237
R1959 SD2_1.n62 SD2_1.t13 1.47236
R1960 SD2_1.n53 SD2_1.n52 1.44171
R1961 SD2_1.n73 SD2_1.t32 1.28985
R1962 SD2_1.n63 SD2_1.n62 1.07211
R1963 SD2_1.n37 SD2_1.n36 1.07199
R1964 SD2_1.n47 SD2_1.n46 1.07199
R1965 SD2_1.n59 SD2_1.n58 1.07199
R1966 SD2_1.n33 SD2_1.n32 1.07053
R1967 SD2_1.n29 SD2_1.n28 0.626751
R1968 SD2_1.n27 SD2_1.n26 0.622777
R1969 SD2_1.n43 SD2_1.n42 0.612573
R1970 SD2_1.n55 SD2_1.n54 0.606132
R1971 SD2_1.n64 SD2_1.n60 0.605265
R1972 SD2_1.n38 SD2_1.n34 0.603102
R1973 SD2_1.n49 SD2_1.n48 0.601395
R1974 SD2_1.n67 SD2_1.n66 0.593475
R1975 SD2_1.n41 SD2_1.n40 0.584536
R1976 SD2_1.n73 SD2_1.n72 0.31735
R1977 SD2_1.n72 SD2_1.n71 0.0635
R1978 SD2_1.n28 SD2_1.n27 0.0264198
R1979 SD2_1.n66 SD2_1.n65 0.0249444
R1980 SD2_1.n40 SD2_1.n39 0.024125
R1981 SD2_1.n42 SD2_1.n41 0.0174125
R1982 SD2_1.n34 SD2_1.n30 0.0172816
R1983 SD2_1.n48 SD2_1.n44 0.0167161
R1984 SD2_1.n54 SD2_1.n50 0.0161504
R1985 SD2_1.n60 SD2_1.n56 0.0144661
R1986 SD2_1.n68 SD2_1.n67 0.0061962
R1987 SD2_1.n39 SD2_1.n38 0.00549888
R1988 SD2_1.n74 SD2_1.n69 0.00543151
R1989 SD2_1.n56 SD2_1.n55 0.005
R1990 SD2_1.n75 SD2_1.n68 0.00441168
R1991 SD2_1.n65 SD2_1.n64 0.00433224
R1992 SD2_1 SD2_1.n75 0.00328222
R1993 SD2_1.n30 SD2_1.n29 0.00275
R1994 SD2_1.n44 SD2_1.n43 0.00275
R1995 SD2_1.n50 SD2_1.n49 0.00275
R1996 ITAIL_SINK.n7 ITAIL_SINK.n6 6.67289
R1997 ITAIL_SINK.n10 ITAIL_SINK.t2 6.13289
R1998 ITAIL_SINK.n9 ITAIL_SINK.n1 3.44202
R1999 ITAIL_SINK.n7 ITAIL_SINK.n5 3.44202
R2000 ITAIL_SINK.n8 ITAIL_SINK.n3 3.40289
R2001 ITAIL_SINK.n3 ITAIL_SINK.t3 2.7305
R2002 ITAIL_SINK.n3 ITAIL_SINK.n2 2.7305
R2003 ITAIL_SINK.n1 ITAIL_SINK.t4 2.7305
R2004 ITAIL_SINK.n1 ITAIL_SINK.n0 2.7305
R2005 ITAIL_SINK.n5 ITAIL_SINK.t5 2.7305
R2006 ITAIL_SINK.n5 ITAIL_SINK.n4 2.7305
R2007 ITAIL_SINK.n8 ITAIL_SINK.n7 0.5405
R2008 ITAIL_SINK.n9 ITAIL_SINK.n8 0.5405
R2009 ITAIL_SINK.n10 ITAIL_SINK.n9 0.5405
R2010 ITAIL_SINK ITAIL_SINK.n10 0.192412
R2011 A2.n2 A2.t13 2.7305
R2012 A2.n2 A2.n1 2.7305
R2013 A2.n27 A2.t1 2.7305
R2014 A2.n27 A2.n26 2.7305
R2015 A2.n22 A2.t9 2.7305
R2016 A2.n22 A2.n21 2.7305
R2017 A2.n16 A2.t6 2.7305
R2018 A2.n16 A2.n15 2.7305
R2019 A2.n8 A2.t8 2.7305
R2020 A2.n8 A2.n7 2.7305
R2021 A2.n13 A2.t12 2.7305
R2022 A2.n13 A2.n12 2.7305
R2023 A2.n5 A2.t5 2.7305
R2024 A2.n5 A2.n4 2.7305
R2025 A2.n36 A2.t2 2.7305
R2026 A2.n36 A2.n35 2.7305
R2027 A2.n3 A2.n2 2.56155
R2028 A2.n6 A2.n5 2.56046
R2029 A2.n14 A2.n13 2.55979
R2030 A2 A2.n39 1.50412
R2031 A2.n24 A2.n23 1.49465
R2032 A2.n29 A2.n28 1.49465
R2033 A2.n10 A2.n9 1.49453
R2034 A2.n18 A2.n17 1.49453
R2035 A2.n28 A2.n27 1.43782
R2036 A2.n9 A2.n8 1.43782
R2037 A2.n23 A2.n22 1.43764
R2038 A2.n17 A2.n16 1.43764
R2039 A2.n38 A2.n36 1.43655
R2040 A2.n10 A2.n6 0.588171
R2041 A2.n18 A2.n14 0.587949
R2042 A2.n3 A2.n0 0.567401
R2043 A2.n29 A2.n25 0.566642
R2044 A2.n24 A2.n20 0.566642
R2045 A2.n33 A2.n32 0.546848
R2046 A2.n34 A2.n3 0.423572
R2047 A2.n19 A2.n11 0.416362
R2048 A2.n31 A2.n30 0.416362
R2049 A2.n20 A2.n19 0.0273831
R2050 A2.n34 A2.n33 0.0273831
R2051 A2.n32 A2.n31 0.0250455
R2052 A2.n31 A2.n24 0.0149265
R2053 A2.n30 A2.n29 0.0149265
R2054 A2.n11 A2.n10 0.0118671
R2055 A2.n19 A2.n18 0.0118671
R2056 A2.n38 A2.n37 0.00291261
R2057 A2.n39 A2.n38 0.00259177
R2058 A2 A2.n34 0.00166883
C0 G_sink_up SD1_1 1.28f
C1 G_sink_dn G1_1 4.2e-19
C2 G1_1 G2_1 0.874f
C3 G_source_dn SD0_1 0.852f
C4 ITAIL_SRC ITAIL_SINK 0.00301f
C5 A1 A2 0.0522f
C6 G_sink_up G_sink_dn 2.32f
C7 ITAIL G2_1 5.61f
C8 G_sink_dn ITAIL_SINK 0.284f
C9 G_sink_up A2 0.18f
C10 G1_2 G1_1 4.36f
C11 SD0_1 SD1_1 0.0712f
C12 G2_1 SD2_1 0.473f
C13 G_sink_dn SD0_1 0.16f
C14 G_sink_up G1_2 0.585f
C15 ITAIL_SINK A2 0.945f
C16 G1_2 ITAIL 0.127f
C17 VDD G_source_dn 4.04f
C18 G1_2 SD2_1 0.118f
C19 VDD ITAIL_SRC 0.802f
C20 G_source_up A1 0.754f
C21 VDD SD1_1 0.848f
C22 SD0_1 G1_2 0.00621f
C23 VDD G_sink_dn 0.0064f
C24 G_source_dn ITAIL_SRC 0.406f
C25 G_source_up G_sink_up 0.0372f
C26 VDD G2_1 0.00603f
C27 G_source_dn SD1_1 0.0433f
C28 VDD A2 0.0289f
C29 A1 G_sink_up 0.00603f
C30 G_source_up ITAIL_SINK 5.02e-19
C31 G_source_dn G_sink_dn 0.32f
C32 G_sink_up G1_1 0.246f
C33 G1_1 ITAIL 0.618f
C34 VDD G1_2 13.9f
C35 G_source_dn A2 0.0015f
C36 G_source_up SD0_1 0.0116f
C37 A1 ITAIL_SINK 1.74e-19
C38 G_sink_dn SD1_1 0.0319f
C39 G1_1 SD2_1 2.49f
C40 G_sink_up ITAIL_SINK 0.182f
C41 ITAIL_SRC A2 4.12e-19
C42 G_source_dn G1_2 0.00217f
C43 SD0_1 G1_1 0.00104f
C44 ITAIL SD2_1 1.02f
C45 G_sink_up SD0_1 0.164f
C46 G_sink_dn A2 0.165f
C47 G1_2 SD1_1 0.376f
C48 VDD G_source_up 8.62f
C49 G_sink_dn G1_2 0.00586f
C50 G1_2 G2_1 0.00451f
C51 VDD A1 0.717f
C52 G_source_up G_source_dn 2.27f
C53 VDD G1_1 9.89f
C54 VDD G_sink_up 0.853f
C55 G_source_up ITAIL_SRC 0.231f
C56 G_source_dn A1 0.219f
C57 VDD ITAIL 0.207f
C58 G_source_up SD1_1 1.84e-20
C59 G_source_dn G1_1 6.12e-19
C60 VDD ITAIL_SINK 0.00102f
C61 G_source_dn G_sink_up 0.484f
C62 G_source_up G_sink_dn 0.00161f
C63 A1 ITAIL_SRC 0.901f
C64 VDD SD2_1 0.0868f
C65 G1_1 SD1_1 0.351f
C66 VDD SD0_1 0.0216f
C67 ITAIL_SRC G_sink_up 3.66e-19
C68 A1 G_sink_dn 0.00133f
C69 G_source_dn ITAIL_SINK 0.00133f
C70 G_source_up A2 0.0185f
.ends

