magic
tech gf180mcuC
magscale 1 10
timestamp 1714558667
<< nwell >>
rect 330 1402 1298 1521
rect 891 1333 1298 1402
rect 932 1313 1028 1333
rect 981 1300 1028 1313
rect 1095 1307 1118 1333
rect 475 998 476 1156
rect 560 953 564 955
rect 529 951 564 953
rect 664 951 686 959
rect 528 940 564 951
rect 529 928 564 940
rect 646 942 686 951
rect 721 942 768 955
rect 646 929 720 942
rect 530 898 564 928
rect 529 894 564 898
rect 530 891 564 894
rect 528 878 564 888
rect 621 882 720 929
rect 646 878 720 882
<< pwell >>
rect 599 785 621 786
rect 832 646 954 812
<< pdiff >>
rect 451 1011 475 1152
rect 451 1000 476 1011
rect 452 998 476 1000
<< psubdiff >>
rect 367 584 963 608
rect 367 534 391 584
rect 813 534 963 584
rect 367 528 963 534
rect 367 515 844 528
<< nsubdiff >>
rect 932 1463 1028 1495
rect 932 1417 955 1463
rect 1001 1417 1028 1463
rect 932 1313 1028 1417
rect 981 1300 1028 1313
rect 1074 1307 1118 1313
rect 1074 1286 1105 1307
<< psubdiffcont >>
rect 391 534 813 584
<< nsubdiffcont >>
rect 955 1417 1001 1463
<< polysilicon >>
rect 504 878 560 954
rect 664 951 720 959
rect 646 938 720 951
rect 646 891 659 938
rect 707 891 720 938
rect 646 878 720 891
rect 488 876 560 878
rect 470 865 560 876
rect 470 818 495 865
rect 543 818 560 865
rect 470 807 560 818
rect 488 805 560 807
rect 504 781 560 805
rect 672 781 720 878
<< polycontact >>
rect 659 891 707 938
rect 495 818 543 865
<< metal1 >>
rect 330 1495 976 1521
rect 330 1463 1028 1495
rect 330 1417 955 1463
rect 1001 1417 1028 1463
rect 330 1402 1028 1417
rect 422 998 479 1402
rect 894 1318 1028 1402
rect 749 1011 897 1058
rect 646 938 720 942
rect 646 929 659 938
rect 621 891 659 929
rect 707 891 720 938
rect 621 882 720 891
rect 646 878 720 882
rect 460 865 544 876
rect 460 818 495 865
rect 543 818 544 865
rect 850 832 897 1011
rect 1214 837 1298 895
rect 460 807 544 818
rect 592 785 897 832
rect 422 629 471 738
rect 592 691 641 785
rect 758 629 807 739
rect 330 608 894 629
rect 330 584 950 608
rect 330 534 391 584
rect 813 544 950 584
rect 813 534 894 544
rect 330 510 894 534
use GF_INV_MAG  GF_INV_MAG_1
timestamp 1714558667
transform 1 0 1012 0 1 706
box -118 -175 286 666
use nmos_3p3_DDNVWA  nmos_3p3_DDNVWA_0
timestamp 1714126980
transform 1 0 700 0 1 715
box -144 -97 144 97
use nmos_3p3_DDNVWA  nmos_3p3_DDNVWA_1
timestamp 1714126980
transform 1 0 532 0 1 715
box -144 -97 144 97
use pmos_3p3_M4YALR  pmos_3p3_M4YALR_0
timestamp 1714126980
transform 1 0 692 0 1 1158
box -202 -290 202 290
use pmos_3p3_M8QNDR  pmos_3p3_M8QNDR_0
timestamp 1714126980
transform 1 0 532 0 1 1158
box -202 -290 202 290
<< labels >>
flabel psubdiffcont 598 561 598 561 0 FreeSans 320 0 0 0 VSS
port 0 nsew
flabel metal1 464 836 464 836 0 FreeSans 320 0 0 0 IN2
port 2 nsew
flabel metal1 634 907 634 907 0 FreeSans 320 0 0 0 IN1
port 3 nsew
flabel metal1 1262 858 1262 858 0 FreeSans 320 0 0 0 OUT
port 4 nsew
<< end >>
