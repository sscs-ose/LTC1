* NGSPICE file created from cap80p_mag_flat.ext - technology: gf180mcuC

.subckt pex_cap80p_mag N P
X0 P.t0 N.t63 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X1 P.t1 N.t62 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X2 P.t2 N.t61 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X3 P.t3 N.t60 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X4 P.t4 N.t59 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X5 P.t5 N.t58 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X6 P.t6 N.t57 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X7 P.t7 N.t56 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X8 P.t8 N.t55 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X9 P.t9 N.t54 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X10 P.t10 N.t53 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X11 P.t11 N.t52 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X12 P.t12 N.t51 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X13 P.t13 N.t50 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X14 P.t14 N.t49 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X15 P.t15 N.t48 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X16 P.t16 N.t47 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X17 P.t17 N.t46 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X18 P.t18 N.t45 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X19 P.t19 N.t44 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X20 P.t20 N.t43 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X21 P.t21 N.t42 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X22 P.t22 N.t41 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X23 P.t23 N.t40 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X24 P.t24 N.t39 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X25 P.t25 N.t38 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X26 P.t26 N.t37 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X27 P.t27 N.t36 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X28 P.t28 N.t35 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X29 P.t29 N.t34 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X30 P.t30 N.t33 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X31 P.t31 N.t32 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X32 P.t32 N.t31 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X33 P.t33 N.t30 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X34 P.t34 N.t29 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X35 P.t35 N.t28 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X36 P.t36 N.t27 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X37 P.t37 N.t26 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X38 P.t38 N.t25 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X39 P.t39 N.t24 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X40 P.t40 N.t23 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X41 P.t41 N.t22 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X42 P.t42 N.t21 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X43 P.t43 N.t20 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X44 P.t44 N.t19 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X45 P.t45 N.t18 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X46 P.t46 N.t17 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X47 P.t47 N.t16 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X48 P.t48 N.t15 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X49 P.t49 N.t14 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X50 P.t50 N.t13 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X51 P.t51 N.t12 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X52 P.t52 N.t11 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X53 P.t53 N.t10 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X54 P.t54 N.t9 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X55 P.t55 N.t8 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X56 P.t56 N.t7 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X57 P.t57 N.t6 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X58 P.t58 N.t5 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X59 P.t59 N.t4 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X60 P.t60 N.t3 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X61 P.t61 N.t2 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X62 P.t62 N.t1 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X63 P.t63 N.t0 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
R0 P P.n76 4.52515
R1 P.n2 P.t4 2.38861
R2 P.n54 P.t22 2.38861
R3 P.n47 P.t3 2.38861
R4 P.n40 P.t57 2.38861
R5 P.n9 P.t16 2.38861
R6 P.n16 P.t5 2.38861
R7 P.n23 P.t29 2.38861
R8 P.n30 P.t46 2.38861
R9 P.n2 P.t62 2.2505
R10 P.n3 P.t42 2.2505
R11 P.n4 P.t36 2.2505
R12 P.n5 P.t10 2.2505
R13 P.n6 P.t24 2.2505
R14 P.n7 P.t27 2.2505
R15 P.n8 P.t6 2.2505
R16 P.n54 P.t18 2.2505
R17 P.n55 P.t56 2.2505
R18 P.n56 P.t52 2.2505
R19 P.n57 P.t30 2.2505
R20 P.n58 P.t40 2.2505
R21 P.n59 P.t0 2.2505
R22 P.n60 P.t19 2.2505
R23 P.n47 P.t1 2.2505
R24 P.n48 P.t41 2.2505
R25 P.n49 P.t35 2.2505
R26 P.n50 P.t9 2.2505
R27 P.n51 P.t23 2.2505
R28 P.n52 P.t17 2.2505
R29 P.n53 P.t2 2.2505
R30 P.n40 P.t53 2.2505
R31 P.n41 P.t31 2.2505
R32 P.n42 P.t28 2.2505
R33 P.n43 P.t61 2.2505
R34 P.n44 P.t8 2.2505
R35 P.n45 P.t20 2.2505
R36 P.n46 P.t38 2.2505
R37 P.n9 P.t14 2.2505
R38 P.n10 P.t50 2.2505
R39 P.n11 P.t48 2.2505
R40 P.n12 P.t21 2.2505
R41 P.n13 P.t34 2.2505
R42 P.n14 P.t7 2.2505
R43 P.n15 P.t39 2.2505
R44 P.n16 P.t63 2.2505
R45 P.n17 P.t43 2.2505
R46 P.n18 P.t37 2.2505
R47 P.n19 P.t11 2.2505
R48 P.n20 P.t25 2.2505
R49 P.n21 P.t33 2.2505
R50 P.n22 P.t13 2.2505
R51 P.n23 P.t26 2.2505
R52 P.n24 P.t59 2.2505
R53 P.n25 P.t55 2.2505
R54 P.n26 P.t32 2.2505
R55 P.n27 P.t45 2.2505
R56 P.n28 P.t60 2.2505
R57 P.n29 P.t47 2.2505
R58 P.n30 P.t44 2.2505
R59 P.n31 P.t15 2.2505
R60 P.n32 P.t12 2.2505
R61 P.n33 P.t49 2.2505
R62 P.n34 P.t58 2.2505
R63 P.n35 P.t54 2.2505
R64 P.n36 P.t51 2.2505
R65 P.n73 P.n72 1.5005
R66 P.n66 P.n65 1.5005
R67 P.n61 P.n60 1.14654
R68 P.n37 P.n36 1.14654
R69 P.n69 P.n68 1.1247
R70 P.n38 P.n37 1.05975
R71 P.n39 P.n38 1.05975
R72 P.n63 P.n39 1.05975
R73 P.n63 P.n62 1.05975
R74 P.n62 P.n61 1.05975
R75 P.n64 P.n63 0.169179
R76 P.n3 P.n2 0.138613
R77 P.n4 P.n3 0.138613
R78 P.n5 P.n4 0.138613
R79 P.n6 P.n5 0.138613
R80 P.n7 P.n6 0.138613
R81 P.n8 P.n7 0.138613
R82 P.n55 P.n54 0.138613
R83 P.n56 P.n55 0.138613
R84 P.n57 P.n56 0.138613
R85 P.n58 P.n57 0.138613
R86 P.n59 P.n58 0.138613
R87 P.n60 P.n59 0.138613
R88 P.n48 P.n47 0.138613
R89 P.n49 P.n48 0.138613
R90 P.n50 P.n49 0.138613
R91 P.n51 P.n50 0.138613
R92 P.n52 P.n51 0.138613
R93 P.n53 P.n52 0.138613
R94 P.n41 P.n40 0.138613
R95 P.n42 P.n41 0.138613
R96 P.n43 P.n42 0.138613
R97 P.n44 P.n43 0.138613
R98 P.n45 P.n44 0.138613
R99 P.n46 P.n45 0.138613
R100 P.n10 P.n9 0.138613
R101 P.n11 P.n10 0.138613
R102 P.n12 P.n11 0.138613
R103 P.n13 P.n12 0.138613
R104 P.n14 P.n13 0.138613
R105 P.n15 P.n14 0.138613
R106 P.n17 P.n16 0.138613
R107 P.n18 P.n17 0.138613
R108 P.n19 P.n18 0.138613
R109 P.n20 P.n19 0.138613
R110 P.n21 P.n20 0.138613
R111 P.n22 P.n21 0.138613
R112 P.n24 P.n23 0.138613
R113 P.n25 P.n24 0.138613
R114 P.n26 P.n25 0.138613
R115 P.n27 P.n26 0.138613
R116 P.n28 P.n27 0.138613
R117 P.n29 P.n28 0.138613
R118 P.n31 P.n30 0.138613
R119 P.n32 P.n31 0.138613
R120 P.n33 P.n32 0.138613
R121 P.n34 P.n33 0.138613
R122 P.n35 P.n34 0.138613
R123 P.n36 P.n35 0.138613
R124 P.n63 P.n8 0.0872924
R125 P.n61 P.n53 0.0872924
R126 P.n62 P.n46 0.0872924
R127 P.n39 P.n15 0.0872924
R128 P.n38 P.n22 0.0872924
R129 P.n37 P.n29 0.0872924
R130 P.n76 P.n75 0.0357703
R131 P.n66 P.n1 0.0350405
R132 P.n72 P.n67 0.0267703
R133 P.n70 P.n69 0.00798833
R134 P.n74 P.n73 0.00341892
R135 P.n71 P.n70 0.00268919
R136 P.n72 P.n71 0.00244595
R137 P P.n0 0.0017973
R138 P.n75 P.n74 0.00171622
R139 P.n73 P.n66 0.00122973
R140 P.n65 P.n64 0.000932432
R141 P.n65 P.n0 0.000824324
R142 N N.n74 4.52418
R143 N.n52 N.t44 3.26618
R144 N.n21 N.t12 3.26618
R145 N.n14 N.t16 3.26618
R146 N.n7 N.t50 3.26618
R147 N.n0 N.t24 3.26618
R148 N.n31 N.t57 3.26618
R149 N.n38 N.t25 3.26618
R150 N.n45 N.t61 3.26618
R151 N.n52 N.t63 2.25486
R152 N.n53 N.t23 2.25486
R153 N.n54 N.t33 2.25486
R154 N.n55 N.t11 2.25486
R155 N.n56 N.t7 2.25486
R156 N.n57 N.t45 2.25486
R157 N.n58 N.t41 2.25486
R158 N.n21 N.t9 2.25486
R159 N.n22 N.t5 2.25486
R160 N.n23 N.t14 2.25486
R161 N.n24 N.t51 2.25486
R162 N.n25 N.t48 2.25486
R163 N.n26 N.t19 2.25486
R164 N.n27 N.t17 2.25486
R165 N.n14 N.t3 2.25486
R166 N.n15 N.t18 2.25486
R167 N.n16 N.t31 2.25486
R168 N.n17 N.t8 2.25486
R169 N.n18 N.t4 2.25486
R170 N.n19 N.t37 2.25486
R171 N.n20 N.t34 2.25486
R172 N.n7 N.t30 2.25486
R173 N.n8 N.t38 2.25486
R174 N.n9 N.t52 2.25486
R175 N.n10 N.t26 2.25486
R176 N.n11 N.t20 2.25486
R177 N.n12 N.t0 2.25486
R178 N.n13 N.t58 2.25486
R179 N.n0 N.t56 2.25486
R180 N.n1 N.t29 2.25486
R181 N.n2 N.t42 2.25486
R182 N.n3 N.t15 2.25486
R183 N.n4 N.t13 2.25486
R184 N.n5 N.t49 2.25486
R185 N.n6 N.t47 2.25486
R186 N.n31 N.t36 2.25486
R187 N.n32 N.t39 2.25486
R188 N.n33 N.t53 2.25486
R189 N.n34 N.t27 2.25486
R190 N.n35 N.t21 2.25486
R191 N.n36 N.t1 2.25486
R192 N.n37 N.t59 2.25486
R193 N.n38 N.t43 2.25486
R194 N.n39 N.t55 2.25486
R195 N.n40 N.t2 2.25486
R196 N.n41 N.t35 2.25486
R197 N.n42 N.t32 2.25486
R198 N.n43 N.t10 2.25486
R199 N.n44 N.t6 2.25486
R200 N.n45 N.t46 2.25486
R201 N.n46 N.t40 2.25486
R202 N.n47 N.t54 2.25486
R203 N.n48 N.t28 2.25486
R204 N.n49 N.t22 2.25486
R205 N.n50 N.t62 2.25486
R206 N.n51 N.t60 2.25486
R207 N.n28 N.n27 1.63171
R208 N.n59 N.n58 1.63033
R209 N.n71 N.n70 1.5005
R210 N.n67 N.n66 1.1247
R211 N.n30 N.n29 1.07514
R212 N.n61 N.n60 1.07514
R213 N.n29 N.n28 1.07476
R214 N.n60 N.n59 1.07438
R215 N.n53 N.n52 1.01182
R216 N.n54 N.n53 1.01182
R217 N.n55 N.n54 1.01182
R218 N.n56 N.n55 1.01182
R219 N.n57 N.n56 1.01182
R220 N.n58 N.n57 1.01182
R221 N.n22 N.n21 1.01182
R222 N.n23 N.n22 1.01182
R223 N.n24 N.n23 1.01182
R224 N.n25 N.n24 1.01182
R225 N.n26 N.n25 1.01182
R226 N.n27 N.n26 1.01182
R227 N.n15 N.n14 1.01182
R228 N.n16 N.n15 1.01182
R229 N.n17 N.n16 1.01182
R230 N.n18 N.n17 1.01182
R231 N.n19 N.n18 1.01182
R232 N.n20 N.n19 1.01182
R233 N.n8 N.n7 1.01182
R234 N.n9 N.n8 1.01182
R235 N.n10 N.n9 1.01182
R236 N.n11 N.n10 1.01182
R237 N.n12 N.n11 1.01182
R238 N.n13 N.n12 1.01182
R239 N.n1 N.n0 1.01182
R240 N.n2 N.n1 1.01182
R241 N.n3 N.n2 1.01182
R242 N.n4 N.n3 1.01182
R243 N.n5 N.n4 1.01182
R244 N.n6 N.n5 1.01182
R245 N.n32 N.n31 1.01182
R246 N.n33 N.n32 1.01182
R247 N.n34 N.n33 1.01182
R248 N.n35 N.n34 1.01182
R249 N.n36 N.n35 1.01182
R250 N.n37 N.n36 1.01182
R251 N.n39 N.n38 1.01182
R252 N.n40 N.n39 1.01182
R253 N.n41 N.n40 1.01182
R254 N.n42 N.n41 1.01182
R255 N.n43 N.n42 1.01182
R256 N.n44 N.n43 1.01182
R257 N.n46 N.n45 1.01182
R258 N.n47 N.n46 1.01182
R259 N.n48 N.n47 1.01182
R260 N.n49 N.n48 1.01182
R261 N.n50 N.n49 1.01182
R262 N.n51 N.n50 1.01182
R263 N.n64 N.n63 0.898925
R264 N.n62 N.n61 0.896194
R265 N.n28 N.n20 0.556878
R266 N.n29 N.n13 0.556878
R267 N.n30 N.n6 0.556878
R268 N.n61 N.n37 0.556878
R269 N.n60 N.n44 0.556878
R270 N.n59 N.n51 0.556878
R271 N.n62 N.n30 0.179065
R272 N.n63 N.n62 0.122988
R273 N.n74 N.n73 0.0347973
R274 N.n70 N.n65 0.0267703
R275 N.n71 N.n64 0.008809
R276 N.n68 N.n67 0.00798833
R277 N.n72 N.n71 0.00463514
R278 N.n69 N.n68 0.00268919
R279 N.n70 N.n69 0.00244595
R280 N.n73 N.n72 0.00147297
R281 N N.n63 0.000932432
C0 N P 0.294p
C1 N VSUBS 0.105p
C2 P VSUBS 0.353p
C3 N.t24 VSUBS 3.73f
C4 N.t56 VSUBS 3.41f
C5 N.n0 VSUBS 1.77f
C6 N.t29 VSUBS 3.41f
C7 N.n1 VSUBS 1.05f
C8 N.t42 VSUBS 3.41f
C9 N.n2 VSUBS 1.05f
C10 N.t15 VSUBS 3.41f
C11 N.n3 VSUBS 1.05f
C12 N.t13 VSUBS 3.41f
C13 N.n4 VSUBS 1.05f
C14 N.t49 VSUBS 3.41f
C15 N.n5 VSUBS 1.05f
C16 N.t47 VSUBS 3.41f
C17 N.n6 VSUBS 0.81f
C18 N.t50 VSUBS 3.73f
C19 N.t30 VSUBS 3.41f
C20 N.n7 VSUBS 1.77f
C21 N.t38 VSUBS 3.41f
C22 N.n8 VSUBS 1.05f
C23 N.t52 VSUBS 3.41f
C24 N.n9 VSUBS 1.05f
C25 N.t26 VSUBS 3.41f
C26 N.n10 VSUBS 1.05f
C27 N.t20 VSUBS 3.41f
C28 N.n11 VSUBS 1.05f
C29 N.t0 VSUBS 3.41f
C30 N.n12 VSUBS 1.05f
C31 N.t58 VSUBS 3.41f
C32 N.n13 VSUBS 0.81f
C33 N.t16 VSUBS 3.73f
C34 N.t3 VSUBS 3.41f
C35 N.n14 VSUBS 1.77f
C36 N.t18 VSUBS 3.41f
C37 N.n15 VSUBS 1.05f
C38 N.t31 VSUBS 3.41f
C39 N.n16 VSUBS 1.05f
C40 N.t8 VSUBS 3.41f
C41 N.n17 VSUBS 1.05f
C42 N.t4 VSUBS 3.41f
C43 N.n18 VSUBS 1.05f
C44 N.t37 VSUBS 3.41f
C45 N.n19 VSUBS 1.05f
C46 N.t34 VSUBS 3.41f
C47 N.n20 VSUBS 0.81f
C48 N.t12 VSUBS 3.73f
C49 N.t9 VSUBS 3.41f
C50 N.n21 VSUBS 1.77f
C51 N.t5 VSUBS 3.41f
C52 N.n22 VSUBS 1.05f
C53 N.t14 VSUBS 3.41f
C54 N.n23 VSUBS 1.05f
C55 N.t51 VSUBS 3.41f
C56 N.n24 VSUBS 1.05f
C57 N.t48 VSUBS 3.41f
C58 N.n25 VSUBS 1.05f
C59 N.t19 VSUBS 3.41f
C60 N.n26 VSUBS 1.05f
C61 N.t17 VSUBS 3.41f
C62 N.n27 VSUBS 1.37f
C63 N.n28 VSUBS 1.65f
C64 N.n29 VSUBS 1.36f
C65 N.n30 VSUBS 0.914f
C66 N.t57 VSUBS 3.73f
C67 N.t36 VSUBS 3.41f
C68 N.n31 VSUBS 1.77f
C69 N.t39 VSUBS 3.41f
C70 N.n32 VSUBS 1.05f
C71 N.t53 VSUBS 3.41f
C72 N.n33 VSUBS 1.05f
C73 N.t27 VSUBS 3.41f
C74 N.n34 VSUBS 1.05f
C75 N.t21 VSUBS 3.41f
C76 N.n35 VSUBS 1.05f
C77 N.t1 VSUBS 3.41f
C78 N.n36 VSUBS 1.05f
C79 N.t59 VSUBS 3.41f
C80 N.n37 VSUBS 0.81f
C81 N.t25 VSUBS 3.73f
C82 N.t43 VSUBS 3.41f
C83 N.n38 VSUBS 1.77f
C84 N.t55 VSUBS 3.41f
C85 N.n39 VSUBS 1.05f
C86 N.t2 VSUBS 3.41f
C87 N.n40 VSUBS 1.05f
C88 N.t35 VSUBS 3.41f
C89 N.n41 VSUBS 1.05f
C90 N.t32 VSUBS 3.41f
C91 N.n42 VSUBS 1.05f
C92 N.t10 VSUBS 3.41f
C93 N.n43 VSUBS 1.05f
C94 N.t6 VSUBS 3.41f
C95 N.n44 VSUBS 0.81f
C96 N.t61 VSUBS 3.73f
C97 N.t46 VSUBS 3.41f
C98 N.n45 VSUBS 1.77f
C99 N.t40 VSUBS 3.41f
C100 N.n46 VSUBS 1.05f
C101 N.t54 VSUBS 3.41f
C102 N.n47 VSUBS 1.05f
C103 N.t28 VSUBS 3.41f
C104 N.n48 VSUBS 1.05f
C105 N.t22 VSUBS 3.41f
C106 N.n49 VSUBS 1.05f
C107 N.t62 VSUBS 3.41f
C108 N.n50 VSUBS 1.05f
C109 N.t60 VSUBS 3.41f
C110 N.n51 VSUBS 0.81f
C111 N.t44 VSUBS 3.73f
C112 N.t63 VSUBS 3.41f
C113 N.n52 VSUBS 1.77f
C114 N.t23 VSUBS 3.41f
C115 N.n53 VSUBS 1.05f
C116 N.t33 VSUBS 3.41f
C117 N.n54 VSUBS 1.05f
C118 N.t11 VSUBS 3.41f
C119 N.n55 VSUBS 1.05f
C120 N.t7 VSUBS 3.41f
C121 N.n56 VSUBS 1.05f
C122 N.t45 VSUBS 3.41f
C123 N.n57 VSUBS 1.05f
C124 N.t41 VSUBS 3.41f
C125 N.n58 VSUBS 1.37f
C126 N.n59 VSUBS 1.65f
C127 N.n60 VSUBS 1.36f
C128 N.n61 VSUBS 1.27f
C129 N.n62 VSUBS 0.6f
C130 N.n63 VSUBS 0.151f
C131 N.n64 VSUBS 0.0603f
C132 N.n65 VSUBS 0.0659f
C133 N.n66 VSUBS 0.325f
C134 N.n67 VSUBS 0.0542f
C135 N.n68 VSUBS 0.0212f
C136 N.n69 VSUBS 0.00289f
C137 N.n70 VSUBS 0.0197f
C138 N.n71 VSUBS 0.0262f
C139 N.n72 VSUBS 0.00357f
C140 N.n73 VSUBS 0.0246f
C141 N.n74 VSUBS 0.0488f
C142 P.n0 VSUBS 2.62e-19
C143 P.n1 VSUBS 0.00603f
C144 P.t6 VSUBS 2.36f
C145 P.t27 VSUBS 2.36f
C146 P.t24 VSUBS 2.36f
C147 P.t10 VSUBS 2.36f
C148 P.t36 VSUBS 2.36f
C149 P.t42 VSUBS 2.36f
C150 P.t62 VSUBS 2.36f
C151 P.t4 VSUBS 2.49f
C152 P.n2 VSUBS 4.3f
C153 P.n3 VSUBS 2.22f
C154 P.n4 VSUBS 2.22f
C155 P.n5 VSUBS 2.22f
C156 P.n6 VSUBS 2.22f
C157 P.n7 VSUBS 2.22f
C158 P.n8 VSUBS 2.09f
C159 P.t39 VSUBS 2.36f
C160 P.t7 VSUBS 2.36f
C161 P.t34 VSUBS 2.36f
C162 P.t21 VSUBS 2.36f
C163 P.t48 VSUBS 2.36f
C164 P.t50 VSUBS 2.36f
C165 P.t14 VSUBS 2.36f
C166 P.t16 VSUBS 2.49f
C167 P.n9 VSUBS 4.3f
C168 P.n10 VSUBS 2.22f
C169 P.n11 VSUBS 2.22f
C170 P.n12 VSUBS 2.22f
C171 P.n13 VSUBS 2.22f
C172 P.n14 VSUBS 2.22f
C173 P.n15 VSUBS 2.09f
C174 P.t13 VSUBS 2.36f
C175 P.t33 VSUBS 2.36f
C176 P.t25 VSUBS 2.36f
C177 P.t11 VSUBS 2.36f
C178 P.t37 VSUBS 2.36f
C179 P.t43 VSUBS 2.36f
C180 P.t63 VSUBS 2.36f
C181 P.t5 VSUBS 2.49f
C182 P.n16 VSUBS 4.3f
C183 P.n17 VSUBS 2.22f
C184 P.n18 VSUBS 2.22f
C185 P.n19 VSUBS 2.22f
C186 P.n20 VSUBS 2.22f
C187 P.n21 VSUBS 2.22f
C188 P.n22 VSUBS 2.09f
C189 P.t47 VSUBS 2.36f
C190 P.t60 VSUBS 2.36f
C191 P.t45 VSUBS 2.36f
C192 P.t32 VSUBS 2.36f
C193 P.t55 VSUBS 2.36f
C194 P.t59 VSUBS 2.36f
C195 P.t26 VSUBS 2.36f
C196 P.t29 VSUBS 2.49f
C197 P.n23 VSUBS 4.3f
C198 P.n24 VSUBS 2.22f
C199 P.n25 VSUBS 2.22f
C200 P.n26 VSUBS 2.22f
C201 P.n27 VSUBS 2.22f
C202 P.n28 VSUBS 2.22f
C203 P.n29 VSUBS 2.09f
C204 P.t51 VSUBS 2.36f
C205 P.t54 VSUBS 2.36f
C206 P.t58 VSUBS 2.36f
C207 P.t49 VSUBS 2.36f
C208 P.t12 VSUBS 2.36f
C209 P.t15 VSUBS 2.36f
C210 P.t44 VSUBS 2.36f
C211 P.t46 VSUBS 2.49f
C212 P.n30 VSUBS 4.3f
C213 P.n31 VSUBS 2.22f
C214 P.n32 VSUBS 2.22f
C215 P.n33 VSUBS 2.22f
C216 P.n34 VSUBS 2.22f
C217 P.n35 VSUBS 2.22f
C218 P.n36 VSUBS 2.27f
C219 P.n37 VSUBS 0.258f
C220 P.n38 VSUBS 0.244f
C221 P.n39 VSUBS 0.244f
C222 P.t38 VSUBS 2.36f
C223 P.t20 VSUBS 2.36f
C224 P.t8 VSUBS 2.36f
C225 P.t61 VSUBS 2.36f
C226 P.t28 VSUBS 2.36f
C227 P.t31 VSUBS 2.36f
C228 P.t53 VSUBS 2.36f
C229 P.t57 VSUBS 2.49f
C230 P.n40 VSUBS 4.3f
C231 P.n41 VSUBS 2.22f
C232 P.n42 VSUBS 2.22f
C233 P.n43 VSUBS 2.22f
C234 P.n44 VSUBS 2.22f
C235 P.n45 VSUBS 2.22f
C236 P.n46 VSUBS 2.09f
C237 P.t2 VSUBS 2.36f
C238 P.t17 VSUBS 2.36f
C239 P.t23 VSUBS 2.36f
C240 P.t9 VSUBS 2.36f
C241 P.t35 VSUBS 2.36f
C242 P.t41 VSUBS 2.36f
C243 P.t1 VSUBS 2.36f
C244 P.t3 VSUBS 2.49f
C245 P.n47 VSUBS 4.3f
C246 P.n48 VSUBS 2.22f
C247 P.n49 VSUBS 2.22f
C248 P.n50 VSUBS 2.22f
C249 P.n51 VSUBS 2.22f
C250 P.n52 VSUBS 2.22f
C251 P.n53 VSUBS 2.09f
C252 P.t19 VSUBS 2.36f
C253 P.t0 VSUBS 2.36f
C254 P.t40 VSUBS 2.36f
C255 P.t30 VSUBS 2.36f
C256 P.t52 VSUBS 2.36f
C257 P.t56 VSUBS 2.36f
C258 P.t18 VSUBS 2.36f
C259 P.t22 VSUBS 2.49f
C260 P.n54 VSUBS 4.3f
C261 P.n55 VSUBS 2.22f
C262 P.n56 VSUBS 2.22f
C263 P.n57 VSUBS 2.22f
C264 P.n58 VSUBS 2.22f
C265 P.n59 VSUBS 2.22f
C266 P.n60 VSUBS 2.27f
C267 P.n61 VSUBS 0.258f
C268 P.n62 VSUBS 0.244f
C269 P.n63 VSUBS 0.253f
C270 P.n64 VSUBS 0.0173f
C271 P.n65 VSUBS 1.22e-19
C272 P.n66 VSUBS 0.00253f
C273 P.n67 VSUBS 0.00674f
C274 P.n68 VSUBS 0.0334f
C275 P.n69 VSUBS 0.00557f
C276 P.n70 VSUBS 0.00218f
C277 P.n71 VSUBS 2.97e-19
C278 P.n72 VSUBS 0.00202f
C279 P.n73 VSUBS 2.62e-19
C280 P.n74 VSUBS 2.97e-19
C281 P.n75 VSUBS 0.00262f
C282 P.n76 VSUBS 0.00509f
.ends

