* NGSPICE file created from MUX_1x8_flat.ext - technology: gf180mcuC

.subckt pex_MUX_1x8 VDD Vout VSS A0 A1 A2 A3 A4 A5 A6 A7 S0 S1 S2 ENA
X0 TG_magic_5.A a_3874_308.t6 TG_GATE_SWITCH_magic_7.B.t61 VDD.t297 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 TG_GATE_SWITCH_magic_1.B a_n4297_n4860.t6 A3.t23 VDD.t2 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 TG_magic_0.A TG_magic_1.CLK TG_GATE_SWITCH_magic_0.B.t34 VSS.t94 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 Vout INVERTER_MUX_1.OUT.t16 TG_magic_0.B.t36 VSS.t138 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X4 INVERTER_MUX_1.OUT S2.t0 VSS.t185 VSS.t35 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X5 A5 a_n4297_n7438.t6 TG_GATE_SWITCH_magic_2.B.t23 VDD.t186 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X6 VSS S1.t0 TG_magic_7.CLK VSS.t16 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X7 TG_GATE_SWITCH_magic_2.B a_n4701_n7438# A5.t35 VSS.t209 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X8 TG_GATE_SWITCH_magic_2.B a_n4297_n7438.t7 A5.t22 VDD.t176 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X9 VSS S2.t1 INVERTER_MUX_1.OUT.t12 VSS.t186 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X10 TG_GATE_SWITCH_magic_6.B a_n2298_n2271# A4.t20 VSS.t41 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X11 TG_magic_0.B a_2061_n2270.t6 TG_magic_0.A.t77 VDD.t13 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X12 TG_GATE_SWITCH_magic_3.B a_5684_1104.t6 TG_magic_5.A.t53 VDD.t238 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X13 TG_magic_0.B a_3817_n991.t6 TG_magic_5.A.t70 VDD.t63 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X14 TG_magic_7.B S1.t1 TG_magic_4.B.t100 VSS.t159 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X15 VDD S0.t0 a_5684_n6152.t3 VDD.t20 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X16 TG_GATE_SWITCH_magic_2.B a_n4297_n7438.t8 A5.t21 VDD.t245 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X17 TG_magic_0.A a_301_308.t6 TG_GATE_SWITCH_magic_6.B.t30 VDD.t83 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X18 A6 a_n4297_300.t6 TG_GATE_SWITCH_magic_3.B.t8 VDD.t77 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X19 TG_GATE_SWITCH_magic_0.B TG_magic_1.CLK TG_magic_0.A.t56 VSS.t93 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X20 TG_GATE_SWITCH_magic_1.B TG_magic_1.CLK TG_magic_4.B.t62 VSS.t74 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X21 a_n2298_307# ENA.t0 VDD.t89 VDD.t88 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X22 TG_magic_4.B a_2061_n4852.t6 TG_magic_7.B.t103 VDD.t15 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X23 Vout S2.t2 TG_magic_7.B.t78 VSS.t23 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X24 TG_magic_5.A a_3874_308.t7 TG_GATE_SWITCH_magic_7.B.t60 VDD.t297 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X25 TG_GATE_SWITCH_magic_1.B a_n4297_n4860.t7 A3.t22 VDD.t2 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X26 TG_GATE_SWITCH_magic_1.B a_n4297_n4860.t8 A3.t21 VDD.t3 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X27 TG_magic_7.B TG_magic_7.CLK TG_magic_2.B.t107 VSS.t225 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X28 TG_GATE_SWITCH_magic_6.B a_n1894_n2271.t6 A4.t27 VDD.t10 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X29 TG_GATE_SWITCH_magic_1.B a_2004_n6151.t6 TG_magic_4.B.t13 VDD.t46 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X30 A5 a_n4701_n7438# TG_GATE_SWITCH_magic_2.B.t59 VSS.t208 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X31 TG_magic_0.B TG_magic_7.CLK TG_magic_0.A.t107 VSS.t226 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X32 TG_magic_5.A a_3874_308.t8 TG_GATE_SWITCH_magic_7.B.t59 VDD.t294 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X33 TG_magic_7.B a_5741_n4853.t6 Vout.t51 VDD.t58 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X34 TG_magic_4.B S0.t1 TG_GATE_SWITCH_magic_5.B.t16 VSS.t128 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X35 TG_magic_0.A S0.t2 TG_GATE_SWITCH_magic_6.B.t27 VSS.t5 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X36 A0 a_n4297_n2278.t6 TG_GATE_SWITCH_magic_0.B.t50 VDD.t18 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X37 VSS TG_magic_1.CLK a_2004_n6151.t5 VSS.t101 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X38 VDD S1.t3 a_3817_n991.t3 VDD.t177 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X39 TG_GATE_SWITCH_magic_2.B a_5684_n6152.t6 TG_magic_2.B.t58 VDD.t287 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X40 A7 a_n2298_n4853# TG_GATE_SWITCH_magic_5.B.t45 VSS.t146 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X41 TG_magic_0.A a_301_308.t7 TG_GATE_SWITCH_magic_6.B.t23 VDD.t83 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X42 VDD S2.t3 INVERTER_MUX_1.OUT.t13 VDD.t203 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X43 A0 a_n4297_n2278.t7 TG_GATE_SWITCH_magic_0.B.t49 VDD.t19 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X44 TG_magic_4.B a_301_n7430.t6 TG_GATE_SWITCH_magic_5.B.t71 VDD.t44 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X45 VDD TG_magic_1.CLK a_2004_n6151.t3 VDD.t125 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X46 A2 a_n1894_307.t6 TG_GATE_SWITCH_magic_7.B.t40 VDD.t106 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X47 TG_GATE_SWITCH_magic_0.B a_2004_1105.t6 TG_magic_0.A.t14 VDD.t69 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X48 TG_GATE_SWITCH_magic_6.B a_n1894_n2271.t7 A4.t28 VDD.t10 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X49 Vout a_5741_n4853.t7 TG_magic_7.B.t107 VDD.t56 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X50 TG_GATE_SWITCH_magic_3.B a_n4297_300.t7 A6.t34 VDD.t174 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X51 TG_magic_0.A a_2061_n2270.t7 TG_magic_0.B.t55 VDD.t14 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X52 TG_GATE_SWITCH_magic_3.B a_n4297_300.t8 A6.t33 VDD.t174 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X53 TG_magic_5.A a_5684_1104.t7 TG_GATE_SWITCH_magic_3.B.t52 VDD.t234 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X54 TG_magic_2.B TG_magic_1.CLK TG_GATE_SWITCH_magic_4.B.t20 VSS.t72 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X55 TG_GATE_SWITCH_magic_6.B a_301_308.t8 TG_magic_0.A.t65 VDD.t79 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X56 a_n4701_n4860# ENA.t1 VDD.t91 VDD.t90 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X57 TG_GATE_SWITCH_magic_2.B a_n4701_n7438# A5.t33 VSS.t207 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X58 TG_magic_2.B a_3874_n7430.t6 TG_GATE_SWITCH_magic_4.B.t0 VDD.t52 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X59 TG_magic_7.B a_2061_n4852.t7 TG_magic_4.B.t72 VDD.t16 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X60 TG_magic_5.A S1.t4 TG_magic_0.B.t37 VSS.t149 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X61 Vout a_5741_n4853.t8 TG_magic_7.B.t104 VDD.t54 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X62 TG_GATE_SWITCH_magic_2.B a_5684_n6152.t7 TG_magic_2.B.t57 VDD.t288 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X63 TG_GATE_SWITCH_magic_0.B TG_magic_1.CLK TG_magic_0.A.t55 VSS.t89 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X64 TG_magic_4.B a_2004_n6151.t7 TG_GATE_SWITCH_magic_1.B.t1 VDD.t47 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X65 TG_magic_7.B a_3817_n4055.t6 TG_magic_2.B.t59 VDD.t65 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X66 Vout a_5741_n4853.t9 TG_magic_7.B.t48 VDD.t57 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X67 TG_magic_0.A a_301_308.t9 TG_GATE_SWITCH_magic_6.B.t2 VDD.t78 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X68 Vout INVERTER_MUX_1.OUT.t17 TG_magic_0.B.t35 VSS.t184 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X69 TG_GATE_SWITCH_magic_0.B a_n4297_n2278.t8 A0.t21 VDD.t2 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X70 TG_GATE_SWITCH_magic_0.B a_n4297_n2278.t9 A0.t20 VDD.t3 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X71 TG_magic_4.B a_2061_n4852.t8 TG_magic_7.B.t49 VDD.t12 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X72 TG_GATE_SWITCH_magic_4.B TG_magic_1.CLK TG_magic_2.B.t68 VSS.t99 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X73 TG_GATE_SWITCH_magic_3.B a_n4297_300.t9 A6.t32 VDD.t174 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X74 TG_GATE_SWITCH_magic_6.B a_301_308.t10 TG_magic_0.A.t16 VDD.t79 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X75 a_n4701_n4860# ENA.t2 VDD.t92 VDD.t90 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X76 TG_GATE_SWITCH_magic_2.B S0.t3 TG_magic_2.B.t11 VSS.t6 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X77 TG_magic_7.B a_5741_n4853.t10 Vout.t0 VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X78 TG_GATE_SWITCH_magic_4.B a_3874_n7430.t7 TG_magic_2.B.t13 VDD.t53 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X79 TG_magic_0.A TG_magic_1.CLK TG_GATE_SWITCH_magic_0.B.t33 VSS.t87 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X80 A0 a_n4701_n2278# TG_GATE_SWITCH_magic_0.B.t16 VSS.t59 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X81 TG_magic_5.A a_3817_n991.t7 TG_magic_0.B.t67 VDD.t66 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X82 TG_magic_7.B a_2061_n4852.t9 TG_magic_4.B.t2 VDD.t16 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X83 TG_magic_0.A a_2004_1105.t7 TG_GATE_SWITCH_magic_0.B.t0 VDD.t59 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X84 TG_magic_4.B S0.t4 TG_GATE_SWITCH_magic_5.B.t15 VSS.t129 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X85 A7 a_n1894_n4853.t6 TG_GATE_SWITCH_magic_5.B.t17 VDD.t39 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X86 TG_GATE_SWITCH_magic_2.B a_5684_n6152.t8 TG_magic_2.B.t56 VDD.t288 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X87 A7 a_n2298_n4853# TG_GATE_SWITCH_magic_5.B.t44 VSS.t143 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X88 Vout a_5741_n4853.t11 TG_magic_7.B.t105 VDD.t57 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X89 TG_magic_4.B a_301_n7430.t7 TG_GATE_SWITCH_magic_5.B.t31 VDD.t40 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X90 TG_GATE_SWITCH_magic_0.B a_n4297_n2278.t10 A0.t19 VDD.t3 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X91 TG_magic_0.A a_2061_n2270.t8 TG_magic_0.B.t61 VDD.t15 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X92 TG_GATE_SWITCH_magic_1.B a_2004_n6151.t8 TG_magic_4.B.t15 VDD.t48 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X93 A1 a_n1894_n7431.t6 TG_GATE_SWITCH_magic_4.B.t67 VDD.t85 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X94 TG_GATE_SWITCH_magic_5.B a_n2298_n4853# A7.t18 VSS.t142 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X95 Vout a_5741_n2271.t6 TG_magic_0.B.t46 VDD.t56 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X96 TG_magic_5.A S0.t5 TG_GATE_SWITCH_magic_3.B.t23 VSS.t7 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X97 TG_magic_0.B a_5741_n2271.t7 Vout.t58 VDD.t58 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X98 TG_magic_2.B a_3817_n4055.t7 TG_magic_7.B.t35 VDD.t67 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X99 TG_magic_5.A TG_magic_1.CLK TG_GATE_SWITCH_magic_7.B.t20 VSS.t88 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X100 TG_magic_2.B TG_magic_1.CLK TG_GATE_SWITCH_magic_4.B.t18 VSS.t98 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X101 VSS TG_magic_1.CLK a_2004_1105.t5 VSS.t84 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X102 A7 a_n1894_n4853.t7 TG_GATE_SWITCH_magic_5.B.t29 VDD.t39 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X103 TG_magic_2.B TG_magic_7.CLK TG_magic_7.B.t84 VSS.t224 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X104 A3 a_n4701_n4860# TG_GATE_SWITCH_magic_1.B.t71 VSS.t204 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X105 TG_magic_5.A a_5684_1104.t8 TG_GATE_SWITCH_magic_3.B.t51 VDD.t239 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X106 TG_GATE_SWITCH_magic_6.B a_301_308.t11 TG_magic_0.A.t17 VDD.t80 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X107 VSS S1.t7 a_3817_n991.t5 VSS.t70 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X108 TG_magic_2.B a_3874_n7430.t8 TG_GATE_SWITCH_magic_4.B.t2 VDD.t68 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X109 a_n4701_300# ENA.t3 VSS.t50 VSS.t49 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X110 a_n4701_n7438# ENA.t4 VSS.t52 VSS.t51 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X111 TG_magic_4.B a_2004_n6151.t9 TG_GATE_SWITCH_magic_1.B.t3 VDD.t47 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X112 TG_magic_2.B S0.t8 TG_GATE_SWITCH_magic_2.B.t7 VSS.t8 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X113 TG_GATE_SWITCH_magic_5.B S0.t9 TG_magic_4.B.t66 VSS.t131 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X114 TG_GATE_SWITCH_magic_7.B TG_magic_1.CLK TG_magic_5.A.t14 VSS.t82 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X115 TG_GATE_SWITCH_magic_6.B a_n2298_n2271# A4.t19 VSS.t45 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X116 TG_magic_2.B a_5684_n6152.t9 TG_GATE_SWITCH_magic_2.B.t39 VDD.t289 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X117 TG_GATE_SWITCH_magic_0.B a_n4701_n2278# A0.t34 VSS.t58 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X118 Vout a_5741_n2271.t8 TG_magic_0.B.t99 VDD.t56 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X119 TG_magic_7.B a_3817_n4055.t8 TG_magic_2.B.t61 VDD.t64 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X120 A6 a_n4701_300# TG_GATE_SWITCH_magic_3.B.t14 VSS.t61 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X121 TG_magic_2.B a_5684_n6152.t10 TG_GATE_SWITCH_magic_2.B.t40 VDD.t290 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X122 TG_GATE_SWITCH_magic_5.B a_301_n7430.t8 TG_magic_4.B.t69 VDD.t45 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X123 TG_magic_0.B INVERTER_MUX_1.OUT.t18 Vout.t40 VSS.t10 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X124 A1 a_n1894_n7431.t7 TG_GATE_SWITCH_magic_4.B.t45 VDD.t246 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X125 a_n4701_n2278# ENA.t5 VDD.t93 VDD.t90 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X126 TG_GATE_SWITCH_magic_4.B a_n1894_n7431.t8 A1.t33 VDD.t87 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X127 TG_magic_5.A a_5684_1104.t9 TG_GATE_SWITCH_magic_3.B.t50 VDD.t239 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X128 TG_magic_0.B a_5741_n2271.t9 Vout.t60 VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X129 Vout a_5741_n2271.t10 TG_magic_0.B.t101 VDD.t54 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X130 TG_magic_0.B a_2061_n2270.t9 TG_magic_0.A.t67 VDD.t16 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X131 TG_magic_0.B a_2061_n2270.t10 TG_magic_0.A.t0 VDD.t11 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X132 TG_magic_4.B TG_magic_1.CLK TG_GATE_SWITCH_magic_1.B.t35 VSS.t97 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X133 TG_magic_4.B S0.t10 TG_GATE_SWITCH_magic_5.B.t13 VSS.t114 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X134 TG_GATE_SWITCH_magic_0.B a_2004_1105.t8 TG_magic_0.A.t37 VDD.t102 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X135 a_n4701_n2278# ENA.t6 VSS.t53 VSS.t49 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X136 A4 a_n2298_n2271# TG_GATE_SWITCH_magic_6.B.t56 VSS.t42 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X137 TG_magic_0.B a_3817_n991.t8 TG_magic_5.A.t52 VDD.t65 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X138 Vout a_5741_n2271.t11 TG_magic_0.B.t102 VDD.t57 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X139 A1 a_n2298_n7431# TG_GATE_SWITCH_magic_4.B.t31 VSS.t146 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X140 TG_magic_7.B S1.t8 TG_magic_4.B.t99 VSS.t152 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X141 TG_magic_0.A a_2061_n2270.t11 TG_magic_0.B.t1 VDD.t12 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X142 TG_magic_7.B TG_magic_7.CLK TG_magic_2.B.t105 VSS.t95 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X143 TG_magic_4.B a_2004_n6151.t10 TG_GATE_SWITCH_magic_1.B.t4 VDD.t49 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X144 TG_magic_4.B a_301_n7430.t9 TG_GATE_SWITCH_magic_5.B.t33 VDD.t42 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X145 TG_GATE_SWITCH_magic_1.B a_2004_n6151.t11 TG_magic_4.B.t18 VDD.t48 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X146 A1 a_n1894_n7431.t9 TG_GATE_SWITCH_magic_4.B.t68 VDD.t246 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X147 TG_magic_0.B a_5741_n2271.t12 Vout.t63 VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X148 a_n2298_n4853# ENA.t7 VSS.t55 VSS.t54 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X149 TG_magic_1.CLK S0.t12 VDD.t163 VDD.t23 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X150 A4 a_n1894_n2271.t8 TG_GATE_SWITCH_magic_6.B.t61 VDD.t39 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X151 TG_GATE_SWITCH_magic_7.B a_n1894_307.t7 A2.t22 VDD.t60 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X152 VSS S1.t9 TG_magic_7.CLK VSS.t16 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X153 Vout INVERTER_MUX_1.OUT.t19 TG_magic_0.B.t34 VSS.t0 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X154 TG_GATE_SWITCH_magic_5.B a_n1894_n4853.t8 A7.t8 VDD.t10 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X155 TG_GATE_SWITCH_magic_0.B TG_magic_1.CLK TG_magic_0.A.t53 VSS.t81 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X156 A1 a_n2298_n7431# TG_GATE_SWITCH_magic_4.B.t30 VSS.t143 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X157 TG_magic_5.A a_3817_n991.t9 TG_magic_0.B.t53 VDD.t67 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X158 TG_GATE_SWITCH_magic_3.B a_n4701_300# A6.t10 VSS.t58 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X159 A6 a_n4297_300.t10 TG_GATE_SWITCH_magic_3.B.t28 VDD.t228 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X160 TG_GATE_SWITCH_magic_4.B a_n2298_n7431# A1.t9 VSS.t142 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X161 TG_magic_5.A S0.t13 TG_GATE_SWITCH_magic_3.B.t24 VSS.t15 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X162 TG_magic_5.A TG_magic_1.CLK TG_GATE_SWITCH_magic_7.B.t19 VSS.t80 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X163 TG_magic_0.A TG_magic_7.CLK TG_magic_0.B.t96 VSS.t213 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X164 TG_magic_5.A a_3874_308.t9 TG_GATE_SWITCH_magic_7.B.t58 VDD.t298 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X165 A7 a_n1894_n4853.t9 TG_GATE_SWITCH_magic_5.B.t28 VDD.t8 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X166 VSS TG_magic_7.CLK a_3817_n4055.t5 VSS.t69 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X167 TG_magic_7.B a_3817_n4055.t9 TG_magic_2.B.t62 VDD.t63 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X168 TG_magic_7.B a_2061_n4852.t10 TG_magic_4.B.t24 VDD.t13 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X169 TG_magic_0.B a_3817_n991.t10 TG_magic_5.A.t50 VDD.t64 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X170 TG_GATE_SWITCH_magic_6.B S0.t14 TG_magic_0.A.t62 VSS.t19 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X171 TG_GATE_SWITCH_magic_5.B a_n1894_n4853.t10 A7.t0 VDD.t7 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X172 VSS S0.t15 a_5684_1104.t2 VSS.t10 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X173 A5 a_n4297_n7438.t9 TG_GATE_SWITCH_magic_2.B.t22 VDD.t186 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X174 TG_GATE_SWITCH_magic_2.B S0.t16 TG_magic_2.B.t9 VSS.t20 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X175 TG_magic_2.B a_3817_n4055.t10 TG_magic_7.B.t2 VDD.t62 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X176 TG_GATE_SWITCH_magic_3.B a_5684_1104.t10 TG_magic_5.A.t57 VDD.t238 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X177 TG_GATE_SWITCH_magic_0.B a_2004_1105.t9 TG_magic_0.A.t38 VDD.t103 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X178 TG_magic_0.A a_301_308.t12 TG_GATE_SWITCH_magic_6.B.t5 VDD.t81 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X179 TG_GATE_SWITCH_magic_4.B a_n1894_n7431.t10 A1.t31 VDD.t299 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X180 TG_magic_7.B a_2061_n4852.t11 TG_magic_4.B.t25 VDD.t13 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X181 A3 a_n4297_n4860.t9 TG_GATE_SWITCH_magic_1.B.t56 VDD.t1 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X182 a_n2298_307# ENA.t8 VDD.t94 VDD.t88 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X183 TG_magic_7.B a_3817_n4055.t11 TG_magic_2.B.t15 VDD.t63 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X184 VSS S2.t4 INVERTER_MUX_1.OUT.t14 VSS.t186 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X185 TG_GATE_SWITCH_magic_3.B a_n4297_300.t11 A6.t30 VDD.t171 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X186 A5 a_n4701_n7438# TG_GATE_SWITCH_magic_2.B.t58 VSS.t208 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X187 A0 a_n4701_n2278# TG_GATE_SWITCH_magic_0.B.t15 VSS.t63 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X188 A5 a_n4297_n7438.t10 TG_GATE_SWITCH_magic_2.B.t21 VDD.t186 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X189 TG_magic_0.B TG_magic_7.CLK TG_magic_0.A.t106 VSS.t226 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X190 TG_magic_4.B S1.t10 TG_magic_7.B.t100 VSS.t155 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X191 TG_GATE_SWITCH_magic_7.B a_3874_308.t10 TG_magic_5.A.t103 VDD.t296 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X192 A5 a_n4297_n7438.t11 TG_GATE_SWITCH_magic_2.B.t20 VDD.t240 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X193 TG_magic_7.B S2.t5 Vout.t54 VSS.t29 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X194 TG_GATE_SWITCH_magic_1.B a_n4701_n4860# A3.t33 VSS.t209 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X195 VSS TG_magic_1.CLK a_2004_n6151.t4 VSS.t101 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X196 VDD TG_magic_1.CLK a_2004_1105.t3 VDD.t122 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X197 TG_GATE_SWITCH_magic_0.B a_2004_1105.t10 TG_magic_0.A.t39 VDD.t103 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X198 A3 a_n4297_n4860.t10 TG_GATE_SWITCH_magic_1.B.t55 VDD.t1 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X199 A3 a_n4297_n4860.t11 TG_GATE_SWITCH_magic_1.B.t54 VDD.t19 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X200 TG_magic_7.B S2.t6 Vout.t55 VSS.t30 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X201 TG_GATE_SWITCH_magic_7.B a_3874_308.t11 TG_magic_5.A.t102 VDD.t295 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X202 A4 a_n1894_n2271.t9 TG_GATE_SWITCH_magic_6.B.t62 VDD.t8 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X203 VDD TG_magic_1.CLK a_2004_n6151.t2 VDD.t125 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X204 a_n2298_n7431# ENA.t9 VSS.t56 VSS.t54 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X205 TG_magic_2.B TG_magic_7.CLK TG_magic_7.B.t83 VSS.t221 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X206 A2 a_n1894_307.t8 TG_GATE_SWITCH_magic_7.B.t14 VDD.t106 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X207 TG_GATE_SWITCH_magic_0.B a_2004_1105.t11 TG_magic_0.A.t40 VDD.t69 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X208 TG_magic_7.CLK S1.t11 VDD.t190 VDD.t25 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X209 TG_GATE_SWITCH_magic_6.B a_301_308.t13 TG_magic_0.A.t19 VDD.t82 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X210 TG_GATE_SWITCH_magic_6.B a_n1894_n2271.t10 A4.t31 VDD.t10 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X211 Vout a_5741_n4853.t12 TG_magic_7.B.t106 VDD.t56 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X212 TG_GATE_SWITCH_magic_1.B a_n4297_n4860.t12 A3.t20 VDD.t17 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X213 TG_magic_5.A a_5684_1104.t11 TG_GATE_SWITCH_magic_3.B.t48 VDD.t234 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X214 TG_GATE_SWITCH_magic_6.B a_n1894_n2271.t11 A4.t32 VDD.t7 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X215 TG_GATE_SWITCH_magic_7.B a_n1894_307.t9 A2.t20 VDD.t61 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X216 TG_magic_0.A a_2004_1105.t12 TG_GATE_SWITCH_magic_0.B.t6 VDD.t104 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X217 TG_magic_1.CLK S0.t17 VSS.t134 VSS.t122 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X218 TG_GATE_SWITCH_magic_2.B a_n4701_n7438# A5.t31 VSS.t207 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X219 VDD TG_magic_1.CLK a_2004_1105.t2 VDD.t122 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X220 a_n2298_n4853# ENA.t10 VDD.t96 VDD.t95 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X221 TG_magic_5.A S1.t12 TG_magic_0.B.t39 VSS.t149 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X222 A4 a_n1894_n2271.t12 TG_GATE_SWITCH_magic_6.B.t65 VDD.t8 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X223 TG_GATE_SWITCH_magic_2.B a_n4297_n7438.t12 A5.t17 VDD.t241 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X224 TG_magic_0.B a_2061_n2270.t12 TG_magic_0.A.t2 VDD.t13 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X225 TG_GATE_SWITCH_magic_7.B a_n2298_307# A2.t35 VSS.t45 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X226 TG_magic_0.B a_3817_n991.t11 TG_magic_5.A.t49 VDD.t63 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X227 A2 a_n1894_307.t10 TG_GATE_SWITCH_magic_7.B.t42 VDD.t189 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X228 TG_GATE_SWITCH_magic_1.B a_n4297_n4860.t13 A3.t19 VDD.t17 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X229 TG_GATE_SWITCH_magic_1.B a_n4297_n4860.t14 A3.t18 VDD.t2 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X230 TG_magic_4.B a_2061_n4852.t12 TG_magic_7.B.t24 VDD.t12 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X231 TG_GATE_SWITCH_magic_4.B TG_magic_1.CLK TG_magic_2.B.t67 VSS.t99 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X232 Vout S2.t7 TG_magic_7.B.t75 VSS.t32 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X233 TG_GATE_SWITCH_magic_6.B a_n1894_n2271.t13 A4.t34 VDD.t7 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X234 TG_GATE_SWITCH_magic_7.B a_n1894_307.t11 A2.t18 VDD.t61 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X235 TG_magic_0.A a_2004_1105.t13 TG_GATE_SWITCH_magic_0.B.t7 VDD.t104 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X236 TG_GATE_SWITCH_magic_7.B TG_magic_1.CLK TG_magic_5.A.t12 VSS.t79 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X237 TG_GATE_SWITCH_magic_3.B S0.t18 TG_magic_5.A.t20 VSS.t21 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X238 VDD S1.t13 TG_magic_7.CLK VDD.t27 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X239 A5 a_n4701_n7438# TG_GATE_SWITCH_magic_2.B.t57 VSS.t206 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X240 TG_GATE_SWITCH_magic_1.B a_n4297_n4860.t15 A3.t17 VDD.t3 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X241 TG_GATE_SWITCH_magic_4.B a_3874_n7430.t9 TG_magic_2.B.t95 VDD.t53 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X242 TG_magic_7.B TG_magic_7.CLK TG_magic_2.B.t103 VSS.t219 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X243 TG_magic_4.B a_2061_n4852.t13 TG_magic_7.B.t25 VDD.t15 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X244 TG_magic_7.B a_5741_n4853.t13 Vout.t21 VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X245 TG_magic_0.A a_2004_1105.t14 TG_GATE_SWITCH_magic_0.B.t8 VDD.t59 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X246 TG_magic_5.A a_3817_n991.t12 TG_magic_0.B.t69 VDD.t62 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X247 VDD S0.t19 a_5684_1104.t3 VDD.t156 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X248 TG_GATE_SWITCH_magic_0.B a_n4701_n2278# A0.t32 VSS.t62 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X249 TG_magic_4.B S0.t20 TG_GATE_SWITCH_magic_5.B.t12 VSS.t129 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X250 VSS S0.t21 TG_magic_1.CLK VSS.t125 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X251 TG_GATE_SWITCH_magic_2.B a_5684_n6152.t11 TG_magic_2.B.t53 VDD.t288 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X252 TG_GATE_SWITCH_magic_1.B a_2004_n6151.t12 TG_magic_4.B.t19 VDD.t50 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X253 TG_magic_0.A S0.t22 TG_GATE_SWITCH_magic_6.B.t29 VSS.t137 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X254 TG_magic_7.B a_5741_n4853.t14 Vout.t22 VDD.t58 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X255 A0 a_n4297_n2278.t11 TG_GATE_SWITCH_magic_0.B.t36 VDD.t1 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X256 A0 a_n4297_n2278.t12 TG_GATE_SWITCH_magic_0.B.t37 VDD.t19 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X257 TG_magic_4.B a_301_n7430.t10 TG_GATE_SWITCH_magic_5.B.t18 VDD.t40 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X258 TG_magic_7.B S1.t14 TG_magic_4.B.t98 VSS.t156 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X259 A2 a_n1894_307.t12 TG_GATE_SWITCH_magic_7.B.t44 VDD.t189 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X260 TG_magic_5.A TG_magic_1.CLK TG_GATE_SWITCH_magic_7.B.t18 VSS.t78 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X261 VDD TG_magic_7.CLK a_3817_n4055.t3 VDD.t177 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X262 TG_GATE_SWITCH_magic_7.B a_3874_308.t12 TG_magic_5.A.t101 VDD.t293 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X263 TG_GATE_SWITCH_magic_7.B a_n2298_307# A2.t34 VSS.t44 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X264 TG_magic_0.A a_2061_n2270.t13 TG_magic_0.B.t3 VDD.t14 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X265 TG_magic_0.B INVERTER_MUX_1.OUT.t20 Vout.t38 VSS.t1 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X266 TG_magic_4.B a_2061_n4852.t14 TG_magic_7.B.t26 VDD.t15 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X267 TG_magic_2.B TG_magic_1.CLK TG_GATE_SWITCH_magic_4.B.t16 VSS.t98 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X268 a_n2298_n2271# ENA.t11 VDD.t97 VDD.t95 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X269 TG_GATE_SWITCH_magic_2.B a_n4701_n7438# A5.t29 VSS.t205 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X270 A4 a_n2298_n2271# TG_GATE_SWITCH_magic_6.B.t55 VSS.t40 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X271 TG_magic_7.B a_5741_n4853.t15 Vout.t23 VDD.t58 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X272 TG_magic_2.B a_3874_n7430.t10 TG_GATE_SWITCH_magic_4.B.t46 VDD.t68 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X273 TG_magic_2.B TG_magic_7.CLK TG_magic_7.B.t82 VSS.t218 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X274 A0 a_n4297_n2278.t13 TG_GATE_SWITCH_magic_0.B.t38 VDD.t19 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X275 a_n4701_n7438# ENA.t12 VSS.t57 VSS.t51 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X276 VSS S0.t25 a_5684_n6152.t5 VSS.t29 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X277 A7 a_n2298_n4853# TG_GATE_SWITCH_magic_5.B.t43 VSS.t141 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X278 TG_magic_4.B a_2004_n6151.t13 TG_GATE_SWITCH_magic_1.B.t7 VDD.t51 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X279 TG_magic_7.B a_3817_n4055.t12 TG_magic_2.B.t16 VDD.t64 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X280 TG_magic_2.B a_3874_n7430.t11 TG_GATE_SWITCH_magic_4.B.t47 VDD.t184 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X281 Vout a_5741_n4853.t16 TG_magic_7.B.t42 VDD.t54 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X282 TG_GATE_SWITCH_magic_7.B a_3874_308.t13 TG_magic_5.A.t100 VDD.t293 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X283 Vout a_5741_n2271.t13 TG_magic_0.B.t104 VDD.t56 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X284 a_n4701_n7438# ENA.t13 VDD.t99 VDD.t98 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X285 TG_GATE_SWITCH_magic_0.B a_n4297_n2278.t14 A0.t15 VDD.t17 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X286 TG_GATE_SWITCH_magic_0.B a_n4297_n2278.t15 A0.t14 VDD.t2 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X287 TG_GATE_SWITCH_magic_2.B a_n4297_n7438.t13 A5.t16 VDD.t245 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X288 TG_magic_7.B a_3817_n4055.t13 TG_magic_2.B.t17 VDD.t65 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X289 a_n2298_n2271# ENA.t14 VDD.t100 VDD.t95 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X290 a_n4701_n4860# ENA.t15 VDD.t101 VDD.t90 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X291 TG_magic_7.B a_5741_n4853.t17 Vout.t25 VDD.t55 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X292 TG_GATE_SWITCH_magic_5.B a_301_n7430.t11 TG_magic_4.B.t4 VDD.t41 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X293 TG_GATE_SWITCH_magic_1.B a_2004_n6151.t14 TG_magic_4.B.t21 VDD.t50 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X294 TG_GATE_SWITCH_magic_2.B S0.t26 TG_magic_2.B.t8 VSS.t113 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X295 TG_magic_4.B S0.t27 TG_GATE_SWITCH_magic_5.B.t11 VSS.t114 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X296 TG_magic_4.B TG_magic_1.CLK TG_GATE_SWITCH_magic_1.B.t34 VSS.t97 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X297 TG_magic_5.A a_3874_308.t14 TG_GATE_SWITCH_magic_7.B.t57 VDD.t294 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X298 TG_GATE_SWITCH_magic_0.B a_2004_1105.t15 TG_magic_0.A.t44 VDD.t102 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X299 TG_GATE_SWITCH_magic_3.B a_5684_1104.t12 TG_magic_5.A.t36 VDD.t235 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X300 a_n4701_n2278# ENA.t16 VSS.t172 VSS.t49 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X301 TG_magic_2.B a_3817_n4055.t14 TG_magic_7.B.t6 VDD.t66 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X302 Vout a_5741_n4853.t18 TG_magic_7.B.t44 VDD.t54 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X303 TG_magic_0.A a_2061_n2270.t14 TG_magic_0.B.t4 VDD.t12 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X304 TG_magic_4.B a_301_n7430.t12 TG_GATE_SWITCH_magic_5.B.t20 VDD.t42 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X305 TG_GATE_SWITCH_magic_0.B a_n4297_n2278.t16 A0.t13 VDD.t2 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X306 TG_magic_4.B a_2004_n6151.t15 TG_GATE_SWITCH_magic_1.B.t9 VDD.t49 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X307 TG_GATE_SWITCH_magic_6.B a_n2298_n2271# A4.t18 VSS.t44 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X308 TG_GATE_SWITCH_magic_5.B a_n2298_n4853# A7.t16 VSS.t140 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X309 A6 a_n4297_300.t12 TG_GATE_SWITCH_magic_3.B.t54 VDD.t75 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X310 TG_magic_7.B a_3817_n4055.t15 TG_magic_2.B.t19 VDD.t65 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X311 A1 a_n1894_n7431.t11 TG_GATE_SWITCH_magic_4.B.t70 VDD.t246 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X312 A6 a_n4297_300.t13 TG_GATE_SWITCH_magic_3.B.t59 VDD.t75 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X313 TG_GATE_SWITCH_magic_3.B a_5684_1104.t13 TG_magic_5.A.t37 VDD.t236 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X314 A6 a_n4701_300# TG_GATE_SWITCH_magic_3.B.t13 VSS.t59 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X315 TG_magic_0.A a_2061_n2270.t15 TG_magic_0.B.t5 VDD.t15 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X316 TG_GATE_SWITCH_magic_4.B a_3874_n7430.t12 TG_magic_2.B.t88 VDD.t185 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X317 TG_GATE_SWITCH_magic_0.B a_n4297_n2278.t17 A0.t12 VDD.t3 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X318 TG_magic_0.B a_5741_n2271.t14 Vout.t65 VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X319 TG_GATE_SWITCH_magic_3.B S0.t28 TG_magic_5.A.t16 VSS.t115 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X320 A2 a_n2298_307# TG_GATE_SWITCH_magic_7.B.t7 VSS.t43 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X321 TG_GATE_SWITCH_magic_7.B a_n1894_307.t13 A2.t16 VDD.t60 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X322 TG_magic_2.B a_3817_n4055.t16 TG_magic_7.B.t8 VDD.t67 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X323 TG_magic_5.A a_3874_308.t15 TG_GATE_SWITCH_magic_7.B.t56 VDD.t294 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X324 TG_magic_0.B S1.t15 TG_magic_5.A.t25 VSS.t157 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X325 TG_magic_0.B a_5741_n2271.t15 Vout.t66 VDD.t58 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X326 A2 a_n2298_307# TG_GATE_SWITCH_magic_7.B.t6 VSS.t42 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X327 VDD S1.t16 a_3817_n991.t2 VDD.t177 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X328 TG_magic_0.A S0.t29 TG_GATE_SWITCH_magic_6.B.t24 VSS.t116 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X329 TG_GATE_SWITCH_magic_3.B a_n4701_300# A6.t8 VSS.t62 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X330 TG_magic_4.B a_2004_n6151.t16 TG_GATE_SWITCH_magic_1.B.t10 VDD.t51 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X331 TG_magic_2.B a_3874_n7430.t13 TG_GATE_SWITCH_magic_4.B.t49 VDD.t184 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X332 A6 a_n4297_300.t14 TG_GATE_SWITCH_magic_3.B.t60 VDD.t75 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X333 TG_magic_2.B a_5684_n6152.t12 TG_GATE_SWITCH_magic_2.B.t42 VDD.t291 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X334 TG_GATE_SWITCH_magic_3.B a_n4701_300# A6.t7 VSS.t58 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X335 TG_GATE_SWITCH_magic_5.B a_n2298_n4853# A7.t15 VSS.t139 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X336 a_n4701_n2278# ENA.t17 VDD.t212 VDD.t90 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X337 TG_magic_0.A a_301_308.t14 TG_GATE_SWITCH_magic_6.B.t7 VDD.t78 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X338 TG_GATE_SWITCH_magic_7.B a_n2298_307# A2.t31 VSS.t41 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X339 TG_magic_0.B a_5741_n2271.t16 Vout.t67 VDD.t55 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X340 TG_magic_2.B a_3817_n4055.t17 TG_magic_7.B.t9 VDD.t67 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X341 TG_GATE_SWITCH_magic_5.B a_301_n7430.t13 TG_magic_4.B.t6 VDD.t41 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X342 TG_magic_0.B a_2061_n2270.t16 TG_magic_0.A.t6 VDD.t16 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X343 TG_GATE_SWITCH_magic_5.B a_301_n7430.t14 TG_magic_4.B.t7 VDD.t43 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X344 TG_magic_2.B a_5684_n6152.t13 TG_GATE_SWITCH_magic_2.B.t43 VDD.t290 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X345 TG_magic_5.A a_3874_308.t16 TG_GATE_SWITCH_magic_7.B.t55 VDD.t298 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X346 VDD S0.t30 TG_magic_1.CLK VDD.t147 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X347 A7 a_n1894_n4853.t11 TG_GATE_SWITCH_magic_5.B.t1 VDD.t8 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X348 TG_GATE_SWITCH_magic_3.B a_n4297_300.t15 A6.t26 VDD.t76 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X349 TG_GATE_SWITCH_magic_3.B a_n4297_300.t16 A6.t25 VDD.t76 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X350 TG_magic_5.A a_5684_1104.t14 TG_GATE_SWITCH_magic_3.B.t45 VDD.t237 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X351 TG_GATE_SWITCH_magic_6.B S0.t31 TG_magic_0.A.t59 VSS.t117 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X352 TG_magic_4.B TG_magic_1.CLK TG_GATE_SWITCH_magic_1.B.t33 VSS.t90 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X353 TG_magic_7.B a_2061_n4852.t15 TG_magic_4.B.t43 VDD.t11 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X354 TG_magic_0.B a_3817_n991.t13 TG_magic_5.A.t68 VDD.t64 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X355 Vout a_5741_n2271.t17 TG_magic_0.B.t11 VDD.t54 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X356 a_n2298_n2271# ENA.t18 VSS.t174 VSS.t173 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X357 TG_GATE_SWITCH_magic_5.B a_n1894_n4853.t12 A7.t2 VDD.t7 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X358 TG_magic_4.B a_2004_n6151.t17 TG_GATE_SWITCH_magic_1.B.t11 VDD.t47 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X359 TG_magic_2.B S0.t32 TG_GATE_SWITCH_magic_2.B.t4 VSS.t118 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X360 A1 a_n2298_n7431# TG_GATE_SWITCH_magic_4.B.t29 VSS.t141 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X361 a_n4701_n2278# ENA.t19 VDD.t213 VDD.t90 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X362 TG_magic_0.B a_3817_n991.t14 TG_magic_5.A.t67 VDD.t65 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X363 TG_GATE_SWITCH_magic_4.B a_3874_n7430.t14 TG_magic_2.B.t90 VDD.t185 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X364 TG_magic_0.A a_301_308.t15 TG_GATE_SWITCH_magic_6.B.t8 VDD.t78 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X365 TG_magic_0.B a_5741_n2271.t18 Vout.t9 VDD.t55 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X366 TG_magic_2.B a_3817_n4055.t18 TG_magic_7.B.t10 VDD.t62 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X367 TG_magic_2.B a_5684_n6152.t14 TG_GATE_SWITCH_magic_2.B.t44 VDD.t290 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X368 TG_magic_0.A a_301_308.t16 TG_GATE_SWITCH_magic_6.B.t9 VDD.t81 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X369 TG_GATE_SWITCH_magic_3.B a_n4297_300.t17 A6.t24 VDD.t76 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X370 TG_magic_5.A a_3817_n991.t15 TG_magic_0.B.t64 VDD.t66 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X371 A7 a_n1894_n4853.t13 TG_GATE_SWITCH_magic_5.B.t3 VDD.t9 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X372 A4 a_n2298_n2271# TG_GATE_SWITCH_magic_6.B.t53 VSS.t43 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X373 TG_magic_2.B S0.t33 TG_GATE_SWITCH_magic_2.B.t5 VSS.t37 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X374 TG_GATE_SWITCH_magic_6.B a_301_308.t17 TG_magic_0.A.t23 VDD.t80 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X375 A0 a_n4701_n2278# TG_GATE_SWITCH_magic_0.B.t14 VSS.t63 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X376 TG_GATE_SWITCH_magic_1.B TG_magic_1.CLK TG_magic_4.B.t58 VSS.t83 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X377 TG_magic_0.A TG_magic_1.CLK TG_GATE_SWITCH_magic_0.B.t32 VSS.t71 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X378 TG_GATE_SWITCH_magic_7.B a_3874_308.t17 TG_magic_5.A.t96 VDD.t296 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X379 TG_GATE_SWITCH_magic_5.B a_n1894_n4853.t14 A7.t4 VDD.t10 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X380 TG_GATE_SWITCH_magic_3.B S0.t34 TG_magic_5.A.t17 VSS.t119 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X381 TG_GATE_SWITCH_magic_1.B a_n4701_n4860# A3.t32 VSS.t209 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X382 A1 a_n1894_n7431.t12 TG_GATE_SWITCH_magic_4.B.t71 VDD.t84 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X383 TG_GATE_SWITCH_magic_1.B a_2004_n6151.t18 TG_magic_4.B.t31 VDD.t48 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X384 TG_GATE_SWITCH_magic_4.B a_n2298_n7431# A1.t7 VSS.t140 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X385 TG_magic_5.A a_3817_n991.t16 TG_magic_0.B.t63 VDD.t67 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X386 TG_GATE_SWITCH_magic_5.B a_301_n7430.t15 TG_magic_4.B.t8 VDD.t43 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X387 TG_magic_0.A TG_magic_7.CLK TG_magic_0.B.t94 VSS.t84 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X388 TG_GATE_SWITCH_magic_7.B a_3874_308.t18 TG_magic_5.A.t95 VDD.t295 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X389 a_n4701_300# ENA.t20 VDD.t215 VDD.t214 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X390 TG_magic_7.CLK S1.t17 VDD.t195 VDD.t25 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X391 TG_magic_0.A a_2004_1105.t16 TG_GATE_SWITCH_magic_0.B.t10 VDD.t105 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X392 TG_GATE_SWITCH_magic_4.B a_n1894_n7431.t13 A1.t28 VDD.t86 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X393 TG_GATE_SWITCH_magic_6.B a_301_308.t18 TG_magic_0.A.t24 VDD.t82 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X394 TG_GATE_SWITCH_magic_6.B a_301_308.t19 TG_magic_0.A.t25 VDD.t80 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X395 A3 a_n4701_n4860# TG_GATE_SWITCH_magic_1.B.t68 VSS.t208 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X396 TG_GATE_SWITCH_magic_5.B a_n1894_n4853.t15 A7.t21 VDD.t10 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X397 TG_GATE_SWITCH_magic_5.B a_n1894_n4853.t16 A7.t22 VDD.t206 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X398 a_n2298_n4853# ENA.t21 VDD.t216 VDD.t95 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X399 Vout S2.t10 TG_magic_7.B.t74 VSS.t39 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X400 TG_magic_4.B S1.t18 TG_magic_7.B.t98 VSS.t101 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X401 a_n2298_307# ENA.t22 VSS.t175 VSS.t173 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X402 VDD S0.t37 TG_magic_1.CLK VDD.t152 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X403 A2 a_n1894_307.t14 TG_GATE_SWITCH_magic_7.B.t46 VDD.t187 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X404 TG_magic_1.CLK S0.t38 VSS.t123 VSS.t122 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X405 A4 a_n1894_n2271.t14 TG_GATE_SWITCH_magic_6.B.t67 VDD.t8 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X406 TG_GATE_SWITCH_magic_2.B a_5684_n6152.t15 TG_magic_2.B.t49 VDD.t292 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X407 TG_magic_0.B a_2061_n2270.t17 TG_magic_0.A.t7 VDD.t11 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X408 A4 a_n1894_n2271.t15 TG_GATE_SWITCH_magic_6.B.t32 VDD.t9 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X409 A3 a_n4297_n4860.t16 TG_GATE_SWITCH_magic_1.B.t49 VDD.t18 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X410 TG_magic_0.B INVERTER_MUX_1.OUT.t21 Vout.t37 VSS.t194 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X411 A2 a_n2298_307# TG_GATE_SWITCH_magic_7.B.t5 VSS.t40 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X412 TG_GATE_SWITCH_magic_6.B a_n1894_n2271.t16 A4.t1 VDD.t7 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X413 VDD S1.t19 TG_magic_7.CLK VDD.t27 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X414 TG_GATE_SWITCH_magic_4.B a_n1894_n7431.t14 A1.t27 VDD.t299 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X415 TG_GATE_SWITCH_magic_6.B S0.t40 TG_magic_0.A.t60 VSS.t124 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X416 TG_GATE_SWITCH_magic_7.B TG_magic_1.CLK TG_magic_5.A.t10 VSS.t70 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X417 A5 a_n4701_n7438# TG_GATE_SWITCH_magic_2.B.t56 VSS.t206 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X418 VDD S0.t41 a_5684_1104.t1 VDD.t156 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X419 TG_magic_5.A a_3817_n991.t17 TG_magic_0.B.t62 VDD.t62 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X420 TG_magic_4.B S1.t20 TG_magic_7.B.t97 VSS.t158 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X421 TG_GATE_SWITCH_magic_1.B a_n4701_n4860# A3.t31 VSS.t207 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X422 TG_GATE_SWITCH_magic_0.B a_n4701_n2278# A0.t30 VSS.t62 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X423 A5 a_n4297_n7438.t14 TG_GATE_SWITCH_magic_2.B.t19 VDD.t175 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X424 TG_GATE_SWITCH_magic_4.B a_3874_n7430.t15 TG_magic_2.B.t91 VDD.t183 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X425 TG_GATE_SWITCH_magic_4.B a_n2298_n7431# A1.t6 VSS.t139 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X426 TG_magic_7.B S2.t11 Vout.t1 VSS.t22 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X427 A4 a_n1894_n2271.t17 TG_GATE_SWITCH_magic_6.B.t34 VDD.t9 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X428 A3 a_n4297_n4860.t17 TG_GATE_SWITCH_magic_1.B.t48 VDD.t18 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X429 A3 a_n4297_n4860.t18 TG_GATE_SWITCH_magic_1.B.t47 VDD.t1 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X430 TG_magic_7.CLK S1.t21 VDD.t198 VDD.t34 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X431 VDD TG_magic_7.CLK a_3817_n4055.t2 VDD.t177 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X432 VSS S0.t42 TG_magic_1.CLK VSS.t125 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X433 TG_GATE_SWITCH_magic_4.B a_n1894_n7431.t15 A1.t26 VDD.t299 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X434 TG_magic_1.CLK S0.t43 VDD.t160 VDD.t159 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X435 A3 a_n4297_n4860.t19 TG_GATE_SWITCH_magic_1.B.t46 VDD.t19 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X436 a_n2298_n7431# ENA.t23 VDD.t218 VDD.t217 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X437 TG_GATE_SWITCH_magic_6.B a_n1894_n2271.t18 A4.t3 VDD.t206 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X438 TG_GATE_SWITCH_magic_7.B a_n1894_307.t15 A2.t14 VDD.t188 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X439 TG_magic_1.CLK S0.t44 VSS.t3 VSS.t2 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X440 TG_GATE_SWITCH_magic_6.B a_n1894_n2271.t19 A4.t4 VDD.t10 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X441 TG_GATE_SWITCH_magic_2.B a_n4701_n7438# A5.t27 VSS.t205 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X442 Vout a_5741_n4853.t19 TG_magic_7.B.t45 VDD.t56 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X443 TG_magic_0.A TG_magic_1.CLK TG_GATE_SWITCH_magic_0.B.t31 VSS.t94 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X444 Vout INVERTER_MUX_1.OUT.t24 TG_magic_0.B.t33 VSS.t138 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X445 TG_GATE_SWITCH_magic_2.B a_n4297_n7438.t15 A5.t14 VDD.t176 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X446 TG_magic_5.A S0.t45 TG_GATE_SWITCH_magic_3.B.t0 VSS.t4 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X447 TG_magic_0.B a_2061_n2270.t18 TG_magic_0.A.t8 VDD.t13 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X448 TG_magic_0.B a_3817_n991.t18 TG_magic_5.A.t73 VDD.t63 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X449 TG_GATE_SWITCH_magic_3.B a_5684_1104.t15 TG_magic_5.A.t39 VDD.t238 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X450 A6 a_n4297_300.t18 TG_GATE_SWITCH_magic_3.B.t64 VDD.t77 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X451 TG_GATE_SWITCH_magic_6.B a_n1894_n2271.t20 A4.t5 VDD.t206 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X452 TG_GATE_SWITCH_magic_1.B a_n4297_n4860.t20 A3.t16 VDD.t17 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X453 TG_GATE_SWITCH_magic_2.B a_n4297_n7438.t16 A5.t13 VDD.t245 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X454 TG_GATE_SWITCH_magic_0.B TG_magic_1.CLK TG_magic_0.A.t50 VSS.t93 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X455 A5 a_n4701_n7438# TG_GATE_SWITCH_magic_2.B.t55 VSS.t204 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X456 a_n2298_307# ENA.t24 VDD.t219 VDD.t88 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X457 a_n2298_n2271# ENA.t25 VDD.t220 VDD.t95 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X458 Vout a_5741_n4853.t20 TG_magic_7.B.t46 VDD.t56 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X459 TG_magic_7.B TG_magic_7.CLK TG_magic_2.B.t101 VSS.t225 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X460 TG_magic_4.B a_2061_n4852.t16 TG_magic_7.B.t28 VDD.t12 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X461 TG_magic_5.A a_3874_308.t19 TG_GATE_SWITCH_magic_7.B.t54 VDD.t297 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X462 TG_GATE_SWITCH_magic_1.B a_n4297_n4860.t21 A3.t15 VDD.t2 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X463 TG_magic_7.B a_5741_n4853.t21 Vout.t29 VDD.t55 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X464 TG_GATE_SWITCH_magic_4.B a_3874_n7430.t16 TG_magic_2.B.t92 VDD.t183 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X465 TG_GATE_SWITCH_magic_1.B a_2004_n6151.t19 TG_magic_4.B.t32 VDD.t46 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X466 TG_GATE_SWITCH_magic_3.B a_5684_1104.t16 TG_magic_5.A.t40 VDD.t235 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X467 TG_GATE_SWITCH_magic_6.B a_n2298_n2271# A4.t17 VSS.t41 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X468 TG_magic_2.B a_3817_n4055.t19 TG_magic_7.B.t11 VDD.t66 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X469 TG_magic_7.B a_5741_n4853.t22 Vout.t43 VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X470 a_n4701_n4860# ENA.t26 VSS.t176 VSS.t51 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X471 A0 a_n4297_n2278.t18 TG_GATE_SWITCH_magic_0.B.t43 VDD.t18 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X472 A0 a_n4297_n2278.t19 TG_GATE_SWITCH_magic_0.B.t44 VDD.t1 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X473 A5 a_n4297_n7438.t17 TG_GATE_SWITCH_magic_2.B.t18 VDD.t240 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X474 TG_GATE_SWITCH_magic_3.B a_5684_1104.t17 TG_magic_5.A.t41 VDD.t238 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X475 TG_magic_7.B S1.t22 TG_magic_4.B.t97 VSS.t159 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X476 TG_magic_0.A a_301_308.t20 TG_GATE_SWITCH_magic_6.B.t13 VDD.t83 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X477 TG_GATE_SWITCH_magic_2.B a_n4297_n7438.t18 A5.t11 VDD.t245 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X478 TG_magic_4.B a_301_n7430.t16 TG_GATE_SWITCH_magic_5.B.t24 VDD.t44 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X479 TG_GATE_SWITCH_magic_3.B a_5684_1104.t18 TG_magic_5.A.t42 VDD.t236 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X480 a_n2298_307# ENA.t27 VDD.t221 VDD.t88 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X481 A6 a_n4701_300# TG_GATE_SWITCH_magic_3.B.t12 VSS.t59 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X482 TG_magic_4.B a_2061_n4852.t17 TG_magic_7.B.t29 VDD.t12 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X483 Vout S2.t12 TG_magic_7.B.t72 VSS.t23 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X484 A2 a_n1894_307.t16 TG_GATE_SWITCH_magic_7.B.t27 VDD.t106 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X485 TG_GATE_SWITCH_magic_0.B a_2004_1105.t17 TG_magic_0.A.t87 VDD.t69 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X486 TG_magic_4.B a_2061_n4852.t18 TG_magic_7.B.t30 VDD.t14 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X487 INVERTER_MUX_1.OUT S2.t13 VDD.t26 VDD.t25 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X488 TG_magic_0.B S1.t23 TG_magic_5.A.t26 VSS.t157 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X489 TG_magic_5.A a_5684_1104.t19 TG_GATE_SWITCH_magic_3.B.t40 VDD.t234 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X490 TG_magic_7.B a_5741_n4853.t23 Vout.t44 VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X491 TG_magic_0.A S0.t46 TG_GATE_SWITCH_magic_6.B.t0 VSS.t5 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X492 A0 a_n4297_n2278.t20 TG_GATE_SWITCH_magic_0.B.t45 VDD.t1 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X493 VDD S1.t25 a_3817_n991.t1 VDD.t177 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X494 TG_GATE_SWITCH_magic_3.B a_n4701_300# A6.t5 VSS.t62 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X495 A7 a_n2298_n4853# TG_GATE_SWITCH_magic_5.B.t42 VSS.t146 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X496 TG_magic_2.B a_3874_n7430.t17 TG_GATE_SWITCH_magic_4.B.t53 VDD.t52 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X497 A0 a_n4297_n2278.t21 TG_GATE_SWITCH_magic_0.B.t46 VDD.t19 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X498 TG_GATE_SWITCH_magic_0.B a_n4297_n2278.t22 A0.t7 VDD.t17 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X499 TG_GATE_SWITCH_magic_2.B a_n4297_n7438.t19 A5.t10 VDD.t241 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X500 VDD S0.t47 a_5684_n6152.t2 VDD.t20 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X501 A2 a_n1894_307.t17 TG_GATE_SWITCH_magic_7.B.t28 VDD.t106 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X502 TG_GATE_SWITCH_magic_0.B a_2004_1105.t18 TG_magic_0.A.t88 VDD.t69 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X503 TG_magic_7.CLK S1.t26 VSS.t161 VSS.t122 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X504 INVERTER_MUX_1.OUT S2.t14 VSS.t25 VSS.t24 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X505 Vout a_5741_n2271.t19 TG_magic_0.B.t13 VDD.t56 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X506 TG_magic_7.B a_3817_n4055.t20 TG_magic_2.B.t24 VDD.t64 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X507 TG_GATE_SWITCH_magic_3.B a_n4297_300.t19 A6.t22 VDD.t174 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X508 TG_GATE_SWITCH_magic_6.B a_301_308.t21 TG_magic_0.A.t27 VDD.t79 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X509 TG_magic_5.A a_5684_1104.t20 TG_GATE_SWITCH_magic_3.B.t39 VDD.t234 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X510 A0 a_n4701_n2278# TG_GATE_SWITCH_magic_0.B.t13 VSS.t61 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X511 TG_GATE_SWITCH_magic_1.B a_2004_n6151.t20 TG_magic_4.B.t33 VDD.t46 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X512 a_n4701_n4860# ENA.t28 VDD.t222 VDD.t90 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X513 TG_GATE_SWITCH_magic_2.B S0.t48 TG_magic_2.B.t5 VSS.t6 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X514 TG_magic_4.B TG_magic_1.CLK TG_GATE_SWITCH_magic_1.B.t32 VSS.t90 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X515 TG_magic_5.A a_5684_1104.t21 TG_GATE_SWITCH_magic_3.B.t38 VDD.t237 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X516 TG_magic_7.B a_2061_n4852.t19 TG_magic_4.B.t47 VDD.t11 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X517 VDD S2.t15 INVERTER_MUX_1.OUT.t2 VDD.t27 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X518 TG_magic_0.A a_2004_1105.t19 TG_GATE_SWITCH_magic_0.B.t57 VDD.t59 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X519 TG_GATE_SWITCH_magic_0.B a_n4297_n2278.t23 A0.t6 VDD.t17 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X520 TG_GATE_SWITCH_magic_2.B a_5684_n6152.t16 TG_magic_2.B.t48 VDD.t287 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X521 TG_magic_4.B a_2004_n6151.t21 TG_GATE_SWITCH_magic_1.B.t15 VDD.t47 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X522 TG_GATE_SWITCH_magic_0.B TG_magic_1.CLK TG_magic_0.A.t49 VSS.t89 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X523 A7 a_n2298_n4853# TG_GATE_SWITCH_magic_5.B.t41 VSS.t143 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X524 TG_magic_4.B a_301_n7430.t17 TG_GATE_SWITCH_magic_5.B.t25 VDD.t44 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X525 Vout INVERTER_MUX_1.OUT.t26 TG_magic_0.B.t32 VSS.t184 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X526 TG_magic_0.A a_2061_n2270.t19 TG_magic_0.B.t9 VDD.t15 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X527 TG_magic_7.B a_3817_n4055.t21 TG_magic_2.B.t25 VDD.t64 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X528 TG_GATE_SWITCH_magic_0.B a_n4297_n2278.t24 A0.t5 VDD.t2 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X529 TG_magic_0.B a_5741_n2271.t20 Vout.t11 VDD.t55 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X530 TG_magic_0.A a_2061_n2270.t20 TG_magic_0.B.t10 VDD.t12 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X531 TG_magic_2.B a_5684_n6152.t17 TG_GATE_SWITCH_magic_2.B.t47 VDD.t290 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X532 TG_GATE_SWITCH_magic_5.B a_n2298_n4853# A7.t12 VSS.t142 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X533 VSS S1.t27 TG_magic_7.CLK VSS.t125 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X534 INVERTER_MUX_1.OUT S2.t16 VDD.t30 VDD.t25 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X535 TG_GATE_SWITCH_magic_1.B TG_magic_1.CLK TG_magic_4.B.t56 VSS.t77 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X536 TG_magic_5.A S0.t49 TG_GATE_SWITCH_magic_3.B.t1 VSS.t7 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X537 VSS S2.t17 INVERTER_MUX_1.OUT.t4 VSS.t26 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X538 TG_magic_5.A TG_magic_1.CLK TG_GATE_SWITCH_magic_7.B.t17 VSS.t88 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X539 TG_magic_5.A a_3817_n991.t19 TG_magic_0.B.t70 VDD.t66 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X540 TG_magic_0.B a_5741_n2271.t21 Vout.t12 VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X541 TG_magic_0.A a_2004_1105.t20 TG_GATE_SWITCH_magic_0.B.t58 VDD.t59 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X542 TG_magic_0.A TG_magic_1.CLK TG_GATE_SWITCH_magic_0.B.t30 VSS.t87 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X543 TG_magic_2.B TG_magic_7.CLK TG_magic_7.B.t81 VSS.t224 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X544 VSS TG_magic_1.CLK a_2004_1105.t4 VSS.t84 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X545 A7 a_n1894_n4853.t17 TG_GATE_SWITCH_magic_5.B.t48 VDD.t9 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X546 TG_GATE_SWITCH_magic_1.B a_2004_n6151.t22 TG_magic_4.B.t35 VDD.t50 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X547 TG_magic_2.B a_3874_n7430.t18 TG_GATE_SWITCH_magic_4.B.t54 VDD.t52 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X548 TG_GATE_SWITCH_magic_1.B TG_magic_1.CLK TG_magic_4.B.t55 VSS.t83 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X549 TG_GATE_SWITCH_magic_0.B a_n4701_n2278# A0.t28 VSS.t60 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X550 TG_GATE_SWITCH_magic_7.B TG_magic_1.CLK TG_magic_5.A.t8 VSS.t82 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X551 TG_GATE_SWITCH_magic_1.B a_2004_n6151.t23 TG_magic_4.B.t36 VDD.t48 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X552 TG_GATE_SWITCH_magic_6.B a_n2298_n2271# A4.t16 VSS.t45 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X553 TG_magic_0.A a_2061_n2270.t21 TG_magic_0.B.t77 VDD.t14 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X554 a_n4701_n7438# ENA.t29 VDD.t223 VDD.t98 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X555 TG_magic_0.A TG_magic_7.CLK TG_magic_0.B.t93 VSS.t84 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X556 TG_GATE_SWITCH_magic_5.B a_301_n7430.t18 TG_magic_4.B.t11 VDD.t45 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X557 TG_magic_2.B a_5684_n6152.t18 TG_GATE_SWITCH_magic_2.B.t48 VDD.t291 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X558 TG_magic_0.A a_2004_1105.t21 TG_GATE_SWITCH_magic_0.B.t59 VDD.t105 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X559 TG_magic_5.A a_5684_1104.t22 TG_GATE_SWITCH_magic_3.B.t37 VDD.t239 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X560 VDD S2.t19 INVERTER_MUX_1.OUT.t5 VDD.t27 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X561 TG_magic_4.B TG_magic_1.CLK TG_GATE_SWITCH_magic_1.B.t31 VSS.t76 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X562 TG_magic_7.B a_2061_n4852.t20 TG_magic_4.B.t48 VDD.t16 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X563 TG_magic_2.B TG_magic_1.CLK TG_GATE_SWITCH_magic_4.B.t15 VSS.t75 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X564 A3 a_n4701_n4860# TG_GATE_SWITCH_magic_1.B.t66 VSS.t208 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X565 A7 a_n1894_n4853.t18 TG_GATE_SWITCH_magic_5.B.t49 VDD.t8 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X566 A4 a_n2298_n2271# TG_GATE_SWITCH_magic_6.B.t50 VSS.t42 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X567 TG_GATE_SWITCH_magic_5.B a_n1894_n4853.t19 A7.t25 VDD.t206 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X568 TG_magic_4.B a_2004_n6151.t24 TG_GATE_SWITCH_magic_1.B.t18 VDD.t51 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X569 TG_GATE_SWITCH_magic_0.B a_2004_1105.t22 TG_magic_0.A.t92 VDD.t102 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X570 TG_magic_5.A S1.t28 TG_magic_0.B.t42 VSS.t164 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X571 Vout a_5741_n4853.t24 TG_magic_7.B.t52 VDD.t57 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X572 TG_magic_2.B a_3874_n7430.t19 TG_GATE_SWITCH_magic_4.B.t34 VDD.t184 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X573 A1 a_n2298_n7431# TG_GATE_SWITCH_magic_4.B.t28 VSS.t146 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X574 TG_magic_2.B S0.t50 TG_GATE_SWITCH_magic_2.B.t1 VSS.t8 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X575 TG_magic_0.B a_3817_n991.t20 TG_magic_5.A.t60 VDD.t64 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X576 TG_magic_0.B a_3817_n991.t21 TG_magic_5.A.t78 VDD.t65 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X577 TG_GATE_SWITCH_magic_5.B S0.t51 TG_magic_4.B.t0 VSS.t9 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X578 TG_GATE_SWITCH_magic_5.B a_n1894_n4853.t20 A7.t26 VDD.t7 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X579 A1 a_n1894_n7431.t16 TG_GATE_SWITCH_magic_4.B.t59 VDD.t85 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X580 TG_magic_2.B a_5684_n6152.t19 TG_GATE_SWITCH_magic_2.B.t49 VDD.t291 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X581 A2 a_n1894_307.t18 TG_GATE_SWITCH_magic_7.B.t29 VDD.t187 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X582 TG_magic_0.B INVERTER_MUX_1.OUT.t27 Vout.t34 VSS.t10 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X583 a_n4701_n2278# ENA.t30 VDD.t224 VDD.t90 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X584 TG_magic_5.A S1.t29 TG_magic_0.B.t43 VSS.t165 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X585 TG_GATE_SWITCH_magic_5.B a_301_n7430.t19 TG_magic_4.B.t12 VDD.t41 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X586 a_n2298_n4853# ENA.t31 VSS.t177 VSS.t54 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X587 TG_magic_2.B a_3817_n4055.t22 TG_magic_7.B.t14 VDD.t62 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X588 TG_magic_0.B a_2061_n2270.t22 TG_magic_0.A.t79 VDD.t11 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X589 A7 a_n1894_n4853.t21 TG_GATE_SWITCH_magic_5.B.t52 VDD.t39 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X590 A7 a_n1894_n4853.t22 TG_GATE_SWITCH_magic_5.B.t53 VDD.t8 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X591 TG_GATE_SWITCH_magic_7.B a_n1894_307.t19 A2.t10 VDD.t60 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X592 TG_GATE_SWITCH_magic_0.B a_2004_1105.t23 TG_magic_0.A.t93 VDD.t102 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X593 TG_GATE_SWITCH_magic_4.B TG_magic_1.CLK TG_magic_2.B.t66 VSS.t73 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X594 TG_magic_7.B S1.t31 TG_magic_4.B.t96 VSS.t152 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X595 TG_GATE_SWITCH_magic_5.B a_n1894_n4853.t23 A7.t29 VDD.t7 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X596 TG_magic_7.B TG_magic_7.CLK TG_magic_2.B.t99 VSS.t95 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X597 TG_GATE_SWITCH_magic_1.B a_n4701_n4860# A3.t30 VSS.t207 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X598 TG_GATE_SWITCH_magic_0.B TG_magic_1.CLK TG_magic_0.A.t47 VSS.t81 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X599 TG_magic_2.B a_5684_n6152.t20 TG_GATE_SWITCH_magic_2.B.t50 VDD.t289 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X600 TG_GATE_SWITCH_magic_4.B a_3874_n7430.t20 TG_magic_2.B.t77 VDD.t185 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X601 TG_magic_5.A a_3817_n991.t22 TG_magic_0.B.t75 VDD.t67 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X602 TG_magic_2.B a_3817_n4055.t23 TG_magic_7.B.t15 VDD.t62 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X603 TG_magic_0.A TG_magic_7.CLK TG_magic_0.B.t92 VSS.t217 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X604 TG_GATE_SWITCH_magic_5.B a_301_n7430.t20 TG_magic_4.B.t84 VDD.t45 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X605 TG_magic_1.CLK S0.t52 VDD.t24 VDD.t23 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X606 TG_magic_0.B S1.t32 TG_magic_5.A.t29 VSS.t91 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X607 A4 a_n1894_n2271.t21 TG_GATE_SWITCH_magic_6.B.t38 VDD.t9 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X608 A6 a_n4297_300.t20 TG_GATE_SWITCH_magic_3.B.t66 VDD.t228 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X609 A6 a_n4297_300.t21 TG_GATE_SWITCH_magic_3.B.t67 VDD.t228 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X610 TG_magic_7.CLK S1.t33 VDD.t202 VDD.t34 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X611 TG_GATE_SWITCH_magic_4.B a_n1894_n7431.t17 A1.t24 VDD.t87 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X612 A1 a_n1894_n7431.t18 TG_GATE_SWITCH_magic_4.B.t61 VDD.t84 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X613 TG_GATE_SWITCH_magic_7.B a_n1894_307.t20 A2.t9 VDD.t60 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X614 TG_GATE_SWITCH_magic_4.B a_n1894_n7431.t19 A1.t22 VDD.t299 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X615 TG_magic_5.A a_3874_308.t20 TG_GATE_SWITCH_magic_7.B.t53 VDD.t298 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X616 TG_GATE_SWITCH_magic_7.B a_n1894_307.t21 A2.t8 VDD.t188 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X617 TG_GATE_SWITCH_magic_4.B a_n1894_n7431.t20 A1.t21 VDD.t86 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X618 A3 a_n4701_n4860# TG_GATE_SWITCH_magic_1.B.t64 VSS.t206 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X619 TG_magic_0.B S1.t34 TG_magic_5.A.t30 VSS.t166 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X620 Vout INVERTER_MUX_1.OUT.t28 TG_magic_0.B.t31 VSS.t0 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X621 VSS TG_magic_7.CLK a_3817_n4055.t4 VSS.t69 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X622 Vout a_5741_n2271.t22 TG_magic_0.B.t16 VDD.t57 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X623 A1 a_n2298_n7431# TG_GATE_SWITCH_magic_4.B.t27 VSS.t143 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X624 VSS S0.t53 a_5684_1104.t0 VSS.t10 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X625 TG_GATE_SWITCH_magic_5.B S0.t54 TG_magic_4.B.t1 VSS.t13 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X626 VDD S1.t35 TG_magic_7.CLK VDD.t203 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X627 A6 a_n4297_300.t22 TG_GATE_SWITCH_magic_3.B.t68 VDD.t228 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X628 TG_magic_1.CLK S0.t55 VSS.t14 VSS.t2 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X629 a_n2298_n4853# ENA.t32 VDD.t225 VDD.t95 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X630 A1 a_n1894_n7431.t21 TG_GATE_SWITCH_magic_4.B.t64 VDD.t84 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X631 TG_GATE_SWITCH_magic_4.B a_n2298_n7431# A1.t3 VSS.t142 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X632 TG_magic_5.A S0.t56 TG_GATE_SWITCH_magic_3.B.t2 VSS.t15 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X633 TG_magic_0.B a_2061_n2270.t23 TG_magic_0.A.t80 VDD.t16 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X634 TG_magic_5.A TG_magic_1.CLK TG_GATE_SWITCH_magic_7.B.t16 VSS.t80 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X635 TG_GATE_SWITCH_magic_5.B a_301_n7430.t21 TG_magic_4.B.t85 VDD.t43 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X636 VSS S0.t57 TG_magic_1.CLK VSS.t16 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X637 A4 a_n1894_n2271.t22 TG_GATE_SWITCH_magic_6.B.t39 VDD.t8 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X638 A4 a_n1894_n2271.t23 TG_GATE_SWITCH_magic_6.B.t40 VDD.t39 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X639 TG_GATE_SWITCH_magic_2.B a_5684_n6152.t21 TG_magic_2.B.t43 VDD.t292 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X640 TG_magic_5.A a_3874_308.t21 TG_GATE_SWITCH_magic_7.B.t52 VDD.t298 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X641 TG_GATE_SWITCH_magic_6.B a_n1894_n2271.t24 A4.t9 VDD.t206 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X642 TG_GATE_SWITCH_magic_4.B a_n1894_n7431.t22 A1.t19 VDD.t86 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X643 TG_magic_0.A a_301_308.t22 TG_GATE_SWITCH_magic_6.B.t15 VDD.t81 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X644 A5 a_n4701_n7438# TG_GATE_SWITCH_magic_2.B.t54 VSS.t204 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X645 TG_magic_0.B TG_magic_7.CLK TG_magic_0.A.t105 VSS.t216 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X646 Vout a_5741_n2271.t23 TG_magic_0.B.t17 VDD.t57 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X647 TG_magic_5.A a_3874_308.t22 TG_GATE_SWITCH_magic_7.B.t51 VDD.t297 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X648 TG_GATE_SWITCH_magic_6.B S0.t58 TG_magic_0.A.t12 VSS.t19 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X649 TG_GATE_SWITCH_magic_3.B a_n4297_300.t23 A6.t18 VDD.t171 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X650 TG_GATE_SWITCH_magic_6.B a_n1894_n2271.t25 A4.t10 VDD.t7 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X651 TG_GATE_SWITCH_magic_3.B a_n4297_300.t24 A6.t17 VDD.t171 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X652 A5 a_n4297_n7438.t20 TG_GATE_SWITCH_magic_2.B.t17 VDD.t186 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X653 TG_GATE_SWITCH_magic_1.B a_n4701_n4860# A3.t29 VSS.t205 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X654 TG_magic_7.CLK S1.t36 VSS.t167 VSS.t122 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X655 TG_GATE_SWITCH_magic_2.B S0.t59 TG_magic_2.B.t3 VSS.t20 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X656 a_n2298_n4853# ENA.t33 VDD.t226 VDD.t95 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X657 a_n4701_n4860# ENA.t34 VSS.t178 VSS.t51 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X658 TG_GATE_SWITCH_magic_7.B a_3874_308.t23 TG_magic_5.A.t90 VDD.t296 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X659 TG_magic_0.B TG_magic_7.CLK TG_magic_0.A.t104 VSS.t215 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X660 TG_magic_5.A a_3817_n991.t23 TG_magic_0.B.t73 VDD.t62 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X661 A3 a_n4297_n4860.t22 TG_GATE_SWITCH_magic_1.B.t43 VDD.t18 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X662 A5 a_n4297_n7438.t21 TG_GATE_SWITCH_magic_2.B.t16 VDD.t240 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X663 TG_magic_7.B S2.t20 Vout.t3 VSS.t29 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X664 TG_GATE_SWITCH_magic_0.B a_2004_1105.t24 TG_magic_0.A.t94 VDD.t103 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X665 A4 a_n1894_n2271.t26 TG_GATE_SWITCH_magic_6.B.t43 VDD.t39 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X666 TG_GATE_SWITCH_magic_2.B a_5684_n6152.t22 TG_magic_2.B.t42 VDD.t292 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X667 TG_magic_0.A a_301_308.t23 TG_GATE_SWITCH_magic_6.B.t16 VDD.t83 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X668 TG_magic_0.A a_301_308.t24 TG_GATE_SWITCH_magic_6.B.t17 VDD.t81 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X669 A3 a_n4297_n4860.t23 TG_GATE_SWITCH_magic_1.B.t42 VDD.t1 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X670 TG_magic_2.B TG_magic_7.CLK TG_magic_7.B.t80 VSS.t221 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X671 TG_GATE_SWITCH_magic_7.B a_3874_308.t24 TG_magic_5.A.t89 VDD.t295 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X672 VDD TG_magic_1.CLK a_2004_n6151.t1 VDD.t125 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X673 VDD TG_magic_7.CLK a_3817_n4055.t1 VDD.t177 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X674 TG_GATE_SWITCH_magic_6.B a_301_308.t25 TG_magic_0.A.t31 VDD.t82 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X675 TG_GATE_SWITCH_magic_3.B a_n4297_300.t25 A6.t16 VDD.t171 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X676 TG_magic_4.B a_2061_n4852.t21 TG_magic_7.B.t33 VDD.t14 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X677 a_n2298_n7431# ENA.t35 VDD.t227 VDD.t217 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X678 TG_GATE_SWITCH_magic_7.B a_3874_308.t25 TG_magic_5.A.t88 VDD.t296 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X679 TG_magic_4.B S1.t37 TG_magic_7.B.t94 VSS.t155 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X680 A5 a_n4297_n7438.t22 TG_GATE_SWITCH_magic_2.B.t15 VDD.t240 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X681 VDD TG_magic_1.CLK a_2004_1105.t1 VDD.t122 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X682 VSS S1.t38 TG_magic_7.CLK VSS.t125 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X683 TG_magic_7.B S2.t21 Vout.t4 VSS.t30 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X684 a_n2298_n7431# ENA.t36 VSS.t179 VSS.t54 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X685 TG_GATE_SWITCH_magic_7.B a_3874_308.t26 TG_magic_5.A.t87 VDD.t295 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X686 VDD TG_magic_7.CLK a_3817_n4055.t0 VDD.t177 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X687 TG_GATE_SWITCH_magic_2.B a_n4297_n7438.t23 A5.t6 VDD.t241 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X688 TG_GATE_SWITCH_magic_6.B a_301_308.t26 TG_magic_0.A.t32 VDD.t82 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X689 A6 a_n4701_300# TG_GATE_SWITCH_magic_3.B.t11 VSS.t63 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X690 TG_magic_7.B a_2061_n4852.t22 TG_magic_4.B.t73 VDD.t13 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X691 TG_magic_7.B a_3817_n4055.t24 TG_magic_2.B.t29 VDD.t63 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X692 a_n2298_n7431# ENA.t37 VDD.t305 VDD.t217 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X693 TG_GATE_SWITCH_magic_1.B a_n4297_n4860.t24 A3.t14 VDD.t17 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X694 TG_GATE_SWITCH_magic_6.B a_301_308.t27 TG_magic_0.A.t33 VDD.t79 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X695 TG_GATE_SWITCH_magic_7.B a_n1894_307.t22 A2.t7 VDD.t61 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X696 TG_magic_0.A a_2004_1105.t25 TG_GATE_SWITCH_magic_0.B.t63 VDD.t104 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X697 TG_GATE_SWITCH_magic_3.B S0.t60 TG_magic_5.A.t3 VSS.t21 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X698 A0 a_n4701_n2278# TG_GATE_SWITCH_magic_0.B.t12 VSS.t61 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X699 TG_GATE_SWITCH_magic_7.B TG_magic_1.CLK TG_magic_5.A.t6 VSS.t79 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X700 a_n2298_n2271# ENA.t38 VDD.t306 VDD.t95 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X701 TG_GATE_SWITCH_magic_1.B a_n4297_n4860.t25 A3.t13 VDD.t3 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X702 TG_GATE_SWITCH_magic_4.B a_3874_n7430.t21 TG_magic_2.B.t78 VDD.t53 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X703 TG_magic_7.B a_5741_n4853.t25 Vout.t46 VDD.t55 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X704 INVERTER_MUX_1.OUT S2.t22 VSS.t31 VSS.t24 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X705 VDD S0.t61 a_5684_1104.t4 VDD.t156 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X706 TG_GATE_SWITCH_magic_3.B a_n4701_300# A6.t3 VSS.t60 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X707 A0 a_n4297_n2278.t25 TG_GATE_SWITCH_magic_0.B.t67 VDD.t18 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X708 A5 a_n4297_n7438.t24 TG_GATE_SWITCH_magic_2.B.t14 VDD.t175 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X709 TG_magic_0.A S0.t62 TG_GATE_SWITCH_magic_6.B.t69 VSS.t137 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X710 TG_GATE_SWITCH_magic_2.B a_n4297_n7438.t25 A5.t4 VDD.t241 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X711 TG_magic_2.B a_3817_n4055.t25 TG_magic_7.B.t17 VDD.t66 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X712 TG_magic_7.B S1.t39 TG_magic_4.B.t95 VSS.t156 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X713 TG_magic_5.A TG_magic_1.CLK TG_GATE_SWITCH_magic_7.B.t15 VSS.t78 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X714 TG_GATE_SWITCH_magic_7.B a_n2298_307# A2.t29 VSS.t45 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X715 VDD TG_magic_1.CLK a_2004_n6151.t0 VDD.t125 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X716 TG_magic_4.B a_301_n7430.t22 TG_GATE_SWITCH_magic_5.B.t59 VDD.t40 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X717 Vout S2.t23 TG_magic_7.B.t69 VSS.t32 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X718 A2 a_n1894_307.t23 TG_GATE_SWITCH_magic_7.B.t34 VDD.t189 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X719 TG_GATE_SWITCH_magic_7.B a_n2298_307# A2.t28 VSS.t44 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X720 TG_GATE_SWITCH_magic_1.B TG_magic_1.CLK TG_magic_4.B.t53 VSS.t77 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X721 INVERTER_MUX_1.OUT S2.t24 VDD.t35 VDD.t34 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X722 TG_GATE_SWITCH_magic_4.B TG_magic_1.CLK TG_magic_2.B.t65 VSS.t69 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X723 TG_magic_0.B INVERTER_MUX_1.OUT.t30 Vout.t32 VSS.t1 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X724 TG_GATE_SWITCH_magic_1.B a_n4297_n4860.t26 A3.t12 VDD.t3 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X725 TG_magic_7.B a_5741_n4853.t26 Vout.t47 VDD.t55 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X726 TG_magic_7.B TG_magic_7.CLK TG_magic_2.B.t97 VSS.t219 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X727 VDD S0.t63 a_5684_1104.t5 VDD.t156 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X728 A0 a_n4297_n2278.t26 TG_GATE_SWITCH_magic_0.B.t68 VDD.t18 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X729 TG_GATE_SWITCH_magic_1.B a_2004_n6151.t25 TG_magic_4.B.t38 VDD.t50 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X730 TG_GATE_SWITCH_magic_4.B a_3874_n7430.t22 TG_magic_2.B.t79 VDD.t183 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X731 TG_magic_2.B a_3817_n4055.t26 TG_magic_7.B.t18 VDD.t66 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X732 TG_magic_2.B a_3874_n7430.t23 TG_GATE_SWITCH_magic_4.B.t38 VDD.t68 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X733 TG_GATE_SWITCH_magic_0.B a_n4701_n2278# A0.t26 VSS.t60 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X734 VSS S2.t25 INVERTER_MUX_1.OUT.t8 VSS.t26 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X735 A0 a_n4297_n2278.t27 TG_GATE_SWITCH_magic_0.B.t69 VDD.t1 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X736 VDD S1.t40 a_3817_n991.t0 VDD.t177 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X737 TG_magic_7.CLK S1.t41 VSS.t180 VSS.t2 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X738 TG_GATE_SWITCH_magic_2.B a_n4297_n7438.t26 A5.t3 VDD.t176 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X739 A7 a_n2298_n4853# TG_GATE_SWITCH_magic_5.B.t40 VSS.t141 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X740 TG_magic_0.A a_2061_n2270.t24 TG_magic_0.B.t80 VDD.t14 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X741 a_n4701_n7438# ENA.t39 VDD.t307 VDD.t98 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X742 INVERTER_MUX_1.OUT S2.t26 VSS.t36 VSS.t35 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X743 TG_GATE_SWITCH_magic_7.B a_3874_308.t27 TG_magic_5.A.t86 VDD.t293 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X744 VDD S0.t65 a_5684_n6152.t1 VDD.t20 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X745 TG_magic_5.A a_5684_1104.t23 TG_GATE_SWITCH_magic_3.B.t36 VDD.t239 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X746 A4 a_n2298_n2271# TG_GATE_SWITCH_magic_6.B.t49 VSS.t40 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X747 TG_GATE_SWITCH_magic_4.B a_3874_n7430.t24 TG_magic_2.B.t81 VDD.t53 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X748 TG_magic_4.B TG_magic_1.CLK TG_GATE_SWITCH_magic_1.B.t30 VSS.t76 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X749 TG_magic_7.B a_2061_n4852.t23 TG_magic_4.B.t74 VDD.t16 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X750 TG_magic_2.B TG_magic_1.CLK TG_GATE_SWITCH_magic_4.B.t12 VSS.t75 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X751 TG_magic_2.B TG_magic_7.CLK TG_magic_7.B.t79 VSS.t218 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X752 TG_GATE_SWITCH_magic_2.B a_5684_n6152.t23 TG_magic_2.B.t41 VDD.t288 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X753 TG_GATE_SWITCH_magic_2.B a_n4701_n7438# A5.t24 VSS.t209 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X754 TG_magic_4.B a_2004_n6151.t26 TG_GATE_SWITCH_magic_1.B.t20 VDD.t51 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X755 VSS S0.t66 a_5684_n6152.t4 VSS.t29 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X756 TG_GATE_SWITCH_magic_3.B a_5684_1104.t24 TG_magic_5.A.t48 VDD.t235 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X757 TG_magic_5.A S1.t42 TG_magic_0.B.t47 VSS.t164 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X758 TG_magic_0.B a_2061_n2270.t25 TG_magic_0.A.t82 VDD.t13 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X759 TG_magic_2.B a_3874_n7430.t25 TG_GATE_SWITCH_magic_4.B.t40 VDD.t184 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X760 TG_magic_7.B a_2061_n4852.t24 TG_magic_4.B.t75 VDD.t11 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X761 Vout a_5741_n4853.t27 TG_magic_7.B.t55 VDD.t57 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X762 TG_magic_0.B a_3817_n991.t24 TG_magic_5.A.t23 VDD.t63 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X763 TG_magic_4.B a_301_n7430.t23 TG_GATE_SWITCH_magic_5.B.t60 VDD.t40 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X764 a_n4701_n7438# ENA.t40 VDD.t308 VDD.t98 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X765 TG_magic_0.A a_2061_n2270.t26 TG_magic_0.B.t82 VDD.t12 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X766 TG_magic_4.B a_301_n7430.t24 TG_GATE_SWITCH_magic_5.B.t61 VDD.t42 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X767 TG_GATE_SWITCH_magic_2.B a_5684_n6152.t24 TG_magic_2.B.t40 VDD.t287 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X768 TG_GATE_SWITCH_magic_5.B S0.t67 TG_magic_4.B.t81 VSS.t9 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X769 TG_GATE_SWITCH_magic_0.B a_n4297_n2278.t28 A0.t1 VDD.t17 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X770 TG_magic_2.B a_5684_n6152.t25 TG_GATE_SWITCH_magic_2.B.t67 VDD.t291 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X771 TG_magic_4.B a_2004_n6151.t27 TG_GATE_SWITCH_magic_1.B.t21 VDD.t49 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X772 VDD S0.t68 a_5684_n6152.t0 VDD.t20 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X773 TG_GATE_SWITCH_magic_5.B a_n2298_n4853# A7.t10 VSS.t140 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X774 TG_magic_5.A S1.t43 TG_magic_0.B.t48 VSS.t165 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X775 TG_magic_4.B a_2061_n4852.t25 TG_magic_7.B.t63 VDD.t15 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X776 INVERTER_MUX_1.OUT S2.t28 VDD.t36 VDD.t34 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X777 TG_GATE_SWITCH_magic_1.B TG_magic_1.CLK TG_magic_4.B.t51 VSS.t74 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X778 TG_GATE_SWITCH_magic_3.B a_5684_1104.t25 TG_magic_5.A.t79 VDD.t236 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X779 TG_GATE_SWITCH_magic_0.B a_n4297_n2278.t29 A0.t0 VDD.t3 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X780 TG_magic_0.B a_5741_n2271.t24 Vout.t15 VDD.t55 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X781 TG_GATE_SWITCH_magic_5.B a_301_n7430.t25 TG_magic_4.B.t89 VDD.t41 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X782 A7 a_n1894_n4853.t24 TG_GATE_SWITCH_magic_5.B.t55 VDD.t39 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X783 A2 a_n2298_307# TG_GATE_SWITCH_magic_7.B.t4 VSS.t43 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X784 TG_GATE_SWITCH_magic_1.B a_2004_n6151.t28 TG_magic_4.B.t41 VDD.t46 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X785 TG_GATE_SWITCH_magic_2.B S0.t69 TG_magic_2.B.t2 VSS.t113 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X786 TG_magic_5.A a_3874_308.t28 TG_GATE_SWITCH_magic_7.B.t50 VDD.t294 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X787 TG_magic_7.B a_5741_n4853.t28 Vout.t49 VDD.t58 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X788 TG_GATE_SWITCH_magic_3.B a_5684_1104.t26 TG_magic_5.A.t80 VDD.t235 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X789 TG_magic_5.A a_3817_n991.t25 TG_magic_0.B.t60 VDD.t66 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X790 TG_magic_7.B a_2061_n4852.t26 TG_magic_4.B.t77 VDD.t11 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X791 TG_magic_2.B a_3874_n7430.t26 TG_GATE_SWITCH_magic_4.B.t41 VDD.t68 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X792 TG_magic_4.B S0.t71 TG_GATE_SWITCH_magic_5.B.t7 VSS.t128 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X793 TG_GATE_SWITCH_magic_4.B TG_magic_1.CLK TG_magic_2.B.t64 VSS.t73 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X794 A7 a_n1894_n4853.t25 TG_GATE_SWITCH_magic_5.B.t56 VDD.t9 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X795 TG_GATE_SWITCH_magic_2.B a_5684_n6152.t26 TG_magic_2.B.t38 VDD.t287 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X796 TG_GATE_SWITCH_magic_6.B a_n2298_n2271# A4.t15 VSS.t44 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X797 TG_magic_4.B a_301_n7430.t26 TG_GATE_SWITCH_magic_5.B.t63 VDD.t44 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X798 A6 a_n4297_300.t26 TG_GATE_SWITCH_magic_3.B.t4 VDD.t75 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X799 TG_GATE_SWITCH_magic_4.B a_3874_n7430.t27 TG_magic_2.B.t84 VDD.t185 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X800 TG_GATE_SWITCH_magic_3.B a_5684_1104.t27 TG_magic_5.A.t81 VDD.t236 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X801 TG_magic_0.A TG_magic_7.CLK TG_magic_0.B.t89 VSS.t217 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X802 TG_GATE_SWITCH_magic_3.B S0.t72 TG_magic_5.A.t74 VSS.t115 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X803 TG_magic_0.B S1.t45 TG_magic_5.A.t33 VSS.t91 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X804 TG_magic_2.B TG_magic_1.CLK TG_GATE_SWITCH_magic_4.B.t10 VSS.t72 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X805 A2 a_n2298_307# TG_GATE_SWITCH_magic_7.B.t3 VSS.t42 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X806 A7 a_n1894_n4853.t26 TG_GATE_SWITCH_magic_5.B.t67 VDD.t9 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X807 VDD S0.t73 TG_magic_1.CLK VDD.t147 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X808 A3 a_n4701_n4860# TG_GATE_SWITCH_magic_1.B.t62 VSS.t206 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X809 TG_magic_5.A a_5684_1104.t28 TG_GATE_SWITCH_magic_3.B.t31 VDD.t237 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X810 TG_GATE_SWITCH_magic_6.B S0.t74 TG_magic_0.A.t75 VSS.t117 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X811 TG_magic_0.A S0.t75 TG_GATE_SWITCH_magic_6.B.t71 VSS.t116 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X812 TG_magic_0.B S1.t46 TG_magic_5.A.t34 VSS.t166 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X813 TG_magic_2.B a_3874_n7430.t28 TG_GATE_SWITCH_magic_4.B.t43 VDD.t52 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X814 Vout a_5741_n4853.t29 TG_magic_7.B.t57 VDD.t54 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X815 TG_magic_0.B a_3817_n991.t26 TG_magic_5.A.t61 VDD.t64 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X816 TG_magic_4.B a_301_n7430.t27 TG_GATE_SWITCH_magic_5.B.t64 VDD.t42 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X817 a_n2298_n2271# ENA.t41 VSS.t231 VSS.t173 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X818 TG_magic_4.B a_2004_n6151.t29 TG_GATE_SWITCH_magic_1.B.t23 VDD.t49 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X819 TG_magic_2.B S0.t76 TG_GATE_SWITCH_magic_2.B.t11 VSS.t118 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X820 TG_GATE_SWITCH_magic_5.B S0.t77 TG_magic_4.B.t83 VSS.t13 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X821 TG_GATE_SWITCH_magic_5.B a_n1894_n4853.t27 A7.t33 VDD.t206 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X822 VDD S1.t47 TG_magic_7.CLK VDD.t203 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X823 TG_magic_7.B a_3817_n4055.t27 TG_magic_2.B.t32 VDD.t65 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X824 A1 a_n1894_n7431.t23 TG_GATE_SWITCH_magic_4.B.t66 VDD.t246 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X825 A1 a_n1894_n7431.t24 TG_GATE_SWITCH_magic_4.B.t3 VDD.t84 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X826 TG_GATE_SWITCH_magic_5.B a_n2298_n4853# A7.t9 VSS.t139 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X827 TG_magic_0.A a_301_308.t28 TG_GATE_SWITCH_magic_6.B.t21 VDD.t78 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X828 TG_GATE_SWITCH_magic_7.B a_n2298_307# A2.t25 VSS.t41 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X829 TG_magic_0.B a_2061_n2270.t27 TG_magic_0.A.t84 VDD.t16 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X830 TG_GATE_SWITCH_magic_5.B a_301_n7430.t28 TG_magic_4.B.t92 VDD.t43 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X831 A1 a_n1894_n7431.t25 TG_GATE_SWITCH_magic_4.B.t4 VDD.t85 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X832 TG_GATE_SWITCH_magic_3.B a_n4297_300.t27 A6.t14 VDD.t76 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X833 TG_magic_0.B a_5741_n2271.t25 Vout.t16 VDD.t58 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X834 TG_GATE_SWITCH_magic_4.B a_n1894_n7431.t26 A1.t15 VDD.t86 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X835 TG_magic_5.A a_5684_1104.t29 TG_GATE_SWITCH_magic_3.B.t30 VDD.t237 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X836 TG_magic_0.B a_2061_n2270.t28 TG_magic_0.A.t85 VDD.t11 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X837 A0 a_n4701_n2278# TG_GATE_SWITCH_magic_0.B.t11 VSS.t59 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X838 TG_magic_0.B TG_magic_7.CLK TG_magic_0.A.t103 VSS.t216 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X839 Vout a_5741_n2271.t26 TG_magic_0.B.t20 VDD.t57 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X840 TG_GATE_SWITCH_magic_5.B a_n1894_n4853.t28 A7.t34 VDD.t206 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X841 A4 a_n2298_n2271# TG_GATE_SWITCH_magic_6.B.t47 VSS.t43 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X842 VSS S0.t78 TG_magic_1.CLK VSS.t16 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X843 A1 a_n2298_n7431# TG_GATE_SWITCH_magic_4.B.t26 VSS.t141 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X844 TG_GATE_SWITCH_magic_1.B a_n4701_n4860# A3.t28 VSS.t205 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X845 TG_magic_0.A TG_magic_1.CLK TG_GATE_SWITCH_magic_0.B.t29 VSS.t71 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X846 TG_magic_0.A a_2061_n2270.t29 TG_magic_0.B.t85 VDD.t15 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X847 TG_magic_0.B TG_magic_7.CLK TG_magic_0.A.t102 VSS.t215 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X848 TG_magic_2.B a_5684_n6152.t27 TG_GATE_SWITCH_magic_2.B.t69 VDD.t289 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X849 TG_GATE_SWITCH_magic_0.B a_2004_1105.t26 TG_magic_0.A.t69 VDD.t103 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X850 A4 a_n1894_n2271.t27 TG_GATE_SWITCH_magic_6.B.t44 VDD.t39 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X851 TG_GATE_SWITCH_magic_2.B a_5684_n6152.t28 TG_magic_2.B.t36 VDD.t292 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X852 A1 a_n1894_n7431.t27 TG_GATE_SWITCH_magic_4.B.t6 VDD.t85 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X853 TG_magic_0.B a_5741_n2271.t27 Vout.t18 VDD.t58 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X854 TG_magic_2.B a_3817_n4055.t28 TG_magic_7.B.t20 VDD.t67 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X855 a_n4701_300# ENA.t42 VDD.t309 VDD.t214 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X856 A4 a_n1894_n2271.t28 TG_GATE_SWITCH_magic_6.B.t45 VDD.t9 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X857 a_n4701_300# ENA.t43 VDD.t310 VDD.t214 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X858 A3 a_n4701_n4860# TG_GATE_SWITCH_magic_1.B.t60 VSS.t204 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X859 TG_magic_0.A a_2004_1105.t27 TG_GATE_SWITCH_magic_0.B.t52 VDD.t105 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X860 TG_GATE_SWITCH_magic_4.B a_n1894_n7431.t28 A1.t13 VDD.t87 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X861 TG_GATE_SWITCH_magic_6.B a_301_308.t29 TG_magic_0.A.t35 VDD.t80 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X862 VSS S1.t48 a_3817_n991.t4 VSS.t70 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X863 Vout a_5741_n2271.t28 TG_magic_0.B.t22 VDD.t54 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X864 TG_magic_2.B S0.t79 TG_GATE_SWITCH_magic_2.B.t9 VSS.t37 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X865 a_n4701_300# ENA.t44 VSS.t232 VSS.t49 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X866 TG_GATE_SWITCH_magic_5.B S0.t80 TG_magic_4.B.t80 VSS.t131 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X867 TG_GATE_SWITCH_magic_3.B S0.t81 TG_magic_5.A.t58 VSS.t119 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X868 TG_magic_2.B a_5684_n6152.t29 TG_GATE_SWITCH_magic_2.B.t71 VDD.t289 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X869 VDD TG_magic_1.CLK a_2004_1105.t0 VDD.t122 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X870 TG_GATE_SWITCH_magic_0.B a_n4701_n2278# A0.t24 VSS.t58 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X871 TG_GATE_SWITCH_magic_4.B a_n2298_n7431# A1.t1 VSS.t140 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X872 A6 a_n4701_300# TG_GATE_SWITCH_magic_3.B.t10 VSS.t61 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X873 TG_magic_4.B S1.t49 TG_magic_7.B.t92 VSS.t101 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X874 TG_GATE_SWITCH_magic_5.B a_301_n7430.t29 TG_magic_4.B.t93 VDD.t45 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X875 a_n2298_307# ENA.t45 VSS.t233 VSS.t173 nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X876 A2 a_n1894_307.t24 TG_GATE_SWITCH_magic_7.B.t35 VDD.t187 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X877 a_n4701_300# ENA.t46 VDD.t311 VDD.t214 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X878 TG_magic_0.A a_2004_1105.t28 TG_GATE_SWITCH_magic_0.B.t53 VDD.t105 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X879 TG_GATE_SWITCH_magic_4.B a_n1894_n7431.t29 A1.t12 VDD.t87 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X880 A6 a_n4701_300# TG_GATE_SWITCH_magic_3.B.t9 VSS.t63 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X881 Vout a_5741_n2271.t29 TG_magic_0.B.t23 VDD.t54 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X882 TG_magic_7.B a_2061_n4852.t27 TG_magic_4.B.t78 VDD.t13 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X883 TG_magic_7.B a_3817_n4055.t29 TG_magic_2.B.t34 VDD.t63 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X884 a_n2298_n7431# ENA.t47 VDD.t312 VDD.t217 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X885 A2 a_n2298_307# TG_GATE_SWITCH_magic_7.B.t2 VSS.t40 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X886 TG_GATE_SWITCH_magic_6.B a_n1894_n2271.t29 A4.t14 VDD.t206 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X887 TG_GATE_SWITCH_magic_7.B a_n1894_307.t25 A2.t4 VDD.t61 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X888 TG_magic_0.A a_2004_1105.t29 TG_GATE_SWITCH_magic_0.B.t54 VDD.t104 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X889 TG_GATE_SWITCH_magic_7.B TG_magic_1.CLK TG_magic_5.A.t4 VSS.t70 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X890 TG_magic_7.CLK S1.t50 VSS.t183 VSS.t2 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X891 TG_magic_0.B a_3817_n991.t27 TG_magic_5.A.t62 VDD.t65 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X892 TG_magic_5.A a_3817_n991.t28 TG_magic_0.B.t74 VDD.t62 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X893 Vout S2.t31 TG_magic_7.B.t68 VSS.t39 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X894 VDD S0.t84 TG_magic_1.CLK VDD.t152 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X895 TG_GATE_SWITCH_magic_3.B a_n4701_300# A6.t0 VSS.t60 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X896 A5 a_n4297_n7438.t27 TG_GATE_SWITCH_magic_2.B.t13 VDD.t175 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X897 A2 a_n1894_307.t26 TG_GATE_SWITCH_magic_7.B.t37 VDD.t187 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X898 TG_GATE_SWITCH_magic_4.B a_n2298_n7431# A1.t0 VSS.t139 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X899 A2 a_n1894_307.t27 TG_GATE_SWITCH_magic_7.B.t38 VDD.t189 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X900 A3 a_n4297_n4860.t27 TG_GATE_SWITCH_magic_1.B.t38 VDD.t18 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X901 TG_magic_0.B INVERTER_MUX_1.OUT.t32 Vout.t31 VSS.t194 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X902 TG_GATE_SWITCH_magic_6.B S0.t85 TG_magic_0.A.t68 VSS.t124 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X903 A3 a_n4297_n4860.t28 TG_GATE_SWITCH_magic_1.B.t37 VDD.t19 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X904 TG_GATE_SWITCH_magic_4.B TG_magic_1.CLK TG_magic_2.B.t63 VSS.t69 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X905 TG_GATE_SWITCH_magic_7.B a_n1894_307.t28 A2.t1 VDD.t188 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X906 TG_GATE_SWITCH_magic_5.B a_n1894_n4853.t29 A7.t35 VDD.t10 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X907 TG_magic_4.B S1.t51 TG_magic_7.B.t91 VSS.t158 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X908 A5 a_n4297_n7438.t28 TG_GATE_SWITCH_magic_2.B.t12 VDD.t175 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X909 TG_magic_4.B a_2061_n4852.t28 TG_magic_7.B.t66 VDD.t14 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X910 TG_magic_5.A a_3817_n991.t29 TG_magic_0.B.t24 VDD.t67 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X911 TG_GATE_SWITCH_magic_4.B a_3874_n7430.t29 TG_magic_2.B.t75 VDD.t183 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X912 TG_magic_7.B S2.t32 Vout.t7 VSS.t22 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X913 TG_GATE_SWITCH_magic_2.B a_n4297_n7438.t29 A5.t0 VDD.t176 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X914 TG_magic_5.A S0.t86 TG_GATE_SWITCH_magic_3.B.t56 VSS.t4 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X915 TG_magic_0.A TG_magic_7.CLK TG_magic_0.B.t86 VSS.t213 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X916 VDD S2.t33 INVERTER_MUX_1.OUT.t15 VDD.t203 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X917 TG_GATE_SWITCH_magic_7.B a_3874_308.t29 TG_magic_5.A.t84 VDD.t293 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X918 A3 a_n4297_n4860.t29 TG_GATE_SWITCH_magic_1.B.t36 VDD.t19 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X919 A6 a_n4297_300.t28 TG_GATE_SWITCH_magic_3.B.t6 VDD.t77 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X920 TG_magic_1.CLK S0.t87 VDD.t252 VDD.t159 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X921 A6 a_n4297_300.t29 TG_GATE_SWITCH_magic_3.B.t7 VDD.t77 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X922 TG_GATE_SWITCH_magic_7.B a_n1894_307.t29 A2.t0 VDD.t188 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X923 TG_magic_4.B a_2061_n4852.t29 TG_magic_7.B.t38 VDD.t14 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
R0 a_3874_308.t15 a_3874_308.n30 40.7345
R1 a_3874_308.n7 a_3874_308.n6 28.094
R2 a_3874_308.n16 a_3874_308.n15 28.094
R3 a_3874_308.n32 a_3874_308.n31 28.094
R4 a_3874_308.n4 a_3874_308.t6 21.9005
R5 a_3874_308.n2 a_3874_308.t20 21.9005
R6 a_3874_308.n1 a_3874_308.t24 21.9005
R7 a_3874_308.n10 a_3874_308.t18 21.9005
R8 a_3874_308.n10 a_3874_308.t11 21.9005
R9 a_3874_308.n22 a_3874_308.t26 21.9005
R10 a_3874_308.n23 a_3874_308.t21 21.9005
R11 a_3874_308.n11 a_3874_308.t9 21.9005
R12 a_3874_308.n11 a_3874_308.t16 21.9005
R13 a_3874_308.n3 a_3874_308.t23 21.9005
R14 a_3874_308.n12 a_3874_308.t17 21.9005
R15 a_3874_308.n12 a_3874_308.t10 21.9005
R16 a_3874_308.n24 a_3874_308.t25 21.9005
R17 a_3874_308.n25 a_3874_308.t7 21.9005
R18 a_3874_308.n13 a_3874_308.t19 21.9005
R19 a_3874_308.n13 a_3874_308.t22 21.9005
R20 a_3874_308.n6 a_3874_308.t14 21.9005
R21 a_3874_308.n15 a_3874_308.t28 21.9005
R22 a_3874_308.n15 a_3874_308.t8 21.9005
R23 a_3874_308.n5 a_3874_308.t12 21.9005
R24 a_3874_308.n14 a_3874_308.t29 21.9005
R25 a_3874_308.n14 a_3874_308.t27 21.9005
R26 a_3874_308.n26 a_3874_308.t13 21.9005
R27 a_3874_308.n31 a_3874_308.t15 21.9005
R28 a_3874_308.n31 a_3874_308.n26 15.8172
R29 a_3874_308.n14 a_3874_308.n13 15.8172
R30 a_3874_308.n26 a_3874_308.n25 15.8172
R31 a_3874_308.n25 a_3874_308.n24 15.8172
R32 a_3874_308.n13 a_3874_308.n12 15.8172
R33 a_3874_308.n12 a_3874_308.n11 15.8172
R34 a_3874_308.n24 a_3874_308.n23 15.8172
R35 a_3874_308.n23 a_3874_308.n22 15.8172
R36 a_3874_308.n11 a_3874_308.n10 15.8172
R37 a_3874_308.n2 a_3874_308.n1 15.8172
R38 a_3874_308.n4 a_3874_308.n3 15.8172
R39 a_3874_308.n3 a_3874_308.n2 15.8172
R40 a_3874_308.n15 a_3874_308.n14 15.8172
R41 a_3874_308.n6 a_3874_308.n5 15.8172
R42 a_3874_308.n5 a_3874_308.n4 15.8172
R43 a_3874_308.n28 a_3874_308.n27 15.1845
R44 a_3874_308.n30 a_3874_308.n29 15.1845
R45 a_3874_308.n29 a_3874_308.n28 15.1845
R46 a_3874_308.n20 a_3874_308.n19 5.44589
R47 a_3874_308.n20 a_3874_308.n18 4.7885
R48 a_3874_308.n7 a_3874_308.n0 4.70615
R49 a_3874_308.n21 a_3874_308.n17 4.4205
R50 a_3874_308.n9 a_3874_308.n8 4.4205
R51 a_3874_308.n34 a_3874_308.n33 4.4205
R52 a_3874_308.n21 a_3874_308.n20 1.1392
R53 a_3874_308.n16 a_3874_308.n9 0.286152
R54 a_3874_308.n33 a_3874_308.n32 0.286152
R55 a_3874_308.n32 a_3874_308.n21 0.282239
R56 a_3874_308.n9 a_3874_308.n7 0.282239
R57 a_3874_308.n33 a_3874_308.n16 0.282239
R58 TG_GATE_SWITCH_magic_7.B.n106 TG_GATE_SWITCH_magic_7.B.n105 6.81159
R59 TG_GATE_SWITCH_magic_7.B.n64 TG_GATE_SWITCH_magic_7.B.n62 5.44589
R60 TG_GATE_SWITCH_magic_7.B.n84 TG_GATE_SWITCH_magic_7.B.n83 5.07789
R61 TG_GATE_SWITCH_magic_7.B.n68 TG_GATE_SWITCH_magic_7.B.t17 4.7885
R62 TG_GATE_SWITCH_magic_7.B.n67 TG_GATE_SWITCH_magic_7.B.t20 4.7885
R63 TG_GATE_SWITCH_magic_7.B.n64 TG_GATE_SWITCH_magic_7.B.n63 4.7885
R64 TG_GATE_SWITCH_magic_7.B.n103 TG_GATE_SWITCH_magic_7.B.t56 4.4205
R65 TG_GATE_SWITCH_magic_7.B.n102 TG_GATE_SWITCH_magic_7.B.t50 4.4205
R66 TG_GATE_SWITCH_magic_7.B.n101 TG_GATE_SWITCH_magic_7.B.t59 4.4205
R67 TG_GATE_SWITCH_magic_7.B.n100 TG_GATE_SWITCH_magic_7.B.t57 4.4205
R68 TG_GATE_SWITCH_magic_7.B.n86 TG_GATE_SWITCH_magic_7.B.n80 4.4205
R69 TG_GATE_SWITCH_magic_7.B.n85 TG_GATE_SWITCH_magic_7.B.n81 4.4205
R70 TG_GATE_SWITCH_magic_7.B.n84 TG_GATE_SWITCH_magic_7.B.n82 4.4205
R71 TG_GATE_SWITCH_magic_7.B.n61 TG_GATE_SWITCH_magic_7.B.n58 3.80789
R72 TG_GATE_SWITCH_magic_7.B.n56 TG_GATE_SWITCH_magic_7.B.n53 3.80789
R73 TG_GATE_SWITCH_magic_7.B.n48 TG_GATE_SWITCH_magic_7.B.n47 3.80789
R74 TG_GATE_SWITCH_magic_7.B.n43 TG_GATE_SWITCH_magic_7.B.n42 3.80789
R75 TG_GATE_SWITCH_magic_7.B.n38 TG_GATE_SWITCH_magic_7.B.n37 3.80789
R76 TG_GATE_SWITCH_magic_7.B.n105 TG_GATE_SWITCH_magic_7.B.n104 3.31029
R77 TG_GATE_SWITCH_magic_7.B.n4 TG_GATE_SWITCH_magic_7.B.n1 3.25789
R78 TG_GATE_SWITCH_magic_7.B.n15 TG_GATE_SWITCH_magic_7.B.n12 3.25789
R79 TG_GATE_SWITCH_magic_7.B.n27 TG_GATE_SWITCH_magic_7.B.n24 3.25789
R80 TG_GATE_SWITCH_magic_7.B.n77 TG_GATE_SWITCH_magic_7.B.n76 3.25789
R81 TG_GATE_SWITCH_magic_7.B.n94 TG_GATE_SWITCH_magic_7.B.n93 3.25789
R82 TG_GATE_SWITCH_magic_7.B.n61 TG_GATE_SWITCH_magic_7.B.n60 3.1505
R83 TG_GATE_SWITCH_magic_7.B.n56 TG_GATE_SWITCH_magic_7.B.n55 3.1505
R84 TG_GATE_SWITCH_magic_7.B.n48 TG_GATE_SWITCH_magic_7.B.n45 3.1505
R85 TG_GATE_SWITCH_magic_7.B.n43 TG_GATE_SWITCH_magic_7.B.n40 3.1505
R86 TG_GATE_SWITCH_magic_7.B.n38 TG_GATE_SWITCH_magic_7.B.n35 3.1505
R87 TG_GATE_SWITCH_magic_7.B.n4 TG_GATE_SWITCH_magic_7.B.n3 2.6005
R88 TG_GATE_SWITCH_magic_7.B.n7 TG_GATE_SWITCH_magic_7.B.n6 2.6005
R89 TG_GATE_SWITCH_magic_7.B.n10 TG_GATE_SWITCH_magic_7.B.n9 2.6005
R90 TG_GATE_SWITCH_magic_7.B.n18 TG_GATE_SWITCH_magic_7.B.n17 2.6005
R91 TG_GATE_SWITCH_magic_7.B.n15 TG_GATE_SWITCH_magic_7.B.n14 2.6005
R92 TG_GATE_SWITCH_magic_7.B.n21 TG_GATE_SWITCH_magic_7.B.n20 2.6005
R93 TG_GATE_SWITCH_magic_7.B.n27 TG_GATE_SWITCH_magic_7.B.n26 2.6005
R94 TG_GATE_SWITCH_magic_7.B.n30 TG_GATE_SWITCH_magic_7.B.n29 2.6005
R95 TG_GATE_SWITCH_magic_7.B.n33 TG_GATE_SWITCH_magic_7.B.n32 2.6005
R96 TG_GATE_SWITCH_magic_7.B.n77 TG_GATE_SWITCH_magic_7.B.n74 2.6005
R97 TG_GATE_SWITCH_magic_7.B.n78 TG_GATE_SWITCH_magic_7.B.n72 2.6005
R98 TG_GATE_SWITCH_magic_7.B.n79 TG_GATE_SWITCH_magic_7.B.n70 2.6005
R99 TG_GATE_SWITCH_magic_7.B.n94 TG_GATE_SWITCH_magic_7.B.n91 2.6005
R100 TG_GATE_SWITCH_magic_7.B.n95 TG_GATE_SWITCH_magic_7.B.n89 2.6005
R101 TG_GATE_SWITCH_magic_7.B.n98 TG_GATE_SWITCH_magic_7.B.n97 2.6005
R102 TG_GATE_SWITCH_magic_7.B.n89 TG_GATE_SWITCH_magic_7.B.t51 1.8205
R103 TG_GATE_SWITCH_magic_7.B.n89 TG_GATE_SWITCH_magic_7.B.n88 1.8205
R104 TG_GATE_SWITCH_magic_7.B.n91 TG_GATE_SWITCH_magic_7.B.t54 1.8205
R105 TG_GATE_SWITCH_magic_7.B.n91 TG_GATE_SWITCH_magic_7.B.n90 1.8205
R106 TG_GATE_SWITCH_magic_7.B.n93 TG_GATE_SWITCH_magic_7.B.t60 1.8205
R107 TG_GATE_SWITCH_magic_7.B.n93 TG_GATE_SWITCH_magic_7.B.n92 1.8205
R108 TG_GATE_SWITCH_magic_7.B.n9 TG_GATE_SWITCH_magic_7.B.t44 1.8205
R109 TG_GATE_SWITCH_magic_7.B.n9 TG_GATE_SWITCH_magic_7.B.n8 1.8205
R110 TG_GATE_SWITCH_magic_7.B.n6 TG_GATE_SWITCH_magic_7.B.t34 1.8205
R111 TG_GATE_SWITCH_magic_7.B.n6 TG_GATE_SWITCH_magic_7.B.n5 1.8205
R112 TG_GATE_SWITCH_magic_7.B.n3 TG_GATE_SWITCH_magic_7.B.t38 1.8205
R113 TG_GATE_SWITCH_magic_7.B.n3 TG_GATE_SWITCH_magic_7.B.n2 1.8205
R114 TG_GATE_SWITCH_magic_7.B.n1 TG_GATE_SWITCH_magic_7.B.t42 1.8205
R115 TG_GATE_SWITCH_magic_7.B.n1 TG_GATE_SWITCH_magic_7.B.n0 1.8205
R116 TG_GATE_SWITCH_magic_7.B.n20 TG_GATE_SWITCH_magic_7.B.t37 1.8205
R117 TG_GATE_SWITCH_magic_7.B.n20 TG_GATE_SWITCH_magic_7.B.n19 1.8205
R118 TG_GATE_SWITCH_magic_7.B.n12 TG_GATE_SWITCH_magic_7.B.t35 1.8205
R119 TG_GATE_SWITCH_magic_7.B.n12 TG_GATE_SWITCH_magic_7.B.n11 1.8205
R120 TG_GATE_SWITCH_magic_7.B.n14 TG_GATE_SWITCH_magic_7.B.t29 1.8205
R121 TG_GATE_SWITCH_magic_7.B.n14 TG_GATE_SWITCH_magic_7.B.n13 1.8205
R122 TG_GATE_SWITCH_magic_7.B.n17 TG_GATE_SWITCH_magic_7.B.t46 1.8205
R123 TG_GATE_SWITCH_magic_7.B.n17 TG_GATE_SWITCH_magic_7.B.n16 1.8205
R124 TG_GATE_SWITCH_magic_7.B.n32 TG_GATE_SWITCH_magic_7.B.t28 1.8205
R125 TG_GATE_SWITCH_magic_7.B.n32 TG_GATE_SWITCH_magic_7.B.n31 1.8205
R126 TG_GATE_SWITCH_magic_7.B.n29 TG_GATE_SWITCH_magic_7.B.t40 1.8205
R127 TG_GATE_SWITCH_magic_7.B.n29 TG_GATE_SWITCH_magic_7.B.n28 1.8205
R128 TG_GATE_SWITCH_magic_7.B.n26 TG_GATE_SWITCH_magic_7.B.t14 1.8205
R129 TG_GATE_SWITCH_magic_7.B.n26 TG_GATE_SWITCH_magic_7.B.n25 1.8205
R130 TG_GATE_SWITCH_magic_7.B.n24 TG_GATE_SWITCH_magic_7.B.t27 1.8205
R131 TG_GATE_SWITCH_magic_7.B.n24 TG_GATE_SWITCH_magic_7.B.n23 1.8205
R132 TG_GATE_SWITCH_magic_7.B.n70 TG_GATE_SWITCH_magic_7.B.t53 1.8205
R133 TG_GATE_SWITCH_magic_7.B.n70 TG_GATE_SWITCH_magic_7.B.n69 1.8205
R134 TG_GATE_SWITCH_magic_7.B.n72 TG_GATE_SWITCH_magic_7.B.t55 1.8205
R135 TG_GATE_SWITCH_magic_7.B.n72 TG_GATE_SWITCH_magic_7.B.n71 1.8205
R136 TG_GATE_SWITCH_magic_7.B.n74 TG_GATE_SWITCH_magic_7.B.t58 1.8205
R137 TG_GATE_SWITCH_magic_7.B.n74 TG_GATE_SWITCH_magic_7.B.n73 1.8205
R138 TG_GATE_SWITCH_magic_7.B.n76 TG_GATE_SWITCH_magic_7.B.t52 1.8205
R139 TG_GATE_SWITCH_magic_7.B.n76 TG_GATE_SWITCH_magic_7.B.n75 1.8205
R140 TG_GATE_SWITCH_magic_7.B.n97 TG_GATE_SWITCH_magic_7.B.t61 1.8205
R141 TG_GATE_SWITCH_magic_7.B.n97 TG_GATE_SWITCH_magic_7.B.n96 1.8205
R142 TG_GATE_SWITCH_magic_7.B.n60 TG_GATE_SWITCH_magic_7.B.t18 1.6385
R143 TG_GATE_SWITCH_magic_7.B.n60 TG_GATE_SWITCH_magic_7.B.n59 1.6385
R144 TG_GATE_SWITCH_magic_7.B.n58 TG_GATE_SWITCH_magic_7.B.t15 1.6385
R145 TG_GATE_SWITCH_magic_7.B.n58 TG_GATE_SWITCH_magic_7.B.n57 1.6385
R146 TG_GATE_SWITCH_magic_7.B.n55 TG_GATE_SWITCH_magic_7.B.t16 1.6385
R147 TG_GATE_SWITCH_magic_7.B.n55 TG_GATE_SWITCH_magic_7.B.n54 1.6385
R148 TG_GATE_SWITCH_magic_7.B.n53 TG_GATE_SWITCH_magic_7.B.t19 1.6385
R149 TG_GATE_SWITCH_magic_7.B.n53 TG_GATE_SWITCH_magic_7.B.n52 1.6385
R150 TG_GATE_SWITCH_magic_7.B.n45 TG_GATE_SWITCH_magic_7.B.t2 1.6385
R151 TG_GATE_SWITCH_magic_7.B.n45 TG_GATE_SWITCH_magic_7.B.n44 1.6385
R152 TG_GATE_SWITCH_magic_7.B.n47 TG_GATE_SWITCH_magic_7.B.t5 1.6385
R153 TG_GATE_SWITCH_magic_7.B.n47 TG_GATE_SWITCH_magic_7.B.n46 1.6385
R154 TG_GATE_SWITCH_magic_7.B.n40 TG_GATE_SWITCH_magic_7.B.t6 1.6385
R155 TG_GATE_SWITCH_magic_7.B.n40 TG_GATE_SWITCH_magic_7.B.n39 1.6385
R156 TG_GATE_SWITCH_magic_7.B.n42 TG_GATE_SWITCH_magic_7.B.t3 1.6385
R157 TG_GATE_SWITCH_magic_7.B.n42 TG_GATE_SWITCH_magic_7.B.n41 1.6385
R158 TG_GATE_SWITCH_magic_7.B.n35 TG_GATE_SWITCH_magic_7.B.t4 1.6385
R159 TG_GATE_SWITCH_magic_7.B.n35 TG_GATE_SWITCH_magic_7.B.n34 1.6385
R160 TG_GATE_SWITCH_magic_7.B.n37 TG_GATE_SWITCH_magic_7.B.t7 1.6385
R161 TG_GATE_SWITCH_magic_7.B.n37 TG_GATE_SWITCH_magic_7.B.n36 1.6385
R162 TG_GATE_SWITCH_magic_7.B.n105 TG_GATE_SWITCH_magic_7.B 1.16794
R163 TG_GATE_SWITCH_magic_7.B.n65 TG_GATE_SWITCH_magic_7.B.n64 0.884196
R164 TG_GATE_SWITCH_magic_7.B.n67 TG_GATE_SWITCH_magic_7.B.n66 0.884196
R165 TG_GATE_SWITCH_magic_7.B.n100 TG_GATE_SWITCH_magic_7.B.n99 0.882239
R166 TG_GATE_SWITCH_magic_7.B.n87 TG_GATE_SWITCH_magic_7.B.n86 0.882239
R167 TG_GATE_SWITCH_magic_7.B.n104 TG_GATE_SWITCH_magic_7.B.n68 0.8105
R168 TG_GATE_SWITCH_magic_7.B.n68 TG_GATE_SWITCH_magic_7.B.n67 0.657891
R169 TG_GATE_SWITCH_magic_7.B.n7 TG_GATE_SWITCH_magic_7.B.n4 0.657891
R170 TG_GATE_SWITCH_magic_7.B.n10 TG_GATE_SWITCH_magic_7.B.n7 0.657891
R171 TG_GATE_SWITCH_magic_7.B.n18 TG_GATE_SWITCH_magic_7.B.n15 0.657891
R172 TG_GATE_SWITCH_magic_7.B.n30 TG_GATE_SWITCH_magic_7.B.n27 0.657891
R173 TG_GATE_SWITCH_magic_7.B.n33 TG_GATE_SWITCH_magic_7.B.n30 0.657891
R174 TG_GATE_SWITCH_magic_7.B.n101 TG_GATE_SWITCH_magic_7.B.n100 0.657891
R175 TG_GATE_SWITCH_magic_7.B.n102 TG_GATE_SWITCH_magic_7.B.n101 0.657891
R176 TG_GATE_SWITCH_magic_7.B.n103 TG_GATE_SWITCH_magic_7.B.n102 0.657891
R177 TG_GATE_SWITCH_magic_7.B.n79 TG_GATE_SWITCH_magic_7.B.n78 0.657891
R178 TG_GATE_SWITCH_magic_7.B.n78 TG_GATE_SWITCH_magic_7.B.n77 0.657891
R179 TG_GATE_SWITCH_magic_7.B.n86 TG_GATE_SWITCH_magic_7.B.n85 0.657891
R180 TG_GATE_SWITCH_magic_7.B.n85 TG_GATE_SWITCH_magic_7.B.n84 0.657891
R181 TG_GATE_SWITCH_magic_7.B.n98 TG_GATE_SWITCH_magic_7.B.n95 0.657891
R182 TG_GATE_SWITCH_magic_7.B.n95 TG_GATE_SWITCH_magic_7.B.n94 0.657891
R183 TG_GATE_SWITCH_magic_7.B.n21 TG_GATE_SWITCH_magic_7.B.n18 0.655976
R184 TG_GATE_SWITCH_magic_7.B.n22 TG_GATE_SWITCH_magic_7.B.n21 0.645657
R185 TG_GATE_SWITCH_magic_7.B.n66 TG_GATE_SWITCH_magic_7.B.n65 0.6005
R186 TG_GATE_SWITCH_magic_7.B.n99 TG_GATE_SWITCH_magic_7.B.n87 0.6005
R187 TG_GATE_SWITCH_magic_7.B.n49 TG_GATE_SWITCH_magic_7.B.n48 0.548416
R188 TG_GATE_SWITCH_magic_7.B.n51 TG_GATE_SWITCH_magic_7.B.n33 0.317366
R189 TG_GATE_SWITCH_magic_7.B.n50 TG_GATE_SWITCH_magic_7.B.n38 0.304838
R190 TG_GATE_SWITCH_magic_7.B.n65 TG_GATE_SWITCH_magic_7.B.n61 0.284196
R191 TG_GATE_SWITCH_magic_7.B.n66 TG_GATE_SWITCH_magic_7.B.n56 0.284196
R192 TG_GATE_SWITCH_magic_7.B.n49 TG_GATE_SWITCH_magic_7.B.n43 0.284196
R193 TG_GATE_SWITCH_magic_7.B.n51 TG_GATE_SWITCH_magic_7.B.n22 0.283032
R194 TG_GATE_SWITCH_magic_7.B.n87 TG_GATE_SWITCH_magic_7.B.n79 0.282239
R195 TG_GATE_SWITCH_magic_7.B.n99 TG_GATE_SWITCH_magic_7.B.n98 0.282239
R196 TG_GATE_SWITCH_magic_7.B.n22 TG_GATE_SWITCH_magic_7.B.n10 0.279866
R197 TG_GATE_SWITCH_magic_7.B.n106 TG_GATE_SWITCH_magic_7.B.n51 0.251024
R198 TG_GATE_SWITCH_magic_7.B.n50 TG_GATE_SWITCH_magic_7.B.n49 0.244078
R199 TG_GATE_SWITCH_magic_7.B.n104 TG_GATE_SWITCH_magic_7.B.n103 0.237239
R200 TG_GATE_SWITCH_magic_7.B.n51 TG_GATE_SWITCH_magic_7.B.n50 0.1355
R201 TG_GATE_SWITCH_magic_7.B TG_GATE_SWITCH_magic_7.B.n106 0.0366932
R202 TG_magic_5.A.n52 TG_magic_5.A.t33 5.44589
R203 TG_magic_5.A.n104 TG_magic_5.A 5.33254
R204 TG_magic_5.A.n95 TG_magic_5.A.t23 5.07789
R205 TG_magic_5.A.n106 TG_magic_5.A.n67 4.7885
R206 TG_magic_5.A.n105 TG_magic_5.A.n68 4.7885
R207 TG_magic_5.A.n52 TG_magic_5.A.t29 4.7885
R208 TG_magic_5.A.n103 TG_magic_5.A.n69 4.4205
R209 TG_magic_5.A.n102 TG_magic_5.A.n70 4.4205
R210 TG_magic_5.A.n101 TG_magic_5.A.n71 4.4205
R211 TG_magic_5.A.n100 TG_magic_5.A.n72 4.4205
R212 TG_magic_5.A.n97 TG_magic_5.A.t73 4.4205
R213 TG_magic_5.A.n96 TG_magic_5.A.t49 4.4205
R214 TG_magic_5.A.n95 TG_magic_5.A.t70 4.4205
R215 TG_magic_5.A.n62 TG_magic_5.A.n61 3.80789
R216 TG_magic_5.A.n57 TG_magic_5.A.n56 3.80789
R217 TG_magic_5.A.n49 TG_magic_5.A.n48 3.80789
R218 TG_magic_5.A.n38 TG_magic_5.A.n37 3.80789
R219 TG_magic_5.A.n43 TG_magic_5.A.n42 3.80789
R220 TG_magic_5.A.n135 TG_magic_5.A.n134 3.80789
R221 TG_magic_5.A.n130 TG_magic_5.A.n129 3.80789
R222 TG_magic_5.A.n125 TG_magic_5.A.n124 3.80789
R223 TG_magic_5.A.n77 TG_magic_5.A.n74 3.25789
R224 TG_magic_5.A.n88 TG_magic_5.A.n85 3.25789
R225 TG_magic_5.A.n15 TG_magic_5.A.n12 3.25789
R226 TG_magic_5.A.n4 TG_magic_5.A.n1 3.25789
R227 TG_magic_5.A.n27 TG_magic_5.A.n24 3.25789
R228 TG_magic_5.A.n114 TG_magic_5.A.n111 3.25789
R229 TG_magic_5.A.n142 TG_magic_5.A.n139 3.25789
R230 TG_magic_5.A.n153 TG_magic_5.A.n150 3.25789
R231 TG_magic_5.A.n62 TG_magic_5.A.n59 3.1505
R232 TG_magic_5.A.n57 TG_magic_5.A.n54 3.1505
R233 TG_magic_5.A.n49 TG_magic_5.A.n46 3.1505
R234 TG_magic_5.A.n38 TG_magic_5.A.n35 3.1505
R235 TG_magic_5.A.n43 TG_magic_5.A.n40 3.1505
R236 TG_magic_5.A.n135 TG_magic_5.A.n132 3.1505
R237 TG_magic_5.A.n130 TG_magic_5.A.n127 3.1505
R238 TG_magic_5.A.n125 TG_magic_5.A.n122 3.1505
R239 TG_magic_5.A.n109 TG_magic_5.A.n108 2.76897
R240 TG_magic_5.A.n77 TG_magic_5.A.n76 2.6005
R241 TG_magic_5.A.n80 TG_magic_5.A.n79 2.6005
R242 TG_magic_5.A.n83 TG_magic_5.A.n82 2.6005
R243 TG_magic_5.A.n88 TG_magic_5.A.n87 2.6005
R244 TG_magic_5.A.n91 TG_magic_5.A.n90 2.6005
R245 TG_magic_5.A.n94 TG_magic_5.A.n93 2.6005
R246 TG_magic_5.A.n15 TG_magic_5.A.n14 2.6005
R247 TG_magic_5.A.n18 TG_magic_5.A.n17 2.6005
R248 TG_magic_5.A.n21 TG_magic_5.A.n20 2.6005
R249 TG_magic_5.A.n4 TG_magic_5.A.n3 2.6005
R250 TG_magic_5.A.n7 TG_magic_5.A.n6 2.6005
R251 TG_magic_5.A.n10 TG_magic_5.A.n9 2.6005
R252 TG_magic_5.A.n27 TG_magic_5.A.n26 2.6005
R253 TG_magic_5.A.n30 TG_magic_5.A.n29 2.6005
R254 TG_magic_5.A.n33 TG_magic_5.A.n32 2.6005
R255 TG_magic_5.A.n114 TG_magic_5.A.n113 2.6005
R256 TG_magic_5.A.n117 TG_magic_5.A.n116 2.6005
R257 TG_magic_5.A.n120 TG_magic_5.A.n119 2.6005
R258 TG_magic_5.A.n145 TG_magic_5.A.n144 2.6005
R259 TG_magic_5.A.n142 TG_magic_5.A.n141 2.6005
R260 TG_magic_5.A.n148 TG_magic_5.A.n147 2.6005
R261 TG_magic_5.A.n153 TG_magic_5.A.n152 2.6005
R262 TG_magic_5.A.n156 TG_magic_5.A.n155 2.6005
R263 TG_magic_5.A.n159 TG_magic_5.A.n158 2.6005
R264 TG_magic_5.A.n108 TG_magic_5.A.n107 2.2505
R265 TG_magic_5.A.n155 TG_magic_5.A.t103 1.8205
R266 TG_magic_5.A.n155 TG_magic_5.A.n154 1.8205
R267 TG_magic_5.A.n152 TG_magic_5.A.t96 1.8205
R268 TG_magic_5.A.n152 TG_magic_5.A.n151 1.8205
R269 TG_magic_5.A.n150 TG_magic_5.A.t90 1.8205
R270 TG_magic_5.A.n150 TG_magic_5.A.n149 1.8205
R271 TG_magic_5.A.n82 TG_magic_5.A.t61 1.8205
R272 TG_magic_5.A.n82 TG_magic_5.A.n81 1.8205
R273 TG_magic_5.A.n79 TG_magic_5.A.t60 1.8205
R274 TG_magic_5.A.n79 TG_magic_5.A.n78 1.8205
R275 TG_magic_5.A.n76 TG_magic_5.A.t68 1.8205
R276 TG_magic_5.A.n76 TG_magic_5.A.n75 1.8205
R277 TG_magic_5.A.n74 TG_magic_5.A.t50 1.8205
R278 TG_magic_5.A.n74 TG_magic_5.A.n73 1.8205
R279 TG_magic_5.A.n93 TG_magic_5.A.t78 1.8205
R280 TG_magic_5.A.n93 TG_magic_5.A.n92 1.8205
R281 TG_magic_5.A.n90 TG_magic_5.A.t67 1.8205
R282 TG_magic_5.A.n90 TG_magic_5.A.n89 1.8205
R283 TG_magic_5.A.n87 TG_magic_5.A.t52 1.8205
R284 TG_magic_5.A.n87 TG_magic_5.A.n86 1.8205
R285 TG_magic_5.A.n85 TG_magic_5.A.t62 1.8205
R286 TG_magic_5.A.n85 TG_magic_5.A.n84 1.8205
R287 TG_magic_5.A.n20 TG_magic_5.A.t41 1.8205
R288 TG_magic_5.A.n20 TG_magic_5.A.n19 1.8205
R289 TG_magic_5.A.n17 TG_magic_5.A.t53 1.8205
R290 TG_magic_5.A.n17 TG_magic_5.A.n16 1.8205
R291 TG_magic_5.A.n14 TG_magic_5.A.t57 1.8205
R292 TG_magic_5.A.n14 TG_magic_5.A.n13 1.8205
R293 TG_magic_5.A.n12 TG_magic_5.A.t39 1.8205
R294 TG_magic_5.A.n12 TG_magic_5.A.n11 1.8205
R295 TG_magic_5.A.n9 TG_magic_5.A.t81 1.8205
R296 TG_magic_5.A.n9 TG_magic_5.A.n8 1.8205
R297 TG_magic_5.A.n6 TG_magic_5.A.t37 1.8205
R298 TG_magic_5.A.n6 TG_magic_5.A.n5 1.8205
R299 TG_magic_5.A.n3 TG_magic_5.A.t42 1.8205
R300 TG_magic_5.A.n3 TG_magic_5.A.n2 1.8205
R301 TG_magic_5.A.n1 TG_magic_5.A.t79 1.8205
R302 TG_magic_5.A.n1 TG_magic_5.A.n0 1.8205
R303 TG_magic_5.A.n32 TG_magic_5.A.t80 1.8205
R304 TG_magic_5.A.n32 TG_magic_5.A.n31 1.8205
R305 TG_magic_5.A.n29 TG_magic_5.A.t36 1.8205
R306 TG_magic_5.A.n29 TG_magic_5.A.n28 1.8205
R307 TG_magic_5.A.n26 TG_magic_5.A.t40 1.8205
R308 TG_magic_5.A.n26 TG_magic_5.A.n25 1.8205
R309 TG_magic_5.A.n24 TG_magic_5.A.t48 1.8205
R310 TG_magic_5.A.n24 TG_magic_5.A.n23 1.8205
R311 TG_magic_5.A.n119 TG_magic_5.A.t87 1.8205
R312 TG_magic_5.A.n119 TG_magic_5.A.n118 1.8205
R313 TG_magic_5.A.n116 TG_magic_5.A.t102 1.8205
R314 TG_magic_5.A.n116 TG_magic_5.A.n115 1.8205
R315 TG_magic_5.A.n113 TG_magic_5.A.t95 1.8205
R316 TG_magic_5.A.n113 TG_magic_5.A.n112 1.8205
R317 TG_magic_5.A.n111 TG_magic_5.A.t89 1.8205
R318 TG_magic_5.A.n111 TG_magic_5.A.n110 1.8205
R319 TG_magic_5.A.n147 TG_magic_5.A.t100 1.8205
R320 TG_magic_5.A.n147 TG_magic_5.A.n146 1.8205
R321 TG_magic_5.A.n139 TG_magic_5.A.t101 1.8205
R322 TG_magic_5.A.n139 TG_magic_5.A.n138 1.8205
R323 TG_magic_5.A.n141 TG_magic_5.A.t84 1.8205
R324 TG_magic_5.A.n141 TG_magic_5.A.n140 1.8205
R325 TG_magic_5.A.n144 TG_magic_5.A.t86 1.8205
R326 TG_magic_5.A.n144 TG_magic_5.A.n143 1.8205
R327 TG_magic_5.A.n158 TG_magic_5.A.t88 1.8205
R328 TG_magic_5.A.n158 TG_magic_5.A.n157 1.8205
R329 TG_magic_5.A.n59 TG_magic_5.A.t25 1.6385
R330 TG_magic_5.A.n59 TG_magic_5.A.n58 1.6385
R331 TG_magic_5.A.n61 TG_magic_5.A.t26 1.6385
R332 TG_magic_5.A.n61 TG_magic_5.A.n60 1.6385
R333 TG_magic_5.A.n54 TG_magic_5.A.t30 1.6385
R334 TG_magic_5.A.n54 TG_magic_5.A.n53 1.6385
R335 TG_magic_5.A.n56 TG_magic_5.A.t34 1.6385
R336 TG_magic_5.A.n56 TG_magic_5.A.n55 1.6385
R337 TG_magic_5.A.n46 TG_magic_5.A.t17 1.6385
R338 TG_magic_5.A.n46 TG_magic_5.A.n45 1.6385
R339 TG_magic_5.A.n48 TG_magic_5.A.t58 1.6385
R340 TG_magic_5.A.n48 TG_magic_5.A.n47 1.6385
R341 TG_magic_5.A.n35 TG_magic_5.A.t3 1.6385
R342 TG_magic_5.A.n35 TG_magic_5.A.n34 1.6385
R343 TG_magic_5.A.n37 TG_magic_5.A.t20 1.6385
R344 TG_magic_5.A.n37 TG_magic_5.A.n36 1.6385
R345 TG_magic_5.A.n40 TG_magic_5.A.t16 1.6385
R346 TG_magic_5.A.n40 TG_magic_5.A.n39 1.6385
R347 TG_magic_5.A.n42 TG_magic_5.A.t74 1.6385
R348 TG_magic_5.A.n42 TG_magic_5.A.n41 1.6385
R349 TG_magic_5.A.n132 TG_magic_5.A.t6 1.6385
R350 TG_magic_5.A.n132 TG_magic_5.A.n131 1.6385
R351 TG_magic_5.A.n134 TG_magic_5.A.t12 1.6385
R352 TG_magic_5.A.n134 TG_magic_5.A.n133 1.6385
R353 TG_magic_5.A.n127 TG_magic_5.A.t8 1.6385
R354 TG_magic_5.A.n127 TG_magic_5.A.n126 1.6385
R355 TG_magic_5.A.n129 TG_magic_5.A.t14 1.6385
R356 TG_magic_5.A.n129 TG_magic_5.A.n128 1.6385
R357 TG_magic_5.A.n122 TG_magic_5.A.t4 1.6385
R358 TG_magic_5.A.n122 TG_magic_5.A.n121 1.6385
R359 TG_magic_5.A.n124 TG_magic_5.A.t10 1.6385
R360 TG_magic_5.A.n124 TG_magic_5.A.n123 1.6385
R361 TG_magic_5.A.n66 TG_magic_5.A.n65 1.44849
R362 TG_magic_5.A.n109 TG_magic_5.A 1.13908
R363 TG_magic_5.A.n98 TG_magic_5.A.n97 0.882239
R364 TG_magic_5.A.n100 TG_magic_5.A.n99 0.882239
R365 TG_magic_5.A.n105 TG_magic_5.A.n104 0.8105
R366 TG_magic_5.A TG_magic_5.A.n109 0.724738
R367 TG_magic_5.A.n80 TG_magic_5.A.n77 0.657891
R368 TG_magic_5.A.n83 TG_magic_5.A.n80 0.657891
R369 TG_magic_5.A.n91 TG_magic_5.A.n88 0.657891
R370 TG_magic_5.A.n94 TG_magic_5.A.n91 0.657891
R371 TG_magic_5.A.n96 TG_magic_5.A.n95 0.657891
R372 TG_magic_5.A.n97 TG_magic_5.A.n96 0.657891
R373 TG_magic_5.A.n103 TG_magic_5.A.n102 0.657891
R374 TG_magic_5.A.n102 TG_magic_5.A.n101 0.657891
R375 TG_magic_5.A.n101 TG_magic_5.A.n100 0.657891
R376 TG_magic_5.A.n106 TG_magic_5.A.n105 0.657891
R377 TG_magic_5.A.n18 TG_magic_5.A.n15 0.657891
R378 TG_magic_5.A.n7 TG_magic_5.A.n4 0.657891
R379 TG_magic_5.A.n10 TG_magic_5.A.n7 0.657891
R380 TG_magic_5.A.n30 TG_magic_5.A.n27 0.657891
R381 TG_magic_5.A.n33 TG_magic_5.A.n30 0.657891
R382 TG_magic_5.A.n117 TG_magic_5.A.n114 0.657891
R383 TG_magic_5.A.n120 TG_magic_5.A.n117 0.657891
R384 TG_magic_5.A.n145 TG_magic_5.A.n142 0.657891
R385 TG_magic_5.A.n156 TG_magic_5.A.n153 0.657891
R386 TG_magic_5.A.n159 TG_magic_5.A.n156 0.657891
R387 TG_magic_5.A.n21 TG_magic_5.A.n18 0.655976
R388 TG_magic_5.A.n148 TG_magic_5.A.n145 0.655976
R389 TG_magic_5.A.n22 TG_magic_5.A.n21 0.646796
R390 TG_magic_5.A.n160 TG_magic_5.A.n148 0.645657
R391 TG_magic_5.A.n99 TG_magic_5.A.n98 0.6005
R392 TG_magic_5.A.n44 TG_magic_5.A.n43 0.548416
R393 TG_magic_5.A.n136 TG_magic_5.A.n135 0.548416
R394 TG_magic_5.A.n64 TG_magic_5.A.n63 0.518782
R395 TG_magic_5.A.n65 TG_magic_5.A.n52 0.496104
R396 TG_magic_5.A.n108 TG_magic_5.A.n66 0.363884
R397 TG_magic_5.A.n51 TG_magic_5.A.n33 0.317366
R398 TG_magic_5.A.n161 TG_magic_5.A.n120 0.317366
R399 TG_magic_5.A.n50 TG_magic_5.A.n49 0.304838
R400 TG_magic_5.A.n137 TG_magic_5.A.n125 0.304838
R401 TG_magic_5.A TG_magic_5.A.n51 0.2873
R402 TG_magic_5.A TG_magic_5.A.n161 0.2873
R403 TG_magic_5.A.n44 TG_magic_5.A.n38 0.284196
R404 TG_magic_5.A.n136 TG_magic_5.A.n130 0.284196
R405 TG_magic_5.A.n161 TG_magic_5.A.n160 0.283032
R406 TG_magic_5.A.n99 TG_magic_5.A.n83 0.282239
R407 TG_magic_5.A.n98 TG_magic_5.A.n94 0.282239
R408 TG_magic_5.A.n51 TG_magic_5.A.n22 0.281892
R409 TG_magic_5.A.n22 TG_magic_5.A.n10 0.279866
R410 TG_magic_5.A.n160 TG_magic_5.A.n159 0.279866
R411 TG_magic_5.A.n50 TG_magic_5.A.n44 0.244078
R412 TG_magic_5.A.n137 TG_magic_5.A.n136 0.244078
R413 TG_magic_5.A.n104 TG_magic_5.A.n103 0.237239
R414 TG_magic_5.A.n65 TG_magic_5.A.n64 0.229487
R415 TG_magic_5.A.n107 TG_magic_5.A.n106 0.211307
R416 TG_magic_5.A.n63 TG_magic_5.A.n62 0.192239
R417 TG_magic_5.A.n64 TG_magic_5.A.n57 0.182457
R418 TG_magic_5.A.n51 TG_magic_5.A.n50 0.1355
R419 TG_magic_5.A.n161 TG_magic_5.A.n137 0.1355
R420 VDD.n783 VDD.n782 327.43
R421 VDD.n390 VDD.t217 73.2007
R422 VDD.n362 VDD.t98 73.2007
R423 VDD.n668 VDD.t88 73.2007
R424 VDD.n680 VDD.t214 73.2007
R425 VDD.n789 VDD.t236 60.5332
R426 VDD.n476 VDD.t287 60.4966
R427 VDD.n437 VDD.t46 60.4966
R428 VDD.n749 VDD.t103 60.4966
R429 VDD.n463 VDD.t52 59.8916
R430 VDD.n424 VDD.t40 59.8916
R431 VDD.n406 VDD.t86 59.8916
R432 VDD.n381 VDD.t241 59.8916
R433 VDD.n717 VDD.t188 59.8916
R434 VDD.n696 VDD.t76 59.8916
R435 VDD.n775 VDD.t297 59.8916
R436 VDD.n736 VDD.t78 59.8916
R437 VDD.n413 VDD.t145 40.6581
R438 VDD.n725 VDD.t150 40.6581
R439 VDD.n410 VDD.t84 40.0531
R440 VDD.n386 VDD.t240 40.0531
R441 VDD.n722 VDD.t106 40.0531
R442 VDD.n673 VDD.t77 40.0531
R443 VDD.n255 VDD.t66 38.634
R444 VDD.n138 VDD.t95 38.634
R445 VDD.n107 VDD.t90 38.634
R446 VDD.n783 VDD.t239 37.5308
R447 VDD.n469 VDD.t289 37.5081
R448 VDD.n451 VDD.t117 37.5081
R449 VDD.n430 VDD.t49 37.5081
R450 VDD.n394 VDD.t166 37.5081
R451 VDD.n369 VDD.t300 37.5081
R452 VDD.n705 VDD.t70 37.5081
R453 VDD.n684 VDD.t112 37.5081
R454 VDD.n763 VDD.t119 37.5081
R455 VDD.n742 VDD.t59 37.5081
R456 VDD.n332 VDD.t183 36.9031
R457 VDD.n463 VDD.t185 36.9031
R458 VDD.n344 VDD.t125 36.9031
R459 VDD.n346 VDD.t45 36.9031
R460 VDD.n424 VDD.t43 36.9031
R461 VDD.n406 VDD.t85 36.9031
R462 VDD.n381 VDD.t175 36.9031
R463 VDD.n717 VDD.t189 36.9031
R464 VDD.n696 VDD.t228 36.9031
R465 VDD.n782 VDD.t295 36.9031
R466 VDD.n775 VDD.t296 36.9031
R467 VDD.n658 VDD.t122 36.9031
R468 VDD.n660 VDD.t82 36.9031
R469 VDD.n736 VDD.t79 36.9031
R470 VDD.n789 VDD.t237 36.3201
R471 VDD.n476 VDD.t290 36.2981
R472 VDD.n437 VDD.t47 36.2981
R473 VDD.n749 VDD.t104 36.2981
R474 VDD.n551 VDD.t159 33.0385
R475 VDD.n240 VDD.t16 31.6097
R476 VDD.n130 VDD.t2 31.6097
R477 VDD.n645 VDD.t234 23.6082
R478 VDD.n478 VDD.t291 23.594
R479 VDD.n439 VDD.t51 23.594
R480 VDD.n751 VDD.t105 23.594
R481 VDD.n461 VDD.t53 22.989
R482 VDD.n422 VDD.t41 22.989
R483 VDD.n404 VDD.t246 22.989
R484 VDD.n379 VDD.t186 22.989
R485 VDD.n715 VDD.t187 22.989
R486 VDD.n694 VDD.t75 22.989
R487 VDD.n773 VDD.t293 22.989
R488 VDD.n734 VDD.t80 22.989
R489 VDD.n229 VDD.t180 22.9462
R490 VDD.n135 VDD.t19 22.6269
R491 VDD.n154 VDD.t7 22.0312
R492 VDD.n572 VDD.t23 21.3909
R493 VDD.n562 VDD.t152 20.3214
R494 VDD.n267 VDD.t4 19.8025
R495 VDD.n246 VDD.t63 19.7962
R496 VDD.n142 VDD.t207 19.7962
R497 VDD.n118 VDD.t107 19.7962
R498 VDD.n32 VDD.t177 19.4769
R499 VDD.n34 VDD.t14 19.4769
R500 VDD.n240 VDD.t12 19.4769
R501 VDD.n130 VDD.t1 19.4769
R502 VDD.n253 VDD.t65 19.1576
R503 VDD.n279 VDD.t57 14.3729
R504 VDD.n457 VDD.t184 13.9146
R505 VDD.n418 VDD.t44 13.9146
R506 VDD.n400 VDD.t87 13.9146
R507 VDD.n375 VDD.t176 13.9146
R508 VDD.n711 VDD.t60 13.9146
R509 VDD.n690 VDD.t174 13.9146
R510 VDD.n769 VDD.t294 13.9146
R511 VDD.n730 VDD.t81 13.9146
R512 VDD.n213 VDD.t27 13.9055
R513 VDD.n442 VDD.t48 13.3096
R514 VDD.n754 VDD.t102 13.3096
R515 VDD.n633 VDD.t238 12.7124
R516 VDD.n488 VDD.t288 12.7047
R517 VDD.n255 VDD.t64 12.4526
R518 VDD.n256 VDD.n254 12.2137
R519 VDD.n241 VDD.n239 12.2137
R520 VDD.n131 VDD.n129 12.2137
R521 VDD.n479 VDD.n477 12.2137
R522 VDD.n464 VDD.n462 12.2137
R523 VDD.n425 VDD.n423 12.2137
R524 VDD.n440 VDD.n438 12.2137
R525 VDD.n407 VDD.n405 12.2137
R526 VDD.n382 VDD.n380 12.2137
R527 VDD.n737 VDD.n735 12.2137
R528 VDD.n752 VDD.n750 12.2137
R529 VDD.n776 VDD.n774 12.2137
R530 VDD.n718 VDD.n716 12.2137
R531 VDD.n697 VDD.n695 12.2137
R532 VDD.n277 VDD.t58 12.1372
R533 VDD.n238 VDD.t15 12.1333
R534 VDD.n152 VDD.t39 12.1333
R535 VDD.n128 VDD.t18 12.1333
R536 VDD.n204 VDD.t34 11.588
R537 VDD.n155 VDD.n153 10.5558
R538 VDD.n280 VDD.n278 9.22945
R539 VDD.n71 VDD.t25 8.618
R540 VDD.n273 VDD.t56 7.3464
R541 VDD.n234 VDD.t11 7.34405
R542 VDD.n148 VDD.t206 7.34405
R543 VDD.n124 VDD.t17 7.34405
R544 VDD.n84 VDD.n83 7.09117
R545 VDD.n258 VDD.t67 7.02477
R546 VDD.n552 VDD.n551 6.3005
R547 VDD.n555 VDD.n554 6.3005
R548 VDD.n554 VDD.n553 6.3005
R549 VDD.n576 VDD.n575 6.3005
R550 VDD.n574 VDD.n573 6.3005
R551 VDD.n573 VDD.n572 6.3005
R552 VDD.n563 VDD.n562 6.3005
R553 VDD.n540 VDD.n539 6.3005
R554 VDD.n571 VDD.n570 6.3005
R555 VDD.n570 VDD.n569 6.3005
R556 VDD.n588 VDD.n587 6.3005
R557 VDD.n587 VDD.n586 6.3005
R558 VDD.n583 VDD.n582 6.3005
R559 VDD.n582 VDD.n581 6.3005
R560 VDD.n591 VDD.n590 6.3005
R561 VDD.n223 VDD.n222 6.3005
R562 VDD.n50 VDD.n49 6.3005
R563 VDD.n212 VDD.n211 6.3005
R564 VDD.n211 VDD.n210 6.3005
R565 VDD.n221 VDD.n220 6.3005
R566 VDD.n52 VDD.n51 6.3005
R567 VDD.n72 VDD.n71 6.3005
R568 VDD.n78 VDD.n77 6.3005
R569 VDD.n77 VDD.n76 6.3005
R570 VDD.n215 VDD.n214 6.3005
R571 VDD.n214 VDD.n213 6.3005
R572 VDD.n198 VDD.n197 6.3005
R573 VDD.n75 VDD.n74 6.3005
R574 VDD.n74 VDD.n73 6.3005
R575 VDD.n206 VDD.n205 6.3005
R576 VDD.n205 VDD.n204 6.3005
R577 VDD.n86 VDD.n85 6.3005
R578 VDD.n169 VDD.n168 6.3005
R579 VDD.n168 VDD.n167 6.3005
R580 VDD.n173 VDD.n172 6.3005
R581 VDD.n171 VDD.n170 6.3005
R582 VDD.n170 VDD.t10 6.3005
R583 VDD.n159 VDD.n158 6.3005
R584 VDD.n158 VDD.n157 6.3005
R585 VDD.n156 VDD.n155 6.3005
R586 VDD.n155 VDD.n154 6.3005
R587 VDD.n280 VDD.n279 6.3005
R588 VDD.n10 VDD.n9 6.3005
R589 VDD.n294 VDD.n293 6.3005
R590 VDD.n298 VDD.n297 6.3005
R591 VDD.n310 VDD.n309 6.3005
R592 VDD.n486 VDD.n485 6.3005
R593 VDD.n484 VDD.n483 6.3005
R594 VDD.n500 VDD.n499 6.3005
R595 VDD.n504 VDD.n503 6.3005
R596 VDD.n517 VDD.n516 6.3005
R597 VDD.n600 VDD.n599 6.3005
R598 VDD.n636 VDD.n635 6.3005
R599 VDD.n616 VDD.n615 6.3005
R600 VDD.n621 VDD.n620 6.3005
R601 VDD.n632 VDD.n631 6.3005
R602 VDD.n226 VDD.n225 6.07044
R603 VDD.n225 VDD.n224 5.76999
R604 VDD.n355 VDD.t305 5.12376
R605 VDD.n538 VDD.n537 5.07789
R606 VDD.n550 VDD.t160 5.07789
R607 VDD.n45 VDD.n43 5.07789
R608 VDD.n48 VDD.n47 5.07789
R609 VDD.n68 VDD.t190 5.07789
R610 VDD.n69 VDD.t26 5.07789
R611 VDD.n101 VDD.t108 5.07789
R612 VDD.n104 VDD.t273 5.07789
R613 VDD.n109 VDD.t213 5.07789
R614 VDD.n112 VDD.t91 5.07789
R615 VDD.n89 VDD.t210 5.07789
R616 VDD.n92 VDD.t254 5.07789
R617 VDD.n95 VDD.t100 5.07789
R618 VDD.n98 VDD.t225 5.07789
R619 VDD.n36 VDD.t280 5.07789
R620 VDD.n39 VDD.t181 5.07789
R621 VDD.n20 VDD.n18 5.07789
R622 VDD.n29 VDD.n28 5.07789
R623 VDD.n12 VDD.t248 5.07789
R624 VDD.n15 VDD.t37 5.07789
R625 VDD.n352 VDD.t168 5.07789
R626 VDD.n359 VDD.t302 5.07789
R627 VDD.n364 VDD.t308 5.07789
R628 VDD.n339 VDD.n337 5.07789
R629 VDD.n348 VDD.t161 5.07789
R630 VDD.n334 VDD.t135 5.07789
R631 VDD.n327 VDD.n325 5.07789
R632 VDD.n677 VDD.t311 5.07789
R633 VDD.n674 VDD.t113 5.07789
R634 VDD.n670 VDD.t221 5.07789
R635 VDD.n665 VDD.t71 5.07789
R636 VDD.n662 VDD.t155 5.07789
R637 VDD.n655 VDD.n654 5.07789
R638 VDD.n648 VDD.t132 5.07789
R639 VDD.n4 VDD.n3 5.07789
R640 VDD.n594 VDD.n593 4.97641
R641 VDD.n185 VDD.n84 4.52963
R642 VDD.n579 VDD.n578 4.5005
R643 VDD.n578 VDD.n577 4.5005
R644 VDD.n561 VDD.n560 4.5005
R645 VDD.n584 VDD.n542 4.5005
R646 VDD.n542 VDD.n541 4.5005
R647 VDD.n558 VDD.n549 4.5005
R648 VDD.n549 VDD.n548 4.5005
R649 VDD.n160 VDD.n88 4.5005
R650 VDD.n88 VDD.n87 4.5005
R651 VDD.n166 VDD.n165 4.5005
R652 VDD.n165 VDD.n164 4.5005
R653 VDD.n176 VDD.n175 4.5005
R654 VDD.n175 VDD.n174 4.5005
R655 VDD.n182 VDD.n181 4.5005
R656 VDD.n181 VDD.n180 4.5005
R657 VDD.n195 VDD.n67 4.5005
R658 VDD.n67 VDD.t203 4.5005
R659 VDD.n209 VDD.n54 4.5005
R660 VDD.n54 VDD.n53 4.5005
R661 VDD.n203 VDD.n56 4.5005
R662 VDD.n56 VDD.n55 4.5005
R663 VDD.n218 VDD.n217 4.5005
R664 VDD.n217 VDD.n216 4.5005
R665 VDD.n296 VDD.n295 4.5005
R666 VDD.n291 VDD.n290 4.5005
R667 VDD.n290 VDD.n289 4.5005
R668 VDD.n307 VDD.n306 4.5005
R669 VDD.n306 VDD.n305 4.5005
R670 VDD.n502 VDD.n501 4.5005
R671 VDD.n497 VDD.n496 4.5005
R672 VDD.n496 VDD.n495 4.5005
R673 VDD.n514 VDD.n513 4.5005
R674 VDD.n513 VDD.n512 4.5005
R675 VDD.n606 VDD.n605 4.5005
R676 VDD.n605 VDD.n604 4.5005
R677 VDD.n618 VDD.n617 4.5005
R678 VDD.n627 VDD.n626 4.5005
R679 VDD.n626 VDD.n625 4.5005
R680 VDD.n538 VDD.n536 4.4205
R681 VDD.n550 VDD.t252 4.4205
R682 VDD.n48 VDD.n46 4.4205
R683 VDD.n45 VDD.n44 4.4205
R684 VDD.n69 VDD.t30 4.4205
R685 VDD.n68 VDD.t195 4.4205
R686 VDD.n106 VDD.t272 4.4205
R687 VDD.n105 VDD.t271 4.4205
R688 VDD.n104 VDD.t274 4.4205
R689 VDD.n103 VDD.t109 4.4205
R690 VDD.n102 VDD.t110 4.4205
R691 VDD.n101 VDD.t111 4.4205
R692 VDD.n114 VDD.t92 4.4205
R693 VDD.n113 VDD.t101 4.4205
R694 VDD.n112 VDD.t222 4.4205
R695 VDD.n111 VDD.t212 4.4205
R696 VDD.n110 VDD.t93 4.4205
R697 VDD.n109 VDD.t224 4.4205
R698 VDD.n94 VDD.t253 4.4205
R699 VDD.n93 VDD.t256 4.4205
R700 VDD.n92 VDD.t255 4.4205
R701 VDD.n91 VDD.t211 4.4205
R702 VDD.n90 VDD.t208 4.4205
R703 VDD.n89 VDD.t209 4.4205
R704 VDD.n100 VDD.t226 4.4205
R705 VDD.n99 VDD.t96 4.4205
R706 VDD.n98 VDD.t216 4.4205
R707 VDD.n97 VDD.t97 4.4205
R708 VDD.n96 VDD.t306 4.4205
R709 VDD.n95 VDD.t220 4.4205
R710 VDD.n41 VDD.t182 4.4205
R711 VDD.n40 VDD.t201 4.4205
R712 VDD.n39 VDD.t231 4.4205
R713 VDD.n38 VDD.t283 4.4205
R714 VDD.n37 VDD.t286 4.4205
R715 VDD.n36 VDD.t275 4.4205
R716 VDD.n31 VDD.n25 4.4205
R717 VDD.n30 VDD.n26 4.4205
R718 VDD.n29 VDD.n27 4.4205
R719 VDD.n24 VDD.n23 4.4205
R720 VDD.n22 VDD.n21 4.4205
R721 VDD.n20 VDD.n19 4.4205
R722 VDD.n17 VDD.t38 4.4205
R723 VDD.n16 VDD.t244 4.4205
R724 VDD.n15 VDD.t31 4.4205
R725 VDD.n14 VDD.t247 4.4205
R726 VDD.n13 VDD.t6 4.4205
R727 VDD.n12 VDD.t5 4.4205
R728 VDD.n354 VDD.t169 4.4205
R729 VDD.n353 VDD.t170 4.4205
R730 VDD.n352 VDD.t167 4.4205
R731 VDD.n358 VDD.t227 4.4205
R732 VDD.n357 VDD.t218 4.4205
R733 VDD.n355 VDD.t312 4.4205
R734 VDD.n361 VDD.t303 4.4205
R735 VDD.n360 VDD.t304 4.4205
R736 VDD.n359 VDD.t301 4.4205
R737 VDD.n366 VDD.t307 4.4205
R738 VDD.n365 VDD.t223 4.4205
R739 VDD.n364 VDD.t99 4.4205
R740 VDD.n343 VDD.n342 4.4205
R741 VDD.n341 VDD.n340 4.4205
R742 VDD.n339 VDD.n338 4.4205
R743 VDD.n350 VDD.t261 4.4205
R744 VDD.n349 VDD.t266 4.4205
R745 VDD.n348 VDD.t146 4.4205
R746 VDD.n336 VDD.t121 4.4205
R747 VDD.n335 VDD.t118 4.4205
R748 VDD.n334 VDD.t134 4.4205
R749 VDD.n331 VDD.n330 4.4205
R750 VDD.n329 VDD.n328 4.4205
R751 VDD.n327 VDD.n326 4.4205
R752 VDD.n679 VDD.t310 4.4205
R753 VDD.n678 VDD.t309 4.4205
R754 VDD.n677 VDD.t215 4.4205
R755 VDD.n676 VDD.t115 4.4205
R756 VDD.n675 VDD.t114 4.4205
R757 VDD.n674 VDD.t116 4.4205
R758 VDD.n672 VDD.t219 4.4205
R759 VDD.n671 VDD.t94 4.4205
R760 VDD.n670 VDD.t89 4.4205
R761 VDD.n667 VDD.t72 4.4205
R762 VDD.n666 VDD.t73 4.4205
R763 VDD.n665 VDD.t74 4.4205
R764 VDD.n664 VDD.t151 4.4205
R765 VDD.n663 VDD.t162 4.4205
R766 VDD.n662 VDD.t249 4.4205
R767 VDD.n657 VDD.n651 4.4205
R768 VDD.n656 VDD.n652 4.4205
R769 VDD.n655 VDD.n653 4.4205
R770 VDD.n650 VDD.t133 4.4205
R771 VDD.n649 VDD.t142 4.4205
R772 VDD.n648 VDD.t120 4.4205
R773 VDD.n6 VDD.n0 4.4205
R774 VDD.n5 VDD.n1 4.4205
R775 VDD.n4 VDD.n2 4.4205
R776 VDD.n541 VDD.t147 4.27857
R777 VDD.n604 VDD.t156 4.23779
R778 VDD.n512 VDD.t20 4.23522
R779 VDD.n87 VDD.t9 4.1512
R780 VDD.n565 VDD.n563 3.8505
R781 VDD.n531 VDD.n530 3.29614
R782 VDD.n547 VDD.n546 3.25789
R783 VDD.n61 VDD.n58 3.25789
R784 VDD.n66 VDD.n65 3.25789
R785 VDD.n566 VDD.n565 3.1505
R786 VDD.n565 VDD.n564 3.1505
R787 VDD.n201 VDD.n200 3.1505
R788 VDD.n200 VDD.n199 3.1505
R789 VDD.n116 VDD.n108 3.1505
R790 VDD.n108 VDD.n107 3.1505
R791 VDD.n134 VDD.n133 3.1505
R792 VDD.n133 VDD.t3 3.1505
R793 VDD.n132 VDD.n131 3.1505
R794 VDD.n131 VDD.n130 3.1505
R795 VDD.n129 VDD.n127 3.1505
R796 VDD.n129 VDD.n128 3.1505
R797 VDD.n126 VDD.n125 3.1505
R798 VDD.n125 VDD.n124 3.1505
R799 VDD.n123 VDD.n122 3.1505
R800 VDD.n122 VDD.n121 3.1505
R801 VDD.n120 VDD.n119 3.1505
R802 VDD.n119 VDD.n118 3.1505
R803 VDD.n136 VDD.n135 3.1505
R804 VDD.n153 VDD.n151 3.1505
R805 VDD.n153 VDD.n152 3.1505
R806 VDD.n150 VDD.n149 3.1505
R807 VDD.n149 VDD.n148 3.1505
R808 VDD.n147 VDD.n146 3.1505
R809 VDD.n146 VDD.n145 3.1505
R810 VDD.n144 VDD.n143 3.1505
R811 VDD.n143 VDD.n142 3.1505
R812 VDD.n140 VDD.n139 3.1505
R813 VDD.n139 VDD.n138 3.1505
R814 VDD.n245 VDD.n35 3.1505
R815 VDD.n35 VDD.n34 3.1505
R816 VDD.n244 VDD.n243 3.1505
R817 VDD.n243 VDD.t13 3.1505
R818 VDD.n242 VDD.n241 3.1505
R819 VDD.n241 VDD.n240 3.1505
R820 VDD.n239 VDD.n237 3.1505
R821 VDD.n239 VDD.n238 3.1505
R822 VDD.n236 VDD.n235 3.1505
R823 VDD.n235 VDD.n234 3.1505
R824 VDD.n233 VDD.n232 3.1505
R825 VDD.n232 VDD.n231 3.1505
R826 VDD.n230 VDD.n229 3.1505
R827 VDD.n264 VDD.n33 3.1505
R828 VDD.n33 VDD.n32 3.1505
R829 VDD.n263 VDD.n262 3.1505
R830 VDD.n262 VDD.n261 3.1505
R831 VDD.n260 VDD.n259 3.1505
R832 VDD.n259 VDD.n258 3.1505
R833 VDD.n257 VDD.n256 3.1505
R834 VDD.n256 VDD.n255 3.1505
R835 VDD.n254 VDD.n252 3.1505
R836 VDD.n254 VDD.n253 3.1505
R837 VDD.n251 VDD.n250 3.1505
R838 VDD.n250 VDD.n249 3.1505
R839 VDD.n248 VDD.n247 3.1505
R840 VDD.n247 VDD.n246 3.1505
R841 VDD.n269 VDD.n268 3.1505
R842 VDD.n268 VDD.n267 3.1505
R843 VDD.n272 VDD.n271 3.1505
R844 VDD.n271 VDD.n270 3.1505
R845 VDD.n275 VDD.n274 3.1505
R846 VDD.n274 VDD.n273 3.1505
R847 VDD.n278 VDD.n276 3.1505
R848 VDD.n278 VDD.n277 3.1505
R849 VDD.n367 VDD.n363 3.1505
R850 VDD.n363 VDD.n362 3.1505
R851 VDD.n385 VDD.n384 3.1505
R852 VDD.n384 VDD.t245 3.1505
R853 VDD.n383 VDD.n382 3.1505
R854 VDD.n382 VDD.n381 3.1505
R855 VDD.n380 VDD.n378 3.1505
R856 VDD.n380 VDD.n379 3.1505
R857 VDD.n377 VDD.n376 3.1505
R858 VDD.n376 VDD.n375 3.1505
R859 VDD.n374 VDD.n373 3.1505
R860 VDD.n373 VDD.n372 3.1505
R861 VDD.n371 VDD.n370 3.1505
R862 VDD.n370 VDD.n369 3.1505
R863 VDD.n387 VDD.n386 3.1505
R864 VDD.n409 VDD.n351 3.1505
R865 VDD.n351 VDD.t299 3.1505
R866 VDD.n408 VDD.n407 3.1505
R867 VDD.n407 VDD.n406 3.1505
R868 VDD.n405 VDD.n403 3.1505
R869 VDD.n405 VDD.n404 3.1505
R870 VDD.n402 VDD.n401 3.1505
R871 VDD.n401 VDD.n400 3.1505
R872 VDD.n399 VDD.n398 3.1505
R873 VDD.n398 VDD.n397 3.1505
R874 VDD.n396 VDD.n395 3.1505
R875 VDD.n395 VDD.n394 3.1505
R876 VDD.n392 VDD.n391 3.1505
R877 VDD.n391 VDD.n390 3.1505
R878 VDD.n411 VDD.n410 3.1505
R879 VDD.n448 VDD.n345 3.1505
R880 VDD.n345 VDD.n344 3.1505
R881 VDD.n447 VDD.n446 3.1505
R882 VDD.n446 VDD.n445 3.1505
R883 VDD.n444 VDD.n443 3.1505
R884 VDD.n443 VDD.n442 3.1505
R885 VDD.n441 VDD.n440 3.1505
R886 VDD.n440 VDD.n439 3.1505
R887 VDD.n438 VDD.n436 3.1505
R888 VDD.n438 VDD.n437 3.1505
R889 VDD.n435 VDD.n434 3.1505
R890 VDD.n434 VDD.n433 3.1505
R891 VDD.n432 VDD.n431 3.1505
R892 VDD.n431 VDD.n430 3.1505
R893 VDD.n429 VDD.n347 3.1505
R894 VDD.n347 VDD.n346 3.1505
R895 VDD.n428 VDD.n427 3.1505
R896 VDD.n427 VDD.t42 3.1505
R897 VDD.n426 VDD.n425 3.1505
R898 VDD.n425 VDD.n424 3.1505
R899 VDD.n423 VDD.n421 3.1505
R900 VDD.n423 VDD.n422 3.1505
R901 VDD.n420 VDD.n419 3.1505
R902 VDD.n419 VDD.n418 3.1505
R903 VDD.n417 VDD.n416 3.1505
R904 VDD.n416 VDD.n415 3.1505
R905 VDD.n414 VDD.n413 3.1505
R906 VDD.n468 VDD.n333 3.1505
R907 VDD.n333 VDD.n332 3.1505
R908 VDD.n467 VDD.n466 3.1505
R909 VDD.n466 VDD.t68 3.1505
R910 VDD.n465 VDD.n464 3.1505
R911 VDD.n464 VDD.n463 3.1505
R912 VDD.n462 VDD.n460 3.1505
R913 VDD.n462 VDD.n461 3.1505
R914 VDD.n459 VDD.n458 3.1505
R915 VDD.n458 VDD.n457 3.1505
R916 VDD.n456 VDD.n455 3.1505
R917 VDD.n455 VDD.n454 3.1505
R918 VDD.n453 VDD.n452 3.1505
R919 VDD.n452 VDD.n451 3.1505
R920 VDD.n471 VDD.n470 3.1505
R921 VDD.n470 VDD.n469 3.1505
R922 VDD.n474 VDD.n473 3.1505
R923 VDD.n473 VDD.n472 3.1505
R924 VDD.n477 VDD.n475 3.1505
R925 VDD.n477 VDD.n476 3.1505
R926 VDD.n480 VDD.n479 3.1505
R927 VDD.n479 VDD.n478 3.1505
R928 VDD.n701 VDD.n673 3.1505
R929 VDD.n700 VDD.n699 3.1505
R930 VDD.n699 VDD.t171 3.1505
R931 VDD.n698 VDD.n697 3.1505
R932 VDD.n697 VDD.n696 3.1505
R933 VDD.n695 VDD.n693 3.1505
R934 VDD.n695 VDD.n694 3.1505
R935 VDD.n692 VDD.n691 3.1505
R936 VDD.n691 VDD.n690 3.1505
R937 VDD.n689 VDD.n688 3.1505
R938 VDD.n688 VDD.n687 3.1505
R939 VDD.n686 VDD.n685 3.1505
R940 VDD.n685 VDD.n684 3.1505
R941 VDD.n682 VDD.n681 3.1505
R942 VDD.n681 VDD.n680 3.1505
R943 VDD.n703 VDD.n669 3.1505
R944 VDD.n669 VDD.n668 3.1505
R945 VDD.n723 VDD.n722 3.1505
R946 VDD.n721 VDD.n720 3.1505
R947 VDD.n720 VDD.t61 3.1505
R948 VDD.n719 VDD.n718 3.1505
R949 VDD.n718 VDD.n717 3.1505
R950 VDD.n716 VDD.n714 3.1505
R951 VDD.n716 VDD.n715 3.1505
R952 VDD.n713 VDD.n712 3.1505
R953 VDD.n712 VDD.n711 3.1505
R954 VDD.n710 VDD.n709 3.1505
R955 VDD.n709 VDD.n708 3.1505
R956 VDD.n707 VDD.n706 3.1505
R957 VDD.n706 VDD.n705 3.1505
R958 VDD.n781 VDD.n780 3.1505
R959 VDD.n782 VDD.n781 3.1505
R960 VDD.n779 VDD.n778 3.1505
R961 VDD.n778 VDD.t298 3.1505
R962 VDD.n777 VDD.n776 3.1505
R963 VDD.n776 VDD.n775 3.1505
R964 VDD.n774 VDD.n772 3.1505
R965 VDD.n774 VDD.n773 3.1505
R966 VDD.n771 VDD.n770 3.1505
R967 VDD.n770 VDD.n769 3.1505
R968 VDD.n768 VDD.n767 3.1505
R969 VDD.n767 VDD.n766 3.1505
R970 VDD.n765 VDD.n764 3.1505
R971 VDD.n764 VDD.n763 3.1505
R972 VDD.n760 VDD.n659 3.1505
R973 VDD.n659 VDD.n658 3.1505
R974 VDD.n759 VDD.n758 3.1505
R975 VDD.n758 VDD.n757 3.1505
R976 VDD.n756 VDD.n755 3.1505
R977 VDD.n755 VDD.n754 3.1505
R978 VDD.n753 VDD.n752 3.1505
R979 VDD.n752 VDD.n751 3.1505
R980 VDD.n750 VDD.n748 3.1505
R981 VDD.n750 VDD.n749 3.1505
R982 VDD.n747 VDD.n746 3.1505
R983 VDD.n746 VDD.n745 3.1505
R984 VDD.n744 VDD.n743 3.1505
R985 VDD.n743 VDD.n742 3.1505
R986 VDD.n741 VDD.n661 3.1505
R987 VDD.n661 VDD.n660 3.1505
R988 VDD.n740 VDD.n739 3.1505
R989 VDD.n739 VDD.t83 3.1505
R990 VDD.n738 VDD.n737 3.1505
R991 VDD.n737 VDD.n736 3.1505
R992 VDD.n735 VDD.n733 3.1505
R993 VDD.n735 VDD.n734 3.1505
R994 VDD.n732 VDD.n731 3.1505
R995 VDD.n731 VDD.n730 3.1505
R996 VDD.n729 VDD.n728 3.1505
R997 VDD.n728 VDD.n727 3.1505
R998 VDD.n726 VDD.n725 3.1505
R999 VDD.n647 VDD.n646 3.1505
R1000 VDD.n646 VDD.n645 3.1505
R1001 VDD.n791 VDD.n790 3.1505
R1002 VDD.n790 VDD.n789 3.1505
R1003 VDD.n788 VDD.n787 3.1505
R1004 VDD.n787 VDD.n786 3.1505
R1005 VDD.n785 VDD.n784 3.1505
R1006 VDD.n784 VDD.n783 3.1505
R1007 VDD.n284 VDD.n10 2.92945
R1008 VDD.n281 VDD.n280 2.92945
R1009 VDD.n490 VDD.n484 2.92945
R1010 VDD.n487 VDD.n486 2.92945
R1011 VDD.n638 VDD.n632 2.92945
R1012 VDD.n637 VDD.n636 2.92945
R1013 VDD.n547 VDD.n544 2.6005
R1014 VDD.n61 VDD.n60 2.6005
R1015 VDD.n66 VDD.n63 2.6005
R1016 VDD.n9 VDD.t0 2.55559
R1017 VDD.n296 VDD.n294 2.48734
R1018 VDD.n502 VDD.n500 2.48734
R1019 VDD.n618 VDD.n616 2.48734
R1020 VDD.n558 VDD.n557 2.363
R1021 VDD.n299 VDD.n298 2.32155
R1022 VDD.n506 VDD.n504 2.32155
R1023 VDD.n622 VDD.n621 2.32155
R1024 VDD.n643 VDD.n642 2.31102
R1025 VDD.n195 VDD.n194 2.2505
R1026 VDD.n322 VDD.n314 2.2505
R1027 VDD.n530 VDD.n522 2.2505
R1028 VDD.n614 VDD.n613 2.2505
R1029 VDD.n596 VDD.n595 2.2505
R1030 VDD.n305 VDD.t55 2.23621
R1031 VDD.n285 VDD.n284 2.1005
R1032 VDD.n284 VDD.n283 2.1005
R1033 VDD.n313 VDD.n312 2.1005
R1034 VDD.n300 VDD.n299 2.1005
R1035 VDD.n299 VDD.t54 2.1005
R1036 VDD.n491 VDD.n490 2.1005
R1037 VDD.n490 VDD.n489 2.1005
R1038 VDD.n506 VDD.n505 2.1005
R1039 VDD.n520 VDD.n519 2.1005
R1040 VDD.n507 VDD.n506 2.1005
R1041 VDD.n602 VDD.n601 2.1005
R1042 VDD.n638 VDD.n634 2.1005
R1043 VDD.n622 VDD.n619 2.1005
R1044 VDD.n623 VDD.n622 2.1005
R1045 VDD.n639 VDD.n638 2.1005
R1046 VDD.n228 VDD.n227 2.04726
R1047 VDD.n544 VDD.t24 1.8205
R1048 VDD.n544 VDD.n543 1.8205
R1049 VDD.n546 VDD.t163 1.8205
R1050 VDD.n546 VDD.n545 1.8205
R1051 VDD.n63 VDD.t36 1.8205
R1052 VDD.n63 VDD.n62 1.8205
R1053 VDD.n65 VDD.t35 1.8205
R1054 VDD.n65 VDD.n64 1.8205
R1055 VDD.n60 VDD.t202 1.8205
R1056 VDD.n60 VDD.n59 1.8205
R1057 VDD.n58 VDD.t198 1.8205
R1058 VDD.n58 VDD.n57 1.8205
R1059 VDD.n175 VDD.n173 1.71366
R1060 VDD.n595 VDD.n594 1.66585
R1061 VDD.n88 VDD.n86 1.65839
R1062 VDD.n594 VDD.n534 1.55581
R1063 VDD.n227 VDD.n226 1.50398
R1064 VDD.n312 VDD.n310 1.27155
R1065 VDD.n519 VDD.n517 1.27155
R1066 VDD.n601 VDD.n600 1.27155
R1067 VDD.n534 VDD.n324 1.14521
R1068 VDD.n593 VDD.n592 1.13368
R1069 VDD.n193 VDD.n185 1.1255
R1070 VDD.n194 VDD.n193 1.07177
R1071 VDD.n200 VDD.n198 1.00582
R1072 VDD.n299 VDD.n296 0.995237
R1073 VDD.n506 VDD.n502 0.995237
R1074 VDD.n622 VDD.n618 0.995237
R1075 VDD.n180 VDD.t8 0.958354
R1076 VDD.n542 VDD.n540 0.8405
R1077 VDD.n358 VDD.n357 0.703756
R1078 VDD.n102 VDD.n101 0.657891
R1079 VDD.n103 VDD.n102 0.657891
R1080 VDD.n106 VDD.n105 0.657891
R1081 VDD.n105 VDD.n104 0.657891
R1082 VDD.n110 VDD.n109 0.657891
R1083 VDD.n111 VDD.n110 0.657891
R1084 VDD.n114 VDD.n113 0.657891
R1085 VDD.n113 VDD.n112 0.657891
R1086 VDD.n90 VDD.n89 0.657891
R1087 VDD.n91 VDD.n90 0.657891
R1088 VDD.n94 VDD.n93 0.657891
R1089 VDD.n93 VDD.n92 0.657891
R1090 VDD.n96 VDD.n95 0.657891
R1091 VDD.n97 VDD.n96 0.657891
R1092 VDD.n100 VDD.n99 0.657891
R1093 VDD.n99 VDD.n98 0.657891
R1094 VDD.n37 VDD.n36 0.657891
R1095 VDD.n38 VDD.n37 0.657891
R1096 VDD.n41 VDD.n40 0.657891
R1097 VDD.n40 VDD.n39 0.657891
R1098 VDD.n22 VDD.n20 0.657891
R1099 VDD.n24 VDD.n22 0.657891
R1100 VDD.n31 VDD.n30 0.657891
R1101 VDD.n30 VDD.n29 0.657891
R1102 VDD.n13 VDD.n12 0.657891
R1103 VDD.n14 VDD.n13 0.657891
R1104 VDD.n17 VDD.n16 0.657891
R1105 VDD.n16 VDD.n15 0.657891
R1106 VDD.n353 VDD.n352 0.657891
R1107 VDD.n354 VDD.n353 0.657891
R1108 VDD.n360 VDD.n359 0.657891
R1109 VDD.n361 VDD.n360 0.657891
R1110 VDD.n365 VDD.n364 0.657891
R1111 VDD.n366 VDD.n365 0.657891
R1112 VDD.n341 VDD.n339 0.657891
R1113 VDD.n343 VDD.n341 0.657891
R1114 VDD.n349 VDD.n348 0.657891
R1115 VDD.n350 VDD.n349 0.657891
R1116 VDD.n335 VDD.n334 0.657891
R1117 VDD.n336 VDD.n335 0.657891
R1118 VDD.n329 VDD.n327 0.657891
R1119 VDD.n331 VDD.n329 0.657891
R1120 VDD.n679 VDD.n678 0.657891
R1121 VDD.n678 VDD.n677 0.657891
R1122 VDD.n676 VDD.n675 0.657891
R1123 VDD.n675 VDD.n674 0.657891
R1124 VDD.n672 VDD.n671 0.657891
R1125 VDD.n671 VDD.n670 0.657891
R1126 VDD.n667 VDD.n666 0.657891
R1127 VDD.n666 VDD.n665 0.657891
R1128 VDD.n664 VDD.n663 0.657891
R1129 VDD.n663 VDD.n662 0.657891
R1130 VDD.n657 VDD.n656 0.657891
R1131 VDD.n656 VDD.n655 0.657891
R1132 VDD.n650 VDD.n649 0.657891
R1133 VDD.n649 VDD.n648 0.657891
R1134 VDD.n6 VDD.n5 0.657891
R1135 VDD.n5 VDD.n4 0.657891
R1136 VDD.n84 VDD.n82 0.620741
R1137 VDD.n634 VDD.n633 0.605827
R1138 VDD.n786 VDD.t235 0.605827
R1139 VDD.n489 VDD.n488 0.605461
R1140 VDD.n472 VDD.t292 0.605461
R1141 VDD.n433 VDD.t50 0.605461
R1142 VDD.n745 VDD.t69 0.605461
R1143 VDD.n367 VDD.n366 0.575987
R1144 VDD.n682 VDD.n679 0.575987
R1145 VDD.n578 VDD.n576 0.5605
R1146 VDD.n565 VDD.n561 0.5605
R1147 VDD.n389 VDD.n358 0.504919
R1148 VDD.n356 VDD.n355 0.502826
R1149 VDD.n82 VDD.n81 0.497868
R1150 VDD.n552 VDD.n550 0.486111
R1151 VDD.n117 VDD.n103 0.472022
R1152 VDD.n117 VDD.n106 0.472022
R1153 VDD.n115 VDD.n111 0.472022
R1154 VDD.n115 VDD.n114 0.472022
R1155 VDD.n141 VDD.n91 0.472022
R1156 VDD.n141 VDD.n94 0.472022
R1157 VDD.n137 VDD.n97 0.472022
R1158 VDD.n137 VDD.n100 0.472022
R1159 VDD.n228 VDD.n38 0.472022
R1160 VDD.n228 VDD.n41 0.472022
R1161 VDD.n265 VDD.n24 0.472022
R1162 VDD.n265 VDD.n31 0.472022
R1163 VDD.n266 VDD.n14 0.472022
R1164 VDD.n266 VDD.n17 0.472022
R1165 VDD.n393 VDD.n354 0.472022
R1166 VDD.n368 VDD.n361 0.472022
R1167 VDD.n449 VDD.n343 0.472022
R1168 VDD.n412 VDD.n350 0.472022
R1169 VDD.n450 VDD.n336 0.472022
R1170 VDD.n521 VDD.n331 0.472022
R1171 VDD.n683 VDD.n676 0.472022
R1172 VDD.n704 VDD.n667 0.472022
R1173 VDD.n761 VDD.n657 0.472022
R1174 VDD.n762 VDD.n650 0.472022
R1175 VDD.n597 VDD.n6 0.472022
R1176 VDD.n724 VDD.n664 0.468109
R1177 VDD.n702 VDD.n672 0.460283
R1178 VDD.n591 VDD.n538 0.4505
R1179 VDD.n567 VDD.n547 0.4505
R1180 VDD.n412 VDD.n411 0.447829
R1181 VDD.n724 VDD.n723 0.443214
R1182 VDD.n219 VDD.n45 0.440717
R1183 VDD.n219 VDD.n48 0.440717
R1184 VDD.n202 VDD.n61 0.440717
R1185 VDD.n202 VDD.n66 0.440717
R1186 VDD.n70 VDD.n68 0.440717
R1187 VDD.n70 VDD.n69 0.440717
R1188 VDD.n137 VDD.n136 0.347792
R1189 VDD.n702 VDD.n701 0.339547
R1190 VDD.n388 VDD.n387 0.327362
R1191 VDD.n283 VDD.n282 0.319887
R1192 VDD.n249 VDD.t62 0.319785
R1193 VDD.n590 VDD.n589 0.309088
R1194 VDD.n471 VDD.n468 0.281105
R1195 VDD.n323 VDD.n322 0.271017
R1196 VDD.n54 VDD.n52 0.268585
R1197 VDD.n266 VDD.n265 0.261967
R1198 VDD.n248 VDD.n245 0.25161
R1199 VDD.n312 VDD.n311 0.234007
R1200 VDD.n762 VDD.n761 0.233259
R1201 VDD.n450 VDD.n449 0.231954
R1202 VDD.n432 VDD.n429 0.224983
R1203 VDD.n744 VDD.n741 0.224983
R1204 VDD.n52 VDD.n50 0.201564
R1205 VDD.n357 VDD.n356 0.20143
R1206 VDD.n519 VDD.n518 0.148469
R1207 VDD.n601 VDD.n598 0.1484
R1208 VDD.n785 VDD 0.144706
R1209 VDD.n780 VDD 0.136899
R1210 VDD.n136 VDD.n134 0.11481
R1211 VDD.n134 VDD.n132 0.11481
R1212 VDD.n127 VDD.n126 0.11481
R1213 VDD.n126 VDD.n123 0.11481
R1214 VDD.n123 VDD.n120 0.11481
R1215 VDD.n151 VDD.n150 0.11481
R1216 VDD.n150 VDD.n147 0.11481
R1217 VDD.n147 VDD.n144 0.11481
R1218 VDD.n245 VDD.n244 0.11481
R1219 VDD.n244 VDD.n242 0.11481
R1220 VDD.n237 VDD.n236 0.11481
R1221 VDD.n236 VDD.n233 0.11481
R1222 VDD.n233 VDD.n230 0.11481
R1223 VDD.n264 VDD.n263 0.11481
R1224 VDD.n263 VDD.n260 0.11481
R1225 VDD.n260 VDD.n257 0.11481
R1226 VDD.n252 VDD.n251 0.11481
R1227 VDD.n251 VDD.n248 0.11481
R1228 VDD.n276 VDD.n275 0.11481
R1229 VDD.n275 VDD.n272 0.11481
R1230 VDD.n272 VDD.n269 0.11481
R1231 VDD.n387 VDD.n385 0.11481
R1232 VDD.n385 VDD.n383 0.11481
R1233 VDD.n378 VDD.n377 0.11481
R1234 VDD.n377 VDD.n374 0.11481
R1235 VDD.n374 VDD.n371 0.11481
R1236 VDD.n411 VDD.n409 0.11481
R1237 VDD.n409 VDD.n408 0.11481
R1238 VDD.n403 VDD.n402 0.11481
R1239 VDD.n402 VDD.n399 0.11481
R1240 VDD.n399 VDD.n396 0.11481
R1241 VDD.n448 VDD.n447 0.11481
R1242 VDD.n447 VDD.n444 0.11481
R1243 VDD.n444 VDD.n441 0.11481
R1244 VDD.n436 VDD.n435 0.11481
R1245 VDD.n435 VDD.n432 0.11481
R1246 VDD.n429 VDD.n428 0.11481
R1247 VDD.n428 VDD.n426 0.11481
R1248 VDD.n421 VDD.n420 0.11481
R1249 VDD.n420 VDD.n417 0.11481
R1250 VDD.n417 VDD.n414 0.11481
R1251 VDD.n468 VDD.n467 0.11481
R1252 VDD.n467 VDD.n465 0.11481
R1253 VDD.n460 VDD.n459 0.11481
R1254 VDD.n459 VDD.n456 0.11481
R1255 VDD.n456 VDD.n453 0.11481
R1256 VDD.n475 VDD.n474 0.11481
R1257 VDD.n474 VDD.n471 0.11481
R1258 VDD.n701 VDD.n700 0.11481
R1259 VDD.n700 VDD.n698 0.11481
R1260 VDD.n693 VDD.n692 0.11481
R1261 VDD.n692 VDD.n689 0.11481
R1262 VDD.n689 VDD.n686 0.11481
R1263 VDD.n723 VDD.n721 0.11481
R1264 VDD.n721 VDD.n719 0.11481
R1265 VDD.n714 VDD.n713 0.11481
R1266 VDD.n713 VDD.n710 0.11481
R1267 VDD.n710 VDD.n707 0.11481
R1268 VDD.n780 VDD.n779 0.11481
R1269 VDD.n779 VDD.n777 0.11481
R1270 VDD.n772 VDD.n771 0.11481
R1271 VDD.n771 VDD.n768 0.11481
R1272 VDD.n768 VDD.n765 0.11481
R1273 VDD.n760 VDD.n759 0.11481
R1274 VDD.n759 VDD.n756 0.11481
R1275 VDD.n756 VDD.n753 0.11481
R1276 VDD.n748 VDD.n747 0.11481
R1277 VDD.n747 VDD.n744 0.11481
R1278 VDD.n741 VDD.n740 0.11481
R1279 VDD.n740 VDD.n738 0.11481
R1280 VDD.n733 VDD.n732 0.11481
R1281 VDD.n732 VDD.n729 0.11481
R1282 VDD.n791 VDD.n788 0.11481
R1283 VDD.n788 VDD.n785 0.11481
R1284 VDD.n556 VDD.n535 0.1148
R1285 VDD.n729 VDD.n726 0.114781
R1286 VDD.n252 VDD 0.114293
R1287 VDD.n436 VDD 0.114293
R1288 VDD.n475 VDD 0.114293
R1289 VDD.n748 VDD 0.114293
R1290 VDD VDD.n791 0.114293
R1291 VDD.n132 VDD 0.113776
R1292 VDD.n242 VDD 0.113776
R1293 VDD.n383 VDD 0.113776
R1294 VDD.n408 VDD 0.113776
R1295 VDD.n426 VDD 0.113776
R1296 VDD.n465 VDD 0.113776
R1297 VDD.n698 VDD 0.113776
R1298 VDD.n719 VDD 0.113776
R1299 VDD.n777 VDD 0.113776
R1300 VDD.n738 VDD 0.113776
R1301 VDD.n117 VDD.n116 0.1055
R1302 VDD.n141 VDD.n140 0.1055
R1303 VDD.n368 VDD.n367 0.1055
R1304 VDD.n393 VDD.n392 0.1055
R1305 VDD.n683 VDD.n682 0.1055
R1306 VDD.n704 VDD.n703 0.104914
R1307 VDD.n116 VDD.n115 0.104466
R1308 VDD.n140 VDD.n137 0.104466
R1309 VDD.n557 VDD.n556 0.104
R1310 VDD.n392 VDD.n389 0.103948
R1311 VDD.n703 VDD.n702 0.101
R1312 VDD.n156 VDD 0.0982586
R1313 VDD.n80 VDD.n79 0.08978
R1314 VDD.n481 VDD.n480 0.0868793
R1315 VDD.n647 VDD.n644 0.0868793
R1316 VDD VDD.n11 0.0858448
R1317 VDD.n194 VDD.n80 0.08546
R1318 VDD.n227 VDD.n42 0.0819014
R1319 VDD.n79 VDD.n42 0.07898
R1320 VDD.n593 VDD.n535 0.073624
R1321 VDD.n534 VDD.n533 0.0577254
R1322 VDD.n319 VDD.n318 0.0563621
R1323 VDD.n527 VDD.n526 0.0563621
R1324 VDD.n613 VDD.n612 0.0563621
R1325 VDD.n284 VDD.n281 0.0557632
R1326 VDD.n490 VDD.n487 0.0557632
R1327 VDD.n638 VDD.n637 0.0557632
R1328 VDD.n189 VDD.n188 0.0551243
R1329 VDD.n322 VDD.n321 0.0548103
R1330 VDD.n530 VDD.n529 0.0548103
R1331 VDD.n193 VDD.n192 0.054604
R1332 VDD.n558 VDD.n555 0.0522986
R1333 VDD.n318 VDD.n317 0.0501552
R1334 VDD.n526 VDD.n525 0.0501552
R1335 VDD.n72 VDD.n70 0.048
R1336 VDD.n190 VDD.n189 0.0462803
R1337 VDD.n584 VDD.n583 0.0419389
R1338 VDD.n559 VDD.n558 0.0406439
R1339 VDD.n555 VDD.n552 0.0406439
R1340 VDD.n206 VDD.n203 0.03925
R1341 VDD.n78 VDD.n75 0.03925
R1342 VDD.n579 VDD.n574 0.0374065
R1343 VDD.n571 VDD.n568 0.0374065
R1344 VDD.n196 VDD.n195 0.037375
R1345 VDD.n75 VDD.n72 0.037375
R1346 VDD.n583 VDD.n580 0.0361115
R1347 VDD.n218 VDD.n215 0.034875
R1348 VDD.n207 VDD.n206 0.034875
R1349 VDD.n588 VDD.n585 0.0348165
R1350 VDD VDD.n559 0.0348165
R1351 VDD.n303 VDD.n302 0.0330862
R1352 VDD.n287 VDD.n286 0.0330862
R1353 VDD.n510 VDD.n509 0.0330862
R1354 VDD.n493 VDD.n492 0.0330862
R1355 VDD.n609 VDD.n608 0.0330862
R1356 VDD.n630 VDD.n629 0.0330862
R1357 VDD.n212 VDD.n209 0.033
R1358 VDD.n219 VDD.n218 0.031125
R1359 VDD.n178 VDD.n177 0.0299828
R1360 VDD.n162 VDD.n161 0.0299828
R1361 VDD.n324 VDD.n7 0.0294655
R1362 VDD.n532 VDD.n531 0.0292534
R1363 VDD.n533 VDD.n532 0.0292534
R1364 VDD.n324 VDD.n323 0.028431
R1365 VDD.n286 VDD.n285 0.0279138
R1366 VDD.n11 VDD.n8 0.0279138
R1367 VDD.n492 VDD.n491 0.0279138
R1368 VDD.n482 VDD.n481 0.0279138
R1369 VDD.n639 VDD.n630 0.0279138
R1370 VDD.n644 VDD.n643 0.0279138
R1371 VDD.n195 VDD.n78 0.027375
R1372 VDD.n169 VDD.n166 0.0263621
R1373 VDD.n183 VDD.n182 0.0258448
R1374 VDD.n160 VDD.n159 0.0253276
R1375 VDD.n176 VDD.n171 0.0248103
R1376 VDD.n592 VDD.n591 0.0244568
R1377 VDD.n185 VDD.n184 0.0242931
R1378 VDD.n203 VDD.n202 0.02425
R1379 VDD.n308 VDD.n307 0.0237759
R1380 VDD.n302 VDD.n301 0.0237759
R1381 VDD.n515 VDD.n514 0.0237759
R1382 VDD.n509 VDD.n508 0.0237759
R1383 VDD.n606 VDD.n603 0.0237759
R1384 VDD.n614 VDD.n609 0.0237759
R1385 VDD.n300 VDD.n292 0.0222241
R1386 VDD.n507 VDD.n498 0.0222241
R1387 VDD.n624 VDD.n623 0.0222241
R1388 VDD.n226 VDD.n223 0.0205
R1389 VDD.n314 VDD.n313 0.0196379
R1390 VDD.n292 VDD.n291 0.0191207
R1391 VDD.n498 VDD.n497 0.0191207
R1392 VDD.n627 VDD.n624 0.0191207
R1393 VDD.n177 VDD.n176 0.0165345
R1394 VDD.n161 VDD.n160 0.0160172
R1395 VDD.n159 VDD.n156 0.0160172
R1396 VDD.n291 VDD.n288 0.0129138
R1397 VDD.n317 VDD.n316 0.0129138
R1398 VDD.n497 VDD.n494 0.0129138
R1399 VDD.n525 VDD.n524 0.0129138
R1400 VDD.n641 VDD.n640 0.0129138
R1401 VDD.n628 VDD.n627 0.0129138
R1402 VDD.n187 VDD.n186 0.0124653
R1403 VDD.n163 VDD.n162 0.0123966
R1404 VDD.n313 VDD.n308 0.0123966
R1405 VDD.n520 VDD.n515 0.0123966
R1406 VDD.n603 VDD.n602 0.0123966
R1407 VDD.n389 VDD.n388 0.0123621
R1408 VDD.n191 VDD.n190 0.0119451
R1409 VDD.n179 VDD.n178 0.0118793
R1410 VDD.n265 VDD.n264 0.0103276
R1411 VDD.n449 VDD.n448 0.0103276
R1412 VDD.n521 VDD.n520 0.0103276
R1413 VDD.n761 VDD.n760 0.0103276
R1414 VDD.n602 VDD.n597 0.0103276
R1415 VDD.n120 VDD.n117 0.00981034
R1416 VDD.n144 VDD.n141 0.00981034
R1417 VDD.n230 VDD.n228 0.00981034
R1418 VDD.n301 VDD.n300 0.00981034
R1419 VDD.n269 VDD.n266 0.00981034
R1420 VDD.n371 VDD.n368 0.00981034
R1421 VDD.n396 VDD.n393 0.00981034
R1422 VDD.n414 VDD.n412 0.00981034
R1423 VDD.n453 VDD.n450 0.00981034
R1424 VDD.n522 VDD.n521 0.00981034
R1425 VDD.n508 VDD.n507 0.00981034
R1426 VDD.n686 VDD.n683 0.00981034
R1427 VDD.n707 VDD.n704 0.00981034
R1428 VDD.n765 VDD.n762 0.00981034
R1429 VDD.n597 VDD.n596 0.00981034
R1430 VDD.n623 VDD.n614 0.00981034
R1431 VDD.n726 VDD.n724 0.00970455
R1432 VDD VDD.n196 0.008625
R1433 VDD.n585 VDD.n584 0.00826978
R1434 VDD.n307 VDD.n304 0.00825862
R1435 VDD.n321 VDD.n320 0.00825862
R1436 VDD.n514 VDD.n511 0.00825862
R1437 VDD.n529 VDD.n528 0.00825862
R1438 VDD.n611 VDD.n610 0.00825862
R1439 VDD.n607 VDD.n606 0.00825862
R1440 VDD.n591 VDD.n588 0.0076223
R1441 VDD.n221 VDD.n219 0.007375
R1442 VDD.n304 VDD.n303 0.0067069
R1443 VDD.n320 VDD.n319 0.0067069
R1444 VDD.n511 VDD.n510 0.0067069
R1445 VDD.n528 VDD.n527 0.0067069
R1446 VDD.n612 VDD.n611 0.0067069
R1447 VDD.n608 VDD.n607 0.0067069
R1448 VDD.n580 VDD.n579 0.00567986
R1449 VDD.n184 VDD.n183 0.00515517
R1450 VDD.n171 VDD.n169 0.00463793
R1451 VDD.n567 VDD.n566 0.00438489
R1452 VDD.n202 VDD.n201 0.00425
R1453 VDD.n192 VDD.n191 0.00362139
R1454 VDD.n182 VDD.n179 0.00360345
R1455 VDD.n188 VDD.n187 0.00310116
R1456 VDD.n166 VDD.n163 0.00308621
R1457 VDD.n209 VDD.n208 0.003
R1458 VDD.n208 VDD.n207 0.002375
R1459 VDD.n288 VDD.n287 0.00205172
R1460 VDD.n316 VDD.n315 0.00205172
R1461 VDD.n494 VDD.n493 0.00205172
R1462 VDD.n524 VDD.n523 0.00205172
R1463 VDD.n642 VDD.n641 0.00205172
R1464 VDD.n629 VDD.n628 0.00205172
R1465 VDD.n568 VDD.n567 0.00179496
R1466 VDD.n566 VDD 0.00179496
R1467 VDD.n223 VDD.n221 0.00175
R1468 VDD.n215 VDD.n212 0.00175
R1469 VDD.n201 VDD 0.00175
R1470 VDD.n127 VDD 0.00153448
R1471 VDD.n151 VDD 0.00153448
R1472 VDD.n237 VDD 0.00153448
R1473 VDD.n276 VDD 0.00153448
R1474 VDD.n378 VDD 0.00153448
R1475 VDD.n403 VDD 0.00153448
R1476 VDD.n421 VDD 0.00153448
R1477 VDD.n460 VDD 0.00153448
R1478 VDD.n693 VDD 0.00153448
R1479 VDD.n714 VDD 0.00153448
R1480 VDD.n772 VDD 0.00153448
R1481 VDD.n733 VDD 0.00153448
R1482 VDD.n574 VDD.n571 0.00114748
R1483 VDD.n257 VDD 0.00101724
R1484 VDD.n285 VDD.n8 0.00101724
R1485 VDD.n441 VDD 0.00101724
R1486 VDD.n491 VDD.n482 0.00101724
R1487 VDD.n480 VDD 0.00101724
R1488 VDD.n753 VDD 0.00101724
R1489 VDD.n643 VDD.n639 0.00101724
R1490 VDD VDD.n647 0.00101724
R1491 a_n4297_n4860.t12 a_n4297_n4860.n30 40.7345
R1492 a_n4297_n4860.n7 a_n4297_n4860.n6 28.094
R1493 a_n4297_n4860.n16 a_n4297_n4860.n15 28.094
R1494 a_n4297_n4860.n32 a_n4297_n4860.n31 28.094
R1495 a_n4297_n4860.n4 a_n4297_n4860.t7 21.9005
R1496 a_n4297_n4860.n2 a_n4297_n4860.t26 21.9005
R1497 a_n4297_n4860.n1 a_n4297_n4860.t29 21.9005
R1498 a_n4297_n4860.n10 a_n4297_n4860.t11 21.9005
R1499 a_n4297_n4860.n10 a_n4297_n4860.t19 21.9005
R1500 a_n4297_n4860.n22 a_n4297_n4860.t28 21.9005
R1501 a_n4297_n4860.n23 a_n4297_n4860.t25 21.9005
R1502 a_n4297_n4860.n11 a_n4297_n4860.t15 21.9005
R1503 a_n4297_n4860.n11 a_n4297_n4860.t8 21.9005
R1504 a_n4297_n4860.n3 a_n4297_n4860.t10 21.9005
R1505 a_n4297_n4860.n12 a_n4297_n4860.t18 21.9005
R1506 a_n4297_n4860.n12 a_n4297_n4860.t23 21.9005
R1507 a_n4297_n4860.n24 a_n4297_n4860.t9 21.9005
R1508 a_n4297_n4860.n25 a_n4297_n4860.t6 21.9005
R1509 a_n4297_n4860.n13 a_n4297_n4860.t21 21.9005
R1510 a_n4297_n4860.n13 a_n4297_n4860.t14 21.9005
R1511 a_n4297_n4860.n6 a_n4297_n4860.t13 21.9005
R1512 a_n4297_n4860.n15 a_n4297_n4860.t24 21.9005
R1513 a_n4297_n4860.n15 a_n4297_n4860.t20 21.9005
R1514 a_n4297_n4860.n5 a_n4297_n4860.t17 21.9005
R1515 a_n4297_n4860.n14 a_n4297_n4860.t22 21.9005
R1516 a_n4297_n4860.n14 a_n4297_n4860.t27 21.9005
R1517 a_n4297_n4860.n26 a_n4297_n4860.t16 21.9005
R1518 a_n4297_n4860.n31 a_n4297_n4860.t12 21.9005
R1519 a_n4297_n4860.n31 a_n4297_n4860.n26 15.8172
R1520 a_n4297_n4860.n14 a_n4297_n4860.n13 15.8172
R1521 a_n4297_n4860.n26 a_n4297_n4860.n25 15.8172
R1522 a_n4297_n4860.n25 a_n4297_n4860.n24 15.8172
R1523 a_n4297_n4860.n13 a_n4297_n4860.n12 15.8172
R1524 a_n4297_n4860.n12 a_n4297_n4860.n11 15.8172
R1525 a_n4297_n4860.n24 a_n4297_n4860.n23 15.8172
R1526 a_n4297_n4860.n23 a_n4297_n4860.n22 15.8172
R1527 a_n4297_n4860.n11 a_n4297_n4860.n10 15.8172
R1528 a_n4297_n4860.n2 a_n4297_n4860.n1 15.8172
R1529 a_n4297_n4860.n4 a_n4297_n4860.n3 15.8172
R1530 a_n4297_n4860.n3 a_n4297_n4860.n2 15.8172
R1531 a_n4297_n4860.n15 a_n4297_n4860.n14 15.8172
R1532 a_n4297_n4860.n6 a_n4297_n4860.n5 15.8172
R1533 a_n4297_n4860.n5 a_n4297_n4860.n4 15.8172
R1534 a_n4297_n4860.n28 a_n4297_n4860.n27 15.1845
R1535 a_n4297_n4860.n30 a_n4297_n4860.n29 15.1845
R1536 a_n4297_n4860.n29 a_n4297_n4860.n28 15.1845
R1537 a_n4297_n4860.n20 a_n4297_n4860.n19 5.44589
R1538 a_n4297_n4860.n20 a_n4297_n4860.n18 4.7885
R1539 a_n4297_n4860.n7 a_n4297_n4860.n0 4.70615
R1540 a_n4297_n4860.n21 a_n4297_n4860.n17 4.4205
R1541 a_n4297_n4860.n9 a_n4297_n4860.n8 4.4205
R1542 a_n4297_n4860.n34 a_n4297_n4860.n33 4.4205
R1543 a_n4297_n4860.n21 a_n4297_n4860.n20 1.1392
R1544 a_n4297_n4860.n16 a_n4297_n4860.n9 0.286152
R1545 a_n4297_n4860.n33 a_n4297_n4860.n32 0.286152
R1546 a_n4297_n4860.n32 a_n4297_n4860.n21 0.282239
R1547 a_n4297_n4860.n9 a_n4297_n4860.n7 0.282239
R1548 a_n4297_n4860.n33 a_n4297_n4860.n16 0.282239
R1549 A3.n47 A3.n45 5.44589
R1550 A3.n26 A3.n25 5.07789
R1551 A3.n51 A3.t29 4.7885
R1552 A3.n50 A3.t28 4.7885
R1553 A3.n47 A3.n46 4.7885
R1554 A3.n31 A3.t19 4.4205
R1555 A3.n32 A3.t16 4.4205
R1556 A3.n33 A3.t14 4.4205
R1557 A3.n34 A3.t20 4.4205
R1558 A3.n28 A3.n22 4.4205
R1559 A3.n27 A3.n23 4.4205
R1560 A3.n26 A3.n24 4.4205
R1561 A3.n44 A3.n41 3.80789
R1562 A3.n39 A3.n36 3.80789
R1563 A3.n8 A3.n7 3.25789
R1564 A3.n19 A3.n18 3.25789
R1565 A3.n44 A3.n43 3.1505
R1566 A3.n39 A3.n38 3.1505
R1567 A3.n8 A3.n5 2.6005
R1568 A3.n9 A3.n3 2.6005
R1569 A3.n10 A3.n1 2.6005
R1570 A3.n19 A3.n16 2.6005
R1571 A3.n20 A3.n14 2.6005
R1572 A3.n21 A3.n12 2.6005
R1573 A3.n1 A3.t22 1.8205
R1574 A3.n1 A3.n0 1.8205
R1575 A3.n3 A3.t18 1.8205
R1576 A3.n3 A3.n2 1.8205
R1577 A3.n5 A3.t15 1.8205
R1578 A3.n5 A3.n4 1.8205
R1579 A3.n7 A3.t23 1.8205
R1580 A3.n7 A3.n6 1.8205
R1581 A3.n12 A3.t12 1.8205
R1582 A3.n12 A3.n11 1.8205
R1583 A3.n14 A3.t21 1.8205
R1584 A3.n14 A3.n13 1.8205
R1585 A3.n16 A3.t17 1.8205
R1586 A3.n16 A3.n15 1.8205
R1587 A3.n18 A3.t13 1.8205
R1588 A3.n18 A3.n17 1.8205
R1589 A3.n43 A3.t32 1.6385
R1590 A3.n43 A3.n42 1.6385
R1591 A3.n41 A3.t33 1.6385
R1592 A3.n41 A3.n40 1.6385
R1593 A3.n38 A3.t30 1.6385
R1594 A3.n38 A3.n37 1.6385
R1595 A3.n36 A3.t31 1.6385
R1596 A3.n36 A3.n35 1.6385
R1597 A3 A3.n52 1.54844
R1598 A3.n48 A3.n47 0.884196
R1599 A3.n50 A3.n49 0.884196
R1600 A3.n29 A3.n28 0.882239
R1601 A3.n31 A3.n30 0.882239
R1602 A3.n10 A3.n9 0.657891
R1603 A3.n9 A3.n8 0.657891
R1604 A3.n21 A3.n20 0.657891
R1605 A3.n20 A3.n19 0.657891
R1606 A3.n28 A3.n27 0.657891
R1607 A3.n27 A3.n26 0.657891
R1608 A3.n32 A3.n31 0.657891
R1609 A3.n33 A3.n32 0.657891
R1610 A3.n34 A3.n33 0.657891
R1611 A3.n51 A3.n50 0.657891
R1612 A3.n52 A3.n51 0.600532
R1613 A3.n30 A3.n29 0.6005
R1614 A3.n49 A3.n48 0.6005
R1615 A3.n48 A3.n44 0.284196
R1616 A3.n49 A3.n39 0.284196
R1617 A3.n30 A3.n10 0.282239
R1618 A3.n29 A3.n21 0.282239
R1619 A3.n52 A3.n34 0.278258
R1620 TG_GATE_SWITCH_magic_1.B.n54 TG_GATE_SWITCH_magic_1.B.n53 8.64842
R1621 TG_GATE_SWITCH_magic_1.B.n10 TG_GATE_SWITCH_magic_1.B.t34 5.44589
R1622 TG_GATE_SWITCH_magic_1.B.n43 TG_GATE_SWITCH_magic_1.B.t4 5.07789
R1623 TG_GATE_SWITCH_magic_1.B.n16 TG_GATE_SWITCH_magic_1.B.n15 4.7885
R1624 TG_GATE_SWITCH_magic_1.B.n14 TG_GATE_SWITCH_magic_1.B.n13 4.7885
R1625 TG_GATE_SWITCH_magic_1.B.n10 TG_GATE_SWITCH_magic_1.B.t35 4.7885
R1626 TG_GATE_SWITCH_magic_1.B.n51 TG_GATE_SWITCH_magic_1.B.n17 4.4205
R1627 TG_GATE_SWITCH_magic_1.B.n50 TG_GATE_SWITCH_magic_1.B.n18 4.4205
R1628 TG_GATE_SWITCH_magic_1.B.n49 TG_GATE_SWITCH_magic_1.B.n19 4.4205
R1629 TG_GATE_SWITCH_magic_1.B.n48 TG_GATE_SWITCH_magic_1.B.n20 4.4205
R1630 TG_GATE_SWITCH_magic_1.B.n45 TG_GATE_SWITCH_magic_1.B.t21 4.4205
R1631 TG_GATE_SWITCH_magic_1.B.n44 TG_GATE_SWITCH_magic_1.B.t23 4.4205
R1632 TG_GATE_SWITCH_magic_1.B.n43 TG_GATE_SWITCH_magic_1.B.t9 4.4205
R1633 TG_GATE_SWITCH_magic_1.B.n9 TG_GATE_SWITCH_magic_1.B.n8 3.80789
R1634 TG_GATE_SWITCH_magic_1.B.n4 TG_GATE_SWITCH_magic_1.B.n3 3.80789
R1635 TG_GATE_SWITCH_magic_1.B.n80 TG_GATE_SWITCH_magic_1.B.n79 3.80789
R1636 TG_GATE_SWITCH_magic_1.B.n75 TG_GATE_SWITCH_magic_1.B.n74 3.80789
R1637 TG_GATE_SWITCH_magic_1.B.n70 TG_GATE_SWITCH_magic_1.B.n69 3.80789
R1638 TG_GATE_SWITCH_magic_1.B.n25 TG_GATE_SWITCH_magic_1.B.n22 3.25789
R1639 TG_GATE_SWITCH_magic_1.B.n36 TG_GATE_SWITCH_magic_1.B.n33 3.25789
R1640 TG_GATE_SWITCH_magic_1.B.n59 TG_GATE_SWITCH_magic_1.B.n56 3.25789
R1641 TG_GATE_SWITCH_magic_1.B.n87 TG_GATE_SWITCH_magic_1.B.n84 3.25789
R1642 TG_GATE_SWITCH_magic_1.B.n98 TG_GATE_SWITCH_magic_1.B.n95 3.25789
R1643 TG_GATE_SWITCH_magic_1.B.n9 TG_GATE_SWITCH_magic_1.B.n6 3.1505
R1644 TG_GATE_SWITCH_magic_1.B.n4 TG_GATE_SWITCH_magic_1.B.n1 3.1505
R1645 TG_GATE_SWITCH_magic_1.B.n80 TG_GATE_SWITCH_magic_1.B.n77 3.1505
R1646 TG_GATE_SWITCH_magic_1.B.n75 TG_GATE_SWITCH_magic_1.B.n72 3.1505
R1647 TG_GATE_SWITCH_magic_1.B.n70 TG_GATE_SWITCH_magic_1.B.n67 3.1505
R1648 TG_GATE_SWITCH_magic_1.B.n53 TG_GATE_SWITCH_magic_1.B 2.8405
R1649 TG_GATE_SWITCH_magic_1.B.n25 TG_GATE_SWITCH_magic_1.B.n24 2.6005
R1650 TG_GATE_SWITCH_magic_1.B.n28 TG_GATE_SWITCH_magic_1.B.n27 2.6005
R1651 TG_GATE_SWITCH_magic_1.B.n31 TG_GATE_SWITCH_magic_1.B.n30 2.6005
R1652 TG_GATE_SWITCH_magic_1.B.n36 TG_GATE_SWITCH_magic_1.B.n35 2.6005
R1653 TG_GATE_SWITCH_magic_1.B.n39 TG_GATE_SWITCH_magic_1.B.n38 2.6005
R1654 TG_GATE_SWITCH_magic_1.B.n42 TG_GATE_SWITCH_magic_1.B.n41 2.6005
R1655 TG_GATE_SWITCH_magic_1.B.n59 TG_GATE_SWITCH_magic_1.B.n58 2.6005
R1656 TG_GATE_SWITCH_magic_1.B.n62 TG_GATE_SWITCH_magic_1.B.n61 2.6005
R1657 TG_GATE_SWITCH_magic_1.B.n65 TG_GATE_SWITCH_magic_1.B.n64 2.6005
R1658 TG_GATE_SWITCH_magic_1.B.n90 TG_GATE_SWITCH_magic_1.B.n89 2.6005
R1659 TG_GATE_SWITCH_magic_1.B.n87 TG_GATE_SWITCH_magic_1.B.n86 2.6005
R1660 TG_GATE_SWITCH_magic_1.B.n93 TG_GATE_SWITCH_magic_1.B.n92 2.6005
R1661 TG_GATE_SWITCH_magic_1.B.n98 TG_GATE_SWITCH_magic_1.B.n97 2.6005
R1662 TG_GATE_SWITCH_magic_1.B.n101 TG_GATE_SWITCH_magic_1.B.n100 2.6005
R1663 TG_GATE_SWITCH_magic_1.B.n104 TG_GATE_SWITCH_magic_1.B.n103 2.6005
R1664 TG_GATE_SWITCH_magic_1.B TG_GATE_SWITCH_magic_1.B.n54 2.37989
R1665 TG_GATE_SWITCH_magic_1.B.n100 TG_GATE_SWITCH_magic_1.B.t42 1.8205
R1666 TG_GATE_SWITCH_magic_1.B.n100 TG_GATE_SWITCH_magic_1.B.n99 1.8205
R1667 TG_GATE_SWITCH_magic_1.B.n97 TG_GATE_SWITCH_magic_1.B.t47 1.8205
R1668 TG_GATE_SWITCH_magic_1.B.n97 TG_GATE_SWITCH_magic_1.B.n96 1.8205
R1669 TG_GATE_SWITCH_magic_1.B.n95 TG_GATE_SWITCH_magic_1.B.t55 1.8205
R1670 TG_GATE_SWITCH_magic_1.B.n95 TG_GATE_SWITCH_magic_1.B.n94 1.8205
R1671 TG_GATE_SWITCH_magic_1.B.n30 TG_GATE_SWITCH_magic_1.B.t7 1.8205
R1672 TG_GATE_SWITCH_magic_1.B.n30 TG_GATE_SWITCH_magic_1.B.n29 1.8205
R1673 TG_GATE_SWITCH_magic_1.B.n27 TG_GATE_SWITCH_magic_1.B.t10 1.8205
R1674 TG_GATE_SWITCH_magic_1.B.n27 TG_GATE_SWITCH_magic_1.B.n26 1.8205
R1675 TG_GATE_SWITCH_magic_1.B.n24 TG_GATE_SWITCH_magic_1.B.t20 1.8205
R1676 TG_GATE_SWITCH_magic_1.B.n24 TG_GATE_SWITCH_magic_1.B.n23 1.8205
R1677 TG_GATE_SWITCH_magic_1.B.n22 TG_GATE_SWITCH_magic_1.B.t18 1.8205
R1678 TG_GATE_SWITCH_magic_1.B.n22 TG_GATE_SWITCH_magic_1.B.n21 1.8205
R1679 TG_GATE_SWITCH_magic_1.B.n41 TG_GATE_SWITCH_magic_1.B.t1 1.8205
R1680 TG_GATE_SWITCH_magic_1.B.n41 TG_GATE_SWITCH_magic_1.B.n40 1.8205
R1681 TG_GATE_SWITCH_magic_1.B.n38 TG_GATE_SWITCH_magic_1.B.t3 1.8205
R1682 TG_GATE_SWITCH_magic_1.B.n38 TG_GATE_SWITCH_magic_1.B.n37 1.8205
R1683 TG_GATE_SWITCH_magic_1.B.n35 TG_GATE_SWITCH_magic_1.B.t15 1.8205
R1684 TG_GATE_SWITCH_magic_1.B.n35 TG_GATE_SWITCH_magic_1.B.n34 1.8205
R1685 TG_GATE_SWITCH_magic_1.B.n33 TG_GATE_SWITCH_magic_1.B.t11 1.8205
R1686 TG_GATE_SWITCH_magic_1.B.n33 TG_GATE_SWITCH_magic_1.B.n32 1.8205
R1687 TG_GATE_SWITCH_magic_1.B.n64 TG_GATE_SWITCH_magic_1.B.t37 1.8205
R1688 TG_GATE_SWITCH_magic_1.B.n64 TG_GATE_SWITCH_magic_1.B.n63 1.8205
R1689 TG_GATE_SWITCH_magic_1.B.n61 TG_GATE_SWITCH_magic_1.B.t46 1.8205
R1690 TG_GATE_SWITCH_magic_1.B.n61 TG_GATE_SWITCH_magic_1.B.n60 1.8205
R1691 TG_GATE_SWITCH_magic_1.B.n58 TG_GATE_SWITCH_magic_1.B.t54 1.8205
R1692 TG_GATE_SWITCH_magic_1.B.n58 TG_GATE_SWITCH_magic_1.B.n57 1.8205
R1693 TG_GATE_SWITCH_magic_1.B.n56 TG_GATE_SWITCH_magic_1.B.t36 1.8205
R1694 TG_GATE_SWITCH_magic_1.B.n56 TG_GATE_SWITCH_magic_1.B.n55 1.8205
R1695 TG_GATE_SWITCH_magic_1.B.n92 TG_GATE_SWITCH_magic_1.B.t49 1.8205
R1696 TG_GATE_SWITCH_magic_1.B.n92 TG_GATE_SWITCH_magic_1.B.n91 1.8205
R1697 TG_GATE_SWITCH_magic_1.B.n84 TG_GATE_SWITCH_magic_1.B.t48 1.8205
R1698 TG_GATE_SWITCH_magic_1.B.n84 TG_GATE_SWITCH_magic_1.B.n83 1.8205
R1699 TG_GATE_SWITCH_magic_1.B.n86 TG_GATE_SWITCH_magic_1.B.t43 1.8205
R1700 TG_GATE_SWITCH_magic_1.B.n86 TG_GATE_SWITCH_magic_1.B.n85 1.8205
R1701 TG_GATE_SWITCH_magic_1.B.n89 TG_GATE_SWITCH_magic_1.B.t38 1.8205
R1702 TG_GATE_SWITCH_magic_1.B.n89 TG_GATE_SWITCH_magic_1.B.n88 1.8205
R1703 TG_GATE_SWITCH_magic_1.B.n103 TG_GATE_SWITCH_magic_1.B.t56 1.8205
R1704 TG_GATE_SWITCH_magic_1.B.n103 TG_GATE_SWITCH_magic_1.B.n102 1.8205
R1705 TG_GATE_SWITCH_magic_1.B.n6 TG_GATE_SWITCH_magic_1.B.t33 1.6385
R1706 TG_GATE_SWITCH_magic_1.B.n6 TG_GATE_SWITCH_magic_1.B.n5 1.6385
R1707 TG_GATE_SWITCH_magic_1.B.n8 TG_GATE_SWITCH_magic_1.B.t32 1.6385
R1708 TG_GATE_SWITCH_magic_1.B.n8 TG_GATE_SWITCH_magic_1.B.n7 1.6385
R1709 TG_GATE_SWITCH_magic_1.B.n1 TG_GATE_SWITCH_magic_1.B.t31 1.6385
R1710 TG_GATE_SWITCH_magic_1.B.n1 TG_GATE_SWITCH_magic_1.B.n0 1.6385
R1711 TG_GATE_SWITCH_magic_1.B.n3 TG_GATE_SWITCH_magic_1.B.t30 1.6385
R1712 TG_GATE_SWITCH_magic_1.B.n3 TG_GATE_SWITCH_magic_1.B.n2 1.6385
R1713 TG_GATE_SWITCH_magic_1.B.n77 TG_GATE_SWITCH_magic_1.B.t60 1.6385
R1714 TG_GATE_SWITCH_magic_1.B.n77 TG_GATE_SWITCH_magic_1.B.n76 1.6385
R1715 TG_GATE_SWITCH_magic_1.B.n79 TG_GATE_SWITCH_magic_1.B.t71 1.6385
R1716 TG_GATE_SWITCH_magic_1.B.n79 TG_GATE_SWITCH_magic_1.B.n78 1.6385
R1717 TG_GATE_SWITCH_magic_1.B.n72 TG_GATE_SWITCH_magic_1.B.t64 1.6385
R1718 TG_GATE_SWITCH_magic_1.B.n72 TG_GATE_SWITCH_magic_1.B.n71 1.6385
R1719 TG_GATE_SWITCH_magic_1.B.n74 TG_GATE_SWITCH_magic_1.B.t62 1.6385
R1720 TG_GATE_SWITCH_magic_1.B.n74 TG_GATE_SWITCH_magic_1.B.n73 1.6385
R1721 TG_GATE_SWITCH_magic_1.B.n67 TG_GATE_SWITCH_magic_1.B.t68 1.6385
R1722 TG_GATE_SWITCH_magic_1.B.n67 TG_GATE_SWITCH_magic_1.B.n66 1.6385
R1723 TG_GATE_SWITCH_magic_1.B.n69 TG_GATE_SWITCH_magic_1.B.t66 1.6385
R1724 TG_GATE_SWITCH_magic_1.B.n69 TG_GATE_SWITCH_magic_1.B.n68 1.6385
R1725 TG_GATE_SWITCH_magic_1.B.n53 TG_GATE_SWITCH_magic_1.B.n52 1.32221
R1726 TG_GATE_SWITCH_magic_1.B.n11 TG_GATE_SWITCH_magic_1.B.n10 0.884196
R1727 TG_GATE_SWITCH_magic_1.B.n14 TG_GATE_SWITCH_magic_1.B.n12 0.884196
R1728 TG_GATE_SWITCH_magic_1.B.n46 TG_GATE_SWITCH_magic_1.B.n45 0.882239
R1729 TG_GATE_SWITCH_magic_1.B.n48 TG_GATE_SWITCH_magic_1.B.n47 0.882239
R1730 TG_GATE_SWITCH_magic_1.B.n52 TG_GATE_SWITCH_magic_1.B.n16 0.8105
R1731 TG_GATE_SWITCH_magic_1.B.n28 TG_GATE_SWITCH_magic_1.B.n25 0.657891
R1732 TG_GATE_SWITCH_magic_1.B.n31 TG_GATE_SWITCH_magic_1.B.n28 0.657891
R1733 TG_GATE_SWITCH_magic_1.B.n39 TG_GATE_SWITCH_magic_1.B.n36 0.657891
R1734 TG_GATE_SWITCH_magic_1.B.n42 TG_GATE_SWITCH_magic_1.B.n39 0.657891
R1735 TG_GATE_SWITCH_magic_1.B.n44 TG_GATE_SWITCH_magic_1.B.n43 0.657891
R1736 TG_GATE_SWITCH_magic_1.B.n45 TG_GATE_SWITCH_magic_1.B.n44 0.657891
R1737 TG_GATE_SWITCH_magic_1.B.n16 TG_GATE_SWITCH_magic_1.B.n14 0.657891
R1738 TG_GATE_SWITCH_magic_1.B.n51 TG_GATE_SWITCH_magic_1.B.n50 0.657891
R1739 TG_GATE_SWITCH_magic_1.B.n50 TG_GATE_SWITCH_magic_1.B.n49 0.657891
R1740 TG_GATE_SWITCH_magic_1.B.n49 TG_GATE_SWITCH_magic_1.B.n48 0.657891
R1741 TG_GATE_SWITCH_magic_1.B.n62 TG_GATE_SWITCH_magic_1.B.n59 0.657891
R1742 TG_GATE_SWITCH_magic_1.B.n65 TG_GATE_SWITCH_magic_1.B.n62 0.657891
R1743 TG_GATE_SWITCH_magic_1.B.n90 TG_GATE_SWITCH_magic_1.B.n87 0.657891
R1744 TG_GATE_SWITCH_magic_1.B.n101 TG_GATE_SWITCH_magic_1.B.n98 0.657891
R1745 TG_GATE_SWITCH_magic_1.B.n104 TG_GATE_SWITCH_magic_1.B.n101 0.657891
R1746 TG_GATE_SWITCH_magic_1.B.n93 TG_GATE_SWITCH_magic_1.B.n90 0.655976
R1747 TG_GATE_SWITCH_magic_1.B.n105 TG_GATE_SWITCH_magic_1.B.n93 0.645657
R1748 TG_GATE_SWITCH_magic_1.B.n47 TG_GATE_SWITCH_magic_1.B.n46 0.6005
R1749 TG_GATE_SWITCH_magic_1.B.n12 TG_GATE_SWITCH_magic_1.B.n11 0.6005
R1750 TG_GATE_SWITCH_magic_1.B.n81 TG_GATE_SWITCH_magic_1.B.n80 0.548416
R1751 TG_GATE_SWITCH_magic_1.B.n106 TG_GATE_SWITCH_magic_1.B.n65 0.317366
R1752 TG_GATE_SWITCH_magic_1.B.n82 TG_GATE_SWITCH_magic_1.B.n70 0.304838
R1753 TG_GATE_SWITCH_magic_1.B.n11 TG_GATE_SWITCH_magic_1.B.n9 0.284196
R1754 TG_GATE_SWITCH_magic_1.B.n12 TG_GATE_SWITCH_magic_1.B.n4 0.284196
R1755 TG_GATE_SWITCH_magic_1.B.n81 TG_GATE_SWITCH_magic_1.B.n75 0.284196
R1756 TG_GATE_SWITCH_magic_1.B.n106 TG_GATE_SWITCH_magic_1.B.n105 0.283032
R1757 TG_GATE_SWITCH_magic_1.B.n47 TG_GATE_SWITCH_magic_1.B.n31 0.282239
R1758 TG_GATE_SWITCH_magic_1.B.n46 TG_GATE_SWITCH_magic_1.B.n42 0.282239
R1759 TG_GATE_SWITCH_magic_1.B.n105 TG_GATE_SWITCH_magic_1.B.n104 0.279866
R1760 TG_GATE_SWITCH_magic_1.B.n82 TG_GATE_SWITCH_magic_1.B.n81 0.244078
R1761 TG_GATE_SWITCH_magic_1.B.n52 TG_GATE_SWITCH_magic_1.B.n51 0.237239
R1762 TG_GATE_SWITCH_magic_1.B.n107 TG_GATE_SWITCH_magic_1.B.n106 0.2009
R1763 TG_GATE_SWITCH_magic_1.B.n106 TG_GATE_SWITCH_magic_1.B.n82 0.1355
R1764 TG_GATE_SWITCH_magic_1.B TG_GATE_SWITCH_magic_1.B.n107 0.0869
R1765 TG_GATE_SWITCH_magic_0.B TG_GATE_SWITCH_magic_0.B.n105 9.68772
R1766 TG_GATE_SWITCH_magic_0.B.n99 TG_GATE_SWITCH_magic_0.B.t29 5.44589
R1767 TG_GATE_SWITCH_magic_0.B.n74 TG_GATE_SWITCH_magic_0.B.t58 5.07789
R1768 TG_GATE_SWITCH_magic_0.B.n103 TG_GATE_SWITCH_magic_0.B.n87 4.7885
R1769 TG_GATE_SWITCH_magic_0.B.n102 TG_GATE_SWITCH_magic_0.B.n88 4.7885
R1770 TG_GATE_SWITCH_magic_0.B.n99 TG_GATE_SWITCH_magic_0.B.t32 4.7885
R1771 TG_GATE_SWITCH_magic_0.B.n80 TG_GATE_SWITCH_magic_0.B.n79 4.4205
R1772 TG_GATE_SWITCH_magic_0.B.n82 TG_GATE_SWITCH_magic_0.B.n81 4.4205
R1773 TG_GATE_SWITCH_magic_0.B.n84 TG_GATE_SWITCH_magic_0.B.n83 4.4205
R1774 TG_GATE_SWITCH_magic_0.B.n86 TG_GATE_SWITCH_magic_0.B.n85 4.4205
R1775 TG_GATE_SWITCH_magic_0.B.n76 TG_GATE_SWITCH_magic_0.B.t57 4.4205
R1776 TG_GATE_SWITCH_magic_0.B.n75 TG_GATE_SWITCH_magic_0.B.t8 4.4205
R1777 TG_GATE_SWITCH_magic_0.B.n74 TG_GATE_SWITCH_magic_0.B.t0 4.4205
R1778 TG_GATE_SWITCH_magic_0.B.n27 TG_GATE_SWITCH_magic_0.B.n24 3.80789
R1779 TG_GATE_SWITCH_magic_0.B.n32 TG_GATE_SWITCH_magic_0.B.n29 3.80789
R1780 TG_GATE_SWITCH_magic_0.B.n93 TG_GATE_SWITCH_magic_0.B.n90 3.80789
R1781 TG_GATE_SWITCH_magic_0.B.n98 TG_GATE_SWITCH_magic_0.B.n95 3.80789
R1782 TG_GATE_SWITCH_magic_0.B.n37 TG_GATE_SWITCH_magic_0.B.n34 3.80789
R1783 TG_GATE_SWITCH_magic_0.B.n71 TG_GATE_SWITCH_magic_0.B.n70 3.25789
R1784 TG_GATE_SWITCH_magic_0.B.n60 TG_GATE_SWITCH_magic_0.B.n59 3.25789
R1785 TG_GATE_SWITCH_magic_0.B.n19 TG_GATE_SWITCH_magic_0.B.n18 3.25789
R1786 TG_GATE_SWITCH_magic_0.B.n8 TG_GATE_SWITCH_magic_0.B.n7 3.25789
R1787 TG_GATE_SWITCH_magic_0.B.n48 TG_GATE_SWITCH_magic_0.B.n47 3.25789
R1788 TG_GATE_SWITCH_magic_0.B.n27 TG_GATE_SWITCH_magic_0.B.n26 3.1505
R1789 TG_GATE_SWITCH_magic_0.B.n32 TG_GATE_SWITCH_magic_0.B.n31 3.1505
R1790 TG_GATE_SWITCH_magic_0.B.n93 TG_GATE_SWITCH_magic_0.B.n92 3.1505
R1791 TG_GATE_SWITCH_magic_0.B.n98 TG_GATE_SWITCH_magic_0.B.n97 3.1505
R1792 TG_GATE_SWITCH_magic_0.B.n37 TG_GATE_SWITCH_magic_0.B.n36 3.1505
R1793 TG_GATE_SWITCH_magic_0.B.n71 TG_GATE_SWITCH_magic_0.B.n68 2.6005
R1794 TG_GATE_SWITCH_magic_0.B.n72 TG_GATE_SWITCH_magic_0.B.n66 2.6005
R1795 TG_GATE_SWITCH_magic_0.B.n73 TG_GATE_SWITCH_magic_0.B.n64 2.6005
R1796 TG_GATE_SWITCH_magic_0.B.n60 TG_GATE_SWITCH_magic_0.B.n57 2.6005
R1797 TG_GATE_SWITCH_magic_0.B.n61 TG_GATE_SWITCH_magic_0.B.n55 2.6005
R1798 TG_GATE_SWITCH_magic_0.B.n62 TG_GATE_SWITCH_magic_0.B.n53 2.6005
R1799 TG_GATE_SWITCH_magic_0.B.n19 TG_GATE_SWITCH_magic_0.B.n16 2.6005
R1800 TG_GATE_SWITCH_magic_0.B.n20 TG_GATE_SWITCH_magic_0.B.n14 2.6005
R1801 TG_GATE_SWITCH_magic_0.B.n21 TG_GATE_SWITCH_magic_0.B.n12 2.6005
R1802 TG_GATE_SWITCH_magic_0.B.n8 TG_GATE_SWITCH_magic_0.B.n5 2.6005
R1803 TG_GATE_SWITCH_magic_0.B.n9 TG_GATE_SWITCH_magic_0.B.n3 2.6005
R1804 TG_GATE_SWITCH_magic_0.B.n10 TG_GATE_SWITCH_magic_0.B.n1 2.6005
R1805 TG_GATE_SWITCH_magic_0.B.n48 TG_GATE_SWITCH_magic_0.B.n45 2.6005
R1806 TG_GATE_SWITCH_magic_0.B.n49 TG_GATE_SWITCH_magic_0.B.n43 2.6005
R1807 TG_GATE_SWITCH_magic_0.B.n50 TG_GATE_SWITCH_magic_0.B.n41 2.6005
R1808 TG_GATE_SWITCH_magic_0.B.n64 TG_GATE_SWITCH_magic_0.B.t6 1.8205
R1809 TG_GATE_SWITCH_magic_0.B.n64 TG_GATE_SWITCH_magic_0.B.n63 1.8205
R1810 TG_GATE_SWITCH_magic_0.B.n66 TG_GATE_SWITCH_magic_0.B.t54 1.8205
R1811 TG_GATE_SWITCH_magic_0.B.n66 TG_GATE_SWITCH_magic_0.B.n65 1.8205
R1812 TG_GATE_SWITCH_magic_0.B.n68 TG_GATE_SWITCH_magic_0.B.t63 1.8205
R1813 TG_GATE_SWITCH_magic_0.B.n68 TG_GATE_SWITCH_magic_0.B.n67 1.8205
R1814 TG_GATE_SWITCH_magic_0.B.n70 TG_GATE_SWITCH_magic_0.B.t7 1.8205
R1815 TG_GATE_SWITCH_magic_0.B.n70 TG_GATE_SWITCH_magic_0.B.n69 1.8205
R1816 TG_GATE_SWITCH_magic_0.B.n53 TG_GATE_SWITCH_magic_0.B.t52 1.8205
R1817 TG_GATE_SWITCH_magic_0.B.n53 TG_GATE_SWITCH_magic_0.B.n52 1.8205
R1818 TG_GATE_SWITCH_magic_0.B.n55 TG_GATE_SWITCH_magic_0.B.t59 1.8205
R1819 TG_GATE_SWITCH_magic_0.B.n55 TG_GATE_SWITCH_magic_0.B.n54 1.8205
R1820 TG_GATE_SWITCH_magic_0.B.n57 TG_GATE_SWITCH_magic_0.B.t10 1.8205
R1821 TG_GATE_SWITCH_magic_0.B.n57 TG_GATE_SWITCH_magic_0.B.n56 1.8205
R1822 TG_GATE_SWITCH_magic_0.B.n59 TG_GATE_SWITCH_magic_0.B.t53 1.8205
R1823 TG_GATE_SWITCH_magic_0.B.n59 TG_GATE_SWITCH_magic_0.B.n58 1.8205
R1824 TG_GATE_SWITCH_magic_0.B.n12 TG_GATE_SWITCH_magic_0.B.t68 1.8205
R1825 TG_GATE_SWITCH_magic_0.B.n12 TG_GATE_SWITCH_magic_0.B.n11 1.8205
R1826 TG_GATE_SWITCH_magic_0.B.n14 TG_GATE_SWITCH_magic_0.B.t50 1.8205
R1827 TG_GATE_SWITCH_magic_0.B.n14 TG_GATE_SWITCH_magic_0.B.n13 1.8205
R1828 TG_GATE_SWITCH_magic_0.B.n16 TG_GATE_SWITCH_magic_0.B.t43 1.8205
R1829 TG_GATE_SWITCH_magic_0.B.n16 TG_GATE_SWITCH_magic_0.B.n15 1.8205
R1830 TG_GATE_SWITCH_magic_0.B.n18 TG_GATE_SWITCH_magic_0.B.t67 1.8205
R1831 TG_GATE_SWITCH_magic_0.B.n18 TG_GATE_SWITCH_magic_0.B.n17 1.8205
R1832 TG_GATE_SWITCH_magic_0.B.n1 TG_GATE_SWITCH_magic_0.B.t45 1.8205
R1833 TG_GATE_SWITCH_magic_0.B.n1 TG_GATE_SWITCH_magic_0.B.n0 1.8205
R1834 TG_GATE_SWITCH_magic_0.B.n3 TG_GATE_SWITCH_magic_0.B.t69 1.8205
R1835 TG_GATE_SWITCH_magic_0.B.n3 TG_GATE_SWITCH_magic_0.B.n2 1.8205
R1836 TG_GATE_SWITCH_magic_0.B.n5 TG_GATE_SWITCH_magic_0.B.t36 1.8205
R1837 TG_GATE_SWITCH_magic_0.B.n5 TG_GATE_SWITCH_magic_0.B.n4 1.8205
R1838 TG_GATE_SWITCH_magic_0.B.n7 TG_GATE_SWITCH_magic_0.B.t44 1.8205
R1839 TG_GATE_SWITCH_magic_0.B.n7 TG_GATE_SWITCH_magic_0.B.n6 1.8205
R1840 TG_GATE_SWITCH_magic_0.B.n41 TG_GATE_SWITCH_magic_0.B.t38 1.8205
R1841 TG_GATE_SWITCH_magic_0.B.n41 TG_GATE_SWITCH_magic_0.B.n40 1.8205
R1842 TG_GATE_SWITCH_magic_0.B.n43 TG_GATE_SWITCH_magic_0.B.t46 1.8205
R1843 TG_GATE_SWITCH_magic_0.B.n43 TG_GATE_SWITCH_magic_0.B.n42 1.8205
R1844 TG_GATE_SWITCH_magic_0.B.n45 TG_GATE_SWITCH_magic_0.B.t49 1.8205
R1845 TG_GATE_SWITCH_magic_0.B.n45 TG_GATE_SWITCH_magic_0.B.n44 1.8205
R1846 TG_GATE_SWITCH_magic_0.B.n47 TG_GATE_SWITCH_magic_0.B.t37 1.8205
R1847 TG_GATE_SWITCH_magic_0.B.n47 TG_GATE_SWITCH_magic_0.B.n46 1.8205
R1848 TG_GATE_SWITCH_magic_0.B.n34 TG_GATE_SWITCH_magic_0.B.t11 1.6385
R1849 TG_GATE_SWITCH_magic_0.B.n34 TG_GATE_SWITCH_magic_0.B.n33 1.6385
R1850 TG_GATE_SWITCH_magic_0.B.n26 TG_GATE_SWITCH_magic_0.B.t14 1.6385
R1851 TG_GATE_SWITCH_magic_0.B.n26 TG_GATE_SWITCH_magic_0.B.n25 1.6385
R1852 TG_GATE_SWITCH_magic_0.B.n24 TG_GATE_SWITCH_magic_0.B.t15 1.6385
R1853 TG_GATE_SWITCH_magic_0.B.n24 TG_GATE_SWITCH_magic_0.B.n23 1.6385
R1854 TG_GATE_SWITCH_magic_0.B.n31 TG_GATE_SWITCH_magic_0.B.t12 1.6385
R1855 TG_GATE_SWITCH_magic_0.B.n31 TG_GATE_SWITCH_magic_0.B.n30 1.6385
R1856 TG_GATE_SWITCH_magic_0.B.n29 TG_GATE_SWITCH_magic_0.B.t13 1.6385
R1857 TG_GATE_SWITCH_magic_0.B.n29 TG_GATE_SWITCH_magic_0.B.n28 1.6385
R1858 TG_GATE_SWITCH_magic_0.B.n92 TG_GATE_SWITCH_magic_0.B.t30 1.6385
R1859 TG_GATE_SWITCH_magic_0.B.n92 TG_GATE_SWITCH_magic_0.B.n91 1.6385
R1860 TG_GATE_SWITCH_magic_0.B.n90 TG_GATE_SWITCH_magic_0.B.t33 1.6385
R1861 TG_GATE_SWITCH_magic_0.B.n90 TG_GATE_SWITCH_magic_0.B.n89 1.6385
R1862 TG_GATE_SWITCH_magic_0.B.n97 TG_GATE_SWITCH_magic_0.B.t34 1.6385
R1863 TG_GATE_SWITCH_magic_0.B.n97 TG_GATE_SWITCH_magic_0.B.n96 1.6385
R1864 TG_GATE_SWITCH_magic_0.B.n95 TG_GATE_SWITCH_magic_0.B.t31 1.6385
R1865 TG_GATE_SWITCH_magic_0.B.n95 TG_GATE_SWITCH_magic_0.B.n94 1.6385
R1866 TG_GATE_SWITCH_magic_0.B.n36 TG_GATE_SWITCH_magic_0.B.t16 1.6385
R1867 TG_GATE_SWITCH_magic_0.B.n36 TG_GATE_SWITCH_magic_0.B.n35 1.6385
R1868 TG_GATE_SWITCH_magic_0.B.n105 TG_GATE_SWITCH_magic_0.B 1.4012
R1869 TG_GATE_SWITCH_magic_0.B.n105 TG_GATE_SWITCH_magic_0.B.n104 1.31163
R1870 TG_GATE_SWITCH_magic_0.B.n100 TG_GATE_SWITCH_magic_0.B.n99 0.884196
R1871 TG_GATE_SWITCH_magic_0.B.n102 TG_GATE_SWITCH_magic_0.B.n101 0.884196
R1872 TG_GATE_SWITCH_magic_0.B.n77 TG_GATE_SWITCH_magic_0.B.n76 0.882239
R1873 TG_GATE_SWITCH_magic_0.B.n80 TG_GATE_SWITCH_magic_0.B.n78 0.882239
R1874 TG_GATE_SWITCH_magic_0.B.n104 TG_GATE_SWITCH_magic_0.B.n103 0.8105
R1875 TG_GATE_SWITCH_magic_0.B.n76 TG_GATE_SWITCH_magic_0.B.n75 0.657891
R1876 TG_GATE_SWITCH_magic_0.B.n75 TG_GATE_SWITCH_magic_0.B.n74 0.657891
R1877 TG_GATE_SWITCH_magic_0.B.n73 TG_GATE_SWITCH_magic_0.B.n72 0.657891
R1878 TG_GATE_SWITCH_magic_0.B.n72 TG_GATE_SWITCH_magic_0.B.n71 0.657891
R1879 TG_GATE_SWITCH_magic_0.B.n62 TG_GATE_SWITCH_magic_0.B.n61 0.657891
R1880 TG_GATE_SWITCH_magic_0.B.n61 TG_GATE_SWITCH_magic_0.B.n60 0.657891
R1881 TG_GATE_SWITCH_magic_0.B.n82 TG_GATE_SWITCH_magic_0.B.n80 0.657891
R1882 TG_GATE_SWITCH_magic_0.B.n84 TG_GATE_SWITCH_magic_0.B.n82 0.657891
R1883 TG_GATE_SWITCH_magic_0.B.n86 TG_GATE_SWITCH_magic_0.B.n84 0.657891
R1884 TG_GATE_SWITCH_magic_0.B.n103 TG_GATE_SWITCH_magic_0.B.n102 0.657891
R1885 TG_GATE_SWITCH_magic_0.B.n20 TG_GATE_SWITCH_magic_0.B.n19 0.657891
R1886 TG_GATE_SWITCH_magic_0.B.n10 TG_GATE_SWITCH_magic_0.B.n9 0.657891
R1887 TG_GATE_SWITCH_magic_0.B.n9 TG_GATE_SWITCH_magic_0.B.n8 0.657891
R1888 TG_GATE_SWITCH_magic_0.B.n50 TG_GATE_SWITCH_magic_0.B.n49 0.657891
R1889 TG_GATE_SWITCH_magic_0.B.n49 TG_GATE_SWITCH_magic_0.B.n48 0.657891
R1890 TG_GATE_SWITCH_magic_0.B.n21 TG_GATE_SWITCH_magic_0.B.n20 0.655976
R1891 TG_GATE_SWITCH_magic_0.B.n22 TG_GATE_SWITCH_magic_0.B.n21 0.645657
R1892 TG_GATE_SWITCH_magic_0.B.n101 TG_GATE_SWITCH_magic_0.B.n100 0.6005
R1893 TG_GATE_SWITCH_magic_0.B.n78 TG_GATE_SWITCH_magic_0.B.n77 0.6005
R1894 TG_GATE_SWITCH_magic_0.B.n38 TG_GATE_SWITCH_magic_0.B.n32 0.548416
R1895 TG_GATE_SWITCH_magic_0.B.n51 TG_GATE_SWITCH_magic_0.B.n50 0.316429
R1896 TG_GATE_SWITCH_magic_0.B.n39 TG_GATE_SWITCH_magic_0.B.n27 0.304838
R1897 TG_GATE_SWITCH_magic_0.B.n101 TG_GATE_SWITCH_magic_0.B.n93 0.284196
R1898 TG_GATE_SWITCH_magic_0.B.n100 TG_GATE_SWITCH_magic_0.B.n98 0.284196
R1899 TG_GATE_SWITCH_magic_0.B.n38 TG_GATE_SWITCH_magic_0.B.n37 0.284196
R1900 TG_GATE_SWITCH_magic_0.B.n51 TG_GATE_SWITCH_magic_0.B.n22 0.283032
R1901 TG_GATE_SWITCH_magic_0.B.n77 TG_GATE_SWITCH_magic_0.B.n73 0.282239
R1902 TG_GATE_SWITCH_magic_0.B.n78 TG_GATE_SWITCH_magic_0.B.n62 0.282239
R1903 TG_GATE_SWITCH_magic_0.B.n22 TG_GATE_SWITCH_magic_0.B.n10 0.279866
R1904 TG_GATE_SWITCH_magic_0.B.n39 TG_GATE_SWITCH_magic_0.B.n38 0.244078
R1905 TG_GATE_SWITCH_magic_0.B TG_GATE_SWITCH_magic_0.B.n51 0.241721
R1906 TG_GATE_SWITCH_magic_0.B.n104 TG_GATE_SWITCH_magic_0.B.n86 0.237239
R1907 TG_GATE_SWITCH_magic_0.B.n51 TG_GATE_SWITCH_magic_0.B.n39 0.136437
R1908 TG_magic_0.A.n106 TG_magic_0.A.n105 5.44589
R1909 TG_magic_0.A.n155 TG_magic_0.A 5.33254
R1910 TG_magic_0.A.n144 TG_magic_0.A.n142 5.07789
R1911 TG_magic_0.A.n106 TG_magic_0.A.n104 4.7885
R1912 TG_magic_0.A.n157 TG_magic_0.A.t107 4.7885
R1913 TG_magic_0.A.n156 TG_magic_0.A.t106 4.7885
R1914 TG_magic_0.A.n154 TG_magic_0.A.t7 4.4205
R1915 TG_magic_0.A.n153 TG_magic_0.A.t79 4.4205
R1916 TG_magic_0.A.n152 TG_magic_0.A.t85 4.4205
R1917 TG_magic_0.A.n151 TG_magic_0.A.t0 4.4205
R1918 TG_magic_0.A.n148 TG_magic_0.A.n147 4.4205
R1919 TG_magic_0.A.n146 TG_magic_0.A.n145 4.4205
R1920 TG_magic_0.A.n144 TG_magic_0.A.n143 4.4205
R1921 TG_magic_0.A.n100 TG_magic_0.A.n99 3.80789
R1922 TG_magic_0.A.n95 TG_magic_0.A.n94 3.80789
R1923 TG_magic_0.A.n90 TG_magic_0.A.n89 3.80789
R1924 TG_magic_0.A.n112 TG_magic_0.A.n111 3.80789
R1925 TG_magic_0.A.n118 TG_magic_0.A.n117 3.80789
R1926 TG_magic_0.A.n49 TG_magic_0.A.n48 3.80789
R1927 TG_magic_0.A.n38 TG_magic_0.A.n37 3.80789
R1928 TG_magic_0.A.n43 TG_magic_0.A.n42 3.80789
R1929 TG_magic_0.A.n15 TG_magic_0.A.n12 3.25789
R1930 TG_magic_0.A.n4 TG_magic_0.A.n1 3.25789
R1931 TG_magic_0.A.n56 TG_magic_0.A.n53 3.25789
R1932 TG_magic_0.A.n67 TG_magic_0.A.n64 3.25789
R1933 TG_magic_0.A.n79 TG_magic_0.A.n76 3.25789
R1934 TG_magic_0.A.n135 TG_magic_0.A.n132 3.25789
R1935 TG_magic_0.A.n124 TG_magic_0.A.n121 3.25789
R1936 TG_magic_0.A.n27 TG_magic_0.A.n24 3.25789
R1937 TG_magic_0.A.n100 TG_magic_0.A.n97 3.1505
R1938 TG_magic_0.A.n95 TG_magic_0.A.n92 3.1505
R1939 TG_magic_0.A.n90 TG_magic_0.A.n87 3.1505
R1940 TG_magic_0.A.n112 TG_magic_0.A.n109 3.1505
R1941 TG_magic_0.A.n118 TG_magic_0.A.n115 3.1505
R1942 TG_magic_0.A.n49 TG_magic_0.A.n46 3.1505
R1943 TG_magic_0.A.n38 TG_magic_0.A.n35 3.1505
R1944 TG_magic_0.A.n43 TG_magic_0.A.n40 3.1505
R1945 TG_magic_0.A.n160 TG_magic_0.A.n159 3.09042
R1946 TG_magic_0.A.n15 TG_magic_0.A.n14 2.6005
R1947 TG_magic_0.A.n18 TG_magic_0.A.n17 2.6005
R1948 TG_magic_0.A.n21 TG_magic_0.A.n20 2.6005
R1949 TG_magic_0.A.n4 TG_magic_0.A.n3 2.6005
R1950 TG_magic_0.A.n7 TG_magic_0.A.n6 2.6005
R1951 TG_magic_0.A.n10 TG_magic_0.A.n9 2.6005
R1952 TG_magic_0.A.n56 TG_magic_0.A.n55 2.6005
R1953 TG_magic_0.A.n59 TG_magic_0.A.n58 2.6005
R1954 TG_magic_0.A.n62 TG_magic_0.A.n61 2.6005
R1955 TG_magic_0.A.n70 TG_magic_0.A.n69 2.6005
R1956 TG_magic_0.A.n67 TG_magic_0.A.n66 2.6005
R1957 TG_magic_0.A.n73 TG_magic_0.A.n72 2.6005
R1958 TG_magic_0.A.n79 TG_magic_0.A.n78 2.6005
R1959 TG_magic_0.A.n82 TG_magic_0.A.n81 2.6005
R1960 TG_magic_0.A.n85 TG_magic_0.A.n84 2.6005
R1961 TG_magic_0.A.n135 TG_magic_0.A.n134 2.6005
R1962 TG_magic_0.A.n138 TG_magic_0.A.n137 2.6005
R1963 TG_magic_0.A.n141 TG_magic_0.A.n140 2.6005
R1964 TG_magic_0.A.n124 TG_magic_0.A.n123 2.6005
R1965 TG_magic_0.A.n127 TG_magic_0.A.n126 2.6005
R1966 TG_magic_0.A.n130 TG_magic_0.A.n129 2.6005
R1967 TG_magic_0.A.n27 TG_magic_0.A.n26 2.6005
R1968 TG_magic_0.A.n30 TG_magic_0.A.n29 2.6005
R1969 TG_magic_0.A.n33 TG_magic_0.A.n32 2.6005
R1970 TG_magic_0.A.n113 TG_magic_0.A.n107 2.59966
R1971 TG_magic_0.A.n159 TG_magic_0.A.n158 2.2505
R1972 TG_magic_0.A.n113 TG_magic_0.A.n112 2.44216
R1973 TG_magic_0.A.n119 TG_magic_0.A.n118 2.44216
R1974 TG_magic_0.A.n20 TG_magic_0.A.t93 1.8205
R1975 TG_magic_0.A.n20 TG_magic_0.A.n19 1.8205
R1976 TG_magic_0.A.n17 TG_magic_0.A.t37 1.8205
R1977 TG_magic_0.A.n17 TG_magic_0.A.n16 1.8205
R1978 TG_magic_0.A.n14 TG_magic_0.A.t44 1.8205
R1979 TG_magic_0.A.n14 TG_magic_0.A.n13 1.8205
R1980 TG_magic_0.A.n12 TG_magic_0.A.t92 1.8205
R1981 TG_magic_0.A.n12 TG_magic_0.A.n11 1.8205
R1982 TG_magic_0.A.n9 TG_magic_0.A.t39 1.8205
R1983 TG_magic_0.A.n9 TG_magic_0.A.n8 1.8205
R1984 TG_magic_0.A.n6 TG_magic_0.A.t94 1.8205
R1985 TG_magic_0.A.n6 TG_magic_0.A.n5 1.8205
R1986 TG_magic_0.A.n3 TG_magic_0.A.t69 1.8205
R1987 TG_magic_0.A.n3 TG_magic_0.A.n2 1.8205
R1988 TG_magic_0.A.n1 TG_magic_0.A.t38 1.8205
R1989 TG_magic_0.A.n1 TG_magic_0.A.n0 1.8205
R1990 TG_magic_0.A.n61 TG_magic_0.A.t16 1.8205
R1991 TG_magic_0.A.n61 TG_magic_0.A.n60 1.8205
R1992 TG_magic_0.A.n58 TG_magic_0.A.t27 1.8205
R1993 TG_magic_0.A.n58 TG_magic_0.A.n57 1.8205
R1994 TG_magic_0.A.n55 TG_magic_0.A.t33 1.8205
R1995 TG_magic_0.A.n55 TG_magic_0.A.n54 1.8205
R1996 TG_magic_0.A.n53 TG_magic_0.A.t65 1.8205
R1997 TG_magic_0.A.n53 TG_magic_0.A.n52 1.8205
R1998 TG_magic_0.A.n72 TG_magic_0.A.t25 1.8205
R1999 TG_magic_0.A.n72 TG_magic_0.A.n71 1.8205
R2000 TG_magic_0.A.n64 TG_magic_0.A.t23 1.8205
R2001 TG_magic_0.A.n64 TG_magic_0.A.n63 1.8205
R2002 TG_magic_0.A.n66 TG_magic_0.A.t17 1.8205
R2003 TG_magic_0.A.n66 TG_magic_0.A.n65 1.8205
R2004 TG_magic_0.A.n69 TG_magic_0.A.t35 1.8205
R2005 TG_magic_0.A.n69 TG_magic_0.A.n68 1.8205
R2006 TG_magic_0.A.n84 TG_magic_0.A.t32 1.8205
R2007 TG_magic_0.A.n84 TG_magic_0.A.n83 1.8205
R2008 TG_magic_0.A.n81 TG_magic_0.A.t19 1.8205
R2009 TG_magic_0.A.n81 TG_magic_0.A.n80 1.8205
R2010 TG_magic_0.A.n78 TG_magic_0.A.t24 1.8205
R2011 TG_magic_0.A.n78 TG_magic_0.A.n77 1.8205
R2012 TG_magic_0.A.n76 TG_magic_0.A.t31 1.8205
R2013 TG_magic_0.A.n76 TG_magic_0.A.n75 1.8205
R2014 TG_magic_0.A.n140 TG_magic_0.A.t8 1.8205
R2015 TG_magic_0.A.n140 TG_magic_0.A.n139 1.8205
R2016 TG_magic_0.A.n137 TG_magic_0.A.t2 1.8205
R2017 TG_magic_0.A.n137 TG_magic_0.A.n136 1.8205
R2018 TG_magic_0.A.n134 TG_magic_0.A.t77 1.8205
R2019 TG_magic_0.A.n134 TG_magic_0.A.n133 1.8205
R2020 TG_magic_0.A.n132 TG_magic_0.A.t82 1.8205
R2021 TG_magic_0.A.n132 TG_magic_0.A.n131 1.8205
R2022 TG_magic_0.A.n129 TG_magic_0.A.t6 1.8205
R2023 TG_magic_0.A.n129 TG_magic_0.A.n128 1.8205
R2024 TG_magic_0.A.n126 TG_magic_0.A.t67 1.8205
R2025 TG_magic_0.A.n126 TG_magic_0.A.n125 1.8205
R2026 TG_magic_0.A.n123 TG_magic_0.A.t84 1.8205
R2027 TG_magic_0.A.n123 TG_magic_0.A.n122 1.8205
R2028 TG_magic_0.A.n121 TG_magic_0.A.t80 1.8205
R2029 TG_magic_0.A.n121 TG_magic_0.A.n120 1.8205
R2030 TG_magic_0.A.n32 TG_magic_0.A.t88 1.8205
R2031 TG_magic_0.A.n32 TG_magic_0.A.n31 1.8205
R2032 TG_magic_0.A.n29 TG_magic_0.A.t14 1.8205
R2033 TG_magic_0.A.n29 TG_magic_0.A.n28 1.8205
R2034 TG_magic_0.A.n26 TG_magic_0.A.t40 1.8205
R2035 TG_magic_0.A.n26 TG_magic_0.A.n25 1.8205
R2036 TG_magic_0.A.n24 TG_magic_0.A.t87 1.8205
R2037 TG_magic_0.A.n24 TG_magic_0.A.n23 1.8205
R2038 TG_magic_0.A.n40 TG_magic_0.A.t47 1.6385
R2039 TG_magic_0.A.n40 TG_magic_0.A.n39 1.6385
R2040 TG_magic_0.A.n97 TG_magic_0.A.t62 1.6385
R2041 TG_magic_0.A.n97 TG_magic_0.A.n96 1.6385
R2042 TG_magic_0.A.n99 TG_magic_0.A.t12 1.6385
R2043 TG_magic_0.A.n99 TG_magic_0.A.n98 1.6385
R2044 TG_magic_0.A.n92 TG_magic_0.A.t75 1.6385
R2045 TG_magic_0.A.n92 TG_magic_0.A.n91 1.6385
R2046 TG_magic_0.A.n94 TG_magic_0.A.t59 1.6385
R2047 TG_magic_0.A.n94 TG_magic_0.A.n93 1.6385
R2048 TG_magic_0.A.n87 TG_magic_0.A.t60 1.6385
R2049 TG_magic_0.A.n87 TG_magic_0.A.n86 1.6385
R2050 TG_magic_0.A.n89 TG_magic_0.A.t68 1.6385
R2051 TG_magic_0.A.n89 TG_magic_0.A.n88 1.6385
R2052 TG_magic_0.A.n109 TG_magic_0.A.t104 1.6385
R2053 TG_magic_0.A.n109 TG_magic_0.A.n108 1.6385
R2054 TG_magic_0.A.n111 TG_magic_0.A.t102 1.6385
R2055 TG_magic_0.A.n111 TG_magic_0.A.n110 1.6385
R2056 TG_magic_0.A.n115 TG_magic_0.A.t105 1.6385
R2057 TG_magic_0.A.n115 TG_magic_0.A.n114 1.6385
R2058 TG_magic_0.A.n117 TG_magic_0.A.t103 1.6385
R2059 TG_magic_0.A.n117 TG_magic_0.A.n116 1.6385
R2060 TG_magic_0.A.n46 TG_magic_0.A.t55 1.6385
R2061 TG_magic_0.A.n46 TG_magic_0.A.n45 1.6385
R2062 TG_magic_0.A.n48 TG_magic_0.A.t49 1.6385
R2063 TG_magic_0.A.n48 TG_magic_0.A.n47 1.6385
R2064 TG_magic_0.A.n35 TG_magic_0.A.t50 1.6385
R2065 TG_magic_0.A.n35 TG_magic_0.A.n34 1.6385
R2066 TG_magic_0.A.n37 TG_magic_0.A.t56 1.6385
R2067 TG_magic_0.A.n37 TG_magic_0.A.n36 1.6385
R2068 TG_magic_0.A.n42 TG_magic_0.A.t53 1.6385
R2069 TG_magic_0.A.n42 TG_magic_0.A.n41 1.6385
R2070 TG_magic_0.A.n149 TG_magic_0.A.n148 0.882239
R2071 TG_magic_0.A.n151 TG_magic_0.A.n150 0.882239
R2072 TG_magic_0.A.n156 TG_magic_0.A.n155 0.8105
R2073 TG_magic_0.A.n18 TG_magic_0.A.n15 0.657891
R2074 TG_magic_0.A.n7 TG_magic_0.A.n4 0.657891
R2075 TG_magic_0.A.n10 TG_magic_0.A.n7 0.657891
R2076 TG_magic_0.A.n59 TG_magic_0.A.n56 0.657891
R2077 TG_magic_0.A.n62 TG_magic_0.A.n59 0.657891
R2078 TG_magic_0.A.n70 TG_magic_0.A.n67 0.657891
R2079 TG_magic_0.A.n82 TG_magic_0.A.n79 0.657891
R2080 TG_magic_0.A.n85 TG_magic_0.A.n82 0.657891
R2081 TG_magic_0.A.n146 TG_magic_0.A.n144 0.657891
R2082 TG_magic_0.A.n148 TG_magic_0.A.n146 0.657891
R2083 TG_magic_0.A.n138 TG_magic_0.A.n135 0.657891
R2084 TG_magic_0.A.n141 TG_magic_0.A.n138 0.657891
R2085 TG_magic_0.A.n127 TG_magic_0.A.n124 0.657891
R2086 TG_magic_0.A.n130 TG_magic_0.A.n127 0.657891
R2087 TG_magic_0.A.n154 TG_magic_0.A.n153 0.657891
R2088 TG_magic_0.A.n153 TG_magic_0.A.n152 0.657891
R2089 TG_magic_0.A.n152 TG_magic_0.A.n151 0.657891
R2090 TG_magic_0.A.n157 TG_magic_0.A.n156 0.657891
R2091 TG_magic_0.A.n30 TG_magic_0.A.n27 0.657891
R2092 TG_magic_0.A.n33 TG_magic_0.A.n30 0.657891
R2093 TG_magic_0.A.n21 TG_magic_0.A.n18 0.655976
R2094 TG_magic_0.A.n73 TG_magic_0.A.n70 0.655976
R2095 TG_magic_0.A.n22 TG_magic_0.A.n21 0.646796
R2096 TG_magic_0.A.n74 TG_magic_0.A.n73 0.645657
R2097 TG_magic_0.A.n150 TG_magic_0.A.n149 0.6005
R2098 TG_magic_0.A.n101 TG_magic_0.A.n100 0.548416
R2099 TG_magic_0.A.n44 TG_magic_0.A.n38 0.548416
R2100 TG_magic_0.A.n119 TG_magic_0.A.n113 0.347488
R2101 TG_magic_0.A.n159 TG_magic_0.A.n119 0.344235
R2102 TG_magic_0.A.n103 TG_magic_0.A.n85 0.317366
R2103 TG_magic_0.A.n51 TG_magic_0.A.n33 0.317366
R2104 TG_magic_0.A.n102 TG_magic_0.A.n90 0.304838
R2105 TG_magic_0.A.n50 TG_magic_0.A.n49 0.304838
R2106 TG_magic_0.A TG_magic_0.A.n103 0.2873
R2107 TG_magic_0.A TG_magic_0.A.n51 0.2873
R2108 TG_magic_0.A.n101 TG_magic_0.A.n95 0.284196
R2109 TG_magic_0.A.n44 TG_magic_0.A.n43 0.284196
R2110 TG_magic_0.A.n103 TG_magic_0.A.n74 0.283032
R2111 TG_magic_0.A.n149 TG_magic_0.A.n141 0.282239
R2112 TG_magic_0.A.n150 TG_magic_0.A.n130 0.282239
R2113 TG_magic_0.A.n51 TG_magic_0.A.n22 0.281892
R2114 TG_magic_0.A.n22 TG_magic_0.A.n10 0.279866
R2115 TG_magic_0.A.n74 TG_magic_0.A.n62 0.279866
R2116 TG_magic_0.A.n102 TG_magic_0.A.n101 0.244078
R2117 TG_magic_0.A.n50 TG_magic_0.A.n44 0.244078
R2118 TG_magic_0.A.n155 TG_magic_0.A.n154 0.237239
R2119 TG_magic_0.A.n158 TG_magic_0.A.n157 0.235158
R2120 TG_magic_0.A.n107 TG_magic_0.A.n106 0.234977
R2121 TG_magic_0.A.n103 TG_magic_0.A.n102 0.1355
R2122 TG_magic_0.A.n51 TG_magic_0.A.n50 0.1355
R2123 TG_magic_0.A TG_magic_0.A.n160 0.0761
R2124 TG_magic_0.A.n160 TG_magic_0.A 0.0605
R2125 VSS.n418 VSS.n417 6.54809e+06
R2126 VSS.n527 VSS.n526 2.57075e+06
R2127 VSS.n363 VSS.t51 23255.7
R2128 VSS.n417 VSS.n416 22086.7
R2129 VSS.n523 VSS.n522 15657.8
R2130 VSS.n66 VSS.n65 13325.2
R2131 VSS.n526 VSS.n525 9158.59
R2132 VSS.n461 VSS.n460 6331.26
R2133 VSS.n526 VSS.n524 5599.06
R2134 VSS.n522 VSS.t122 1313.37
R2135 VSS.t49 VSS.n363 685.898
R2136 VSS.n524 VSS.n523 359.269
R2137 VSS.n416 VSS.t173 323.719
R2138 VSS.t140 VSS.t146 256.411
R2139 VSS.n462 VSS.n461 234.763
R2140 VSS.n336 VSS.n335 225.963
R2141 VSS.n419 VSS.n418 201.846
R2142 VSS.t51 VSS.n362 193.911
R2143 VSS.n364 VSS.t49 193.911
R2144 VSS.n327 VSS.t54 193.911
R2145 VSS.n341 VSS.t207 158.655
R2146 VSS.n380 VSS.t60 158.655
R2147 VSS.n403 VSS.t44 158.655
R2148 VSS.n457 VSS.t116 158.655
R2149 VSS.n534 VSS.t129 149.374
R2150 VSS.n145 VSS.n144 133.013
R2151 VSS.n460 VSS.t131 132.776
R2152 VSS.t218 VSS.t72 123.397
R2153 VSS.t75 VSS.t221 123.397
R2154 VSS.t83 VSS.t159 123.397
R2155 VSS.t156 VSS.t74 123.397
R2156 VSS.t6 VSS.t23 123.397
R2157 VSS.t39 VSS.t113 123.397
R2158 VSS.t115 VSS.t138 123.397
R2159 VSS.t184 VSS.t21 123.397
R2160 VSS.t149 VSS.t80 123.397
R2161 VSS.t88 VSS.t165 123.397
R2162 VSS.t93 VSS.t216 123.397
R2163 VSS.t226 VSS.t81 123.397
R2164 VSS.t5 VSS.n462 115.385
R2165 VSS.n454 VSS.t19 106.743
R2166 VSS.n353 VSS.t210 99.3595
R2167 VSS.n368 VSS.t64 99.3595
R2168 VSS.n391 VSS.t46 99.3595
R2169 VSS.n323 VSS.t144 99.3595
R2170 VSS.n9 VSS.t95 99.3595
R2171 VSS.n17 VSS.t97 99.3595
R2172 VSS.n1 VSS.t37 99.3595
R2173 VSS.n81 VSS.t4 99.3595
R2174 VSS.n101 VSS.t91 99.3595
R2175 VSS.n121 VSS.t71 99.3595
R2176 VSS.n336 VSS.t208 97.7569
R2177 VSS.n341 VSS.t206 97.7569
R2178 VSS.n175 VSS.t63 97.7569
R2179 VSS.n380 VSS.t59 97.7569
R2180 VSS.n403 VSS.t42 97.7569
R2181 VSS.n574 VSS.t69 97.7569
R2182 VSS.n569 VSS.t73 97.7569
R2183 VSS.n556 VSS.t101 97.7569
R2184 VSS.n551 VSS.t158 97.7569
R2185 VSS.n60 VSS.t29 97.7569
R2186 VSS.n55 VSS.t22 97.7569
R2187 VSS.n66 VSS.t10 97.7569
R2188 VSS.n45 VSS.t194 97.7569
R2189 VSS.n86 VSS.t70 97.7569
R2190 VSS.n39 VSS.t82 97.7569
R2191 VSS.n106 VSS.t84 97.7569
R2192 VSS.n33 VSS.t217 97.7569
R2193 VSS.n125 VSS.t124 97.7569
R2194 VSS.n457 VSS.t117 97.7569
R2195 VSS.n7 VSS.t219 96.1543
R2196 VSS.n15 VSS.t90 96.1543
R2197 VSS.n583 VSS.t118 96.1543
R2198 VSS.n75 VSS.t7 96.1543
R2199 VSS.n95 VSS.t166 96.1543
R2200 VSS.n115 VSS.t94 96.1543
R2201 VSS.n534 VSS.t13 92.0386
R2202 VSS.n487 VSS.t2 85.5972
R2203 VSS.n214 VSS.t142 67.3082
R2204 VSS.n567 VSS.t225 62.5005
R2205 VSS.n549 VSS.t76 62.5005
R2206 VSS.n53 VSS.t8 62.5005
R2207 VSS.n73 VSS.t15 62.5005
R2208 VSS.n93 VSS.t157 62.5005
R2209 VSS.n113 VSS.t87 62.5005
R2210 VSS.n345 VSS.t204 60.8979
R2211 VSS.n377 VSS.t61 60.8979
R2212 VSS.n400 VSS.t40 60.8979
R2213 VSS.n567 VSS.t99 60.8979
R2214 VSS.n549 VSS.t155 60.8979
R2215 VSS.n53 VSS.t30 60.8979
R2216 VSS.n73 VSS.t1 60.8979
R2217 VSS.n93 VSS.t79 60.8979
R2218 VSS.n113 VSS.t213 60.8979
R2219 VSS.n452 VSS.t137 58.9893
R2220 VSS.n416 VSS.n415 58.0362
R2221 VSS.n335 VSS.n334 58.0362
R2222 VSS.t122 VSS.n521 53.4984
R2223 VSS.n24 VSS.t26 45.2651
R2224 VSS.n527 VSS.t9 39.2298
R2225 VSS.n347 VSS.t205 36.8595
R2226 VSS.n375 VSS.t62 36.8595
R2227 VSS.n398 VSS.t41 36.8595
R2228 VSS.n317 VSS.t140 36.8595
R2229 VSS.n7 VSS.t75 36.8595
R2230 VSS.n15 VSS.t156 36.8595
R2231 VSS.n583 VSS.t39 36.8595
R2232 VSS.n75 VSS.t184 36.8595
R2233 VSS.n95 VSS.t88 36.8595
R2234 VSS.n115 VSS.t226 36.8595
R2235 VSS.n569 VSS.t218 35.2569
R2236 VSS.n551 VSS.t83 35.2569
R2237 VSS.n55 VSS.t6 35.2569
R2238 VSS.n45 VSS.t115 35.2569
R2239 VSS.n39 VSS.t149 35.2569
R2240 VSS.n33 VSS.t93 35.2569
R2241 VSS.n149 VSS.t43 20.8338
R2242 VSS.n205 VSS.t141 19.2313
R2243 VSS.n28 VSS.t16 18.7248
R2244 VSS.n528 VSS.n527 18.1064
R2245 VSS.n22 VSS.t128 18.1064
R2246 VSS.n259 VSS.t186 13.5799
R2247 VSS.n271 VSS.t24 13.5799
R2248 VSS.n56 VSS.n54 13.5707
R2249 VSS.n74 VSS.n46 13.5707
R2250 VSS.n76 VSS.n74 13.5707
R2251 VSS.n94 VSS.n40 13.5707
R2252 VSS.n96 VSS.n94 13.5707
R2253 VSS.n114 VSS.n34 13.5707
R2254 VSS.n116 VSS.n114 13.5707
R2255 VSS.n570 VSS.n568 13.5707
R2256 VSS.n568 VSS.n8 13.5707
R2257 VSS.n552 VSS.n550 13.5707
R2258 VSS.n550 VSS.n16 13.5707
R2259 VSS.n401 VSS.n399 13.5707
R2260 VSS.n348 VSS.n346 13.5707
R2261 VSS.n378 VSS.n376 13.5707
R2262 VSS.n455 VSS.n453 13.4479
R2263 VSS.n428 VSS.t120 11.2365
R2264 VSS.n237 VSS.t35 9.05343
R2265 VSS.n253 VSS.n252 7.5446
R2266 VSS.n249 VSS.n247 6.88824
R2267 VSS.n218 VSS.t31 6.88824
R2268 VSS.n468 VSS.n466 6.88824
R2269 VSS.n471 VSS.n470 6.88824
R2270 VSS.n516 VSS.t123 6.88824
R2271 VSS.n517 VSS.t161 6.88824
R2272 VSS.n146 VSS.n145 6.47389
R2273 VSS.n249 VSS.n248 6.4265
R2274 VSS.n218 VSS.t25 6.4265
R2275 VSS.n471 VSS.n469 6.4265
R2276 VSS.n468 VSS.n467 6.4265
R2277 VSS.n517 VSS.t167 6.4265
R2278 VSS.n516 VSS.t134 6.4265
R2279 VSS.n291 VSS.n290 6.05549
R2280 VSS.n37 VSS.n35 5.44589
R2281 VSS.n139 VSS.t121 5.44589
R2282 VSS.n6 VSS.n4 5.44589
R2283 VSS.n11 VSS.t96 5.44589
R2284 VSS.n19 VSS.t160 5.44589
R2285 VSS.n217 VSS.t110 5.44589
R2286 VSS.n14 VSS.n13 5.44589
R2287 VSS.n184 VSS.t200 5.44589
R2288 VSS.n185 VSS.t147 5.44589
R2289 VSS.n330 VSS.t55 5.44589
R2290 VSS.n332 VSS.t56 5.44589
R2291 VSS.n182 VSS.t212 5.44589
R2292 VSS.n183 VSS.t229 5.44589
R2293 VSS.n357 VSS.t176 5.44589
R2294 VSS.n358 VSS.t57 5.44589
R2295 VSS.n177 VSS.t67 5.44589
R2296 VSS.n178 VSS.t65 5.44589
R2297 VSS.n179 VSS.t50 5.44589
R2298 VSS.n180 VSS.t172 5.44589
R2299 VSS.n173 VSS.t233 5.44589
R2300 VSS.n174 VSS.t231 5.44589
R2301 VSS.n171 VSS.t47 5.44589
R2302 VSS.n172 VSS.t171 5.44589
R2303 VSS.n32 VSS.t214 5.44589
R2304 VSS.n38 VSS.t92 5.44589
R2305 VSS.n43 VSS.n42 5.44589
R2306 VSS.n49 VSS.n47 5.44589
R2307 VSS.n44 VSS.t195 5.44589
R2308 VSS.n3 VSS.t191 5.44589
R2309 VSS.n52 VSS.n51 5.44589
R2310 VSS.n493 VSS.t125 5.35029
R2311 VSS.n520 VSS.n31 5.23127
R2312 VSS.n27 VSS.n25 5.2198
R2313 VSS.n167 VSS.n166 5.2005
R2314 VSS.n166 VSS.n165 5.2005
R2315 VSS.n159 VSS.n158 5.2005
R2316 VSS.n158 VSS.n157 5.2005
R2317 VSS.n151 VSS.n150 5.2005
R2318 VSS.n150 VSS.n149 5.2005
R2319 VSS.n141 VSS.n140 5.2005
R2320 VSS.n160 VSS.t45 5.2005
R2321 VSS.n213 VSS.n212 5.2005
R2322 VSS.n212 VSS.n211 5.2005
R2323 VSS.n204 VSS.n203 5.2005
R2324 VSS.n203 VSS.n202 5.2005
R2325 VSS.n299 VSS.n298 5.2005
R2326 VSS.n298 VSS.n297 5.2005
R2327 VSS.n302 VSS.n301 5.2005
R2328 VSS.n301 VSS.n300 5.2005
R2329 VSS.n188 VSS.n187 5.2005
R2330 VSS.n187 VSS.n186 5.2005
R2331 VSS.n196 VSS.n195 5.2005
R2332 VSS.n195 VSS.n194 5.2005
R2333 VSS.n193 VSS.n192 5.2005
R2334 VSS.n192 VSS.t139 5.2005
R2335 VSS.n210 VSS.n209 5.2005
R2336 VSS.n209 VSS.n208 5.2005
R2337 VSS.n252 VSS.n251 5.2005
R2338 VSS.n533 VSS.n532 5.2005
R2339 VSS.n532 VSS.n531 5.2005
R2340 VSS.n283 VSS.n282 5.2005
R2341 VSS.n282 VSS.n281 5.2005
R2342 VSS.n273 VSS.n272 5.2005
R2343 VSS.n272 VSS.n271 5.2005
R2344 VSS.n236 VSS.n235 5.2005
R2345 VSS.n235 VSS.n234 5.2005
R2346 VSS.n25 VSS.n24 5.2005
R2347 VSS.n530 VSS.n529 5.2005
R2348 VSS.n529 VSS.n528 5.2005
R2349 VSS.n21 VSS.n20 5.2005
R2350 VSS.n255 VSS.n254 5.2005
R2351 VSS.n254 VSS.n253 5.2005
R2352 VSS.n264 VSS.n263 5.2005
R2353 VSS.n263 VSS.n262 5.2005
R2354 VSS.n261 VSS.n260 5.2005
R2355 VSS.n260 VSS.n259 5.2005
R2356 VSS.n279 VSS.n278 5.2005
R2357 VSS.n278 VSS.n277 5.2005
R2358 VSS.n498 VSS.n497 5.2005
R2359 VSS.n497 VSS.n496 5.2005
R2360 VSS.n31 VSS.n30 5.2005
R2361 VSS.n486 VSS.n485 5.2005
R2362 VSS.n485 VSS.n484 5.2005
R2363 VSS.n29 VSS.n28 5.2005
R2364 VSS.n492 VSS.n491 5.2005
R2365 VSS.n491 VSS.n490 5.2005
R2366 VSS.n520 VSS.n519 5.2005
R2367 VSS.n521 VSS.n520 5.2005
R2368 VSS.n510 VSS.n509 5.2005
R2369 VSS.n502 VSS.n501 5.2005
R2370 VSS.n501 VSS.n500 5.2005
R2371 VSS.n424 VSS.n423 5.2005
R2372 VSS.n423 VSS.n422 5.2005
R2373 VSS.n447 VSS.n446 5.2005
R2374 VSS.n446 VSS.n445 5.2005
R2375 VSS.n438 VSS.n437 5.2005
R2376 VSS.n437 VSS.n436 5.2005
R2377 VSS.n453 VSS.n452 5.2005
R2378 VSS.n430 VSS.n429 5.2005
R2379 VSS.n429 VSS.n428 5.2005
R2380 VSS.n31 VSS.n29 5.0005
R2381 VSS.n451 VSS.n130 4.85138
R2382 VSS.n294 VSS.t143 4.80819
R2383 VSS.n37 VSS.n36 4.7885
R2384 VSS.n139 VSS.t198 4.7885
R2385 VSS.n6 VSS.n5 4.7885
R2386 VSS.n11 VSS.t100 4.7885
R2387 VSS.n19 VSS.t148 4.7885
R2388 VSS.n217 VSS.t130 4.7885
R2389 VSS.n14 VSS.n12 4.7885
R2390 VSS.n185 VSS.t145 4.7885
R2391 VSS.n184 VSS.t199 4.7885
R2392 VSS.n330 VSS.t177 4.7885
R2393 VSS.n332 VSS.t179 4.7885
R2394 VSS.n183 VSS.t230 4.7885
R2395 VSS.n182 VSS.t211 4.7885
R2396 VSS.n358 VSS.t52 4.7885
R2397 VSS.n357 VSS.t178 4.7885
R2398 VSS.n178 VSS.t66 4.7885
R2399 VSS.n177 VSS.t68 4.7885
R2400 VSS.n180 VSS.t53 4.7885
R2401 VSS.n179 VSS.t232 4.7885
R2402 VSS.n174 VSS.t174 4.7885
R2403 VSS.n173 VSS.t175 4.7885
R2404 VSS.n172 VSS.t170 4.7885
R2405 VSS.n171 VSS.t48 4.7885
R2406 VSS.n32 VSS.t220 4.7885
R2407 VSS.n38 VSS.t106 4.7885
R2408 VSS.n43 VSS.n41 4.7885
R2409 VSS.n49 VSS.n48 4.7885
R2410 VSS.n44 VSS.t201 4.7885
R2411 VSS.n3 VSS.t38 4.7885
R2412 VSS.n52 VSS.n50 4.7885
R2413 VSS.n529 VSS.n27 4.66717
R2414 VSS.n163 VSS.n162 4.5005
R2415 VSS.n162 VSS.n161 4.5005
R2416 VSS.n143 VSS.n142 4.5005
R2417 VSS.n154 VSS.n153 4.5005
R2418 VSS.n153 VSS.n152 4.5005
R2419 VSS.n170 VSS.n169 4.5005
R2420 VSS.n169 VSS.n168 4.5005
R2421 VSS.n207 VSS.n206 4.5005
R2422 VSS.n206 VSS.n205 4.5005
R2423 VSS.n289 VSS.n288 4.5005
R2424 VSS.n296 VSS.n295 4.5005
R2425 VSS.n295 VSS.n294 4.5005
R2426 VSS.n191 VSS.n190 4.5005
R2427 VSS.n190 VSS.n189 4.5005
R2428 VSS.n199 VSS.n198 4.5005
R2429 VSS.n198 VSS.n197 4.5005
R2430 VSS.n216 VSS.n215 4.5005
R2431 VSS.n215 VSS.n214 4.5005
R2432 VSS.n276 VSS.n275 4.5005
R2433 VSS.n275 VSS.n274 4.5005
R2434 VSS.n23 VSS.n22 4.5005
R2435 VSS.n220 VSS.n27 4.5005
R2436 VSS.n27 VSS.n26 4.5005
R2437 VSS.n239 VSS.n238 4.5005
R2438 VSS.n238 VSS.n237 4.5005
R2439 VSS.n258 VSS.n257 4.5005
R2440 VSS.n257 VSS.n256 4.5005
R2441 VSS.n268 VSS.n267 4.5005
R2442 VSS.n267 VSS.n266 4.5005
R2443 VSS.n286 VSS.n285 4.5005
R2444 VSS.n285 VSS.n284 4.5005
R2445 VSS.n505 VSS.n504 4.5005
R2446 VSS.n504 VSS.n503 4.5005
R2447 VSS.n495 VSS.n494 4.5005
R2448 VSS.n494 VSS.n493 4.5005
R2449 VSS.n489 VSS.n488 4.5005
R2450 VSS.n488 VSS.n487 4.5005
R2451 VSS.n513 VSS.n512 4.5005
R2452 VSS.n512 VSS.n511 4.5005
R2453 VSS.n440 VSS.n439 4.5005
R2454 VSS.n435 VSS.n434 4.5005
R2455 VSS.n434 VSS.n433 4.5005
R2456 VSS.n130 VSS.n129 4.5005
R2457 VSS.n136 VSS.n135 4.5005
R2458 VSS.n421 VSS.n420 4.5005
R2459 VSS.n420 VSS.n419 4.5005
R2460 VSS.n246 VSS.n243 3.61224
R2461 VSS.n476 VSS.n473 3.61224
R2462 VSS.n481 VSS.n480 3.61224
R2463 VSS.n245 VSS.t36 3.2765
R2464 VSS.n245 VSS.n244 3.2765
R2465 VSS.n243 VSS.t185 3.2765
R2466 VSS.n243 VSS.n242 3.2765
R2467 VSS.n478 VSS.t183 3.2765
R2468 VSS.n478 VSS.n477 3.2765
R2469 VSS.n480 VSS.t180 3.2765
R2470 VSS.n480 VSS.n479 3.2765
R2471 VSS.n475 VSS.t3 3.2765
R2472 VSS.n475 VSS.n474 3.2765
R2473 VSS.n473 VSS.t14 3.2765
R2474 VSS.n473 VSS.n472 3.2765
R2475 VSS.n246 VSS.n245 3.1505
R2476 VSS.n476 VSS.n475 3.1505
R2477 VSS.n481 VSS.n478 3.1505
R2478 VSS.n25 VSS.n23 3.00927
R2479 VSS.n64 VSS 2.94101
R2480 VSS.n340 VSS.n339 2.6005
R2481 VSS.n339 VSS.t209 2.6005
R2482 VSS.n343 VSS.n342 2.6005
R2483 VSS.n342 VSS.n341 2.6005
R2484 VSS.n346 VSS.n344 2.6005
R2485 VSS.n346 VSS.n345 2.6005
R2486 VSS.n349 VSS.n348 2.6005
R2487 VSS.n348 VSS.n347 2.6005
R2488 VSS.n352 VSS.n351 2.6005
R2489 VSS.n351 VSS.n350 2.6005
R2490 VSS.n355 VSS.n354 2.6005
R2491 VSS.n354 VSS.n353 2.6005
R2492 VSS.n361 VSS.n360 2.6005
R2493 VSS.n362 VSS.n361 2.6005
R2494 VSS.n338 VSS.n337 2.6005
R2495 VSS.n337 VSS.n336 2.6005
R2496 VSS.n385 VSS.n176 2.6005
R2497 VSS.n176 VSS.n175 2.6005
R2498 VSS.n384 VSS.n383 2.6005
R2499 VSS.n383 VSS.t58 2.6005
R2500 VSS.n382 VSS.n381 2.6005
R2501 VSS.n381 VSS.n380 2.6005
R2502 VSS.n379 VSS.n378 2.6005
R2503 VSS.n378 VSS.n377 2.6005
R2504 VSS.n376 VSS.n374 2.6005
R2505 VSS.n376 VSS.n375 2.6005
R2506 VSS.n373 VSS.n372 2.6005
R2507 VSS.n372 VSS.n371 2.6005
R2508 VSS.n370 VSS.n369 2.6005
R2509 VSS.n369 VSS.n368 2.6005
R2510 VSS.n366 VSS.n365 2.6005
R2511 VSS.n365 VSS.n364 2.6005
R2512 VSS.n405 VSS.n404 2.6005
R2513 VSS.n404 VSS.n403 2.6005
R2514 VSS.n402 VSS.n401 2.6005
R2515 VSS.n401 VSS.n400 2.6005
R2516 VSS.n399 VSS.n397 2.6005
R2517 VSS.n399 VSS.n398 2.6005
R2518 VSS.n396 VSS.n395 2.6005
R2519 VSS.n395 VSS.n394 2.6005
R2520 VSS.n393 VSS.n392 2.6005
R2521 VSS.n392 VSS.n391 2.6005
R2522 VSS.n389 VSS.n388 2.6005
R2523 VSS.n388 VSS.n387 2.6005
R2524 VSS.n329 VSS.n328 2.6005
R2525 VSS.n328 VSS.n327 2.6005
R2526 VSS.n325 VSS.n324 2.6005
R2527 VSS.n324 VSS.n323 2.6005
R2528 VSS.n322 VSS.n321 2.6005
R2529 VSS.n321 VSS.n320 2.6005
R2530 VSS.n319 VSS.n318 2.6005
R2531 VSS.n318 VSS.n317 2.6005
R2532 VSS.n316 VSS.n315 2.6005
R2533 VSS.n315 VSS.n314 2.6005
R2534 VSS.n541 VSS.n540 2.6005
R2535 VSS.n540 VSS.n539 2.6005
R2536 VSS.n538 VSS.n537 2.6005
R2537 VSS.n537 VSS.t114 2.6005
R2538 VSS.n536 VSS.n535 2.6005
R2539 VSS.n535 VSS.n534 2.6005
R2540 VSS.n543 VSS.n18 2.6005
R2541 VSS.n18 VSS.n17 2.6005
R2542 VSS.n555 VSS.n554 2.6005
R2543 VSS.n554 VSS.t152 2.6005
R2544 VSS.n553 VSS.n552 2.6005
R2545 VSS.n552 VSS.n551 2.6005
R2546 VSS.n550 VSS.n548 2.6005
R2547 VSS.n550 VSS.n549 2.6005
R2548 VSS.n547 VSS.n16 2.6005
R2549 VSS.n16 VSS.n15 2.6005
R2550 VSS.n546 VSS.n545 2.6005
R2551 VSS.n545 VSS.n544 2.6005
R2552 VSS.n558 VSS.n557 2.6005
R2553 VSS.n557 VSS.n556 2.6005
R2554 VSS.n561 VSS.n10 2.6005
R2555 VSS.n10 VSS.n9 2.6005
R2556 VSS.n573 VSS.n572 2.6005
R2557 VSS.n572 VSS.t98 2.6005
R2558 VSS.n571 VSS.n570 2.6005
R2559 VSS.n570 VSS.n569 2.6005
R2560 VSS.n568 VSS.n566 2.6005
R2561 VSS.n568 VSS.n567 2.6005
R2562 VSS.n565 VSS.n8 2.6005
R2563 VSS.n8 VSS.n7 2.6005
R2564 VSS.n564 VSS.n563 2.6005
R2565 VSS.n563 VSS.n562 2.6005
R2566 VSS.n576 VSS.n575 2.6005
R2567 VSS.n575 VSS.n574 2.6005
R2568 VSS.n426 VSS.n138 2.6005
R2569 VSS.n138 VSS.n137 2.6005
R2570 VSS.n108 VSS.n107 2.6005
R2571 VSS.n107 VSS.n106 2.6005
R2572 VSS.n110 VSS.n109 2.6005
R2573 VSS.n109 VSS.t215 2.6005
R2574 VSS.n111 VSS.n34 2.6005
R2575 VSS.n34 VSS.n33 2.6005
R2576 VSS.n114 VSS.n112 2.6005
R2577 VSS.n114 VSS.n113 2.6005
R2578 VSS.n117 VSS.n116 2.6005
R2579 VSS.n116 VSS.n115 2.6005
R2580 VSS.n120 VSS.n119 2.6005
R2581 VSS.n119 VSS.n118 2.6005
R2582 VSS.n123 VSS.n122 2.6005
R2583 VSS.n122 VSS.n121 2.6005
R2584 VSS.n127 VSS.n126 2.6005
R2585 VSS.n126 VSS.n125 2.6005
R2586 VSS.n464 VSS.n463 2.6005
R2587 VSS.n463 VSS.t5 2.6005
R2588 VSS.n459 VSS.n458 2.6005
R2589 VSS.n458 VSS.n457 2.6005
R2590 VSS.n456 VSS.n455 2.6005
R2591 VSS.n455 VSS.n454 2.6005
R2592 VSS.n451 VSS.n128 2.6005
R2593 VSS.n451 VSS.n450 2.6005
R2594 VSS.n443 VSS.n442 2.6005
R2595 VSS.n442 VSS.n441 2.6005
R2596 VSS.n88 VSS.n87 2.6005
R2597 VSS.n87 VSS.n86 2.6005
R2598 VSS.n90 VSS.n89 2.6005
R2599 VSS.n89 VSS.t78 2.6005
R2600 VSS.n91 VSS.n40 2.6005
R2601 VSS.n40 VSS.n39 2.6005
R2602 VSS.n94 VSS.n92 2.6005
R2603 VSS.n94 VSS.n93 2.6005
R2604 VSS.n97 VSS.n96 2.6005
R2605 VSS.n96 VSS.n95 2.6005
R2606 VSS.n100 VSS.n99 2.6005
R2607 VSS.n99 VSS.n98 2.6005
R2608 VSS.n103 VSS.n102 2.6005
R2609 VSS.n102 VSS.n101 2.6005
R2610 VSS.n68 VSS.n67 2.6005
R2611 VSS.n67 VSS.n66 2.6005
R2612 VSS.n70 VSS.n69 2.6005
R2613 VSS.n69 VSS.t0 2.6005
R2614 VSS.n71 VSS.n46 2.6005
R2615 VSS.n46 VSS.n45 2.6005
R2616 VSS.n74 VSS.n72 2.6005
R2617 VSS.n74 VSS.n73 2.6005
R2618 VSS.n77 VSS.n76 2.6005
R2619 VSS.n76 VSS.n75 2.6005
R2620 VSS.n80 VSS.n79 2.6005
R2621 VSS.n79 VSS.n78 2.6005
R2622 VSS.n83 VSS.n82 2.6005
R2623 VSS.n82 VSS.n81 2.6005
R2624 VSS.n579 VSS.n2 2.6005
R2625 VSS.n2 VSS.n1 2.6005
R2626 VSS.n59 VSS.n58 2.6005
R2627 VSS.n58 VSS.t32 2.6005
R2628 VSS.n57 VSS.n56 2.6005
R2629 VSS.n56 VSS.n55 2.6005
R2630 VSS.n54 VSS.n0 2.6005
R2631 VSS.n54 VSS.n53 2.6005
R2632 VSS.n585 VSS.n584 2.6005
R2633 VSS.n584 VSS.n583 2.6005
R2634 VSS.n582 VSS.n581 2.6005
R2635 VSS.n581 VSS.n580 2.6005
R2636 VSS.n62 VSS.n61 2.6005
R2637 VSS.n61 VSS.n60 2.6005
R2638 VSS.n506 VSS.n465 2.5504
R2639 VSS.n303 VSS.n291 2.02106
R2640 VSS.n147 VSS.n146 1.83012
R2641 VSS.n513 VSS.n508 1.60615
R2642 VSS.n562 VSS.t224 1.60306
R2643 VSS.n544 VSS.t77 1.60306
R2644 VSS.n580 VSS.t20 1.60306
R2645 VSS.n78 VSS.t119 1.60306
R2646 VSS.n98 VSS.t164 1.60306
R2647 VSS.n118 VSS.t89 1.60306
R2648 VSS.n271 VSS.t109 1.50932
R2649 VSS.n304 VSS.n303 1.5005
R2650 VSS.n512 VSS.n510 1.30819
R2651 VSS.n448 VSS.n134 1.18011
R2652 VSS.n313 VSS.n312 1.17928
R2653 VSS.n421 VSS.n414 1.13085
R2654 VSS.n506 VSS.n505 1.12905
R2655 VSS.n146 VSS.n143 1.09698
R2656 VSS.n230 VSS.n229 0.954617
R2657 VSS.n407 VSS.n406 0.950603
R2658 VSS.n287 VSS.n286 0.906347
R2659 VSS.n291 VSS.n289 0.738188
R2660 VSS.n23 VSS.n21 0.675939
R2661 VSS.n331 VSS.n330 0.520309
R2662 VSS.n333 VSS.n332 0.506013
R2663 VSS.n162 VSS.n160 0.491728
R2664 VSS.n105 VSS.n37 0.468109
R2665 VSS.n425 VSS.n139 0.468109
R2666 VSS.n577 VSS.n6 0.468109
R2667 VSS.n560 VSS.n11 0.468109
R2668 VSS.n542 VSS.n19 0.468109
R2669 VSS.n280 VSS.n217 0.468109
R2670 VSS.n559 VSS.n14 0.468109
R2671 VSS.n326 VSS.n184 0.468109
R2672 VSS.n326 VSS.n185 0.468109
R2673 VSS.n356 VSS.n182 0.468109
R2674 VSS.n356 VSS.n183 0.468109
R2675 VSS.n359 VSS.n357 0.468109
R2676 VSS.n359 VSS.n358 0.468109
R2677 VSS.n367 VSS.n177 0.468109
R2678 VSS.n367 VSS.n178 0.468109
R2679 VSS.n181 VSS.n179 0.468109
R2680 VSS.n181 VSS.n180 0.468109
R2681 VSS.n386 VSS.n173 0.468109
R2682 VSS.n390 VSS.n171 0.468109
R2683 VSS.n390 VSS.n172 0.468109
R2684 VSS.n124 VSS.n32 0.468109
R2685 VSS.n104 VSS.n38 0.468109
R2686 VSS.n85 VSS.n43 0.468109
R2687 VSS.n64 VSS.n49 0.468109
R2688 VSS.n84 VSS.n44 0.468109
R2689 VSS.n578 VSS.n3 0.468109
R2690 VSS.n63 VSS.n52 0.468109
R2691 VSS.n250 VSS.n249 0.462042
R2692 VSS.n386 VSS.n174 0.460283
R2693 VSS.n138 VSS.n136 0.430325
R2694 VSS.n143 VSS.n141 0.430325
R2695 VSS.n414 VSS.n411 0.392577
R2696 VSS.n304 VSS.n287 0.371885
R2697 VSS.n442 VSS.n440 0.368921
R2698 VSS.n219 VSS.n218 0.368157
R2699 VSS.n265 VSS.n219 0.36433
R2700 VSS.n386 VSS.n385 0.340076
R2701 VSS.n338 VSS.n333 0.277362
R2702 VSS.n85 VSS.n84 0.261967
R2703 VSS.n578 VSS.n577 0.261178
R2704 VSS.n250 VSS.n246 0.254848
R2705 VSS.n499 VSS.n468 0.254848
R2706 VSS.n499 VSS.n471 0.254848
R2707 VSS.n483 VSS.n476 0.254848
R2708 VSS.n483 VSS.n481 0.254848
R2709 VSS.n518 VSS.n516 0.254848
R2710 VSS.n518 VSS.n517 0.254848
R2711 VSS.n560 VSS.n559 0.233875
R2712 VSS.n105 VSS.n104 0.232588
R2713 VSS.n542 VSS.n541 0.215672
R2714 VSS.n127 VSS.n124 0.215672
R2715 VSS.n453 VSS.n451 0.123307
R2716 VSS.n576 VSS.n573 0.11481
R2717 VSS.n573 VSS.n571 0.11481
R2718 VSS.n565 VSS.n564 0.11481
R2719 VSS.n564 VSS.n561 0.11481
R2720 VSS.n558 VSS.n555 0.11481
R2721 VSS.n555 VSS.n553 0.11481
R2722 VSS.n547 VSS.n546 0.11481
R2723 VSS.n546 VSS.n543 0.11481
R2724 VSS.n541 VSS.n538 0.11481
R2725 VSS.n538 VSS.n536 0.11481
R2726 VSS.n322 VSS.n319 0.11481
R2727 VSS.n325 VSS.n322 0.11481
R2728 VSS.n340 VSS.n338 0.11481
R2729 VSS.n343 VSS.n340 0.11481
R2730 VSS.n344 VSS.n343 0.11481
R2731 VSS.n352 VSS.n349 0.11481
R2732 VSS.n355 VSS.n352 0.11481
R2733 VSS.n385 VSS.n384 0.11481
R2734 VSS.n384 VSS.n382 0.11481
R2735 VSS.n382 VSS.n379 0.11481
R2736 VSS.n374 VSS.n373 0.11481
R2737 VSS.n373 VSS.n370 0.11481
R2738 VSS.n405 VSS.n402 0.11481
R2739 VSS.n397 VSS.n396 0.11481
R2740 VSS.n396 VSS.n393 0.11481
R2741 VSS.n110 VSS.n108 0.11481
R2742 VSS.n111 VSS.n110 0.11481
R2743 VSS.n120 VSS.n117 0.11481
R2744 VSS.n123 VSS.n120 0.11481
R2745 VSS.n464 VSS.n459 0.11481
R2746 VSS.n459 VSS.n456 0.11481
R2747 VSS.n90 VSS.n88 0.11481
R2748 VSS.n91 VSS.n90 0.11481
R2749 VSS.n100 VSS.n97 0.11481
R2750 VSS.n103 VSS.n100 0.11481
R2751 VSS.n70 VSS.n68 0.11481
R2752 VSS.n71 VSS.n70 0.11481
R2753 VSS.n80 VSS.n77 0.11481
R2754 VSS.n83 VSS.n80 0.11481
R2755 VSS.n62 VSS.n59 0.11481
R2756 VSS.n59 VSS.n57 0.11481
R2757 VSS.n585 VSS.n582 0.11481
R2758 VSS.n582 VSS.n579 0.11481
R2759 VSS.n536 VSS.n533 0.112741
R2760 VSS.n507 VSS.n506 0.111264
R2761 VSS VSS.n565 0.11119
R2762 VSS VSS.n547 0.11119
R2763 VSS.n319 VSS 0.11119
R2764 VSS.n349 VSS 0.11119
R2765 VSS.n374 VSS 0.11119
R2766 VSS.n397 VSS 0.11119
R2767 VSS.n117 VSS 0.11119
R2768 VSS.n97 VSS 0.11119
R2769 VSS.n77 VSS 0.11119
R2770 VSS VSS.n585 0.11119
R2771 VSS.n571 VSS 0.110672
R2772 VSS.n553 VSS 0.110672
R2773 VSS VSS.n111 0.110672
R2774 VSS VSS.n91 0.110672
R2775 VSS VSS.n71 0.110672
R2776 VSS.n57 VSS 0.110672
R2777 VSS.n131 VSS 0.110155
R2778 VSS.n329 VSS.n326 0.1055
R2779 VSS.n360 VSS.n356 0.1055
R2780 VSS.n367 VSS.n366 0.1055
R2781 VSS.n390 VSS.n389 0.1055
R2782 VSS.n465 VSS.n464 0.1055
R2783 VSS.n360 VSS.n359 0.104466
R2784 VSS.n366 VSS.n181 0.104466
R2785 VSS.n389 VSS.n386 0.102827
R2786 VSS.n508 VSS.n507 0.102239
R2787 VSS VSS.n63 0.0905
R2788 VSS.n331 VSS.n329 0.0899828
R2789 VSS VSS.n219 0.0833777
R2790 VSS.n316 VSS.n313 0.0825347
R2791 VSS.n406 VSS.n405 0.0654462
R2792 VSS.n519 VSS.n518 0.062569
R2793 VSS.n413 VSS.n412 0.0557273
R2794 VSS.n408 VSS.n407 0.0552159
R2795 VSS.n414 VSS.n413 0.0547659
R2796 VSS.n226 VSS.n225 0.0538898
R2797 VSS.n222 VSS.n221 0.0538898
R2798 VSS.n305 VSS.n304 0.0538898
R2799 VSS.n309 VSS.n308 0.0538898
R2800 VSS.n229 VSS.n228 0.0447373
R2801 VSS.n225 VSS.n224 0.0447373
R2802 VSS.n308 VSS.n307 0.0447373
R2803 VSS.n312 VSS.n311 0.0447373
R2804 VSS.n498 VSS.n495 0.044569
R2805 VSS.n411 VSS.n410 0.0439659
R2806 VSS.n134 VSS.n133 0.0434545
R2807 VSS.n489 VSS.n486 0.0427069
R2808 VSS.n519 VSS.n515 0.0427069
R2809 VSS.n450 VSS.n449 0.0413621
R2810 VSS.n495 VSS.n492 0.0408448
R2811 VSS.n492 VSS.n489 0.0408448
R2812 VSS.n515 VSS.n514 0.0408448
R2813 VSS.n514 VSS.n513 0.0402241
R2814 VSS.n220 VSS 0.0361897
R2815 VSS.n448 VSS.n447 0.0352265
R2816 VSS.n231 VSS.n230 0.0350052
R2817 VSS.n255 VSS.n241 0.0299828
R2818 VSS.n273 VSS.n270 0.0299828
R2819 VSS.n204 VSS.n201 0.0299828
R2820 VSS.n159 VSS.n156 0.0299828
R2821 VSS.n431 VSS.n430 0.0299828
R2822 VSS.n486 VSS.n483 0.0278103
R2823 VSS.n505 VSS.n502 0.0271897
R2824 VSS.n216 VSS.n213 0.0268793
R2825 VSS.n447 VSS.n444 0.0268793
R2826 VSS.n430 VSS.n427 0.0268793
R2827 VSS.n299 VSS.n296 0.0263621
R2828 VSS.n199 VSS.n196 0.0263621
R2829 VSS.n163 VSS.n159 0.0263621
R2830 VSS.n232 VSS.n231 0.0258448
R2831 VSS.n210 VSS.n207 0.0258448
R2832 VSS.n443 VSS.n438 0.0258448
R2833 VSS.n258 VSS.n255 0.0253276
R2834 VSS.n276 VSS.n273 0.0253276
R2835 VSS.n193 VSS.n191 0.0253276
R2836 VSS.n151 VSS.n148 0.0253276
R2837 VSS.n303 VSS.n302 0.0248103
R2838 VSS.n167 VSS.n164 0.0248103
R2839 VSS.n236 VSS.n233 0.0232586
R2840 VSS.n264 VSS.n261 0.0227414
R2841 VSS.n286 VSS.n283 0.017569
R2842 VSS.n239 VSS.n236 0.0170517
R2843 VSS.n265 VSS.n264 0.0165345
R2844 VSS.n191 VSS.n188 0.0160172
R2845 VSS.n207 VSS.n204 0.0160172
R2846 VSS.n154 VSS.n151 0.0160172
R2847 VSS.n170 VSS.n167 0.0160172
R2848 VSS.n425 VSS.n424 0.0160172
R2849 VSS.n424 VSS.n421 0.0160172
R2850 VSS.n438 VSS.n435 0.0155
R2851 VSS.n435 VSS.n432 0.0139483
R2852 VSS.n133 VSS.n132 0.0137955
R2853 VSS.n155 VSS.n154 0.013431
R2854 VSS.n410 VSS.n409 0.0132841
R2855 VSS.n283 VSS.n280 0.0129138
R2856 VSS.n449 VSS.n448 0.0127046
R2857 VSS.n240 VSS.n239 0.0123966
R2858 VSS.n269 VSS.n268 0.0123966
R2859 VSS.n293 VSS.n292 0.0123966
R2860 VSS.n201 VSS.n200 0.0123966
R2861 VSS.n228 VSS.n227 0.0121949
R2862 VSS.n224 VSS.n223 0.0121949
R2863 VSS.n307 VSS.n306 0.0121949
R2864 VSS.n311 VSS.n310 0.0121949
R2865 VSS.n406 VSS.n170 0.0120024
R2866 VSS.n230 VSS.n220 0.011929
R2867 VSS.n577 VSS.n576 0.0103276
R2868 VSS.n559 VSS.n558 0.0103276
R2869 VSS.n108 VSS.n105 0.0103276
R2870 VSS.n88 VSS.n85 0.0103276
R2871 VSS.n68 VSS.n64 0.0103276
R2872 VSS.n63 VSS.n62 0.0103276
R2873 VSS.n561 VSS.n560 0.00981034
R2874 VSS.n543 VSS.n542 0.00981034
R2875 VSS.n280 VSS.n279 0.00981034
R2876 VSS.n326 VSS.n325 0.00981034
R2877 VSS.n356 VSS.n355 0.00981034
R2878 VSS.n370 VSS.n367 0.00981034
R2879 VSS.n393 VSS.n390 0.00981034
R2880 VSS.n124 VSS.n123 0.00981034
R2881 VSS.n465 VSS.n127 0.00981034
R2882 VSS.n426 VSS.n425 0.00981034
R2883 VSS.n104 VSS.n103 0.00981034
R2884 VSS.n84 VSS.n83 0.00981034
R2885 VSS.n579 VSS.n578 0.00981034
R2886 VSS.n251 VSS 0.0076223
R2887 VSS.n482 VSS 0.00732759
R2888 VSS.n279 VSS.n276 0.00722414
R2889 VSS.n261 VSS.n258 0.0067069
R2890 VSS.n313 VSS.n216 0.00626092
R2891 VSS.n233 VSS.n232 0.00618966
R2892 VSS.n333 VSS.n331 0.0053
R2893 VSS.n499 VSS.n498 0.00484483
R2894 VSS.n566 VSS 0.00463793
R2895 VSS.n548 VSS 0.00463793
R2896 VSS.n302 VSS.n299 0.00463793
R2897 VSS.n164 VSS.n163 0.00463793
R2898 VSS.n112 VSS 0.00463793
R2899 VSS.n92 VSS 0.00463793
R2900 VSS.n72 VSS 0.00463793
R2901 VSS VSS.n0 0.00463793
R2902 VSS.n251 VSS.n250 0.00438489
R2903 VSS.n483 VSS.n482 0.00422414
R2904 VSS.n513 VSS 0.00422414
R2905 VSS.n566 VSS 0.00412069
R2906 VSS.n548 VSS 0.00412069
R2907 VSS.n530 VSS 0.00412069
R2908 VSS.n196 VSS.n193 0.00412069
R2909 VSS VSS.n316 0.00412069
R2910 VSS.n344 VSS 0.00412069
R2911 VSS.n379 VSS 0.00412069
R2912 VSS.n148 VSS.n147 0.00412069
R2913 VSS.n402 VSS 0.00412069
R2914 VSS.n112 VSS 0.00412069
R2915 VSS.n456 VSS 0.00412069
R2916 VSS.n427 VSS.n426 0.00412069
R2917 VSS.n92 VSS 0.00412069
R2918 VSS.n72 VSS 0.00412069
R2919 VSS VSS.n0 0.00412069
R2920 VSS.n213 VSS.n210 0.00360345
R2921 VSS.n444 VSS.n443 0.00360345
R2922 VSS.n241 VSS.n240 0.00308621
R2923 VSS.n270 VSS.n269 0.00308621
R2924 VSS.n296 VSS.n293 0.00308621
R2925 VSS.n200 VSS.n199 0.00308621
R2926 VSS.n227 VSS.n226 0.00304237
R2927 VSS.n223 VSS.n222 0.00304237
R2928 VSS.n306 VSS.n305 0.00304237
R2929 VSS.n310 VSS.n309 0.00304237
R2930 VSS.n533 VSS.n530 0.00256897
R2931 VSS.n502 VSS.n499 0.00236207
R2932 VSS.n156 VSS.n155 0.00205172
R2933 VSS.n409 VSS.n408 0.00203409
R2934 VSS.n450 VSS.n131 0.00153448
R2935 VSS.n432 VSS.n431 0.00153448
R2936 VSS.n268 VSS.n265 0.00101724
R2937 INVERTER_MUX_1.OUT.n0 INVERTER_MUX_1.OUT.t33 68.1773
R2938 INVERTER_MUX_1.OUT.n11 INVERTER_MUX_1.OUT.n10 52.5344
R2939 INVERTER_MUX_1.OUT.n12 INVERTER_MUX_1.OUT.t25 47.0594
R2940 INVERTER_MUX_1.OUT.t31 INVERTER_MUX_1.OUT.t23 43.8005
R2941 INVERTER_MUX_1.OUT.t29 INVERTER_MUX_1.OUT.t31 43.8005
R2942 INVERTER_MUX_1.OUT.t25 INVERTER_MUX_1.OUT.t29 43.8005
R2943 INVERTER_MUX_1.OUT.t27 INVERTER_MUX_1.OUT.n4 33.763
R2944 INVERTER_MUX_1.OUT.n9 INVERTER_MUX_1.OUT.t20 21.9005
R2945 INVERTER_MUX_1.OUT.n9 INVERTER_MUX_1.OUT.t30 21.9005
R2946 INVERTER_MUX_1.OUT.n8 INVERTER_MUX_1.OUT.t16 21.9005
R2947 INVERTER_MUX_1.OUT.n8 INVERTER_MUX_1.OUT.t24 21.9005
R2948 INVERTER_MUX_1.OUT.n7 INVERTER_MUX_1.OUT.t32 21.9005
R2949 INVERTER_MUX_1.OUT.n7 INVERTER_MUX_1.OUT.t21 21.9005
R2950 INVERTER_MUX_1.OUT.n6 INVERTER_MUX_1.OUT.t28 21.9005
R2951 INVERTER_MUX_1.OUT.n6 INVERTER_MUX_1.OUT.t19 21.9005
R2952 INVERTER_MUX_1.OUT.n5 INVERTER_MUX_1.OUT.t18 21.9005
R2953 INVERTER_MUX_1.OUT.n5 INVERTER_MUX_1.OUT.t27 21.9005
R2954 INVERTER_MUX_1.OUT.n4 INVERTER_MUX_1.OUT.n3 20.8576
R2955 INVERTER_MUX_1.OUT.n3 INVERTER_MUX_1.OUT.n2 20.8576
R2956 INVERTER_MUX_1.OUT.n2 INVERTER_MUX_1.OUT.n1 20.8576
R2957 INVERTER_MUX_1.OUT.n1 INVERTER_MUX_1.OUT.n0 20.8576
R2958 INVERTER_MUX_1.OUT.n10 INVERTER_MUX_1.OUT.n9 19.4672
R2959 INVERTER_MUX_1.OUT.n12 INVERTER_MUX_1.OUT.t22 19.4237
R2960 INVERTER_MUX_1.OUT.n10 INVERTER_MUX_1.OUT.t17 18.2505
R2961 INVERTER_MUX_1.OUT.n11 INVERTER_MUX_1.OUT.t33 18.2505
R2962 INVERTER_MUX_1.OUT.n10 INVERTER_MUX_1.OUT.t26 18.2505
R2963 INVERTER_MUX_1.OUT.t22 INVERTER_MUX_1.OUT.n11 18.2505
R2964 INVERTER_MUX_1.OUT.n9 INVERTER_MUX_1.OUT.n8 15.8172
R2965 INVERTER_MUX_1.OUT.n8 INVERTER_MUX_1.OUT.n7 15.8172
R2966 INVERTER_MUX_1.OUT.n7 INVERTER_MUX_1.OUT.n6 15.8172
R2967 INVERTER_MUX_1.OUT.n6 INVERTER_MUX_1.OUT.n5 15.8172
R2968 INVERTER_MUX_1.OUT.n1 INVERTER_MUX_1.OUT.t20 15.6434
R2969 INVERTER_MUX_1.OUT.n2 INVERTER_MUX_1.OUT.t16 15.6434
R2970 INVERTER_MUX_1.OUT.n3 INVERTER_MUX_1.OUT.t32 15.6434
R2971 INVERTER_MUX_1.OUT.n4 INVERTER_MUX_1.OUT.t28 15.6434
R2972 INVERTER_MUX_1.OUT.n0 INVERTER_MUX_1.OUT.t26 15.6434
R2973 INVERTER_MUX_1.OUT INVERTER_MUX_1.OUT.n12 8.63236
R2974 INVERTER_MUX_1.OUT.n27 INVERTER_MUX_1.OUT.n26 3.61224
R2975 INVERTER_MUX_1.OUT.n22 INVERTER_MUX_1.OUT.n21 3.61224
R2976 INVERTER_MUX_1.OUT.n24 INVERTER_MUX_1.OUT.t14 3.2765
R2977 INVERTER_MUX_1.OUT.n24 INVERTER_MUX_1.OUT.n23 3.2765
R2978 INVERTER_MUX_1.OUT.n26 INVERTER_MUX_1.OUT.t12 3.2765
R2979 INVERTER_MUX_1.OUT.n26 INVERTER_MUX_1.OUT.n25 3.2765
R2980 INVERTER_MUX_1.OUT.n19 INVERTER_MUX_1.OUT.t8 3.2765
R2981 INVERTER_MUX_1.OUT.n19 INVERTER_MUX_1.OUT.n18 3.2765
R2982 INVERTER_MUX_1.OUT.n21 INVERTER_MUX_1.OUT.t4 3.2765
R2983 INVERTER_MUX_1.OUT.n21 INVERTER_MUX_1.OUT.n20 3.2765
R2984 INVERTER_MUX_1.OUT.n17 INVERTER_MUX_1.OUT.n14 3.25789
R2985 INVERTER_MUX_1.OUT.n32 INVERTER_MUX_1.OUT.n29 3.25789
R2986 INVERTER_MUX_1.OUT.n27 INVERTER_MUX_1.OUT.n24 3.1505
R2987 INVERTER_MUX_1.OUT.n22 INVERTER_MUX_1.OUT.n19 3.1505
R2988 INVERTER_MUX_1.OUT.n17 INVERTER_MUX_1.OUT.n16 2.6005
R2989 INVERTER_MUX_1.OUT.n32 INVERTER_MUX_1.OUT.n31 2.6005
R2990 INVERTER_MUX_1.OUT.n29 INVERTER_MUX_1.OUT.t13 1.8205
R2991 INVERTER_MUX_1.OUT.n29 INVERTER_MUX_1.OUT.n28 1.8205
R2992 INVERTER_MUX_1.OUT.n16 INVERTER_MUX_1.OUT.t2 1.8205
R2993 INVERTER_MUX_1.OUT.n16 INVERTER_MUX_1.OUT.n15 1.8205
R2994 INVERTER_MUX_1.OUT.n14 INVERTER_MUX_1.OUT.t5 1.8205
R2995 INVERTER_MUX_1.OUT.n14 INVERTER_MUX_1.OUT.n13 1.8205
R2996 INVERTER_MUX_1.OUT.n31 INVERTER_MUX_1.OUT.t15 1.8205
R2997 INVERTER_MUX_1.OUT.n31 INVERTER_MUX_1.OUT.n30 1.8205
R2998 INVERTER_MUX_1.OUT.n34 INVERTER_MUX_1.OUT.n33 0.626587
R2999 INVERTER_MUX_1.OUT.n34 INVERTER_MUX_1.OUT.n17 0.427022
R3000 INVERTER_MUX_1.OUT.n33 INVERTER_MUX_1.OUT.n32 0.427022
R3001 INVERTER_MUX_1.OUT INVERTER_MUX_1.OUT.n34 0.278778
R3002 INVERTER_MUX_1.OUT.n33 INVERTER_MUX_1.OUT.n27 0.26463
R3003 INVERTER_MUX_1.OUT.n34 INVERTER_MUX_1.OUT.n22 0.26463
R3004 TG_magic_0.B.n64 TG_magic_0.B.n63 5.44589
R3005 TG_magic_0.B.n93 TG_magic_0.B.n91 5.07789
R3006 TG_magic_0.B.n68 TG_magic_0.B.t35 4.7885
R3007 TG_magic_0.B.n67 TG_magic_0.B.t32 4.7885
R3008 TG_magic_0.B.n64 TG_magic_0.B.n62 4.7885
R3009 TG_magic_0.B.n103 TG_magic_0.B.t99 4.4205
R3010 TG_magic_0.B.n102 TG_magic_0.B.t104 4.4205
R3011 TG_magic_0.B.n101 TG_magic_0.B.t13 4.4205
R3012 TG_magic_0.B.n100 TG_magic_0.B.t46 4.4205
R3013 TG_magic_0.B.n97 TG_magic_0.B.n96 4.4205
R3014 TG_magic_0.B.n95 TG_magic_0.B.n94 4.4205
R3015 TG_magic_0.B.n93 TG_magic_0.B.n92 4.4205
R3016 TG_magic_0.B.n134 TG_magic_0.B.n131 3.80789
R3017 TG_magic_0.B.n139 TG_magic_0.B.n136 3.80789
R3018 TG_magic_0.B.n32 TG_magic_0.B.n29 3.80789
R3019 TG_magic_0.B.n27 TG_magic_0.B.n24 3.80789
R3020 TG_magic_0.B.n38 TG_magic_0.B.n35 3.80789
R3021 TG_magic_0.B.n56 TG_magic_0.B.n55 3.80789
R3022 TG_magic_0.B.n61 TG_magic_0.B.n60 3.80789
R3023 TG_magic_0.B.n144 TG_magic_0.B.n141 3.80789
R3024 TG_magic_0.B.n8 TG_magic_0.B.n7 3.25789
R3025 TG_magic_0.B.n19 TG_magic_0.B.n18 3.25789
R3026 TG_magic_0.B.n48 TG_magic_0.B.n47 3.25789
R3027 TG_magic_0.B.n84 TG_magic_0.B.n81 3.25789
R3028 TG_magic_0.B.n73 TG_magic_0.B.n70 3.25789
R3029 TG_magic_0.B.n126 TG_magic_0.B.n125 3.25789
R3030 TG_magic_0.B.n115 TG_magic_0.B.n114 3.25789
R3031 TG_magic_0.B.n155 TG_magic_0.B.n154 3.25789
R3032 TG_magic_0.B.n134 TG_magic_0.B.n133 3.1505
R3033 TG_magic_0.B.n139 TG_magic_0.B.n138 3.1505
R3034 TG_magic_0.B.n32 TG_magic_0.B.n31 3.1505
R3035 TG_magic_0.B.n27 TG_magic_0.B.n26 3.1505
R3036 TG_magic_0.B.n38 TG_magic_0.B.n37 3.1505
R3037 TG_magic_0.B.n56 TG_magic_0.B.n53 3.1505
R3038 TG_magic_0.B.n61 TG_magic_0.B.n58 3.1505
R3039 TG_magic_0.B.n144 TG_magic_0.B.n143 3.1505
R3040 TG_magic_0.B.n106 TG_magic_0.B.n105 2.8437
R3041 TG_magic_0.B.n8 TG_magic_0.B.n5 2.6005
R3042 TG_magic_0.B.n9 TG_magic_0.B.n3 2.6005
R3043 TG_magic_0.B.n10 TG_magic_0.B.n1 2.6005
R3044 TG_magic_0.B.n19 TG_magic_0.B.n16 2.6005
R3045 TG_magic_0.B.n20 TG_magic_0.B.n14 2.6005
R3046 TG_magic_0.B.n21 TG_magic_0.B.n12 2.6005
R3047 TG_magic_0.B.n48 TG_magic_0.B.n45 2.6005
R3048 TG_magic_0.B.n49 TG_magic_0.B.n43 2.6005
R3049 TG_magic_0.B.n50 TG_magic_0.B.n41 2.6005
R3050 TG_magic_0.B.n84 TG_magic_0.B.n83 2.6005
R3051 TG_magic_0.B.n87 TG_magic_0.B.n86 2.6005
R3052 TG_magic_0.B.n90 TG_magic_0.B.n89 2.6005
R3053 TG_magic_0.B.n73 TG_magic_0.B.n72 2.6005
R3054 TG_magic_0.B.n76 TG_magic_0.B.n75 2.6005
R3055 TG_magic_0.B.n79 TG_magic_0.B.n78 2.6005
R3056 TG_magic_0.B.n126 TG_magic_0.B.n123 2.6005
R3057 TG_magic_0.B.n127 TG_magic_0.B.n121 2.6005
R3058 TG_magic_0.B.n128 TG_magic_0.B.n119 2.6005
R3059 TG_magic_0.B.n115 TG_magic_0.B.n112 2.6005
R3060 TG_magic_0.B.n116 TG_magic_0.B.n110 2.6005
R3061 TG_magic_0.B.n117 TG_magic_0.B.n108 2.6005
R3062 TG_magic_0.B.n155 TG_magic_0.B.n152 2.6005
R3063 TG_magic_0.B.n156 TG_magic_0.B.n150 2.6005
R3064 TG_magic_0.B.n157 TG_magic_0.B.n148 2.6005
R3065 TG_magic_0.B.n1 TG_magic_0.B.t64 1.8205
R3066 TG_magic_0.B.n1 TG_magic_0.B.n0 1.8205
R3067 TG_magic_0.B.n3 TG_magic_0.B.t70 1.8205
R3068 TG_magic_0.B.n3 TG_magic_0.B.n2 1.8205
R3069 TG_magic_0.B.n5 TG_magic_0.B.t60 1.8205
R3070 TG_magic_0.B.n5 TG_magic_0.B.n4 1.8205
R3071 TG_magic_0.B.n7 TG_magic_0.B.t67 1.8205
R3072 TG_magic_0.B.n7 TG_magic_0.B.n6 1.8205
R3073 TG_magic_0.B.n12 TG_magic_0.B.t24 1.8205
R3074 TG_magic_0.B.n12 TG_magic_0.B.n11 1.8205
R3075 TG_magic_0.B.n14 TG_magic_0.B.t53 1.8205
R3076 TG_magic_0.B.n14 TG_magic_0.B.n13 1.8205
R3077 TG_magic_0.B.n16 TG_magic_0.B.t63 1.8205
R3078 TG_magic_0.B.n16 TG_magic_0.B.n15 1.8205
R3079 TG_magic_0.B.n18 TG_magic_0.B.t75 1.8205
R3080 TG_magic_0.B.n18 TG_magic_0.B.n17 1.8205
R3081 TG_magic_0.B.n41 TG_magic_0.B.t69 1.8205
R3082 TG_magic_0.B.n41 TG_magic_0.B.n40 1.8205
R3083 TG_magic_0.B.n43 TG_magic_0.B.t62 1.8205
R3084 TG_magic_0.B.n43 TG_magic_0.B.n42 1.8205
R3085 TG_magic_0.B.n45 TG_magic_0.B.t73 1.8205
R3086 TG_magic_0.B.n45 TG_magic_0.B.n44 1.8205
R3087 TG_magic_0.B.n47 TG_magic_0.B.t74 1.8205
R3088 TG_magic_0.B.n47 TG_magic_0.B.n46 1.8205
R3089 TG_magic_0.B.n89 TG_magic_0.B.t22 1.8205
R3090 TG_magic_0.B.n89 TG_magic_0.B.n88 1.8205
R3091 TG_magic_0.B.n86 TG_magic_0.B.t11 1.8205
R3092 TG_magic_0.B.n86 TG_magic_0.B.n85 1.8205
R3093 TG_magic_0.B.n83 TG_magic_0.B.t101 1.8205
R3094 TG_magic_0.B.n83 TG_magic_0.B.n82 1.8205
R3095 TG_magic_0.B.n81 TG_magic_0.B.t23 1.8205
R3096 TG_magic_0.B.n81 TG_magic_0.B.n80 1.8205
R3097 TG_magic_0.B.n78 TG_magic_0.B.t16 1.8205
R3098 TG_magic_0.B.n78 TG_magic_0.B.n77 1.8205
R3099 TG_magic_0.B.n75 TG_magic_0.B.t102 1.8205
R3100 TG_magic_0.B.n75 TG_magic_0.B.n74 1.8205
R3101 TG_magic_0.B.n72 TG_magic_0.B.t20 1.8205
R3102 TG_magic_0.B.n72 TG_magic_0.B.n71 1.8205
R3103 TG_magic_0.B.n70 TG_magic_0.B.t17 1.8205
R3104 TG_magic_0.B.n70 TG_magic_0.B.n69 1.8205
R3105 TG_magic_0.B.n119 TG_magic_0.B.t85 1.8205
R3106 TG_magic_0.B.n119 TG_magic_0.B.n118 1.8205
R3107 TG_magic_0.B.n121 TG_magic_0.B.t61 1.8205
R3108 TG_magic_0.B.n121 TG_magic_0.B.n120 1.8205
R3109 TG_magic_0.B.n123 TG_magic_0.B.t5 1.8205
R3110 TG_magic_0.B.n123 TG_magic_0.B.n122 1.8205
R3111 TG_magic_0.B.n125 TG_magic_0.B.t9 1.8205
R3112 TG_magic_0.B.n125 TG_magic_0.B.n124 1.8205
R3113 TG_magic_0.B.n108 TG_magic_0.B.t1 1.8205
R3114 TG_magic_0.B.n108 TG_magic_0.B.n107 1.8205
R3115 TG_magic_0.B.n110 TG_magic_0.B.t4 1.8205
R3116 TG_magic_0.B.n110 TG_magic_0.B.n109 1.8205
R3117 TG_magic_0.B.n112 TG_magic_0.B.t10 1.8205
R3118 TG_magic_0.B.n112 TG_magic_0.B.n111 1.8205
R3119 TG_magic_0.B.n114 TG_magic_0.B.t82 1.8205
R3120 TG_magic_0.B.n114 TG_magic_0.B.n113 1.8205
R3121 TG_magic_0.B.n148 TG_magic_0.B.t77 1.8205
R3122 TG_magic_0.B.n148 TG_magic_0.B.n147 1.8205
R3123 TG_magic_0.B.n150 TG_magic_0.B.t80 1.8205
R3124 TG_magic_0.B.n150 TG_magic_0.B.n149 1.8205
R3125 TG_magic_0.B.n152 TG_magic_0.B.t55 1.8205
R3126 TG_magic_0.B.n152 TG_magic_0.B.n151 1.8205
R3127 TG_magic_0.B.n154 TG_magic_0.B.t3 1.8205
R3128 TG_magic_0.B.n154 TG_magic_0.B.n153 1.8205
R3129 TG_magic_0.B.n143 TG_magic_0.B.t96 1.6385
R3130 TG_magic_0.B.n143 TG_magic_0.B.n142 1.6385
R3131 TG_magic_0.B.n133 TG_magic_0.B.t93 1.6385
R3132 TG_magic_0.B.n133 TG_magic_0.B.n132 1.6385
R3133 TG_magic_0.B.n131 TG_magic_0.B.t94 1.6385
R3134 TG_magic_0.B.n131 TG_magic_0.B.n130 1.6385
R3135 TG_magic_0.B.n138 TG_magic_0.B.t89 1.6385
R3136 TG_magic_0.B.n138 TG_magic_0.B.n137 1.6385
R3137 TG_magic_0.B.n136 TG_magic_0.B.t92 1.6385
R3138 TG_magic_0.B.n136 TG_magic_0.B.n135 1.6385
R3139 TG_magic_0.B.n31 TG_magic_0.B.t39 1.6385
R3140 TG_magic_0.B.n31 TG_magic_0.B.n30 1.6385
R3141 TG_magic_0.B.n29 TG_magic_0.B.t37 1.6385
R3142 TG_magic_0.B.n29 TG_magic_0.B.n28 1.6385
R3143 TG_magic_0.B.n26 TG_magic_0.B.t48 1.6385
R3144 TG_magic_0.B.n26 TG_magic_0.B.n25 1.6385
R3145 TG_magic_0.B.n24 TG_magic_0.B.t43 1.6385
R3146 TG_magic_0.B.n24 TG_magic_0.B.n23 1.6385
R3147 TG_magic_0.B.n37 TG_magic_0.B.t47 1.6385
R3148 TG_magic_0.B.n37 TG_magic_0.B.n36 1.6385
R3149 TG_magic_0.B.n35 TG_magic_0.B.t42 1.6385
R3150 TG_magic_0.B.n35 TG_magic_0.B.n34 1.6385
R3151 TG_magic_0.B.n53 TG_magic_0.B.t36 1.6385
R3152 TG_magic_0.B.n53 TG_magic_0.B.n52 1.6385
R3153 TG_magic_0.B.n55 TG_magic_0.B.t33 1.6385
R3154 TG_magic_0.B.n55 TG_magic_0.B.n54 1.6385
R3155 TG_magic_0.B.n58 TG_magic_0.B.t31 1.6385
R3156 TG_magic_0.B.n58 TG_magic_0.B.n57 1.6385
R3157 TG_magic_0.B.n60 TG_magic_0.B.t34 1.6385
R3158 TG_magic_0.B.n60 TG_magic_0.B.n59 1.6385
R3159 TG_magic_0.B.n141 TG_magic_0.B.t86 1.6385
R3160 TG_magic_0.B.n141 TG_magic_0.B.n140 1.6385
R3161 TG_magic_0.B.n105 TG_magic_0.B.n104 1.49583
R3162 TG_magic_0.B.n105 TG_magic_0.B 1.16766
R3163 TG_magic_0.B.n65 TG_magic_0.B.n64 0.884196
R3164 TG_magic_0.B.n67 TG_magic_0.B.n66 0.884196
R3165 TG_magic_0.B.n98 TG_magic_0.B.n97 0.882239
R3166 TG_magic_0.B.n100 TG_magic_0.B.n99 0.882239
R3167 TG_magic_0.B.n104 TG_magic_0.B.n68 0.8105
R3168 TG_magic_0.B.n10 TG_magic_0.B.n9 0.657891
R3169 TG_magic_0.B.n9 TG_magic_0.B.n8 0.657891
R3170 TG_magic_0.B.n20 TG_magic_0.B.n19 0.657891
R3171 TG_magic_0.B.n50 TG_magic_0.B.n49 0.657891
R3172 TG_magic_0.B.n49 TG_magic_0.B.n48 0.657891
R3173 TG_magic_0.B.n95 TG_magic_0.B.n93 0.657891
R3174 TG_magic_0.B.n97 TG_magic_0.B.n95 0.657891
R3175 TG_magic_0.B.n87 TG_magic_0.B.n84 0.657891
R3176 TG_magic_0.B.n90 TG_magic_0.B.n87 0.657891
R3177 TG_magic_0.B.n76 TG_magic_0.B.n73 0.657891
R3178 TG_magic_0.B.n79 TG_magic_0.B.n76 0.657891
R3179 TG_magic_0.B.n68 TG_magic_0.B.n67 0.657891
R3180 TG_magic_0.B.n103 TG_magic_0.B.n102 0.657891
R3181 TG_magic_0.B.n102 TG_magic_0.B.n101 0.657891
R3182 TG_magic_0.B.n101 TG_magic_0.B.n100 0.657891
R3183 TG_magic_0.B.n127 TG_magic_0.B.n126 0.657891
R3184 TG_magic_0.B.n117 TG_magic_0.B.n116 0.657891
R3185 TG_magic_0.B.n116 TG_magic_0.B.n115 0.657891
R3186 TG_magic_0.B.n157 TG_magic_0.B.n156 0.657891
R3187 TG_magic_0.B.n156 TG_magic_0.B.n155 0.657891
R3188 TG_magic_0.B.n21 TG_magic_0.B.n20 0.655976
R3189 TG_magic_0.B.n128 TG_magic_0.B.n127 0.655976
R3190 TG_magic_0.B.n22 TG_magic_0.B.n21 0.646796
R3191 TG_magic_0.B.n129 TG_magic_0.B.n128 0.645657
R3192 TG_magic_0.B.n99 TG_magic_0.B.n98 0.6005
R3193 TG_magic_0.B.n66 TG_magic_0.B.n65 0.6005
R3194 TG_magic_0.B.n33 TG_magic_0.B.n32 0.548416
R3195 TG_magic_0.B.n145 TG_magic_0.B.n144 0.548416
R3196 TG_magic_0.B.n51 TG_magic_0.B.n50 0.316429
R3197 TG_magic_0.B.n158 TG_magic_0.B.n157 0.316429
R3198 TG_magic_0.B.n146 TG_magic_0.B.n134 0.304838
R3199 TG_magic_0.B.n39 TG_magic_0.B.n38 0.304838
R3200 TG_magic_0.B TG_magic_0.B.n51 0.2873
R3201 TG_magic_0.B TG_magic_0.B.n158 0.2873
R3202 TG_magic_0.B.n145 TG_magic_0.B.n139 0.284196
R3203 TG_magic_0.B.n33 TG_magic_0.B.n27 0.284196
R3204 TG_magic_0.B.n66 TG_magic_0.B.n56 0.284196
R3205 TG_magic_0.B.n65 TG_magic_0.B.n61 0.284196
R3206 TG_magic_0.B.n158 TG_magic_0.B.n129 0.283032
R3207 TG_magic_0.B.n98 TG_magic_0.B.n90 0.282239
R3208 TG_magic_0.B.n99 TG_magic_0.B.n79 0.282239
R3209 TG_magic_0.B.n51 TG_magic_0.B.n22 0.281892
R3210 TG_magic_0.B.n22 TG_magic_0.B.n10 0.279866
R3211 TG_magic_0.B.n129 TG_magic_0.B.n117 0.279866
R3212 TG_magic_0.B.n39 TG_magic_0.B.n33 0.244078
R3213 TG_magic_0.B.n146 TG_magic_0.B.n145 0.244078
R3214 TG_magic_0.B.n104 TG_magic_0.B.n103 0.237239
R3215 TG_magic_0.B.n51 TG_magic_0.B.n39 0.136437
R3216 TG_magic_0.B.n158 TG_magic_0.B.n146 0.136437
R3217 TG_magic_0.B TG_magic_0.B.n106 0.0893
R3218 TG_magic_0.B.n106 TG_magic_0.B 0.0725
R3219 Vout.n4 Vout.n1 3.80789
R3220 Vout.n9 Vout.n6 3.80789
R3221 Vout.n15 Vout.n12 3.80789
R3222 Vout.n97 Vout.n96 3.80789
R3223 Vout.n92 Vout.n91 3.80789
R3224 Vout.n103 Vout.n102 3.80789
R3225 Vout.n36 Vout.n35 3.25789
R3226 Vout.n25 Vout.n24 3.25789
R3227 Vout.n48 Vout.n47 3.25789
R3228 Vout.n57 Vout.n54 3.25789
R3229 Vout.n68 Vout.n65 3.25789
R3230 Vout.n80 Vout.n77 3.25789
R3231 Vout.n4 Vout.n3 3.1505
R3232 Vout.n9 Vout.n8 3.1505
R3233 Vout.n15 Vout.n14 3.1505
R3234 Vout.n97 Vout.n94 3.1505
R3235 Vout.n92 Vout.n89 3.1505
R3236 Vout.n103 Vout.n100 3.1505
R3237 Vout.n36 Vout.n33 2.6005
R3238 Vout.n37 Vout.n31 2.6005
R3239 Vout.n38 Vout.n29 2.6005
R3240 Vout.n25 Vout.n22 2.6005
R3241 Vout.n26 Vout.n20 2.6005
R3242 Vout.n27 Vout.n18 2.6005
R3243 Vout.n48 Vout.n45 2.6005
R3244 Vout.n49 Vout.n43 2.6005
R3245 Vout.n50 Vout.n41 2.6005
R3246 Vout.n57 Vout.n56 2.6005
R3247 Vout.n60 Vout.n59 2.6005
R3248 Vout.n63 Vout.n62 2.6005
R3249 Vout.n68 Vout.n67 2.6005
R3250 Vout.n71 Vout.n70 2.6005
R3251 Vout.n74 Vout.n73 2.6005
R3252 Vout.n80 Vout.n79 2.6005
R3253 Vout.n83 Vout.n82 2.6005
R3254 Vout.n86 Vout.n85 2.6005
R3255 Vout.n29 Vout.t18 1.8205
R3256 Vout.n29 Vout.n28 1.8205
R3257 Vout.n31 Vout.t58 1.8205
R3258 Vout.n31 Vout.n30 1.8205
R3259 Vout.n33 Vout.t66 1.8205
R3260 Vout.n33 Vout.n32 1.8205
R3261 Vout.n35 Vout.t16 1.8205
R3262 Vout.n35 Vout.n34 1.8205
R3263 Vout.n18 Vout.t63 1.8205
R3264 Vout.n18 Vout.n17 1.8205
R3265 Vout.n20 Vout.t65 1.8205
R3266 Vout.n20 Vout.n19 1.8205
R3267 Vout.n22 Vout.t12 1.8205
R3268 Vout.n22 Vout.n21 1.8205
R3269 Vout.n24 Vout.t60 1.8205
R3270 Vout.n24 Vout.n23 1.8205
R3271 Vout.n41 Vout.t9 1.8205
R3272 Vout.n41 Vout.n40 1.8205
R3273 Vout.n43 Vout.t11 1.8205
R3274 Vout.n43 Vout.n42 1.8205
R3275 Vout.n45 Vout.t15 1.8205
R3276 Vout.n45 Vout.n44 1.8205
R3277 Vout.n47 Vout.t67 1.8205
R3278 Vout.n47 Vout.n46 1.8205
R3279 Vout.n62 Vout.t43 1.8205
R3280 Vout.n62 Vout.n61 1.8205
R3281 Vout.n59 Vout.t21 1.8205
R3282 Vout.n59 Vout.n58 1.8205
R3283 Vout.n56 Vout.t0 1.8205
R3284 Vout.n56 Vout.n55 1.8205
R3285 Vout.n54 Vout.t44 1.8205
R3286 Vout.n54 Vout.n53 1.8205
R3287 Vout.n73 Vout.t22 1.8205
R3288 Vout.n73 Vout.n72 1.8205
R3289 Vout.n70 Vout.t51 1.8205
R3290 Vout.n70 Vout.n69 1.8205
R3291 Vout.n67 Vout.t49 1.8205
R3292 Vout.n67 Vout.n66 1.8205
R3293 Vout.n65 Vout.t23 1.8205
R3294 Vout.n65 Vout.n64 1.8205
R3295 Vout.n85 Vout.t46 1.8205
R3296 Vout.n85 Vout.n84 1.8205
R3297 Vout.n82 Vout.t29 1.8205
R3298 Vout.n82 Vout.n81 1.8205
R3299 Vout.n79 Vout.t25 1.8205
R3300 Vout.n79 Vout.n78 1.8205
R3301 Vout.n77 Vout.t47 1.8205
R3302 Vout.n77 Vout.n76 1.8205
R3303 Vout.n3 Vout.t37 1.6385
R3304 Vout.n3 Vout.n2 1.6385
R3305 Vout.n1 Vout.t31 1.6385
R3306 Vout.n1 Vout.n0 1.6385
R3307 Vout.n6 Vout.t38 1.6385
R3308 Vout.n6 Vout.n5 1.6385
R3309 Vout.n8 Vout.t32 1.6385
R3310 Vout.n8 Vout.n7 1.6385
R3311 Vout.n14 Vout.t40 1.6385
R3312 Vout.n14 Vout.n13 1.6385
R3313 Vout.n12 Vout.t34 1.6385
R3314 Vout.n12 Vout.n11 1.6385
R3315 Vout.n94 Vout.t4 1.6385
R3316 Vout.n94 Vout.n93 1.6385
R3317 Vout.n96 Vout.t55 1.6385
R3318 Vout.n96 Vout.n95 1.6385
R3319 Vout.n89 Vout.t7 1.6385
R3320 Vout.n89 Vout.n88 1.6385
R3321 Vout.n91 Vout.t1 1.6385
R3322 Vout.n91 Vout.n90 1.6385
R3323 Vout.n100 Vout.t54 1.6385
R3324 Vout.n100 Vout.n99 1.6385
R3325 Vout.n102 Vout.t3 1.6385
R3326 Vout.n102 Vout.n101 1.6385
R3327 Vout.n37 Vout.n36 0.657891
R3328 Vout.n27 Vout.n26 0.657891
R3329 Vout.n26 Vout.n25 0.657891
R3330 Vout.n50 Vout.n49 0.657891
R3331 Vout.n49 Vout.n48 0.657891
R3332 Vout.n60 Vout.n57 0.657891
R3333 Vout.n63 Vout.n60 0.657891
R3334 Vout.n71 Vout.n68 0.657891
R3335 Vout.n83 Vout.n80 0.657891
R3336 Vout.n86 Vout.n83 0.657891
R3337 Vout.n38 Vout.n37 0.655976
R3338 Vout.n74 Vout.n71 0.655976
R3339 Vout.n39 Vout.n38 0.645657
R3340 Vout.n75 Vout.n74 0.645657
R3341 Vout.n10 Vout.n9 0.548416
R3342 Vout.n98 Vout.n97 0.548416
R3343 Vout.n104 Vout.n103 0.310609
R3344 Vout.n16 Vout.n15 0.309196
R3345 Vout.n87 Vout.n86 0.299432
R3346 Vout.n51 Vout.n50 0.297594
R3347 Vout.n10 Vout.n4 0.284196
R3348 Vout.n98 Vout.n92 0.284196
R3349 Vout.n39 Vout.n27 0.279866
R3350 Vout.n75 Vout.n63 0.279866
R3351 Vout.n87 Vout.n75 0.182778
R3352 Vout.n51 Vout.n39 0.166829
R3353 Vout.n104 Vout.n98 0.131784
R3354 Vout.n16 Vout.n10 0.120225
R3355 Vout Vout.n105 0.08654
R3356 Vout Vout.n52 0.0822871
R3357 Vout.n105 Vout.n104 0.0552826
R3358 Vout.n52 Vout.n16 0.0482273
R3359 Vout.n52 Vout.n51 0.0432273
R3360 Vout.n105 Vout.n87 0.0430543
R3361 S2.n12 S2.t27 68.1773
R3362 S2.n16 S2.n15 52.5344
R3363 S2.n17 S2.t29 47.0594
R3364 S2.t9 S2.t30 43.8005
R3365 S2.t18 S2.t9 43.8005
R3366 S2.t29 S2.t18 43.8005
R3367 S2.t15 S2.t19 43.8005
R3368 S2.t24 S2.t28 43.8005
R3369 S2.t33 S2.t3 43.8005
R3370 S2.t13 S2.t16 43.8005
R3371 S2.n9 S2.t20 33.763
R3372 S2.t25 S2.t17 30.7648
R3373 S2.t0 S2.t26 30.7648
R3374 S2.t4 S2.t1 30.7648
R3375 S2.t22 S2.t14 30.7648
R3376 S2.n0 S2.t25 30.3737
R3377 S2.n1 S2.t0 30.3737
R3378 S2.n2 S2.t4 30.3737
R3379 S2.n8 S2.t5 21.9005
R3380 S2.t20 S2.n8 21.9005
R3381 S2.n7 S2.t23 21.9005
R3382 S2.n7 S2.t7 21.9005
R3383 S2.n6 S2.t32 21.9005
R3384 S2.n6 S2.t11 21.9005
R3385 S2.n5 S2.t12 21.9005
R3386 S2.t2 S2.n5 21.9005
R3387 S2.n14 S2.t21 21.9005
R3388 S2.n14 S2.t6 21.9005
R3389 S2.n0 S2.t15 21.6398
R3390 S2.n1 S2.t24 21.6398
R3391 S2.n2 S2.t33 21.6398
R3392 S2.n3 S2.t13 21.6398
R3393 S2.n10 S2.n9 20.8576
R3394 S2.n11 S2.n10 20.8576
R3395 S2.n13 S2.n11 20.8576
R3396 S2.n13 S2.n12 20.8576
R3397 S2.n15 S2.n14 19.4672
R3398 S2.n17 S2.t8 19.4237
R3399 S2.n16 S2.t27 18.2505
R3400 S2.n15 S2.t10 18.2505
R3401 S2.n15 S2.t31 18.2505
R3402 S2.t8 S2.n16 18.2505
R3403 S2.n4 S2.t22 17.7827
R3404 S2.n1 S2.n0 17.255
R3405 S2.n2 S2.n1 17.255
R3406 S2.n3 S2.n2 17.255
R3407 S2.n8 S2.n7 15.8172
R3408 S2.n7 S2.n6 15.8172
R3409 S2.n6 S2.n5 15.8172
R3410 S2.n14 S2.n5 15.8172
R3411 S2.n9 S2.t7 15.6434
R3412 S2.n10 S2.t11 15.6434
R3413 S2.n11 S2.t2 15.6434
R3414 S2.t6 S2.n13 15.6434
R3415 S2.n12 S2.t10 15.6434
R3416 S2.n18 S2 9.47615
R3417 S2 S2.n17 8.63236
R3418 S2.n4 S2.n3 8.06475
R3419 S2 S2.n4 4.24369
R3420 S2 S2.n18 1.79166
R3421 S2.n18 S2 1.44502
R3422 a_n4297_n7438.t7 a_n4297_n7438.n19 40.7345
R3423 a_n4297_n7438.n24 a_n4297_n7438.n5 28.094
R3424 a_n4297_n7438.n21 a_n4297_n7438.n20 28.094
R3425 a_n4297_n7438.n32 a_n4297_n7438.n31 28.094
R3426 a_n4297_n7438.n26 a_n4297_n7438.t21 21.9005
R3427 a_n4297_n7438.n26 a_n4297_n7438.t17 21.9005
R3428 a_n4297_n7438.n0 a_n4297_n7438.t11 21.9005
R3429 a_n4297_n7438.n11 a_n4297_n7438.t22 21.9005
R3430 a_n4297_n7438.n12 a_n4297_n7438.t18 21.9005
R3431 a_n4297_n7438.n1 a_n4297_n7438.t8 21.9005
R3432 a_n4297_n7438.n27 a_n4297_n7438.t13 21.9005
R3433 a_n4297_n7438.n27 a_n4297_n7438.t16 21.9005
R3434 a_n4297_n7438.n28 a_n4297_n7438.t27 21.9005
R3435 a_n4297_n7438.n28 a_n4297_n7438.t24 21.9005
R3436 a_n4297_n7438.n2 a_n4297_n7438.t14 21.9005
R3437 a_n4297_n7438.n13 a_n4297_n7438.t28 21.9005
R3438 a_n4297_n7438.n14 a_n4297_n7438.t25 21.9005
R3439 a_n4297_n7438.n3 a_n4297_n7438.t12 21.9005
R3440 a_n4297_n7438.n29 a_n4297_n7438.t19 21.9005
R3441 a_n4297_n7438.n29 a_n4297_n7438.t23 21.9005
R3442 a_n4297_n7438.n30 a_n4297_n7438.t9 21.9005
R3443 a_n4297_n7438.n30 a_n4297_n7438.t6 21.9005
R3444 a_n4297_n7438.n4 a_n4297_n7438.t20 21.9005
R3445 a_n4297_n7438.n15 a_n4297_n7438.t10 21.9005
R3446 a_n4297_n7438.n20 a_n4297_n7438.t7 21.9005
R3447 a_n4297_n7438.n5 a_n4297_n7438.t15 21.9005
R3448 a_n4297_n7438.n31 a_n4297_n7438.t26 21.9005
R3449 a_n4297_n7438.n31 a_n4297_n7438.t29 21.9005
R3450 a_n4297_n7438.n20 a_n4297_n7438.n15 15.8172
R3451 a_n4297_n7438.n5 a_n4297_n7438.n4 15.8172
R3452 a_n4297_n7438.n4 a_n4297_n7438.n3 15.8172
R3453 a_n4297_n7438.n15 a_n4297_n7438.n14 15.8172
R3454 a_n4297_n7438.n14 a_n4297_n7438.n13 15.8172
R3455 a_n4297_n7438.n3 a_n4297_n7438.n2 15.8172
R3456 a_n4297_n7438.n2 a_n4297_n7438.n1 15.8172
R3457 a_n4297_n7438.n13 a_n4297_n7438.n12 15.8172
R3458 a_n4297_n7438.n12 a_n4297_n7438.n11 15.8172
R3459 a_n4297_n7438.n1 a_n4297_n7438.n0 15.8172
R3460 a_n4297_n7438.n27 a_n4297_n7438.n26 15.8172
R3461 a_n4297_n7438.n29 a_n4297_n7438.n28 15.8172
R3462 a_n4297_n7438.n28 a_n4297_n7438.n27 15.8172
R3463 a_n4297_n7438.n31 a_n4297_n7438.n30 15.8172
R3464 a_n4297_n7438.n30 a_n4297_n7438.n29 15.8172
R3465 a_n4297_n7438.n17 a_n4297_n7438.n16 15.1845
R3466 a_n4297_n7438.n19 a_n4297_n7438.n18 15.1845
R3467 a_n4297_n7438.n18 a_n4297_n7438.n17 15.1845
R3468 a_n4297_n7438.n8 a_n4297_n7438.n6 5.44589
R3469 a_n4297_n7438.n8 a_n4297_n7438.n7 4.7885
R3470 a_n4297_n7438.n32 a_n4297_n7438.n25 4.70615
R3471 a_n4297_n7438.n23 a_n4297_n7438.n22 4.4205
R3472 a_n4297_n7438.n10 a_n4297_n7438.n9 4.4205
R3473 a_n4297_n7438.n34 a_n4297_n7438.n33 4.4205
R3474 a_n4297_n7438.n10 a_n4297_n7438.n8 1.1392
R3475 a_n4297_n7438.n23 a_n4297_n7438.n21 0.286152
R3476 a_n4297_n7438.n33 a_n4297_n7438.n24 0.286152
R3477 a_n4297_n7438.n21 a_n4297_n7438.n10 0.282239
R3478 a_n4297_n7438.n24 a_n4297_n7438.n23 0.282239
R3479 a_n4297_n7438.n33 a_n4297_n7438.n32 0.282239
R3480 TG_GATE_SWITCH_magic_2.B.n54 TG_GATE_SWITCH_magic_2.B.n53 9.66506
R3481 TG_GATE_SWITCH_magic_2.B.n10 TG_GATE_SWITCH_magic_2.B.t5 5.44589
R3482 TG_GATE_SWITCH_magic_2.B.n43 TG_GATE_SWITCH_magic_2.B.t71 5.07789
R3483 TG_GATE_SWITCH_magic_2.B.n16 TG_GATE_SWITCH_magic_2.B.n15 4.7885
R3484 TG_GATE_SWITCH_magic_2.B.n14 TG_GATE_SWITCH_magic_2.B.n13 4.7885
R3485 TG_GATE_SWITCH_magic_2.B.n10 TG_GATE_SWITCH_magic_2.B.t9 4.7885
R3486 TG_GATE_SWITCH_magic_2.B.n51 TG_GATE_SWITCH_magic_2.B.n17 4.4205
R3487 TG_GATE_SWITCH_magic_2.B.n50 TG_GATE_SWITCH_magic_2.B.n18 4.4205
R3488 TG_GATE_SWITCH_magic_2.B.n49 TG_GATE_SWITCH_magic_2.B.n19 4.4205
R3489 TG_GATE_SWITCH_magic_2.B.n48 TG_GATE_SWITCH_magic_2.B.n20 4.4205
R3490 TG_GATE_SWITCH_magic_2.B.n45 TG_GATE_SWITCH_magic_2.B.t69 4.4205
R3491 TG_GATE_SWITCH_magic_2.B.n44 TG_GATE_SWITCH_magic_2.B.t50 4.4205
R3492 TG_GATE_SWITCH_magic_2.B.n43 TG_GATE_SWITCH_magic_2.B.t39 4.4205
R3493 TG_GATE_SWITCH_magic_2.B.n9 TG_GATE_SWITCH_magic_2.B.n8 3.80789
R3494 TG_GATE_SWITCH_magic_2.B.n4 TG_GATE_SWITCH_magic_2.B.n3 3.80789
R3495 TG_GATE_SWITCH_magic_2.B.n59 TG_GATE_SWITCH_magic_2.B.n56 3.80789
R3496 TG_GATE_SWITCH_magic_2.B.n64 TG_GATE_SWITCH_magic_2.B.n61 3.80789
R3497 TG_GATE_SWITCH_magic_2.B.n69 TG_GATE_SWITCH_magic_2.B.n66 3.80789
R3498 TG_GATE_SWITCH_magic_2.B.n25 TG_GATE_SWITCH_magic_2.B.n22 3.25789
R3499 TG_GATE_SWITCH_magic_2.B.n36 TG_GATE_SWITCH_magic_2.B.n33 3.25789
R3500 TG_GATE_SWITCH_magic_2.B.n80 TG_GATE_SWITCH_magic_2.B.n79 3.25789
R3501 TG_GATE_SWITCH_magic_2.B.n91 TG_GATE_SWITCH_magic_2.B.n90 3.25789
R3502 TG_GATE_SWITCH_magic_2.B.n102 TG_GATE_SWITCH_magic_2.B.n99 3.25789
R3503 TG_GATE_SWITCH_magic_2.B.n9 TG_GATE_SWITCH_magic_2.B.n6 3.1505
R3504 TG_GATE_SWITCH_magic_2.B.n4 TG_GATE_SWITCH_magic_2.B.n1 3.1505
R3505 TG_GATE_SWITCH_magic_2.B.n59 TG_GATE_SWITCH_magic_2.B.n58 3.1505
R3506 TG_GATE_SWITCH_magic_2.B.n64 TG_GATE_SWITCH_magic_2.B.n63 3.1505
R3507 TG_GATE_SWITCH_magic_2.B.n69 TG_GATE_SWITCH_magic_2.B.n68 3.1505
R3508 TG_GATE_SWITCH_magic_2.B.n25 TG_GATE_SWITCH_magic_2.B.n24 2.6005
R3509 TG_GATE_SWITCH_magic_2.B.n28 TG_GATE_SWITCH_magic_2.B.n27 2.6005
R3510 TG_GATE_SWITCH_magic_2.B.n31 TG_GATE_SWITCH_magic_2.B.n30 2.6005
R3511 TG_GATE_SWITCH_magic_2.B.n36 TG_GATE_SWITCH_magic_2.B.n35 2.6005
R3512 TG_GATE_SWITCH_magic_2.B.n39 TG_GATE_SWITCH_magic_2.B.n38 2.6005
R3513 TG_GATE_SWITCH_magic_2.B.n42 TG_GATE_SWITCH_magic_2.B.n41 2.6005
R3514 TG_GATE_SWITCH_magic_2.B.n80 TG_GATE_SWITCH_magic_2.B.n77 2.6005
R3515 TG_GATE_SWITCH_magic_2.B.n81 TG_GATE_SWITCH_magic_2.B.n75 2.6005
R3516 TG_GATE_SWITCH_magic_2.B.n82 TG_GATE_SWITCH_magic_2.B.n73 2.6005
R3517 TG_GATE_SWITCH_magic_2.B.n91 TG_GATE_SWITCH_magic_2.B.n88 2.6005
R3518 TG_GATE_SWITCH_magic_2.B.n92 TG_GATE_SWITCH_magic_2.B.n86 2.6005
R3519 TG_GATE_SWITCH_magic_2.B.n93 TG_GATE_SWITCH_magic_2.B.n84 2.6005
R3520 TG_GATE_SWITCH_magic_2.B.n104 TG_GATE_SWITCH_magic_2.B.n95 2.6005
R3521 TG_GATE_SWITCH_magic_2.B.n103 TG_GATE_SWITCH_magic_2.B.n97 2.6005
R3522 TG_GATE_SWITCH_magic_2.B.n102 TG_GATE_SWITCH_magic_2.B.n101 2.6005
R3523 TG_GATE_SWITCH_magic_2.B TG_GATE_SWITCH_magic_2.B.n54 2.32408
R3524 TG_GATE_SWITCH_magic_2.B.n97 TG_GATE_SWITCH_magic_2.B.t17 1.8205
R3525 TG_GATE_SWITCH_magic_2.B.n97 TG_GATE_SWITCH_magic_2.B.n96 1.8205
R3526 TG_GATE_SWITCH_magic_2.B.n99 TG_GATE_SWITCH_magic_2.B.t22 1.8205
R3527 TG_GATE_SWITCH_magic_2.B.n99 TG_GATE_SWITCH_magic_2.B.n98 1.8205
R3528 TG_GATE_SWITCH_magic_2.B.n95 TG_GATE_SWITCH_magic_2.B.t21 1.8205
R3529 TG_GATE_SWITCH_magic_2.B.n95 TG_GATE_SWITCH_magic_2.B.n94 1.8205
R3530 TG_GATE_SWITCH_magic_2.B.n30 TG_GATE_SWITCH_magic_2.B.t48 1.8205
R3531 TG_GATE_SWITCH_magic_2.B.n30 TG_GATE_SWITCH_magic_2.B.n29 1.8205
R3532 TG_GATE_SWITCH_magic_2.B.n27 TG_GATE_SWITCH_magic_2.B.t42 1.8205
R3533 TG_GATE_SWITCH_magic_2.B.n27 TG_GATE_SWITCH_magic_2.B.n26 1.8205
R3534 TG_GATE_SWITCH_magic_2.B.n24 TG_GATE_SWITCH_magic_2.B.t67 1.8205
R3535 TG_GATE_SWITCH_magic_2.B.n24 TG_GATE_SWITCH_magic_2.B.n23 1.8205
R3536 TG_GATE_SWITCH_magic_2.B.n22 TG_GATE_SWITCH_magic_2.B.t49 1.8205
R3537 TG_GATE_SWITCH_magic_2.B.n22 TG_GATE_SWITCH_magic_2.B.n21 1.8205
R3538 TG_GATE_SWITCH_magic_2.B.n41 TG_GATE_SWITCH_magic_2.B.t43 1.8205
R3539 TG_GATE_SWITCH_magic_2.B.n41 TG_GATE_SWITCH_magic_2.B.n40 1.8205
R3540 TG_GATE_SWITCH_magic_2.B.n38 TG_GATE_SWITCH_magic_2.B.t40 1.8205
R3541 TG_GATE_SWITCH_magic_2.B.n38 TG_GATE_SWITCH_magic_2.B.n37 1.8205
R3542 TG_GATE_SWITCH_magic_2.B.n35 TG_GATE_SWITCH_magic_2.B.t47 1.8205
R3543 TG_GATE_SWITCH_magic_2.B.n35 TG_GATE_SWITCH_magic_2.B.n34 1.8205
R3544 TG_GATE_SWITCH_magic_2.B.n33 TG_GATE_SWITCH_magic_2.B.t44 1.8205
R3545 TG_GATE_SWITCH_magic_2.B.n33 TG_GATE_SWITCH_magic_2.B.n32 1.8205
R3546 TG_GATE_SWITCH_magic_2.B.n73 TG_GATE_SWITCH_magic_2.B.t15 1.8205
R3547 TG_GATE_SWITCH_magic_2.B.n73 TG_GATE_SWITCH_magic_2.B.n72 1.8205
R3548 TG_GATE_SWITCH_magic_2.B.n75 TG_GATE_SWITCH_magic_2.B.t20 1.8205
R3549 TG_GATE_SWITCH_magic_2.B.n75 TG_GATE_SWITCH_magic_2.B.n74 1.8205
R3550 TG_GATE_SWITCH_magic_2.B.n77 TG_GATE_SWITCH_magic_2.B.t18 1.8205
R3551 TG_GATE_SWITCH_magic_2.B.n77 TG_GATE_SWITCH_magic_2.B.n76 1.8205
R3552 TG_GATE_SWITCH_magic_2.B.n79 TG_GATE_SWITCH_magic_2.B.t16 1.8205
R3553 TG_GATE_SWITCH_magic_2.B.n79 TG_GATE_SWITCH_magic_2.B.n78 1.8205
R3554 TG_GATE_SWITCH_magic_2.B.n84 TG_GATE_SWITCH_magic_2.B.t12 1.8205
R3555 TG_GATE_SWITCH_magic_2.B.n84 TG_GATE_SWITCH_magic_2.B.n83 1.8205
R3556 TG_GATE_SWITCH_magic_2.B.n86 TG_GATE_SWITCH_magic_2.B.t19 1.8205
R3557 TG_GATE_SWITCH_magic_2.B.n86 TG_GATE_SWITCH_magic_2.B.n85 1.8205
R3558 TG_GATE_SWITCH_magic_2.B.n88 TG_GATE_SWITCH_magic_2.B.t14 1.8205
R3559 TG_GATE_SWITCH_magic_2.B.n88 TG_GATE_SWITCH_magic_2.B.n87 1.8205
R3560 TG_GATE_SWITCH_magic_2.B.n90 TG_GATE_SWITCH_magic_2.B.t13 1.8205
R3561 TG_GATE_SWITCH_magic_2.B.n90 TG_GATE_SWITCH_magic_2.B.n89 1.8205
R3562 TG_GATE_SWITCH_magic_2.B.n101 TG_GATE_SWITCH_magic_2.B.t23 1.8205
R3563 TG_GATE_SWITCH_magic_2.B.n101 TG_GATE_SWITCH_magic_2.B.n100 1.8205
R3564 TG_GATE_SWITCH_magic_2.B.n53 TG_GATE_SWITCH_magic_2.B.n52 1.80703
R3565 TG_GATE_SWITCH_magic_2.B.n6 TG_GATE_SWITCH_magic_2.B.t4 1.6385
R3566 TG_GATE_SWITCH_magic_2.B.n6 TG_GATE_SWITCH_magic_2.B.n5 1.6385
R3567 TG_GATE_SWITCH_magic_2.B.n8 TG_GATE_SWITCH_magic_2.B.t11 1.6385
R3568 TG_GATE_SWITCH_magic_2.B.n8 TG_GATE_SWITCH_magic_2.B.n7 1.6385
R3569 TG_GATE_SWITCH_magic_2.B.n1 TG_GATE_SWITCH_magic_2.B.t1 1.6385
R3570 TG_GATE_SWITCH_magic_2.B.n1 TG_GATE_SWITCH_magic_2.B.n0 1.6385
R3571 TG_GATE_SWITCH_magic_2.B.n3 TG_GATE_SWITCH_magic_2.B.t7 1.6385
R3572 TG_GATE_SWITCH_magic_2.B.n3 TG_GATE_SWITCH_magic_2.B.n2 1.6385
R3573 TG_GATE_SWITCH_magic_2.B.n58 TG_GATE_SWITCH_magic_2.B.t58 1.6385
R3574 TG_GATE_SWITCH_magic_2.B.n58 TG_GATE_SWITCH_magic_2.B.n57 1.6385
R3575 TG_GATE_SWITCH_magic_2.B.n56 TG_GATE_SWITCH_magic_2.B.t59 1.6385
R3576 TG_GATE_SWITCH_magic_2.B.n56 TG_GATE_SWITCH_magic_2.B.n55 1.6385
R3577 TG_GATE_SWITCH_magic_2.B.n63 TG_GATE_SWITCH_magic_2.B.t56 1.6385
R3578 TG_GATE_SWITCH_magic_2.B.n63 TG_GATE_SWITCH_magic_2.B.n62 1.6385
R3579 TG_GATE_SWITCH_magic_2.B.n61 TG_GATE_SWITCH_magic_2.B.t57 1.6385
R3580 TG_GATE_SWITCH_magic_2.B.n61 TG_GATE_SWITCH_magic_2.B.n60 1.6385
R3581 TG_GATE_SWITCH_magic_2.B.n66 TG_GATE_SWITCH_magic_2.B.t55 1.6385
R3582 TG_GATE_SWITCH_magic_2.B.n66 TG_GATE_SWITCH_magic_2.B.n65 1.6385
R3583 TG_GATE_SWITCH_magic_2.B.n68 TG_GATE_SWITCH_magic_2.B.t54 1.6385
R3584 TG_GATE_SWITCH_magic_2.B.n68 TG_GATE_SWITCH_magic_2.B.n67 1.6385
R3585 TG_GATE_SWITCH_magic_2.B.n53 TG_GATE_SWITCH_magic_2.B 1.16601
R3586 TG_GATE_SWITCH_magic_2.B.n11 TG_GATE_SWITCH_magic_2.B.n10 0.884196
R3587 TG_GATE_SWITCH_magic_2.B.n14 TG_GATE_SWITCH_magic_2.B.n12 0.884196
R3588 TG_GATE_SWITCH_magic_2.B.n46 TG_GATE_SWITCH_magic_2.B.n45 0.882239
R3589 TG_GATE_SWITCH_magic_2.B.n48 TG_GATE_SWITCH_magic_2.B.n47 0.882239
R3590 TG_GATE_SWITCH_magic_2.B.n52 TG_GATE_SWITCH_magic_2.B.n16 0.8105
R3591 TG_GATE_SWITCH_magic_2.B.n28 TG_GATE_SWITCH_magic_2.B.n25 0.657891
R3592 TG_GATE_SWITCH_magic_2.B.n31 TG_GATE_SWITCH_magic_2.B.n28 0.657891
R3593 TG_GATE_SWITCH_magic_2.B.n39 TG_GATE_SWITCH_magic_2.B.n36 0.657891
R3594 TG_GATE_SWITCH_magic_2.B.n42 TG_GATE_SWITCH_magic_2.B.n39 0.657891
R3595 TG_GATE_SWITCH_magic_2.B.n44 TG_GATE_SWITCH_magic_2.B.n43 0.657891
R3596 TG_GATE_SWITCH_magic_2.B.n45 TG_GATE_SWITCH_magic_2.B.n44 0.657891
R3597 TG_GATE_SWITCH_magic_2.B.n16 TG_GATE_SWITCH_magic_2.B.n14 0.657891
R3598 TG_GATE_SWITCH_magic_2.B.n51 TG_GATE_SWITCH_magic_2.B.n50 0.657891
R3599 TG_GATE_SWITCH_magic_2.B.n50 TG_GATE_SWITCH_magic_2.B.n49 0.657891
R3600 TG_GATE_SWITCH_magic_2.B.n49 TG_GATE_SWITCH_magic_2.B.n48 0.657891
R3601 TG_GATE_SWITCH_magic_2.B.n82 TG_GATE_SWITCH_magic_2.B.n81 0.657891
R3602 TG_GATE_SWITCH_magic_2.B.n81 TG_GATE_SWITCH_magic_2.B.n80 0.657891
R3603 TG_GATE_SWITCH_magic_2.B.n93 TG_GATE_SWITCH_magic_2.B.n92 0.657891
R3604 TG_GATE_SWITCH_magic_2.B.n92 TG_GATE_SWITCH_magic_2.B.n91 0.657891
R3605 TG_GATE_SWITCH_magic_2.B.n103 TG_GATE_SWITCH_magic_2.B.n102 0.657891
R3606 TG_GATE_SWITCH_magic_2.B.n104 TG_GATE_SWITCH_magic_2.B.n103 0.655976
R3607 TG_GATE_SWITCH_magic_2.B.n105 TG_GATE_SWITCH_magic_2.B.n104 0.645657
R3608 TG_GATE_SWITCH_magic_2.B.n47 TG_GATE_SWITCH_magic_2.B.n46 0.6005
R3609 TG_GATE_SWITCH_magic_2.B.n12 TG_GATE_SWITCH_magic_2.B.n11 0.6005
R3610 TG_GATE_SWITCH_magic_2.B.n70 TG_GATE_SWITCH_magic_2.B.n69 0.548416
R3611 TG_GATE_SWITCH_magic_2.B.n106 TG_GATE_SWITCH_magic_2.B.n82 0.316429
R3612 TG_GATE_SWITCH_magic_2.B.n71 TG_GATE_SWITCH_magic_2.B.n59 0.304838
R3613 TG_GATE_SWITCH_magic_2.B.n11 TG_GATE_SWITCH_magic_2.B.n9 0.284196
R3614 TG_GATE_SWITCH_magic_2.B.n12 TG_GATE_SWITCH_magic_2.B.n4 0.284196
R3615 TG_GATE_SWITCH_magic_2.B.n70 TG_GATE_SWITCH_magic_2.B.n64 0.284196
R3616 TG_GATE_SWITCH_magic_2.B.n106 TG_GATE_SWITCH_magic_2.B.n105 0.283032
R3617 TG_GATE_SWITCH_magic_2.B.n47 TG_GATE_SWITCH_magic_2.B.n31 0.282239
R3618 TG_GATE_SWITCH_magic_2.B.n46 TG_GATE_SWITCH_magic_2.B.n42 0.282239
R3619 TG_GATE_SWITCH_magic_2.B.n105 TG_GATE_SWITCH_magic_2.B.n93 0.279866
R3620 TG_GATE_SWITCH_magic_2.B.n71 TG_GATE_SWITCH_magic_2.B.n70 0.244078
R3621 TG_GATE_SWITCH_magic_2.B.n52 TG_GATE_SWITCH_magic_2.B.n51 0.237239
R3622 TG_GATE_SWITCH_magic_2.B.n107 TG_GATE_SWITCH_magic_2.B.n106 0.2033
R3623 TG_GATE_SWITCH_magic_2.B.n106 TG_GATE_SWITCH_magic_2.B.n71 0.136437
R3624 TG_GATE_SWITCH_magic_2.B TG_GATE_SWITCH_magic_2.B.n107 0.0845
R3625 A5.n47 A5.n46 5.44589
R3626 A5.n24 A5.n22 5.07789
R3627 A5.n50 A5.t29 4.7885
R3628 A5.n51 A5.t27 4.7885
R3629 A5.n47 A5.n45 4.7885
R3630 A5.n34 A5.t22 4.4205
R3631 A5.n33 A5.t14 4.4205
R3632 A5.n32 A5.t3 4.4205
R3633 A5.n31 A5.t0 4.4205
R3634 A5.n28 A5.n27 4.4205
R3635 A5.n26 A5.n25 4.4205
R3636 A5.n24 A5.n23 4.4205
R3637 A5.n39 A5.n38 3.80789
R3638 A5.n44 A5.n43 3.80789
R3639 A5.n15 A5.n12 3.25789
R3640 A5.n4 A5.n1 3.25789
R3641 A5.n39 A5.n36 3.1505
R3642 A5.n44 A5.n41 3.1505
R3643 A5.n15 A5.n14 2.6005
R3644 A5.n18 A5.n17 2.6005
R3645 A5.n21 A5.n20 2.6005
R3646 A5.n4 A5.n3 2.6005
R3647 A5.n7 A5.n6 2.6005
R3648 A5.n10 A5.n9 2.6005
R3649 A5.n20 A5.t13 1.8205
R3650 A5.n20 A5.n19 1.8205
R3651 A5.n17 A5.t16 1.8205
R3652 A5.n17 A5.n16 1.8205
R3653 A5.n14 A5.t21 1.8205
R3654 A5.n14 A5.n13 1.8205
R3655 A5.n12 A5.t11 1.8205
R3656 A5.n12 A5.n11 1.8205
R3657 A5.n9 A5.t6 1.8205
R3658 A5.n9 A5.n8 1.8205
R3659 A5.n6 A5.t10 1.8205
R3660 A5.n6 A5.n5 1.8205
R3661 A5.n3 A5.t17 1.8205
R3662 A5.n3 A5.n2 1.8205
R3663 A5.n1 A5.t4 1.8205
R3664 A5.n1 A5.n0 1.8205
R3665 A5.n36 A5.t33 1.6385
R3666 A5.n36 A5.n35 1.6385
R3667 A5.n38 A5.t31 1.6385
R3668 A5.n38 A5.n37 1.6385
R3669 A5.n41 A5.t24 1.6385
R3670 A5.n41 A5.n40 1.6385
R3671 A5.n43 A5.t35 1.6385
R3672 A5.n43 A5.n42 1.6385
R3673 A5 A5.n52 1.54838
R3674 A5.n48 A5.n47 0.884196
R3675 A5.n50 A5.n49 0.884196
R3676 A5.n29 A5.n28 0.882239
R3677 A5.n31 A5.n30 0.882239
R3678 A5.n51 A5.n50 0.657891
R3679 A5.n26 A5.n24 0.657891
R3680 A5.n28 A5.n26 0.657891
R3681 A5.n18 A5.n15 0.657891
R3682 A5.n21 A5.n18 0.657891
R3683 A5.n7 A5.n4 0.657891
R3684 A5.n10 A5.n7 0.657891
R3685 A5.n34 A5.n33 0.657891
R3686 A5.n33 A5.n32 0.657891
R3687 A5.n32 A5.n31 0.657891
R3688 A5.n49 A5.n48 0.6005
R3689 A5.n30 A5.n29 0.6005
R3690 A5.n52 A5.n51 0.60042
R3691 A5.n49 A5.n39 0.284196
R3692 A5.n48 A5.n44 0.284196
R3693 A5.n29 A5.n21 0.282239
R3694 A5.n30 A5.n10 0.282239
R3695 A5.n52 A5.n34 0.277389
R3696 S1.n1 S1.t48 68.1773
R3697 S1.n20 S1.t2 68.1773
R3698 S1.n11 S1.n10 52.5344
R3699 S1.n24 S1.n23 52.5344
R3700 S1.n12 S1.t16 47.0594
R3701 S1.n25 S1.t5 47.0594
R3702 S1.t40 S1.t3 43.8005
R3703 S1.t25 S1.t40 43.8005
R3704 S1.t16 S1.t25 43.8005
R3705 S1.t30 S1.t6 43.8005
R3706 S1.t44 S1.t30 43.8005
R3707 S1.t5 S1.t44 43.8005
R3708 S1.t13 S1.t19 43.8005
R3709 S1.t21 S1.t33 43.8005
R3710 S1.t35 S1.t47 43.8005
R3711 S1.t11 S1.t17 43.8005
R3712 S1.n5 S1.t32 33.8934
R3713 S1.n17 S1.t49 33.763
R3714 S1.t26 S1.t36 30.7648
R3715 S1.t27 S1.t38 30.7648
R3716 S1.t41 S1.t50 30.7648
R3717 S1.t0 S1.t9 30.7648
R3718 S1.n27 S1.t27 30.3737
R3719 S1.n28 S1.t41 30.3737
R3720 S1.n29 S1.t0 30.3737
R3721 S1.t32 S1.n4 21.9005
R3722 S1.n4 S1.t45 21.9005
R3723 S1.n3 S1.t28 21.9005
R3724 S1.n3 S1.t42 21.9005
R3725 S1.n2 S1.t34 21.9005
R3726 S1.n2 S1.t46 21.9005
R3727 S1.t29 S1.n0 21.9005
R3728 S1.n0 S1.t43 21.9005
R3729 S1.n9 S1.t23 21.9005
R3730 S1.n9 S1.t15 21.9005
R3731 S1.n16 S1.t18 21.9005
R3732 S1.t49 S1.n16 21.9005
R3733 S1.n15 S1.t31 21.9005
R3734 S1.n15 S1.t8 21.9005
R3735 S1.n14 S1.t51 21.9005
R3736 S1.n14 S1.t20 21.9005
R3737 S1.n13 S1.t22 21.9005
R3738 S1.t1 S1.n13 21.9005
R3739 S1.n22 S1.t37 21.9005
R3740 S1.n22 S1.t10 21.9005
R3741 S1.n27 S1.t13 21.6398
R3742 S1.n28 S1.t21 21.6398
R3743 S1.n29 S1.t35 21.6398
R3744 S1.n30 S1.t11 21.6398
R3745 S1.n8 S1.n1 20.8576
R3746 S1.n8 S1.n7 20.8576
R3747 S1.n7 S1.n6 20.8576
R3748 S1.n6 S1.n5 20.8576
R3749 S1.n18 S1.n17 20.8576
R3750 S1.n19 S1.n18 20.8576
R3751 S1.n21 S1.n19 20.8576
R3752 S1.n21 S1.n20 20.8576
R3753 S1.n10 S1.n9 19.4672
R3754 S1.n23 S1.n22 19.4672
R3755 S1.n12 S1.t7 19.4237
R3756 S1.n25 S1.t24 19.4237
R3757 S1.n10 S1.t12 18.2505
R3758 S1.n11 S1.t48 18.2505
R3759 S1.n10 S1.t4 18.2505
R3760 S1.t7 S1.n11 18.2505
R3761 S1.n24 S1.t2 18.2505
R3762 S1.n23 S1.t39 18.2505
R3763 S1.n23 S1.t14 18.2505
R3764 S1.t24 S1.n24 18.2505
R3765 S1.n31 S1.t26 17.8543
R3766 S1.n28 S1.n27 17.255
R3767 S1.n29 S1.n28 17.255
R3768 S1.n30 S1.n29 17.255
R3769 S1.n4 S1.n3 15.8172
R3770 S1.n3 S1.n2 15.8172
R3771 S1.n2 S1.n0 15.8172
R3772 S1.n9 S1.n0 15.8172
R3773 S1.n16 S1.n15 15.8172
R3774 S1.n15 S1.n14 15.8172
R3775 S1.n14 S1.n13 15.8172
R3776 S1.n22 S1.n13 15.8172
R3777 S1.n5 S1.t28 15.6434
R3778 S1.n6 S1.t34 15.6434
R3779 S1.n7 S1.t29 15.6434
R3780 S1.t15 S1.n8 15.6434
R3781 S1.n1 S1.t4 15.6434
R3782 S1.n17 S1.t8 15.6434
R3783 S1.n18 S1.t20 15.6434
R3784 S1.n19 S1.t1 15.6434
R3785 S1.t10 S1.n21 15.6434
R3786 S1.n20 S1.t39 15.6434
R3787 S1.n26 S1 10.5832
R3788 S1 S1.n25 8.63236
R3789 S1 S1.n12 8.62829
R3790 S1.n31 S1.n30 7.99318
R3791 S1.n26 S1 5.35201
R3792 S1 S1.n31 4.24427
R3793 S1.n32 S1.n26 2.93261
R3794 S1.n34 S1.n33 2.37219
R3795 S1 S1.n34 2.28599
R3796 S1.n32 S1 1.23201
R3797 S1.n33 S1.n32 0.303526
R3798 S1 S1.n33 0.12219
R3799 A4.n47 A4.n46 5.44589
R3800 A4.n24 A4.n22 5.07789
R3801 A4.n50 A4.t17 4.7885
R3802 A4.n51 A4.t20 4.7885
R3803 A4.n47 A4.n45 4.7885
R3804 A4.n34 A4.t5 4.4205
R3805 A4.n33 A4.t9 4.4205
R3806 A4.n32 A4.t14 4.4205
R3807 A4.n31 A4.t3 4.4205
R3808 A4.n28 A4.n27 4.4205
R3809 A4.n26 A4.n25 4.4205
R3810 A4.n24 A4.n23 4.4205
R3811 A4.n39 A4.n38 3.80789
R3812 A4.n44 A4.n43 3.80789
R3813 A4.n15 A4.n12 3.25789
R3814 A4.n4 A4.n1 3.25789
R3815 A4.n39 A4.n36 3.1505
R3816 A4.n44 A4.n41 3.1505
R3817 A4.n53 A4 3.10602
R3818 A4.n15 A4.n14 2.6005
R3819 A4.n18 A4.n17 2.6005
R3820 A4.n21 A4.n20 2.6005
R3821 A4.n4 A4.n3 2.6005
R3822 A4.n7 A4.n6 2.6005
R3823 A4.n10 A4.n9 2.6005
R3824 A4.n20 A4.t27 1.8205
R3825 A4.n20 A4.n19 1.8205
R3826 A4.n17 A4.t4 1.8205
R3827 A4.n17 A4.n16 1.8205
R3828 A4.n14 A4.t31 1.8205
R3829 A4.n14 A4.n13 1.8205
R3830 A4.n12 A4.t28 1.8205
R3831 A4.n12 A4.n11 1.8205
R3832 A4.n9 A4.t32 1.8205
R3833 A4.n9 A4.n8 1.8205
R3834 A4.n6 A4.t10 1.8205
R3835 A4.n6 A4.n5 1.8205
R3836 A4.n3 A4.t1 1.8205
R3837 A4.n3 A4.n2 1.8205
R3838 A4.n1 A4.t34 1.8205
R3839 A4.n1 A4.n0 1.8205
R3840 A4.n36 A4.t15 1.6385
R3841 A4.n36 A4.n35 1.6385
R3842 A4.n38 A4.t18 1.6385
R3843 A4.n38 A4.n37 1.6385
R3844 A4.n41 A4.t19 1.6385
R3845 A4.n41 A4.n40 1.6385
R3846 A4.n43 A4.t16 1.6385
R3847 A4.n43 A4.n42 1.6385
R3848 A4.n53 A4.n52 1.35968
R3849 A4.n48 A4.n47 0.884196
R3850 A4.n50 A4.n49 0.884196
R3851 A4.n29 A4.n28 0.882239
R3852 A4.n31 A4.n30 0.882239
R3853 A4.n51 A4.n50 0.657891
R3854 A4.n26 A4.n24 0.657891
R3855 A4.n28 A4.n26 0.657891
R3856 A4.n18 A4.n15 0.657891
R3857 A4.n21 A4.n18 0.657891
R3858 A4.n7 A4.n4 0.657891
R3859 A4.n10 A4.n7 0.657891
R3860 A4.n34 A4.n33 0.657891
R3861 A4.n33 A4.n32 0.657891
R3862 A4.n32 A4.n31 0.657891
R3863 A4.n49 A4.n48 0.6005
R3864 A4.n30 A4.n29 0.6005
R3865 A4.n52 A4.n51 0.60042
R3866 A4.n49 A4.n39 0.284196
R3867 A4.n48 A4.n44 0.284196
R3868 A4.n29 A4.n21 0.282239
R3869 A4.n30 A4.n10 0.282239
R3870 A4.n52 A4.n34 0.277389
R3871 A4 A4.n53 0.189193
R3872 TG_GATE_SWITCH_magic_6.B.n48 TG_GATE_SWITCH_magic_6.B.n46 5.44589
R3873 TG_GATE_SWITCH_magic_6.B.n27 TG_GATE_SWITCH_magic_6.B.n26 5.07789
R3874 TG_GATE_SWITCH_magic_6.B.n52 TG_GATE_SWITCH_magic_6.B.t69 4.7885
R3875 TG_GATE_SWITCH_magic_6.B.n51 TG_GATE_SWITCH_magic_6.B.t29 4.7885
R3876 TG_GATE_SWITCH_magic_6.B.n48 TG_GATE_SWITCH_magic_6.B.n47 4.7885
R3877 TG_GATE_SWITCH_magic_6.B.n32 TG_GATE_SWITCH_magic_6.B.t15 4.4205
R3878 TG_GATE_SWITCH_magic_6.B.n33 TG_GATE_SWITCH_magic_6.B.t9 4.4205
R3879 TG_GATE_SWITCH_magic_6.B.n34 TG_GATE_SWITCH_magic_6.B.t5 4.4205
R3880 TG_GATE_SWITCH_magic_6.B.n35 TG_GATE_SWITCH_magic_6.B.t17 4.4205
R3881 TG_GATE_SWITCH_magic_6.B.n29 TG_GATE_SWITCH_magic_6.B.n23 4.4205
R3882 TG_GATE_SWITCH_magic_6.B.n28 TG_GATE_SWITCH_magic_6.B.n24 4.4205
R3883 TG_GATE_SWITCH_magic_6.B.n27 TG_GATE_SWITCH_magic_6.B.n25 4.4205
R3884 TG_GATE_SWITCH_magic_6.B.n83 TG_GATE_SWITCH_magic_6.B.n80 3.80789
R3885 TG_GATE_SWITCH_magic_6.B.n88 TG_GATE_SWITCH_magic_6.B.n85 3.80789
R3886 TG_GATE_SWITCH_magic_6.B.n45 TG_GATE_SWITCH_magic_6.B.n42 3.80789
R3887 TG_GATE_SWITCH_magic_6.B.n40 TG_GATE_SWITCH_magic_6.B.n37 3.80789
R3888 TG_GATE_SWITCH_magic_6.B.n93 TG_GATE_SWITCH_magic_6.B.n90 3.80789
R3889 TG_GATE_SWITCH_magic_6.B.n9 TG_GATE_SWITCH_magic_6.B.n8 3.25789
R3890 TG_GATE_SWITCH_magic_6.B.n20 TG_GATE_SWITCH_magic_6.B.n19 3.25789
R3891 TG_GATE_SWITCH_magic_6.B.n75 TG_GATE_SWITCH_magic_6.B.n74 3.25789
R3892 TG_GATE_SWITCH_magic_6.B.n64 TG_GATE_SWITCH_magic_6.B.n63 3.25789
R3893 TG_GATE_SWITCH_magic_6.B.n104 TG_GATE_SWITCH_magic_6.B.n103 3.25789
R3894 TG_GATE_SWITCH_magic_6.B.n55 TG_GATE_SWITCH_magic_6.B.n54 3.21114
R3895 TG_GATE_SWITCH_magic_6.B.n83 TG_GATE_SWITCH_magic_6.B.n82 3.1505
R3896 TG_GATE_SWITCH_magic_6.B.n88 TG_GATE_SWITCH_magic_6.B.n87 3.1505
R3897 TG_GATE_SWITCH_magic_6.B.n45 TG_GATE_SWITCH_magic_6.B.n44 3.1505
R3898 TG_GATE_SWITCH_magic_6.B.n40 TG_GATE_SWITCH_magic_6.B.n39 3.1505
R3899 TG_GATE_SWITCH_magic_6.B.n93 TG_GATE_SWITCH_magic_6.B.n92 3.1505
R3900 TG_GATE_SWITCH_magic_6.B.n9 TG_GATE_SWITCH_magic_6.B.n6 2.6005
R3901 TG_GATE_SWITCH_magic_6.B.n10 TG_GATE_SWITCH_magic_6.B.n4 2.6005
R3902 TG_GATE_SWITCH_magic_6.B.n11 TG_GATE_SWITCH_magic_6.B.n2 2.6005
R3903 TG_GATE_SWITCH_magic_6.B.n20 TG_GATE_SWITCH_magic_6.B.n17 2.6005
R3904 TG_GATE_SWITCH_magic_6.B.n21 TG_GATE_SWITCH_magic_6.B.n15 2.6005
R3905 TG_GATE_SWITCH_magic_6.B.n22 TG_GATE_SWITCH_magic_6.B.n13 2.6005
R3906 TG_GATE_SWITCH_magic_6.B.n75 TG_GATE_SWITCH_magic_6.B.n72 2.6005
R3907 TG_GATE_SWITCH_magic_6.B.n76 TG_GATE_SWITCH_magic_6.B.n70 2.6005
R3908 TG_GATE_SWITCH_magic_6.B.n77 TG_GATE_SWITCH_magic_6.B.n68 2.6005
R3909 TG_GATE_SWITCH_magic_6.B.n64 TG_GATE_SWITCH_magic_6.B.n61 2.6005
R3910 TG_GATE_SWITCH_magic_6.B.n65 TG_GATE_SWITCH_magic_6.B.n59 2.6005
R3911 TG_GATE_SWITCH_magic_6.B.n66 TG_GATE_SWITCH_magic_6.B.n57 2.6005
R3912 TG_GATE_SWITCH_magic_6.B.n104 TG_GATE_SWITCH_magic_6.B.n101 2.6005
R3913 TG_GATE_SWITCH_magic_6.B.n105 TG_GATE_SWITCH_magic_6.B.n99 2.6005
R3914 TG_GATE_SWITCH_magic_6.B.n106 TG_GATE_SWITCH_magic_6.B.n97 2.6005
R3915 TG_GATE_SWITCH_magic_6.B.n108 TG_GATE_SWITCH_magic_6.B.n55 2.32083
R3916 TG_GATE_SWITCH_magic_6.B.n54 TG_GATE_SWITCH_magic_6.B.n0 2.25155
R3917 TG_GATE_SWITCH_magic_6.B.n2 TG_GATE_SWITCH_magic_6.B.t7 1.8205
R3918 TG_GATE_SWITCH_magic_6.B.n2 TG_GATE_SWITCH_magic_6.B.n1 1.8205
R3919 TG_GATE_SWITCH_magic_6.B.n4 TG_GATE_SWITCH_magic_6.B.t2 1.8205
R3920 TG_GATE_SWITCH_magic_6.B.n4 TG_GATE_SWITCH_magic_6.B.n3 1.8205
R3921 TG_GATE_SWITCH_magic_6.B.n6 TG_GATE_SWITCH_magic_6.B.t21 1.8205
R3922 TG_GATE_SWITCH_magic_6.B.n6 TG_GATE_SWITCH_magic_6.B.n5 1.8205
R3923 TG_GATE_SWITCH_magic_6.B.n8 TG_GATE_SWITCH_magic_6.B.t8 1.8205
R3924 TG_GATE_SWITCH_magic_6.B.n8 TG_GATE_SWITCH_magic_6.B.n7 1.8205
R3925 TG_GATE_SWITCH_magic_6.B.n13 TG_GATE_SWITCH_magic_6.B.t30 1.8205
R3926 TG_GATE_SWITCH_magic_6.B.n13 TG_GATE_SWITCH_magic_6.B.n12 1.8205
R3927 TG_GATE_SWITCH_magic_6.B.n15 TG_GATE_SWITCH_magic_6.B.t16 1.8205
R3928 TG_GATE_SWITCH_magic_6.B.n15 TG_GATE_SWITCH_magic_6.B.n14 1.8205
R3929 TG_GATE_SWITCH_magic_6.B.n17 TG_GATE_SWITCH_magic_6.B.t13 1.8205
R3930 TG_GATE_SWITCH_magic_6.B.n17 TG_GATE_SWITCH_magic_6.B.n16 1.8205
R3931 TG_GATE_SWITCH_magic_6.B.n19 TG_GATE_SWITCH_magic_6.B.t23 1.8205
R3932 TG_GATE_SWITCH_magic_6.B.n19 TG_GATE_SWITCH_magic_6.B.n18 1.8205
R3933 TG_GATE_SWITCH_magic_6.B.n68 TG_GATE_SWITCH_magic_6.B.t43 1.8205
R3934 TG_GATE_SWITCH_magic_6.B.n68 TG_GATE_SWITCH_magic_6.B.n67 1.8205
R3935 TG_GATE_SWITCH_magic_6.B.n70 TG_GATE_SWITCH_magic_6.B.t44 1.8205
R3936 TG_GATE_SWITCH_magic_6.B.n70 TG_GATE_SWITCH_magic_6.B.n69 1.8205
R3937 TG_GATE_SWITCH_magic_6.B.n72 TG_GATE_SWITCH_magic_6.B.t61 1.8205
R3938 TG_GATE_SWITCH_magic_6.B.n72 TG_GATE_SWITCH_magic_6.B.n71 1.8205
R3939 TG_GATE_SWITCH_magic_6.B.n74 TG_GATE_SWITCH_magic_6.B.t40 1.8205
R3940 TG_GATE_SWITCH_magic_6.B.n74 TG_GATE_SWITCH_magic_6.B.n73 1.8205
R3941 TG_GATE_SWITCH_magic_6.B.n57 TG_GATE_SWITCH_magic_6.B.t34 1.8205
R3942 TG_GATE_SWITCH_magic_6.B.n57 TG_GATE_SWITCH_magic_6.B.n56 1.8205
R3943 TG_GATE_SWITCH_magic_6.B.n59 TG_GATE_SWITCH_magic_6.B.t38 1.8205
R3944 TG_GATE_SWITCH_magic_6.B.n59 TG_GATE_SWITCH_magic_6.B.n58 1.8205
R3945 TG_GATE_SWITCH_magic_6.B.n61 TG_GATE_SWITCH_magic_6.B.t45 1.8205
R3946 TG_GATE_SWITCH_magic_6.B.n61 TG_GATE_SWITCH_magic_6.B.n60 1.8205
R3947 TG_GATE_SWITCH_magic_6.B.n63 TG_GATE_SWITCH_magic_6.B.t32 1.8205
R3948 TG_GATE_SWITCH_magic_6.B.n63 TG_GATE_SWITCH_magic_6.B.n62 1.8205
R3949 TG_GATE_SWITCH_magic_6.B.n97 TG_GATE_SWITCH_magic_6.B.t65 1.8205
R3950 TG_GATE_SWITCH_magic_6.B.n97 TG_GATE_SWITCH_magic_6.B.n96 1.8205
R3951 TG_GATE_SWITCH_magic_6.B.n99 TG_GATE_SWITCH_magic_6.B.t67 1.8205
R3952 TG_GATE_SWITCH_magic_6.B.n99 TG_GATE_SWITCH_magic_6.B.n98 1.8205
R3953 TG_GATE_SWITCH_magic_6.B.n101 TG_GATE_SWITCH_magic_6.B.t39 1.8205
R3954 TG_GATE_SWITCH_magic_6.B.n101 TG_GATE_SWITCH_magic_6.B.n100 1.8205
R3955 TG_GATE_SWITCH_magic_6.B.n103 TG_GATE_SWITCH_magic_6.B.t62 1.8205
R3956 TG_GATE_SWITCH_magic_6.B.n103 TG_GATE_SWITCH_magic_6.B.n102 1.8205
R3957 TG_GATE_SWITCH_magic_6.B.n90 TG_GATE_SWITCH_magic_6.B.t49 1.6385
R3958 TG_GATE_SWITCH_magic_6.B.n90 TG_GATE_SWITCH_magic_6.B.n89 1.6385
R3959 TG_GATE_SWITCH_magic_6.B.n82 TG_GATE_SWITCH_magic_6.B.t47 1.6385
R3960 TG_GATE_SWITCH_magic_6.B.n82 TG_GATE_SWITCH_magic_6.B.n81 1.6385
R3961 TG_GATE_SWITCH_magic_6.B.n80 TG_GATE_SWITCH_magic_6.B.t53 1.6385
R3962 TG_GATE_SWITCH_magic_6.B.n80 TG_GATE_SWITCH_magic_6.B.n79 1.6385
R3963 TG_GATE_SWITCH_magic_6.B.n87 TG_GATE_SWITCH_magic_6.B.t50 1.6385
R3964 TG_GATE_SWITCH_magic_6.B.n87 TG_GATE_SWITCH_magic_6.B.n86 1.6385
R3965 TG_GATE_SWITCH_magic_6.B.n85 TG_GATE_SWITCH_magic_6.B.t56 1.6385
R3966 TG_GATE_SWITCH_magic_6.B.n85 TG_GATE_SWITCH_magic_6.B.n84 1.6385
R3967 TG_GATE_SWITCH_magic_6.B.n44 TG_GATE_SWITCH_magic_6.B.t0 1.6385
R3968 TG_GATE_SWITCH_magic_6.B.n44 TG_GATE_SWITCH_magic_6.B.n43 1.6385
R3969 TG_GATE_SWITCH_magic_6.B.n42 TG_GATE_SWITCH_magic_6.B.t27 1.6385
R3970 TG_GATE_SWITCH_magic_6.B.n42 TG_GATE_SWITCH_magic_6.B.n41 1.6385
R3971 TG_GATE_SWITCH_magic_6.B.n39 TG_GATE_SWITCH_magic_6.B.t71 1.6385
R3972 TG_GATE_SWITCH_magic_6.B.n39 TG_GATE_SWITCH_magic_6.B.n38 1.6385
R3973 TG_GATE_SWITCH_magic_6.B.n37 TG_GATE_SWITCH_magic_6.B.t24 1.6385
R3974 TG_GATE_SWITCH_magic_6.B.n37 TG_GATE_SWITCH_magic_6.B.n36 1.6385
R3975 TG_GATE_SWITCH_magic_6.B.n92 TG_GATE_SWITCH_magic_6.B.t55 1.6385
R3976 TG_GATE_SWITCH_magic_6.B.n92 TG_GATE_SWITCH_magic_6.B.n91 1.6385
R3977 TG_GATE_SWITCH_magic_6.B.n54 TG_GATE_SWITCH_magic_6.B.n53 1.51805
R3978 TG_GATE_SWITCH_magic_6.B.n49 TG_GATE_SWITCH_magic_6.B.n48 0.884196
R3979 TG_GATE_SWITCH_magic_6.B.n51 TG_GATE_SWITCH_magic_6.B.n50 0.884196
R3980 TG_GATE_SWITCH_magic_6.B.n30 TG_GATE_SWITCH_magic_6.B.n29 0.882239
R3981 TG_GATE_SWITCH_magic_6.B.n32 TG_GATE_SWITCH_magic_6.B.n31 0.882239
R3982 TG_GATE_SWITCH_magic_6.B.n53 TG_GATE_SWITCH_magic_6.B.n52 0.8105
R3983 TG_GATE_SWITCH_magic_6.B.n11 TG_GATE_SWITCH_magic_6.B.n10 0.657891
R3984 TG_GATE_SWITCH_magic_6.B.n10 TG_GATE_SWITCH_magic_6.B.n9 0.657891
R3985 TG_GATE_SWITCH_magic_6.B.n22 TG_GATE_SWITCH_magic_6.B.n21 0.657891
R3986 TG_GATE_SWITCH_magic_6.B.n21 TG_GATE_SWITCH_magic_6.B.n20 0.657891
R3987 TG_GATE_SWITCH_magic_6.B.n29 TG_GATE_SWITCH_magic_6.B.n28 0.657891
R3988 TG_GATE_SWITCH_magic_6.B.n28 TG_GATE_SWITCH_magic_6.B.n27 0.657891
R3989 TG_GATE_SWITCH_magic_6.B.n33 TG_GATE_SWITCH_magic_6.B.n32 0.657891
R3990 TG_GATE_SWITCH_magic_6.B.n34 TG_GATE_SWITCH_magic_6.B.n33 0.657891
R3991 TG_GATE_SWITCH_magic_6.B.n35 TG_GATE_SWITCH_magic_6.B.n34 0.657891
R3992 TG_GATE_SWITCH_magic_6.B.n52 TG_GATE_SWITCH_magic_6.B.n51 0.657891
R3993 TG_GATE_SWITCH_magic_6.B.n76 TG_GATE_SWITCH_magic_6.B.n75 0.657891
R3994 TG_GATE_SWITCH_magic_6.B.n66 TG_GATE_SWITCH_magic_6.B.n65 0.657891
R3995 TG_GATE_SWITCH_magic_6.B.n65 TG_GATE_SWITCH_magic_6.B.n64 0.657891
R3996 TG_GATE_SWITCH_magic_6.B.n106 TG_GATE_SWITCH_magic_6.B.n105 0.657891
R3997 TG_GATE_SWITCH_magic_6.B.n105 TG_GATE_SWITCH_magic_6.B.n104 0.657891
R3998 TG_GATE_SWITCH_magic_6.B.n77 TG_GATE_SWITCH_magic_6.B.n76 0.655976
R3999 TG_GATE_SWITCH_magic_6.B.n78 TG_GATE_SWITCH_magic_6.B.n77 0.645657
R4000 TG_GATE_SWITCH_magic_6.B.n50 TG_GATE_SWITCH_magic_6.B.n49 0.6005
R4001 TG_GATE_SWITCH_magic_6.B.n31 TG_GATE_SWITCH_magic_6.B.n30 0.6005
R4002 TG_GATE_SWITCH_magic_6.B.n94 TG_GATE_SWITCH_magic_6.B.n93 0.548416
R4003 TG_GATE_SWITCH_magic_6.B.n107 TG_GATE_SWITCH_magic_6.B.n106 0.316429
R4004 TG_GATE_SWITCH_magic_6.B.n95 TG_GATE_SWITCH_magic_6.B.n83 0.304838
R4005 TG_GATE_SWITCH_magic_6.B.n94 TG_GATE_SWITCH_magic_6.B.n88 0.284196
R4006 TG_GATE_SWITCH_magic_6.B.n49 TG_GATE_SWITCH_magic_6.B.n45 0.284196
R4007 TG_GATE_SWITCH_magic_6.B.n50 TG_GATE_SWITCH_magic_6.B.n40 0.284196
R4008 TG_GATE_SWITCH_magic_6.B.n107 TG_GATE_SWITCH_magic_6.B.n78 0.283032
R4009 TG_GATE_SWITCH_magic_6.B.n31 TG_GATE_SWITCH_magic_6.B.n11 0.282239
R4010 TG_GATE_SWITCH_magic_6.B.n30 TG_GATE_SWITCH_magic_6.B.n22 0.282239
R4011 TG_GATE_SWITCH_magic_6.B.n78 TG_GATE_SWITCH_magic_6.B.n66 0.279866
R4012 TG_GATE_SWITCH_magic_6.B.n95 TG_GATE_SWITCH_magic_6.B.n94 0.244078
R4013 TG_GATE_SWITCH_magic_6.B.n53 TG_GATE_SWITCH_magic_6.B.n35 0.237239
R4014 TG_GATE_SWITCH_magic_6.B.n108 TG_GATE_SWITCH_magic_6.B.n107 0.2201
R4015 TG_GATE_SWITCH_magic_6.B.n107 TG_GATE_SWITCH_magic_6.B.n95 0.136437
R4016 TG_GATE_SWITCH_magic_6.B TG_GATE_SWITCH_magic_6.B.n108 0.0677
R4017 TG_GATE_SWITCH_magic_6.B.n0 TG_GATE_SWITCH_magic_6.B 0.0244241
R4018 a_2061_n2270.t17 a_2061_n2270.n19 40.7345
R4019 a_2061_n2270.n24 a_2061_n2270.n5 28.094
R4020 a_2061_n2270.n21 a_2061_n2270.n20 28.094
R4021 a_2061_n2270.n32 a_2061_n2270.n31 28.094
R4022 a_2061_n2270.n26 a_2061_n2270.t13 21.9005
R4023 a_2061_n2270.n26 a_2061_n2270.t7 21.9005
R4024 a_2061_n2270.n0 a_2061_n2270.t24 21.9005
R4025 a_2061_n2270.n11 a_2061_n2270.t21 21.9005
R4026 a_2061_n2270.n12 a_2061_n2270.t25 21.9005
R4027 a_2061_n2270.n1 a_2061_n2270.t6 21.9005
R4028 a_2061_n2270.n27 a_2061_n2270.t12 21.9005
R4029 a_2061_n2270.n27 a_2061_n2270.t18 21.9005
R4030 a_2061_n2270.n28 a_2061_n2270.t26 21.9005
R4031 a_2061_n2270.n28 a_2061_n2270.t20 21.9005
R4032 a_2061_n2270.n2 a_2061_n2270.t14 21.9005
R4033 a_2061_n2270.n13 a_2061_n2270.t11 21.9005
R4034 a_2061_n2270.n14 a_2061_n2270.t23 21.9005
R4035 a_2061_n2270.n3 a_2061_n2270.t27 21.9005
R4036 a_2061_n2270.n29 a_2061_n2270.t9 21.9005
R4037 a_2061_n2270.n29 a_2061_n2270.t16 21.9005
R4038 a_2061_n2270.n30 a_2061_n2270.t19 21.9005
R4039 a_2061_n2270.n30 a_2061_n2270.t15 21.9005
R4040 a_2061_n2270.n4 a_2061_n2270.t8 21.9005
R4041 a_2061_n2270.n15 a_2061_n2270.t29 21.9005
R4042 a_2061_n2270.n20 a_2061_n2270.t17 21.9005
R4043 a_2061_n2270.n5 a_2061_n2270.t22 21.9005
R4044 a_2061_n2270.n31 a_2061_n2270.t28 21.9005
R4045 a_2061_n2270.n31 a_2061_n2270.t10 21.9005
R4046 a_2061_n2270.n20 a_2061_n2270.n15 15.8172
R4047 a_2061_n2270.n5 a_2061_n2270.n4 15.8172
R4048 a_2061_n2270.n4 a_2061_n2270.n3 15.8172
R4049 a_2061_n2270.n15 a_2061_n2270.n14 15.8172
R4050 a_2061_n2270.n14 a_2061_n2270.n13 15.8172
R4051 a_2061_n2270.n3 a_2061_n2270.n2 15.8172
R4052 a_2061_n2270.n2 a_2061_n2270.n1 15.8172
R4053 a_2061_n2270.n13 a_2061_n2270.n12 15.8172
R4054 a_2061_n2270.n12 a_2061_n2270.n11 15.8172
R4055 a_2061_n2270.n1 a_2061_n2270.n0 15.8172
R4056 a_2061_n2270.n27 a_2061_n2270.n26 15.8172
R4057 a_2061_n2270.n29 a_2061_n2270.n28 15.8172
R4058 a_2061_n2270.n28 a_2061_n2270.n27 15.8172
R4059 a_2061_n2270.n31 a_2061_n2270.n30 15.8172
R4060 a_2061_n2270.n30 a_2061_n2270.n29 15.8172
R4061 a_2061_n2270.n17 a_2061_n2270.n16 15.1845
R4062 a_2061_n2270.n19 a_2061_n2270.n18 15.1845
R4063 a_2061_n2270.n18 a_2061_n2270.n17 15.1845
R4064 a_2061_n2270.n8 a_2061_n2270.n6 5.44589
R4065 a_2061_n2270.n8 a_2061_n2270.n7 4.7885
R4066 a_2061_n2270.n32 a_2061_n2270.n25 4.70615
R4067 a_2061_n2270.n23 a_2061_n2270.n22 4.4205
R4068 a_2061_n2270.n10 a_2061_n2270.n9 4.4205
R4069 a_2061_n2270.n34 a_2061_n2270.n33 4.4205
R4070 a_2061_n2270.n10 a_2061_n2270.n8 1.1392
R4071 a_2061_n2270.n23 a_2061_n2270.n21 0.286152
R4072 a_2061_n2270.n33 a_2061_n2270.n24 0.286152
R4073 a_2061_n2270.n21 a_2061_n2270.n10 0.282239
R4074 a_2061_n2270.n24 a_2061_n2270.n23 0.282239
R4075 a_2061_n2270.n33 a_2061_n2270.n32 0.282239
R4076 a_5684_1104.t17 a_5684_1104.n17 40.7345
R4077 a_5684_1104.n19 a_5684_1104.n18 28.094
R4078 a_5684_1104.n6 a_5684_1104.n5 28.094
R4079 a_5684_1104.n27 a_5684_1104.n26 28.094
R4080 a_5684_1104.n5 a_5684_1104.t15 21.9005
R4081 a_5684_1104.n5 a_5684_1104.t10 21.9005
R4082 a_5684_1104.n3 a_5684_1104.t25 21.9005
R4083 a_5684_1104.n1 a_5684_1104.t24 21.9005
R4084 a_5684_1104.n0 a_5684_1104.t8 21.9005
R4085 a_5684_1104.n0 a_5684_1104.t23 21.9005
R4086 a_5684_1104.n21 a_5684_1104.t22 21.9005
R4087 a_5684_1104.n9 a_5684_1104.t9 21.9005
R4088 a_5684_1104.n10 a_5684_1104.t26 21.9005
R4089 a_5684_1104.n22 a_5684_1104.t12 21.9005
R4090 a_5684_1104.n1 a_5684_1104.t16 21.9005
R4091 a_5684_1104.n2 a_5684_1104.t28 21.9005
R4092 a_5684_1104.n2 a_5684_1104.t21 21.9005
R4093 a_5684_1104.n23 a_5684_1104.t14 21.9005
R4094 a_5684_1104.n11 a_5684_1104.t29 21.9005
R4095 a_5684_1104.n12 a_5684_1104.t27 21.9005
R4096 a_5684_1104.n24 a_5684_1104.t13 21.9005
R4097 a_5684_1104.n3 a_5684_1104.t18 21.9005
R4098 a_5684_1104.n4 a_5684_1104.t19 21.9005
R4099 a_5684_1104.n4 a_5684_1104.t11 21.9005
R4100 a_5684_1104.n25 a_5684_1104.t7 21.9005
R4101 a_5684_1104.n13 a_5684_1104.t20 21.9005
R4102 a_5684_1104.n18 a_5684_1104.t17 21.9005
R4103 a_5684_1104.n26 a_5684_1104.t6 21.9005
R4104 a_5684_1104.n18 a_5684_1104.n13 15.8172
R4105 a_5684_1104.n26 a_5684_1104.n25 15.8172
R4106 a_5684_1104.n25 a_5684_1104.n24 15.8172
R4107 a_5684_1104.n13 a_5684_1104.n12 15.8172
R4108 a_5684_1104.n12 a_5684_1104.n11 15.8172
R4109 a_5684_1104.n24 a_5684_1104.n23 15.8172
R4110 a_5684_1104.n23 a_5684_1104.n22 15.8172
R4111 a_5684_1104.n11 a_5684_1104.n10 15.8172
R4112 a_5684_1104.n10 a_5684_1104.n9 15.8172
R4113 a_5684_1104.n22 a_5684_1104.n21 15.8172
R4114 a_5684_1104.n1 a_5684_1104.n0 15.8172
R4115 a_5684_1104.n2 a_5684_1104.n1 15.8172
R4116 a_5684_1104.n3 a_5684_1104.n2 15.8172
R4117 a_5684_1104.n4 a_5684_1104.n3 15.8172
R4118 a_5684_1104.n5 a_5684_1104.n4 15.8172
R4119 a_5684_1104.n15 a_5684_1104.n14 15.1845
R4120 a_5684_1104.n16 a_5684_1104.n15 15.1845
R4121 a_5684_1104.n17 a_5684_1104.n16 15.1845
R4122 a_5684_1104.n7 a_5684_1104.t2 5.44589
R4123 a_5684_1104.n7 a_5684_1104.t0 4.7885
R4124 a_5684_1104.n6 a_5684_1104.t4 4.70615
R4125 a_5684_1104.n8 a_5684_1104.t5 4.4205
R4126 a_5684_1104.n20 a_5684_1104.t3 4.4205
R4127 a_5684_1104.t1 a_5684_1104.n28 4.4205
R4128 a_5684_1104.n8 a_5684_1104.n7 1.1392
R4129 a_5684_1104.n20 a_5684_1104.n19 0.286152
R4130 a_5684_1104.n28 a_5684_1104.n27 0.286152
R4131 a_5684_1104.n27 a_5684_1104.n20 0.282239
R4132 a_5684_1104.n19 a_5684_1104.n8 0.282239
R4133 a_5684_1104.n28 a_5684_1104.n6 0.282239
R4134 TG_GATE_SWITCH_magic_3.B.n106 TG_GATE_SWITCH_magic_3.B.n105 10.8777
R4135 TG_GATE_SWITCH_magic_3.B.n64 TG_GATE_SWITCH_magic_3.B.t56 5.44589
R4136 TG_GATE_SWITCH_magic_3.B.n91 TG_GATE_SWITCH_magic_3.B.t50 5.07789
R4137 TG_GATE_SWITCH_magic_3.B.n68 TG_GATE_SWITCH_magic_3.B.n52 4.7885
R4138 TG_GATE_SWITCH_magic_3.B.n67 TG_GATE_SWITCH_magic_3.B.n53 4.7885
R4139 TG_GATE_SWITCH_magic_3.B.n64 TG_GATE_SWITCH_magic_3.B.t0 4.7885
R4140 TG_GATE_SWITCH_magic_3.B.n103 TG_GATE_SWITCH_magic_3.B.n102 4.4205
R4141 TG_GATE_SWITCH_magic_3.B.n99 TG_GATE_SWITCH_magic_3.B.n98 4.4205
R4142 TG_GATE_SWITCH_magic_3.B.n97 TG_GATE_SWITCH_magic_3.B.n96 4.4205
R4143 TG_GATE_SWITCH_magic_3.B.n93 TG_GATE_SWITCH_magic_3.B.t51 4.4205
R4144 TG_GATE_SWITCH_magic_3.B.n92 TG_GATE_SWITCH_magic_3.B.t36 4.4205
R4145 TG_GATE_SWITCH_magic_3.B.n91 TG_GATE_SWITCH_magic_3.B.t37 4.4205
R4146 TG_GATE_SWITCH_magic_3.B.n101 TG_GATE_SWITCH_magic_3.B.n100 4.4205
R4147 TG_GATE_SWITCH_magic_3.B.n58 TG_GATE_SWITCH_magic_3.B.n55 3.80789
R4148 TG_GATE_SWITCH_magic_3.B.n63 TG_GATE_SWITCH_magic_3.B.n60 3.80789
R4149 TG_GATE_SWITCH_magic_3.B.n48 TG_GATE_SWITCH_magic_3.B.n47 3.80789
R4150 TG_GATE_SWITCH_magic_3.B.n43 TG_GATE_SWITCH_magic_3.B.n42 3.80789
R4151 TG_GATE_SWITCH_magic_3.B.n38 TG_GATE_SWITCH_magic_3.B.n37 3.80789
R4152 TG_GATE_SWITCH_magic_3.B.n88 TG_GATE_SWITCH_magic_3.B.n87 3.25789
R4153 TG_GATE_SWITCH_magic_3.B.n77 TG_GATE_SWITCH_magic_3.B.n76 3.25789
R4154 TG_GATE_SWITCH_magic_3.B.n4 TG_GATE_SWITCH_magic_3.B.n1 3.25789
R4155 TG_GATE_SWITCH_magic_3.B.n15 TG_GATE_SWITCH_magic_3.B.n12 3.25789
R4156 TG_GATE_SWITCH_magic_3.B.n27 TG_GATE_SWITCH_magic_3.B.n24 3.25789
R4157 TG_GATE_SWITCH_magic_3.B.n58 TG_GATE_SWITCH_magic_3.B.n57 3.1505
R4158 TG_GATE_SWITCH_magic_3.B.n63 TG_GATE_SWITCH_magic_3.B.n62 3.1505
R4159 TG_GATE_SWITCH_magic_3.B.n48 TG_GATE_SWITCH_magic_3.B.n45 3.1505
R4160 TG_GATE_SWITCH_magic_3.B.n43 TG_GATE_SWITCH_magic_3.B.n40 3.1505
R4161 TG_GATE_SWITCH_magic_3.B.n38 TG_GATE_SWITCH_magic_3.B.n35 3.1505
R4162 TG_GATE_SWITCH_magic_3.B.n88 TG_GATE_SWITCH_magic_3.B.n85 2.6005
R4163 TG_GATE_SWITCH_magic_3.B.n89 TG_GATE_SWITCH_magic_3.B.n83 2.6005
R4164 TG_GATE_SWITCH_magic_3.B.n90 TG_GATE_SWITCH_magic_3.B.n81 2.6005
R4165 TG_GATE_SWITCH_magic_3.B.n77 TG_GATE_SWITCH_magic_3.B.n74 2.6005
R4166 TG_GATE_SWITCH_magic_3.B.n78 TG_GATE_SWITCH_magic_3.B.n72 2.6005
R4167 TG_GATE_SWITCH_magic_3.B.n79 TG_GATE_SWITCH_magic_3.B.n70 2.6005
R4168 TG_GATE_SWITCH_magic_3.B.n4 TG_GATE_SWITCH_magic_3.B.n3 2.6005
R4169 TG_GATE_SWITCH_magic_3.B.n7 TG_GATE_SWITCH_magic_3.B.n6 2.6005
R4170 TG_GATE_SWITCH_magic_3.B.n10 TG_GATE_SWITCH_magic_3.B.n9 2.6005
R4171 TG_GATE_SWITCH_magic_3.B.n18 TG_GATE_SWITCH_magic_3.B.n17 2.6005
R4172 TG_GATE_SWITCH_magic_3.B.n15 TG_GATE_SWITCH_magic_3.B.n14 2.6005
R4173 TG_GATE_SWITCH_magic_3.B.n21 TG_GATE_SWITCH_magic_3.B.n20 2.6005
R4174 TG_GATE_SWITCH_magic_3.B.n27 TG_GATE_SWITCH_magic_3.B.n26 2.6005
R4175 TG_GATE_SWITCH_magic_3.B.n30 TG_GATE_SWITCH_magic_3.B.n29 2.6005
R4176 TG_GATE_SWITCH_magic_3.B.n33 TG_GATE_SWITCH_magic_3.B.n32 2.6005
R4177 TG_GATE_SWITCH_magic_3.B.n81 TG_GATE_SWITCH_magic_3.B.t31 1.8205
R4178 TG_GATE_SWITCH_magic_3.B.n81 TG_GATE_SWITCH_magic_3.B.n80 1.8205
R4179 TG_GATE_SWITCH_magic_3.B.n83 TG_GATE_SWITCH_magic_3.B.t38 1.8205
R4180 TG_GATE_SWITCH_magic_3.B.n83 TG_GATE_SWITCH_magic_3.B.n82 1.8205
R4181 TG_GATE_SWITCH_magic_3.B.n85 TG_GATE_SWITCH_magic_3.B.t45 1.8205
R4182 TG_GATE_SWITCH_magic_3.B.n85 TG_GATE_SWITCH_magic_3.B.n84 1.8205
R4183 TG_GATE_SWITCH_magic_3.B.n87 TG_GATE_SWITCH_magic_3.B.t30 1.8205
R4184 TG_GATE_SWITCH_magic_3.B.n87 TG_GATE_SWITCH_magic_3.B.n86 1.8205
R4185 TG_GATE_SWITCH_magic_3.B.n70 TG_GATE_SWITCH_magic_3.B.t40 1.8205
R4186 TG_GATE_SWITCH_magic_3.B.n70 TG_GATE_SWITCH_magic_3.B.n69 1.8205
R4187 TG_GATE_SWITCH_magic_3.B.n72 TG_GATE_SWITCH_magic_3.B.t48 1.8205
R4188 TG_GATE_SWITCH_magic_3.B.n72 TG_GATE_SWITCH_magic_3.B.n71 1.8205
R4189 TG_GATE_SWITCH_magic_3.B.n74 TG_GATE_SWITCH_magic_3.B.t52 1.8205
R4190 TG_GATE_SWITCH_magic_3.B.n74 TG_GATE_SWITCH_magic_3.B.n73 1.8205
R4191 TG_GATE_SWITCH_magic_3.B.n76 TG_GATE_SWITCH_magic_3.B.t39 1.8205
R4192 TG_GATE_SWITCH_magic_3.B.n76 TG_GATE_SWITCH_magic_3.B.n75 1.8205
R4193 TG_GATE_SWITCH_magic_3.B.n9 TG_GATE_SWITCH_magic_3.B.t68 1.8205
R4194 TG_GATE_SWITCH_magic_3.B.n9 TG_GATE_SWITCH_magic_3.B.n8 1.8205
R4195 TG_GATE_SWITCH_magic_3.B.n6 TG_GATE_SWITCH_magic_3.B.t28 1.8205
R4196 TG_GATE_SWITCH_magic_3.B.n6 TG_GATE_SWITCH_magic_3.B.n5 1.8205
R4197 TG_GATE_SWITCH_magic_3.B.n3 TG_GATE_SWITCH_magic_3.B.t67 1.8205
R4198 TG_GATE_SWITCH_magic_3.B.n3 TG_GATE_SWITCH_magic_3.B.n2 1.8205
R4199 TG_GATE_SWITCH_magic_3.B.n1 TG_GATE_SWITCH_magic_3.B.t66 1.8205
R4200 TG_GATE_SWITCH_magic_3.B.n1 TG_GATE_SWITCH_magic_3.B.n0 1.8205
R4201 TG_GATE_SWITCH_magic_3.B.n20 TG_GATE_SWITCH_magic_3.B.t60 1.8205
R4202 TG_GATE_SWITCH_magic_3.B.n20 TG_GATE_SWITCH_magic_3.B.n19 1.8205
R4203 TG_GATE_SWITCH_magic_3.B.n12 TG_GATE_SWITCH_magic_3.B.t59 1.8205
R4204 TG_GATE_SWITCH_magic_3.B.n12 TG_GATE_SWITCH_magic_3.B.n11 1.8205
R4205 TG_GATE_SWITCH_magic_3.B.n14 TG_GATE_SWITCH_magic_3.B.t54 1.8205
R4206 TG_GATE_SWITCH_magic_3.B.n14 TG_GATE_SWITCH_magic_3.B.n13 1.8205
R4207 TG_GATE_SWITCH_magic_3.B.n17 TG_GATE_SWITCH_magic_3.B.t4 1.8205
R4208 TG_GATE_SWITCH_magic_3.B.n17 TG_GATE_SWITCH_magic_3.B.n16 1.8205
R4209 TG_GATE_SWITCH_magic_3.B.n32 TG_GATE_SWITCH_magic_3.B.t8 1.8205
R4210 TG_GATE_SWITCH_magic_3.B.n32 TG_GATE_SWITCH_magic_3.B.n31 1.8205
R4211 TG_GATE_SWITCH_magic_3.B.n29 TG_GATE_SWITCH_magic_3.B.t64 1.8205
R4212 TG_GATE_SWITCH_magic_3.B.n29 TG_GATE_SWITCH_magic_3.B.n28 1.8205
R4213 TG_GATE_SWITCH_magic_3.B.n26 TG_GATE_SWITCH_magic_3.B.t6 1.8205
R4214 TG_GATE_SWITCH_magic_3.B.n26 TG_GATE_SWITCH_magic_3.B.n25 1.8205
R4215 TG_GATE_SWITCH_magic_3.B.n24 TG_GATE_SWITCH_magic_3.B.t7 1.8205
R4216 TG_GATE_SWITCH_magic_3.B.n24 TG_GATE_SWITCH_magic_3.B.n23 1.8205
R4217 TG_GATE_SWITCH_magic_3.B.n57 TG_GATE_SWITCH_magic_3.B.t2 1.6385
R4218 TG_GATE_SWITCH_magic_3.B.n57 TG_GATE_SWITCH_magic_3.B.n56 1.6385
R4219 TG_GATE_SWITCH_magic_3.B.n55 TG_GATE_SWITCH_magic_3.B.t24 1.6385
R4220 TG_GATE_SWITCH_magic_3.B.n55 TG_GATE_SWITCH_magic_3.B.n54 1.6385
R4221 TG_GATE_SWITCH_magic_3.B.n62 TG_GATE_SWITCH_magic_3.B.t23 1.6385
R4222 TG_GATE_SWITCH_magic_3.B.n62 TG_GATE_SWITCH_magic_3.B.n61 1.6385
R4223 TG_GATE_SWITCH_magic_3.B.n60 TG_GATE_SWITCH_magic_3.B.t1 1.6385
R4224 TG_GATE_SWITCH_magic_3.B.n60 TG_GATE_SWITCH_magic_3.B.n59 1.6385
R4225 TG_GATE_SWITCH_magic_3.B.n45 TG_GATE_SWITCH_magic_3.B.t14 1.6385
R4226 TG_GATE_SWITCH_magic_3.B.n45 TG_GATE_SWITCH_magic_3.B.n44 1.6385
R4227 TG_GATE_SWITCH_magic_3.B.n47 TG_GATE_SWITCH_magic_3.B.t10 1.6385
R4228 TG_GATE_SWITCH_magic_3.B.n47 TG_GATE_SWITCH_magic_3.B.n46 1.6385
R4229 TG_GATE_SWITCH_magic_3.B.n40 TG_GATE_SWITCH_magic_3.B.t12 1.6385
R4230 TG_GATE_SWITCH_magic_3.B.n40 TG_GATE_SWITCH_magic_3.B.n39 1.6385
R4231 TG_GATE_SWITCH_magic_3.B.n42 TG_GATE_SWITCH_magic_3.B.t13 1.6385
R4232 TG_GATE_SWITCH_magic_3.B.n42 TG_GATE_SWITCH_magic_3.B.n41 1.6385
R4233 TG_GATE_SWITCH_magic_3.B.n35 TG_GATE_SWITCH_magic_3.B.t9 1.6385
R4234 TG_GATE_SWITCH_magic_3.B.n35 TG_GATE_SWITCH_magic_3.B.n34 1.6385
R4235 TG_GATE_SWITCH_magic_3.B.n37 TG_GATE_SWITCH_magic_3.B.t11 1.6385
R4236 TG_GATE_SWITCH_magic_3.B.n37 TG_GATE_SWITCH_magic_3.B.n36 1.6385
R4237 TG_GATE_SWITCH_magic_3.B.n105 TG_GATE_SWITCH_magic_3.B.n104 1.53161
R4238 TG_GATE_SWITCH_magic_3.B.n105 TG_GATE_SWITCH_magic_3.B 1.19982
R4239 TG_GATE_SWITCH_magic_3.B.n65 TG_GATE_SWITCH_magic_3.B.n64 0.884196
R4240 TG_GATE_SWITCH_magic_3.B.n67 TG_GATE_SWITCH_magic_3.B.n66 0.884196
R4241 TG_GATE_SWITCH_magic_3.B.n94 TG_GATE_SWITCH_magic_3.B.n93 0.882239
R4242 TG_GATE_SWITCH_magic_3.B.n97 TG_GATE_SWITCH_magic_3.B.n95 0.882239
R4243 TG_GATE_SWITCH_magic_3.B.n104 TG_GATE_SWITCH_magic_3.B.n68 0.8105
R4244 TG_GATE_SWITCH_magic_3.B.n93 TG_GATE_SWITCH_magic_3.B.n92 0.657891
R4245 TG_GATE_SWITCH_magic_3.B.n92 TG_GATE_SWITCH_magic_3.B.n91 0.657891
R4246 TG_GATE_SWITCH_magic_3.B.n90 TG_GATE_SWITCH_magic_3.B.n89 0.657891
R4247 TG_GATE_SWITCH_magic_3.B.n89 TG_GATE_SWITCH_magic_3.B.n88 0.657891
R4248 TG_GATE_SWITCH_magic_3.B.n79 TG_GATE_SWITCH_magic_3.B.n78 0.657891
R4249 TG_GATE_SWITCH_magic_3.B.n78 TG_GATE_SWITCH_magic_3.B.n77 0.657891
R4250 TG_GATE_SWITCH_magic_3.B.n68 TG_GATE_SWITCH_magic_3.B.n67 0.657891
R4251 TG_GATE_SWITCH_magic_3.B.n7 TG_GATE_SWITCH_magic_3.B.n4 0.657891
R4252 TG_GATE_SWITCH_magic_3.B.n10 TG_GATE_SWITCH_magic_3.B.n7 0.657891
R4253 TG_GATE_SWITCH_magic_3.B.n18 TG_GATE_SWITCH_magic_3.B.n15 0.657891
R4254 TG_GATE_SWITCH_magic_3.B.n30 TG_GATE_SWITCH_magic_3.B.n27 0.657891
R4255 TG_GATE_SWITCH_magic_3.B.n33 TG_GATE_SWITCH_magic_3.B.n30 0.657891
R4256 TG_GATE_SWITCH_magic_3.B.n99 TG_GATE_SWITCH_magic_3.B.n97 0.657891
R4257 TG_GATE_SWITCH_magic_3.B.n101 TG_GATE_SWITCH_magic_3.B.n99 0.657891
R4258 TG_GATE_SWITCH_magic_3.B.n103 TG_GATE_SWITCH_magic_3.B.n101 0.657891
R4259 TG_GATE_SWITCH_magic_3.B.n21 TG_GATE_SWITCH_magic_3.B.n18 0.655976
R4260 TG_GATE_SWITCH_magic_3.B.n22 TG_GATE_SWITCH_magic_3.B.n21 0.645657
R4261 TG_GATE_SWITCH_magic_3.B.n95 TG_GATE_SWITCH_magic_3.B.n94 0.6005
R4262 TG_GATE_SWITCH_magic_3.B.n66 TG_GATE_SWITCH_magic_3.B.n65 0.6005
R4263 TG_GATE_SWITCH_magic_3.B.n49 TG_GATE_SWITCH_magic_3.B.n48 0.548416
R4264 TG_GATE_SWITCH_magic_3.B.n51 TG_GATE_SWITCH_magic_3.B.n33 0.317366
R4265 TG_GATE_SWITCH_magic_3.B.n50 TG_GATE_SWITCH_magic_3.B.n38 0.304838
R4266 TG_GATE_SWITCH_magic_3.B.n66 TG_GATE_SWITCH_magic_3.B.n58 0.284196
R4267 TG_GATE_SWITCH_magic_3.B.n65 TG_GATE_SWITCH_magic_3.B.n63 0.284196
R4268 TG_GATE_SWITCH_magic_3.B.n49 TG_GATE_SWITCH_magic_3.B.n43 0.284196
R4269 TG_GATE_SWITCH_magic_3.B.n51 TG_GATE_SWITCH_magic_3.B.n22 0.283032
R4270 TG_GATE_SWITCH_magic_3.B.n94 TG_GATE_SWITCH_magic_3.B.n90 0.282239
R4271 TG_GATE_SWITCH_magic_3.B.n95 TG_GATE_SWITCH_magic_3.B.n79 0.282239
R4272 TG_GATE_SWITCH_magic_3.B.n22 TG_GATE_SWITCH_magic_3.B.n10 0.279866
R4273 TG_GATE_SWITCH_magic_3.B.n106 TG_GATE_SWITCH_magic_3.B.n51 0.255514
R4274 TG_GATE_SWITCH_magic_3.B.n50 TG_GATE_SWITCH_magic_3.B.n49 0.244078
R4275 TG_GATE_SWITCH_magic_3.B.n104 TG_GATE_SWITCH_magic_3.B.n103 0.237239
R4276 TG_GATE_SWITCH_magic_3.B.n51 TG_GATE_SWITCH_magic_3.B.n50 0.1355
R4277 TG_GATE_SWITCH_magic_3.B TG_GATE_SWITCH_magic_3.B.n106 0.0324516
R4278 a_3817_n991.t29 a_3817_n991.n16 40.7345
R4279 a_3817_n991.n20 a_3817_n991.n5 28.094
R4280 a_3817_n991.n18 a_3817_n991.n17 28.094
R4281 a_3817_n991.n28 a_3817_n991.n27 28.094
R4282 a_3817_n991.n22 a_3817_n991.t18 21.9005
R4283 a_3817_n991.n22 a_3817_n991.t11 21.9005
R4284 a_3817_n991.n0 a_3817_n991.t6 21.9005
R4285 a_3817_n991.n8 a_3817_n991.t24 21.9005
R4286 a_3817_n991.n9 a_3817_n991.t12 21.9005
R4287 a_3817_n991.n1 a_3817_n991.t17 21.9005
R4288 a_3817_n991.n23 a_3817_n991.t23 21.9005
R4289 a_3817_n991.n23 a_3817_n991.t28 21.9005
R4290 a_3817_n991.n24 a_3817_n991.t21 21.9005
R4291 a_3817_n991.n24 a_3817_n991.t14 21.9005
R4292 a_3817_n991.n2 a_3817_n991.t8 21.9005
R4293 a_3817_n991.n10 a_3817_n991.t27 21.9005
R4294 a_3817_n991.n11 a_3817_n991.t15 21.9005
R4295 a_3817_n991.n3 a_3817_n991.t19 21.9005
R4296 a_3817_n991.n25 a_3817_n991.t25 21.9005
R4297 a_3817_n991.n25 a_3817_n991.t7 21.9005
R4298 a_3817_n991.n26 a_3817_n991.t26 21.9005
R4299 a_3817_n991.n26 a_3817_n991.t20 21.9005
R4300 a_3817_n991.n4 a_3817_n991.t13 21.9005
R4301 a_3817_n991.n12 a_3817_n991.t10 21.9005
R4302 a_3817_n991.n17 a_3817_n991.t29 21.9005
R4303 a_3817_n991.n5 a_3817_n991.t9 21.9005
R4304 a_3817_n991.n27 a_3817_n991.t16 21.9005
R4305 a_3817_n991.n27 a_3817_n991.t22 21.9005
R4306 a_3817_n991.n17 a_3817_n991.n12 15.8172
R4307 a_3817_n991.n5 a_3817_n991.n4 15.8172
R4308 a_3817_n991.n4 a_3817_n991.n3 15.8172
R4309 a_3817_n991.n12 a_3817_n991.n11 15.8172
R4310 a_3817_n991.n11 a_3817_n991.n10 15.8172
R4311 a_3817_n991.n3 a_3817_n991.n2 15.8172
R4312 a_3817_n991.n2 a_3817_n991.n1 15.8172
R4313 a_3817_n991.n10 a_3817_n991.n9 15.8172
R4314 a_3817_n991.n9 a_3817_n991.n8 15.8172
R4315 a_3817_n991.n1 a_3817_n991.n0 15.8172
R4316 a_3817_n991.n23 a_3817_n991.n22 15.8172
R4317 a_3817_n991.n24 a_3817_n991.n23 15.8172
R4318 a_3817_n991.n25 a_3817_n991.n24 15.8172
R4319 a_3817_n991.n26 a_3817_n991.n25 15.8172
R4320 a_3817_n991.n27 a_3817_n991.n26 15.8172
R4321 a_3817_n991.n14 a_3817_n991.n13 15.1845
R4322 a_3817_n991.n15 a_3817_n991.n14 15.1845
R4323 a_3817_n991.n16 a_3817_n991.n15 15.1845
R4324 a_3817_n991.n6 a_3817_n991.t4 5.44589
R4325 a_3817_n991.n6 a_3817_n991.t5 4.7885
R4326 a_3817_n991.t3 a_3817_n991.n28 4.70615
R4327 a_3817_n991.n19 a_3817_n991.t1 4.4205
R4328 a_3817_n991.n21 a_3817_n991.t0 4.4205
R4329 a_3817_n991.n7 a_3817_n991.t2 4.4205
R4330 a_3817_n991.n7 a_3817_n991.n6 1.1392
R4331 a_3817_n991.n21 a_3817_n991.n20 0.286152
R4332 a_3817_n991.n19 a_3817_n991.n18 0.286152
R4333 a_3817_n991.n28 a_3817_n991.n21 0.282239
R4334 a_3817_n991.n18 a_3817_n991.n7 0.282239
R4335 a_3817_n991.n20 a_3817_n991.n19 0.282239
R4336 TG_magic_4.B.n114 TG_magic_4.B.n112 5.44589
R4337 TG_magic_4.B.n162 TG_magic_4.B 5.33254
R4338 TG_magic_4.B.n153 TG_magic_4.B.n152 5.07789
R4339 TG_magic_4.B.n163 TG_magic_4.B.t98 4.7885
R4340 TG_magic_4.B.n114 TG_magic_4.B.n113 4.7885
R4341 TG_magic_4.B.n158 TG_magic_4.B.t77 4.4205
R4342 TG_magic_4.B.n159 TG_magic_4.B.t43 4.4205
R4343 TG_magic_4.B.n160 TG_magic_4.B.t47 4.4205
R4344 TG_magic_4.B.n161 TG_magic_4.B.t75 4.4205
R4345 TG_magic_4.B.n155 TG_magic_4.B.n149 4.4205
R4346 TG_magic_4.B.n154 TG_magic_4.B.n150 4.4205
R4347 TG_magic_4.B.n153 TG_magic_4.B.n151 4.4205
R4348 TG_magic_4.B.n110 TG_magic_4.B.n109 3.86778
R4349 TG_magic_4.B.n29 TG_magic_4.B.n26 3.80789
R4350 TG_magic_4.B.n40 TG_magic_4.B.n37 3.80789
R4351 TG_magic_4.B.n81 TG_magic_4.B.n78 3.80789
R4352 TG_magic_4.B.n86 TG_magic_4.B.n83 3.80789
R4353 TG_magic_4.B.n91 TG_magic_4.B.n88 3.80789
R4354 TG_magic_4.B.n120 TG_magic_4.B.n117 3.80789
R4355 TG_magic_4.B.n34 TG_magic_4.B.n31 3.80789
R4356 TG_magic_4.B.n10 TG_magic_4.B.n9 3.25789
R4357 TG_magic_4.B.n21 TG_magic_4.B.n20 3.25789
R4358 TG_magic_4.B.n73 TG_magic_4.B.n72 3.25789
R4359 TG_magic_4.B.n62 TG_magic_4.B.n61 3.25789
R4360 TG_magic_4.B.n102 TG_magic_4.B.n101 3.25789
R4361 TG_magic_4.B.n135 TG_magic_4.B.n134 3.25789
R4362 TG_magic_4.B.n146 TG_magic_4.B.n145 3.25789
R4363 TG_magic_4.B.n50 TG_magic_4.B.n49 3.25789
R4364 TG_magic_4.B.n167 TG_magic_4.B.n0 3.18617
R4365 TG_magic_4.B.n29 TG_magic_4.B.n28 3.1505
R4366 TG_magic_4.B.n40 TG_magic_4.B.n39 3.1505
R4367 TG_magic_4.B.n81 TG_magic_4.B.n80 3.1505
R4368 TG_magic_4.B.n86 TG_magic_4.B.n85 3.1505
R4369 TG_magic_4.B.n91 TG_magic_4.B.n90 3.1505
R4370 TG_magic_4.B.n120 TG_magic_4.B.n119 3.1505
R4371 TG_magic_4.B.n34 TG_magic_4.B.n33 3.1505
R4372 TG_magic_4.B.n164 TG_magic_4.B.t95 3.02839
R4373 TG_magic_4.B.n123 TG_magic_4.B.n115 2.60595
R4374 TG_magic_4.B.n10 TG_magic_4.B.n7 2.6005
R4375 TG_magic_4.B.n11 TG_magic_4.B.n5 2.6005
R4376 TG_magic_4.B.n12 TG_magic_4.B.n3 2.6005
R4377 TG_magic_4.B.n21 TG_magic_4.B.n18 2.6005
R4378 TG_magic_4.B.n22 TG_magic_4.B.n16 2.6005
R4379 TG_magic_4.B.n23 TG_magic_4.B.n14 2.6005
R4380 TG_magic_4.B.n73 TG_magic_4.B.n70 2.6005
R4381 TG_magic_4.B.n74 TG_magic_4.B.n68 2.6005
R4382 TG_magic_4.B.n75 TG_magic_4.B.n66 2.6005
R4383 TG_magic_4.B.n62 TG_magic_4.B.n59 2.6005
R4384 TG_magic_4.B.n63 TG_magic_4.B.n57 2.6005
R4385 TG_magic_4.B.n64 TG_magic_4.B.n55 2.6005
R4386 TG_magic_4.B.n102 TG_magic_4.B.n99 2.6005
R4387 TG_magic_4.B.n103 TG_magic_4.B.n97 2.6005
R4388 TG_magic_4.B.n104 TG_magic_4.B.n95 2.6005
R4389 TG_magic_4.B.n135 TG_magic_4.B.n132 2.6005
R4390 TG_magic_4.B.n136 TG_magic_4.B.n130 2.6005
R4391 TG_magic_4.B.n137 TG_magic_4.B.n128 2.6005
R4392 TG_magic_4.B.n146 TG_magic_4.B.n143 2.6005
R4393 TG_magic_4.B.n147 TG_magic_4.B.n141 2.6005
R4394 TG_magic_4.B.n148 TG_magic_4.B.n139 2.6005
R4395 TG_magic_4.B.n50 TG_magic_4.B.n47 2.6005
R4396 TG_magic_4.B.n51 TG_magic_4.B.n45 2.6005
R4397 TG_magic_4.B.n52 TG_magic_4.B.n43 2.6005
R4398 TG_magic_4.B.n0 TG_magic_4.B.n166 2.25068
R4399 TG_magic_4.B.n123 TG_magic_4.B.n122 2.2505
R4400 TG_magic_4.B.n1 TG_magic_4.B.n125 2.25002
R4401 TG_magic_4.B.n1 TG_magic_4.B.n111 2.24533
R4402 TG_magic_4.B.n3 TG_magic_4.B.t41 1.8205
R4403 TG_magic_4.B.n3 TG_magic_4.B.n2 1.8205
R4404 TG_magic_4.B.n5 TG_magic_4.B.t13 1.8205
R4405 TG_magic_4.B.n5 TG_magic_4.B.n4 1.8205
R4406 TG_magic_4.B.n7 TG_magic_4.B.t33 1.8205
R4407 TG_magic_4.B.n7 TG_magic_4.B.n6 1.8205
R4408 TG_magic_4.B.n9 TG_magic_4.B.t32 1.8205
R4409 TG_magic_4.B.n9 TG_magic_4.B.n8 1.8205
R4410 TG_magic_4.B.n14 TG_magic_4.B.t31 1.8205
R4411 TG_magic_4.B.n14 TG_magic_4.B.n13 1.8205
R4412 TG_magic_4.B.n16 TG_magic_4.B.t36 1.8205
R4413 TG_magic_4.B.n16 TG_magic_4.B.n15 1.8205
R4414 TG_magic_4.B.n18 TG_magic_4.B.t18 1.8205
R4415 TG_magic_4.B.n18 TG_magic_4.B.n17 1.8205
R4416 TG_magic_4.B.n20 TG_magic_4.B.t15 1.8205
R4417 TG_magic_4.B.n20 TG_magic_4.B.n19 1.8205
R4418 TG_magic_4.B.n66 TG_magic_4.B.t12 1.8205
R4419 TG_magic_4.B.n66 TG_magic_4.B.n65 1.8205
R4420 TG_magic_4.B.n68 TG_magic_4.B.t89 1.8205
R4421 TG_magic_4.B.n68 TG_magic_4.B.n67 1.8205
R4422 TG_magic_4.B.n70 TG_magic_4.B.t6 1.8205
R4423 TG_magic_4.B.n70 TG_magic_4.B.n69 1.8205
R4424 TG_magic_4.B.n72 TG_magic_4.B.t4 1.8205
R4425 TG_magic_4.B.n72 TG_magic_4.B.n71 1.8205
R4426 TG_magic_4.B.n55 TG_magic_4.B.t85 1.8205
R4427 TG_magic_4.B.n55 TG_magic_4.B.n54 1.8205
R4428 TG_magic_4.B.n57 TG_magic_4.B.t92 1.8205
R4429 TG_magic_4.B.n57 TG_magic_4.B.n56 1.8205
R4430 TG_magic_4.B.n59 TG_magic_4.B.t8 1.8205
R4431 TG_magic_4.B.n59 TG_magic_4.B.n58 1.8205
R4432 TG_magic_4.B.n61 TG_magic_4.B.t7 1.8205
R4433 TG_magic_4.B.n61 TG_magic_4.B.n60 1.8205
R4434 TG_magic_4.B.n95 TG_magic_4.B.t93 1.8205
R4435 TG_magic_4.B.n95 TG_magic_4.B.n94 1.8205
R4436 TG_magic_4.B.n97 TG_magic_4.B.t69 1.8205
R4437 TG_magic_4.B.n97 TG_magic_4.B.n96 1.8205
R4438 TG_magic_4.B.n99 TG_magic_4.B.t84 1.8205
R4439 TG_magic_4.B.n99 TG_magic_4.B.n98 1.8205
R4440 TG_magic_4.B.n101 TG_magic_4.B.t11 1.8205
R4441 TG_magic_4.B.n101 TG_magic_4.B.n100 1.8205
R4442 TG_magic_4.B.n128 TG_magic_4.B.t2 1.8205
R4443 TG_magic_4.B.n128 TG_magic_4.B.n127 1.8205
R4444 TG_magic_4.B.n130 TG_magic_4.B.t48 1.8205
R4445 TG_magic_4.B.n130 TG_magic_4.B.n129 1.8205
R4446 TG_magic_4.B.n132 TG_magic_4.B.t74 1.8205
R4447 TG_magic_4.B.n132 TG_magic_4.B.n131 1.8205
R4448 TG_magic_4.B.n134 TG_magic_4.B.t72 1.8205
R4449 TG_magic_4.B.n134 TG_magic_4.B.n133 1.8205
R4450 TG_magic_4.B.n139 TG_magic_4.B.t25 1.8205
R4451 TG_magic_4.B.n139 TG_magic_4.B.n138 1.8205
R4452 TG_magic_4.B.n141 TG_magic_4.B.t73 1.8205
R4453 TG_magic_4.B.n141 TG_magic_4.B.n140 1.8205
R4454 TG_magic_4.B.n143 TG_magic_4.B.t78 1.8205
R4455 TG_magic_4.B.n143 TG_magic_4.B.n142 1.8205
R4456 TG_magic_4.B.n145 TG_magic_4.B.t24 1.8205
R4457 TG_magic_4.B.n145 TG_magic_4.B.n144 1.8205
R4458 TG_magic_4.B.n43 TG_magic_4.B.t35 1.8205
R4459 TG_magic_4.B.n43 TG_magic_4.B.n42 1.8205
R4460 TG_magic_4.B.n45 TG_magic_4.B.t38 1.8205
R4461 TG_magic_4.B.n45 TG_magic_4.B.n44 1.8205
R4462 TG_magic_4.B.n47 TG_magic_4.B.t21 1.8205
R4463 TG_magic_4.B.n47 TG_magic_4.B.n46 1.8205
R4464 TG_magic_4.B.n49 TG_magic_4.B.t19 1.8205
R4465 TG_magic_4.B.n49 TG_magic_4.B.n48 1.8205
R4466 TG_magic_4.B.n110 TG_magic_4.B.n107 1.81712
R4467 TG_magic_4.B.n31 TG_magic_4.B.t51 1.6385
R4468 TG_magic_4.B.n31 TG_magic_4.B.n30 1.6385
R4469 TG_magic_4.B.n28 TG_magic_4.B.t55 1.6385
R4470 TG_magic_4.B.n28 TG_magic_4.B.n27 1.6385
R4471 TG_magic_4.B.n26 TG_magic_4.B.t58 1.6385
R4472 TG_magic_4.B.n26 TG_magic_4.B.n25 1.6385
R4473 TG_magic_4.B.n39 TG_magic_4.B.t53 1.6385
R4474 TG_magic_4.B.n39 TG_magic_4.B.n38 1.6385
R4475 TG_magic_4.B.n37 TG_magic_4.B.t56 1.6385
R4476 TG_magic_4.B.n37 TG_magic_4.B.n36 1.6385
R4477 TG_magic_4.B.n80 TG_magic_4.B.t66 1.6385
R4478 TG_magic_4.B.n80 TG_magic_4.B.n79 1.6385
R4479 TG_magic_4.B.n78 TG_magic_4.B.t80 1.6385
R4480 TG_magic_4.B.n78 TG_magic_4.B.n77 1.6385
R4481 TG_magic_4.B.n85 TG_magic_4.B.t83 1.6385
R4482 TG_magic_4.B.n85 TG_magic_4.B.n84 1.6385
R4483 TG_magic_4.B.n83 TG_magic_4.B.t1 1.6385
R4484 TG_magic_4.B.n83 TG_magic_4.B.n82 1.6385
R4485 TG_magic_4.B.n90 TG_magic_4.B.t81 1.6385
R4486 TG_magic_4.B.n90 TG_magic_4.B.n89 1.6385
R4487 TG_magic_4.B.n88 TG_magic_4.B.t0 1.6385
R4488 TG_magic_4.B.n88 TG_magic_4.B.n87 1.6385
R4489 TG_magic_4.B.n107 TG_magic_4.B.t100 1.6385
R4490 TG_magic_4.B.n107 TG_magic_4.B.n106 1.6385
R4491 TG_magic_4.B.n109 TG_magic_4.B.t97 1.6385
R4492 TG_magic_4.B.n109 TG_magic_4.B.n108 1.6385
R4493 TG_magic_4.B.n119 TG_magic_4.B.t99 1.6385
R4494 TG_magic_4.B.n119 TG_magic_4.B.n118 1.6385
R4495 TG_magic_4.B.n117 TG_magic_4.B.t96 1.6385
R4496 TG_magic_4.B.n117 TG_magic_4.B.n116 1.6385
R4497 TG_magic_4.B.n33 TG_magic_4.B.t62 1.6385
R4498 TG_magic_4.B.n33 TG_magic_4.B.n32 1.6385
R4499 TG_magic_4.B.n156 TG_magic_4.B.n155 0.882239
R4500 TG_magic_4.B.n158 TG_magic_4.B.n157 0.882239
R4501 TG_magic_4.B.n163 TG_magic_4.B.n162 0.8105
R4502 TG_magic_4.B.n164 TG_magic_4.B.n163 0.745261
R4503 TG_magic_4.B.n12 TG_magic_4.B.n11 0.657891
R4504 TG_magic_4.B.n11 TG_magic_4.B.n10 0.657891
R4505 TG_magic_4.B.n22 TG_magic_4.B.n21 0.657891
R4506 TG_magic_4.B.n74 TG_magic_4.B.n73 0.657891
R4507 TG_magic_4.B.n64 TG_magic_4.B.n63 0.657891
R4508 TG_magic_4.B.n63 TG_magic_4.B.n62 0.657891
R4509 TG_magic_4.B.n104 TG_magic_4.B.n103 0.657891
R4510 TG_magic_4.B.n103 TG_magic_4.B.n102 0.657891
R4511 TG_magic_4.B.n137 TG_magic_4.B.n136 0.657891
R4512 TG_magic_4.B.n136 TG_magic_4.B.n135 0.657891
R4513 TG_magic_4.B.n148 TG_magic_4.B.n147 0.657891
R4514 TG_magic_4.B.n147 TG_magic_4.B.n146 0.657891
R4515 TG_magic_4.B.n155 TG_magic_4.B.n154 0.657891
R4516 TG_magic_4.B.n154 TG_magic_4.B.n153 0.657891
R4517 TG_magic_4.B.n159 TG_magic_4.B.n158 0.657891
R4518 TG_magic_4.B.n160 TG_magic_4.B.n159 0.657891
R4519 TG_magic_4.B.n161 TG_magic_4.B.n160 0.657891
R4520 TG_magic_4.B.n52 TG_magic_4.B.n51 0.657891
R4521 TG_magic_4.B.n51 TG_magic_4.B.n50 0.657891
R4522 TG_magic_4.B.n23 TG_magic_4.B.n22 0.655976
R4523 TG_magic_4.B.n75 TG_magic_4.B.n74 0.655976
R4524 TG_magic_4.B.n24 TG_magic_4.B.n23 0.646796
R4525 TG_magic_4.B.n76 TG_magic_4.B.n75 0.645657
R4526 TG_magic_4.B.n157 TG_magic_4.B.n156 0.6005
R4527 TG_magic_4.B.n35 TG_magic_4.B.n29 0.548416
R4528 TG_magic_4.B.n92 TG_magic_4.B.n91 0.548416
R4529 TG_magic_4.B.n1 TG_magic_4.B.n123 0.338918
R4530 TG_magic_4.B.n105 TG_magic_4.B.n104 0.316429
R4531 TG_magic_4.B.n53 TG_magic_4.B.n52 0.316429
R4532 TG_magic_4.B.n0 TG_magic_4.B.n126 0.308702
R4533 TG_magic_4.B.n41 TG_magic_4.B.n40 0.304838
R4534 TG_magic_4.B.n93 TG_magic_4.B.n81 0.304838
R4535 TG_magic_4.B TG_magic_4.B.n105 0.2873
R4536 TG_magic_4.B TG_magic_4.B.n53 0.2873
R4537 TG_magic_4.B.n92 TG_magic_4.B.n86 0.284196
R4538 TG_magic_4.B.n35 TG_magic_4.B.n34 0.284196
R4539 TG_magic_4.B.n105 TG_magic_4.B.n76 0.283032
R4540 TG_magic_4.B.n157 TG_magic_4.B.n137 0.282239
R4541 TG_magic_4.B.n156 TG_magic_4.B.n148 0.282239
R4542 TG_magic_4.B.n53 TG_magic_4.B.n24 0.281892
R4543 TG_magic_4.B.n24 TG_magic_4.B.n12 0.279866
R4544 TG_magic_4.B.n76 TG_magic_4.B.n64 0.279866
R4545 TG_magic_4.B.n93 TG_magic_4.B.n92 0.244078
R4546 TG_magic_4.B.n41 TG_magic_4.B.n35 0.244078
R4547 TG_magic_4.B.n162 TG_magic_4.B.n161 0.237239
R4548 TG_magic_4.B.n115 TG_magic_4.B.n114 0.218422
R4549 TG_magic_4.B.n122 TG_magic_4.B.n120 0.203127
R4550 TG_magic_4.B.n105 TG_magic_4.B.n93 0.136437
R4551 TG_magic_4.B.n53 TG_magic_4.B.n41 0.136437
R4552 TG_magic_4.B.n111 TG_magic_4.B.n110 0.0902293
R4553 TG_magic_4.B.n165 TG_magic_4.B.n164 0.0754787
R4554 TG_magic_4.B.n167 TG_magic_4.B 0.0689
R4555 TG_magic_4.B TG_magic_4.B.n167 0.0677
R4556 TG_magic_4.B.n125 TG_magic_4.B.n124 0.0587165
R4557 TG_magic_4.B.n122 TG_magic_4.B.n121 0.0513235
R4558 TG_magic_4.B.n126 TG_magic_4.B.n1 0.0379187
R4559 TG_magic_4.B.n166 TG_magic_4.B.n165 0.0350713
R4560 TG_magic_7.B.n94 TG_magic_7.B.n92 5.44589
R4561 TG_magic_7.B.n78 TG_magic_7.B.n77 5.07789
R4562 TG_magic_7.B.n94 TG_magic_7.B.n93 4.7885
R4563 TG_magic_7.B.n103 TG_magic_7.B.t68 4.7885
R4564 TG_magic_7.B.n102 TG_magic_7.B.t74 4.7885
R4565 TG_magic_7.B.n86 TG_magic_7.B.t45 4.4205
R4566 TG_magic_7.B.n85 TG_magic_7.B.t106 4.4205
R4567 TG_magic_7.B.n84 TG_magic_7.B.t107 4.4205
R4568 TG_magic_7.B.n83 TG_magic_7.B.t46 4.4205
R4569 TG_magic_7.B.n80 TG_magic_7.B.n74 4.4205
R4570 TG_magic_7.B.n79 TG_magic_7.B.n75 4.4205
R4571 TG_magic_7.B.n78 TG_magic_7.B.n76 4.4205
R4572 TG_magic_7.B.n91 TG_magic_7.B.n88 3.80789
R4573 TG_magic_7.B.n49 TG_magic_7.B.n48 3.80789
R4574 TG_magic_7.B.n38 TG_magic_7.B.n37 3.80789
R4575 TG_magic_7.B.n43 TG_magic_7.B.n42 3.80789
R4576 TG_magic_7.B.n155 TG_magic_7.B.n154 3.80789
R4577 TG_magic_7.B.n150 TG_magic_7.B.n149 3.80789
R4578 TG_magic_7.B.n145 TG_magic_7.B.n144 3.80789
R4579 TG_magic_7.B.n100 TG_magic_7.B.n97 3.80789
R4580 TG_magic_7.B.n60 TG_magic_7.B.n59 3.25789
R4581 TG_magic_7.B.n71 TG_magic_7.B.n70 3.25789
R4582 TG_magic_7.B.n15 TG_magic_7.B.n12 3.25789
R4583 TG_magic_7.B.n4 TG_magic_7.B.n1 3.25789
R4584 TG_magic_7.B.n27 TG_magic_7.B.n24 3.25789
R4585 TG_magic_7.B.n111 TG_magic_7.B.n108 3.25789
R4586 TG_magic_7.B.n122 TG_magic_7.B.n119 3.25789
R4587 TG_magic_7.B.n134 TG_magic_7.B.n131 3.25789
R4588 TG_magic_7.B.n91 TG_magic_7.B.n90 3.1505
R4589 TG_magic_7.B.n49 TG_magic_7.B.n46 3.1505
R4590 TG_magic_7.B.n38 TG_magic_7.B.n35 3.1505
R4591 TG_magic_7.B.n43 TG_magic_7.B.n40 3.1505
R4592 TG_magic_7.B.n155 TG_magic_7.B.n152 3.1505
R4593 TG_magic_7.B.n150 TG_magic_7.B.n147 3.1505
R4594 TG_magic_7.B.n145 TG_magic_7.B.n142 3.1505
R4595 TG_magic_7.B.n100 TG_magic_7.B.n99 3.1505
R4596 TG_magic_7.B.n106 TG_magic_7.B.n105 2.81987
R4597 TG_magic_7.B.n60 TG_magic_7.B.n57 2.6005
R4598 TG_magic_7.B.n61 TG_magic_7.B.n55 2.6005
R4599 TG_magic_7.B.n62 TG_magic_7.B.n53 2.6005
R4600 TG_magic_7.B.n71 TG_magic_7.B.n68 2.6005
R4601 TG_magic_7.B.n72 TG_magic_7.B.n66 2.6005
R4602 TG_magic_7.B.n73 TG_magic_7.B.n64 2.6005
R4603 TG_magic_7.B.n15 TG_magic_7.B.n14 2.6005
R4604 TG_magic_7.B.n18 TG_magic_7.B.n17 2.6005
R4605 TG_magic_7.B.n21 TG_magic_7.B.n20 2.6005
R4606 TG_magic_7.B.n4 TG_magic_7.B.n3 2.6005
R4607 TG_magic_7.B.n7 TG_magic_7.B.n6 2.6005
R4608 TG_magic_7.B.n10 TG_magic_7.B.n9 2.6005
R4609 TG_magic_7.B.n27 TG_magic_7.B.n26 2.6005
R4610 TG_magic_7.B.n30 TG_magic_7.B.n29 2.6005
R4611 TG_magic_7.B.n33 TG_magic_7.B.n32 2.6005
R4612 TG_magic_7.B.n111 TG_magic_7.B.n110 2.6005
R4613 TG_magic_7.B.n114 TG_magic_7.B.n113 2.6005
R4614 TG_magic_7.B.n117 TG_magic_7.B.n116 2.6005
R4615 TG_magic_7.B.n125 TG_magic_7.B.n124 2.6005
R4616 TG_magic_7.B.n122 TG_magic_7.B.n121 2.6005
R4617 TG_magic_7.B.n128 TG_magic_7.B.n127 2.6005
R4618 TG_magic_7.B.n134 TG_magic_7.B.n133 2.6005
R4619 TG_magic_7.B.n137 TG_magic_7.B.n136 2.6005
R4620 TG_magic_7.B.n140 TG_magic_7.B.n139 2.6005
R4621 TG_magic_7.B.n53 TG_magic_7.B.t105 1.8205
R4622 TG_magic_7.B.n53 TG_magic_7.B.n52 1.8205
R4623 TG_magic_7.B.n55 TG_magic_7.B.t52 1.8205
R4624 TG_magic_7.B.n55 TG_magic_7.B.n54 1.8205
R4625 TG_magic_7.B.n57 TG_magic_7.B.t55 1.8205
R4626 TG_magic_7.B.n57 TG_magic_7.B.n56 1.8205
R4627 TG_magic_7.B.n59 TG_magic_7.B.t48 1.8205
R4628 TG_magic_7.B.n59 TG_magic_7.B.n58 1.8205
R4629 TG_magic_7.B.n64 TG_magic_7.B.t44 1.8205
R4630 TG_magic_7.B.n64 TG_magic_7.B.n63 1.8205
R4631 TG_magic_7.B.n66 TG_magic_7.B.t57 1.8205
R4632 TG_magic_7.B.n66 TG_magic_7.B.n65 1.8205
R4633 TG_magic_7.B.n68 TG_magic_7.B.t104 1.8205
R4634 TG_magic_7.B.n68 TG_magic_7.B.n67 1.8205
R4635 TG_magic_7.B.n70 TG_magic_7.B.t42 1.8205
R4636 TG_magic_7.B.n70 TG_magic_7.B.n69 1.8205
R4637 TG_magic_7.B.n20 TG_magic_7.B.t8 1.8205
R4638 TG_magic_7.B.n20 TG_magic_7.B.n19 1.8205
R4639 TG_magic_7.B.n17 TG_magic_7.B.t35 1.8205
R4640 TG_magic_7.B.n17 TG_magic_7.B.n16 1.8205
R4641 TG_magic_7.B.n14 TG_magic_7.B.t20 1.8205
R4642 TG_magic_7.B.n14 TG_magic_7.B.n13 1.8205
R4643 TG_magic_7.B.n12 TG_magic_7.B.t9 1.8205
R4644 TG_magic_7.B.n12 TG_magic_7.B.n11 1.8205
R4645 TG_magic_7.B.n9 TG_magic_7.B.t17 1.8205
R4646 TG_magic_7.B.n9 TG_magic_7.B.n8 1.8205
R4647 TG_magic_7.B.n6 TG_magic_7.B.t11 1.8205
R4648 TG_magic_7.B.n6 TG_magic_7.B.n5 1.8205
R4649 TG_magic_7.B.n3 TG_magic_7.B.t6 1.8205
R4650 TG_magic_7.B.n3 TG_magic_7.B.n2 1.8205
R4651 TG_magic_7.B.n1 TG_magic_7.B.t18 1.8205
R4652 TG_magic_7.B.n1 TG_magic_7.B.n0 1.8205
R4653 TG_magic_7.B.n32 TG_magic_7.B.t14 1.8205
R4654 TG_magic_7.B.n32 TG_magic_7.B.n31 1.8205
R4655 TG_magic_7.B.n29 TG_magic_7.B.t10 1.8205
R4656 TG_magic_7.B.n29 TG_magic_7.B.n28 1.8205
R4657 TG_magic_7.B.n26 TG_magic_7.B.t2 1.8205
R4658 TG_magic_7.B.n26 TG_magic_7.B.n25 1.8205
R4659 TG_magic_7.B.n24 TG_magic_7.B.t15 1.8205
R4660 TG_magic_7.B.n24 TG_magic_7.B.n23 1.8205
R4661 TG_magic_7.B.n116 TG_magic_7.B.t28 1.8205
R4662 TG_magic_7.B.n116 TG_magic_7.B.n115 1.8205
R4663 TG_magic_7.B.n113 TG_magic_7.B.t24 1.8205
R4664 TG_magic_7.B.n113 TG_magic_7.B.n112 1.8205
R4665 TG_magic_7.B.n110 TG_magic_7.B.t49 1.8205
R4666 TG_magic_7.B.n110 TG_magic_7.B.n109 1.8205
R4667 TG_magic_7.B.n108 TG_magic_7.B.t29 1.8205
R4668 TG_magic_7.B.n108 TG_magic_7.B.n107 1.8205
R4669 TG_magic_7.B.n127 TG_magic_7.B.t25 1.8205
R4670 TG_magic_7.B.n127 TG_magic_7.B.n126 1.8205
R4671 TG_magic_7.B.n119 TG_magic_7.B.t26 1.8205
R4672 TG_magic_7.B.n119 TG_magic_7.B.n118 1.8205
R4673 TG_magic_7.B.n121 TG_magic_7.B.t63 1.8205
R4674 TG_magic_7.B.n121 TG_magic_7.B.n120 1.8205
R4675 TG_magic_7.B.n124 TG_magic_7.B.t103 1.8205
R4676 TG_magic_7.B.n124 TG_magic_7.B.n123 1.8205
R4677 TG_magic_7.B.n139 TG_magic_7.B.t66 1.8205
R4678 TG_magic_7.B.n139 TG_magic_7.B.n138 1.8205
R4679 TG_magic_7.B.n136 TG_magic_7.B.t33 1.8205
R4680 TG_magic_7.B.n136 TG_magic_7.B.n135 1.8205
R4681 TG_magic_7.B.n133 TG_magic_7.B.t30 1.8205
R4682 TG_magic_7.B.n133 TG_magic_7.B.n132 1.8205
R4683 TG_magic_7.B.n131 TG_magic_7.B.t38 1.8205
R4684 TG_magic_7.B.n131 TG_magic_7.B.n130 1.8205
R4685 TG_magic_7.B.n97 TG_magic_7.B.t72 1.6385
R4686 TG_magic_7.B.n97 TG_magic_7.B.n96 1.6385
R4687 TG_magic_7.B.n90 TG_magic_7.B.t75 1.6385
R4688 TG_magic_7.B.n90 TG_magic_7.B.n89 1.6385
R4689 TG_magic_7.B.n88 TG_magic_7.B.t69 1.6385
R4690 TG_magic_7.B.n88 TG_magic_7.B.n87 1.6385
R4691 TG_magic_7.B.n46 TG_magic_7.B.t84 1.6385
R4692 TG_magic_7.B.n46 TG_magic_7.B.n45 1.6385
R4693 TG_magic_7.B.n48 TG_magic_7.B.t81 1.6385
R4694 TG_magic_7.B.n48 TG_magic_7.B.n47 1.6385
R4695 TG_magic_7.B.n35 TG_magic_7.B.t83 1.6385
R4696 TG_magic_7.B.n35 TG_magic_7.B.n34 1.6385
R4697 TG_magic_7.B.n37 TG_magic_7.B.t80 1.6385
R4698 TG_magic_7.B.n37 TG_magic_7.B.n36 1.6385
R4699 TG_magic_7.B.n40 TG_magic_7.B.t79 1.6385
R4700 TG_magic_7.B.n40 TG_magic_7.B.n39 1.6385
R4701 TG_magic_7.B.n42 TG_magic_7.B.t82 1.6385
R4702 TG_magic_7.B.n42 TG_magic_7.B.n41 1.6385
R4703 TG_magic_7.B.n152 TG_magic_7.B.t94 1.6385
R4704 TG_magic_7.B.n152 TG_magic_7.B.n151 1.6385
R4705 TG_magic_7.B.n154 TG_magic_7.B.t100 1.6385
R4706 TG_magic_7.B.n154 TG_magic_7.B.n153 1.6385
R4707 TG_magic_7.B.n147 TG_magic_7.B.t91 1.6385
R4708 TG_magic_7.B.n147 TG_magic_7.B.n146 1.6385
R4709 TG_magic_7.B.n149 TG_magic_7.B.t97 1.6385
R4710 TG_magic_7.B.n149 TG_magic_7.B.n148 1.6385
R4711 TG_magic_7.B.n142 TG_magic_7.B.t98 1.6385
R4712 TG_magic_7.B.n142 TG_magic_7.B.n141 1.6385
R4713 TG_magic_7.B.n144 TG_magic_7.B.t92 1.6385
R4714 TG_magic_7.B.n144 TG_magic_7.B.n143 1.6385
R4715 TG_magic_7.B.n99 TG_magic_7.B.t78 1.6385
R4716 TG_magic_7.B.n99 TG_magic_7.B.n98 1.6385
R4717 TG_magic_7.B.n105 TG_magic_7.B.n104 1.53097
R4718 TG_magic_7.B.n105 TG_magic_7.B 1.18827
R4719 TG_magic_7.B.n95 TG_magic_7.B.n94 0.884196
R4720 TG_magic_7.B.n102 TG_magic_7.B.n101 0.884196
R4721 TG_magic_7.B.n81 TG_magic_7.B.n80 0.882239
R4722 TG_magic_7.B.n83 TG_magic_7.B.n82 0.882239
R4723 TG_magic_7.B.n104 TG_magic_7.B.n103 0.8105
R4724 TG_magic_7.B.n62 TG_magic_7.B.n61 0.657891
R4725 TG_magic_7.B.n61 TG_magic_7.B.n60 0.657891
R4726 TG_magic_7.B.n73 TG_magic_7.B.n72 0.657891
R4727 TG_magic_7.B.n72 TG_magic_7.B.n71 0.657891
R4728 TG_magic_7.B.n80 TG_magic_7.B.n79 0.657891
R4729 TG_magic_7.B.n79 TG_magic_7.B.n78 0.657891
R4730 TG_magic_7.B.n84 TG_magic_7.B.n83 0.657891
R4731 TG_magic_7.B.n85 TG_magic_7.B.n84 0.657891
R4732 TG_magic_7.B.n86 TG_magic_7.B.n85 0.657891
R4733 TG_magic_7.B.n18 TG_magic_7.B.n15 0.657891
R4734 TG_magic_7.B.n7 TG_magic_7.B.n4 0.657891
R4735 TG_magic_7.B.n10 TG_magic_7.B.n7 0.657891
R4736 TG_magic_7.B.n30 TG_magic_7.B.n27 0.657891
R4737 TG_magic_7.B.n33 TG_magic_7.B.n30 0.657891
R4738 TG_magic_7.B.n114 TG_magic_7.B.n111 0.657891
R4739 TG_magic_7.B.n117 TG_magic_7.B.n114 0.657891
R4740 TG_magic_7.B.n125 TG_magic_7.B.n122 0.657891
R4741 TG_magic_7.B.n137 TG_magic_7.B.n134 0.657891
R4742 TG_magic_7.B.n140 TG_magic_7.B.n137 0.657891
R4743 TG_magic_7.B.n103 TG_magic_7.B.n102 0.657891
R4744 TG_magic_7.B.n21 TG_magic_7.B.n18 0.655976
R4745 TG_magic_7.B.n128 TG_magic_7.B.n125 0.655976
R4746 TG_magic_7.B.n22 TG_magic_7.B.n21 0.646796
R4747 TG_magic_7.B.n129 TG_magic_7.B.n128 0.645657
R4748 TG_magic_7.B.n82 TG_magic_7.B.n81 0.6005
R4749 TG_magic_7.B.n101 TG_magic_7.B.n95 0.6005
R4750 TG_magic_7.B.n44 TG_magic_7.B.n43 0.548416
R4751 TG_magic_7.B.n156 TG_magic_7.B.n155 0.548416
R4752 TG_magic_7.B.n51 TG_magic_7.B.n33 0.317366
R4753 TG_magic_7.B.n158 TG_magic_7.B.n140 0.317366
R4754 TG_magic_7.B.n50 TG_magic_7.B.n49 0.304838
R4755 TG_magic_7.B.n157 TG_magic_7.B.n145 0.304838
R4756 TG_magic_7.B TG_magic_7.B.n158 0.2873
R4757 TG_magic_7.B TG_magic_7.B.n51 0.2873
R4758 TG_magic_7.B.n95 TG_magic_7.B.n91 0.284196
R4759 TG_magic_7.B.n44 TG_magic_7.B.n38 0.284196
R4760 TG_magic_7.B.n156 TG_magic_7.B.n150 0.284196
R4761 TG_magic_7.B.n101 TG_magic_7.B.n100 0.284196
R4762 TG_magic_7.B.n158 TG_magic_7.B.n129 0.283032
R4763 TG_magic_7.B.n82 TG_magic_7.B.n62 0.282239
R4764 TG_magic_7.B.n81 TG_magic_7.B.n73 0.282239
R4765 TG_magic_7.B.n51 TG_magic_7.B.n22 0.281892
R4766 TG_magic_7.B.n22 TG_magic_7.B.n10 0.279866
R4767 TG_magic_7.B.n129 TG_magic_7.B.n117 0.279866
R4768 TG_magic_7.B.n50 TG_magic_7.B.n44 0.244078
R4769 TG_magic_7.B.n157 TG_magic_7.B.n156 0.244078
R4770 TG_magic_7.B.n104 TG_magic_7.B.n86 0.237239
R4771 TG_magic_7.B.n51 TG_magic_7.B.n50 0.1355
R4772 TG_magic_7.B.n158 TG_magic_7.B.n157 0.1355
R4773 TG_magic_7.B TG_magic_7.B.n106 0.1229
R4774 TG_magic_7.B.n106 TG_magic_7.B 0.0749
R4775 S0.n31 S0.t15 68.1773
R4776 S0.n25 S0.t82 68.1773
R4777 S0.n42 S0.n41 52.5344
R4778 S0.n29 S0.n28 52.5344
R4779 S0.n57 S0.n56 52.5344
R4780 S0.n11 S0.n10 52.5344
R4781 S0.n43 S0.t63 47.0594
R4782 S0.n30 S0.t39 47.0594
R4783 S0.n58 S0.t68 47.0594
R4784 S0.n12 S0.t7 47.0594
R4785 S0.t73 S0.t30 43.8005
R4786 S0.t12 S0.t52 43.8005
R4787 S0.t37 S0.t84 43.8005
R4788 S0.t43 S0.t87 43.8005
R4789 S0.t41 S0.t61 43.8005
R4790 S0.t19 S0.t41 43.8005
R4791 S0.t63 S0.t19 43.8005
R4792 S0.t11 S0.t36 43.8005
R4793 S0.t83 S0.t11 43.8005
R4794 S0.t39 S0.t83 43.8005
R4795 S0.t47 S0.t65 43.8005
R4796 S0.t0 S0.t47 43.8005
R4797 S0.t68 S0.t0 43.8005
R4798 S0.t70 S0.t64 43.8005
R4799 S0.t24 S0.t70 43.8005
R4800 S0.t7 S0.t24 43.8005
R4801 S0.t45 S0.n35 33.8934
R4802 S0.n22 S0.t85 33.763
R4803 S0.t42 S0.t21 30.7648
R4804 S0.t55 S0.t44 30.7648
R4805 S0.t78 S0.t57 30.7648
R4806 S0.t38 S0.t17 30.7648
R4807 S0.n13 S0.t42 30.3737
R4808 S0.n14 S0.t55 30.3737
R4809 S0.n15 S0.t78 30.3737
R4810 S0.n40 S0.t13 21.9005
R4811 S0.n40 S0.t56 21.9005
R4812 S0.n39 S0.t60 21.9005
R4813 S0.n39 S0.t18 21.9005
R4814 S0.n38 S0.t49 21.9005
R4815 S0.n38 S0.t5 21.9005
R4816 S0.n37 S0.t34 21.9005
R4817 S0.n37 S0.t81 21.9005
R4818 S0.n36 S0.t86 21.9005
R4819 S0.n36 S0.t45 21.9005
R4820 S0.n21 S0.t40 21.9005
R4821 S0.t85 S0.n21 21.9005
R4822 S0.n20 S0.t2 21.9005
R4823 S0.n20 S0.t46 21.9005
R4824 S0.n19 S0.t74 21.9005
R4825 S0.n19 S0.t31 21.9005
R4826 S0.n18 S0.t29 21.9005
R4827 S0.t75 S0.n18 21.9005
R4828 S0.n27 S0.t14 21.9005
R4829 S0.n27 S0.t58 21.9005
R4830 S0.n48 S0.t79 21.9005
R4831 S0.n48 S0.t33 21.9005
R4832 S0.n50 S0.t59 21.9005
R4833 S0.n50 S0.t16 21.9005
R4834 S0.n52 S0.t32 21.9005
R4835 S0.n52 S0.t76 21.9005
R4836 S0.n54 S0.t69 21.9005
R4837 S0.n54 S0.t26 21.9005
R4838 S0.n55 S0.t8 21.9005
R4839 S0.n55 S0.t50 21.9005
R4840 S0.n9 S0.t51 21.9005
R4841 S0.n9 S0.t67 21.9005
R4842 S0.n8 S0.t4 21.9005
R4843 S0.n8 S0.t20 21.9005
R4844 S0.n7 S0.t54 21.9005
R4845 S0.n7 S0.t77 21.9005
R4846 S0.n6 S0.t10 21.9005
R4847 S0.n6 S0.t27 21.9005
R4848 S0.n5 S0.t9 21.9005
R4849 S0.n5 S0.t80 21.9005
R4850 S0.n13 S0.t73 21.6398
R4851 S0.n14 S0.t12 21.6398
R4852 S0.n15 S0.t37 21.6398
R4853 S0.n16 S0.t43 21.6398
R4854 S0.n32 S0.n31 20.8576
R4855 S0.n33 S0.n32 20.8576
R4856 S0.n34 S0.n33 20.8576
R4857 S0.n35 S0.n34 20.8576
R4858 S0.n23 S0.n22 20.8576
R4859 S0.n24 S0.n23 20.8576
R4860 S0.n26 S0.n24 20.8576
R4861 S0.n26 S0.n25 20.8576
R4862 S0.n47 S0.n46 20.8576
R4863 S0.n1 S0.n0 20.8576
R4864 S0.n41 S0.n40 19.4672
R4865 S0.n28 S0.n27 19.4672
R4866 S0.n56 S0.n55 19.4672
R4867 S0.n10 S0.n9 19.4672
R4868 S0.n43 S0.t53 19.4237
R4869 S0.n30 S0.t35 19.4237
R4870 S0.n58 S0.t25 19.4237
R4871 S0.n12 S0.t23 19.4237
R4872 S0.n42 S0.t15 18.2505
R4873 S0.n41 S0.t72 18.2505
R4874 S0.n41 S0.t28 18.2505
R4875 S0.t53 S0.n42 18.2505
R4876 S0.n29 S0.t82 18.2505
R4877 S0.n28 S0.t22 18.2505
R4878 S0.n28 S0.t62 18.2505
R4879 S0.t35 S0.n29 18.2505
R4880 S0.n56 S0.t48 18.2505
R4881 S0.n57 S0.t66 18.2505
R4882 S0.n56 S0.t3 18.2505
R4883 S0.t25 S0.n57 18.2505
R4884 S0.n10 S0.t1 18.2505
R4885 S0.n11 S0.t6 18.2505
R4886 S0.n10 S0.t71 18.2505
R4887 S0.t23 S0.n11 18.2505
R4888 S0.n17 S0.t38 17.7827
R4889 S0.n14 S0.n13 17.255
R4890 S0.n15 S0.n14 17.255
R4891 S0.n16 S0.n15 17.255
R4892 S0.n40 S0.n39 15.8172
R4893 S0.n39 S0.n38 15.8172
R4894 S0.n38 S0.n37 15.8172
R4895 S0.n37 S0.n36 15.8172
R4896 S0.n21 S0.n20 15.8172
R4897 S0.n20 S0.n19 15.8172
R4898 S0.n19 S0.n18 15.8172
R4899 S0.n27 S0.n18 15.8172
R4900 S0.n50 S0.n48 15.8172
R4901 S0.n52 S0.n50 15.8172
R4902 S0.n54 S0.n52 15.8172
R4903 S0.n55 S0.n54 15.8172
R4904 S0.n9 S0.n8 15.8172
R4905 S0.n8 S0.n7 15.8172
R4906 S0.n7 S0.n6 15.8172
R4907 S0.n6 S0.n5 15.8172
R4908 S0.n32 S0.t56 15.6434
R4909 S0.n33 S0.t18 15.6434
R4910 S0.n34 S0.t5 15.6434
R4911 S0.n35 S0.t81 15.6434
R4912 S0.n31 S0.t72 15.6434
R4913 S0.n22 S0.t46 15.6434
R4914 S0.n23 S0.t31 15.6434
R4915 S0.n24 S0.t75 15.6434
R4916 S0.t58 S0.n26 15.6434
R4917 S0.n25 S0.t22 15.6434
R4918 S0.t59 S0.n49 15.6434
R4919 S0.t32 S0.n51 15.6434
R4920 S0.t69 S0.n53 15.6434
R4921 S0.t3 S0.n47 15.6434
R4922 S0.t4 S0.n2 15.6434
R4923 S0.t54 S0.n3 15.6434
R4924 S0.t10 S0.n4 15.6434
R4925 S0.t71 S0.n1 15.6434
R4926 S0.n44 S0 14.8438
R4927 S0 S0.n30 8.63236
R4928 S0 S0.n12 8.63236
R4929 S0 S0.n43 8.63011
R4930 S0.n59 S0.n58 8.59261
R4931 S0.n60 S0.n59 8.2322
R4932 S0.n17 S0.n16 8.06475
R4933 S0.n60 S0.n45 7.19405
R4934 S0 S0.n17 4.24369
R4935 S0 S0.n44 2.56189
R4936 S0 S0.n60 0.485265
R4937 S0.n44 S0 0.440704
R4938 S0.n45 S0 0.247147
R4939 S0.n45 S0 0.182052
R4940 S0.n59 S0 0.00343915
R4941 a_5684_n6152.t8 a_5684_n6152.n10 40.7345
R4942 a_5684_n6152.n19 a_5684_n6152.n18 28.094
R4943 a_5684_n6152.n12 a_5684_n6152.n11 28.094
R4944 a_5684_n6152.n27 a_5684_n6152.n26 28.094
R4945 a_5684_n6152.n26 a_5684_n6152.t11 21.9005
R4946 a_5684_n6152.n11 a_5684_n6152.t8 21.9005
R4947 a_5684_n6152.n2 a_5684_n6152.t29 21.9005
R4948 a_5684_n6152.n21 a_5684_n6152.t9 21.9005
R4949 a_5684_n6152.n21 a_5684_n6152.t20 21.9005
R4950 a_5684_n6152.n13 a_5684_n6152.t27 21.9005
R4951 a_5684_n6152.n14 a_5684_n6152.t21 21.9005
R4952 a_5684_n6152.n22 a_5684_n6152.t15 21.9005
R4953 a_5684_n6152.n22 a_5684_n6152.t28 21.9005
R4954 a_5684_n6152.n3 a_5684_n6152.t22 21.9005
R4955 a_5684_n6152.n4 a_5684_n6152.t14 21.9005
R4956 a_5684_n6152.n23 a_5684_n6152.t17 21.9005
R4957 a_5684_n6152.n23 a_5684_n6152.t10 21.9005
R4958 a_5684_n6152.n15 a_5684_n6152.t13 21.9005
R4959 a_5684_n6152.n16 a_5684_n6152.t24 21.9005
R4960 a_5684_n6152.n24 a_5684_n6152.t16 21.9005
R4961 a_5684_n6152.n24 a_5684_n6152.t6 21.9005
R4962 a_5684_n6152.n5 a_5684_n6152.t26 21.9005
R4963 a_5684_n6152.n6 a_5684_n6152.t19 21.9005
R4964 a_5684_n6152.n25 a_5684_n6152.t25 21.9005
R4965 a_5684_n6152.n25 a_5684_n6152.t12 21.9005
R4966 a_5684_n6152.n17 a_5684_n6152.t18 21.9005
R4967 a_5684_n6152.n18 a_5684_n6152.t7 21.9005
R4968 a_5684_n6152.n26 a_5684_n6152.t23 21.9005
R4969 a_5684_n6152.n26 a_5684_n6152.n25 15.8172
R4970 a_5684_n6152.n11 a_5684_n6152.n6 15.8172
R4971 a_5684_n6152.n6 a_5684_n6152.n5 15.8172
R4972 a_5684_n6152.n25 a_5684_n6152.n24 15.8172
R4973 a_5684_n6152.n24 a_5684_n6152.n23 15.8172
R4974 a_5684_n6152.n5 a_5684_n6152.n4 15.8172
R4975 a_5684_n6152.n4 a_5684_n6152.n3 15.8172
R4976 a_5684_n6152.n23 a_5684_n6152.n22 15.8172
R4977 a_5684_n6152.n22 a_5684_n6152.n21 15.8172
R4978 a_5684_n6152.n3 a_5684_n6152.n2 15.8172
R4979 a_5684_n6152.n14 a_5684_n6152.n13 15.8172
R4980 a_5684_n6152.n15 a_5684_n6152.n14 15.8172
R4981 a_5684_n6152.n16 a_5684_n6152.n15 15.8172
R4982 a_5684_n6152.n17 a_5684_n6152.n16 15.8172
R4983 a_5684_n6152.n18 a_5684_n6152.n17 15.8172
R4984 a_5684_n6152.n8 a_5684_n6152.n7 15.1845
R4985 a_5684_n6152.n9 a_5684_n6152.n8 15.1845
R4986 a_5684_n6152.n10 a_5684_n6152.n9 15.1845
R4987 a_5684_n6152.n0 a_5684_n6152.t4 5.44589
R4988 a_5684_n6152.n0 a_5684_n6152.t5 4.7885
R4989 a_5684_n6152.n19 a_5684_n6152.t1 4.70615
R4990 a_5684_n6152.n1 a_5684_n6152.t0 4.4205
R4991 a_5684_n6152.n20 a_5684_n6152.t2 4.4205
R4992 a_5684_n6152.t3 a_5684_n6152.n28 4.4205
R4993 a_5684_n6152.n1 a_5684_n6152.n0 1.1392
R4994 a_5684_n6152.n27 a_5684_n6152.n20 0.286152
R4995 a_5684_n6152.n28 a_5684_n6152.n12 0.286152
R4996 a_5684_n6152.n12 a_5684_n6152.n1 0.282239
R4997 a_5684_n6152.n20 a_5684_n6152.n19 0.282239
R4998 a_5684_n6152.n28 a_5684_n6152.n27 0.282239
R4999 a_301_308.t24 a_301_308.n22 40.7345
R5000 a_301_308.n24 a_301_308.n23 28.094
R5001 a_301_308.n7 a_301_308.n6 28.094
R5002 a_301_308.n32 a_301_308.n31 28.094
R5003 a_301_308.n4 a_301_308.t14 21.9005
R5004 a_301_308.n2 a_301_308.t6 21.9005
R5005 a_301_308.n1 a_301_308.t25 21.9005
R5006 a_301_308.n1 a_301_308.t18 21.9005
R5007 a_301_308.n26 a_301_308.t13 21.9005
R5008 a_301_308.n14 a_301_308.t26 21.9005
R5009 a_301_308.n15 a_301_308.t7 21.9005
R5010 a_301_308.n27 a_301_308.t20 21.9005
R5011 a_301_308.n2 a_301_308.t23 21.9005
R5012 a_301_308.n3 a_301_308.t8 21.9005
R5013 a_301_308.n3 a_301_308.t27 21.9005
R5014 a_301_308.n28 a_301_308.t21 21.9005
R5015 a_301_308.n16 a_301_308.t10 21.9005
R5016 a_301_308.n17 a_301_308.t15 21.9005
R5017 a_301_308.n29 a_301_308.t28 21.9005
R5018 a_301_308.n4 a_301_308.t9 21.9005
R5019 a_301_308.n6 a_301_308.t22 21.9005
R5020 a_301_308.n6 a_301_308.t16 21.9005
R5021 a_301_308.n5 a_301_308.t17 21.9005
R5022 a_301_308.n5 a_301_308.t11 21.9005
R5023 a_301_308.n30 a_301_308.t29 21.9005
R5024 a_301_308.n18 a_301_308.t19 21.9005
R5025 a_301_308.n23 a_301_308.t24 21.9005
R5026 a_301_308.n31 a_301_308.t12 21.9005
R5027 a_301_308.n23 a_301_308.n18 15.8172
R5028 a_301_308.n31 a_301_308.n30 15.8172
R5029 a_301_308.n30 a_301_308.n29 15.8172
R5030 a_301_308.n18 a_301_308.n17 15.8172
R5031 a_301_308.n17 a_301_308.n16 15.8172
R5032 a_301_308.n29 a_301_308.n28 15.8172
R5033 a_301_308.n28 a_301_308.n27 15.8172
R5034 a_301_308.n16 a_301_308.n15 15.8172
R5035 a_301_308.n15 a_301_308.n14 15.8172
R5036 a_301_308.n27 a_301_308.n26 15.8172
R5037 a_301_308.n2 a_301_308.n1 15.8172
R5038 a_301_308.n4 a_301_308.n3 15.8172
R5039 a_301_308.n3 a_301_308.n2 15.8172
R5040 a_301_308.n6 a_301_308.n5 15.8172
R5041 a_301_308.n5 a_301_308.n4 15.8172
R5042 a_301_308.n20 a_301_308.n19 15.1845
R5043 a_301_308.n22 a_301_308.n21 15.1845
R5044 a_301_308.n21 a_301_308.n20 15.1845
R5045 a_301_308.n12 a_301_308.n11 5.44589
R5046 a_301_308.n12 a_301_308.n10 4.7885
R5047 a_301_308.n7 a_301_308.n0 4.70615
R5048 a_301_308.n13 a_301_308.n9 4.4205
R5049 a_301_308.n25 a_301_308.n8 4.4205
R5050 a_301_308.n34 a_301_308.n33 4.4205
R5051 a_301_308.n13 a_301_308.n12 1.1392
R5052 a_301_308.n25 a_301_308.n24 0.286152
R5053 a_301_308.n33 a_301_308.n32 0.286152
R5054 a_301_308.n32 a_301_308.n25 0.282239
R5055 a_301_308.n24 a_301_308.n13 0.282239
R5056 a_301_308.n33 a_301_308.n7 0.282239
R5057 a_n4297_300.t9 a_n4297_300.n30 40.7345
R5058 a_n4297_300.n7 a_n4297_300.n6 28.094
R5059 a_n4297_300.n16 a_n4297_300.n15 28.094
R5060 a_n4297_300.n32 a_n4297_300.n31 28.094
R5061 a_n4297_300.n4 a_n4297_300.t15 21.9005
R5062 a_n4297_300.n2 a_n4297_300.t24 21.9005
R5063 a_n4297_300.n1 a_n4297_300.t29 21.9005
R5064 a_n4297_300.n10 a_n4297_300.t28 21.9005
R5065 a_n4297_300.n10 a_n4297_300.t18 21.9005
R5066 a_n4297_300.n22 a_n4297_300.t6 21.9005
R5067 a_n4297_300.n23 a_n4297_300.t25 21.9005
R5068 a_n4297_300.n11 a_n4297_300.t11 21.9005
R5069 a_n4297_300.n11 a_n4297_300.t23 21.9005
R5070 a_n4297_300.n3 a_n4297_300.t20 21.9005
R5071 a_n4297_300.n12 a_n4297_300.t21 21.9005
R5072 a_n4297_300.n12 a_n4297_300.t10 21.9005
R5073 a_n4297_300.n24 a_n4297_300.t22 21.9005
R5074 a_n4297_300.n25 a_n4297_300.t17 21.9005
R5075 a_n4297_300.n13 a_n4297_300.t27 21.9005
R5076 a_n4297_300.n13 a_n4297_300.t16 21.9005
R5077 a_n4297_300.n6 a_n4297_300.t8 21.9005
R5078 a_n4297_300.n15 a_n4297_300.t19 21.9005
R5079 a_n4297_300.n15 a_n4297_300.t7 21.9005
R5080 a_n4297_300.n5 a_n4297_300.t13 21.9005
R5081 a_n4297_300.n14 a_n4297_300.t12 21.9005
R5082 a_n4297_300.n14 a_n4297_300.t26 21.9005
R5083 a_n4297_300.n26 a_n4297_300.t14 21.9005
R5084 a_n4297_300.n31 a_n4297_300.t9 21.9005
R5085 a_n4297_300.n31 a_n4297_300.n26 15.8172
R5086 a_n4297_300.n14 a_n4297_300.n13 15.8172
R5087 a_n4297_300.n26 a_n4297_300.n25 15.8172
R5088 a_n4297_300.n25 a_n4297_300.n24 15.8172
R5089 a_n4297_300.n13 a_n4297_300.n12 15.8172
R5090 a_n4297_300.n12 a_n4297_300.n11 15.8172
R5091 a_n4297_300.n24 a_n4297_300.n23 15.8172
R5092 a_n4297_300.n23 a_n4297_300.n22 15.8172
R5093 a_n4297_300.n11 a_n4297_300.n10 15.8172
R5094 a_n4297_300.n2 a_n4297_300.n1 15.8172
R5095 a_n4297_300.n4 a_n4297_300.n3 15.8172
R5096 a_n4297_300.n3 a_n4297_300.n2 15.8172
R5097 a_n4297_300.n15 a_n4297_300.n14 15.8172
R5098 a_n4297_300.n6 a_n4297_300.n5 15.8172
R5099 a_n4297_300.n5 a_n4297_300.n4 15.8172
R5100 a_n4297_300.n28 a_n4297_300.n27 15.1845
R5101 a_n4297_300.n30 a_n4297_300.n29 15.1845
R5102 a_n4297_300.n29 a_n4297_300.n28 15.1845
R5103 a_n4297_300.n20 a_n4297_300.n19 5.44589
R5104 a_n4297_300.n20 a_n4297_300.n18 4.7885
R5105 a_n4297_300.n7 a_n4297_300.n0 4.70615
R5106 a_n4297_300.n21 a_n4297_300.n17 4.4205
R5107 a_n4297_300.n9 a_n4297_300.n8 4.4205
R5108 a_n4297_300.n34 a_n4297_300.n33 4.4205
R5109 a_n4297_300.n21 a_n4297_300.n20 1.1392
R5110 a_n4297_300.n16 a_n4297_300.n9 0.286152
R5111 a_n4297_300.n33 a_n4297_300.n32 0.286152
R5112 a_n4297_300.n32 a_n4297_300.n21 0.282239
R5113 a_n4297_300.n9 a_n4297_300.n7 0.282239
R5114 a_n4297_300.n33 a_n4297_300.n16 0.282239
R5115 A6.n47 A6.n45 5.44589
R5116 A6.n26 A6.n25 5.07789
R5117 A6.n51 A6.t5 4.7885
R5118 A6.n50 A6.t8 4.7885
R5119 A6.n47 A6.n46 4.7885
R5120 A6.n31 A6.t33 4.4205
R5121 A6.n32 A6.t34 4.4205
R5122 A6.n33 A6.t22 4.4205
R5123 A6.n34 A6.t32 4.4205
R5124 A6.n28 A6.n22 4.4205
R5125 A6.n27 A6.n23 4.4205
R5126 A6.n26 A6.n24 4.4205
R5127 A6.n44 A6.n41 3.80789
R5128 A6.n39 A6.n36 3.80789
R5129 A6.n8 A6.n7 3.25789
R5130 A6.n19 A6.n18 3.25789
R5131 A6.n44 A6.n43 3.1505
R5132 A6.n39 A6.n38 3.1505
R5133 A6.n8 A6.n5 2.6005
R5134 A6.n9 A6.n3 2.6005
R5135 A6.n10 A6.n1 2.6005
R5136 A6.n19 A6.n16 2.6005
R5137 A6.n20 A6.n14 2.6005
R5138 A6.n21 A6.n12 2.6005
R5139 A6.n1 A6.t26 1.8205
R5140 A6.n1 A6.n0 1.8205
R5141 A6.n3 A6.t25 1.8205
R5142 A6.n3 A6.n2 1.8205
R5143 A6.n5 A6.t14 1.8205
R5144 A6.n5 A6.n4 1.8205
R5145 A6.n7 A6.t24 1.8205
R5146 A6.n7 A6.n6 1.8205
R5147 A6.n12 A6.t17 1.8205
R5148 A6.n12 A6.n11 1.8205
R5149 A6.n14 A6.t18 1.8205
R5150 A6.n14 A6.n13 1.8205
R5151 A6.n16 A6.t30 1.8205
R5152 A6.n16 A6.n15 1.8205
R5153 A6.n18 A6.t16 1.8205
R5154 A6.n18 A6.n17 1.8205
R5155 A6.n43 A6.t10 1.6385
R5156 A6.n43 A6.n42 1.6385
R5157 A6.n41 A6.t7 1.6385
R5158 A6.n41 A6.n40 1.6385
R5159 A6.n38 A6.t3 1.6385
R5160 A6.n38 A6.n37 1.6385
R5161 A6.n36 A6.t0 1.6385
R5162 A6.n36 A6.n35 1.6385
R5163 A6 A6.n52 1.54844
R5164 A6.n48 A6.n47 0.884196
R5165 A6.n50 A6.n49 0.884196
R5166 A6.n29 A6.n28 0.882239
R5167 A6.n31 A6.n30 0.882239
R5168 A6.n10 A6.n9 0.657891
R5169 A6.n9 A6.n8 0.657891
R5170 A6.n21 A6.n20 0.657891
R5171 A6.n20 A6.n19 0.657891
R5172 A6.n28 A6.n27 0.657891
R5173 A6.n27 A6.n26 0.657891
R5174 A6.n32 A6.n31 0.657891
R5175 A6.n33 A6.n32 0.657891
R5176 A6.n34 A6.n33 0.657891
R5177 A6.n51 A6.n50 0.657891
R5178 A6.n52 A6.n51 0.600532
R5179 A6.n30 A6.n29 0.6005
R5180 A6.n49 A6.n48 0.6005
R5181 A6.n48 A6.n44 0.284196
R5182 A6.n49 A6.n39 0.284196
R5183 A6.n30 A6.n10 0.282239
R5184 A6.n29 A6.n21 0.282239
R5185 A6.n52 A6.n34 0.278258
R5186 ENA.n4 ENA.t27 44.713
R5187 ENA.n3 ENA.t46 44.713
R5188 ENA.n0 ENA.t19 44.713
R5189 ENA.n14 ENA.t14 44.713
R5190 ENA.n24 ENA.t1 44.713
R5191 ENA.n27 ENA.t32 44.713
R5192 ENA.n37 ENA.t37 44.713
R5193 ENA.n45 ENA.t40 44.713
R5194 ENA.t45 ENA.t22 43.8005
R5195 ENA.t8 ENA.t24 43.8005
R5196 ENA.t0 ENA.t8 43.8005
R5197 ENA.t27 ENA.t0 43.8005
R5198 ENA.t3 ENA.t44 43.8005
R5199 ENA.t42 ENA.t43 43.8005
R5200 ENA.t20 ENA.t42 43.8005
R5201 ENA.t46 ENA.t20 43.8005
R5202 ENA.t5 ENA.t17 43.8005
R5203 ENA.t30 ENA.t5 43.8005
R5204 ENA.t19 ENA.t30 43.8005
R5205 ENA.t16 ENA.t6 43.8005
R5206 ENA.t38 ENA.t11 43.8005
R5207 ENA.t25 ENA.t38 43.8005
R5208 ENA.t14 ENA.t25 43.8005
R5209 ENA.t41 ENA.t18 43.8005
R5210 ENA.t26 ENA.t34 43.8005
R5211 ENA.t15 ENA.t2 43.8005
R5212 ENA.t28 ENA.t15 43.8005
R5213 ENA.t1 ENA.t28 43.8005
R5214 ENA.t7 ENA.t31 43.8005
R5215 ENA.t10 ENA.t33 43.8005
R5216 ENA.t21 ENA.t10 43.8005
R5217 ENA.t32 ENA.t21 43.8005
R5218 ENA.t23 ENA.t35 43.8005
R5219 ENA.t47 ENA.t23 43.8005
R5220 ENA.t37 ENA.t47 43.8005
R5221 ENA.t9 ENA.t36 43.8005
R5222 ENA.t29 ENA.t39 43.8005
R5223 ENA.t13 ENA.t29 43.8005
R5224 ENA.t40 ENA.t13 43.8005
R5225 ENA.t12 ENA.t4 43.8005
R5226 ENA.n4 ENA.t45 20.7273
R5227 ENA.n3 ENA.t3 20.7273
R5228 ENA.n0 ENA.t16 20.7273
R5229 ENA.n14 ENA.t41 20.7273
R5230 ENA.n24 ENA.t26 20.7273
R5231 ENA.n27 ENA.t7 20.7273
R5232 ENA.n37 ENA.t9 20.7273
R5233 ENA.n45 ENA.t12 20.7273
R5234 ENA ENA.n13 8.0005
R5235 ENA.n25 ENA.n24 6.09337
R5236 ENA.n8 ENA.n3 6.04485
R5237 ENA.n5 ENA.n4 6.0288
R5238 ENA.n47 ENA.n45 5.80834
R5239 ENA.n15 ENA.n14 5.6366
R5240 ENA.n28 ENA.n27 5.07708
R5241 ENA.n38 ENA.n37 5.07708
R5242 ENA.n1 ENA.n0 5.07642
R5243 ENA ENA.n55 4.89473
R5244 ENA.n11 ENA.n10 4.5005
R5245 ENA.n8 ENA.n7 4.5005
R5246 ENA.n17 ENA.n13 4.5005
R5247 ENA.n18 ENA.n17 3.36698
R5248 ENA.n20 ENA.n19 3.11702
R5249 ENA.n47 ENA.n46 2.97306
R5250 ENA.n41 ENA.n36 2.81699
R5251 ENA.n32 ENA.n31 2.66698
R5252 ENA.n33 ENA.n32 2.58104
R5253 ENA.n42 ENA.n41 2.57371
R5254 ENA.n12 ENA.n11 2.37035
R5255 ENA.n6 ENA 2.28422
R5256 ENA.n7 ENA.n6 2.27686
R5257 ENA.n52 ENA.n44 2.26755
R5258 ENA.n53 ENA.n35 2.26592
R5259 ENA.n9 ENA.n2 2.2505
R5260 ENA.n34 ENA 2.2505
R5261 ENA.n53 ENA.n52 2.08841
R5262 ENA ENA.n12 1.27356
R5263 ENA.n6 ENA.n5 1.19179
R5264 ENA.n21 ENA.n1 1.05063
R5265 ENA.n40 ENA.n38 1.04974
R5266 ENA.n30 ENA.n28 1.04299
R5267 ENA.n18 ENA 0.954762
R5268 ENA.n55 ENA.n54 0.593375
R5269 ENA.n16 ENA.n15 0.406055
R5270 ENA.n49 ENA.n47 0.263268
R5271 ENA.n52 ENA.n51 0.104841
R5272 ENA.n54 ENA.n26 0.068
R5273 ENA.n20 ENA.n18 0.0430568
R5274 ENA ENA.n5 0.0381415
R5275 ENA.n26 ENA.n25 0.026375
R5276 ENA.n54 ENA.n53 0.02525
R5277 ENA.n51 ENA.n50 0.0237418
R5278 ENA.n34 ENA.n33 0.01925
R5279 ENA.n11 ENA.n2 0.0167931
R5280 ENA.n10 ENA.n9 0.0159918
R5281 ENA.n16 ENA 0.0159545
R5282 ENA.n43 ENA.n42 0.01475
R5283 ENA.n50 ENA.n49 0.0133571
R5284 ENA.n39 ENA 0.0127255
R5285 ENA.n10 ENA 0.0115656
R5286 ENA.n40 ENA.n39 0.0114212
R5287 ENA.n29 ENA 0.0111893
R5288 ENA.n30 ENA.n29 0.0111847
R5289 ENA.n49 ENA.n48 0.0108228
R5290 ENA ENA.n22 0.00999612
R5291 ENA.n41 ENA.n40 0.00963044
R5292 ENA.n21 ENA.n20 0.00907143
R5293 ENA.n48 ENA 0.00787592
R5294 ENA.n22 ENA.n21 0.00656755
R5295 ENA.n17 ENA.n16 0.00595455
R5296 ENA.n7 ENA.n2 0.00593103
R5297 ENA.n9 ENA.n8 0.00566393
R5298 ENA.n12 ENA 0.00566393
R5299 ENA.n44 ENA.n43 0.005
R5300 ENA.n55 ENA.n23 0.005
R5301 ENA.n32 ENA.n30 0.0041
R5302 ENA ENA.n23 0.003875
R5303 ENA.n35 ENA.n34 0.00275
R5304 ENA ENA.n26 0.00275
R5305 a_2061_n4852.t24 a_2061_n4852.n27 40.7345
R5306 a_2061_n4852.n7 a_2061_n4852.n6 28.094
R5307 a_2061_n4852.n16 a_2061_n4852.n15 28.094
R5308 a_2061_n4852.n29 a_2061_n4852.n28 28.094
R5309 a_2061_n4852.n4 a_2061_n4852.t9 21.9005
R5310 a_2061_n4852.n2 a_2061_n4852.t11 21.9005
R5311 a_2061_n4852.n1 a_2061_n4852.t29 21.9005
R5312 a_2061_n4852.n10 a_2061_n4852.t18 21.9005
R5313 a_2061_n4852.n19 a_2061_n4852.t21 21.9005
R5314 a_2061_n4852.n19 a_2061_n4852.t28 21.9005
R5315 a_2061_n4852.n20 a_2061_n4852.t10 21.9005
R5316 a_2061_n4852.n20 a_2061_n4852.t27 21.9005
R5317 a_2061_n4852.n11 a_2061_n4852.t22 21.9005
R5318 a_2061_n4852.n3 a_2061_n4852.t17 21.9005
R5319 a_2061_n4852.n12 a_2061_n4852.t8 21.9005
R5320 a_2061_n4852.n21 a_2061_n4852.t12 21.9005
R5321 a_2061_n4852.n21 a_2061_n4852.t16 21.9005
R5322 a_2061_n4852.n22 a_2061_n4852.t7 21.9005
R5323 a_2061_n4852.n22 a_2061_n4852.t23 21.9005
R5324 a_2061_n4852.n13 a_2061_n4852.t20 21.9005
R5325 a_2061_n4852.n6 a_2061_n4852.t26 21.9005
R5326 a_2061_n4852.n28 a_2061_n4852.t19 21.9005
R5327 a_2061_n4852.n15 a_2061_n4852.t15 21.9005
R5328 a_2061_n4852.n5 a_2061_n4852.t14 21.9005
R5329 a_2061_n4852.n14 a_2061_n4852.t25 21.9005
R5330 a_2061_n4852.n23 a_2061_n4852.t6 21.9005
R5331 a_2061_n4852.n23 a_2061_n4852.t13 21.9005
R5332 a_2061_n4852.n28 a_2061_n4852.t24 21.9005
R5333 a_2061_n4852.n28 a_2061_n4852.n23 15.8172
R5334 a_2061_n4852.n14 a_2061_n4852.n13 15.8172
R5335 a_2061_n4852.n23 a_2061_n4852.n22 15.8172
R5336 a_2061_n4852.n22 a_2061_n4852.n21 15.8172
R5337 a_2061_n4852.n13 a_2061_n4852.n12 15.8172
R5338 a_2061_n4852.n12 a_2061_n4852.n11 15.8172
R5339 a_2061_n4852.n21 a_2061_n4852.n20 15.8172
R5340 a_2061_n4852.n20 a_2061_n4852.n19 15.8172
R5341 a_2061_n4852.n11 a_2061_n4852.n10 15.8172
R5342 a_2061_n4852.n2 a_2061_n4852.n1 15.8172
R5343 a_2061_n4852.n4 a_2061_n4852.n3 15.8172
R5344 a_2061_n4852.n3 a_2061_n4852.n2 15.8172
R5345 a_2061_n4852.n15 a_2061_n4852.n14 15.8172
R5346 a_2061_n4852.n6 a_2061_n4852.n5 15.8172
R5347 a_2061_n4852.n5 a_2061_n4852.n4 15.8172
R5348 a_2061_n4852.n25 a_2061_n4852.n24 15.1845
R5349 a_2061_n4852.n27 a_2061_n4852.n26 15.1845
R5350 a_2061_n4852.n26 a_2061_n4852.n25 15.1845
R5351 a_2061_n4852.n32 a_2061_n4852.n31 5.44589
R5352 a_2061_n4852.n32 a_2061_n4852.n30 4.7885
R5353 a_2061_n4852.n7 a_2061_n4852.n0 4.70615
R5354 a_2061_n4852.n18 a_2061_n4852.n17 4.4205
R5355 a_2061_n4852.n9 a_2061_n4852.n8 4.4205
R5356 a_2061_n4852.n34 a_2061_n4852.n33 4.4205
R5357 a_2061_n4852.n33 a_2061_n4852.n32 1.1392
R5358 a_2061_n4852.n16 a_2061_n4852.n9 0.286152
R5359 a_2061_n4852.n29 a_2061_n4852.n18 0.286152
R5360 a_2061_n4852.n9 a_2061_n4852.n7 0.282239
R5361 a_2061_n4852.n18 a_2061_n4852.n16 0.282239
R5362 a_2061_n4852.n33 a_2061_n4852.n29 0.282239
R5363 TG_magic_2.B.n104 TG_magic_2.B.t99 5.44589
R5364 TG_magic_2.B.n155 TG_magic_2.B 5.33254
R5365 TG_magic_2.B.n142 TG_magic_2.B.t62 5.07789
R5366 TG_magic_2.B.n157 TG_magic_2.B.n156 4.7885
R5367 TG_magic_2.B.n159 TG_magic_2.B.n158 4.7885
R5368 TG_magic_2.B.n104 TG_magic_2.B.t105 4.7885
R5369 TG_magic_2.B.n148 TG_magic_2.B.n147 4.4205
R5370 TG_magic_2.B.n150 TG_magic_2.B.n149 4.4205
R5371 TG_magic_2.B.n152 TG_magic_2.B.n151 4.4205
R5372 TG_magic_2.B.n154 TG_magic_2.B.n153 4.4205
R5373 TG_magic_2.B.n144 TG_magic_2.B.t15 4.4205
R5374 TG_magic_2.B.n143 TG_magic_2.B.t29 4.4205
R5375 TG_magic_2.B.n142 TG_magic_2.B.t34 4.4205
R5376 TG_magic_2.B.n79 TG_magic_2.B.n76 3.80789
R5377 TG_magic_2.B.n84 TG_magic_2.B.n81 3.80789
R5378 TG_magic_2.B.n89 TG_magic_2.B.n86 3.80789
R5379 TG_magic_2.B.n117 TG_magic_2.B.n114 3.80789
R5380 TG_magic_2.B.n110 TG_magic_2.B.n107 3.80789
R5381 TG_magic_2.B.n9 TG_magic_2.B.n6 3.80789
R5382 TG_magic_2.B.n4 TG_magic_2.B.n1 3.80789
R5383 TG_magic_2.B.n15 TG_magic_2.B.n12 3.80789
R5384 TG_magic_2.B.n71 TG_magic_2.B.n70 3.25789
R5385 TG_magic_2.B.n60 TG_magic_2.B.n59 3.25789
R5386 TG_magic_2.B.n100 TG_magic_2.B.n99 3.25789
R5387 TG_magic_2.B.n139 TG_magic_2.B.n138 3.25789
R5388 TG_magic_2.B.n128 TG_magic_2.B.n127 3.25789
R5389 TG_magic_2.B.n25 TG_magic_2.B.n24 3.25789
R5390 TG_magic_2.B.n36 TG_magic_2.B.n35 3.25789
R5391 TG_magic_2.B.n45 TG_magic_2.B.n44 3.25789
R5392 TG_magic_2.B.n79 TG_magic_2.B.n78 3.1505
R5393 TG_magic_2.B.n84 TG_magic_2.B.n83 3.1505
R5394 TG_magic_2.B.n89 TG_magic_2.B.n88 3.1505
R5395 TG_magic_2.B.n117 TG_magic_2.B.n116 3.1505
R5396 TG_magic_2.B.n110 TG_magic_2.B.n109 3.1505
R5397 TG_magic_2.B.n9 TG_magic_2.B.n8 3.1505
R5398 TG_magic_2.B.n4 TG_magic_2.B.n3 3.1505
R5399 TG_magic_2.B.n15 TG_magic_2.B.n14 3.1505
R5400 TG_magic_2.B.n164 TG_magic_2.B.n163 2.88408
R5401 TG_magic_2.B.n112 TG_magic_2.B.n105 2.70652
R5402 TG_magic_2.B.n71 TG_magic_2.B.n68 2.6005
R5403 TG_magic_2.B.n72 TG_magic_2.B.n66 2.6005
R5404 TG_magic_2.B.n73 TG_magic_2.B.n64 2.6005
R5405 TG_magic_2.B.n60 TG_magic_2.B.n57 2.6005
R5406 TG_magic_2.B.n61 TG_magic_2.B.n55 2.6005
R5407 TG_magic_2.B.n62 TG_magic_2.B.n53 2.6005
R5408 TG_magic_2.B.n100 TG_magic_2.B.n97 2.6005
R5409 TG_magic_2.B.n101 TG_magic_2.B.n95 2.6005
R5410 TG_magic_2.B.n102 TG_magic_2.B.n93 2.6005
R5411 TG_magic_2.B.n139 TG_magic_2.B.n136 2.6005
R5412 TG_magic_2.B.n140 TG_magic_2.B.n134 2.6005
R5413 TG_magic_2.B.n141 TG_magic_2.B.n132 2.6005
R5414 TG_magic_2.B.n128 TG_magic_2.B.n125 2.6005
R5415 TG_magic_2.B.n129 TG_magic_2.B.n123 2.6005
R5416 TG_magic_2.B.n130 TG_magic_2.B.n121 2.6005
R5417 TG_magic_2.B.n25 TG_magic_2.B.n22 2.6005
R5418 TG_magic_2.B.n26 TG_magic_2.B.n20 2.6005
R5419 TG_magic_2.B.n27 TG_magic_2.B.n18 2.6005
R5420 TG_magic_2.B.n36 TG_magic_2.B.n33 2.6005
R5421 TG_magic_2.B.n37 TG_magic_2.B.n31 2.6005
R5422 TG_magic_2.B.n38 TG_magic_2.B.n29 2.6005
R5423 TG_magic_2.B.n45 TG_magic_2.B.n42 2.6005
R5424 TG_magic_2.B.n49 TG_magic_2.B.n40 2.6005
R5425 TG_magic_2.B.n48 TG_magic_2.B.n47 2.6005
R5426 TG_magic_2.B.n112 TG_magic_2.B.n111 2.2505
R5427 TG_magic_2.B.n119 TG_magic_2.B.n118 2.2505
R5428 TG_magic_2.B.n163 TG_magic_2.B.n162 2.2505
R5429 TG_magic_2.B.n40 TG_magic_2.B.t38 1.8205
R5430 TG_magic_2.B.n40 TG_magic_2.B.n39 1.8205
R5431 TG_magic_2.B.n42 TG_magic_2.B.t48 1.8205
R5432 TG_magic_2.B.n42 TG_magic_2.B.n41 1.8205
R5433 TG_magic_2.B.n44 TG_magic_2.B.t40 1.8205
R5434 TG_magic_2.B.n44 TG_magic_2.B.n43 1.8205
R5435 TG_magic_2.B.n64 TG_magic_2.B.t13 1.8205
R5436 TG_magic_2.B.n64 TG_magic_2.B.n63 1.8205
R5437 TG_magic_2.B.n66 TG_magic_2.B.t95 1.8205
R5438 TG_magic_2.B.n66 TG_magic_2.B.n65 1.8205
R5439 TG_magic_2.B.n68 TG_magic_2.B.t81 1.8205
R5440 TG_magic_2.B.n68 TG_magic_2.B.n67 1.8205
R5441 TG_magic_2.B.n70 TG_magic_2.B.t78 1.8205
R5442 TG_magic_2.B.n70 TG_magic_2.B.n69 1.8205
R5443 TG_magic_2.B.n53 TG_magic_2.B.t77 1.8205
R5444 TG_magic_2.B.n53 TG_magic_2.B.n52 1.8205
R5445 TG_magic_2.B.n55 TG_magic_2.B.t84 1.8205
R5446 TG_magic_2.B.n55 TG_magic_2.B.n54 1.8205
R5447 TG_magic_2.B.n57 TG_magic_2.B.t90 1.8205
R5448 TG_magic_2.B.n57 TG_magic_2.B.n56 1.8205
R5449 TG_magic_2.B.n59 TG_magic_2.B.t88 1.8205
R5450 TG_magic_2.B.n59 TG_magic_2.B.n58 1.8205
R5451 TG_magic_2.B.n93 TG_magic_2.B.t79 1.8205
R5452 TG_magic_2.B.n93 TG_magic_2.B.n92 1.8205
R5453 TG_magic_2.B.n95 TG_magic_2.B.t75 1.8205
R5454 TG_magic_2.B.n95 TG_magic_2.B.n94 1.8205
R5455 TG_magic_2.B.n97 TG_magic_2.B.t92 1.8205
R5456 TG_magic_2.B.n97 TG_magic_2.B.n96 1.8205
R5457 TG_magic_2.B.n99 TG_magic_2.B.t91 1.8205
R5458 TG_magic_2.B.n99 TG_magic_2.B.n98 1.8205
R5459 TG_magic_2.B.n132 TG_magic_2.B.t19 1.8205
R5460 TG_magic_2.B.n132 TG_magic_2.B.n131 1.8205
R5461 TG_magic_2.B.n134 TG_magic_2.B.t32 1.8205
R5462 TG_magic_2.B.n134 TG_magic_2.B.n133 1.8205
R5463 TG_magic_2.B.n136 TG_magic_2.B.t59 1.8205
R5464 TG_magic_2.B.n136 TG_magic_2.B.n135 1.8205
R5465 TG_magic_2.B.n138 TG_magic_2.B.t17 1.8205
R5466 TG_magic_2.B.n138 TG_magic_2.B.n137 1.8205
R5467 TG_magic_2.B.n121 TG_magic_2.B.t25 1.8205
R5468 TG_magic_2.B.n121 TG_magic_2.B.n120 1.8205
R5469 TG_magic_2.B.n123 TG_magic_2.B.t61 1.8205
R5470 TG_magic_2.B.n123 TG_magic_2.B.n122 1.8205
R5471 TG_magic_2.B.n125 TG_magic_2.B.t16 1.8205
R5472 TG_magic_2.B.n125 TG_magic_2.B.n124 1.8205
R5473 TG_magic_2.B.n127 TG_magic_2.B.t24 1.8205
R5474 TG_magic_2.B.n127 TG_magic_2.B.n126 1.8205
R5475 TG_magic_2.B.n18 TG_magic_2.B.t42 1.8205
R5476 TG_magic_2.B.n18 TG_magic_2.B.n17 1.8205
R5477 TG_magic_2.B.n20 TG_magic_2.B.t36 1.8205
R5478 TG_magic_2.B.n20 TG_magic_2.B.n19 1.8205
R5479 TG_magic_2.B.n22 TG_magic_2.B.t49 1.8205
R5480 TG_magic_2.B.n22 TG_magic_2.B.n21 1.8205
R5481 TG_magic_2.B.n24 TG_magic_2.B.t43 1.8205
R5482 TG_magic_2.B.n24 TG_magic_2.B.n23 1.8205
R5483 TG_magic_2.B.n29 TG_magic_2.B.t56 1.8205
R5484 TG_magic_2.B.n29 TG_magic_2.B.n28 1.8205
R5485 TG_magic_2.B.n31 TG_magic_2.B.t53 1.8205
R5486 TG_magic_2.B.n31 TG_magic_2.B.n30 1.8205
R5487 TG_magic_2.B.n33 TG_magic_2.B.t41 1.8205
R5488 TG_magic_2.B.n33 TG_magic_2.B.n32 1.8205
R5489 TG_magic_2.B.n35 TG_magic_2.B.t57 1.8205
R5490 TG_magic_2.B.n35 TG_magic_2.B.n34 1.8205
R5491 TG_magic_2.B.n47 TG_magic_2.B.t58 1.8205
R5492 TG_magic_2.B.n47 TG_magic_2.B.n46 1.8205
R5493 TG_magic_2.B.n78 TG_magic_2.B.t63 1.6385
R5494 TG_magic_2.B.n78 TG_magic_2.B.n77 1.6385
R5495 TG_magic_2.B.n76 TG_magic_2.B.t65 1.6385
R5496 TG_magic_2.B.n76 TG_magic_2.B.n75 1.6385
R5497 TG_magic_2.B.n83 TG_magic_2.B.t64 1.6385
R5498 TG_magic_2.B.n83 TG_magic_2.B.n82 1.6385
R5499 TG_magic_2.B.n81 TG_magic_2.B.t66 1.6385
R5500 TG_magic_2.B.n81 TG_magic_2.B.n80 1.6385
R5501 TG_magic_2.B.n88 TG_magic_2.B.t67 1.6385
R5502 TG_magic_2.B.n88 TG_magic_2.B.n87 1.6385
R5503 TG_magic_2.B.n86 TG_magic_2.B.t68 1.6385
R5504 TG_magic_2.B.n86 TG_magic_2.B.n85 1.6385
R5505 TG_magic_2.B.n116 TG_magic_2.B.t101 1.6385
R5506 TG_magic_2.B.n116 TG_magic_2.B.n115 1.6385
R5507 TG_magic_2.B.n114 TG_magic_2.B.t107 1.6385
R5508 TG_magic_2.B.n114 TG_magic_2.B.n113 1.6385
R5509 TG_magic_2.B.n109 TG_magic_2.B.t103 1.6385
R5510 TG_magic_2.B.n109 TG_magic_2.B.n108 1.6385
R5511 TG_magic_2.B.n107 TG_magic_2.B.t97 1.6385
R5512 TG_magic_2.B.n107 TG_magic_2.B.n106 1.6385
R5513 TG_magic_2.B.n8 TG_magic_2.B.t5 1.6385
R5514 TG_magic_2.B.n8 TG_magic_2.B.n7 1.6385
R5515 TG_magic_2.B.n6 TG_magic_2.B.t11 1.6385
R5516 TG_magic_2.B.n6 TG_magic_2.B.n5 1.6385
R5517 TG_magic_2.B.n3 TG_magic_2.B.t8 1.6385
R5518 TG_magic_2.B.n3 TG_magic_2.B.n2 1.6385
R5519 TG_magic_2.B.n1 TG_magic_2.B.t2 1.6385
R5520 TG_magic_2.B.n1 TG_magic_2.B.n0 1.6385
R5521 TG_magic_2.B.n14 TG_magic_2.B.t9 1.6385
R5522 TG_magic_2.B.n14 TG_magic_2.B.n13 1.6385
R5523 TG_magic_2.B.n12 TG_magic_2.B.t3 1.6385
R5524 TG_magic_2.B.n12 TG_magic_2.B.n11 1.6385
R5525 TG_magic_2.B.n145 TG_magic_2.B.n144 0.882239
R5526 TG_magic_2.B.n148 TG_magic_2.B.n146 0.882239
R5527 TG_magic_2.B.n157 TG_magic_2.B.n155 0.8105
R5528 TG_magic_2.B.n72 TG_magic_2.B.n71 0.657891
R5529 TG_magic_2.B.n62 TG_magic_2.B.n61 0.657891
R5530 TG_magic_2.B.n61 TG_magic_2.B.n60 0.657891
R5531 TG_magic_2.B.n102 TG_magic_2.B.n101 0.657891
R5532 TG_magic_2.B.n101 TG_magic_2.B.n100 0.657891
R5533 TG_magic_2.B.n144 TG_magic_2.B.n143 0.657891
R5534 TG_magic_2.B.n143 TG_magic_2.B.n142 0.657891
R5535 TG_magic_2.B.n141 TG_magic_2.B.n140 0.657891
R5536 TG_magic_2.B.n140 TG_magic_2.B.n139 0.657891
R5537 TG_magic_2.B.n130 TG_magic_2.B.n129 0.657891
R5538 TG_magic_2.B.n129 TG_magic_2.B.n128 0.657891
R5539 TG_magic_2.B.n150 TG_magic_2.B.n148 0.657891
R5540 TG_magic_2.B.n152 TG_magic_2.B.n150 0.657891
R5541 TG_magic_2.B.n154 TG_magic_2.B.n152 0.657891
R5542 TG_magic_2.B.n159 TG_magic_2.B.n157 0.657891
R5543 TG_magic_2.B.n27 TG_magic_2.B.n26 0.657891
R5544 TG_magic_2.B.n26 TG_magic_2.B.n25 0.657891
R5545 TG_magic_2.B.n37 TG_magic_2.B.n36 0.657891
R5546 TG_magic_2.B.n49 TG_magic_2.B.n48 0.657891
R5547 TG_magic_2.B.n48 TG_magic_2.B.n45 0.657891
R5548 TG_magic_2.B.n73 TG_magic_2.B.n72 0.655976
R5549 TG_magic_2.B.n38 TG_magic_2.B.n37 0.655976
R5550 TG_magic_2.B.n50 TG_magic_2.B.n38 0.646796
R5551 TG_magic_2.B.n74 TG_magic_2.B.n73 0.645657
R5552 TG_magic_2.B.n146 TG_magic_2.B.n145 0.6005
R5553 TG_magic_2.B.n90 TG_magic_2.B.n89 0.548416
R5554 TG_magic_2.B.n10 TG_magic_2.B.n9 0.548416
R5555 TG_magic_2.B.n162 TG_magic_2.B.n161 0.516295
R5556 TG_magic_2.B.n119 TG_magic_2.B.n112 0.469375
R5557 TG_magic_2.B.n163 TG_magic_2.B.n119 0.468521
R5558 TG_magic_2.B.n161 TG_magic_2.B.n160 0.448625
R5559 TG_magic_2.B.n103 TG_magic_2.B.n102 0.316429
R5560 TG_magic_2.B.n51 TG_magic_2.B.n27 0.316429
R5561 TG_magic_2.B.n91 TG_magic_2.B.n79 0.304838
R5562 TG_magic_2.B.n16 TG_magic_2.B.n15 0.304838
R5563 TG_magic_2.B TG_magic_2.B.n103 0.2873
R5564 TG_magic_2.B TG_magic_2.B.n51 0.287174
R5565 TG_magic_2.B.n90 TG_magic_2.B.n84 0.284196
R5566 TG_magic_2.B.n10 TG_magic_2.B.n4 0.284196
R5567 TG_magic_2.B.n103 TG_magic_2.B.n74 0.283032
R5568 TG_magic_2.B.n145 TG_magic_2.B.n141 0.282239
R5569 TG_magic_2.B.n146 TG_magic_2.B.n130 0.282239
R5570 TG_magic_2.B.n51 TG_magic_2.B.n50 0.281892
R5571 TG_magic_2.B.n74 TG_magic_2.B.n62 0.279866
R5572 TG_magic_2.B.n50 TG_magic_2.B.n49 0.279866
R5573 TG_magic_2.B.n91 TG_magic_2.B.n90 0.244078
R5574 TG_magic_2.B.n16 TG_magic_2.B.n10 0.244078
R5575 TG_magic_2.B.n155 TG_magic_2.B.n154 0.237239
R5576 TG_magic_2.B.n105 TG_magic_2.B.n104 0.214935
R5577 TG_magic_2.B.n162 TG_magic_2.B.n159 0.206468
R5578 TG_magic_2.B.n111 TG_magic_2.B.n110 0.200307
R5579 TG_magic_2.B.n118 TG_magic_2.B.n117 0.198664
R5580 TG_magic_2.B TG_magic_2.B.n164 0.146158
R5581 TG_magic_2.B.n103 TG_magic_2.B.n91 0.136437
R5582 TG_magic_2.B.n51 TG_magic_2.B.n16 0.136437
R5583 TG_magic_2.B.n164 TG_magic_2.B 0.107932
R5584 a_n1894_n2271.t20 a_n1894_n2271.n19 40.7345
R5585 a_n1894_n2271.n24 a_n1894_n2271.n5 28.094
R5586 a_n1894_n2271.n21 a_n1894_n2271.n20 28.094
R5587 a_n1894_n2271.n33 a_n1894_n2271.n32 28.094
R5588 a_n1894_n2271.n27 a_n1894_n2271.t9 21.9005
R5589 a_n1894_n2271.n27 a_n1894_n2271.t22 21.9005
R5590 a_n1894_n2271.n0 a_n1894_n2271.t14 21.9005
R5591 a_n1894_n2271.n11 a_n1894_n2271.t12 21.9005
R5592 a_n1894_n2271.n12 a_n1894_n2271.t7 21.9005
R5593 a_n1894_n2271.n1 a_n1894_n2271.t10 21.9005
R5594 a_n1894_n2271.n28 a_n1894_n2271.t19 21.9005
R5595 a_n1894_n2271.n28 a_n1894_n2271.t6 21.9005
R5596 a_n1894_n2271.n29 a_n1894_n2271.t15 21.9005
R5597 a_n1894_n2271.n29 a_n1894_n2271.t28 21.9005
R5598 a_n1894_n2271.n2 a_n1894_n2271.t21 21.9005
R5599 a_n1894_n2271.n13 a_n1894_n2271.t17 21.9005
R5600 a_n1894_n2271.n14 a_n1894_n2271.t13 21.9005
R5601 a_n1894_n2271.n3 a_n1894_n2271.t16 21.9005
R5602 a_n1894_n2271.n30 a_n1894_n2271.t25 21.9005
R5603 a_n1894_n2271.n30 a_n1894_n2271.t11 21.9005
R5604 a_n1894_n2271.n31 a_n1894_n2271.t23 21.9005
R5605 a_n1894_n2271.n31 a_n1894_n2271.t8 21.9005
R5606 a_n1894_n2271.n4 a_n1894_n2271.t27 21.9005
R5607 a_n1894_n2271.n15 a_n1894_n2271.t26 21.9005
R5608 a_n1894_n2271.n20 a_n1894_n2271.t20 21.9005
R5609 a_n1894_n2271.n5 a_n1894_n2271.t24 21.9005
R5610 a_n1894_n2271.n32 a_n1894_n2271.t29 21.9005
R5611 a_n1894_n2271.n32 a_n1894_n2271.t18 21.9005
R5612 a_n1894_n2271.n20 a_n1894_n2271.n15 15.8172
R5613 a_n1894_n2271.n5 a_n1894_n2271.n4 15.8172
R5614 a_n1894_n2271.n4 a_n1894_n2271.n3 15.8172
R5615 a_n1894_n2271.n15 a_n1894_n2271.n14 15.8172
R5616 a_n1894_n2271.n14 a_n1894_n2271.n13 15.8172
R5617 a_n1894_n2271.n3 a_n1894_n2271.n2 15.8172
R5618 a_n1894_n2271.n2 a_n1894_n2271.n1 15.8172
R5619 a_n1894_n2271.n13 a_n1894_n2271.n12 15.8172
R5620 a_n1894_n2271.n12 a_n1894_n2271.n11 15.8172
R5621 a_n1894_n2271.n1 a_n1894_n2271.n0 15.8172
R5622 a_n1894_n2271.n28 a_n1894_n2271.n27 15.8172
R5623 a_n1894_n2271.n30 a_n1894_n2271.n29 15.8172
R5624 a_n1894_n2271.n29 a_n1894_n2271.n28 15.8172
R5625 a_n1894_n2271.n32 a_n1894_n2271.n31 15.8172
R5626 a_n1894_n2271.n31 a_n1894_n2271.n30 15.8172
R5627 a_n1894_n2271.n17 a_n1894_n2271.n16 15.1845
R5628 a_n1894_n2271.n19 a_n1894_n2271.n18 15.1845
R5629 a_n1894_n2271.n18 a_n1894_n2271.n17 15.1845
R5630 a_n1894_n2271.n8 a_n1894_n2271.n6 5.44589
R5631 a_n1894_n2271.n8 a_n1894_n2271.n7 4.7885
R5632 a_n1894_n2271.n34 a_n1894_n2271.n33 4.70615
R5633 a_n1894_n2271.n23 a_n1894_n2271.n22 4.4205
R5634 a_n1894_n2271.n26 a_n1894_n2271.n25 4.4205
R5635 a_n1894_n2271.n10 a_n1894_n2271.n9 4.4205
R5636 a_n1894_n2271.n10 a_n1894_n2271.n8 1.1392
R5637 a_n1894_n2271.n26 a_n1894_n2271.n24 0.286152
R5638 a_n1894_n2271.n23 a_n1894_n2271.n21 0.286152
R5639 a_n1894_n2271.n33 a_n1894_n2271.n26 0.282239
R5640 a_n1894_n2271.n21 a_n1894_n2271.n10 0.282239
R5641 a_n1894_n2271.n24 a_n1894_n2271.n23 0.282239
R5642 a_2004_n6151.t18 a_2004_n6151.n25 40.7345
R5643 a_2004_n6151.n15 a_2004_n6151.n6 28.094
R5644 a_2004_n6151.n13 a_2004_n6151.n12 28.094
R5645 a_2004_n6151.n27 a_2004_n6151.n26 28.094
R5646 a_2004_n6151.n26 a_2004_n6151.t18 21.9005
R5647 a_2004_n6151.n17 a_2004_n6151.t10 21.9005
R5648 a_2004_n6151.n17 a_2004_n6151.t15 21.9005
R5649 a_2004_n6151.n1 a_2004_n6151.t29 21.9005
R5650 a_2004_n6151.n7 a_2004_n6151.t27 21.9005
R5651 a_2004_n6151.n8 a_2004_n6151.t12 21.9005
R5652 a_2004_n6151.n2 a_2004_n6151.t14 21.9005
R5653 a_2004_n6151.n18 a_2004_n6151.t25 21.9005
R5654 a_2004_n6151.n18 a_2004_n6151.t22 21.9005
R5655 a_2004_n6151.n19 a_2004_n6151.t17 21.9005
R5656 a_2004_n6151.n19 a_2004_n6151.t21 21.9005
R5657 a_2004_n6151.n3 a_2004_n6151.t9 21.9005
R5658 a_2004_n6151.n9 a_2004_n6151.t7 21.9005
R5659 a_2004_n6151.n10 a_2004_n6151.t19 21.9005
R5660 a_2004_n6151.n4 a_2004_n6151.t20 21.9005
R5661 a_2004_n6151.n20 a_2004_n6151.t6 21.9005
R5662 a_2004_n6151.n20 a_2004_n6151.t28 21.9005
R5663 a_2004_n6151.n21 a_2004_n6151.t24 21.9005
R5664 a_2004_n6151.n21 a_2004_n6151.t26 21.9005
R5665 a_2004_n6151.n5 a_2004_n6151.t16 21.9005
R5666 a_2004_n6151.n11 a_2004_n6151.t13 21.9005
R5667 a_2004_n6151.n12 a_2004_n6151.t8 21.9005
R5668 a_2004_n6151.n6 a_2004_n6151.t11 21.9005
R5669 a_2004_n6151.n26 a_2004_n6151.t23 21.9005
R5670 a_2004_n6151.n6 a_2004_n6151.n5 15.8172
R5671 a_2004_n6151.n26 a_2004_n6151.n21 15.8172
R5672 a_2004_n6151.n21 a_2004_n6151.n20 15.8172
R5673 a_2004_n6151.n5 a_2004_n6151.n4 15.8172
R5674 a_2004_n6151.n4 a_2004_n6151.n3 15.8172
R5675 a_2004_n6151.n20 a_2004_n6151.n19 15.8172
R5676 a_2004_n6151.n19 a_2004_n6151.n18 15.8172
R5677 a_2004_n6151.n3 a_2004_n6151.n2 15.8172
R5678 a_2004_n6151.n2 a_2004_n6151.n1 15.8172
R5679 a_2004_n6151.n18 a_2004_n6151.n17 15.8172
R5680 a_2004_n6151.n8 a_2004_n6151.n7 15.8172
R5681 a_2004_n6151.n9 a_2004_n6151.n8 15.8172
R5682 a_2004_n6151.n10 a_2004_n6151.n9 15.8172
R5683 a_2004_n6151.n11 a_2004_n6151.n10 15.8172
R5684 a_2004_n6151.n12 a_2004_n6151.n11 15.8172
R5685 a_2004_n6151.n23 a_2004_n6151.n22 15.1845
R5686 a_2004_n6151.n24 a_2004_n6151.n23 15.1845
R5687 a_2004_n6151.n25 a_2004_n6151.n24 15.1845
R5688 a_2004_n6151.n0 a_2004_n6151.t5 5.44589
R5689 a_2004_n6151.n0 a_2004_n6151.t4 4.7885
R5690 a_2004_n6151.n13 a_2004_n6151.t1 4.70615
R5691 a_2004_n6151.n14 a_2004_n6151.t0 4.4205
R5692 a_2004_n6151.n16 a_2004_n6151.t2 4.4205
R5693 a_2004_n6151.t3 a_2004_n6151.n28 4.4205
R5694 a_2004_n6151.n28 a_2004_n6151.n0 1.1392
R5695 a_2004_n6151.n27 a_2004_n6151.n16 0.286152
R5696 a_2004_n6151.n15 a_2004_n6151.n14 0.286152
R5697 a_2004_n6151.n16 a_2004_n6151.n15 0.282239
R5698 a_2004_n6151.n14 a_2004_n6151.n13 0.282239
R5699 a_2004_n6151.n28 a_2004_n6151.n27 0.282239
R5700 a_5741_n4853.t19 a_5741_n4853.n22 40.7345
R5701 a_5741_n4853.n24 a_5741_n4853.n23 28.094
R5702 a_5741_n4853.n7 a_5741_n4853.n6 28.094
R5703 a_5741_n4853.n32 a_5741_n4853.n31 28.094
R5704 a_5741_n4853.n4 a_5741_n4853.t11 21.9005
R5705 a_5741_n4853.n2 a_5741_n4853.t18 21.9005
R5706 a_5741_n4853.n1 a_5741_n4853.t26 21.9005
R5707 a_5741_n4853.n1 a_5741_n4853.t17 21.9005
R5708 a_5741_n4853.n26 a_5741_n4853.t21 21.9005
R5709 a_5741_n4853.n14 a_5741_n4853.t25 21.9005
R5710 a_5741_n4853.n15 a_5741_n4853.t16 21.9005
R5711 a_5741_n4853.n27 a_5741_n4853.t8 21.9005
R5712 a_5741_n4853.n2 a_5741_n4853.t29 21.9005
R5713 a_5741_n4853.n3 a_5741_n4853.t23 21.9005
R5714 a_5741_n4853.n3 a_5741_n4853.t10 21.9005
R5715 a_5741_n4853.n28 a_5741_n4853.t13 21.9005
R5716 a_5741_n4853.n16 a_5741_n4853.t22 21.9005
R5717 a_5741_n4853.n17 a_5741_n4853.t9 21.9005
R5718 a_5741_n4853.n29 a_5741_n4853.t27 21.9005
R5719 a_5741_n4853.n4 a_5741_n4853.t24 21.9005
R5720 a_5741_n4853.n6 a_5741_n4853.t20 21.9005
R5721 a_5741_n4853.n6 a_5741_n4853.t7 21.9005
R5722 a_5741_n4853.n5 a_5741_n4853.t15 21.9005
R5723 a_5741_n4853.n5 a_5741_n4853.t28 21.9005
R5724 a_5741_n4853.n30 a_5741_n4853.t6 21.9005
R5725 a_5741_n4853.n18 a_5741_n4853.t14 21.9005
R5726 a_5741_n4853.n23 a_5741_n4853.t19 21.9005
R5727 a_5741_n4853.n31 a_5741_n4853.t12 21.9005
R5728 a_5741_n4853.n23 a_5741_n4853.n18 15.8172
R5729 a_5741_n4853.n31 a_5741_n4853.n30 15.8172
R5730 a_5741_n4853.n30 a_5741_n4853.n29 15.8172
R5731 a_5741_n4853.n18 a_5741_n4853.n17 15.8172
R5732 a_5741_n4853.n17 a_5741_n4853.n16 15.8172
R5733 a_5741_n4853.n29 a_5741_n4853.n28 15.8172
R5734 a_5741_n4853.n28 a_5741_n4853.n27 15.8172
R5735 a_5741_n4853.n16 a_5741_n4853.n15 15.8172
R5736 a_5741_n4853.n15 a_5741_n4853.n14 15.8172
R5737 a_5741_n4853.n27 a_5741_n4853.n26 15.8172
R5738 a_5741_n4853.n2 a_5741_n4853.n1 15.8172
R5739 a_5741_n4853.n4 a_5741_n4853.n3 15.8172
R5740 a_5741_n4853.n3 a_5741_n4853.n2 15.8172
R5741 a_5741_n4853.n6 a_5741_n4853.n5 15.8172
R5742 a_5741_n4853.n5 a_5741_n4853.n4 15.8172
R5743 a_5741_n4853.n20 a_5741_n4853.n19 15.1845
R5744 a_5741_n4853.n22 a_5741_n4853.n21 15.1845
R5745 a_5741_n4853.n21 a_5741_n4853.n20 15.1845
R5746 a_5741_n4853.n12 a_5741_n4853.n11 5.44589
R5747 a_5741_n4853.n12 a_5741_n4853.n10 4.7885
R5748 a_5741_n4853.n7 a_5741_n4853.n0 4.70615
R5749 a_5741_n4853.n13 a_5741_n4853.n9 4.4205
R5750 a_5741_n4853.n25 a_5741_n4853.n8 4.4205
R5751 a_5741_n4853.n34 a_5741_n4853.n33 4.4205
R5752 a_5741_n4853.n13 a_5741_n4853.n12 1.1392
R5753 a_5741_n4853.n25 a_5741_n4853.n24 0.286152
R5754 a_5741_n4853.n33 a_5741_n4853.n32 0.286152
R5755 a_5741_n4853.n32 a_5741_n4853.n25 0.282239
R5756 a_5741_n4853.n24 a_5741_n4853.n13 0.282239
R5757 a_5741_n4853.n33 a_5741_n4853.n7 0.282239
R5758 TG_GATE_SWITCH_magic_5.B.n99 TG_GATE_SWITCH_magic_5.B.n98 5.44589
R5759 TG_GATE_SWITCH_magic_5.B.n76 TG_GATE_SWITCH_magic_5.B.n74 5.07789
R5760 TG_GATE_SWITCH_magic_5.B.n102 TG_GATE_SWITCH_magic_5.B.t7 4.7885
R5761 TG_GATE_SWITCH_magic_5.B.n99 TG_GATE_SWITCH_magic_5.B.n97 4.7885
R5762 TG_GATE_SWITCH_magic_5.B.n103 TG_GATE_SWITCH_magic_5.B.t16 4.7885
R5763 TG_GATE_SWITCH_magic_5.B.n86 TG_GATE_SWITCH_magic_5.B.t63 4.4205
R5764 TG_GATE_SWITCH_magic_5.B.n85 TG_GATE_SWITCH_magic_5.B.t71 4.4205
R5765 TG_GATE_SWITCH_magic_5.B.n84 TG_GATE_SWITCH_magic_5.B.t25 4.4205
R5766 TG_GATE_SWITCH_magic_5.B.n83 TG_GATE_SWITCH_magic_5.B.t24 4.4205
R5767 TG_GATE_SWITCH_magic_5.B.n80 TG_GATE_SWITCH_magic_5.B.n79 4.4205
R5768 TG_GATE_SWITCH_magic_5.B.n78 TG_GATE_SWITCH_magic_5.B.n77 4.4205
R5769 TG_GATE_SWITCH_magic_5.B.n76 TG_GATE_SWITCH_magic_5.B.n75 4.4205
R5770 TG_GATE_SWITCH_magic_5.B.n106 TG_GATE_SWITCH_magic_5.B.n105 4.26515
R5771 TG_GATE_SWITCH_magic_5.B.n91 TG_GATE_SWITCH_magic_5.B.n90 3.80789
R5772 TG_GATE_SWITCH_magic_5.B.n96 TG_GATE_SWITCH_magic_5.B.n95 3.80789
R5773 TG_GATE_SWITCH_magic_5.B.n48 TG_GATE_SWITCH_magic_5.B.n47 3.80789
R5774 TG_GATE_SWITCH_magic_5.B.n43 TG_GATE_SWITCH_magic_5.B.n42 3.80789
R5775 TG_GATE_SWITCH_magic_5.B.n38 TG_GATE_SWITCH_magic_5.B.n37 3.80789
R5776 TG_GATE_SWITCH_magic_5.B.n67 TG_GATE_SWITCH_magic_5.B.n64 3.25789
R5777 TG_GATE_SWITCH_magic_5.B.n56 TG_GATE_SWITCH_magic_5.B.n53 3.25789
R5778 TG_GATE_SWITCH_magic_5.B.n4 TG_GATE_SWITCH_magic_5.B.n1 3.25789
R5779 TG_GATE_SWITCH_magic_5.B.n15 TG_GATE_SWITCH_magic_5.B.n12 3.25789
R5780 TG_GATE_SWITCH_magic_5.B.n27 TG_GATE_SWITCH_magic_5.B.n24 3.25789
R5781 TG_GATE_SWITCH_magic_5.B.n91 TG_GATE_SWITCH_magic_5.B.n88 3.1505
R5782 TG_GATE_SWITCH_magic_5.B.n96 TG_GATE_SWITCH_magic_5.B.n93 3.1505
R5783 TG_GATE_SWITCH_magic_5.B.n48 TG_GATE_SWITCH_magic_5.B.n45 3.1505
R5784 TG_GATE_SWITCH_magic_5.B.n43 TG_GATE_SWITCH_magic_5.B.n40 3.1505
R5785 TG_GATE_SWITCH_magic_5.B.n38 TG_GATE_SWITCH_magic_5.B.n35 3.1505
R5786 TG_GATE_SWITCH_magic_5.B.n67 TG_GATE_SWITCH_magic_5.B.n66 2.6005
R5787 TG_GATE_SWITCH_magic_5.B.n70 TG_GATE_SWITCH_magic_5.B.n69 2.6005
R5788 TG_GATE_SWITCH_magic_5.B.n73 TG_GATE_SWITCH_magic_5.B.n72 2.6005
R5789 TG_GATE_SWITCH_magic_5.B.n56 TG_GATE_SWITCH_magic_5.B.n55 2.6005
R5790 TG_GATE_SWITCH_magic_5.B.n59 TG_GATE_SWITCH_magic_5.B.n58 2.6005
R5791 TG_GATE_SWITCH_magic_5.B.n62 TG_GATE_SWITCH_magic_5.B.n61 2.6005
R5792 TG_GATE_SWITCH_magic_5.B.n4 TG_GATE_SWITCH_magic_5.B.n3 2.6005
R5793 TG_GATE_SWITCH_magic_5.B.n7 TG_GATE_SWITCH_magic_5.B.n6 2.6005
R5794 TG_GATE_SWITCH_magic_5.B.n10 TG_GATE_SWITCH_magic_5.B.n9 2.6005
R5795 TG_GATE_SWITCH_magic_5.B.n18 TG_GATE_SWITCH_magic_5.B.n17 2.6005
R5796 TG_GATE_SWITCH_magic_5.B.n15 TG_GATE_SWITCH_magic_5.B.n14 2.6005
R5797 TG_GATE_SWITCH_magic_5.B.n21 TG_GATE_SWITCH_magic_5.B.n20 2.6005
R5798 TG_GATE_SWITCH_magic_5.B.n27 TG_GATE_SWITCH_magic_5.B.n26 2.6005
R5799 TG_GATE_SWITCH_magic_5.B.n30 TG_GATE_SWITCH_magic_5.B.n29 2.6005
R5800 TG_GATE_SWITCH_magic_5.B.n33 TG_GATE_SWITCH_magic_5.B.n32 2.6005
R5801 TG_GATE_SWITCH_magic_5.B.n72 TG_GATE_SWITCH_magic_5.B.t61 1.8205
R5802 TG_GATE_SWITCH_magic_5.B.n72 TG_GATE_SWITCH_magic_5.B.n71 1.8205
R5803 TG_GATE_SWITCH_magic_5.B.n69 TG_GATE_SWITCH_magic_5.B.t64 1.8205
R5804 TG_GATE_SWITCH_magic_5.B.n69 TG_GATE_SWITCH_magic_5.B.n68 1.8205
R5805 TG_GATE_SWITCH_magic_5.B.n66 TG_GATE_SWITCH_magic_5.B.t20 1.8205
R5806 TG_GATE_SWITCH_magic_5.B.n66 TG_GATE_SWITCH_magic_5.B.n65 1.8205
R5807 TG_GATE_SWITCH_magic_5.B.n64 TG_GATE_SWITCH_magic_5.B.t33 1.8205
R5808 TG_GATE_SWITCH_magic_5.B.n64 TG_GATE_SWITCH_magic_5.B.n63 1.8205
R5809 TG_GATE_SWITCH_magic_5.B.n61 TG_GATE_SWITCH_magic_5.B.t59 1.8205
R5810 TG_GATE_SWITCH_magic_5.B.n61 TG_GATE_SWITCH_magic_5.B.n60 1.8205
R5811 TG_GATE_SWITCH_magic_5.B.n58 TG_GATE_SWITCH_magic_5.B.t60 1.8205
R5812 TG_GATE_SWITCH_magic_5.B.n58 TG_GATE_SWITCH_magic_5.B.n57 1.8205
R5813 TG_GATE_SWITCH_magic_5.B.n55 TG_GATE_SWITCH_magic_5.B.t18 1.8205
R5814 TG_GATE_SWITCH_magic_5.B.n55 TG_GATE_SWITCH_magic_5.B.n54 1.8205
R5815 TG_GATE_SWITCH_magic_5.B.n53 TG_GATE_SWITCH_magic_5.B.t31 1.8205
R5816 TG_GATE_SWITCH_magic_5.B.n53 TG_GATE_SWITCH_magic_5.B.n52 1.8205
R5817 TG_GATE_SWITCH_magic_5.B.n9 TG_GATE_SWITCH_magic_5.B.t56 1.8205
R5818 TG_GATE_SWITCH_magic_5.B.n9 TG_GATE_SWITCH_magic_5.B.n8 1.8205
R5819 TG_GATE_SWITCH_magic_5.B.n6 TG_GATE_SWITCH_magic_5.B.t48 1.8205
R5820 TG_GATE_SWITCH_magic_5.B.n6 TG_GATE_SWITCH_magic_5.B.n5 1.8205
R5821 TG_GATE_SWITCH_magic_5.B.n3 TG_GATE_SWITCH_magic_5.B.t3 1.8205
R5822 TG_GATE_SWITCH_magic_5.B.n3 TG_GATE_SWITCH_magic_5.B.n2 1.8205
R5823 TG_GATE_SWITCH_magic_5.B.n1 TG_GATE_SWITCH_magic_5.B.t67 1.8205
R5824 TG_GATE_SWITCH_magic_5.B.n1 TG_GATE_SWITCH_magic_5.B.n0 1.8205
R5825 TG_GATE_SWITCH_magic_5.B.n20 TG_GATE_SWITCH_magic_5.B.t17 1.8205
R5826 TG_GATE_SWITCH_magic_5.B.n20 TG_GATE_SWITCH_magic_5.B.n19 1.8205
R5827 TG_GATE_SWITCH_magic_5.B.n12 TG_GATE_SWITCH_magic_5.B.t29 1.8205
R5828 TG_GATE_SWITCH_magic_5.B.n12 TG_GATE_SWITCH_magic_5.B.n11 1.8205
R5829 TG_GATE_SWITCH_magic_5.B.n14 TG_GATE_SWITCH_magic_5.B.t52 1.8205
R5830 TG_GATE_SWITCH_magic_5.B.n14 TG_GATE_SWITCH_magic_5.B.n13 1.8205
R5831 TG_GATE_SWITCH_magic_5.B.n17 TG_GATE_SWITCH_magic_5.B.t55 1.8205
R5832 TG_GATE_SWITCH_magic_5.B.n17 TG_GATE_SWITCH_magic_5.B.n16 1.8205
R5833 TG_GATE_SWITCH_magic_5.B.n32 TG_GATE_SWITCH_magic_5.B.t49 1.8205
R5834 TG_GATE_SWITCH_magic_5.B.n32 TG_GATE_SWITCH_magic_5.B.n31 1.8205
R5835 TG_GATE_SWITCH_magic_5.B.n29 TG_GATE_SWITCH_magic_5.B.t1 1.8205
R5836 TG_GATE_SWITCH_magic_5.B.n29 TG_GATE_SWITCH_magic_5.B.n28 1.8205
R5837 TG_GATE_SWITCH_magic_5.B.n26 TG_GATE_SWITCH_magic_5.B.t28 1.8205
R5838 TG_GATE_SWITCH_magic_5.B.n26 TG_GATE_SWITCH_magic_5.B.n25 1.8205
R5839 TG_GATE_SWITCH_magic_5.B.n24 TG_GATE_SWITCH_magic_5.B.t53 1.8205
R5840 TG_GATE_SWITCH_magic_5.B.n24 TG_GATE_SWITCH_magic_5.B.n23 1.8205
R5841 TG_GATE_SWITCH_magic_5.B.n88 TG_GATE_SWITCH_magic_5.B.t15 1.6385
R5842 TG_GATE_SWITCH_magic_5.B.n88 TG_GATE_SWITCH_magic_5.B.n87 1.6385
R5843 TG_GATE_SWITCH_magic_5.B.n90 TG_GATE_SWITCH_magic_5.B.t12 1.6385
R5844 TG_GATE_SWITCH_magic_5.B.n90 TG_GATE_SWITCH_magic_5.B.n89 1.6385
R5845 TG_GATE_SWITCH_magic_5.B.n93 TG_GATE_SWITCH_magic_5.B.t13 1.6385
R5846 TG_GATE_SWITCH_magic_5.B.n93 TG_GATE_SWITCH_magic_5.B.n92 1.6385
R5847 TG_GATE_SWITCH_magic_5.B.n95 TG_GATE_SWITCH_magic_5.B.t11 1.6385
R5848 TG_GATE_SWITCH_magic_5.B.n95 TG_GATE_SWITCH_magic_5.B.n94 1.6385
R5849 TG_GATE_SWITCH_magic_5.B.n45 TG_GATE_SWITCH_magic_5.B.t42 1.6385
R5850 TG_GATE_SWITCH_magic_5.B.n45 TG_GATE_SWITCH_magic_5.B.n44 1.6385
R5851 TG_GATE_SWITCH_magic_5.B.n47 TG_GATE_SWITCH_magic_5.B.t45 1.6385
R5852 TG_GATE_SWITCH_magic_5.B.n47 TG_GATE_SWITCH_magic_5.B.n46 1.6385
R5853 TG_GATE_SWITCH_magic_5.B.n40 TG_GATE_SWITCH_magic_5.B.t43 1.6385
R5854 TG_GATE_SWITCH_magic_5.B.n40 TG_GATE_SWITCH_magic_5.B.n39 1.6385
R5855 TG_GATE_SWITCH_magic_5.B.n42 TG_GATE_SWITCH_magic_5.B.t40 1.6385
R5856 TG_GATE_SWITCH_magic_5.B.n42 TG_GATE_SWITCH_magic_5.B.n41 1.6385
R5857 TG_GATE_SWITCH_magic_5.B.n35 TG_GATE_SWITCH_magic_5.B.t44 1.6385
R5858 TG_GATE_SWITCH_magic_5.B.n35 TG_GATE_SWITCH_magic_5.B.n34 1.6385
R5859 TG_GATE_SWITCH_magic_5.B.n37 TG_GATE_SWITCH_magic_5.B.t41 1.6385
R5860 TG_GATE_SWITCH_magic_5.B.n37 TG_GATE_SWITCH_magic_5.B.n36 1.6385
R5861 TG_GATE_SWITCH_magic_5.B.n105 TG_GATE_SWITCH_magic_5.B.n104 1.56655
R5862 TG_GATE_SWITCH_magic_5.B.n105 TG_GATE_SWITCH_magic_5.B 1.16233
R5863 TG_GATE_SWITCH_magic_5.B.n100 TG_GATE_SWITCH_magic_5.B.n99 0.884196
R5864 TG_GATE_SWITCH_magic_5.B.n102 TG_GATE_SWITCH_magic_5.B.n101 0.884196
R5865 TG_GATE_SWITCH_magic_5.B.n81 TG_GATE_SWITCH_magic_5.B.n80 0.882239
R5866 TG_GATE_SWITCH_magic_5.B.n83 TG_GATE_SWITCH_magic_5.B.n82 0.882239
R5867 TG_GATE_SWITCH_magic_5.B.n104 TG_GATE_SWITCH_magic_5.B.n103 0.8105
R5868 TG_GATE_SWITCH_magic_5.B.n78 TG_GATE_SWITCH_magic_5.B.n76 0.657891
R5869 TG_GATE_SWITCH_magic_5.B.n80 TG_GATE_SWITCH_magic_5.B.n78 0.657891
R5870 TG_GATE_SWITCH_magic_5.B.n70 TG_GATE_SWITCH_magic_5.B.n67 0.657891
R5871 TG_GATE_SWITCH_magic_5.B.n73 TG_GATE_SWITCH_magic_5.B.n70 0.657891
R5872 TG_GATE_SWITCH_magic_5.B.n59 TG_GATE_SWITCH_magic_5.B.n56 0.657891
R5873 TG_GATE_SWITCH_magic_5.B.n62 TG_GATE_SWITCH_magic_5.B.n59 0.657891
R5874 TG_GATE_SWITCH_magic_5.B.n86 TG_GATE_SWITCH_magic_5.B.n85 0.657891
R5875 TG_GATE_SWITCH_magic_5.B.n85 TG_GATE_SWITCH_magic_5.B.n84 0.657891
R5876 TG_GATE_SWITCH_magic_5.B.n84 TG_GATE_SWITCH_magic_5.B.n83 0.657891
R5877 TG_GATE_SWITCH_magic_5.B.n7 TG_GATE_SWITCH_magic_5.B.n4 0.657891
R5878 TG_GATE_SWITCH_magic_5.B.n10 TG_GATE_SWITCH_magic_5.B.n7 0.657891
R5879 TG_GATE_SWITCH_magic_5.B.n18 TG_GATE_SWITCH_magic_5.B.n15 0.657891
R5880 TG_GATE_SWITCH_magic_5.B.n30 TG_GATE_SWITCH_magic_5.B.n27 0.657891
R5881 TG_GATE_SWITCH_magic_5.B.n33 TG_GATE_SWITCH_magic_5.B.n30 0.657891
R5882 TG_GATE_SWITCH_magic_5.B.n103 TG_GATE_SWITCH_magic_5.B.n102 0.657891
R5883 TG_GATE_SWITCH_magic_5.B.n21 TG_GATE_SWITCH_magic_5.B.n18 0.655976
R5884 TG_GATE_SWITCH_magic_5.B.n22 TG_GATE_SWITCH_magic_5.B.n21 0.645657
R5885 TG_GATE_SWITCH_magic_5.B.n101 TG_GATE_SWITCH_magic_5.B.n100 0.6005
R5886 TG_GATE_SWITCH_magic_5.B.n82 TG_GATE_SWITCH_magic_5.B.n81 0.6005
R5887 TG_GATE_SWITCH_magic_5.B.n49 TG_GATE_SWITCH_magic_5.B.n48 0.548416
R5888 TG_GATE_SWITCH_magic_5.B.n51 TG_GATE_SWITCH_magic_5.B.n33 0.317366
R5889 TG_GATE_SWITCH_magic_5.B.n50 TG_GATE_SWITCH_magic_5.B.n38 0.304838
R5890 TG_GATE_SWITCH_magic_5.B.n101 TG_GATE_SWITCH_magic_5.B.n91 0.284196
R5891 TG_GATE_SWITCH_magic_5.B.n100 TG_GATE_SWITCH_magic_5.B.n96 0.284196
R5892 TG_GATE_SWITCH_magic_5.B.n49 TG_GATE_SWITCH_magic_5.B.n43 0.284196
R5893 TG_GATE_SWITCH_magic_5.B.n51 TG_GATE_SWITCH_magic_5.B.n22 0.283032
R5894 TG_GATE_SWITCH_magic_5.B.n81 TG_GATE_SWITCH_magic_5.B.n73 0.282239
R5895 TG_GATE_SWITCH_magic_5.B.n82 TG_GATE_SWITCH_magic_5.B.n62 0.282239
R5896 TG_GATE_SWITCH_magic_5.B.n22 TG_GATE_SWITCH_magic_5.B.n10 0.279866
R5897 TG_GATE_SWITCH_magic_5.B.n50 TG_GATE_SWITCH_magic_5.B.n49 0.244078
R5898 TG_GATE_SWITCH_magic_5.B.n104 TG_GATE_SWITCH_magic_5.B.n86 0.237239
R5899 TG_GATE_SWITCH_magic_5.B.n106 TG_GATE_SWITCH_magic_5.B.n51 0.228729
R5900 TG_GATE_SWITCH_magic_5.B.n51 TG_GATE_SWITCH_magic_5.B.n50 0.1355
R5901 TG_GATE_SWITCH_magic_5.B TG_GATE_SWITCH_magic_5.B.n106 0.0554087
R5902 a_n4297_n2278.t23 a_n4297_n2278.n13 40.7345
R5903 a_n4297_n2278.n15 a_n4297_n2278.n14 28.094
R5904 a_n4297_n2278.n24 a_n4297_n2278.n23 28.094
R5905 a_n4297_n2278.n32 a_n4297_n2278.n31 28.094
R5906 a_n4297_n2278.n5 a_n4297_n2278.t13 21.9005
R5907 a_n4297_n2278.n26 a_n4297_n2278.t21 21.9005
R5908 a_n4297_n2278.n26 a_n4297_n2278.t7 21.9005
R5909 a_n4297_n2278.n18 a_n4297_n2278.t12 21.9005
R5910 a_n4297_n2278.n19 a_n4297_n2278.t9 21.9005
R5911 a_n4297_n2278.n27 a_n4297_n2278.t29 21.9005
R5912 a_n4297_n2278.n27 a_n4297_n2278.t17 21.9005
R5913 a_n4297_n2278.n6 a_n4297_n2278.t10 21.9005
R5914 a_n4297_n2278.n7 a_n4297_n2278.t20 21.9005
R5915 a_n4297_n2278.n28 a_n4297_n2278.t27 21.9005
R5916 a_n4297_n2278.n28 a_n4297_n2278.t11 21.9005
R5917 a_n4297_n2278.n20 a_n4297_n2278.t19 21.9005
R5918 a_n4297_n2278.n21 a_n4297_n2278.t15 21.9005
R5919 a_n4297_n2278.n29 a_n4297_n2278.t8 21.9005
R5920 a_n4297_n2278.n29 a_n4297_n2278.t24 21.9005
R5921 a_n4297_n2278.n8 a_n4297_n2278.t16 21.9005
R5922 a_n4297_n2278.n31 a_n4297_n2278.t28 21.9005
R5923 a_n4297_n2278.n14 a_n4297_n2278.t23 21.9005
R5924 a_n4297_n2278.n9 a_n4297_n2278.t26 21.9005
R5925 a_n4297_n2278.n30 a_n4297_n2278.t6 21.9005
R5926 a_n4297_n2278.n30 a_n4297_n2278.t18 21.9005
R5927 a_n4297_n2278.n22 a_n4297_n2278.t25 21.9005
R5928 a_n4297_n2278.n23 a_n4297_n2278.t22 21.9005
R5929 a_n4297_n2278.n31 a_n4297_n2278.t14 21.9005
R5930 a_n4297_n2278.n31 a_n4297_n2278.n30 15.8172
R5931 a_n4297_n2278.n9 a_n4297_n2278.n8 15.8172
R5932 a_n4297_n2278.n30 a_n4297_n2278.n29 15.8172
R5933 a_n4297_n2278.n29 a_n4297_n2278.n28 15.8172
R5934 a_n4297_n2278.n8 a_n4297_n2278.n7 15.8172
R5935 a_n4297_n2278.n7 a_n4297_n2278.n6 15.8172
R5936 a_n4297_n2278.n28 a_n4297_n2278.n27 15.8172
R5937 a_n4297_n2278.n27 a_n4297_n2278.n26 15.8172
R5938 a_n4297_n2278.n6 a_n4297_n2278.n5 15.8172
R5939 a_n4297_n2278.n20 a_n4297_n2278.n19 15.8172
R5940 a_n4297_n2278.n19 a_n4297_n2278.n18 15.8172
R5941 a_n4297_n2278.n22 a_n4297_n2278.n21 15.8172
R5942 a_n4297_n2278.n21 a_n4297_n2278.n20 15.8172
R5943 a_n4297_n2278.n14 a_n4297_n2278.n9 15.8172
R5944 a_n4297_n2278.n23 a_n4297_n2278.n22 15.8172
R5945 a_n4297_n2278.n12 a_n4297_n2278.n11 15.1845
R5946 a_n4297_n2278.n11 a_n4297_n2278.n10 15.1845
R5947 a_n4297_n2278.n13 a_n4297_n2278.n12 15.1845
R5948 a_n4297_n2278.n2 a_n4297_n2278.n0 5.44589
R5949 a_n4297_n2278.n2 a_n4297_n2278.n1 4.7885
R5950 a_n4297_n2278.n24 a_n4297_n2278.n17 4.70615
R5951 a_n4297_n2278.n4 a_n4297_n2278.n3 4.4205
R5952 a_n4297_n2278.n25 a_n4297_n2278.n16 4.4205
R5953 a_n4297_n2278.n34 a_n4297_n2278.n33 4.4205
R5954 a_n4297_n2278.n4 a_n4297_n2278.n2 1.1392
R5955 a_n4297_n2278.n32 a_n4297_n2278.n25 0.286152
R5956 a_n4297_n2278.n33 a_n4297_n2278.n15 0.286152
R5957 a_n4297_n2278.n15 a_n4297_n2278.n4 0.282239
R5958 a_n4297_n2278.n25 a_n4297_n2278.n24 0.282239
R5959 a_n4297_n2278.n33 a_n4297_n2278.n32 0.282239
R5960 A0.n47 A0.n46 5.44589
R5961 A0.n24 A0.n22 5.07789
R5962 A0.n50 A0.t32 4.7885
R5963 A0.n51 A0.t30 4.7885
R5964 A0.n47 A0.n45 4.7885
R5965 A0.n34 A0.t6 4.4205
R5966 A0.n33 A0.t1 4.4205
R5967 A0.n32 A0.t15 4.4205
R5968 A0.n31 A0.t7 4.4205
R5969 A0.n28 A0.n27 4.4205
R5970 A0.n26 A0.n25 4.4205
R5971 A0.n24 A0.n23 4.4205
R5972 A0.n39 A0.n38 3.80789
R5973 A0.n44 A0.n43 3.80789
R5974 A0.n15 A0.n12 3.25789
R5975 A0.n4 A0.n1 3.25789
R5976 A0.n39 A0.n36 3.1505
R5977 A0.n44 A0.n41 3.1505
R5978 A0.n15 A0.n14 2.6005
R5979 A0.n18 A0.n17 2.6005
R5980 A0.n21 A0.n20 2.6005
R5981 A0.n4 A0.n3 2.6005
R5982 A0.n7 A0.n6 2.6005
R5983 A0.n10 A0.n9 2.6005
R5984 A0.n20 A0.t20 1.8205
R5985 A0.n20 A0.n19 1.8205
R5986 A0.n17 A0.t0 1.8205
R5987 A0.n17 A0.n16 1.8205
R5988 A0.n14 A0.t12 1.8205
R5989 A0.n14 A0.n13 1.8205
R5990 A0.n12 A0.t19 1.8205
R5991 A0.n12 A0.n11 1.8205
R5992 A0.n9 A0.t14 1.8205
R5993 A0.n9 A0.n8 1.8205
R5994 A0.n6 A0.t21 1.8205
R5995 A0.n6 A0.n5 1.8205
R5996 A0.n3 A0.t5 1.8205
R5997 A0.n3 A0.n2 1.8205
R5998 A0.n1 A0.t13 1.8205
R5999 A0.n1 A0.n0 1.8205
R6000 A0.n36 A0.t28 1.6385
R6001 A0.n36 A0.n35 1.6385
R6002 A0.n38 A0.t26 1.6385
R6003 A0.n38 A0.n37 1.6385
R6004 A0.n41 A0.t24 1.6385
R6005 A0.n41 A0.n40 1.6385
R6006 A0.n43 A0.t34 1.6385
R6007 A0.n43 A0.n42 1.6385
R6008 A0 A0.n52 1.54838
R6009 A0.n48 A0.n47 0.884196
R6010 A0.n50 A0.n49 0.884196
R6011 A0.n29 A0.n28 0.882239
R6012 A0.n31 A0.n30 0.882239
R6013 A0.n51 A0.n50 0.657891
R6014 A0.n26 A0.n24 0.657891
R6015 A0.n28 A0.n26 0.657891
R6016 A0.n18 A0.n15 0.657891
R6017 A0.n21 A0.n18 0.657891
R6018 A0.n7 A0.n4 0.657891
R6019 A0.n10 A0.n7 0.657891
R6020 A0.n34 A0.n33 0.657891
R6021 A0.n33 A0.n32 0.657891
R6022 A0.n32 A0.n31 0.657891
R6023 A0.n49 A0.n48 0.6005
R6024 A0.n30 A0.n29 0.6005
R6025 A0.n52 A0.n51 0.60042
R6026 A0.n49 A0.n39 0.284196
R6027 A0.n48 A0.n44 0.284196
R6028 A0.n29 A0.n21 0.282239
R6029 A0.n30 A0.n10 0.282239
R6030 A0.n52 A0.n34 0.277389
R6031 A7.n47 A7.n45 5.44589
R6032 A7.n26 A7.n25 5.07789
R6033 A7.n51 A7.t16 4.7885
R6034 A7.n50 A7.t10 4.7885
R6035 A7.n47 A7.n46 4.7885
R6036 A7.n31 A7.t34 4.4205
R6037 A7.n32 A7.t22 4.4205
R6038 A7.n33 A7.t25 4.4205
R6039 A7.n34 A7.t33 4.4205
R6040 A7.n28 A7.n22 4.4205
R6041 A7.n27 A7.n23 4.4205
R6042 A7.n26 A7.n24 4.4205
R6043 A7.n53 A7 3.97587
R6044 A7.n44 A7.n41 3.80789
R6045 A7.n39 A7.n36 3.80789
R6046 A7.n8 A7.n7 3.25789
R6047 A7.n19 A7.n18 3.25789
R6048 A7.n44 A7.n43 3.1505
R6049 A7.n39 A7.n38 3.1505
R6050 A7.n8 A7.n5 2.6005
R6051 A7.n9 A7.n3 2.6005
R6052 A7.n10 A7.n1 2.6005
R6053 A7.n19 A7.n16 2.6005
R6054 A7.n20 A7.n14 2.6005
R6055 A7.n21 A7.n12 2.6005
R6056 A7.n1 A7.t29 1.8205
R6057 A7.n1 A7.n0 1.8205
R6058 A7.n3 A7.t0 1.8205
R6059 A7.n3 A7.n2 1.8205
R6060 A7.n5 A7.t2 1.8205
R6061 A7.n5 A7.n4 1.8205
R6062 A7.n7 A7.t26 1.8205
R6063 A7.n7 A7.n6 1.8205
R6064 A7.n12 A7.t21 1.8205
R6065 A7.n12 A7.n11 1.8205
R6066 A7.n14 A7.t35 1.8205
R6067 A7.n14 A7.n13 1.8205
R6068 A7.n16 A7.t8 1.8205
R6069 A7.n16 A7.n15 1.8205
R6070 A7.n18 A7.t4 1.8205
R6071 A7.n18 A7.n17 1.8205
R6072 A7.n43 A7.t15 1.6385
R6073 A7.n43 A7.n42 1.6385
R6074 A7.n41 A7.t9 1.6385
R6075 A7.n41 A7.n40 1.6385
R6076 A7.n38 A7.t12 1.6385
R6077 A7.n38 A7.n37 1.6385
R6078 A7.n36 A7.t18 1.6385
R6079 A7.n36 A7.n35 1.6385
R6080 A7.n53 A7.n52 1.36282
R6081 A7.n48 A7.n47 0.884196
R6082 A7.n50 A7.n49 0.884196
R6083 A7.n29 A7.n28 0.882239
R6084 A7.n31 A7.n30 0.882239
R6085 A7.n10 A7.n9 0.657891
R6086 A7.n9 A7.n8 0.657891
R6087 A7.n21 A7.n20 0.657891
R6088 A7.n20 A7.n19 0.657891
R6089 A7.n28 A7.n27 0.657891
R6090 A7.n27 A7.n26 0.657891
R6091 A7.n32 A7.n31 0.657891
R6092 A7.n33 A7.n32 0.657891
R6093 A7.n34 A7.n33 0.657891
R6094 A7.n51 A7.n50 0.657891
R6095 A7.n52 A7.n51 0.600532
R6096 A7.n30 A7.n29 0.6005
R6097 A7.n49 A7.n48 0.6005
R6098 A7.n48 A7.n44 0.284196
R6099 A7.n49 A7.n39 0.284196
R6100 A7.n30 A7.n10 0.282239
R6101 A7.n29 A7.n21 0.282239
R6102 A7.n52 A7.n34 0.278258
R6103 A7 A7.n53 0.186125
R6104 a_301_n7430.t26 a_301_n7430.n30 40.7345
R6105 a_301_n7430.n20 a_301_n7430.n9 28.094
R6106 a_301_n7430.n18 a_301_n7430.n17 28.094
R6107 a_301_n7430.n32 a_301_n7430.n31 28.094
R6108 a_301_n7430.n22 a_301_n7430.t29 21.9005
R6109 a_301_n7430.n22 a_301_n7430.t8 21.9005
R6110 a_301_n7430.n4 a_301_n7430.t20 21.9005
R6111 a_301_n7430.n12 a_301_n7430.t18 21.9005
R6112 a_301_n7430.n13 a_301_n7430.t24 21.9005
R6113 a_301_n7430.n5 a_301_n7430.t27 21.9005
R6114 a_301_n7430.n23 a_301_n7430.t12 21.9005
R6115 a_301_n7430.n23 a_301_n7430.t9 21.9005
R6116 a_301_n7430.n24 a_301_n7430.t21 21.9005
R6117 a_301_n7430.n24 a_301_n7430.t28 21.9005
R6118 a_301_n7430.n6 a_301_n7430.t15 21.9005
R6119 a_301_n7430.n14 a_301_n7430.t14 21.9005
R6120 a_301_n7430.n15 a_301_n7430.t22 21.9005
R6121 a_301_n7430.n7 a_301_n7430.t23 21.9005
R6122 a_301_n7430.n25 a_301_n7430.t10 21.9005
R6123 a_301_n7430.n25 a_301_n7430.t7 21.9005
R6124 a_301_n7430.n31 a_301_n7430.t26 21.9005
R6125 a_301_n7430.n26 a_301_n7430.t19 21.9005
R6126 a_301_n7430.n26 a_301_n7430.t25 21.9005
R6127 a_301_n7430.n8 a_301_n7430.t13 21.9005
R6128 a_301_n7430.n16 a_301_n7430.t11 21.9005
R6129 a_301_n7430.n17 a_301_n7430.t16 21.9005
R6130 a_301_n7430.n9 a_301_n7430.t17 21.9005
R6131 a_301_n7430.n31 a_301_n7430.t6 21.9005
R6132 a_301_n7430.n9 a_301_n7430.n8 15.8172
R6133 a_301_n7430.n31 a_301_n7430.n26 15.8172
R6134 a_301_n7430.n26 a_301_n7430.n25 15.8172
R6135 a_301_n7430.n8 a_301_n7430.n7 15.8172
R6136 a_301_n7430.n7 a_301_n7430.n6 15.8172
R6137 a_301_n7430.n25 a_301_n7430.n24 15.8172
R6138 a_301_n7430.n24 a_301_n7430.n23 15.8172
R6139 a_301_n7430.n6 a_301_n7430.n5 15.8172
R6140 a_301_n7430.n5 a_301_n7430.n4 15.8172
R6141 a_301_n7430.n23 a_301_n7430.n22 15.8172
R6142 a_301_n7430.n14 a_301_n7430.n13 15.8172
R6143 a_301_n7430.n13 a_301_n7430.n12 15.8172
R6144 a_301_n7430.n16 a_301_n7430.n15 15.8172
R6145 a_301_n7430.n15 a_301_n7430.n14 15.8172
R6146 a_301_n7430.n17 a_301_n7430.n16 15.8172
R6147 a_301_n7430.n29 a_301_n7430.n28 15.1845
R6148 a_301_n7430.n28 a_301_n7430.n27 15.1845
R6149 a_301_n7430.n30 a_301_n7430.n29 15.1845
R6150 a_301_n7430.n2 a_301_n7430.n0 5.44589
R6151 a_301_n7430.n2 a_301_n7430.n1 4.7885
R6152 a_301_n7430.n18 a_301_n7430.n11 4.70615
R6153 a_301_n7430.n19 a_301_n7430.n10 4.4205
R6154 a_301_n7430.n21 a_301_n7430.n3 4.4205
R6155 a_301_n7430.n34 a_301_n7430.n33 4.4205
R6156 a_301_n7430.n33 a_301_n7430.n2 1.1392
R6157 a_301_n7430.n32 a_301_n7430.n21 0.286152
R6158 a_301_n7430.n20 a_301_n7430.n19 0.286152
R6159 a_301_n7430.n21 a_301_n7430.n20 0.282239
R6160 a_301_n7430.n19 a_301_n7430.n18 0.282239
R6161 a_301_n7430.n33 a_301_n7430.n32 0.282239
R6162 a_n1894_307.t20 a_n1894_307.n30 40.7345
R6163 a_n1894_307.n7 a_n1894_307.n6 28.094
R6164 a_n1894_307.n16 a_n1894_307.n15 28.094
R6165 a_n1894_307.n32 a_n1894_307.n31 28.094
R6166 a_n1894_307.n4 a_n1894_307.t28 21.9005
R6167 a_n1894_307.n2 a_n1894_307.t9 21.9005
R6168 a_n1894_307.n1 a_n1894_307.t16 21.9005
R6169 a_n1894_307.n10 a_n1894_307.t8 21.9005
R6170 a_n1894_307.n10 a_n1894_307.t6 21.9005
R6171 a_n1894_307.n22 a_n1894_307.t17 21.9005
R6172 a_n1894_307.n23 a_n1894_307.t11 21.9005
R6173 a_n1894_307.n11 a_n1894_307.t22 21.9005
R6174 a_n1894_307.n11 a_n1894_307.t25 21.9005
R6175 a_n1894_307.n3 a_n1894_307.t10 21.9005
R6176 a_n1894_307.n12 a_n1894_307.t27 21.9005
R6177 a_n1894_307.n12 a_n1894_307.t23 21.9005
R6178 a_n1894_307.n24 a_n1894_307.t12 21.9005
R6179 a_n1894_307.n25 a_n1894_307.t29 21.9005
R6180 a_n1894_307.n13 a_n1894_307.t15 21.9005
R6181 a_n1894_307.n13 a_n1894_307.t21 21.9005
R6182 a_n1894_307.n6 a_n1894_307.t19 21.9005
R6183 a_n1894_307.n15 a_n1894_307.t7 21.9005
R6184 a_n1894_307.n15 a_n1894_307.t13 21.9005
R6185 a_n1894_307.n5 a_n1894_307.t24 21.9005
R6186 a_n1894_307.n14 a_n1894_307.t18 21.9005
R6187 a_n1894_307.n14 a_n1894_307.t14 21.9005
R6188 a_n1894_307.n26 a_n1894_307.t26 21.9005
R6189 a_n1894_307.n31 a_n1894_307.t20 21.9005
R6190 a_n1894_307.n31 a_n1894_307.n26 15.8172
R6191 a_n1894_307.n14 a_n1894_307.n13 15.8172
R6192 a_n1894_307.n26 a_n1894_307.n25 15.8172
R6193 a_n1894_307.n25 a_n1894_307.n24 15.8172
R6194 a_n1894_307.n13 a_n1894_307.n12 15.8172
R6195 a_n1894_307.n12 a_n1894_307.n11 15.8172
R6196 a_n1894_307.n24 a_n1894_307.n23 15.8172
R6197 a_n1894_307.n23 a_n1894_307.n22 15.8172
R6198 a_n1894_307.n11 a_n1894_307.n10 15.8172
R6199 a_n1894_307.n2 a_n1894_307.n1 15.8172
R6200 a_n1894_307.n4 a_n1894_307.n3 15.8172
R6201 a_n1894_307.n3 a_n1894_307.n2 15.8172
R6202 a_n1894_307.n15 a_n1894_307.n14 15.8172
R6203 a_n1894_307.n6 a_n1894_307.n5 15.8172
R6204 a_n1894_307.n5 a_n1894_307.n4 15.8172
R6205 a_n1894_307.n28 a_n1894_307.n27 15.1845
R6206 a_n1894_307.n30 a_n1894_307.n29 15.1845
R6207 a_n1894_307.n29 a_n1894_307.n28 15.1845
R6208 a_n1894_307.n20 a_n1894_307.n19 5.44589
R6209 a_n1894_307.n20 a_n1894_307.n18 4.7885
R6210 a_n1894_307.n7 a_n1894_307.n0 4.70615
R6211 a_n1894_307.n21 a_n1894_307.n17 4.4205
R6212 a_n1894_307.n9 a_n1894_307.n8 4.4205
R6213 a_n1894_307.n34 a_n1894_307.n33 4.4205
R6214 a_n1894_307.n21 a_n1894_307.n20 1.1392
R6215 a_n1894_307.n16 a_n1894_307.n9 0.286152
R6216 a_n1894_307.n33 a_n1894_307.n32 0.286152
R6217 a_n1894_307.n32 a_n1894_307.n21 0.282239
R6218 a_n1894_307.n9 a_n1894_307.n7 0.282239
R6219 a_n1894_307.n33 a_n1894_307.n16 0.282239
R6220 A2.n47 A2.n45 5.44589
R6221 A2.n26 A2.n25 5.07789
R6222 A2.n51 A2.t31 4.7885
R6223 A2.n50 A2.t25 4.7885
R6224 A2.n47 A2.n46 4.7885
R6225 A2.n31 A2.t10 4.4205
R6226 A2.n32 A2.t16 4.4205
R6227 A2.n33 A2.t22 4.4205
R6228 A2.n34 A2.t9 4.4205
R6229 A2.n28 A2.n22 4.4205
R6230 A2.n27 A2.n23 4.4205
R6231 A2.n26 A2.n24 4.4205
R6232 A2.n44 A2.n41 3.80789
R6233 A2.n39 A2.n36 3.80789
R6234 A2.n53 A2 3.25827
R6235 A2.n8 A2.n7 3.25789
R6236 A2.n19 A2.n18 3.25789
R6237 A2.n44 A2.n43 3.1505
R6238 A2.n39 A2.n38 3.1505
R6239 A2.n8 A2.n5 2.6005
R6240 A2.n9 A2.n3 2.6005
R6241 A2.n10 A2.n1 2.6005
R6242 A2.n19 A2.n16 2.6005
R6243 A2.n20 A2.n14 2.6005
R6244 A2.n21 A2.n12 2.6005
R6245 A2.n1 A2.t1 1.8205
R6246 A2.n1 A2.n0 1.8205
R6247 A2.n3 A2.t8 1.8205
R6248 A2.n3 A2.n2 1.8205
R6249 A2.n5 A2.t14 1.8205
R6250 A2.n5 A2.n4 1.8205
R6251 A2.n7 A2.t0 1.8205
R6252 A2.n7 A2.n6 1.8205
R6253 A2.n12 A2.t20 1.8205
R6254 A2.n12 A2.n11 1.8205
R6255 A2.n14 A2.t4 1.8205
R6256 A2.n14 A2.n13 1.8205
R6257 A2.n16 A2.t7 1.8205
R6258 A2.n16 A2.n15 1.8205
R6259 A2.n18 A2.t18 1.8205
R6260 A2.n18 A2.n17 1.8205
R6261 A2.n43 A2.t29 1.6385
R6262 A2.n43 A2.n42 1.6385
R6263 A2.n41 A2.t35 1.6385
R6264 A2.n41 A2.n40 1.6385
R6265 A2.n38 A2.t34 1.6385
R6266 A2.n38 A2.n37 1.6385
R6267 A2.n36 A2.t28 1.6385
R6268 A2.n36 A2.n35 1.6385
R6269 A2.n53 A2.n52 1.32907
R6270 A2.n48 A2.n47 0.884196
R6271 A2.n50 A2.n49 0.884196
R6272 A2.n29 A2.n28 0.882239
R6273 A2.n31 A2.n30 0.882239
R6274 A2.n10 A2.n9 0.657891
R6275 A2.n9 A2.n8 0.657891
R6276 A2.n21 A2.n20 0.657891
R6277 A2.n20 A2.n19 0.657891
R6278 A2.n28 A2.n27 0.657891
R6279 A2.n27 A2.n26 0.657891
R6280 A2.n32 A2.n31 0.657891
R6281 A2.n33 A2.n32 0.657891
R6282 A2.n34 A2.n33 0.657891
R6283 A2.n51 A2.n50 0.657891
R6284 A2.n52 A2.n51 0.600532
R6285 A2.n30 A2.n29 0.6005
R6286 A2.n49 A2.n48 0.6005
R6287 A2.n48 A2.n44 0.284196
R6288 A2.n49 A2.n39 0.284196
R6289 A2.n30 A2.n10 0.282239
R6290 A2.n29 A2.n21 0.282239
R6291 A2.n52 A2.n34 0.278258
R6292 A2 A2.n53 0.219875
R6293 a_2004_1105.t23 a_2004_1105.n16 40.7345
R6294 a_2004_1105.n20 a_2004_1105.n5 28.094
R6295 a_2004_1105.n18 a_2004_1105.n17 28.094
R6296 a_2004_1105.n28 a_2004_1105.n27 28.094
R6297 a_2004_1105.n27 a_2004_1105.t22 21.9005
R6298 a_2004_1105.n25 a_2004_1105.t9 21.9005
R6299 a_2004_1105.n23 a_2004_1105.t17 21.9005
R6300 a_2004_1105.n22 a_2004_1105.t19 21.9005
R6301 a_2004_1105.n22 a_2004_1105.t14 21.9005
R6302 a_2004_1105.n0 a_2004_1105.t7 21.9005
R6303 a_2004_1105.n8 a_2004_1105.t20 21.9005
R6304 a_2004_1105.n9 a_2004_1105.t18 21.9005
R6305 a_2004_1105.n1 a_2004_1105.t6 21.9005
R6306 a_2004_1105.n23 a_2004_1105.t11 21.9005
R6307 a_2004_1105.n24 a_2004_1105.t12 21.9005
R6308 a_2004_1105.n24 a_2004_1105.t29 21.9005
R6309 a_2004_1105.n2 a_2004_1105.t25 21.9005
R6310 a_2004_1105.n10 a_2004_1105.t13 21.9005
R6311 a_2004_1105.n11 a_2004_1105.t10 21.9005
R6312 a_2004_1105.n3 a_2004_1105.t24 21.9005
R6313 a_2004_1105.n25 a_2004_1105.t26 21.9005
R6314 a_2004_1105.n26 a_2004_1105.t27 21.9005
R6315 a_2004_1105.n26 a_2004_1105.t21 21.9005
R6316 a_2004_1105.n4 a_2004_1105.t16 21.9005
R6317 a_2004_1105.n12 a_2004_1105.t28 21.9005
R6318 a_2004_1105.n17 a_2004_1105.t23 21.9005
R6319 a_2004_1105.n5 a_2004_1105.t8 21.9005
R6320 a_2004_1105.n27 a_2004_1105.t15 21.9005
R6321 a_2004_1105.n17 a_2004_1105.n12 15.8172
R6322 a_2004_1105.n5 a_2004_1105.n4 15.8172
R6323 a_2004_1105.n4 a_2004_1105.n3 15.8172
R6324 a_2004_1105.n12 a_2004_1105.n11 15.8172
R6325 a_2004_1105.n11 a_2004_1105.n10 15.8172
R6326 a_2004_1105.n3 a_2004_1105.n2 15.8172
R6327 a_2004_1105.n2 a_2004_1105.n1 15.8172
R6328 a_2004_1105.n10 a_2004_1105.n9 15.8172
R6329 a_2004_1105.n9 a_2004_1105.n8 15.8172
R6330 a_2004_1105.n1 a_2004_1105.n0 15.8172
R6331 a_2004_1105.n23 a_2004_1105.n22 15.8172
R6332 a_2004_1105.n24 a_2004_1105.n23 15.8172
R6333 a_2004_1105.n25 a_2004_1105.n24 15.8172
R6334 a_2004_1105.n26 a_2004_1105.n25 15.8172
R6335 a_2004_1105.n27 a_2004_1105.n26 15.8172
R6336 a_2004_1105.n14 a_2004_1105.n13 15.1845
R6337 a_2004_1105.n15 a_2004_1105.n14 15.1845
R6338 a_2004_1105.n16 a_2004_1105.n15 15.1845
R6339 a_2004_1105.n6 a_2004_1105.t5 5.44589
R6340 a_2004_1105.n6 a_2004_1105.t4 4.7885
R6341 a_2004_1105.t3 a_2004_1105.n28 4.70615
R6342 a_2004_1105.n7 a_2004_1105.t2 4.4205
R6343 a_2004_1105.n19 a_2004_1105.t1 4.4205
R6344 a_2004_1105.n21 a_2004_1105.t0 4.4205
R6345 a_2004_1105.n7 a_2004_1105.n6 1.1392
R6346 a_2004_1105.n21 a_2004_1105.n20 0.286152
R6347 a_2004_1105.n19 a_2004_1105.n18 0.286152
R6348 a_2004_1105.n28 a_2004_1105.n21 0.282239
R6349 a_2004_1105.n20 a_2004_1105.n19 0.282239
R6350 a_2004_1105.n18 a_2004_1105.n7 0.282239
R6351 TG_GATE_SWITCH_magic_4.B.n106 TG_GATE_SWITCH_magic_4.B.n52 5.6895
R6352 TG_GATE_SWITCH_magic_4.B.n95 TG_GATE_SWITCH_magic_4.B.n94 5.44589
R6353 TG_GATE_SWITCH_magic_4.B.n77 TG_GATE_SWITCH_magic_4.B.n75 5.07789
R6354 TG_GATE_SWITCH_magic_4.B.n104 TG_GATE_SWITCH_magic_4.B.t12 4.7885
R6355 TG_GATE_SWITCH_magic_4.B.n103 TG_GATE_SWITCH_magic_4.B.t15 4.7885
R6356 TG_GATE_SWITCH_magic_4.B.n95 TG_GATE_SWITCH_magic_4.B.n93 4.7885
R6357 TG_GATE_SWITCH_magic_4.B.n87 TG_GATE_SWITCH_magic_4.B.t34 4.4205
R6358 TG_GATE_SWITCH_magic_4.B.n86 TG_GATE_SWITCH_magic_4.B.t40 4.4205
R6359 TG_GATE_SWITCH_magic_4.B.n85 TG_GATE_SWITCH_magic_4.B.t49 4.4205
R6360 TG_GATE_SWITCH_magic_4.B.n84 TG_GATE_SWITCH_magic_4.B.t47 4.4205
R6361 TG_GATE_SWITCH_magic_4.B.n81 TG_GATE_SWITCH_magic_4.B.n80 4.4205
R6362 TG_GATE_SWITCH_magic_4.B.n79 TG_GATE_SWITCH_magic_4.B.n78 4.4205
R6363 TG_GATE_SWITCH_magic_4.B.n77 TG_GATE_SWITCH_magic_4.B.n76 4.4205
R6364 TG_GATE_SWITCH_magic_4.B.n27 TG_GATE_SWITCH_magic_4.B.n24 3.80789
R6365 TG_GATE_SWITCH_magic_4.B.n32 TG_GATE_SWITCH_magic_4.B.n29 3.80789
R6366 TG_GATE_SWITCH_magic_4.B.n37 TG_GATE_SWITCH_magic_4.B.n34 3.80789
R6367 TG_GATE_SWITCH_magic_4.B.n92 TG_GATE_SWITCH_magic_4.B.n91 3.80789
R6368 TG_GATE_SWITCH_magic_4.B.n101 TG_GATE_SWITCH_magic_4.B.n100 3.80789
R6369 TG_GATE_SWITCH_magic_4.B.n68 TG_GATE_SWITCH_magic_4.B.n65 3.25789
R6370 TG_GATE_SWITCH_magic_4.B.n57 TG_GATE_SWITCH_magic_4.B.n54 3.25789
R6371 TG_GATE_SWITCH_magic_4.B.n19 TG_GATE_SWITCH_magic_4.B.n18 3.25789
R6372 TG_GATE_SWITCH_magic_4.B.n8 TG_GATE_SWITCH_magic_4.B.n7 3.25789
R6373 TG_GATE_SWITCH_magic_4.B.n48 TG_GATE_SWITCH_magic_4.B.n47 3.25789
R6374 TG_GATE_SWITCH_magic_4.B.n27 TG_GATE_SWITCH_magic_4.B.n26 3.1505
R6375 TG_GATE_SWITCH_magic_4.B.n32 TG_GATE_SWITCH_magic_4.B.n31 3.1505
R6376 TG_GATE_SWITCH_magic_4.B.n37 TG_GATE_SWITCH_magic_4.B.n36 3.1505
R6377 TG_GATE_SWITCH_magic_4.B.n92 TG_GATE_SWITCH_magic_4.B.n89 3.1505
R6378 TG_GATE_SWITCH_magic_4.B.n101 TG_GATE_SWITCH_magic_4.B.n98 3.1505
R6379 TG_GATE_SWITCH_magic_4.B.n68 TG_GATE_SWITCH_magic_4.B.n67 2.6005
R6380 TG_GATE_SWITCH_magic_4.B.n71 TG_GATE_SWITCH_magic_4.B.n70 2.6005
R6381 TG_GATE_SWITCH_magic_4.B.n74 TG_GATE_SWITCH_magic_4.B.n73 2.6005
R6382 TG_GATE_SWITCH_magic_4.B.n57 TG_GATE_SWITCH_magic_4.B.n56 2.6005
R6383 TG_GATE_SWITCH_magic_4.B.n60 TG_GATE_SWITCH_magic_4.B.n59 2.6005
R6384 TG_GATE_SWITCH_magic_4.B.n63 TG_GATE_SWITCH_magic_4.B.n62 2.6005
R6385 TG_GATE_SWITCH_magic_4.B.n19 TG_GATE_SWITCH_magic_4.B.n16 2.6005
R6386 TG_GATE_SWITCH_magic_4.B.n20 TG_GATE_SWITCH_magic_4.B.n14 2.6005
R6387 TG_GATE_SWITCH_magic_4.B.n21 TG_GATE_SWITCH_magic_4.B.n12 2.6005
R6388 TG_GATE_SWITCH_magic_4.B.n8 TG_GATE_SWITCH_magic_4.B.n5 2.6005
R6389 TG_GATE_SWITCH_magic_4.B.n9 TG_GATE_SWITCH_magic_4.B.n3 2.6005
R6390 TG_GATE_SWITCH_magic_4.B.n10 TG_GATE_SWITCH_magic_4.B.n1 2.6005
R6391 TG_GATE_SWITCH_magic_4.B.n48 TG_GATE_SWITCH_magic_4.B.n45 2.6005
R6392 TG_GATE_SWITCH_magic_4.B.n49 TG_GATE_SWITCH_magic_4.B.n43 2.6005
R6393 TG_GATE_SWITCH_magic_4.B.n50 TG_GATE_SWITCH_magic_4.B.n41 2.6005
R6394 TG_GATE_SWITCH_magic_4.B.n73 TG_GATE_SWITCH_magic_4.B.t38 1.8205
R6395 TG_GATE_SWITCH_magic_4.B.n73 TG_GATE_SWITCH_magic_4.B.n72 1.8205
R6396 TG_GATE_SWITCH_magic_4.B.n70 TG_GATE_SWITCH_magic_4.B.t41 1.8205
R6397 TG_GATE_SWITCH_magic_4.B.n70 TG_GATE_SWITCH_magic_4.B.n69 1.8205
R6398 TG_GATE_SWITCH_magic_4.B.n67 TG_GATE_SWITCH_magic_4.B.t46 1.8205
R6399 TG_GATE_SWITCH_magic_4.B.n67 TG_GATE_SWITCH_magic_4.B.n66 1.8205
R6400 TG_GATE_SWITCH_magic_4.B.n65 TG_GATE_SWITCH_magic_4.B.t2 1.8205
R6401 TG_GATE_SWITCH_magic_4.B.n65 TG_GATE_SWITCH_magic_4.B.n64 1.8205
R6402 TG_GATE_SWITCH_magic_4.B.n62 TG_GATE_SWITCH_magic_4.B.t53 1.8205
R6403 TG_GATE_SWITCH_magic_4.B.n62 TG_GATE_SWITCH_magic_4.B.n61 1.8205
R6404 TG_GATE_SWITCH_magic_4.B.n59 TG_GATE_SWITCH_magic_4.B.t54 1.8205
R6405 TG_GATE_SWITCH_magic_4.B.n59 TG_GATE_SWITCH_magic_4.B.n58 1.8205
R6406 TG_GATE_SWITCH_magic_4.B.n56 TG_GATE_SWITCH_magic_4.B.t0 1.8205
R6407 TG_GATE_SWITCH_magic_4.B.n56 TG_GATE_SWITCH_magic_4.B.n55 1.8205
R6408 TG_GATE_SWITCH_magic_4.B.n54 TG_GATE_SWITCH_magic_4.B.t43 1.8205
R6409 TG_GATE_SWITCH_magic_4.B.n54 TG_GATE_SWITCH_magic_4.B.n53 1.8205
R6410 TG_GATE_SWITCH_magic_4.B.n12 TG_GATE_SWITCH_magic_4.B.t68 1.8205
R6411 TG_GATE_SWITCH_magic_4.B.n12 TG_GATE_SWITCH_magic_4.B.n11 1.8205
R6412 TG_GATE_SWITCH_magic_4.B.n14 TG_GATE_SWITCH_magic_4.B.t70 1.8205
R6413 TG_GATE_SWITCH_magic_4.B.n14 TG_GATE_SWITCH_magic_4.B.n13 1.8205
R6414 TG_GATE_SWITCH_magic_4.B.n16 TG_GATE_SWITCH_magic_4.B.t66 1.8205
R6415 TG_GATE_SWITCH_magic_4.B.n16 TG_GATE_SWITCH_magic_4.B.n15 1.8205
R6416 TG_GATE_SWITCH_magic_4.B.n18 TG_GATE_SWITCH_magic_4.B.t45 1.8205
R6417 TG_GATE_SWITCH_magic_4.B.n18 TG_GATE_SWITCH_magic_4.B.n17 1.8205
R6418 TG_GATE_SWITCH_magic_4.B.n1 TG_GATE_SWITCH_magic_4.B.t6 1.8205
R6419 TG_GATE_SWITCH_magic_4.B.n1 TG_GATE_SWITCH_magic_4.B.n0 1.8205
R6420 TG_GATE_SWITCH_magic_4.B.n3 TG_GATE_SWITCH_magic_4.B.t67 1.8205
R6421 TG_GATE_SWITCH_magic_4.B.n3 TG_GATE_SWITCH_magic_4.B.n2 1.8205
R6422 TG_GATE_SWITCH_magic_4.B.n5 TG_GATE_SWITCH_magic_4.B.t59 1.8205
R6423 TG_GATE_SWITCH_magic_4.B.n5 TG_GATE_SWITCH_magic_4.B.n4 1.8205
R6424 TG_GATE_SWITCH_magic_4.B.n7 TG_GATE_SWITCH_magic_4.B.t4 1.8205
R6425 TG_GATE_SWITCH_magic_4.B.n7 TG_GATE_SWITCH_magic_4.B.n6 1.8205
R6426 TG_GATE_SWITCH_magic_4.B.n41 TG_GATE_SWITCH_magic_4.B.t64 1.8205
R6427 TG_GATE_SWITCH_magic_4.B.n41 TG_GATE_SWITCH_magic_4.B.n40 1.8205
R6428 TG_GATE_SWITCH_magic_4.B.n43 TG_GATE_SWITCH_magic_4.B.t3 1.8205
R6429 TG_GATE_SWITCH_magic_4.B.n43 TG_GATE_SWITCH_magic_4.B.n42 1.8205
R6430 TG_GATE_SWITCH_magic_4.B.n45 TG_GATE_SWITCH_magic_4.B.t71 1.8205
R6431 TG_GATE_SWITCH_magic_4.B.n45 TG_GATE_SWITCH_magic_4.B.n44 1.8205
R6432 TG_GATE_SWITCH_magic_4.B.n47 TG_GATE_SWITCH_magic_4.B.t61 1.8205
R6433 TG_GATE_SWITCH_magic_4.B.n47 TG_GATE_SWITCH_magic_4.B.n46 1.8205
R6434 TG_GATE_SWITCH_magic_4.B.n98 TG_GATE_SWITCH_magic_4.B.t10 1.6385
R6435 TG_GATE_SWITCH_magic_4.B.n98 TG_GATE_SWITCH_magic_4.B.n97 1.6385
R6436 TG_GATE_SWITCH_magic_4.B.n26 TG_GATE_SWITCH_magic_4.B.t30 1.6385
R6437 TG_GATE_SWITCH_magic_4.B.n26 TG_GATE_SWITCH_magic_4.B.n25 1.6385
R6438 TG_GATE_SWITCH_magic_4.B.n24 TG_GATE_SWITCH_magic_4.B.t27 1.6385
R6439 TG_GATE_SWITCH_magic_4.B.n24 TG_GATE_SWITCH_magic_4.B.n23 1.6385
R6440 TG_GATE_SWITCH_magic_4.B.n31 TG_GATE_SWITCH_magic_4.B.t29 1.6385
R6441 TG_GATE_SWITCH_magic_4.B.n31 TG_GATE_SWITCH_magic_4.B.n30 1.6385
R6442 TG_GATE_SWITCH_magic_4.B.n29 TG_GATE_SWITCH_magic_4.B.t26 1.6385
R6443 TG_GATE_SWITCH_magic_4.B.n29 TG_GATE_SWITCH_magic_4.B.n28 1.6385
R6444 TG_GATE_SWITCH_magic_4.B.n34 TG_GATE_SWITCH_magic_4.B.t31 1.6385
R6445 TG_GATE_SWITCH_magic_4.B.n34 TG_GATE_SWITCH_magic_4.B.n33 1.6385
R6446 TG_GATE_SWITCH_magic_4.B.n36 TG_GATE_SWITCH_magic_4.B.t28 1.6385
R6447 TG_GATE_SWITCH_magic_4.B.n36 TG_GATE_SWITCH_magic_4.B.n35 1.6385
R6448 TG_GATE_SWITCH_magic_4.B.n89 TG_GATE_SWITCH_magic_4.B.t18 1.6385
R6449 TG_GATE_SWITCH_magic_4.B.n89 TG_GATE_SWITCH_magic_4.B.n88 1.6385
R6450 TG_GATE_SWITCH_magic_4.B.n91 TG_GATE_SWITCH_magic_4.B.t16 1.6385
R6451 TG_GATE_SWITCH_magic_4.B.n91 TG_GATE_SWITCH_magic_4.B.n90 1.6385
R6452 TG_GATE_SWITCH_magic_4.B.n100 TG_GATE_SWITCH_magic_4.B.t20 1.6385
R6453 TG_GATE_SWITCH_magic_4.B.n100 TG_GATE_SWITCH_magic_4.B.n99 1.6385
R6454 TG_GATE_SWITCH_magic_4.B.n106 TG_GATE_SWITCH_magic_4.B.n105 1.58607
R6455 TG_GATE_SWITCH_magic_4.B TG_GATE_SWITCH_magic_4.B.n106 1.17023
R6456 TG_GATE_SWITCH_magic_4.B.n103 TG_GATE_SWITCH_magic_4.B.n102 0.884196
R6457 TG_GATE_SWITCH_magic_4.B.n96 TG_GATE_SWITCH_magic_4.B.n95 0.884196
R6458 TG_GATE_SWITCH_magic_4.B.n82 TG_GATE_SWITCH_magic_4.B.n81 0.882239
R6459 TG_GATE_SWITCH_magic_4.B.n84 TG_GATE_SWITCH_magic_4.B.n83 0.882239
R6460 TG_GATE_SWITCH_magic_4.B.n105 TG_GATE_SWITCH_magic_4.B.n104 0.8105
R6461 TG_GATE_SWITCH_magic_4.B.n79 TG_GATE_SWITCH_magic_4.B.n77 0.657891
R6462 TG_GATE_SWITCH_magic_4.B.n81 TG_GATE_SWITCH_magic_4.B.n79 0.657891
R6463 TG_GATE_SWITCH_magic_4.B.n71 TG_GATE_SWITCH_magic_4.B.n68 0.657891
R6464 TG_GATE_SWITCH_magic_4.B.n74 TG_GATE_SWITCH_magic_4.B.n71 0.657891
R6465 TG_GATE_SWITCH_magic_4.B.n60 TG_GATE_SWITCH_magic_4.B.n57 0.657891
R6466 TG_GATE_SWITCH_magic_4.B.n63 TG_GATE_SWITCH_magic_4.B.n60 0.657891
R6467 TG_GATE_SWITCH_magic_4.B.n87 TG_GATE_SWITCH_magic_4.B.n86 0.657891
R6468 TG_GATE_SWITCH_magic_4.B.n86 TG_GATE_SWITCH_magic_4.B.n85 0.657891
R6469 TG_GATE_SWITCH_magic_4.B.n85 TG_GATE_SWITCH_magic_4.B.n84 0.657891
R6470 TG_GATE_SWITCH_magic_4.B.n20 TG_GATE_SWITCH_magic_4.B.n19 0.657891
R6471 TG_GATE_SWITCH_magic_4.B.n10 TG_GATE_SWITCH_magic_4.B.n9 0.657891
R6472 TG_GATE_SWITCH_magic_4.B.n9 TG_GATE_SWITCH_magic_4.B.n8 0.657891
R6473 TG_GATE_SWITCH_magic_4.B.n50 TG_GATE_SWITCH_magic_4.B.n49 0.657891
R6474 TG_GATE_SWITCH_magic_4.B.n49 TG_GATE_SWITCH_magic_4.B.n48 0.657891
R6475 TG_GATE_SWITCH_magic_4.B.n104 TG_GATE_SWITCH_magic_4.B.n103 0.657891
R6476 TG_GATE_SWITCH_magic_4.B.n21 TG_GATE_SWITCH_magic_4.B.n20 0.655976
R6477 TG_GATE_SWITCH_magic_4.B.n22 TG_GATE_SWITCH_magic_4.B.n21 0.645657
R6478 TG_GATE_SWITCH_magic_4.B.n83 TG_GATE_SWITCH_magic_4.B.n82 0.6005
R6479 TG_GATE_SWITCH_magic_4.B.n102 TG_GATE_SWITCH_magic_4.B.n96 0.6005
R6480 TG_GATE_SWITCH_magic_4.B.n38 TG_GATE_SWITCH_magic_4.B.n37 0.548416
R6481 TG_GATE_SWITCH_magic_4.B.n51 TG_GATE_SWITCH_magic_4.B.n50 0.316429
R6482 TG_GATE_SWITCH_magic_4.B.n39 TG_GATE_SWITCH_magic_4.B.n27 0.304838
R6483 TG_GATE_SWITCH_magic_4.B.n38 TG_GATE_SWITCH_magic_4.B.n32 0.284196
R6484 TG_GATE_SWITCH_magic_4.B.n96 TG_GATE_SWITCH_magic_4.B.n92 0.284196
R6485 TG_GATE_SWITCH_magic_4.B.n102 TG_GATE_SWITCH_magic_4.B.n101 0.284196
R6486 TG_GATE_SWITCH_magic_4.B.n51 TG_GATE_SWITCH_magic_4.B.n22 0.283032
R6487 TG_GATE_SWITCH_magic_4.B.n82 TG_GATE_SWITCH_magic_4.B.n74 0.282239
R6488 TG_GATE_SWITCH_magic_4.B.n83 TG_GATE_SWITCH_magic_4.B.n63 0.282239
R6489 TG_GATE_SWITCH_magic_4.B.n22 TG_GATE_SWITCH_magic_4.B.n10 0.279866
R6490 TG_GATE_SWITCH_magic_4.B.n52 TG_GATE_SWITCH_magic_4.B.n51 0.245695
R6491 TG_GATE_SWITCH_magic_4.B.n39 TG_GATE_SWITCH_magic_4.B.n38 0.244078
R6492 TG_GATE_SWITCH_magic_4.B.n105 TG_GATE_SWITCH_magic_4.B.n87 0.237239
R6493 TG_GATE_SWITCH_magic_4.B.n51 TG_GATE_SWITCH_magic_4.B.n39 0.136437
R6494 TG_GATE_SWITCH_magic_4.B.n52 TG_GATE_SWITCH_magic_4.B 0.0416746
R6495 a_3874_n7430.t19 a_3874_n7430.n30 40.7345
R6496 a_3874_n7430.n20 a_3874_n7430.n9 28.094
R6497 a_3874_n7430.n18 a_3874_n7430.n17 28.094
R6498 a_3874_n7430.n32 a_3874_n7430.n31 28.094
R6499 a_3874_n7430.n22 a_3874_n7430.t22 21.9005
R6500 a_3874_n7430.n22 a_3874_n7430.t29 21.9005
R6501 a_3874_n7430.n4 a_3874_n7430.t16 21.9005
R6502 a_3874_n7430.n12 a_3874_n7430.t15 21.9005
R6503 a_3874_n7430.n13 a_3874_n7430.t23 21.9005
R6504 a_3874_n7430.n5 a_3874_n7430.t26 21.9005
R6505 a_3874_n7430.n23 a_3874_n7430.t10 21.9005
R6506 a_3874_n7430.n23 a_3874_n7430.t8 21.9005
R6507 a_3874_n7430.n24 a_3874_n7430.t20 21.9005
R6508 a_3874_n7430.n24 a_3874_n7430.t27 21.9005
R6509 a_3874_n7430.n6 a_3874_n7430.t14 21.9005
R6510 a_3874_n7430.n14 a_3874_n7430.t12 21.9005
R6511 a_3874_n7430.n15 a_3874_n7430.t17 21.9005
R6512 a_3874_n7430.n7 a_3874_n7430.t18 21.9005
R6513 a_3874_n7430.n25 a_3874_n7430.t6 21.9005
R6514 a_3874_n7430.n25 a_3874_n7430.t28 21.9005
R6515 a_3874_n7430.n31 a_3874_n7430.t19 21.9005
R6516 a_3874_n7430.n26 a_3874_n7430.t7 21.9005
R6517 a_3874_n7430.n26 a_3874_n7430.t9 21.9005
R6518 a_3874_n7430.n8 a_3874_n7430.t24 21.9005
R6519 a_3874_n7430.n16 a_3874_n7430.t21 21.9005
R6520 a_3874_n7430.n17 a_3874_n7430.t11 21.9005
R6521 a_3874_n7430.n9 a_3874_n7430.t13 21.9005
R6522 a_3874_n7430.n31 a_3874_n7430.t25 21.9005
R6523 a_3874_n7430.n9 a_3874_n7430.n8 15.8172
R6524 a_3874_n7430.n31 a_3874_n7430.n26 15.8172
R6525 a_3874_n7430.n26 a_3874_n7430.n25 15.8172
R6526 a_3874_n7430.n8 a_3874_n7430.n7 15.8172
R6527 a_3874_n7430.n7 a_3874_n7430.n6 15.8172
R6528 a_3874_n7430.n25 a_3874_n7430.n24 15.8172
R6529 a_3874_n7430.n24 a_3874_n7430.n23 15.8172
R6530 a_3874_n7430.n6 a_3874_n7430.n5 15.8172
R6531 a_3874_n7430.n5 a_3874_n7430.n4 15.8172
R6532 a_3874_n7430.n23 a_3874_n7430.n22 15.8172
R6533 a_3874_n7430.n14 a_3874_n7430.n13 15.8172
R6534 a_3874_n7430.n13 a_3874_n7430.n12 15.8172
R6535 a_3874_n7430.n16 a_3874_n7430.n15 15.8172
R6536 a_3874_n7430.n15 a_3874_n7430.n14 15.8172
R6537 a_3874_n7430.n17 a_3874_n7430.n16 15.8172
R6538 a_3874_n7430.n29 a_3874_n7430.n28 15.1845
R6539 a_3874_n7430.n28 a_3874_n7430.n27 15.1845
R6540 a_3874_n7430.n30 a_3874_n7430.n29 15.1845
R6541 a_3874_n7430.n2 a_3874_n7430.n0 5.44589
R6542 a_3874_n7430.n2 a_3874_n7430.n1 4.7885
R6543 a_3874_n7430.n18 a_3874_n7430.n11 4.70615
R6544 a_3874_n7430.n19 a_3874_n7430.n10 4.4205
R6545 a_3874_n7430.n21 a_3874_n7430.n3 4.4205
R6546 a_3874_n7430.n34 a_3874_n7430.n33 4.4205
R6547 a_3874_n7430.n33 a_3874_n7430.n2 1.1392
R6548 a_3874_n7430.n32 a_3874_n7430.n21 0.286152
R6549 a_3874_n7430.n20 a_3874_n7430.n19 0.286152
R6550 a_3874_n7430.n21 a_3874_n7430.n20 0.282239
R6551 a_3874_n7430.n19 a_3874_n7430.n18 0.282239
R6552 a_3874_n7430.n33 a_3874_n7430.n32 0.282239
R6553 a_3817_n4055.t16 a_3817_n4055.n17 40.7345
R6554 a_3817_n4055.n19 a_3817_n4055.n18 28.094
R6555 a_3817_n4055.n6 a_3817_n4055.n5 28.094
R6556 a_3817_n4055.n27 a_3817_n4055.n26 28.094
R6557 a_3817_n4055.n5 a_3817_n4055.t17 21.9005
R6558 a_3817_n4055.n5 a_3817_n4055.t28 21.9005
R6559 a_3817_n4055.n3 a_3817_n4055.t26 21.9005
R6560 a_3817_n4055.n1 a_3817_n4055.t23 21.9005
R6561 a_3817_n4055.n0 a_3817_n4055.t11 21.9005
R6562 a_3817_n4055.n0 a_3817_n4055.t24 21.9005
R6563 a_3817_n4055.n21 a_3817_n4055.t29 21.9005
R6564 a_3817_n4055.n9 a_3817_n4055.t9 21.9005
R6565 a_3817_n4055.n10 a_3817_n4055.t22 21.9005
R6566 a_3817_n4055.n22 a_3817_n4055.t18 21.9005
R6567 a_3817_n4055.n1 a_3817_n4055.t10 21.9005
R6568 a_3817_n4055.n2 a_3817_n4055.t15 21.9005
R6569 a_3817_n4055.n2 a_3817_n4055.t27 21.9005
R6570 a_3817_n4055.n23 a_3817_n4055.t6 21.9005
R6571 a_3817_n4055.n11 a_3817_n4055.t13 21.9005
R6572 a_3817_n4055.n12 a_3817_n4055.t25 21.9005
R6573 a_3817_n4055.n24 a_3817_n4055.t19 21.9005
R6574 a_3817_n4055.n3 a_3817_n4055.t14 21.9005
R6575 a_3817_n4055.n4 a_3817_n4055.t21 21.9005
R6576 a_3817_n4055.n4 a_3817_n4055.t8 21.9005
R6577 a_3817_n4055.n25 a_3817_n4055.t12 21.9005
R6578 a_3817_n4055.n13 a_3817_n4055.t20 21.9005
R6579 a_3817_n4055.n18 a_3817_n4055.t16 21.9005
R6580 a_3817_n4055.n26 a_3817_n4055.t7 21.9005
R6581 a_3817_n4055.n18 a_3817_n4055.n13 15.8172
R6582 a_3817_n4055.n26 a_3817_n4055.n25 15.8172
R6583 a_3817_n4055.n25 a_3817_n4055.n24 15.8172
R6584 a_3817_n4055.n13 a_3817_n4055.n12 15.8172
R6585 a_3817_n4055.n12 a_3817_n4055.n11 15.8172
R6586 a_3817_n4055.n24 a_3817_n4055.n23 15.8172
R6587 a_3817_n4055.n23 a_3817_n4055.n22 15.8172
R6588 a_3817_n4055.n11 a_3817_n4055.n10 15.8172
R6589 a_3817_n4055.n10 a_3817_n4055.n9 15.8172
R6590 a_3817_n4055.n22 a_3817_n4055.n21 15.8172
R6591 a_3817_n4055.n1 a_3817_n4055.n0 15.8172
R6592 a_3817_n4055.n2 a_3817_n4055.n1 15.8172
R6593 a_3817_n4055.n3 a_3817_n4055.n2 15.8172
R6594 a_3817_n4055.n4 a_3817_n4055.n3 15.8172
R6595 a_3817_n4055.n5 a_3817_n4055.n4 15.8172
R6596 a_3817_n4055.n15 a_3817_n4055.n14 15.1845
R6597 a_3817_n4055.n16 a_3817_n4055.n15 15.1845
R6598 a_3817_n4055.n17 a_3817_n4055.n16 15.1845
R6599 a_3817_n4055.n7 a_3817_n4055.t4 5.44589
R6600 a_3817_n4055.n7 a_3817_n4055.t5 4.7885
R6601 a_3817_n4055.n6 a_3817_n4055.t0 4.70615
R6602 a_3817_n4055.n8 a_3817_n4055.t1 4.4205
R6603 a_3817_n4055.n20 a_3817_n4055.t2 4.4205
R6604 a_3817_n4055.t3 a_3817_n4055.n28 4.4205
R6605 a_3817_n4055.n8 a_3817_n4055.n7 1.1392
R6606 a_3817_n4055.n20 a_3817_n4055.n19 0.286152
R6607 a_3817_n4055.n28 a_3817_n4055.n27 0.286152
R6608 a_3817_n4055.n27 a_3817_n4055.n20 0.282239
R6609 a_3817_n4055.n19 a_3817_n4055.n8 0.282239
R6610 a_3817_n4055.n28 a_3817_n4055.n6 0.282239
R6611 a_n1894_n4853.t27 a_n1894_n4853.n22 40.7345
R6612 a_n1894_n4853.n24 a_n1894_n4853.n23 28.094
R6613 a_n1894_n4853.n7 a_n1894_n4853.n6 28.094
R6614 a_n1894_n4853.n32 a_n1894_n4853.n31 28.094
R6615 a_n1894_n4853.n4 a_n1894_n4853.t23 21.9005
R6616 a_n1894_n4853.n2 a_n1894_n4853.t15 21.9005
R6617 a_n1894_n4853.n1 a_n1894_n4853.t22 21.9005
R6618 a_n1894_n4853.n1 a_n1894_n4853.t9 21.9005
R6619 a_n1894_n4853.n26 a_n1894_n4853.t11 21.9005
R6620 a_n1894_n4853.n14 a_n1894_n4853.t18 21.9005
R6621 a_n1894_n4853.n15 a_n1894_n4853.t14 21.9005
R6622 a_n1894_n4853.n27 a_n1894_n4853.t8 21.9005
R6623 a_n1894_n4853.n2 a_n1894_n4853.t29 21.9005
R6624 a_n1894_n4853.n3 a_n1894_n4853.t26 21.9005
R6625 a_n1894_n4853.n3 a_n1894_n4853.t13 21.9005
R6626 a_n1894_n4853.n28 a_n1894_n4853.t17 21.9005
R6627 a_n1894_n4853.n16 a_n1894_n4853.t25 21.9005
R6628 a_n1894_n4853.n17 a_n1894_n4853.t20 21.9005
R6629 a_n1894_n4853.n29 a_n1894_n4853.t12 21.9005
R6630 a_n1894_n4853.n4 a_n1894_n4853.t10 21.9005
R6631 a_n1894_n4853.n6 a_n1894_n4853.t28 21.9005
R6632 a_n1894_n4853.n6 a_n1894_n4853.t16 21.9005
R6633 a_n1894_n4853.n5 a_n1894_n4853.t7 21.9005
R6634 a_n1894_n4853.n5 a_n1894_n4853.t21 21.9005
R6635 a_n1894_n4853.n30 a_n1894_n4853.t24 21.9005
R6636 a_n1894_n4853.n18 a_n1894_n4853.t6 21.9005
R6637 a_n1894_n4853.n23 a_n1894_n4853.t27 21.9005
R6638 a_n1894_n4853.n31 a_n1894_n4853.t19 21.9005
R6639 a_n1894_n4853.n23 a_n1894_n4853.n18 15.8172
R6640 a_n1894_n4853.n31 a_n1894_n4853.n30 15.8172
R6641 a_n1894_n4853.n30 a_n1894_n4853.n29 15.8172
R6642 a_n1894_n4853.n18 a_n1894_n4853.n17 15.8172
R6643 a_n1894_n4853.n17 a_n1894_n4853.n16 15.8172
R6644 a_n1894_n4853.n29 a_n1894_n4853.n28 15.8172
R6645 a_n1894_n4853.n28 a_n1894_n4853.n27 15.8172
R6646 a_n1894_n4853.n16 a_n1894_n4853.n15 15.8172
R6647 a_n1894_n4853.n15 a_n1894_n4853.n14 15.8172
R6648 a_n1894_n4853.n27 a_n1894_n4853.n26 15.8172
R6649 a_n1894_n4853.n2 a_n1894_n4853.n1 15.8172
R6650 a_n1894_n4853.n4 a_n1894_n4853.n3 15.8172
R6651 a_n1894_n4853.n3 a_n1894_n4853.n2 15.8172
R6652 a_n1894_n4853.n6 a_n1894_n4853.n5 15.8172
R6653 a_n1894_n4853.n5 a_n1894_n4853.n4 15.8172
R6654 a_n1894_n4853.n20 a_n1894_n4853.n19 15.1845
R6655 a_n1894_n4853.n22 a_n1894_n4853.n21 15.1845
R6656 a_n1894_n4853.n21 a_n1894_n4853.n20 15.1845
R6657 a_n1894_n4853.n12 a_n1894_n4853.n11 5.44589
R6658 a_n1894_n4853.n12 a_n1894_n4853.n10 4.7885
R6659 a_n1894_n4853.n7 a_n1894_n4853.n0 4.70615
R6660 a_n1894_n4853.n13 a_n1894_n4853.n9 4.4205
R6661 a_n1894_n4853.n25 a_n1894_n4853.n8 4.4205
R6662 a_n1894_n4853.n34 a_n1894_n4853.n33 4.4205
R6663 a_n1894_n4853.n13 a_n1894_n4853.n12 1.1392
R6664 a_n1894_n4853.n25 a_n1894_n4853.n24 0.286152
R6665 a_n1894_n4853.n33 a_n1894_n4853.n32 0.286152
R6666 a_n1894_n4853.n32 a_n1894_n4853.n25 0.282239
R6667 a_n1894_n4853.n24 a_n1894_n4853.n13 0.282239
R6668 a_n1894_n4853.n33 a_n1894_n4853.n7 0.282239
R6669 a_n1894_n7431.t29 a_n1894_n7431.n19 40.7345
R6670 a_n1894_n7431.n24 a_n1894_n7431.n5 28.094
R6671 a_n1894_n7431.n21 a_n1894_n7431.n20 28.094
R6672 a_n1894_n7431.n32 a_n1894_n7431.n31 28.094
R6673 a_n1894_n7431.n26 a_n1894_n7431.t18 21.9005
R6674 a_n1894_n7431.n26 a_n1894_n7431.t12 21.9005
R6675 a_n1894_n7431.n0 a_n1894_n7431.t24 21.9005
R6676 a_n1894_n7431.n11 a_n1894_n7431.t21 21.9005
R6677 a_n1894_n7431.n12 a_n1894_n7431.t15 21.9005
R6678 a_n1894_n7431.n1 a_n1894_n7431.t19 21.9005
R6679 a_n1894_n7431.n27 a_n1894_n7431.t10 21.9005
R6680 a_n1894_n7431.n27 a_n1894_n7431.t14 21.9005
R6681 a_n1894_n7431.n28 a_n1894_n7431.t25 21.9005
R6682 a_n1894_n7431.n28 a_n1894_n7431.t16 21.9005
R6683 a_n1894_n7431.n2 a_n1894_n7431.t6 21.9005
R6684 a_n1894_n7431.n13 a_n1894_n7431.t27 21.9005
R6685 a_n1894_n7431.n14 a_n1894_n7431.t22 21.9005
R6686 a_n1894_n7431.n3 a_n1894_n7431.t26 21.9005
R6687 a_n1894_n7431.n29 a_n1894_n7431.t13 21.9005
R6688 a_n1894_n7431.n29 a_n1894_n7431.t20 21.9005
R6689 a_n1894_n7431.n30 a_n1894_n7431.t7 21.9005
R6690 a_n1894_n7431.n30 a_n1894_n7431.t23 21.9005
R6691 a_n1894_n7431.n4 a_n1894_n7431.t11 21.9005
R6692 a_n1894_n7431.n15 a_n1894_n7431.t9 21.9005
R6693 a_n1894_n7431.n20 a_n1894_n7431.t29 21.9005
R6694 a_n1894_n7431.n5 a_n1894_n7431.t8 21.9005
R6695 a_n1894_n7431.n31 a_n1894_n7431.t17 21.9005
R6696 a_n1894_n7431.n31 a_n1894_n7431.t28 21.9005
R6697 a_n1894_n7431.n20 a_n1894_n7431.n15 15.8172
R6698 a_n1894_n7431.n5 a_n1894_n7431.n4 15.8172
R6699 a_n1894_n7431.n4 a_n1894_n7431.n3 15.8172
R6700 a_n1894_n7431.n15 a_n1894_n7431.n14 15.8172
R6701 a_n1894_n7431.n14 a_n1894_n7431.n13 15.8172
R6702 a_n1894_n7431.n3 a_n1894_n7431.n2 15.8172
R6703 a_n1894_n7431.n2 a_n1894_n7431.n1 15.8172
R6704 a_n1894_n7431.n13 a_n1894_n7431.n12 15.8172
R6705 a_n1894_n7431.n12 a_n1894_n7431.n11 15.8172
R6706 a_n1894_n7431.n1 a_n1894_n7431.n0 15.8172
R6707 a_n1894_n7431.n27 a_n1894_n7431.n26 15.8172
R6708 a_n1894_n7431.n29 a_n1894_n7431.n28 15.8172
R6709 a_n1894_n7431.n28 a_n1894_n7431.n27 15.8172
R6710 a_n1894_n7431.n31 a_n1894_n7431.n30 15.8172
R6711 a_n1894_n7431.n30 a_n1894_n7431.n29 15.8172
R6712 a_n1894_n7431.n17 a_n1894_n7431.n16 15.1845
R6713 a_n1894_n7431.n19 a_n1894_n7431.n18 15.1845
R6714 a_n1894_n7431.n18 a_n1894_n7431.n17 15.1845
R6715 a_n1894_n7431.n8 a_n1894_n7431.n6 5.44589
R6716 a_n1894_n7431.n8 a_n1894_n7431.n7 4.7885
R6717 a_n1894_n7431.n32 a_n1894_n7431.n25 4.70615
R6718 a_n1894_n7431.n23 a_n1894_n7431.n22 4.4205
R6719 a_n1894_n7431.n10 a_n1894_n7431.n9 4.4205
R6720 a_n1894_n7431.n34 a_n1894_n7431.n33 4.4205
R6721 a_n1894_n7431.n10 a_n1894_n7431.n8 1.1392
R6722 a_n1894_n7431.n23 a_n1894_n7431.n21 0.286152
R6723 a_n1894_n7431.n33 a_n1894_n7431.n24 0.286152
R6724 a_n1894_n7431.n21 a_n1894_n7431.n10 0.282239
R6725 a_n1894_n7431.n24 a_n1894_n7431.n23 0.282239
R6726 a_n1894_n7431.n33 a_n1894_n7431.n32 0.282239
R6727 A1.n47 A1.n46 5.44589
R6728 A1.n24 A1.n22 5.07789
R6729 A1.n50 A1.t1 4.7885
R6730 A1.n51 A1.t7 4.7885
R6731 A1.n47 A1.n45 4.7885
R6732 A1.n34 A1.t12 4.4205
R6733 A1.n33 A1.t33 4.4205
R6734 A1.n32 A1.t24 4.4205
R6735 A1.n31 A1.t13 4.4205
R6736 A1.n28 A1.n27 4.4205
R6737 A1.n26 A1.n25 4.4205
R6738 A1.n24 A1.n23 4.4205
R6739 A1.n53 A1 4.04383
R6740 A1.n39 A1.n38 3.80789
R6741 A1.n44 A1.n43 3.80789
R6742 A1.n15 A1.n12 3.25789
R6743 A1.n4 A1.n1 3.25789
R6744 A1.n39 A1.n36 3.1505
R6745 A1.n44 A1.n41 3.1505
R6746 A1.n15 A1.n14 2.6005
R6747 A1.n18 A1.n17 2.6005
R6748 A1.n21 A1.n20 2.6005
R6749 A1.n4 A1.n3 2.6005
R6750 A1.n7 A1.n6 2.6005
R6751 A1.n10 A1.n9 2.6005
R6752 A1.n20 A1.t27 1.8205
R6753 A1.n20 A1.n19 1.8205
R6754 A1.n17 A1.t31 1.8205
R6755 A1.n17 A1.n16 1.8205
R6756 A1.n14 A1.t22 1.8205
R6757 A1.n14 A1.n13 1.8205
R6758 A1.n12 A1.t26 1.8205
R6759 A1.n12 A1.n11 1.8205
R6760 A1.n9 A1.t21 1.8205
R6761 A1.n9 A1.n8 1.8205
R6762 A1.n6 A1.t28 1.8205
R6763 A1.n6 A1.n5 1.8205
R6764 A1.n3 A1.t15 1.8205
R6765 A1.n3 A1.n2 1.8205
R6766 A1.n1 A1.t19 1.8205
R6767 A1.n1 A1.n0 1.8205
R6768 A1.n36 A1.t3 1.6385
R6769 A1.n36 A1.n35 1.6385
R6770 A1.n38 A1.t9 1.6385
R6771 A1.n38 A1.n37 1.6385
R6772 A1.n41 A1.t6 1.6385
R6773 A1.n41 A1.n40 1.6385
R6774 A1.n43 A1.t0 1.6385
R6775 A1.n43 A1.n42 1.6385
R6776 A1.n53 A1.n52 1.36224
R6777 A1.n48 A1.n47 0.884196
R6778 A1.n50 A1.n49 0.884196
R6779 A1.n29 A1.n28 0.882239
R6780 A1.n31 A1.n30 0.882239
R6781 A1.n51 A1.n50 0.657891
R6782 A1.n26 A1.n24 0.657891
R6783 A1.n28 A1.n26 0.657891
R6784 A1.n18 A1.n15 0.657891
R6785 A1.n21 A1.n18 0.657891
R6786 A1.n7 A1.n4 0.657891
R6787 A1.n10 A1.n7 0.657891
R6788 A1.n34 A1.n33 0.657891
R6789 A1.n33 A1.n32 0.657891
R6790 A1.n32 A1.n31 0.657891
R6791 A1.n49 A1.n48 0.6005
R6792 A1.n30 A1.n29 0.6005
R6793 A1.n52 A1.n51 0.60042
R6794 A1.n49 A1.n39 0.284196
R6795 A1.n48 A1.n44 0.284196
R6796 A1.n29 A1.n21 0.282239
R6797 A1.n30 A1.n10 0.282239
R6798 A1.n52 A1.n34 0.277389
R6799 A1 A1.n53 0.186636
R6800 a_5741_n2271.t8 a_5741_n2271.n19 40.7345
R6801 a_5741_n2271.n24 a_5741_n2271.n5 28.094
R6802 a_5741_n2271.n21 a_5741_n2271.n20 28.094
R6803 a_5741_n2271.n33 a_5741_n2271.n32 28.094
R6804 a_5741_n2271.n27 a_5741_n2271.t16 21.9005
R6805 a_5741_n2271.n27 a_5741_n2271.t24 21.9005
R6806 a_5741_n2271.n0 a_5741_n2271.t20 21.9005
R6807 a_5741_n2271.n11 a_5741_n2271.t18 21.9005
R6808 a_5741_n2271.n12 a_5741_n2271.t29 21.9005
R6809 a_5741_n2271.n1 a_5741_n2271.t10 21.9005
R6810 a_5741_n2271.n28 a_5741_n2271.t17 21.9005
R6811 a_5741_n2271.n28 a_5741_n2271.t28 21.9005
R6812 a_5741_n2271.n29 a_5741_n2271.t9 21.9005
R6813 a_5741_n2271.n29 a_5741_n2271.t21 21.9005
R6814 a_5741_n2271.n2 a_5741_n2271.t14 21.9005
R6815 a_5741_n2271.n13 a_5741_n2271.t12 21.9005
R6816 a_5741_n2271.n14 a_5741_n2271.t23 21.9005
R6817 a_5741_n2271.n3 a_5741_n2271.t26 21.9005
R6818 a_5741_n2271.n30 a_5741_n2271.t11 21.9005
R6819 a_5741_n2271.n30 a_5741_n2271.t22 21.9005
R6820 a_5741_n2271.n31 a_5741_n2271.t25 21.9005
R6821 a_5741_n2271.n31 a_5741_n2271.t15 21.9005
R6822 a_5741_n2271.n4 a_5741_n2271.t7 21.9005
R6823 a_5741_n2271.n15 a_5741_n2271.t27 21.9005
R6824 a_5741_n2271.n20 a_5741_n2271.t8 21.9005
R6825 a_5741_n2271.n5 a_5741_n2271.t13 21.9005
R6826 a_5741_n2271.n32 a_5741_n2271.t19 21.9005
R6827 a_5741_n2271.n32 a_5741_n2271.t6 21.9005
R6828 a_5741_n2271.n20 a_5741_n2271.n15 15.8172
R6829 a_5741_n2271.n5 a_5741_n2271.n4 15.8172
R6830 a_5741_n2271.n4 a_5741_n2271.n3 15.8172
R6831 a_5741_n2271.n15 a_5741_n2271.n14 15.8172
R6832 a_5741_n2271.n14 a_5741_n2271.n13 15.8172
R6833 a_5741_n2271.n3 a_5741_n2271.n2 15.8172
R6834 a_5741_n2271.n2 a_5741_n2271.n1 15.8172
R6835 a_5741_n2271.n13 a_5741_n2271.n12 15.8172
R6836 a_5741_n2271.n12 a_5741_n2271.n11 15.8172
R6837 a_5741_n2271.n1 a_5741_n2271.n0 15.8172
R6838 a_5741_n2271.n28 a_5741_n2271.n27 15.8172
R6839 a_5741_n2271.n30 a_5741_n2271.n29 15.8172
R6840 a_5741_n2271.n29 a_5741_n2271.n28 15.8172
R6841 a_5741_n2271.n32 a_5741_n2271.n31 15.8172
R6842 a_5741_n2271.n31 a_5741_n2271.n30 15.8172
R6843 a_5741_n2271.n17 a_5741_n2271.n16 15.1845
R6844 a_5741_n2271.n19 a_5741_n2271.n18 15.1845
R6845 a_5741_n2271.n18 a_5741_n2271.n17 15.1845
R6846 a_5741_n2271.n8 a_5741_n2271.n6 5.44589
R6847 a_5741_n2271.n8 a_5741_n2271.n7 4.7885
R6848 a_5741_n2271.n34 a_5741_n2271.n33 4.70615
R6849 a_5741_n2271.n23 a_5741_n2271.n22 4.4205
R6850 a_5741_n2271.n26 a_5741_n2271.n25 4.4205
R6851 a_5741_n2271.n10 a_5741_n2271.n9 4.4205
R6852 a_5741_n2271.n10 a_5741_n2271.n8 1.1392
R6853 a_5741_n2271.n26 a_5741_n2271.n24 0.286152
R6854 a_5741_n2271.n23 a_5741_n2271.n21 0.286152
R6855 a_5741_n2271.n33 a_5741_n2271.n26 0.282239
R6856 a_5741_n2271.n21 a_5741_n2271.n10 0.282239
R6857 a_5741_n2271.n24 a_5741_n2271.n23 0.282239
C0 ENA A5 0.493f
C1 TG_magic_0.A S0 0.453f
C2 a_n4701_n4860# VDD 1.27f
C3 TG_magic_7.B Vout 4.92f
C4 TG_magic_7.B VDD 2.21f
C5 a_n2298_n2271# A2 0.00501f
C6 TG_GATE_SWITCH_magic_6.B A4 4.94f
C7 S0 A1 0.0542f
C8 a_n4701_300# TG_GATE_SWITCH_magic_3.B 0.175f
C9 VDD A7 1.95f
C10 TG_magic_7.CLK TG_magic_4.B 0.255f
C11 TG_magic_1.CLK TG_magic_0.A 0.666f
C12 a_n2298_307# TG_GATE_SWITCH_magic_6.B 0.0247f
C13 VDD A4 1.69f
C14 a_n4701_n2278# A2 0.0176f
C15 TG_GATE_SWITCH_magic_0.B a_n2298_n2271# 0.0258f
C16 ENA A6 0.581f
C17 a_n2298_307# VDD 1.27f
C18 S0 A2 0.0527f
C19 TG_magic_7.CLK TG_magic_0.B 0.175f
C20 TG_GATE_SWITCH_magic_0.B a_n4701_n2278# 0.194f
C21 TG_GATE_SWITCH_magic_1.B TG_GATE_SWITCH_magic_5.B 0.462f
C22 TG_GATE_SWITCH_magic_2.B VDD 3.91f
C23 TG_GATE_SWITCH_magic_0.B S0 0.353f
C24 ENA A1 0.772f
C25 TG_GATE_SWITCH_magic_5.B TG_magic_4.B 5.09f
C26 a_n4701_300# VDD 1.27f
C27 TG_magic_2.B Vout 2.99e-19
C28 TG_magic_5.A TG_magic_0.B 5.35f
C29 TG_magic_2.B VDD 1.78f
C30 Vout S2 0.184f
C31 a_n2298_n2271# A0 4.03e-20
C32 TG_GATE_SWITCH_magic_6.B S1 0.0878f
C33 VDD S2 1.4f
C34 TG_magic_7.CLK TG_magic_7.B 0.885f
C35 INVERTER_MUX_1.OUT TG_magic_4.B 0.0122f
C36 TG_magic_1.CLK TG_GATE_SWITCH_magic_0.B 0.343f
C37 TG_GATE_SWITCH_magic_4.B A1 4.98f
C38 S1 Vout 0.00182f
C39 VDD S1 2.52f
C40 a_n2298_n4853# TG_GATE_SWITCH_magic_5.B 0.195f
C41 a_n2298_n2271# a_n2298_n4853# 0.00174f
C42 TG_GATE_SWITCH_magic_1.B S0 0.341f
C43 TG_magic_7.CLK A4 7.7e-20
C44 a_n4701_n2278# A0 0.378f
C45 a_n2298_n7431# VDD 1.27f
C46 ENA A2 1.05f
C47 TG_magic_5.A TG_magic_7.B 0.0014f
C48 INVERTER_MUX_1.OUT a_n2298_n4853# 1.84e-20
C49 TG_magic_4.B S0 0.668f
C50 INVERTER_MUX_1.OUT TG_magic_0.B 0.567f
C51 TG_magic_1.CLK TG_GATE_SWITCH_magic_1.B 0.342f
C52 S0 A0 0.101f
C53 a_n4701_n7438# VDD 1.27f
C54 TG_magic_1.CLK TG_magic_4.B 0.606f
C55 TG_GATE_SWITCH_magic_0.B ENA 0.507f
C56 a_n2298_n4853# S0 5.65e-19
C57 TG_GATE_SWITCH_magic_5.B A7 4.96f
C58 a_n2298_n2271# A7 5.21e-19
C59 TG_magic_0.B S0 0.00263f
C60 INVERTER_MUX_1.OUT TG_magic_7.B 8.56e-19
C61 TG_magic_7.CLK TG_magic_2.B 0.66f
C62 a_n4701_n2278# a_n4701_n4860# 0.00174f
C63 INVERTER_MUX_1.OUT A7 5.31e-20
C64 a_n2298_n2271# A4 0.458f
C65 TG_GATE_SWITCH_magic_1.B ENA 0.526f
C66 TG_magic_1.CLK TG_magic_0.B 0.0897f
C67 a_n4701_n2278# A7 0.00111f
C68 TG_magic_7.CLK S2 0.99f
C69 a_n2298_307# a_n2298_n2271# 0.0482f
C70 ENA A3 0.68f
C71 TG_magic_7.CLK S1 3.94f
C72 a_n4701_n2278# A4 0.0431f
C73 TG_magic_7.B S0 0.0107f
C74 TG_GATE_SWITCH_magic_3.B TG_GATE_SWITCH_magic_6.B 0.206f
C75 S0 A7 0.149f
C76 TG_GATE_SWITCH_magic_1.B TG_GATE_SWITCH_magic_4.B 0.953f
C77 ENA A0 0.703f
C78 TG_magic_4.B TG_GATE_SWITCH_magic_4.B 0.19f
C79 S0 A4 1.34f
C80 TG_GATE_SWITCH_magic_3.B VDD 4.14f
C81 TG_magic_1.CLK TG_magic_7.B 0.0937f
C82 a_n2298_n4853# ENA 0.178f
C83 TG_magic_5.A S1 0.665f
C84 TG_GATE_SWITCH_magic_5.B TG_GATE_SWITCH_magic_2.B 0.204f
C85 a_n2298_307# S0 0.00513f
C86 TG_magic_1.CLK A4 5.39e-22
C87 TG_GATE_SWITCH_magic_5.B S2 0.268f
C88 A5 A1 0.217f
C89 a_n4701_300# a_n4701_n2278# 0.0482f
C90 TG_GATE_SWITCH_magic_5.B S1 0.00476f
C91 INVERTER_MUX_1.OUT S2 0.42f
C92 a_n2298_n2271# S1 0.038f
C93 TG_GATE_SWITCH_magic_7.B TG_magic_0.A 0.175f
C94 a_n4701_n4860# ENA 0.324f
C95 TG_GATE_SWITCH_magic_5.B a_n2298_n7431# 0.0251f
C96 TG_GATE_SWITCH_magic_2.B S0 0.636f
C97 INVERTER_MUX_1.OUT S1 3.07f
C98 ENA A7 0.353f
C99 TG_GATE_SWITCH_magic_6.B VDD 1.83f
C100 TG_magic_2.B S0 0.694f
C101 a_n4701_n2278# S1 0.0382f
C102 S0 S2 0.656f
C103 ENA A4 0.424f
C104 VDD Vout 2.94f
C105 TG_magic_1.CLK TG_GATE_SWITCH_magic_2.B 0.0206f
C106 TG_magic_1.CLK TG_magic_2.B 0.247f
C107 S0 S1 1.02f
C108 a_n2298_307# ENA 0.176f
C109 TG_magic_1.CLK S2 0.754f
C110 TG_GATE_SWITCH_magic_7.B A2 4.98f
C111 a_n2298_n7431# S0 0.00673f
C112 TG_magic_1.CLK S1 0.222f
C113 A6 A2 0.235f
C114 TG_GATE_SWITCH_magic_3.B TG_magic_5.A 5.17f
C115 TG_GATE_SWITCH_magic_7.B TG_GATE_SWITCH_magic_0.B 1.06f
C116 TG_GATE_SWITCH_magic_2.B ENA 0.335f
C117 a_n4701_300# ENA 0.269f
C118 TG_GATE_SWITCH_magic_1.B A5 0.0442f
C119 TG_GATE_SWITCH_magic_0.B A6 0.0424f
C120 ENA S2 0.615f
C121 TG_GATE_SWITCH_magic_6.B TG_magic_7.CLK 3.4e-19
C122 TG_GATE_SWITCH_magic_2.B TG_GATE_SWITCH_magic_4.B 1.08f
C123 TG_magic_2.B TG_GATE_SWITCH_magic_4.B 5.07f
C124 ENA S1 0.0622f
C125 TG_magic_7.CLK Vout 0.00172f
C126 TG_magic_7.CLK VDD 2.05f
C127 TG_GATE_SWITCH_magic_4.B S2 0.00247f
C128 a_n2298_n7431# ENA 0.172f
C129 TG_GATE_SWITCH_magic_3.B INVERTER_MUX_1.OUT 0.00166f
C130 TG_magic_0.A TG_GATE_SWITCH_magic_0.B 5.35f
C131 a_n4701_n7438# ENA 0.294f
C132 a_n2298_n7431# TG_GATE_SWITCH_magic_4.B 0.174f
C133 TG_magic_5.A Vout 2.05e-19
C134 TG_magic_5.A VDD 2.21f
C135 TG_GATE_SWITCH_magic_3.B S0 0.573f
C136 TG_GATE_SWITCH_magic_6.B a_n2298_n2271# 0.198f
C137 TG_GATE_SWITCH_magic_1.B A1 0.241f
C138 a_n4701_n4860# A5 0.00143f
C139 TG_magic_1.CLK TG_GATE_SWITCH_magic_3.B 0.0213f
C140 A3 A1 0.0136f
C141 TG_GATE_SWITCH_magic_5.B VDD 1.62f
C142 TG_GATE_SWITCH_magic_0.B A2 0.273f
C143 a_n2298_n2271# VDD 1.27f
C144 INVERTER_MUX_1.OUT Vout 0.185f
C145 INVERTER_MUX_1.OUT VDD 1.87f
C146 a_n4701_n2278# VDD 1.27f
C147 TG_GATE_SWITCH_magic_6.B S0 0.781f
C148 a_n2298_n4853# A1 0.00381f
C149 TG_magic_0.A TG_magic_0.B 4.99f
C150 S0 Vout 0.00876f
C151 TG_GATE_SWITCH_magic_3.B ENA 0.306f
C152 VDD S0 6.58f
C153 a_n2298_307# TG_GATE_SWITCH_magic_7.B 0.174f
C154 TG_magic_1.CLK TG_GATE_SWITCH_magic_6.B 0.013f
C155 TG_magic_5.A TG_magic_7.CLK 5.14e-19
C156 A2 A0 0.0212f
C157 TG_magic_1.CLK VDD 3.76f
C158 TG_GATE_SWITCH_magic_2.B A5 5.01f
C159 a_n2298_307# A6 4.24e-19
C160 a_n4701_n4860# A1 0.0142f
C161 S2 A5 0.00688f
C162 TG_GATE_SWITCH_magic_0.B A0 4.94f
C163 TG_magic_7.CLK TG_GATE_SWITCH_magic_5.B 2.45e-19
C164 TG_GATE_SWITCH_magic_6.B ENA 0.00116f
C165 TG_magic_7.CLK INVERTER_MUX_1.OUT 0.459f
C166 TG_GATE_SWITCH_magic_1.B A3 4.94f
C167 a_n2298_307# TG_magic_0.A 4.79e-22
C168 TG_GATE_SWITCH_magic_1.B TG_magic_4.B 5.35f
C169 a_n2298_n7431# A5 4.03e-20
C170 a_n4701_300# A6 0.396f
C171 VDD ENA 4.51f
C172 TG_GATE_SWITCH_magic_7.B S1 0.00166f
C173 a_n4701_n7438# A5 0.405f
C174 TG_magic_5.A INVERTER_MUX_1.OUT 0.257f
C175 TG_magic_7.CLK S0 0.0232f
C176 a_n2298_n4853# TG_GATE_SWITCH_magic_1.B 0.024f
C177 TG_GATE_SWITCH_magic_4.B VDD 2.1f
C178 A2 A4 0.014f
C179 a_n2298_n4853# A3 4.24e-19
C180 TG_GATE_SWITCH_magic_2.B A1 0.409f
C181 TG_magic_1.CLK TG_magic_7.CLK 3.25f
C182 TG_GATE_SWITCH_magic_0.B A7 0.00201f
C183 a_n2298_307# A2 0.532f
C184 TG_magic_5.A S0 0.461f
C185 INVERTER_MUX_1.OUT TG_GATE_SWITCH_magic_5.B 0.00322f
C186 S2 A1 0.165f
C187 TG_GATE_SWITCH_magic_0.B A4 0.181f
C188 a_n4701_n2278# a_n2298_n2271# 2.53e-19
C189 TG_magic_0.A S1 0.268f
C190 a_n4701_n4860# TG_GATE_SWITCH_magic_1.B 0.192f
C191 TG_magic_1.CLK TG_magic_5.A 0.235f
C192 a_n2298_307# TG_GATE_SWITCH_magic_0.B 0.0578f
C193 TG_GATE_SWITCH_magic_1.B A7 0.199f
C194 a_n4701_n4860# A3 0.377f
C195 a_n2298_n7431# A1 0.502f
C196 TG_GATE_SWITCH_magic_5.B S0 0.693f
C197 A3 A7 0.305f
C198 a_n2298_n2271# S0 0.046f
C199 TG_magic_4.B TG_magic_7.B 4.98f
C200 a_n4701_300# A2 0.146f
C201 INVERTER_MUX_1.OUT S0 0.0658f
C202 A0 A7 0.00395f
C203 a_n4701_n7438# A1 0.133f
C204 TG_magic_1.CLK TG_GATE_SWITCH_magic_5.B 0.00555f
C205 TG_magic_1.CLK a_n2298_n2271# 1.32e-19
C206 a_n4701_n2278# S0 0.0328f
C207 a_n4701_n4860# a_n2298_n4853# 3.22e-19
C208 a_n4701_300# TG_GATE_SWITCH_magic_0.B 0.017f
C209 A0 A4 0.296f
C210 TG_magic_7.CLK TG_GATE_SWITCH_magic_4.B 0.00166f
C211 a_n2298_n4853# A7 0.481f
C212 TG_magic_1.CLK INVERTER_MUX_1.OUT 0.635f
C213 TG_GATE_SWITCH_magic_3.B TG_GATE_SWITCH_magic_7.B 0.978f
C214 TG_magic_0.B TG_magic_7.B 0.00132f
C215 TG_GATE_SWITCH_magic_0.B S1 0.0864f
C216 TG_GATE_SWITCH_magic_1.B TG_GATE_SWITCH_magic_2.B 0.442f
C217 TG_GATE_SWITCH_magic_3.B A6 5.03f
C218 TG_magic_1.CLK S0 0.755f
C219 TG_GATE_SWITCH_magic_5.B ENA 0.00106f
C220 TG_magic_4.B TG_GATE_SWITCH_magic_2.B 0.104f
C221 a_n2298_n2271# ENA 0.18f
C222 TG_GATE_SWITCH_magic_1.B S2 0.158f
C223 a_n4701_n4860# A7 0.0654f
C224 TG_magic_4.B TG_magic_2.B 0.186f
C225 A3 S2 0.147f
C226 VDD A5 1.53f
C227 a_n4701_300# A0 0.00143f
C228 TG_magic_4.B S2 0.0558f
C229 TG_GATE_SWITCH_magic_1.B S1 0.008f
C230 TG_GATE_SWITCH_magic_3.B TG_magic_0.A 0.111f
C231 TG_GATE_SWITCH_magic_7.B TG_GATE_SWITCH_magic_6.B 0.285f
C232 a_n4701_n2278# ENA 0.359f
C233 TG_GATE_SWITCH_magic_5.B TG_GATE_SWITCH_magic_4.B 0.299f
C234 S1 A3 0.0115f
C235 TG_GATE_SWITCH_magic_1.B a_n2298_n7431# 0.0561f
C236 TG_magic_4.B S1 0.384f
C237 TG_GATE_SWITCH_magic_7.B VDD 2.36f
C238 TG_magic_4.B a_n2298_n7431# 2.4e-22
C239 A0 S1 0.137f
C240 TG_magic_0.B TG_magic_2.B 0.00159f
C241 ENA S0 0.0467f
C242 a_n2298_n4853# S2 0.12f
C243 TG_GATE_SWITCH_magic_1.B a_n4701_n7438# 0.017f
C244 TG_magic_0.B S2 1.13e-19
C245 a_n2298_307# A4 0.0034f
C246 VDD A6 1.53f
C247 a_n4701_n7438# A3 0.00143f
C248 a_n2298_n4853# S1 0.00431f
C249 TG_GATE_SWITCH_magic_4.B S0 0.234f
C250 TG_magic_0.B S1 0.878f
C251 TG_GATE_SWITCH_magic_3.B A2 0.426f
C252 a_n2298_n4853# a_n2298_n7431# 0.0482f
C253 TG_GATE_SWITCH_magic_6.B TG_magic_0.A 5.12f
C254 TG_magic_7.B TG_GATE_SWITCH_magic_2.B 0.001f
C255 TG_magic_7.B TG_magic_2.B 5.36f
C256 TG_magic_1.CLK TG_GATE_SWITCH_magic_4.B 0.419f
C257 a_n4701_n4860# S2 0.1f
C258 TG_magic_0.A VDD 2.23f
C259 TG_magic_7.B S2 0.582f
C260 TG_GATE_SWITCH_magic_3.B TG_GATE_SWITCH_magic_0.B 0.433f
C261 A7 S2 0.257f
C262 VDD A1 1.49f
C263 a_n4701_n4860# S1 0.00367f
C264 TG_magic_7.B S1 0.173f
C265 S1 A7 0.12f
C266 a_n4701_300# a_n2298_307# 3.22e-19
C267 a_n2298_n7431# A7 0.00143f
C268 TG_GATE_SWITCH_magic_6.B A2 0.0365f
C269 A4 S1 0.15f
C270 a_n4701_n4860# a_n4701_n7438# 0.0482f
C271 VDD A2 1.5f
C272 TG_GATE_SWITCH_magic_6.B TG_GATE_SWITCH_magic_0.B 0.465f
C273 TG_GATE_SWITCH_magic_7.B TG_magic_5.A 5.14f
C274 TG_magic_2.B TG_GATE_SWITCH_magic_2.B 5.18f
C275 TG_GATE_SWITCH_magic_2.B S2 0.00485f
C276 TG_GATE_SWITCH_magic_0.B VDD 2.28f
C277 TG_magic_2.B S2 0.245f
C278 TG_GATE_SWITCH_magic_3.B TG_magic_0.B 9.58e-19
C279 TG_magic_0.A TG_magic_7.CLK 0.37f
C280 TG_magic_2.B S1 4.79e-19
C281 a_n2298_n7431# TG_GATE_SWITCH_magic_2.B 0.0575f
C282 S1 S2 0.0964f
C283 TG_GATE_SWITCH_magic_1.B VDD 1.98f
C284 a_n2298_n7431# S2 0.00981f
C285 TG_magic_0.A TG_magic_5.A 0.18f
C286 a_n4701_n7438# TG_GATE_SWITCH_magic_2.B 0.175f
C287 VDD A3 1.5f
C288 TG_magic_4.B VDD 1.77f
C289 VDD A0 1.49f
C290 a_n4701_n7438# S2 0.00948f
C291 a_n4701_n2278# A6 0.00143f
C292 TG_GATE_SWITCH_magic_7.B S0 0.156f
C293 a_n2298_n4853# VDD 1.27f
C294 TG_GATE_SWITCH_magic_5.B A1 0.039f
C295 TG_magic_0.B Vout 4.92f
C296 a_n2298_307# TG_GATE_SWITCH_magic_3.B 0.0563f
C297 TG_magic_1.CLK TG_GATE_SWITCH_magic_7.B 0.363f
C298 a_n4701_n7438# a_n2298_n7431# 2.53e-19
C299 TG_magic_0.B VDD 2.38f
C300 TG_GATE_SWITCH_magic_0.B TG_magic_7.CLK 0.00166f
C301 TG_magic_0.A INVERTER_MUX_1.OUT 0.0649f
.ends

