magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -3754 -2190 3754 2190
<< nwell >>
rect -1754 -190 1754 190
<< pmos >>
rect -1580 -60 -1480 60
rect -1376 -60 -1276 60
rect -1172 -60 -1072 60
rect -968 -60 -868 60
rect -764 -60 -664 60
rect -560 -60 -460 60
rect -356 -60 -256 60
rect -152 -60 -52 60
rect 52 -60 152 60
rect 256 -60 356 60
rect 460 -60 560 60
rect 664 -60 764 60
rect 868 -60 968 60
rect 1072 -60 1172 60
rect 1276 -60 1376 60
rect 1480 -60 1580 60
<< pdiff >>
rect -1668 23 -1580 60
rect -1668 -23 -1655 23
rect -1609 -23 -1580 23
rect -1668 -60 -1580 -23
rect -1480 23 -1376 60
rect -1480 -23 -1451 23
rect -1405 -23 -1376 23
rect -1480 -60 -1376 -23
rect -1276 23 -1172 60
rect -1276 -23 -1247 23
rect -1201 -23 -1172 23
rect -1276 -60 -1172 -23
rect -1072 23 -968 60
rect -1072 -23 -1043 23
rect -997 -23 -968 23
rect -1072 -60 -968 -23
rect -868 23 -764 60
rect -868 -23 -839 23
rect -793 -23 -764 23
rect -868 -60 -764 -23
rect -664 23 -560 60
rect -664 -23 -635 23
rect -589 -23 -560 23
rect -664 -60 -560 -23
rect -460 23 -356 60
rect -460 -23 -431 23
rect -385 -23 -356 23
rect -460 -60 -356 -23
rect -256 23 -152 60
rect -256 -23 -227 23
rect -181 -23 -152 23
rect -256 -60 -152 -23
rect -52 23 52 60
rect -52 -23 -23 23
rect 23 -23 52 23
rect -52 -60 52 -23
rect 152 23 256 60
rect 152 -23 181 23
rect 227 -23 256 23
rect 152 -60 256 -23
rect 356 23 460 60
rect 356 -23 385 23
rect 431 -23 460 23
rect 356 -60 460 -23
rect 560 23 664 60
rect 560 -23 589 23
rect 635 -23 664 23
rect 560 -60 664 -23
rect 764 23 868 60
rect 764 -23 793 23
rect 839 -23 868 23
rect 764 -60 868 -23
rect 968 23 1072 60
rect 968 -23 997 23
rect 1043 -23 1072 23
rect 968 -60 1072 -23
rect 1172 23 1276 60
rect 1172 -23 1201 23
rect 1247 -23 1276 23
rect 1172 -60 1276 -23
rect 1376 23 1480 60
rect 1376 -23 1405 23
rect 1451 -23 1480 23
rect 1376 -60 1480 -23
rect 1580 23 1668 60
rect 1580 -23 1609 23
rect 1655 -23 1668 23
rect 1580 -60 1668 -23
<< pdiffc >>
rect -1655 -23 -1609 23
rect -1451 -23 -1405 23
rect -1247 -23 -1201 23
rect -1043 -23 -997 23
rect -839 -23 -793 23
rect -635 -23 -589 23
rect -431 -23 -385 23
rect -227 -23 -181 23
rect -23 -23 23 23
rect 181 -23 227 23
rect 385 -23 431 23
rect 589 -23 635 23
rect 793 -23 839 23
rect 997 -23 1043 23
rect 1201 -23 1247 23
rect 1405 -23 1451 23
rect 1609 -23 1655 23
<< polysilicon >>
rect -1580 60 -1480 104
rect -1376 60 -1276 104
rect -1172 60 -1072 104
rect -968 60 -868 104
rect -764 60 -664 104
rect -560 60 -460 104
rect -356 60 -256 104
rect -152 60 -52 104
rect 52 60 152 104
rect 256 60 356 104
rect 460 60 560 104
rect 664 60 764 104
rect 868 60 968 104
rect 1072 60 1172 104
rect 1276 60 1376 104
rect 1480 60 1580 104
rect -1580 -104 -1480 -60
rect -1376 -104 -1276 -60
rect -1172 -104 -1072 -60
rect -968 -104 -868 -60
rect -764 -104 -664 -60
rect -560 -104 -460 -60
rect -356 -104 -256 -60
rect -152 -104 -52 -60
rect 52 -104 152 -60
rect 256 -104 356 -60
rect 460 -104 560 -60
rect 664 -104 764 -60
rect 868 -104 968 -60
rect 1072 -104 1172 -60
rect 1276 -104 1376 -60
rect 1480 -104 1580 -60
<< metal1 >>
rect -1655 23 -1609 58
rect -1655 -58 -1609 -23
rect -1451 23 -1405 58
rect -1451 -58 -1405 -23
rect -1247 23 -1201 58
rect -1247 -58 -1201 -23
rect -1043 23 -997 58
rect -1043 -58 -997 -23
rect -839 23 -793 58
rect -839 -58 -793 -23
rect -635 23 -589 58
rect -635 -58 -589 -23
rect -431 23 -385 58
rect -431 -58 -385 -23
rect -227 23 -181 58
rect -227 -58 -181 -23
rect -23 23 23 58
rect -23 -58 23 -23
rect 181 23 227 58
rect 181 -58 227 -23
rect 385 23 431 58
rect 385 -58 431 -23
rect 589 23 635 58
rect 589 -58 635 -23
rect 793 23 839 58
rect 793 -58 839 -23
rect 997 23 1043 58
rect 997 -58 1043 -23
rect 1201 23 1247 58
rect 1201 -58 1247 -23
rect 1405 23 1451 58
rect 1405 -58 1451 -23
rect 1609 23 1655 58
rect 1609 -58 1655 -23
<< end >>
