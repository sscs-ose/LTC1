* NGSPICE file created from mux_8x1_ibr_flat.ext - technology: gf180mcuC

.subckt pex_mux_8x1_ibr VDD VSS S1 S0 OUT S2 I0 I7 I3 I2 I5 I1 I4 I6
X0 mux_4x1_ibr_0.mux_2x1_ibr_2.I1 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 VDD.t42 VDD.t41 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1 mux_2x1_ibr_0.nand2_ibr_1.IN2 S2.t0 a_3615_1307# VSS.t29 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2 VDD mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_4x1_ibr_0.mux_2x1_ibr_2.I1 VDD.t110 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 S1.t0 a_2490_n1395# VSS.t23 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X4 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 S1.t1 VDD.t31 VDD.t30 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X5 VDD mux_2x1_ibr_0.I0 mux_2x1_ibr_0.nand2_ibr_2.OUT VDD.t88 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X6 mux_2x1_ibr_0.nand2_ibr_1.IN2 mux_2x1_ibr_0.I1 VDD.t50 VDD.t49 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X7 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 VDD.t87 VDD.t86 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X8 mux_2x1_ibr_0.nand2_ibr_2.OUT mux_2x1_ibr_0.I0 a_4178_707# VSS.t11 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X9 a_1927_707# mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 VSS.t48 VSS.t33 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X10 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 S0.t0 VDD.t37 VDD.t36 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X11 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 VDD.t1 VDD.t0 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X12 VDD S1.t2 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 VDD.t32 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X13 a_3053_707# mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 VSS.t1 VSS.t0 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X14 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 VDD.t43 VDD.t0 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X15 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 S0.t1 a_238_n1395# VSS.t30 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X16 a_1927_n1395# mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 VSS.t6 VSS.t5 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X17 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 VDD.t29 VDD.t28 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X18 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 S0.t2 VDD.t70 VDD.t69 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X19 VDD mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT VDD.t81 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X20 VDD I4.t0 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT VDD.t64 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X21 a_1927_1307# mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 VSS.t34 VSS.t33 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X22 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT I4.t1 a_801_707# VSS.t36 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X23 VDD S0.t3 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 VDD.t71 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X24 a_1364_n1395# I3.t0 VSS.t62 VSS.t61 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X25 mux_4x1_ibr_1.mux_2x1_ibr_2.I1 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 VDD.t7 VDD.t6 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X26 mux_4x1_ibr_0.mux_2x1_ibr_2.I1 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT a_1927_1307# VSS.t42 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X27 VDD S1.t3 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 VDD.t94 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X28 VDD I6.t0 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT VDD.t38 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X29 VDD mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_4x1_ibr_0.mux_2x1_ibr_2.I0 VDD.t44 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X30 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 S0.t4 VDD.t75 VDD.t74 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X31 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT I6.t1 a_1927_707# VSS.t42 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X32 VDD mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT VDD.t81 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X33 VDD S0.t5 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 VDD.t51 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X34 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT mux_4x1_ibr_0.mux_2x1_ibr_2.I0 a_3053_707# VSS.t21 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X35 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 mux_4x1_ibr_0.mux_2x1_ibr_2.I1 VDD.t9 VDD.t8 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X36 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 I3.t1 VDD.t109 VDD.t108 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X37 a_3615_1307# mux_2x1_ibr_0.I1 VSS.t38 VSS.t37 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X38 a_1927_n795# mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 VSS.t56 VSS.t5 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X39 a_238_n1395# I1.t0 VSS.t32 VSS.t31 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X40 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT I2.t0 a_1927_n795# VSS.t26 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X41 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 S1.t4 VSS.t50 VSS.t49 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X42 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 I1.t1 VDD.t60 VDD.t59 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X43 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 S0.t6 VSS.t40 VSS.t39 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X44 mux_2x1_ibr_0.I0 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT a_3053_n1395# VSS.t45 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X45 VDD S0.t7 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 VDD.t54 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X46 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 S0.t8 VSS.t59 VSS.t58 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X47 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 S1.t5 a_2490_1307# VSS.t51 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X48 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT a_801_1307# VSS.t36 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X49 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 I7.t0 VDD.t100 VDD.t99 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X50 mux_2x1_ibr_0.I1 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 VDD.t3 VDD.t2 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X51 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 S1.t6 VDD.t85 VDD.t84 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X52 a_2490_1307# mux_4x1_ibr_0.mux_2x1_ibr_2.I1 VSS.t8 VSS.t7 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X53 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 S0.t9 a_238_1307# VSS.t60 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X54 VDD mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT mux_2x1_ibr_0.I0 VDD.t78 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X55 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 S0.t10 VDD.t107 VDD.t106 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X56 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 VDD.t105 VDD.t104 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X57 VDD mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT mux_2x1_ibr_0.I1 VDD.t25 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X58 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 I5.t0 VDD.t19 VDD.t18 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X59 a_2490_n1395# mux_4x1_ibr_1.mux_2x1_ibr_2.I1 VSS.t55 VSS.t54 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X60 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 S0.t11 VSS.t15 VSS.t14 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X61 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 VDD.t103 VDD.t86 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X62 mux_2x1_ibr_0.nand2_ibr_2.IN2 S2.t1 VDD.t48 VDD.t47 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X63 VDD mux_2x1_ibr_0.nand2_ibr_2.OUT OUT.t0 VDD.t15 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X64 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT I0.t0 a_801_n795# VSS.t20 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X65 OUT mux_2x1_ibr_0.nand2_ibr_1.IN2 VDD.t58 VDD.t57 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X66 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 mux_4x1_ibr_1.mux_2x1_ibr_2.I1 VDD.t102 VDD.t101 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X67 VDD I2.t1 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT VDD.t38 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X68 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 S0.t12 a_1364_1307# VSS.t16 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X69 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 S0.t13 a_1364_n1395# VSS.t17 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X70 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT a_801_n1395# VSS.t20 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X71 a_1364_1307# I7.t1 VSS.t53 VSS.t52 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X72 a_3053_1307# mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 VSS.t2 VSS.t0 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X73 VDD S0.t14 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 VDD.t61 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X74 VDD mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_4x1_ibr_1.mux_2x1_ibr_2.I0 VDD.t22 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X75 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 VDD.t35 VDD.t28 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X76 a_801_1307# mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 VSS.t57 VSS.t24 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X77 a_3053_n1395# mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 VSS.t4 VSS.t3 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X78 a_801_707# mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 VSS.t25 VSS.t24 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X79 mux_2x1_ibr_0.I1 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT a_3053_1307# VSS.t21 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X80 VDD S2.t2 mux_2x1_ibr_0.nand2_ibr_1.IN2 VDD.t10 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X81 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 S1.t7 VSS.t47 VSS.t46 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X82 a_238_1307# I5.t1 VSS.t13 VSS.t12 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X83 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 S0.t15 VSS.t44 VSS.t43 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X84 OUT mux_2x1_ibr_0.nand2_ibr_2.OUT a_4178_1307# VSS.t11 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X85 mux_2x1_ibr_0.I0 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 VDD.t5 VDD.t4 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X86 mux_4x1_ibr_1.mux_2x1_ibr_2.I1 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT a_1927_n1395# VSS.t26 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X87 a_3053_n795# mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 VSS.t35 VSS.t3 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X88 a_4178_1307# mux_2x1_ibr_0.nand2_ibr_1.IN2 VSS.t41 VSS.t18 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X89 VDD I0.t1 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT VDD.t64 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X90 mux_2x1_ibr_0.nand2_ibr_2.IN2 S2.t3 VSS.t28 VSS.t27 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X91 a_801_n1395# mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 VSS.t10 VSS.t9 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X92 a_801_n795# mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 VSS.t22 VSS.t9 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X93 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT mux_4x1_ibr_1.mux_2x1_ibr_2.I0 a_3053_n795# VSS.t45 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X94 mux_2x1_ibr_0.nand2_ibr_2.OUT mux_2x1_ibr_0.nand2_ibr_2.IN2 VDD.t21 VDD.t20 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X95 VDD mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_4x1_ibr_1.mux_2x1_ibr_2.I1 VDD.t91 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X96 a_4178_707# mux_2x1_ibr_0.nand2_ibr_2.IN2 VSS.t19 VSS.t18 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X97 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 VDD.t14 VDD.t13 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
R0 VDD.t57 VDD.t10 763.259
R1 VDD.t2 VDD.t94 763.259
R2 VDD.t110 VDD.t8 763.259
R3 VDD.t41 VDD.t54 763.259
R4 VDD.t44 VDD.t99 763.259
R5 VDD.t51 VDD.t104 763.259
R6 VDD.t4 VDD.t32 763.259
R7 VDD.t91 VDD.t101 763.259
R8 VDD.t61 VDD.t6 763.259
R9 VDD.t22 VDD.t108 763.259
R10 VDD.t71 VDD.t13 763.259
R11 VDD.t25 VDD.t49 761.365
R12 VDD.n53 VDD.t20 386.348
R13 VDD.n67 VDD.t84 365.673
R14 VDD.n117 VDD.t69 365.673
R15 VDD.n38 VDD.t106 365.673
R16 VDD.n53 VDD.t47 362.409
R17 VDD.n68 VDD.t30 360.012
R18 VDD.n115 VDD.t36 360.012
R19 VDD.n37 VDD.t74 360.012
R20 VDD.n117 VDD.n116 322.221
R21 VDD.n74 VDD.n53 319.75
R22 VDD.n67 VDD.n66 319.733
R23 VDD.n118 VDD.n117 319.733
R24 VDD.n39 VDD.n38 319.733
R25 VDD.n79 VDD.t15 193.183
R26 VDD.n87 VDD.t10 193.183
R27 VDD.n88 VDD.t25 193.183
R28 VDD.n96 VDD.t94 193.183
R29 VDD.n97 VDD.t110 193.183
R30 VDD.n106 VDD.t54 193.183
R31 VDD.n107 VDD.t44 193.183
R32 VDD.n108 VDD.t51 193.183
R33 VDD.n52 VDD.t88 193.183
R34 VDD.n6 VDD.t78 193.183
R35 VDD.n16 VDD.t32 193.183
R36 VDD.n17 VDD.t91 193.183
R37 VDD.n18 VDD.t61 193.183
R38 VDD.n20 VDD.t22 193.183
R39 VDD.n24 VDD.t71 193.183
R40 VDD.t0 VDD.n69 192.236
R41 VDD.n114 VDD.t28 192.236
R42 VDD.n36 VDD.t86 192.236
R43 VDD.n79 VDD.t57 109.849
R44 VDD.t49 VDD.n87 109.849
R45 VDD.n88 VDD.t2 109.849
R46 VDD.t8 VDD.n96 109.849
R47 VDD.n97 VDD.t41 109.849
R48 VDD.t99 VDD.n106 109.849
R49 VDD.t104 VDD.n107 109.849
R50 VDD.n108 VDD.t18 109.849
R51 VDD.t20 VDD.n52 109.849
R52 VDD.n6 VDD.t4 109.849
R53 VDD.t101 VDD.n16 109.849
R54 VDD.t6 VDD.n17 109.849
R55 VDD.t108 VDD.n18 109.849
R56 VDD.t13 VDD.n20 109.849
R57 VDD.n24 VDD.t59 109.849
R58 VDD.n70 VDD.t81 96.5914
R59 VDD.n43 VDD.t64 96.5914
R60 VDD.n0 VDD.t38 96.5914
R61 VDD.n70 VDD.t0 54.9247
R62 VDD.t28 VDD.n43 54.9247
R63 VDD.t86 VDD.n0 54.9247
R64 VDD.n58 VDD 18.0631
R65 VDD.n75 VDD 11.7877
R66 VDD.n25 VDD.n24 6.3005
R67 VDD.n28 VDD.n20 6.3005
R68 VDD.n31 VDD.n18 6.3005
R69 VDD.n17 VDD.n2 6.3005
R70 VDD.n16 VDD.n15 6.3005
R71 VDD.n7 VDD.n6 6.3005
R72 VDD.n52 VDD.n51 6.3005
R73 VDD.n80 VDD.n79 6.3005
R74 VDD.n87 VDD.n86 6.3005
R75 VDD.n89 VDD.n88 6.3005
R76 VDD.n96 VDD.n95 6.3005
R77 VDD.n98 VDD.n97 6.3005
R78 VDD.n106 VDD.n105 6.3005
R79 VDD.n107 VDD.n44 6.3005
R80 VDD.n109 VDD.n108 6.3005
R81 VDD VDD.n5 5.23855
R82 VDD VDD.n50 5.23855
R83 VDD VDD.n78 5.23855
R84 VDD.n109 VDD.t19 5.21701
R85 VDD.n25 VDD.t60 5.21701
R86 VDD.n118 VDD.t70 5.19258
R87 VDD.n116 VDD.t37 5.19258
R88 VDD.n73 VDD.t48 5.1858
R89 VDD.n65 VDD.t85 5.14703
R90 VDD.n60 VDD.t31 5.14703
R91 VDD.n124 VDD.t75 5.14703
R92 VDD.n40 VDD.t107 5.14703
R93 VDD.n104 VDD.t100 5.13746
R94 VDD.n94 VDD.t9 5.13746
R95 VDD.n85 VDD.t50 5.13746
R96 VDD.n14 VDD.t102 5.13746
R97 VDD.n30 VDD.t109 5.13746
R98 VDD.n63 VDD.n61 5.13287
R99 VDD.n63 VDD.n62 5.13287
R100 VDD.n110 VDD.n45 5.13287
R101 VDD.n103 VDD.n102 5.13287
R102 VDD.n101 VDD.n46 5.13287
R103 VDD.n93 VDD.n92 5.13287
R104 VDD.n91 VDD.n47 5.13287
R105 VDD.n84 VDD.n83 5.13287
R106 VDD.n82 VDD.n49 5.13287
R107 VDD.n72 VDD.n54 5.13287
R108 VDD.n72 VDD.n55 5.13287
R109 VDD.n11 VDD.n4 5.13287
R110 VDD.n13 VDD.n12 5.13287
R111 VDD.n32 VDD.n3 5.13287
R112 VDD.n29 VDD.n19 5.13287
R113 VDD.n122 VDD.n41 5.13287
R114 VDD.n122 VDD.n42 5.13287
R115 VDD.n26 VDD.n23 5.13287
R116 VDD.n112 VDD.t105 3.91303
R117 VDD.n48 VDD.t3 3.91303
R118 VDD.n99 VDD.t42 3.91303
R119 VDD.n77 VDD.t58 3.91303
R120 VDD.n34 VDD.t7 3.9128
R121 VDD.n22 VDD.t14 3.9128
R122 VDD.n9 VDD.t5 3.91277
R123 VDD.n9 VDD.n8 3.87701
R124 VDD.n22 VDD.n21 3.87649
R125 VDD.n113 VDD.n112 3.87623
R126 VDD.n56 VDD.n48 3.87623
R127 VDD.n99 VDD.n1 3.87623
R128 VDD.n35 VDD.n34 3.87585
R129 VDD.n77 VDD.n76 3.87523
R130 VDD.n1 VDD.t87 3.51093
R131 VDD.n76 VDD.t21 3.51093
R132 VDD.n113 VDD.t35 3.51093
R133 VDD.n56 VDD.t1 3.51093
R134 VDD.n21 VDD.t29 3.51079
R135 VDD.n8 VDD.t43 3.51063
R136 VDD.n35 VDD.t103 3.51063
R137 VDD.n73 VDD.n72 3.45802
R138 VDD.n71 VDD.n70 3.15287
R139 VDD.n121 VDD.n43 3.1505
R140 VDD.n128 VDD.n0 3.1505
R141 VDD.n69 VDD.n68 0.939698
R142 VDD.n115 VDD.n114 0.939698
R143 VDD.n37 VDD.n36 0.939698
R144 VDD.n119 VDD 0.412255
R145 VDD.n126 VDD 0.412255
R146 VDD.n126 VDD 0.412255
R147 VDD VDD.n58 0.411896
R148 VDD.n119 VDD 0.411255
R149 VDD.n127 VDD.n35 0.273886
R150 VDD.n120 VDD.n113 0.272927
R151 VDD.n57 VDD.n56 0.272927
R152 VDD.n76 VDD.n75 0.272927
R153 VDD.n127 VDD.n1 0.272927
R154 VDD.n112 VDD.n111 0.22389
R155 VDD.n90 VDD.n48 0.22389
R156 VDD.n81 VDD.n77 0.22389
R157 VDD.n100 VDD.n99 0.22389
R158 VDD.n34 VDD.n33 0.22353
R159 VDD.n27 VDD.n22 0.22353
R160 VDD.n10 VDD.n9 0.223424
R161 VDD.n65 VDD.n64 0.176707
R162 VDD.n64 VDD.n60 0.143461
R163 VDD.n14 VDD.n13 0.141016
R164 VDD.n30 VDD.n29 0.141016
R165 VDD.n94 VDD.n93 0.141016
R166 VDD.n104 VDD.n103 0.141016
R167 VDD.n85 VDD.n84 0.140435
R168 VDD.n123 VDD.n40 0.139013
R169 VDD.n124 VDD.n123 0.139013
R170 VDD VDD.n11 0.106177
R171 VDD.n13 VDD 0.106177
R172 VDD.n32 VDD 0.106177
R173 VDD.n29 VDD 0.106177
R174 VDD.n26 VDD 0.106177
R175 VDD VDD.n82 0.106177
R176 VDD.n84 VDD 0.106177
R177 VDD VDD.n91 0.106177
R178 VDD.n93 VDD 0.106177
R179 VDD VDD.n101 0.106177
R180 VDD.n103 VDD 0.106177
R181 VDD.n110 VDD 0.106177
R182 VDD.n10 VDD.n7 0.0800484
R183 VDD.n15 VDD.n14 0.0800484
R184 VDD.n33 VDD.n2 0.0800484
R185 VDD.n28 VDD.n27 0.0800484
R186 VDD.n75 VDD.n51 0.0800484
R187 VDD.n81 VDD.n80 0.0800484
R188 VDD.n86 VDD.n85 0.0800484
R189 VDD.n90 VDD.n89 0.0800484
R190 VDD.n95 VDD.n94 0.0800484
R191 VDD.n100 VDD.n98 0.0800484
R192 VDD.n111 VDD.n44 0.0800484
R193 VDD VDD.n30 0.0788871
R194 VDD VDD.n104 0.0788871
R195 VDD VDD.n10 0.0713387
R196 VDD.n33 VDD 0.0713387
R197 VDD.n27 VDD 0.0713387
R198 VDD VDD.n81 0.0713387
R199 VDD VDD.n90 0.0713387
R200 VDD VDD.n100 0.0713387
R201 VDD.n111 VDD 0.0713387
R202 VDD.n11 VDD 0.0701774
R203 VDD VDD.n32 0.0701774
R204 VDD VDD.n26 0.0701774
R205 VDD.n82 VDD 0.0701774
R206 VDD.n91 VDD 0.0701774
R207 VDD.n101 VDD 0.0701774
R208 VDD VDD.n110 0.0701774
R209 VDD.n122 VDD 0.0533387
R210 VDD.n72 VDD 0.0533387
R211 VDD.n63 VDD 0.0513065
R212 VDD.n66 VDD.n65 0.0460556
R213 VDD.n60 VDD.n59 0.0460556
R214 VDD.n40 VDD.n39 0.0460556
R215 VDD.n125 VDD.n124 0.0460556
R216 VDD.n121 VDD.n120 0.0402742
R217 VDD.n71 VDD.n57 0.0402742
R218 VDD.n128 VDD.n127 0.0402742
R219 VDD.n123 VDD.n122 0.0338871
R220 VDD.n64 VDD.n63 0.0318548
R221 VDD.n58 VDD.n57 0.0239437
R222 VDD.n120 VDD.n119 0.0225645
R223 VDD.n127 VDD.n126 0.0225645
R224 VDD.n68 VDD.n67 0.00925055
R225 VDD.n117 VDD.n115 0.00925055
R226 VDD.n38 VDD.n37 0.00925055
R227 VDD.n74 VDD.n73 0.00883333
R228 VDD.n7 VDD 0.00166129
R229 VDD.n15 VDD 0.00166129
R230 VDD VDD.n2 0.00166129
R231 VDD VDD.n31 0.00166129
R232 VDD.n31 VDD 0.00166129
R233 VDD VDD.n28 0.00166129
R234 VDD VDD.n25 0.00166129
R235 VDD.n51 VDD 0.00166129
R236 VDD.n80 VDD 0.00166129
R237 VDD.n86 VDD 0.00166129
R238 VDD.n89 VDD 0.00166129
R239 VDD.n95 VDD 0.00166129
R240 VDD.n98 VDD 0.00166129
R241 VDD.n105 VDD 0.00166129
R242 VDD.n105 VDD 0.00166129
R243 VDD VDD.n44 0.00166129
R244 VDD VDD.n109 0.00166129
R245 VDD VDD.n121 0.00108064
R246 VDD VDD.n71 0.00108064
R247 VDD VDD.n128 0.00108064
R248 VDD.n66 VDD 0.00105556
R249 VDD.n59 VDD 0.00105556
R250 VDD.n116 VDD 0.00105556
R251 VDD VDD.n118 0.00105556
R252 VDD.n39 VDD 0.00105556
R253 VDD VDD.n125 0.00105556
R254 VDD VDD.n74 0.00105556
R255 S2.n1 S2.t0 31.528
R256 S2.n0 S2.t1 25.7638
R257 S2.n1 S2.t2 15.3826
R258 S2.n0 S2.t3 13.2969
R259 S2.n2 S2.n1 7.62851
R260 S2.n5 S2 2.26613
R261 S2.n6 S2.n4 2.2505
R262 S2.n3 S2.n2 2.2324
R263 S2.n6 S2.n0 2.11815
R264 S2.n2 S2 0.107918
R265 S2.n4 S2.n3 0.0289694
R266 S2.n6 S2.n5 0.00563331
R267 S2 S2.n4 0.00233673
R268 S2.n5 S2 0.00193332
R269 S2 S2.n6 0.00142783
R270 VSS.n37 VSS.n36 28802.9
R271 VSS.t12 VSS.t31 23952.8
R272 VSS.t45 VSS.n25 21804.7
R273 VSS.t54 VSS.t26 1483.3
R274 VSS.t5 VSS.t17 1483.3
R275 VSS.t61 VSS.t20 1483.3
R276 VSS.t9 VSS.t30 1483.3
R277 VSS.t29 VSS.t18 1483.3
R278 VSS.t0 VSS.t51 1483.3
R279 VSS.t52 VSS.t36 1483.3
R280 VSS.t60 VSS.t24 1483.3
R281 VSS.t37 VSS.t21 1479.61
R282 VSS.t23 VSS.t3 1367.44
R283 VSS.n12 VSS.t11 353.341
R284 VSS.n36 VSS.n35 349.661
R285 VSS.n58 VSS.n57 349.661
R286 VSS.n38 VSS.n37 349.661
R287 VSS.n47 VSS.n6 349.661
R288 VSS.n25 VSS.n24 345.981
R289 VSS.n27 VSS.t45 298.279
R290 VSS.n29 VSS.t54 235.561
R291 VSS.n35 VSS.t5 235.561
R292 VSS.n59 VSS.t61 235.561
R293 VSS.n57 VSS.t9 235.561
R294 VSS.t31 VSS.n49 235.561
R295 VSS.t18 VSS.n12 235.561
R296 VSS.n14 VSS.t37 235.561
R297 VSS.n24 VSS.t0 235.561
R298 VSS.n17 VSS.t7 235.561
R299 VSS.n38 VSS.t33 235.561
R300 VSS.n43 VSS.t52 235.561
R301 VSS.t24 VSS.n47 235.561
R302 VSS.n50 VSS.t12 235.561
R303 VSS.t3 VSS.n27 198.853
R304 VSS.n54 VSS.t40 9.34566
R305 VSS.n9 VSS.t28 9.34566
R306 VSS.n21 VSS.t47 9.34566
R307 VSS.n40 VSS.t44 9.34566
R308 VSS.n4 VSS.t59 9.34566
R309 VSS.n7 VSS.t50 9.34566
R310 VSS.n32 VSS.t15 9.34566
R311 VSS.n25 VSS.t21 7.36177
R312 VSS.n3 VSS.t22 7.19156
R313 VSS.n3 VSS.t10 7.19156
R314 VSS.n11 VSS.t41 7.19156
R315 VSS.n11 VSS.t19 7.19156
R316 VSS.n16 VSS.t38 7.19156
R317 VSS.n19 VSS.t2 7.19156
R318 VSS.n19 VSS.t1 7.19156
R319 VSS.n20 VSS.t8 7.19156
R320 VSS.n39 VSS.t34 7.19156
R321 VSS.n39 VSS.t48 7.19156
R322 VSS.n45 VSS.t53 7.19156
R323 VSS.n46 VSS.t57 7.19156
R324 VSS.n46 VSS.t25 7.19156
R325 VSS.n52 VSS.t13 7.19156
R326 VSS.n53 VSS.t32 7.19156
R327 VSS.n26 VSS.t35 7.19156
R328 VSS.n26 VSS.t4 7.19156
R329 VSS.n31 VSS.t55 7.19156
R330 VSS.n34 VSS.t56 7.19156
R331 VSS.n34 VSS.t6 7.19156
R332 VSS.n0 VSS.t62 7.19156
R333 VSS.t49 VSS.t23 3.68113
R334 VSS.n36 VSS.t26 3.68113
R335 VSS.t17 VSS.t14 3.68113
R336 VSS.t20 VSS.n58 3.68113
R337 VSS.t30 VSS.t39 3.68113
R338 VSS.t27 VSS.t29 3.68113
R339 VSS.t51 VSS.t46 3.68113
R340 VSS.n37 VSS.t42 3.68113
R341 VSS.t43 VSS.t16 3.68113
R342 VSS.t36 VSS.n6 3.68113
R343 VSS.t58 VSS.t60 3.68113
R344 VSS.n60 VSS.n1 3.37613
R345 VSS.n30 VSS.n28 3.37613
R346 VSS.n15 VSS.n13 3.37613
R347 VSS.n23 VSS.n18 3.37613
R348 VSS.n44 VSS.n42 3.37613
R349 VSS.n51 VSS.n48 3.37613
R350 VSS.n56 VSS.n2 3.37613
R351 VSS.n57 VSS 2.6035
R352 VSS.n47 VSS 2.6035
R353 VSS VSS.n38 2.6035
R354 VSS.n24 VSS 2.6035
R355 VSS.n12 VSS 2.6035
R356 VSS.n35 VSS 2.6035
R357 VSS.n27 VSS 2.60269
R358 VSS.n56 VSS.n55 2.6005
R359 VSS.t39 VSS.n56 2.6005
R360 VSS VSS.n2 2.6005
R361 VSS.n49 VSS.n2 2.6005
R362 VSS VSS.n51 2.6005
R363 VSS.n51 VSS.n50 2.6005
R364 VSS VSS.n44 2.6005
R365 VSS.n44 VSS.n43 2.6005
R366 VSS VSS.n18 2.6005
R367 VSS.n18 VSS.n17 2.6005
R368 VSS VSS.n15 2.6005
R369 VSS.n15 VSS.n14 2.6005
R370 VSS.n13 VSS.n10 2.6005
R371 VSS.n13 VSS.t27 2.6005
R372 VSS.n23 VSS.n22 2.6005
R373 VSS.t46 VSS.n23 2.6005
R374 VSS.n42 VSS.n41 2.6005
R375 VSS.n42 VSS.t43 2.6005
R376 VSS.n48 VSS.n5 2.6005
R377 VSS.n48 VSS.t58 2.6005
R378 VSS.n28 VSS.n8 2.6005
R379 VSS.n28 VSS.t49 2.6005
R380 VSS VSS.n30 2.6005
R381 VSS.n30 VSS.n29 2.6005
R382 VSS.n33 VSS.n1 2.6005
R383 VSS.t14 VSS.n1 2.6005
R384 VSS VSS.n60 2.6005
R385 VSS.n60 VSS.n59 2.6005
R386 VSS.n55 VSS.n3 0.131017
R387 VSS.n11 VSS.n10 0.131017
R388 VSS.n22 VSS.n19 0.131017
R389 VSS.n41 VSS.n39 0.131017
R390 VSS.n46 VSS.n5 0.131017
R391 VSS.n26 VSS.n8 0.131017
R392 VSS.n34 VSS.n33 0.131017
R393 VSS.n3 VSS 0.0595367
R394 VSS VSS.n11 0.0595367
R395 VSS.n19 VSS 0.0595367
R396 VSS.n39 VSS 0.0595367
R397 VSS VSS.n46 0.0595367
R398 VSS VSS.n26 0.0595367
R399 VSS VSS.n34 0.0595367
R400 VSS.n16 VSS 0.0569474
R401 VSS VSS.n20 0.0569474
R402 VSS.n45 VSS 0.0569474
R403 VSS.n52 VSS 0.0569474
R404 VSS VSS.n53 0.0569474
R405 VSS.n31 VSS 0.0569474
R406 VSS VSS.n0 0.0569474
R407 VSS VSS.n9 0.0340526
R408 VSS VSS.n21 0.0340526
R409 VSS VSS.n40 0.0340526
R410 VSS VSS.n4 0.0340526
R411 VSS VSS.n54 0.0340526
R412 VSS VSS.n7 0.0340526
R413 VSS VSS.n32 0.0320789
R414 VSS VSS.n16 0.0158947
R415 VSS.n20 VSS 0.0158947
R416 VSS VSS.n45 0.0158947
R417 VSS VSS.n52 0.0158947
R418 VSS.n53 VSS 0.0158947
R419 VSS VSS.n31 0.0158947
R420 VSS VSS.n0 0.0158947
R421 VSS VSS.n9 0.00405263
R422 VSS.n21 VSS 0.00405263
R423 VSS VSS.n4 0.00405263
R424 VSS.n54 VSS 0.00405263
R425 VSS VSS.n7 0.00405263
R426 VSS.n40 VSS 0.00247368
R427 VSS.n32 VSS 0.00247368
R428 VSS.n10 VSS 0.000894737
R429 VSS.n22 VSS 0.000894737
R430 VSS.n41 VSS 0.000894737
R431 VSS.n5 VSS 0.000894737
R432 VSS.n55 VSS 0.000894737
R433 VSS.n8 VSS 0.000894737
R434 VSS.n33 VSS 0.000894737
R435 S1.n0 S1.t5 31.528
R436 S1.n4 S1.t0 31.528
R437 S1.n12 S1.t6 25.7638
R438 S1.n2 S1.t1 25.7638
R439 S1.n0 S1.t3 15.3826
R440 S1.n4 S1.t2 15.3826
R441 S1.n12 S1.t7 13.2969
R442 S1.n2 S1.t4 13.2969
R443 S1.n17 S1.n0 7.62076
R444 S1.n5 S1.n4 7.62076
R445 S1.n11 S1.n10 6.90126
R446 S1.n7 S1.n6 4.54699
R447 S1.n16 S1.n15 4.54699
R448 S1.n14 S1 4.52833
R449 S1.n8 S1 4.52833
R450 S1.n13 S1.n11 2.25478
R451 S1.n10 S1.n3 2.25386
R452 S1.n9 S1.n3 2.2505
R453 S1.n13 S1.n1 2.2505
R454 S1.n13 S1.n12 2.11815
R455 S1.n3 S1.n2 2.11815
R456 S1.n8 S1.n7 1.33991
R457 S1.n16 S1.n14 1.33848
R458 S1.n7 S1.n5 1.12145
R459 S1.n17 S1.n16 1.12145
R460 S1.n6 S1 0.0780197
R461 S1.n15 S1 0.0780197
R462 S1.n6 S1 0.0359098
R463 S1.n15 S1 0.032959
R464 S1.n9 S1.n8 0.0289694
R465 S1.n14 S1.n1 0.0289694
R466 S1.n11 S1 0.0169815
R467 S1.n10 S1 0.0160631
R468 S1 S1.n9 0.00233673
R469 S1 S1.n1 0.00233673
R470 S1 S1.n5 0.00197541
R471 S1 S1.n17 0.00197541
R472 S1 S1.n13 0.00142783
R473 S1 S1.n3 0.00142783
R474 S0.n0 S0.t9 31.528
R475 S0.n20 S0.t1 31.528
R476 S0.n12 S0.t13 31.528
R477 S0.n2 S0.t12 31.528
R478 S0.n29 S0.t2 25.7638
R479 S0.n10 S0.t0 25.7638
R480 S0.n15 S0.t4 25.7638
R481 S0.n5 S0.t10 25.7638
R482 S0.n0 S0.t5 15.3826
R483 S0.n20 S0.t3 15.3826
R484 S0.n12 S0.t14 15.3826
R485 S0.n2 S0.t7 15.3826
R486 S0.n29 S0.t8 13.2969
R487 S0.n10 S0.t6 13.2969
R488 S0.n15 S0.t11 13.2969
R489 S0.n5 S0.t15 13.2969
R490 S0.n13 S0.n12 7.6291
R491 S0.n3 S0.n2 7.6289
R492 S0.n1 S0.n0 7.62076
R493 S0.n21 S0.n20 7.62076
R494 S0.n19 S0 4.53443
R495 S0.n35 S0 4.53443
R496 S0.n32 S0 4.52853
R497 S0.n31 S0 4.52833
R498 S0.n25 S0 4.52833
R499 S0.n17 S0 4.52833
R500 S0.n7 S0 4.52833
R501 S0.n30 S0.n28 2.25478
R502 S0.n27 S0.n11 2.25386
R503 S0.n26 S0.n11 2.2505
R504 S0.n30 S0.n9 2.2505
R505 S0.n33 S0.n8 2.19776
R506 S0.n23 S0.n18 2.19633
R507 S0.n30 S0.n29 2.11815
R508 S0.n11 S0.n10 2.11815
R509 S0.n16 S0.n15 2.11815
R510 S0.n6 S0.n5 2.11815
R511 S0.n28 S0.n27 1.87738
R512 S0.n22 S0.n21 1.5005
R513 S0.n34 S0.n1 1.5005
R514 S0.n25 S0.n24 1.31185
R515 S0.n32 S0.n31 1.31042
R516 S0.n18 S0.n17 1.2853
R517 S0.n8 S0.n7 1.28387
R518 S0.n6 S0.n4 1.13046
R519 S0.n16 S0.n14 1.13
R520 S0.n8 S0.n3 0.948428
R521 S0.n18 S0.n13 0.948389
R522 S0.n13 S0 0.109321
R523 S0.n3 S0 0.108522
R524 S0 S0.n35 0.0780742
R525 S0.n19 S0 0.0780197
R526 S0.n21 S0.n19 0.0373852
R527 S0.n35 S0.n1 0.0373852
R528 S0.n24 S0.n23 0.0359098
R529 S0.n33 S0.n32 0.0359098
R530 S0.n17 S0.n14 0.0303837
R531 S0.n7 S0.n4 0.0303834
R532 S0.n26 S0.n25 0.0289694
R533 S0.n31 S0.n9 0.0289694
R534 S0.n28 S0 0.0169815
R535 S0.n27 S0 0.0160631
R536 S0 S0.n1 0.00935246
R537 S0.n22 S0 0.00345082
R538 S0 S0.n34 0.00345082
R539 S0 S0.n26 0.00233673
R540 S0 S0.n9 0.00233673
R541 S0.n23 S0.n22 0.00197541
R542 S0.n34 S0.n33 0.00197541
R543 S0.n4 S0 0.00192201
R544 S0.n14 S0 0.00192164
R545 S0 S0.n30 0.00142783
R546 S0 S0.n11 0.00142783
R547 S0 S0.n16 0.00142783
R548 S0 S0.n6 0.00142783
R549 I4.n0 I4.t1 31.528
R550 I4.n0 I4.t0 15.3826
R551 I4 I4.n0 8.74076
R552 I3.n0 I3.t1 30.9379
R553 I3.n0 I3.t0 21.6422
R554 I3 I3.n0 4.0005
R555 I6.n0 I6.t1 31.528
R556 I6.n0 I6.t0 15.3826
R557 I6.n1 I6.n0 8.74076
R558 I6.n1 I6 0.116616
R559 I6 I6.n1 0.00202542
R560 I1.n0 I1.t1 30.9379
R561 I1.n0 I1.t0 21.6422
R562 I1 I1.n0 4.005
R563 I2.n0 I2.t0 31.528
R564 I2.n0 I2.t1 15.3826
R565 I2.n1 I2.n0 8.74076
R566 I2.n1 I2 0.00197541
R567 I2 I2.n1 0.00197541
R568 I7.n0 I7.t0 30.9379
R569 I7.n0 I7.t1 21.6422
R570 I7 I7.n0 4.0005
R571 I5.n0 I5.t0 30.9379
R572 I5.n0 I5.t1 21.6422
R573 I5 I5.n0 4.005
R574 OUT OUT.n2 7.15141
R575 OUT.n3 OUT.n1 3.2163
R576 OUT.n1 OUT.t0 2.2755
R577 OUT.n1 OUT.n0 2.2755
R578 OUT OUT.n3 0.0537653
R579 OUT.n3 OUT 0.0119545
R580 I0.n0 I0.t0 31.528
R581 I0.n0 I0.t1 15.3826
R582 I0 I0.n0 8.74076
C0 I4 S0 0.00512f
C1 mux_2x1_ibr_0.nand2_ibr_1.IN2 a_4178_1307# 0.00372f
C2 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT 0.0241f
C3 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 VDD 0.405f
C4 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 I6 1.04e-19
C5 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT a_2490_n1395# 9.43e-19
C6 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT S0 0.00112f
C7 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.63f
C8 I0 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 3e-19
C9 S0 a_1364_1307# 0.0151f
C10 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 0.285f
C11 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 S1 0.00266f
C12 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 I0 0.0148f
C13 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 a_1364_n1395# 0.00211f
C14 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT a_1927_n1395# 0.00949f
C15 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT VDD 0.664f
C16 mux_2x1_ibr_0.nand2_ibr_2.OUT VDD 0.635f
C17 a_801_707# mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.0964f
C18 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 S1 4.51e-21
C19 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 VDD 0.405f
C20 a_1927_707# S1 2.15e-19
C21 mux_2x1_ibr_0.I1 S0 6.5e-20
C22 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 S0 0.207f
C23 I0 S0 0.00507f
C24 S0 a_1364_n1395# 0.0151f
C25 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.053f
C26 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 a_801_n1395# 0.069f
C27 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 a_801_1307# 0.00372f
C28 a_801_n1395# mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.00372f
C29 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.00212f
C30 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.053f
C31 a_4178_707# VDD 0.00444f
C32 a_801_707# S0 6.89e-19
C33 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_4x1_ibr_0.mux_2x1_ibr_2.I1 0.328f
C34 S0 a_801_n1395# 9.5e-19
C35 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.0189f
C36 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 I2 0.0036f
C37 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.0102f
C38 a_238_n1395# mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.069f
C39 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT VDD 0.664f
C40 VDD mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.461f
C41 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 S0 0.136f
C42 S0 a_238_n1395# 0.0144f
C43 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 a_3053_n795# 0.00372f
C44 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 S0 0.378f
C45 a_1927_707# S0 2.62e-19
C46 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.12f
C47 a_1927_n795# VDD 0.00444f
C48 S2 a_3615_1307# 0.0144f
C49 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT a_2490_1307# 9.43e-19
C50 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 S0 0.162f
C51 mux_2x1_ibr_0.I0 mux_2x1_ibr_0.nand2_ibr_2.IN2 0.051f
C52 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT 0.0112f
C53 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.0102f
C54 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT a_1927_1307# 0.00949f
C55 mux_2x1_ibr_0.I0 mux_2x1_ibr_0.I1 2.74e-20
C56 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_2x1_ibr_0.I0 0.0073f
C57 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 a_801_n795# 1.5e-19
C58 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT VDD 0.634f
C59 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 a_3053_707# 0.00375f
C60 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 a_801_1307# 0.069f
C61 I6 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT 0.202f
C62 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 9.55e-20
C63 a_801_n795# S0 6.89e-19
C64 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.0048f
C65 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.00212f
C66 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT 0.0241f
C67 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 S0 0.162f
C68 VDD mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.462f
C69 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT a_3615_1307# 9.46e-19
C70 mux_2x1_ibr_0.nand2_ibr_2.IN2 S2 0.136f
C71 S1 mux_4x1_ibr_1.mux_2x1_ibr_2.I1 0.0593f
C72 I4 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.0036f
C73 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT a_3053_1307# 0.00949f
C74 mux_2x1_ibr_0.I1 S2 0.0594f
C75 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 S2 0.00519f
C76 OUT a_4178_1307# 0.069f
C77 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT 0.053f
C78 a_1927_707# mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT 0.0964f
C79 VDD mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.46f
C80 I6 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.0473f
C81 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_4x1_ibr_1.mux_2x1_ibr_2.I1 0.00147f
C82 a_2490_n1395# mux_4x1_ibr_1.mux_2x1_ibr_2.I1 0.00372f
C83 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.0189f
C84 S0 mux_4x1_ibr_1.mux_2x1_ibr_2.I1 0.0109f
C85 a_1927_n795# I2 0.00293f
C86 mux_2x1_ibr_0.nand2_ibr_2.IN2 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT 0.0113f
C87 mux_2x1_ibr_0.nand2_ibr_2.OUT mux_2x1_ibr_0.nand2_ibr_2.IN2 0.12f
C88 I6 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 0.0036f
C89 a_1927_n1395# mux_4x1_ibr_1.mux_2x1_ibr_2.I1 0.069f
C90 mux_2x1_ibr_0.nand2_ibr_1.IN2 OUT 0.109f
C91 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT I4 3e-19
C92 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 S1 0.0863f
C93 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT mux_2x1_ibr_0.I1 0.329f
C94 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT 0.25f
C95 mux_2x1_ibr_0.nand2_ibr_2.OUT mux_4x1_ibr_0.mux_2x1_ibr_2.I0 3.46e-19
C96 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 0.0646f
C97 a_4178_707# mux_2x1_ibr_0.nand2_ibr_2.IN2 0.00372f
C98 a_2490_n1395# S1 0.0144f
C99 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.00216f
C100 S0 S1 0.00413f
C101 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.0106f
C102 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.00212f
C103 a_1927_707# mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.00372f
C104 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 a_3053_n1395# 2.44e-19
C105 mux_4x1_ibr_0.mux_2x1_ibr_2.I1 VDD 0.423f
C106 VDD mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.456f
C107 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.109f
C108 S0 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.0532f
C109 I0 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.202f
C110 mux_4x1_ibr_0.mux_2x1_ibr_2.I1 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.11f
C111 VDD a_3615_1307# 3.14e-19
C112 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 a_2490_n1395# 1.04e-19
C113 a_1927_n795# mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT 0.0964f
C114 I2 VDD 0.261f
C115 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT a_3053_n795# 0.0964f
C116 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 S0 0.207f
C117 S0 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.368f
C118 VDD a_238_1307# 3.14e-19
C119 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT a_801_n1395# 0.00949f
C120 VDD a_3053_1307# 0.00444f
C121 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 a_1927_n1395# 2.44e-19
C122 VDD a_3053_n795# 0.00444f
C123 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 a_3053_1307# 0.00372f
C124 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.0112f
C125 VDD a_2490_1307# 3.14e-19
C126 mux_2x1_ibr_0.nand2_ibr_1.IN2 S2 0.341f
C127 I4 VDD 0.258f
C128 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 a_2490_1307# 0.069f
C129 VDD a_1927_1307# 0.00444f
C130 mux_2x1_ibr_0.nand2_ibr_2.OUT a_4178_1307# 0.00949f
C131 mux_2x1_ibr_0.I0 S1 0.0118f
C132 a_1927_n795# mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.00372f
C133 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT VDD 0.665f
C134 VDD a_1364_1307# 3.14e-19
C135 mux_2x1_ibr_0.nand2_ibr_2.IN2 VDD 0.402f
C136 a_3053_707# S1 2.62e-19
C137 I6 VDD 0.258f
C138 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 S1 0.16f
C139 mux_2x1_ibr_0.I1 VDD 0.423f
C140 mux_2x1_ibr_0.I0 a_3053_n1395# 0.069f
C141 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 VDD 1.41f
C142 I0 VDD 0.258f
C143 VDD a_1364_n1395# 3.14e-19
C144 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT S1 0.113f
C145 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_2x1_ibr_0.I0 0.0449f
C146 mux_2x1_ibr_0.I1 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.109f
C147 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.00154f
C148 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT a_801_1307# 0.00949f
C149 a_801_707# VDD 0.00444f
C150 a_801_n795# mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.0964f
C151 mux_2x1_ibr_0.nand2_ibr_1.IN2 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT 0.0106f
C152 mux_2x1_ibr_0.nand2_ibr_1.IN2 mux_2x1_ibr_0.nand2_ibr_2.OUT 0.053f
C153 VDD a_801_n1395# 0.00444f
C154 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 0.0646f
C155 mux_2x1_ibr_0.I0 S0 6.5e-20
C156 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.053f
C157 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.12f
C158 S0 a_801_1307# 9.5e-19
C159 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 VDD 0.405f
C160 S2 S1 0.0018f
C161 VDD a_238_n1395# 3.14e-19
C162 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 VDD 0.46f
C163 a_1927_707# VDD 0.00444f
C164 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT S0 0.00113f
C165 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 a_238_1307# 0.069f
C166 a_1364_n1395# mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.069f
C167 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 S1 0.00266f
C168 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 VDD 0.404f
C169 mux_4x1_ibr_0.mux_2x1_ibr_2.I1 a_2490_1307# 0.00372f
C170 OUT mux_2x1_ibr_0.I0 1.49e-19
C171 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.00212f
C172 a_4178_1307# VDD 0.00444f
C173 mux_4x1_ibr_0.mux_2x1_ibr_2.I1 a_1927_1307# 0.069f
C174 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT S1 0.00228f
C175 mux_2x1_ibr_0.nand2_ibr_2.OUT S1 1.54e-19
C176 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.0112f
C177 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 S1 0.16f
C178 a_801_n795# VDD 0.00444f
C179 mux_4x1_ibr_1.mux_2x1_ibr_2.I1 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.11f
C180 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 9.55e-20
C181 I6 mux_4x1_ibr_0.mux_2x1_ibr_2.I1 1.36e-19
C182 I2 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT 0.203f
C183 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 VDD 0.404f
C184 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 S0 0.136f
C185 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 mux_2x1_ibr_0.I0 3.43e-19
C186 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_4x1_ibr_0.mux_2x1_ibr_2.I1 0.00147f
C187 I2 I6 0.00246f
C188 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.109f
C189 mux_2x1_ibr_0.I1 a_3615_1307# 0.00372f
C190 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 9.55e-20
C191 S1 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.342f
C192 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 I2 1.04e-19
C193 mux_2x1_ibr_0.nand2_ibr_1.IN2 VDD 0.461f
C194 OUT S2 0.00946f
C195 mux_2x1_ibr_0.I1 a_3053_1307# 0.069f
C196 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 a_3053_1307# 2.44e-19
C197 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.00342f
C198 a_1927_n795# S1 2.15e-19
C199 a_3053_n1395# mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.00372f
C200 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 mux_4x1_ibr_0.mux_2x1_ibr_2.I1 0.109f
C201 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.63f
C202 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.00154f
C203 mux_2x1_ibr_0.I0 S2 4.25e-19
C204 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.053f
C205 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 a_2490_1307# 1.04e-19
C206 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 I2 0.0473f
C207 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 I4 0.0148f
C208 I0 I4 0.00246f
C209 a_2490_n1395# mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.069f
C210 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT S0 0.0532f
C211 a_3053_707# S2 2.16e-19
C212 S0 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 4.45e-19
C213 VDD mux_4x1_ibr_1.mux_2x1_ibr_2.I1 0.423f
C214 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 a_1927_1307# 2.44e-19
C215 I4 a_801_707# 0.00293f
C216 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 a_1927_n795# 8.2e-19
C217 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.00212f
C218 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT S1 0.00227f
C219 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 a_1364_1307# 0.00211f
C220 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_2x1_ibr_0.nand2_ibr_2.IN2 0.00494f
C221 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 I6 0.01f
C222 a_1927_n795# S0 2.62e-19
C223 mux_2x1_ibr_0.nand2_ibr_2.OUT OUT 0.303f
C224 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_2x1_ibr_0.I1 5.19e-19
C225 VDD S1 1.58f
C226 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT a_3053_n1395# 0.00949f
C227 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 a_1927_1307# 0.00372f
C228 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT 0.12f
C229 S1 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.342f
C230 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 a_801_707# 1.5e-19
C231 mux_2x1_ibr_0.nand2_ibr_2.OUT mux_2x1_ibr_0.I0 0.234f
C232 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT 0.25f
C233 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT 0.12f
C234 mux_4x1_ibr_1.mux_2x1_ibr_2.I1 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.109f
C235 a_3053_707# mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT 0.0964f
C236 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 a_1364_1307# 0.069f
C237 a_3053_n1395# VDD 0.00444f
C238 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 a_3053_707# 0.00372f
C239 VDD mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.664f
C240 I6 a_1927_707# 0.00293f
C241 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 I4 0.0473f
C242 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 0.00216f
C243 mux_2x1_ibr_0.I0 a_4178_707# 0.00293f
C244 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 VDD 1.36f
C245 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 9.55e-20
C246 VDD mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.456f
C247 I0 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.0036f
C248 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.0169f
C249 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT 0.0112f
C250 a_2490_n1395# VDD 3.14e-19
C251 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 a_1927_707# 8.2e-19
C252 VDD S0 3.48f
C253 mux_2x1_ibr_0.I0 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.11f
C254 S1 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 4.51e-21
C255 mux_2x1_ibr_0.nand2_ibr_1.IN2 a_3615_1307# 0.069f
C256 S0 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 4.45e-19
C257 a_1927_n1395# VDD 0.00444f
C258 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.00212f
C259 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT S2 0.109f
C260 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.0048f
C261 mux_2x1_ibr_0.nand2_ibr_2.OUT S2 4.46e-19
C262 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 S2 3.66e-19
C263 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 a_801_707# 0.00372f
C264 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.0169f
C265 a_4178_707# S2 2.62e-19
C266 S0 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.378f
C267 a_801_n795# I0 0.00293f
C268 I2 mux_4x1_ibr_1.mux_2x1_ibr_2.I1 1.36e-19
C269 OUT VDD 0.234f
C270 a_1927_n1395# mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.00372f
C271 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT mux_2x1_ibr_0.I0 0.419f
C272 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 I0 0.0473f
C273 mux_4x1_ibr_0.mux_2x1_ibr_2.I1 S1 0.0593f
C274 mux_2x1_ibr_0.nand2_ibr_1.IN2 mux_2x1_ibr_0.nand2_ibr_2.IN2 0.00212f
C275 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT 0.12f
C276 mux_2x1_ibr_0.I0 VDD 1.44f
C277 mux_2x1_ibr_0.nand2_ibr_1.IN2 mux_2x1_ibr_0.I1 0.11f
C278 I2 S1 0.00826f
C279 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT 0.12f
C280 a_3053_707# VDD 0.00444f
C281 VDD a_801_1307# 0.00444f
C282 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 VDD 0.405f
C283 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.053f
C284 S1 a_3053_n795# 2.62e-19
C285 mux_2x1_ibr_0.nand2_ibr_2.OUT a_4178_707# 0.0964f
C286 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT VDD 0.665f
C287 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_4x1_ibr_1.mux_2x1_ibr_2.I1 0.328f
C288 mux_4x1_ibr_0.mux_2x1_ibr_2.I1 S0 0.0109f
C289 S1 a_2490_1307# 0.0144f
C290 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 I2 0.01f
C291 S0 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.368f
C292 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.0106f
C293 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.00216f
C294 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 a_3053_n795# 0.00375f
C295 S0 a_238_1307# 0.0144f
C296 S2 VDD 0.596f
C297 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT S1 0.113f
C298 I4 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.202f
C299 mux_2x1_ibr_0.nand2_ibr_2.IN2 S1 2.44e-19
C300 I6 S1 0.00831f
C301 S2 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 4.52e-21
C302 mux_2x1_ibr_0.I1 S1 0.00946f
C303 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 S1 0.0874f
C304 a_801_n795# mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.00372f
C305 a_3053_n1395# VSS 0.0676f
C306 a_2490_n1395# VSS 0.0676f
C307 a_1927_n1395# VSS 0.0676f
C308 a_1364_n1395# VSS 0.0676f
C309 a_801_n1395# VSS 0.0676f
C310 a_238_n1395# VSS 0.0678f
C311 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 VSS 0.412f
C312 mux_4x1_ibr_1.mux_2x1_ibr_2.I1 VSS 0.416f
C313 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 VSS 0.412f
C314 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 VSS 0.435f
C315 a_3053_n795# VSS 0.0676f
C316 a_1927_n795# VSS 0.0676f
C317 a_801_n795# VSS 0.0676f
C318 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT VSS 0.598f
C319 mux_4x1_ibr_1.mux_2x1_ibr_2.I0 VSS 0.771f
C320 mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 VSS 0.416f
C321 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT VSS 0.489f
C322 I2 VSS 0.226f
C323 mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 VSS 0.417f
C324 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT VSS 0.43f
C325 I0 VSS 0.226f
C326 mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 VSS 0.436f
C327 a_4178_707# VSS 0.0676f
C328 mux_2x1_ibr_0.I0 VSS 1.4f
C329 mux_2x1_ibr_0.nand2_ibr_2.IN2 VSS 0.422f
C330 a_3053_707# VSS 0.0676f
C331 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 VSS 0.417f
C332 a_1927_707# VSS 0.0676f
C333 I6 VSS 0.226f
C334 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 VSS 0.417f
C335 a_801_707# VSS 0.0676f
C336 I4 VSS 0.226f
C337 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 VSS 0.436f
C338 a_4178_1307# VSS 0.0676f
C339 a_3615_1307# VSS 0.0676f
C340 a_3053_1307# VSS 0.0676f
C341 a_2490_1307# VSS 0.0676f
C342 a_1927_1307# VSS 0.0676f
C343 a_1364_1307# VSS 0.0676f
C344 a_801_1307# VSS 0.0676f
C345 a_238_1307# VSS 0.0678f
C346 OUT VSS 0.14f
C347 mux_4x1_ibr_0.mux_2x1_ibr_2.I0 VSS 0.714f
C348 mux_2x1_ibr_0.nand2_ibr_2.OUT VSS 0.653f
C349 mux_2x1_ibr_0.nand2_ibr_1.IN2 VSS 0.412f
C350 S2 VSS 0.714f
C351 mux_2x1_ibr_0.I1 VSS 0.416f
C352 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT VSS 0.489f
C353 mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 VSS 0.412f
C354 S1 VSS 1.53f
C355 mux_4x1_ibr_0.mux_2x1_ibr_2.I1 VSS 0.416f
C356 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT VSS 0.489f
C357 mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 VSS 0.412f
C358 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT VSS 0.43f
C359 mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 VSS 0.435f
C360 S0 VSS 3.98f
C361 VDD VSS 27.8f
C362 S0.t5 VSS 0.0227f
C363 S0.t9 VSS 0.0284f
C364 S0.n0 VSS 0.0671f
C365 S0.n1 VSS 0.0171f
C366 S0.t7 VSS 0.0227f
C367 S0.t12 VSS 0.0284f
C368 S0.n2 VSS 0.0672f
C369 S0.n3 VSS 0.0353f
C370 S0.n4 VSS 0.00656f
C371 S0.t15 VSS 0.00827f
C372 S0.t10 VSS 0.0329f
C373 S0.n5 VSS 0.0535f
C374 S0.n6 VSS 0.0184f
C375 S0.n7 VSS 0.131f
C376 S0.n8 VSS 0.325f
C377 S0.n9 VSS 0.00689f
C378 S0.t0 VSS 0.0329f
C379 S0.t6 VSS 0.00827f
C380 S0.n10 VSS 0.0535f
C381 S0.n11 VSS 0.0184f
C382 S0.t14 VSS 0.0227f
C383 S0.t13 VSS 0.0284f
C384 S0.n12 VSS 0.0672f
C385 S0.n13 VSS 0.0352f
C386 S0.n14 VSS 0.00656f
C387 S0.t4 VSS 0.0329f
C388 S0.t11 VSS 0.00827f
C389 S0.n15 VSS 0.0535f
C390 S0.n16 VSS 0.0184f
C391 S0.n17 VSS 0.131f
C392 S0.n18 VSS 0.325f
C393 S0.n19 VSS 0.00965f
C394 S0.t3 VSS 0.0227f
C395 S0.t1 VSS 0.0284f
C396 S0.n20 VSS 0.0671f
C397 S0.n21 VSS 0.0274f
C398 S0.n22 VSS 3.88e-19
C399 S0.n23 VSS 0.19f
C400 S0.n24 VSS 0.134f
C401 S0.n25 VSS 0.133f
C402 S0.n26 VSS 0.00689f
C403 S0.n27 VSS 0.189f
C404 S0.n28 VSS 0.189f
C405 S0.t8 VSS 0.00827f
C406 S0.t2 VSS 0.0329f
C407 S0.n29 VSS 0.0535f
C408 S0.n30 VSS 0.0184f
C409 S0.n31 VSS 0.133f
C410 S0.n32 VSS 0.134f
C411 S0.n33 VSS 0.19f
C412 S0.n34 VSS 3.88e-19
C413 S0.n35 VSS 0.00964f
C414 VDD.t38 VSS 0.0685f
C415 VDD.n0 VSS 0.0327f
C416 VDD.t87 VSS 0.00199f
C417 VDD.n1 VSS 0.0166f
C418 VDD.t103 VSS 0.00199f
C419 VDD.n2 VSS 0.00814f
C420 VDD.n3 VSS 0.00263f
C421 VDD.t32 VSS 0.0347f
C422 VDD.n4 VSS 0.00263f
C423 VDD.n5 VSS 0.00289f
C424 VDD.t78 VSS 0.0343f
C425 VDD.t4 VSS 0.0317f
C426 VDD.n6 VSS 0.0163f
C427 VDD.n7 VSS 0.00814f
C428 VDD.t5 VSS 0.00216f
C429 VDD.t43 VSS 0.00199f
C430 VDD.n8 VSS 0.0166f
C431 VDD.n9 VSS 0.0183f
C432 VDD.n10 VSS 0.00644f
C433 VDD.n11 VSS 0.0105f
C434 VDD.t102 VSS 0.00263f
C435 VDD.n12 VSS 0.00263f
C436 VDD.n13 VSS 0.013f
C437 VDD.n14 VSS 0.0121f
C438 VDD.n15 VSS 0.00814f
C439 VDD.n16 VSS 0.0163f
C440 VDD.t101 VSS 0.0317f
C441 VDD.t91 VSS 0.0347f
C442 VDD.n17 VSS 0.0163f
C443 VDD.t6 VSS 0.0317f
C444 VDD.t61 VSS 0.0347f
C445 VDD.n18 VSS 0.0163f
C446 VDD.t109 VSS 0.00263f
C447 VDD.n19 VSS 0.00263f
C448 VDD.t108 VSS 0.0317f
C449 VDD.t22 VSS 0.0347f
C450 VDD.n20 VSS 0.0163f
C451 VDD.t14 VSS 0.00216f
C452 VDD.t29 VSS 0.00199f
C453 VDD.n21 VSS 0.0166f
C454 VDD.n22 VSS 0.0183f
C455 VDD.n23 VSS 0.00263f
C456 VDD.t13 VSS 0.0317f
C457 VDD.t71 VSS 0.0347f
C458 VDD.t59 VSS 0.0316f
C459 VDD.n24 VSS 0.0163f
C460 VDD.t60 VSS 0.00282f
C461 VDD.n25 VSS 0.0202f
C462 VDD.n26 VSS 0.0105f
C463 VDD.n27 VSS 0.00644f
C464 VDD.n28 VSS 0.00814f
C465 VDD.n29 VSS 0.013f
C466 VDD.n30 VSS 0.012f
C467 VDD.n31 VSS 0.00542f
C468 VDD.n32 VSS 0.0105f
C469 VDD.n33 VSS 0.00644f
C470 VDD.t7 VSS 0.00216f
C471 VDD.n34 VSS 0.0183f
C472 VDD.n35 VSS 0.0166f
C473 VDD.t75 VSS 0.00264f
C474 VDD.t107 VSS 0.00264f
C475 VDD.t86 VSS 0.0359f
C476 VDD.n36 VSS 0.0283f
C477 VDD.t74 VSS 0.0295f
C478 VDD.t106 VSS 0.0296f
C479 VDD.n38 VSS 0.0294f
C480 VDD.n39 VSS 0.0217f
C481 VDD.n40 VSS 0.0124f
C482 VDD.n41 VSS 0.00263f
C483 VDD.n42 VSS 0.00263f
C484 VDD.t64 VSS 0.0685f
C485 VDD.n43 VSS 0.0327f
C486 VDD.t35 VSS 0.00199f
C487 VDD.t105 VSS 0.00216f
C488 VDD.n44 VSS 0.00814f
C489 VDD.n45 VSS 0.00263f
C490 VDD.t54 VSS 0.0347f
C491 VDD.n46 VSS 0.00263f
C492 VDD.t94 VSS 0.0347f
C493 VDD.n47 VSS 0.00263f
C494 VDD.t3 VSS 0.00216f
C495 VDD.n48 VSS 0.0183f
C496 VDD.t10 VSS 0.0347f
C497 VDD.n49 VSS 0.00263f
C498 VDD.t58 VSS 0.00216f
C499 VDD.t21 VSS 0.00199f
C500 VDD.n50 VSS 0.00289f
C501 VDD.n51 VSS 0.00814f
C502 VDD.t47 VSS 0.0296f
C503 VDD.t88 VSS 0.0343f
C504 VDD.n52 VSS 0.0163f
C505 VDD.t20 VSS 0.018f
C506 VDD.n53 VSS 0.0288f
C507 VDD.t48 VSS 0.00269f
C508 VDD.n54 VSS 0.00263f
C509 VDD.n55 VSS 0.00263f
C510 VDD.t1 VSS 0.00199f
C511 VDD.n56 VSS 0.0166f
C512 VDD.n57 VSS 0.0114f
C513 VDD.t81 VSS 0.0685f
C514 VDD.t84 VSS 0.0296f
C515 VDD.t85 VSS 0.00264f
C516 VDD.t31 VSS 0.00264f
C517 VDD.n58 VSS 0.00773f
C518 VDD.n59 VSS 0.0217f
C519 VDD.n60 VSS 0.0126f
C520 VDD.n61 VSS 0.00263f
C521 VDD.n62 VSS 0.00263f
C522 VDD.n63 VSS 0.0203f
C523 VDD.n64 VSS 0.026f
C524 VDD.n65 VSS 0.0158f
C525 VDD.n66 VSS 0.0217f
C526 VDD.n67 VSS 0.0294f
C527 VDD.t30 VSS 0.0295f
C528 VDD.n69 VSS 0.0283f
C529 VDD.t0 VSS 0.0359f
C530 VDD.n70 VSS 0.0327f
C531 VDD.n71 VSS 0.0163f
C532 VDD.n72 VSS 0.0259f
C533 VDD.n73 VSS 0.0252f
C534 VDD.n74 VSS 0.0203f
C535 VDD.n75 VSS 0.00949f
C536 VDD.n76 VSS 0.0166f
C537 VDD.n77 VSS 0.0183f
C538 VDD.n78 VSS 0.00289f
C539 VDD.t15 VSS 0.0343f
C540 VDD.t57 VSS 0.0317f
C541 VDD.n79 VSS 0.0163f
C542 VDD.n80 VSS 0.00814f
C543 VDD.n81 VSS 0.00644f
C544 VDD.n82 VSS 0.0105f
C545 VDD.t50 VSS 0.00263f
C546 VDD.n83 VSS 0.00263f
C547 VDD.n84 VSS 0.013f
C548 VDD.n85 VSS 0.0121f
C549 VDD.n86 VSS 0.00814f
C550 VDD.n87 VSS 0.0163f
C551 VDD.t49 VSS 0.0316f
C552 VDD.t25 VSS 0.0346f
C553 VDD.t2 VSS 0.0317f
C554 VDD.n88 VSS 0.0163f
C555 VDD.n89 VSS 0.00814f
C556 VDD.n90 VSS 0.00644f
C557 VDD.n91 VSS 0.0105f
C558 VDD.t9 VSS 0.00263f
C559 VDD.n92 VSS 0.00263f
C560 VDD.n93 VSS 0.013f
C561 VDD.n94 VSS 0.0121f
C562 VDD.n95 VSS 0.00814f
C563 VDD.n96 VSS 0.0163f
C564 VDD.t8 VSS 0.0317f
C565 VDD.t110 VSS 0.0347f
C566 VDD.t41 VSS 0.0317f
C567 VDD.n97 VSS 0.0163f
C568 VDD.n98 VSS 0.00814f
C569 VDD.t42 VSS 0.00216f
C570 VDD.n99 VSS 0.0183f
C571 VDD.n100 VSS 0.00644f
C572 VDD.n101 VSS 0.0105f
C573 VDD.t100 VSS 0.00263f
C574 VDD.n102 VSS 0.00263f
C575 VDD.n103 VSS 0.013f
C576 VDD.n104 VSS 0.012f
C577 VDD.n105 VSS 0.00542f
C578 VDD.n106 VSS 0.0163f
C579 VDD.t99 VSS 0.0317f
C580 VDD.t44 VSS 0.0347f
C581 VDD.n107 VSS 0.0163f
C582 VDD.t104 VSS 0.0317f
C583 VDD.t51 VSS 0.0347f
C584 VDD.t18 VSS 0.0316f
C585 VDD.n108 VSS 0.0163f
C586 VDD.t19 VSS 0.00282f
C587 VDD.n109 VSS 0.0202f
C588 VDD.n110 VSS 0.0105f
C589 VDD.n111 VSS 0.00644f
C590 VDD.n112 VSS 0.0183f
C591 VDD.n113 VSS 0.0166f
C592 VDD.t69 VSS 0.0296f
C593 VDD.t28 VSS 0.0359f
C594 VDD.n114 VSS 0.0283f
C595 VDD.t36 VSS 0.0295f
C596 VDD.t37 VSS 0.00274f
C597 VDD.n116 VSS 0.0331f
C598 VDD.n117 VSS 0.0294f
C599 VDD.t70 VSS 0.00274f
C600 VDD.n118 VSS 0.033f
C601 VDD.n119 VSS 0.00812f
C602 VDD.n120 VSS 0.0111f
C603 VDD.n121 VSS 0.0163f
C604 VDD.n122 VSS 0.0209f
C605 VDD.n123 VSS 0.0292f
C606 VDD.n124 VSS 0.0124f
C607 VDD.n125 VSS 0.0217f
C608 VDD.n126 VSS 0.00812f
C609 VDD.n127 VSS 0.0111f
C610 VDD.n128 VSS 0.0163f
.ends

