* NGSPICE file created from Local_Enc_v2_flat.ext - technology: gf180mcuC

.subckt Local_Enc_v2_flat Q Ri-1 Ri Ci VDD VSS QB
X0 NAND_9.B NAND_13.B VDD.t39 VDD.t38 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X1 a_305_1140# NAND_9.B VSS.t19 VSS.t18 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X2 a_305_3086# Ci.t0 VSS.t14 VSS.t13 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X3 a_305_6005# NAND_13.B VSS.t22 VSS.t21 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X4 QB NAND_3.B VDD.t1 VDD.t0 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X5 NAND_13.B NAND_1.B a_305_6981# VSS.t6 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X6 NAND_13.A NAND_12.B VDD.t6 VDD.t5 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X7 NAND_13.A NAND_12.A a_305_5030# VSS.t10 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X8 Q NAND_9.B VDD.t34 VDD.t33 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X9 VDD Ri-1.t0 NAND_1.B VDD.t40 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X10 NAND_13.B NAND_1.B VDD.t11 VDD.t10 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X11 a_305_2111# NAND_9.B VSS.t17 VSS.t16 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X12 VDD Ri.t0 NAND_12.A VDD.t14 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X13 a_305_165# NAND_3.B VSS.t1 VSS.t0 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X14 VDD NAND_9.B NAND_3.B VDD.t30 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X15 NAND_1.B Ri-1.t1 a_305_7966# VSS.t24 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X16 a_305_6981# NAND_1.B VSS.t5 VSS.t4 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X17 a_305_5030# NAND_12.B VSS.t3 VSS.t2 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X18 VDD Ci.t1 NAND_12.B VDD.t2 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X19 VDD Q.t3 QB.t1 VDD.t35 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X20 NAND_1.B Ri-1.t2 VDD.t44 VDD.t43 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X21 NAND_12.A Ri.t1 VDD.t18 VDD.t17 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X22 NAND_12.A Ri.t2 a_305_4056# VSS.t7 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X23 VDD NAND_13.A NAND_9.B VDD.t25 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X24 NAND_3.B NAND_9.B VDD.t29 VDD.t28 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X25 NAND_3.B NAND_9.B a_305_1140# VSS.t15 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X26 a_305_7966# Ri-1.t3 VSS.t26 VSS.t25 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X27 NAND_9.B NAND_13.A a_305_6005# VSS.t12 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X28 NAND_12.B Ci.t2 VDD.t13 VDD.t12 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X29 NAND_12.B Ci.t3 a_305_3086# VSS.t23 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X30 QB Q.t4 a_305_165# VSS.t20 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X31 VDD QB.t3 Q.t0 VDD.t22 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X32 VDD NAND_12.A NAND_13.A VDD.t19 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X33 VDD NAND_1.B NAND_13.B VDD.t7 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X34 a_305_4056# Ri.t3 VSS.t9 VSS.t8 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X35 Q QB.t4 a_305_2111# VSS.t11 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
R0 VDD.n1 VDD.t40 178.431
R1 VDD.n4 VDD.t7 178.431
R2 VDD.n8 VDD.t25 178.431
R3 VDD.n12 VDD.t19 178.431
R4 VDD.n16 VDD.t14 178.431
R5 VDD.n20 VDD.t2 178.431
R6 VDD.n24 VDD.t22 178.431
R7 VDD.n28 VDD.t30 178.431
R8 VDD.n32 VDD.t35 178.431
R9 VDD.n1 VDD.t43 135.294
R10 VDD.n4 VDD.t10 135.294
R11 VDD.n8 VDD.t38 135.294
R12 VDD.n12 VDD.t5 135.294
R13 VDD.n16 VDD.t17 135.294
R14 VDD.n20 VDD.t12 135.294
R15 VDD.n24 VDD.t33 135.294
R16 VDD.n28 VDD.t28 135.294
R17 VDD.n32 VDD.t0 135.294
R18 VDD.n5 VDD.n3 6.69527
R19 VDD.n9 VDD.n7 6.69527
R20 VDD.n13 VDD.n11 6.69527
R21 VDD.n17 VDD.n15 6.69527
R22 VDD.n21 VDD.n19 6.69527
R23 VDD.n25 VDD.n23 6.69527
R24 VDD.n29 VDD.n27 6.69527
R25 VDD.n33 VDD.n31 6.69527
R26 VDD.n2 VDD.n0 6.69527
R27 VDD.n6 VDD.t11 6.55815
R28 VDD.n10 VDD.t39 6.55815
R29 VDD.n14 VDD.t6 6.55815
R30 VDD.n18 VDD.t18 6.55815
R31 VDD.n22 VDD.t13 6.55815
R32 VDD.n26 VDD.t34 6.55815
R33 VDD.n30 VDD.t29 6.55815
R34 VDD.n34 VDD.t1 6.55815
R35 VDD.n42 VDD.t44 6.55815
R36 VDD.n5 VDD.n4 6.3005
R37 VDD.n9 VDD.n8 6.3005
R38 VDD.n13 VDD.n12 6.3005
R39 VDD.n17 VDD.n16 6.3005
R40 VDD.n21 VDD.n20 6.3005
R41 VDD.n25 VDD.n24 6.3005
R42 VDD.n29 VDD.n28 6.3005
R43 VDD.n33 VDD.n32 6.3005
R44 VDD.n2 VDD.n1 6.3005
R45 VDD.n35 VDD.n34 4.83679
R46 VDD VDD.n41 4.76956
R47 VDD.n40 VDD.n10 3.30864
R48 VDD.n41 VDD.n6 3.30818
R49 VDD.n39 VDD.n14 3.30724
R50 VDD.n38 VDD.n18 3.30677
R51 VDD.n37 VDD.n22 3.30677
R52 VDD.n36 VDD.n26 3.30677
R53 VDD.n35 VDD.n30 3.30631
R54 VDD.n39 VDD.n38 1.56955
R55 VDD.n36 VDD.n35 1.54914
R56 VDD.n40 VDD.n39 1.53098
R57 VDD.n41 VDD.n40 1.52295
R58 VDD.n38 VDD.n37 1.51604
R59 VDD.n37 VDD.n36 1.46348
R60 VDD.n6 VDD 0.0893
R61 VDD.n10 VDD 0.0893
R62 VDD.n14 VDD 0.0893
R63 VDD.n18 VDD 0.0893
R64 VDD.n22 VDD 0.0893
R65 VDD.n26 VDD 0.0893
R66 VDD.n30 VDD 0.0893
R67 VDD.n34 VDD 0.0893
R68 VDD VDD.n42 0.0893
R69 VDD.n42 VDD 0.0701
R70 VDD VDD.n5 0.0017
R71 VDD VDD.n9 0.0017
R72 VDD VDD.n13 0.0017
R73 VDD VDD.n17 0.0017
R74 VDD VDD.n21 0.0017
R75 VDD VDD.n25 0.0017
R76 VDD VDD.n29 0.0017
R77 VDD VDD.n33 0.0017
R78 VDD VDD.n2 0.0017
R79 VSS.t24 VSS.n1 6936.85
R80 VSS.n3 VSS.t25 6157.22
R81 VSS.n1 VSS.n0 4206.85
R82 VSS.t7 VSS.n32 2819.02
R83 VSS.t11 VSS.n20 2812.91
R84 VSS.t10 VSS.n38 2794.72
R85 VSS.t23 VSS.n26 2788.71
R86 VSS.t15 VSS.n14 2788.71
R87 VSS.t8 VSS.n33 1427.17
R88 VSS.t16 VSS.n21 1424.08
R89 VSS.t2 VSS.n39 1414.87
R90 VSS.t13 VSS.n27 1411.83
R91 VSS.t21 VSS.n7 1411.83
R92 VSS.t18 VSS.n15 1411.83
R93 VSS.t4 VSS.n3 1408.8
R94 VSS.n11 VSS.t20 682.1
R95 VSS.n11 VSS.t0 601.852
R96 VSS.n34 VSS.t7 600.543
R97 VSS.n22 VSS.t11 599.241
R98 VSS.n40 VSS.t10 595.366
R99 VSS.n28 VSS.t23 594.087
R100 VSS.n8 VSS.t12 594.087
R101 VSS.n16 VSS.t15 594.087
R102 VSS.n4 VSS.t6 592.812
R103 VSS.n2 VSS.t24 581.58
R104 VSS.n34 VSS.t8 529.891
R105 VSS.n22 VSS.t16 528.742
R106 VSS.n40 VSS.t2 525.323
R107 VSS.n28 VSS.t13 524.194
R108 VSS.n8 VSS.t21 524.194
R109 VSS.n16 VSS.t18 524.194
R110 VSS.n4 VSS.t4 523.069
R111 VSS.t25 VSS.n2 513.159
R112 VSS.n24 VSS.t17 6.65541
R113 VSS.n30 VSS.t14 6.65541
R114 VSS.n36 VSS.t9 6.65541
R115 VSS.n42 VSS.t3 6.65541
R116 VSS.n10 VSS.t22 6.65541
R117 VSS.n6 VSS.t5 6.65541
R118 VSS.n13 VSS.t1 6.65541
R119 VSS.n18 VSS.t19 6.65541
R120 VSS.n46 VSS.t26 6.65541
R121 VSS.n23 VSS.n22 5.2005
R122 VSS.n29 VSS.n28 5.2005
R123 VSS.n35 VSS.n34 5.2005
R124 VSS.n41 VSS.n40 5.2005
R125 VSS.n9 VSS.n8 5.2005
R126 VSS.n17 VSS.n16 5.2005
R127 VSS.n12 VSS.n11 5.2005
R128 VSS.n5 VSS.n4 5.2005
R129 VSS.n47 VSS.n2 5.2005
R130 VSS.n19 VSS.n13 4.69005
R131 VSS VSS.n45 4.35564
R132 VSS.n25 VSS.n24 3.04452
R133 VSS.n19 VSS.n18 3.04452
R134 VSS.n31 VSS.n30 3.0433
R135 VSS.n37 VSS.n36 3.0433
R136 VSS.n44 VSS.n10 3.0433
R137 VSS.n43 VSS.n42 3.04289
R138 VSS.n45 VSS.n6 3.04289
R139 VSS.n45 VSS.n44 1.55259
R140 VSS.n31 VSS.n25 1.55119
R141 VSS.n25 VSS.n19 1.52708
R142 VSS.n44 VSS.n43 1.52661
R143 VSS.n37 VSS.n31 1.52574
R144 VSS.n43 VSS.n37 1.52273
R145 VSS.n46 VSS 0.216546
R146 VSS.n24 VSS.n23 0.142847
R147 VSS.n30 VSS.n29 0.142847
R148 VSS.n36 VSS.n35 0.142847
R149 VSS.n42 VSS.n41 0.142847
R150 VSS.n10 VSS.n9 0.142847
R151 VSS.n6 VSS.n5 0.142847
R152 VSS.n13 VSS.n12 0.142847
R153 VSS.n18 VSS.n17 0.142847
R154 VSS.n47 VSS.n46 0.142847
R155 VSS.n23 VSS 0.00141837
R156 VSS.n29 VSS 0.00141837
R157 VSS.n35 VSS 0.00141837
R158 VSS.n41 VSS 0.00141837
R159 VSS.n9 VSS 0.00141837
R160 VSS.n5 VSS 0.00141837
R161 VSS.n12 VSS 0.00141837
R162 VSS.n17 VSS 0.00141837
R163 VSS VSS.n47 0.00141837
R164 Ci.n0 Ci.t1 28.2228
R165 Ci.n1 Ci.t0 26.9784
R166 Ci.n1 Ci.t2 14.7248
R167 Ci.n0 Ci.t3 14.4701
R168 Ci Ci.n0 4.53357
R169 Ci Ci.n1 4.18544
R170 QB.n0 QB.t3 28.2228
R171 QB.n0 QB.t4 14.4701
R172 QB.n5 QB.n2 6.8765
R173 QB QB.n0 4.52271
R174 QB.n4 QB.t1 3.6405
R175 QB.n4 QB.n3 3.6405
R176 QB.n5 QB.n4 3.08447
R177 QB.n1 QB 2.25992
R178 QB QB.n1 0.725894
R179 QB QB.n5 0.17463
R180 Q.n0 Q.t3 28.2228
R181 Q.n0 Q.t4 14.4701
R182 Q.n5 Q.n2 6.8765
R183 Q Q.n0 4.53357
R184 Q.n4 Q.t0 3.6405
R185 Q.n4 Q.n3 3.6405
R186 Q.n5 Q.n4 3.08447
R187 Q.n1 Q 2.2656
R188 Q Q.n1 0.340471
R189 Q Q.n5 0.17463
R190 Ri-1.n0 Ri-1.t0 28.2228
R191 Ri-1.n1 Ri-1.t3 26.9784
R192 Ri-1.n1 Ri-1.t2 14.7248
R193 Ri-1.n0 Ri-1.t1 14.4701
R194 Ri-1 Ri-1.n0 4.53357
R195 Ri-1 Ri-1.n1 4.18544
R196 Ri.n0 Ri.t0 28.2228
R197 Ri.n1 Ri.t3 26.9784
R198 Ri.n1 Ri.t1 14.7248
R199 Ri.n0 Ri.t2 14.4701
R200 Ri Ri.n0 4.53357
R201 Ri Ri.n1 4.18544
C0 a_305_6005# NAND_13.B 0.00521f
C1 a_305_165# QB 0.0419f
C2 a_305_6981# NAND_13.A 3.37e-19
C3 NAND_1.B NAND_13.A 0.0045f
C4 QB Ci 0.00223f
C5 a_305_165# Q 0.0812f
C6 NAND_12.B NAND_9.B 0.618f
C7 a_305_1140# NAND_3.B 0.0442f
C8 NAND_12.B NAND_12.A 0.625f
C9 Ci Q 1.17e-19
C10 a_305_3086# QB 5.71e-20
C11 VDD NAND_13.A 0.425f
C12 NAND_9.B NAND_12.A 0.0342f
C13 a_305_4056# Ri 0.0852f
C14 VDD QB 0.428f
C15 a_305_5030# Ri 5.72e-20
C16 NAND_12.B Ci 0.237f
C17 VDD Q 0.48f
C18 a_305_6005# NAND_13.A 0.0857f
C19 QB NAND_3.B 0.155f
C20 a_305_5030# NAND_13.B 2.42e-19
C21 NAND_1.B a_305_7966# 0.0455f
C22 NAND_12.B a_305_3086# 0.0419f
C23 NAND_9.B Ci 0.0159f
C24 NAND_13.B NAND_13.A 0.31f
C25 NAND_12.A Ci 2.21e-20
C26 NAND_3.B Q 0.785f
C27 NAND_9.B NAND_1.B 1.76e-19
C28 VDD a_305_7966# 4.39e-19
C29 NAND_12.B VDD 0.575f
C30 NAND_9.B a_305_3086# 0.00221f
C31 NAND_9.B VDD 1.07f
C32 VDD NAND_12.A 0.459f
C33 a_305_7966# Ri-1 0.0852f
C34 a_305_6005# NAND_12.B 4.92e-19
C35 a_305_1140# QB 0.0033f
C36 NAND_12.B Ri 0.0173f
C37 a_305_5030# NAND_13.A 0.0419f
C38 NAND_9.B NAND_3.B 0.242f
C39 NAND_1.B a_305_6981# 0.0864f
C40 a_305_3086# Ci 0.0852f
C41 a_305_1140# Q 2.69e-19
C42 a_305_6005# NAND_9.B 0.0419f
C43 NAND_12.B NAND_13.B 0.0374f
C44 NAND_9.B Ri 0.00203f
C45 a_305_6005# NAND_12.A 3.42e-19
C46 NAND_12.A Ri 0.241f
C47 VDD Ci 0.369f
C48 NAND_9.B NAND_13.B 0.0708f
C49 a_305_165# NAND_3.B 0.00517f
C50 NAND_12.A NAND_13.B 0.00164f
C51 NAND_1.B VDD 0.784f
C52 NAND_12.B a_305_4056# 0.00207f
C53 Ci Ri 0.0048f
C54 QB Q 0.806f
C55 NAND_1.B Ri-1 0.256f
C56 NAND_9.B a_305_1140# 0.0855f
C57 QB a_305_2111# 0.0816f
C58 NAND_12.B a_305_5030# 0.00994f
C59 NAND_9.B a_305_4056# 3.08e-19
C60 NAND_12.B NAND_13.A 0.0793f
C61 NAND_13.B a_305_6981# 0.0455f
C62 NAND_12.A a_305_4056# 0.0421f
C63 a_305_2111# Q 0.0432f
C64 VDD NAND_3.B 0.609f
C65 NAND_9.B a_305_5030# 9.56e-21
C66 VDD Ri-1 0.373f
C67 NAND_1.B NAND_13.B 0.354f
C68 NAND_12.A a_305_5030# 0.0868f
C69 VDD Ri 0.369f
C70 NAND_9.B NAND_13.A 0.494f
C71 NAND_12.A NAND_13.A 0.255f
C72 NAND_12.B Q 0.00934f
C73 VDD NAND_13.B 0.631f
C74 NAND_9.B QB 0.769f
C75 a_305_4056# Ci 5.77e-20
C76 NAND_9.B Q 0.151f
C77 NAND_9.B a_305_2111# 0.00687f
C78 NAND_13.B Ri-1 1.14e-19
C79 a_305_165# VSS 0.0989f
C80 a_305_1140# VSS 0.0983f
C81 NAND_3.B VSS 0.717f
C82 a_305_2111# VSS 0.0983f
C83 Q VSS 1.36f
C84 QB VSS 1.7f
C85 a_305_3086# VSS 0.0989f
C86 Ci VSS 0.605f
C87 a_305_4056# VSS 0.0989f
C88 Ri VSS 0.605f
C89 a_305_5030# VSS 0.0983f
C90 NAND_12.A VSS 0.705f
C91 NAND_12.B VSS 0.961f
C92 a_305_6005# VSS 0.0989f
C93 NAND_9.B VSS 2.51f
C94 NAND_13.A VSS 0.795f
C95 a_305_6981# VSS 0.0989f
C96 NAND_13.B VSS 0.827f
C97 a_305_7966# VSS 0.0983f
C98 NAND_1.B VSS 1.26f
C99 Ri-1 VSS 0.602f
C100 VDD VSS 20.1f
.ends

