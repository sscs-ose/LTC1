magic
tech gf180mcuC
magscale 1 10
timestamp 1693455138
<< error_s >>
rect -24043 -23291 -23831 -23281
rect -3429 -23291 -3217 -23281
<< metal1 >>
rect -22857 -43714 -22497 -43673
rect -22857 -43854 -22794 -43714
rect -22565 -43854 -22497 -43714
rect -22857 -43908 -22497 -43854
<< via1 >>
rect -22794 -43854 -22565 -43714
<< metal2 >>
rect -22857 -43714 -22497 -43673
rect -22857 -43854 -22794 -43714
rect -22565 -43854 -22497 -43714
rect -22857 -43908 -22497 -43854
<< via2 >>
rect -22794 -43854 -22565 -43714
<< metal3 >>
rect -22857 -43714 -22497 -43673
rect -22857 -43854 -22794 -43714
rect -22565 -43854 -22497 -43714
rect -22857 -43908 -22497 -43854
<< via3 >>
rect -22794 -43854 -22565 -43714
<< metal4 >>
rect -22751 -43673 -22631 -43411
rect -22857 -43714 -22497 -43673
rect -22857 -43854 -22794 -43714
rect -22565 -43854 -22497 -43714
rect -22857 -43908 -22497 -43854
<< metal5 >>
rect -24005 -2735 -23915 -2345
rect -24457 -2825 -23338 -2735
rect -24457 -3133 -24367 -2825
rect -23428 -3136 -23338 -2825
rect -25719 -23519 -25384 -22927
rect -23981 -23192 -23893 -23114
rect -3367 -23192 -3279 -23114
rect -23981 -23280 -3279 -23192
rect -23981 -23348 -23893 -23280
rect -3367 -23348 -3279 -23280
rect -24561 -43659 -24408 -43330
rect -23422 -43659 -23269 -43331
rect -24561 -43812 -23269 -43659
use mim_2p0fF_Q6YL6H  mim_2p0fF_Q6YL6H_0
timestamp 1693455138
transform 1 0 -23764 0 1 -23231
box -20547 -20300 20547 20300
<< labels >>
flabel via3 -22691 -43785 -22691 -43785 0 FreeSans 800 0 0 0 N
port 1 nsew
<< end >>
