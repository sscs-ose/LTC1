magic
tech gf180mcuC
magscale 1 10
timestamp 1691496637
<< nwell >>
rect 75 8206 639 8716
rect 75 7221 639 7731
rect 75 6245 639 6755
rect 75 5270 639 5780
rect 75 4296 639 4806
rect 75 3326 639 3836
rect 75 2351 639 2861
rect 75 1380 639 1890
rect 75 405 639 915
<< pwell >>
rect 366 8178 426 8179
rect 366 8134 429 8178
rect 137 7898 577 8134
rect 366 7193 426 7194
rect 366 7149 429 7193
rect 137 6913 577 7149
rect 366 6217 426 6218
rect 366 6173 429 6217
rect 137 5937 577 6173
rect 366 5242 426 5243
rect 366 5198 429 5242
rect 137 4962 577 5198
rect 366 4268 426 4269
rect 366 4224 429 4268
rect 137 3988 577 4224
rect 366 3298 426 3299
rect 366 3254 429 3298
rect 137 3018 577 3254
rect 366 2323 426 2324
rect 366 2279 429 2323
rect 137 2043 577 2279
rect 366 1352 426 1353
rect 366 1308 429 1352
rect 137 1072 577 1308
rect 366 377 426 378
rect 366 333 429 377
rect 137 97 577 333
<< nmos >>
rect 249 7966 305 8066
rect 409 7966 465 8066
rect 249 6981 305 7081
rect 409 6981 465 7081
rect 249 6005 305 6105
rect 409 6005 465 6105
rect 249 5030 305 5130
rect 409 5030 465 5130
rect 249 4056 305 4156
rect 409 4056 465 4156
rect 249 3086 305 3186
rect 409 3086 465 3186
rect 249 2111 305 2211
rect 409 2111 465 2211
rect 249 1140 305 1240
rect 409 1140 465 1240
rect 249 165 305 265
rect 409 165 465 265
<< pmos >>
rect 249 8336 305 8436
rect 409 8336 465 8436
rect 249 7351 305 7451
rect 409 7351 465 7451
rect 249 6375 305 6475
rect 409 6375 465 6475
rect 249 5400 305 5500
rect 409 5400 465 5500
rect 249 4426 305 4526
rect 409 4426 465 4526
rect 249 3456 305 3556
rect 409 3456 465 3556
rect 249 2481 305 2581
rect 409 2481 465 2581
rect 249 1510 305 1610
rect 409 1510 465 1610
rect 249 535 305 635
rect 409 535 465 635
<< ndiff >>
rect 161 8053 249 8066
rect 161 7979 174 8053
rect 220 7979 249 8053
rect 161 7966 249 7979
rect 305 8053 409 8066
rect 305 7979 334 8053
rect 380 7979 409 8053
rect 305 7966 409 7979
rect 465 8053 553 8066
rect 465 7979 494 8053
rect 540 7979 553 8053
rect 465 7966 553 7979
rect 161 7068 249 7081
rect 161 6994 174 7068
rect 220 6994 249 7068
rect 161 6981 249 6994
rect 305 7068 409 7081
rect 305 6994 334 7068
rect 380 6994 409 7068
rect 305 6981 409 6994
rect 465 7068 553 7081
rect 465 6994 494 7068
rect 540 6994 553 7068
rect 465 6981 553 6994
rect 161 6092 249 6105
rect 161 6018 174 6092
rect 220 6018 249 6092
rect 161 6005 249 6018
rect 305 6092 409 6105
rect 305 6018 334 6092
rect 380 6018 409 6092
rect 305 6005 409 6018
rect 465 6092 553 6105
rect 465 6018 494 6092
rect 540 6018 553 6092
rect 465 6005 553 6018
rect 161 5117 249 5130
rect 161 5043 174 5117
rect 220 5043 249 5117
rect 161 5030 249 5043
rect 305 5117 409 5130
rect 305 5043 334 5117
rect 380 5043 409 5117
rect 305 5030 409 5043
rect 465 5117 553 5130
rect 465 5043 494 5117
rect 540 5043 553 5117
rect 465 5030 553 5043
rect 161 4143 249 4156
rect 161 4069 174 4143
rect 220 4069 249 4143
rect 161 4056 249 4069
rect 305 4143 409 4156
rect 305 4069 334 4143
rect 380 4069 409 4143
rect 305 4056 409 4069
rect 465 4143 553 4156
rect 465 4069 494 4143
rect 540 4069 553 4143
rect 465 4056 553 4069
rect 161 3173 249 3186
rect 161 3099 174 3173
rect 220 3099 249 3173
rect 161 3086 249 3099
rect 305 3173 409 3186
rect 305 3099 334 3173
rect 380 3099 409 3173
rect 305 3086 409 3099
rect 465 3173 553 3186
rect 465 3099 494 3173
rect 540 3099 553 3173
rect 465 3086 553 3099
rect 161 2198 249 2211
rect 161 2124 174 2198
rect 220 2124 249 2198
rect 161 2111 249 2124
rect 305 2198 409 2211
rect 305 2124 334 2198
rect 380 2124 409 2198
rect 305 2111 409 2124
rect 465 2198 553 2211
rect 465 2124 494 2198
rect 540 2124 553 2198
rect 465 2111 553 2124
rect 161 1227 249 1240
rect 161 1153 174 1227
rect 220 1153 249 1227
rect 161 1140 249 1153
rect 305 1227 409 1240
rect 305 1153 334 1227
rect 380 1153 409 1227
rect 305 1140 409 1153
rect 465 1227 553 1240
rect 465 1153 494 1227
rect 540 1153 553 1227
rect 465 1140 553 1153
rect 161 252 249 265
rect 161 178 174 252
rect 220 178 249 252
rect 161 165 249 178
rect 305 252 409 265
rect 305 178 334 252
rect 380 178 409 252
rect 305 165 409 178
rect 465 252 553 265
rect 465 178 494 252
rect 540 178 553 252
rect 465 165 553 178
<< pdiff >>
rect 161 8423 249 8436
rect 161 8349 174 8423
rect 220 8349 249 8423
rect 161 8336 249 8349
rect 305 8423 409 8436
rect 305 8349 334 8423
rect 380 8349 409 8423
rect 305 8336 409 8349
rect 465 8423 553 8436
rect 465 8349 494 8423
rect 540 8349 553 8423
rect 465 8336 553 8349
rect 161 7438 249 7451
rect 161 7364 174 7438
rect 220 7364 249 7438
rect 161 7351 249 7364
rect 305 7438 409 7451
rect 305 7364 334 7438
rect 380 7364 409 7438
rect 305 7351 409 7364
rect 465 7438 553 7451
rect 465 7364 494 7438
rect 540 7364 553 7438
rect 465 7351 553 7364
rect 161 6462 249 6475
rect 161 6388 174 6462
rect 220 6388 249 6462
rect 161 6375 249 6388
rect 305 6462 409 6475
rect 305 6388 334 6462
rect 380 6388 409 6462
rect 305 6375 409 6388
rect 465 6462 553 6475
rect 465 6388 494 6462
rect 540 6388 553 6462
rect 465 6375 553 6388
rect 161 5487 249 5500
rect 161 5413 174 5487
rect 220 5413 249 5487
rect 161 5400 249 5413
rect 305 5487 409 5500
rect 305 5413 334 5487
rect 380 5413 409 5487
rect 305 5400 409 5413
rect 465 5487 553 5500
rect 465 5413 494 5487
rect 540 5413 553 5487
rect 465 5400 553 5413
rect 161 4513 249 4526
rect 161 4439 174 4513
rect 220 4439 249 4513
rect 161 4426 249 4439
rect 305 4513 409 4526
rect 305 4439 334 4513
rect 380 4439 409 4513
rect 305 4426 409 4439
rect 465 4513 553 4526
rect 465 4439 494 4513
rect 540 4439 553 4513
rect 465 4426 553 4439
rect 161 3543 249 3556
rect 161 3469 174 3543
rect 220 3469 249 3543
rect 161 3456 249 3469
rect 305 3543 409 3556
rect 305 3469 334 3543
rect 380 3469 409 3543
rect 305 3456 409 3469
rect 465 3543 553 3556
rect 465 3469 494 3543
rect 540 3469 553 3543
rect 465 3456 553 3469
rect 161 2568 249 2581
rect 161 2494 174 2568
rect 220 2494 249 2568
rect 161 2481 249 2494
rect 305 2568 409 2581
rect 305 2494 334 2568
rect 380 2494 409 2568
rect 305 2481 409 2494
rect 465 2568 553 2581
rect 465 2494 494 2568
rect 540 2494 553 2568
rect 465 2481 553 2494
rect 161 1597 249 1610
rect 161 1523 174 1597
rect 220 1523 249 1597
rect 161 1510 249 1523
rect 305 1597 409 1610
rect 305 1523 334 1597
rect 380 1523 409 1597
rect 305 1510 409 1523
rect 465 1597 553 1610
rect 465 1523 494 1597
rect 540 1523 553 1597
rect 465 1510 553 1523
rect 161 622 249 635
rect 161 548 174 622
rect 220 548 249 622
rect 161 535 249 548
rect 305 622 409 635
rect 305 548 334 622
rect 380 548 409 622
rect 305 535 409 548
rect 465 622 553 635
rect 465 548 494 622
rect 540 548 553 622
rect 465 535 553 548
<< ndiffc >>
rect 174 7979 220 8053
rect 334 7979 380 8053
rect 494 7979 540 8053
rect 174 6994 220 7068
rect 334 6994 380 7068
rect 494 6994 540 7068
rect 174 6018 220 6092
rect 334 6018 380 6092
rect 494 6018 540 6092
rect 174 5043 220 5117
rect 334 5043 380 5117
rect 494 5043 540 5117
rect 174 4069 220 4143
rect 334 4069 380 4143
rect 494 4069 540 4143
rect 174 3099 220 3173
rect 334 3099 380 3173
rect 494 3099 540 3173
rect 174 2124 220 2198
rect 334 2124 380 2198
rect 494 2124 540 2198
rect 174 1153 220 1227
rect 334 1153 380 1227
rect 494 1153 540 1227
rect 174 178 220 252
rect 334 178 380 252
rect 494 178 540 252
<< pdiffc >>
rect 174 8349 220 8423
rect 334 8349 380 8423
rect 494 8349 540 8423
rect 174 7364 220 7438
rect 334 7364 380 7438
rect 494 7364 540 7438
rect 174 6388 220 6462
rect 334 6388 380 6462
rect 494 6388 540 6462
rect 174 5413 220 5487
rect 334 5413 380 5487
rect 494 5413 540 5487
rect 174 4439 220 4513
rect 334 4439 380 4513
rect 494 4439 540 4513
rect 174 3469 220 3543
rect 334 3469 380 3543
rect 494 3469 540 3543
rect 174 2494 220 2568
rect 334 2494 380 2568
rect 494 2494 540 2568
rect 174 1523 220 1597
rect 334 1523 380 1597
rect 494 1523 540 1597
rect 174 548 220 622
rect 334 548 380 622
rect 494 548 540 622
<< psubdiff >>
rect 87 7872 641 7888
rect 87 7824 118 7872
rect 587 7824 641 7872
rect 87 7806 641 7824
rect 87 6887 641 6903
rect 87 6839 118 6887
rect 587 6839 641 6887
rect 87 6821 641 6839
rect 87 5911 641 5927
rect 87 5863 118 5911
rect 587 5863 641 5911
rect 87 5845 641 5863
rect 87 4936 641 4952
rect 87 4888 118 4936
rect 587 4888 641 4936
rect 87 4870 641 4888
rect 87 3962 641 3978
rect 87 3914 118 3962
rect 587 3914 641 3962
rect 87 3896 641 3914
rect 87 2992 641 3008
rect 87 2944 118 2992
rect 587 2944 641 2992
rect 87 2926 641 2944
rect 87 2017 641 2033
rect 87 1969 118 2017
rect 587 1969 641 2017
rect 87 1951 641 1969
rect 87 1046 641 1062
rect 87 998 118 1046
rect 587 998 641 1046
rect 87 980 641 998
rect 87 71 641 87
rect 87 23 118 71
rect 587 23 641 71
rect 87 5 641 23
<< nsubdiff >>
rect 153 8670 559 8690
rect 153 8614 190 8670
rect 502 8614 559 8670
rect 153 8593 559 8614
rect 153 7685 559 7705
rect 153 7629 190 7685
rect 502 7629 559 7685
rect 153 7608 559 7629
rect 153 6709 559 6729
rect 153 6653 190 6709
rect 502 6653 559 6709
rect 153 6632 559 6653
rect 153 5734 559 5754
rect 153 5678 190 5734
rect 502 5678 559 5734
rect 153 5657 559 5678
rect 153 4760 559 4780
rect 153 4704 190 4760
rect 502 4704 559 4760
rect 153 4683 559 4704
rect 153 3790 559 3810
rect 153 3734 190 3790
rect 502 3734 559 3790
rect 153 3713 559 3734
rect 153 2815 559 2835
rect 153 2759 190 2815
rect 502 2759 559 2815
rect 153 2738 559 2759
rect 153 1844 559 1864
rect 153 1788 190 1844
rect 502 1788 559 1844
rect 153 1767 559 1788
rect 153 869 559 889
rect 153 813 190 869
rect 502 813 559 869
rect 153 792 559 813
<< psubdiffcont >>
rect 118 7824 587 7872
rect 118 6839 587 6887
rect 118 5863 587 5911
rect 118 4888 587 4936
rect 118 3914 587 3962
rect 118 2944 587 2992
rect 118 1969 587 2017
rect 118 998 587 1046
rect 118 23 587 71
<< nsubdiffcont >>
rect 190 8614 502 8670
rect 190 7629 502 7685
rect 190 6653 502 6709
rect 190 5678 502 5734
rect 190 4704 502 4760
rect 190 3734 502 3790
rect 190 2759 502 2815
rect 190 1788 502 1844
rect 190 813 502 869
<< polysilicon >>
rect 249 8436 305 8480
rect 409 8436 465 8480
rect 249 8292 305 8336
rect 175 8278 305 8292
rect 175 8219 189 8278
rect 252 8219 305 8278
rect 175 8204 305 8219
rect 249 8066 305 8204
rect 409 8191 465 8336
rect 353 8178 465 8191
rect 353 8119 366 8178
rect 429 8119 465 8178
rect 353 8106 465 8119
rect 409 8066 465 8106
rect 249 7922 305 7966
rect 409 7922 465 7966
rect 249 7451 305 7495
rect 409 7451 465 7495
rect 249 7307 305 7351
rect 175 7293 305 7307
rect 175 7234 189 7293
rect 252 7234 305 7293
rect 175 7219 305 7234
rect 249 7081 305 7219
rect 409 7206 465 7351
rect 353 7193 465 7206
rect 353 7134 366 7193
rect 429 7134 465 7193
rect 353 7121 465 7134
rect 409 7081 465 7121
rect 249 6937 305 6981
rect 409 6937 465 6981
rect 249 6475 305 6519
rect 409 6475 465 6519
rect 249 6331 305 6375
rect 175 6317 305 6331
rect 175 6258 189 6317
rect 252 6258 305 6317
rect 175 6243 305 6258
rect 249 6105 305 6243
rect 409 6230 465 6375
rect 353 6217 465 6230
rect 353 6158 366 6217
rect 429 6158 465 6217
rect 353 6145 465 6158
rect 409 6105 465 6145
rect 249 5961 305 6005
rect 409 5961 465 6005
rect 249 5500 305 5544
rect 409 5500 465 5544
rect 249 5356 305 5400
rect 175 5342 305 5356
rect 175 5283 189 5342
rect 252 5283 305 5342
rect 175 5268 305 5283
rect 249 5130 305 5268
rect 409 5255 465 5400
rect 353 5242 465 5255
rect 353 5183 366 5242
rect 429 5183 465 5242
rect 353 5170 465 5183
rect 409 5130 465 5170
rect 249 4986 305 5030
rect 409 4986 465 5030
rect 249 4526 305 4570
rect 409 4526 465 4570
rect 249 4382 305 4426
rect 175 4368 305 4382
rect 175 4309 189 4368
rect 252 4309 305 4368
rect 175 4294 305 4309
rect 249 4156 305 4294
rect 409 4281 465 4426
rect 353 4268 465 4281
rect 353 4209 366 4268
rect 429 4209 465 4268
rect 353 4196 465 4209
rect 409 4156 465 4196
rect 249 4012 305 4056
rect 409 4012 465 4056
rect 249 3556 305 3600
rect 409 3556 465 3600
rect 249 3412 305 3456
rect 175 3398 305 3412
rect 175 3339 189 3398
rect 252 3339 305 3398
rect 175 3324 305 3339
rect 249 3186 305 3324
rect 409 3311 465 3456
rect 353 3298 465 3311
rect 353 3239 366 3298
rect 429 3239 465 3298
rect 353 3226 465 3239
rect 409 3186 465 3226
rect 249 3042 305 3086
rect 409 3042 465 3086
rect 249 2581 305 2625
rect 409 2581 465 2625
rect 249 2437 305 2481
rect 175 2423 305 2437
rect 175 2364 189 2423
rect 252 2364 305 2423
rect 175 2349 305 2364
rect 249 2211 305 2349
rect 409 2336 465 2481
rect 353 2323 465 2336
rect 353 2264 366 2323
rect 429 2264 465 2323
rect 353 2251 465 2264
rect 409 2211 465 2251
rect 249 2067 305 2111
rect 409 2067 465 2111
rect 249 1610 305 1654
rect 409 1610 465 1654
rect 249 1466 305 1510
rect 175 1452 305 1466
rect 175 1393 189 1452
rect 252 1393 305 1452
rect 175 1378 305 1393
rect 249 1240 305 1378
rect 409 1365 465 1510
rect 353 1352 465 1365
rect 353 1293 366 1352
rect 429 1293 465 1352
rect 353 1280 465 1293
rect 409 1240 465 1280
rect 249 1096 305 1140
rect 409 1096 465 1140
rect 249 635 305 679
rect 409 635 465 679
rect 249 491 305 535
rect 175 477 305 491
rect 175 418 189 477
rect 252 418 305 477
rect 175 403 305 418
rect 249 265 305 403
rect 409 390 465 535
rect 353 377 465 390
rect 353 318 366 377
rect 429 318 465 377
rect 353 305 465 318
rect 409 265 465 305
rect 249 121 305 165
rect 409 121 465 165
<< polycontact >>
rect 189 8219 252 8278
rect 366 8119 429 8178
rect 189 7234 252 7293
rect 366 7134 429 7193
rect 189 6258 252 6317
rect 366 6158 429 6217
rect 189 5283 252 5342
rect 366 5183 429 5242
rect 189 4309 252 4368
rect 366 4209 429 4268
rect 189 3339 252 3398
rect 366 3239 429 3298
rect 189 2364 252 2423
rect 366 2264 429 2323
rect 189 1393 252 1452
rect 366 1293 429 1352
rect 189 418 252 477
rect 366 318 429 377
<< metal1 >>
rect -590 8663 -510 8677
rect 75 8670 639 8716
rect 75 8663 190 8670
rect -590 8662 190 8663
rect -590 8608 -576 8662
rect -522 8614 190 8662
rect 502 8614 639 8670
rect -522 8608 639 8614
rect -590 8607 639 8608
rect -590 8598 -510 8607
rect 75 8566 639 8607
rect 171 8423 222 8566
rect 171 8349 174 8423
rect 220 8349 222 8423
rect 171 8347 222 8349
rect 334 8423 380 8434
rect 174 8338 220 8347
rect 334 8296 380 8349
rect 494 8423 540 8566
rect 494 8338 540 8349
rect 608 8296 694 8306
rect 334 8292 443 8296
rect 608 8292 624 8296
rect 175 8278 264 8292
rect 175 8250 189 8278
rect 74 8219 189 8250
rect 252 8219 264 8278
rect 334 8250 624 8292
rect 410 8246 624 8250
rect 74 8204 264 8219
rect 76 8156 122 8204
rect 355 8178 440 8189
rect 355 8156 366 8178
rect 76 8119 366 8156
rect 429 8119 440 8178
rect 76 8110 440 8119
rect 174 8053 220 8064
rect 334 8063 380 8064
rect 174 7899 220 7979
rect 321 8053 388 8063
rect 321 7979 334 8053
rect 380 7979 388 8053
rect 321 7965 388 7979
rect 494 8053 540 8246
rect 608 8242 624 8246
rect 678 8242 694 8296
rect 608 8231 694 8242
rect 494 7968 540 7979
rect -409 7870 -330 7883
rect 51 7872 667 7899
rect 51 7870 118 7872
rect -409 7814 -397 7870
rect -341 7824 118 7870
rect 587 7824 667 7872
rect -341 7814 667 7824
rect -409 7808 -330 7814
rect 51 7801 667 7814
rect -591 7687 -511 7699
rect 75 7687 639 7731
rect -591 7631 -577 7687
rect -521 7685 639 7687
rect -521 7631 190 7685
rect -591 7620 -511 7631
rect 75 7629 190 7631
rect 502 7629 639 7685
rect 75 7581 639 7629
rect 171 7438 222 7581
rect 171 7364 174 7438
rect 220 7364 222 7438
rect 171 7362 222 7364
rect 334 7438 380 7449
rect 174 7353 220 7362
rect 334 7311 380 7364
rect 494 7438 540 7581
rect 494 7353 540 7364
rect 600 7311 680 7323
rect 334 7307 443 7311
rect 600 7307 613 7311
rect 175 7293 264 7307
rect 49 7265 127 7267
rect 175 7265 189 7293
rect 49 7263 189 7265
rect 49 7207 61 7263
rect 117 7234 189 7263
rect 252 7234 264 7293
rect 334 7265 613 7307
rect 410 7261 613 7265
rect 117 7219 264 7234
rect 117 7207 127 7219
rect 49 7196 127 7207
rect 76 7171 127 7196
rect 355 7193 440 7204
rect 355 7171 366 7193
rect 76 7134 366 7171
rect 429 7134 440 7193
rect 76 7125 440 7134
rect 174 7068 220 7079
rect 334 7078 380 7079
rect 174 6914 220 6994
rect 321 7068 388 7078
rect 321 6994 334 7068
rect 380 6994 388 7068
rect 321 6980 388 6994
rect 494 7068 540 7261
rect 600 7257 613 7261
rect 667 7257 680 7311
rect 600 7252 680 7257
rect 494 6983 540 6994
rect -407 6898 -328 6909
rect 51 6898 667 6914
rect -407 6842 -397 6898
rect -341 6887 667 6898
rect -341 6842 118 6887
rect -407 6834 -328 6842
rect 51 6839 118 6842
rect 587 6839 667 6887
rect 51 6816 667 6839
rect -592 6716 -512 6728
rect 75 6716 639 6755
rect -592 6660 -577 6716
rect -521 6709 639 6716
rect -521 6660 190 6709
rect -592 6649 -512 6660
rect 75 6653 190 6660
rect 502 6653 639 6709
rect 75 6605 639 6653
rect 171 6462 222 6605
rect 171 6388 174 6462
rect 220 6388 222 6462
rect 171 6386 222 6388
rect 334 6462 380 6473
rect 174 6377 220 6386
rect 334 6335 380 6388
rect 494 6462 540 6605
rect 494 6377 540 6388
rect 873 6335 953 6347
rect 334 6331 443 6335
rect 873 6331 886 6335
rect 43 6312 127 6320
rect 43 6256 55 6312
rect 111 6289 127 6312
rect 175 6317 264 6331
rect 175 6289 189 6317
rect 111 6258 189 6289
rect 252 6258 264 6317
rect 334 6289 886 6331
rect 410 6285 886 6289
rect 111 6256 264 6258
rect 43 6243 264 6256
rect 352 6217 440 6228
rect 352 6216 366 6217
rect 352 6195 365 6216
rect 76 6160 365 6195
rect 76 6158 366 6160
rect 429 6158 440 6217
rect 76 6149 440 6158
rect 174 6092 220 6103
rect 334 6102 380 6103
rect 174 5938 220 6018
rect 321 6092 388 6102
rect 321 6018 334 6092
rect 380 6018 388 6092
rect 321 6004 388 6018
rect 494 6092 540 6285
rect 873 6281 886 6285
rect 940 6281 953 6335
rect 873 6277 953 6281
rect 494 6007 540 6018
rect -408 5911 -329 5920
rect 51 5911 667 5938
rect -408 5855 -397 5911
rect -341 5863 118 5911
rect 587 5863 667 5911
rect -341 5855 667 5863
rect -408 5845 -329 5855
rect 51 5840 667 5855
rect -589 5740 -509 5752
rect 75 5740 639 5780
rect -589 5684 -577 5740
rect -521 5734 639 5740
rect -521 5684 190 5734
rect -589 5673 -509 5684
rect 75 5678 190 5684
rect 502 5678 639 5734
rect 75 5630 639 5678
rect 171 5487 222 5630
rect 171 5413 174 5487
rect 220 5413 222 5487
rect 171 5411 222 5413
rect 334 5487 380 5498
rect 174 5402 220 5411
rect 334 5360 380 5413
rect 494 5487 540 5630
rect 494 5402 540 5413
rect 692 5360 780 5373
rect 334 5356 443 5360
rect 692 5356 703 5360
rect 23 5333 103 5344
rect 23 5277 37 5333
rect 93 5314 103 5333
rect 175 5342 264 5356
rect 175 5314 189 5342
rect 93 5283 189 5314
rect 252 5283 264 5342
rect 334 5314 703 5356
rect 410 5310 703 5314
rect 93 5277 264 5283
rect 23 5269 264 5277
rect 74 5268 264 5269
rect 351 5253 439 5254
rect 351 5244 440 5253
rect 351 5220 362 5244
rect 418 5242 440 5244
rect 76 5188 362 5220
rect 76 5183 366 5188
rect 429 5183 440 5242
rect 76 5174 440 5183
rect 174 5117 220 5128
rect 334 5127 380 5128
rect 174 4963 220 5043
rect 321 5117 388 5127
rect 321 5043 334 5117
rect 380 5043 388 5117
rect 321 5029 388 5043
rect 494 5117 540 5310
rect 692 5306 703 5310
rect 757 5306 780 5360
rect 692 5297 780 5306
rect 494 5032 540 5043
rect -407 4939 -328 4950
rect 51 4939 667 4963
rect -407 4883 -397 4939
rect -341 4936 667 4939
rect -341 4888 118 4936
rect 587 4888 667 4936
rect -341 4883 667 4888
rect -407 4875 -328 4883
rect 51 4865 667 4883
rect 75 4760 639 4806
rect -588 4740 -508 4752
rect 75 4740 190 4760
rect -588 4684 -577 4740
rect -521 4704 190 4740
rect 502 4704 639 4760
rect -521 4684 639 4704
rect -588 4673 -508 4684
rect 75 4656 639 4684
rect 171 4513 222 4656
rect 171 4439 174 4513
rect 220 4439 222 4513
rect 171 4437 222 4439
rect 334 4513 380 4524
rect 174 4428 220 4437
rect 334 4386 380 4439
rect 494 4513 540 4656
rect 494 4428 540 4439
rect 574 4386 662 4396
rect 334 4382 443 4386
rect 574 4382 588 4386
rect 175 4368 264 4382
rect 175 4340 189 4368
rect 74 4309 189 4340
rect 252 4309 264 4368
rect 334 4340 588 4382
rect 410 4336 588 4340
rect 74 4294 264 4309
rect 494 4332 588 4336
rect 642 4332 662 4386
rect 494 4324 662 4332
rect 76 4246 122 4294
rect 355 4268 440 4279
rect 355 4246 366 4268
rect 76 4209 366 4246
rect 429 4209 440 4268
rect 76 4200 440 4209
rect 174 4143 220 4154
rect 334 4153 380 4154
rect 174 3989 220 4069
rect 321 4143 388 4153
rect 321 4069 334 4143
rect 380 4069 388 4143
rect 321 4055 388 4069
rect 494 4143 540 4324
rect 494 4058 540 4069
rect -408 3970 -329 3981
rect 51 3970 667 3989
rect -408 3914 -397 3970
rect -341 3962 667 3970
rect -341 3914 118 3962
rect 587 3914 667 3962
rect -408 3906 -329 3914
rect 51 3891 667 3914
rect 75 3790 639 3836
rect -588 3773 -508 3786
rect 75 3773 190 3790
rect -588 3717 -577 3773
rect -521 3734 190 3773
rect 502 3734 639 3790
rect -521 3717 639 3734
rect -588 3707 -508 3717
rect 75 3686 639 3717
rect 171 3543 222 3686
rect 171 3469 174 3543
rect 220 3469 222 3543
rect 171 3467 222 3469
rect 334 3543 380 3554
rect 174 3458 220 3467
rect 334 3416 380 3469
rect 494 3543 540 3686
rect 494 3458 540 3469
rect 735 3416 815 3427
rect 334 3412 443 3416
rect 735 3412 745 3416
rect 175 3398 264 3412
rect 175 3370 189 3398
rect 74 3339 189 3370
rect 252 3339 264 3398
rect 334 3370 745 3412
rect 410 3366 745 3370
rect 74 3324 264 3339
rect 76 3276 122 3324
rect 355 3298 440 3309
rect 355 3276 366 3298
rect 76 3239 366 3276
rect 429 3239 440 3298
rect 76 3230 440 3239
rect 174 3173 220 3184
rect 334 3183 380 3184
rect 174 3019 220 3099
rect 321 3173 388 3183
rect 321 3099 334 3173
rect 380 3099 388 3173
rect 321 3085 388 3099
rect 494 3173 540 3366
rect 735 3362 745 3366
rect 799 3362 815 3416
rect 735 3352 815 3362
rect 494 3088 540 3099
rect -408 3000 -329 3008
rect 51 3000 667 3019
rect -408 2944 -397 3000
rect -341 2992 667 3000
rect -341 2944 118 2992
rect 587 2944 667 2992
rect -408 2933 -329 2944
rect 51 2921 667 2944
rect -588 2839 -508 2852
rect 75 2839 639 2861
rect -588 2783 -577 2839
rect -521 2815 639 2839
rect -521 2783 190 2815
rect -588 2773 -508 2783
rect 75 2759 190 2783
rect 502 2759 639 2815
rect 75 2711 639 2759
rect 171 2568 222 2711
rect 171 2494 174 2568
rect 220 2494 222 2568
rect 171 2492 222 2494
rect 334 2568 380 2579
rect 174 2483 220 2492
rect 334 2441 380 2494
rect 494 2568 540 2711
rect 494 2483 540 2494
rect 761 2441 848 2457
rect 334 2437 443 2441
rect 761 2437 776 2441
rect 175 2423 264 2437
rect -63 2406 16 2417
rect -63 2350 -52 2406
rect 4 2395 16 2406
rect 175 2395 189 2423
rect 4 2364 189 2395
rect 252 2364 264 2423
rect 334 2395 776 2437
rect 410 2391 776 2395
rect 4 2350 264 2364
rect -63 2349 264 2350
rect -63 2338 16 2349
rect 355 2323 440 2334
rect 355 2301 366 2323
rect -237 2281 -156 2292
rect -237 2225 -224 2281
rect -168 2274 -156 2281
rect 76 2274 366 2301
rect -168 2264 366 2274
rect 429 2264 440 2323
rect -168 2255 440 2264
rect -168 2228 122 2255
rect -168 2225 -156 2228
rect -237 2218 -156 2225
rect 174 2198 220 2209
rect 334 2208 380 2209
rect 174 2044 220 2124
rect 321 2198 388 2208
rect 321 2124 334 2198
rect 380 2124 388 2198
rect 321 2110 388 2124
rect 494 2198 540 2391
rect 761 2387 776 2391
rect 830 2387 848 2441
rect 761 2381 848 2387
rect 494 2113 540 2124
rect -411 2013 -332 2022
rect 51 2017 667 2044
rect 51 2013 118 2017
rect -411 1957 -397 2013
rect -341 1969 118 2013
rect 587 1969 667 2017
rect -341 1957 667 1969
rect -411 1947 -332 1957
rect 51 1946 667 1957
rect -587 1852 -507 1864
rect 75 1852 639 1890
rect -587 1796 -577 1852
rect -521 1844 639 1852
rect -521 1796 190 1844
rect -587 1785 -507 1796
rect 75 1788 190 1796
rect 502 1788 639 1844
rect 75 1740 639 1788
rect 171 1597 222 1740
rect 171 1523 174 1597
rect 220 1523 222 1597
rect 171 1521 222 1523
rect 334 1597 380 1608
rect 174 1512 220 1521
rect 334 1470 380 1523
rect 494 1597 540 1740
rect 494 1512 540 1523
rect 334 1466 443 1470
rect 175 1452 264 1466
rect 175 1424 189 1452
rect -63 1394 13 1404
rect 74 1394 189 1424
rect -63 1338 -52 1394
rect 4 1393 189 1394
rect 252 1393 264 1452
rect 334 1424 639 1466
rect 410 1420 639 1424
rect 4 1378 264 1393
rect 4 1338 122 1378
rect -63 1328 13 1338
rect 76 1330 122 1338
rect 355 1352 440 1363
rect 355 1330 366 1352
rect 76 1293 366 1330
rect 429 1293 440 1352
rect 76 1284 440 1293
rect 174 1227 220 1238
rect 334 1237 380 1238
rect 174 1073 220 1153
rect 321 1227 388 1237
rect 321 1153 334 1227
rect 380 1153 388 1227
rect 321 1139 388 1153
rect 494 1227 540 1420
rect 587 1212 669 1225
rect 587 1208 600 1212
rect 540 1162 600 1208
rect 587 1158 600 1162
rect 654 1158 669 1212
rect 587 1153 669 1158
rect 494 1142 540 1153
rect -411 1041 -332 1051
rect 51 1046 667 1073
rect 51 1041 118 1046
rect -411 985 -397 1041
rect -341 998 118 1041
rect 587 998 667 1046
rect -341 985 667 998
rect -411 976 -332 985
rect 51 975 667 985
rect -587 876 -507 888
rect 75 876 639 915
rect -587 820 -577 876
rect -521 869 639 876
rect -521 820 190 869
rect -587 809 -507 820
rect 75 813 190 820
rect 502 813 639 869
rect 75 765 639 813
rect 171 622 222 765
rect 171 548 174 622
rect 220 548 222 622
rect 171 546 222 548
rect 334 622 380 633
rect 174 537 220 546
rect 334 495 380 548
rect 494 622 540 765
rect 494 537 540 548
rect 955 495 1033 504
rect 334 491 443 495
rect 955 491 966 495
rect 175 477 264 491
rect 42 464 124 475
rect 42 408 54 464
rect 110 449 124 464
rect 175 449 189 477
rect 110 418 189 449
rect 252 418 264 477
rect 334 449 966 491
rect 410 445 966 449
rect 110 408 264 418
rect 42 403 264 408
rect 355 377 440 388
rect -121 355 -45 357
rect 355 355 366 377
rect -121 346 366 355
rect -121 290 -110 346
rect -54 318 366 346
rect 429 318 440 377
rect -54 309 440 318
rect -54 290 -45 309
rect -121 281 -45 290
rect 174 252 220 263
rect 334 262 380 263
rect 174 98 220 178
rect 321 252 388 262
rect 321 178 334 252
rect 380 178 388 252
rect 321 164 388 178
rect 494 252 540 445
rect 955 441 966 445
rect 1020 441 1033 495
rect 955 430 1033 441
rect 494 167 540 178
rect -408 77 -329 85
rect -408 23 -396 77
rect -342 73 -329 77
rect 51 73 667 98
rect -342 71 667 73
rect -342 27 118 71
rect -342 23 -329 27
rect -408 10 -329 23
rect 51 23 118 27
rect 587 23 667 71
rect 51 0 667 23
<< via1 >>
rect -576 8608 -522 8662
rect 624 8242 678 8296
rect -397 7814 -341 7870
rect -577 7631 -521 7687
rect 61 7207 117 7263
rect 613 7257 667 7311
rect -397 6842 -341 6898
rect -577 6660 -521 6716
rect 55 6256 111 6312
rect 365 6160 366 6216
rect 366 6160 421 6216
rect 886 6281 940 6335
rect -397 5855 -341 5911
rect -577 5684 -521 5740
rect 37 5277 93 5333
rect 362 5242 418 5244
rect 362 5188 366 5242
rect 366 5188 418 5242
rect 703 5306 757 5360
rect -397 4883 -341 4939
rect -577 4684 -521 4740
rect 588 4332 642 4386
rect -397 3914 -341 3970
rect -577 3717 -521 3773
rect 745 3362 799 3416
rect -397 2944 -341 3000
rect -577 2783 -521 2839
rect -52 2350 4 2406
rect -224 2225 -168 2281
rect 776 2387 830 2441
rect -397 1957 -341 2013
rect -577 1796 -521 1852
rect -52 1338 4 1394
rect 600 1158 654 1212
rect -397 985 -341 1041
rect -577 820 -521 876
rect 54 408 110 464
rect -110 290 -54 346
rect 966 441 1020 495
rect -396 23 -342 77
<< metal2 >>
rect -590 8662 -510 8677
rect -590 8608 -576 8662
rect -522 8608 -510 8662
rect -590 8598 -510 8608
rect -577 7699 -521 8598
rect 608 8296 694 8306
rect 608 8242 624 8296
rect 678 8242 694 8296
rect 608 8231 694 8242
rect -409 7870 -330 7883
rect -409 7814 -397 7870
rect -341 7814 -330 7870
rect -409 7808 -330 7814
rect -591 7687 -511 7699
rect -591 7631 -577 7687
rect -521 7631 -511 7687
rect -591 7620 -511 7631
rect -577 6728 -521 7620
rect -397 6909 -341 7808
rect 46 7550 132 7564
rect 623 7558 679 8231
rect 46 7494 61 7550
rect 117 7494 132 7550
rect 46 7489 132 7494
rect 610 7550 696 7558
rect 610 7494 623 7550
rect 679 7494 696 7550
rect 61 7267 117 7489
rect 610 7483 696 7494
rect 600 7311 680 7323
rect 49 7263 127 7267
rect 49 7207 61 7263
rect 117 7207 127 7263
rect 600 7257 613 7311
rect 667 7257 680 7311
rect 600 7252 680 7257
rect 49 7196 127 7207
rect -407 6898 -328 6909
rect -407 6842 -397 6898
rect -341 6842 -328 6898
rect -407 6834 -328 6842
rect -592 6716 -512 6728
rect -592 6660 -577 6716
rect -521 6660 -512 6716
rect -592 6649 -512 6660
rect -577 5752 -521 6649
rect -397 5920 -341 6834
rect 44 6568 114 6578
rect 612 6574 668 7252
rect 44 6512 55 6568
rect 111 6512 114 6568
rect 44 6507 114 6512
rect 606 6568 676 6574
rect 606 6512 612 6568
rect 668 6512 676 6568
rect 55 6320 111 6507
rect 606 6503 676 6512
rect 873 6335 953 6347
rect 43 6312 127 6320
rect 43 6256 55 6312
rect 111 6256 127 6312
rect 873 6281 886 6335
rect 940 6281 953 6335
rect 873 6277 953 6281
rect 43 6243 127 6256
rect 352 6216 440 6228
rect 352 6160 365 6216
rect 421 6160 758 6216
rect 352 6152 440 6160
rect -408 5911 -329 5920
rect -408 5855 -397 5911
rect -341 5855 -329 5911
rect -408 5845 -329 5855
rect -589 5740 -509 5752
rect -589 5684 -577 5740
rect -521 5684 -509 5740
rect -589 5673 -509 5684
rect -577 4752 -521 5673
rect -397 4950 -341 5845
rect 702 5373 758 6160
rect 692 5360 780 5373
rect 23 5333 103 5344
rect 23 5277 37 5333
rect 93 5277 103 5333
rect 692 5306 703 5360
rect 757 5306 780 5360
rect 692 5297 780 5306
rect 23 5269 103 5277
rect 37 5055 93 5269
rect 351 5244 439 5253
rect 351 5188 362 5244
rect 418 5188 643 5244
rect 351 5176 439 5188
rect 25 5046 105 5055
rect 25 4990 37 5046
rect 93 4990 105 5046
rect 25 4980 105 4990
rect -407 4939 -328 4950
rect -407 4883 -397 4939
rect -341 4883 -328 4939
rect -407 4875 -328 4883
rect -588 4740 -508 4752
rect -588 4684 -577 4740
rect -521 4684 -508 4740
rect -588 4673 -508 4684
rect -577 3786 -521 4673
rect -397 3981 -341 4875
rect 587 4396 643 5188
rect 738 5046 818 5060
rect 738 4990 744 5046
rect 800 4990 818 5046
rect 738 4985 818 4990
rect 574 4386 662 4396
rect 574 4332 588 4386
rect 642 4332 662 4386
rect 574 4324 662 4332
rect -408 3970 -329 3981
rect -408 3914 -397 3970
rect -341 3914 -329 3970
rect -408 3906 -329 3914
rect -588 3773 -508 3786
rect -588 3717 -577 3773
rect -521 3717 -508 3773
rect -588 3707 -508 3717
rect -577 2852 -521 3707
rect -397 3008 -341 3906
rect 744 3427 800 4985
rect 735 3416 815 3427
rect 735 3362 745 3416
rect 799 3362 815 3416
rect 735 3352 815 3362
rect -408 3000 -329 3008
rect -408 2944 -397 3000
rect -341 2944 -329 3000
rect -408 2933 -329 2944
rect -588 2839 -508 2852
rect -588 2783 -577 2839
rect -521 2783 -508 2839
rect -588 2773 -508 2783
rect -577 1864 -521 2773
rect -397 2022 -341 2933
rect -65 2707 13 2721
rect 885 2711 941 6277
rect -65 2651 -52 2707
rect 4 2651 13 2707
rect -65 2644 13 2651
rect 878 2707 952 2711
rect 878 2651 885 2707
rect 941 2651 952 2707
rect -52 2417 4 2644
rect 878 2641 952 2651
rect 761 2441 848 2457
rect -63 2406 16 2417
rect -63 2350 -52 2406
rect 4 2350 16 2406
rect 761 2387 776 2441
rect 830 2387 848 2441
rect 761 2381 848 2387
rect -63 2338 16 2350
rect -237 2281 -156 2292
rect -237 2225 -224 2281
rect -168 2225 -156 2281
rect -237 2218 -156 2225
rect -411 2013 -332 2022
rect -411 1957 -397 2013
rect -341 1957 -332 2013
rect -411 1947 -332 1957
rect -587 1852 -507 1864
rect -587 1796 -577 1852
rect -521 1796 -507 1852
rect -587 1785 -507 1796
rect -577 888 -521 1785
rect -397 1051 -341 1947
rect -224 1129 -168 2218
rect -52 1404 4 2338
rect -63 1394 13 1404
rect -63 1338 -52 1394
rect 4 1338 13 1394
rect -63 1328 13 1338
rect 587 1212 669 1225
rect 587 1158 600 1212
rect 654 1158 669 1212
rect 587 1153 669 1158
rect -235 1122 -157 1129
rect -235 1066 -224 1122
rect -168 1066 -157 1122
rect -235 1055 -157 1066
rect -411 1041 -332 1051
rect -411 985 -397 1041
rect -341 985 -332 1041
rect -411 976 -332 985
rect -587 876 -507 888
rect -587 820 -577 876
rect -521 820 -507 876
rect -587 809 -507 820
rect -397 85 -341 976
rect -120 944 -44 955
rect -120 888 -110 944
rect -54 888 -44 944
rect -120 879 -44 888
rect -110 357 -54 879
rect 39 746 117 757
rect 599 753 655 1153
rect 775 954 831 2381
rect 953 1122 1031 1132
rect 953 1066 965 1122
rect 1021 1066 1031 1122
rect 953 1058 1031 1066
rect 766 944 842 954
rect 766 888 775 944
rect 831 888 842 944
rect 766 878 842 888
rect 39 690 54 746
rect 110 690 117 746
rect 39 685 117 690
rect 592 746 670 753
rect 592 690 599 746
rect 655 690 670 746
rect 54 475 110 685
rect 592 681 670 690
rect 965 504 1021 1058
rect 955 495 1033 504
rect 42 464 124 475
rect 42 408 54 464
rect 110 408 124 464
rect 955 441 966 495
rect 1020 441 1033 495
rect 955 430 1033 441
rect 42 403 124 408
rect -121 346 -45 357
rect -121 290 -110 346
rect -54 290 -45 346
rect -121 281 -45 290
rect -408 77 -329 85
rect -408 23 -396 77
rect -342 23 -329 77
rect -408 10 -329 23
<< via2 >>
rect 61 7494 117 7550
rect 623 7494 679 7550
rect 55 6512 111 6568
rect 612 6512 668 6568
rect 37 4990 93 5046
rect 744 4990 800 5046
rect -52 2651 4 2707
rect 885 2651 941 2707
rect -224 1066 -168 1122
rect -110 888 -54 944
rect 965 1066 1021 1122
rect 775 888 831 944
rect 54 690 110 746
rect 599 690 655 746
<< metal3 >>
rect 46 7550 132 7564
rect 610 7550 696 7558
rect 46 7494 61 7550
rect 117 7494 623 7550
rect 679 7494 696 7550
rect 46 7489 132 7494
rect 610 7483 696 7494
rect 44 6568 114 6578
rect 606 6568 676 6574
rect 44 6512 55 6568
rect 111 6512 612 6568
rect 668 6512 677 6568
rect 44 6507 114 6512
rect 606 6503 676 6512
rect 25 5046 105 5055
rect 738 5046 818 5060
rect 25 4990 37 5046
rect 93 4990 744 5046
rect 800 4990 818 5046
rect 25 4980 105 4990
rect 738 4985 818 4990
rect -65 2707 13 2721
rect 878 2707 952 2711
rect -65 2651 -52 2707
rect 4 2651 885 2707
rect 941 2651 952 2707
rect -65 2644 13 2651
rect 878 2641 952 2651
rect -235 1122 -157 1129
rect 953 1122 1031 1132
rect -235 1066 -224 1122
rect -168 1066 965 1122
rect 1021 1066 1031 1122
rect -235 1055 -157 1066
rect 953 1058 1031 1066
rect -120 944 -44 955
rect 766 944 842 954
rect -120 888 -110 944
rect -54 888 775 944
rect 831 888 842 944
rect -120 879 -44 888
rect 766 878 842 888
rect 39 746 117 757
rect 592 746 670 753
rect 39 690 54 746
rect 110 690 599 746
rect 655 690 670 746
rect 39 685 117 690
rect 592 681 670 690
<< labels >>
flabel via1 990 473 990 473 0 FreeSans 480 0 0 0 QB
port 0 nsew
flabel via1 792 2412 792 2412 0 FreeSans 480 0 0 0 Q
port 1 nsew
flabel metal1 90 8176 90 8176 0 FreeSans 480 0 0 0 Ri-1
port 2 nsew
flabel metal1 93 4257 93 4257 0 FreeSans 480 0 0 0 Ri
port 3 nsew
flabel metal1 93 3298 93 3298 0 FreeSans 480 0 0 0 Ci
port 4 nsew
flabel metal1 80 8650 80 8650 0 FreeSans 480 0 0 0 VDD
port 5 nsew
flabel metal1 0 7850 0 7850 0 FreeSans 480 0 0 0 VSS
port 6 nsew
flabel nsubdiffcont 344 8642 344 8642 0 FreeSans 320 0 0 0 NAND_14.VDD
flabel psubdiffcont 353 7850 353 7850 0 FreeSans 320 0 0 0 NAND_14.VSS
flabel metal1 104 8228 104 8228 0 FreeSans 480 0 0 0 NAND_14.B
flabel metal1 107 8130 107 8130 0 FreeSans 480 0 0 0 NAND_14.A
flabel metal1 606 8274 606 8274 0 FreeSans 480 0 0 0 NAND_14.OUT
flabel nsubdiffcont 344 6681 344 6681 0 FreeSans 320 0 0 0 NAND_13.VDD
flabel psubdiffcont 353 5889 353 5889 0 FreeSans 320 0 0 0 NAND_13.VSS
flabel metal1 104 6267 104 6267 0 FreeSans 480 0 0 0 NAND_13.B
flabel metal1 107 6169 107 6169 0 FreeSans 480 0 0 0 NAND_13.A
flabel metal1 606 6313 606 6313 0 FreeSans 480 0 0 0 NAND_13.OUT
flabel nsubdiffcont 344 5706 344 5706 0 FreeSans 320 0 0 0 NAND_12.VDD
flabel psubdiffcont 353 4914 353 4914 0 FreeSans 320 0 0 0 NAND_12.VSS
flabel metal1 104 5292 104 5292 0 FreeSans 480 0 0 0 NAND_12.B
flabel metal1 107 5194 107 5194 0 FreeSans 480 0 0 0 NAND_12.A
flabel metal1 606 5338 606 5338 0 FreeSans 480 0 0 0 NAND_12.OUT
flabel nsubdiffcont 344 4732 344 4732 0 FreeSans 320 0 0 0 NAND_11.VDD
flabel psubdiffcont 353 3940 353 3940 0 FreeSans 320 0 0 0 NAND_11.VSS
flabel metal1 104 4318 104 4318 0 FreeSans 480 0 0 0 NAND_11.B
flabel metal1 107 4220 107 4220 0 FreeSans 480 0 0 0 NAND_11.A
flabel metal1 606 4364 606 4364 0 FreeSans 480 0 0 0 NAND_11.OUT
flabel nsubdiffcont 344 2787 344 2787 0 FreeSans 320 0 0 0 NAND_9.VDD
flabel psubdiffcont 353 1995 353 1995 0 FreeSans 320 0 0 0 NAND_9.VSS
flabel metal1 104 2373 104 2373 0 FreeSans 480 0 0 0 NAND_9.B
flabel metal1 107 2275 107 2275 0 FreeSans 480 0 0 0 NAND_9.A
flabel metal1 606 2419 606 2419 0 FreeSans 480 0 0 0 NAND_9.OUT
flabel nsubdiffcont 344 841 344 841 0 FreeSans 320 0 0 0 NAND_3.VDD
flabel psubdiffcont 353 49 353 49 0 FreeSans 320 0 0 0 NAND_3.VSS
flabel metal1 104 427 104 427 0 FreeSans 480 0 0 0 NAND_3.B
flabel metal1 107 329 107 329 0 FreeSans 480 0 0 0 NAND_3.A
flabel metal1 606 473 606 473 0 FreeSans 480 0 0 0 NAND_3.OUT
flabel nsubdiffcont 344 1816 344 1816 0 FreeSans 320 0 0 0 NAND_2.VDD
flabel psubdiffcont 353 1024 353 1024 0 FreeSans 320 0 0 0 NAND_2.VSS
flabel metal1 104 1402 104 1402 0 FreeSans 480 0 0 0 NAND_2.B
flabel metal1 107 1304 107 1304 0 FreeSans 480 0 0 0 NAND_2.A
flabel metal1 606 1448 606 1448 0 FreeSans 480 0 0 0 NAND_2.OUT
flabel nsubdiffcont 344 7657 344 7657 0 FreeSans 320 0 0 0 NAND_1.VDD
flabel psubdiffcont 353 6865 353 6865 0 FreeSans 320 0 0 0 NAND_1.VSS
flabel metal1 104 7243 104 7243 0 FreeSans 480 0 0 0 NAND_1.B
flabel metal1 107 7145 107 7145 0 FreeSans 480 0 0 0 NAND_1.A
flabel metal1 606 7289 606 7289 0 FreeSans 480 0 0 0 NAND_1.OUT
flabel nsubdiffcont 344 3762 344 3762 0 FreeSans 320 0 0 0 NAND_0.VDD
flabel psubdiffcont 353 2970 353 2970 0 FreeSans 320 0 0 0 NAND_0.VSS
flabel metal1 104 3348 104 3348 0 FreeSans 480 0 0 0 NAND_0.B
flabel metal1 107 3250 107 3250 0 FreeSans 480 0 0 0 NAND_0.A
flabel metal1 606 3394 606 3394 0 FreeSans 480 0 0 0 NAND_0.OUT
<< end >>
