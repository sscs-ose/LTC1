magic
tech gf180mcuD
magscale 1 10
timestamp 1713971361
<< checkpaint >>
rect 1309 -2332 11664 7505
<< nwell >>
rect 5819 4436 5892 4509
<< pwell >>
rect 6177 -246 6262 2045
<< metal1 >>
rect 4540 5489 4618 5505
rect 4454 5486 4618 5489
rect 4454 5434 4552 5486
rect 4604 5434 4618 5486
rect 4454 5431 4618 5434
rect 4540 5418 4618 5431
rect 6035 4845 9234 4971
rect 4464 3875 4561 3903
rect 4386 3861 4561 3875
rect 4386 3809 4487 3861
rect 4539 3809 4561 3861
rect 4386 3795 4561 3809
rect 4464 3774 4561 3795
rect 3854 2429 3963 2485
rect 3854 2377 3885 2429
rect 3937 2377 3963 2429
rect 4218 2395 4406 2581
rect 3854 2358 3963 2377
rect 8730 2250 9484 2306
rect 3516 1989 3820 2007
rect 3502 1987 3820 1989
rect 3502 1985 3531 1987
rect 3475 1935 3531 1985
rect 3583 1935 3648 1987
rect 3700 1985 3820 1987
rect 3700 1935 3821 1985
rect 3475 1929 3821 1935
rect 3516 1910 3820 1929
rect 3334 -60 3839 -25
rect 6499 -59 9291 36
rect 3309 -65 3839 -60
rect 3309 -117 3380 -65
rect 3432 -117 3523 -65
rect 3575 -117 3839 -65
rect 3309 -121 3839 -117
rect 3334 -134 3839 -121
<< via1 >>
rect 4552 5434 4604 5486
rect 4487 3809 4539 3861
rect 3885 2377 3937 2429
rect 3531 1935 3583 1987
rect 3648 1935 3700 1987
rect 3380 -117 3432 -65
rect 3523 -117 3575 -65
<< metal2 >>
rect 4540 5486 4626 5505
rect 4540 5434 4552 5486
rect 4604 5437 4626 5486
rect 4604 5434 5814 5437
rect 4540 5418 5814 5434
rect 4556 5379 5814 5418
rect 5756 4533 5814 5379
rect 5729 4511 5825 4533
rect 5729 4455 5757 4511
rect 5813 4455 5825 4511
rect 5729 4436 5825 4455
rect 4464 3861 4561 3903
rect 4464 3809 4487 3861
rect 4539 3809 4561 3861
rect 4464 3774 4561 3809
rect 4471 3035 4551 3774
rect 4195 2493 4434 2615
rect 3854 2462 3963 2485
rect 4195 2462 4287 2493
rect 3822 2437 4287 2462
rect 4343 2462 4434 2493
rect 4343 2437 4881 2462
rect 3822 2429 4881 2437
rect 3822 2377 3885 2429
rect 3937 2377 4881 2429
rect 5756 2400 5814 4436
rect 3822 2354 4881 2377
rect 3516 1989 3820 2007
rect 3516 1933 3529 1989
rect 3585 1933 3646 1989
rect 3702 1933 3820 1989
rect 3516 1910 3820 1933
rect 3334 -63 3839 -25
rect 3334 -119 3378 -63
rect 3434 -119 3521 -63
rect 3577 -119 3839 -63
rect 3334 -134 3839 -119
<< via2 >>
rect 5757 4455 5813 4511
rect 4287 2437 4343 2493
rect 3529 1987 3585 1989
rect 3529 1935 3531 1987
rect 3531 1935 3583 1987
rect 3583 1935 3585 1987
rect 3529 1933 3585 1935
rect 3646 1987 3702 1989
rect 3646 1935 3648 1987
rect 3648 1935 3700 1987
rect 3700 1935 3702 1987
rect 3646 1933 3702 1935
rect 3378 -65 3434 -63
rect 3378 -117 3380 -65
rect 3380 -117 3432 -65
rect 3432 -117 3434 -65
rect 3378 -119 3434 -117
rect 3521 -65 3577 -63
rect 3521 -117 3523 -65
rect 3523 -117 3575 -65
rect 3575 -117 3577 -65
rect 3521 -119 3577 -117
<< metal3 >>
rect 5729 4519 5825 4533
rect 5729 4511 5937 4519
rect 5729 4455 5757 4511
rect 5813 4455 5937 4511
rect 5729 4446 5937 4455
rect 5729 4436 5892 4446
rect 5412 2844 5503 3411
rect 4770 2753 5503 2844
rect 4195 2567 4434 2615
rect 4770 2567 4861 2753
rect 4195 2493 4861 2567
rect 4195 2437 4287 2493
rect 4343 2476 4861 2493
rect 4343 2437 4434 2476
rect 4195 2375 4434 2437
rect 3516 1989 3820 2007
rect 3516 1933 3529 1989
rect 3585 1933 3646 1989
rect 3702 1933 3820 1989
rect 3516 1910 3820 1933
rect 3334 -63 3839 -25
rect 3334 -119 3378 -63
rect 3434 -119 3521 -63
rect 3577 -119 3901 -63
rect 3334 -134 3839 -119
use NMOS_Pairs  NMOS_Pairs_0
timestamp 1713971361
transform 1 0 4485 0 1 -292
box -791 -40 5078 2784
use VCTRL_mag  VCTRL_mag_0
timestamp 1713185578
transform 1 0 2760 0 1 3772
box 1436 -1269 6904 1605
<< labels >>
flabel metal1 s 3901 2453 3901 2453 0 FreeSans 2500 0 0 0 OUT
port 1 nsew
flabel metal1 s 3658 1952 3658 1952 0 FreeSans 2500 0 0 0 IN
port 2 nsew
flabel metal1 s 4491 5463 4491 5463 0 FreeSans 2500 0 0 0 OUTB
port 3 nsew
flabel metal1 s 9450 2273 9450 2273 0 FreeSans 2500 0 0 0 VCTRL2
port 4 nsew
flabel metal1 s 7684 4936 7684 4936 0 FreeSans 2500 0 0 0 VDD
port 5 nsew
flabel metal1 s 7594 -25 7594 -25 0 FreeSans 2500 0 0 0 VSS
port 6 nsew
flabel metal1 s 4424 3829 4424 3829 0 FreeSans 2500 0 0 0 VCTRL
port 7 nsew
flabel metal1 s 3314 -83 3314 -83 0 FreeSans 2500 0 0 0 INB
port 8 nsew
<< end >>
