magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1478 -1046 1478 1046
<< metal1 >>
rect -478 40 478 46
rect -478 14 -472 40
rect -446 14 -418 40
rect -392 14 -364 40
rect -338 14 -310 40
rect -284 14 -256 40
rect -230 14 -202 40
rect -176 14 -148 40
rect -122 14 -94 40
rect -68 14 -40 40
rect -14 14 14 40
rect 40 14 68 40
rect 94 14 122 40
rect 148 14 176 40
rect 202 14 230 40
rect 256 14 284 40
rect 310 14 338 40
rect 364 14 392 40
rect 418 14 446 40
rect 472 14 478 40
rect -478 -14 478 14
rect -478 -40 -472 -14
rect -446 -40 -418 -14
rect -392 -40 -364 -14
rect -338 -40 -310 -14
rect -284 -40 -256 -14
rect -230 -40 -202 -14
rect -176 -40 -148 -14
rect -122 -40 -94 -14
rect -68 -40 -40 -14
rect -14 -40 14 -14
rect 40 -40 68 -14
rect 94 -40 122 -14
rect 148 -40 176 -14
rect 202 -40 230 -14
rect 256 -40 284 -14
rect 310 -40 338 -14
rect 364 -40 392 -14
rect 418 -40 446 -14
rect 472 -40 478 -14
rect -478 -46 478 -40
<< via1 >>
rect -472 14 -446 40
rect -418 14 -392 40
rect -364 14 -338 40
rect -310 14 -284 40
rect -256 14 -230 40
rect -202 14 -176 40
rect -148 14 -122 40
rect -94 14 -68 40
rect -40 14 -14 40
rect 14 14 40 40
rect 68 14 94 40
rect 122 14 148 40
rect 176 14 202 40
rect 230 14 256 40
rect 284 14 310 40
rect 338 14 364 40
rect 392 14 418 40
rect 446 14 472 40
rect -472 -40 -446 -14
rect -418 -40 -392 -14
rect -364 -40 -338 -14
rect -310 -40 -284 -14
rect -256 -40 -230 -14
rect -202 -40 -176 -14
rect -148 -40 -122 -14
rect -94 -40 -68 -14
rect -40 -40 -14 -14
rect 14 -40 40 -14
rect 68 -40 94 -14
rect 122 -40 148 -14
rect 176 -40 202 -14
rect 230 -40 256 -14
rect 284 -40 310 -14
rect 338 -40 364 -14
rect 392 -40 418 -14
rect 446 -40 472 -14
<< metal2 >>
rect -478 40 478 46
rect -478 14 -472 40
rect -446 14 -418 40
rect -392 14 -364 40
rect -338 14 -310 40
rect -284 14 -256 40
rect -230 14 -202 40
rect -176 14 -148 40
rect -122 14 -94 40
rect -68 14 -40 40
rect -14 14 14 40
rect 40 14 68 40
rect 94 14 122 40
rect 148 14 176 40
rect 202 14 230 40
rect 256 14 284 40
rect 310 14 338 40
rect 364 14 392 40
rect 418 14 446 40
rect 472 14 478 40
rect -478 -14 478 14
rect -478 -40 -472 -14
rect -446 -40 -418 -14
rect -392 -40 -364 -14
rect -338 -40 -310 -14
rect -284 -40 -256 -14
rect -230 -40 -202 -14
rect -176 -40 -148 -14
rect -122 -40 -94 -14
rect -68 -40 -40 -14
rect -14 -40 14 -14
rect 40 -40 68 -14
rect 94 -40 122 -14
rect 148 -40 176 -14
rect 202 -40 230 -14
rect 256 -40 284 -14
rect 310 -40 338 -14
rect 364 -40 392 -14
rect 418 -40 446 -14
rect 472 -40 478 -14
rect -478 -46 478 -40
<< end >>
