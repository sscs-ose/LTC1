magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1046 -1046 1046 1046
<< metal1 >>
rect -46 40 46 46
rect -46 14 -40 40
rect -14 14 14 40
rect 40 14 46 40
rect -46 -14 46 14
rect -46 -40 -40 -14
rect -14 -40 14 -14
rect 40 -40 46 -14
rect -46 -46 46 -40
<< via1 >>
rect -40 14 -14 40
rect 14 14 40 40
rect -40 -40 -14 -14
rect 14 -40 40 -14
<< metal2 >>
rect -46 40 46 46
rect -46 14 -40 40
rect -14 14 14 40
rect 40 14 46 40
rect -46 -14 46 14
rect -46 -40 -40 -14
rect -14 -40 14 -14
rect 40 -40 46 -14
rect -46 -46 46 -40
<< end >>
