magic
tech gf180mcuC
magscale 1 10
timestamp 1699271742
<< nwell >>
rect -350 3294 1462 3508
<< psubdiff >>
rect -279 -193 1391 -180
rect -279 -239 -266 -193
rect -220 -239 -172 -193
rect -126 -239 -78 -193
rect -32 -239 16 -193
rect 62 -239 110 -193
rect 156 -239 204 -193
rect 250 -239 298 -193
rect 344 -239 392 -193
rect 438 -239 486 -193
rect 532 -239 580 -193
rect 626 -239 674 -193
rect 720 -239 768 -193
rect 814 -239 862 -193
rect 908 -239 956 -193
rect 1002 -239 1050 -193
rect 1096 -239 1144 -193
rect 1190 -239 1238 -193
rect 1284 -239 1332 -193
rect 1378 -239 1391 -193
rect -279 -252 1391 -239
<< nsubdiff >>
rect -326 3471 1438 3484
rect -326 3425 -313 3471
rect -267 3425 -219 3471
rect -173 3425 -125 3471
rect -79 3425 -31 3471
rect 15 3425 63 3471
rect 109 3425 157 3471
rect 203 3425 251 3471
rect 297 3425 345 3471
rect 391 3425 439 3471
rect 485 3425 533 3471
rect 579 3425 627 3471
rect 673 3425 721 3471
rect 767 3425 815 3471
rect 861 3425 909 3471
rect 955 3425 1003 3471
rect 1049 3425 1097 3471
rect 1143 3425 1191 3471
rect 1237 3425 1285 3471
rect 1331 3425 1379 3471
rect 1425 3425 1438 3471
rect -326 3412 1438 3425
<< psubdiffcont >>
rect -266 -239 -220 -193
rect -172 -239 -126 -193
rect -78 -239 -32 -193
rect 16 -239 62 -193
rect 110 -239 156 -193
rect 204 -239 250 -193
rect 298 -239 344 -193
rect 392 -239 438 -193
rect 486 -239 532 -193
rect 580 -239 626 -193
rect 674 -239 720 -193
rect 768 -239 814 -193
rect 862 -239 908 -193
rect 956 -239 1002 -193
rect 1050 -239 1096 -193
rect 1144 -239 1190 -193
rect 1238 -239 1284 -193
rect 1332 -239 1378 -193
<< nsubdiffcont >>
rect -313 3425 -267 3471
rect -219 3425 -173 3471
rect -125 3425 -79 3471
rect -31 3425 15 3471
rect 63 3425 109 3471
rect 157 3425 203 3471
rect 251 3425 297 3471
rect 345 3425 391 3471
rect 439 3425 485 3471
rect 533 3425 579 3471
rect 627 3425 673 3471
rect 721 3425 767 3471
rect 815 3425 861 3471
rect 909 3425 955 3471
rect 1003 3425 1049 3471
rect 1097 3425 1143 3471
rect 1191 3425 1237 3471
rect 1285 3425 1331 3471
rect 1379 3425 1425 3471
<< polysilicon >>
rect 112 3184 1288 3240
rect -176 1856 -120 2634
rect 112 2630 168 2640
rect 272 2630 328 2640
rect 432 2630 488 2640
rect 592 2630 648 2640
rect 752 2630 808 2640
rect 912 2630 968 2640
rect 1072 2630 1128 2640
rect 1232 2630 1288 2640
rect 112 2569 1288 2630
rect 112 1990 168 2569
rect 272 1990 328 2569
rect 432 1990 488 2569
rect 592 1990 648 2569
rect 752 1990 808 2569
rect 912 1990 968 2569
rect 1072 1990 1128 2569
rect 1232 1990 1288 2569
rect 112 1929 1288 1990
rect 112 1862 168 1929
rect 272 1862 328 1929
rect 432 1862 488 1929
rect 592 1862 648 1929
rect 752 1862 808 1929
rect 912 1862 968 1929
rect 1072 1862 1128 1929
rect 1232 1862 1288 1929
rect -296 1260 -224 1268
rect -176 1260 -120 1368
rect 112 1348 168 1368
rect -296 1255 -120 1260
rect -296 1209 -283 1255
rect -237 1209 -120 1255
rect -296 1204 -120 1209
rect -72 1270 0 1278
rect 112 1276 1128 1348
rect 112 1270 168 1276
rect -72 1265 168 1270
rect -72 1219 -59 1265
rect -13 1219 168 1265
rect -72 1214 168 1219
rect -72 1206 0 1214
rect -296 1196 -224 1204
rect -176 804 -120 1204
rect 112 804 168 840
rect 272 804 328 840
rect 432 804 488 840
rect 592 804 648 840
rect 752 804 808 840
rect 912 804 968 840
rect 1072 804 1128 840
rect 1232 804 1288 840
rect -176 744 1288 804
rect -176 411 -120 744
rect 112 411 168 744
rect 272 411 328 744
rect 432 411 488 744
rect 592 411 648 744
rect 752 411 808 744
rect 912 411 968 744
rect 1072 411 1128 744
rect 1232 411 1288 744
rect -176 351 1288 411
rect -176 318 -120 351
rect 112 312 168 351
rect 272 312 328 351
rect 432 312 488 351
rect 592 312 648 351
rect 752 312 808 351
rect 912 312 968 351
rect 1072 312 1128 351
rect 1232 312 1288 351
rect -176 -8 1288 48
<< polycontact >>
rect -283 1209 -237 1255
rect -59 1219 -13 1265
<< metal1 >>
rect -350 3471 1462 3504
rect -350 3425 -313 3471
rect -267 3425 -219 3471
rect -173 3425 -125 3471
rect -79 3425 -31 3471
rect 15 3425 63 3471
rect 109 3425 157 3471
rect 203 3425 251 3471
rect 297 3425 345 3471
rect 391 3425 439 3471
rect 485 3425 533 3471
rect 579 3425 627 3471
rect 673 3425 721 3471
rect 767 3425 815 3471
rect 861 3425 909 3471
rect 955 3425 1003 3471
rect 1049 3425 1097 3471
rect 1143 3425 1191 3471
rect 1237 3425 1285 3471
rect 1331 3425 1379 3471
rect 1425 3425 1462 3471
rect -350 3392 1462 3425
rect -251 1831 -205 3392
rect 37 3300 1363 3346
rect -91 1276 -45 2729
rect 37 2338 83 3300
rect 997 3254 1043 3300
rect 1162 3254 1208 3300
rect 1317 3254 1363 3300
rect 197 3208 883 3254
rect 13 2323 112 2338
rect 13 2253 28 2323
rect 96 2253 112 2323
rect 13 2239 112 2253
rect 37 1348 83 2239
rect 197 1850 243 3208
rect 357 2338 403 2708
rect 328 2323 427 2338
rect 328 2253 343 2323
rect 411 2253 427 2323
rect 328 2239 427 2253
rect 169 1680 268 1695
rect 169 1610 184 1680
rect 252 1610 268 1680
rect 169 1596 268 1610
rect 357 1348 403 2239
rect 517 1849 563 3208
rect 677 2338 723 2719
rect 648 2323 747 2338
rect 648 2253 663 2323
rect 731 2253 747 2323
rect 648 2239 747 2253
rect 489 1680 588 1695
rect 489 1610 504 1680
rect 572 1610 588 1680
rect 489 1596 588 1610
rect 677 1348 723 2239
rect 837 1849 883 3208
rect 997 3208 1363 3254
rect 997 2338 1043 3208
rect 968 2323 1067 2338
rect 968 2253 983 2323
rect 1051 2253 1067 2323
rect 968 2239 1067 2253
rect 997 1850 1043 2239
rect 1157 1695 1203 2720
rect 1317 2338 1363 3208
rect 1288 2323 1387 2338
rect 1288 2253 1303 2323
rect 1371 2253 1387 2323
rect 1288 2239 1387 2253
rect 809 1680 908 1695
rect 809 1610 824 1680
rect 892 1610 908 1680
rect 809 1596 908 1610
rect 1129 1680 1228 1695
rect 1129 1610 1144 1680
rect 1212 1610 1228 1680
rect 1129 1596 1228 1610
rect 37 1302 723 1348
rect -294 1255 -226 1266
rect -339 1209 -283 1255
rect -237 1209 -226 1255
rect -294 1198 -226 1209
rect -91 1265 -2 1276
rect -91 1219 -59 1265
rect -13 1219 -2 1265
rect -91 1208 -2 1219
rect -251 -160 -205 870
rect -91 305 -45 1208
rect 180 1180 226 1302
rect 320 1180 366 1302
rect 461 1180 507 1302
rect 580 1180 626 1302
rect 677 1180 723 1302
rect 37 1134 723 1180
rect 37 305 83 1134
rect 37 -68 83 98
rect 197 24 243 853
rect 357 303 403 1134
rect 517 24 563 854
rect 677 300 723 1134
rect 837 1230 883 1454
rect 1157 1230 1203 1596
rect 1317 1425 1363 2239
rect 1317 1379 1471 1425
rect 837 1184 1306 1230
rect 837 24 883 1184
rect 197 -22 883 24
rect 997 24 1043 853
rect 1157 305 1203 1184
rect 1317 24 1363 854
rect 997 -22 1363 24
rect 997 -68 1043 -22
rect 37 -114 1043 -68
rect -288 -193 1400 -160
rect -288 -239 -266 -193
rect -220 -239 -172 -193
rect -126 -239 -78 -193
rect -32 -239 16 -193
rect 62 -239 110 -193
rect 156 -239 204 -193
rect 250 -239 298 -193
rect 344 -239 392 -193
rect 438 -239 486 -193
rect 532 -239 580 -193
rect 626 -239 674 -193
rect 720 -239 768 -193
rect 814 -239 862 -193
rect 908 -239 956 -193
rect 1002 -239 1050 -193
rect 1096 -239 1144 -193
rect 1190 -239 1238 -193
rect 1284 -239 1332 -193
rect 1378 -239 1400 -193
rect -288 -272 1400 -239
<< via1 >>
rect 28 2253 96 2323
rect 343 2253 411 2323
rect 184 1610 252 1680
rect 663 2253 731 2323
rect 504 1610 572 1680
rect 983 2253 1051 2323
rect 1303 2253 1371 2323
rect 824 1610 892 1680
rect 1144 1610 1212 1680
<< metal2 >>
rect 5 2323 1397 2346
rect 5 2253 28 2323
rect 96 2253 343 2323
rect 411 2253 663 2323
rect 731 2253 983 2323
rect 1051 2253 1303 2323
rect 1371 2253 1397 2323
rect 5 2232 1397 2253
rect 162 1680 1232 1707
rect 162 1610 184 1680
rect 252 1610 504 1680
rect 572 1610 824 1680
rect 892 1610 1144 1680
rect 1212 1610 1232 1680
rect 162 1582 1232 1610
use nmos_3p3_RZHRT2  nmos_3p3_RZHRT2_0
timestamp 1692335619
transform 1 0 700 0 1 579
box -700 -579 700 579
use nmos_3p3_Y4JRT2  nmos_3p3_Y4JRT2_0
timestamp 1692335619
transform 1 0 -148 0 1 579
box -140 -579 140 579
use pmos_3p3_M6SUKR  pmos_3p3_M6SUKR_1
timestamp 1692335619
transform 1 0 700 0 1 2278
box -762 -1016 762 1016
use pmos_3p3_METUKR  pmos_3p3_METUKR_0
timestamp 1692335619
transform 1 0 -148 0 1 2278
box -202 -1016 202 1016
<< labels >>
flabel metal1 561 -216 561 -216 0 FreeSans 320 0 0 0 VSS
port 1 nsew
flabel nsubdiffcont 462 3448 462 3448 0 FreeSans 320 0 0 0 VDD
port 2 nsew
flabel polycontact -22 1239 -22 1239 0 FreeSans 640 0 0 0 CLKB
port 6 nsew
flabel metal1 1278 1204 1278 1204 0 FreeSans 640 0 0 0 VIN
port 7 nsew
flabel metal1 1433 1404 1433 1404 0 FreeSans 640 0 0 0 VOUT
port 8 nsew
flabel metal1 -318 1232 -318 1232 0 FreeSans 640 0 0 0 CLK
port 9 nsew
<< end >>
