magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1646 1019 1646
<< metal2 >>
rect -19 641 19 646
rect -19 613 -14 641
rect 14 613 19 641
rect -19 575 19 613
rect -19 547 -14 575
rect 14 547 19 575
rect -19 509 19 547
rect -19 481 -14 509
rect 14 481 19 509
rect -19 443 19 481
rect -19 415 -14 443
rect 14 415 19 443
rect -19 377 19 415
rect -19 349 -14 377
rect 14 349 19 377
rect -19 311 19 349
rect -19 283 -14 311
rect 14 283 19 311
rect -19 245 19 283
rect -19 217 -14 245
rect 14 217 19 245
rect -19 179 19 217
rect -19 151 -14 179
rect 14 151 19 179
rect -19 113 19 151
rect -19 85 -14 113
rect 14 85 19 113
rect -19 47 19 85
rect -19 19 -14 47
rect 14 19 19 47
rect -19 -19 19 19
rect -19 -47 -14 -19
rect 14 -47 19 -19
rect -19 -85 19 -47
rect -19 -113 -14 -85
rect 14 -113 19 -85
rect -19 -151 19 -113
rect -19 -179 -14 -151
rect 14 -179 19 -151
rect -19 -217 19 -179
rect -19 -245 -14 -217
rect 14 -245 19 -217
rect -19 -283 19 -245
rect -19 -311 -14 -283
rect 14 -311 19 -283
rect -19 -349 19 -311
rect -19 -377 -14 -349
rect 14 -377 19 -349
rect -19 -415 19 -377
rect -19 -443 -14 -415
rect 14 -443 19 -415
rect -19 -481 19 -443
rect -19 -509 -14 -481
rect 14 -509 19 -481
rect -19 -547 19 -509
rect -19 -575 -14 -547
rect 14 -575 19 -547
rect -19 -613 19 -575
rect -19 -641 -14 -613
rect 14 -641 19 -613
rect -19 -646 19 -641
<< via2 >>
rect -14 613 14 641
rect -14 547 14 575
rect -14 481 14 509
rect -14 415 14 443
rect -14 349 14 377
rect -14 283 14 311
rect -14 217 14 245
rect -14 151 14 179
rect -14 85 14 113
rect -14 19 14 47
rect -14 -47 14 -19
rect -14 -113 14 -85
rect -14 -179 14 -151
rect -14 -245 14 -217
rect -14 -311 14 -283
rect -14 -377 14 -349
rect -14 -443 14 -415
rect -14 -509 14 -481
rect -14 -575 14 -547
rect -14 -641 14 -613
<< metal3 >>
rect -19 641 19 646
rect -19 613 -14 641
rect 14 613 19 641
rect -19 575 19 613
rect -19 547 -14 575
rect 14 547 19 575
rect -19 509 19 547
rect -19 481 -14 509
rect 14 481 19 509
rect -19 443 19 481
rect -19 415 -14 443
rect 14 415 19 443
rect -19 377 19 415
rect -19 349 -14 377
rect 14 349 19 377
rect -19 311 19 349
rect -19 283 -14 311
rect 14 283 19 311
rect -19 245 19 283
rect -19 217 -14 245
rect 14 217 19 245
rect -19 179 19 217
rect -19 151 -14 179
rect 14 151 19 179
rect -19 113 19 151
rect -19 85 -14 113
rect 14 85 19 113
rect -19 47 19 85
rect -19 19 -14 47
rect 14 19 19 47
rect -19 -19 19 19
rect -19 -47 -14 -19
rect 14 -47 19 -19
rect -19 -85 19 -47
rect -19 -113 -14 -85
rect 14 -113 19 -85
rect -19 -151 19 -113
rect -19 -179 -14 -151
rect 14 -179 19 -151
rect -19 -217 19 -179
rect -19 -245 -14 -217
rect 14 -245 19 -217
rect -19 -283 19 -245
rect -19 -311 -14 -283
rect 14 -311 19 -283
rect -19 -349 19 -311
rect -19 -377 -14 -349
rect 14 -377 19 -349
rect -19 -415 19 -377
rect -19 -443 -14 -415
rect 14 -443 19 -415
rect -19 -481 19 -443
rect -19 -509 -14 -481
rect 14 -509 19 -481
rect -19 -547 19 -509
rect -19 -575 -14 -547
rect 14 -575 19 -547
rect -19 -613 19 -575
rect -19 -641 -14 -613
rect 14 -641 19 -613
rect -19 -646 19 -641
<< end >>
