magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1643 1019 1643
<< metal1 >>
rect -19 637 19 643
rect -19 -637 -13 637
rect 13 -637 19 637
rect -19 -643 19 -637
<< via1 >>
rect -13 -637 13 637
<< metal2 >>
rect -19 637 19 643
rect -19 -637 -13 637
rect 13 -637 19 637
rect -19 -643 19 -637
<< end >>
