magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1331 -1019 1331 1019
<< metal1 >>
rect -331 13 331 19
rect -331 -13 -325 13
rect 325 -13 331 13
rect -331 -19 331 -13
<< via1 >>
rect -325 -13 325 13
<< metal2 >>
rect -331 13 331 19
rect -331 -13 -325 13
rect 325 -13 331 13
rect -331 -19 331 -13
<< end >>
