** sch_path: /home/shahid/GF180Projects/Tapeout/Xschem/MUX_8x1/muxWnonovpclkTB.sch
**.subckt muxWnonovpclkTB OUT
*.opin OUT
V1 IN1 GND 900m
.save i(v1)
V2 IN2 GND 700m
.save i(v2)
V3 IN3 GND 400m
.save i(v3)
V4 IN4 GND 100m
.save i(v4)
V6 IN5 GND 0
.save i(v6)
V7 IN6 GND 400m
.save i(v7)
V8 IN7 GND 700m
.save i(v8)
V9 IN8 GND 900m
.save i(v9)
V10 VDD VSS 3.3
.save i(v10)
V11 A1 VSS pulse(3.3 0 0 100p 100p 5u 10u)
.save i(v11)
V12 B1 VSS pulse(3.3 0 0 100p 100p 10u 20u)0
.save i(v12)
V13 C1 VSS pulse(3.3 0 0 100p 100p 20u 40u)3.3
.save i(v13)
V14 VSS GND 0
.save i(v14)
V5 EN GND 3.3
.save i(v5)
R1 OUT GND 10k m=1
x1 VSS VDD IN1 IN2 IN3 B1 IN4 OUT IN5 C1 IN6 IN7 IN8 A1 EN pex_MUX_8x1_Layout
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.include pex_MUX_8x1_Layout.spice
.control
set color0 = white
set color1 = black
save all
*dc v10 0 3.3 0.1
tran 100n 40u
*plot v(IN1) v(IN2)+4 v(IN3)+8 v(IN4)+12 v(IN5)+16 v(IN6)+20 v(IN7)+24 v(IN8)+28 v(OUT)+32
plot v(OUT)
plot v(A1) v(B1)+3.5 v(C1)+7
*write test_nfet_03v3.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
