magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2495 -9745 2495 9745
<< psubdiff >>
rect -495 7723 495 7745
rect -495 -7723 -473 7723
rect 473 -7723 495 7723
rect -495 -7745 495 -7723
<< psubdiffcont >>
rect -473 -7723 473 7723
<< metal1 >>
rect -484 7723 484 7734
rect -484 -7723 -473 7723
rect 473 -7723 484 7723
rect -484 -7734 484 -7723
<< end >>
