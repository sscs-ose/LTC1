magic
tech gf180mcuC
magscale 1 10
timestamp 1694610567
<< nwell >>
rect -4904 -386 4904 386
<< nsubdiff >>
rect -4880 290 4880 362
rect -4880 -290 -4808 290
rect 4808 -290 4880 290
rect -4880 -362 4880 -290
<< polysilicon >>
rect -4720 189 -4520 202
rect -4720 143 -4707 189
rect -4533 143 -4520 189
rect -4720 100 -4520 143
rect -4720 -143 -4520 -100
rect -4720 -189 -4707 -143
rect -4533 -189 -4520 -143
rect -4720 -202 -4520 -189
rect -4440 189 -4240 202
rect -4440 143 -4427 189
rect -4253 143 -4240 189
rect -4440 100 -4240 143
rect -4440 -143 -4240 -100
rect -4440 -189 -4427 -143
rect -4253 -189 -4240 -143
rect -4440 -202 -4240 -189
rect -4160 189 -3960 202
rect -4160 143 -4147 189
rect -3973 143 -3960 189
rect -4160 100 -3960 143
rect -4160 -143 -3960 -100
rect -4160 -189 -4147 -143
rect -3973 -189 -3960 -143
rect -4160 -202 -3960 -189
rect -3880 189 -3680 202
rect -3880 143 -3867 189
rect -3693 143 -3680 189
rect -3880 100 -3680 143
rect -3880 -143 -3680 -100
rect -3880 -189 -3867 -143
rect -3693 -189 -3680 -143
rect -3880 -202 -3680 -189
rect -3600 189 -3400 202
rect -3600 143 -3587 189
rect -3413 143 -3400 189
rect -3600 100 -3400 143
rect -3600 -143 -3400 -100
rect -3600 -189 -3587 -143
rect -3413 -189 -3400 -143
rect -3600 -202 -3400 -189
rect -3320 189 -3120 202
rect -3320 143 -3307 189
rect -3133 143 -3120 189
rect -3320 100 -3120 143
rect -3320 -143 -3120 -100
rect -3320 -189 -3307 -143
rect -3133 -189 -3120 -143
rect -3320 -202 -3120 -189
rect -3040 189 -2840 202
rect -3040 143 -3027 189
rect -2853 143 -2840 189
rect -3040 100 -2840 143
rect -3040 -143 -2840 -100
rect -3040 -189 -3027 -143
rect -2853 -189 -2840 -143
rect -3040 -202 -2840 -189
rect -2760 189 -2560 202
rect -2760 143 -2747 189
rect -2573 143 -2560 189
rect -2760 100 -2560 143
rect -2760 -143 -2560 -100
rect -2760 -189 -2747 -143
rect -2573 -189 -2560 -143
rect -2760 -202 -2560 -189
rect -2480 189 -2280 202
rect -2480 143 -2467 189
rect -2293 143 -2280 189
rect -2480 100 -2280 143
rect -2480 -143 -2280 -100
rect -2480 -189 -2467 -143
rect -2293 -189 -2280 -143
rect -2480 -202 -2280 -189
rect -2200 189 -2000 202
rect -2200 143 -2187 189
rect -2013 143 -2000 189
rect -2200 100 -2000 143
rect -2200 -143 -2000 -100
rect -2200 -189 -2187 -143
rect -2013 -189 -2000 -143
rect -2200 -202 -2000 -189
rect -1920 189 -1720 202
rect -1920 143 -1907 189
rect -1733 143 -1720 189
rect -1920 100 -1720 143
rect -1920 -143 -1720 -100
rect -1920 -189 -1907 -143
rect -1733 -189 -1720 -143
rect -1920 -202 -1720 -189
rect -1640 189 -1440 202
rect -1640 143 -1627 189
rect -1453 143 -1440 189
rect -1640 100 -1440 143
rect -1640 -143 -1440 -100
rect -1640 -189 -1627 -143
rect -1453 -189 -1440 -143
rect -1640 -202 -1440 -189
rect -1360 189 -1160 202
rect -1360 143 -1347 189
rect -1173 143 -1160 189
rect -1360 100 -1160 143
rect -1360 -143 -1160 -100
rect -1360 -189 -1347 -143
rect -1173 -189 -1160 -143
rect -1360 -202 -1160 -189
rect -1080 189 -880 202
rect -1080 143 -1067 189
rect -893 143 -880 189
rect -1080 100 -880 143
rect -1080 -143 -880 -100
rect -1080 -189 -1067 -143
rect -893 -189 -880 -143
rect -1080 -202 -880 -189
rect -800 189 -600 202
rect -800 143 -787 189
rect -613 143 -600 189
rect -800 100 -600 143
rect -800 -143 -600 -100
rect -800 -189 -787 -143
rect -613 -189 -600 -143
rect -800 -202 -600 -189
rect -520 189 -320 202
rect -520 143 -507 189
rect -333 143 -320 189
rect -520 100 -320 143
rect -520 -143 -320 -100
rect -520 -189 -507 -143
rect -333 -189 -320 -143
rect -520 -202 -320 -189
rect -240 189 -40 202
rect -240 143 -227 189
rect -53 143 -40 189
rect -240 100 -40 143
rect -240 -143 -40 -100
rect -240 -189 -227 -143
rect -53 -189 -40 -143
rect -240 -202 -40 -189
rect 40 189 240 202
rect 40 143 53 189
rect 227 143 240 189
rect 40 100 240 143
rect 40 -143 240 -100
rect 40 -189 53 -143
rect 227 -189 240 -143
rect 40 -202 240 -189
rect 320 189 520 202
rect 320 143 333 189
rect 507 143 520 189
rect 320 100 520 143
rect 320 -143 520 -100
rect 320 -189 333 -143
rect 507 -189 520 -143
rect 320 -202 520 -189
rect 600 189 800 202
rect 600 143 613 189
rect 787 143 800 189
rect 600 100 800 143
rect 600 -143 800 -100
rect 600 -189 613 -143
rect 787 -189 800 -143
rect 600 -202 800 -189
rect 880 189 1080 202
rect 880 143 893 189
rect 1067 143 1080 189
rect 880 100 1080 143
rect 880 -143 1080 -100
rect 880 -189 893 -143
rect 1067 -189 1080 -143
rect 880 -202 1080 -189
rect 1160 189 1360 202
rect 1160 143 1173 189
rect 1347 143 1360 189
rect 1160 100 1360 143
rect 1160 -143 1360 -100
rect 1160 -189 1173 -143
rect 1347 -189 1360 -143
rect 1160 -202 1360 -189
rect 1440 189 1640 202
rect 1440 143 1453 189
rect 1627 143 1640 189
rect 1440 100 1640 143
rect 1440 -143 1640 -100
rect 1440 -189 1453 -143
rect 1627 -189 1640 -143
rect 1440 -202 1640 -189
rect 1720 189 1920 202
rect 1720 143 1733 189
rect 1907 143 1920 189
rect 1720 100 1920 143
rect 1720 -143 1920 -100
rect 1720 -189 1733 -143
rect 1907 -189 1920 -143
rect 1720 -202 1920 -189
rect 2000 189 2200 202
rect 2000 143 2013 189
rect 2187 143 2200 189
rect 2000 100 2200 143
rect 2000 -143 2200 -100
rect 2000 -189 2013 -143
rect 2187 -189 2200 -143
rect 2000 -202 2200 -189
rect 2280 189 2480 202
rect 2280 143 2293 189
rect 2467 143 2480 189
rect 2280 100 2480 143
rect 2280 -143 2480 -100
rect 2280 -189 2293 -143
rect 2467 -189 2480 -143
rect 2280 -202 2480 -189
rect 2560 189 2760 202
rect 2560 143 2573 189
rect 2747 143 2760 189
rect 2560 100 2760 143
rect 2560 -143 2760 -100
rect 2560 -189 2573 -143
rect 2747 -189 2760 -143
rect 2560 -202 2760 -189
rect 2840 189 3040 202
rect 2840 143 2853 189
rect 3027 143 3040 189
rect 2840 100 3040 143
rect 2840 -143 3040 -100
rect 2840 -189 2853 -143
rect 3027 -189 3040 -143
rect 2840 -202 3040 -189
rect 3120 189 3320 202
rect 3120 143 3133 189
rect 3307 143 3320 189
rect 3120 100 3320 143
rect 3120 -143 3320 -100
rect 3120 -189 3133 -143
rect 3307 -189 3320 -143
rect 3120 -202 3320 -189
rect 3400 189 3600 202
rect 3400 143 3413 189
rect 3587 143 3600 189
rect 3400 100 3600 143
rect 3400 -143 3600 -100
rect 3400 -189 3413 -143
rect 3587 -189 3600 -143
rect 3400 -202 3600 -189
rect 3680 189 3880 202
rect 3680 143 3693 189
rect 3867 143 3880 189
rect 3680 100 3880 143
rect 3680 -143 3880 -100
rect 3680 -189 3693 -143
rect 3867 -189 3880 -143
rect 3680 -202 3880 -189
rect 3960 189 4160 202
rect 3960 143 3973 189
rect 4147 143 4160 189
rect 3960 100 4160 143
rect 3960 -143 4160 -100
rect 3960 -189 3973 -143
rect 4147 -189 4160 -143
rect 3960 -202 4160 -189
rect 4240 189 4440 202
rect 4240 143 4253 189
rect 4427 143 4440 189
rect 4240 100 4440 143
rect 4240 -143 4440 -100
rect 4240 -189 4253 -143
rect 4427 -189 4440 -143
rect 4240 -202 4440 -189
rect 4520 189 4720 202
rect 4520 143 4533 189
rect 4707 143 4720 189
rect 4520 100 4720 143
rect 4520 -143 4720 -100
rect 4520 -189 4533 -143
rect 4707 -189 4720 -143
rect 4520 -202 4720 -189
<< polycontact >>
rect -4707 143 -4533 189
rect -4707 -189 -4533 -143
rect -4427 143 -4253 189
rect -4427 -189 -4253 -143
rect -4147 143 -3973 189
rect -4147 -189 -3973 -143
rect -3867 143 -3693 189
rect -3867 -189 -3693 -143
rect -3587 143 -3413 189
rect -3587 -189 -3413 -143
rect -3307 143 -3133 189
rect -3307 -189 -3133 -143
rect -3027 143 -2853 189
rect -3027 -189 -2853 -143
rect -2747 143 -2573 189
rect -2747 -189 -2573 -143
rect -2467 143 -2293 189
rect -2467 -189 -2293 -143
rect -2187 143 -2013 189
rect -2187 -189 -2013 -143
rect -1907 143 -1733 189
rect -1907 -189 -1733 -143
rect -1627 143 -1453 189
rect -1627 -189 -1453 -143
rect -1347 143 -1173 189
rect -1347 -189 -1173 -143
rect -1067 143 -893 189
rect -1067 -189 -893 -143
rect -787 143 -613 189
rect -787 -189 -613 -143
rect -507 143 -333 189
rect -507 -189 -333 -143
rect -227 143 -53 189
rect -227 -189 -53 -143
rect 53 143 227 189
rect 53 -189 227 -143
rect 333 143 507 189
rect 333 -189 507 -143
rect 613 143 787 189
rect 613 -189 787 -143
rect 893 143 1067 189
rect 893 -189 1067 -143
rect 1173 143 1347 189
rect 1173 -189 1347 -143
rect 1453 143 1627 189
rect 1453 -189 1627 -143
rect 1733 143 1907 189
rect 1733 -189 1907 -143
rect 2013 143 2187 189
rect 2013 -189 2187 -143
rect 2293 143 2467 189
rect 2293 -189 2467 -143
rect 2573 143 2747 189
rect 2573 -189 2747 -143
rect 2853 143 3027 189
rect 2853 -189 3027 -143
rect 3133 143 3307 189
rect 3133 -189 3307 -143
rect 3413 143 3587 189
rect 3413 -189 3587 -143
rect 3693 143 3867 189
rect 3693 -189 3867 -143
rect 3973 143 4147 189
rect 3973 -189 4147 -143
rect 4253 143 4427 189
rect 4253 -189 4427 -143
rect 4533 143 4707 189
rect 4533 -189 4707 -143
<< ppolyres >>
rect -4720 -100 -4520 100
rect -4440 -100 -4240 100
rect -4160 -100 -3960 100
rect -3880 -100 -3680 100
rect -3600 -100 -3400 100
rect -3320 -100 -3120 100
rect -3040 -100 -2840 100
rect -2760 -100 -2560 100
rect -2480 -100 -2280 100
rect -2200 -100 -2000 100
rect -1920 -100 -1720 100
rect -1640 -100 -1440 100
rect -1360 -100 -1160 100
rect -1080 -100 -880 100
rect -800 -100 -600 100
rect -520 -100 -320 100
rect -240 -100 -40 100
rect 40 -100 240 100
rect 320 -100 520 100
rect 600 -100 800 100
rect 880 -100 1080 100
rect 1160 -100 1360 100
rect 1440 -100 1640 100
rect 1720 -100 1920 100
rect 2000 -100 2200 100
rect 2280 -100 2480 100
rect 2560 -100 2760 100
rect 2840 -100 3040 100
rect 3120 -100 3320 100
rect 3400 -100 3600 100
rect 3680 -100 3880 100
rect 3960 -100 4160 100
rect 4240 -100 4440 100
rect 4520 -100 4720 100
<< metal1 >>
rect -4718 143 -4707 189
rect -4533 143 -4522 189
rect -4438 143 -4427 189
rect -4253 143 -4242 189
rect -4158 143 -4147 189
rect -3973 143 -3962 189
rect -3878 143 -3867 189
rect -3693 143 -3682 189
rect -3598 143 -3587 189
rect -3413 143 -3402 189
rect -3318 143 -3307 189
rect -3133 143 -3122 189
rect -3038 143 -3027 189
rect -2853 143 -2842 189
rect -2758 143 -2747 189
rect -2573 143 -2562 189
rect -2478 143 -2467 189
rect -2293 143 -2282 189
rect -2198 143 -2187 189
rect -2013 143 -2002 189
rect -1918 143 -1907 189
rect -1733 143 -1722 189
rect -1638 143 -1627 189
rect -1453 143 -1442 189
rect -1358 143 -1347 189
rect -1173 143 -1162 189
rect -1078 143 -1067 189
rect -893 143 -882 189
rect -798 143 -787 189
rect -613 143 -602 189
rect -518 143 -507 189
rect -333 143 -322 189
rect -238 143 -227 189
rect -53 143 -42 189
rect 42 143 53 189
rect 227 143 238 189
rect 322 143 333 189
rect 507 143 518 189
rect 602 143 613 189
rect 787 143 798 189
rect 882 143 893 189
rect 1067 143 1078 189
rect 1162 143 1173 189
rect 1347 143 1358 189
rect 1442 143 1453 189
rect 1627 143 1638 189
rect 1722 143 1733 189
rect 1907 143 1918 189
rect 2002 143 2013 189
rect 2187 143 2198 189
rect 2282 143 2293 189
rect 2467 143 2478 189
rect 2562 143 2573 189
rect 2747 143 2758 189
rect 2842 143 2853 189
rect 3027 143 3038 189
rect 3122 143 3133 189
rect 3307 143 3318 189
rect 3402 143 3413 189
rect 3587 143 3598 189
rect 3682 143 3693 189
rect 3867 143 3878 189
rect 3962 143 3973 189
rect 4147 143 4158 189
rect 4242 143 4253 189
rect 4427 143 4438 189
rect 4522 143 4533 189
rect 4707 143 4718 189
rect -4718 -189 -4707 -143
rect -4533 -189 -4522 -143
rect -4438 -189 -4427 -143
rect -4253 -189 -4242 -143
rect -4158 -189 -4147 -143
rect -3973 -189 -3962 -143
rect -3878 -189 -3867 -143
rect -3693 -189 -3682 -143
rect -3598 -189 -3587 -143
rect -3413 -189 -3402 -143
rect -3318 -189 -3307 -143
rect -3133 -189 -3122 -143
rect -3038 -189 -3027 -143
rect -2853 -189 -2842 -143
rect -2758 -189 -2747 -143
rect -2573 -189 -2562 -143
rect -2478 -189 -2467 -143
rect -2293 -189 -2282 -143
rect -2198 -189 -2187 -143
rect -2013 -189 -2002 -143
rect -1918 -189 -1907 -143
rect -1733 -189 -1722 -143
rect -1638 -189 -1627 -143
rect -1453 -189 -1442 -143
rect -1358 -189 -1347 -143
rect -1173 -189 -1162 -143
rect -1078 -189 -1067 -143
rect -893 -189 -882 -143
rect -798 -189 -787 -143
rect -613 -189 -602 -143
rect -518 -189 -507 -143
rect -333 -189 -322 -143
rect -238 -189 -227 -143
rect -53 -189 -42 -143
rect 42 -189 53 -143
rect 227 -189 238 -143
rect 322 -189 333 -143
rect 507 -189 518 -143
rect 602 -189 613 -143
rect 787 -189 798 -143
rect 882 -189 893 -143
rect 1067 -189 1078 -143
rect 1162 -189 1173 -143
rect 1347 -189 1358 -143
rect 1442 -189 1453 -143
rect 1627 -189 1638 -143
rect 1722 -189 1733 -143
rect 1907 -189 1918 -143
rect 2002 -189 2013 -143
rect 2187 -189 2198 -143
rect 2282 -189 2293 -143
rect 2467 -189 2478 -143
rect 2562 -189 2573 -143
rect 2747 -189 2758 -143
rect 2842 -189 2853 -143
rect 3027 -189 3038 -143
rect 3122 -189 3133 -143
rect 3307 -189 3318 -143
rect 3402 -189 3413 -143
rect 3587 -189 3598 -143
rect 3682 -189 3693 -143
rect 3867 -189 3878 -143
rect 3962 -189 3973 -143
rect 4147 -189 4158 -143
rect 4242 -189 4253 -143
rect 4427 -189 4438 -143
rect 4522 -189 4533 -143
rect 4707 -189 4718 -143
<< properties >>
string FIXED_BBOX -4844 -326 4844 326
string gencell ppolyf_u
string library gf180mcu
string parameters w 1.0 l 1.0 m 1 nx 34 wmin 0.80 lmin 1.00 rho 315 val 338.709 dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0
<< end >>
