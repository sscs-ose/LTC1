magic
tech gf180mcuC
magscale 1 10
timestamp 1693830637
<< nwell >>
rect -3258 1140 3962 1350
rect -3256 760 3954 1140
<< pwell >>
rect -538 2159 2322 2415
rect -538 1785 2510 2041
rect -2069 0 -1670 256
rect -860 0 -852 256
rect -324 0 -316 256
rect 8 0 16 256
rect 544 0 552 256
rect 876 0 884 256
rect 1412 94 1420 256
rect -2069 -326 -1659 -70
rect -861 -325 -852 -70
rect -324 -326 -316 -70
rect 8 -326 16 -70
rect 544 -326 552 -70
rect 876 -326 884 -70
rect 1343 -326 1599 94
rect 2231 0 2620 256
rect 2227 -326 2620 -70
<< psubdiff >>
rect -3789 3833 -3630 3855
rect -3789 3712 -3763 3833
rect -3652 3712 -3630 3833
rect -3789 3684 -3630 3712
rect -3422 3838 -3263 3860
rect -3422 3717 -3396 3838
rect -3285 3717 -3263 3838
rect -3422 3689 -3263 3717
rect -2963 3838 -2804 3860
rect -2963 3717 -2937 3838
rect -2826 3717 -2804 3838
rect -2963 3689 -2804 3717
rect -2733 3838 -2574 3860
rect -2733 3717 -2707 3838
rect -2596 3717 -2574 3838
rect -2733 3689 -2574 3717
rect -2503 3838 -2344 3860
rect -2503 3717 -2477 3838
rect -2366 3717 -2344 3838
rect -2503 3689 -2344 3717
rect -2273 3838 -2114 3860
rect -2273 3717 -2247 3838
rect -2136 3717 -2114 3838
rect -2273 3689 -2114 3717
rect -2043 3838 -1884 3860
rect -2043 3717 -2017 3838
rect -1906 3717 -1884 3838
rect -2043 3689 -1884 3717
rect -1813 3838 -1654 3860
rect -1813 3717 -1787 3838
rect -1676 3717 -1654 3838
rect -1813 3689 -1654 3717
rect -1583 3838 -1424 3860
rect -1583 3717 -1557 3838
rect -1446 3717 -1424 3838
rect -1583 3689 -1424 3717
rect -1353 3838 -1194 3860
rect -1353 3717 -1327 3838
rect -1216 3717 -1194 3838
rect -1353 3689 -1194 3717
rect -1123 3838 -964 3860
rect -1123 3717 -1097 3838
rect -986 3717 -964 3838
rect -1123 3689 -964 3717
rect -893 3838 -734 3860
rect -893 3717 -867 3838
rect -756 3717 -734 3838
rect -893 3689 -734 3717
rect -663 3838 -504 3860
rect -663 3717 -637 3838
rect -526 3717 -504 3838
rect -663 3689 -504 3717
rect -433 3838 -274 3860
rect -433 3717 -407 3838
rect -296 3717 -274 3838
rect -433 3689 -274 3717
rect -203 3838 -44 3860
rect -203 3717 -177 3838
rect -66 3717 -44 3838
rect -203 3689 -44 3717
rect 27 3838 186 3860
rect 27 3717 53 3838
rect 164 3717 186 3838
rect 27 3689 186 3717
rect 257 3838 416 3860
rect 257 3717 283 3838
rect 394 3717 416 3838
rect 257 3689 416 3717
rect 487 3838 646 3860
rect 487 3717 513 3838
rect 624 3717 646 3838
rect 487 3689 646 3717
rect 717 3838 876 3860
rect 717 3717 743 3838
rect 854 3717 876 3838
rect 717 3689 876 3717
rect 947 3838 1106 3860
rect 947 3717 973 3838
rect 1084 3717 1106 3838
rect 947 3689 1106 3717
rect 1177 3838 1336 3860
rect 1177 3717 1203 3838
rect 1314 3717 1336 3838
rect 1177 3689 1336 3717
rect 1407 3838 1566 3860
rect 1407 3717 1433 3838
rect 1544 3717 1566 3838
rect 1407 3689 1566 3717
rect 1637 3838 1796 3860
rect 1637 3717 1663 3838
rect 1774 3717 1796 3838
rect 1637 3689 1796 3717
rect 1867 3838 2026 3860
rect 1867 3717 1893 3838
rect 2004 3717 2026 3838
rect 1867 3689 2026 3717
rect 2097 3838 2256 3860
rect 2097 3717 2123 3838
rect 2234 3717 2256 3838
rect 2097 3689 2256 3717
rect 2327 3838 2486 3860
rect 2327 3717 2353 3838
rect 2464 3717 2486 3838
rect 2327 3689 2486 3717
rect 2557 3838 2716 3860
rect 2557 3717 2583 3838
rect 2694 3717 2716 3838
rect 2557 3689 2716 3717
rect 2787 3838 2946 3860
rect 2787 3717 2813 3838
rect 2924 3717 2946 3838
rect 2787 3689 2946 3717
rect 3017 3838 3176 3860
rect 3017 3717 3043 3838
rect 3154 3717 3176 3838
rect 3017 3689 3176 3717
rect 3247 3838 3406 3860
rect 3247 3717 3273 3838
rect 3384 3717 3406 3838
rect 3247 3689 3406 3717
rect 3477 3838 3636 3860
rect 3477 3717 3503 3838
rect 3614 3717 3636 3838
rect 3477 3689 3636 3717
rect 3715 3838 3874 3860
rect 3715 3717 3741 3838
rect 3852 3717 3874 3838
rect 3715 3689 3874 3717
rect 3945 3838 4104 3860
rect 3945 3717 3971 3838
rect 4082 3717 4104 3838
rect 3945 3689 4104 3717
rect 4175 3838 4334 3860
rect 4175 3717 4201 3838
rect 4312 3717 4334 3838
rect 4175 3689 4334 3717
rect -3789 3603 -3630 3625
rect -3789 3482 -3763 3603
rect -3652 3482 -3630 3603
rect -3789 3454 -3630 3482
rect 4187 3474 4346 3496
rect -3789 3373 -3630 3395
rect -3789 3252 -3763 3373
rect -3652 3252 -3630 3373
rect -3789 3224 -3630 3252
rect 4187 3353 4213 3474
rect 4324 3353 4346 3474
rect 4187 3325 4346 3353
rect -3789 3143 -3630 3165
rect 4187 3244 4346 3266
rect -3789 3022 -3763 3143
rect -3652 3022 -3630 3143
rect 4187 3123 4213 3244
rect 4324 3123 4346 3244
rect 4187 3095 4346 3123
rect -3789 2994 -3630 3022
rect 4187 3014 4346 3036
rect -3789 2913 -3630 2935
rect -3789 2792 -3763 2913
rect -3652 2792 -3630 2913
rect 4187 2893 4213 3014
rect 4324 2893 4346 3014
rect 4187 2865 4346 2893
rect -3789 2764 -3630 2792
rect 4187 2784 4346 2806
rect -2215 2735 -2056 2757
rect -3789 2683 -3630 2705
rect -3789 2562 -3763 2683
rect -3652 2562 -3630 2683
rect -2215 2614 -2189 2735
rect -2078 2614 -2056 2735
rect -2215 2586 -2056 2614
rect -1995 2735 -1836 2757
rect -1995 2614 -1969 2735
rect -1858 2614 -1836 2735
rect -1995 2586 -1836 2614
rect -1775 2735 -1616 2757
rect -1775 2614 -1749 2735
rect -1638 2614 -1616 2735
rect -1775 2586 -1616 2614
rect -1555 2735 -1396 2757
rect -1555 2614 -1529 2735
rect -1418 2614 -1396 2735
rect -1555 2586 -1396 2614
rect -1335 2735 -1176 2757
rect -1335 2614 -1309 2735
rect -1198 2614 -1176 2735
rect -1335 2586 -1176 2614
rect -1115 2735 -956 2757
rect -1115 2614 -1089 2735
rect -978 2614 -956 2735
rect -1115 2586 -956 2614
rect -895 2735 -736 2757
rect -895 2614 -869 2735
rect -758 2614 -736 2735
rect -895 2586 -736 2614
rect -675 2735 -516 2757
rect -675 2614 -649 2735
rect -538 2614 -516 2735
rect -675 2586 -516 2614
rect -455 2735 -296 2757
rect -455 2614 -429 2735
rect -318 2614 -296 2735
rect -455 2586 -296 2614
rect -235 2735 -76 2757
rect -235 2614 -209 2735
rect -98 2614 -76 2735
rect -235 2586 -76 2614
rect -15 2735 144 2757
rect -15 2614 11 2735
rect 122 2614 144 2735
rect -15 2586 144 2614
rect 205 2735 364 2757
rect 205 2614 231 2735
rect 342 2614 364 2735
rect 205 2586 364 2614
rect 425 2735 584 2757
rect 425 2614 451 2735
rect 562 2614 584 2735
rect 425 2586 584 2614
rect 645 2735 804 2757
rect 645 2614 671 2735
rect 782 2614 804 2735
rect 645 2586 804 2614
rect 865 2735 1024 2757
rect 865 2614 891 2735
rect 1002 2614 1024 2735
rect 865 2586 1024 2614
rect 1085 2735 1244 2757
rect 1085 2614 1111 2735
rect 1222 2614 1244 2735
rect 1085 2586 1244 2614
rect 1305 2735 1464 2757
rect 1305 2614 1331 2735
rect 1442 2614 1464 2735
rect 1305 2586 1464 2614
rect 1525 2735 1684 2757
rect 1525 2614 1551 2735
rect 1662 2614 1684 2735
rect 1525 2586 1684 2614
rect 1745 2735 1904 2757
rect 1745 2614 1771 2735
rect 1882 2614 1904 2735
rect 1745 2586 1904 2614
rect 1965 2735 2124 2757
rect 1965 2614 1991 2735
rect 2102 2614 2124 2735
rect 1965 2586 2124 2614
rect 2185 2735 2344 2757
rect 2185 2614 2211 2735
rect 2322 2614 2344 2735
rect 2185 2586 2344 2614
rect 2405 2735 2564 2757
rect 2405 2614 2431 2735
rect 2542 2614 2564 2735
rect 2405 2586 2564 2614
rect 2625 2735 2784 2757
rect 2625 2614 2651 2735
rect 2762 2614 2784 2735
rect 2625 2586 2784 2614
rect 2845 2735 3004 2757
rect 2845 2614 2871 2735
rect 2982 2614 3004 2735
rect 4187 2663 4213 2784
rect 4324 2663 4346 2784
rect 4187 2635 4346 2663
rect 2845 2586 3004 2614
rect -3789 2534 -3630 2562
rect 4187 2554 4346 2576
rect -3789 2453 -3630 2475
rect -3789 2332 -3763 2453
rect -3652 2332 -3630 2453
rect 4187 2433 4213 2554
rect 4324 2433 4346 2554
rect 4187 2405 4346 2433
rect -3789 2304 -3630 2332
rect 4187 2324 4346 2346
rect -3789 2223 -3630 2245
rect -3789 2102 -3763 2223
rect -3652 2102 -3630 2223
rect 4187 2203 4213 2324
rect 4324 2203 4346 2324
rect -3789 2074 -3630 2102
rect 4187 2175 4346 2203
rect 4187 2094 4346 2116
rect -3789 1993 -3630 2015
rect -3789 1872 -3763 1993
rect -3652 1872 -3630 1993
rect 4187 1973 4213 2094
rect 4324 1973 4346 2094
rect 4187 1945 4346 1973
rect -3789 1844 -3630 1872
rect 4187 1864 4346 1886
rect -3789 1763 -3630 1785
rect -3789 1642 -3763 1763
rect -3652 1642 -3630 1763
rect 4187 1743 4213 1864
rect 4324 1743 4346 1864
rect 4187 1715 4346 1743
rect -3789 1614 -3630 1642
rect -2231 1619 -2072 1641
rect -3789 1533 -3630 1555
rect -3789 1412 -3763 1533
rect -3652 1412 -3630 1533
rect -2231 1498 -2205 1619
rect -2094 1498 -2072 1619
rect -2231 1470 -2072 1498
rect -2011 1619 -1852 1641
rect -2011 1498 -1985 1619
rect -1874 1498 -1852 1619
rect -2011 1470 -1852 1498
rect -1791 1619 -1632 1641
rect -1791 1498 -1765 1619
rect -1654 1498 -1632 1619
rect -1791 1470 -1632 1498
rect -1571 1619 -1412 1641
rect -1571 1498 -1545 1619
rect -1434 1498 -1412 1619
rect -1571 1470 -1412 1498
rect -1351 1619 -1192 1641
rect -1351 1498 -1325 1619
rect -1214 1498 -1192 1619
rect -1351 1470 -1192 1498
rect -1131 1619 -972 1641
rect -1131 1498 -1105 1619
rect -994 1498 -972 1619
rect -1131 1470 -972 1498
rect -911 1619 -752 1641
rect -911 1498 -885 1619
rect -774 1498 -752 1619
rect -911 1470 -752 1498
rect -691 1619 -532 1641
rect -691 1498 -665 1619
rect -554 1498 -532 1619
rect -691 1470 -532 1498
rect -471 1619 -312 1641
rect -471 1498 -445 1619
rect -334 1498 -312 1619
rect -471 1470 -312 1498
rect -251 1619 -92 1641
rect -251 1498 -225 1619
rect -114 1498 -92 1619
rect -251 1470 -92 1498
rect -31 1619 128 1641
rect -31 1498 -5 1619
rect 106 1498 128 1619
rect -31 1470 128 1498
rect 189 1619 348 1641
rect 189 1498 215 1619
rect 326 1498 348 1619
rect 189 1470 348 1498
rect 409 1619 568 1641
rect 409 1498 435 1619
rect 546 1498 568 1619
rect 409 1470 568 1498
rect 629 1619 788 1641
rect 629 1498 655 1619
rect 766 1498 788 1619
rect 629 1470 788 1498
rect 849 1619 1008 1641
rect 849 1498 875 1619
rect 986 1498 1008 1619
rect 849 1470 1008 1498
rect 1069 1619 1228 1641
rect 1069 1498 1095 1619
rect 1206 1498 1228 1619
rect 1069 1470 1228 1498
rect 1289 1619 1448 1641
rect 1289 1498 1315 1619
rect 1426 1498 1448 1619
rect 1289 1470 1448 1498
rect 1509 1619 1668 1641
rect 1509 1498 1535 1619
rect 1646 1498 1668 1619
rect 1509 1470 1668 1498
rect 1729 1619 1888 1641
rect 1729 1498 1755 1619
rect 1866 1498 1888 1619
rect 1729 1470 1888 1498
rect 1949 1619 2108 1641
rect 1949 1498 1975 1619
rect 2086 1498 2108 1619
rect 1949 1470 2108 1498
rect 2169 1619 2328 1641
rect 2169 1498 2195 1619
rect 2306 1498 2328 1619
rect 2169 1470 2328 1498
rect 2389 1619 2548 1641
rect 2389 1498 2415 1619
rect 2526 1498 2548 1619
rect 2389 1470 2548 1498
rect 2609 1619 2768 1641
rect 2609 1498 2635 1619
rect 2746 1498 2768 1619
rect 2609 1470 2768 1498
rect 2829 1619 2988 1641
rect 2829 1498 2855 1619
rect 2966 1498 2988 1619
rect 2829 1470 2988 1498
rect 4187 1634 4346 1656
rect 4187 1513 4213 1634
rect 4324 1513 4346 1634
rect 4187 1485 4346 1513
rect -3789 1384 -3630 1412
rect 4187 1404 4346 1426
rect -3789 1303 -3630 1325
rect -3789 1182 -3763 1303
rect -3652 1182 -3630 1303
rect 4187 1283 4213 1404
rect 4324 1283 4346 1404
rect 4187 1255 4346 1283
rect -3789 1154 -3630 1182
rect 4187 1174 4346 1196
rect -3789 1073 -3630 1095
rect -3789 952 -3763 1073
rect -3652 952 -3630 1073
rect 4187 1053 4213 1174
rect 4324 1053 4346 1174
rect 4187 1025 4346 1053
rect -3789 924 -3630 952
rect 4187 944 4346 966
rect -3789 843 -3630 865
rect -3789 722 -3763 843
rect -3652 722 -3630 843
rect 4187 823 4213 944
rect 4324 823 4346 944
rect 4187 795 4346 823
rect -3789 694 -3630 722
rect 4187 714 4346 736
rect -3789 613 -3630 635
rect -3789 492 -3763 613
rect -3652 492 -3630 613
rect 4187 593 4213 714
rect 4324 593 4346 714
rect 4187 565 4346 593
rect -3789 464 -3630 492
rect -876 511 1629 537
rect -876 436 -801 511
rect 1521 436 1629 511
rect -876 413 1629 436
rect 4187 484 4346 506
rect -3789 383 -3630 405
rect -3789 262 -3763 383
rect -3652 262 -3630 383
rect 4187 363 4213 484
rect 4324 363 4346 484
rect 4187 335 4346 363
rect -3789 234 -3630 262
rect -3789 153 -3630 175
rect -3789 32 -3763 153
rect -3652 32 -3630 153
rect -3789 4 -3630 32
rect -3789 -77 -3630 -55
rect -3789 -198 -3763 -77
rect -3652 -198 -3630 -77
rect -3789 -226 -3630 -198
rect -3789 -307 -3630 -285
rect -3789 -428 -3763 -307
rect -3652 -428 -3630 -307
rect 4187 254 4346 276
rect 4187 133 4213 254
rect 4324 133 4346 254
rect 4187 105 4346 133
rect 4187 24 4346 46
rect 4187 -97 4213 24
rect 4324 -97 4346 24
rect 4187 -125 4346 -97
rect 4187 -206 4346 -184
rect 4187 -327 4213 -206
rect 4324 -327 4346 -206
rect 4187 -355 4346 -327
rect -3789 -456 -3630 -428
rect 4187 -436 4346 -414
rect 4187 -557 4213 -436
rect 4324 -557 4346 -436
rect 4187 -585 4346 -557
rect -3733 -623 -3574 -601
rect -3733 -744 -3707 -623
rect -3596 -744 -3574 -623
rect -3733 -772 -3574 -744
rect -3503 -623 -3344 -601
rect -3503 -744 -3477 -623
rect -3366 -744 -3344 -623
rect -3503 -772 -3344 -744
rect -3273 -623 -3114 -601
rect -3273 -744 -3247 -623
rect -3136 -744 -3114 -623
rect -3273 -772 -3114 -744
rect -3043 -623 -2884 -601
rect -3043 -744 -3017 -623
rect -2906 -744 -2884 -623
rect -3043 -772 -2884 -744
rect -2813 -623 -2654 -601
rect -2813 -744 -2787 -623
rect -2676 -744 -2654 -623
rect -2813 -772 -2654 -744
rect -2583 -623 -2424 -601
rect -2583 -744 -2557 -623
rect -2446 -744 -2424 -623
rect -2583 -772 -2424 -744
rect -2353 -623 -2194 -601
rect -2353 -744 -2327 -623
rect -2216 -744 -2194 -623
rect -2353 -772 -2194 -744
rect -2123 -623 -1964 -601
rect -2123 -744 -2097 -623
rect -1986 -744 -1964 -623
rect -2123 -772 -1964 -744
rect -1893 -623 -1734 -601
rect -1893 -744 -1867 -623
rect -1756 -744 -1734 -623
rect -1893 -772 -1734 -744
rect -1663 -623 -1504 -601
rect -1663 -744 -1637 -623
rect -1526 -744 -1504 -623
rect -1663 -772 -1504 -744
rect -1433 -623 -1274 -601
rect -1433 -744 -1407 -623
rect -1296 -744 -1274 -623
rect -1433 -772 -1274 -744
rect -1203 -623 -1044 -601
rect -1203 -744 -1177 -623
rect -1066 -744 -1044 -623
rect -1203 -772 -1044 -744
rect -973 -623 -814 -601
rect -973 -744 -947 -623
rect -836 -744 -814 -623
rect -973 -772 -814 -744
rect -743 -623 -584 -601
rect -743 -744 -717 -623
rect -606 -744 -584 -623
rect -743 -772 -584 -744
rect -513 -623 -354 -601
rect -513 -744 -487 -623
rect -376 -744 -354 -623
rect -513 -772 -354 -744
rect -283 -623 -124 -601
rect -283 -744 -257 -623
rect -146 -744 -124 -623
rect -283 -772 -124 -744
rect -53 -623 106 -601
rect -53 -744 -27 -623
rect 84 -744 106 -623
rect -53 -772 106 -744
rect 177 -623 336 -601
rect 177 -744 203 -623
rect 314 -744 336 -623
rect 177 -772 336 -744
rect 407 -623 566 -601
rect 407 -744 433 -623
rect 544 -744 566 -623
rect 407 -772 566 -744
rect 637 -623 796 -601
rect 637 -744 663 -623
rect 774 -744 796 -623
rect 637 -772 796 -744
rect 867 -623 1026 -601
rect 867 -744 893 -623
rect 1004 -744 1026 -623
rect 867 -772 1026 -744
rect 1097 -623 1256 -601
rect 1097 -744 1123 -623
rect 1234 -744 1256 -623
rect 1097 -772 1256 -744
rect 1327 -623 1486 -601
rect 1327 -744 1353 -623
rect 1464 -744 1486 -623
rect 1327 -772 1486 -744
rect 1557 -623 1716 -601
rect 1557 -744 1583 -623
rect 1694 -744 1716 -623
rect 1557 -772 1716 -744
rect 1787 -623 1946 -601
rect 1787 -744 1813 -623
rect 1924 -744 1946 -623
rect 1787 -772 1946 -744
rect 2017 -623 2176 -601
rect 2017 -744 2043 -623
rect 2154 -744 2176 -623
rect 2017 -772 2176 -744
rect 2247 -623 2406 -601
rect 2247 -744 2273 -623
rect 2384 -744 2406 -623
rect 2247 -772 2406 -744
rect 2477 -623 2636 -601
rect 2477 -744 2503 -623
rect 2614 -744 2636 -623
rect 2477 -772 2636 -744
rect 2707 -623 2866 -601
rect 2707 -744 2733 -623
rect 2844 -744 2866 -623
rect 2707 -772 2866 -744
rect 2937 -623 3096 -601
rect 2937 -744 2963 -623
rect 3074 -744 3096 -623
rect 2937 -772 3096 -744
rect 3167 -623 3326 -601
rect 3167 -744 3193 -623
rect 3304 -744 3326 -623
rect 3167 -772 3326 -744
rect 3397 -623 3556 -601
rect 3397 -744 3423 -623
rect 3534 -744 3556 -623
rect 3397 -772 3556 -744
rect 3627 -623 3786 -601
rect 3627 -744 3653 -623
rect 3764 -744 3786 -623
rect 3627 -772 3786 -744
rect 3857 -623 4016 -601
rect 3857 -744 3883 -623
rect 3994 -744 4016 -623
rect 3857 -772 4016 -744
<< nsubdiff >>
rect -3039 1295 -2922 1309
rect -3039 1202 -3025 1295
rect -2937 1202 -2922 1295
rect -3039 1186 -2922 1202
rect -2829 1295 -2712 1309
rect -2829 1202 -2815 1295
rect -2727 1202 -2712 1295
rect -2829 1186 -2712 1202
rect -2619 1295 -2502 1309
rect -2619 1202 -2605 1295
rect -2517 1202 -2502 1295
rect -2619 1186 -2502 1202
rect -2409 1295 -2292 1309
rect -2409 1202 -2395 1295
rect -2307 1202 -2292 1295
rect -2409 1186 -2292 1202
rect -2199 1295 -2082 1309
rect -2199 1202 -2185 1295
rect -2097 1202 -2082 1295
rect -2199 1186 -2082 1202
rect -1989 1295 -1872 1309
rect -1989 1202 -1975 1295
rect -1887 1202 -1872 1295
rect -1989 1186 -1872 1202
rect -1779 1295 -1662 1309
rect -1779 1202 -1765 1295
rect -1677 1202 -1662 1295
rect -1779 1186 -1662 1202
rect -1569 1295 -1452 1309
rect -1569 1202 -1555 1295
rect -1467 1202 -1452 1295
rect -1569 1186 -1452 1202
rect -1348 1295 -1231 1309
rect -1348 1202 -1334 1295
rect -1246 1202 -1231 1295
rect -1348 1186 -1231 1202
rect -1138 1295 -1021 1309
rect -1138 1202 -1124 1295
rect -1036 1202 -1021 1295
rect -1138 1186 -1021 1202
rect -928 1295 -811 1309
rect -928 1202 -914 1295
rect -826 1202 -811 1295
rect -928 1186 -811 1202
rect -718 1295 -601 1309
rect -718 1202 -704 1295
rect -616 1202 -601 1295
rect -718 1186 -601 1202
rect -508 1295 -391 1309
rect -508 1202 -494 1295
rect -406 1202 -391 1295
rect -508 1186 -391 1202
rect -298 1295 -181 1309
rect -298 1202 -284 1295
rect -196 1202 -181 1295
rect -298 1186 -181 1202
rect -88 1295 29 1309
rect -88 1202 -74 1295
rect 14 1202 29 1295
rect -88 1186 29 1202
rect 122 1295 239 1309
rect 122 1202 136 1295
rect 224 1202 239 1295
rect 122 1186 239 1202
rect 332 1295 449 1309
rect 332 1202 346 1295
rect 434 1202 449 1295
rect 332 1186 449 1202
rect 542 1295 659 1309
rect 542 1202 556 1295
rect 644 1202 659 1295
rect 542 1186 659 1202
rect 752 1295 869 1309
rect 752 1202 766 1295
rect 854 1202 869 1295
rect 752 1186 869 1202
rect 962 1295 1079 1309
rect 962 1202 976 1295
rect 1064 1202 1079 1295
rect 962 1186 1079 1202
rect 1172 1295 1289 1309
rect 1172 1202 1186 1295
rect 1274 1202 1289 1295
rect 1172 1186 1289 1202
rect 1382 1295 1499 1309
rect 1382 1202 1396 1295
rect 1484 1202 1499 1295
rect 1382 1186 1499 1202
rect 1592 1295 1709 1309
rect 1592 1202 1606 1295
rect 1694 1202 1709 1295
rect 1592 1186 1709 1202
rect 1802 1295 1919 1309
rect 1802 1202 1816 1295
rect 1904 1202 1919 1295
rect 1802 1186 1919 1202
rect 2076 1295 2193 1309
rect 2076 1202 2090 1295
rect 2178 1202 2193 1295
rect 2076 1186 2193 1202
rect 2286 1295 2403 1309
rect 2286 1202 2300 1295
rect 2388 1202 2403 1295
rect 2286 1186 2403 1202
rect 2496 1295 2613 1309
rect 2496 1202 2510 1295
rect 2598 1202 2613 1295
rect 2496 1186 2613 1202
rect 2706 1295 2823 1309
rect 2706 1202 2720 1295
rect 2808 1202 2823 1295
rect 2706 1186 2823 1202
rect 2916 1295 3033 1309
rect 2916 1202 2930 1295
rect 3018 1202 3033 1295
rect 2916 1186 3033 1202
rect 3126 1295 3243 1309
rect 3126 1202 3140 1295
rect 3228 1202 3243 1295
rect 3126 1186 3243 1202
rect 3336 1295 3453 1309
rect 3336 1202 3350 1295
rect 3438 1202 3453 1295
rect 3336 1186 3453 1202
rect 3546 1295 3663 1309
rect 3546 1202 3560 1295
rect 3648 1202 3663 1295
rect 3546 1186 3663 1202
rect 3756 1295 3873 1309
rect 3756 1202 3770 1295
rect 3858 1202 3873 1295
rect 3756 1186 3873 1202
<< psubdiffcont >>
rect -3763 3712 -3652 3833
rect -3396 3717 -3285 3838
rect -2937 3717 -2826 3838
rect -2707 3717 -2596 3838
rect -2477 3717 -2366 3838
rect -2247 3717 -2136 3838
rect -2017 3717 -1906 3838
rect -1787 3717 -1676 3838
rect -1557 3717 -1446 3838
rect -1327 3717 -1216 3838
rect -1097 3717 -986 3838
rect -867 3717 -756 3838
rect -637 3717 -526 3838
rect -407 3717 -296 3838
rect -177 3717 -66 3838
rect 53 3717 164 3838
rect 283 3717 394 3838
rect 513 3717 624 3838
rect 743 3717 854 3838
rect 973 3717 1084 3838
rect 1203 3717 1314 3838
rect 1433 3717 1544 3838
rect 1663 3717 1774 3838
rect 1893 3717 2004 3838
rect 2123 3717 2234 3838
rect 2353 3717 2464 3838
rect 2583 3717 2694 3838
rect 2813 3717 2924 3838
rect 3043 3717 3154 3838
rect 3273 3717 3384 3838
rect 3503 3717 3614 3838
rect 3741 3717 3852 3838
rect 3971 3717 4082 3838
rect 4201 3717 4312 3838
rect -3763 3482 -3652 3603
rect -3763 3252 -3652 3373
rect 4213 3353 4324 3474
rect -3763 3022 -3652 3143
rect 4213 3123 4324 3244
rect -3763 2792 -3652 2913
rect 4213 2893 4324 3014
rect -3763 2562 -3652 2683
rect -2189 2614 -2078 2735
rect -1969 2614 -1858 2735
rect -1749 2614 -1638 2735
rect -1529 2614 -1418 2735
rect -1309 2614 -1198 2735
rect -1089 2614 -978 2735
rect -869 2614 -758 2735
rect -649 2614 -538 2735
rect -429 2614 -318 2735
rect -209 2614 -98 2735
rect 11 2614 122 2735
rect 231 2614 342 2735
rect 451 2614 562 2735
rect 671 2614 782 2735
rect 891 2614 1002 2735
rect 1111 2614 1222 2735
rect 1331 2614 1442 2735
rect 1551 2614 1662 2735
rect 1771 2614 1882 2735
rect 1991 2614 2102 2735
rect 2211 2614 2322 2735
rect 2431 2614 2542 2735
rect 2651 2614 2762 2735
rect 2871 2614 2982 2735
rect 4213 2663 4324 2784
rect -3763 2332 -3652 2453
rect 4213 2433 4324 2554
rect -3763 2102 -3652 2223
rect 4213 2203 4324 2324
rect -3763 1872 -3652 1993
rect 4213 1973 4324 2094
rect -3763 1642 -3652 1763
rect 4213 1743 4324 1864
rect -3763 1412 -3652 1533
rect -2205 1498 -2094 1619
rect -1985 1498 -1874 1619
rect -1765 1498 -1654 1619
rect -1545 1498 -1434 1619
rect -1325 1498 -1214 1619
rect -1105 1498 -994 1619
rect -885 1498 -774 1619
rect -665 1498 -554 1619
rect -445 1498 -334 1619
rect -225 1498 -114 1619
rect -5 1498 106 1619
rect 215 1498 326 1619
rect 435 1498 546 1619
rect 655 1498 766 1619
rect 875 1498 986 1619
rect 1095 1498 1206 1619
rect 1315 1498 1426 1619
rect 1535 1498 1646 1619
rect 1755 1498 1866 1619
rect 1975 1498 2086 1619
rect 2195 1498 2306 1619
rect 2415 1498 2526 1619
rect 2635 1498 2746 1619
rect 2855 1498 2966 1619
rect 4213 1513 4324 1634
rect -3763 1182 -3652 1303
rect 4213 1283 4324 1404
rect -3763 952 -3652 1073
rect 4213 1053 4324 1174
rect -3763 722 -3652 843
rect 4213 823 4324 944
rect -3763 492 -3652 613
rect 4213 593 4324 714
rect -801 436 1521 511
rect -3763 262 -3652 383
rect 4213 363 4324 484
rect -3763 32 -3652 153
rect -3763 -198 -3652 -77
rect -3763 -428 -3652 -307
rect 4213 133 4324 254
rect 4213 -97 4324 24
rect 4213 -327 4324 -206
rect 4213 -557 4324 -436
rect -3707 -744 -3596 -623
rect -3477 -744 -3366 -623
rect -3247 -744 -3136 -623
rect -3017 -744 -2906 -623
rect -2787 -744 -2676 -623
rect -2557 -744 -2446 -623
rect -2327 -744 -2216 -623
rect -2097 -744 -1986 -623
rect -1867 -744 -1756 -623
rect -1637 -744 -1526 -623
rect -1407 -744 -1296 -623
rect -1177 -744 -1066 -623
rect -947 -744 -836 -623
rect -717 -744 -606 -623
rect -487 -744 -376 -623
rect -257 -744 -146 -623
rect -27 -744 84 -623
rect 203 -744 314 -623
rect 433 -744 544 -623
rect 663 -744 774 -623
rect 893 -744 1004 -623
rect 1123 -744 1234 -623
rect 1353 -744 1464 -623
rect 1583 -744 1694 -623
rect 1813 -744 1924 -623
rect 2043 -744 2154 -623
rect 2273 -744 2384 -623
rect 2503 -744 2614 -623
rect 2733 -744 2844 -623
rect 2963 -744 3074 -623
rect 3193 -744 3304 -623
rect 3423 -744 3534 -623
rect 3653 -744 3764 -623
rect 3883 -744 3994 -623
<< nsubdiffcont >>
rect -3025 1202 -2937 1295
rect -2815 1202 -2727 1295
rect -2605 1202 -2517 1295
rect -2395 1202 -2307 1295
rect -2185 1202 -2097 1295
rect -1975 1202 -1887 1295
rect -1765 1202 -1677 1295
rect -1555 1202 -1467 1295
rect -1334 1202 -1246 1295
rect -1124 1202 -1036 1295
rect -914 1202 -826 1295
rect -704 1202 -616 1295
rect -494 1202 -406 1295
rect -284 1202 -196 1295
rect -74 1202 14 1295
rect 136 1202 224 1295
rect 346 1202 434 1295
rect 556 1202 644 1295
rect 766 1202 854 1295
rect 976 1202 1064 1295
rect 1186 1202 1274 1295
rect 1396 1202 1484 1295
rect 1606 1202 1694 1295
rect 1816 1202 1904 1295
rect 2090 1202 2178 1295
rect 2300 1202 2388 1295
rect 2510 1202 2598 1295
rect 2720 1202 2808 1295
rect 2930 1202 3018 1295
rect 3140 1202 3228 1295
rect 3350 1202 3438 1295
rect 3560 1202 3648 1295
rect 3770 1202 3858 1295
<< polysilicon >>
rect -2850 3630 3574 3644
rect -2850 3558 -2836 3630
rect -2764 3608 3574 3630
rect -2764 3558 -2750 3608
rect -2850 3515 -2750 3558
rect -2238 3538 -2138 3608
rect -2034 3538 -1934 3608
rect -1422 3538 -1322 3608
rect -1218 3538 -1118 3608
rect -606 3538 -506 3608
rect -402 3538 -302 3608
rect 210 3538 310 3608
rect 414 3538 514 3608
rect 1026 3538 1126 3608
rect 1230 3538 1330 3608
rect 1842 3538 1942 3608
rect 2046 3538 2146 3608
rect 2658 3538 2758 3608
rect 2862 3538 2962 3608
rect 3474 3538 3574 3608
rect -3160 3267 -3058 3288
rect -3160 3210 -3132 3267
rect -3077 3250 -3058 3267
rect -2646 3250 -2546 3356
rect -2442 3250 -2342 3356
rect -1830 3250 -1730 3356
rect -1626 3250 -1526 3356
rect -1014 3250 -914 3356
rect -810 3250 -710 3356
rect -198 3250 -98 3356
rect 6 3250 106 3356
rect 618 3250 718 3356
rect 822 3250 922 3356
rect 1434 3250 1534 3355
rect 1638 3250 1738 3356
rect 2250 3250 2350 3356
rect 2454 3250 2554 3356
rect 3066 3250 3166 3356
rect 3270 3250 3370 3356
rect -3077 3214 3574 3250
rect -3077 3210 -3058 3214
rect -3160 3176 -3058 3210
rect -2850 3144 -2750 3214
rect -2238 3144 -2138 3214
rect -2034 3144 -1934 3214
rect -1422 3144 -1322 3214
rect -1218 3144 -1118 3214
rect -606 3144 -506 3214
rect -402 3144 -302 3214
rect 210 3144 310 3214
rect 414 3144 514 3214
rect 1026 3144 1126 3214
rect 1230 3144 1330 3214
rect 1842 3144 1942 3214
rect 2046 3144 2146 3214
rect 2658 3144 2758 3214
rect 2862 3144 2962 3214
rect 3474 3144 3574 3214
rect -2646 2916 -2546 2936
rect -2646 2844 -2632 2916
rect -2560 2866 -2546 2916
rect -2442 2866 -2342 2936
rect -1830 2866 -1730 2936
rect -1626 2866 -1526 2936
rect -1014 2866 -914 2936
rect -810 2866 -710 2936
rect -198 2866 -98 2936
rect 6 2866 106 2936
rect 618 2866 718 2936
rect 822 2866 922 2936
rect 1434 2866 1534 2936
rect 1638 2866 1738 2936
rect 2250 2866 2350 2936
rect 2454 2866 2554 2936
rect 3066 2866 3166 2936
rect 3270 2916 3370 2936
rect 3270 2866 3284 2916
rect -2560 2844 3284 2866
rect 3356 2844 3370 2916
rect -2646 2830 3370 2844
rect -2107 2495 -2014 2510
rect -2107 2444 -2089 2495
rect -2037 2493 -2014 2495
rect -414 2493 -326 2504
rect 371 2498 486 2517
rect 371 2493 389 2498
rect -2037 2490 389 2493
rect -2037 2457 -400 2490
rect -2037 2444 -2006 2457
rect -2107 2427 -2006 2444
rect -2106 2391 -2006 2427
rect -1494 2391 -1394 2457
rect -1290 2391 -1190 2457
rect -678 2391 -578 2457
rect -414 2430 -400 2457
rect -340 2457 389 2490
rect -340 2430 -238 2457
rect -414 2416 -238 2430
rect -338 2391 -238 2416
rect 274 2441 389 2457
rect 459 2493 486 2498
rect 459 2479 2951 2493
rect 459 2457 1191 2479
rect 459 2441 578 2457
rect 274 2426 578 2441
rect 274 2391 374 2426
rect 478 2391 578 2426
rect 1090 2407 1191 2457
rect 1263 2457 2865 2479
rect 1263 2407 1277 2457
rect 1090 2393 1277 2407
rect 1090 2391 1190 2393
rect 1423 2391 1523 2457
rect 2035 2391 2135 2457
rect 2239 2391 2339 2457
rect 2851 2407 2865 2457
rect 2937 2407 2951 2479
rect 2851 2391 2951 2407
rect -2567 2119 -2474 2135
rect -2567 2059 -2552 2119
rect -2492 2108 -2474 2119
rect -1902 2108 -1802 2199
rect -1698 2108 -1598 2198
rect -1086 2108 -986 2198
rect -882 2108 -782 2199
rect -134 2158 -34 2183
rect -134 2108 -120 2158
rect -2492 2086 -120 2108
rect -48 2108 -34 2158
rect 70 2108 170 2183
rect 682 2158 782 2183
rect 682 2108 696 2158
rect -48 2086 696 2108
rect 768 2108 782 2158
rect 886 2108 986 2183
rect 1627 2108 1727 2183
rect 1831 2108 1931 2184
rect 2443 2108 2543 2183
rect 2647 2108 2747 2184
rect 768 2086 2951 2108
rect -2492 2072 2951 2086
rect -2492 2059 -2474 2072
rect -2567 2041 -2474 2059
rect -2106 2017 -2006 2072
rect -1494 2017 -1394 2072
rect -1290 2017 -1190 2072
rect -678 2017 -578 2072
rect -338 2017 -238 2072
rect 274 2017 373 2072
rect 478 2017 577 2072
rect 1090 2017 1189 2072
rect 1423 2017 1523 2072
rect 2035 2017 2135 2072
rect 2239 2017 2339 2072
rect 2851 2017 2951 2072
rect -1902 1783 -1802 1809
rect -1920 1759 -1802 1783
rect -1920 1709 -1903 1759
rect -1854 1744 -1802 1759
rect -1698 1744 -1598 1845
rect -1086 1744 -986 1845
rect -882 1744 -782 1844
rect -134 1772 -34 1809
rect 70 1772 170 1809
rect -134 1757 170 1772
rect -134 1744 -14 1757
rect -1854 1709 -14 1744
rect -1920 1708 -14 1709
rect -1920 1692 -1832 1708
rect -37 1704 -14 1708
rect 45 1744 170 1757
rect 682 1781 782 1809
rect 886 1781 986 1809
rect 682 1764 986 1781
rect 682 1744 799 1764
rect 45 1708 799 1744
rect 45 1704 74 1708
rect -37 1689 74 1704
rect 779 1706 799 1708
rect 866 1744 986 1764
rect 1627 1744 1727 1809
rect 1831 1744 1931 1809
rect 2443 1744 2543 1809
rect 2647 1744 2747 1810
rect 866 1708 2747 1744
rect 866 1706 892 1708
rect 779 1687 892 1706
rect 3688 1141 3788 1142
rect -3084 1127 3788 1141
rect -3084 1104 -1202 1127
rect -3084 1054 -2984 1104
rect -2472 1054 -2372 1104
rect -2268 1054 -2168 1104
rect -1656 1054 -1556 1104
rect -1216 1055 -1202 1104
rect -1130 1104 1858 1127
rect -1130 1055 -1116 1104
rect -1216 1041 -1116 1055
rect -604 1054 -504 1104
rect -400 1054 -300 1104
rect 212 1054 312 1104
rect 416 1054 516 1104
rect 1028 1054 1128 1104
rect 1232 1054 1332 1104
rect 1844 1055 1858 1104
rect 1930 1104 3788 1127
rect 1930 1055 1944 1104
rect 1844 1041 1944 1055
rect 2260 1054 2360 1104
rect 2872 1054 2972 1104
rect 3076 1054 3176 1104
rect 3688 1054 3788 1104
rect -2880 790 -2780 846
rect -2676 790 -2576 883
rect -2064 790 -1964 882
rect -1860 790 -1760 881
rect -1012 839 -912 853
rect -1012 790 -998 839
rect -2880 767 -998 790
rect -926 790 -912 839
rect -808 790 -708 846
rect -196 790 -96 846
rect 8 790 108 846
rect 620 790 720 846
rect 824 790 924 846
rect 1436 790 1536 846
rect 1640 839 1740 853
rect 1640 790 1654 839
rect -926 767 1654 790
rect 1726 790 1740 839
rect 2464 790 2564 878
rect 2668 790 2768 878
rect 3280 790 3380 878
rect 3484 790 3584 878
rect 1726 767 3584 790
rect -2880 753 3584 767
rect -2637 288 3188 324
rect -2637 -193 -2537 288
rect -2433 -353 -2333 77
rect -2229 -353 -2129 221
rect -2025 -220 -1925 288
rect -1684 232 -1584 288
rect -1072 232 -972 288
rect -740 232 -640 288
rect -204 283 764 288
rect -204 188 -104 283
rect 663 229 764 283
rect 1200 280 3188 288
rect 1200 232 1300 280
rect 1532 232 1632 280
rect 2144 232 2244 280
rect -204 24 137 27
rect -1684 -94 -1584 24
rect -1480 -94 -1380 24
rect -1276 -94 -1176 24
rect -1072 -94 -972 24
rect -740 -94 -640 24
rect -536 -94 -436 24
rect -204 -4 228 24
rect -204 -42 109 -4
rect 45 -61 109 -42
rect 175 -61 228 -4
rect 45 -79 228 -61
rect 128 -94 228 -79
rect 332 -9 432 24
rect 332 -81 346 -9
rect 403 -81 432 -9
rect 332 -94 432 -81
rect 996 -94 1096 24
rect 1200 -94 1300 24
rect 1532 -94 1632 24
rect 1736 -94 1836 24
rect 1940 -94 2040 24
rect 2144 -94 2244 24
rect 332 -95 417 -94
rect 2476 -117 2576 280
rect -1480 -353 -1380 -301
rect -1276 -353 -1176 -302
rect -536 -353 -436 -302
rect -2433 -354 -436 -353
rect -204 -354 -104 -302
rect 332 -354 432 -302
rect -2433 -356 432 -354
rect 664 -356 764 -302
rect 996 -352 1096 -302
rect 1736 -352 1836 -302
rect 1940 -352 2040 -302
rect 2680 -352 2780 60
rect 2884 -352 2984 92
rect 3088 -112 3188 280
rect 996 -356 2984 -352
rect -2433 -399 2984 -356
<< polycontact >>
rect -2836 3558 -2764 3630
rect -3132 3210 -3077 3267
rect -2632 2844 -2560 2916
rect 3284 2844 3356 2916
rect -2089 2444 -2037 2495
rect -400 2430 -340 2490
rect 389 2441 459 2498
rect 1191 2407 1263 2479
rect 2865 2407 2937 2479
rect -2552 2059 -2492 2119
rect -120 2086 -48 2158
rect 696 2086 768 2158
rect -1903 1709 -1854 1759
rect -14 1704 45 1757
rect 799 1706 866 1764
rect -1202 1055 -1130 1127
rect 1858 1055 1930 1127
rect -998 767 -926 839
rect 1654 767 1726 839
rect 109 -61 175 -4
rect 346 -81 403 -9
<< metal1 >>
rect -3789 3838 4358 3860
rect -3789 3833 -3396 3838
rect -3789 3712 -3763 3833
rect -3652 3717 -3396 3833
rect -3285 3717 -2937 3838
rect -2826 3717 -2707 3838
rect -2596 3717 -2477 3838
rect -2366 3717 -2247 3838
rect -2136 3717 -2017 3838
rect -1906 3717 -1787 3838
rect -1676 3717 -1557 3838
rect -1446 3717 -1327 3838
rect -1216 3717 -1097 3838
rect -986 3717 -867 3838
rect -756 3717 -637 3838
rect -526 3717 -407 3838
rect -296 3717 -177 3838
rect -66 3717 53 3838
rect 164 3717 283 3838
rect 394 3717 513 3838
rect 624 3717 743 3838
rect 854 3717 973 3838
rect 1084 3717 1203 3838
rect 1314 3717 1433 3838
rect 1544 3717 1663 3838
rect 1774 3717 1893 3838
rect 2004 3717 2123 3838
rect 2234 3717 2353 3838
rect 2464 3717 2583 3838
rect 2694 3717 2813 3838
rect 2924 3717 3043 3838
rect 3154 3717 3273 3838
rect 3384 3717 3503 3838
rect 3614 3817 3741 3838
rect 3667 3739 3741 3817
rect 3614 3717 3741 3739
rect 3852 3717 3971 3838
rect 4082 3717 4201 3838
rect 4312 3717 4358 3838
rect -3652 3712 4358 3717
rect -3789 3689 4358 3712
rect -3789 3603 -3618 3689
rect -3789 3482 -3763 3603
rect -3652 3482 -3618 3603
rect -2845 3630 -2755 3639
rect -2845 3558 -2836 3630
rect -2764 3558 -2755 3630
rect -2845 3549 -2755 3558
rect -2517 3483 -2471 3689
rect -1701 3492 -1655 3689
rect -885 3492 -839 3689
rect -69 3492 -23 3689
rect 747 3492 793 3689
rect 1563 3492 1609 3689
rect 2379 3492 2425 3689
rect 3195 3492 3241 3689
rect -3789 3373 -3618 3482
rect -2740 3462 -2654 3477
rect -2740 3405 -2727 3462
rect -2670 3405 -2654 3462
rect -2740 3394 -2654 3405
rect -2334 3464 -2248 3479
rect -2334 3407 -2321 3464
rect -2264 3407 -2248 3464
rect -2334 3396 -2248 3407
rect -1929 3465 -1843 3480
rect -1929 3408 -1916 3465
rect -1859 3408 -1843 3465
rect -1929 3397 -1843 3408
rect -1523 3461 -1437 3476
rect -1523 3404 -1510 3461
rect -1453 3404 -1437 3461
rect -1523 3393 -1437 3404
rect -1112 3467 -1026 3482
rect -1112 3410 -1099 3467
rect -1042 3410 -1026 3467
rect -1112 3399 -1026 3410
rect -704 3464 -618 3479
rect -704 3407 -691 3464
rect -634 3407 -618 3464
rect -704 3396 -618 3407
rect -294 3466 -208 3481
rect -294 3409 -281 3466
rect -224 3409 -208 3466
rect -294 3398 -208 3409
rect 115 3467 201 3482
rect 115 3410 128 3467
rect 185 3410 201 3467
rect 115 3399 201 3410
rect 521 3467 607 3482
rect 521 3410 534 3467
rect 591 3410 607 3467
rect 521 3399 607 3410
rect 930 3465 1016 3480
rect 930 3408 943 3465
rect 1000 3408 1016 3465
rect 930 3397 1016 3408
rect 1336 3470 1422 3485
rect 1336 3413 1349 3470
rect 1406 3413 1422 3470
rect 1336 3402 1422 3413
rect 1749 3470 1835 3485
rect 1749 3413 1762 3470
rect 1819 3413 1835 3470
rect 1749 3402 1835 3413
rect 2153 3467 2239 3482
rect 2153 3410 2166 3467
rect 2223 3410 2239 3467
rect 2153 3399 2239 3410
rect 2560 3465 2646 3480
rect 2560 3408 2573 3465
rect 2630 3408 2646 3465
rect 2560 3397 2646 3408
rect 2968 3464 3054 3479
rect 2968 3407 2981 3464
rect 3038 3407 3054 3464
rect 2968 3396 3054 3407
rect 3377 3464 3463 3479
rect 3377 3407 3390 3464
rect 3447 3407 3463 3464
rect 3377 3396 3463 3407
rect 4187 3474 4358 3689
rect -3789 3252 -3763 3373
rect -3652 3252 -3618 3373
rect -2925 3317 -2879 3376
rect -2109 3317 -2063 3377
rect -1293 3317 -1247 3377
rect -477 3317 -431 3377
rect 339 3317 385 3376
rect 1155 3317 1201 3376
rect 1971 3317 2017 3377
rect 2787 3317 2833 3377
rect 3603 3317 3649 3377
rect 4187 3353 4213 3474
rect 4324 3353 4358 3474
rect -3789 3143 -3618 3252
rect -3160 3267 -3058 3288
rect -3160 3210 -3132 3267
rect -3077 3210 -3058 3267
rect -2925 3229 3826 3317
rect 4187 3244 4358 3353
rect -3160 3176 -3058 3210
rect -3789 3022 -3763 3143
rect -3652 3022 -3618 3143
rect -3789 2913 -3618 3022
rect -3789 2792 -3763 2913
rect -3652 2792 -3618 2913
rect -3789 2683 -3618 2792
rect -3789 2562 -3763 2683
rect -3652 2562 -3618 2683
rect -3789 2453 -3618 2562
rect -3789 2332 -3763 2453
rect -3652 2332 -3618 2453
rect -3789 2223 -3618 2332
rect -3789 2102 -3763 2223
rect -3652 2102 -3618 2223
rect -3789 1993 -3618 2102
rect -3152 2118 -3078 3176
rect -2517 3098 -2471 3229
rect -1701 3098 -1655 3229
rect -885 3098 -839 3229
rect -69 3098 -23 3229
rect 747 3098 793 3229
rect 1563 3098 1609 3229
rect 2379 3098 2425 3229
rect 3195 3098 3241 3229
rect 4187 3123 4213 3244
rect 4324 3123 4358 3244
rect -2742 3073 -2656 3088
rect -2742 3016 -2729 3073
rect -2672 3016 -2656 3073
rect -2742 3005 -2656 3016
rect -2335 3073 -2249 3088
rect -2335 3016 -2322 3073
rect -2265 3016 -2249 3073
rect -2335 3005 -2249 3016
rect -1929 3071 -1843 3086
rect -1929 3014 -1916 3071
rect -1859 3014 -1843 3071
rect -1929 3003 -1843 3014
rect -1520 3073 -1434 3088
rect -1520 3016 -1507 3073
rect -1450 3016 -1434 3073
rect -1520 3005 -1434 3016
rect -1113 3069 -1027 3084
rect -1113 3012 -1100 3069
rect -1043 3012 -1027 3069
rect -1113 3001 -1027 3012
rect -706 3072 -620 3087
rect -706 3015 -693 3072
rect -636 3015 -620 3072
rect -706 3004 -620 3015
rect -296 3073 -210 3088
rect -296 3016 -283 3073
rect -226 3016 -210 3073
rect -296 3005 -210 3016
rect 114 3070 200 3085
rect 114 3013 127 3070
rect 184 3013 200 3070
rect 114 3002 200 3013
rect 521 3069 607 3084
rect 521 3012 534 3069
rect 591 3012 607 3069
rect 521 3001 607 3012
rect 930 3071 1016 3086
rect 930 3014 943 3071
rect 1000 3014 1016 3071
rect 930 3003 1016 3014
rect 1336 3076 1422 3091
rect 1336 3019 1349 3076
rect 1406 3019 1422 3076
rect 1336 3008 1422 3019
rect 1744 3074 1830 3089
rect 1744 3017 1757 3074
rect 1814 3017 1830 3074
rect 1744 3006 1830 3017
rect 2153 3073 2239 3088
rect 2153 3016 2166 3073
rect 2223 3016 2239 3073
rect 2153 3005 2239 3016
rect 2561 3072 2647 3087
rect 2561 3015 2574 3072
rect 2631 3015 2647 3072
rect 2561 3004 2647 3015
rect 2970 3075 3056 3090
rect 2970 3018 2983 3075
rect 3040 3018 3056 3075
rect 2970 3007 3056 3018
rect 3378 3072 3464 3087
rect 3378 3015 3391 3072
rect 3448 3015 3464 3072
rect 3378 3004 3464 3015
rect 4187 3014 4358 3123
rect -2925 2695 -2879 2982
rect -2641 2916 -2551 2925
rect -2641 2844 -2632 2916
rect -2560 2844 -2551 2916
rect -2641 2835 -2551 2844
rect -2109 2757 -2063 2982
rect -1293 2757 -1247 2982
rect -477 2757 -431 2982
rect 339 2757 385 2982
rect 1155 2757 1201 2982
rect 1971 2757 2017 2982
rect 2787 2757 2833 2982
rect 3275 2916 3365 2925
rect 3275 2844 3284 2916
rect 3356 2844 3365 2916
rect 3275 2835 3365 2844
rect -2215 2735 3060 2757
rect 3603 2739 3649 2982
rect 4187 2893 4213 3014
rect 4324 2893 4358 3014
rect 4187 2784 4358 2893
rect -2215 2698 -2189 2735
rect -2370 2695 -2189 2698
rect -2925 2649 -2189 2695
rect -2370 2626 -2189 2649
rect -2567 2119 -2474 2135
rect -2567 2118 -2552 2119
rect -3152 2059 -2552 2118
rect -2492 2059 -2474 2119
rect -3152 2044 -2474 2059
rect -2567 2041 -2474 2044
rect -3789 1872 -3763 1993
rect -3652 1872 -3618 1993
rect -3789 1763 -3618 1872
rect -3789 1642 -3763 1763
rect -3652 1642 -3618 1763
rect -3789 1533 -3618 1642
rect -2370 1613 -2298 2626
rect -2215 2614 -2189 2626
rect -2078 2614 -1969 2735
rect -1858 2614 -1749 2735
rect -1638 2614 -1529 2735
rect -1418 2614 -1309 2735
rect -1198 2614 -1089 2735
rect -978 2614 -869 2735
rect -758 2614 -649 2735
rect -538 2614 -429 2735
rect -318 2614 -209 2735
rect -98 2614 11 2735
rect 122 2614 231 2735
rect 342 2614 451 2735
rect 562 2614 671 2735
rect 782 2614 891 2735
rect 1002 2614 1111 2735
rect 1222 2614 1331 2735
rect 1442 2614 1551 2735
rect 1662 2614 1771 2735
rect 1882 2614 1991 2735
rect 2102 2614 2211 2735
rect 2322 2614 2431 2735
rect 2542 2614 2651 2735
rect 2762 2614 2871 2735
rect 2982 2717 3060 2735
rect 3572 2717 3689 2739
rect 2982 2716 3689 2717
rect 2982 2640 3590 2716
rect 3666 2640 3689 2716
rect 2982 2639 3689 2640
rect 2982 2614 3060 2639
rect 3572 2627 3689 2639
rect 4187 2663 4213 2784
rect 4324 2663 4358 2784
rect -2215 2586 3060 2614
rect -2107 2495 -2014 2510
rect -2107 2494 -2089 2495
rect -2107 2438 -2091 2494
rect -2037 2494 -2014 2495
rect -2035 2438 -2014 2494
rect -2107 2427 -2014 2438
rect -1773 2345 -1727 2586
rect -957 2345 -911 2586
rect -419 2499 -343 2502
rect -578 2485 -489 2496
rect -578 2431 -561 2485
rect -507 2482 -489 2485
rect -419 2493 -331 2499
rect -419 2482 -410 2493
rect -354 2490 -331 2493
rect -507 2437 -410 2482
rect -507 2433 -400 2437
rect -507 2431 -489 2433
rect -578 2424 -489 2431
rect -419 2430 -400 2433
rect -340 2430 -331 2490
rect -419 2421 -331 2430
rect -419 2417 -343 2421
rect -1998 2323 -1913 2336
rect -1998 2270 -1984 2323
rect -1927 2270 -1913 2323
rect -1998 2255 -1913 2270
rect -1590 2317 -1505 2330
rect -1590 2264 -1576 2317
rect -1519 2264 -1505 2317
rect -1590 2249 -1505 2264
rect -1184 2321 -1099 2334
rect -1184 2268 -1170 2321
rect -1113 2268 -1099 2321
rect -1184 2253 -1099 2268
rect -777 2317 -692 2330
rect -777 2264 -763 2317
rect -706 2264 -692 2317
rect -777 2249 -692 2264
rect -2181 2169 -2135 2238
rect -414 2237 -365 2417
rect -5 2345 41 2586
rect 371 2498 486 2517
rect 371 2441 389 2498
rect 459 2441 486 2498
rect 371 2426 486 2441
rect 403 2345 449 2426
rect 811 2345 857 2586
rect 1182 2479 1272 2488
rect 1182 2407 1191 2479
rect 1263 2407 1272 2479
rect 1182 2398 1272 2407
rect 1219 2345 1265 2398
rect 1756 2345 1802 2586
rect 2572 2345 2618 2586
rect 4187 2554 4358 2663
rect 2856 2479 2946 2488
rect 2856 2407 2865 2479
rect 2937 2407 2946 2479
rect 2856 2398 2946 2407
rect 4187 2433 4213 2554
rect 4324 2433 4358 2554
rect -226 2312 -149 2325
rect -226 2255 -214 2312
rect -162 2255 -149 2312
rect -226 2244 -149 2255
rect 179 2313 256 2326
rect 179 2256 191 2313
rect 243 2256 256 2313
rect 179 2245 256 2256
rect 587 2322 664 2335
rect 587 2265 599 2322
rect 651 2265 664 2322
rect 587 2254 664 2265
rect 993 2317 1070 2330
rect 993 2260 1005 2317
rect 1057 2260 1070 2317
rect 993 2249 1070 2260
rect 1529 2318 1614 2331
rect 1529 2265 1543 2318
rect 1600 2265 1614 2318
rect 1529 2250 1614 2265
rect 1937 2319 2022 2332
rect 1937 2266 1951 2319
rect 2008 2266 2022 2319
rect 1937 2251 2022 2266
rect 2347 2322 2432 2335
rect 2347 2269 2361 2322
rect 2418 2269 2432 2322
rect 2347 2254 2432 2269
rect 2752 2322 2837 2335
rect 2752 2269 2766 2322
rect 2823 2269 2837 2322
rect 2752 2254 2837 2269
rect 4187 2324 4358 2433
rect -1365 2169 -1319 2233
rect -2206 2147 -882 2169
rect -2206 2093 -961 2147
rect -907 2143 -882 2147
rect -549 2143 -503 2233
rect 1348 2169 1394 2233
rect 2164 2169 2210 2233
rect 2980 2169 3026 2229
rect 4187 2203 4213 2324
rect 4324 2203 4358 2324
rect 1332 2167 3198 2169
rect -907 2097 -503 2143
rect -129 2158 -39 2167
rect -907 2093 -882 2097
rect -2206 2072 -882 2093
rect -129 2086 -120 2158
rect -48 2086 -39 2158
rect -129 2077 -39 2086
rect 687 2158 777 2167
rect 687 2086 696 2158
rect 768 2086 777 2158
rect 687 2077 777 2086
rect 1330 2148 3198 2167
rect 1330 2092 1352 2148
rect 1408 2092 3198 2148
rect 1330 2072 3198 2092
rect 4187 2094 4358 2203
rect -1773 1971 -1727 2072
rect -980 2070 -883 2072
rect 1330 2070 1427 2072
rect -957 1971 -911 2070
rect 1756 1971 1802 2072
rect 2572 1971 2618 2072
rect 4187 1973 4213 2094
rect 4324 1973 4358 2094
rect -1998 1949 -1913 1962
rect -1998 1896 -1984 1949
rect -1927 1896 -1913 1949
rect -1998 1881 -1913 1896
rect -1591 1945 -1506 1958
rect -1591 1892 -1577 1945
rect -1520 1892 -1506 1945
rect -1591 1877 -1506 1892
rect -1184 1944 -1099 1957
rect -1184 1891 -1170 1944
rect -1113 1891 -1099 1944
rect -1184 1876 -1099 1891
rect -777 1944 -692 1957
rect -777 1891 -763 1944
rect -706 1891 -692 1944
rect -777 1876 -692 1891
rect -226 1944 -149 1957
rect -226 1887 -214 1944
rect -162 1887 -149 1944
rect -226 1876 -149 1887
rect 173 1947 250 1960
rect 173 1890 185 1947
rect 237 1890 250 1947
rect 173 1879 250 1890
rect 585 1942 662 1955
rect 585 1885 597 1942
rect 649 1885 662 1942
rect 585 1874 662 1885
rect 993 1940 1070 1953
rect 993 1883 1005 1940
rect 1057 1883 1070 1940
rect 993 1872 1070 1883
rect 1526 1942 1611 1955
rect 1526 1889 1540 1942
rect 1597 1889 1611 1942
rect 1526 1874 1611 1889
rect 1937 1946 2022 1959
rect 1937 1893 1951 1946
rect 2008 1893 2022 1946
rect 1937 1878 2022 1893
rect 2345 1946 2430 1959
rect 2345 1893 2359 1946
rect 2416 1893 2430 1946
rect 2345 1878 2430 1893
rect 2756 1948 2841 1961
rect 2756 1895 2770 1948
rect 2827 1895 2841 1948
rect 2756 1880 2841 1895
rect 4187 1864 4358 1973
rect -2181 1641 -2135 1858
rect -1924 1762 -1832 1783
rect -1924 1699 -1912 1762
rect -1851 1699 -1832 1762
rect -1924 1689 -1832 1699
rect -1365 1641 -1319 1855
rect -549 1641 -503 1855
rect -413 1641 -367 1857
rect -6 1780 41 1855
rect -17 1772 41 1780
rect -37 1771 74 1772
rect -37 1715 -16 1771
rect 40 1757 74 1771
rect -37 1704 -14 1715
rect 45 1704 74 1757
rect -37 1689 74 1704
rect 403 1641 449 1855
rect 811 1781 857 1855
rect 779 1764 892 1781
rect 779 1758 799 1764
rect 866 1758 892 1764
rect 779 1706 798 1758
rect 874 1706 892 1758
rect 779 1687 892 1706
rect 1219 1641 1265 1855
rect 1348 1641 1394 1855
rect 2164 1641 2210 1855
rect 2980 1641 3026 1855
rect 4187 1743 4213 1864
rect 4324 1743 4358 1864
rect -2231 1619 3044 1641
rect -2231 1613 -2205 1619
rect -2370 1541 -2205 1613
rect -3789 1412 -3763 1533
rect -3652 1412 -3618 1533
rect -2231 1498 -2205 1541
rect -2094 1498 -1985 1619
rect -1874 1498 -1765 1619
rect -1654 1498 -1545 1619
rect -1434 1498 -1325 1619
rect -1214 1498 -1105 1619
rect -994 1498 -885 1619
rect -774 1498 -665 1619
rect -554 1498 -445 1619
rect -334 1498 -225 1619
rect -114 1498 -5 1619
rect 106 1498 215 1619
rect 326 1498 435 1619
rect 546 1498 655 1619
rect 766 1498 875 1619
rect 986 1498 1095 1619
rect 1206 1498 1315 1619
rect 1426 1498 1535 1619
rect 1646 1498 1755 1619
rect 1866 1498 1975 1619
rect 2086 1498 2195 1619
rect 2306 1498 2415 1619
rect 2526 1498 2635 1619
rect 2746 1498 2855 1619
rect 2966 1604 3044 1619
rect 4187 1634 4358 1743
rect 4187 1604 4213 1634
rect 2966 1526 4213 1604
rect 2966 1498 3044 1526
rect -2231 1470 3044 1498
rect 4187 1513 4213 1526
rect 4324 1513 4358 1634
rect -3789 1303 -3618 1412
rect 4187 1404 4358 1513
rect -3789 1182 -3763 1303
rect -3652 1182 -3618 1303
rect -3258 1295 3962 1350
rect -3258 1202 -3025 1295
rect -2937 1202 -2815 1295
rect -2727 1202 -2605 1295
rect -2517 1202 -2395 1295
rect -2307 1202 -2185 1295
rect -2097 1202 -1975 1295
rect -1887 1202 -1765 1295
rect -1677 1202 -1555 1295
rect -1467 1202 -1334 1295
rect -1246 1268 -1124 1295
rect -1227 1214 -1124 1268
rect -1246 1202 -1124 1214
rect -1036 1202 -914 1295
rect -826 1202 -704 1295
rect -616 1202 -494 1295
rect -406 1202 -284 1295
rect -196 1202 -74 1295
rect 14 1202 136 1295
rect 224 1290 346 1295
rect 224 1236 329 1290
rect 224 1202 346 1236
rect 434 1202 556 1295
rect 644 1202 766 1295
rect 854 1202 976 1295
rect 1064 1278 1186 1295
rect 1064 1224 1157 1278
rect 1064 1202 1186 1224
rect 1274 1202 1396 1295
rect 1484 1202 1606 1295
rect 1694 1202 1816 1295
rect 1904 1278 2090 1295
rect 1904 1224 1977 1278
rect 2030 1224 2090 1278
rect 1904 1202 2090 1224
rect 2178 1202 2300 1295
rect 2388 1202 2510 1295
rect 2598 1202 2720 1295
rect 2808 1202 2930 1295
rect 3018 1202 3140 1295
rect 3228 1202 3350 1295
rect 3438 1202 3560 1295
rect 3648 1202 3770 1295
rect 3858 1202 3962 1295
rect -3258 1186 3962 1202
rect 4187 1283 4213 1404
rect 4324 1283 4358 1404
rect -3789 1073 -3618 1182
rect -3789 952 -3763 1073
rect -3652 952 -3618 1073
rect -3159 1008 -3113 1186
rect -2343 1008 -2297 1186
rect -1750 1000 -1660 1010
rect -1527 1008 -1481 1186
rect -1198 1136 -1152 1138
rect -1211 1127 -1121 1136
rect -1211 1055 -1202 1127
rect -1130 1109 -1121 1127
rect 1849 1127 1939 1136
rect 1849 1109 1858 1127
rect -1130 1063 1858 1109
rect -1130 1055 -1041 1063
rect -1211 1046 -1041 1055
rect -1087 1006 -1041 1046
rect -679 1008 -633 1063
rect -271 1008 -225 1063
rect 137 1008 183 1063
rect 545 1008 591 1063
rect 953 1008 999 1063
rect 1361 1008 1407 1063
rect 1769 1055 1858 1063
rect 1930 1055 1939 1127
rect 1769 1046 1939 1055
rect 1769 1008 1815 1046
rect 2185 1008 2231 1186
rect 3001 1008 3047 1186
rect 3817 1008 3863 1186
rect 4187 1174 4358 1283
rect 4187 1053 4213 1174
rect 4324 1053 4358 1174
rect -3789 843 -3618 952
rect -2979 985 -2898 995
rect -2979 932 -2968 985
rect -2915 932 -2898 985
rect -2979 919 -2898 932
rect -2562 990 -2481 1000
rect -2562 937 -2551 990
rect -2498 937 -2481 990
rect -2562 924 -2481 937
rect -2152 990 -2071 1000
rect -2152 937 -2141 990
rect -2088 937 -2071 990
rect -2152 924 -2071 937
rect -1750 930 -1740 1000
rect -1670 930 -1660 1000
rect -1750 920 -1660 930
rect -1303 970 -1224 983
rect -1303 916 -1291 970
rect -1238 916 -1224 970
rect -1303 904 -1224 916
rect -499 970 -420 983
rect -499 916 -487 970
rect -434 916 -420 970
rect 320 972 399 985
rect -499 904 -420 916
rect -3789 722 -3763 843
rect -3652 722 -3618 843
rect -2751 837 -2705 892
rect -1935 837 -1889 892
rect -883 848 -837 895
rect -1007 839 -837 848
rect -1011 838 -998 839
rect -3789 613 -3618 722
rect -3789 492 -3763 613
rect -3652 492 -3618 613
rect -3150 816 -1125 837
rect -3150 812 -2925 816
rect -3150 758 -3112 812
rect -3058 762 -2925 812
rect -2871 762 -1125 816
rect -1011 782 -1002 838
rect -926 828 -837 839
rect -67 828 -21 938
rect 320 918 332 972
rect 385 918 399 972
rect 1135 973 1214 986
rect 320 906 399 918
rect 749 828 795 938
rect 1135 919 1147 973
rect 1200 919 1214 973
rect 1135 907 1214 919
rect 1955 974 2034 987
rect 1955 920 1967 974
rect 2020 920 2034 974
rect 1955 908 2034 920
rect 2373 983 2454 993
rect 2373 930 2384 983
rect 2437 930 2454 983
rect 2373 917 2454 930
rect 2780 981 2861 991
rect 2780 928 2791 981
rect 2844 928 2861 981
rect 2780 915 2861 928
rect 3187 981 3268 991
rect 3187 928 3198 981
rect 3251 928 3268 981
rect 3187 915 3268 928
rect 3592 981 3673 991
rect 3592 928 3603 981
rect 3656 928 3673 981
rect 3592 915 3673 928
rect 4187 944 4358 1053
rect 1565 848 1611 892
rect 1565 839 1735 848
rect 1565 828 1654 839
rect -926 782 1654 828
rect -1011 781 -998 782
rect -3058 758 -1125 762
rect -1007 767 -998 781
rect -926 767 -917 782
rect -1007 758 -917 767
rect 1645 767 1654 782
rect 1726 767 1735 839
rect 1645 758 1735 767
rect 2593 842 2639 892
rect 3409 842 3455 892
rect 2593 796 3455 842
rect 4187 823 4213 944
rect 4324 823 4358 944
rect -3150 733 -1125 758
rect 2593 757 3453 796
rect -3150 707 -1047 733
rect 2593 707 2653 757
rect -3150 697 2653 707
rect -3150 684 -2797 697
rect -3150 653 -2800 684
rect -1253 657 2653 697
rect 4187 714 4358 823
rect -3150 651 -2888 653
rect -3150 597 -3121 651
rect -3067 599 -2888 651
rect -2834 599 -2800 653
rect -3067 597 -2800 599
rect -3150 570 -2800 597
rect -2730 600 -2646 615
rect -2730 546 -2716 600
rect -2662 546 -2646 600
rect 3185 601 3269 618
rect -2730 532 -2646 546
rect -2392 564 -1034 565
rect -967 564 -919 565
rect -151 564 -100 565
rect 664 564 718 565
rect 1484 564 1532 565
rect 1711 564 2913 565
rect -3789 383 -3618 492
rect -3789 262 -3763 383
rect -3652 262 -3618 383
rect -3789 153 -3618 262
rect -3789 32 -3763 153
rect -3652 32 -3618 153
rect -3789 -77 -3618 32
rect -3789 -198 -3763 -77
rect -3652 -198 -3618 -77
rect -3789 -307 -3618 -198
rect -3789 -428 -3763 -307
rect -3652 -428 -3618 -307
rect -2712 -320 -2666 532
rect -2392 511 2913 564
rect 3185 545 3198 601
rect 3254 545 3269 601
rect 3185 535 3269 545
rect 4187 593 4213 714
rect 4324 593 4358 714
rect -2392 436 -801 511
rect 1521 461 2913 511
rect 3025 461 3117 472
rect 1521 460 3166 461
rect 1521 436 3033 460
rect -2392 381 3033 436
rect -2508 9 -2462 70
rect -2525 -4 -2450 9
rect -2525 -58 -2512 -4
rect -2458 -58 -2450 -4
rect -2525 -68 -2450 -58
rect -2508 -140 -2462 -68
rect -2304 -140 -2258 381
rect -1776 259 -1695 271
rect -1776 205 -1762 259
rect -1708 205 -1695 259
rect -1776 193 -1695 205
rect -2100 9 -2054 70
rect -2115 -3 -2040 9
rect -2115 -57 -2104 -3
rect -2050 -57 -2040 -3
rect -2115 -69 -2040 -57
rect -2100 -140 -2054 -69
rect -1896 -320 -1850 70
rect -2712 -366 -1850 -320
rect -1760 -317 -1711 193
rect -1559 -7 -1503 190
rect -1568 -16 -1494 -7
rect -1568 -72 -1559 -16
rect -1503 -72 -1494 -16
rect -1568 -80 -1494 -72
rect -1560 -81 -1502 -80
rect -1559 -261 -1503 -81
rect -1354 -261 -1298 381
rect -1152 -4 -1097 186
rect -1158 -16 -1085 -4
rect -1158 -72 -1150 -16
rect -1094 -72 -1085 -16
rect -1158 -81 -1085 -72
rect -1152 -260 -1097 -81
rect -948 -317 -894 187
rect -1760 -366 -894 -317
rect -818 -404 -766 191
rect -615 -9 -562 190
rect -625 -26 -545 -9
rect -625 -80 -615 -26
rect -561 -80 -545 -26
rect -625 -94 -545 -80
rect -615 -263 -562 -94
rect -3789 -601 -3618 -428
rect -833 -412 -751 -404
rect -833 -466 -819 -412
rect -765 -466 -751 -412
rect -833 -476 -751 -466
rect -408 -522 -358 381
rect 37 320 108 332
rect 37 266 49 320
rect 103 266 108 320
rect 37 253 108 266
rect -283 -268 -231 188
rect -81 16 -25 190
rect 52 72 99 253
rect 255 70 306 187
rect -92 13 -22 16
rect -92 -41 -80 13
rect -26 -41 -22 13
rect -92 -55 -22 -41
rect 46 -4 186 8
rect 46 -61 109 -4
rect 175 -61 186 -4
rect 46 -78 186 -61
rect 254 -9 412 0
rect -298 -271 -218 -268
rect -298 -325 -284 -271
rect -230 -325 -218 -271
rect -298 -331 -218 -325
rect -81 -323 -29 -135
rect 46 -258 103 -78
rect 254 -81 346 -9
rect 403 -81 412 -9
rect 254 -90 412 -81
rect 254 -259 305 -90
rect 458 -323 516 381
rect 580 18 643 193
rect 576 14 650 18
rect 576 -42 583 14
rect 639 -42 650 14
rect 576 -55 650 -42
rect 585 -323 638 -131
rect 791 -258 841 223
rect -81 -369 638 -323
rect 785 -270 858 -258
rect 917 -264 972 381
rect 1118 -32 1175 190
rect 1099 -41 1180 -32
rect 1099 -97 1115 -41
rect 1171 -97 1180 -41
rect 1099 -106 1180 -97
rect 1118 -260 1175 -106
rect 785 -326 789 -270
rect 845 -326 858 -270
rect 785 -339 858 -326
rect -81 -370 -28 -369
rect 1325 -372 1376 209
rect 1453 -301 1505 192
rect 1658 15 1710 189
rect 1644 10 1725 15
rect 1644 -46 1657 10
rect 1713 -46 1725 10
rect 1644 -55 1725 -46
rect 1658 -262 1710 -55
rect 1861 -258 1913 381
rect 2809 380 3033 381
rect 3113 380 3166 460
rect 2809 379 3166 380
rect 2268 260 2341 273
rect 2268 204 2278 260
rect 2334 204 2341 260
rect 2065 23 2117 188
rect 2268 185 2341 204
rect 2059 10 2132 23
rect 2059 -46 2067 10
rect 2123 -46 2132 10
rect 2059 -58 2132 -46
rect 2065 -263 2117 -58
rect 1453 -337 1589 -301
rect 2270 -337 2321 185
rect 1453 -353 2321 -337
rect 2401 -304 2447 70
rect 2605 6 2651 70
rect 2591 -5 2663 6
rect 2591 -59 2601 -5
rect 2655 -59 2663 -5
rect 2591 -68 2663 -59
rect 2605 -140 2651 -68
rect 2809 -140 2855 379
rect 3025 372 3117 379
rect 3013 5 3059 70
rect 3000 -4 3072 5
rect 3000 -58 3009 -4
rect 3063 -58 3072 -4
rect 3000 -69 3072 -58
rect 3013 -140 3059 -69
rect 3217 -304 3263 535
rect 4187 484 4358 593
rect 3344 461 3448 472
rect 4187 461 4213 484
rect 3311 379 3354 461
rect 3436 379 4213 461
rect 3344 370 3448 379
rect 2401 -350 3263 -304
rect 4187 363 4213 379
rect 4324 363 4358 484
rect 4187 254 4358 363
rect 4187 133 4213 254
rect 4324 133 4358 254
rect 4187 24 4358 133
rect 4187 -97 4213 24
rect 4324 -97 4358 24
rect 4187 -206 4358 -97
rect 4187 -327 4213 -206
rect 4324 -327 4358 -206
rect 1325 -382 1409 -372
rect 1325 -438 1341 -382
rect 1397 -438 1409 -382
rect 1537 -389 2321 -353
rect 1325 -439 1409 -438
rect 4187 -436 4358 -327
rect 4187 -557 4213 -436
rect 4324 -557 4358 -436
rect 4187 -601 4358 -557
rect -3789 -623 4358 -601
rect -3789 -744 -3707 -623
rect -3596 -744 -3477 -623
rect -3366 -744 -3247 -623
rect -3136 -744 -3017 -623
rect -2906 -744 -2787 -623
rect -2676 -744 -2557 -623
rect -2446 -744 -2327 -623
rect -2216 -744 -2097 -623
rect -1986 -744 -1867 -623
rect -1756 -744 -1637 -623
rect -1526 -744 -1407 -623
rect -1296 -744 -1177 -623
rect -1066 -744 -947 -623
rect -836 -744 -717 -623
rect -606 -744 -487 -623
rect -376 -744 -257 -623
rect -146 -744 -27 -623
rect 84 -744 203 -623
rect 314 -744 433 -623
rect 544 -744 663 -623
rect 774 -744 893 -623
rect 1004 -744 1123 -623
rect 1234 -744 1353 -623
rect 1464 -744 1583 -623
rect 1694 -744 1813 -623
rect 1924 -744 2043 -623
rect 2154 -744 2273 -623
rect 2384 -744 2503 -623
rect 2614 -744 2733 -623
rect 2844 -744 2963 -623
rect 3074 -744 3193 -623
rect 3304 -744 3423 -623
rect 3534 -744 3653 -623
rect 3764 -744 3883 -623
rect 3994 -744 4358 -623
rect -3789 -772 4358 -744
<< via1 >>
rect 3589 3739 3614 3817
rect 3614 3739 3667 3817
rect -2829 3566 -2772 3622
rect -2727 3405 -2670 3462
rect -2321 3407 -2264 3464
rect -1916 3408 -1859 3465
rect -1510 3404 -1453 3461
rect -1099 3410 -1042 3467
rect -691 3407 -634 3464
rect -281 3409 -224 3466
rect 128 3410 185 3467
rect 534 3410 591 3467
rect 943 3408 1000 3465
rect 1349 3413 1406 3470
rect 1762 3413 1819 3470
rect 2166 3410 2223 3467
rect 2573 3408 2630 3465
rect 2981 3407 3038 3464
rect 3390 3407 3447 3464
rect -2729 3016 -2672 3073
rect -2322 3016 -2265 3073
rect -1916 3014 -1859 3071
rect -1507 3016 -1450 3073
rect -1100 3012 -1043 3069
rect -693 3015 -636 3072
rect -283 3016 -226 3073
rect 127 3013 184 3070
rect 534 3012 591 3069
rect 943 3014 1000 3071
rect 1349 3019 1406 3076
rect 1757 3017 1814 3074
rect 2166 3016 2223 3073
rect 2574 3015 2631 3072
rect 2983 3018 3040 3075
rect 3391 3015 3448 3072
rect -2629 2848 -2570 2907
rect 3291 2851 3346 2905
rect 3590 2640 3666 2716
rect -2091 2444 -2089 2494
rect -2089 2444 -2037 2495
rect -2037 2444 -2035 2494
rect -2091 2438 -2035 2444
rect -561 2431 -507 2485
rect -410 2490 -354 2493
rect -410 2437 -400 2490
rect -400 2437 -354 2490
rect -1984 2270 -1927 2323
rect -1576 2264 -1519 2317
rect -1170 2268 -1113 2321
rect -763 2264 -706 2317
rect 2874 2416 2929 2471
rect -214 2255 -162 2312
rect 191 2256 243 2313
rect 599 2265 651 2322
rect 1005 2260 1057 2317
rect 1543 2265 1600 2318
rect 1951 2266 2008 2319
rect 2361 2269 2418 2322
rect 2766 2269 2823 2322
rect -961 2093 -907 2147
rect -108 2092 -52 2148
rect 702 2092 758 2148
rect 1352 2092 1408 2148
rect -1984 1896 -1927 1949
rect -1577 1892 -1520 1945
rect -1170 1891 -1113 1944
rect -763 1891 -706 1944
rect -214 1887 -162 1944
rect 185 1890 237 1947
rect 597 1885 649 1942
rect 1005 1883 1057 1940
rect 1540 1889 1597 1942
rect 1951 1893 2008 1946
rect 2359 1893 2416 1946
rect 2770 1895 2827 1948
rect -1912 1759 -1851 1762
rect -1912 1709 -1903 1759
rect -1903 1709 -1854 1759
rect -1854 1709 -1851 1759
rect -1912 1699 -1851 1709
rect -16 1757 40 1771
rect -16 1715 -14 1757
rect -14 1715 40 1757
rect 798 1706 799 1758
rect 799 1706 866 1758
rect 866 1706 874 1758
rect -1280 1214 -1246 1268
rect -1246 1214 -1227 1268
rect -479 1216 -426 1270
rect 329 1236 346 1290
rect 346 1236 382 1290
rect 1157 1224 1186 1278
rect 1186 1224 1210 1278
rect 1977 1224 2030 1278
rect -2968 932 -2915 985
rect -2551 937 -2498 990
rect -2141 937 -2088 990
rect -1740 930 -1670 1000
rect -1291 916 -1238 970
rect -487 916 -434 970
rect -3112 758 -3058 812
rect -2925 762 -2871 816
rect -1002 782 -998 838
rect -998 782 -946 838
rect 332 918 385 972
rect 1147 919 1200 973
rect 1967 920 2020 974
rect 2384 930 2437 983
rect 2791 928 2844 981
rect 3198 928 3251 981
rect 3603 928 3656 981
rect 1667 778 1723 834
rect -3121 597 -3067 651
rect -2888 599 -2834 653
rect -2716 546 -2662 600
rect 3198 545 3254 601
rect -2512 -58 -2458 -4
rect -1762 205 -1708 259
rect -2104 -57 -2050 -3
rect -1559 -72 -1503 -16
rect -1150 -72 -1094 -16
rect -615 -80 -561 -26
rect -819 -466 -765 -412
rect 49 266 103 320
rect -80 -41 -26 13
rect -284 -325 -230 -271
rect 583 -42 639 14
rect 1115 -97 1171 -41
rect 789 -326 845 -270
rect 1657 -46 1713 10
rect 3033 380 3113 460
rect 2278 204 2334 260
rect 2067 -46 2123 10
rect 2601 -59 2655 -5
rect 3009 -58 3063 -4
rect 3354 379 3436 461
rect 1341 -438 1397 -382
<< metal2 >>
rect 3580 3817 3674 3833
rect 3580 3739 3589 3817
rect 3667 3739 3674 3817
rect 3580 3725 3674 3739
rect -2909 3622 -2755 3639
rect -2909 3566 -2829 3622
rect -2772 3566 -2755 3622
rect -2909 3549 -2755 3566
rect -2909 2932 -2818 3549
rect -2740 3462 -2654 3477
rect -2740 3405 -2727 3462
rect -2670 3458 -2654 3462
rect -2334 3464 -2248 3479
rect -2334 3458 -2321 3464
rect -2670 3407 -2321 3458
rect -2264 3458 -2248 3464
rect -1929 3465 -1843 3480
rect -1929 3458 -1916 3465
rect -2264 3408 -1916 3458
rect -1859 3458 -1843 3465
rect -1523 3461 -1437 3476
rect -1523 3458 -1510 3461
rect -1859 3408 -1510 3458
rect -2264 3407 -1510 3408
rect -2670 3405 -1510 3407
rect -2740 3404 -1510 3405
rect -1453 3458 -1437 3461
rect -1112 3467 -1026 3482
rect -1112 3458 -1099 3467
rect -1453 3410 -1099 3458
rect -1042 3458 -1026 3467
rect -704 3464 -618 3479
rect -704 3458 -691 3464
rect -1042 3410 -691 3458
rect -1453 3407 -691 3410
rect -634 3458 -618 3464
rect -294 3466 -208 3481
rect -294 3458 -281 3466
rect -634 3409 -281 3458
rect -224 3458 -208 3466
rect 115 3467 201 3482
rect 115 3458 128 3467
rect -224 3410 128 3458
rect 185 3458 201 3467
rect 521 3467 607 3482
rect 521 3458 534 3467
rect 185 3410 534 3458
rect 591 3458 607 3467
rect 930 3465 1016 3480
rect 930 3458 943 3465
rect 591 3410 943 3458
rect -224 3409 943 3410
rect -634 3408 943 3409
rect 1000 3458 1016 3465
rect 1336 3470 1422 3485
rect 1336 3458 1349 3470
rect 1000 3413 1349 3458
rect 1406 3458 1422 3470
rect 1749 3470 1835 3485
rect 1749 3458 1762 3470
rect 1406 3413 1762 3458
rect 1819 3458 1835 3470
rect 2153 3467 2239 3482
rect 2153 3458 2166 3467
rect 1819 3413 2166 3458
rect 1000 3410 2166 3413
rect 2223 3458 2239 3467
rect 2560 3465 2646 3480
rect 2560 3458 2573 3465
rect 2223 3410 2573 3458
rect 1000 3408 2573 3410
rect 2630 3458 2646 3465
rect 2968 3464 3054 3479
rect 2968 3458 2981 3464
rect 2630 3408 2981 3458
rect -634 3407 2981 3408
rect 3038 3458 3054 3464
rect 3377 3464 3463 3479
rect 3377 3458 3390 3464
rect 3038 3407 3390 3458
rect 3447 3407 3463 3464
rect -1453 3404 3463 3407
rect -2740 3402 3463 3404
rect -2740 3394 -2654 3402
rect -2334 3396 -2248 3402
rect -1929 3397 -1843 3402
rect -2733 3088 -2677 3394
rect -2323 3088 -2267 3396
rect -2742 3073 -2656 3088
rect -2742 3016 -2729 3073
rect -2672 3016 -2656 3073
rect -2742 3005 -2656 3016
rect -2335 3073 -2249 3088
rect -1918 3086 -1862 3397
rect -1523 3393 -1437 3402
rect -1112 3399 -1026 3402
rect -1508 3088 -1452 3393
rect -2335 3016 -2322 3073
rect -2265 3016 -2249 3073
rect -2335 3005 -2249 3016
rect -1929 3071 -1843 3086
rect -1929 3014 -1916 3071
rect -1859 3014 -1843 3071
rect -1929 3003 -1843 3014
rect -1520 3073 -1434 3088
rect -1101 3084 -1045 3399
rect -704 3396 -618 3402
rect -294 3398 -208 3402
rect 115 3399 201 3402
rect 521 3399 607 3402
rect -695 3087 -639 3396
rect -282 3088 -226 3398
rect -1520 3016 -1507 3073
rect -1450 3016 -1434 3073
rect -1520 3005 -1434 3016
rect -1113 3069 -1027 3084
rect -1113 3012 -1100 3069
rect -1043 3012 -1027 3069
rect -1113 3001 -1027 3012
rect -706 3072 -620 3087
rect -706 3015 -693 3072
rect -636 3015 -620 3072
rect -706 3004 -620 3015
rect -296 3073 -210 3088
rect 119 3085 175 3399
rect -296 3016 -283 3073
rect -226 3016 -210 3073
rect -296 3005 -210 3016
rect 114 3070 200 3085
rect 529 3084 585 3399
rect 930 3397 1016 3402
rect 936 3086 992 3397
rect 1347 3091 1403 3402
rect 114 3013 127 3070
rect 184 3013 200 3070
rect 114 3002 200 3013
rect 521 3069 607 3084
rect 521 3012 534 3069
rect 591 3012 607 3069
rect 521 3001 607 3012
rect 930 3071 1016 3086
rect 930 3014 943 3071
rect 1000 3014 1016 3071
rect 930 3003 1016 3014
rect 1336 3076 1422 3091
rect 1754 3089 1810 3402
rect 2153 3399 2239 3402
rect 1336 3019 1349 3076
rect 1406 3019 1422 3076
rect 1336 3008 1422 3019
rect 1744 3074 1830 3089
rect 2165 3088 2221 3399
rect 2560 3397 2646 3402
rect 1744 3017 1757 3074
rect 1814 3017 1830 3074
rect 1744 3006 1830 3017
rect 2153 3073 2239 3088
rect 2576 3087 2632 3397
rect 2968 3396 3054 3402
rect 3377 3396 3463 3402
rect 2983 3090 3039 3396
rect 2153 3016 2166 3073
rect 2223 3016 2239 3073
rect 2153 3005 2239 3016
rect 2561 3072 2647 3087
rect 2561 3015 2574 3072
rect 2631 3015 2647 3072
rect 2561 3004 2647 3015
rect 2970 3075 3056 3090
rect 3397 3087 3453 3396
rect 2970 3018 2983 3075
rect 3040 3018 3056 3075
rect 2970 3007 3056 3018
rect 3378 3072 3464 3087
rect 3378 3015 3391 3072
rect 3448 3015 3464 3072
rect 3378 3004 3464 3015
rect -2909 2907 -2551 2932
rect 3317 2925 3395 2926
rect -2909 2848 -2629 2907
rect -2570 2848 -2551 2907
rect -2909 2841 -2551 2848
rect -2647 2835 -2551 2841
rect 3275 2905 3395 2925
rect 3275 2851 3291 2905
rect 3346 2851 3395 2905
rect 3275 2835 3395 2851
rect -2647 2503 -2556 2835
rect -773 2622 1599 2678
rect -2107 2503 -2014 2510
rect -2647 2495 -2014 2503
rect -2647 2494 -2089 2495
rect -2037 2494 -2014 2495
rect -2647 2438 -2091 2494
rect -2035 2438 -2014 2494
rect -2647 2412 -2014 2438
rect -2256 1782 -2104 2412
rect -1998 2330 -1913 2336
rect -1184 2330 -1099 2334
rect -773 2330 -717 2622
rect -581 2493 -343 2502
rect -581 2485 -410 2493
rect -581 2431 -561 2485
rect -507 2437 -410 2485
rect -354 2437 -343 2493
rect -507 2431 -343 2437
rect -581 2417 -343 2431
rect -1998 2323 -692 2330
rect -1998 2270 -1984 2323
rect -1927 2321 -692 2323
rect -1927 2317 -1170 2321
rect -1927 2274 -1576 2317
rect -1927 2270 -1913 2274
rect -1998 2255 -1913 2270
rect -1590 2264 -1576 2274
rect -1519 2274 -1170 2317
rect -1519 2264 -1505 2274
rect -1980 1962 -1924 2255
rect -1590 2249 -1505 2264
rect -1184 2268 -1170 2274
rect -1113 2317 -692 2321
rect -1113 2274 -763 2317
rect -1113 2268 -1099 2274
rect -1184 2253 -1099 2268
rect -777 2264 -763 2274
rect -706 2264 -692 2317
rect -1998 1949 -1913 1962
rect -1577 1958 -1521 2249
rect -1998 1896 -1984 1949
rect -1927 1896 -1913 1949
rect -1998 1881 -1913 1896
rect -1591 1945 -1506 1958
rect -1176 1957 -1120 2253
rect -777 2249 -692 2264
rect -980 2148 -883 2167
rect -980 2092 -962 2148
rect -906 2092 -883 2148
rect -980 2070 -883 2092
rect -773 1957 -717 2249
rect -1591 1892 -1577 1945
rect -1520 1892 -1506 1945
rect -1591 1877 -1506 1892
rect -1184 1944 -1099 1957
rect -1184 1891 -1170 1944
rect -1113 1891 -1099 1944
rect -1184 1876 -1099 1891
rect -777 1944 -692 1957
rect -777 1891 -763 1944
rect -706 1891 -692 1944
rect -777 1876 -692 1891
rect -1924 1782 -1832 1783
rect -3355 1762 -1802 1782
rect -3355 1699 -1912 1762
rect -1851 1699 -1802 1762
rect -3355 1611 -1802 1699
rect -581 1737 -354 2417
rect -226 2317 -149 2325
rect 179 2317 256 2326
rect 587 2322 664 2335
rect 1543 2331 1599 2622
rect 2856 2484 2946 2488
rect 3290 2484 3395 2835
rect 3589 2739 3667 3725
rect 3572 2716 3689 2739
rect 3572 2640 3590 2716
rect 3666 2640 3689 2716
rect 3572 2627 3689 2640
rect 2856 2471 3395 2484
rect 2856 2416 2874 2471
rect 2929 2416 3395 2471
rect 2856 2406 3395 2416
rect 2856 2398 2946 2406
rect 587 2317 599 2322
rect -226 2313 599 2317
rect -226 2312 191 2313
rect -226 2255 -214 2312
rect -162 2261 191 2312
rect -162 2255 -149 2261
rect -226 2244 -149 2255
rect 179 2256 191 2261
rect 243 2265 599 2313
rect 651 2317 664 2322
rect 993 2317 1070 2330
rect 651 2265 1005 2317
rect 243 2261 1005 2265
rect 243 2256 256 2261
rect 179 2245 256 2256
rect 587 2254 664 2261
rect 991 2260 1005 2261
rect 1057 2260 1070 2317
rect -209 2170 -153 2244
rect -209 2148 -40 2170
rect -209 2092 -108 2148
rect -52 2092 -40 2148
rect -209 2080 -40 2092
rect -209 1957 -153 2080
rect 182 1960 238 2245
rect 602 2166 658 2254
rect 991 2249 1070 2260
rect 1529 2318 1614 2331
rect 1529 2265 1543 2318
rect 1600 2316 1614 2318
rect 1937 2319 2022 2332
rect 1937 2316 1951 2319
rect 1600 2266 1951 2316
rect 2008 2315 2022 2319
rect 2347 2322 2432 2335
rect 2347 2315 2361 2322
rect 2008 2269 2361 2315
rect 2418 2314 2432 2322
rect 2752 2322 2837 2335
rect 2752 2314 2766 2322
rect 2418 2269 2766 2314
rect 2823 2269 2837 2322
rect 2008 2266 2837 2269
rect 1600 2265 2837 2266
rect 1529 2257 2837 2265
rect 1529 2250 1614 2257
rect 1937 2251 2022 2257
rect 2347 2254 2432 2257
rect 2752 2254 2837 2257
rect 602 2148 776 2166
rect 602 2092 702 2148
rect 758 2092 776 2148
rect 602 2078 776 2092
rect -226 1944 -149 1957
rect -226 1887 -214 1944
rect -162 1887 -149 1944
rect -226 1876 -149 1887
rect 173 1947 250 1960
rect 602 1955 658 2078
rect 173 1890 185 1947
rect 237 1890 250 1947
rect 173 1879 250 1890
rect 585 1942 662 1955
rect 585 1885 597 1942
rect 649 1885 662 1942
rect 585 1874 662 1885
rect 991 1953 1047 2249
rect 1330 2148 1427 2167
rect 1330 2092 1352 2148
rect 1408 2092 1427 2148
rect 1330 2070 1427 2092
rect 1544 1955 1602 2250
rect 1944 1959 2000 2251
rect 2366 1959 2422 2254
rect 2769 1961 2825 2254
rect 991 1940 1070 1953
rect 991 1883 1005 1940
rect 1057 1883 1070 1940
rect 991 1877 1070 1883
rect 993 1872 1070 1877
rect 1526 1942 1611 1955
rect 1526 1889 1540 1942
rect 1597 1889 1611 1942
rect 1526 1874 1611 1889
rect 1937 1946 2022 1959
rect 1937 1893 1951 1946
rect 2008 1893 2022 1946
rect 1937 1878 2022 1893
rect 2345 1946 2430 1959
rect 2345 1893 2359 1946
rect 2416 1893 2430 1946
rect 2345 1878 2430 1893
rect 2756 1948 2841 1961
rect 2756 1895 2770 1948
rect 2827 1895 2841 1948
rect 2756 1880 2841 1895
rect -37 1779 73 1785
rect 780 1779 888 1780
rect -54 1771 941 1779
rect -54 1737 -16 1771
rect -581 1715 -16 1737
rect 40 1758 941 1771
rect 40 1715 798 1758
rect -581 1706 798 1715
rect 874 1706 941 1758
rect -581 1611 941 1706
rect -3355 1495 941 1611
rect -3355 836 -3068 1495
rect -1728 1361 2446 1417
rect -1728 1010 -1672 1361
rect 317 1290 396 1303
rect -1292 1268 -1213 1281
rect -1292 1222 -1280 1268
rect -1296 1214 -1280 1222
rect -1227 1214 -1213 1268
rect -1296 1202 -1213 1214
rect -491 1270 -412 1283
rect -491 1216 -479 1270
rect -426 1216 -412 1270
rect 317 1236 329 1290
rect 382 1236 396 1290
rect 317 1224 396 1236
rect 1145 1278 1224 1291
rect 1145 1224 1157 1278
rect 1210 1224 1224 1278
rect -491 1204 -412 1216
rect -1750 1000 -1660 1010
rect -2979 986 -2898 995
rect -2562 990 -2481 1000
rect -2562 986 -2551 990
rect -2979 985 -2551 986
rect -2979 932 -2968 985
rect -2915 937 -2551 985
rect -2498 986 -2481 990
rect -2152 990 -2071 1000
rect -2152 986 -2141 990
rect -2498 937 -2141 986
rect -2088 986 -2071 990
rect -1750 986 -1740 1000
rect -2088 937 -1740 986
rect -2915 932 -1740 937
rect -2979 930 -1740 932
rect -1670 930 -1660 1000
rect -1296 983 -1232 1202
rect -488 983 -424 1204
rect 329 985 393 1224
rect 1145 1212 1224 1224
rect 1965 1278 2044 1291
rect 1965 1224 1977 1278
rect 2030 1224 2044 1278
rect 1965 1212 2044 1224
rect 1149 986 1213 1212
rect 1971 987 2035 1212
rect 2390 993 2446 1361
rect -2979 919 -2898 930
rect -2562 924 -2481 930
rect -2152 924 -2071 930
rect -1750 920 -1660 930
rect -1303 970 -1224 983
rect -1303 916 -1291 970
rect -1238 916 -1224 970
rect -1303 904 -1224 916
rect -499 970 -420 983
rect -499 916 -487 970
rect -434 916 -420 970
rect -499 904 -420 916
rect 320 972 399 985
rect 320 918 332 972
rect 385 918 399 972
rect 320 906 399 918
rect 1135 973 1214 986
rect 1135 919 1147 973
rect 1200 919 1214 973
rect 1135 907 1214 919
rect 1955 984 2035 987
rect 1955 974 2034 984
rect 1955 920 1967 974
rect 2020 920 2034 974
rect 1955 908 2034 920
rect 2373 983 2454 993
rect 2373 930 2384 983
rect 2437 980 2454 983
rect 2780 981 2861 991
rect 2780 980 2791 981
rect 2437 930 2791 980
rect 2373 928 2791 930
rect 2844 980 2861 981
rect 3187 981 3268 991
rect 3187 980 3198 981
rect 2844 928 3198 980
rect 3251 980 3268 981
rect 3592 981 3673 991
rect 3592 980 3603 981
rect 3251 928 3603 980
rect 3656 928 3673 981
rect 2373 924 3673 928
rect 2373 917 2454 924
rect 2780 915 2861 924
rect 3187 915 3268 924
rect 3592 915 3673 924
rect -1012 838 -912 847
rect -3355 816 -2810 836
rect -3355 812 -2925 816
rect -3355 758 -3112 812
rect -3058 762 -2925 812
rect -2871 762 -2810 816
rect -3058 758 -2810 762
rect -3355 653 -2810 758
rect -1012 782 -1002 838
rect -946 782 -912 838
rect -1012 753 -912 782
rect 1638 834 1738 849
rect 1638 778 1667 834
rect 1723 778 1738 834
rect 1638 755 1738 778
rect -3355 651 -2888 653
rect -3355 597 -3121 651
rect -3067 599 -2888 651
rect -2834 599 -2810 653
rect -3067 597 -2810 599
rect -3355 576 -2810 597
rect -2730 601 -2646 615
rect -1002 601 -946 753
rect 1667 601 1723 755
rect 3185 601 3269 618
rect -2730 600 3198 601
rect -3355 571 -3068 576
rect -2730 546 -2716 600
rect -2662 546 3198 600
rect -2730 545 3198 546
rect 3254 545 3269 601
rect -2730 532 -2646 545
rect 3185 535 3269 545
rect 2140 476 2265 484
rect 2140 460 2153 476
rect -1747 404 2153 460
rect -1747 271 -1691 404
rect 2140 389 2153 404
rect 2240 460 2265 476
rect 3025 461 3117 472
rect 3344 461 3448 472
rect 3025 460 3354 461
rect 2240 389 2317 460
rect 2140 378 2317 389
rect -1776 259 -1691 271
rect -1776 205 -1762 259
rect -1708 205 -1691 259
rect 37 321 108 332
rect 2010 321 2078 331
rect 37 320 2012 321
rect 37 266 49 320
rect 103 266 2012 320
rect 37 265 2012 266
rect 2068 265 2078 321
rect 37 253 108 265
rect 2010 255 2078 265
rect 2261 273 2317 378
rect 3025 380 3033 460
rect 3113 380 3354 460
rect 3025 379 3354 380
rect 3436 379 3448 461
rect 3025 372 3117 379
rect 3344 370 3448 379
rect 2261 260 2341 273
rect -1776 198 -1691 205
rect 2261 204 2278 260
rect 2334 204 2343 260
rect -1776 193 -1695 198
rect 2261 187 2341 204
rect 2268 185 2341 187
rect -907 90 1713 146
rect -2525 -2 -2450 9
rect -2115 -2 -2040 9
rect -2525 -3 -2040 -2
rect -2525 -4 -2104 -3
rect -2525 -58 -2512 -4
rect -2458 -57 -2104 -4
rect -2050 -57 -2040 -3
rect -2458 -58 -2040 -57
rect -2525 -68 -2450 -58
rect -2115 -69 -2040 -58
rect -1568 -16 -1494 -7
rect -1158 -16 -1085 -4
rect -907 -16 -851 90
rect -92 14 -22 16
rect 575 14 651 18
rect 1657 15 1713 90
rect -92 13 583 14
rect -2113 -573 -2057 -69
rect -1568 -72 -1559 -16
rect -1503 -72 -1150 -16
rect -1094 -72 -851 -16
rect -625 -25 -545 -9
rect -625 -26 -350 -25
rect -1568 -81 -1494 -72
rect -1158 -81 -1085 -72
rect -625 -80 -615 -26
rect -561 -80 -350 -26
rect -92 -41 -80 13
rect -26 -41 583 13
rect -92 -42 583 -41
rect 639 -42 651 14
rect 1647 10 1725 15
rect 2059 10 2132 23
rect 1099 -41 1180 -32
rect -92 -55 -22 -42
rect 575 -55 651 -42
rect -625 -81 -350 -80
rect -625 -94 -545 -81
rect -406 -128 -350 -81
rect 837 -97 1115 -41
rect 1171 -97 1180 -41
rect 1647 -46 1657 10
rect 1713 -46 2067 10
rect 2123 -46 2132 10
rect 2591 -4 2663 6
rect 3000 -4 3072 5
rect 2591 -5 3009 -4
rect 2591 -15 2601 -5
rect 1647 -55 1725 -46
rect 2059 -58 2132 -46
rect 837 -128 893 -97
rect 1099 -106 1180 -97
rect 2574 -59 2601 -15
rect 2655 -58 3009 -5
rect 3063 -58 3072 -4
rect 2655 -59 3072 -58
rect 2574 -60 3072 -59
rect 2574 -68 2663 -60
rect -406 -184 893 -128
rect -300 -270 -216 -258
rect 785 -270 858 -258
rect -300 -271 789 -270
rect -300 -325 -284 -271
rect -230 -325 789 -271
rect -300 -326 789 -325
rect 845 -326 858 -270
rect -300 -342 -216 -326
rect 785 -339 858 -326
rect 1325 -382 1409 -372
rect -827 -412 -753 -404
rect -827 -466 -819 -412
rect -765 -417 -753 -412
rect 1325 -417 1341 -382
rect -765 -438 1341 -417
rect 1397 -417 1409 -382
rect 2273 -417 2345 -407
rect 1397 -438 2283 -417
rect -765 -466 2283 -438
rect -827 -473 2283 -466
rect 2339 -473 2345 -417
rect -827 -481 -753 -473
rect 2273 -486 2345 -473
rect 2574 -573 2630 -68
rect 3000 -69 3072 -60
rect -2113 -629 2630 -573
<< via2 >>
rect -962 2147 -906 2148
rect -962 2093 -961 2147
rect -961 2093 -907 2147
rect -907 2093 -906 2147
rect -962 2092 -906 2093
rect 1352 2092 1408 2148
rect 2153 389 2240 476
rect 2012 265 2068 321
rect 583 -42 639 14
rect 2283 -473 2339 -417
<< metal3 >>
rect -980 2148 -883 2167
rect 1330 2148 1427 2167
rect -980 2092 -962 2148
rect -906 2092 1352 2148
rect 1408 2092 1427 2148
rect -980 2070 -883 2092
rect 1330 2070 1427 2092
rect 583 25 639 565
rect 2153 484 2240 485
rect 2140 476 2265 484
rect 2140 389 2153 476
rect 2240 471 2265 476
rect 2240 401 2490 471
rect 2240 389 2265 401
rect 2140 378 2265 389
rect 2010 321 2078 331
rect 2010 265 2012 321
rect 2068 265 2490 321
rect 2010 255 2078 265
rect 574 14 652 25
rect 574 -42 583 14
rect 639 -42 652 14
rect 574 -54 652 -42
rect 574 -55 651 -54
rect 2273 -417 2345 -407
rect 2273 -473 2283 -417
rect 2339 -473 2495 -417
rect 2273 -486 2345 -473
use nmos_3p3_9NPLV7  nmos_3p3_9NPLV7_0
timestamp 1693373438
transform 1 0 362 0 1 3434
box -3324 -128 3324 128
use nmos_3p3_9NPLV7  nmos_3p3_9NPLV7_1
timestamp 1693373438
transform 1 0 362 0 1 3040
box -3324 -128 3324 128
use nmos_3p3_AJEA3B  nmos_3p3_AJEA3B_0
timestamp 1693304636
transform 1 0 2187 0 1 2287
box -876 -128 876 128
use nmos_3p3_AJEA3B  nmos_3p3_AJEA3B_1
timestamp 1693304636
transform 1 0 2187 0 1 1913
box -876 -128 876 128
use nmos_3p3_AJEA3B  nmos_3p3_AJEA3B_2
timestamp 1693304636
transform 1 0 -1342 0 1 2287
box -876 -128 876 128
use nmos_3p3_AJEA3B  nmos_3p3_AJEA3B_3
timestamp 1693304636
transform 1 0 -1342 0 1 1913
box -876 -128 876 128
use nmos_3p3_AJEA3B  nmos_3p3_AJEA3B_4
timestamp 1693304636
transform 1 0 426 0 1 2287
box -876 -128 876 128
use nmos_3p3_AJEA3B  nmos_3p3_AJEA3B_5
timestamp 1693304636
transform 1 0 426 0 1 1913
box -876 -128 876 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_0
timestamp 1692803904
transform 1 0 382 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_1
timestamp 1692803904
transform 1 0 178 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_2
timestamp 1692803904
transform 1 0 382 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_3
timestamp 1692803904
transform 1 0 178 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_4
timestamp 1692803904
transform 1 0 1046 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_5
timestamp 1692803904
transform 1 0 -154 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_6
timestamp 1692803904
transform 1 0 714 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_7
timestamp 1692803904
transform 1 0 -154 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_8
timestamp 1692803904
transform 1 0 714 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_9
timestamp 1692803904
transform 1 0 1046 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_10
timestamp 1692803904
transform 1 0 1250 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_11
timestamp 1692803904
transform 1 0 1250 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_12
timestamp 1692803904
transform 1 0 2194 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_13
timestamp 1692803904
transform 1 0 -486 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_14
timestamp 1692803904
transform 1 0 -486 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_15
timestamp 1692803904
transform 1 0 -690 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_16
timestamp 1692803904
transform 1 0 -690 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_17
timestamp 1692803904
transform 1 0 1990 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_18
timestamp 1692803904
transform 1 0 1786 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_19
timestamp 1692803904
transform 1 0 1582 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_20
timestamp 1692803904
transform 1 0 -1022 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_21
timestamp 1692803904
transform 1 0 -1226 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_22
timestamp 1692803904
transform 1 0 -1430 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_23
timestamp 1692803904
transform 1 0 2526 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_24
timestamp 1692803904
transform 1 0 -1634 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_25
timestamp 1692803904
transform 1 0 -1975 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_26
timestamp 1692803904
transform 1 0 2526 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_27
timestamp 1692803904
transform 1 0 -1634 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_28
timestamp 1692803904
transform 1 0 -1430 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_29
timestamp 1692803904
transform 1 0 -1226 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_30
timestamp 1692803904
transform 1 0 -1022 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_31
timestamp 1692803904
transform 1 0 1582 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_32
timestamp 1692803904
transform 1 0 1786 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_33
timestamp 1692803904
transform 1 0 1990 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_34
timestamp 1692803904
transform 1 0 2194 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_35
timestamp 1692803904
transform 1 0 -1975 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_36
timestamp 1692803904
transform 1 0 2730 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_37
timestamp 1692803904
transform 1 0 2730 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_38
timestamp 1692803904
transform 1 0 -2587 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_39
timestamp 1692803904
transform 1 0 -2587 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_40
timestamp 1692803904
transform 1 0 -2179 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_41
timestamp 1692803904
transform 1 0 -2383 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_42
timestamp 1692803904
transform 1 0 -2179 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_43
timestamp 1692803904
transform 1 0 -2383 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_44
timestamp 1692803904
transform 1 0 3138 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_45
timestamp 1692803904
transform 1 0 2934 0 1 128
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_46
timestamp 1692803904
transform 1 0 3138 0 1 -198
box -162 -128 162 128
use nmos_3p3_MGEA3B  nmos_3p3_MGEA3B_47
timestamp 1692803904
transform 1 0 2934 0 1 -198
box -162 -128 162 128
use pmos_3p3_DVJ9E7  pmos_3p3_DVJ9E7_0
timestamp 1693295468
transform 1 0 364 0 1 950
box -1754 -190 1754 190
use pmos_3p3_KYXSLM  pmos_3p3_KYXSLM_0
timestamp 1693295468
transform 1 0 3024 0 1 950
box -938 -190 938 190
use pmos_3p3_KYXSLM  pmos_3p3_KYXSLM_1
timestamp 1693295468
transform 1 0 -2320 0 1 950
box -938 -190 938 190
<< labels >>
flabel psubdiffcont -2150 2670 -2150 2670 0 FreeSans 320 0 0 0 VSS
port 0 nsew
flabel via1 2790 1920 2790 1920 0 FreeSans 320 0 0 0 SD0_1
port 4 nsew
flabel nsubdiffcont -1330 1240 -1330 1240 0 FreeSans 320 0 0 0 VDD
port 5 nsew
flabel polycontact -1160 1090 -1160 1090 0 FreeSans 320 0 0 0 G1_1
port 6 nsew
flabel polycontact -970 810 -970 810 0 FreeSans 320 0 0 0 G1_2
port 7 nsew
flabel via1 -1710 960 -1710 960 0 FreeSans 320 0 0 0 SD1_1
port 8 nsew
flabel via1 -2080 -30 -2080 -30 0 FreeSans 320 0 0 0 SD2_1
port 9 nsew
flabel polysilicon 70 -50 70 -50 0 FreeSans 320 0 0 0 ITAIL
port 10 nsew
flabel polycontact 380 -50 380 -50 0 FreeSans 320 0 0 0 G2_1
port 11 nsew
flabel metal1 280 160 280 160 0 FreeSans 320 0 0 0 SD2_2
port 12 nsew
flabel metal1 -60 170 -60 170 0 FreeSans 320 0 0 0 OUT_2
port 13 nsew
flabel metal1 70 170 70 170 0 FreeSans 320 0 0 0 OUT_1
port 14 nsew
flabel metal1 -260 -30 -260 -30 0 FreeSans 320 0 0 0 SD2_3
port 15 nsew
flabel via1 -590 -40 -590 -40 0 FreeSans 320 0 0 0 SD2_4
port 16 nsew
flabel metal1 -800 160 -800 160 0 FreeSans 320 0 0 0 OUT_3
port 17 nsew
flabel metal1 -930 -210 -930 -210 0 FreeSans 320 0 0 0 OUT_4
port 18 nsew
flabel via1 -1120 -40 -1120 -40 0 FreeSans 320 0 0 0 SD2_5
port 19 nsew
flabel via1 -190 2280 -190 2280 0 FreeSans 320 0 0 0 SD0_2
port 21 nsew
flabel metal1 3150 2110 3150 2110 0 FreeSans 320 0 0 0 OUT_5
port 22 nsew
flabel polycontact -2060 2470 -2060 2470 0 FreeSans 320 0 0 0 ITAIL_1
port 1 nsew
flabel via1 -2295 3441 -2295 3441 0 FreeSans 320 0 0 0 SD3_1
port 23 nsew
flabel metal1 3756 3277 3756 3277 0 FreeSans 320 0 0 0 OUT_6
port 24 nsew
<< end >>
