magic
tech gf180mcuC
magscale 1 10
timestamp 1693568990
<< nwell >>
rect -282 -530 282 530
<< pmos >>
rect -108 -400 -52 400
rect 52 -400 108 400
<< pdiff >>
rect -196 387 -108 400
rect -196 -387 -183 387
rect -137 -387 -108 387
rect -196 -400 -108 -387
rect -52 387 52 400
rect -52 -387 -23 387
rect 23 -387 52 387
rect -52 -400 52 -387
rect 108 387 196 400
rect 108 -387 137 387
rect 183 -387 196 387
rect 108 -400 196 -387
<< pdiffc >>
rect -183 -387 -137 387
rect -23 -387 23 387
rect 137 -387 183 387
<< polysilicon >>
rect -108 400 -52 444
rect 52 400 108 444
rect -108 -444 -52 -400
rect 52 -444 108 -400
<< metal1 >>
rect -183 387 -137 398
rect -183 -398 -137 -387
rect -23 387 23 398
rect -23 -398 23 -387
rect 137 387 183 398
rect 137 -398 183 -387
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 4 l 0.280 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
