magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -3244 -2180 3244 2180
<< nwell >>
rect -1244 -180 1244 180
<< pmos >>
rect -1070 -50 -970 50
rect -866 -50 -766 50
rect -662 -50 -562 50
rect -458 -50 -358 50
rect -254 -50 -154 50
rect -50 -50 50 50
rect 154 -50 254 50
rect 358 -50 458 50
rect 562 -50 662 50
rect 766 -50 866 50
rect 970 -50 1070 50
<< pdiff >>
rect -1158 23 -1070 50
rect -1158 -23 -1145 23
rect -1099 -23 -1070 23
rect -1158 -50 -1070 -23
rect -970 23 -866 50
rect -970 -23 -941 23
rect -895 -23 -866 23
rect -970 -50 -866 -23
rect -766 23 -662 50
rect -766 -23 -737 23
rect -691 -23 -662 23
rect -766 -50 -662 -23
rect -562 23 -458 50
rect -562 -23 -533 23
rect -487 -23 -458 23
rect -562 -50 -458 -23
rect -358 23 -254 50
rect -358 -23 -329 23
rect -283 -23 -254 23
rect -358 -50 -254 -23
rect -154 23 -50 50
rect -154 -23 -125 23
rect -79 -23 -50 23
rect -154 -50 -50 -23
rect 50 23 154 50
rect 50 -23 79 23
rect 125 -23 154 23
rect 50 -50 154 -23
rect 254 23 358 50
rect 254 -23 283 23
rect 329 -23 358 23
rect 254 -50 358 -23
rect 458 23 562 50
rect 458 -23 487 23
rect 533 -23 562 23
rect 458 -50 562 -23
rect 662 23 766 50
rect 662 -23 691 23
rect 737 -23 766 23
rect 662 -50 766 -23
rect 866 23 970 50
rect 866 -23 895 23
rect 941 -23 970 23
rect 866 -50 970 -23
rect 1070 23 1158 50
rect 1070 -23 1099 23
rect 1145 -23 1158 23
rect 1070 -50 1158 -23
<< pdiffc >>
rect -1145 -23 -1099 23
rect -941 -23 -895 23
rect -737 -23 -691 23
rect -533 -23 -487 23
rect -329 -23 -283 23
rect -125 -23 -79 23
rect 79 -23 125 23
rect 283 -23 329 23
rect 487 -23 533 23
rect 691 -23 737 23
rect 895 -23 941 23
rect 1099 -23 1145 23
<< polysilicon >>
rect -1070 50 -970 94
rect -866 50 -766 94
rect -662 50 -562 94
rect -458 50 -358 94
rect -254 50 -154 94
rect -50 50 50 94
rect 154 50 254 94
rect 358 50 458 94
rect 562 50 662 94
rect 766 50 866 94
rect 970 50 1070 94
rect -1070 -94 -970 -50
rect -866 -94 -766 -50
rect -662 -94 -562 -50
rect -458 -94 -358 -50
rect -254 -94 -154 -50
rect -50 -94 50 -50
rect 154 -94 254 -50
rect 358 -94 458 -50
rect 562 -94 662 -50
rect 766 -94 866 -50
rect 970 -94 1070 -50
<< metal1 >>
rect -1145 23 -1099 48
rect -1145 -48 -1099 -23
rect -941 23 -895 48
rect -941 -48 -895 -23
rect -737 23 -691 48
rect -737 -48 -691 -23
rect -533 23 -487 48
rect -533 -48 -487 -23
rect -329 23 -283 48
rect -329 -48 -283 -23
rect -125 23 -79 48
rect -125 -48 -79 -23
rect 79 23 125 48
rect 79 -48 125 -23
rect 283 23 329 48
rect 283 -48 329 -23
rect 487 23 533 48
rect 487 -48 533 -23
rect 691 23 737 48
rect 691 -48 737 -23
rect 895 23 941 48
rect 895 -48 941 -23
rect 1099 23 1145 48
rect 1099 -48 1145 -23
<< end >>
