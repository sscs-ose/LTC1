magic
tech gf180mcuD
magscale 1 10
timestamp 1713971515
<< checkpaint >>
rect -2155 -7517 35192 7581
<< nwell >>
rect 6246 3962 6974 5113
rect 14428 4186 14814 5113
rect 28910 4324 29071 4351
rect 28910 4244 29236 4324
rect 25194 3999 25577 4053
rect 25196 3473 25577 3999
rect 28910 3296 29071 4244
rect 30855 3296 30999 4351
rect 7592 126 8320 1277
rect 14484 127 14870 1054
rect 20992 127 21302 1225
rect 22371 127 22557 1225
rect 23442 127 23562 1225
rect 29740 151 29921 224
rect 7592 -4482 8325 -3940
rect 7592 -4510 8366 -4482
rect 1020 -5090 1022 -4935
rect 7592 -5090 8325 -4510
rect 14490 -5090 14808 -4163
<< pwell >>
rect 21754 3156 21850 3516
rect 28848 2911 29133 3271
rect 30793 2911 31063 3271
rect 20992 1301 21268 1618
<< psubdiff >>
rect 28832 2846 29127 2864
rect 28832 2800 28940 2846
rect 28986 2800 29127 2846
rect 28832 2783 29127 2800
<< nsubdiff >>
rect 29062 4307 29236 4324
rect 29062 4261 29104 4307
rect 29150 4261 29236 4307
rect 29062 4244 29236 4261
rect 29740 151 29921 224
<< psubdiffcont >>
rect 28940 2800 28986 2846
<< nsubdiffcont >>
rect 29104 4261 29150 4307
<< metal1 >>
rect -16 5504 23455 5565
rect -16 4098 45 5504
rect 6710 5358 22787 5409
rect 917 5251 998 5252
rect 917 5237 6481 5251
rect 917 5185 931 5237
rect 983 5185 6481 5237
rect 917 5172 6481 5185
rect 917 5171 998 5172
rect 6402 4464 6481 5172
rect 6170 4385 6481 4464
rect 917 4212 994 4226
rect 917 4160 931 4212
rect 983 4160 994 4212
rect 6710 4163 6761 5358
rect 14647 5215 14723 5227
rect 14647 5163 14659 5215
rect 14711 5163 14723 5215
rect 14647 5151 14723 5163
rect 19564 5220 19644 5231
rect 22342 5220 22425 5232
rect 19564 5219 22425 5220
rect 19564 5167 19578 5219
rect 19630 5173 22357 5219
rect 19630 5167 19644 5173
rect 22307 5167 22357 5173
rect 22409 5167 22425 5219
rect 19564 5155 19644 5167
rect 22342 5155 22425 5167
rect 22554 5082 22628 5088
rect 22211 5074 22628 5082
rect 22211 5022 22560 5074
rect 22612 5022 22628 5074
rect 22211 5015 22628 5022
rect 22554 5008 22628 5015
rect 14519 4809 14703 4856
rect 22736 4341 22787 5358
rect 22607 4328 22787 4341
rect 22607 4276 22620 4328
rect 22672 4276 22787 4328
rect 22607 4273 22787 4276
rect 22607 4264 22686 4273
rect 23394 4264 23455 5504
rect 23587 5535 25213 5581
rect 23587 4912 23633 5535
rect 23957 5458 24023 5465
rect 23957 5406 23964 5458
rect 24016 5406 24023 5458
rect 24607 5460 24663 5462
rect 24607 5408 24609 5460
rect 24661 5408 24663 5460
rect 24607 5406 24663 5408
rect 23957 5399 24023 5406
rect 23587 4860 23832 4912
rect 24792 4911 25012 4968
rect 23673 4385 23842 4452
rect 24705 4391 24776 4422
rect 24701 4385 24780 4391
rect 23389 4250 23466 4264
rect 13547 4216 13625 4229
rect 13547 4213 13560 4216
rect 13501 4164 13560 4213
rect 13612 4164 13625 4216
rect 917 4146 994 4160
rect 6703 4001 6761 4163
rect 13547 4152 13625 4164
rect 15580 4215 15651 4227
rect 15580 4163 15592 4215
rect 15644 4163 15651 4215
rect 23389 4198 23401 4250
rect 23453 4198 23466 4250
rect 23389 4184 23466 4198
rect 15580 4151 15651 4163
rect 22277 4166 22350 4178
rect 22277 4165 22768 4166
rect 22277 4113 22290 4165
rect 22342 4113 22768 4165
rect 22277 4112 22768 4113
rect 22277 4100 22350 4112
rect 863 2949 885 3024
rect 6703 2648 6750 4001
rect 14844 3706 14899 3707
rect 14254 3703 14309 3704
rect 14254 3651 14255 3703
rect 14307 3651 14309 3703
rect 14844 3654 14845 3706
rect 14897 3654 14899 3706
rect 22244 3088 22311 3100
rect 7062 2654 7139 2667
rect 7062 2648 7074 2654
rect 6703 2602 7074 2648
rect 7126 2602 7139 2654
rect 6703 2601 7139 2602
rect 7062 2589 7139 2601
rect 944 2279 1023 2294
rect 944 2227 957 2279
rect 1009 2227 1023 2279
rect 944 2217 1023 2227
rect 7289 2169 7337 3084
rect 22244 3082 22257 3088
rect 13601 3018 13674 3030
rect 13601 2966 13609 3018
rect 13661 2966 13674 3018
rect 13601 2954 13674 2966
rect 15562 3021 15638 3034
rect 15562 2969 15574 3021
rect 15626 2969 15638 3021
rect 15562 2956 15638 2969
rect 19220 2729 19298 2743
rect 19220 2677 19234 2729
rect 19286 2677 19298 2729
rect 19220 2664 19298 2677
rect 19826 2706 19903 2719
rect 19235 2467 19281 2664
rect 19826 2654 19838 2706
rect 19890 2704 19903 2706
rect 21531 2707 21609 2719
rect 21531 2704 21544 2707
rect 19890 2657 21544 2704
rect 19890 2654 19903 2657
rect 19826 2642 19903 2654
rect 21531 2655 21544 2657
rect 21596 2655 21609 2707
rect 21531 2643 21609 2655
rect 19395 2469 19474 2483
rect 19395 2467 19408 2469
rect 19235 2421 19408 2467
rect 19395 2417 19408 2421
rect 19460 2417 19474 2469
rect 19395 2404 19474 2417
rect 13676 2215 13713 2290
rect 15524 2215 15557 2290
rect 8237 2078 8309 2087
rect 9563 2078 9642 2085
rect 8237 2073 9642 2078
rect 8237 2021 8250 2073
rect 8302 2072 9642 2073
rect 8302 2021 9576 2072
rect 8237 2020 9576 2021
rect 9628 2020 9642 2072
rect 8237 2018 9642 2020
rect 8237 2007 8309 2018
rect 9563 2007 9642 2018
rect 21883 1770 21936 1771
rect 21935 1718 21936 1770
rect 21996 1748 22063 3065
rect 22185 3036 22257 3082
rect 22309 3036 22311 3088
rect 22244 3024 22311 3036
rect 22357 3089 22417 4028
rect 22714 3577 22768 4112
rect 23673 4134 23723 4385
rect 24701 4333 24714 4385
rect 24766 4333 24780 4385
rect 24701 4328 24780 4333
rect 24705 4301 24776 4328
rect 24956 4243 25011 4911
rect 25167 4421 25213 5535
rect 25333 5461 25409 5474
rect 25333 5409 25345 5461
rect 25397 5409 25409 5461
rect 25333 5396 25409 5409
rect 25346 4561 25394 5396
rect 25346 4513 27373 4561
rect 25167 4375 26994 4421
rect 24956 4188 25510 4243
rect 23673 4084 25325 4134
rect 23198 3601 23252 3602
rect 23198 3549 23199 3601
rect 23251 3549 23252 3601
rect 23640 3390 23703 3538
rect 25275 3428 25325 4084
rect 23409 3327 23703 3390
rect 22357 3040 22710 3089
rect 22199 2713 22270 2721
rect 22357 2713 22417 3040
rect 22199 2708 22417 2713
rect 22199 2656 22211 2708
rect 22263 2656 22417 2708
rect 22199 2653 22417 2656
rect 22199 2644 22270 2653
rect 22457 2073 22560 2159
rect 21344 1590 21426 1604
rect 165 1589 221 1590
rect 165 1537 167 1589
rect 219 1537 221 1589
rect 21344 1538 21359 1590
rect 21411 1538 21426 1590
rect 21344 1525 21426 1538
rect 21358 1479 21411 1525
rect 21313 1426 21411 1479
rect 7779 1247 7855 1261
rect 21313 1248 21366 1426
rect 22235 1262 22313 1274
rect 7779 1245 7792 1247
rect 7764 1198 7792 1245
rect 7779 1195 7792 1198
rect 7844 1195 7855 1247
rect 22235 1210 22248 1262
rect 22300 1210 22313 1262
rect 22235 1198 22313 1210
rect 7779 1181 7855 1195
rect 940 1081 1011 1096
rect 940 1029 944 1081
rect 996 1029 1011 1081
rect 940 1016 1011 1029
rect 13575 1089 13649 1102
rect 13575 1037 13584 1089
rect 13636 1037 13649 1089
rect 13575 1024 13649 1037
rect 15602 1088 15679 1102
rect 15602 1036 15615 1088
rect 15667 1036 15679 1088
rect 15602 1022 15679 1036
rect 8308 836 8382 854
rect 8302 821 8382 836
rect 8302 769 8314 821
rect 8366 769 8382 821
rect 8302 755 8382 769
rect 8302 754 8379 755
rect 8037 633 8117 646
rect 8037 581 8051 633
rect 8103 581 8117 633
rect 8037 568 8117 581
rect 594 162 598 214
rect 650 162 654 214
rect 0 -1201 47 74
rect 6694 13 6775 19
rect 8053 13 8101 568
rect 20845 478 20924 860
rect 21206 717 21262 794
rect 20845 399 21141 478
rect 6694 6 8101 13
rect 6694 -46 6708 6
rect 6760 -35 8101 6
rect 6760 -46 6775 -35
rect 6694 -59 6775 -46
rect 597 -135 654 -132
rect 597 -187 599 -135
rect 651 -187 654 -135
rect 597 -189 654 -187
rect 6192 -752 6260 -751
rect 6170 -765 6263 -752
rect 6170 -817 6201 -765
rect 6253 -817 6263 -765
rect 6170 -831 6263 -817
rect 943 -1022 1026 -1014
rect 943 -1074 958 -1022
rect 1010 -1074 1026 -1022
rect 943 -1088 1026 -1074
rect 6712 -1221 6760 -59
rect 9749 -183 9834 233
rect 21062 102 21141 399
rect 22233 213 22287 214
rect 19011 90 21141 102
rect 19001 82 21141 90
rect 19001 30 19014 82
rect 19066 30 21141 82
rect 19001 23 21141 30
rect 19001 16 19078 23
rect 21768 -172 21850 199
rect 22233 161 22234 213
rect 22286 161 22287 213
rect 13551 -1003 13627 -988
rect 13551 -1055 13562 -1003
rect 13614 -1055 13627 -1003
rect 13551 -1069 13627 -1055
rect 15597 -996 15677 -984
rect 15597 -1048 15611 -996
rect 15663 -1048 15677 -996
rect 15597 -1060 15677 -1048
rect 22457 -1154 22503 2073
rect 23409 1819 23472 3327
rect 25455 2715 25510 4188
rect 25563 3464 25609 4375
rect 26148 3516 26649 3559
rect 26148 3511 26437 3516
rect 26425 3464 26437 3511
rect 26489 3511 26649 3516
rect 26489 3464 26503 3511
rect 25563 3418 25906 3464
rect 26425 3451 26503 3464
rect 26559 2967 26623 2973
rect 26559 2915 26565 2967
rect 26617 2915 26623 2967
rect 26559 2909 26623 2915
rect 26588 2728 26672 2735
rect 26546 2719 26672 2728
rect 26546 2715 26604 2719
rect 25455 2667 26604 2715
rect 26656 2667 26672 2719
rect 26948 2720 26994 4375
rect 27325 4279 27373 4513
rect 28817 4307 29236 4324
rect 28817 4261 29104 4307
rect 29150 4261 29236 4307
rect 28817 4248 29236 4261
rect 30753 4248 31108 4324
rect 28826 4244 29236 4248
rect 28889 3788 28968 3801
rect 28889 3736 28902 3788
rect 28954 3736 28968 3788
rect 30857 3786 30933 3798
rect 28889 3724 28968 3736
rect 29042 3737 29157 3784
rect 30857 3775 30869 3786
rect 29042 3583 29089 3737
rect 30852 3734 30869 3775
rect 30921 3734 30933 3786
rect 30852 3729 30933 3734
rect 30990 3737 31085 3784
rect 29011 3569 29089 3583
rect 30990 3721 31084 3737
rect 32780 3729 32928 3775
rect 30990 3582 31037 3721
rect 29011 3517 29024 3569
rect 29076 3517 29089 3569
rect 29011 3510 29089 3517
rect 30892 3569 31037 3582
rect 30892 3517 30906 3569
rect 30958 3517 31037 3569
rect 30892 3510 31037 3517
rect 29011 3504 29084 3510
rect 32878 3036 32928 3729
rect 32878 2986 33192 3036
rect 27328 2846 27381 2847
rect 27380 2794 27381 2846
rect 27328 2793 27381 2794
rect 28832 2846 29234 2864
rect 28832 2800 28940 2846
rect 28986 2800 29234 2846
rect 28832 2783 29234 2800
rect 30775 2783 31086 2864
rect 26948 2674 33051 2720
rect 25455 2660 26672 2667
rect 26546 2659 26672 2660
rect 26588 2652 26672 2659
rect 23560 2168 23672 2269
rect 23579 1906 23626 2168
rect 23744 2038 23803 2039
rect 23744 1986 23747 2038
rect 23799 1986 23803 2038
rect 23744 1985 23803 1986
rect 23579 1859 24815 1906
rect 23746 1779 23805 1780
rect 23746 1727 23749 1779
rect 23801 1727 23805 1779
rect 23746 1726 23805 1727
rect 23615 1301 23786 1318
rect 23615 1249 23703 1301
rect 23755 1249 23786 1301
rect 24768 1259 24815 1859
rect 25106 1690 25152 2029
rect 33005 1956 33051 2674
rect 25467 1692 25547 1705
rect 25467 1690 25481 1692
rect 25106 1644 25481 1690
rect 25467 1640 25481 1644
rect 25533 1640 25547 1692
rect 25467 1628 25547 1640
rect 25484 1418 25530 1628
rect 27610 1535 27687 1548
rect 27610 1483 27622 1535
rect 27674 1483 27687 1535
rect 27610 1470 27687 1483
rect 25484 1372 25757 1418
rect 23615 1234 23786 1249
rect 24576 1212 24815 1259
rect 23420 729 23502 781
rect 22750 215 22804 216
rect 22750 163 22751 215
rect 22803 163 22804 215
rect 23420 106 23473 729
rect 24474 214 24553 224
rect 24474 162 24490 214
rect 24542 213 24553 214
rect 24542 162 26818 213
rect 24474 157 26818 162
rect 24474 153 24553 157
rect 22636 51 23473 106
rect 22434 -1169 22519 -1154
rect 22434 -1221 22451 -1169
rect 22503 -1221 22519 -1169
rect 22434 -1235 22519 -1221
rect 173 -1491 243 -1478
rect 173 -1543 177 -1491
rect 229 -1543 243 -1491
rect 22636 -1507 22691 51
rect 28450 4 28527 15
rect 22871 1 28527 4
rect 22871 -51 28459 1
rect 28511 -51 28527 1
rect 22871 -55 28527 -51
rect 22871 -765 22930 -55
rect 28450 -65 28527 -55
rect 28992 -187 29040 215
rect 29740 151 29921 224
rect 33142 47 33192 2986
rect 29586 -3 33192 47
rect 22871 -824 23237 -765
rect 28410 -1010 28493 -996
rect 28410 -1062 28425 -1010
rect 28477 -1062 28493 -1010
rect 28410 -1078 28493 -1062
rect 173 -1547 243 -1543
rect 14320 -1516 14377 -1514
rect 14320 -1568 14322 -1516
rect 14374 -1568 14377 -1516
rect 14862 -1515 14919 -1513
rect 14862 -1567 14864 -1515
rect 14916 -1567 14919 -1515
rect 14862 -1568 14919 -1567
rect 22271 -1562 22691 -1507
rect 14320 -1569 14377 -1568
rect 13683 -2087 13761 -2073
rect 13683 -2139 13695 -2087
rect 13747 -2139 13761 -2087
rect 867 -2267 884 -2192
rect 966 -2937 1047 -2923
rect 966 -2989 980 -2937
rect 1032 -2989 1047 -2937
rect 966 -2998 1047 -2989
rect 7119 -3053 7187 -2144
rect 13683 -2151 13761 -2139
rect 13695 -2197 13745 -2151
rect 13543 -2247 13745 -2197
rect 15586 -2188 15668 -2176
rect 15586 -2240 15600 -2188
rect 15652 -2198 15668 -2188
rect 15652 -2240 15789 -2198
rect 15586 -2244 15789 -2240
rect 15586 -2252 15668 -2244
rect 19136 -2487 19214 -2474
rect 10405 -2503 10483 -2490
rect 10405 -2555 10418 -2503
rect 10470 -2555 10483 -2503
rect 19136 -2539 19149 -2487
rect 19201 -2539 19214 -2487
rect 19136 -2552 19214 -2539
rect 10405 -2567 10483 -2555
rect 8224 -3151 8300 -3137
rect 8224 -3203 8236 -3151
rect 8288 -3154 8300 -3151
rect 10421 -3154 10468 -2567
rect 13686 -3002 13705 -2927
rect 15521 -3002 15552 -2927
rect 8288 -3201 10468 -3154
rect 19150 -3183 19201 -2552
rect 22271 -2721 22326 -1562
rect 22508 -1868 22594 -1854
rect 22508 -1920 22525 -1868
rect 22577 -1920 22594 -1868
rect 22508 -1934 22594 -1920
rect 21346 -2776 22326 -2721
rect 20887 -3171 20963 -3158
rect 20887 -3183 20899 -3171
rect 8288 -3203 8300 -3201
rect 8224 -3216 8300 -3203
rect 19150 -3223 20899 -3183
rect 20951 -3223 20963 -3171
rect 19150 -3234 20963 -3223
rect 20887 -3236 20963 -3234
rect 20930 -3368 20931 -3316
rect 20983 -3368 20984 -3316
rect 7781 -3965 7860 -3952
rect 7781 -4017 7793 -3965
rect 7845 -4017 7860 -3965
rect 7781 -4018 7860 -4017
rect 7781 -4024 7854 -4018
rect 959 -4142 1030 -4129
rect 959 -4194 966 -4142
rect 1018 -4194 1030 -4142
rect 959 -4206 1030 -4194
rect 7799 -5117 7854 -4024
rect 14519 -4026 14703 -3980
rect 13580 -4121 13649 -4103
rect 13580 -4173 13591 -4121
rect 13643 -4173 13649 -4121
rect 15592 -4132 15664 -4117
rect 13580 -4190 13649 -4173
rect 14490 -4155 14577 -4140
rect 14490 -4207 14507 -4155
rect 14559 -4207 14577 -4155
rect 15592 -4184 15606 -4132
rect 15658 -4184 15664 -4132
rect 15592 -4198 15664 -4184
rect 14490 -4222 14577 -4207
rect 8300 -4363 8373 -4362
rect 8300 -4377 8378 -4363
rect 8300 -4429 8312 -4377
rect 8364 -4429 8378 -4377
rect 8300 -4442 8378 -4429
rect 20837 -4377 20906 -4361
rect 20837 -4429 20844 -4377
rect 20896 -4429 20906 -4377
rect 21346 -4380 21401 -2776
rect 22526 -2881 22578 -1934
rect 23007 -2123 23093 -2109
rect 23007 -2175 23024 -2123
rect 23076 -2125 23093 -2123
rect 23076 -2171 24929 -2125
rect 23076 -2175 23093 -2171
rect 23007 -2189 23093 -2175
rect 24883 -2659 24929 -2171
rect 28519 -2267 28548 -2192
rect 24872 -2672 24951 -2659
rect 24872 -2724 24885 -2672
rect 24937 -2724 24951 -2672
rect 24872 -2737 24951 -2724
rect 8300 -4444 8373 -4442
rect 20837 -4447 20906 -4429
rect 21267 -4435 21401 -4380
rect 21605 -2933 22578 -2881
rect 15633 -5064 15762 -4987
rect 21267 -5117 21322 -4435
rect 7799 -5172 21324 -5117
rect 961 -5266 1037 -5262
rect 961 -5274 14319 -5266
rect 961 -5326 973 -5274
rect 1025 -5318 14319 -5274
rect 1025 -5326 1037 -5318
rect 961 -5338 1037 -5326
rect 14267 -5465 14319 -5318
rect 14544 -5301 14621 -5287
rect 14544 -5353 14556 -5301
rect 14608 -5303 14621 -5301
rect 21357 -5302 21434 -5289
rect 21357 -5303 21369 -5302
rect 14608 -5353 21369 -5303
rect 14544 -5367 14621 -5353
rect 21357 -5354 21369 -5353
rect 21421 -5354 21434 -5302
rect 21357 -5366 21434 -5354
rect 21605 -5465 21657 -2933
rect 28409 -2944 28484 -2929
rect 28409 -2996 28417 -2944
rect 28469 -2996 28484 -2944
rect 28409 -3009 28484 -2996
rect 21902 -3065 21903 -3013
rect 21955 -3065 21956 -3013
rect 29586 -3550 29636 -3
rect 29367 -3600 29636 -3550
rect 28407 -4138 28483 -4124
rect 28407 -4190 28419 -4138
rect 28471 -4190 28483 -4138
rect 28407 -4203 28483 -4190
rect 21761 -5301 21837 -5289
rect 21761 -5353 21773 -5301
rect 21825 -5303 21837 -5301
rect 29586 -5303 29636 -3600
rect 21825 -5353 29636 -5303
rect 21761 -5365 21837 -5353
rect 14267 -5517 21657 -5465
<< via1 >>
rect 931 5185 983 5237
rect 931 4160 983 4212
rect 14659 5163 14711 5215
rect 19578 5167 19630 5219
rect 22357 5167 22409 5219
rect 22560 5022 22612 5074
rect 22620 4276 22672 4328
rect 23964 5406 24016 5458
rect 24609 5408 24661 5460
rect 13560 4164 13612 4216
rect 15592 4163 15644 4215
rect 23401 4198 23453 4250
rect 22290 4113 22342 4165
rect 14255 3651 14307 3703
rect 14845 3654 14897 3706
rect 7074 2602 7126 2654
rect 957 2227 1009 2279
rect 13609 2966 13661 3018
rect 15574 2969 15626 3021
rect 19234 2677 19286 2729
rect 19838 2654 19890 2706
rect 21544 2655 21596 2707
rect 19408 2417 19460 2469
rect 8250 2021 8302 2073
rect 9576 2020 9628 2072
rect 21883 1718 21935 1770
rect 22257 3036 22309 3088
rect 24714 4333 24766 4385
rect 25345 5409 25397 5461
rect 24942 3956 24994 4008
rect 23199 3549 23251 3601
rect 22211 2656 22263 2708
rect 167 1537 219 1589
rect 21359 1538 21411 1590
rect 7792 1195 7844 1247
rect 22248 1210 22300 1262
rect 944 1029 996 1081
rect 13584 1037 13636 1089
rect 15615 1036 15667 1088
rect 8314 769 8366 821
rect 8051 581 8103 633
rect 598 162 650 214
rect 6708 -46 6760 6
rect 599 -187 651 -135
rect 6201 -817 6253 -765
rect 958 -1074 1010 -1022
rect 19014 30 19066 82
rect 22234 161 22286 213
rect 13562 -1055 13614 -1003
rect 15611 -1048 15663 -996
rect 25760 3946 25812 3998
rect 26437 3464 26489 3516
rect 26565 2915 26617 2967
rect 26604 2667 26656 2719
rect 28902 3736 28954 3788
rect 30869 3734 30921 3786
rect 29024 3517 29076 3569
rect 30906 3517 30958 3569
rect 27328 2794 27380 2846
rect 23747 1986 23799 2038
rect 23749 1727 23801 1779
rect 23703 1249 23755 1301
rect 25481 1640 25533 1692
rect 27622 1483 27674 1535
rect 22751 163 22803 215
rect 24490 162 24542 214
rect 22451 -1221 22503 -1169
rect 177 -1543 229 -1491
rect 28459 -51 28511 1
rect 28425 -1062 28477 -1010
rect 14322 -1568 14374 -1516
rect 14864 -1567 14916 -1515
rect 13695 -2139 13747 -2087
rect 980 -2989 1032 -2937
rect 15600 -2240 15652 -2188
rect 10418 -2555 10470 -2503
rect 19149 -2539 19201 -2487
rect 8236 -3203 8288 -3151
rect 22525 -1920 22577 -1868
rect 20899 -3223 20951 -3171
rect 20931 -3368 20983 -3316
rect 7793 -4017 7845 -3965
rect 966 -4194 1018 -4142
rect 13591 -4173 13643 -4121
rect 14507 -4207 14559 -4155
rect 15606 -4184 15658 -4132
rect 8312 -4429 8364 -4377
rect 20844 -4429 20896 -4377
rect 23024 -2175 23076 -2123
rect 24885 -2724 24937 -2672
rect 973 -5326 1025 -5274
rect 14556 -5353 14608 -5301
rect 21369 -5354 21421 -5302
rect 28417 -2996 28469 -2944
rect 21903 -3065 21955 -3013
rect 28419 -4190 28471 -4138
rect 21773 -5353 21825 -5301
<< metal2 >>
rect 6467 5463 22089 5523
rect 23950 5466 24029 5469
rect 24594 5466 24676 5469
rect 25333 5466 25409 5474
rect 917 5237 998 5252
rect 917 5185 931 5237
rect 983 5185 998 5237
rect 917 5171 998 5185
rect 926 4226 988 5171
rect 917 4212 994 4226
rect 917 4160 931 4212
rect 983 4160 994 4212
rect 917 4146 994 4160
rect 944 2283 1023 2294
rect 944 2227 956 2283
rect 1012 2227 1023 2283
rect 944 2217 1023 2227
rect 6467 2120 6527 5463
rect 6849 5296 21170 5357
rect 6849 2515 6910 5296
rect 14647 5224 14723 5227
rect 14647 5215 18329 5224
rect 19564 5223 19644 5231
rect 14647 5163 14659 5215
rect 14711 5165 18329 5215
rect 14711 5163 14723 5165
rect 14647 5151 14723 5163
rect 18270 4698 18329 5165
rect 18687 5219 19644 5223
rect 18687 5167 19578 5219
rect 19630 5167 19644 5219
rect 18687 5164 19644 5167
rect 18687 4698 18746 5164
rect 19564 5155 19644 5164
rect 18270 4639 18746 4698
rect 13547 4218 13625 4229
rect 13547 4162 13558 4218
rect 13614 4162 13625 4218
rect 15580 4215 15651 4227
rect 13547 4152 13625 4162
rect 15573 4163 15592 4215
rect 15644 4163 15651 4215
rect 15573 4151 15651 4163
rect 14242 3709 14321 3716
rect 14840 3709 14911 3718
rect 14242 3706 14911 3709
rect 14242 3703 14845 3706
rect 14242 3651 14255 3703
rect 14307 3654 14845 3703
rect 14897 3654 14911 3706
rect 14307 3653 14911 3654
rect 14307 3651 14321 3653
rect 14242 3639 14321 3651
rect 14840 3639 14911 3653
rect 15573 3034 15629 4151
rect 13585 3020 13674 3030
rect 15562 3021 15638 3034
rect 15562 3020 15574 3021
rect 13559 3019 15574 3020
rect 13559 2964 13596 3019
rect 13652 3018 15574 3019
rect 13661 2969 15574 3018
rect 15626 2969 15638 3021
rect 13661 2966 15638 2969
rect 13585 2963 13596 2964
rect 13652 2964 15638 2966
rect 13652 2963 13674 2964
rect 13585 2954 13674 2963
rect 15562 2956 15638 2964
rect 13585 2953 13664 2954
rect 16726 2777 16801 2787
rect 13776 2725 13852 2735
rect 13776 2669 13786 2725
rect 13842 2721 13852 2725
rect 19220 2729 19298 2743
rect 19220 2721 19234 2729
rect 13842 2677 19234 2721
rect 19286 2677 19298 2729
rect 13842 2669 19298 2677
rect 7062 2663 7139 2667
rect 13776 2665 19298 2669
rect 7062 2654 8300 2663
rect 13776 2659 13852 2665
rect 19220 2664 19298 2665
rect 19826 2706 19903 2719
rect 7062 2602 7074 2654
rect 7126 2602 8300 2654
rect 19826 2654 19838 2706
rect 19890 2654 19903 2706
rect 19826 2642 19903 2654
rect 7062 2594 8300 2602
rect 7062 2589 7139 2594
rect 6849 2454 7851 2515
rect 6467 2060 7391 2120
rect 153 1592 233 1602
rect -1 1589 233 1592
rect -1 1537 167 1589
rect 219 1537 233 1589
rect -1 1536 233 1537
rect -1 -1487 55 1536
rect 153 1525 233 1536
rect 917 1085 1011 1096
rect 917 1029 944 1085
rect 1000 1029 1011 1085
rect 917 1015 1011 1029
rect 7331 636 7391 2060
rect 7790 1261 7851 2454
rect 8231 2087 8300 2594
rect 19395 2472 19474 2483
rect 19833 2472 19891 2642
rect 19395 2469 19891 2472
rect 19395 2417 19408 2469
rect 19460 2417 19891 2469
rect 19395 2414 19891 2417
rect 19395 2404 19474 2414
rect 8231 2073 8309 2087
rect 8231 2047 8250 2073
rect 8237 2021 8250 2047
rect 8302 2021 8309 2073
rect 8237 2007 8309 2021
rect 9563 2077 9642 2085
rect 9563 2072 10928 2077
rect 9563 2020 9576 2072
rect 9628 2020 10928 2072
rect 9563 2014 10928 2020
rect 9563 2007 9642 2014
rect 7779 1247 7855 1261
rect 7779 1195 7792 1247
rect 7844 1195 7855 1247
rect 7779 1181 7855 1195
rect 10865 1122 10928 2014
rect 12717 1655 14723 1718
rect 12717 1122 12780 1655
rect 10865 1059 12780 1122
rect 13572 1089 13653 1115
rect 13572 1037 13584 1089
rect 13636 1037 13653 1089
rect 13572 1027 13653 1037
rect 13575 1024 13653 1027
rect 8302 821 8379 836
rect 8302 769 8314 821
rect 8366 769 8379 821
rect 8302 754 8379 769
rect 8037 637 8117 646
rect 7989 636 8117 637
rect 7331 633 8117 636
rect 7331 581 8051 633
rect 8103 581 8117 633
rect 7331 576 8117 581
rect 8037 568 8117 576
rect 582 214 667 226
rect 582 162 598 214
rect 650 162 667 214
rect 582 155 667 162
rect 594 -125 654 155
rect 8311 89 8369 754
rect 10124 132 11292 190
rect 10124 89 10182 132
rect 905 -29 3543 44
rect 8311 31 10182 89
rect 11234 69 11292 132
rect 13595 69 13653 1024
rect 6694 8 6775 19
rect 11234 11 13653 69
rect 585 -135 666 -125
rect 585 -187 599 -135
rect 651 -187 666 -135
rect 585 -194 666 -187
rect 913 -985 986 -29
rect 3470 -160 3543 -29
rect 4120 -75 6318 -2
rect 6694 -48 6706 8
rect 6762 -48 6775 8
rect 6694 -59 6775 -48
rect 14660 -54 14723 1655
rect 15602 1088 15679 1102
rect 15602 1036 15615 1088
rect 15667 1036 15679 1088
rect 15602 1022 15679 1036
rect 15609 23 15668 1022
rect 21109 795 21170 5296
rect 22029 2903 22089 5463
rect 23658 5458 24048 5466
rect 23658 5406 23964 5458
rect 24016 5406 24048 5458
rect 23658 5400 24048 5406
rect 24594 5461 25409 5466
rect 24594 5460 25345 5461
rect 24594 5408 24609 5460
rect 24661 5409 25345 5460
rect 25397 5409 25409 5461
rect 24661 5408 25409 5409
rect 24594 5401 25409 5408
rect 24594 5400 24676 5401
rect 22342 5219 22425 5232
rect 22342 5167 22357 5219
rect 22409 5167 22425 5219
rect 22342 5155 22425 5167
rect 22349 4535 22419 5155
rect 22554 5080 22628 5088
rect 23658 5080 23724 5400
rect 23945 5387 24048 5400
rect 25333 5396 25409 5401
rect 22554 5074 23724 5080
rect 22554 5022 22560 5074
rect 22612 5022 23724 5074
rect 22554 5014 23724 5022
rect 22554 5008 22628 5014
rect 22342 4465 30929 4535
rect 24701 4386 24780 4391
rect 23195 4385 24780 4386
rect 22607 4328 22686 4341
rect 22607 4276 22620 4328
rect 22672 4276 22686 4328
rect 22607 4264 22686 4276
rect 23195 4333 24714 4385
rect 24766 4333 24780 4385
rect 23195 4328 24780 4333
rect 23195 4327 24747 4328
rect 22617 4220 22677 4264
rect 22277 4166 22350 4178
rect 22267 4165 22350 4166
rect 22267 4113 22290 4165
rect 22342 4113 22350 4165
rect 22267 4100 22350 4113
rect 22267 3100 22334 4100
rect 22621 3837 22677 4220
rect 22244 3088 22334 3100
rect 22244 3036 22257 3088
rect 22309 3036 22334 3088
rect 22244 3024 22334 3036
rect 22403 3781 22677 3837
rect 21355 2843 22089 2903
rect 21355 1604 21415 2843
rect 21531 2711 21609 2719
rect 22199 2711 22270 2721
rect 21531 2708 22270 2711
rect 21531 2707 22211 2708
rect 21531 2655 21544 2707
rect 21596 2656 22211 2707
rect 22263 2656 22270 2708
rect 21596 2655 22270 2656
rect 21531 2653 22270 2655
rect 21531 2643 21609 2653
rect 22199 2644 22270 2653
rect 22403 2623 22459 3781
rect 23195 3601 23254 4327
rect 23389 4258 23466 4264
rect 23389 4250 28962 4258
rect 23389 4198 23401 4250
rect 23453 4198 28962 4250
rect 23389 4190 28962 4198
rect 23389 4184 23466 4190
rect 24930 4009 25006 4020
rect 25748 4009 25824 4010
rect 24930 4008 25824 4009
rect 24930 3956 24942 4008
rect 24994 3998 25824 4008
rect 24994 3956 25760 3998
rect 24930 3951 25760 3956
rect 24930 3944 25006 3951
rect 23195 3599 23199 3601
rect 23186 3549 23199 3599
rect 23251 3599 23254 3601
rect 23251 3549 23264 3599
rect 23186 3537 23264 3549
rect 23506 3011 24200 3069
rect 22403 2567 22609 2623
rect 23506 2376 23564 3011
rect 22243 2318 23564 2376
rect 21874 1770 21945 1784
rect 21874 1718 21883 1770
rect 21935 1718 21945 1770
rect 21874 1707 21945 1718
rect 21344 1590 21426 1604
rect 21344 1538 21359 1590
rect 21411 1538 21426 1590
rect 21344 1525 21426 1538
rect 21877 1120 21940 1707
rect 22243 1320 22301 2318
rect 23732 2038 23815 2051
rect 23732 1986 23747 2038
rect 23799 1986 23815 2038
rect 23732 1984 23815 1986
rect 23735 1983 23809 1984
rect 23743 1790 23806 1983
rect 23735 1779 23817 1790
rect 23735 1727 23749 1779
rect 23801 1727 23817 1779
rect 23735 1714 23817 1727
rect 23743 1627 23806 1714
rect 22455 1564 23806 1627
rect 22243 1274 22304 1320
rect 22235 1262 22313 1274
rect 22235 1210 22248 1262
rect 22300 1210 22313 1262
rect 22235 1198 22313 1210
rect 22455 1120 22518 1564
rect 23615 1312 23786 1318
rect 21877 1057 22518 1120
rect 23407 1301 23786 1312
rect 23407 1250 23703 1301
rect 21109 717 21313 795
rect 22741 222 22819 227
rect 22222 215 22819 222
rect 22222 213 22751 215
rect 18222 137 18848 196
rect 22222 161 22234 213
rect 22286 163 22751 213
rect 22803 163 22819 215
rect 22286 161 22819 163
rect 22222 155 22819 161
rect 22222 153 22815 155
rect 22222 150 22300 153
rect 18222 23 18281 137
rect 18789 83 18848 137
rect 19001 83 19082 98
rect 18789 82 19082 83
rect 18789 30 19014 82
rect 19066 30 19082 82
rect 18789 24 19082 30
rect 15609 -36 18281 23
rect 19001 16 19082 24
rect 23407 9 23469 1250
rect 23615 1249 23703 1250
rect 23755 1249 23786 1301
rect 23615 1234 23786 1249
rect 25321 224 25379 3951
rect 25748 3946 25760 3951
rect 25812 3946 25824 3998
rect 25748 3934 25824 3946
rect 28894 3801 28962 4190
rect 26431 3730 27811 3799
rect 26431 3578 26500 3730
rect 27742 3579 27811 3730
rect 28889 3788 28968 3801
rect 30859 3798 30929 4465
rect 28889 3736 28902 3788
rect 28954 3736 28968 3788
rect 28889 3724 28968 3736
rect 30857 3786 30933 3798
rect 30857 3734 30869 3786
rect 30921 3734 30933 3786
rect 30857 3729 30933 3734
rect 29011 3579 29089 3583
rect 30892 3579 30972 3582
rect 26425 3516 26503 3578
rect 26425 3464 26437 3516
rect 26489 3464 26503 3516
rect 27742 3569 30972 3579
rect 27742 3517 29024 3569
rect 29076 3517 30906 3569
rect 30958 3517 30972 3569
rect 27742 3510 30972 3517
rect 29011 3504 29089 3510
rect 26425 3451 26503 3464
rect 25475 2967 26778 2985
rect 25475 2921 26565 2967
rect 25475 1705 25539 2921
rect 26547 2915 26565 2921
rect 26617 2921 26778 2967
rect 26617 2915 26635 2921
rect 26547 2897 26635 2915
rect 26714 2851 26778 2921
rect 27316 2851 27393 2859
rect 26714 2846 27393 2851
rect 26714 2794 27328 2846
rect 27380 2794 27393 2846
rect 26714 2787 27393 2794
rect 27316 2780 27393 2787
rect 26588 2719 26672 2735
rect 26588 2667 26604 2719
rect 26656 2667 26672 2719
rect 26588 2652 26672 2667
rect 25467 1692 25547 1705
rect 25467 1640 25481 1692
rect 25533 1640 25547 1692
rect 25467 1628 25547 1640
rect 26601 1541 26660 2652
rect 29789 2156 29846 2157
rect 29845 2100 29846 2156
rect 27610 1541 27687 1548
rect 26601 1535 27687 1541
rect 26601 1483 27622 1535
rect 27674 1483 27687 1535
rect 26601 1482 27687 1483
rect 27563 1478 27687 1482
rect 27610 1470 27687 1478
rect 24474 214 25379 224
rect 24474 162 24490 214
rect 24542 166 25379 214
rect 24542 162 24557 166
rect 24474 153 24557 162
rect 15258 -54 15321 -48
rect 4120 -160 4193 -75
rect 3470 -233 4193 -160
rect 6245 -546 6318 -75
rect 14660 -117 15321 -54
rect 15258 -174 15321 -117
rect 22956 -53 23469 9
rect 28450 1 28527 15
rect 28450 -51 28459 1
rect 28511 -51 28527 1
rect 15258 -237 15669 -174
rect 6190 -619 6318 -546
rect 6190 -765 6263 -619
rect 6190 -817 6201 -765
rect 6253 -817 6263 -765
rect 6190 -830 6263 -817
rect 15606 -984 15669 -237
rect 913 -1022 1023 -985
rect 913 -1072 958 -1022
rect 943 -1074 958 -1072
rect 1010 -1074 1023 -1022
rect 13551 -1003 13627 -988
rect 13551 -1055 13562 -1003
rect 13614 -1055 13627 -1003
rect 13551 -1069 13627 -1055
rect 15597 -996 15677 -984
rect 15597 -1048 15611 -996
rect 15663 -1048 15677 -996
rect 15597 -1060 15677 -1048
rect 943 -1088 1023 -1074
rect 173 -1487 243 -1478
rect -1 -1491 245 -1487
rect -1 -1543 177 -1491
rect 229 -1543 245 -1491
rect 164 -1556 245 -1543
rect 10405 -2503 10483 -2498
rect 10405 -2555 10418 -2503
rect 10470 -2505 10483 -2503
rect 13567 -2505 13623 -1069
rect 22434 -1169 22519 -1154
rect 22434 -1221 22451 -1169
rect 22503 -1221 22519 -1169
rect 22434 -1235 22519 -1221
rect 14308 -1513 14389 -1502
rect 14850 -1513 14931 -1501
rect 14308 -1515 14931 -1513
rect 14308 -1516 14864 -1515
rect 14308 -1568 14322 -1516
rect 14374 -1567 14864 -1516
rect 14916 -1567 14931 -1515
rect 22445 -1516 22501 -1235
rect 14374 -1568 14931 -1567
rect 14308 -1570 14931 -1568
rect 14308 -1581 14389 -1570
rect 14850 -1580 14931 -1570
rect 22306 -1572 22501 -1516
rect 13683 -2078 13761 -2073
rect 15381 -2078 15444 -2077
rect 13683 -2084 15647 -2078
rect 13683 -2140 13694 -2084
rect 13750 -2140 15647 -2084
rect 13683 -2141 15647 -2140
rect 13683 -2151 13761 -2141
rect 10470 -2555 13623 -2505
rect 15381 -2496 15444 -2141
rect 15584 -2176 15647 -2141
rect 22306 -2121 22362 -1572
rect 22508 -1868 22594 -1854
rect 22956 -1868 23018 -53
rect 28450 -65 28527 -51
rect 28457 -111 28525 -65
rect 28467 -994 28525 -111
rect 28410 -1004 28525 -994
rect 28388 -1010 28525 -1004
rect 28388 -1062 28425 -1010
rect 28477 -1062 28525 -1010
rect 28410 -1078 28493 -1062
rect 22508 -1920 22525 -1868
rect 22577 -1920 23018 -1868
rect 22508 -1930 23018 -1920
rect 22508 -1934 22594 -1930
rect 23007 -2121 23093 -2109
rect 22306 -2123 23093 -2121
rect 22306 -2175 23024 -2123
rect 23076 -2175 23093 -2123
rect 15584 -2182 15668 -2176
rect 22306 -2177 23093 -2175
rect 15584 -2188 15706 -2182
rect 15584 -2240 15600 -2188
rect 15652 -2240 15706 -2188
rect 23007 -2189 23093 -2177
rect 15584 -2245 15706 -2240
rect 15586 -2252 15668 -2245
rect 19136 -2487 19214 -2474
rect 19136 -2496 19149 -2487
rect 15381 -2539 19149 -2496
rect 19201 -2539 19214 -2487
rect 15381 -2552 19214 -2539
rect 10405 -2561 13623 -2555
rect 24872 -2672 24951 -2659
rect 24872 -2724 24885 -2672
rect 24937 -2724 24951 -2672
rect 24872 -2737 24951 -2724
rect 966 -2935 1047 -2923
rect 966 -2991 978 -2935
rect 1034 -2991 1047 -2935
rect 966 -2998 1047 -2991
rect 21890 -3011 21968 -3001
rect 21706 -3013 21968 -3011
rect 21706 -3065 21903 -3013
rect 21955 -3065 21968 -3013
rect 21706 -3069 21968 -3065
rect 8224 -3147 8300 -3137
rect 7783 -3151 8300 -3147
rect 7783 -3203 8236 -3151
rect 8288 -3203 8300 -3151
rect 20888 -3158 20965 -3157
rect 7783 -3204 8300 -3203
rect 7783 -3952 7840 -3204
rect 8224 -3216 8300 -3204
rect 20887 -3168 20965 -3158
rect 20887 -3224 20898 -3168
rect 20954 -3224 20965 -3168
rect 20887 -3235 20965 -3224
rect 20887 -3236 20963 -3235
rect 20918 -3309 20996 -3304
rect 21706 -3309 21764 -3069
rect 21890 -3077 21968 -3069
rect 20918 -3316 21764 -3309
rect 20918 -3368 20931 -3316
rect 20983 -3367 21764 -3316
rect 20983 -3368 20996 -3367
rect 20918 -3380 20996 -3368
rect 7781 -3965 7860 -3952
rect 7781 -4017 7793 -3965
rect 7845 -4017 7860 -3965
rect 7781 -4018 7860 -4017
rect 7781 -4024 7854 -4018
rect 7783 -4103 7840 -4024
rect 13580 -4108 13659 -4104
rect 13580 -4121 13674 -4108
rect 15592 -4121 15664 -4117
rect 959 -4142 1025 -4129
rect 959 -4194 966 -4142
rect 1018 -4194 1025 -4142
rect 13580 -4173 13591 -4121
rect 13643 -4173 13674 -4121
rect 15587 -4132 15664 -4121
rect 14513 -4140 14569 -4136
rect 13580 -4190 13674 -4173
rect 13592 -4191 13674 -4190
rect 959 -4206 1025 -4194
rect 966 -5262 1022 -4206
rect 8300 -4377 8373 -4362
rect 8300 -4429 8312 -4377
rect 8364 -4429 8373 -4377
rect 8300 -4444 8373 -4429
rect 8301 -5136 8366 -4444
rect 13609 -5136 13674 -4191
rect 14490 -4155 14577 -4140
rect 14490 -4207 14507 -4155
rect 14559 -4207 14577 -4155
rect 14490 -4222 14577 -4207
rect 15587 -4184 15606 -4132
rect 15658 -4184 15664 -4132
rect 15587 -4198 15664 -4184
rect 8301 -5201 13674 -5136
rect 961 -5274 1037 -5262
rect 961 -5326 973 -5274
rect 1025 -5326 1037 -5274
rect 961 -5338 1037 -5326
rect 14513 -5287 14569 -4222
rect 15587 -5153 15648 -4198
rect 20837 -4377 20906 -4361
rect 20837 -4429 20844 -4377
rect 20896 -4429 20906 -4377
rect 20837 -4447 20906 -4429
rect 20841 -4791 20902 -4447
rect 20841 -4852 20940 -4791
rect 20879 -5153 20940 -4852
rect 15587 -5214 20940 -5153
rect 24877 -5272 24933 -2737
rect 28409 -2940 28484 -2929
rect 28409 -2996 28417 -2940
rect 28473 -2996 28484 -2940
rect 28409 -3009 28484 -2996
rect 28407 -4131 28483 -4124
rect 28407 -4138 28509 -4131
rect 28407 -4190 28419 -4138
rect 28471 -4190 28509 -4138
rect 28407 -4203 28509 -4190
rect 28453 -5272 28509 -4203
rect 14513 -5301 14621 -5287
rect 14513 -5353 14556 -5301
rect 14608 -5353 14621 -5301
rect 14513 -5358 14621 -5353
rect 14544 -5367 14621 -5358
rect 21357 -5297 21434 -5289
rect 21761 -5297 21837 -5289
rect 21357 -5301 21837 -5297
rect 21357 -5302 21773 -5301
rect 21357 -5354 21369 -5302
rect 21421 -5353 21773 -5302
rect 21825 -5353 21837 -5301
rect 24877 -5328 28509 -5272
rect 21421 -5354 21837 -5353
rect 21357 -5356 21837 -5354
rect 21357 -5366 21434 -5356
rect 21761 -5365 21837 -5356
<< via2 >>
rect 956 2279 1012 2283
rect 956 2227 957 2279
rect 957 2227 1009 2279
rect 1009 2227 1012 2279
rect 13558 4216 13614 4218
rect 13558 4164 13560 4216
rect 13560 4164 13612 4216
rect 13612 4164 13614 4216
rect 13558 4162 13614 4164
rect 13596 3018 13652 3019
rect 13596 2966 13609 3018
rect 13609 2966 13652 3018
rect 13596 2963 13652 2966
rect 13786 2669 13842 2725
rect 944 1081 1000 1085
rect 944 1029 996 1081
rect 996 1029 1000 1081
rect 6706 6 6762 8
rect 6706 -46 6708 6
rect 6708 -46 6760 6
rect 6760 -46 6762 6
rect 6706 -48 6762 -46
rect 29789 2100 29845 2156
rect 13694 -2087 13750 -2084
rect 13694 -2139 13695 -2087
rect 13695 -2139 13747 -2087
rect 13747 -2139 13750 -2087
rect 13694 -2140 13750 -2139
rect 978 -2937 1034 -2935
rect 978 -2989 980 -2937
rect 980 -2989 1032 -2937
rect 1032 -2989 1034 -2937
rect 978 -2991 1034 -2989
rect 20898 -3171 20954 -3168
rect 20898 -3223 20899 -3171
rect 20899 -3223 20951 -3171
rect 20951 -3223 20954 -3171
rect 20898 -3224 20954 -3223
rect 28417 -2944 28473 -2940
rect 28417 -2996 28469 -2944
rect 28469 -2996 28473 -2944
<< metal3 >>
rect 13547 4219 13625 4229
rect 13516 4218 13845 4219
rect 13516 4162 13558 4218
rect 13614 4162 13845 4218
rect 13516 4160 13845 4162
rect 13547 4152 13625 4160
rect 13585 3019 13664 3030
rect 13585 2963 13596 3019
rect 13652 2963 13664 3019
rect 13585 2953 13664 2963
rect 13595 2744 13662 2953
rect 848 2677 13662 2744
rect 13786 2735 13845 4160
rect 848 2625 915 2677
rect -155 2558 915 2625
rect -155 -2925 -88 2558
rect 848 2293 915 2558
rect 13595 2571 13662 2677
rect 13776 2725 13852 2735
rect 13776 2669 13786 2725
rect 13842 2669 13852 2725
rect 13776 2659 13852 2669
rect 13595 2504 13757 2571
rect 848 2283 1029 2293
rect 848 2227 956 2283
rect 1012 2227 1029 2283
rect 848 2226 1029 2227
rect 917 1085 1011 1096
rect 917 1029 944 1085
rect 1000 1029 1011 1085
rect 917 1015 1011 1029
rect 917 9 977 1015
rect 6694 9 6775 19
rect 917 8 6775 9
rect 917 -48 6706 8
rect 6762 -48 6775 8
rect 917 -51 6775 -48
rect 6694 -59 6775 -51
rect 13690 -2073 13757 2504
rect 29794 2167 29851 2188
rect 29779 2156 29852 2167
rect 29779 2100 29789 2156
rect 29845 2100 29852 2156
rect 29779 2090 29852 2100
rect 13683 -2084 13761 -2073
rect 13683 -2140 13694 -2084
rect 13750 -2140 13761 -2084
rect 13683 -2151 13761 -2140
rect 966 -2925 1047 -2923
rect -155 -2935 1063 -2925
rect -155 -2991 978 -2935
rect 1034 -2991 1063 -2935
rect 28409 -2940 28484 -2929
rect 28409 -2943 28417 -2940
rect -155 -2992 1063 -2991
rect 966 -2998 1047 -2992
rect 28393 -2996 28417 -2943
rect 28473 -2943 28484 -2940
rect 28473 -2996 28596 -2943
rect 28393 -3000 28596 -2996
rect 28409 -3009 28596 -3000
rect 20888 -3167 20965 -3157
rect 28539 -3167 28596 -3009
rect 29794 -3167 29851 2090
rect 20888 -3168 29851 -3167
rect 20888 -3224 20898 -3168
rect 20954 -3224 29851 -3168
rect 20888 -3235 20965 -3224
use 3_inp_AND_magic  3_inp_AND_magic_0
timestamp 1713349043
transform 1 0 23744 0 1 3517
box -184 -1564 1665 536
use 3_inp_NOR  3_inp_NOR_0
timestamp 1713185578
transform 1 0 22550 0 -1 652
box -79 -2959 921 525
use buffer_magic  buffer_magic_0
timestamp 1713185578
transform 1 0 30999 0 1 3772
box 0 -989 1784 579
use buffer_magic  buffer_magic_1
timestamp 1713185578
transform 1 0 27126 0 1 3772
box 0 -989 1784 579
use buffer_magic  buffer_magic_2
timestamp 1713185578
transform 1 0 29071 0 1 3772
box 0 -989 1784 579
use DFF_magic  DFF_magic_0
timestamp 1713971515
transform 1 0 27541 0 1 866
box -2075 -819 5510 1706
use inverter_magic  inverter_magic_0
timestamp 1713185578
transform 1 0 25577 0 1 3473
box 0 -569 1108 580
use MDFF  MDFF_0
timestamp 1713277963
transform 1 0 6012 0 1 3477
box -6012 -8693 1961 -3553
use MDFF  MDFF_1
timestamp 1713277963
transform 1 0 20668 0 -1 -8671
box -6012 -8693 1961 -3553
use MDFF  MDFF_3
timestamp 1713277963
transform 1 0 6012 0 1 8693
box -6012 -8693 1961 -3553
use MDFF  MDFF_4
timestamp 1713277963
transform -1 0 8554 0 -1 -8671
box -6012 -8693 1961 -3553
use MDFF  MDFF_5
timestamp 1713277963
transform -1 0 8554 0 -1 -3454
box -6012 -8693 1961 -3553
use MDFF  MDFF_6
timestamp 1713277963
transform 1 0 20668 0 -1 -3454
box -6012 -8693 1961 -3553
use MDFF  MDFF_7
timestamp 1713277963
transform -1 0 23401 0 1 3477
box -6012 -8693 1961 -3553
use NAND_magic  NAND_magic_0
timestamp 1713185578
transform 1 0 23762 0 1 4959
box -14 -744 1108 536
use NOR_gate  NOR_gate_0
timestamp 1713185578
transform 1 0 21248 0 -1 795
box -72 -1005 1136 668
use NOR_gate  NOR_gate_1
timestamp 1713185578
transform 1 0 23537 0 -1 795
box -72 -1005 1136 668
<< labels >>
flabel nsubdiffcont 29127 4284 29127 4284 0 FreeSans 750 0 0 0 VDD
flabel psubdiffcont 28963 2824 28963 2824 0 FreeSans 750 0 0 0 VSS
flabel metal1 s 22386 3918 22386 3918 0 FreeSans 750 0 0 0 Q1
port 1 nsew
flabel metal1 s 15544 2250 15544 2250 0 FreeSans 750 0 0 0 D2_1
port 2 nsew
flabel metal1 s 6730 4120 6730 4120 0 FreeSans 750 0 0 0 Q2
port 3 nsew
flabel metal1 s 13693 2253 13693 2253 0 FreeSans 750 0 0 0 D2_2
port 4 nsew
flabel metal1 s 22483 -1060 22483 -1060 0 FreeSans 750 0 0 0 Q3
port 5 nsew
flabel metal1 s 15545 -2969 15545 -2969 0 FreeSans 750 0 0 0 D2_3
port 6 nsew
flabel metal1 s 21633 -3882 21633 -3882 0 FreeSans 750 0 0 0 Q4
port 7 nsew
flabel metal1 s 28540 -2228 28540 -2228 0 FreeSans 750 0 0 0 D2_4
port 8 nsew
flabel metal1 s 7827 -4093 7827 -4093 0 FreeSans 750 0 0 0 Q5
port 9 nsew
flabel metal1 s 870 -2229 870 -2229 0 FreeSans 750 0 0 0 D2_5
port 10 nsew
flabel metal1 s 6734 -1116 6734 -1116 0 FreeSans 750 0 0 0 Q6
port 11 nsew
flabel metal1 s 13696 -2961 13696 -2961 0 FreeSans 750 0 0 0 D2_6
port 12 nsew
flabel metal1 s 7769 1221 7769 1221 0 FreeSans 750 0 0 0 Q7
port 13 nsew
flabel metal1 s 871 2982 871 2982 0 FreeSans 750 0 0 0 D2_7
port 14 nsew
flabel metal1 s 19167 -2918 19167 -2918 0 FreeSans 750 0 0 0 G-CLK
port 15 nsew
flabel metal1 s 26593 3532 26593 3532 0 FreeSans 750 0 0 0 LD
port 16 nsew
<< end >>
