magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2088 -2044 2228 3044
<< mvnmos >>
rect 0 0 140 1000
<< mvndiff >>
rect -88 987 0 1000
rect -88 941 -75 987
rect -29 941 0 987
rect -88 884 0 941
rect -88 838 -75 884
rect -29 838 0 884
rect -88 781 0 838
rect -88 735 -75 781
rect -29 735 0 781
rect -88 678 0 735
rect -88 632 -75 678
rect -29 632 0 678
rect -88 575 0 632
rect -88 529 -75 575
rect -29 529 0 575
rect -88 472 0 529
rect -88 426 -75 472
rect -29 426 0 472
rect -88 369 0 426
rect -88 323 -75 369
rect -29 323 0 369
rect -88 266 0 323
rect -88 220 -75 266
rect -29 220 0 266
rect -88 163 0 220
rect -88 117 -75 163
rect -29 117 0 163
rect -88 59 0 117
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 140 987 228 1000
rect 140 941 169 987
rect 215 941 228 987
rect 140 884 228 941
rect 140 838 169 884
rect 215 838 228 884
rect 140 781 228 838
rect 140 735 169 781
rect 215 735 228 781
rect 140 678 228 735
rect 140 632 169 678
rect 215 632 228 678
rect 140 575 228 632
rect 140 529 169 575
rect 215 529 228 575
rect 140 472 228 529
rect 140 426 169 472
rect 215 426 228 472
rect 140 369 228 426
rect 140 323 169 369
rect 215 323 228 369
rect 140 266 228 323
rect 140 220 169 266
rect 215 220 228 266
rect 140 163 228 220
rect 140 117 169 163
rect 215 117 228 163
rect 140 59 228 117
rect 140 13 169 59
rect 215 13 228 59
rect 140 0 228 13
<< mvndiffc >>
rect -75 941 -29 987
rect -75 838 -29 884
rect -75 735 -29 781
rect -75 632 -29 678
rect -75 529 -29 575
rect -75 426 -29 472
rect -75 323 -29 369
rect -75 220 -29 266
rect -75 117 -29 163
rect -75 13 -29 59
rect 169 941 215 987
rect 169 838 215 884
rect 169 735 215 781
rect 169 632 215 678
rect 169 529 215 575
rect 169 426 215 472
rect 169 323 215 369
rect 169 220 215 266
rect 169 117 215 163
rect 169 13 215 59
<< polysilicon >>
rect 0 1000 140 1044
rect 0 -44 140 0
<< metal1 >>
rect -75 987 -29 1000
rect -75 884 -29 941
rect -75 781 -29 838
rect -75 678 -29 735
rect -75 575 -29 632
rect -75 472 -29 529
rect -75 369 -29 426
rect -75 266 -29 323
rect -75 163 -29 220
rect -75 59 -29 117
rect -75 0 -29 13
rect 169 987 215 1000
rect 169 884 215 941
rect 169 781 215 838
rect 169 678 215 735
rect 169 575 215 632
rect 169 472 215 529
rect 169 369 215 426
rect 169 266 215 323
rect 169 163 215 220
rect 169 59 215 117
rect 169 0 215 13
<< labels >>
rlabel metal1 192 500 192 500 4 D
rlabel metal1 -52 500 -52 500 4 S
<< end >>
