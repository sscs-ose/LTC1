magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2032 11097 3032 71968
<< psubdiff >>
rect 0 69778 1000 69968
rect 0 13287 93 69778
rect 907 13287 1000 69778
rect 0 13097 1000 13287
<< metal1 >>
rect -32 69789 1032 69957
rect -32 13276 14 69789
rect 82 63646 918 64954
rect 82 49240 918 50548
rect 986 13276 1032 69789
rect -32 13108 1032 13276
<< metal2 >>
rect 0 63600 1000 65000
rect 0 49200 1000 50600
<< metal3 >>
rect 0 63600 1000 65000
rect 0 49200 1000 50600
use M1_PSUB_CDNS_690335831656  M1_PSUB_CDNS_690335831656_0
timestamp 1713338890
transform 1 0 952 0 1 41524
box -45 -28395 45 28395
use M1_PSUB_CDNS_690335831656  M1_PSUB_CDNS_690335831656_1
timestamp 1713338890
transform -1 0 48 0 1 41524
box -45 -28395 45 28395
use M1_PSUB_CDNS_6903358316578  M1_PSUB_CDNS_6903358316578_0
timestamp 1713338890
transform 1 0 501 0 1 69873
box -345 -95 345 95
use M1_PSUB_CDNS_6903358316578  M1_PSUB_CDNS_6903358316578_1
timestamp 1713338890
transform 1 0 501 0 -1 13192
box -345 -95 345 95
use M2_M1_CDNS_69033583165699  M2_M1_CDNS_69033583165699_0
timestamp 1713338890
transform 1 0 506 0 1 64300
box -286 -534 286 534
use M2_M1_CDNS_69033583165699  M2_M1_CDNS_69033583165699_1
timestamp 1713338890
transform 1 0 498 0 1 49894
box -286 -534 286 534
use M3_M2_CDNS_69033583165698  M3_M2_CDNS_69033583165698_0
timestamp 1713338890
transform 1 0 506 0 1 64300
box -286 -534 286 534
use M3_M2_CDNS_69033583165698  M3_M2_CDNS_69033583165698_1
timestamp 1713338890
transform 1 0 498 0 1 49894
box -286 -534 286 534
use POLY_SUB_FILL_3  POLY_SUB_FILL_3_0
array 0 0 0 0 96 574
timestamp 1713338890
transform 1 0 187 0 1 13813
box -127 -235 772 615
<< labels >>
rlabel metal3 s 498 64258 498 64258 4 VSS
port 1 nsew
rlabel metal3 s 510 50023 510 50023 4 VSS
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1000 70000
<< end >>
