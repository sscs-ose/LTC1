magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -2501 -1019 2501 1019
<< metal1 >>
rect -1501 13 1501 19
rect -1501 -13 -1495 13
rect -1469 -13 -1419 13
rect -1393 -13 -1343 13
rect -1317 -13 -1267 13
rect -1241 -13 -1191 13
rect -1165 -13 -1115 13
rect -1089 -13 -1039 13
rect -1013 -13 -963 13
rect -937 -13 -887 13
rect -861 -13 -811 13
rect -785 -13 -735 13
rect -709 -13 -659 13
rect -633 -13 -583 13
rect -557 -13 -507 13
rect -481 -13 -431 13
rect -405 -13 -355 13
rect -329 -13 -279 13
rect -253 -13 -203 13
rect -177 -13 -127 13
rect -101 -13 -51 13
rect -25 -13 25 13
rect 51 -13 101 13
rect 127 -13 177 13
rect 203 -13 253 13
rect 279 -13 329 13
rect 355 -13 405 13
rect 431 -13 481 13
rect 507 -13 557 13
rect 583 -13 633 13
rect 659 -13 709 13
rect 735 -13 785 13
rect 811 -13 861 13
rect 887 -13 937 13
rect 963 -13 1013 13
rect 1039 -13 1089 13
rect 1115 -13 1165 13
rect 1191 -13 1241 13
rect 1267 -13 1317 13
rect 1343 -13 1393 13
rect 1419 -13 1469 13
rect 1495 -13 1501 13
rect -1501 -19 1501 -13
<< via1 >>
rect -1495 -13 -1469 13
rect -1419 -13 -1393 13
rect -1343 -13 -1317 13
rect -1267 -13 -1241 13
rect -1191 -13 -1165 13
rect -1115 -13 -1089 13
rect -1039 -13 -1013 13
rect -963 -13 -937 13
rect -887 -13 -861 13
rect -811 -13 -785 13
rect -735 -13 -709 13
rect -659 -13 -633 13
rect -583 -13 -557 13
rect -507 -13 -481 13
rect -431 -13 -405 13
rect -355 -13 -329 13
rect -279 -13 -253 13
rect -203 -13 -177 13
rect -127 -13 -101 13
rect -51 -13 -25 13
rect 25 -13 51 13
rect 101 -13 127 13
rect 177 -13 203 13
rect 253 -13 279 13
rect 329 -13 355 13
rect 405 -13 431 13
rect 481 -13 507 13
rect 557 -13 583 13
rect 633 -13 659 13
rect 709 -13 735 13
rect 785 -13 811 13
rect 861 -13 887 13
rect 937 -13 963 13
rect 1013 -13 1039 13
rect 1089 -13 1115 13
rect 1165 -13 1191 13
rect 1241 -13 1267 13
rect 1317 -13 1343 13
rect 1393 -13 1419 13
rect 1469 -13 1495 13
<< metal2 >>
rect -1501 13 1501 19
rect -1501 -13 -1495 13
rect -1469 -13 -1419 13
rect -1393 -13 -1343 13
rect -1317 -13 -1267 13
rect -1241 -13 -1191 13
rect -1165 -13 -1115 13
rect -1089 -13 -1039 13
rect -1013 -13 -963 13
rect -937 -13 -887 13
rect -861 -13 -811 13
rect -785 -13 -735 13
rect -709 -13 -659 13
rect -633 -13 -583 13
rect -557 -13 -507 13
rect -481 -13 -431 13
rect -405 -13 -355 13
rect -329 -13 -279 13
rect -253 -13 -203 13
rect -177 -13 -127 13
rect -101 -13 -51 13
rect -25 -13 25 13
rect 51 -13 101 13
rect 127 -13 177 13
rect 203 -13 253 13
rect 279 -13 329 13
rect 355 -13 405 13
rect 431 -13 481 13
rect 507 -13 557 13
rect 583 -13 633 13
rect 659 -13 709 13
rect 735 -13 785 13
rect 811 -13 861 13
rect 887 -13 937 13
rect 963 -13 1013 13
rect 1039 -13 1089 13
rect 1115 -13 1165 13
rect 1191 -13 1241 13
rect 1267 -13 1317 13
rect 1343 -13 1393 13
rect 1419 -13 1469 13
rect 1495 -13 1501 13
rect -1501 -19 1501 -13
<< end >>
