magic
tech gf180mcuC
magscale 1 10
timestamp 1693477706
<< nwell >>
rect -60 908 881 1080
<< psubdiff >>
rect -229 1208 1036 1236
rect -229 1206 -56 1208
rect -229 1142 -212 1206
rect -142 1144 -56 1206
rect 14 1144 69 1208
rect 139 1144 194 1208
rect 264 1144 319 1208
rect 389 1144 444 1208
rect 514 1144 569 1208
rect 639 1144 694 1208
rect 764 1144 819 1208
rect 889 1144 944 1208
rect 1014 1144 1036 1208
rect -142 1142 1036 1144
rect -229 1119 1036 1142
rect -229 997 -120 1119
rect -229 933 -211 997
rect -141 933 -120 997
rect 927 1005 1036 1119
rect -229 862 -120 933
rect 927 942 947 1005
rect 1016 942 1036 1005
rect -229 798 -211 862
rect -141 798 -120 862
rect -229 727 -120 798
rect -229 663 -211 727
rect -141 663 -120 727
rect -229 592 -120 663
rect -229 528 -211 592
rect -141 528 -120 592
rect -229 457 -120 528
rect -229 393 -211 457
rect -141 393 -120 457
rect -229 322 -120 393
rect -229 258 -211 322
rect -141 258 -120 322
rect -229 187 -120 258
rect 927 870 1036 942
rect 927 807 947 870
rect 1016 807 1036 870
rect 927 735 1036 807
rect 927 672 947 735
rect 1016 672 1036 735
rect 927 600 1036 672
rect 927 537 947 600
rect 1016 537 1036 600
rect 927 465 1036 537
rect 927 402 947 465
rect 1016 402 1036 465
rect 927 330 1036 402
rect 927 267 947 330
rect 1016 267 1036 330
rect -229 123 -211 187
rect -141 123 -120 187
rect -229 52 -120 123
rect 927 195 1036 267
rect 927 132 947 195
rect 1016 132 1036 195
rect -229 -12 -211 52
rect -141 -12 -120 52
rect -229 -83 -120 -12
rect -229 -147 -211 -83
rect -141 -147 -120 -83
rect -229 -218 -120 -147
rect -229 -282 -211 -218
rect -141 -282 -120 -218
rect -229 -321 -120 -282
rect 927 60 1036 132
rect 927 -3 947 60
rect 1016 -3 1036 60
rect 927 -75 1036 -3
rect 927 -138 947 -75
rect 1016 -138 1036 -75
rect 927 -210 1036 -138
rect 927 -273 947 -210
rect 1016 -273 1036 -210
rect 927 -321 1036 -273
rect -229 -345 1036 -321
rect -229 -349 947 -345
rect -229 -412 -208 -349
rect -139 -412 -83 -349
rect -14 -412 42 -349
rect 111 -412 167 -349
rect 236 -412 292 -349
rect 361 -412 417 -349
rect 486 -412 542 -349
rect 611 -412 667 -349
rect 736 -412 792 -349
rect 861 -408 947 -349
rect 1016 -408 1036 -345
rect 861 -412 1036 -408
rect -229 -438 1036 -412
<< nsubdiff >>
rect -9 972 823 986
rect -9 922 11 972
rect 60 922 112 972
rect 161 922 213 972
rect 262 922 314 972
rect 363 922 415 972
rect 464 922 516 972
rect 565 922 617 972
rect 666 922 718 972
rect 767 922 823 972
rect -9 908 823 922
<< psubdiffcont >>
rect -212 1142 -142 1206
rect -56 1144 14 1208
rect 69 1144 139 1208
rect 194 1144 264 1208
rect 319 1144 389 1208
rect 444 1144 514 1208
rect 569 1144 639 1208
rect 694 1144 764 1208
rect 819 1144 889 1208
rect 944 1144 1014 1208
rect -211 933 -141 997
rect 947 942 1016 1005
rect -211 798 -141 862
rect -211 663 -141 727
rect -211 528 -141 592
rect -211 393 -141 457
rect -211 258 -141 322
rect 947 807 1016 870
rect 947 672 1016 735
rect 947 537 1016 600
rect 947 402 1016 465
rect 947 267 1016 330
rect -211 123 -141 187
rect 947 132 1016 195
rect -211 -12 -141 52
rect -211 -147 -141 -83
rect -211 -282 -141 -218
rect 947 -3 1016 60
rect 947 -138 1016 -75
rect 947 -273 1016 -210
rect -208 -412 -139 -349
rect -83 -412 -14 -349
rect 42 -412 111 -349
rect 167 -412 236 -349
rect 292 -412 361 -349
rect 417 -412 486 -349
rect 542 -412 611 -349
rect 667 -412 736 -349
rect 792 -412 861 -349
rect 947 -408 1016 -345
<< nsubdiffcont >>
rect 11 922 60 972
rect 112 922 161 972
rect 213 922 262 972
rect 314 922 363 972
rect 415 922 464 972
rect 516 922 565 972
rect 617 922 666 972
rect 718 922 767 972
<< polysilicon >>
rect 114 216 184 247
rect 51 203 184 216
rect 51 148 66 203
rect 123 197 184 203
rect 288 197 358 246
rect 462 197 532 245
rect 636 197 706 241
rect 123 148 706 197
rect 51 144 706 148
rect 51 134 184 144
rect 114 103 184 134
rect 288 102 358 144
rect 462 101 532 144
rect 636 97 706 144
<< polycontact >>
rect 66 148 123 203
<< metal1 >>
rect -229 1208 1036 1236
rect -229 1206 -56 1208
rect -229 1142 -212 1206
rect -142 1144 -56 1206
rect 14 1144 69 1208
rect 139 1144 194 1208
rect 264 1144 319 1208
rect 389 1144 444 1208
rect 514 1144 569 1208
rect 639 1144 694 1208
rect 764 1144 819 1208
rect 889 1144 944 1208
rect 1014 1144 1036 1208
rect -142 1142 1036 1144
rect -229 1119 1036 1142
rect -229 997 -120 1119
rect -229 933 -211 997
rect -141 933 -120 997
rect 927 1005 1036 1119
rect -229 862 -120 933
rect -9 972 823 986
rect -9 922 11 972
rect 60 922 112 972
rect 161 922 213 972
rect 262 922 314 972
rect 363 922 415 972
rect 464 922 516 972
rect 565 922 617 972
rect 666 922 718 972
rect 767 922 823 972
rect -9 908 823 922
rect 927 942 947 1005
rect 1016 942 1036 1005
rect -229 798 -211 862
rect -141 798 -120 862
rect 39 825 85 908
rect 387 829 433 908
rect 735 827 781 908
rect 927 870 1036 942
rect -229 727 -120 798
rect -229 663 -211 727
rect -141 663 -120 727
rect -229 592 -120 663
rect -229 528 -211 592
rect -141 528 -120 592
rect -229 457 -120 528
rect -229 393 -211 457
rect -141 393 -120 457
rect -229 322 -120 393
rect -229 258 -211 322
rect -141 258 -120 322
rect 927 807 947 870
rect 1016 807 1036 870
rect 927 735 1036 807
rect 927 672 947 735
rect 1016 672 1036 735
rect 927 600 1036 672
rect 927 537 947 600
rect 1016 537 1036 600
rect 927 465 1036 537
rect 927 402 947 465
rect 1016 402 1036 465
rect 927 330 1036 402
rect -229 187 -120 258
rect 51 203 134 216
rect 51 198 66 203
rect -229 123 -211 187
rect -141 123 -120 187
rect 7 152 66 198
rect 51 148 66 152
rect 123 148 134 203
rect 51 134 134 148
rect 213 190 259 302
rect 561 190 607 293
rect 927 267 947 330
rect 1016 267 1036 330
rect 927 195 1036 267
rect 213 144 766 190
rect -229 52 -120 123
rect -229 -12 -211 52
rect -141 -12 -120 52
rect 213 45 259 144
rect 561 36 607 144
rect 927 132 947 195
rect 1016 132 1036 195
rect 927 60 1036 132
rect -229 -83 -120 -12
rect -229 -147 -211 -83
rect -141 -147 -120 -83
rect -229 -218 -120 -147
rect 927 -3 947 60
rect 1016 -3 1036 60
rect 927 -75 1036 -3
rect 927 -138 947 -75
rect 1016 -138 1036 -75
rect -229 -282 -211 -218
rect -141 -282 -120 -218
rect -229 -321 -120 -282
rect 39 -321 85 -194
rect 387 -321 433 -188
rect 735 -321 781 -194
rect 927 -210 1036 -138
rect 927 -273 947 -210
rect 1016 -273 1036 -210
rect 927 -321 1036 -273
rect -229 -345 1036 -321
rect -229 -349 947 -345
rect -229 -412 -208 -349
rect -139 -412 -83 -349
rect -14 -412 42 -349
rect 111 -412 167 -349
rect 236 -412 292 -349
rect 361 -412 417 -349
rect 486 -412 542 -349
rect 611 -412 667 -349
rect 736 -412 792 -349
rect 861 -408 947 -349
rect 1016 -408 1036 -345
rect 861 -412 1036 -408
rect -229 -438 1036 -412
use nmos_3p3_S7UZWU  nmos_3p3_S7UZWU_0
timestamp 1693477706
transform 1 0 410 0 1 -78
box -408 -208 408 208
use pmos_3p3_MD4UPK  pmos_3p3_MD4UPK_0
timestamp 1693477706
transform 1 0 410 0 1 562
box -470 -410 470 410
<< labels >>
flabel metal1 277 937 277 937 0 FreeSans 320 0 0 0 VDD
port 0 nsew
flabel metal1 30 173 30 173 0 FreeSans 320 0 0 0 IN
port 1 nsew
flabel metal1 736 167 736 167 0 FreeSans 320 0 0 0 OUT
port 2 nsew
flabel metal1 403 -309 403 -309 0 FreeSans 320 0 0 0 VSS
port 4 nsew
<< end >>
