magic
tech gf180mcuC
magscale 1 10
timestamp 1692950850
<< nwell >>
rect -817 1943 -712 1945
rect -3723 1885 -2663 1906
rect -817 1905 243 1943
<< psubdiff >>
rect -4178 4062 2072 4075
rect -4178 4006 -4129 4062
rect -4074 4006 -3979 4062
rect -3924 4006 -3829 4062
rect -3774 4006 -3679 4062
rect -3624 4006 -3529 4062
rect -3474 4006 -3379 4062
rect -3324 4006 -3229 4062
rect -3174 4006 -3079 4062
rect -3024 4006 -2929 4062
rect -2874 4006 -2779 4062
rect -2724 4006 -2629 4062
rect -2574 4006 -2479 4062
rect -2424 4006 -2329 4062
rect -2274 4006 -2179 4062
rect -2124 4006 -2029 4062
rect -1974 4006 -1879 4062
rect -1824 4006 -1729 4062
rect -1674 4006 -1579 4062
rect -1524 4006 -1429 4062
rect -1374 4006 -1279 4062
rect -1224 4006 -1129 4062
rect -1074 4006 -979 4062
rect -924 4006 -829 4062
rect -774 4006 -679 4062
rect -624 4006 -529 4062
rect -474 4006 -379 4062
rect -324 4006 -229 4062
rect -174 4006 -79 4062
rect -24 4006 71 4062
rect 126 4006 221 4062
rect 276 4006 371 4062
rect 426 4006 521 4062
rect 576 4006 671 4062
rect 726 4006 821 4062
rect 876 4006 971 4062
rect 1026 4006 1121 4062
rect 1176 4006 1271 4062
rect 1326 4006 1421 4062
rect 1476 4006 1571 4062
rect 1626 4006 1721 4062
rect 1776 4006 1871 4062
rect 1926 4035 2072 4062
rect 1926 4006 2000 4035
rect -4178 3985 2000 4006
rect -4178 3955 -4088 3985
rect -4178 3899 -4162 3955
rect -4107 3899 -4088 3955
rect -4178 3805 -4088 3899
rect -4178 3749 -4162 3805
rect -4107 3749 -4088 3805
rect -4178 3655 -4088 3749
rect -4178 3599 -4162 3655
rect -4107 3599 -4088 3655
rect -4178 3505 -4088 3599
rect -4178 3449 -4162 3505
rect -4107 3449 -4088 3505
rect -4178 3355 -4088 3449
rect -4178 3299 -4162 3355
rect -4107 3299 -4088 3355
rect -4178 3205 -4088 3299
rect -4178 3149 -4162 3205
rect -4107 3149 -4088 3205
rect -4178 3055 -4088 3149
rect -4178 2999 -4162 3055
rect -4107 2999 -4088 3055
rect -4178 2905 -4088 2999
rect -4178 2849 -4162 2905
rect -4107 2849 -4088 2905
rect -4178 2755 -4088 2849
rect -4178 2699 -4162 2755
rect -4107 2699 -4088 2755
rect -4178 2605 -4088 2699
rect -4178 2549 -4162 2605
rect -4107 2549 -4088 2605
rect -4178 2455 -4088 2549
rect -4178 2399 -4162 2455
rect -4107 2399 -4088 2455
rect -4178 2305 -4088 2399
rect -4178 2249 -4162 2305
rect -4107 2249 -4088 2305
rect -4178 2155 -4088 2249
rect -4178 2099 -4162 2155
rect -4107 2099 -4088 2155
rect -4178 2005 -4088 2099
rect -4178 1949 -4162 2005
rect -4107 1949 -4088 2005
rect -4178 1855 -4088 1949
rect -4178 1799 -4162 1855
rect -4107 1799 -4088 1855
rect -4178 1705 -4088 1799
rect -4178 1649 -4162 1705
rect -4107 1649 -4088 1705
rect -4178 1555 -4088 1649
rect -4178 1499 -4162 1555
rect -4107 1499 -4088 1555
rect -4178 1405 -4088 1499
rect -4178 1349 -4162 1405
rect -4107 1349 -4088 1405
rect -4178 1255 -4088 1349
rect -4178 1199 -4162 1255
rect -4107 1199 -4088 1255
rect -4178 1105 -4088 1199
rect -4178 1049 -4162 1105
rect -4107 1049 -4088 1105
rect -4178 955 -4088 1049
rect -4178 899 -4162 955
rect -4107 899 -4088 955
rect -4178 805 -4088 899
rect -4178 749 -4162 805
rect -4107 749 -4088 805
rect -4178 655 -4088 749
rect -4178 599 -4162 655
rect -4107 599 -4088 655
rect -4178 505 -4088 599
rect -4178 449 -4162 505
rect -4107 449 -4088 505
rect -4178 355 -4088 449
rect -4178 299 -4162 355
rect -4107 299 -4088 355
rect -4178 205 -4088 299
rect -4178 149 -4162 205
rect -4107 149 -4088 205
rect -4178 55 -4088 149
rect -4178 -1 -4162 55
rect -4107 -1 -4088 55
rect -4178 -115 -4088 -1
rect 1982 3979 2000 3985
rect 2055 3979 2072 4035
rect 1982 3885 2072 3979
rect 1982 3829 2000 3885
rect 2055 3829 2072 3885
rect 1982 3735 2072 3829
rect 1982 3679 2000 3735
rect 2055 3679 2072 3735
rect 1982 3585 2072 3679
rect 1982 3529 2000 3585
rect 2055 3529 2072 3585
rect 1982 3435 2072 3529
rect 1982 3379 2000 3435
rect 2055 3379 2072 3435
rect 1982 3285 2072 3379
rect 1982 3229 2000 3285
rect 2055 3229 2072 3285
rect 1982 3135 2072 3229
rect 1982 3079 2000 3135
rect 2055 3079 2072 3135
rect 1982 2985 2072 3079
rect 1982 2929 2000 2985
rect 2055 2929 2072 2985
rect 1982 2835 2072 2929
rect 1982 2779 2000 2835
rect 2055 2779 2072 2835
rect 1982 2685 2072 2779
rect 1982 2629 2000 2685
rect 2055 2629 2072 2685
rect 1982 2535 2072 2629
rect 1982 2479 2000 2535
rect 2055 2479 2072 2535
rect 1982 2385 2072 2479
rect 1982 2329 2000 2385
rect 2055 2329 2072 2385
rect 1982 2235 2072 2329
rect 1982 2179 2000 2235
rect 2055 2179 2072 2235
rect 1982 2085 2072 2179
rect 1982 2029 2000 2085
rect 2055 2029 2072 2085
rect 1982 1935 2072 2029
rect 1982 1879 2000 1935
rect 2055 1879 2072 1935
rect 1982 1785 2072 1879
rect 1982 1729 2000 1785
rect 2055 1729 2072 1785
rect 1982 1635 2072 1729
rect 1982 1579 2000 1635
rect 2055 1579 2072 1635
rect 1982 1485 2072 1579
rect 1982 1429 2000 1485
rect 2055 1429 2072 1485
rect 1982 1335 2072 1429
rect 1982 1279 2000 1335
rect 2055 1279 2072 1335
rect 1982 1185 2072 1279
rect 1982 1129 2000 1185
rect 2055 1129 2072 1185
rect 1982 1035 2072 1129
rect 1982 979 2000 1035
rect 2055 979 2072 1035
rect 1982 885 2072 979
rect 1982 829 2000 885
rect 2055 829 2072 885
rect 1982 735 2072 829
rect 1982 679 2000 735
rect 2055 679 2072 735
rect 1982 585 2072 679
rect 1982 529 2000 585
rect 2055 529 2072 585
rect 1982 435 2072 529
rect 1982 379 2000 435
rect 2055 379 2072 435
rect 1982 285 2072 379
rect 1982 229 2000 285
rect 2055 229 2072 285
rect 1982 135 2072 229
rect 1982 79 2000 135
rect 2055 79 2072 135
rect 1982 -15 2072 79
rect 1982 -71 2000 -15
rect 2055 -71 2072 -15
rect 1982 -115 2072 -71
rect -4178 -131 2072 -115
rect -4178 -187 -4062 -131
rect -4007 -187 -3912 -131
rect -3857 -187 -3762 -131
rect -3707 -187 -3612 -131
rect -3557 -187 -3462 -131
rect -3407 -187 -3312 -131
rect -3257 -187 -3162 -131
rect -3107 -187 -3012 -131
rect -2957 -187 -2862 -131
rect -2807 -187 -2712 -131
rect -2657 -187 -2562 -131
rect -2507 -187 -2412 -131
rect -2357 -187 -2262 -131
rect -2207 -187 -2112 -131
rect -2057 -187 -1962 -131
rect -1907 -187 -1812 -131
rect -1757 -187 -1662 -131
rect -1607 -187 -1512 -131
rect -1457 -187 -1362 -131
rect -1307 -187 -1212 -131
rect -1157 -187 -1062 -131
rect -1007 -187 -912 -131
rect -857 -187 -762 -131
rect -707 -187 -612 -131
rect -557 -187 -462 -131
rect -407 -187 -312 -131
rect -257 -187 -162 -131
rect -107 -187 -12 -131
rect 43 -187 138 -131
rect 193 -187 288 -131
rect 343 -187 438 -131
rect 493 -187 588 -131
rect 643 -187 738 -131
rect 793 -187 888 -131
rect 943 -187 1038 -131
rect 1093 -187 1188 -131
rect 1243 -187 1338 -131
rect 1393 -187 1488 -131
rect 1543 -187 1638 -131
rect 1693 -187 1788 -131
rect 1843 -187 1938 -131
rect 1993 -187 2072 -131
rect -4178 -205 2072 -187
<< psubdiffcont >>
rect -4129 4006 -4074 4062
rect -3979 4006 -3924 4062
rect -3829 4006 -3774 4062
rect -3679 4006 -3624 4062
rect -3529 4006 -3474 4062
rect -3379 4006 -3324 4062
rect -3229 4006 -3174 4062
rect -3079 4006 -3024 4062
rect -2929 4006 -2874 4062
rect -2779 4006 -2724 4062
rect -2629 4006 -2574 4062
rect -2479 4006 -2424 4062
rect -2329 4006 -2274 4062
rect -2179 4006 -2124 4062
rect -2029 4006 -1974 4062
rect -1879 4006 -1824 4062
rect -1729 4006 -1674 4062
rect -1579 4006 -1524 4062
rect -1429 4006 -1374 4062
rect -1279 4006 -1224 4062
rect -1129 4006 -1074 4062
rect -979 4006 -924 4062
rect -829 4006 -774 4062
rect -679 4006 -624 4062
rect -529 4006 -474 4062
rect -379 4006 -324 4062
rect -229 4006 -174 4062
rect -79 4006 -24 4062
rect 71 4006 126 4062
rect 221 4006 276 4062
rect 371 4006 426 4062
rect 521 4006 576 4062
rect 671 4006 726 4062
rect 821 4006 876 4062
rect 971 4006 1026 4062
rect 1121 4006 1176 4062
rect 1271 4006 1326 4062
rect 1421 4006 1476 4062
rect 1571 4006 1626 4062
rect 1721 4006 1776 4062
rect 1871 4006 1926 4062
rect -4162 3899 -4107 3955
rect -4162 3749 -4107 3805
rect -4162 3599 -4107 3655
rect -4162 3449 -4107 3505
rect -4162 3299 -4107 3355
rect -4162 3149 -4107 3205
rect -4162 2999 -4107 3055
rect -4162 2849 -4107 2905
rect -4162 2699 -4107 2755
rect -4162 2549 -4107 2605
rect -4162 2399 -4107 2455
rect -4162 2249 -4107 2305
rect -4162 2099 -4107 2155
rect -4162 1949 -4107 2005
rect -4162 1799 -4107 1855
rect -4162 1649 -4107 1705
rect -4162 1499 -4107 1555
rect -4162 1349 -4107 1405
rect -4162 1199 -4107 1255
rect -4162 1049 -4107 1105
rect -4162 899 -4107 955
rect -4162 749 -4107 805
rect -4162 599 -4107 655
rect -4162 449 -4107 505
rect -4162 299 -4107 355
rect -4162 149 -4107 205
rect -4162 -1 -4107 55
rect 2000 3979 2055 4035
rect 2000 3829 2055 3885
rect 2000 3679 2055 3735
rect 2000 3529 2055 3585
rect 2000 3379 2055 3435
rect 2000 3229 2055 3285
rect 2000 3079 2055 3135
rect 2000 2929 2055 2985
rect 2000 2779 2055 2835
rect 2000 2629 2055 2685
rect 2000 2479 2055 2535
rect 2000 2329 2055 2385
rect 2000 2179 2055 2235
rect 2000 2029 2055 2085
rect 2000 1879 2055 1935
rect 2000 1729 2055 1785
rect 2000 1579 2055 1635
rect 2000 1429 2055 1485
rect 2000 1279 2055 1335
rect 2000 1129 2055 1185
rect 2000 979 2055 1035
rect 2000 829 2055 885
rect 2000 679 2055 735
rect 2000 529 2055 585
rect 2000 379 2055 435
rect 2000 229 2055 285
rect 2000 79 2055 135
rect 2000 -71 2055 -15
rect -4062 -187 -4007 -131
rect -3912 -187 -3857 -131
rect -3762 -187 -3707 -131
rect -3612 -187 -3557 -131
rect -3462 -187 -3407 -131
rect -3312 -187 -3257 -131
rect -3162 -187 -3107 -131
rect -3012 -187 -2957 -131
rect -2862 -187 -2807 -131
rect -2712 -187 -2657 -131
rect -2562 -187 -2507 -131
rect -2412 -187 -2357 -131
rect -2262 -187 -2207 -131
rect -2112 -187 -2057 -131
rect -1962 -187 -1907 -131
rect -1812 -187 -1757 -131
rect -1662 -187 -1607 -131
rect -1512 -187 -1457 -131
rect -1362 -187 -1307 -131
rect -1212 -187 -1157 -131
rect -1062 -187 -1007 -131
rect -912 -187 -857 -131
rect -762 -187 -707 -131
rect -612 -187 -557 -131
rect -462 -187 -407 -131
rect -312 -187 -257 -131
rect -162 -187 -107 -131
rect -12 -187 43 -131
rect 138 -187 193 -131
rect 288 -187 343 -131
rect 438 -187 493 -131
rect 588 -187 643 -131
rect 738 -187 793 -131
rect 888 -187 943 -131
rect 1038 -187 1093 -131
rect 1188 -187 1243 -131
rect 1338 -187 1393 -131
rect 1488 -187 1543 -131
rect 1638 -187 1693 -131
rect 1788 -187 1843 -131
rect 1938 -187 1993 -131
<< metal1 >>
rect -4189 4062 2082 4087
rect -4189 4006 -4129 4062
rect -4074 4006 -3979 4062
rect -3924 4006 -3829 4062
rect -3774 4006 -3679 4062
rect -3624 4006 -3529 4062
rect -3474 4006 -3379 4062
rect -3324 4006 -3229 4062
rect -3174 4006 -3079 4062
rect -3024 4006 -2929 4062
rect -2874 4006 -2779 4062
rect -2724 4006 -2629 4062
rect -2574 4006 -2479 4062
rect -2424 4006 -2329 4062
rect -2274 4006 -2179 4062
rect -2124 4006 -2029 4062
rect -1974 4006 -1879 4062
rect -1824 4006 -1729 4062
rect -1674 4006 -1579 4062
rect -1524 4006 -1429 4062
rect -1374 4006 -1279 4062
rect -1224 4006 -1129 4062
rect -1074 4006 -979 4062
rect -924 4006 -829 4062
rect -774 4006 -679 4062
rect -624 4006 -529 4062
rect -474 4006 -379 4062
rect -324 4006 -229 4062
rect -174 4006 -79 4062
rect -24 4006 71 4062
rect 126 4006 221 4062
rect 276 4006 371 4062
rect 426 4006 521 4062
rect 576 4006 671 4062
rect 726 4006 821 4062
rect 876 4006 971 4062
rect 1026 4006 1121 4062
rect 1176 4006 1271 4062
rect 1326 4006 1421 4062
rect 1476 4006 1571 4062
rect 1626 4006 1721 4062
rect 1776 4006 1871 4062
rect 1926 4035 2082 4062
rect 1926 4006 2000 4035
rect -4189 3979 2000 4006
rect 2055 3979 2082 4035
rect -4189 3964 2082 3979
rect -4189 3955 -4066 3964
rect -4189 3899 -4162 3955
rect -4107 3899 -4066 3955
rect -4189 3805 -4066 3899
rect -4189 3749 -4162 3805
rect -4107 3749 -4066 3805
rect 1959 3885 2082 3964
rect 1959 3829 2000 3885
rect 2055 3829 2082 3885
rect -2506 3792 -2420 3801
rect -4189 3655 -4066 3749
rect -2580 3736 -2495 3792
rect -2439 3736 -2420 3792
rect -2506 3733 -2420 3736
rect 1959 3735 2082 3829
rect -4189 3599 -4162 3655
rect -4107 3599 -4066 3655
rect -2780 3609 -2240 3668
rect -4189 3505 -4066 3599
rect -1299 3642 -759 3701
rect 93 3648 633 3707
rect 1959 3679 2000 3735
rect 2055 3679 2082 3735
rect -4189 3449 -4162 3505
rect -4107 3449 -4066 3505
rect -4189 3355 -4066 3449
rect -4189 3299 -4162 3355
rect -4107 3299 -4066 3355
rect 1959 3585 2082 3679
rect 1959 3529 2000 3585
rect 2055 3529 2082 3585
rect 1959 3435 2082 3529
rect 1959 3379 2000 3435
rect 2055 3379 2082 3435
rect -1224 3325 -1116 3335
rect 489 3333 574 3346
rect 489 3332 709 3333
rect -4189 3205 -4066 3299
rect -1323 3324 -827 3325
rect -4189 3149 -4162 3205
rect -4107 3149 -4066 3205
rect -3721 3187 -3618 3233
rect -2652 3224 -2233 3270
rect -1323 3254 -1209 3324
rect -1139 3254 -827 3324
rect 489 3262 502 3332
rect 572 3262 709 3332
rect 1959 3285 2082 3379
rect 489 3261 709 3262
rect 489 3259 574 3261
rect -1323 3253 -827 3254
rect -1224 3241 -1116 3253
rect 1588 3232 1858 3278
rect 1959 3229 2000 3285
rect 2055 3229 2082 3285
rect -4189 3055 -4066 3149
rect -4189 2999 -4162 3055
rect -4107 2999 -4066 3055
rect -4189 2905 -4066 2999
rect -4189 2849 -4162 2905
rect -4107 2849 -4066 2905
rect -4189 2755 -4066 2849
rect 1959 3135 2082 3229
rect 1959 3079 2000 3135
rect 2055 3079 2082 3135
rect 1959 2985 2082 3079
rect 1959 2929 2000 2985
rect 2055 2929 2082 2985
rect 1959 2835 2082 2929
rect 1959 2779 2000 2835
rect 2055 2779 2082 2835
rect -4189 2699 -4162 2755
rect -4107 2699 -4066 2755
rect -1144 2732 -1068 2748
rect -4189 2605 -4066 2699
rect -4189 2549 -4162 2605
rect -4107 2549 -4066 2605
rect -4189 2455 -4066 2549
rect -4189 2399 -4162 2455
rect -4107 2399 -4066 2455
rect -4189 2305 -4066 2399
rect -4189 2249 -4162 2305
rect -4107 2249 -4066 2305
rect -4189 2155 -4066 2249
rect -4189 2099 -4162 2155
rect -4107 2099 -4066 2155
rect -4189 2005 -4066 2099
rect -4189 1949 -4162 2005
rect -4107 1949 -4066 2005
rect -4189 1855 -4066 1949
rect -4189 1799 -4162 1855
rect -4107 1799 -4066 1855
rect -4189 1705 -4066 1799
rect -4189 1649 -4162 1705
rect -4107 1649 -4066 1705
rect -4189 1555 -4066 1649
rect -4189 1499 -4162 1555
rect -4107 1499 -4066 1555
rect -4189 1405 -4066 1499
rect -4189 1349 -4162 1405
rect -4107 1349 -4066 1405
rect -4189 1255 -4066 1349
rect -4189 1199 -4162 1255
rect -4107 1199 -4066 1255
rect -4189 1105 -4066 1199
rect -4189 1049 -4162 1105
rect -4107 1049 -4066 1105
rect -3945 1880 -3848 2722
rect -2363 2643 -2264 2674
rect -1144 2669 -1135 2732
rect -1072 2669 -1068 2732
rect -1144 2658 -1068 2669
rect -738 2730 -652 2744
rect -738 2673 -725 2730
rect -663 2673 -652 2730
rect -738 2659 -652 2673
rect -2363 2587 -2340 2643
rect -2281 2587 -2264 2643
rect -2363 2560 -2264 2587
rect -2666 2389 -2358 2444
rect -2413 2176 -2358 2389
rect -2413 2163 -2314 2176
rect -3765 2088 -3583 2113
rect -2413 2109 -2378 2163
rect -2324 2109 -2314 2163
rect -2413 2108 -2314 2109
rect -2380 2097 -2314 2108
rect -3765 2032 -3736 2088
rect -3677 2032 -3583 2088
rect -3765 2011 -3583 2032
rect -2509 2015 -2424 2029
rect -2509 1961 -2494 2015
rect -2440 1961 -2424 2015
rect -2509 1958 -2424 1961
rect -3723 1885 -2663 1906
rect -3945 1822 -3925 1880
rect -3868 1822 -3848 1880
rect -3945 1167 -3848 1822
rect -2495 1407 -2440 1958
rect -1134 1932 -1071 2658
rect -2327 1880 -2250 1909
rect -1293 1887 -1071 1932
rect -817 1943 -712 1945
rect -817 1910 -367 1943
rect -308 1910 243 1943
rect -817 1905 243 1910
rect 324 1911 421 2761
rect 1959 2685 2082 2779
rect 1959 2629 2000 2685
rect 2055 2629 2082 2685
rect 1959 2535 2082 2629
rect 1959 2479 2000 2535
rect 2055 2479 2082 2535
rect 1959 2385 2082 2479
rect 1959 2329 2000 2385
rect 2055 2329 2082 2385
rect 1959 2235 2082 2329
rect 1959 2179 2000 2235
rect 2055 2179 2082 2235
rect 1959 2085 2082 2179
rect 1959 2029 2000 2085
rect 2055 2029 2082 2085
rect 1753 1964 1854 1968
rect 1753 1940 1765 1964
rect -1293 1886 -1087 1887
rect -2327 1822 -2320 1880
rect -2262 1822 -2250 1880
rect -2327 1807 -2250 1822
rect -2666 1352 -2440 1407
rect -3945 1070 -3753 1167
rect -4189 955 -4066 1049
rect -1133 1033 -1087 1886
rect 324 1839 688 1911
rect 1600 1894 1765 1940
rect 1743 1892 1765 1894
rect 1837 1892 1854 1964
rect 1743 1879 1854 1892
rect 1959 1935 2082 2029
rect 1959 1879 2000 1935
rect 2055 1879 2082 1935
rect -908 1437 -833 1449
rect -908 1372 -907 1437
rect -842 1372 -833 1437
rect -908 1359 -833 1372
rect 324 1188 421 1839
rect 273 1091 421 1188
rect 1743 1067 1815 1879
rect -4189 899 -4162 955
rect -4107 899 -4066 955
rect -4189 805 -4066 899
rect -4189 749 -4162 805
rect -4107 749 -4066 805
rect -4189 655 -4066 749
rect -4189 599 -4162 655
rect -4107 599 -4066 655
rect -2465 958 -2263 1004
rect -1283 987 -1087 1033
rect 563 1007 615 1018
rect 361 961 615 1007
rect 1570 995 1815 1067
rect 1959 1785 2082 1879
rect 1959 1729 2000 1785
rect 2055 1729 2082 1785
rect 1959 1635 2082 1729
rect 1959 1579 2000 1635
rect 2055 1579 2082 1635
rect 1959 1485 2082 1579
rect 1959 1429 2000 1485
rect 2055 1429 2082 1485
rect 1959 1335 2082 1429
rect 1959 1279 2000 1335
rect 2055 1279 2082 1335
rect 1959 1185 2082 1279
rect 1959 1129 2000 1185
rect 2055 1129 2082 1185
rect 1959 1035 2082 1129
rect -4189 505 -4066 599
rect -4189 449 -4162 505
rect -4107 449 -4066 505
rect -4189 355 -4066 449
rect -4189 299 -4162 355
rect -4107 299 -4066 355
rect -4189 205 -4066 299
rect -4189 149 -4162 205
rect -4107 149 -4066 205
rect -4189 55 -4066 149
rect -4189 -1 -4162 55
rect -4107 -1 -4066 55
rect -4189 -99 -4066 -1
rect -3722 559 -3618 605
rect -3722 35 -3676 559
rect -2465 35 -2419 958
rect 361 626 407 961
rect 563 957 615 961
rect 1959 979 2000 1035
rect 2055 979 2082 1035
rect 138 580 407 626
rect 1959 885 2082 979
rect 1959 829 2000 885
rect 2055 829 2082 885
rect 1959 735 2082 829
rect 1959 679 2000 735
rect 2055 679 2082 735
rect 1959 585 2082 679
rect 1959 529 2000 585
rect 2055 529 2082 585
rect 1959 435 2082 529
rect 1959 379 2000 435
rect 2055 379 2082 435
rect 1959 285 2082 379
rect 1959 229 2000 285
rect 2055 229 2082 285
rect -3722 -11 -2419 35
rect 1959 135 2082 229
rect 1959 79 2000 135
rect 2055 79 2082 135
rect 1959 -15 2082 79
rect 1959 -71 2000 -15
rect 2055 -71 2082 -15
rect 1959 -99 2082 -71
rect -4189 -131 2082 -99
rect -4189 -187 -4062 -131
rect -4007 -187 -3912 -131
rect -3857 -187 -3762 -131
rect -3707 -187 -3612 -131
rect -3557 -187 -3462 -131
rect -3407 -187 -3312 -131
rect -3257 -187 -3162 -131
rect -3107 -187 -3012 -131
rect -2957 -187 -2862 -131
rect -2807 -187 -2712 -131
rect -2657 -187 -2562 -131
rect -2507 -187 -2412 -131
rect -2357 -187 -2262 -131
rect -2207 -187 -2112 -131
rect -2057 -187 -1962 -131
rect -1907 -187 -1812 -131
rect -1757 -187 -1662 -131
rect -1607 -187 -1512 -131
rect -1457 -187 -1362 -131
rect -1307 -187 -1212 -131
rect -1157 -187 -1062 -131
rect -1007 -187 -912 -131
rect -857 -187 -762 -131
rect -707 -187 -612 -131
rect -557 -187 -462 -131
rect -407 -187 -312 -131
rect -257 -187 -162 -131
rect -107 -187 -12 -131
rect 43 -187 138 -131
rect 193 -187 288 -131
rect 343 -187 438 -131
rect 493 -187 588 -131
rect 643 -187 738 -131
rect 793 -187 888 -131
rect 943 -187 1038 -131
rect 1093 -187 1188 -131
rect 1243 -187 1338 -131
rect 1393 -187 1488 -131
rect 1543 -187 1638 -131
rect 1693 -187 1788 -131
rect 1843 -187 1938 -131
rect 1993 -187 2082 -131
rect -4189 -221 2082 -187
rect -3706 -222 2082 -221
<< via1 >>
rect -2495 3736 -2439 3792
rect -2895 3617 -2836 3673
rect -2046 3593 -1987 3649
rect 874 3599 933 3655
rect -1209 3254 -1139 3324
rect 502 3262 572 3332
rect -1135 2669 -1072 2732
rect -725 2673 -663 2730
rect -2340 2587 -2281 2643
rect -1461 2575 -1402 2631
rect -2378 2109 -2324 2163
rect -3736 2032 -3677 2088
rect -2494 1961 -2440 2015
rect -3925 1822 -3868 1880
rect -367 1910 -308 1966
rect 628 2462 687 2518
rect -2320 1822 -2262 1880
rect -1979 1435 -1920 1491
rect 1765 1892 1837 1964
rect -907 1372 -842 1437
rect 918 1433 977 1489
rect -2891 116 -2832 172
rect -1441 345 -1382 401
rect 678 346 737 402
rect -674 150 -615 206
<< metal2 >>
rect -2506 3792 -1138 3801
rect -2506 3736 -2495 3792
rect -2439 3745 -1138 3792
rect -2439 3736 -2420 3745
rect -2506 3733 -2420 3736
rect -2907 3675 -2822 3685
rect -2907 3615 -2897 3675
rect -2834 3615 -2822 3675
rect -2907 3603 -2822 3615
rect -3757 2090 -3649 2109
rect -3757 2030 -3738 2090
rect -3675 2030 -3649 2090
rect -3757 2016 -3649 2030
rect -2495 2029 -2439 3733
rect -2058 3651 -1973 3661
rect -2058 3591 -2048 3651
rect -1985 3591 -1973 3651
rect -2058 3579 -1973 3591
rect -1210 3335 -1138 3745
rect 862 3657 947 3667
rect 862 3597 872 3657
rect 935 3597 947 3657
rect 862 3585 947 3597
rect -1224 3324 -1116 3335
rect -1224 3254 -1209 3324
rect -1139 3254 -1116 3324
rect 489 3332 574 3346
rect 489 3262 502 3332
rect 572 3262 574 3332
rect 489 3259 574 3262
rect -1224 3241 -1116 3254
rect -1144 2732 -1068 2748
rect -738 2732 -652 2744
rect -2363 2645 -2264 2674
rect -1144 2669 -1135 2732
rect -1072 2730 -652 2732
rect -1072 2673 -725 2730
rect -663 2673 -652 2730
rect -1072 2669 -652 2673
rect -1144 2658 -1068 2669
rect -738 2659 -652 2669
rect 501 2658 573 3259
rect -2363 2585 -2342 2645
rect -2279 2585 -2264 2645
rect -2363 2560 -2264 2585
rect -1473 2633 -1388 2643
rect -1473 2573 -1463 2633
rect -1400 2573 -1388 2633
rect 501 2586 1837 2658
rect -1473 2561 -1388 2573
rect 616 2520 701 2530
rect 616 2460 626 2520
rect 689 2460 701 2520
rect 616 2448 701 2460
rect -2380 2167 -2314 2176
rect -2380 2163 -939 2167
rect -2380 2109 -2378 2163
rect -2324 2109 -939 2163
rect -2380 2102 -939 2109
rect -2380 2097 -2314 2102
rect -2509 2015 -2424 2029
rect -2509 1961 -2494 2015
rect -2440 1961 -2424 2015
rect -2509 1958 -2424 1961
rect -3941 1880 -3865 1892
rect -2327 1880 -2250 1909
rect -3941 1822 -3925 1880
rect -3868 1822 -2320 1880
rect -2262 1822 -2250 1880
rect -3941 1811 -3865 1822
rect -2327 1807 -2250 1822
rect -1991 1493 -1906 1503
rect -1991 1433 -1981 1493
rect -1918 1433 -1906 1493
rect -1991 1421 -1906 1433
rect -1004 1449 -939 2102
rect -379 1968 -294 1978
rect 1765 1968 1837 2586
rect -379 1908 -369 1968
rect -306 1908 -294 1968
rect -379 1896 -294 1908
rect 1753 1964 1854 1968
rect 1753 1892 1765 1964
rect 1837 1892 1854 1964
rect 1753 1879 1854 1892
rect 906 1491 991 1501
rect -1004 1437 -833 1449
rect -1004 1372 -907 1437
rect -842 1372 -833 1437
rect 906 1431 916 1491
rect 979 1431 991 1491
rect 906 1419 991 1431
rect -912 1359 -833 1372
rect -1453 403 -1368 413
rect -1453 343 -1443 403
rect -1380 343 -1368 403
rect -1453 331 -1368 343
rect 666 404 751 414
rect 666 344 676 404
rect 739 344 751 404
rect 666 332 751 344
rect -686 208 -601 218
rect -2903 174 -2818 184
rect -2903 114 -2893 174
rect -2830 114 -2818 174
rect -686 148 -676 208
rect -613 148 -601 208
rect -686 136 -601 148
rect -2903 102 -2818 114
<< via2 >>
rect -2897 3673 -2834 3675
rect -2897 3617 -2895 3673
rect -2895 3617 -2836 3673
rect -2836 3617 -2834 3673
rect -2897 3615 -2834 3617
rect -3738 2088 -3675 2090
rect -3738 2032 -3736 2088
rect -3736 2032 -3677 2088
rect -3677 2032 -3675 2088
rect -3738 2030 -3675 2032
rect -2048 3649 -1985 3651
rect -2048 3593 -2046 3649
rect -2046 3593 -1987 3649
rect -1987 3593 -1985 3649
rect -2048 3591 -1985 3593
rect 872 3655 935 3657
rect 872 3599 874 3655
rect 874 3599 933 3655
rect 933 3599 935 3655
rect 872 3597 935 3599
rect -2342 2643 -2279 2645
rect -2342 2587 -2340 2643
rect -2340 2587 -2281 2643
rect -2281 2587 -2279 2643
rect -2342 2585 -2279 2587
rect -1463 2631 -1400 2633
rect -1463 2575 -1461 2631
rect -1461 2575 -1402 2631
rect -1402 2575 -1400 2631
rect -1463 2573 -1400 2575
rect 626 2518 689 2520
rect 626 2462 628 2518
rect 628 2462 687 2518
rect 687 2462 689 2518
rect 626 2460 689 2462
rect -1981 1491 -1918 1493
rect -1981 1435 -1979 1491
rect -1979 1435 -1920 1491
rect -1920 1435 -1918 1491
rect -1981 1433 -1918 1435
rect -369 1966 -306 1968
rect -369 1910 -367 1966
rect -367 1910 -308 1966
rect -308 1910 -306 1966
rect -369 1908 -306 1910
rect 916 1489 979 1491
rect 916 1433 918 1489
rect 918 1433 977 1489
rect 977 1433 979 1489
rect 916 1431 979 1433
rect -1443 401 -1380 403
rect -1443 345 -1441 401
rect -1441 345 -1382 401
rect -1382 345 -1380 401
rect -1443 343 -1380 345
rect 676 402 739 404
rect 676 346 678 402
rect 678 346 737 402
rect 737 346 739 402
rect 676 344 739 346
rect -2893 172 -2830 174
rect -2893 116 -2891 172
rect -2891 116 -2832 172
rect -2832 116 -2830 172
rect -2893 114 -2830 116
rect -676 206 -613 208
rect -676 150 -674 206
rect -674 150 -615 206
rect -615 150 -613 206
rect -676 148 -613 150
<< metal3 >>
rect -2907 3675 -2822 3685
rect -2907 3615 -2897 3675
rect -2834 3615 -2822 3675
rect 862 3665 947 3667
rect -2907 3603 -2822 3615
rect -2058 3651 -1973 3661
rect -2058 3591 -2048 3651
rect -1985 3634 -1973 3651
rect 862 3657 961 3665
rect -1985 3591 -1918 3634
rect -2058 3574 -1918 3591
rect 862 3597 872 3657
rect 935 3597 961 3657
rect 862 3585 961 3597
rect -2363 2646 -2264 2674
rect -3506 2645 -2264 2646
rect -3506 2585 -2342 2645
rect -2279 2585 -2264 2645
rect -3757 2090 -3649 2109
rect -3757 2030 -3738 2090
rect -3675 2086 -3649 2090
rect -3506 2086 -3445 2585
rect -2363 2560 -2264 2585
rect -3675 2030 -3444 2086
rect -3757 2025 -3444 2030
rect -3757 2016 -3649 2025
rect -3506 2020 -3445 2025
rect -1978 1503 -1918 3574
rect -1473 2633 -1388 2643
rect -1473 2606 -1463 2633
rect -1477 2573 -1463 2606
rect -1400 2573 -1388 2633
rect -1477 2561 -1388 2573
rect -1477 1982 -1414 2561
rect 616 2520 701 2530
rect 616 2460 626 2520
rect 689 2460 701 2520
rect 616 2448 701 2460
rect 624 1982 687 2448
rect -1477 1968 687 1982
rect -1477 1919 -369 1968
rect -1991 1493 -1906 1503
rect -1991 1433 -1981 1493
rect -1918 1433 -1906 1493
rect -1991 1421 -1906 1433
rect -2903 174 -2818 184
rect -2903 114 -2893 174
rect -2830 173 -2818 174
rect -1978 173 -1918 1421
rect -1477 413 -1414 1919
rect -379 1908 -369 1919
rect -306 1919 687 1968
rect -306 1908 -294 1919
rect -379 1896 -294 1908
rect 624 414 687 1919
rect 901 1501 961 3585
rect 901 1491 991 1501
rect 901 1431 916 1491
rect 979 1431 991 1491
rect 901 1419 991 1431
rect -1477 403 -1368 413
rect -1477 343 -1443 403
rect -1380 343 -1368 403
rect -1477 337 -1368 343
rect -1453 331 -1368 337
rect 624 404 751 414
rect 624 344 676 404
rect 739 344 751 404
rect 624 332 751 344
rect -686 208 -601 218
rect -686 173 -676 208
rect -2830 148 -676 173
rect -613 173 -601 208
rect 901 173 961 1419
rect -613 148 961 173
rect -2830 114 961 148
rect -2903 113 961 114
rect -2903 102 -2818 113
use INV_2  INV_2_0
timestamp 1692626060
transform -1 0 -1216 0 -1 3226
box 21 -485 1081 648
use INV_2  INV_2_1
timestamp 1692626060
transform 1 0 -2318 0 1 1930
box 21 -485 1081 648
use INV_2  INV_2_2
timestamp 1692626060
transform 1 0 575 0 -1 3234
box 21 -485 1081 648
use INV_2  INV_2_3
timestamp 1692626060
transform 1 0 575 0 1 1938
box 21 -485 1081 648
use INV_2  INV_2_4
timestamp 1692626060
transform -1 0 1677 0 -1 968
box 21 -485 1081 648
use INV_2  INV_2_5
timestamp 1692626060
transform -1 0 -1216 0 -1 960
box 21 -485 1081 648
use Tr_Gate  Tr_Gate_0 ~/GF180Projects/Layout/Magic/VCO1/Tr_Gate
timestamp 1691796835
transform 1 0 -817 0 1 1343
box -53 -1233 1187 569
use Tr_Gate  Tr_Gate_1
timestamp 1691796835
transform 1 0 -817 0 -1 2509
box -53 -1233 1187 569
use Tr_Gate  Tr_Gate_2
timestamp 1691796835
transform -1 0 -2663 0 -1 2470
box -53 -1233 1187 569
use Tr_Gate  Tr_Gate_3
timestamp 1691796835
transform -1 0 -2663 0 1 1322
box -53 -1233 1187 569
<< labels >>
flabel metal1 -3700 3207 -3699 3208 0 FreeSans 800 0 0 0 D
port 0 nsew
flabel via1 1813 1916 1813 1916 0 FreeSans 800 0 0 0 Q
port 2 nsew
flabel metal1 1835 3254 1835 3254 0 FreeSans 800 0 0 0 Q-
port 3 nsew
flabel metal1 324 3679 324 3679 0 FreeSans 800 0 0 0 VSS
port 4 nsew
flabel metal1 -3762 2064 -3762 2064 0 FreeSans 800 0 0 0 VDD
port 5 nsew
flabel metal1 -2550 3766 -2550 3766 0 FreeSans 800 0 0 0 CLK
port 1 nsew
<< end >>
