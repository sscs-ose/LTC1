magic
tech gf180mcuD
magscale 1 5
timestamp 1713185578
<< checkpaint >>
rect -19705 -19480 19705 19480
<< mimcap >>
rect -18645 18284 -15545 18390
rect -18645 15596 -18553 18284
rect -15637 15596 -15545 18284
rect -18645 15490 -15545 15596
rect -15238 18284 -12138 18390
rect -15238 15596 -15146 18284
rect -12230 15596 -12138 18284
rect -15238 15490 -12138 15596
rect -11831 18284 -8731 18390
rect -11831 15596 -11739 18284
rect -8823 15596 -8731 18284
rect -11831 15490 -8731 15596
rect -8424 18284 -5324 18390
rect -8424 15596 -8332 18284
rect -5416 15596 -5324 18284
rect -8424 15490 -5324 15596
rect -5017 18284 -1917 18390
rect -5017 15596 -4925 18284
rect -2009 15596 -1917 18284
rect -5017 15490 -1917 15596
rect -1610 18284 1490 18390
rect -1610 15596 -1518 18284
rect 1398 15596 1490 18284
rect -1610 15490 1490 15596
rect 1797 18284 4897 18390
rect 1797 15596 1889 18284
rect 4805 15596 4897 18284
rect 1797 15490 4897 15596
rect 5204 18284 8304 18390
rect 5204 15596 5296 18284
rect 8212 15596 8304 18284
rect 5204 15490 8304 15596
rect 8611 18284 11711 18390
rect 8611 15596 8703 18284
rect 11619 15596 11711 18284
rect 8611 15490 11711 15596
rect 12018 18284 15118 18390
rect 12018 15596 12110 18284
rect 15026 15596 15118 18284
rect 12018 15490 15118 15596
rect 15425 18284 18525 18390
rect 15425 15596 15517 18284
rect 18433 15596 18525 18284
rect 15425 15490 18525 15596
rect -18645 15204 -15545 15310
rect -18645 12516 -18553 15204
rect -15637 12516 -15545 15204
rect -18645 12410 -15545 12516
rect -15238 15204 -12138 15310
rect -15238 12516 -15146 15204
rect -12230 12516 -12138 15204
rect -15238 12410 -12138 12516
rect -11831 15204 -8731 15310
rect -11831 12516 -11739 15204
rect -8823 12516 -8731 15204
rect -11831 12410 -8731 12516
rect -8424 15204 -5324 15310
rect -8424 12516 -8332 15204
rect -5416 12516 -5324 15204
rect -8424 12410 -5324 12516
rect -5017 15204 -1917 15310
rect -5017 12516 -4925 15204
rect -2009 12516 -1917 15204
rect -5017 12410 -1917 12516
rect -1610 15204 1490 15310
rect -1610 12516 -1518 15204
rect 1398 12516 1490 15204
rect -1610 12410 1490 12516
rect 1797 15204 4897 15310
rect 1797 12516 1889 15204
rect 4805 12516 4897 15204
rect 1797 12410 4897 12516
rect 5204 15204 8304 15310
rect 5204 12516 5296 15204
rect 8212 12516 8304 15204
rect 5204 12410 8304 12516
rect 8611 15204 11711 15310
rect 8611 12516 8703 15204
rect 11619 12516 11711 15204
rect 8611 12410 11711 12516
rect 12018 15204 15118 15310
rect 12018 12516 12110 15204
rect 15026 12516 15118 15204
rect 12018 12410 15118 12516
rect 15425 15204 18525 15310
rect 15425 12516 15517 15204
rect 18433 12516 18525 15204
rect 15425 12410 18525 12516
rect -18645 12124 -15545 12230
rect -18645 9436 -18553 12124
rect -15637 9436 -15545 12124
rect -18645 9330 -15545 9436
rect -15238 12124 -12138 12230
rect -15238 9436 -15146 12124
rect -12230 9436 -12138 12124
rect -15238 9330 -12138 9436
rect -11831 12124 -8731 12230
rect -11831 9436 -11739 12124
rect -8823 9436 -8731 12124
rect -11831 9330 -8731 9436
rect -8424 12124 -5324 12230
rect -8424 9436 -8332 12124
rect -5416 9436 -5324 12124
rect -8424 9330 -5324 9436
rect -5017 12124 -1917 12230
rect -5017 9436 -4925 12124
rect -2009 9436 -1917 12124
rect -5017 9330 -1917 9436
rect -1610 12124 1490 12230
rect -1610 9436 -1518 12124
rect 1398 9436 1490 12124
rect -1610 9330 1490 9436
rect 1797 12124 4897 12230
rect 1797 9436 1889 12124
rect 4805 9436 4897 12124
rect 1797 9330 4897 9436
rect 5204 12124 8304 12230
rect 5204 9436 5296 12124
rect 8212 9436 8304 12124
rect 5204 9330 8304 9436
rect 8611 12124 11711 12230
rect 8611 9436 8703 12124
rect 11619 9436 11711 12124
rect 8611 9330 11711 9436
rect 12018 12124 15118 12230
rect 12018 9436 12110 12124
rect 15026 9436 15118 12124
rect 12018 9330 15118 9436
rect 15425 12124 18525 12230
rect 15425 9436 15517 12124
rect 18433 9436 18525 12124
rect 15425 9330 18525 9436
rect -18645 9044 -15545 9150
rect -18645 6356 -18553 9044
rect -15637 6356 -15545 9044
rect -18645 6250 -15545 6356
rect -15238 9044 -12138 9150
rect -15238 6356 -15146 9044
rect -12230 6356 -12138 9044
rect -15238 6250 -12138 6356
rect -11831 9044 -8731 9150
rect -11831 6356 -11739 9044
rect -8823 6356 -8731 9044
rect -11831 6250 -8731 6356
rect -8424 9044 -5324 9150
rect -8424 6356 -8332 9044
rect -5416 6356 -5324 9044
rect -8424 6250 -5324 6356
rect -5017 9044 -1917 9150
rect -5017 6356 -4925 9044
rect -2009 6356 -1917 9044
rect -5017 6250 -1917 6356
rect -1610 9044 1490 9150
rect -1610 6356 -1518 9044
rect 1398 6356 1490 9044
rect -1610 6250 1490 6356
rect 1797 9044 4897 9150
rect 1797 6356 1889 9044
rect 4805 6356 4897 9044
rect 1797 6250 4897 6356
rect 5204 9044 8304 9150
rect 5204 6356 5296 9044
rect 8212 6356 8304 9044
rect 5204 6250 8304 6356
rect 8611 9044 11711 9150
rect 8611 6356 8703 9044
rect 11619 6356 11711 9044
rect 8611 6250 11711 6356
rect 12018 9044 15118 9150
rect 12018 6356 12110 9044
rect 15026 6356 15118 9044
rect 12018 6250 15118 6356
rect 15425 9044 18525 9150
rect 15425 6356 15517 9044
rect 18433 6356 18525 9044
rect 15425 6250 18525 6356
rect -18645 5964 -15545 6070
rect -18645 3276 -18553 5964
rect -15637 3276 -15545 5964
rect -18645 3170 -15545 3276
rect -15238 5964 -12138 6070
rect -15238 3276 -15146 5964
rect -12230 3276 -12138 5964
rect -15238 3170 -12138 3276
rect -11831 5964 -8731 6070
rect -11831 3276 -11739 5964
rect -8823 3276 -8731 5964
rect -11831 3170 -8731 3276
rect -8424 5964 -5324 6070
rect -8424 3276 -8332 5964
rect -5416 3276 -5324 5964
rect -8424 3170 -5324 3276
rect -5017 5964 -1917 6070
rect -5017 3276 -4925 5964
rect -2009 3276 -1917 5964
rect -5017 3170 -1917 3276
rect -1610 5964 1490 6070
rect -1610 3276 -1518 5964
rect 1398 3276 1490 5964
rect -1610 3170 1490 3276
rect 1797 5964 4897 6070
rect 1797 3276 1889 5964
rect 4805 3276 4897 5964
rect 1797 3170 4897 3276
rect 5204 5964 8304 6070
rect 5204 3276 5296 5964
rect 8212 3276 8304 5964
rect 5204 3170 8304 3276
rect 8611 5964 11711 6070
rect 8611 3276 8703 5964
rect 11619 3276 11711 5964
rect 8611 3170 11711 3276
rect 12018 5964 15118 6070
rect 12018 3276 12110 5964
rect 15026 3276 15118 5964
rect 12018 3170 15118 3276
rect 15425 5964 18525 6070
rect 15425 3276 15517 5964
rect 18433 3276 18525 5964
rect 15425 3170 18525 3276
rect -18645 2884 -15545 2990
rect -18645 196 -18553 2884
rect -15637 196 -15545 2884
rect -18645 90 -15545 196
rect -15238 2884 -12138 2990
rect -15238 196 -15146 2884
rect -12230 196 -12138 2884
rect -15238 90 -12138 196
rect -11831 2884 -8731 2990
rect -11831 196 -11739 2884
rect -8823 196 -8731 2884
rect -11831 90 -8731 196
rect -8424 2884 -5324 2990
rect -8424 196 -8332 2884
rect -5416 196 -5324 2884
rect -8424 90 -5324 196
rect -5017 2884 -1917 2990
rect -5017 196 -4925 2884
rect -2009 196 -1917 2884
rect -5017 90 -1917 196
rect -1610 2884 1490 2990
rect -1610 196 -1518 2884
rect 1398 196 1490 2884
rect -1610 90 1490 196
rect 1797 2884 4897 2990
rect 1797 196 1889 2884
rect 4805 196 4897 2884
rect 1797 90 4897 196
rect 5204 2884 8304 2990
rect 5204 196 5296 2884
rect 8212 196 8304 2884
rect 5204 90 8304 196
rect 8611 2884 11711 2990
rect 8611 196 8703 2884
rect 11619 196 11711 2884
rect 8611 90 11711 196
rect 12018 2884 15118 2990
rect 12018 196 12110 2884
rect 15026 196 15118 2884
rect 12018 90 15118 196
rect 15425 2884 18525 2990
rect 15425 196 15517 2884
rect 18433 196 18525 2884
rect 15425 90 18525 196
rect -18645 -196 -15545 -90
rect -18645 -2884 -18553 -196
rect -15637 -2884 -15545 -196
rect -18645 -2990 -15545 -2884
rect -15238 -196 -12138 -90
rect -15238 -2884 -15146 -196
rect -12230 -2884 -12138 -196
rect -15238 -2990 -12138 -2884
rect -11831 -196 -8731 -90
rect -11831 -2884 -11739 -196
rect -8823 -2884 -8731 -196
rect -11831 -2990 -8731 -2884
rect -8424 -196 -5324 -90
rect -8424 -2884 -8332 -196
rect -5416 -2884 -5324 -196
rect -8424 -2990 -5324 -2884
rect -5017 -196 -1917 -90
rect -5017 -2884 -4925 -196
rect -2009 -2884 -1917 -196
rect -5017 -2990 -1917 -2884
rect -1610 -196 1490 -90
rect -1610 -2884 -1518 -196
rect 1398 -2884 1490 -196
rect -1610 -2990 1490 -2884
rect 1797 -196 4897 -90
rect 1797 -2884 1889 -196
rect 4805 -2884 4897 -196
rect 1797 -2990 4897 -2884
rect 5204 -196 8304 -90
rect 5204 -2884 5296 -196
rect 8212 -2884 8304 -196
rect 5204 -2990 8304 -2884
rect 8611 -196 11711 -90
rect 8611 -2884 8703 -196
rect 11619 -2884 11711 -196
rect 8611 -2990 11711 -2884
rect 12018 -196 15118 -90
rect 12018 -2884 12110 -196
rect 15026 -2884 15118 -196
rect 12018 -2990 15118 -2884
rect 15425 -196 18525 -90
rect 15425 -2884 15517 -196
rect 18433 -2884 18525 -196
rect 15425 -2990 18525 -2884
rect -18645 -3276 -15545 -3170
rect -18645 -5964 -18553 -3276
rect -15637 -5964 -15545 -3276
rect -18645 -6070 -15545 -5964
rect -15238 -3276 -12138 -3170
rect -15238 -5964 -15146 -3276
rect -12230 -5964 -12138 -3276
rect -15238 -6070 -12138 -5964
rect -11831 -3276 -8731 -3170
rect -11831 -5964 -11739 -3276
rect -8823 -5964 -8731 -3276
rect -11831 -6070 -8731 -5964
rect -8424 -3276 -5324 -3170
rect -8424 -5964 -8332 -3276
rect -5416 -5964 -5324 -3276
rect -8424 -6070 -5324 -5964
rect -5017 -3276 -1917 -3170
rect -5017 -5964 -4925 -3276
rect -2009 -5964 -1917 -3276
rect -5017 -6070 -1917 -5964
rect -1610 -3276 1490 -3170
rect -1610 -5964 -1518 -3276
rect 1398 -5964 1490 -3276
rect -1610 -6070 1490 -5964
rect 1797 -3276 4897 -3170
rect 1797 -5964 1889 -3276
rect 4805 -5964 4897 -3276
rect 1797 -6070 4897 -5964
rect 5204 -3276 8304 -3170
rect 5204 -5964 5296 -3276
rect 8212 -5964 8304 -3276
rect 5204 -6070 8304 -5964
rect 8611 -3276 11711 -3170
rect 8611 -5964 8703 -3276
rect 11619 -5964 11711 -3276
rect 8611 -6070 11711 -5964
rect 12018 -3276 15118 -3170
rect 12018 -5964 12110 -3276
rect 15026 -5964 15118 -3276
rect 12018 -6070 15118 -5964
rect 15425 -3276 18525 -3170
rect 15425 -5964 15517 -3276
rect 18433 -5964 18525 -3276
rect 15425 -6070 18525 -5964
rect -18645 -6356 -15545 -6250
rect -18645 -9044 -18553 -6356
rect -15637 -9044 -15545 -6356
rect -18645 -9150 -15545 -9044
rect -15238 -6356 -12138 -6250
rect -15238 -9044 -15146 -6356
rect -12230 -9044 -12138 -6356
rect -15238 -9150 -12138 -9044
rect -11831 -6356 -8731 -6250
rect -11831 -9044 -11739 -6356
rect -8823 -9044 -8731 -6356
rect -11831 -9150 -8731 -9044
rect -8424 -6356 -5324 -6250
rect -8424 -9044 -8332 -6356
rect -5416 -9044 -5324 -6356
rect -8424 -9150 -5324 -9044
rect -5017 -6356 -1917 -6250
rect -5017 -9044 -4925 -6356
rect -2009 -9044 -1917 -6356
rect -5017 -9150 -1917 -9044
rect -1610 -6356 1490 -6250
rect -1610 -9044 -1518 -6356
rect 1398 -9044 1490 -6356
rect -1610 -9150 1490 -9044
rect 1797 -6356 4897 -6250
rect 1797 -9044 1889 -6356
rect 4805 -9044 4897 -6356
rect 1797 -9150 4897 -9044
rect 5204 -6356 8304 -6250
rect 5204 -9044 5296 -6356
rect 8212 -9044 8304 -6356
rect 5204 -9150 8304 -9044
rect 8611 -6356 11711 -6250
rect 8611 -9044 8703 -6356
rect 11619 -9044 11711 -6356
rect 8611 -9150 11711 -9044
rect 12018 -6356 15118 -6250
rect 12018 -9044 12110 -6356
rect 15026 -9044 15118 -6356
rect 12018 -9150 15118 -9044
rect 15425 -6356 18525 -6250
rect 15425 -9044 15517 -6356
rect 18433 -9044 18525 -6356
rect 15425 -9150 18525 -9044
rect -18645 -9436 -15545 -9330
rect -18645 -12124 -18553 -9436
rect -15637 -12124 -15545 -9436
rect -18645 -12230 -15545 -12124
rect -15238 -9436 -12138 -9330
rect -15238 -12124 -15146 -9436
rect -12230 -12124 -12138 -9436
rect -15238 -12230 -12138 -12124
rect -11831 -9436 -8731 -9330
rect -11831 -12124 -11739 -9436
rect -8823 -12124 -8731 -9436
rect -11831 -12230 -8731 -12124
rect -8424 -9436 -5324 -9330
rect -8424 -12124 -8332 -9436
rect -5416 -12124 -5324 -9436
rect -8424 -12230 -5324 -12124
rect -5017 -9436 -1917 -9330
rect -5017 -12124 -4925 -9436
rect -2009 -12124 -1917 -9436
rect -5017 -12230 -1917 -12124
rect -1610 -9436 1490 -9330
rect -1610 -12124 -1518 -9436
rect 1398 -12124 1490 -9436
rect -1610 -12230 1490 -12124
rect 1797 -9436 4897 -9330
rect 1797 -12124 1889 -9436
rect 4805 -12124 4897 -9436
rect 1797 -12230 4897 -12124
rect 5204 -9436 8304 -9330
rect 5204 -12124 5296 -9436
rect 8212 -12124 8304 -9436
rect 5204 -12230 8304 -12124
rect 8611 -9436 11711 -9330
rect 8611 -12124 8703 -9436
rect 11619 -12124 11711 -9436
rect 8611 -12230 11711 -12124
rect 12018 -9436 15118 -9330
rect 12018 -12124 12110 -9436
rect 15026 -12124 15118 -9436
rect 12018 -12230 15118 -12124
rect 15425 -9436 18525 -9330
rect 15425 -12124 15517 -9436
rect 18433 -12124 18525 -9436
rect 15425 -12230 18525 -12124
rect -18645 -12516 -15545 -12410
rect -18645 -15204 -18553 -12516
rect -15637 -15204 -15545 -12516
rect -18645 -15310 -15545 -15204
rect -15238 -12516 -12138 -12410
rect -15238 -15204 -15146 -12516
rect -12230 -15204 -12138 -12516
rect -15238 -15310 -12138 -15204
rect -11831 -12516 -8731 -12410
rect -11831 -15204 -11739 -12516
rect -8823 -15204 -8731 -12516
rect -11831 -15310 -8731 -15204
rect -8424 -12516 -5324 -12410
rect -8424 -15204 -8332 -12516
rect -5416 -15204 -5324 -12516
rect -8424 -15310 -5324 -15204
rect -5017 -12516 -1917 -12410
rect -5017 -15204 -4925 -12516
rect -2009 -15204 -1917 -12516
rect -5017 -15310 -1917 -15204
rect -1610 -12516 1490 -12410
rect -1610 -15204 -1518 -12516
rect 1398 -15204 1490 -12516
rect -1610 -15310 1490 -15204
rect 1797 -12516 4897 -12410
rect 1797 -15204 1889 -12516
rect 4805 -15204 4897 -12516
rect 1797 -15310 4897 -15204
rect 5204 -12516 8304 -12410
rect 5204 -15204 5296 -12516
rect 8212 -15204 8304 -12516
rect 5204 -15310 8304 -15204
rect 8611 -12516 11711 -12410
rect 8611 -15204 8703 -12516
rect 11619 -15204 11711 -12516
rect 8611 -15310 11711 -15204
rect 12018 -12516 15118 -12410
rect 12018 -15204 12110 -12516
rect 15026 -15204 15118 -12516
rect 12018 -15310 15118 -15204
rect 15425 -12516 18525 -12410
rect 15425 -15204 15517 -12516
rect 18433 -15204 18525 -12516
rect 15425 -15310 18525 -15204
rect -18645 -15596 -15545 -15490
rect -18645 -18284 -18553 -15596
rect -15637 -18284 -15545 -15596
rect -18645 -18390 -15545 -18284
rect -15238 -15596 -12138 -15490
rect -15238 -18284 -15146 -15596
rect -12230 -18284 -12138 -15596
rect -15238 -18390 -12138 -18284
rect -11831 -15596 -8731 -15490
rect -11831 -18284 -11739 -15596
rect -8823 -18284 -8731 -15596
rect -11831 -18390 -8731 -18284
rect -8424 -15596 -5324 -15490
rect -8424 -18284 -8332 -15596
rect -5416 -18284 -5324 -15596
rect -8424 -18390 -5324 -18284
rect -5017 -15596 -1917 -15490
rect -5017 -18284 -4925 -15596
rect -2009 -18284 -1917 -15596
rect -5017 -18390 -1917 -18284
rect -1610 -15596 1490 -15490
rect -1610 -18284 -1518 -15596
rect 1398 -18284 1490 -15596
rect -1610 -18390 1490 -18284
rect 1797 -15596 4897 -15490
rect 1797 -18284 1889 -15596
rect 4805 -18284 4897 -15596
rect 1797 -18390 4897 -18284
rect 5204 -15596 8304 -15490
rect 5204 -18284 5296 -15596
rect 8212 -18284 8304 -15596
rect 5204 -18390 8304 -18284
rect 8611 -15596 11711 -15490
rect 8611 -18284 8703 -15596
rect 11619 -18284 11711 -15596
rect 8611 -18390 11711 -18284
rect 12018 -15596 15118 -15490
rect 12018 -18284 12110 -15596
rect 15026 -18284 15118 -15596
rect 12018 -18390 15118 -18284
rect 15425 -15596 18525 -15490
rect 15425 -18284 15517 -15596
rect 18433 -18284 18525 -15596
rect 15425 -18390 18525 -18284
<< mimcapcontact >>
rect -18553 15596 -15637 18284
rect -15146 15596 -12230 18284
rect -11739 15596 -8823 18284
rect -8332 15596 -5416 18284
rect -4925 15596 -2009 18284
rect -1518 15596 1398 18284
rect 1889 15596 4805 18284
rect 5296 15596 8212 18284
rect 8703 15596 11619 18284
rect 12110 15596 15026 18284
rect 15517 15596 18433 18284
rect -18553 12516 -15637 15204
rect -15146 12516 -12230 15204
rect -11739 12516 -8823 15204
rect -8332 12516 -5416 15204
rect -4925 12516 -2009 15204
rect -1518 12516 1398 15204
rect 1889 12516 4805 15204
rect 5296 12516 8212 15204
rect 8703 12516 11619 15204
rect 12110 12516 15026 15204
rect 15517 12516 18433 15204
rect -18553 9436 -15637 12124
rect -15146 9436 -12230 12124
rect -11739 9436 -8823 12124
rect -8332 9436 -5416 12124
rect -4925 9436 -2009 12124
rect -1518 9436 1398 12124
rect 1889 9436 4805 12124
rect 5296 9436 8212 12124
rect 8703 9436 11619 12124
rect 12110 9436 15026 12124
rect 15517 9436 18433 12124
rect -18553 6356 -15637 9044
rect -15146 6356 -12230 9044
rect -11739 6356 -8823 9044
rect -8332 6356 -5416 9044
rect -4925 6356 -2009 9044
rect -1518 6356 1398 9044
rect 1889 6356 4805 9044
rect 5296 6356 8212 9044
rect 8703 6356 11619 9044
rect 12110 6356 15026 9044
rect 15517 6356 18433 9044
rect -18553 3276 -15637 5964
rect -15146 3276 -12230 5964
rect -11739 3276 -8823 5964
rect -8332 3276 -5416 5964
rect -4925 3276 -2009 5964
rect -1518 3276 1398 5964
rect 1889 3276 4805 5964
rect 5296 3276 8212 5964
rect 8703 3276 11619 5964
rect 12110 3276 15026 5964
rect 15517 3276 18433 5964
rect -18553 196 -15637 2884
rect -15146 196 -12230 2884
rect -11739 196 -8823 2884
rect -8332 196 -5416 2884
rect -4925 196 -2009 2884
rect -1518 196 1398 2884
rect 1889 196 4805 2884
rect 5296 196 8212 2884
rect 8703 196 11619 2884
rect 12110 196 15026 2884
rect 15517 196 18433 2884
rect -18553 -2884 -15637 -196
rect -15146 -2884 -12230 -196
rect -11739 -2884 -8823 -196
rect -8332 -2884 -5416 -196
rect -4925 -2884 -2009 -196
rect -1518 -2884 1398 -196
rect 1889 -2884 4805 -196
rect 5296 -2884 8212 -196
rect 8703 -2884 11619 -196
rect 12110 -2884 15026 -196
rect 15517 -2884 18433 -196
rect -18553 -5964 -15637 -3276
rect -15146 -5964 -12230 -3276
rect -11739 -5964 -8823 -3276
rect -8332 -5964 -5416 -3276
rect -4925 -5964 -2009 -3276
rect -1518 -5964 1398 -3276
rect 1889 -5964 4805 -3276
rect 5296 -5964 8212 -3276
rect 8703 -5964 11619 -3276
rect 12110 -5964 15026 -3276
rect 15517 -5964 18433 -3276
rect -18553 -9044 -15637 -6356
rect -15146 -9044 -12230 -6356
rect -11739 -9044 -8823 -6356
rect -8332 -9044 -5416 -6356
rect -4925 -9044 -2009 -6356
rect -1518 -9044 1398 -6356
rect 1889 -9044 4805 -6356
rect 5296 -9044 8212 -6356
rect 8703 -9044 11619 -6356
rect 12110 -9044 15026 -6356
rect 15517 -9044 18433 -6356
rect -18553 -12124 -15637 -9436
rect -15146 -12124 -12230 -9436
rect -11739 -12124 -8823 -9436
rect -8332 -12124 -5416 -9436
rect -4925 -12124 -2009 -9436
rect -1518 -12124 1398 -9436
rect 1889 -12124 4805 -9436
rect 5296 -12124 8212 -9436
rect 8703 -12124 11619 -9436
rect 12110 -12124 15026 -9436
rect 15517 -12124 18433 -9436
rect -18553 -15204 -15637 -12516
rect -15146 -15204 -12230 -12516
rect -11739 -15204 -8823 -12516
rect -8332 -15204 -5416 -12516
rect -4925 -15204 -2009 -12516
rect -1518 -15204 1398 -12516
rect 1889 -15204 4805 -12516
rect 5296 -15204 8212 -12516
rect 8703 -15204 11619 -12516
rect 12110 -15204 15026 -12516
rect 15517 -15204 18433 -12516
rect -18553 -18284 -15637 -15596
rect -15146 -18284 -12230 -15596
rect -11739 -18284 -8823 -15596
rect -8332 -18284 -5416 -15596
rect -4925 -18284 -2009 -15596
rect -1518 -18284 1398 -15596
rect 1889 -18284 4805 -15596
rect 5296 -18284 8212 -15596
rect 8703 -18284 11619 -15596
rect 12110 -18284 15026 -15596
rect 15517 -18284 18433 -15596
<< metal4 >>
rect -18705 18410 -15365 18450
rect -18705 18390 -15432 18410
rect -18705 15490 -18645 18390
rect -15545 15490 -15432 18390
rect -18705 15470 -15432 15490
rect -15404 15470 -15365 18410
rect -18705 15430 -15365 15470
rect -15298 18410 -11958 18450
rect -15298 18390 -12025 18410
rect -15298 15490 -15238 18390
rect -12138 15490 -12025 18390
rect -15298 15470 -12025 15490
rect -11997 15470 -11958 18410
rect -15298 15430 -11958 15470
rect -11891 18410 -8551 18450
rect -11891 18390 -8618 18410
rect -11891 15490 -11831 18390
rect -8731 15490 -8618 18390
rect -11891 15470 -8618 15490
rect -8590 15470 -8551 18410
rect -11891 15430 -8551 15470
rect -8484 18410 -5144 18450
rect -8484 18390 -5211 18410
rect -8484 15490 -8424 18390
rect -5324 15490 -5211 18390
rect -8484 15470 -5211 15490
rect -5183 15470 -5144 18410
rect -8484 15430 -5144 15470
rect -5077 18410 -1737 18450
rect -5077 18390 -1804 18410
rect -5077 15490 -5017 18390
rect -1917 15490 -1804 18390
rect -5077 15470 -1804 15490
rect -1776 15470 -1737 18410
rect -5077 15430 -1737 15470
rect -1670 18410 1670 18450
rect -1670 18390 1603 18410
rect -1670 15490 -1610 18390
rect 1490 15490 1603 18390
rect -1670 15470 1603 15490
rect 1631 15470 1670 18410
rect -1670 15430 1670 15470
rect 1737 18410 5077 18450
rect 1737 18390 5010 18410
rect 1737 15490 1797 18390
rect 4897 15490 5010 18390
rect 1737 15470 5010 15490
rect 5038 15470 5077 18410
rect 1737 15430 5077 15470
rect 5144 18410 8484 18450
rect 5144 18390 8417 18410
rect 5144 15490 5204 18390
rect 8304 15490 8417 18390
rect 5144 15470 8417 15490
rect 8445 15470 8484 18410
rect 5144 15430 8484 15470
rect 8551 18410 11891 18450
rect 8551 18390 11824 18410
rect 8551 15490 8611 18390
rect 11711 15490 11824 18390
rect 8551 15470 11824 15490
rect 11852 15470 11891 18410
rect 8551 15430 11891 15470
rect 11958 18410 15298 18450
rect 11958 18390 15231 18410
rect 11958 15490 12018 18390
rect 15118 15490 15231 18390
rect 11958 15470 15231 15490
rect 15259 15470 15298 18410
rect 11958 15430 15298 15470
rect 15365 18410 18705 18450
rect 15365 18390 18638 18410
rect 15365 15490 15425 18390
rect 18525 15490 18638 18390
rect 15365 15470 18638 15490
rect 18666 15470 18705 18410
rect 15365 15430 18705 15470
rect -18705 15330 -15365 15370
rect -18705 15310 -15432 15330
rect -18705 12410 -18645 15310
rect -15545 12410 -15432 15310
rect -18705 12390 -15432 12410
rect -15404 12390 -15365 15330
rect -18705 12350 -15365 12390
rect -15298 15330 -11958 15370
rect -15298 15310 -12025 15330
rect -15298 12410 -15238 15310
rect -12138 12410 -12025 15310
rect -15298 12390 -12025 12410
rect -11997 12390 -11958 15330
rect -15298 12350 -11958 12390
rect -11891 15330 -8551 15370
rect -11891 15310 -8618 15330
rect -11891 12410 -11831 15310
rect -8731 12410 -8618 15310
rect -11891 12390 -8618 12410
rect -8590 12390 -8551 15330
rect -11891 12350 -8551 12390
rect -8484 15330 -5144 15370
rect -8484 15310 -5211 15330
rect -8484 12410 -8424 15310
rect -5324 12410 -5211 15310
rect -8484 12390 -5211 12410
rect -5183 12390 -5144 15330
rect -8484 12350 -5144 12390
rect -5077 15330 -1737 15370
rect -5077 15310 -1804 15330
rect -5077 12410 -5017 15310
rect -1917 12410 -1804 15310
rect -5077 12390 -1804 12410
rect -1776 12390 -1737 15330
rect -5077 12350 -1737 12390
rect -1670 15330 1670 15370
rect -1670 15310 1603 15330
rect -1670 12410 -1610 15310
rect 1490 12410 1603 15310
rect -1670 12390 1603 12410
rect 1631 12390 1670 15330
rect -1670 12350 1670 12390
rect 1737 15330 5077 15370
rect 1737 15310 5010 15330
rect 1737 12410 1797 15310
rect 4897 12410 5010 15310
rect 1737 12390 5010 12410
rect 5038 12390 5077 15330
rect 1737 12350 5077 12390
rect 5144 15330 8484 15370
rect 5144 15310 8417 15330
rect 5144 12410 5204 15310
rect 8304 12410 8417 15310
rect 5144 12390 8417 12410
rect 8445 12390 8484 15330
rect 5144 12350 8484 12390
rect 8551 15330 11891 15370
rect 8551 15310 11824 15330
rect 8551 12410 8611 15310
rect 11711 12410 11824 15310
rect 8551 12390 11824 12410
rect 11852 12390 11891 15330
rect 8551 12350 11891 12390
rect 11958 15330 15298 15370
rect 11958 15310 15231 15330
rect 11958 12410 12018 15310
rect 15118 12410 15231 15310
rect 11958 12390 15231 12410
rect 15259 12390 15298 15330
rect 11958 12350 15298 12390
rect 15365 15330 18705 15370
rect 15365 15310 18638 15330
rect 15365 12410 15425 15310
rect 18525 12410 18638 15310
rect 15365 12390 18638 12410
rect 18666 12390 18705 15330
rect 15365 12350 18705 12390
rect -18705 12250 -15365 12290
rect -18705 12230 -15432 12250
rect -18705 9330 -18645 12230
rect -15545 9330 -15432 12230
rect -18705 9310 -15432 9330
rect -15404 9310 -15365 12250
rect -18705 9270 -15365 9310
rect -15298 12250 -11958 12290
rect -15298 12230 -12025 12250
rect -15298 9330 -15238 12230
rect -12138 9330 -12025 12230
rect -15298 9310 -12025 9330
rect -11997 9310 -11958 12250
rect -15298 9270 -11958 9310
rect -11891 12250 -8551 12290
rect -11891 12230 -8618 12250
rect -11891 9330 -11831 12230
rect -8731 9330 -8618 12230
rect -11891 9310 -8618 9330
rect -8590 9310 -8551 12250
rect -11891 9270 -8551 9310
rect -8484 12250 -5144 12290
rect -8484 12230 -5211 12250
rect -8484 9330 -8424 12230
rect -5324 9330 -5211 12230
rect -8484 9310 -5211 9330
rect -5183 9310 -5144 12250
rect -8484 9270 -5144 9310
rect -5077 12250 -1737 12290
rect -5077 12230 -1804 12250
rect -5077 9330 -5017 12230
rect -1917 9330 -1804 12230
rect -5077 9310 -1804 9330
rect -1776 9310 -1737 12250
rect -5077 9270 -1737 9310
rect -1670 12250 1670 12290
rect -1670 12230 1603 12250
rect -1670 9330 -1610 12230
rect 1490 9330 1603 12230
rect -1670 9310 1603 9330
rect 1631 9310 1670 12250
rect -1670 9270 1670 9310
rect 1737 12250 5077 12290
rect 1737 12230 5010 12250
rect 1737 9330 1797 12230
rect 4897 9330 5010 12230
rect 1737 9310 5010 9330
rect 5038 9310 5077 12250
rect 1737 9270 5077 9310
rect 5144 12250 8484 12290
rect 5144 12230 8417 12250
rect 5144 9330 5204 12230
rect 8304 9330 8417 12230
rect 5144 9310 8417 9330
rect 8445 9310 8484 12250
rect 5144 9270 8484 9310
rect 8551 12250 11891 12290
rect 8551 12230 11824 12250
rect 8551 9330 8611 12230
rect 11711 9330 11824 12230
rect 8551 9310 11824 9330
rect 11852 9310 11891 12250
rect 8551 9270 11891 9310
rect 11958 12250 15298 12290
rect 11958 12230 15231 12250
rect 11958 9330 12018 12230
rect 15118 9330 15231 12230
rect 11958 9310 15231 9330
rect 15259 9310 15298 12250
rect 11958 9270 15298 9310
rect 15365 12250 18705 12290
rect 15365 12230 18638 12250
rect 15365 9330 15425 12230
rect 18525 9330 18638 12230
rect 15365 9310 18638 9330
rect 18666 9310 18705 12250
rect 15365 9270 18705 9310
rect -18705 9170 -15365 9210
rect -18705 9150 -15432 9170
rect -18705 6250 -18645 9150
rect -15545 6250 -15432 9150
rect -18705 6230 -15432 6250
rect -15404 6230 -15365 9170
rect -18705 6190 -15365 6230
rect -15298 9170 -11958 9210
rect -15298 9150 -12025 9170
rect -15298 6250 -15238 9150
rect -12138 6250 -12025 9150
rect -15298 6230 -12025 6250
rect -11997 6230 -11958 9170
rect -15298 6190 -11958 6230
rect -11891 9170 -8551 9210
rect -11891 9150 -8618 9170
rect -11891 6250 -11831 9150
rect -8731 6250 -8618 9150
rect -11891 6230 -8618 6250
rect -8590 6230 -8551 9170
rect -11891 6190 -8551 6230
rect -8484 9170 -5144 9210
rect -8484 9150 -5211 9170
rect -8484 6250 -8424 9150
rect -5324 6250 -5211 9150
rect -8484 6230 -5211 6250
rect -5183 6230 -5144 9170
rect -8484 6190 -5144 6230
rect -5077 9170 -1737 9210
rect -5077 9150 -1804 9170
rect -5077 6250 -5017 9150
rect -1917 6250 -1804 9150
rect -5077 6230 -1804 6250
rect -1776 6230 -1737 9170
rect -5077 6190 -1737 6230
rect -1670 9170 1670 9210
rect -1670 9150 1603 9170
rect -1670 6250 -1610 9150
rect 1490 6250 1603 9150
rect -1670 6230 1603 6250
rect 1631 6230 1670 9170
rect -1670 6190 1670 6230
rect 1737 9170 5077 9210
rect 1737 9150 5010 9170
rect 1737 6250 1797 9150
rect 4897 6250 5010 9150
rect 1737 6230 5010 6250
rect 5038 6230 5077 9170
rect 1737 6190 5077 6230
rect 5144 9170 8484 9210
rect 5144 9150 8417 9170
rect 5144 6250 5204 9150
rect 8304 6250 8417 9150
rect 5144 6230 8417 6250
rect 8445 6230 8484 9170
rect 5144 6190 8484 6230
rect 8551 9170 11891 9210
rect 8551 9150 11824 9170
rect 8551 6250 8611 9150
rect 11711 6250 11824 9150
rect 8551 6230 11824 6250
rect 11852 6230 11891 9170
rect 8551 6190 11891 6230
rect 11958 9170 15298 9210
rect 11958 9150 15231 9170
rect 11958 6250 12018 9150
rect 15118 6250 15231 9150
rect 11958 6230 15231 6250
rect 15259 6230 15298 9170
rect 11958 6190 15298 6230
rect 15365 9170 18705 9210
rect 15365 9150 18638 9170
rect 15365 6250 15425 9150
rect 18525 6250 18638 9150
rect 15365 6230 18638 6250
rect 18666 6230 18705 9170
rect 15365 6190 18705 6230
rect -18705 6090 -15365 6130
rect -18705 6070 -15432 6090
rect -18705 3170 -18645 6070
rect -15545 3170 -15432 6070
rect -18705 3150 -15432 3170
rect -15404 3150 -15365 6090
rect -18705 3110 -15365 3150
rect -15298 6090 -11958 6130
rect -15298 6070 -12025 6090
rect -15298 3170 -15238 6070
rect -12138 3170 -12025 6070
rect -15298 3150 -12025 3170
rect -11997 3150 -11958 6090
rect -15298 3110 -11958 3150
rect -11891 6090 -8551 6130
rect -11891 6070 -8618 6090
rect -11891 3170 -11831 6070
rect -8731 3170 -8618 6070
rect -11891 3150 -8618 3170
rect -8590 3150 -8551 6090
rect -11891 3110 -8551 3150
rect -8484 6090 -5144 6130
rect -8484 6070 -5211 6090
rect -8484 3170 -8424 6070
rect -5324 3170 -5211 6070
rect -8484 3150 -5211 3170
rect -5183 3150 -5144 6090
rect -8484 3110 -5144 3150
rect -5077 6090 -1737 6130
rect -5077 6070 -1804 6090
rect -5077 3170 -5017 6070
rect -1917 3170 -1804 6070
rect -5077 3150 -1804 3170
rect -1776 3150 -1737 6090
rect -5077 3110 -1737 3150
rect -1670 6090 1670 6130
rect -1670 6070 1603 6090
rect -1670 3170 -1610 6070
rect 1490 3170 1603 6070
rect -1670 3150 1603 3170
rect 1631 3150 1670 6090
rect -1670 3110 1670 3150
rect 1737 6090 5077 6130
rect 1737 6070 5010 6090
rect 1737 3170 1797 6070
rect 4897 3170 5010 6070
rect 1737 3150 5010 3170
rect 5038 3150 5077 6090
rect 1737 3110 5077 3150
rect 5144 6090 8484 6130
rect 5144 6070 8417 6090
rect 5144 3170 5204 6070
rect 8304 3170 8417 6070
rect 5144 3150 8417 3170
rect 8445 3150 8484 6090
rect 5144 3110 8484 3150
rect 8551 6090 11891 6130
rect 8551 6070 11824 6090
rect 8551 3170 8611 6070
rect 11711 3170 11824 6070
rect 8551 3150 11824 3170
rect 11852 3150 11891 6090
rect 8551 3110 11891 3150
rect 11958 6090 15298 6130
rect 11958 6070 15231 6090
rect 11958 3170 12018 6070
rect 15118 3170 15231 6070
rect 11958 3150 15231 3170
rect 15259 3150 15298 6090
rect 11958 3110 15298 3150
rect 15365 6090 18705 6130
rect 15365 6070 18638 6090
rect 15365 3170 15425 6070
rect 18525 3170 18638 6070
rect 15365 3150 18638 3170
rect 18666 3150 18705 6090
rect 15365 3110 18705 3150
rect -18705 3010 -15365 3050
rect -18705 2990 -15432 3010
rect -18705 90 -18645 2990
rect -15545 90 -15432 2990
rect -18705 70 -15432 90
rect -15404 70 -15365 3010
rect -18705 30 -15365 70
rect -15298 3010 -11958 3050
rect -15298 2990 -12025 3010
rect -15298 90 -15238 2990
rect -12138 90 -12025 2990
rect -15298 70 -12025 90
rect -11997 70 -11958 3010
rect -15298 30 -11958 70
rect -11891 3010 -8551 3050
rect -11891 2990 -8618 3010
rect -11891 90 -11831 2990
rect -8731 90 -8618 2990
rect -11891 70 -8618 90
rect -8590 70 -8551 3010
rect -11891 30 -8551 70
rect -8484 3010 -5144 3050
rect -8484 2990 -5211 3010
rect -8484 90 -8424 2990
rect -5324 90 -5211 2990
rect -8484 70 -5211 90
rect -5183 70 -5144 3010
rect -8484 30 -5144 70
rect -5077 3010 -1737 3050
rect -5077 2990 -1804 3010
rect -5077 90 -5017 2990
rect -1917 90 -1804 2990
rect -5077 70 -1804 90
rect -1776 70 -1737 3010
rect -5077 30 -1737 70
rect -1670 3010 1670 3050
rect -1670 2990 1603 3010
rect -1670 90 -1610 2990
rect 1490 90 1603 2990
rect -1670 70 1603 90
rect 1631 70 1670 3010
rect -1670 30 1670 70
rect 1737 3010 5077 3050
rect 1737 2990 5010 3010
rect 1737 90 1797 2990
rect 4897 90 5010 2990
rect 1737 70 5010 90
rect 5038 70 5077 3010
rect 1737 30 5077 70
rect 5144 3010 8484 3050
rect 5144 2990 8417 3010
rect 5144 90 5204 2990
rect 8304 90 8417 2990
rect 5144 70 8417 90
rect 8445 70 8484 3010
rect 5144 30 8484 70
rect 8551 3010 11891 3050
rect 8551 2990 11824 3010
rect 8551 90 8611 2990
rect 11711 90 11824 2990
rect 8551 70 11824 90
rect 11852 70 11891 3010
rect 8551 30 11891 70
rect 11958 3010 15298 3050
rect 11958 2990 15231 3010
rect 11958 90 12018 2990
rect 15118 90 15231 2990
rect 11958 70 15231 90
rect 15259 70 15298 3010
rect 11958 30 15298 70
rect 15365 3010 18705 3050
rect 15365 2990 18638 3010
rect 15365 90 15425 2990
rect 18525 90 18638 2990
rect 15365 70 18638 90
rect 18666 70 18705 3010
rect 15365 30 18705 70
rect -18705 -70 -15365 -30
rect -18705 -90 -15432 -70
rect -18705 -2990 -18645 -90
rect -15545 -2990 -15432 -90
rect -18705 -3010 -15432 -2990
rect -15404 -3010 -15365 -70
rect -18705 -3050 -15365 -3010
rect -15298 -70 -11958 -30
rect -15298 -90 -12025 -70
rect -15298 -2990 -15238 -90
rect -12138 -2990 -12025 -90
rect -15298 -3010 -12025 -2990
rect -11997 -3010 -11958 -70
rect -15298 -3050 -11958 -3010
rect -11891 -70 -8551 -30
rect -11891 -90 -8618 -70
rect -11891 -2990 -11831 -90
rect -8731 -2990 -8618 -90
rect -11891 -3010 -8618 -2990
rect -8590 -3010 -8551 -70
rect -11891 -3050 -8551 -3010
rect -8484 -70 -5144 -30
rect -8484 -90 -5211 -70
rect -8484 -2990 -8424 -90
rect -5324 -2990 -5211 -90
rect -8484 -3010 -5211 -2990
rect -5183 -3010 -5144 -70
rect -8484 -3050 -5144 -3010
rect -5077 -70 -1737 -30
rect -5077 -90 -1804 -70
rect -5077 -2990 -5017 -90
rect -1917 -2990 -1804 -90
rect -5077 -3010 -1804 -2990
rect -1776 -3010 -1737 -70
rect -5077 -3050 -1737 -3010
rect -1670 -70 1670 -30
rect -1670 -90 1603 -70
rect -1670 -2990 -1610 -90
rect 1490 -2990 1603 -90
rect -1670 -3010 1603 -2990
rect 1631 -3010 1670 -70
rect -1670 -3050 1670 -3010
rect 1737 -70 5077 -30
rect 1737 -90 5010 -70
rect 1737 -2990 1797 -90
rect 4897 -2990 5010 -90
rect 1737 -3010 5010 -2990
rect 5038 -3010 5077 -70
rect 1737 -3050 5077 -3010
rect 5144 -70 8484 -30
rect 5144 -90 8417 -70
rect 5144 -2990 5204 -90
rect 8304 -2990 8417 -90
rect 5144 -3010 8417 -2990
rect 8445 -3010 8484 -70
rect 5144 -3050 8484 -3010
rect 8551 -70 11891 -30
rect 8551 -90 11824 -70
rect 8551 -2990 8611 -90
rect 11711 -2990 11824 -90
rect 8551 -3010 11824 -2990
rect 11852 -3010 11891 -70
rect 8551 -3050 11891 -3010
rect 11958 -70 15298 -30
rect 11958 -90 15231 -70
rect 11958 -2990 12018 -90
rect 15118 -2990 15231 -90
rect 11958 -3010 15231 -2990
rect 15259 -3010 15298 -70
rect 11958 -3050 15298 -3010
rect 15365 -70 18705 -30
rect 15365 -90 18638 -70
rect 15365 -2990 15425 -90
rect 18525 -2990 18638 -90
rect 15365 -3010 18638 -2990
rect 18666 -3010 18705 -70
rect 15365 -3050 18705 -3010
rect -18705 -3150 -15365 -3110
rect -18705 -3170 -15432 -3150
rect -18705 -6070 -18645 -3170
rect -15545 -6070 -15432 -3170
rect -18705 -6090 -15432 -6070
rect -15404 -6090 -15365 -3150
rect -18705 -6130 -15365 -6090
rect -15298 -3150 -11958 -3110
rect -15298 -3170 -12025 -3150
rect -15298 -6070 -15238 -3170
rect -12138 -6070 -12025 -3170
rect -15298 -6090 -12025 -6070
rect -11997 -6090 -11958 -3150
rect -15298 -6130 -11958 -6090
rect -11891 -3150 -8551 -3110
rect -11891 -3170 -8618 -3150
rect -11891 -6070 -11831 -3170
rect -8731 -6070 -8618 -3170
rect -11891 -6090 -8618 -6070
rect -8590 -6090 -8551 -3150
rect -11891 -6130 -8551 -6090
rect -8484 -3150 -5144 -3110
rect -8484 -3170 -5211 -3150
rect -8484 -6070 -8424 -3170
rect -5324 -6070 -5211 -3170
rect -8484 -6090 -5211 -6070
rect -5183 -6090 -5144 -3150
rect -8484 -6130 -5144 -6090
rect -5077 -3150 -1737 -3110
rect -5077 -3170 -1804 -3150
rect -5077 -6070 -5017 -3170
rect -1917 -6070 -1804 -3170
rect -5077 -6090 -1804 -6070
rect -1776 -6090 -1737 -3150
rect -5077 -6130 -1737 -6090
rect -1670 -3150 1670 -3110
rect -1670 -3170 1603 -3150
rect -1670 -6070 -1610 -3170
rect 1490 -6070 1603 -3170
rect -1670 -6090 1603 -6070
rect 1631 -6090 1670 -3150
rect -1670 -6130 1670 -6090
rect 1737 -3150 5077 -3110
rect 1737 -3170 5010 -3150
rect 1737 -6070 1797 -3170
rect 4897 -6070 5010 -3170
rect 1737 -6090 5010 -6070
rect 5038 -6090 5077 -3150
rect 1737 -6130 5077 -6090
rect 5144 -3150 8484 -3110
rect 5144 -3170 8417 -3150
rect 5144 -6070 5204 -3170
rect 8304 -6070 8417 -3170
rect 5144 -6090 8417 -6070
rect 8445 -6090 8484 -3150
rect 5144 -6130 8484 -6090
rect 8551 -3150 11891 -3110
rect 8551 -3170 11824 -3150
rect 8551 -6070 8611 -3170
rect 11711 -6070 11824 -3170
rect 8551 -6090 11824 -6070
rect 11852 -6090 11891 -3150
rect 8551 -6130 11891 -6090
rect 11958 -3150 15298 -3110
rect 11958 -3170 15231 -3150
rect 11958 -6070 12018 -3170
rect 15118 -6070 15231 -3170
rect 11958 -6090 15231 -6070
rect 15259 -6090 15298 -3150
rect 11958 -6130 15298 -6090
rect 15365 -3150 18705 -3110
rect 15365 -3170 18638 -3150
rect 15365 -6070 15425 -3170
rect 18525 -6070 18638 -3170
rect 15365 -6090 18638 -6070
rect 18666 -6090 18705 -3150
rect 15365 -6130 18705 -6090
rect -18705 -6230 -15365 -6190
rect -18705 -6250 -15432 -6230
rect -18705 -9150 -18645 -6250
rect -15545 -9150 -15432 -6250
rect -18705 -9170 -15432 -9150
rect -15404 -9170 -15365 -6230
rect -18705 -9210 -15365 -9170
rect -15298 -6230 -11958 -6190
rect -15298 -6250 -12025 -6230
rect -15298 -9150 -15238 -6250
rect -12138 -9150 -12025 -6250
rect -15298 -9170 -12025 -9150
rect -11997 -9170 -11958 -6230
rect -15298 -9210 -11958 -9170
rect -11891 -6230 -8551 -6190
rect -11891 -6250 -8618 -6230
rect -11891 -9150 -11831 -6250
rect -8731 -9150 -8618 -6250
rect -11891 -9170 -8618 -9150
rect -8590 -9170 -8551 -6230
rect -11891 -9210 -8551 -9170
rect -8484 -6230 -5144 -6190
rect -8484 -6250 -5211 -6230
rect -8484 -9150 -8424 -6250
rect -5324 -9150 -5211 -6250
rect -8484 -9170 -5211 -9150
rect -5183 -9170 -5144 -6230
rect -8484 -9210 -5144 -9170
rect -5077 -6230 -1737 -6190
rect -5077 -6250 -1804 -6230
rect -5077 -9150 -5017 -6250
rect -1917 -9150 -1804 -6250
rect -5077 -9170 -1804 -9150
rect -1776 -9170 -1737 -6230
rect -5077 -9210 -1737 -9170
rect -1670 -6230 1670 -6190
rect -1670 -6250 1603 -6230
rect -1670 -9150 -1610 -6250
rect 1490 -9150 1603 -6250
rect -1670 -9170 1603 -9150
rect 1631 -9170 1670 -6230
rect -1670 -9210 1670 -9170
rect 1737 -6230 5077 -6190
rect 1737 -6250 5010 -6230
rect 1737 -9150 1797 -6250
rect 4897 -9150 5010 -6250
rect 1737 -9170 5010 -9150
rect 5038 -9170 5077 -6230
rect 1737 -9210 5077 -9170
rect 5144 -6230 8484 -6190
rect 5144 -6250 8417 -6230
rect 5144 -9150 5204 -6250
rect 8304 -9150 8417 -6250
rect 5144 -9170 8417 -9150
rect 8445 -9170 8484 -6230
rect 5144 -9210 8484 -9170
rect 8551 -6230 11891 -6190
rect 8551 -6250 11824 -6230
rect 8551 -9150 8611 -6250
rect 11711 -9150 11824 -6250
rect 8551 -9170 11824 -9150
rect 11852 -9170 11891 -6230
rect 8551 -9210 11891 -9170
rect 11958 -6230 15298 -6190
rect 11958 -6250 15231 -6230
rect 11958 -9150 12018 -6250
rect 15118 -9150 15231 -6250
rect 11958 -9170 15231 -9150
rect 15259 -9170 15298 -6230
rect 11958 -9210 15298 -9170
rect 15365 -6230 18705 -6190
rect 15365 -6250 18638 -6230
rect 15365 -9150 15425 -6250
rect 18525 -9150 18638 -6250
rect 15365 -9170 18638 -9150
rect 18666 -9170 18705 -6230
rect 15365 -9210 18705 -9170
rect -18705 -9310 -15365 -9270
rect -18705 -9330 -15432 -9310
rect -18705 -12230 -18645 -9330
rect -15545 -12230 -15432 -9330
rect -18705 -12250 -15432 -12230
rect -15404 -12250 -15365 -9310
rect -18705 -12290 -15365 -12250
rect -15298 -9310 -11958 -9270
rect -15298 -9330 -12025 -9310
rect -15298 -12230 -15238 -9330
rect -12138 -12230 -12025 -9330
rect -15298 -12250 -12025 -12230
rect -11997 -12250 -11958 -9310
rect -15298 -12290 -11958 -12250
rect -11891 -9310 -8551 -9270
rect -11891 -9330 -8618 -9310
rect -11891 -12230 -11831 -9330
rect -8731 -12230 -8618 -9330
rect -11891 -12250 -8618 -12230
rect -8590 -12250 -8551 -9310
rect -11891 -12290 -8551 -12250
rect -8484 -9310 -5144 -9270
rect -8484 -9330 -5211 -9310
rect -8484 -12230 -8424 -9330
rect -5324 -12230 -5211 -9330
rect -8484 -12250 -5211 -12230
rect -5183 -12250 -5144 -9310
rect -8484 -12290 -5144 -12250
rect -5077 -9310 -1737 -9270
rect -5077 -9330 -1804 -9310
rect -5077 -12230 -5017 -9330
rect -1917 -12230 -1804 -9330
rect -5077 -12250 -1804 -12230
rect -1776 -12250 -1737 -9310
rect -5077 -12290 -1737 -12250
rect -1670 -9310 1670 -9270
rect -1670 -9330 1603 -9310
rect -1670 -12230 -1610 -9330
rect 1490 -12230 1603 -9330
rect -1670 -12250 1603 -12230
rect 1631 -12250 1670 -9310
rect -1670 -12290 1670 -12250
rect 1737 -9310 5077 -9270
rect 1737 -9330 5010 -9310
rect 1737 -12230 1797 -9330
rect 4897 -12230 5010 -9330
rect 1737 -12250 5010 -12230
rect 5038 -12250 5077 -9310
rect 1737 -12290 5077 -12250
rect 5144 -9310 8484 -9270
rect 5144 -9330 8417 -9310
rect 5144 -12230 5204 -9330
rect 8304 -12230 8417 -9330
rect 5144 -12250 8417 -12230
rect 8445 -12250 8484 -9310
rect 5144 -12290 8484 -12250
rect 8551 -9310 11891 -9270
rect 8551 -9330 11824 -9310
rect 8551 -12230 8611 -9330
rect 11711 -12230 11824 -9330
rect 8551 -12250 11824 -12230
rect 11852 -12250 11891 -9310
rect 8551 -12290 11891 -12250
rect 11958 -9310 15298 -9270
rect 11958 -9330 15231 -9310
rect 11958 -12230 12018 -9330
rect 15118 -12230 15231 -9330
rect 11958 -12250 15231 -12230
rect 15259 -12250 15298 -9310
rect 11958 -12290 15298 -12250
rect 15365 -9310 18705 -9270
rect 15365 -9330 18638 -9310
rect 15365 -12230 15425 -9330
rect 18525 -12230 18638 -9330
rect 15365 -12250 18638 -12230
rect 18666 -12250 18705 -9310
rect 15365 -12290 18705 -12250
rect -18705 -12390 -15365 -12350
rect -18705 -12410 -15432 -12390
rect -18705 -15310 -18645 -12410
rect -15545 -15310 -15432 -12410
rect -18705 -15330 -15432 -15310
rect -15404 -15330 -15365 -12390
rect -18705 -15370 -15365 -15330
rect -15298 -12390 -11958 -12350
rect -15298 -12410 -12025 -12390
rect -15298 -15310 -15238 -12410
rect -12138 -15310 -12025 -12410
rect -15298 -15330 -12025 -15310
rect -11997 -15330 -11958 -12390
rect -15298 -15370 -11958 -15330
rect -11891 -12390 -8551 -12350
rect -11891 -12410 -8618 -12390
rect -11891 -15310 -11831 -12410
rect -8731 -15310 -8618 -12410
rect -11891 -15330 -8618 -15310
rect -8590 -15330 -8551 -12390
rect -11891 -15370 -8551 -15330
rect -8484 -12390 -5144 -12350
rect -8484 -12410 -5211 -12390
rect -8484 -15310 -8424 -12410
rect -5324 -15310 -5211 -12410
rect -8484 -15330 -5211 -15310
rect -5183 -15330 -5144 -12390
rect -8484 -15370 -5144 -15330
rect -5077 -12390 -1737 -12350
rect -5077 -12410 -1804 -12390
rect -5077 -15310 -5017 -12410
rect -1917 -15310 -1804 -12410
rect -5077 -15330 -1804 -15310
rect -1776 -15330 -1737 -12390
rect -5077 -15370 -1737 -15330
rect -1670 -12390 1670 -12350
rect -1670 -12410 1603 -12390
rect -1670 -15310 -1610 -12410
rect 1490 -15310 1603 -12410
rect -1670 -15330 1603 -15310
rect 1631 -15330 1670 -12390
rect -1670 -15370 1670 -15330
rect 1737 -12390 5077 -12350
rect 1737 -12410 5010 -12390
rect 1737 -15310 1797 -12410
rect 4897 -15310 5010 -12410
rect 1737 -15330 5010 -15310
rect 5038 -15330 5077 -12390
rect 1737 -15370 5077 -15330
rect 5144 -12390 8484 -12350
rect 5144 -12410 8417 -12390
rect 5144 -15310 5204 -12410
rect 8304 -15310 8417 -12410
rect 5144 -15330 8417 -15310
rect 8445 -15330 8484 -12390
rect 5144 -15370 8484 -15330
rect 8551 -12390 11891 -12350
rect 8551 -12410 11824 -12390
rect 8551 -15310 8611 -12410
rect 11711 -15310 11824 -12410
rect 8551 -15330 11824 -15310
rect 11852 -15330 11891 -12390
rect 8551 -15370 11891 -15330
rect 11958 -12390 15298 -12350
rect 11958 -12410 15231 -12390
rect 11958 -15310 12018 -12410
rect 15118 -15310 15231 -12410
rect 11958 -15330 15231 -15310
rect 15259 -15330 15298 -12390
rect 11958 -15370 15298 -15330
rect 15365 -12390 18705 -12350
rect 15365 -12410 18638 -12390
rect 15365 -15310 15425 -12410
rect 18525 -15310 18638 -12410
rect 15365 -15330 18638 -15310
rect 18666 -15330 18705 -12390
rect 15365 -15370 18705 -15330
rect -18705 -15470 -15365 -15430
rect -18705 -15490 -15432 -15470
rect -18705 -18390 -18645 -15490
rect -15545 -18390 -15432 -15490
rect -18705 -18410 -15432 -18390
rect -15404 -18410 -15365 -15470
rect -18705 -18450 -15365 -18410
rect -15298 -15470 -11958 -15430
rect -15298 -15490 -12025 -15470
rect -15298 -18390 -15238 -15490
rect -12138 -18390 -12025 -15490
rect -15298 -18410 -12025 -18390
rect -11997 -18410 -11958 -15470
rect -15298 -18450 -11958 -18410
rect -11891 -15470 -8551 -15430
rect -11891 -15490 -8618 -15470
rect -11891 -18390 -11831 -15490
rect -8731 -18390 -8618 -15490
rect -11891 -18410 -8618 -18390
rect -8590 -18410 -8551 -15470
rect -11891 -18450 -8551 -18410
rect -8484 -15470 -5144 -15430
rect -8484 -15490 -5211 -15470
rect -8484 -18390 -8424 -15490
rect -5324 -18390 -5211 -15490
rect -8484 -18410 -5211 -18390
rect -5183 -18410 -5144 -15470
rect -8484 -18450 -5144 -18410
rect -5077 -15470 -1737 -15430
rect -5077 -15490 -1804 -15470
rect -5077 -18390 -5017 -15490
rect -1917 -18390 -1804 -15490
rect -5077 -18410 -1804 -18390
rect -1776 -18410 -1737 -15470
rect -5077 -18450 -1737 -18410
rect -1670 -15470 1670 -15430
rect -1670 -15490 1603 -15470
rect -1670 -18390 -1610 -15490
rect 1490 -18390 1603 -15490
rect -1670 -18410 1603 -18390
rect 1631 -18410 1670 -15470
rect -1670 -18450 1670 -18410
rect 1737 -15470 5077 -15430
rect 1737 -15490 5010 -15470
rect 1737 -18390 1797 -15490
rect 4897 -18390 5010 -15490
rect 1737 -18410 5010 -18390
rect 5038 -18410 5077 -15470
rect 1737 -18450 5077 -18410
rect 5144 -15470 8484 -15430
rect 5144 -15490 8417 -15470
rect 5144 -18390 5204 -15490
rect 8304 -18390 8417 -15490
rect 5144 -18410 8417 -18390
rect 8445 -18410 8484 -15470
rect 5144 -18450 8484 -18410
rect 8551 -15470 11891 -15430
rect 8551 -15490 11824 -15470
rect 8551 -18390 8611 -15490
rect 11711 -18390 11824 -15490
rect 8551 -18410 11824 -18390
rect 11852 -18410 11891 -15470
rect 8551 -18450 11891 -18410
rect 11958 -15470 15298 -15430
rect 11958 -15490 15231 -15470
rect 11958 -18390 12018 -15490
rect 15118 -18390 15231 -15490
rect 11958 -18410 15231 -18390
rect 15259 -18410 15298 -15470
rect 11958 -18450 15298 -18410
rect 15365 -15470 18705 -15430
rect 15365 -15490 18638 -15470
rect 15365 -18390 15425 -15490
rect 18525 -18390 18638 -15490
rect 15365 -18410 18638 -18390
rect 18666 -18410 18705 -15470
rect 15365 -18450 18705 -18410
<< via4 >>
rect -15432 15470 -15404 18410
rect -12025 15470 -11997 18410
rect -8618 15470 -8590 18410
rect -5211 15470 -5183 18410
rect -1804 15470 -1776 18410
rect 1603 15470 1631 18410
rect 5010 15470 5038 18410
rect 8417 15470 8445 18410
rect 11824 15470 11852 18410
rect 15231 15470 15259 18410
rect 18638 15470 18666 18410
rect -15432 12390 -15404 15330
rect -12025 12390 -11997 15330
rect -8618 12390 -8590 15330
rect -5211 12390 -5183 15330
rect -1804 12390 -1776 15330
rect 1603 12390 1631 15330
rect 5010 12390 5038 15330
rect 8417 12390 8445 15330
rect 11824 12390 11852 15330
rect 15231 12390 15259 15330
rect 18638 12390 18666 15330
rect -15432 9310 -15404 12250
rect -12025 9310 -11997 12250
rect -8618 9310 -8590 12250
rect -5211 9310 -5183 12250
rect -1804 9310 -1776 12250
rect 1603 9310 1631 12250
rect 5010 9310 5038 12250
rect 8417 9310 8445 12250
rect 11824 9310 11852 12250
rect 15231 9310 15259 12250
rect 18638 9310 18666 12250
rect -15432 6230 -15404 9170
rect -12025 6230 -11997 9170
rect -8618 6230 -8590 9170
rect -5211 6230 -5183 9170
rect -1804 6230 -1776 9170
rect 1603 6230 1631 9170
rect 5010 6230 5038 9170
rect 8417 6230 8445 9170
rect 11824 6230 11852 9170
rect 15231 6230 15259 9170
rect 18638 6230 18666 9170
rect -15432 3150 -15404 6090
rect -12025 3150 -11997 6090
rect -8618 3150 -8590 6090
rect -5211 3150 -5183 6090
rect -1804 3150 -1776 6090
rect 1603 3150 1631 6090
rect 5010 3150 5038 6090
rect 8417 3150 8445 6090
rect 11824 3150 11852 6090
rect 15231 3150 15259 6090
rect 18638 3150 18666 6090
rect -15432 70 -15404 3010
rect -12025 70 -11997 3010
rect -8618 70 -8590 3010
rect -5211 70 -5183 3010
rect -1804 70 -1776 3010
rect 1603 70 1631 3010
rect 5010 70 5038 3010
rect 8417 70 8445 3010
rect 11824 70 11852 3010
rect 15231 70 15259 3010
rect 18638 70 18666 3010
rect -15432 -3010 -15404 -70
rect -12025 -3010 -11997 -70
rect -8618 -3010 -8590 -70
rect -5211 -3010 -5183 -70
rect -1804 -3010 -1776 -70
rect 1603 -3010 1631 -70
rect 5010 -3010 5038 -70
rect 8417 -3010 8445 -70
rect 11824 -3010 11852 -70
rect 15231 -3010 15259 -70
rect 18638 -3010 18666 -70
rect -15432 -6090 -15404 -3150
rect -12025 -6090 -11997 -3150
rect -8618 -6090 -8590 -3150
rect -5211 -6090 -5183 -3150
rect -1804 -6090 -1776 -3150
rect 1603 -6090 1631 -3150
rect 5010 -6090 5038 -3150
rect 8417 -6090 8445 -3150
rect 11824 -6090 11852 -3150
rect 15231 -6090 15259 -3150
rect 18638 -6090 18666 -3150
rect -15432 -9170 -15404 -6230
rect -12025 -9170 -11997 -6230
rect -8618 -9170 -8590 -6230
rect -5211 -9170 -5183 -6230
rect -1804 -9170 -1776 -6230
rect 1603 -9170 1631 -6230
rect 5010 -9170 5038 -6230
rect 8417 -9170 8445 -6230
rect 11824 -9170 11852 -6230
rect 15231 -9170 15259 -6230
rect 18638 -9170 18666 -6230
rect -15432 -12250 -15404 -9310
rect -12025 -12250 -11997 -9310
rect -8618 -12250 -8590 -9310
rect -5211 -12250 -5183 -9310
rect -1804 -12250 -1776 -9310
rect 1603 -12250 1631 -9310
rect 5010 -12250 5038 -9310
rect 8417 -12250 8445 -9310
rect 11824 -12250 11852 -9310
rect 15231 -12250 15259 -9310
rect 18638 -12250 18666 -9310
rect -15432 -15330 -15404 -12390
rect -12025 -15330 -11997 -12390
rect -8618 -15330 -8590 -12390
rect -5211 -15330 -5183 -12390
rect -1804 -15330 -1776 -12390
rect 1603 -15330 1631 -12390
rect 5010 -15330 5038 -12390
rect 8417 -15330 8445 -12390
rect 11824 -15330 11852 -12390
rect 15231 -15330 15259 -12390
rect 18638 -15330 18666 -12390
rect -15432 -18410 -15404 -15470
rect -12025 -18410 -11997 -15470
rect -8618 -18410 -8590 -15470
rect -5211 -18410 -5183 -15470
rect -1804 -18410 -1776 -15470
rect 1603 -18410 1631 -15470
rect 5010 -18410 5038 -15470
rect 8417 -18410 8445 -15470
rect 11824 -18410 11852 -15470
rect 15231 -18410 15259 -15470
rect 18638 -18410 18666 -15470
<< metal5 >>
rect -17148 18350 -17042 18480
rect -15471 18410 -15365 18480
rect -18605 18284 -15585 18350
rect -18605 15596 -18553 18284
rect -15637 15596 -15585 18284
rect -18605 15530 -15585 15596
rect -17148 15270 -17042 15530
rect -15471 15470 -15432 18410
rect -15404 15470 -15365 18410
rect -13741 18350 -13635 18480
rect -12064 18410 -11958 18480
rect -15198 18284 -12178 18350
rect -15198 15596 -15146 18284
rect -12230 15596 -12178 18284
rect -15198 15530 -12178 15596
rect -15471 15330 -15365 15470
rect -18605 15204 -15585 15270
rect -18605 12516 -18553 15204
rect -15637 12516 -15585 15204
rect -18605 12450 -15585 12516
rect -17148 12190 -17042 12450
rect -15471 12390 -15432 15330
rect -15404 12390 -15365 15330
rect -13741 15270 -13635 15530
rect -12064 15470 -12025 18410
rect -11997 15470 -11958 18410
rect -10334 18350 -10228 18480
rect -8657 18410 -8551 18480
rect -11791 18284 -8771 18350
rect -11791 15596 -11739 18284
rect -8823 15596 -8771 18284
rect -11791 15530 -8771 15596
rect -12064 15330 -11958 15470
rect -15198 15204 -12178 15270
rect -15198 12516 -15146 15204
rect -12230 12516 -12178 15204
rect -15198 12450 -12178 12516
rect -15471 12250 -15365 12390
rect -18605 12124 -15585 12190
rect -18605 9436 -18553 12124
rect -15637 9436 -15585 12124
rect -18605 9370 -15585 9436
rect -17148 9110 -17042 9370
rect -15471 9310 -15432 12250
rect -15404 9310 -15365 12250
rect -13741 12190 -13635 12450
rect -12064 12390 -12025 15330
rect -11997 12390 -11958 15330
rect -10334 15270 -10228 15530
rect -8657 15470 -8618 18410
rect -8590 15470 -8551 18410
rect -6927 18350 -6821 18480
rect -5250 18410 -5144 18480
rect -8384 18284 -5364 18350
rect -8384 15596 -8332 18284
rect -5416 15596 -5364 18284
rect -8384 15530 -5364 15596
rect -8657 15330 -8551 15470
rect -11791 15204 -8771 15270
rect -11791 12516 -11739 15204
rect -8823 12516 -8771 15204
rect -11791 12450 -8771 12516
rect -12064 12250 -11958 12390
rect -15198 12124 -12178 12190
rect -15198 9436 -15146 12124
rect -12230 9436 -12178 12124
rect -15198 9370 -12178 9436
rect -15471 9170 -15365 9310
rect -18605 9044 -15585 9110
rect -18605 6356 -18553 9044
rect -15637 6356 -15585 9044
rect -18605 6290 -15585 6356
rect -17148 6030 -17042 6290
rect -15471 6230 -15432 9170
rect -15404 6230 -15365 9170
rect -13741 9110 -13635 9370
rect -12064 9310 -12025 12250
rect -11997 9310 -11958 12250
rect -10334 12190 -10228 12450
rect -8657 12390 -8618 15330
rect -8590 12390 -8551 15330
rect -6927 15270 -6821 15530
rect -5250 15470 -5211 18410
rect -5183 15470 -5144 18410
rect -3520 18350 -3414 18480
rect -1843 18410 -1737 18480
rect -4977 18284 -1957 18350
rect -4977 15596 -4925 18284
rect -2009 15596 -1957 18284
rect -4977 15530 -1957 15596
rect -5250 15330 -5144 15470
rect -8384 15204 -5364 15270
rect -8384 12516 -8332 15204
rect -5416 12516 -5364 15204
rect -8384 12450 -5364 12516
rect -8657 12250 -8551 12390
rect -11791 12124 -8771 12190
rect -11791 9436 -11739 12124
rect -8823 9436 -8771 12124
rect -11791 9370 -8771 9436
rect -12064 9170 -11958 9310
rect -15198 9044 -12178 9110
rect -15198 6356 -15146 9044
rect -12230 6356 -12178 9044
rect -15198 6290 -12178 6356
rect -15471 6090 -15365 6230
rect -18605 5964 -15585 6030
rect -18605 3276 -18553 5964
rect -15637 3276 -15585 5964
rect -18605 3210 -15585 3276
rect -17148 2950 -17042 3210
rect -15471 3150 -15432 6090
rect -15404 3150 -15365 6090
rect -13741 6030 -13635 6290
rect -12064 6230 -12025 9170
rect -11997 6230 -11958 9170
rect -10334 9110 -10228 9370
rect -8657 9310 -8618 12250
rect -8590 9310 -8551 12250
rect -6927 12190 -6821 12450
rect -5250 12390 -5211 15330
rect -5183 12390 -5144 15330
rect -3520 15270 -3414 15530
rect -1843 15470 -1804 18410
rect -1776 15470 -1737 18410
rect -113 18350 -7 18480
rect 1564 18410 1670 18480
rect -1570 18284 1450 18350
rect -1570 15596 -1518 18284
rect 1398 15596 1450 18284
rect -1570 15530 1450 15596
rect -1843 15330 -1737 15470
rect -4977 15204 -1957 15270
rect -4977 12516 -4925 15204
rect -2009 12516 -1957 15204
rect -4977 12450 -1957 12516
rect -5250 12250 -5144 12390
rect -8384 12124 -5364 12190
rect -8384 9436 -8332 12124
rect -5416 9436 -5364 12124
rect -8384 9370 -5364 9436
rect -8657 9170 -8551 9310
rect -11791 9044 -8771 9110
rect -11791 6356 -11739 9044
rect -8823 6356 -8771 9044
rect -11791 6290 -8771 6356
rect -12064 6090 -11958 6230
rect -15198 5964 -12178 6030
rect -15198 3276 -15146 5964
rect -12230 3276 -12178 5964
rect -15198 3210 -12178 3276
rect -15471 3010 -15365 3150
rect -18605 2884 -15585 2950
rect -18605 196 -18553 2884
rect -15637 196 -15585 2884
rect -18605 130 -15585 196
rect -17148 -130 -17042 130
rect -15471 70 -15432 3010
rect -15404 70 -15365 3010
rect -13741 2950 -13635 3210
rect -12064 3150 -12025 6090
rect -11997 3150 -11958 6090
rect -10334 6030 -10228 6290
rect -8657 6230 -8618 9170
rect -8590 6230 -8551 9170
rect -6927 9110 -6821 9370
rect -5250 9310 -5211 12250
rect -5183 9310 -5144 12250
rect -3520 12190 -3414 12450
rect -1843 12390 -1804 15330
rect -1776 12390 -1737 15330
rect -113 15270 -7 15530
rect 1564 15470 1603 18410
rect 1631 15470 1670 18410
rect 3294 18350 3400 18480
rect 4971 18410 5077 18480
rect 1837 18284 4857 18350
rect 1837 15596 1889 18284
rect 4805 15596 4857 18284
rect 1837 15530 4857 15596
rect 1564 15330 1670 15470
rect -1570 15204 1450 15270
rect -1570 12516 -1518 15204
rect 1398 12516 1450 15204
rect -1570 12450 1450 12516
rect -1843 12250 -1737 12390
rect -4977 12124 -1957 12190
rect -4977 9436 -4925 12124
rect -2009 9436 -1957 12124
rect -4977 9370 -1957 9436
rect -5250 9170 -5144 9310
rect -8384 9044 -5364 9110
rect -8384 6356 -8332 9044
rect -5416 6356 -5364 9044
rect -8384 6290 -5364 6356
rect -8657 6090 -8551 6230
rect -11791 5964 -8771 6030
rect -11791 3276 -11739 5964
rect -8823 3276 -8771 5964
rect -11791 3210 -8771 3276
rect -12064 3010 -11958 3150
rect -15198 2884 -12178 2950
rect -15198 196 -15146 2884
rect -12230 196 -12178 2884
rect -15198 130 -12178 196
rect -15471 -70 -15365 70
rect -18605 -196 -15585 -130
rect -18605 -2884 -18553 -196
rect -15637 -2884 -15585 -196
rect -18605 -2950 -15585 -2884
rect -17148 -3210 -17042 -2950
rect -15471 -3010 -15432 -70
rect -15404 -3010 -15365 -70
rect -13741 -130 -13635 130
rect -12064 70 -12025 3010
rect -11997 70 -11958 3010
rect -10334 2950 -10228 3210
rect -8657 3150 -8618 6090
rect -8590 3150 -8551 6090
rect -6927 6030 -6821 6290
rect -5250 6230 -5211 9170
rect -5183 6230 -5144 9170
rect -3520 9110 -3414 9370
rect -1843 9310 -1804 12250
rect -1776 9310 -1737 12250
rect -113 12190 -7 12450
rect 1564 12390 1603 15330
rect 1631 12390 1670 15330
rect 3294 15270 3400 15530
rect 4971 15470 5010 18410
rect 5038 15470 5077 18410
rect 6701 18350 6807 18480
rect 8378 18410 8484 18480
rect 5244 18284 8264 18350
rect 5244 15596 5296 18284
rect 8212 15596 8264 18284
rect 5244 15530 8264 15596
rect 4971 15330 5077 15470
rect 1837 15204 4857 15270
rect 1837 12516 1889 15204
rect 4805 12516 4857 15204
rect 1837 12450 4857 12516
rect 1564 12250 1670 12390
rect -1570 12124 1450 12190
rect -1570 9436 -1518 12124
rect 1398 9436 1450 12124
rect -1570 9370 1450 9436
rect -1843 9170 -1737 9310
rect -4977 9044 -1957 9110
rect -4977 6356 -4925 9044
rect -2009 6356 -1957 9044
rect -4977 6290 -1957 6356
rect -5250 6090 -5144 6230
rect -8384 5964 -5364 6030
rect -8384 3276 -8332 5964
rect -5416 3276 -5364 5964
rect -8384 3210 -5364 3276
rect -8657 3010 -8551 3150
rect -11791 2884 -8771 2950
rect -11791 196 -11739 2884
rect -8823 196 -8771 2884
rect -11791 130 -8771 196
rect -12064 -70 -11958 70
rect -15198 -196 -12178 -130
rect -15198 -2884 -15146 -196
rect -12230 -2884 -12178 -196
rect -15198 -2950 -12178 -2884
rect -15471 -3150 -15365 -3010
rect -18605 -3276 -15585 -3210
rect -18605 -5964 -18553 -3276
rect -15637 -5964 -15585 -3276
rect -18605 -6030 -15585 -5964
rect -17148 -6290 -17042 -6030
rect -15471 -6090 -15432 -3150
rect -15404 -6090 -15365 -3150
rect -13741 -3210 -13635 -2950
rect -12064 -3010 -12025 -70
rect -11997 -3010 -11958 -70
rect -10334 -130 -10228 130
rect -8657 70 -8618 3010
rect -8590 70 -8551 3010
rect -6927 2950 -6821 3210
rect -5250 3150 -5211 6090
rect -5183 3150 -5144 6090
rect -3520 6030 -3414 6290
rect -1843 6230 -1804 9170
rect -1776 6230 -1737 9170
rect -113 9110 -7 9370
rect 1564 9310 1603 12250
rect 1631 9310 1670 12250
rect 3294 12190 3400 12450
rect 4971 12390 5010 15330
rect 5038 12390 5077 15330
rect 6701 15270 6807 15530
rect 8378 15470 8417 18410
rect 8445 15470 8484 18410
rect 10108 18350 10214 18480
rect 11785 18410 11891 18480
rect 8651 18284 11671 18350
rect 8651 15596 8703 18284
rect 11619 15596 11671 18284
rect 8651 15530 11671 15596
rect 8378 15330 8484 15470
rect 5244 15204 8264 15270
rect 5244 12516 5296 15204
rect 8212 12516 8264 15204
rect 5244 12450 8264 12516
rect 4971 12250 5077 12390
rect 1837 12124 4857 12190
rect 1837 9436 1889 12124
rect 4805 9436 4857 12124
rect 1837 9370 4857 9436
rect 1564 9170 1670 9310
rect -1570 9044 1450 9110
rect -1570 6356 -1518 9044
rect 1398 6356 1450 9044
rect -1570 6290 1450 6356
rect -1843 6090 -1737 6230
rect -4977 5964 -1957 6030
rect -4977 3276 -4925 5964
rect -2009 3276 -1957 5964
rect -4977 3210 -1957 3276
rect -5250 3010 -5144 3150
rect -8384 2884 -5364 2950
rect -8384 196 -8332 2884
rect -5416 196 -5364 2884
rect -8384 130 -5364 196
rect -8657 -70 -8551 70
rect -11791 -196 -8771 -130
rect -11791 -2884 -11739 -196
rect -8823 -2884 -8771 -196
rect -11791 -2950 -8771 -2884
rect -12064 -3150 -11958 -3010
rect -15198 -3276 -12178 -3210
rect -15198 -5964 -15146 -3276
rect -12230 -5964 -12178 -3276
rect -15198 -6030 -12178 -5964
rect -15471 -6230 -15365 -6090
rect -18605 -6356 -15585 -6290
rect -18605 -9044 -18553 -6356
rect -15637 -9044 -15585 -6356
rect -18605 -9110 -15585 -9044
rect -17148 -9370 -17042 -9110
rect -15471 -9170 -15432 -6230
rect -15404 -9170 -15365 -6230
rect -13741 -6290 -13635 -6030
rect -12064 -6090 -12025 -3150
rect -11997 -6090 -11958 -3150
rect -10334 -3210 -10228 -2950
rect -8657 -3010 -8618 -70
rect -8590 -3010 -8551 -70
rect -6927 -130 -6821 130
rect -5250 70 -5211 3010
rect -5183 70 -5144 3010
rect -3520 2950 -3414 3210
rect -1843 3150 -1804 6090
rect -1776 3150 -1737 6090
rect -113 6030 -7 6290
rect 1564 6230 1603 9170
rect 1631 6230 1670 9170
rect 3294 9110 3400 9370
rect 4971 9310 5010 12250
rect 5038 9310 5077 12250
rect 6701 12190 6807 12450
rect 8378 12390 8417 15330
rect 8445 12390 8484 15330
rect 10108 15270 10214 15530
rect 11785 15470 11824 18410
rect 11852 15470 11891 18410
rect 13515 18350 13621 18480
rect 15192 18410 15298 18480
rect 12058 18284 15078 18350
rect 12058 15596 12110 18284
rect 15026 15596 15078 18284
rect 12058 15530 15078 15596
rect 11785 15330 11891 15470
rect 8651 15204 11671 15270
rect 8651 12516 8703 15204
rect 11619 12516 11671 15204
rect 8651 12450 11671 12516
rect 8378 12250 8484 12390
rect 5244 12124 8264 12190
rect 5244 9436 5296 12124
rect 8212 9436 8264 12124
rect 5244 9370 8264 9436
rect 4971 9170 5077 9310
rect 1837 9044 4857 9110
rect 1837 6356 1889 9044
rect 4805 6356 4857 9044
rect 1837 6290 4857 6356
rect 1564 6090 1670 6230
rect -1570 5964 1450 6030
rect -1570 3276 -1518 5964
rect 1398 3276 1450 5964
rect -1570 3210 1450 3276
rect -1843 3010 -1737 3150
rect -4977 2884 -1957 2950
rect -4977 196 -4925 2884
rect -2009 196 -1957 2884
rect -4977 130 -1957 196
rect -5250 -70 -5144 70
rect -8384 -196 -5364 -130
rect -8384 -2884 -8332 -196
rect -5416 -2884 -5364 -196
rect -8384 -2950 -5364 -2884
rect -8657 -3150 -8551 -3010
rect -11791 -3276 -8771 -3210
rect -11791 -5964 -11739 -3276
rect -8823 -5964 -8771 -3276
rect -11791 -6030 -8771 -5964
rect -12064 -6230 -11958 -6090
rect -15198 -6356 -12178 -6290
rect -15198 -9044 -15146 -6356
rect -12230 -9044 -12178 -6356
rect -15198 -9110 -12178 -9044
rect -15471 -9310 -15365 -9170
rect -18605 -9436 -15585 -9370
rect -18605 -12124 -18553 -9436
rect -15637 -12124 -15585 -9436
rect -18605 -12190 -15585 -12124
rect -17148 -12450 -17042 -12190
rect -15471 -12250 -15432 -9310
rect -15404 -12250 -15365 -9310
rect -13741 -9370 -13635 -9110
rect -12064 -9170 -12025 -6230
rect -11997 -9170 -11958 -6230
rect -10334 -6290 -10228 -6030
rect -8657 -6090 -8618 -3150
rect -8590 -6090 -8551 -3150
rect -6927 -3210 -6821 -2950
rect -5250 -3010 -5211 -70
rect -5183 -3010 -5144 -70
rect -3520 -130 -3414 130
rect -1843 70 -1804 3010
rect -1776 70 -1737 3010
rect -113 2950 -7 3210
rect 1564 3150 1603 6090
rect 1631 3150 1670 6090
rect 3294 6030 3400 6290
rect 4971 6230 5010 9170
rect 5038 6230 5077 9170
rect 6701 9110 6807 9370
rect 8378 9310 8417 12250
rect 8445 9310 8484 12250
rect 10108 12190 10214 12450
rect 11785 12390 11824 15330
rect 11852 12390 11891 15330
rect 13515 15270 13621 15530
rect 15192 15470 15231 18410
rect 15259 15470 15298 18410
rect 16922 18350 17028 18480
rect 18599 18410 18705 18480
rect 15465 18284 18485 18350
rect 15465 15596 15517 18284
rect 18433 15596 18485 18284
rect 15465 15530 18485 15596
rect 15192 15330 15298 15470
rect 12058 15204 15078 15270
rect 12058 12516 12110 15204
rect 15026 12516 15078 15204
rect 12058 12450 15078 12516
rect 11785 12250 11891 12390
rect 8651 12124 11671 12190
rect 8651 9436 8703 12124
rect 11619 9436 11671 12124
rect 8651 9370 11671 9436
rect 8378 9170 8484 9310
rect 5244 9044 8264 9110
rect 5244 6356 5296 9044
rect 8212 6356 8264 9044
rect 5244 6290 8264 6356
rect 4971 6090 5077 6230
rect 1837 5964 4857 6030
rect 1837 3276 1889 5964
rect 4805 3276 4857 5964
rect 1837 3210 4857 3276
rect 1564 3010 1670 3150
rect -1570 2884 1450 2950
rect -1570 196 -1518 2884
rect 1398 196 1450 2884
rect -1570 130 1450 196
rect -1843 -70 -1737 70
rect -4977 -196 -1957 -130
rect -4977 -2884 -4925 -196
rect -2009 -2884 -1957 -196
rect -4977 -2950 -1957 -2884
rect -5250 -3150 -5144 -3010
rect -8384 -3276 -5364 -3210
rect -8384 -5964 -8332 -3276
rect -5416 -5964 -5364 -3276
rect -8384 -6030 -5364 -5964
rect -8657 -6230 -8551 -6090
rect -11791 -6356 -8771 -6290
rect -11791 -9044 -11739 -6356
rect -8823 -9044 -8771 -6356
rect -11791 -9110 -8771 -9044
rect -12064 -9310 -11958 -9170
rect -15198 -9436 -12178 -9370
rect -15198 -12124 -15146 -9436
rect -12230 -12124 -12178 -9436
rect -15198 -12190 -12178 -12124
rect -15471 -12390 -15365 -12250
rect -18605 -12516 -15585 -12450
rect -18605 -15204 -18553 -12516
rect -15637 -15204 -15585 -12516
rect -18605 -15270 -15585 -15204
rect -17148 -15530 -17042 -15270
rect -15471 -15330 -15432 -12390
rect -15404 -15330 -15365 -12390
rect -13741 -12450 -13635 -12190
rect -12064 -12250 -12025 -9310
rect -11997 -12250 -11958 -9310
rect -10334 -9370 -10228 -9110
rect -8657 -9170 -8618 -6230
rect -8590 -9170 -8551 -6230
rect -6927 -6290 -6821 -6030
rect -5250 -6090 -5211 -3150
rect -5183 -6090 -5144 -3150
rect -3520 -3210 -3414 -2950
rect -1843 -3010 -1804 -70
rect -1776 -3010 -1737 -70
rect -113 -130 -7 130
rect 1564 70 1603 3010
rect 1631 70 1670 3010
rect 3294 2950 3400 3210
rect 4971 3150 5010 6090
rect 5038 3150 5077 6090
rect 6701 6030 6807 6290
rect 8378 6230 8417 9170
rect 8445 6230 8484 9170
rect 10108 9110 10214 9370
rect 11785 9310 11824 12250
rect 11852 9310 11891 12250
rect 13515 12190 13621 12450
rect 15192 12390 15231 15330
rect 15259 12390 15298 15330
rect 16922 15270 17028 15530
rect 18599 15470 18638 18410
rect 18666 15470 18705 18410
rect 18599 15330 18705 15470
rect 15465 15204 18485 15270
rect 15465 12516 15517 15204
rect 18433 12516 18485 15204
rect 15465 12450 18485 12516
rect 15192 12250 15298 12390
rect 12058 12124 15078 12190
rect 12058 9436 12110 12124
rect 15026 9436 15078 12124
rect 12058 9370 15078 9436
rect 11785 9170 11891 9310
rect 8651 9044 11671 9110
rect 8651 6356 8703 9044
rect 11619 6356 11671 9044
rect 8651 6290 11671 6356
rect 8378 6090 8484 6230
rect 5244 5964 8264 6030
rect 5244 3276 5296 5964
rect 8212 3276 8264 5964
rect 5244 3210 8264 3276
rect 4971 3010 5077 3150
rect 1837 2884 4857 2950
rect 1837 196 1889 2884
rect 4805 196 4857 2884
rect 1837 130 4857 196
rect 1564 -70 1670 70
rect -1570 -196 1450 -130
rect -1570 -2884 -1518 -196
rect 1398 -2884 1450 -196
rect -1570 -2950 1450 -2884
rect -1843 -3150 -1737 -3010
rect -4977 -3276 -1957 -3210
rect -4977 -5964 -4925 -3276
rect -2009 -5964 -1957 -3276
rect -4977 -6030 -1957 -5964
rect -5250 -6230 -5144 -6090
rect -8384 -6356 -5364 -6290
rect -8384 -9044 -8332 -6356
rect -5416 -9044 -5364 -6356
rect -8384 -9110 -5364 -9044
rect -8657 -9310 -8551 -9170
rect -11791 -9436 -8771 -9370
rect -11791 -12124 -11739 -9436
rect -8823 -12124 -8771 -9436
rect -11791 -12190 -8771 -12124
rect -12064 -12390 -11958 -12250
rect -15198 -12516 -12178 -12450
rect -15198 -15204 -15146 -12516
rect -12230 -15204 -12178 -12516
rect -15198 -15270 -12178 -15204
rect -15471 -15470 -15365 -15330
rect -18605 -15596 -15585 -15530
rect -18605 -18284 -18553 -15596
rect -15637 -18284 -15585 -15596
rect -18605 -18350 -15585 -18284
rect -17148 -18480 -17042 -18350
rect -15471 -18410 -15432 -15470
rect -15404 -18410 -15365 -15470
rect -13741 -15530 -13635 -15270
rect -12064 -15330 -12025 -12390
rect -11997 -15330 -11958 -12390
rect -10334 -12450 -10228 -12190
rect -8657 -12250 -8618 -9310
rect -8590 -12250 -8551 -9310
rect -6927 -9370 -6821 -9110
rect -5250 -9170 -5211 -6230
rect -5183 -9170 -5144 -6230
rect -3520 -6290 -3414 -6030
rect -1843 -6090 -1804 -3150
rect -1776 -6090 -1737 -3150
rect -113 -3210 -7 -2950
rect 1564 -3010 1603 -70
rect 1631 -3010 1670 -70
rect 3294 -130 3400 130
rect 4971 70 5010 3010
rect 5038 70 5077 3010
rect 6701 2950 6807 3210
rect 8378 3150 8417 6090
rect 8445 3150 8484 6090
rect 10108 6030 10214 6290
rect 11785 6230 11824 9170
rect 11852 6230 11891 9170
rect 13515 9110 13621 9370
rect 15192 9310 15231 12250
rect 15259 9310 15298 12250
rect 16922 12190 17028 12450
rect 18599 12390 18638 15330
rect 18666 12390 18705 15330
rect 18599 12250 18705 12390
rect 15465 12124 18485 12190
rect 15465 9436 15517 12124
rect 18433 9436 18485 12124
rect 15465 9370 18485 9436
rect 15192 9170 15298 9310
rect 12058 9044 15078 9110
rect 12058 6356 12110 9044
rect 15026 6356 15078 9044
rect 12058 6290 15078 6356
rect 11785 6090 11891 6230
rect 8651 5964 11671 6030
rect 8651 3276 8703 5964
rect 11619 3276 11671 5964
rect 8651 3210 11671 3276
rect 8378 3010 8484 3150
rect 5244 2884 8264 2950
rect 5244 196 5296 2884
rect 8212 196 8264 2884
rect 5244 130 8264 196
rect 4971 -70 5077 70
rect 1837 -196 4857 -130
rect 1837 -2884 1889 -196
rect 4805 -2884 4857 -196
rect 1837 -2950 4857 -2884
rect 1564 -3150 1670 -3010
rect -1570 -3276 1450 -3210
rect -1570 -5964 -1518 -3276
rect 1398 -5964 1450 -3276
rect -1570 -6030 1450 -5964
rect -1843 -6230 -1737 -6090
rect -4977 -6356 -1957 -6290
rect -4977 -9044 -4925 -6356
rect -2009 -9044 -1957 -6356
rect -4977 -9110 -1957 -9044
rect -5250 -9310 -5144 -9170
rect -8384 -9436 -5364 -9370
rect -8384 -12124 -8332 -9436
rect -5416 -12124 -5364 -9436
rect -8384 -12190 -5364 -12124
rect -8657 -12390 -8551 -12250
rect -11791 -12516 -8771 -12450
rect -11791 -15204 -11739 -12516
rect -8823 -15204 -8771 -12516
rect -11791 -15270 -8771 -15204
rect -12064 -15470 -11958 -15330
rect -15198 -15596 -12178 -15530
rect -15198 -18284 -15146 -15596
rect -12230 -18284 -12178 -15596
rect -15198 -18350 -12178 -18284
rect -15471 -18480 -15365 -18410
rect -13741 -18480 -13635 -18350
rect -12064 -18410 -12025 -15470
rect -11997 -18410 -11958 -15470
rect -10334 -15530 -10228 -15270
rect -8657 -15330 -8618 -12390
rect -8590 -15330 -8551 -12390
rect -6927 -12450 -6821 -12190
rect -5250 -12250 -5211 -9310
rect -5183 -12250 -5144 -9310
rect -3520 -9370 -3414 -9110
rect -1843 -9170 -1804 -6230
rect -1776 -9170 -1737 -6230
rect -113 -6290 -7 -6030
rect 1564 -6090 1603 -3150
rect 1631 -6090 1670 -3150
rect 3294 -3210 3400 -2950
rect 4971 -3010 5010 -70
rect 5038 -3010 5077 -70
rect 6701 -130 6807 130
rect 8378 70 8417 3010
rect 8445 70 8484 3010
rect 10108 2950 10214 3210
rect 11785 3150 11824 6090
rect 11852 3150 11891 6090
rect 13515 6030 13621 6290
rect 15192 6230 15231 9170
rect 15259 6230 15298 9170
rect 16922 9110 17028 9370
rect 18599 9310 18638 12250
rect 18666 9310 18705 12250
rect 18599 9170 18705 9310
rect 15465 9044 18485 9110
rect 15465 6356 15517 9044
rect 18433 6356 18485 9044
rect 15465 6290 18485 6356
rect 15192 6090 15298 6230
rect 12058 5964 15078 6030
rect 12058 3276 12110 5964
rect 15026 3276 15078 5964
rect 12058 3210 15078 3276
rect 11785 3010 11891 3150
rect 8651 2884 11671 2950
rect 8651 196 8703 2884
rect 11619 196 11671 2884
rect 8651 130 11671 196
rect 8378 -70 8484 70
rect 5244 -196 8264 -130
rect 5244 -2884 5296 -196
rect 8212 -2884 8264 -196
rect 5244 -2950 8264 -2884
rect 4971 -3150 5077 -3010
rect 1837 -3276 4857 -3210
rect 1837 -5964 1889 -3276
rect 4805 -5964 4857 -3276
rect 1837 -6030 4857 -5964
rect 1564 -6230 1670 -6090
rect -1570 -6356 1450 -6290
rect -1570 -9044 -1518 -6356
rect 1398 -9044 1450 -6356
rect -1570 -9110 1450 -9044
rect -1843 -9310 -1737 -9170
rect -4977 -9436 -1957 -9370
rect -4977 -12124 -4925 -9436
rect -2009 -12124 -1957 -9436
rect -4977 -12190 -1957 -12124
rect -5250 -12390 -5144 -12250
rect -8384 -12516 -5364 -12450
rect -8384 -15204 -8332 -12516
rect -5416 -15204 -5364 -12516
rect -8384 -15270 -5364 -15204
rect -8657 -15470 -8551 -15330
rect -11791 -15596 -8771 -15530
rect -11791 -18284 -11739 -15596
rect -8823 -18284 -8771 -15596
rect -11791 -18350 -8771 -18284
rect -12064 -18480 -11958 -18410
rect -10334 -18480 -10228 -18350
rect -8657 -18410 -8618 -15470
rect -8590 -18410 -8551 -15470
rect -6927 -15530 -6821 -15270
rect -5250 -15330 -5211 -12390
rect -5183 -15330 -5144 -12390
rect -3520 -12450 -3414 -12190
rect -1843 -12250 -1804 -9310
rect -1776 -12250 -1737 -9310
rect -113 -9370 -7 -9110
rect 1564 -9170 1603 -6230
rect 1631 -9170 1670 -6230
rect 3294 -6290 3400 -6030
rect 4971 -6090 5010 -3150
rect 5038 -6090 5077 -3150
rect 6701 -3210 6807 -2950
rect 8378 -3010 8417 -70
rect 8445 -3010 8484 -70
rect 10108 -130 10214 130
rect 11785 70 11824 3010
rect 11852 70 11891 3010
rect 13515 2950 13621 3210
rect 15192 3150 15231 6090
rect 15259 3150 15298 6090
rect 16922 6030 17028 6290
rect 18599 6230 18638 9170
rect 18666 6230 18705 9170
rect 18599 6090 18705 6230
rect 15465 5964 18485 6030
rect 15465 3276 15517 5964
rect 18433 3276 18485 5964
rect 15465 3210 18485 3276
rect 15192 3010 15298 3150
rect 12058 2884 15078 2950
rect 12058 196 12110 2884
rect 15026 196 15078 2884
rect 12058 130 15078 196
rect 11785 -70 11891 70
rect 8651 -196 11671 -130
rect 8651 -2884 8703 -196
rect 11619 -2884 11671 -196
rect 8651 -2950 11671 -2884
rect 8378 -3150 8484 -3010
rect 5244 -3276 8264 -3210
rect 5244 -5964 5296 -3276
rect 8212 -5964 8264 -3276
rect 5244 -6030 8264 -5964
rect 4971 -6230 5077 -6090
rect 1837 -6356 4857 -6290
rect 1837 -9044 1889 -6356
rect 4805 -9044 4857 -6356
rect 1837 -9110 4857 -9044
rect 1564 -9310 1670 -9170
rect -1570 -9436 1450 -9370
rect -1570 -12124 -1518 -9436
rect 1398 -12124 1450 -9436
rect -1570 -12190 1450 -12124
rect -1843 -12390 -1737 -12250
rect -4977 -12516 -1957 -12450
rect -4977 -15204 -4925 -12516
rect -2009 -15204 -1957 -12516
rect -4977 -15270 -1957 -15204
rect -5250 -15470 -5144 -15330
rect -8384 -15596 -5364 -15530
rect -8384 -18284 -8332 -15596
rect -5416 -18284 -5364 -15596
rect -8384 -18350 -5364 -18284
rect -8657 -18480 -8551 -18410
rect -6927 -18480 -6821 -18350
rect -5250 -18410 -5211 -15470
rect -5183 -18410 -5144 -15470
rect -3520 -15530 -3414 -15270
rect -1843 -15330 -1804 -12390
rect -1776 -15330 -1737 -12390
rect -113 -12450 -7 -12190
rect 1564 -12250 1603 -9310
rect 1631 -12250 1670 -9310
rect 3294 -9370 3400 -9110
rect 4971 -9170 5010 -6230
rect 5038 -9170 5077 -6230
rect 6701 -6290 6807 -6030
rect 8378 -6090 8417 -3150
rect 8445 -6090 8484 -3150
rect 10108 -3210 10214 -2950
rect 11785 -3010 11824 -70
rect 11852 -3010 11891 -70
rect 13515 -130 13621 130
rect 15192 70 15231 3010
rect 15259 70 15298 3010
rect 16922 2950 17028 3210
rect 18599 3150 18638 6090
rect 18666 3150 18705 6090
rect 18599 3010 18705 3150
rect 15465 2884 18485 2950
rect 15465 196 15517 2884
rect 18433 196 18485 2884
rect 15465 130 18485 196
rect 15192 -70 15298 70
rect 12058 -196 15078 -130
rect 12058 -2884 12110 -196
rect 15026 -2884 15078 -196
rect 12058 -2950 15078 -2884
rect 11785 -3150 11891 -3010
rect 8651 -3276 11671 -3210
rect 8651 -5964 8703 -3276
rect 11619 -5964 11671 -3276
rect 8651 -6030 11671 -5964
rect 8378 -6230 8484 -6090
rect 5244 -6356 8264 -6290
rect 5244 -9044 5296 -6356
rect 8212 -9044 8264 -6356
rect 5244 -9110 8264 -9044
rect 4971 -9310 5077 -9170
rect 1837 -9436 4857 -9370
rect 1837 -12124 1889 -9436
rect 4805 -12124 4857 -9436
rect 1837 -12190 4857 -12124
rect 1564 -12390 1670 -12250
rect -1570 -12516 1450 -12450
rect -1570 -15204 -1518 -12516
rect 1398 -15204 1450 -12516
rect -1570 -15270 1450 -15204
rect -1843 -15470 -1737 -15330
rect -4977 -15596 -1957 -15530
rect -4977 -18284 -4925 -15596
rect -2009 -18284 -1957 -15596
rect -4977 -18350 -1957 -18284
rect -5250 -18480 -5144 -18410
rect -3520 -18480 -3414 -18350
rect -1843 -18410 -1804 -15470
rect -1776 -18410 -1737 -15470
rect -113 -15530 -7 -15270
rect 1564 -15330 1603 -12390
rect 1631 -15330 1670 -12390
rect 3294 -12450 3400 -12190
rect 4971 -12250 5010 -9310
rect 5038 -12250 5077 -9310
rect 6701 -9370 6807 -9110
rect 8378 -9170 8417 -6230
rect 8445 -9170 8484 -6230
rect 10108 -6290 10214 -6030
rect 11785 -6090 11824 -3150
rect 11852 -6090 11891 -3150
rect 13515 -3210 13621 -2950
rect 15192 -3010 15231 -70
rect 15259 -3010 15298 -70
rect 16922 -130 17028 130
rect 18599 70 18638 3010
rect 18666 70 18705 3010
rect 18599 -70 18705 70
rect 15465 -196 18485 -130
rect 15465 -2884 15517 -196
rect 18433 -2884 18485 -196
rect 15465 -2950 18485 -2884
rect 15192 -3150 15298 -3010
rect 12058 -3276 15078 -3210
rect 12058 -5964 12110 -3276
rect 15026 -5964 15078 -3276
rect 12058 -6030 15078 -5964
rect 11785 -6230 11891 -6090
rect 8651 -6356 11671 -6290
rect 8651 -9044 8703 -6356
rect 11619 -9044 11671 -6356
rect 8651 -9110 11671 -9044
rect 8378 -9310 8484 -9170
rect 5244 -9436 8264 -9370
rect 5244 -12124 5296 -9436
rect 8212 -12124 8264 -9436
rect 5244 -12190 8264 -12124
rect 4971 -12390 5077 -12250
rect 1837 -12516 4857 -12450
rect 1837 -15204 1889 -12516
rect 4805 -15204 4857 -12516
rect 1837 -15270 4857 -15204
rect 1564 -15470 1670 -15330
rect -1570 -15596 1450 -15530
rect -1570 -18284 -1518 -15596
rect 1398 -18284 1450 -15596
rect -1570 -18350 1450 -18284
rect -1843 -18480 -1737 -18410
rect -113 -18480 -7 -18350
rect 1564 -18410 1603 -15470
rect 1631 -18410 1670 -15470
rect 3294 -15530 3400 -15270
rect 4971 -15330 5010 -12390
rect 5038 -15330 5077 -12390
rect 6701 -12450 6807 -12190
rect 8378 -12250 8417 -9310
rect 8445 -12250 8484 -9310
rect 10108 -9370 10214 -9110
rect 11785 -9170 11824 -6230
rect 11852 -9170 11891 -6230
rect 13515 -6290 13621 -6030
rect 15192 -6090 15231 -3150
rect 15259 -6090 15298 -3150
rect 16922 -3210 17028 -2950
rect 18599 -3010 18638 -70
rect 18666 -3010 18705 -70
rect 18599 -3150 18705 -3010
rect 15465 -3276 18485 -3210
rect 15465 -5964 15517 -3276
rect 18433 -5964 18485 -3276
rect 15465 -6030 18485 -5964
rect 15192 -6230 15298 -6090
rect 12058 -6356 15078 -6290
rect 12058 -9044 12110 -6356
rect 15026 -9044 15078 -6356
rect 12058 -9110 15078 -9044
rect 11785 -9310 11891 -9170
rect 8651 -9436 11671 -9370
rect 8651 -12124 8703 -9436
rect 11619 -12124 11671 -9436
rect 8651 -12190 11671 -12124
rect 8378 -12390 8484 -12250
rect 5244 -12516 8264 -12450
rect 5244 -15204 5296 -12516
rect 8212 -15204 8264 -12516
rect 5244 -15270 8264 -15204
rect 4971 -15470 5077 -15330
rect 1837 -15596 4857 -15530
rect 1837 -18284 1889 -15596
rect 4805 -18284 4857 -15596
rect 1837 -18350 4857 -18284
rect 1564 -18480 1670 -18410
rect 3294 -18480 3400 -18350
rect 4971 -18410 5010 -15470
rect 5038 -18410 5077 -15470
rect 6701 -15530 6807 -15270
rect 8378 -15330 8417 -12390
rect 8445 -15330 8484 -12390
rect 10108 -12450 10214 -12190
rect 11785 -12250 11824 -9310
rect 11852 -12250 11891 -9310
rect 13515 -9370 13621 -9110
rect 15192 -9170 15231 -6230
rect 15259 -9170 15298 -6230
rect 16922 -6290 17028 -6030
rect 18599 -6090 18638 -3150
rect 18666 -6090 18705 -3150
rect 18599 -6230 18705 -6090
rect 15465 -6356 18485 -6290
rect 15465 -9044 15517 -6356
rect 18433 -9044 18485 -6356
rect 15465 -9110 18485 -9044
rect 15192 -9310 15298 -9170
rect 12058 -9436 15078 -9370
rect 12058 -12124 12110 -9436
rect 15026 -12124 15078 -9436
rect 12058 -12190 15078 -12124
rect 11785 -12390 11891 -12250
rect 8651 -12516 11671 -12450
rect 8651 -15204 8703 -12516
rect 11619 -15204 11671 -12516
rect 8651 -15270 11671 -15204
rect 8378 -15470 8484 -15330
rect 5244 -15596 8264 -15530
rect 5244 -18284 5296 -15596
rect 8212 -18284 8264 -15596
rect 5244 -18350 8264 -18284
rect 4971 -18480 5077 -18410
rect 6701 -18480 6807 -18350
rect 8378 -18410 8417 -15470
rect 8445 -18410 8484 -15470
rect 10108 -15530 10214 -15270
rect 11785 -15330 11824 -12390
rect 11852 -15330 11891 -12390
rect 13515 -12450 13621 -12190
rect 15192 -12250 15231 -9310
rect 15259 -12250 15298 -9310
rect 16922 -9370 17028 -9110
rect 18599 -9170 18638 -6230
rect 18666 -9170 18705 -6230
rect 18599 -9310 18705 -9170
rect 15465 -9436 18485 -9370
rect 15465 -12124 15517 -9436
rect 18433 -12124 18485 -9436
rect 15465 -12190 18485 -12124
rect 15192 -12390 15298 -12250
rect 12058 -12516 15078 -12450
rect 12058 -15204 12110 -12516
rect 15026 -15204 15078 -12516
rect 12058 -15270 15078 -15204
rect 11785 -15470 11891 -15330
rect 8651 -15596 11671 -15530
rect 8651 -18284 8703 -15596
rect 11619 -18284 11671 -15596
rect 8651 -18350 11671 -18284
rect 8378 -18480 8484 -18410
rect 10108 -18480 10214 -18350
rect 11785 -18410 11824 -15470
rect 11852 -18410 11891 -15470
rect 13515 -15530 13621 -15270
rect 15192 -15330 15231 -12390
rect 15259 -15330 15298 -12390
rect 16922 -12450 17028 -12190
rect 18599 -12250 18638 -9310
rect 18666 -12250 18705 -9310
rect 18599 -12390 18705 -12250
rect 15465 -12516 18485 -12450
rect 15465 -15204 15517 -12516
rect 18433 -15204 18485 -12516
rect 15465 -15270 18485 -15204
rect 15192 -15470 15298 -15330
rect 12058 -15596 15078 -15530
rect 12058 -18284 12110 -15596
rect 15026 -18284 15078 -15596
rect 12058 -18350 15078 -18284
rect 11785 -18480 11891 -18410
rect 13515 -18480 13621 -18350
rect 15192 -18410 15231 -15470
rect 15259 -18410 15298 -15470
rect 16922 -15530 17028 -15270
rect 18599 -15330 18638 -12390
rect 18666 -15330 18705 -12390
rect 18599 -15470 18705 -15330
rect 15465 -15596 18485 -15530
rect 15465 -18284 15517 -15596
rect 18433 -18284 18485 -15596
rect 15465 -18350 18485 -18284
rect 15192 -18480 15298 -18410
rect 16922 -18480 17028 -18350
rect 18599 -18410 18638 -15470
rect 18666 -18410 18705 -15470
rect 18599 -18480 18705 -18410
<< properties >>
string FIXED_BBOX 15365 15430 18585 18450
<< end >>
