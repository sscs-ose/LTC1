magic
tech gf180mcuD
magscale 1 10
timestamp 1713277963
<< checkpaint >>
rect -3637 -2810 4187 3564
<< nwell >>
rect -1604 1453 -712 1536
rect -1287 1438 -968 1453
rect -1287 1433 -1028 1438
<< pwell >>
rect -650 591 -427 612
rect -775 406 -427 591
rect 766 -421 891 -222
rect 1442 -421 1538 -61
<< psubdiff >>
rect -1229 120 -1098 145
rect -1229 74 -1180 120
rect -1134 74 -1098 120
rect -1229 50 -1098 74
<< nsubdiff >>
rect -1287 1499 -968 1512
rect -1287 1453 -1270 1499
rect -1130 1453 -968 1499
rect -1287 1438 -968 1453
<< psubdiffcont >>
rect -1180 74 -1134 120
<< nsubdiffcont >>
rect -1270 1453 -1130 1499
<< polysilicon >>
rect -1430 1007 -886 1055
rect -1430 651 -1318 710
rect -1430 605 -1404 651
rect -1358 613 -1318 651
rect -1358 605 -886 613
rect -1430 567 -886 605
rect -998 263 -886 289
rect -998 217 -962 263
rect -916 217 -886 263
rect -998 200 -886 217
<< polycontact >>
rect -1404 605 -1358 651
rect -962 217 -916 263
<< metal1 >>
rect -1508 1499 -778 1513
rect -1508 1453 -1270 1499
rect -1130 1498 -778 1499
rect -1130 1495 -529 1498
rect -1130 1453 -590 1495
rect -1508 1443 -590 1453
rect -538 1443 -529 1495
rect 692 1446 957 1496
rect -1508 1441 -529 1443
rect -1508 1439 -530 1441
rect -1508 1433 -778 1439
rect -1505 741 -1459 1433
rect -1426 660 -1335 672
rect -1637 651 -1335 660
rect -1637 605 -1404 651
rect -1358 605 -1335 651
rect -1637 597 -1335 605
rect -1426 586 -1335 597
rect -1289 652 -1243 1321
rect -1073 741 -1027 1433
rect -857 1050 -811 1321
rect -857 982 -707 1050
rect 766 1009 873 1055
rect 729 1006 873 1009
rect -857 652 -811 982
rect 827 845 873 1006
rect -1289 604 -811 652
rect -1505 146 -1459 521
rect -1289 301 -1243 604
rect -1073 146 -1027 521
rect -857 301 -811 604
rect -724 587 -558 636
rect 392 459 462 462
rect 392 407 401 459
rect 453 407 462 459
rect 392 405 462 407
rect 641 460 711 463
rect 641 408 650 460
rect 702 408 711 460
rect 1914 417 2187 464
rect 641 406 711 408
rect -599 303 -529 306
rect -980 263 -899 277
rect -980 217 -962 263
rect -916 249 -899 263
rect -599 251 -590 303
rect -538 251 -529 303
rect -599 249 -529 251
rect -916 217 -691 249
rect -980 203 -691 217
rect -1531 120 -790 146
rect -1531 74 -1180 120
rect -1134 74 -790 120
rect -1531 49 -790 74
rect -991 -737 -931 49
rect -738 -144 -691 203
rect 818 -77 941 13
rect 818 -138 869 -77
rect -746 -212 -574 -144
rect 768 -184 869 -138
rect 768 -185 827 -184
rect -715 -607 -559 -558
rect 920 -725 979 -520
rect 671 -730 979 -725
rect 392 -734 462 -731
rect -991 -788 -603 -737
rect 392 -786 401 -734
rect 453 -786 462 -734
rect 392 -788 462 -786
rect 641 -733 979 -730
rect 641 -785 650 -733
rect 702 -785 979 -733
rect 641 -787 979 -785
rect 671 -788 979 -787
rect 671 -790 965 -788
<< via1 >>
rect -590 1443 -538 1495
rect 401 407 453 459
rect 650 408 702 460
rect -590 251 -538 303
rect 401 -786 453 -734
rect 650 -785 702 -733
<< metal2 >>
rect -601 1495 -527 1510
rect -601 1443 -590 1495
rect -538 1443 -527 1495
rect -601 1431 -527 1443
rect -599 476 -529 1431
rect -602 316 -529 476
rect 390 459 465 474
rect 390 407 401 459
rect 453 407 465 459
rect 390 392 465 407
rect 639 460 715 475
rect 639 408 650 460
rect 702 408 715 460
rect 639 392 715 408
rect -602 303 -527 316
rect -602 251 -590 303
rect -538 251 -527 303
rect -602 237 -527 251
rect 392 -718 462 392
rect 641 -125 711 392
rect 641 -215 708 -125
rect 641 -718 711 -215
rect 390 -734 465 -718
rect 390 -786 401 -734
rect 453 -786 465 -734
rect 390 -800 465 -786
rect 639 -733 713 -718
rect 639 -785 650 -733
rect 702 -785 713 -733
rect 639 -799 713 -785
use AND2_magic  AND2_magic_0
timestamp 1713185578
transform 1 0 -747 0 1 990
box 35 -598 1575 546
use AND2_magic  AND2_magic_1
timestamp 1713185578
transform 1 0 -747 0 1 -204
box 35 -598 1575 546
use nmos_3p3_G2UGVV  nmos_3p3_G2UGVV_0
timestamp 1713185578
transform 1 0 -1158 0 1 411
box -384 -180 384 180
use OR_magic  OR_magic_0
timestamp 1713277963
transform 1 0 828 0 1 925
box 0 -1478 1136 611
use pmos_3p3_VRCSD7  pmos_3p3_VRCSD7_0
timestamp 1713185578
transform 1 0 -1158 0 1 1031
box -446 -422 446 422
<< labels >>
flabel psubdiffcont -1157 98 -1157 98 0 FreeSans 750 0 0 0 VSS
flabel metal1 s -701 611 -701 611 0 FreeSans 750 0 0 0 IN1
port 1 nsew
flabel metal1 s -701 -588 -701 -588 0 FreeSans 750 0 0 0 IN2
port 2 nsew
flabel metal1 s 2142 436 2142 436 0 FreeSans 750 0 0 0 VOUT
port 3 nsew
flabel metal1 s -1530 626 -1530 626 0 FreeSans 750 0 0 0 SEL
port 4 nsew
flabel metal1 s -1001 1478 -1001 1478 0 FreeSans 1250 0 0 0 VDD
port 5 nsew
<< end >>
