magic
tech gf180mcuC
magscale 1 10
timestamp 1693477706
<< nwell >>
rect 1151 1068 2091 1226
rect 1598 1036 1644 1068
rect 1946 1036 1992 1068
<< psubdiff >>
rect 1017 1319 2227 1332
rect 1017 1266 1031 1319
rect 1083 1266 1192 1319
rect 1244 1266 1353 1319
rect 1405 1266 1514 1319
rect 1566 1266 1675 1319
rect 1727 1266 1836 1319
rect 1888 1266 1997 1319
rect 2049 1266 2158 1319
rect 2210 1266 2227 1319
rect 1017 1250 2227 1266
rect 1017 1158 1096 1250
rect 1017 1105 1031 1158
rect 1083 1105 1096 1158
rect 2148 1158 2227 1250
rect 2148 1105 2162 1158
rect 2214 1105 2227 1158
rect 1017 997 1096 1105
rect 1017 944 1031 997
rect 1083 944 1096 997
rect 1017 836 1096 944
rect 2148 997 2227 1105
rect 2148 944 2162 997
rect 2214 944 2227 997
rect 1017 783 1031 836
rect 1083 783 1096 836
rect 1017 675 1096 783
rect 2148 836 2227 944
rect 2148 783 2162 836
rect 2214 783 2227 836
rect 1017 622 1031 675
rect 1083 622 1096 675
rect 1017 515 1096 622
rect 1017 462 1031 515
rect 1083 462 1096 515
rect 1017 430 1096 462
rect 2148 675 2227 783
rect 2148 622 2162 675
rect 2214 622 2227 675
rect 2148 515 2227 622
rect 2148 462 2162 515
rect 2214 462 2227 515
rect 2148 430 2227 462
rect 1017 414 2227 430
rect 1017 361 1032 414
rect 1084 361 1193 414
rect 1245 361 1354 414
rect 1406 361 1515 414
rect 1567 361 1676 414
rect 1728 361 1837 414
rect 1889 361 1998 414
rect 2050 361 2159 414
rect 2211 361 2227 414
rect 1017 348 2227 361
<< nsubdiff >>
rect 1329 1167 1920 1181
rect 1329 1166 1451 1167
rect 1329 1119 1347 1166
rect 1393 1120 1451 1166
rect 1497 1120 1558 1167
rect 1604 1166 1920 1167
rect 1604 1120 1663 1166
rect 1393 1119 1663 1120
rect 1709 1165 1920 1166
rect 1709 1119 1784 1165
rect 1329 1118 1784 1119
rect 1830 1118 1920 1165
rect 1329 1105 1920 1118
<< psubdiffcont >>
rect 1031 1266 1083 1319
rect 1192 1266 1244 1319
rect 1353 1266 1405 1319
rect 1514 1266 1566 1319
rect 1675 1266 1727 1319
rect 1836 1266 1888 1319
rect 1997 1266 2049 1319
rect 2158 1266 2210 1319
rect 1031 1105 1083 1158
rect 2162 1105 2214 1158
rect 1031 944 1083 997
rect 2162 944 2214 997
rect 1031 783 1083 836
rect 2162 783 2214 836
rect 1031 622 1083 675
rect 1031 462 1083 515
rect 2162 622 2214 675
rect 2162 462 2214 515
rect 1032 361 1084 414
rect 1193 361 1245 414
rect 1354 361 1406 414
rect 1515 361 1567 414
rect 1676 361 1728 414
rect 1837 361 1889 414
rect 1998 361 2050 414
rect 2159 361 2211 414
<< nsubdiffcont >>
rect 1347 1119 1393 1166
rect 1451 1120 1497 1167
rect 1558 1120 1604 1167
rect 1663 1119 1709 1166
rect 1784 1118 1830 1165
<< polysilicon >>
rect 1325 878 1395 894
rect 1259 876 1395 878
rect 1499 876 1569 894
rect 1673 876 1743 894
rect 1847 876 1917 894
rect 1259 859 1917 876
rect 1259 809 1272 859
rect 1321 809 1917 859
rect 1259 801 1917 809
rect 1259 796 1395 801
rect 1325 761 1395 796
rect 1499 761 1569 801
rect 1673 761 1743 801
rect 1847 761 1917 801
<< polycontact >>
rect 1272 809 1321 859
<< metal1 >>
rect 1017 1319 2227 1332
rect 1017 1266 1031 1319
rect 1083 1266 1192 1319
rect 1244 1266 1353 1319
rect 1405 1266 1514 1319
rect 1566 1266 1675 1319
rect 1727 1266 1836 1319
rect 1888 1266 1997 1319
rect 2049 1266 2158 1319
rect 2210 1266 2227 1319
rect 1017 1250 2227 1266
rect 1017 1158 1096 1250
rect 1017 1105 1031 1158
rect 1083 1105 1096 1158
rect 1017 997 1096 1105
rect 1249 1167 1992 1181
rect 1249 1166 1451 1167
rect 1249 1119 1347 1166
rect 1393 1120 1451 1166
rect 1497 1120 1558 1167
rect 1604 1166 1992 1167
rect 1604 1120 1663 1166
rect 1393 1119 1663 1120
rect 1709 1165 1992 1166
rect 1709 1119 1784 1165
rect 1249 1118 1784 1119
rect 1830 1118 1992 1165
rect 1249 1105 1992 1118
rect 1249 1036 1296 1105
rect 1598 1036 1644 1105
rect 1946 1036 1992 1105
rect 2148 1158 2227 1250
rect 2148 1105 2162 1158
rect 2214 1105 2227 1158
rect 1017 944 1031 997
rect 1083 944 1096 997
rect 1017 836 1096 944
rect 2148 997 2227 1105
rect 2148 944 2162 997
rect 2214 944 2227 997
rect 1258 863 1329 866
rect 1017 783 1031 836
rect 1083 783 1096 836
rect 1154 859 1329 863
rect 1154 809 1272 859
rect 1321 809 1329 859
rect 1154 803 1329 809
rect 1258 798 1329 803
rect 1424 836 1470 940
rect 1772 836 1818 940
rect 2148 836 2227 944
rect 1017 675 1096 783
rect 1424 790 2004 836
rect 1424 715 1470 790
rect 1772 715 1818 790
rect 2148 783 2162 836
rect 2214 783 2227 836
rect 1017 622 1031 675
rect 1083 622 1096 675
rect 1017 515 1096 622
rect 2148 675 2227 783
rect 2148 622 2162 675
rect 2214 622 2227 675
rect 1017 462 1031 515
rect 1083 462 1096 515
rect 1017 430 1096 462
rect 1250 430 1296 519
rect 1598 430 1644 521
rect 1946 430 1992 519
rect 2148 515 2227 622
rect 2148 462 2162 515
rect 2214 462 2227 515
rect 2148 430 2227 462
rect 1017 414 2227 430
rect 1017 361 1032 414
rect 1084 361 1193 414
rect 1245 361 1354 414
rect 1406 361 1515 414
rect 1567 361 1676 414
rect 1728 361 1837 414
rect 1889 361 1998 414
rect 2050 361 2159 414
rect 2211 361 2227 414
rect 1017 348 2227 361
use nmos_3p3_VDSZE6  nmos_3p3_VDSZE6_0
timestamp 1693477706
transform 1 0 1621 0 1 617
box -408 -168 408 168
use pmos_3p3_HDJZPK  pmos_3p3_HDJZPK_0
timestamp 1693477706
transform 1 0 1621 0 1 988
box -470 -180 470 180
<< labels >>
flabel metal1 1984 810 1984 810 0 FreeSans 640 0 0 0 OUT
port 1 nsew
flabel metal1 1621 1140 1621 1140 0 FreeSans 640 0 0 0 VDD
port 3 nsew
flabel metal1 1163 825 1163 825 0 FreeSans 640 0 0 0 IN
port 0 nsew
flabel metal1 1270 450 1270 450 0 FreeSans 640 0 0 0 VSS
port 4 nsew
<< end >>
