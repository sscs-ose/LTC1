magic
tech gf180mcuC
magscale 1 10
timestamp 1714543819
<< nwell >>
rect 5305 1636 5343 1716
rect 4684 323 4750 387
rect 5729 318 6019 329
rect 6030 318 6092 383
<< pwell >>
rect 1545 904 2949 1008
rect 1545 675 2961 904
rect 7988 681 9404 910
<< psubdiff >>
rect 3886 -942 3898 -914
<< nsubdiff >>
rect 5305 1636 5343 1716
<< metal1 >>
rect 5177 3368 5362 3382
rect 5177 3316 5190 3368
rect 5242 3316 5296 3368
rect 5348 3316 5362 3368
rect 5177 3302 5362 3316
rect 2881 3080 3400 3179
rect 5226 2968 5311 3302
rect 5177 2954 5362 2968
rect 5177 2902 5190 2954
rect 5242 2902 5296 2954
rect 5348 2902 5362 2954
rect 5177 2888 5362 2902
rect 3501 2741 6585 2822
rect 500 2549 685 2563
rect 500 2497 514 2549
rect 566 2497 620 2549
rect 672 2497 685 2549
rect 500 2483 685 2497
rect 6937 2549 7122 2563
rect 6937 2497 6951 2549
rect 7003 2497 7057 2549
rect 7109 2497 7122 2549
rect 6937 2483 7122 2497
rect 4347 2426 4427 2439
rect 4347 2374 4361 2426
rect 4413 2374 4427 2426
rect 5232 2417 5312 2430
rect 4347 2320 4427 2374
rect 4347 2268 4361 2320
rect 4413 2268 4427 2320
rect 4654 2364 4839 2378
rect 4654 2312 4668 2364
rect 4720 2312 4774 2364
rect 4826 2312 4839 2364
rect 4654 2298 4839 2312
rect 5232 2365 5246 2417
rect 5298 2365 5312 2417
rect 5232 2311 5312 2365
rect 4347 2254 4427 2268
rect 5232 2259 5246 2311
rect 5298 2259 5312 2311
rect 5532 2375 5717 2389
rect 5532 2323 5546 2375
rect 5598 2323 5652 2375
rect 5704 2323 5717 2375
rect 5532 2309 5717 2323
rect 5232 2245 5312 2259
rect 466 1941 651 1955
rect 466 1889 480 1941
rect 532 1889 586 1941
rect 638 1889 651 1941
rect 466 1875 651 1889
rect 6935 1937 7120 1951
rect 6935 1885 6949 1937
rect 7001 1885 7055 1937
rect 7107 1885 7120 1937
rect 6935 1871 7120 1885
rect 3500 1760 6583 1850
rect 490 1284 878 1321
rect 490 1226 681 1284
rect 739 1226 878 1284
rect 490 1213 878 1226
rect 2891 1284 2970 1298
rect 2891 1226 2903 1284
rect 2961 1226 2970 1284
rect 2891 1213 2970 1226
rect 7108 1285 7191 1299
rect 9402 1298 9784 1328
rect 7108 1227 7124 1285
rect 7182 1227 7191 1285
rect 7108 1215 7191 1227
rect 9340 1284 9784 1298
rect 9340 1226 9346 1284
rect 9404 1226 9784 1284
rect 9340 1213 9784 1226
rect 9402 1197 9784 1213
rect 4296 1180 4481 1194
rect 4296 1128 4310 1180
rect 4362 1128 4416 1180
rect 4468 1128 4481 1180
rect 4296 1114 4481 1128
rect 4678 1169 4863 1183
rect 4678 1117 4692 1169
rect 4744 1117 4798 1169
rect 4850 1117 4863 1169
rect 4678 1103 4863 1117
rect 5213 1176 5398 1190
rect 5213 1124 5227 1176
rect 5279 1124 5333 1176
rect 5385 1124 5398 1176
rect 5213 1110 5398 1124
rect 5586 1169 5771 1183
rect 5586 1117 5600 1169
rect 5652 1117 5706 1169
rect 5758 1117 5771 1169
rect 5586 1103 5771 1117
rect 3497 527 6582 644
rect 3512 526 3988 527
rect 5117 526 5320 527
rect 4684 382 4770 393
rect 1683 354 1868 368
rect 1683 302 1697 354
rect 1749 302 1803 354
rect 1855 302 1868 354
rect 1683 288 1868 302
rect 2549 354 2734 368
rect 2549 302 2563 354
rect 2615 302 2669 354
rect 2721 302 2734 354
rect 4684 330 4696 382
rect 4748 330 4770 382
rect 4684 321 4770 330
rect 6025 379 6099 406
rect 6025 327 6031 379
rect 6083 327 6099 379
rect 6025 310 6099 327
rect 8124 351 8309 365
rect 2549 288 2734 302
rect 8124 299 8138 351
rect 8190 299 8244 351
rect 8296 299 8309 351
rect 8124 285 8309 299
rect 8982 351 9167 365
rect 8982 299 8996 351
rect 9048 299 9102 351
rect 9154 299 9167 351
rect 8982 285 9167 299
rect 3910 -391 4095 -377
rect 3910 -443 3924 -391
rect 3976 -443 4030 -391
rect 4082 -443 4095 -391
rect 5254 -391 5439 -377
rect 3910 -457 4095 -443
rect 4703 -448 4837 -401
rect 5254 -443 5268 -391
rect 5320 -443 5374 -391
rect 5426 -443 5439 -391
rect 5254 -457 5439 -443
rect 6033 -449 6167 -402
rect 3499 -1031 6583 -914
rect 478 -1190 663 -1176
rect 478 -1242 492 -1190
rect 544 -1242 598 -1190
rect 650 -1242 663 -1190
rect 6906 -1192 7091 -1178
rect 478 -1256 663 -1242
rect 5729 -1245 5809 -1232
rect 5729 -1270 5743 -1245
rect 5703 -1297 5743 -1270
rect 5795 -1297 5809 -1245
rect 6906 -1244 6920 -1192
rect 6972 -1244 7026 -1192
rect 7078 -1244 7091 -1192
rect 6906 -1258 7091 -1244
rect 5703 -1351 5809 -1297
rect 5703 -1403 5743 -1351
rect 5795 -1403 5809 -1351
rect 5703 -1417 5809 -1403
rect 4572 -1594 4757 -1580
rect 4572 -1646 4586 -1594
rect 4638 -1646 4692 -1594
rect 4744 -1646 4757 -1594
rect 4572 -1660 4757 -1646
rect 5328 -1616 5513 -1602
rect 5328 -1668 5342 -1616
rect 5394 -1668 5448 -1616
rect 5500 -1668 5513 -1616
rect 5328 -1682 5513 -1668
rect 464 -1800 649 -1786
rect 464 -1852 478 -1800
rect 530 -1852 584 -1800
rect 636 -1852 649 -1800
rect 464 -1866 649 -1852
rect 3497 -2110 5636 -2030
rect 5703 -2325 5783 -1417
rect 6905 -1809 7090 -1795
rect 6905 -1861 6919 -1809
rect 6971 -1861 7025 -1809
rect 7077 -1861 7090 -1809
rect 6905 -1875 7090 -1861
rect 5703 -2377 5717 -2325
rect 5769 -2377 5783 -2325
rect 5703 -2431 5783 -2377
rect 667 -2454 742 -2440
rect 667 -2512 681 -2454
rect 739 -2512 742 -2454
rect 667 -2525 742 -2512
rect 2898 -2454 2973 -2441
rect 2898 -2512 2903 -2454
rect 2961 -2512 2973 -2454
rect 5703 -2483 5717 -2431
rect 5769 -2483 5783 -2431
rect 5703 -2497 5783 -2483
rect 7107 -2454 7185 -2440
rect 2898 -2526 2973 -2512
rect 7107 -2512 7124 -2454
rect 7182 -2512 7185 -2454
rect 7107 -2525 7185 -2512
rect 9342 -2454 9417 -2440
rect 9342 -2512 9346 -2454
rect 9404 -2512 9417 -2454
rect 9342 -2525 9417 -2512
rect 5698 -2633 5778 -2620
rect 4570 -2673 4755 -2659
rect 5698 -2671 5712 -2633
rect 4570 -2725 4584 -2673
rect 4636 -2725 4690 -2673
rect 4742 -2725 4755 -2673
rect 4570 -2739 4755 -2725
rect 5328 -2696 5513 -2682
rect 5328 -2748 5342 -2696
rect 5394 -2748 5448 -2696
rect 5500 -2748 5513 -2696
rect 5328 -2762 5513 -2748
rect 5692 -2685 5712 -2671
rect 5764 -2671 5778 -2633
rect 6015 -2635 6095 -2622
rect 6015 -2671 6029 -2635
rect 5764 -2685 6029 -2671
rect 5692 -2687 6029 -2685
rect 6081 -2687 6095 -2635
rect 5692 -2739 6095 -2687
rect 5692 -2772 5712 -2739
rect 5698 -2791 5712 -2772
rect 5764 -2741 6095 -2739
rect 5764 -2772 6029 -2741
rect 5764 -2791 5778 -2772
rect 5698 -2805 5778 -2791
rect 6015 -2793 6029 -2772
rect 6081 -2793 6095 -2741
rect 6015 -2807 6095 -2793
rect 3500 -3187 6582 -3106
rect 1681 -3380 1866 -3366
rect 1681 -3432 1695 -3380
rect 1747 -3432 1801 -3380
rect 1853 -3432 1866 -3380
rect 1681 -3446 1866 -3432
rect 2539 -3386 2724 -3372
rect 2539 -3438 2553 -3386
rect 2605 -3438 2659 -3386
rect 2711 -3438 2724 -3386
rect 2539 -3452 2724 -3438
rect 8118 -3385 8303 -3371
rect 8118 -3437 8132 -3385
rect 8184 -3437 8238 -3385
rect 8290 -3437 8303 -3385
rect 8118 -3451 8303 -3437
rect 8984 -3384 9169 -3370
rect 8984 -3436 8998 -3384
rect 9050 -3436 9104 -3384
rect 9156 -3436 9169 -3384
rect 8984 -3450 9169 -3436
rect 3494 -3734 6579 -3600
<< via1 >>
rect 5190 3316 5242 3368
rect 5296 3316 5348 3368
rect 5190 2902 5242 2954
rect 5296 2902 5348 2954
rect 4682 2611 4734 2663
rect 5555 2614 5607 2666
rect 514 2497 566 2549
rect 620 2497 672 2549
rect 6951 2497 7003 2549
rect 7057 2497 7109 2549
rect 4361 2374 4413 2426
rect 4361 2268 4413 2320
rect 4668 2312 4720 2364
rect 4774 2312 4826 2364
rect 5246 2365 5298 2417
rect 5246 2259 5298 2311
rect 5546 2323 5598 2375
rect 5652 2323 5704 2375
rect 480 1889 532 1941
rect 586 1889 638 1941
rect 6949 1885 7001 1937
rect 7055 1885 7107 1937
rect 387 1654 440 1707
rect 4751 1630 4803 1682
rect 5653 1629 5705 1681
rect 6712 1671 6764 1723
rect 9761 1662 9813 1714
rect 681 1226 739 1284
rect 2903 1226 2961 1284
rect 7124 1227 7182 1285
rect 9346 1226 9404 1284
rect 4310 1128 4362 1180
rect 4416 1128 4468 1180
rect 4692 1117 4744 1169
rect 4798 1117 4850 1169
rect 5227 1124 5279 1176
rect 5333 1124 5385 1176
rect 5600 1117 5652 1169
rect 5706 1117 5758 1169
rect 1697 302 1749 354
rect 1803 302 1855 354
rect 2563 302 2615 354
rect 2669 302 2721 354
rect 4696 330 4748 382
rect 6031 327 6083 379
rect 8138 299 8190 351
rect 8244 299 8296 351
rect 8996 299 9048 351
rect 9102 299 9154 351
rect 3924 -443 3976 -391
rect 4030 -443 4082 -391
rect 5268 -443 5320 -391
rect 5374 -443 5426 -391
rect 385 -635 437 -583
rect 3229 -635 3281 -583
rect 9764 -646 9816 -594
rect 492 -1242 544 -1190
rect 598 -1242 650 -1190
rect 4675 -1341 4727 -1289
rect 5743 -1297 5795 -1245
rect 6920 -1244 6972 -1192
rect 7026 -1244 7078 -1192
rect 5743 -1403 5795 -1351
rect 4586 -1646 4638 -1594
rect 4692 -1646 4744 -1594
rect 5342 -1668 5394 -1616
rect 5448 -1668 5500 -1616
rect 478 -1852 530 -1800
rect 584 -1852 636 -1800
rect 6919 -1861 6971 -1809
rect 7025 -1861 7077 -1809
rect 6709 -2033 6761 -1981
rect 5336 -2418 5388 -2366
rect 5717 -2377 5769 -2325
rect 681 -2512 739 -2454
rect 2903 -2512 2961 -2454
rect 5717 -2483 5769 -2431
rect 7124 -2512 7182 -2454
rect 9346 -2512 9404 -2454
rect 4584 -2725 4636 -2673
rect 4690 -2725 4742 -2673
rect 5342 -2748 5394 -2696
rect 5448 -2748 5500 -2696
rect 5712 -2685 5764 -2633
rect 6029 -2687 6081 -2635
rect 5712 -2791 5764 -2739
rect 6029 -2793 6081 -2741
rect 1695 -3432 1747 -3380
rect 1801 -3432 1853 -3380
rect 2553 -3438 2605 -3386
rect 2659 -3438 2711 -3386
rect 8132 -3437 8184 -3385
rect 8238 -3437 8290 -3385
rect 8998 -3436 9050 -3384
rect 9104 -3436 9156 -3384
<< metal2 >>
rect 3332 3368 6521 3408
rect 3332 3316 5190 3368
rect 5242 3316 5296 3368
rect 5348 3316 6521 3368
rect 3332 3259 6521 3316
rect -5 2549 686 2572
rect -5 2497 514 2549
rect 566 2497 620 2549
rect 672 2497 686 2549
rect -5 2468 686 2497
rect -5 -3627 99 2468
rect 195 1941 652 1964
rect 195 1889 480 1941
rect 532 1889 586 1941
rect 638 1889 652 1941
rect 195 1860 652 1889
rect 195 -3364 299 1860
rect 372 1707 451 1721
rect 372 1654 387 1707
rect 440 1654 451 1707
rect 372 -583 451 1654
rect 666 1284 749 1298
rect 666 1226 681 1284
rect 739 1226 749 1284
rect 666 1214 749 1226
rect 2891 1284 2970 1298
rect 2891 1226 2903 1284
rect 2961 1226 2970 1284
rect 2891 1213 2970 1226
rect 1683 354 1868 368
rect 1683 302 1697 354
rect 1749 302 1803 354
rect 1855 302 1868 354
rect 1683 288 1868 302
rect 2549 354 2734 368
rect 2549 302 2563 354
rect 2615 302 2669 354
rect 2721 343 2734 354
rect 3332 343 3481 3259
rect 3844 3045 6296 3194
rect 3844 1004 3993 3045
rect 4327 2428 4430 3045
rect 5177 2954 5362 2968
rect 5177 2902 5190 2954
rect 5242 2902 5296 2954
rect 5348 2902 5362 2954
rect 5177 2888 5362 2902
rect 4670 2663 5084 2684
rect 4670 2611 4682 2663
rect 4734 2611 5084 2663
rect 4670 2598 5084 2611
rect 4347 2426 4427 2428
rect 4347 2374 4361 2426
rect 4413 2374 4427 2426
rect 4347 2320 4427 2374
rect 4347 2268 4361 2320
rect 4413 2268 4427 2320
rect 4652 2364 4910 2392
rect 4652 2312 4668 2364
rect 4720 2312 4774 2364
rect 4826 2312 4910 2364
rect 4652 2283 4910 2312
rect 4347 2254 4427 2268
rect 4809 1955 4910 2283
rect 4191 1854 4910 1955
rect 4191 1216 4292 1854
rect 4998 1700 5084 2598
rect 5219 2419 5322 2888
rect 5543 2666 6059 2677
rect 5543 2614 5555 2666
rect 5607 2614 6059 2666
rect 5543 2591 6059 2614
rect 5232 2417 5312 2419
rect 5232 2365 5246 2417
rect 5298 2365 5312 2417
rect 5232 2311 5312 2365
rect 5232 2259 5246 2311
rect 5298 2259 5312 2311
rect 5531 2375 5790 2401
rect 5531 2323 5546 2375
rect 5598 2323 5652 2375
rect 5704 2323 5790 2375
rect 5531 2295 5790 2323
rect 5232 2245 5312 2259
rect 5182 1936 5240 1937
rect 5704 1936 5790 2295
rect 5182 1850 5790 1936
rect 4737 1682 5110 1700
rect 4737 1630 4751 1682
rect 4803 1630 5110 1682
rect 4737 1614 5110 1630
rect 4191 1194 4476 1216
rect 4191 1180 4481 1194
rect 4680 1183 4928 1196
rect 4191 1128 4310 1180
rect 4362 1128 4416 1180
rect 4468 1128 4481 1180
rect 4191 1115 4481 1128
rect 4296 1114 4481 1115
rect 4678 1169 4928 1183
rect 4678 1117 4692 1169
rect 4744 1117 4798 1169
rect 4850 1117 4928 1169
rect 4678 1103 4928 1117
rect 4680 1091 4928 1103
rect 2721 302 3481 343
rect 2549 288 3481 302
rect 1715 -61 1864 288
rect 2552 194 3481 288
rect 3559 855 3993 1004
rect 3559 -58 3708 855
rect 4823 634 4928 1091
rect 3440 -61 3708 -58
rect 1715 -207 3708 -61
rect 3852 529 4928 634
rect 1715 -210 3542 -207
rect 3852 -377 3957 529
rect 5024 409 5110 1614
rect 5182 1204 5240 1850
rect 5973 1739 6059 2591
rect 6147 1982 6296 3045
rect 6372 2600 6521 3259
rect 6372 2549 7123 2600
rect 6372 2497 6951 2549
rect 7003 2497 7057 2549
rect 7109 2497 7123 2549
rect 6372 2451 7123 2497
rect 6147 1937 7139 1982
rect 6147 1885 6949 1937
rect 7001 1885 7055 1937
rect 7107 1885 7139 1937
rect 6147 1833 7139 1885
rect 5639 1723 6774 1739
rect 5639 1681 6712 1723
rect 5639 1629 5653 1681
rect 5705 1671 6712 1681
rect 6764 1671 6774 1723
rect 5705 1653 6774 1671
rect 9749 1714 10078 1737
rect 9749 1662 9761 1714
rect 9813 1662 10078 1714
rect 5705 1629 5725 1653
rect 5639 1609 5725 1629
rect 5182 1190 5395 1204
rect 5724 1202 5828 1204
rect 5182 1176 5398 1190
rect 5182 1124 5227 1176
rect 5279 1124 5333 1176
rect 5385 1124 5398 1176
rect 5182 1118 5398 1124
rect 5213 1110 5398 1118
rect 5586 1169 5828 1202
rect 5586 1117 5600 1169
rect 5652 1117 5706 1169
rect 5758 1117 5828 1169
rect 5586 1089 5828 1117
rect 5724 712 5828 1089
rect 4662 382 5110 409
rect 4662 330 4696 382
rect 4748 330 5110 382
rect 4662 323 5110 330
rect 5210 608 5828 712
rect 4684 321 4770 323
rect 3852 -391 4095 -377
rect 3852 -443 3924 -391
rect 3976 -443 4030 -391
rect 4082 -443 4095 -391
rect 3852 -457 4095 -443
rect 3852 -458 3957 -457
rect 372 -635 385 -583
rect 437 -635 451 -583
rect 372 -649 451 -635
rect 3215 -583 3845 -568
rect 3215 -635 3229 -583
rect 3281 -635 3845 -583
rect 3215 -649 3845 -635
rect 3764 -957 3845 -649
rect 4975 -579 5061 323
rect 5210 -353 5283 608
rect 6013 405 6099 1653
rect 9749 1651 10078 1662
rect 7108 1285 7191 1299
rect 7108 1227 7124 1285
rect 7182 1227 7191 1285
rect 7108 1215 7191 1227
rect 9340 1284 9419 1298
rect 9340 1226 9346 1284
rect 9404 1226 9419 1284
rect 9340 1213 9419 1226
rect 5647 379 6099 405
rect 5647 327 6031 379
rect 6083 327 6099 379
rect 5647 318 6099 327
rect 6492 365 8128 366
rect 6492 351 8309 365
rect 5210 -391 5440 -353
rect 5210 -443 5268 -391
rect 5320 -443 5374 -391
rect 5426 -443 5440 -391
rect 5210 -457 5440 -443
rect 5647 -579 5733 318
rect 4975 -665 5733 -579
rect 6492 299 8138 351
rect 8190 299 8244 351
rect 8296 299 8309 351
rect 6492 285 8309 299
rect 8982 351 9167 365
rect 8982 299 8996 351
rect 9048 299 9102 351
rect 9154 299 9167 351
rect 8982 285 9167 299
rect 6492 260 8273 285
rect 3764 -1038 4747 -957
rect 478 -1190 4377 -1123
rect 478 -1242 492 -1190
rect 544 -1242 598 -1190
rect 650 -1227 4377 -1190
rect 650 -1242 663 -1227
rect 478 -1256 663 -1242
rect 4103 -1323 4196 -1320
rect 362 -1411 4196 -1323
rect 362 -1778 450 -1411
rect 362 -1786 647 -1778
rect 362 -1800 649 -1786
rect 362 -1852 478 -1800
rect 530 -1852 584 -1800
rect 636 -1852 649 -1800
rect 362 -1866 649 -1852
rect 362 -1873 647 -1866
rect 667 -2454 742 -2440
rect 667 -2512 681 -2454
rect 739 -2512 742 -2454
rect 667 -2525 742 -2512
rect 2898 -2454 2973 -2441
rect 2898 -2512 2903 -2454
rect 2961 -2512 2973 -2454
rect 2898 -2526 2973 -2512
rect 4103 -2658 4196 -1411
rect 4273 -1562 4377 -1227
rect 4666 -1270 4747 -1038
rect 5729 -1245 5809 -1232
rect 5729 -1270 5743 -1245
rect 4666 -1289 5743 -1270
rect 4666 -1341 4675 -1289
rect 4727 -1297 5743 -1289
rect 5795 -1270 5809 -1245
rect 5795 -1297 6335 -1270
rect 4727 -1341 6335 -1297
rect 4666 -1351 6335 -1341
rect 5729 -1403 5743 -1351
rect 5795 -1403 5809 -1351
rect 5729 -1417 5809 -1403
rect 4273 -1594 4757 -1562
rect 4273 -1646 4586 -1594
rect 4638 -1646 4692 -1594
rect 4744 -1646 4757 -1594
rect 4273 -1666 4757 -1646
rect 5328 -1616 5945 -1590
rect 5328 -1668 5342 -1616
rect 5394 -1668 5448 -1616
rect 5500 -1668 5945 -1616
rect 5328 -1694 5945 -1668
rect 5703 -2325 5783 -2312
rect 5703 -2349 5717 -2325
rect 5321 -2366 5717 -2349
rect 5321 -2418 5336 -2366
rect 5388 -2377 5717 -2366
rect 5769 -2377 5783 -2325
rect 5388 -2418 5783 -2377
rect 5321 -2430 5783 -2418
rect 5703 -2431 5783 -2430
rect 5703 -2483 5717 -2431
rect 5769 -2483 5783 -2431
rect 5703 -2497 5783 -2483
rect 5698 -2633 5778 -2620
rect 4103 -2673 4757 -2658
rect 5698 -2671 5712 -2633
rect 4103 -2725 4584 -2673
rect 4636 -2725 4690 -2673
rect 4742 -2725 4757 -2673
rect 4103 -2751 4757 -2725
rect 5325 -2685 5712 -2671
rect 5764 -2685 5778 -2633
rect 5325 -2696 5778 -2685
rect 5325 -2748 5342 -2696
rect 5394 -2748 5448 -2696
rect 5500 -2739 5778 -2696
rect 5500 -2748 5712 -2739
rect 5325 -2772 5712 -2748
rect 5698 -2791 5712 -2772
rect 5764 -2791 5778 -2739
rect 5698 -2805 5778 -2791
rect 195 -3366 1827 -3364
rect 195 -3380 1866 -3366
rect 195 -3432 1695 -3380
rect 1747 -3432 1801 -3380
rect 1853 -3432 1866 -3380
rect 195 -3446 1866 -3432
rect 2539 -3386 2724 -3372
rect 2539 -3438 2553 -3386
rect 2605 -3438 2659 -3386
rect 2711 -3438 2724 -3386
rect 195 -3468 1827 -3446
rect 2539 -3452 2724 -3438
rect 2543 -3627 2647 -3452
rect -5 -3731 2647 -3627
rect 5841 -3623 5945 -1694
rect 6254 -1961 6335 -1351
rect 6492 -1778 6598 260
rect 9009 -61 9115 285
rect 6668 -167 9115 -61
rect 6668 -1160 6774 -167
rect 9992 -579 10078 1651
rect 9741 -594 10078 -579
rect 9741 -646 9764 -594
rect 9816 -646 10078 -594
rect 9741 -665 10078 -646
rect 6668 -1192 7095 -1160
rect 6668 -1244 6920 -1192
rect 6972 -1244 7026 -1192
rect 7078 -1244 7095 -1192
rect 6668 -1266 7095 -1244
rect 6492 -1795 7089 -1778
rect 6492 -1809 7090 -1795
rect 6492 -1861 6919 -1809
rect 6971 -1861 7025 -1809
rect 7077 -1861 7090 -1809
rect 6492 -1875 7090 -1861
rect 6492 -1884 7089 -1875
rect 6254 -1981 6780 -1961
rect 6254 -2033 6709 -1981
rect 6761 -2033 6780 -1981
rect 6254 -2042 6780 -2033
rect 7107 -2454 7185 -2440
rect 7107 -2512 7124 -2454
rect 7182 -2512 7185 -2454
rect 7107 -2525 7185 -2512
rect 9342 -2454 9417 -2440
rect 9342 -2512 9346 -2454
rect 9404 -2512 9417 -2454
rect 9342 -2525 9417 -2512
rect 6015 -2635 6095 -2622
rect 6015 -2687 6029 -2635
rect 6081 -2673 6095 -2635
rect 6081 -2687 6244 -2673
rect 6015 -2741 6244 -2687
rect 6015 -2793 6029 -2741
rect 6081 -2793 6244 -2741
rect 6015 -2807 6244 -2793
rect 6144 -3375 6244 -2807
rect 8118 -3375 8303 -3371
rect 6144 -3385 8303 -3375
rect 6144 -3437 8132 -3385
rect 8184 -3437 8238 -3385
rect 8290 -3437 8303 -3385
rect 6144 -3451 8303 -3437
rect 8984 -3384 9169 -3370
rect 8984 -3436 8998 -3384
rect 9050 -3436 9104 -3384
rect 9156 -3436 9169 -3384
rect 8984 -3450 9169 -3436
rect 6144 -3475 8302 -3451
rect 9011 -3623 9115 -3450
rect 5841 -3727 9115 -3623
<< via2 >>
rect 681 1226 739 1284
rect 2903 1226 2961 1284
rect 7124 1227 7182 1285
rect 9346 1226 9404 1284
rect 681 -2512 739 -2454
rect 2903 -2512 2961 -2454
rect 7124 -2512 7182 -2454
rect 9346 -2512 9404 -2454
<< metal3 >>
rect 2867 1500 9445 1634
rect 633 1303 767 1304
rect 633 1284 775 1303
rect 633 1226 681 1284
rect 739 1226 775 1284
rect 633 962 775 1226
rect 2867 1284 3001 1500
rect 2867 1226 2903 1284
rect 2961 1226 3001 1284
rect 2867 1200 3001 1226
rect 7086 1285 7220 1306
rect 7086 1227 7124 1285
rect 7182 1227 7220 1285
rect 7086 962 7220 1227
rect 633 828 7220 962
rect 9311 1284 9445 1500
rect 9311 1226 9346 1284
rect 9404 1226 9445 1284
rect 633 -2454 767 828
rect 9311 -2109 9445 1226
rect 633 -2512 681 -2454
rect 739 -2512 767 -2454
rect 633 -2774 767 -2512
rect 2871 -2243 9448 -2109
rect 2871 -2454 3005 -2243
rect 2871 -2512 2903 -2454
rect 2961 -2512 3005 -2454
rect 2871 -2546 3005 -2512
rect 7085 -2454 7219 -2431
rect 7085 -2512 7124 -2454
rect 7182 -2512 7219 -2454
rect 7085 -2774 7219 -2512
rect 9311 -2454 9448 -2243
rect 9311 -2512 9346 -2454
rect 9404 -2512 9448 -2454
rect 9311 -2534 9448 -2512
rect 9314 -2538 9448 -2534
rect 633 -2908 7219 -2774
use Delay_Cell_mag  Delay_Cell_mag_0
timestamp 1714462644
transform 1 0 6674 0 1 -999
box -231 -2739 3409 681
use Delay_Cell_mag  Delay_Cell_mag_1
timestamp 1714462644
transform 1 0 231 0 1 2739
box -231 -2739 3409 681
use Delay_Cell_mag  Delay_Cell_mag_2
timestamp 1714462644
transform 1 0 231 0 1 -999
box -231 -2739 3409 681
use Delay_Cell_mag  Delay_Cell_mag_3
timestamp 1714462644
transform 1 0 6674 0 1 2740
box -231 -2739 3409 681
use GF_INV1  GF_INV1_0
timestamp 1714543819
transform 1 0 5292 0 1 1979
box -231 -55 589 842
use GF_INV1  GF_INV1_1
timestamp 1714543819
transform 1 0 4416 0 1 1978
box -231 -55 589 842
use GF_INV4  GF_INV4_0
timestamp 1714492828
transform 1 0 5207 0 1 1199
box -146 -481 701 650
use GF_INV4  GF_INV4_1
timestamp 1714492828
transform 1 0 4304 0 1 1199
box -146 -481 701 650
use GF_INV16  GF_INV16_1
timestamp 1714491929
transform 1 0 3969 0 1 -593
box -208 -438 1036 1236
use GF_INV16  GF_INV16_2
timestamp 1714491929
transform 1 0 5290 0 1 -593
box -208 -438 1036 1236
use Stage_INV  Stage_INV_0
timestamp 1714537808
transform 1 0 3411 0 1 -2459
box 1017 348 2227 1332
use Stage_INV  Stage_INV_1
timestamp 1714537808
transform 1 0 3411 0 1 -3536
box 1017 348 2227 1332
<< labels >>
flabel metal1 4977 -3671 4977 -3671 0 FreeSans 1600 0 0 0 VSS
port 0 nsew
flabel metal1 524 1266 524 1266 0 FreeSans 1600 0 0 0 EN
port 1 nsew
flabel metal1 9716 1266 9716 1266 0 FreeSans 1600 0 0 0 VCONT
port 2 nsew
flabel metal1 6136 -430 6136 -430 0 FreeSans 1600 0 0 0 OUT
port 3 nsew
flabel metal1 4788 -423 4788 -423 0 FreeSans 1600 0 0 0 OUTB
port 4 nsew
flabel metal1 3067 3132 3067 3132 0 FreeSans 1600 0 0 0 VDD
port 6 nsew
<< end >>
