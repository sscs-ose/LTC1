magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1019 1019 1019
<< metal1 >>
rect -19 13 19 19
rect -19 -13 -13 13
rect 13 -13 19 13
rect -19 -19 19 -13
<< via1 >>
rect -13 -13 13 13
<< metal2 >>
rect -19 13 19 19
rect -19 -13 -13 13
rect 13 -13 19 13
rect -19 -19 19 -13
<< end >>
